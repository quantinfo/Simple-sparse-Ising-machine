//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [37:0] counter;
initial counter = 38'b0;
reg [15:0] solution;
reg [15:0] solution_check;
wire [15:0] solution_set;
initial solution_check = 16'b1101101101011001;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
reg [0:495] InitCond;
reg run;
wire [275:0] LFSRcolor0;
wire [367:0] LFSRcolor1;
wire [275:0] LFSRcolor2;
wire [45:0] LFSRcolor3;
wire [183:0] LFSRcolor4;
reg [277:0] BiasedRNG;       //For I=+/-1 cases
reg [217:0] UnbiasedRNG;   //For I=0 cases
reg [0:519] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[176] = 1'b1;
initial m[243] = 1'b0;
initial m[253] = 1'b0;
initial m[268] = 1'b1;
initial m[288] = 1'b1;
initial m[313] = 1'b0;
initial m[343] = 1'b1;
initial m[378] = 1'b0;
initial m[413] = 1'b1;
initial m[443] = 1'b1;
initial m[468] = 1'b0;
initial m[488] = 1'b1;
initial m[503] = 1'b1;
initial m[513] = 1'b0;
initial m[518] = 1'b1;
initial m[519] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[242] = 1'b0;
initial m[252] = 1'b0;
initial m[267] = 1'b0;
initial m[287] = 1'b0;
initial m[312] = 1'b0;
initial m[342] = 1'b0;
initial m[377] = 1'b0;
initial m[380] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
//To control whether the system runs or resets using VIO and counter:
always @(posedge sample_clk) begin
    if (reset) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 16'b0;
        failure = 1'b0;
        solution_check = solution_set;
        m[176] = solution_set[0];
        m[243] = solution_set[1];
        m[253] = solution_set[2];
        m[268] = solution_set[3];
        m[288] = solution_set[4];
        m[313] = solution_set[5];
        m[343] = solution_set[6];
        m[378] = solution_set[7];
        m[413] = solution_set[8];
        m[443] = solution_set[9];
        m[468] = solution_set[10];
        m[488] = solution_set[11];
        m[503] = solution_set[12];
        m[513] = solution_set[13];
        m[518] = solution_set[14];
        m[519] = solution_set[15];
    end else if (solution_flag) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 16'b0;
        failure = 1'b0;
    end else if (counter < 38'b11111111111111111111111111111111111111) begin
        if (counter == 1) begin
            InitCond[0] = UnbiasedRNG[0];
            InitCond[1] = UnbiasedRNG[1];
            InitCond[2] = UnbiasedRNG[2];
            InitCond[3] = UnbiasedRNG[3];
            InitCond[4] = UnbiasedRNG[4];
            InitCond[5] = UnbiasedRNG[5];
            InitCond[6] = UnbiasedRNG[6];
            InitCond[7] = UnbiasedRNG[7];
            InitCond[8] = UnbiasedRNG[8];
            InitCond[9] = UnbiasedRNG[9];
            InitCond[10] = UnbiasedRNG[10];
            InitCond[11] = UnbiasedRNG[11];
            InitCond[12] = UnbiasedRNG[12];
            InitCond[13] = UnbiasedRNG[13];
            InitCond[14] = UnbiasedRNG[14];
            InitCond[15] = UnbiasedRNG[15];
            InitCond[16] = UnbiasedRNG[16];
            InitCond[17] = UnbiasedRNG[17];
            InitCond[18] = UnbiasedRNG[18];
            InitCond[19] = UnbiasedRNG[19];
            InitCond[20] = UnbiasedRNG[20];
            InitCond[21] = UnbiasedRNG[21];
            InitCond[22] = UnbiasedRNG[22];
            InitCond[23] = UnbiasedRNG[23];
            InitCond[24] = UnbiasedRNG[24];
            InitCond[25] = UnbiasedRNG[25];
            InitCond[26] = UnbiasedRNG[26];
            InitCond[27] = UnbiasedRNG[27];
            InitCond[28] = UnbiasedRNG[28];
            InitCond[29] = UnbiasedRNG[29];
            InitCond[30] = UnbiasedRNG[30];
            InitCond[31] = UnbiasedRNG[31];
            InitCond[32] = UnbiasedRNG[32];
            InitCond[33] = UnbiasedRNG[33];
            InitCond[34] = UnbiasedRNG[34];
            InitCond[35] = UnbiasedRNG[35];
            InitCond[36] = UnbiasedRNG[36];
            InitCond[37] = UnbiasedRNG[37];
            InitCond[38] = UnbiasedRNG[38];
            InitCond[39] = UnbiasedRNG[39];
            InitCond[40] = UnbiasedRNG[40];
            InitCond[41] = UnbiasedRNG[41];
            InitCond[42] = UnbiasedRNG[42];
            InitCond[43] = UnbiasedRNG[43];
            InitCond[44] = UnbiasedRNG[44];
            InitCond[45] = UnbiasedRNG[45];
            InitCond[46] = UnbiasedRNG[46];
            InitCond[47] = UnbiasedRNG[47];
            InitCond[48] = UnbiasedRNG[48];
            InitCond[49] = UnbiasedRNG[49];
            InitCond[50] = UnbiasedRNG[50];
            InitCond[51] = UnbiasedRNG[51];
            InitCond[52] = UnbiasedRNG[52];
            InitCond[53] = UnbiasedRNG[53];
            InitCond[54] = UnbiasedRNG[54];
            InitCond[55] = UnbiasedRNG[55];
            InitCond[56] = UnbiasedRNG[56];
            InitCond[57] = UnbiasedRNG[57];
            InitCond[58] = UnbiasedRNG[58];
            InitCond[59] = UnbiasedRNG[59];
            InitCond[60] = UnbiasedRNG[60];
            InitCond[61] = UnbiasedRNG[61];
            InitCond[62] = UnbiasedRNG[62];
            InitCond[63] = UnbiasedRNG[63];
            InitCond[64] = UnbiasedRNG[64];
            InitCond[65] = UnbiasedRNG[65];
            InitCond[66] = UnbiasedRNG[66];
            InitCond[67] = UnbiasedRNG[67];
            InitCond[68] = UnbiasedRNG[68];
            InitCond[69] = UnbiasedRNG[69];
            InitCond[70] = UnbiasedRNG[70];
            InitCond[71] = UnbiasedRNG[71];
            InitCond[72] = UnbiasedRNG[72];
            InitCond[73] = UnbiasedRNG[73];
            InitCond[74] = UnbiasedRNG[74];
            InitCond[75] = UnbiasedRNG[75];
            InitCond[76] = UnbiasedRNG[76];
            InitCond[77] = UnbiasedRNG[77];
            InitCond[78] = UnbiasedRNG[78];
            InitCond[79] = UnbiasedRNG[79];
            InitCond[80] = UnbiasedRNG[80];
            InitCond[81] = UnbiasedRNG[81];
            InitCond[82] = UnbiasedRNG[82];
            InitCond[83] = UnbiasedRNG[83];
            InitCond[84] = UnbiasedRNG[84];
            InitCond[85] = UnbiasedRNG[85];
            InitCond[86] = UnbiasedRNG[86];
            InitCond[87] = UnbiasedRNG[87];
            InitCond[88] = UnbiasedRNG[88];
            InitCond[89] = UnbiasedRNG[89];
            InitCond[90] = UnbiasedRNG[90];
            InitCond[91] = UnbiasedRNG[91];
            InitCond[92] = UnbiasedRNG[92];
            InitCond[93] = UnbiasedRNG[93];
            InitCond[94] = UnbiasedRNG[94];
            InitCond[95] = UnbiasedRNG[95];
            InitCond[96] = UnbiasedRNG[96];
            InitCond[97] = UnbiasedRNG[97];
            InitCond[98] = UnbiasedRNG[98];
            InitCond[99] = UnbiasedRNG[99];
            InitCond[100] = UnbiasedRNG[100];
            InitCond[101] = UnbiasedRNG[101];
            InitCond[102] = UnbiasedRNG[102];
            InitCond[103] = UnbiasedRNG[103];
            InitCond[104] = UnbiasedRNG[104];
            InitCond[105] = UnbiasedRNG[105];
            InitCond[106] = UnbiasedRNG[106];
            InitCond[107] = UnbiasedRNG[107];
            InitCond[108] = UnbiasedRNG[108];
            InitCond[109] = UnbiasedRNG[109];
            InitCond[110] = UnbiasedRNG[110];
            InitCond[111] = UnbiasedRNG[111];
            InitCond[112] = UnbiasedRNG[112];
            InitCond[113] = UnbiasedRNG[113];
            InitCond[114] = UnbiasedRNG[114];
            InitCond[115] = UnbiasedRNG[115];
            InitCond[116] = UnbiasedRNG[116];
            InitCond[117] = UnbiasedRNG[117];
            InitCond[118] = UnbiasedRNG[118];
            InitCond[119] = UnbiasedRNG[119];
            InitCond[120] = UnbiasedRNG[120];
            InitCond[121] = UnbiasedRNG[121];
            InitCond[122] = UnbiasedRNG[122];
            InitCond[123] = UnbiasedRNG[123];
            InitCond[124] = UnbiasedRNG[124];
            InitCond[125] = UnbiasedRNG[125];
            InitCond[126] = UnbiasedRNG[126];
            InitCond[127] = UnbiasedRNG[127];
            InitCond[128] = UnbiasedRNG[128];
            InitCond[129] = UnbiasedRNG[129];
            InitCond[130] = UnbiasedRNG[130];
            InitCond[131] = UnbiasedRNG[131];
            InitCond[132] = UnbiasedRNG[132];
            InitCond[133] = UnbiasedRNG[133];
            InitCond[134] = UnbiasedRNG[134];
            InitCond[135] = UnbiasedRNG[135];
            InitCond[136] = UnbiasedRNG[136];
            InitCond[137] = UnbiasedRNG[137];
            InitCond[138] = UnbiasedRNG[138];
            InitCond[139] = UnbiasedRNG[139];
            InitCond[140] = UnbiasedRNG[140];
            InitCond[141] = UnbiasedRNG[141];
            InitCond[142] = UnbiasedRNG[142];
            InitCond[143] = UnbiasedRNG[143];
            InitCond[144] = UnbiasedRNG[144];
            InitCond[145] = UnbiasedRNG[145];
            InitCond[146] = UnbiasedRNG[146];
            InitCond[147] = UnbiasedRNG[147];
            InitCond[148] = UnbiasedRNG[148];
            InitCond[149] = UnbiasedRNG[149];
            InitCond[150] = UnbiasedRNG[150];
            InitCond[151] = UnbiasedRNG[151];
            InitCond[152] = UnbiasedRNG[152];
            InitCond[153] = UnbiasedRNG[153];
            InitCond[154] = UnbiasedRNG[154];
            InitCond[155] = UnbiasedRNG[155];
            InitCond[156] = UnbiasedRNG[156];
            InitCond[157] = UnbiasedRNG[157];
            InitCond[158] = UnbiasedRNG[158];
            InitCond[159] = UnbiasedRNG[159];
            InitCond[160] = UnbiasedRNG[160];
            InitCond[161] = UnbiasedRNG[161];
            InitCond[162] = UnbiasedRNG[162];
            InitCond[163] = UnbiasedRNG[163];
            InitCond[164] = UnbiasedRNG[164];
            InitCond[165] = UnbiasedRNG[165];
            InitCond[166] = UnbiasedRNG[166];
            InitCond[167] = UnbiasedRNG[167];
            InitCond[168] = UnbiasedRNG[168];
            InitCond[169] = UnbiasedRNG[169];
            InitCond[170] = UnbiasedRNG[170];
            InitCond[171] = UnbiasedRNG[171];
            InitCond[172] = UnbiasedRNG[172];
            InitCond[173] = UnbiasedRNG[173];
            InitCond[174] = UnbiasedRNG[174];
            InitCond[175] = UnbiasedRNG[175];
            InitCond[176] = UnbiasedRNG[176];
            InitCond[177] = UnbiasedRNG[177];
            InitCond[178] = UnbiasedRNG[178];
            InitCond[179] = UnbiasedRNG[179];
            InitCond[180] = UnbiasedRNG[180];
            InitCond[181] = UnbiasedRNG[181];
            InitCond[182] = UnbiasedRNG[182];
            InitCond[183] = UnbiasedRNG[183];
            InitCond[184] = UnbiasedRNG[184];
            InitCond[185] = UnbiasedRNG[185];
            InitCond[186] = UnbiasedRNG[186];
            InitCond[187] = UnbiasedRNG[187];
            InitCond[188] = UnbiasedRNG[188];
            InitCond[189] = UnbiasedRNG[189];
            InitCond[190] = UnbiasedRNG[190];
            InitCond[191] = UnbiasedRNG[191];
            InitCond[192] = UnbiasedRNG[192];
            InitCond[193] = UnbiasedRNG[193];
            InitCond[194] = UnbiasedRNG[194];
            InitCond[195] = UnbiasedRNG[195];
            InitCond[196] = UnbiasedRNG[196];
            InitCond[197] = UnbiasedRNG[197];
            InitCond[198] = UnbiasedRNG[198];
            InitCond[199] = UnbiasedRNG[199];
            InitCond[200] = UnbiasedRNG[200];
            InitCond[201] = UnbiasedRNG[201];
            InitCond[202] = UnbiasedRNG[202];
            InitCond[203] = UnbiasedRNG[203];
            InitCond[204] = UnbiasedRNG[204];
            InitCond[205] = UnbiasedRNG[205];
            InitCond[206] = UnbiasedRNG[206];
            InitCond[207] = UnbiasedRNG[207];
            InitCond[208] = UnbiasedRNG[208];
            InitCond[209] = UnbiasedRNG[209];
            InitCond[210] = UnbiasedRNG[210];
            InitCond[211] = UnbiasedRNG[211];
            InitCond[212] = UnbiasedRNG[212];
            InitCond[213] = UnbiasedRNG[213];
            InitCond[214] = UnbiasedRNG[214];
            InitCond[215] = UnbiasedRNG[215];
            InitCond[216] = UnbiasedRNG[216];
            InitCond[217] = UnbiasedRNG[217];
        end
        else if (counter == 2) begin
            InitCond[218] = UnbiasedRNG[0];
            InitCond[219] = UnbiasedRNG[1];
            InitCond[220] = UnbiasedRNG[2];
            InitCond[221] = UnbiasedRNG[3];
            InitCond[222] = UnbiasedRNG[4];
            InitCond[223] = UnbiasedRNG[5];
            InitCond[224] = UnbiasedRNG[6];
            InitCond[225] = UnbiasedRNG[7];
            InitCond[226] = UnbiasedRNG[8];
            InitCond[227] = UnbiasedRNG[9];
            InitCond[228] = UnbiasedRNG[10];
            InitCond[229] = UnbiasedRNG[11];
            InitCond[230] = UnbiasedRNG[12];
            InitCond[231] = UnbiasedRNG[13];
            InitCond[232] = UnbiasedRNG[14];
            InitCond[233] = UnbiasedRNG[15];
            InitCond[234] = UnbiasedRNG[16];
            InitCond[235] = UnbiasedRNG[17];
            InitCond[236] = UnbiasedRNG[18];
            InitCond[237] = UnbiasedRNG[19];
            InitCond[238] = UnbiasedRNG[20];
            InitCond[239] = UnbiasedRNG[21];
            InitCond[240] = UnbiasedRNG[22];
            InitCond[241] = UnbiasedRNG[23];
            InitCond[242] = UnbiasedRNG[24];
            InitCond[243] = UnbiasedRNG[25];
            InitCond[244] = UnbiasedRNG[26];
            InitCond[245] = UnbiasedRNG[27];
            InitCond[246] = UnbiasedRNG[28];
            InitCond[247] = UnbiasedRNG[29];
            InitCond[248] = UnbiasedRNG[30];
            InitCond[249] = UnbiasedRNG[31];
            InitCond[250] = UnbiasedRNG[32];
            InitCond[251] = UnbiasedRNG[33];
            InitCond[252] = UnbiasedRNG[34];
            InitCond[253] = UnbiasedRNG[35];
            InitCond[254] = UnbiasedRNG[36];
            InitCond[255] = UnbiasedRNG[37];
            InitCond[256] = UnbiasedRNG[38];
            InitCond[257] = UnbiasedRNG[39];
            InitCond[258] = UnbiasedRNG[40];
            InitCond[259] = UnbiasedRNG[41];
            InitCond[260] = UnbiasedRNG[42];
            InitCond[261] = UnbiasedRNG[43];
            InitCond[262] = UnbiasedRNG[44];
            InitCond[263] = UnbiasedRNG[45];
            InitCond[264] = UnbiasedRNG[46];
            InitCond[265] = UnbiasedRNG[47];
            InitCond[266] = UnbiasedRNG[48];
            InitCond[267] = UnbiasedRNG[49];
            InitCond[268] = UnbiasedRNG[50];
            InitCond[269] = UnbiasedRNG[51];
            InitCond[270] = UnbiasedRNG[52];
            InitCond[271] = UnbiasedRNG[53];
            InitCond[272] = UnbiasedRNG[54];
            InitCond[273] = UnbiasedRNG[55];
            InitCond[274] = UnbiasedRNG[56];
            InitCond[275] = UnbiasedRNG[57];
            InitCond[276] = UnbiasedRNG[58];
            InitCond[277] = UnbiasedRNG[59];
            InitCond[278] = UnbiasedRNG[60];
            InitCond[279] = UnbiasedRNG[61];
            InitCond[280] = UnbiasedRNG[62];
            InitCond[281] = UnbiasedRNG[63];
            InitCond[282] = UnbiasedRNG[64];
            InitCond[283] = UnbiasedRNG[65];
            InitCond[284] = UnbiasedRNG[66];
            InitCond[285] = UnbiasedRNG[67];
            InitCond[286] = UnbiasedRNG[68];
            InitCond[287] = UnbiasedRNG[69];
            InitCond[288] = UnbiasedRNG[70];
            InitCond[289] = UnbiasedRNG[71];
            InitCond[290] = UnbiasedRNG[72];
            InitCond[291] = UnbiasedRNG[73];
            InitCond[292] = UnbiasedRNG[74];
            InitCond[293] = UnbiasedRNG[75];
            InitCond[294] = UnbiasedRNG[76];
            InitCond[295] = UnbiasedRNG[77];
            InitCond[296] = UnbiasedRNG[78];
            InitCond[297] = UnbiasedRNG[79];
            InitCond[298] = UnbiasedRNG[80];
            InitCond[299] = UnbiasedRNG[81];
            InitCond[300] = UnbiasedRNG[82];
            InitCond[301] = UnbiasedRNG[83];
            InitCond[302] = UnbiasedRNG[84];
            InitCond[303] = UnbiasedRNG[85];
            InitCond[304] = UnbiasedRNG[86];
            InitCond[305] = UnbiasedRNG[87];
            InitCond[306] = UnbiasedRNG[88];
            InitCond[307] = UnbiasedRNG[89];
            InitCond[308] = UnbiasedRNG[90];
            InitCond[309] = UnbiasedRNG[91];
            InitCond[310] = UnbiasedRNG[92];
            InitCond[311] = UnbiasedRNG[93];
            InitCond[312] = UnbiasedRNG[94];
            InitCond[313] = UnbiasedRNG[95];
            InitCond[314] = UnbiasedRNG[96];
            InitCond[315] = UnbiasedRNG[97];
            InitCond[316] = UnbiasedRNG[98];
            InitCond[317] = UnbiasedRNG[99];
            InitCond[318] = UnbiasedRNG[100];
            InitCond[319] = UnbiasedRNG[101];
            InitCond[320] = UnbiasedRNG[102];
            InitCond[321] = UnbiasedRNG[103];
            InitCond[322] = UnbiasedRNG[104];
            InitCond[323] = UnbiasedRNG[105];
            InitCond[324] = UnbiasedRNG[106];
            InitCond[325] = UnbiasedRNG[107];
            InitCond[326] = UnbiasedRNG[108];
            InitCond[327] = UnbiasedRNG[109];
            InitCond[328] = UnbiasedRNG[110];
            InitCond[329] = UnbiasedRNG[111];
            InitCond[330] = UnbiasedRNG[112];
            InitCond[331] = UnbiasedRNG[113];
            InitCond[332] = UnbiasedRNG[114];
            InitCond[333] = UnbiasedRNG[115];
            InitCond[334] = UnbiasedRNG[116];
            InitCond[335] = UnbiasedRNG[117];
            InitCond[336] = UnbiasedRNG[118];
            InitCond[337] = UnbiasedRNG[119];
            InitCond[338] = UnbiasedRNG[120];
            InitCond[339] = UnbiasedRNG[121];
            InitCond[340] = UnbiasedRNG[122];
            InitCond[341] = UnbiasedRNG[123];
            InitCond[342] = UnbiasedRNG[124];
            InitCond[343] = UnbiasedRNG[125];
            InitCond[344] = UnbiasedRNG[126];
            InitCond[345] = UnbiasedRNG[127];
            InitCond[346] = UnbiasedRNG[128];
            InitCond[347] = UnbiasedRNG[129];
            InitCond[348] = UnbiasedRNG[130];
            InitCond[349] = UnbiasedRNG[131];
            InitCond[350] = UnbiasedRNG[132];
            InitCond[351] = UnbiasedRNG[133];
            InitCond[352] = UnbiasedRNG[134];
            InitCond[353] = UnbiasedRNG[135];
            InitCond[354] = UnbiasedRNG[136];
            InitCond[355] = UnbiasedRNG[137];
            InitCond[356] = UnbiasedRNG[138];
            InitCond[357] = UnbiasedRNG[139];
            InitCond[358] = UnbiasedRNG[140];
            InitCond[359] = UnbiasedRNG[141];
            InitCond[360] = UnbiasedRNG[142];
            InitCond[361] = UnbiasedRNG[143];
            InitCond[362] = UnbiasedRNG[144];
            InitCond[363] = UnbiasedRNG[145];
            InitCond[364] = UnbiasedRNG[146];
            InitCond[365] = UnbiasedRNG[147];
            InitCond[366] = UnbiasedRNG[148];
            InitCond[367] = UnbiasedRNG[149];
            InitCond[368] = UnbiasedRNG[150];
            InitCond[369] = UnbiasedRNG[151];
            InitCond[370] = UnbiasedRNG[152];
            InitCond[371] = UnbiasedRNG[153];
            InitCond[372] = UnbiasedRNG[154];
            InitCond[373] = UnbiasedRNG[155];
            InitCond[374] = UnbiasedRNG[156];
            InitCond[375] = UnbiasedRNG[157];
            InitCond[376] = UnbiasedRNG[158];
            InitCond[377] = UnbiasedRNG[159];
            InitCond[378] = UnbiasedRNG[160];
            InitCond[379] = UnbiasedRNG[161];
            InitCond[380] = UnbiasedRNG[162];
            InitCond[381] = UnbiasedRNG[163];
            InitCond[382] = UnbiasedRNG[164];
            InitCond[383] = UnbiasedRNG[165];
            InitCond[384] = UnbiasedRNG[166];
            InitCond[385] = UnbiasedRNG[167];
            InitCond[386] = UnbiasedRNG[168];
            InitCond[387] = UnbiasedRNG[169];
            InitCond[388] = UnbiasedRNG[170];
            InitCond[389] = UnbiasedRNG[171];
            InitCond[390] = UnbiasedRNG[172];
            InitCond[391] = UnbiasedRNG[173];
            InitCond[392] = UnbiasedRNG[174];
            InitCond[393] = UnbiasedRNG[175];
            InitCond[394] = UnbiasedRNG[176];
            InitCond[395] = UnbiasedRNG[177];
            InitCond[396] = UnbiasedRNG[178];
            InitCond[397] = UnbiasedRNG[179];
            InitCond[398] = UnbiasedRNG[180];
            InitCond[399] = UnbiasedRNG[181];
            InitCond[400] = UnbiasedRNG[182];
            InitCond[401] = UnbiasedRNG[183];
            InitCond[402] = UnbiasedRNG[184];
            InitCond[403] = UnbiasedRNG[185];
            InitCond[404] = UnbiasedRNG[186];
            InitCond[405] = UnbiasedRNG[187];
            InitCond[406] = UnbiasedRNG[188];
            InitCond[407] = UnbiasedRNG[189];
            InitCond[408] = UnbiasedRNG[190];
            InitCond[409] = UnbiasedRNG[191];
            InitCond[410] = UnbiasedRNG[192];
            InitCond[411] = UnbiasedRNG[193];
            InitCond[412] = UnbiasedRNG[194];
            InitCond[413] = UnbiasedRNG[195];
            InitCond[414] = UnbiasedRNG[196];
            InitCond[415] = UnbiasedRNG[197];
            InitCond[416] = UnbiasedRNG[198];
            InitCond[417] = UnbiasedRNG[199];
            InitCond[418] = UnbiasedRNG[200];
            InitCond[419] = UnbiasedRNG[201];
            InitCond[420] = UnbiasedRNG[202];
            InitCond[421] = UnbiasedRNG[203];
            InitCond[422] = UnbiasedRNG[204];
            InitCond[423] = UnbiasedRNG[205];
            InitCond[424] = UnbiasedRNG[206];
            InitCond[425] = UnbiasedRNG[207];
            InitCond[426] = UnbiasedRNG[208];
            InitCond[427] = UnbiasedRNG[209];
            InitCond[428] = UnbiasedRNG[210];
            InitCond[429] = UnbiasedRNG[211];
            InitCond[430] = UnbiasedRNG[212];
            InitCond[431] = UnbiasedRNG[213];
            InitCond[432] = UnbiasedRNG[214];
            InitCond[433] = UnbiasedRNG[215];
            InitCond[434] = UnbiasedRNG[216];
            InitCond[435] = UnbiasedRNG[217];
        end
        else if (counter == 3) begin
            InitCond[436] = UnbiasedRNG[0];
            InitCond[437] = UnbiasedRNG[1];
            InitCond[438] = UnbiasedRNG[2];
            InitCond[439] = UnbiasedRNG[3];
            InitCond[440] = UnbiasedRNG[4];
            InitCond[441] = UnbiasedRNG[5];
            InitCond[442] = UnbiasedRNG[6];
            InitCond[443] = UnbiasedRNG[7];
            InitCond[444] = UnbiasedRNG[8];
            InitCond[445] = UnbiasedRNG[9];
            InitCond[446] = UnbiasedRNG[10];
            InitCond[447] = UnbiasedRNG[11];
            InitCond[448] = UnbiasedRNG[12];
            InitCond[449] = UnbiasedRNG[13];
            InitCond[450] = UnbiasedRNG[14];
            InitCond[451] = UnbiasedRNG[15];
            InitCond[452] = UnbiasedRNG[16];
            InitCond[453] = UnbiasedRNG[17];
            InitCond[454] = UnbiasedRNG[18];
            InitCond[455] = UnbiasedRNG[19];
            InitCond[456] = UnbiasedRNG[20];
            InitCond[457] = UnbiasedRNG[21];
            InitCond[458] = UnbiasedRNG[22];
            InitCond[459] = UnbiasedRNG[23];
            InitCond[460] = UnbiasedRNG[24];
            InitCond[461] = UnbiasedRNG[25];
            InitCond[462] = UnbiasedRNG[26];
            InitCond[463] = UnbiasedRNG[27];
            InitCond[464] = UnbiasedRNG[28];
            InitCond[465] = UnbiasedRNG[29];
            InitCond[466] = UnbiasedRNG[30];
            InitCond[467] = UnbiasedRNG[31];
            InitCond[468] = UnbiasedRNG[32];
            InitCond[469] = UnbiasedRNG[33];
            InitCond[470] = UnbiasedRNG[34];
            InitCond[471] = UnbiasedRNG[35];
            InitCond[472] = UnbiasedRNG[36];
            InitCond[473] = UnbiasedRNG[37];
            InitCond[474] = UnbiasedRNG[38];
            InitCond[475] = UnbiasedRNG[39];
            InitCond[476] = UnbiasedRNG[40];
            InitCond[477] = UnbiasedRNG[41];
            InitCond[478] = UnbiasedRNG[42];
            InitCond[479] = UnbiasedRNG[43];
            InitCond[480] = UnbiasedRNG[44];
            InitCond[481] = UnbiasedRNG[45];
            InitCond[482] = UnbiasedRNG[46];
            InitCond[483] = UnbiasedRNG[47];
            InitCond[484] = UnbiasedRNG[48];
            InitCond[485] = UnbiasedRNG[49];
            InitCond[486] = UnbiasedRNG[50];
            InitCond[487] = UnbiasedRNG[51];
            InitCond[488] = UnbiasedRNG[52];
            InitCond[489] = UnbiasedRNG[53];
            InitCond[490] = UnbiasedRNG[54];
            InitCond[491] = UnbiasedRNG[55];
            InitCond[492] = UnbiasedRNG[56];
            InitCond[493] = UnbiasedRNG[57];
            InitCond[494] = UnbiasedRNG[58];
            InitCond[495] = UnbiasedRNG[59];
        end
        else if (counter==5)
            run = 1'b1;
        counter = counter+38'b1;
        solution = {m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[15],m[14],m[13],m[12],m[11],m[10],m[9],m[8]};
    end else begin 
        counter = 38'b0;
        failure = 1'b1;
        run = 1'b0;
    end
end

//To measure on only the last step using ILA:
always @(negedge sample_clk) begin
    if (solution_flag)
        solution_flag = 1'b0;
    else if ((run & (solution == solution_check)) | failure)
        solution_flag = 1'b1;
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = run?((((m[16]&~m[17])|(~m[16]&m[17]))&UnbiasedRNG[0])|((m[16]&m[17]))):InitCond[0];
    m[1] = run?((((m[18]&~m[19])|(~m[18]&m[19]))&UnbiasedRNG[1])|((m[18]&m[19]))):InitCond[1];
    m[2] = run?((((m[20]&~m[21])|(~m[20]&m[21]))&UnbiasedRNG[2])|((m[20]&m[21]))):InitCond[2];
    m[3] = run?((((m[22]&~m[23])|(~m[22]&m[23]))&UnbiasedRNG[3])|((m[22]&m[23]))):InitCond[3];
    m[4] = run?((((m[24]&~m[25])|(~m[24]&m[25]))&UnbiasedRNG[4])|((m[24]&m[25]))):InitCond[4];
    m[5] = run?((((m[26]&~m[27])|(~m[26]&m[27]))&UnbiasedRNG[5])|((m[26]&m[27]))):InitCond[5];
    m[6] = run?((((m[28]&~m[29])|(~m[28]&m[29]))&UnbiasedRNG[6])|((m[28]&m[29]))):InitCond[6];
    m[7] = run?((((m[30]&~m[31])|(~m[30]&m[31]))&UnbiasedRNG[7])|((m[30]&m[31]))):InitCond[7];
    m[8] = run?((((m[32]&~m[33])|(~m[32]&m[33]))&UnbiasedRNG[8])|((m[32]&m[33]))):InitCond[8];
    m[9] = run?((((m[34]&~m[35])|(~m[34]&m[35]))&UnbiasedRNG[9])|((m[34]&m[35]))):InitCond[9];
    m[10] = run?((((m[36]&~m[37])|(~m[36]&m[37]))&UnbiasedRNG[10])|((m[36]&m[37]))):InitCond[10];
    m[11] = run?((((m[38]&~m[39])|(~m[38]&m[39]))&UnbiasedRNG[11])|((m[38]&m[39]))):InitCond[11];
    m[12] = run?((((m[40]&~m[41])|(~m[40]&m[41]))&UnbiasedRNG[12])|((m[40]&m[41]))):InitCond[12];
    m[13] = run?((((m[42]&~m[43])|(~m[42]&m[43]))&UnbiasedRNG[13])|((m[42]&m[43]))):InitCond[13];
    m[14] = run?((((m[44]&~m[45])|(~m[44]&m[45]))&UnbiasedRNG[14])|((m[44]&m[45]))):InitCond[14];
    m[15] = run?((((m[46]&~m[47])|(~m[46]&m[47]))&UnbiasedRNG[15])|((m[46]&m[47]))):InitCond[15];
    m[48] = run?((((~m[16]&~m[112]&~m[176])|(m[16]&m[112]&~m[176]))&BiasedRNG[0])|(((m[16]&~m[112]&~m[176])|(~m[16]&m[112]&m[176]))&~BiasedRNG[0])|((~m[16]&~m[112]&m[176])|(m[16]&~m[112]&m[176])|(m[16]&m[112]&m[176]))):InitCond[16];
    m[49] = run?((((~m[16]&~m[120]&~m[184])|(m[16]&m[120]&~m[184]))&BiasedRNG[1])|(((m[16]&~m[120]&~m[184])|(~m[16]&m[120]&m[184]))&~BiasedRNG[1])|((~m[16]&~m[120]&m[184])|(m[16]&~m[120]&m[184])|(m[16]&m[120]&m[184]))):InitCond[17];
    m[50] = run?((((~m[16]&~m[128]&~m[192])|(m[16]&m[128]&~m[192]))&BiasedRNG[2])|(((m[16]&~m[128]&~m[192])|(~m[16]&m[128]&m[192]))&~BiasedRNG[2])|((~m[16]&~m[128]&m[192])|(m[16]&~m[128]&m[192])|(m[16]&m[128]&m[192]))):InitCond[18];
    m[51] = run?((((~m[16]&~m[136]&~m[200])|(m[16]&m[136]&~m[200]))&BiasedRNG[3])|(((m[16]&~m[136]&~m[200])|(~m[16]&m[136]&m[200]))&~BiasedRNG[3])|((~m[16]&~m[136]&m[200])|(m[16]&~m[136]&m[200])|(m[16]&m[136]&m[200]))):InitCond[19];
    m[52] = run?((((~m[17]&~m[144]&~m[208])|(m[17]&m[144]&~m[208]))&BiasedRNG[4])|(((m[17]&~m[144]&~m[208])|(~m[17]&m[144]&m[208]))&~BiasedRNG[4])|((~m[17]&~m[144]&m[208])|(m[17]&~m[144]&m[208])|(m[17]&m[144]&m[208]))):InitCond[20];
    m[53] = run?((((~m[17]&~m[152]&~m[216])|(m[17]&m[152]&~m[216]))&BiasedRNG[5])|(((m[17]&~m[152]&~m[216])|(~m[17]&m[152]&m[216]))&~BiasedRNG[5])|((~m[17]&~m[152]&m[216])|(m[17]&~m[152]&m[216])|(m[17]&m[152]&m[216]))):InitCond[21];
    m[54] = run?((((~m[17]&~m[160]&~m[224])|(m[17]&m[160]&~m[224]))&BiasedRNG[6])|(((m[17]&~m[160]&~m[224])|(~m[17]&m[160]&m[224]))&~BiasedRNG[6])|((~m[17]&~m[160]&m[224])|(m[17]&~m[160]&m[224])|(m[17]&m[160]&m[224]))):InitCond[22];
    m[55] = run?((((~m[17]&~m[168]&~m[232])|(m[17]&m[168]&~m[232]))&BiasedRNG[7])|(((m[17]&~m[168]&~m[232])|(~m[17]&m[168]&m[232]))&~BiasedRNG[7])|((~m[17]&~m[168]&m[232])|(m[17]&~m[168]&m[232])|(m[17]&m[168]&m[232]))):InitCond[23];
    m[56] = run?((((~m[18]&~m[113]&~m[177])|(m[18]&m[113]&~m[177]))&BiasedRNG[8])|(((m[18]&~m[113]&~m[177])|(~m[18]&m[113]&m[177]))&~BiasedRNG[8])|((~m[18]&~m[113]&m[177])|(m[18]&~m[113]&m[177])|(m[18]&m[113]&m[177]))):InitCond[24];
    m[57] = run?((((~m[18]&~m[121]&~m[185])|(m[18]&m[121]&~m[185]))&BiasedRNG[9])|(((m[18]&~m[121]&~m[185])|(~m[18]&m[121]&m[185]))&~BiasedRNG[9])|((~m[18]&~m[121]&m[185])|(m[18]&~m[121]&m[185])|(m[18]&m[121]&m[185]))):InitCond[25];
    m[58] = run?((((~m[18]&~m[129]&~m[193])|(m[18]&m[129]&~m[193]))&BiasedRNG[10])|(((m[18]&~m[129]&~m[193])|(~m[18]&m[129]&m[193]))&~BiasedRNG[10])|((~m[18]&~m[129]&m[193])|(m[18]&~m[129]&m[193])|(m[18]&m[129]&m[193]))):InitCond[26];
    m[59] = run?((((~m[18]&~m[137]&~m[201])|(m[18]&m[137]&~m[201]))&BiasedRNG[11])|(((m[18]&~m[137]&~m[201])|(~m[18]&m[137]&m[201]))&~BiasedRNG[11])|((~m[18]&~m[137]&m[201])|(m[18]&~m[137]&m[201])|(m[18]&m[137]&m[201]))):InitCond[27];
    m[60] = run?((((~m[19]&~m[145]&~m[209])|(m[19]&m[145]&~m[209]))&BiasedRNG[12])|(((m[19]&~m[145]&~m[209])|(~m[19]&m[145]&m[209]))&~BiasedRNG[12])|((~m[19]&~m[145]&m[209])|(m[19]&~m[145]&m[209])|(m[19]&m[145]&m[209]))):InitCond[28];
    m[61] = run?((((~m[19]&~m[153]&~m[217])|(m[19]&m[153]&~m[217]))&BiasedRNG[13])|(((m[19]&~m[153]&~m[217])|(~m[19]&m[153]&m[217]))&~BiasedRNG[13])|((~m[19]&~m[153]&m[217])|(m[19]&~m[153]&m[217])|(m[19]&m[153]&m[217]))):InitCond[29];
    m[62] = run?((((~m[19]&~m[161]&~m[225])|(m[19]&m[161]&~m[225]))&BiasedRNG[14])|(((m[19]&~m[161]&~m[225])|(~m[19]&m[161]&m[225]))&~BiasedRNG[14])|((~m[19]&~m[161]&m[225])|(m[19]&~m[161]&m[225])|(m[19]&m[161]&m[225]))):InitCond[30];
    m[63] = run?((((~m[19]&~m[169]&~m[233])|(m[19]&m[169]&~m[233]))&BiasedRNG[15])|(((m[19]&~m[169]&~m[233])|(~m[19]&m[169]&m[233]))&~BiasedRNG[15])|((~m[19]&~m[169]&m[233])|(m[19]&~m[169]&m[233])|(m[19]&m[169]&m[233]))):InitCond[31];
    m[64] = run?((((~m[20]&~m[114]&~m[178])|(m[20]&m[114]&~m[178]))&BiasedRNG[16])|(((m[20]&~m[114]&~m[178])|(~m[20]&m[114]&m[178]))&~BiasedRNG[16])|((~m[20]&~m[114]&m[178])|(m[20]&~m[114]&m[178])|(m[20]&m[114]&m[178]))):InitCond[32];
    m[65] = run?((((~m[20]&~m[122]&~m[186])|(m[20]&m[122]&~m[186]))&BiasedRNG[17])|(((m[20]&~m[122]&~m[186])|(~m[20]&m[122]&m[186]))&~BiasedRNG[17])|((~m[20]&~m[122]&m[186])|(m[20]&~m[122]&m[186])|(m[20]&m[122]&m[186]))):InitCond[33];
    m[66] = run?((((~m[20]&~m[130]&~m[194])|(m[20]&m[130]&~m[194]))&BiasedRNG[18])|(((m[20]&~m[130]&~m[194])|(~m[20]&m[130]&m[194]))&~BiasedRNG[18])|((~m[20]&~m[130]&m[194])|(m[20]&~m[130]&m[194])|(m[20]&m[130]&m[194]))):InitCond[34];
    m[67] = run?((((~m[20]&~m[138]&~m[202])|(m[20]&m[138]&~m[202]))&BiasedRNG[19])|(((m[20]&~m[138]&~m[202])|(~m[20]&m[138]&m[202]))&~BiasedRNG[19])|((~m[20]&~m[138]&m[202])|(m[20]&~m[138]&m[202])|(m[20]&m[138]&m[202]))):InitCond[35];
    m[68] = run?((((~m[21]&~m[146]&~m[210])|(m[21]&m[146]&~m[210]))&BiasedRNG[20])|(((m[21]&~m[146]&~m[210])|(~m[21]&m[146]&m[210]))&~BiasedRNG[20])|((~m[21]&~m[146]&m[210])|(m[21]&~m[146]&m[210])|(m[21]&m[146]&m[210]))):InitCond[36];
    m[69] = run?((((~m[21]&~m[154]&~m[218])|(m[21]&m[154]&~m[218]))&BiasedRNG[21])|(((m[21]&~m[154]&~m[218])|(~m[21]&m[154]&m[218]))&~BiasedRNG[21])|((~m[21]&~m[154]&m[218])|(m[21]&~m[154]&m[218])|(m[21]&m[154]&m[218]))):InitCond[37];
    m[70] = run?((((~m[21]&~m[162]&~m[226])|(m[21]&m[162]&~m[226]))&BiasedRNG[22])|(((m[21]&~m[162]&~m[226])|(~m[21]&m[162]&m[226]))&~BiasedRNG[22])|((~m[21]&~m[162]&m[226])|(m[21]&~m[162]&m[226])|(m[21]&m[162]&m[226]))):InitCond[38];
    m[71] = run?((((~m[21]&~m[170]&~m[234])|(m[21]&m[170]&~m[234]))&BiasedRNG[23])|(((m[21]&~m[170]&~m[234])|(~m[21]&m[170]&m[234]))&~BiasedRNG[23])|((~m[21]&~m[170]&m[234])|(m[21]&~m[170]&m[234])|(m[21]&m[170]&m[234]))):InitCond[39];
    m[72] = run?((((~m[22]&~m[115]&~m[179])|(m[22]&m[115]&~m[179]))&BiasedRNG[24])|(((m[22]&~m[115]&~m[179])|(~m[22]&m[115]&m[179]))&~BiasedRNG[24])|((~m[22]&~m[115]&m[179])|(m[22]&~m[115]&m[179])|(m[22]&m[115]&m[179]))):InitCond[40];
    m[73] = run?((((~m[22]&~m[123]&~m[187])|(m[22]&m[123]&~m[187]))&BiasedRNG[25])|(((m[22]&~m[123]&~m[187])|(~m[22]&m[123]&m[187]))&~BiasedRNG[25])|((~m[22]&~m[123]&m[187])|(m[22]&~m[123]&m[187])|(m[22]&m[123]&m[187]))):InitCond[41];
    m[74] = run?((((~m[22]&~m[131]&~m[195])|(m[22]&m[131]&~m[195]))&BiasedRNG[26])|(((m[22]&~m[131]&~m[195])|(~m[22]&m[131]&m[195]))&~BiasedRNG[26])|((~m[22]&~m[131]&m[195])|(m[22]&~m[131]&m[195])|(m[22]&m[131]&m[195]))):InitCond[42];
    m[75] = run?((((~m[22]&~m[139]&~m[203])|(m[22]&m[139]&~m[203]))&BiasedRNG[27])|(((m[22]&~m[139]&~m[203])|(~m[22]&m[139]&m[203]))&~BiasedRNG[27])|((~m[22]&~m[139]&m[203])|(m[22]&~m[139]&m[203])|(m[22]&m[139]&m[203]))):InitCond[43];
    m[76] = run?((((~m[23]&~m[147]&~m[211])|(m[23]&m[147]&~m[211]))&BiasedRNG[28])|(((m[23]&~m[147]&~m[211])|(~m[23]&m[147]&m[211]))&~BiasedRNG[28])|((~m[23]&~m[147]&m[211])|(m[23]&~m[147]&m[211])|(m[23]&m[147]&m[211]))):InitCond[44];
    m[77] = run?((((~m[23]&~m[155]&~m[219])|(m[23]&m[155]&~m[219]))&BiasedRNG[29])|(((m[23]&~m[155]&~m[219])|(~m[23]&m[155]&m[219]))&~BiasedRNG[29])|((~m[23]&~m[155]&m[219])|(m[23]&~m[155]&m[219])|(m[23]&m[155]&m[219]))):InitCond[45];
    m[78] = run?((((~m[23]&~m[163]&~m[227])|(m[23]&m[163]&~m[227]))&BiasedRNG[30])|(((m[23]&~m[163]&~m[227])|(~m[23]&m[163]&m[227]))&~BiasedRNG[30])|((~m[23]&~m[163]&m[227])|(m[23]&~m[163]&m[227])|(m[23]&m[163]&m[227]))):InitCond[46];
    m[79] = run?((((~m[23]&~m[171]&~m[235])|(m[23]&m[171]&~m[235]))&BiasedRNG[31])|(((m[23]&~m[171]&~m[235])|(~m[23]&m[171]&m[235]))&~BiasedRNG[31])|((~m[23]&~m[171]&m[235])|(m[23]&~m[171]&m[235])|(m[23]&m[171]&m[235]))):InitCond[47];
    m[80] = run?((((~m[24]&~m[116]&~m[180])|(m[24]&m[116]&~m[180]))&BiasedRNG[32])|(((m[24]&~m[116]&~m[180])|(~m[24]&m[116]&m[180]))&~BiasedRNG[32])|((~m[24]&~m[116]&m[180])|(m[24]&~m[116]&m[180])|(m[24]&m[116]&m[180]))):InitCond[48];
    m[81] = run?((((~m[24]&~m[124]&~m[188])|(m[24]&m[124]&~m[188]))&BiasedRNG[33])|(((m[24]&~m[124]&~m[188])|(~m[24]&m[124]&m[188]))&~BiasedRNG[33])|((~m[24]&~m[124]&m[188])|(m[24]&~m[124]&m[188])|(m[24]&m[124]&m[188]))):InitCond[49];
    m[82] = run?((((~m[24]&~m[132]&~m[196])|(m[24]&m[132]&~m[196]))&BiasedRNG[34])|(((m[24]&~m[132]&~m[196])|(~m[24]&m[132]&m[196]))&~BiasedRNG[34])|((~m[24]&~m[132]&m[196])|(m[24]&~m[132]&m[196])|(m[24]&m[132]&m[196]))):InitCond[50];
    m[83] = run?((((~m[24]&~m[140]&~m[204])|(m[24]&m[140]&~m[204]))&BiasedRNG[35])|(((m[24]&~m[140]&~m[204])|(~m[24]&m[140]&m[204]))&~BiasedRNG[35])|((~m[24]&~m[140]&m[204])|(m[24]&~m[140]&m[204])|(m[24]&m[140]&m[204]))):InitCond[51];
    m[84] = run?((((~m[25]&~m[148]&~m[212])|(m[25]&m[148]&~m[212]))&BiasedRNG[36])|(((m[25]&~m[148]&~m[212])|(~m[25]&m[148]&m[212]))&~BiasedRNG[36])|((~m[25]&~m[148]&m[212])|(m[25]&~m[148]&m[212])|(m[25]&m[148]&m[212]))):InitCond[52];
    m[85] = run?((((~m[25]&~m[156]&~m[220])|(m[25]&m[156]&~m[220]))&BiasedRNG[37])|(((m[25]&~m[156]&~m[220])|(~m[25]&m[156]&m[220]))&~BiasedRNG[37])|((~m[25]&~m[156]&m[220])|(m[25]&~m[156]&m[220])|(m[25]&m[156]&m[220]))):InitCond[53];
    m[86] = run?((((~m[25]&~m[164]&~m[228])|(m[25]&m[164]&~m[228]))&BiasedRNG[38])|(((m[25]&~m[164]&~m[228])|(~m[25]&m[164]&m[228]))&~BiasedRNG[38])|((~m[25]&~m[164]&m[228])|(m[25]&~m[164]&m[228])|(m[25]&m[164]&m[228]))):InitCond[54];
    m[87] = run?((((~m[25]&~m[172]&~m[236])|(m[25]&m[172]&~m[236]))&BiasedRNG[39])|(((m[25]&~m[172]&~m[236])|(~m[25]&m[172]&m[236]))&~BiasedRNG[39])|((~m[25]&~m[172]&m[236])|(m[25]&~m[172]&m[236])|(m[25]&m[172]&m[236]))):InitCond[55];
    m[88] = run?((((~m[26]&~m[117]&~m[181])|(m[26]&m[117]&~m[181]))&BiasedRNG[40])|(((m[26]&~m[117]&~m[181])|(~m[26]&m[117]&m[181]))&~BiasedRNG[40])|((~m[26]&~m[117]&m[181])|(m[26]&~m[117]&m[181])|(m[26]&m[117]&m[181]))):InitCond[56];
    m[89] = run?((((~m[26]&~m[125]&~m[189])|(m[26]&m[125]&~m[189]))&BiasedRNG[41])|(((m[26]&~m[125]&~m[189])|(~m[26]&m[125]&m[189]))&~BiasedRNG[41])|((~m[26]&~m[125]&m[189])|(m[26]&~m[125]&m[189])|(m[26]&m[125]&m[189]))):InitCond[57];
    m[90] = run?((((~m[26]&~m[133]&~m[197])|(m[26]&m[133]&~m[197]))&BiasedRNG[42])|(((m[26]&~m[133]&~m[197])|(~m[26]&m[133]&m[197]))&~BiasedRNG[42])|((~m[26]&~m[133]&m[197])|(m[26]&~m[133]&m[197])|(m[26]&m[133]&m[197]))):InitCond[58];
    m[91] = run?((((~m[26]&~m[141]&~m[205])|(m[26]&m[141]&~m[205]))&BiasedRNG[43])|(((m[26]&~m[141]&~m[205])|(~m[26]&m[141]&m[205]))&~BiasedRNG[43])|((~m[26]&~m[141]&m[205])|(m[26]&~m[141]&m[205])|(m[26]&m[141]&m[205]))):InitCond[59];
    m[92] = run?((((~m[27]&~m[149]&~m[213])|(m[27]&m[149]&~m[213]))&BiasedRNG[44])|(((m[27]&~m[149]&~m[213])|(~m[27]&m[149]&m[213]))&~BiasedRNG[44])|((~m[27]&~m[149]&m[213])|(m[27]&~m[149]&m[213])|(m[27]&m[149]&m[213]))):InitCond[60];
    m[93] = run?((((~m[27]&~m[157]&~m[221])|(m[27]&m[157]&~m[221]))&BiasedRNG[45])|(((m[27]&~m[157]&~m[221])|(~m[27]&m[157]&m[221]))&~BiasedRNG[45])|((~m[27]&~m[157]&m[221])|(m[27]&~m[157]&m[221])|(m[27]&m[157]&m[221]))):InitCond[61];
    m[94] = run?((((~m[27]&~m[165]&~m[229])|(m[27]&m[165]&~m[229]))&BiasedRNG[46])|(((m[27]&~m[165]&~m[229])|(~m[27]&m[165]&m[229]))&~BiasedRNG[46])|((~m[27]&~m[165]&m[229])|(m[27]&~m[165]&m[229])|(m[27]&m[165]&m[229]))):InitCond[62];
    m[95] = run?((((~m[27]&~m[173]&~m[237])|(m[27]&m[173]&~m[237]))&BiasedRNG[47])|(((m[27]&~m[173]&~m[237])|(~m[27]&m[173]&m[237]))&~BiasedRNG[47])|((~m[27]&~m[173]&m[237])|(m[27]&~m[173]&m[237])|(m[27]&m[173]&m[237]))):InitCond[63];
    m[96] = run?((((~m[28]&~m[118]&~m[182])|(m[28]&m[118]&~m[182]))&BiasedRNG[48])|(((m[28]&~m[118]&~m[182])|(~m[28]&m[118]&m[182]))&~BiasedRNG[48])|((~m[28]&~m[118]&m[182])|(m[28]&~m[118]&m[182])|(m[28]&m[118]&m[182]))):InitCond[64];
    m[97] = run?((((~m[28]&~m[126]&~m[190])|(m[28]&m[126]&~m[190]))&BiasedRNG[49])|(((m[28]&~m[126]&~m[190])|(~m[28]&m[126]&m[190]))&~BiasedRNG[49])|((~m[28]&~m[126]&m[190])|(m[28]&~m[126]&m[190])|(m[28]&m[126]&m[190]))):InitCond[65];
    m[98] = run?((((~m[28]&~m[134]&~m[198])|(m[28]&m[134]&~m[198]))&BiasedRNG[50])|(((m[28]&~m[134]&~m[198])|(~m[28]&m[134]&m[198]))&~BiasedRNG[50])|((~m[28]&~m[134]&m[198])|(m[28]&~m[134]&m[198])|(m[28]&m[134]&m[198]))):InitCond[66];
    m[99] = run?((((~m[28]&~m[142]&~m[206])|(m[28]&m[142]&~m[206]))&BiasedRNG[51])|(((m[28]&~m[142]&~m[206])|(~m[28]&m[142]&m[206]))&~BiasedRNG[51])|((~m[28]&~m[142]&m[206])|(m[28]&~m[142]&m[206])|(m[28]&m[142]&m[206]))):InitCond[67];
    m[100] = run?((((~m[29]&~m[150]&~m[214])|(m[29]&m[150]&~m[214]))&BiasedRNG[52])|(((m[29]&~m[150]&~m[214])|(~m[29]&m[150]&m[214]))&~BiasedRNG[52])|((~m[29]&~m[150]&m[214])|(m[29]&~m[150]&m[214])|(m[29]&m[150]&m[214]))):InitCond[68];
    m[101] = run?((((~m[29]&~m[158]&~m[222])|(m[29]&m[158]&~m[222]))&BiasedRNG[53])|(((m[29]&~m[158]&~m[222])|(~m[29]&m[158]&m[222]))&~BiasedRNG[53])|((~m[29]&~m[158]&m[222])|(m[29]&~m[158]&m[222])|(m[29]&m[158]&m[222]))):InitCond[69];
    m[102] = run?((((~m[29]&~m[166]&~m[230])|(m[29]&m[166]&~m[230]))&BiasedRNG[54])|(((m[29]&~m[166]&~m[230])|(~m[29]&m[166]&m[230]))&~BiasedRNG[54])|((~m[29]&~m[166]&m[230])|(m[29]&~m[166]&m[230])|(m[29]&m[166]&m[230]))):InitCond[70];
    m[103] = run?((((~m[29]&~m[174]&~m[238])|(m[29]&m[174]&~m[238]))&BiasedRNG[55])|(((m[29]&~m[174]&~m[238])|(~m[29]&m[174]&m[238]))&~BiasedRNG[55])|((~m[29]&~m[174]&m[238])|(m[29]&~m[174]&m[238])|(m[29]&m[174]&m[238]))):InitCond[71];
    m[104] = run?((((~m[30]&~m[119]&~m[183])|(m[30]&m[119]&~m[183]))&BiasedRNG[56])|(((m[30]&~m[119]&~m[183])|(~m[30]&m[119]&m[183]))&~BiasedRNG[56])|((~m[30]&~m[119]&m[183])|(m[30]&~m[119]&m[183])|(m[30]&m[119]&m[183]))):InitCond[72];
    m[105] = run?((((~m[30]&~m[127]&~m[191])|(m[30]&m[127]&~m[191]))&BiasedRNG[57])|(((m[30]&~m[127]&~m[191])|(~m[30]&m[127]&m[191]))&~BiasedRNG[57])|((~m[30]&~m[127]&m[191])|(m[30]&~m[127]&m[191])|(m[30]&m[127]&m[191]))):InitCond[73];
    m[106] = run?((((~m[30]&~m[135]&~m[199])|(m[30]&m[135]&~m[199]))&BiasedRNG[58])|(((m[30]&~m[135]&~m[199])|(~m[30]&m[135]&m[199]))&~BiasedRNG[58])|((~m[30]&~m[135]&m[199])|(m[30]&~m[135]&m[199])|(m[30]&m[135]&m[199]))):InitCond[74];
    m[107] = run?((((~m[30]&~m[143]&~m[207])|(m[30]&m[143]&~m[207]))&BiasedRNG[59])|(((m[30]&~m[143]&~m[207])|(~m[30]&m[143]&m[207]))&~BiasedRNG[59])|((~m[30]&~m[143]&m[207])|(m[30]&~m[143]&m[207])|(m[30]&m[143]&m[207]))):InitCond[75];
    m[108] = run?((((~m[31]&~m[151]&~m[215])|(m[31]&m[151]&~m[215]))&BiasedRNG[60])|(((m[31]&~m[151]&~m[215])|(~m[31]&m[151]&m[215]))&~BiasedRNG[60])|((~m[31]&~m[151]&m[215])|(m[31]&~m[151]&m[215])|(m[31]&m[151]&m[215]))):InitCond[76];
    m[109] = run?((((~m[31]&~m[159]&~m[223])|(m[31]&m[159]&~m[223]))&BiasedRNG[61])|(((m[31]&~m[159]&~m[223])|(~m[31]&m[159]&m[223]))&~BiasedRNG[61])|((~m[31]&~m[159]&m[223])|(m[31]&~m[159]&m[223])|(m[31]&m[159]&m[223]))):InitCond[77];
    m[110] = run?((((~m[31]&~m[167]&~m[231])|(m[31]&m[167]&~m[231]))&BiasedRNG[62])|(((m[31]&~m[167]&~m[231])|(~m[31]&m[167]&m[231]))&~BiasedRNG[62])|((~m[31]&~m[167]&m[231])|(m[31]&~m[167]&m[231])|(m[31]&m[167]&m[231]))):InitCond[78];
    m[111] = run?((((~m[31]&~m[175]&~m[239])|(m[31]&m[175]&~m[239]))&BiasedRNG[63])|(((m[31]&~m[175]&~m[239])|(~m[31]&m[175]&m[239]))&~BiasedRNG[63])|((~m[31]&~m[175]&m[239])|(m[31]&~m[175]&m[239])|(m[31]&m[175]&m[239]))):InitCond[79];
    m[240] = run?((((m[177]&~m[241]&~m[242]&~m[243]&~m[244])|(~m[177]&~m[241]&~m[242]&m[243]&~m[244])|(m[177]&m[241]&~m[242]&m[243]&~m[244])|(m[177]&~m[241]&m[242]&m[243]&~m[244])|(~m[177]&m[241]&~m[242]&~m[243]&m[244])|(~m[177]&~m[241]&m[242]&~m[243]&m[244])|(m[177]&m[241]&m[242]&~m[243]&m[244])|(~m[177]&m[241]&m[242]&m[243]&m[244]))&UnbiasedRNG[16])|((m[177]&~m[241]&~m[242]&m[243]&~m[244])|(~m[177]&~m[241]&~m[242]&~m[243]&m[244])|(m[177]&~m[241]&~m[242]&~m[243]&m[244])|(m[177]&m[241]&~m[242]&~m[243]&m[244])|(m[177]&~m[241]&m[242]&~m[243]&m[244])|(~m[177]&~m[241]&~m[242]&m[243]&m[244])|(m[177]&~m[241]&~m[242]&m[243]&m[244])|(~m[177]&m[241]&~m[242]&m[243]&m[244])|(m[177]&m[241]&~m[242]&m[243]&m[244])|(~m[177]&~m[241]&m[242]&m[243]&m[244])|(m[177]&~m[241]&m[242]&m[243]&m[244])|(m[177]&m[241]&m[242]&m[243]&m[244]))):InitCond[80];
    m[245] = run?((((m[178]&~m[246]&~m[247]&~m[248]&~m[249])|(~m[178]&~m[246]&~m[247]&m[248]&~m[249])|(m[178]&m[246]&~m[247]&m[248]&~m[249])|(m[178]&~m[246]&m[247]&m[248]&~m[249])|(~m[178]&m[246]&~m[247]&~m[248]&m[249])|(~m[178]&~m[246]&m[247]&~m[248]&m[249])|(m[178]&m[246]&m[247]&~m[248]&m[249])|(~m[178]&m[246]&m[247]&m[248]&m[249]))&UnbiasedRNG[17])|((m[178]&~m[246]&~m[247]&m[248]&~m[249])|(~m[178]&~m[246]&~m[247]&~m[248]&m[249])|(m[178]&~m[246]&~m[247]&~m[248]&m[249])|(m[178]&m[246]&~m[247]&~m[248]&m[249])|(m[178]&~m[246]&m[247]&~m[248]&m[249])|(~m[178]&~m[246]&~m[247]&m[248]&m[249])|(m[178]&~m[246]&~m[247]&m[248]&m[249])|(~m[178]&m[246]&~m[247]&m[248]&m[249])|(m[178]&m[246]&~m[247]&m[248]&m[249])|(~m[178]&~m[246]&m[247]&m[248]&m[249])|(m[178]&~m[246]&m[247]&m[248]&m[249])|(m[178]&m[246]&m[247]&m[248]&m[249]))):InitCond[81];
    m[250] = run?((((m[248]&~m[251]&~m[252]&~m[253]&~m[254])|(~m[248]&~m[251]&~m[252]&m[253]&~m[254])|(m[248]&m[251]&~m[252]&m[253]&~m[254])|(m[248]&~m[251]&m[252]&m[253]&~m[254])|(~m[248]&m[251]&~m[252]&~m[253]&m[254])|(~m[248]&~m[251]&m[252]&~m[253]&m[254])|(m[248]&m[251]&m[252]&~m[253]&m[254])|(~m[248]&m[251]&m[252]&m[253]&m[254]))&UnbiasedRNG[18])|((m[248]&~m[251]&~m[252]&m[253]&~m[254])|(~m[248]&~m[251]&~m[252]&~m[253]&m[254])|(m[248]&~m[251]&~m[252]&~m[253]&m[254])|(m[248]&m[251]&~m[252]&~m[253]&m[254])|(m[248]&~m[251]&m[252]&~m[253]&m[254])|(~m[248]&~m[251]&~m[252]&m[253]&m[254])|(m[248]&~m[251]&~m[252]&m[253]&m[254])|(~m[248]&m[251]&~m[252]&m[253]&m[254])|(m[248]&m[251]&~m[252]&m[253]&m[254])|(~m[248]&~m[251]&m[252]&m[253]&m[254])|(m[248]&~m[251]&m[252]&m[253]&m[254])|(m[248]&m[251]&m[252]&m[253]&m[254]))):InitCond[82];
    m[255] = run?((((m[179]&~m[256]&~m[257]&~m[258]&~m[259])|(~m[179]&~m[256]&~m[257]&m[258]&~m[259])|(m[179]&m[256]&~m[257]&m[258]&~m[259])|(m[179]&~m[256]&m[257]&m[258]&~m[259])|(~m[179]&m[256]&~m[257]&~m[258]&m[259])|(~m[179]&~m[256]&m[257]&~m[258]&m[259])|(m[179]&m[256]&m[257]&~m[258]&m[259])|(~m[179]&m[256]&m[257]&m[258]&m[259]))&UnbiasedRNG[19])|((m[179]&~m[256]&~m[257]&m[258]&~m[259])|(~m[179]&~m[256]&~m[257]&~m[258]&m[259])|(m[179]&~m[256]&~m[257]&~m[258]&m[259])|(m[179]&m[256]&~m[257]&~m[258]&m[259])|(m[179]&~m[256]&m[257]&~m[258]&m[259])|(~m[179]&~m[256]&~m[257]&m[258]&m[259])|(m[179]&~m[256]&~m[257]&m[258]&m[259])|(~m[179]&m[256]&~m[257]&m[258]&m[259])|(m[179]&m[256]&~m[257]&m[258]&m[259])|(~m[179]&~m[256]&m[257]&m[258]&m[259])|(m[179]&~m[256]&m[257]&m[258]&m[259])|(m[179]&m[256]&m[257]&m[258]&m[259]))):InitCond[83];
    m[260] = run?((((m[258]&~m[261]&~m[262]&~m[263]&~m[264])|(~m[258]&~m[261]&~m[262]&m[263]&~m[264])|(m[258]&m[261]&~m[262]&m[263]&~m[264])|(m[258]&~m[261]&m[262]&m[263]&~m[264])|(~m[258]&m[261]&~m[262]&~m[263]&m[264])|(~m[258]&~m[261]&m[262]&~m[263]&m[264])|(m[258]&m[261]&m[262]&~m[263]&m[264])|(~m[258]&m[261]&m[262]&m[263]&m[264]))&UnbiasedRNG[20])|((m[258]&~m[261]&~m[262]&m[263]&~m[264])|(~m[258]&~m[261]&~m[262]&~m[263]&m[264])|(m[258]&~m[261]&~m[262]&~m[263]&m[264])|(m[258]&m[261]&~m[262]&~m[263]&m[264])|(m[258]&~m[261]&m[262]&~m[263]&m[264])|(~m[258]&~m[261]&~m[262]&m[263]&m[264])|(m[258]&~m[261]&~m[262]&m[263]&m[264])|(~m[258]&m[261]&~m[262]&m[263]&m[264])|(m[258]&m[261]&~m[262]&m[263]&m[264])|(~m[258]&~m[261]&m[262]&m[263]&m[264])|(m[258]&~m[261]&m[262]&m[263]&m[264])|(m[258]&m[261]&m[262]&m[263]&m[264]))):InitCond[84];
    m[265] = run?((((m[263]&~m[266]&~m[267]&~m[268]&~m[269])|(~m[263]&~m[266]&~m[267]&m[268]&~m[269])|(m[263]&m[266]&~m[267]&m[268]&~m[269])|(m[263]&~m[266]&m[267]&m[268]&~m[269])|(~m[263]&m[266]&~m[267]&~m[268]&m[269])|(~m[263]&~m[266]&m[267]&~m[268]&m[269])|(m[263]&m[266]&m[267]&~m[268]&m[269])|(~m[263]&m[266]&m[267]&m[268]&m[269]))&UnbiasedRNG[21])|((m[263]&~m[266]&~m[267]&m[268]&~m[269])|(~m[263]&~m[266]&~m[267]&~m[268]&m[269])|(m[263]&~m[266]&~m[267]&~m[268]&m[269])|(m[263]&m[266]&~m[267]&~m[268]&m[269])|(m[263]&~m[266]&m[267]&~m[268]&m[269])|(~m[263]&~m[266]&~m[267]&m[268]&m[269])|(m[263]&~m[266]&~m[267]&m[268]&m[269])|(~m[263]&m[266]&~m[267]&m[268]&m[269])|(m[263]&m[266]&~m[267]&m[268]&m[269])|(~m[263]&~m[266]&m[267]&m[268]&m[269])|(m[263]&~m[266]&m[267]&m[268]&m[269])|(m[263]&m[266]&m[267]&m[268]&m[269]))):InitCond[85];
    m[270] = run?((((m[180]&~m[271]&~m[272]&~m[273]&~m[274])|(~m[180]&~m[271]&~m[272]&m[273]&~m[274])|(m[180]&m[271]&~m[272]&m[273]&~m[274])|(m[180]&~m[271]&m[272]&m[273]&~m[274])|(~m[180]&m[271]&~m[272]&~m[273]&m[274])|(~m[180]&~m[271]&m[272]&~m[273]&m[274])|(m[180]&m[271]&m[272]&~m[273]&m[274])|(~m[180]&m[271]&m[272]&m[273]&m[274]))&UnbiasedRNG[22])|((m[180]&~m[271]&~m[272]&m[273]&~m[274])|(~m[180]&~m[271]&~m[272]&~m[273]&m[274])|(m[180]&~m[271]&~m[272]&~m[273]&m[274])|(m[180]&m[271]&~m[272]&~m[273]&m[274])|(m[180]&~m[271]&m[272]&~m[273]&m[274])|(~m[180]&~m[271]&~m[272]&m[273]&m[274])|(m[180]&~m[271]&~m[272]&m[273]&m[274])|(~m[180]&m[271]&~m[272]&m[273]&m[274])|(m[180]&m[271]&~m[272]&m[273]&m[274])|(~m[180]&~m[271]&m[272]&m[273]&m[274])|(m[180]&~m[271]&m[272]&m[273]&m[274])|(m[180]&m[271]&m[272]&m[273]&m[274]))):InitCond[86];
    m[275] = run?((((m[273]&~m[276]&~m[277]&~m[278]&~m[279])|(~m[273]&~m[276]&~m[277]&m[278]&~m[279])|(m[273]&m[276]&~m[277]&m[278]&~m[279])|(m[273]&~m[276]&m[277]&m[278]&~m[279])|(~m[273]&m[276]&~m[277]&~m[278]&m[279])|(~m[273]&~m[276]&m[277]&~m[278]&m[279])|(m[273]&m[276]&m[277]&~m[278]&m[279])|(~m[273]&m[276]&m[277]&m[278]&m[279]))&UnbiasedRNG[23])|((m[273]&~m[276]&~m[277]&m[278]&~m[279])|(~m[273]&~m[276]&~m[277]&~m[278]&m[279])|(m[273]&~m[276]&~m[277]&~m[278]&m[279])|(m[273]&m[276]&~m[277]&~m[278]&m[279])|(m[273]&~m[276]&m[277]&~m[278]&m[279])|(~m[273]&~m[276]&~m[277]&m[278]&m[279])|(m[273]&~m[276]&~m[277]&m[278]&m[279])|(~m[273]&m[276]&~m[277]&m[278]&m[279])|(m[273]&m[276]&~m[277]&m[278]&m[279])|(~m[273]&~m[276]&m[277]&m[278]&m[279])|(m[273]&~m[276]&m[277]&m[278]&m[279])|(m[273]&m[276]&m[277]&m[278]&m[279]))):InitCond[87];
    m[280] = run?((((m[278]&~m[281]&~m[282]&~m[283]&~m[284])|(~m[278]&~m[281]&~m[282]&m[283]&~m[284])|(m[278]&m[281]&~m[282]&m[283]&~m[284])|(m[278]&~m[281]&m[282]&m[283]&~m[284])|(~m[278]&m[281]&~m[282]&~m[283]&m[284])|(~m[278]&~m[281]&m[282]&~m[283]&m[284])|(m[278]&m[281]&m[282]&~m[283]&m[284])|(~m[278]&m[281]&m[282]&m[283]&m[284]))&UnbiasedRNG[24])|((m[278]&~m[281]&~m[282]&m[283]&~m[284])|(~m[278]&~m[281]&~m[282]&~m[283]&m[284])|(m[278]&~m[281]&~m[282]&~m[283]&m[284])|(m[278]&m[281]&~m[282]&~m[283]&m[284])|(m[278]&~m[281]&m[282]&~m[283]&m[284])|(~m[278]&~m[281]&~m[282]&m[283]&m[284])|(m[278]&~m[281]&~m[282]&m[283]&m[284])|(~m[278]&m[281]&~m[282]&m[283]&m[284])|(m[278]&m[281]&~m[282]&m[283]&m[284])|(~m[278]&~m[281]&m[282]&m[283]&m[284])|(m[278]&~m[281]&m[282]&m[283]&m[284])|(m[278]&m[281]&m[282]&m[283]&m[284]))):InitCond[88];
    m[285] = run?((((m[283]&~m[286]&~m[287]&~m[288]&~m[289])|(~m[283]&~m[286]&~m[287]&m[288]&~m[289])|(m[283]&m[286]&~m[287]&m[288]&~m[289])|(m[283]&~m[286]&m[287]&m[288]&~m[289])|(~m[283]&m[286]&~m[287]&~m[288]&m[289])|(~m[283]&~m[286]&m[287]&~m[288]&m[289])|(m[283]&m[286]&m[287]&~m[288]&m[289])|(~m[283]&m[286]&m[287]&m[288]&m[289]))&UnbiasedRNG[25])|((m[283]&~m[286]&~m[287]&m[288]&~m[289])|(~m[283]&~m[286]&~m[287]&~m[288]&m[289])|(m[283]&~m[286]&~m[287]&~m[288]&m[289])|(m[283]&m[286]&~m[287]&~m[288]&m[289])|(m[283]&~m[286]&m[287]&~m[288]&m[289])|(~m[283]&~m[286]&~m[287]&m[288]&m[289])|(m[283]&~m[286]&~m[287]&m[288]&m[289])|(~m[283]&m[286]&~m[287]&m[288]&m[289])|(m[283]&m[286]&~m[287]&m[288]&m[289])|(~m[283]&~m[286]&m[287]&m[288]&m[289])|(m[283]&~m[286]&m[287]&m[288]&m[289])|(m[283]&m[286]&m[287]&m[288]&m[289]))):InitCond[89];
    m[290] = run?((((m[181]&~m[291]&~m[292]&~m[293]&~m[294])|(~m[181]&~m[291]&~m[292]&m[293]&~m[294])|(m[181]&m[291]&~m[292]&m[293]&~m[294])|(m[181]&~m[291]&m[292]&m[293]&~m[294])|(~m[181]&m[291]&~m[292]&~m[293]&m[294])|(~m[181]&~m[291]&m[292]&~m[293]&m[294])|(m[181]&m[291]&m[292]&~m[293]&m[294])|(~m[181]&m[291]&m[292]&m[293]&m[294]))&UnbiasedRNG[26])|((m[181]&~m[291]&~m[292]&m[293]&~m[294])|(~m[181]&~m[291]&~m[292]&~m[293]&m[294])|(m[181]&~m[291]&~m[292]&~m[293]&m[294])|(m[181]&m[291]&~m[292]&~m[293]&m[294])|(m[181]&~m[291]&m[292]&~m[293]&m[294])|(~m[181]&~m[291]&~m[292]&m[293]&m[294])|(m[181]&~m[291]&~m[292]&m[293]&m[294])|(~m[181]&m[291]&~m[292]&m[293]&m[294])|(m[181]&m[291]&~m[292]&m[293]&m[294])|(~m[181]&~m[291]&m[292]&m[293]&m[294])|(m[181]&~m[291]&m[292]&m[293]&m[294])|(m[181]&m[291]&m[292]&m[293]&m[294]))):InitCond[90];
    m[295] = run?((((m[293]&~m[296]&~m[297]&~m[298]&~m[299])|(~m[293]&~m[296]&~m[297]&m[298]&~m[299])|(m[293]&m[296]&~m[297]&m[298]&~m[299])|(m[293]&~m[296]&m[297]&m[298]&~m[299])|(~m[293]&m[296]&~m[297]&~m[298]&m[299])|(~m[293]&~m[296]&m[297]&~m[298]&m[299])|(m[293]&m[296]&m[297]&~m[298]&m[299])|(~m[293]&m[296]&m[297]&m[298]&m[299]))&UnbiasedRNG[27])|((m[293]&~m[296]&~m[297]&m[298]&~m[299])|(~m[293]&~m[296]&~m[297]&~m[298]&m[299])|(m[293]&~m[296]&~m[297]&~m[298]&m[299])|(m[293]&m[296]&~m[297]&~m[298]&m[299])|(m[293]&~m[296]&m[297]&~m[298]&m[299])|(~m[293]&~m[296]&~m[297]&m[298]&m[299])|(m[293]&~m[296]&~m[297]&m[298]&m[299])|(~m[293]&m[296]&~m[297]&m[298]&m[299])|(m[293]&m[296]&~m[297]&m[298]&m[299])|(~m[293]&~m[296]&m[297]&m[298]&m[299])|(m[293]&~m[296]&m[297]&m[298]&m[299])|(m[293]&m[296]&m[297]&m[298]&m[299]))):InitCond[91];
    m[300] = run?((((m[298]&~m[301]&~m[302]&~m[303]&~m[304])|(~m[298]&~m[301]&~m[302]&m[303]&~m[304])|(m[298]&m[301]&~m[302]&m[303]&~m[304])|(m[298]&~m[301]&m[302]&m[303]&~m[304])|(~m[298]&m[301]&~m[302]&~m[303]&m[304])|(~m[298]&~m[301]&m[302]&~m[303]&m[304])|(m[298]&m[301]&m[302]&~m[303]&m[304])|(~m[298]&m[301]&m[302]&m[303]&m[304]))&UnbiasedRNG[28])|((m[298]&~m[301]&~m[302]&m[303]&~m[304])|(~m[298]&~m[301]&~m[302]&~m[303]&m[304])|(m[298]&~m[301]&~m[302]&~m[303]&m[304])|(m[298]&m[301]&~m[302]&~m[303]&m[304])|(m[298]&~m[301]&m[302]&~m[303]&m[304])|(~m[298]&~m[301]&~m[302]&m[303]&m[304])|(m[298]&~m[301]&~m[302]&m[303]&m[304])|(~m[298]&m[301]&~m[302]&m[303]&m[304])|(m[298]&m[301]&~m[302]&m[303]&m[304])|(~m[298]&~m[301]&m[302]&m[303]&m[304])|(m[298]&~m[301]&m[302]&m[303]&m[304])|(m[298]&m[301]&m[302]&m[303]&m[304]))):InitCond[92];
    m[305] = run?((((m[303]&~m[306]&~m[307]&~m[308]&~m[309])|(~m[303]&~m[306]&~m[307]&m[308]&~m[309])|(m[303]&m[306]&~m[307]&m[308]&~m[309])|(m[303]&~m[306]&m[307]&m[308]&~m[309])|(~m[303]&m[306]&~m[307]&~m[308]&m[309])|(~m[303]&~m[306]&m[307]&~m[308]&m[309])|(m[303]&m[306]&m[307]&~m[308]&m[309])|(~m[303]&m[306]&m[307]&m[308]&m[309]))&UnbiasedRNG[29])|((m[303]&~m[306]&~m[307]&m[308]&~m[309])|(~m[303]&~m[306]&~m[307]&~m[308]&m[309])|(m[303]&~m[306]&~m[307]&~m[308]&m[309])|(m[303]&m[306]&~m[307]&~m[308]&m[309])|(m[303]&~m[306]&m[307]&~m[308]&m[309])|(~m[303]&~m[306]&~m[307]&m[308]&m[309])|(m[303]&~m[306]&~m[307]&m[308]&m[309])|(~m[303]&m[306]&~m[307]&m[308]&m[309])|(m[303]&m[306]&~m[307]&m[308]&m[309])|(~m[303]&~m[306]&m[307]&m[308]&m[309])|(m[303]&~m[306]&m[307]&m[308]&m[309])|(m[303]&m[306]&m[307]&m[308]&m[309]))):InitCond[93];
    m[310] = run?((((m[308]&~m[311]&~m[312]&~m[313]&~m[314])|(~m[308]&~m[311]&~m[312]&m[313]&~m[314])|(m[308]&m[311]&~m[312]&m[313]&~m[314])|(m[308]&~m[311]&m[312]&m[313]&~m[314])|(~m[308]&m[311]&~m[312]&~m[313]&m[314])|(~m[308]&~m[311]&m[312]&~m[313]&m[314])|(m[308]&m[311]&m[312]&~m[313]&m[314])|(~m[308]&m[311]&m[312]&m[313]&m[314]))&UnbiasedRNG[30])|((m[308]&~m[311]&~m[312]&m[313]&~m[314])|(~m[308]&~m[311]&~m[312]&~m[313]&m[314])|(m[308]&~m[311]&~m[312]&~m[313]&m[314])|(m[308]&m[311]&~m[312]&~m[313]&m[314])|(m[308]&~m[311]&m[312]&~m[313]&m[314])|(~m[308]&~m[311]&~m[312]&m[313]&m[314])|(m[308]&~m[311]&~m[312]&m[313]&m[314])|(~m[308]&m[311]&~m[312]&m[313]&m[314])|(m[308]&m[311]&~m[312]&m[313]&m[314])|(~m[308]&~m[311]&m[312]&m[313]&m[314])|(m[308]&~m[311]&m[312]&m[313]&m[314])|(m[308]&m[311]&m[312]&m[313]&m[314]))):InitCond[94];
    m[315] = run?((((m[182]&~m[316]&~m[317]&~m[318]&~m[319])|(~m[182]&~m[316]&~m[317]&m[318]&~m[319])|(m[182]&m[316]&~m[317]&m[318]&~m[319])|(m[182]&~m[316]&m[317]&m[318]&~m[319])|(~m[182]&m[316]&~m[317]&~m[318]&m[319])|(~m[182]&~m[316]&m[317]&~m[318]&m[319])|(m[182]&m[316]&m[317]&~m[318]&m[319])|(~m[182]&m[316]&m[317]&m[318]&m[319]))&UnbiasedRNG[31])|((m[182]&~m[316]&~m[317]&m[318]&~m[319])|(~m[182]&~m[316]&~m[317]&~m[318]&m[319])|(m[182]&~m[316]&~m[317]&~m[318]&m[319])|(m[182]&m[316]&~m[317]&~m[318]&m[319])|(m[182]&~m[316]&m[317]&~m[318]&m[319])|(~m[182]&~m[316]&~m[317]&m[318]&m[319])|(m[182]&~m[316]&~m[317]&m[318]&m[319])|(~m[182]&m[316]&~m[317]&m[318]&m[319])|(m[182]&m[316]&~m[317]&m[318]&m[319])|(~m[182]&~m[316]&m[317]&m[318]&m[319])|(m[182]&~m[316]&m[317]&m[318]&m[319])|(m[182]&m[316]&m[317]&m[318]&m[319]))):InitCond[95];
    m[320] = run?((((m[318]&~m[321]&~m[322]&~m[323]&~m[324])|(~m[318]&~m[321]&~m[322]&m[323]&~m[324])|(m[318]&m[321]&~m[322]&m[323]&~m[324])|(m[318]&~m[321]&m[322]&m[323]&~m[324])|(~m[318]&m[321]&~m[322]&~m[323]&m[324])|(~m[318]&~m[321]&m[322]&~m[323]&m[324])|(m[318]&m[321]&m[322]&~m[323]&m[324])|(~m[318]&m[321]&m[322]&m[323]&m[324]))&UnbiasedRNG[32])|((m[318]&~m[321]&~m[322]&m[323]&~m[324])|(~m[318]&~m[321]&~m[322]&~m[323]&m[324])|(m[318]&~m[321]&~m[322]&~m[323]&m[324])|(m[318]&m[321]&~m[322]&~m[323]&m[324])|(m[318]&~m[321]&m[322]&~m[323]&m[324])|(~m[318]&~m[321]&~m[322]&m[323]&m[324])|(m[318]&~m[321]&~m[322]&m[323]&m[324])|(~m[318]&m[321]&~m[322]&m[323]&m[324])|(m[318]&m[321]&~m[322]&m[323]&m[324])|(~m[318]&~m[321]&m[322]&m[323]&m[324])|(m[318]&~m[321]&m[322]&m[323]&m[324])|(m[318]&m[321]&m[322]&m[323]&m[324]))):InitCond[96];
    m[325] = run?((((m[323]&~m[326]&~m[327]&~m[328]&~m[329])|(~m[323]&~m[326]&~m[327]&m[328]&~m[329])|(m[323]&m[326]&~m[327]&m[328]&~m[329])|(m[323]&~m[326]&m[327]&m[328]&~m[329])|(~m[323]&m[326]&~m[327]&~m[328]&m[329])|(~m[323]&~m[326]&m[327]&~m[328]&m[329])|(m[323]&m[326]&m[327]&~m[328]&m[329])|(~m[323]&m[326]&m[327]&m[328]&m[329]))&UnbiasedRNG[33])|((m[323]&~m[326]&~m[327]&m[328]&~m[329])|(~m[323]&~m[326]&~m[327]&~m[328]&m[329])|(m[323]&~m[326]&~m[327]&~m[328]&m[329])|(m[323]&m[326]&~m[327]&~m[328]&m[329])|(m[323]&~m[326]&m[327]&~m[328]&m[329])|(~m[323]&~m[326]&~m[327]&m[328]&m[329])|(m[323]&~m[326]&~m[327]&m[328]&m[329])|(~m[323]&m[326]&~m[327]&m[328]&m[329])|(m[323]&m[326]&~m[327]&m[328]&m[329])|(~m[323]&~m[326]&m[327]&m[328]&m[329])|(m[323]&~m[326]&m[327]&m[328]&m[329])|(m[323]&m[326]&m[327]&m[328]&m[329]))):InitCond[97];
    m[330] = run?((((m[328]&~m[331]&~m[332]&~m[333]&~m[334])|(~m[328]&~m[331]&~m[332]&m[333]&~m[334])|(m[328]&m[331]&~m[332]&m[333]&~m[334])|(m[328]&~m[331]&m[332]&m[333]&~m[334])|(~m[328]&m[331]&~m[332]&~m[333]&m[334])|(~m[328]&~m[331]&m[332]&~m[333]&m[334])|(m[328]&m[331]&m[332]&~m[333]&m[334])|(~m[328]&m[331]&m[332]&m[333]&m[334]))&UnbiasedRNG[34])|((m[328]&~m[331]&~m[332]&m[333]&~m[334])|(~m[328]&~m[331]&~m[332]&~m[333]&m[334])|(m[328]&~m[331]&~m[332]&~m[333]&m[334])|(m[328]&m[331]&~m[332]&~m[333]&m[334])|(m[328]&~m[331]&m[332]&~m[333]&m[334])|(~m[328]&~m[331]&~m[332]&m[333]&m[334])|(m[328]&~m[331]&~m[332]&m[333]&m[334])|(~m[328]&m[331]&~m[332]&m[333]&m[334])|(m[328]&m[331]&~m[332]&m[333]&m[334])|(~m[328]&~m[331]&m[332]&m[333]&m[334])|(m[328]&~m[331]&m[332]&m[333]&m[334])|(m[328]&m[331]&m[332]&m[333]&m[334]))):InitCond[98];
    m[335] = run?((((m[333]&~m[336]&~m[337]&~m[338]&~m[339])|(~m[333]&~m[336]&~m[337]&m[338]&~m[339])|(m[333]&m[336]&~m[337]&m[338]&~m[339])|(m[333]&~m[336]&m[337]&m[338]&~m[339])|(~m[333]&m[336]&~m[337]&~m[338]&m[339])|(~m[333]&~m[336]&m[337]&~m[338]&m[339])|(m[333]&m[336]&m[337]&~m[338]&m[339])|(~m[333]&m[336]&m[337]&m[338]&m[339]))&UnbiasedRNG[35])|((m[333]&~m[336]&~m[337]&m[338]&~m[339])|(~m[333]&~m[336]&~m[337]&~m[338]&m[339])|(m[333]&~m[336]&~m[337]&~m[338]&m[339])|(m[333]&m[336]&~m[337]&~m[338]&m[339])|(m[333]&~m[336]&m[337]&~m[338]&m[339])|(~m[333]&~m[336]&~m[337]&m[338]&m[339])|(m[333]&~m[336]&~m[337]&m[338]&m[339])|(~m[333]&m[336]&~m[337]&m[338]&m[339])|(m[333]&m[336]&~m[337]&m[338]&m[339])|(~m[333]&~m[336]&m[337]&m[338]&m[339])|(m[333]&~m[336]&m[337]&m[338]&m[339])|(m[333]&m[336]&m[337]&m[338]&m[339]))):InitCond[99];
    m[340] = run?((((m[338]&~m[341]&~m[342]&~m[343]&~m[344])|(~m[338]&~m[341]&~m[342]&m[343]&~m[344])|(m[338]&m[341]&~m[342]&m[343]&~m[344])|(m[338]&~m[341]&m[342]&m[343]&~m[344])|(~m[338]&m[341]&~m[342]&~m[343]&m[344])|(~m[338]&~m[341]&m[342]&~m[343]&m[344])|(m[338]&m[341]&m[342]&~m[343]&m[344])|(~m[338]&m[341]&m[342]&m[343]&m[344]))&UnbiasedRNG[36])|((m[338]&~m[341]&~m[342]&m[343]&~m[344])|(~m[338]&~m[341]&~m[342]&~m[343]&m[344])|(m[338]&~m[341]&~m[342]&~m[343]&m[344])|(m[338]&m[341]&~m[342]&~m[343]&m[344])|(m[338]&~m[341]&m[342]&~m[343]&m[344])|(~m[338]&~m[341]&~m[342]&m[343]&m[344])|(m[338]&~m[341]&~m[342]&m[343]&m[344])|(~m[338]&m[341]&~m[342]&m[343]&m[344])|(m[338]&m[341]&~m[342]&m[343]&m[344])|(~m[338]&~m[341]&m[342]&m[343]&m[344])|(m[338]&~m[341]&m[342]&m[343]&m[344])|(m[338]&m[341]&m[342]&m[343]&m[344]))):InitCond[100];
    m[345] = run?((((m[183]&~m[346]&~m[347]&~m[348]&~m[349])|(~m[183]&~m[346]&~m[347]&m[348]&~m[349])|(m[183]&m[346]&~m[347]&m[348]&~m[349])|(m[183]&~m[346]&m[347]&m[348]&~m[349])|(~m[183]&m[346]&~m[347]&~m[348]&m[349])|(~m[183]&~m[346]&m[347]&~m[348]&m[349])|(m[183]&m[346]&m[347]&~m[348]&m[349])|(~m[183]&m[346]&m[347]&m[348]&m[349]))&UnbiasedRNG[37])|((m[183]&~m[346]&~m[347]&m[348]&~m[349])|(~m[183]&~m[346]&~m[347]&~m[348]&m[349])|(m[183]&~m[346]&~m[347]&~m[348]&m[349])|(m[183]&m[346]&~m[347]&~m[348]&m[349])|(m[183]&~m[346]&m[347]&~m[348]&m[349])|(~m[183]&~m[346]&~m[347]&m[348]&m[349])|(m[183]&~m[346]&~m[347]&m[348]&m[349])|(~m[183]&m[346]&~m[347]&m[348]&m[349])|(m[183]&m[346]&~m[347]&m[348]&m[349])|(~m[183]&~m[346]&m[347]&m[348]&m[349])|(m[183]&~m[346]&m[347]&m[348]&m[349])|(m[183]&m[346]&m[347]&m[348]&m[349]))):InitCond[101];
    m[350] = run?((((m[348]&~m[351]&~m[352]&~m[353]&~m[354])|(~m[348]&~m[351]&~m[352]&m[353]&~m[354])|(m[348]&m[351]&~m[352]&m[353]&~m[354])|(m[348]&~m[351]&m[352]&m[353]&~m[354])|(~m[348]&m[351]&~m[352]&~m[353]&m[354])|(~m[348]&~m[351]&m[352]&~m[353]&m[354])|(m[348]&m[351]&m[352]&~m[353]&m[354])|(~m[348]&m[351]&m[352]&m[353]&m[354]))&UnbiasedRNG[38])|((m[348]&~m[351]&~m[352]&m[353]&~m[354])|(~m[348]&~m[351]&~m[352]&~m[353]&m[354])|(m[348]&~m[351]&~m[352]&~m[353]&m[354])|(m[348]&m[351]&~m[352]&~m[353]&m[354])|(m[348]&~m[351]&m[352]&~m[353]&m[354])|(~m[348]&~m[351]&~m[352]&m[353]&m[354])|(m[348]&~m[351]&~m[352]&m[353]&m[354])|(~m[348]&m[351]&~m[352]&m[353]&m[354])|(m[348]&m[351]&~m[352]&m[353]&m[354])|(~m[348]&~m[351]&m[352]&m[353]&m[354])|(m[348]&~m[351]&m[352]&m[353]&m[354])|(m[348]&m[351]&m[352]&m[353]&m[354]))):InitCond[102];
    m[355] = run?((((m[353]&~m[356]&~m[357]&~m[358]&~m[359])|(~m[353]&~m[356]&~m[357]&m[358]&~m[359])|(m[353]&m[356]&~m[357]&m[358]&~m[359])|(m[353]&~m[356]&m[357]&m[358]&~m[359])|(~m[353]&m[356]&~m[357]&~m[358]&m[359])|(~m[353]&~m[356]&m[357]&~m[358]&m[359])|(m[353]&m[356]&m[357]&~m[358]&m[359])|(~m[353]&m[356]&m[357]&m[358]&m[359]))&UnbiasedRNG[39])|((m[353]&~m[356]&~m[357]&m[358]&~m[359])|(~m[353]&~m[356]&~m[357]&~m[358]&m[359])|(m[353]&~m[356]&~m[357]&~m[358]&m[359])|(m[353]&m[356]&~m[357]&~m[358]&m[359])|(m[353]&~m[356]&m[357]&~m[358]&m[359])|(~m[353]&~m[356]&~m[357]&m[358]&m[359])|(m[353]&~m[356]&~m[357]&m[358]&m[359])|(~m[353]&m[356]&~m[357]&m[358]&m[359])|(m[353]&m[356]&~m[357]&m[358]&m[359])|(~m[353]&~m[356]&m[357]&m[358]&m[359])|(m[353]&~m[356]&m[357]&m[358]&m[359])|(m[353]&m[356]&m[357]&m[358]&m[359]))):InitCond[103];
    m[360] = run?((((m[358]&~m[361]&~m[362]&~m[363]&~m[364])|(~m[358]&~m[361]&~m[362]&m[363]&~m[364])|(m[358]&m[361]&~m[362]&m[363]&~m[364])|(m[358]&~m[361]&m[362]&m[363]&~m[364])|(~m[358]&m[361]&~m[362]&~m[363]&m[364])|(~m[358]&~m[361]&m[362]&~m[363]&m[364])|(m[358]&m[361]&m[362]&~m[363]&m[364])|(~m[358]&m[361]&m[362]&m[363]&m[364]))&UnbiasedRNG[40])|((m[358]&~m[361]&~m[362]&m[363]&~m[364])|(~m[358]&~m[361]&~m[362]&~m[363]&m[364])|(m[358]&~m[361]&~m[362]&~m[363]&m[364])|(m[358]&m[361]&~m[362]&~m[363]&m[364])|(m[358]&~m[361]&m[362]&~m[363]&m[364])|(~m[358]&~m[361]&~m[362]&m[363]&m[364])|(m[358]&~m[361]&~m[362]&m[363]&m[364])|(~m[358]&m[361]&~m[362]&m[363]&m[364])|(m[358]&m[361]&~m[362]&m[363]&m[364])|(~m[358]&~m[361]&m[362]&m[363]&m[364])|(m[358]&~m[361]&m[362]&m[363]&m[364])|(m[358]&m[361]&m[362]&m[363]&m[364]))):InitCond[104];
    m[365] = run?((((m[363]&~m[366]&~m[367]&~m[368]&~m[369])|(~m[363]&~m[366]&~m[367]&m[368]&~m[369])|(m[363]&m[366]&~m[367]&m[368]&~m[369])|(m[363]&~m[366]&m[367]&m[368]&~m[369])|(~m[363]&m[366]&~m[367]&~m[368]&m[369])|(~m[363]&~m[366]&m[367]&~m[368]&m[369])|(m[363]&m[366]&m[367]&~m[368]&m[369])|(~m[363]&m[366]&m[367]&m[368]&m[369]))&UnbiasedRNG[41])|((m[363]&~m[366]&~m[367]&m[368]&~m[369])|(~m[363]&~m[366]&~m[367]&~m[368]&m[369])|(m[363]&~m[366]&~m[367]&~m[368]&m[369])|(m[363]&m[366]&~m[367]&~m[368]&m[369])|(m[363]&~m[366]&m[367]&~m[368]&m[369])|(~m[363]&~m[366]&~m[367]&m[368]&m[369])|(m[363]&~m[366]&~m[367]&m[368]&m[369])|(~m[363]&m[366]&~m[367]&m[368]&m[369])|(m[363]&m[366]&~m[367]&m[368]&m[369])|(~m[363]&~m[366]&m[367]&m[368]&m[369])|(m[363]&~m[366]&m[367]&m[368]&m[369])|(m[363]&m[366]&m[367]&m[368]&m[369]))):InitCond[105];
    m[370] = run?((((m[368]&~m[371]&~m[372]&~m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&m[373]&~m[374])|(m[368]&m[371]&~m[372]&m[373]&~m[374])|(m[368]&~m[371]&m[372]&m[373]&~m[374])|(~m[368]&m[371]&~m[372]&~m[373]&m[374])|(~m[368]&~m[371]&m[372]&~m[373]&m[374])|(m[368]&m[371]&m[372]&~m[373]&m[374])|(~m[368]&m[371]&m[372]&m[373]&m[374]))&UnbiasedRNG[42])|((m[368]&~m[371]&~m[372]&m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&m[372]&~m[373]&m[374])|(~m[368]&~m[371]&~m[372]&m[373]&m[374])|(m[368]&~m[371]&~m[372]&m[373]&m[374])|(~m[368]&m[371]&~m[372]&m[373]&m[374])|(m[368]&m[371]&~m[372]&m[373]&m[374])|(~m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&m[371]&m[372]&m[373]&m[374]))):InitCond[106];
    m[375] = run?((((m[373]&~m[376]&~m[377]&~m[378]&~m[379])|(~m[373]&~m[376]&~m[377]&m[378]&~m[379])|(m[373]&m[376]&~m[377]&m[378]&~m[379])|(m[373]&~m[376]&m[377]&m[378]&~m[379])|(~m[373]&m[376]&~m[377]&~m[378]&m[379])|(~m[373]&~m[376]&m[377]&~m[378]&m[379])|(m[373]&m[376]&m[377]&~m[378]&m[379])|(~m[373]&m[376]&m[377]&m[378]&m[379]))&UnbiasedRNG[43])|((m[373]&~m[376]&~m[377]&m[378]&~m[379])|(~m[373]&~m[376]&~m[377]&~m[378]&m[379])|(m[373]&~m[376]&~m[377]&~m[378]&m[379])|(m[373]&m[376]&~m[377]&~m[378]&m[379])|(m[373]&~m[376]&m[377]&~m[378]&m[379])|(~m[373]&~m[376]&~m[377]&m[378]&m[379])|(m[373]&~m[376]&~m[377]&m[378]&m[379])|(~m[373]&m[376]&~m[377]&m[378]&m[379])|(m[373]&m[376]&~m[377]&m[378]&m[379])|(~m[373]&~m[376]&m[377]&m[378]&m[379])|(m[373]&~m[376]&m[377]&m[378]&m[379])|(m[373]&m[376]&m[377]&m[378]&m[379]))):InitCond[107];
    m[385] = run?((((m[383]&~m[386]&~m[387]&~m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&m[388]&~m[389])|(m[383]&m[386]&~m[387]&m[388]&~m[389])|(m[383]&~m[386]&m[387]&m[388]&~m[389])|(~m[383]&m[386]&~m[387]&~m[388]&m[389])|(~m[383]&~m[386]&m[387]&~m[388]&m[389])|(m[383]&m[386]&m[387]&~m[388]&m[389])|(~m[383]&m[386]&m[387]&m[388]&m[389]))&UnbiasedRNG[44])|((m[383]&~m[386]&~m[387]&m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&m[387]&~m[388]&m[389])|(~m[383]&~m[386]&~m[387]&m[388]&m[389])|(m[383]&~m[386]&~m[387]&m[388]&m[389])|(~m[383]&m[386]&~m[387]&m[388]&m[389])|(m[383]&m[386]&~m[387]&m[388]&m[389])|(~m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&m[386]&m[387]&m[388]&m[389]))):InitCond[108];
    m[390] = run?((((m[388]&~m[391]&~m[392]&~m[393]&~m[394])|(~m[388]&~m[391]&~m[392]&m[393]&~m[394])|(m[388]&m[391]&~m[392]&m[393]&~m[394])|(m[388]&~m[391]&m[392]&m[393]&~m[394])|(~m[388]&m[391]&~m[392]&~m[393]&m[394])|(~m[388]&~m[391]&m[392]&~m[393]&m[394])|(m[388]&m[391]&m[392]&~m[393]&m[394])|(~m[388]&m[391]&m[392]&m[393]&m[394]))&UnbiasedRNG[45])|((m[388]&~m[391]&~m[392]&m[393]&~m[394])|(~m[388]&~m[391]&~m[392]&~m[393]&m[394])|(m[388]&~m[391]&~m[392]&~m[393]&m[394])|(m[388]&m[391]&~m[392]&~m[393]&m[394])|(m[388]&~m[391]&m[392]&~m[393]&m[394])|(~m[388]&~m[391]&~m[392]&m[393]&m[394])|(m[388]&~m[391]&~m[392]&m[393]&m[394])|(~m[388]&m[391]&~m[392]&m[393]&m[394])|(m[388]&m[391]&~m[392]&m[393]&m[394])|(~m[388]&~m[391]&m[392]&m[393]&m[394])|(m[388]&~m[391]&m[392]&m[393]&m[394])|(m[388]&m[391]&m[392]&m[393]&m[394]))):InitCond[109];
    m[395] = run?((((m[393]&~m[396]&~m[397]&~m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&m[398]&~m[399])|(m[393]&m[396]&~m[397]&m[398]&~m[399])|(m[393]&~m[396]&m[397]&m[398]&~m[399])|(~m[393]&m[396]&~m[397]&~m[398]&m[399])|(~m[393]&~m[396]&m[397]&~m[398]&m[399])|(m[393]&m[396]&m[397]&~m[398]&m[399])|(~m[393]&m[396]&m[397]&m[398]&m[399]))&UnbiasedRNG[46])|((m[393]&~m[396]&~m[397]&m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&m[397]&~m[398]&m[399])|(~m[393]&~m[396]&~m[397]&m[398]&m[399])|(m[393]&~m[396]&~m[397]&m[398]&m[399])|(~m[393]&m[396]&~m[397]&m[398]&m[399])|(m[393]&m[396]&~m[397]&m[398]&m[399])|(~m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&m[396]&m[397]&m[398]&m[399]))):InitCond[110];
    m[400] = run?((((m[398]&~m[401]&~m[402]&~m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&m[403]&~m[404])|(m[398]&m[401]&~m[402]&m[403]&~m[404])|(m[398]&~m[401]&m[402]&m[403]&~m[404])|(~m[398]&m[401]&~m[402]&~m[403]&m[404])|(~m[398]&~m[401]&m[402]&~m[403]&m[404])|(m[398]&m[401]&m[402]&~m[403]&m[404])|(~m[398]&m[401]&m[402]&m[403]&m[404]))&UnbiasedRNG[47])|((m[398]&~m[401]&~m[402]&m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&m[402]&~m[403]&m[404])|(~m[398]&~m[401]&~m[402]&m[403]&m[404])|(m[398]&~m[401]&~m[402]&m[403]&m[404])|(~m[398]&m[401]&~m[402]&m[403]&m[404])|(m[398]&m[401]&~m[402]&m[403]&m[404])|(~m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&m[401]&m[402]&m[403]&m[404]))):InitCond[111];
    m[405] = run?((((m[403]&~m[406]&~m[407]&~m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&m[408]&~m[409])|(m[403]&m[406]&~m[407]&m[408]&~m[409])|(m[403]&~m[406]&m[407]&m[408]&~m[409])|(~m[403]&m[406]&~m[407]&~m[408]&m[409])|(~m[403]&~m[406]&m[407]&~m[408]&m[409])|(m[403]&m[406]&m[407]&~m[408]&m[409])|(~m[403]&m[406]&m[407]&m[408]&m[409]))&UnbiasedRNG[48])|((m[403]&~m[406]&~m[407]&m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&m[407]&~m[408]&m[409])|(~m[403]&~m[406]&~m[407]&m[408]&m[409])|(m[403]&~m[406]&~m[407]&m[408]&m[409])|(~m[403]&m[406]&~m[407]&m[408]&m[409])|(m[403]&m[406]&~m[407]&m[408]&m[409])|(~m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&m[406]&m[407]&m[408]&m[409]))):InitCond[112];
    m[410] = run?((((m[408]&~m[411]&~m[412]&~m[413]&~m[414])|(~m[408]&~m[411]&~m[412]&m[413]&~m[414])|(m[408]&m[411]&~m[412]&m[413]&~m[414])|(m[408]&~m[411]&m[412]&m[413]&~m[414])|(~m[408]&m[411]&~m[412]&~m[413]&m[414])|(~m[408]&~m[411]&m[412]&~m[413]&m[414])|(m[408]&m[411]&m[412]&~m[413]&m[414])|(~m[408]&m[411]&m[412]&m[413]&m[414]))&UnbiasedRNG[49])|((m[408]&~m[411]&~m[412]&m[413]&~m[414])|(~m[408]&~m[411]&~m[412]&~m[413]&m[414])|(m[408]&~m[411]&~m[412]&~m[413]&m[414])|(m[408]&m[411]&~m[412]&~m[413]&m[414])|(m[408]&~m[411]&m[412]&~m[413]&m[414])|(~m[408]&~m[411]&~m[412]&m[413]&m[414])|(m[408]&~m[411]&~m[412]&m[413]&m[414])|(~m[408]&m[411]&~m[412]&m[413]&m[414])|(m[408]&m[411]&~m[412]&m[413]&m[414])|(~m[408]&~m[411]&m[412]&m[413]&m[414])|(m[408]&~m[411]&m[412]&m[413]&m[414])|(m[408]&m[411]&m[412]&m[413]&m[414]))):InitCond[113];
    m[415] = run?((((m[384]&~m[416]&~m[417]&~m[418]&~m[419])|(~m[384]&~m[416]&~m[417]&m[418]&~m[419])|(m[384]&m[416]&~m[417]&m[418]&~m[419])|(m[384]&~m[416]&m[417]&m[418]&~m[419])|(~m[384]&m[416]&~m[417]&~m[418]&m[419])|(~m[384]&~m[416]&m[417]&~m[418]&m[419])|(m[384]&m[416]&m[417]&~m[418]&m[419])|(~m[384]&m[416]&m[417]&m[418]&m[419]))&UnbiasedRNG[50])|((m[384]&~m[416]&~m[417]&m[418]&~m[419])|(~m[384]&~m[416]&~m[417]&~m[418]&m[419])|(m[384]&~m[416]&~m[417]&~m[418]&m[419])|(m[384]&m[416]&~m[417]&~m[418]&m[419])|(m[384]&~m[416]&m[417]&~m[418]&m[419])|(~m[384]&~m[416]&~m[417]&m[418]&m[419])|(m[384]&~m[416]&~m[417]&m[418]&m[419])|(~m[384]&m[416]&~m[417]&m[418]&m[419])|(m[384]&m[416]&~m[417]&m[418]&m[419])|(~m[384]&~m[416]&m[417]&m[418]&m[419])|(m[384]&~m[416]&m[417]&m[418]&m[419])|(m[384]&m[416]&m[417]&m[418]&m[419]))):InitCond[114];
    m[420] = run?((((m[418]&~m[421]&~m[422]&~m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&m[423]&~m[424])|(m[418]&m[421]&~m[422]&m[423]&~m[424])|(m[418]&~m[421]&m[422]&m[423]&~m[424])|(~m[418]&m[421]&~m[422]&~m[423]&m[424])|(~m[418]&~m[421]&m[422]&~m[423]&m[424])|(m[418]&m[421]&m[422]&~m[423]&m[424])|(~m[418]&m[421]&m[422]&m[423]&m[424]))&UnbiasedRNG[51])|((m[418]&~m[421]&~m[422]&m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&m[422]&~m[423]&m[424])|(~m[418]&~m[421]&~m[422]&m[423]&m[424])|(m[418]&~m[421]&~m[422]&m[423]&m[424])|(~m[418]&m[421]&~m[422]&m[423]&m[424])|(m[418]&m[421]&~m[422]&m[423]&m[424])|(~m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&m[421]&m[422]&m[423]&m[424]))):InitCond[115];
    m[425] = run?((((m[423]&~m[426]&~m[427]&~m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&m[428]&~m[429])|(m[423]&m[426]&~m[427]&m[428]&~m[429])|(m[423]&~m[426]&m[427]&m[428]&~m[429])|(~m[423]&m[426]&~m[427]&~m[428]&m[429])|(~m[423]&~m[426]&m[427]&~m[428]&m[429])|(m[423]&m[426]&m[427]&~m[428]&m[429])|(~m[423]&m[426]&m[427]&m[428]&m[429]))&UnbiasedRNG[52])|((m[423]&~m[426]&~m[427]&m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&m[427]&~m[428]&m[429])|(~m[423]&~m[426]&~m[427]&m[428]&m[429])|(m[423]&~m[426]&~m[427]&m[428]&m[429])|(~m[423]&m[426]&~m[427]&m[428]&m[429])|(m[423]&m[426]&~m[427]&m[428]&m[429])|(~m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&m[426]&m[427]&m[428]&m[429]))):InitCond[116];
    m[430] = run?((((m[428]&~m[431]&~m[432]&~m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&m[433]&~m[434])|(m[428]&m[431]&~m[432]&m[433]&~m[434])|(m[428]&~m[431]&m[432]&m[433]&~m[434])|(~m[428]&m[431]&~m[432]&~m[433]&m[434])|(~m[428]&~m[431]&m[432]&~m[433]&m[434])|(m[428]&m[431]&m[432]&~m[433]&m[434])|(~m[428]&m[431]&m[432]&m[433]&m[434]))&UnbiasedRNG[53])|((m[428]&~m[431]&~m[432]&m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&m[432]&~m[433]&m[434])|(~m[428]&~m[431]&~m[432]&m[433]&m[434])|(m[428]&~m[431]&~m[432]&m[433]&m[434])|(~m[428]&m[431]&~m[432]&m[433]&m[434])|(m[428]&m[431]&~m[432]&m[433]&m[434])|(~m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&m[431]&m[432]&m[433]&m[434]))):InitCond[117];
    m[435] = run?((((m[433]&~m[436]&~m[437]&~m[438]&~m[439])|(~m[433]&~m[436]&~m[437]&m[438]&~m[439])|(m[433]&m[436]&~m[437]&m[438]&~m[439])|(m[433]&~m[436]&m[437]&m[438]&~m[439])|(~m[433]&m[436]&~m[437]&~m[438]&m[439])|(~m[433]&~m[436]&m[437]&~m[438]&m[439])|(m[433]&m[436]&m[437]&~m[438]&m[439])|(~m[433]&m[436]&m[437]&m[438]&m[439]))&UnbiasedRNG[54])|((m[433]&~m[436]&~m[437]&m[438]&~m[439])|(~m[433]&~m[436]&~m[437]&~m[438]&m[439])|(m[433]&~m[436]&~m[437]&~m[438]&m[439])|(m[433]&m[436]&~m[437]&~m[438]&m[439])|(m[433]&~m[436]&m[437]&~m[438]&m[439])|(~m[433]&~m[436]&~m[437]&m[438]&m[439])|(m[433]&~m[436]&~m[437]&m[438]&m[439])|(~m[433]&m[436]&~m[437]&m[438]&m[439])|(m[433]&m[436]&~m[437]&m[438]&m[439])|(~m[433]&~m[436]&m[437]&m[438]&m[439])|(m[433]&~m[436]&m[437]&m[438]&m[439])|(m[433]&m[436]&m[437]&m[438]&m[439]))):InitCond[118];
    m[440] = run?((((m[438]&~m[441]&~m[442]&~m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&m[443]&~m[444])|(m[438]&m[441]&~m[442]&m[443]&~m[444])|(m[438]&~m[441]&m[442]&m[443]&~m[444])|(~m[438]&m[441]&~m[442]&~m[443]&m[444])|(~m[438]&~m[441]&m[442]&~m[443]&m[444])|(m[438]&m[441]&m[442]&~m[443]&m[444])|(~m[438]&m[441]&m[442]&m[443]&m[444]))&UnbiasedRNG[55])|((m[438]&~m[441]&~m[442]&m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&m[442]&~m[443]&m[444])|(~m[438]&~m[441]&~m[442]&m[443]&m[444])|(m[438]&~m[441]&~m[442]&m[443]&m[444])|(~m[438]&m[441]&~m[442]&m[443]&m[444])|(m[438]&m[441]&~m[442]&m[443]&m[444])|(~m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&m[441]&m[442]&m[443]&m[444]))):InitCond[119];
    m[445] = run?((((m[419]&~m[446]&~m[447]&~m[448]&~m[449])|(~m[419]&~m[446]&~m[447]&m[448]&~m[449])|(m[419]&m[446]&~m[447]&m[448]&~m[449])|(m[419]&~m[446]&m[447]&m[448]&~m[449])|(~m[419]&m[446]&~m[447]&~m[448]&m[449])|(~m[419]&~m[446]&m[447]&~m[448]&m[449])|(m[419]&m[446]&m[447]&~m[448]&m[449])|(~m[419]&m[446]&m[447]&m[448]&m[449]))&UnbiasedRNG[56])|((m[419]&~m[446]&~m[447]&m[448]&~m[449])|(~m[419]&~m[446]&~m[447]&~m[448]&m[449])|(m[419]&~m[446]&~m[447]&~m[448]&m[449])|(m[419]&m[446]&~m[447]&~m[448]&m[449])|(m[419]&~m[446]&m[447]&~m[448]&m[449])|(~m[419]&~m[446]&~m[447]&m[448]&m[449])|(m[419]&~m[446]&~m[447]&m[448]&m[449])|(~m[419]&m[446]&~m[447]&m[448]&m[449])|(m[419]&m[446]&~m[447]&m[448]&m[449])|(~m[419]&~m[446]&m[447]&m[448]&m[449])|(m[419]&~m[446]&m[447]&m[448]&m[449])|(m[419]&m[446]&m[447]&m[448]&m[449]))):InitCond[120];
    m[450] = run?((((m[448]&~m[451]&~m[452]&~m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&m[453]&~m[454])|(m[448]&m[451]&~m[452]&m[453]&~m[454])|(m[448]&~m[451]&m[452]&m[453]&~m[454])|(~m[448]&m[451]&~m[452]&~m[453]&m[454])|(~m[448]&~m[451]&m[452]&~m[453]&m[454])|(m[448]&m[451]&m[452]&~m[453]&m[454])|(~m[448]&m[451]&m[452]&m[453]&m[454]))&UnbiasedRNG[57])|((m[448]&~m[451]&~m[452]&m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&m[452]&~m[453]&m[454])|(~m[448]&~m[451]&~m[452]&m[453]&m[454])|(m[448]&~m[451]&~m[452]&m[453]&m[454])|(~m[448]&m[451]&~m[452]&m[453]&m[454])|(m[448]&m[451]&~m[452]&m[453]&m[454])|(~m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&m[451]&m[452]&m[453]&m[454]))):InitCond[121];
    m[455] = run?((((m[453]&~m[456]&~m[457]&~m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&m[458]&~m[459])|(m[453]&m[456]&~m[457]&m[458]&~m[459])|(m[453]&~m[456]&m[457]&m[458]&~m[459])|(~m[453]&m[456]&~m[457]&~m[458]&m[459])|(~m[453]&~m[456]&m[457]&~m[458]&m[459])|(m[453]&m[456]&m[457]&~m[458]&m[459])|(~m[453]&m[456]&m[457]&m[458]&m[459]))&UnbiasedRNG[58])|((m[453]&~m[456]&~m[457]&m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&m[457]&~m[458]&m[459])|(~m[453]&~m[456]&~m[457]&m[458]&m[459])|(m[453]&~m[456]&~m[457]&m[458]&m[459])|(~m[453]&m[456]&~m[457]&m[458]&m[459])|(m[453]&m[456]&~m[457]&m[458]&m[459])|(~m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&m[456]&m[457]&m[458]&m[459]))):InitCond[122];
    m[460] = run?((((m[458]&~m[461]&~m[462]&~m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&m[463]&~m[464])|(m[458]&m[461]&~m[462]&m[463]&~m[464])|(m[458]&~m[461]&m[462]&m[463]&~m[464])|(~m[458]&m[461]&~m[462]&~m[463]&m[464])|(~m[458]&~m[461]&m[462]&~m[463]&m[464])|(m[458]&m[461]&m[462]&~m[463]&m[464])|(~m[458]&m[461]&m[462]&m[463]&m[464]))&UnbiasedRNG[59])|((m[458]&~m[461]&~m[462]&m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&m[462]&~m[463]&m[464])|(~m[458]&~m[461]&~m[462]&m[463]&m[464])|(m[458]&~m[461]&~m[462]&m[463]&m[464])|(~m[458]&m[461]&~m[462]&m[463]&m[464])|(m[458]&m[461]&~m[462]&m[463]&m[464])|(~m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&m[461]&m[462]&m[463]&m[464]))):InitCond[123];
    m[465] = run?((((m[463]&~m[466]&~m[467]&~m[468]&~m[469])|(~m[463]&~m[466]&~m[467]&m[468]&~m[469])|(m[463]&m[466]&~m[467]&m[468]&~m[469])|(m[463]&~m[466]&m[467]&m[468]&~m[469])|(~m[463]&m[466]&~m[467]&~m[468]&m[469])|(~m[463]&~m[466]&m[467]&~m[468]&m[469])|(m[463]&m[466]&m[467]&~m[468]&m[469])|(~m[463]&m[466]&m[467]&m[468]&m[469]))&UnbiasedRNG[60])|((m[463]&~m[466]&~m[467]&m[468]&~m[469])|(~m[463]&~m[466]&~m[467]&~m[468]&m[469])|(m[463]&~m[466]&~m[467]&~m[468]&m[469])|(m[463]&m[466]&~m[467]&~m[468]&m[469])|(m[463]&~m[466]&m[467]&~m[468]&m[469])|(~m[463]&~m[466]&~m[467]&m[468]&m[469])|(m[463]&~m[466]&~m[467]&m[468]&m[469])|(~m[463]&m[466]&~m[467]&m[468]&m[469])|(m[463]&m[466]&~m[467]&m[468]&m[469])|(~m[463]&~m[466]&m[467]&m[468]&m[469])|(m[463]&~m[466]&m[467]&m[468]&m[469])|(m[463]&m[466]&m[467]&m[468]&m[469]))):InitCond[124];
    m[470] = run?((((m[449]&~m[471]&~m[472]&~m[473]&~m[474])|(~m[449]&~m[471]&~m[472]&m[473]&~m[474])|(m[449]&m[471]&~m[472]&m[473]&~m[474])|(m[449]&~m[471]&m[472]&m[473]&~m[474])|(~m[449]&m[471]&~m[472]&~m[473]&m[474])|(~m[449]&~m[471]&m[472]&~m[473]&m[474])|(m[449]&m[471]&m[472]&~m[473]&m[474])|(~m[449]&m[471]&m[472]&m[473]&m[474]))&UnbiasedRNG[61])|((m[449]&~m[471]&~m[472]&m[473]&~m[474])|(~m[449]&~m[471]&~m[472]&~m[473]&m[474])|(m[449]&~m[471]&~m[472]&~m[473]&m[474])|(m[449]&m[471]&~m[472]&~m[473]&m[474])|(m[449]&~m[471]&m[472]&~m[473]&m[474])|(~m[449]&~m[471]&~m[472]&m[473]&m[474])|(m[449]&~m[471]&~m[472]&m[473]&m[474])|(~m[449]&m[471]&~m[472]&m[473]&m[474])|(m[449]&m[471]&~m[472]&m[473]&m[474])|(~m[449]&~m[471]&m[472]&m[473]&m[474])|(m[449]&~m[471]&m[472]&m[473]&m[474])|(m[449]&m[471]&m[472]&m[473]&m[474]))):InitCond[125];
    m[475] = run?((((m[473]&~m[476]&~m[477]&~m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&m[478]&~m[479])|(m[473]&m[476]&~m[477]&m[478]&~m[479])|(m[473]&~m[476]&m[477]&m[478]&~m[479])|(~m[473]&m[476]&~m[477]&~m[478]&m[479])|(~m[473]&~m[476]&m[477]&~m[478]&m[479])|(m[473]&m[476]&m[477]&~m[478]&m[479])|(~m[473]&m[476]&m[477]&m[478]&m[479]))&UnbiasedRNG[62])|((m[473]&~m[476]&~m[477]&m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&m[477]&~m[478]&m[479])|(~m[473]&~m[476]&~m[477]&m[478]&m[479])|(m[473]&~m[476]&~m[477]&m[478]&m[479])|(~m[473]&m[476]&~m[477]&m[478]&m[479])|(m[473]&m[476]&~m[477]&m[478]&m[479])|(~m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&m[476]&m[477]&m[478]&m[479]))):InitCond[126];
    m[480] = run?((((m[478]&~m[481]&~m[482]&~m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&m[483]&~m[484])|(m[478]&m[481]&~m[482]&m[483]&~m[484])|(m[478]&~m[481]&m[482]&m[483]&~m[484])|(~m[478]&m[481]&~m[482]&~m[483]&m[484])|(~m[478]&~m[481]&m[482]&~m[483]&m[484])|(m[478]&m[481]&m[482]&~m[483]&m[484])|(~m[478]&m[481]&m[482]&m[483]&m[484]))&UnbiasedRNG[63])|((m[478]&~m[481]&~m[482]&m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&m[482]&~m[483]&m[484])|(~m[478]&~m[481]&~m[482]&m[483]&m[484])|(m[478]&~m[481]&~m[482]&m[483]&m[484])|(~m[478]&m[481]&~m[482]&m[483]&m[484])|(m[478]&m[481]&~m[482]&m[483]&m[484])|(~m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&m[481]&m[482]&m[483]&m[484]))):InitCond[127];
    m[485] = run?((((m[483]&~m[486]&~m[487]&~m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&m[488]&~m[489])|(m[483]&m[486]&~m[487]&m[488]&~m[489])|(m[483]&~m[486]&m[487]&m[488]&~m[489])|(~m[483]&m[486]&~m[487]&~m[488]&m[489])|(~m[483]&~m[486]&m[487]&~m[488]&m[489])|(m[483]&m[486]&m[487]&~m[488]&m[489])|(~m[483]&m[486]&m[487]&m[488]&m[489]))&UnbiasedRNG[64])|((m[483]&~m[486]&~m[487]&m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&m[487]&~m[488]&m[489])|(~m[483]&~m[486]&~m[487]&m[488]&m[489])|(m[483]&~m[486]&~m[487]&m[488]&m[489])|(~m[483]&m[486]&~m[487]&m[488]&m[489])|(m[483]&m[486]&~m[487]&m[488]&m[489])|(~m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&m[486]&m[487]&m[488]&m[489]))):InitCond[128];
    m[490] = run?((((m[474]&~m[491]&~m[492]&~m[493]&~m[494])|(~m[474]&~m[491]&~m[492]&m[493]&~m[494])|(m[474]&m[491]&~m[492]&m[493]&~m[494])|(m[474]&~m[491]&m[492]&m[493]&~m[494])|(~m[474]&m[491]&~m[492]&~m[493]&m[494])|(~m[474]&~m[491]&m[492]&~m[493]&m[494])|(m[474]&m[491]&m[492]&~m[493]&m[494])|(~m[474]&m[491]&m[492]&m[493]&m[494]))&UnbiasedRNG[65])|((m[474]&~m[491]&~m[492]&m[493]&~m[494])|(~m[474]&~m[491]&~m[492]&~m[493]&m[494])|(m[474]&~m[491]&~m[492]&~m[493]&m[494])|(m[474]&m[491]&~m[492]&~m[493]&m[494])|(m[474]&~m[491]&m[492]&~m[493]&m[494])|(~m[474]&~m[491]&~m[492]&m[493]&m[494])|(m[474]&~m[491]&~m[492]&m[493]&m[494])|(~m[474]&m[491]&~m[492]&m[493]&m[494])|(m[474]&m[491]&~m[492]&m[493]&m[494])|(~m[474]&~m[491]&m[492]&m[493]&m[494])|(m[474]&~m[491]&m[492]&m[493]&m[494])|(m[474]&m[491]&m[492]&m[493]&m[494]))):InitCond[129];
    m[495] = run?((((m[493]&~m[496]&~m[497]&~m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&m[498]&~m[499])|(m[493]&m[496]&~m[497]&m[498]&~m[499])|(m[493]&~m[496]&m[497]&m[498]&~m[499])|(~m[493]&m[496]&~m[497]&~m[498]&m[499])|(~m[493]&~m[496]&m[497]&~m[498]&m[499])|(m[493]&m[496]&m[497]&~m[498]&m[499])|(~m[493]&m[496]&m[497]&m[498]&m[499]))&UnbiasedRNG[66])|((m[493]&~m[496]&~m[497]&m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&m[497]&~m[498]&m[499])|(~m[493]&~m[496]&~m[497]&m[498]&m[499])|(m[493]&~m[496]&~m[497]&m[498]&m[499])|(~m[493]&m[496]&~m[497]&m[498]&m[499])|(m[493]&m[496]&~m[497]&m[498]&m[499])|(~m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&m[496]&m[497]&m[498]&m[499]))):InitCond[130];
    m[500] = run?((((m[498]&~m[501]&~m[502]&~m[503]&~m[504])|(~m[498]&~m[501]&~m[502]&m[503]&~m[504])|(m[498]&m[501]&~m[502]&m[503]&~m[504])|(m[498]&~m[501]&m[502]&m[503]&~m[504])|(~m[498]&m[501]&~m[502]&~m[503]&m[504])|(~m[498]&~m[501]&m[502]&~m[503]&m[504])|(m[498]&m[501]&m[502]&~m[503]&m[504])|(~m[498]&m[501]&m[502]&m[503]&m[504]))&UnbiasedRNG[67])|((m[498]&~m[501]&~m[502]&m[503]&~m[504])|(~m[498]&~m[501]&~m[502]&~m[503]&m[504])|(m[498]&~m[501]&~m[502]&~m[503]&m[504])|(m[498]&m[501]&~m[502]&~m[503]&m[504])|(m[498]&~m[501]&m[502]&~m[503]&m[504])|(~m[498]&~m[501]&~m[502]&m[503]&m[504])|(m[498]&~m[501]&~m[502]&m[503]&m[504])|(~m[498]&m[501]&~m[502]&m[503]&m[504])|(m[498]&m[501]&~m[502]&m[503]&m[504])|(~m[498]&~m[501]&m[502]&m[503]&m[504])|(m[498]&~m[501]&m[502]&m[503]&m[504])|(m[498]&m[501]&m[502]&m[503]&m[504]))):InitCond[131];
    m[505] = run?((((m[494]&~m[506]&~m[507]&~m[508]&~m[509])|(~m[494]&~m[506]&~m[507]&m[508]&~m[509])|(m[494]&m[506]&~m[507]&m[508]&~m[509])|(m[494]&~m[506]&m[507]&m[508]&~m[509])|(~m[494]&m[506]&~m[507]&~m[508]&m[509])|(~m[494]&~m[506]&m[507]&~m[508]&m[509])|(m[494]&m[506]&m[507]&~m[508]&m[509])|(~m[494]&m[506]&m[507]&m[508]&m[509]))&UnbiasedRNG[68])|((m[494]&~m[506]&~m[507]&m[508]&~m[509])|(~m[494]&~m[506]&~m[507]&~m[508]&m[509])|(m[494]&~m[506]&~m[507]&~m[508]&m[509])|(m[494]&m[506]&~m[507]&~m[508]&m[509])|(m[494]&~m[506]&m[507]&~m[508]&m[509])|(~m[494]&~m[506]&~m[507]&m[508]&m[509])|(m[494]&~m[506]&~m[507]&m[508]&m[509])|(~m[494]&m[506]&~m[507]&m[508]&m[509])|(m[494]&m[506]&~m[507]&m[508]&m[509])|(~m[494]&~m[506]&m[507]&m[508]&m[509])|(m[494]&~m[506]&m[507]&m[508]&m[509])|(m[494]&m[506]&m[507]&m[508]&m[509]))):InitCond[132];
    m[510] = run?((((m[508]&~m[511]&~m[512]&~m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&m[513]&~m[514])|(m[508]&m[511]&~m[512]&m[513]&~m[514])|(m[508]&~m[511]&m[512]&m[513]&~m[514])|(~m[508]&m[511]&~m[512]&~m[513]&m[514])|(~m[508]&~m[511]&m[512]&~m[513]&m[514])|(m[508]&m[511]&m[512]&~m[513]&m[514])|(~m[508]&m[511]&m[512]&m[513]&m[514]))&UnbiasedRNG[69])|((m[508]&~m[511]&~m[512]&m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&m[512]&~m[513]&m[514])|(~m[508]&~m[511]&~m[512]&m[513]&m[514])|(m[508]&~m[511]&~m[512]&m[513]&m[514])|(~m[508]&m[511]&~m[512]&m[513]&m[514])|(m[508]&m[511]&~m[512]&m[513]&m[514])|(~m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&m[511]&m[512]&m[513]&m[514]))):InitCond[133];
    m[515] = run?((((m[509]&~m[516]&~m[517]&~m[518]&~m[519])|(~m[509]&~m[516]&~m[517]&m[518]&~m[519])|(m[509]&m[516]&~m[517]&m[518]&~m[519])|(m[509]&~m[516]&m[517]&m[518]&~m[519])|(~m[509]&m[516]&~m[517]&~m[518]&m[519])|(~m[509]&~m[516]&m[517]&~m[518]&m[519])|(m[509]&m[516]&m[517]&~m[518]&m[519])|(~m[509]&m[516]&m[517]&m[518]&m[519]))&UnbiasedRNG[70])|((m[509]&~m[516]&~m[517]&m[518]&~m[519])|(~m[509]&~m[516]&~m[517]&~m[518]&m[519])|(m[509]&~m[516]&~m[517]&~m[518]&m[519])|(m[509]&m[516]&~m[517]&~m[518]&m[519])|(m[509]&~m[516]&m[517]&~m[518]&m[519])|(~m[509]&~m[516]&~m[517]&m[518]&m[519])|(m[509]&~m[516]&~m[517]&m[518]&m[519])|(~m[509]&m[516]&~m[517]&m[518]&m[519])|(m[509]&m[516]&~m[517]&m[518]&m[519])|(~m[509]&~m[516]&m[517]&m[518]&m[519])|(m[509]&~m[516]&m[517]&m[518]&m[519])|(m[509]&m[516]&m[517]&m[518]&m[519]))):InitCond[134];
end

always @(posedge color1_clk) begin
    m[16] = run?((((m[0]&m[48]&~m[49]&~m[50]&~m[51])|(m[0]&~m[48]&m[49]&~m[50]&~m[51])|(~m[0]&m[48]&m[49]&~m[50]&~m[51])|(m[0]&~m[48]&~m[49]&m[50]&~m[51])|(~m[0]&m[48]&~m[49]&m[50]&~m[51])|(~m[0]&~m[48]&m[49]&m[50]&~m[51])|(m[0]&~m[48]&~m[49]&~m[50]&m[51])|(~m[0]&m[48]&~m[49]&~m[50]&m[51])|(~m[0]&~m[48]&m[49]&~m[50]&m[51])|(~m[0]&~m[48]&~m[49]&m[50]&m[51]))&BiasedRNG[64])|(((m[0]&m[48]&m[49]&~m[50]&~m[51])|(m[0]&m[48]&~m[49]&m[50]&~m[51])|(m[0]&~m[48]&m[49]&m[50]&~m[51])|(~m[0]&m[48]&m[49]&m[50]&~m[51])|(m[0]&m[48]&~m[49]&~m[50]&m[51])|(m[0]&~m[48]&m[49]&~m[50]&m[51])|(~m[0]&m[48]&m[49]&~m[50]&m[51])|(m[0]&~m[48]&~m[49]&m[50]&m[51])|(~m[0]&m[48]&~m[49]&m[50]&m[51])|(~m[0]&~m[48]&m[49]&m[50]&m[51]))&~BiasedRNG[64])|((m[0]&m[48]&m[49]&m[50]&~m[51])|(m[0]&m[48]&m[49]&~m[50]&m[51])|(m[0]&m[48]&~m[49]&m[50]&m[51])|(m[0]&~m[48]&m[49]&m[50]&m[51])|(~m[0]&m[48]&m[49]&m[50]&m[51])|(m[0]&m[48]&m[49]&m[50]&m[51]))):InitCond[135];
    m[17] = run?((((m[0]&m[52]&~m[53]&~m[54]&~m[55])|(m[0]&~m[52]&m[53]&~m[54]&~m[55])|(~m[0]&m[52]&m[53]&~m[54]&~m[55])|(m[0]&~m[52]&~m[53]&m[54]&~m[55])|(~m[0]&m[52]&~m[53]&m[54]&~m[55])|(~m[0]&~m[52]&m[53]&m[54]&~m[55])|(m[0]&~m[52]&~m[53]&~m[54]&m[55])|(~m[0]&m[52]&~m[53]&~m[54]&m[55])|(~m[0]&~m[52]&m[53]&~m[54]&m[55])|(~m[0]&~m[52]&~m[53]&m[54]&m[55]))&BiasedRNG[65])|(((m[0]&m[52]&m[53]&~m[54]&~m[55])|(m[0]&m[52]&~m[53]&m[54]&~m[55])|(m[0]&~m[52]&m[53]&m[54]&~m[55])|(~m[0]&m[52]&m[53]&m[54]&~m[55])|(m[0]&m[52]&~m[53]&~m[54]&m[55])|(m[0]&~m[52]&m[53]&~m[54]&m[55])|(~m[0]&m[52]&m[53]&~m[54]&m[55])|(m[0]&~m[52]&~m[53]&m[54]&m[55])|(~m[0]&m[52]&~m[53]&m[54]&m[55])|(~m[0]&~m[52]&m[53]&m[54]&m[55]))&~BiasedRNG[65])|((m[0]&m[52]&m[53]&m[54]&~m[55])|(m[0]&m[52]&m[53]&~m[54]&m[55])|(m[0]&m[52]&~m[53]&m[54]&m[55])|(m[0]&~m[52]&m[53]&m[54]&m[55])|(~m[0]&m[52]&m[53]&m[54]&m[55])|(m[0]&m[52]&m[53]&m[54]&m[55]))):InitCond[136];
    m[18] = run?((((m[1]&m[56]&~m[57]&~m[58]&~m[59])|(m[1]&~m[56]&m[57]&~m[58]&~m[59])|(~m[1]&m[56]&m[57]&~m[58]&~m[59])|(m[1]&~m[56]&~m[57]&m[58]&~m[59])|(~m[1]&m[56]&~m[57]&m[58]&~m[59])|(~m[1]&~m[56]&m[57]&m[58]&~m[59])|(m[1]&~m[56]&~m[57]&~m[58]&m[59])|(~m[1]&m[56]&~m[57]&~m[58]&m[59])|(~m[1]&~m[56]&m[57]&~m[58]&m[59])|(~m[1]&~m[56]&~m[57]&m[58]&m[59]))&BiasedRNG[66])|(((m[1]&m[56]&m[57]&~m[58]&~m[59])|(m[1]&m[56]&~m[57]&m[58]&~m[59])|(m[1]&~m[56]&m[57]&m[58]&~m[59])|(~m[1]&m[56]&m[57]&m[58]&~m[59])|(m[1]&m[56]&~m[57]&~m[58]&m[59])|(m[1]&~m[56]&m[57]&~m[58]&m[59])|(~m[1]&m[56]&m[57]&~m[58]&m[59])|(m[1]&~m[56]&~m[57]&m[58]&m[59])|(~m[1]&m[56]&~m[57]&m[58]&m[59])|(~m[1]&~m[56]&m[57]&m[58]&m[59]))&~BiasedRNG[66])|((m[1]&m[56]&m[57]&m[58]&~m[59])|(m[1]&m[56]&m[57]&~m[58]&m[59])|(m[1]&m[56]&~m[57]&m[58]&m[59])|(m[1]&~m[56]&m[57]&m[58]&m[59])|(~m[1]&m[56]&m[57]&m[58]&m[59])|(m[1]&m[56]&m[57]&m[58]&m[59]))):InitCond[137];
    m[19] = run?((((m[1]&m[60]&~m[61]&~m[62]&~m[63])|(m[1]&~m[60]&m[61]&~m[62]&~m[63])|(~m[1]&m[60]&m[61]&~m[62]&~m[63])|(m[1]&~m[60]&~m[61]&m[62]&~m[63])|(~m[1]&m[60]&~m[61]&m[62]&~m[63])|(~m[1]&~m[60]&m[61]&m[62]&~m[63])|(m[1]&~m[60]&~m[61]&~m[62]&m[63])|(~m[1]&m[60]&~m[61]&~m[62]&m[63])|(~m[1]&~m[60]&m[61]&~m[62]&m[63])|(~m[1]&~m[60]&~m[61]&m[62]&m[63]))&BiasedRNG[67])|(((m[1]&m[60]&m[61]&~m[62]&~m[63])|(m[1]&m[60]&~m[61]&m[62]&~m[63])|(m[1]&~m[60]&m[61]&m[62]&~m[63])|(~m[1]&m[60]&m[61]&m[62]&~m[63])|(m[1]&m[60]&~m[61]&~m[62]&m[63])|(m[1]&~m[60]&m[61]&~m[62]&m[63])|(~m[1]&m[60]&m[61]&~m[62]&m[63])|(m[1]&~m[60]&~m[61]&m[62]&m[63])|(~m[1]&m[60]&~m[61]&m[62]&m[63])|(~m[1]&~m[60]&m[61]&m[62]&m[63]))&~BiasedRNG[67])|((m[1]&m[60]&m[61]&m[62]&~m[63])|(m[1]&m[60]&m[61]&~m[62]&m[63])|(m[1]&m[60]&~m[61]&m[62]&m[63])|(m[1]&~m[60]&m[61]&m[62]&m[63])|(~m[1]&m[60]&m[61]&m[62]&m[63])|(m[1]&m[60]&m[61]&m[62]&m[63]))):InitCond[138];
    m[20] = run?((((m[2]&m[64]&~m[65]&~m[66]&~m[67])|(m[2]&~m[64]&m[65]&~m[66]&~m[67])|(~m[2]&m[64]&m[65]&~m[66]&~m[67])|(m[2]&~m[64]&~m[65]&m[66]&~m[67])|(~m[2]&m[64]&~m[65]&m[66]&~m[67])|(~m[2]&~m[64]&m[65]&m[66]&~m[67])|(m[2]&~m[64]&~m[65]&~m[66]&m[67])|(~m[2]&m[64]&~m[65]&~m[66]&m[67])|(~m[2]&~m[64]&m[65]&~m[66]&m[67])|(~m[2]&~m[64]&~m[65]&m[66]&m[67]))&BiasedRNG[68])|(((m[2]&m[64]&m[65]&~m[66]&~m[67])|(m[2]&m[64]&~m[65]&m[66]&~m[67])|(m[2]&~m[64]&m[65]&m[66]&~m[67])|(~m[2]&m[64]&m[65]&m[66]&~m[67])|(m[2]&m[64]&~m[65]&~m[66]&m[67])|(m[2]&~m[64]&m[65]&~m[66]&m[67])|(~m[2]&m[64]&m[65]&~m[66]&m[67])|(m[2]&~m[64]&~m[65]&m[66]&m[67])|(~m[2]&m[64]&~m[65]&m[66]&m[67])|(~m[2]&~m[64]&m[65]&m[66]&m[67]))&~BiasedRNG[68])|((m[2]&m[64]&m[65]&m[66]&~m[67])|(m[2]&m[64]&m[65]&~m[66]&m[67])|(m[2]&m[64]&~m[65]&m[66]&m[67])|(m[2]&~m[64]&m[65]&m[66]&m[67])|(~m[2]&m[64]&m[65]&m[66]&m[67])|(m[2]&m[64]&m[65]&m[66]&m[67]))):InitCond[139];
    m[21] = run?((((m[2]&m[68]&~m[69]&~m[70]&~m[71])|(m[2]&~m[68]&m[69]&~m[70]&~m[71])|(~m[2]&m[68]&m[69]&~m[70]&~m[71])|(m[2]&~m[68]&~m[69]&m[70]&~m[71])|(~m[2]&m[68]&~m[69]&m[70]&~m[71])|(~m[2]&~m[68]&m[69]&m[70]&~m[71])|(m[2]&~m[68]&~m[69]&~m[70]&m[71])|(~m[2]&m[68]&~m[69]&~m[70]&m[71])|(~m[2]&~m[68]&m[69]&~m[70]&m[71])|(~m[2]&~m[68]&~m[69]&m[70]&m[71]))&BiasedRNG[69])|(((m[2]&m[68]&m[69]&~m[70]&~m[71])|(m[2]&m[68]&~m[69]&m[70]&~m[71])|(m[2]&~m[68]&m[69]&m[70]&~m[71])|(~m[2]&m[68]&m[69]&m[70]&~m[71])|(m[2]&m[68]&~m[69]&~m[70]&m[71])|(m[2]&~m[68]&m[69]&~m[70]&m[71])|(~m[2]&m[68]&m[69]&~m[70]&m[71])|(m[2]&~m[68]&~m[69]&m[70]&m[71])|(~m[2]&m[68]&~m[69]&m[70]&m[71])|(~m[2]&~m[68]&m[69]&m[70]&m[71]))&~BiasedRNG[69])|((m[2]&m[68]&m[69]&m[70]&~m[71])|(m[2]&m[68]&m[69]&~m[70]&m[71])|(m[2]&m[68]&~m[69]&m[70]&m[71])|(m[2]&~m[68]&m[69]&m[70]&m[71])|(~m[2]&m[68]&m[69]&m[70]&m[71])|(m[2]&m[68]&m[69]&m[70]&m[71]))):InitCond[140];
    m[22] = run?((((m[3]&m[72]&~m[73]&~m[74]&~m[75])|(m[3]&~m[72]&m[73]&~m[74]&~m[75])|(~m[3]&m[72]&m[73]&~m[74]&~m[75])|(m[3]&~m[72]&~m[73]&m[74]&~m[75])|(~m[3]&m[72]&~m[73]&m[74]&~m[75])|(~m[3]&~m[72]&m[73]&m[74]&~m[75])|(m[3]&~m[72]&~m[73]&~m[74]&m[75])|(~m[3]&m[72]&~m[73]&~m[74]&m[75])|(~m[3]&~m[72]&m[73]&~m[74]&m[75])|(~m[3]&~m[72]&~m[73]&m[74]&m[75]))&BiasedRNG[70])|(((m[3]&m[72]&m[73]&~m[74]&~m[75])|(m[3]&m[72]&~m[73]&m[74]&~m[75])|(m[3]&~m[72]&m[73]&m[74]&~m[75])|(~m[3]&m[72]&m[73]&m[74]&~m[75])|(m[3]&m[72]&~m[73]&~m[74]&m[75])|(m[3]&~m[72]&m[73]&~m[74]&m[75])|(~m[3]&m[72]&m[73]&~m[74]&m[75])|(m[3]&~m[72]&~m[73]&m[74]&m[75])|(~m[3]&m[72]&~m[73]&m[74]&m[75])|(~m[3]&~m[72]&m[73]&m[74]&m[75]))&~BiasedRNG[70])|((m[3]&m[72]&m[73]&m[74]&~m[75])|(m[3]&m[72]&m[73]&~m[74]&m[75])|(m[3]&m[72]&~m[73]&m[74]&m[75])|(m[3]&~m[72]&m[73]&m[74]&m[75])|(~m[3]&m[72]&m[73]&m[74]&m[75])|(m[3]&m[72]&m[73]&m[74]&m[75]))):InitCond[141];
    m[23] = run?((((m[3]&m[76]&~m[77]&~m[78]&~m[79])|(m[3]&~m[76]&m[77]&~m[78]&~m[79])|(~m[3]&m[76]&m[77]&~m[78]&~m[79])|(m[3]&~m[76]&~m[77]&m[78]&~m[79])|(~m[3]&m[76]&~m[77]&m[78]&~m[79])|(~m[3]&~m[76]&m[77]&m[78]&~m[79])|(m[3]&~m[76]&~m[77]&~m[78]&m[79])|(~m[3]&m[76]&~m[77]&~m[78]&m[79])|(~m[3]&~m[76]&m[77]&~m[78]&m[79])|(~m[3]&~m[76]&~m[77]&m[78]&m[79]))&BiasedRNG[71])|(((m[3]&m[76]&m[77]&~m[78]&~m[79])|(m[3]&m[76]&~m[77]&m[78]&~m[79])|(m[3]&~m[76]&m[77]&m[78]&~m[79])|(~m[3]&m[76]&m[77]&m[78]&~m[79])|(m[3]&m[76]&~m[77]&~m[78]&m[79])|(m[3]&~m[76]&m[77]&~m[78]&m[79])|(~m[3]&m[76]&m[77]&~m[78]&m[79])|(m[3]&~m[76]&~m[77]&m[78]&m[79])|(~m[3]&m[76]&~m[77]&m[78]&m[79])|(~m[3]&~m[76]&m[77]&m[78]&m[79]))&~BiasedRNG[71])|((m[3]&m[76]&m[77]&m[78]&~m[79])|(m[3]&m[76]&m[77]&~m[78]&m[79])|(m[3]&m[76]&~m[77]&m[78]&m[79])|(m[3]&~m[76]&m[77]&m[78]&m[79])|(~m[3]&m[76]&m[77]&m[78]&m[79])|(m[3]&m[76]&m[77]&m[78]&m[79]))):InitCond[142];
    m[24] = run?((((m[4]&m[80]&~m[81]&~m[82]&~m[83])|(m[4]&~m[80]&m[81]&~m[82]&~m[83])|(~m[4]&m[80]&m[81]&~m[82]&~m[83])|(m[4]&~m[80]&~m[81]&m[82]&~m[83])|(~m[4]&m[80]&~m[81]&m[82]&~m[83])|(~m[4]&~m[80]&m[81]&m[82]&~m[83])|(m[4]&~m[80]&~m[81]&~m[82]&m[83])|(~m[4]&m[80]&~m[81]&~m[82]&m[83])|(~m[4]&~m[80]&m[81]&~m[82]&m[83])|(~m[4]&~m[80]&~m[81]&m[82]&m[83]))&BiasedRNG[72])|(((m[4]&m[80]&m[81]&~m[82]&~m[83])|(m[4]&m[80]&~m[81]&m[82]&~m[83])|(m[4]&~m[80]&m[81]&m[82]&~m[83])|(~m[4]&m[80]&m[81]&m[82]&~m[83])|(m[4]&m[80]&~m[81]&~m[82]&m[83])|(m[4]&~m[80]&m[81]&~m[82]&m[83])|(~m[4]&m[80]&m[81]&~m[82]&m[83])|(m[4]&~m[80]&~m[81]&m[82]&m[83])|(~m[4]&m[80]&~m[81]&m[82]&m[83])|(~m[4]&~m[80]&m[81]&m[82]&m[83]))&~BiasedRNG[72])|((m[4]&m[80]&m[81]&m[82]&~m[83])|(m[4]&m[80]&m[81]&~m[82]&m[83])|(m[4]&m[80]&~m[81]&m[82]&m[83])|(m[4]&~m[80]&m[81]&m[82]&m[83])|(~m[4]&m[80]&m[81]&m[82]&m[83])|(m[4]&m[80]&m[81]&m[82]&m[83]))):InitCond[143];
    m[25] = run?((((m[4]&m[84]&~m[85]&~m[86]&~m[87])|(m[4]&~m[84]&m[85]&~m[86]&~m[87])|(~m[4]&m[84]&m[85]&~m[86]&~m[87])|(m[4]&~m[84]&~m[85]&m[86]&~m[87])|(~m[4]&m[84]&~m[85]&m[86]&~m[87])|(~m[4]&~m[84]&m[85]&m[86]&~m[87])|(m[4]&~m[84]&~m[85]&~m[86]&m[87])|(~m[4]&m[84]&~m[85]&~m[86]&m[87])|(~m[4]&~m[84]&m[85]&~m[86]&m[87])|(~m[4]&~m[84]&~m[85]&m[86]&m[87]))&BiasedRNG[73])|(((m[4]&m[84]&m[85]&~m[86]&~m[87])|(m[4]&m[84]&~m[85]&m[86]&~m[87])|(m[4]&~m[84]&m[85]&m[86]&~m[87])|(~m[4]&m[84]&m[85]&m[86]&~m[87])|(m[4]&m[84]&~m[85]&~m[86]&m[87])|(m[4]&~m[84]&m[85]&~m[86]&m[87])|(~m[4]&m[84]&m[85]&~m[86]&m[87])|(m[4]&~m[84]&~m[85]&m[86]&m[87])|(~m[4]&m[84]&~m[85]&m[86]&m[87])|(~m[4]&~m[84]&m[85]&m[86]&m[87]))&~BiasedRNG[73])|((m[4]&m[84]&m[85]&m[86]&~m[87])|(m[4]&m[84]&m[85]&~m[86]&m[87])|(m[4]&m[84]&~m[85]&m[86]&m[87])|(m[4]&~m[84]&m[85]&m[86]&m[87])|(~m[4]&m[84]&m[85]&m[86]&m[87])|(m[4]&m[84]&m[85]&m[86]&m[87]))):InitCond[144];
    m[26] = run?((((m[5]&m[88]&~m[89]&~m[90]&~m[91])|(m[5]&~m[88]&m[89]&~m[90]&~m[91])|(~m[5]&m[88]&m[89]&~m[90]&~m[91])|(m[5]&~m[88]&~m[89]&m[90]&~m[91])|(~m[5]&m[88]&~m[89]&m[90]&~m[91])|(~m[5]&~m[88]&m[89]&m[90]&~m[91])|(m[5]&~m[88]&~m[89]&~m[90]&m[91])|(~m[5]&m[88]&~m[89]&~m[90]&m[91])|(~m[5]&~m[88]&m[89]&~m[90]&m[91])|(~m[5]&~m[88]&~m[89]&m[90]&m[91]))&BiasedRNG[74])|(((m[5]&m[88]&m[89]&~m[90]&~m[91])|(m[5]&m[88]&~m[89]&m[90]&~m[91])|(m[5]&~m[88]&m[89]&m[90]&~m[91])|(~m[5]&m[88]&m[89]&m[90]&~m[91])|(m[5]&m[88]&~m[89]&~m[90]&m[91])|(m[5]&~m[88]&m[89]&~m[90]&m[91])|(~m[5]&m[88]&m[89]&~m[90]&m[91])|(m[5]&~m[88]&~m[89]&m[90]&m[91])|(~m[5]&m[88]&~m[89]&m[90]&m[91])|(~m[5]&~m[88]&m[89]&m[90]&m[91]))&~BiasedRNG[74])|((m[5]&m[88]&m[89]&m[90]&~m[91])|(m[5]&m[88]&m[89]&~m[90]&m[91])|(m[5]&m[88]&~m[89]&m[90]&m[91])|(m[5]&~m[88]&m[89]&m[90]&m[91])|(~m[5]&m[88]&m[89]&m[90]&m[91])|(m[5]&m[88]&m[89]&m[90]&m[91]))):InitCond[145];
    m[27] = run?((((m[5]&m[92]&~m[93]&~m[94]&~m[95])|(m[5]&~m[92]&m[93]&~m[94]&~m[95])|(~m[5]&m[92]&m[93]&~m[94]&~m[95])|(m[5]&~m[92]&~m[93]&m[94]&~m[95])|(~m[5]&m[92]&~m[93]&m[94]&~m[95])|(~m[5]&~m[92]&m[93]&m[94]&~m[95])|(m[5]&~m[92]&~m[93]&~m[94]&m[95])|(~m[5]&m[92]&~m[93]&~m[94]&m[95])|(~m[5]&~m[92]&m[93]&~m[94]&m[95])|(~m[5]&~m[92]&~m[93]&m[94]&m[95]))&BiasedRNG[75])|(((m[5]&m[92]&m[93]&~m[94]&~m[95])|(m[5]&m[92]&~m[93]&m[94]&~m[95])|(m[5]&~m[92]&m[93]&m[94]&~m[95])|(~m[5]&m[92]&m[93]&m[94]&~m[95])|(m[5]&m[92]&~m[93]&~m[94]&m[95])|(m[5]&~m[92]&m[93]&~m[94]&m[95])|(~m[5]&m[92]&m[93]&~m[94]&m[95])|(m[5]&~m[92]&~m[93]&m[94]&m[95])|(~m[5]&m[92]&~m[93]&m[94]&m[95])|(~m[5]&~m[92]&m[93]&m[94]&m[95]))&~BiasedRNG[75])|((m[5]&m[92]&m[93]&m[94]&~m[95])|(m[5]&m[92]&m[93]&~m[94]&m[95])|(m[5]&m[92]&~m[93]&m[94]&m[95])|(m[5]&~m[92]&m[93]&m[94]&m[95])|(~m[5]&m[92]&m[93]&m[94]&m[95])|(m[5]&m[92]&m[93]&m[94]&m[95]))):InitCond[146];
    m[28] = run?((((m[6]&m[96]&~m[97]&~m[98]&~m[99])|(m[6]&~m[96]&m[97]&~m[98]&~m[99])|(~m[6]&m[96]&m[97]&~m[98]&~m[99])|(m[6]&~m[96]&~m[97]&m[98]&~m[99])|(~m[6]&m[96]&~m[97]&m[98]&~m[99])|(~m[6]&~m[96]&m[97]&m[98]&~m[99])|(m[6]&~m[96]&~m[97]&~m[98]&m[99])|(~m[6]&m[96]&~m[97]&~m[98]&m[99])|(~m[6]&~m[96]&m[97]&~m[98]&m[99])|(~m[6]&~m[96]&~m[97]&m[98]&m[99]))&BiasedRNG[76])|(((m[6]&m[96]&m[97]&~m[98]&~m[99])|(m[6]&m[96]&~m[97]&m[98]&~m[99])|(m[6]&~m[96]&m[97]&m[98]&~m[99])|(~m[6]&m[96]&m[97]&m[98]&~m[99])|(m[6]&m[96]&~m[97]&~m[98]&m[99])|(m[6]&~m[96]&m[97]&~m[98]&m[99])|(~m[6]&m[96]&m[97]&~m[98]&m[99])|(m[6]&~m[96]&~m[97]&m[98]&m[99])|(~m[6]&m[96]&~m[97]&m[98]&m[99])|(~m[6]&~m[96]&m[97]&m[98]&m[99]))&~BiasedRNG[76])|((m[6]&m[96]&m[97]&m[98]&~m[99])|(m[6]&m[96]&m[97]&~m[98]&m[99])|(m[6]&m[96]&~m[97]&m[98]&m[99])|(m[6]&~m[96]&m[97]&m[98]&m[99])|(~m[6]&m[96]&m[97]&m[98]&m[99])|(m[6]&m[96]&m[97]&m[98]&m[99]))):InitCond[147];
    m[29] = run?((((m[6]&m[100]&~m[101]&~m[102]&~m[103])|(m[6]&~m[100]&m[101]&~m[102]&~m[103])|(~m[6]&m[100]&m[101]&~m[102]&~m[103])|(m[6]&~m[100]&~m[101]&m[102]&~m[103])|(~m[6]&m[100]&~m[101]&m[102]&~m[103])|(~m[6]&~m[100]&m[101]&m[102]&~m[103])|(m[6]&~m[100]&~m[101]&~m[102]&m[103])|(~m[6]&m[100]&~m[101]&~m[102]&m[103])|(~m[6]&~m[100]&m[101]&~m[102]&m[103])|(~m[6]&~m[100]&~m[101]&m[102]&m[103]))&BiasedRNG[77])|(((m[6]&m[100]&m[101]&~m[102]&~m[103])|(m[6]&m[100]&~m[101]&m[102]&~m[103])|(m[6]&~m[100]&m[101]&m[102]&~m[103])|(~m[6]&m[100]&m[101]&m[102]&~m[103])|(m[6]&m[100]&~m[101]&~m[102]&m[103])|(m[6]&~m[100]&m[101]&~m[102]&m[103])|(~m[6]&m[100]&m[101]&~m[102]&m[103])|(m[6]&~m[100]&~m[101]&m[102]&m[103])|(~m[6]&m[100]&~m[101]&m[102]&m[103])|(~m[6]&~m[100]&m[101]&m[102]&m[103]))&~BiasedRNG[77])|((m[6]&m[100]&m[101]&m[102]&~m[103])|(m[6]&m[100]&m[101]&~m[102]&m[103])|(m[6]&m[100]&~m[101]&m[102]&m[103])|(m[6]&~m[100]&m[101]&m[102]&m[103])|(~m[6]&m[100]&m[101]&m[102]&m[103])|(m[6]&m[100]&m[101]&m[102]&m[103]))):InitCond[148];
    m[30] = run?((((m[7]&m[104]&~m[105]&~m[106]&~m[107])|(m[7]&~m[104]&m[105]&~m[106]&~m[107])|(~m[7]&m[104]&m[105]&~m[106]&~m[107])|(m[7]&~m[104]&~m[105]&m[106]&~m[107])|(~m[7]&m[104]&~m[105]&m[106]&~m[107])|(~m[7]&~m[104]&m[105]&m[106]&~m[107])|(m[7]&~m[104]&~m[105]&~m[106]&m[107])|(~m[7]&m[104]&~m[105]&~m[106]&m[107])|(~m[7]&~m[104]&m[105]&~m[106]&m[107])|(~m[7]&~m[104]&~m[105]&m[106]&m[107]))&BiasedRNG[78])|(((m[7]&m[104]&m[105]&~m[106]&~m[107])|(m[7]&m[104]&~m[105]&m[106]&~m[107])|(m[7]&~m[104]&m[105]&m[106]&~m[107])|(~m[7]&m[104]&m[105]&m[106]&~m[107])|(m[7]&m[104]&~m[105]&~m[106]&m[107])|(m[7]&~m[104]&m[105]&~m[106]&m[107])|(~m[7]&m[104]&m[105]&~m[106]&m[107])|(m[7]&~m[104]&~m[105]&m[106]&m[107])|(~m[7]&m[104]&~m[105]&m[106]&m[107])|(~m[7]&~m[104]&m[105]&m[106]&m[107]))&~BiasedRNG[78])|((m[7]&m[104]&m[105]&m[106]&~m[107])|(m[7]&m[104]&m[105]&~m[106]&m[107])|(m[7]&m[104]&~m[105]&m[106]&m[107])|(m[7]&~m[104]&m[105]&m[106]&m[107])|(~m[7]&m[104]&m[105]&m[106]&m[107])|(m[7]&m[104]&m[105]&m[106]&m[107]))):InitCond[149];
    m[31] = run?((((m[7]&m[108]&~m[109]&~m[110]&~m[111])|(m[7]&~m[108]&m[109]&~m[110]&~m[111])|(~m[7]&m[108]&m[109]&~m[110]&~m[111])|(m[7]&~m[108]&~m[109]&m[110]&~m[111])|(~m[7]&m[108]&~m[109]&m[110]&~m[111])|(~m[7]&~m[108]&m[109]&m[110]&~m[111])|(m[7]&~m[108]&~m[109]&~m[110]&m[111])|(~m[7]&m[108]&~m[109]&~m[110]&m[111])|(~m[7]&~m[108]&m[109]&~m[110]&m[111])|(~m[7]&~m[108]&~m[109]&m[110]&m[111]))&BiasedRNG[79])|(((m[7]&m[108]&m[109]&~m[110]&~m[111])|(m[7]&m[108]&~m[109]&m[110]&~m[111])|(m[7]&~m[108]&m[109]&m[110]&~m[111])|(~m[7]&m[108]&m[109]&m[110]&~m[111])|(m[7]&m[108]&~m[109]&~m[110]&m[111])|(m[7]&~m[108]&m[109]&~m[110]&m[111])|(~m[7]&m[108]&m[109]&~m[110]&m[111])|(m[7]&~m[108]&~m[109]&m[110]&m[111])|(~m[7]&m[108]&~m[109]&m[110]&m[111])|(~m[7]&~m[108]&m[109]&m[110]&m[111]))&~BiasedRNG[79])|((m[7]&m[108]&m[109]&m[110]&~m[111])|(m[7]&m[108]&m[109]&~m[110]&m[111])|(m[7]&m[108]&~m[109]&m[110]&m[111])|(m[7]&~m[108]&m[109]&m[110]&m[111])|(~m[7]&m[108]&m[109]&m[110]&m[111])|(m[7]&m[108]&m[109]&m[110]&m[111]))):InitCond[150];
    m[32] = run?((((m[8]&m[112]&~m[113]&~m[114]&~m[115])|(m[8]&~m[112]&m[113]&~m[114]&~m[115])|(~m[8]&m[112]&m[113]&~m[114]&~m[115])|(m[8]&~m[112]&~m[113]&m[114]&~m[115])|(~m[8]&m[112]&~m[113]&m[114]&~m[115])|(~m[8]&~m[112]&m[113]&m[114]&~m[115])|(m[8]&~m[112]&~m[113]&~m[114]&m[115])|(~m[8]&m[112]&~m[113]&~m[114]&m[115])|(~m[8]&~m[112]&m[113]&~m[114]&m[115])|(~m[8]&~m[112]&~m[113]&m[114]&m[115]))&BiasedRNG[80])|(((m[8]&m[112]&m[113]&~m[114]&~m[115])|(m[8]&m[112]&~m[113]&m[114]&~m[115])|(m[8]&~m[112]&m[113]&m[114]&~m[115])|(~m[8]&m[112]&m[113]&m[114]&~m[115])|(m[8]&m[112]&~m[113]&~m[114]&m[115])|(m[8]&~m[112]&m[113]&~m[114]&m[115])|(~m[8]&m[112]&m[113]&~m[114]&m[115])|(m[8]&~m[112]&~m[113]&m[114]&m[115])|(~m[8]&m[112]&~m[113]&m[114]&m[115])|(~m[8]&~m[112]&m[113]&m[114]&m[115]))&~BiasedRNG[80])|((m[8]&m[112]&m[113]&m[114]&~m[115])|(m[8]&m[112]&m[113]&~m[114]&m[115])|(m[8]&m[112]&~m[113]&m[114]&m[115])|(m[8]&~m[112]&m[113]&m[114]&m[115])|(~m[8]&m[112]&m[113]&m[114]&m[115])|(m[8]&m[112]&m[113]&m[114]&m[115]))):InitCond[151];
    m[33] = run?((((m[8]&m[116]&~m[117]&~m[118]&~m[119])|(m[8]&~m[116]&m[117]&~m[118]&~m[119])|(~m[8]&m[116]&m[117]&~m[118]&~m[119])|(m[8]&~m[116]&~m[117]&m[118]&~m[119])|(~m[8]&m[116]&~m[117]&m[118]&~m[119])|(~m[8]&~m[116]&m[117]&m[118]&~m[119])|(m[8]&~m[116]&~m[117]&~m[118]&m[119])|(~m[8]&m[116]&~m[117]&~m[118]&m[119])|(~m[8]&~m[116]&m[117]&~m[118]&m[119])|(~m[8]&~m[116]&~m[117]&m[118]&m[119]))&BiasedRNG[81])|(((m[8]&m[116]&m[117]&~m[118]&~m[119])|(m[8]&m[116]&~m[117]&m[118]&~m[119])|(m[8]&~m[116]&m[117]&m[118]&~m[119])|(~m[8]&m[116]&m[117]&m[118]&~m[119])|(m[8]&m[116]&~m[117]&~m[118]&m[119])|(m[8]&~m[116]&m[117]&~m[118]&m[119])|(~m[8]&m[116]&m[117]&~m[118]&m[119])|(m[8]&~m[116]&~m[117]&m[118]&m[119])|(~m[8]&m[116]&~m[117]&m[118]&m[119])|(~m[8]&~m[116]&m[117]&m[118]&m[119]))&~BiasedRNG[81])|((m[8]&m[116]&m[117]&m[118]&~m[119])|(m[8]&m[116]&m[117]&~m[118]&m[119])|(m[8]&m[116]&~m[117]&m[118]&m[119])|(m[8]&~m[116]&m[117]&m[118]&m[119])|(~m[8]&m[116]&m[117]&m[118]&m[119])|(m[8]&m[116]&m[117]&m[118]&m[119]))):InitCond[152];
    m[34] = run?((((m[9]&m[120]&~m[121]&~m[122]&~m[123])|(m[9]&~m[120]&m[121]&~m[122]&~m[123])|(~m[9]&m[120]&m[121]&~m[122]&~m[123])|(m[9]&~m[120]&~m[121]&m[122]&~m[123])|(~m[9]&m[120]&~m[121]&m[122]&~m[123])|(~m[9]&~m[120]&m[121]&m[122]&~m[123])|(m[9]&~m[120]&~m[121]&~m[122]&m[123])|(~m[9]&m[120]&~m[121]&~m[122]&m[123])|(~m[9]&~m[120]&m[121]&~m[122]&m[123])|(~m[9]&~m[120]&~m[121]&m[122]&m[123]))&BiasedRNG[82])|(((m[9]&m[120]&m[121]&~m[122]&~m[123])|(m[9]&m[120]&~m[121]&m[122]&~m[123])|(m[9]&~m[120]&m[121]&m[122]&~m[123])|(~m[9]&m[120]&m[121]&m[122]&~m[123])|(m[9]&m[120]&~m[121]&~m[122]&m[123])|(m[9]&~m[120]&m[121]&~m[122]&m[123])|(~m[9]&m[120]&m[121]&~m[122]&m[123])|(m[9]&~m[120]&~m[121]&m[122]&m[123])|(~m[9]&m[120]&~m[121]&m[122]&m[123])|(~m[9]&~m[120]&m[121]&m[122]&m[123]))&~BiasedRNG[82])|((m[9]&m[120]&m[121]&m[122]&~m[123])|(m[9]&m[120]&m[121]&~m[122]&m[123])|(m[9]&m[120]&~m[121]&m[122]&m[123])|(m[9]&~m[120]&m[121]&m[122]&m[123])|(~m[9]&m[120]&m[121]&m[122]&m[123])|(m[9]&m[120]&m[121]&m[122]&m[123]))):InitCond[153];
    m[35] = run?((((m[9]&m[124]&~m[125]&~m[126]&~m[127])|(m[9]&~m[124]&m[125]&~m[126]&~m[127])|(~m[9]&m[124]&m[125]&~m[126]&~m[127])|(m[9]&~m[124]&~m[125]&m[126]&~m[127])|(~m[9]&m[124]&~m[125]&m[126]&~m[127])|(~m[9]&~m[124]&m[125]&m[126]&~m[127])|(m[9]&~m[124]&~m[125]&~m[126]&m[127])|(~m[9]&m[124]&~m[125]&~m[126]&m[127])|(~m[9]&~m[124]&m[125]&~m[126]&m[127])|(~m[9]&~m[124]&~m[125]&m[126]&m[127]))&BiasedRNG[83])|(((m[9]&m[124]&m[125]&~m[126]&~m[127])|(m[9]&m[124]&~m[125]&m[126]&~m[127])|(m[9]&~m[124]&m[125]&m[126]&~m[127])|(~m[9]&m[124]&m[125]&m[126]&~m[127])|(m[9]&m[124]&~m[125]&~m[126]&m[127])|(m[9]&~m[124]&m[125]&~m[126]&m[127])|(~m[9]&m[124]&m[125]&~m[126]&m[127])|(m[9]&~m[124]&~m[125]&m[126]&m[127])|(~m[9]&m[124]&~m[125]&m[126]&m[127])|(~m[9]&~m[124]&m[125]&m[126]&m[127]))&~BiasedRNG[83])|((m[9]&m[124]&m[125]&m[126]&~m[127])|(m[9]&m[124]&m[125]&~m[126]&m[127])|(m[9]&m[124]&~m[125]&m[126]&m[127])|(m[9]&~m[124]&m[125]&m[126]&m[127])|(~m[9]&m[124]&m[125]&m[126]&m[127])|(m[9]&m[124]&m[125]&m[126]&m[127]))):InitCond[154];
    m[36] = run?((((m[10]&m[128]&~m[129]&~m[130]&~m[131])|(m[10]&~m[128]&m[129]&~m[130]&~m[131])|(~m[10]&m[128]&m[129]&~m[130]&~m[131])|(m[10]&~m[128]&~m[129]&m[130]&~m[131])|(~m[10]&m[128]&~m[129]&m[130]&~m[131])|(~m[10]&~m[128]&m[129]&m[130]&~m[131])|(m[10]&~m[128]&~m[129]&~m[130]&m[131])|(~m[10]&m[128]&~m[129]&~m[130]&m[131])|(~m[10]&~m[128]&m[129]&~m[130]&m[131])|(~m[10]&~m[128]&~m[129]&m[130]&m[131]))&BiasedRNG[84])|(((m[10]&m[128]&m[129]&~m[130]&~m[131])|(m[10]&m[128]&~m[129]&m[130]&~m[131])|(m[10]&~m[128]&m[129]&m[130]&~m[131])|(~m[10]&m[128]&m[129]&m[130]&~m[131])|(m[10]&m[128]&~m[129]&~m[130]&m[131])|(m[10]&~m[128]&m[129]&~m[130]&m[131])|(~m[10]&m[128]&m[129]&~m[130]&m[131])|(m[10]&~m[128]&~m[129]&m[130]&m[131])|(~m[10]&m[128]&~m[129]&m[130]&m[131])|(~m[10]&~m[128]&m[129]&m[130]&m[131]))&~BiasedRNG[84])|((m[10]&m[128]&m[129]&m[130]&~m[131])|(m[10]&m[128]&m[129]&~m[130]&m[131])|(m[10]&m[128]&~m[129]&m[130]&m[131])|(m[10]&~m[128]&m[129]&m[130]&m[131])|(~m[10]&m[128]&m[129]&m[130]&m[131])|(m[10]&m[128]&m[129]&m[130]&m[131]))):InitCond[155];
    m[37] = run?((((m[10]&m[132]&~m[133]&~m[134]&~m[135])|(m[10]&~m[132]&m[133]&~m[134]&~m[135])|(~m[10]&m[132]&m[133]&~m[134]&~m[135])|(m[10]&~m[132]&~m[133]&m[134]&~m[135])|(~m[10]&m[132]&~m[133]&m[134]&~m[135])|(~m[10]&~m[132]&m[133]&m[134]&~m[135])|(m[10]&~m[132]&~m[133]&~m[134]&m[135])|(~m[10]&m[132]&~m[133]&~m[134]&m[135])|(~m[10]&~m[132]&m[133]&~m[134]&m[135])|(~m[10]&~m[132]&~m[133]&m[134]&m[135]))&BiasedRNG[85])|(((m[10]&m[132]&m[133]&~m[134]&~m[135])|(m[10]&m[132]&~m[133]&m[134]&~m[135])|(m[10]&~m[132]&m[133]&m[134]&~m[135])|(~m[10]&m[132]&m[133]&m[134]&~m[135])|(m[10]&m[132]&~m[133]&~m[134]&m[135])|(m[10]&~m[132]&m[133]&~m[134]&m[135])|(~m[10]&m[132]&m[133]&~m[134]&m[135])|(m[10]&~m[132]&~m[133]&m[134]&m[135])|(~m[10]&m[132]&~m[133]&m[134]&m[135])|(~m[10]&~m[132]&m[133]&m[134]&m[135]))&~BiasedRNG[85])|((m[10]&m[132]&m[133]&m[134]&~m[135])|(m[10]&m[132]&m[133]&~m[134]&m[135])|(m[10]&m[132]&~m[133]&m[134]&m[135])|(m[10]&~m[132]&m[133]&m[134]&m[135])|(~m[10]&m[132]&m[133]&m[134]&m[135])|(m[10]&m[132]&m[133]&m[134]&m[135]))):InitCond[156];
    m[38] = run?((((m[11]&m[136]&~m[137]&~m[138]&~m[139])|(m[11]&~m[136]&m[137]&~m[138]&~m[139])|(~m[11]&m[136]&m[137]&~m[138]&~m[139])|(m[11]&~m[136]&~m[137]&m[138]&~m[139])|(~m[11]&m[136]&~m[137]&m[138]&~m[139])|(~m[11]&~m[136]&m[137]&m[138]&~m[139])|(m[11]&~m[136]&~m[137]&~m[138]&m[139])|(~m[11]&m[136]&~m[137]&~m[138]&m[139])|(~m[11]&~m[136]&m[137]&~m[138]&m[139])|(~m[11]&~m[136]&~m[137]&m[138]&m[139]))&BiasedRNG[86])|(((m[11]&m[136]&m[137]&~m[138]&~m[139])|(m[11]&m[136]&~m[137]&m[138]&~m[139])|(m[11]&~m[136]&m[137]&m[138]&~m[139])|(~m[11]&m[136]&m[137]&m[138]&~m[139])|(m[11]&m[136]&~m[137]&~m[138]&m[139])|(m[11]&~m[136]&m[137]&~m[138]&m[139])|(~m[11]&m[136]&m[137]&~m[138]&m[139])|(m[11]&~m[136]&~m[137]&m[138]&m[139])|(~m[11]&m[136]&~m[137]&m[138]&m[139])|(~m[11]&~m[136]&m[137]&m[138]&m[139]))&~BiasedRNG[86])|((m[11]&m[136]&m[137]&m[138]&~m[139])|(m[11]&m[136]&m[137]&~m[138]&m[139])|(m[11]&m[136]&~m[137]&m[138]&m[139])|(m[11]&~m[136]&m[137]&m[138]&m[139])|(~m[11]&m[136]&m[137]&m[138]&m[139])|(m[11]&m[136]&m[137]&m[138]&m[139]))):InitCond[157];
    m[39] = run?((((m[11]&m[140]&~m[141]&~m[142]&~m[143])|(m[11]&~m[140]&m[141]&~m[142]&~m[143])|(~m[11]&m[140]&m[141]&~m[142]&~m[143])|(m[11]&~m[140]&~m[141]&m[142]&~m[143])|(~m[11]&m[140]&~m[141]&m[142]&~m[143])|(~m[11]&~m[140]&m[141]&m[142]&~m[143])|(m[11]&~m[140]&~m[141]&~m[142]&m[143])|(~m[11]&m[140]&~m[141]&~m[142]&m[143])|(~m[11]&~m[140]&m[141]&~m[142]&m[143])|(~m[11]&~m[140]&~m[141]&m[142]&m[143]))&BiasedRNG[87])|(((m[11]&m[140]&m[141]&~m[142]&~m[143])|(m[11]&m[140]&~m[141]&m[142]&~m[143])|(m[11]&~m[140]&m[141]&m[142]&~m[143])|(~m[11]&m[140]&m[141]&m[142]&~m[143])|(m[11]&m[140]&~m[141]&~m[142]&m[143])|(m[11]&~m[140]&m[141]&~m[142]&m[143])|(~m[11]&m[140]&m[141]&~m[142]&m[143])|(m[11]&~m[140]&~m[141]&m[142]&m[143])|(~m[11]&m[140]&~m[141]&m[142]&m[143])|(~m[11]&~m[140]&m[141]&m[142]&m[143]))&~BiasedRNG[87])|((m[11]&m[140]&m[141]&m[142]&~m[143])|(m[11]&m[140]&m[141]&~m[142]&m[143])|(m[11]&m[140]&~m[141]&m[142]&m[143])|(m[11]&~m[140]&m[141]&m[142]&m[143])|(~m[11]&m[140]&m[141]&m[142]&m[143])|(m[11]&m[140]&m[141]&m[142]&m[143]))):InitCond[158];
    m[40] = run?((((m[12]&m[144]&~m[145]&~m[146]&~m[147])|(m[12]&~m[144]&m[145]&~m[146]&~m[147])|(~m[12]&m[144]&m[145]&~m[146]&~m[147])|(m[12]&~m[144]&~m[145]&m[146]&~m[147])|(~m[12]&m[144]&~m[145]&m[146]&~m[147])|(~m[12]&~m[144]&m[145]&m[146]&~m[147])|(m[12]&~m[144]&~m[145]&~m[146]&m[147])|(~m[12]&m[144]&~m[145]&~m[146]&m[147])|(~m[12]&~m[144]&m[145]&~m[146]&m[147])|(~m[12]&~m[144]&~m[145]&m[146]&m[147]))&BiasedRNG[88])|(((m[12]&m[144]&m[145]&~m[146]&~m[147])|(m[12]&m[144]&~m[145]&m[146]&~m[147])|(m[12]&~m[144]&m[145]&m[146]&~m[147])|(~m[12]&m[144]&m[145]&m[146]&~m[147])|(m[12]&m[144]&~m[145]&~m[146]&m[147])|(m[12]&~m[144]&m[145]&~m[146]&m[147])|(~m[12]&m[144]&m[145]&~m[146]&m[147])|(m[12]&~m[144]&~m[145]&m[146]&m[147])|(~m[12]&m[144]&~m[145]&m[146]&m[147])|(~m[12]&~m[144]&m[145]&m[146]&m[147]))&~BiasedRNG[88])|((m[12]&m[144]&m[145]&m[146]&~m[147])|(m[12]&m[144]&m[145]&~m[146]&m[147])|(m[12]&m[144]&~m[145]&m[146]&m[147])|(m[12]&~m[144]&m[145]&m[146]&m[147])|(~m[12]&m[144]&m[145]&m[146]&m[147])|(m[12]&m[144]&m[145]&m[146]&m[147]))):InitCond[159];
    m[41] = run?((((m[12]&m[148]&~m[149]&~m[150]&~m[151])|(m[12]&~m[148]&m[149]&~m[150]&~m[151])|(~m[12]&m[148]&m[149]&~m[150]&~m[151])|(m[12]&~m[148]&~m[149]&m[150]&~m[151])|(~m[12]&m[148]&~m[149]&m[150]&~m[151])|(~m[12]&~m[148]&m[149]&m[150]&~m[151])|(m[12]&~m[148]&~m[149]&~m[150]&m[151])|(~m[12]&m[148]&~m[149]&~m[150]&m[151])|(~m[12]&~m[148]&m[149]&~m[150]&m[151])|(~m[12]&~m[148]&~m[149]&m[150]&m[151]))&BiasedRNG[89])|(((m[12]&m[148]&m[149]&~m[150]&~m[151])|(m[12]&m[148]&~m[149]&m[150]&~m[151])|(m[12]&~m[148]&m[149]&m[150]&~m[151])|(~m[12]&m[148]&m[149]&m[150]&~m[151])|(m[12]&m[148]&~m[149]&~m[150]&m[151])|(m[12]&~m[148]&m[149]&~m[150]&m[151])|(~m[12]&m[148]&m[149]&~m[150]&m[151])|(m[12]&~m[148]&~m[149]&m[150]&m[151])|(~m[12]&m[148]&~m[149]&m[150]&m[151])|(~m[12]&~m[148]&m[149]&m[150]&m[151]))&~BiasedRNG[89])|((m[12]&m[148]&m[149]&m[150]&~m[151])|(m[12]&m[148]&m[149]&~m[150]&m[151])|(m[12]&m[148]&~m[149]&m[150]&m[151])|(m[12]&~m[148]&m[149]&m[150]&m[151])|(~m[12]&m[148]&m[149]&m[150]&m[151])|(m[12]&m[148]&m[149]&m[150]&m[151]))):InitCond[160];
    m[42] = run?((((m[13]&m[152]&~m[153]&~m[154]&~m[155])|(m[13]&~m[152]&m[153]&~m[154]&~m[155])|(~m[13]&m[152]&m[153]&~m[154]&~m[155])|(m[13]&~m[152]&~m[153]&m[154]&~m[155])|(~m[13]&m[152]&~m[153]&m[154]&~m[155])|(~m[13]&~m[152]&m[153]&m[154]&~m[155])|(m[13]&~m[152]&~m[153]&~m[154]&m[155])|(~m[13]&m[152]&~m[153]&~m[154]&m[155])|(~m[13]&~m[152]&m[153]&~m[154]&m[155])|(~m[13]&~m[152]&~m[153]&m[154]&m[155]))&BiasedRNG[90])|(((m[13]&m[152]&m[153]&~m[154]&~m[155])|(m[13]&m[152]&~m[153]&m[154]&~m[155])|(m[13]&~m[152]&m[153]&m[154]&~m[155])|(~m[13]&m[152]&m[153]&m[154]&~m[155])|(m[13]&m[152]&~m[153]&~m[154]&m[155])|(m[13]&~m[152]&m[153]&~m[154]&m[155])|(~m[13]&m[152]&m[153]&~m[154]&m[155])|(m[13]&~m[152]&~m[153]&m[154]&m[155])|(~m[13]&m[152]&~m[153]&m[154]&m[155])|(~m[13]&~m[152]&m[153]&m[154]&m[155]))&~BiasedRNG[90])|((m[13]&m[152]&m[153]&m[154]&~m[155])|(m[13]&m[152]&m[153]&~m[154]&m[155])|(m[13]&m[152]&~m[153]&m[154]&m[155])|(m[13]&~m[152]&m[153]&m[154]&m[155])|(~m[13]&m[152]&m[153]&m[154]&m[155])|(m[13]&m[152]&m[153]&m[154]&m[155]))):InitCond[161];
    m[43] = run?((((m[13]&m[156]&~m[157]&~m[158]&~m[159])|(m[13]&~m[156]&m[157]&~m[158]&~m[159])|(~m[13]&m[156]&m[157]&~m[158]&~m[159])|(m[13]&~m[156]&~m[157]&m[158]&~m[159])|(~m[13]&m[156]&~m[157]&m[158]&~m[159])|(~m[13]&~m[156]&m[157]&m[158]&~m[159])|(m[13]&~m[156]&~m[157]&~m[158]&m[159])|(~m[13]&m[156]&~m[157]&~m[158]&m[159])|(~m[13]&~m[156]&m[157]&~m[158]&m[159])|(~m[13]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[91])|(((m[13]&m[156]&m[157]&~m[158]&~m[159])|(m[13]&m[156]&~m[157]&m[158]&~m[159])|(m[13]&~m[156]&m[157]&m[158]&~m[159])|(~m[13]&m[156]&m[157]&m[158]&~m[159])|(m[13]&m[156]&~m[157]&~m[158]&m[159])|(m[13]&~m[156]&m[157]&~m[158]&m[159])|(~m[13]&m[156]&m[157]&~m[158]&m[159])|(m[13]&~m[156]&~m[157]&m[158]&m[159])|(~m[13]&m[156]&~m[157]&m[158]&m[159])|(~m[13]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[91])|((m[13]&m[156]&m[157]&m[158]&~m[159])|(m[13]&m[156]&m[157]&~m[158]&m[159])|(m[13]&m[156]&~m[157]&m[158]&m[159])|(m[13]&~m[156]&m[157]&m[158]&m[159])|(~m[13]&m[156]&m[157]&m[158]&m[159])|(m[13]&m[156]&m[157]&m[158]&m[159]))):InitCond[162];
    m[44] = run?((((m[14]&m[160]&~m[161]&~m[162]&~m[163])|(m[14]&~m[160]&m[161]&~m[162]&~m[163])|(~m[14]&m[160]&m[161]&~m[162]&~m[163])|(m[14]&~m[160]&~m[161]&m[162]&~m[163])|(~m[14]&m[160]&~m[161]&m[162]&~m[163])|(~m[14]&~m[160]&m[161]&m[162]&~m[163])|(m[14]&~m[160]&~m[161]&~m[162]&m[163])|(~m[14]&m[160]&~m[161]&~m[162]&m[163])|(~m[14]&~m[160]&m[161]&~m[162]&m[163])|(~m[14]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[92])|(((m[14]&m[160]&m[161]&~m[162]&~m[163])|(m[14]&m[160]&~m[161]&m[162]&~m[163])|(m[14]&~m[160]&m[161]&m[162]&~m[163])|(~m[14]&m[160]&m[161]&m[162]&~m[163])|(m[14]&m[160]&~m[161]&~m[162]&m[163])|(m[14]&~m[160]&m[161]&~m[162]&m[163])|(~m[14]&m[160]&m[161]&~m[162]&m[163])|(m[14]&~m[160]&~m[161]&m[162]&m[163])|(~m[14]&m[160]&~m[161]&m[162]&m[163])|(~m[14]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[92])|((m[14]&m[160]&m[161]&m[162]&~m[163])|(m[14]&m[160]&m[161]&~m[162]&m[163])|(m[14]&m[160]&~m[161]&m[162]&m[163])|(m[14]&~m[160]&m[161]&m[162]&m[163])|(~m[14]&m[160]&m[161]&m[162]&m[163])|(m[14]&m[160]&m[161]&m[162]&m[163]))):InitCond[163];
    m[45] = run?((((m[14]&m[164]&~m[165]&~m[166]&~m[167])|(m[14]&~m[164]&m[165]&~m[166]&~m[167])|(~m[14]&m[164]&m[165]&~m[166]&~m[167])|(m[14]&~m[164]&~m[165]&m[166]&~m[167])|(~m[14]&m[164]&~m[165]&m[166]&~m[167])|(~m[14]&~m[164]&m[165]&m[166]&~m[167])|(m[14]&~m[164]&~m[165]&~m[166]&m[167])|(~m[14]&m[164]&~m[165]&~m[166]&m[167])|(~m[14]&~m[164]&m[165]&~m[166]&m[167])|(~m[14]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[93])|(((m[14]&m[164]&m[165]&~m[166]&~m[167])|(m[14]&m[164]&~m[165]&m[166]&~m[167])|(m[14]&~m[164]&m[165]&m[166]&~m[167])|(~m[14]&m[164]&m[165]&m[166]&~m[167])|(m[14]&m[164]&~m[165]&~m[166]&m[167])|(m[14]&~m[164]&m[165]&~m[166]&m[167])|(~m[14]&m[164]&m[165]&~m[166]&m[167])|(m[14]&~m[164]&~m[165]&m[166]&m[167])|(~m[14]&m[164]&~m[165]&m[166]&m[167])|(~m[14]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[93])|((m[14]&m[164]&m[165]&m[166]&~m[167])|(m[14]&m[164]&m[165]&~m[166]&m[167])|(m[14]&m[164]&~m[165]&m[166]&m[167])|(m[14]&~m[164]&m[165]&m[166]&m[167])|(~m[14]&m[164]&m[165]&m[166]&m[167])|(m[14]&m[164]&m[165]&m[166]&m[167]))):InitCond[164];
    m[46] = run?((((m[15]&m[168]&~m[169]&~m[170]&~m[171])|(m[15]&~m[168]&m[169]&~m[170]&~m[171])|(~m[15]&m[168]&m[169]&~m[170]&~m[171])|(m[15]&~m[168]&~m[169]&m[170]&~m[171])|(~m[15]&m[168]&~m[169]&m[170]&~m[171])|(~m[15]&~m[168]&m[169]&m[170]&~m[171])|(m[15]&~m[168]&~m[169]&~m[170]&m[171])|(~m[15]&m[168]&~m[169]&~m[170]&m[171])|(~m[15]&~m[168]&m[169]&~m[170]&m[171])|(~m[15]&~m[168]&~m[169]&m[170]&m[171]))&BiasedRNG[94])|(((m[15]&m[168]&m[169]&~m[170]&~m[171])|(m[15]&m[168]&~m[169]&m[170]&~m[171])|(m[15]&~m[168]&m[169]&m[170]&~m[171])|(~m[15]&m[168]&m[169]&m[170]&~m[171])|(m[15]&m[168]&~m[169]&~m[170]&m[171])|(m[15]&~m[168]&m[169]&~m[170]&m[171])|(~m[15]&m[168]&m[169]&~m[170]&m[171])|(m[15]&~m[168]&~m[169]&m[170]&m[171])|(~m[15]&m[168]&~m[169]&m[170]&m[171])|(~m[15]&~m[168]&m[169]&m[170]&m[171]))&~BiasedRNG[94])|((m[15]&m[168]&m[169]&m[170]&~m[171])|(m[15]&m[168]&m[169]&~m[170]&m[171])|(m[15]&m[168]&~m[169]&m[170]&m[171])|(m[15]&~m[168]&m[169]&m[170]&m[171])|(~m[15]&m[168]&m[169]&m[170]&m[171])|(m[15]&m[168]&m[169]&m[170]&m[171]))):InitCond[165];
    m[47] = run?((((m[15]&m[172]&~m[173]&~m[174]&~m[175])|(m[15]&~m[172]&m[173]&~m[174]&~m[175])|(~m[15]&m[172]&m[173]&~m[174]&~m[175])|(m[15]&~m[172]&~m[173]&m[174]&~m[175])|(~m[15]&m[172]&~m[173]&m[174]&~m[175])|(~m[15]&~m[172]&m[173]&m[174]&~m[175])|(m[15]&~m[172]&~m[173]&~m[174]&m[175])|(~m[15]&m[172]&~m[173]&~m[174]&m[175])|(~m[15]&~m[172]&m[173]&~m[174]&m[175])|(~m[15]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[95])|(((m[15]&m[172]&m[173]&~m[174]&~m[175])|(m[15]&m[172]&~m[173]&m[174]&~m[175])|(m[15]&~m[172]&m[173]&m[174]&~m[175])|(~m[15]&m[172]&m[173]&m[174]&~m[175])|(m[15]&m[172]&~m[173]&~m[174]&m[175])|(m[15]&~m[172]&m[173]&~m[174]&m[175])|(~m[15]&m[172]&m[173]&~m[174]&m[175])|(m[15]&~m[172]&~m[173]&m[174]&m[175])|(~m[15]&m[172]&~m[173]&m[174]&m[175])|(~m[15]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[95])|((m[15]&m[172]&m[173]&m[174]&~m[175])|(m[15]&m[172]&m[173]&~m[174]&m[175])|(m[15]&m[172]&~m[173]&m[174]&m[175])|(m[15]&~m[172]&m[173]&m[174]&m[175])|(~m[15]&m[172]&m[173]&m[174]&m[175])|(m[15]&m[172]&m[173]&m[174]&m[175]))):InitCond[166];
    m[177] = run?((((m[56]&~m[113]&m[240])|(~m[56]&m[113]&m[240]))&BiasedRNG[96])|(((m[56]&m[113]&~m[240]))&~BiasedRNG[96])|((m[56]&m[113]&m[240]))):InitCond[167];
    m[178] = run?((((m[64]&~m[114]&m[245])|(~m[64]&m[114]&m[245]))&BiasedRNG[97])|(((m[64]&m[114]&~m[245]))&~BiasedRNG[97])|((m[64]&m[114]&m[245]))):InitCond[168];
    m[179] = run?((((m[72]&~m[115]&m[255])|(~m[72]&m[115]&m[255]))&BiasedRNG[98])|(((m[72]&m[115]&~m[255]))&~BiasedRNG[98])|((m[72]&m[115]&m[255]))):InitCond[169];
    m[180] = run?((((m[80]&~m[116]&m[270])|(~m[80]&m[116]&m[270]))&BiasedRNG[99])|(((m[80]&m[116]&~m[270]))&~BiasedRNG[99])|((m[80]&m[116]&m[270]))):InitCond[170];
    m[181] = run?((((m[88]&~m[117]&m[290])|(~m[88]&m[117]&m[290]))&BiasedRNG[100])|(((m[88]&m[117]&~m[290]))&~BiasedRNG[100])|((m[88]&m[117]&m[290]))):InitCond[171];
    m[182] = run?((((m[96]&~m[118]&m[315])|(~m[96]&m[118]&m[315]))&BiasedRNG[101])|(((m[96]&m[118]&~m[315]))&~BiasedRNG[101])|((m[96]&m[118]&m[315]))):InitCond[172];
    m[183] = run?((((m[104]&~m[119]&m[345])|(~m[104]&m[119]&m[345]))&BiasedRNG[102])|(((m[104]&m[119]&~m[345]))&~BiasedRNG[102])|((m[104]&m[119]&m[345]))):InitCond[173];
    m[184] = run?((((m[49]&~m[120]&m[241])|(~m[49]&m[120]&m[241]))&BiasedRNG[103])|(((m[49]&m[120]&~m[241]))&~BiasedRNG[103])|((m[49]&m[120]&m[241]))):InitCond[174];
    m[185] = run?((((m[57]&~m[121]&m[246])|(~m[57]&m[121]&m[246]))&BiasedRNG[104])|(((m[57]&m[121]&~m[246]))&~BiasedRNG[104])|((m[57]&m[121]&m[246]))):InitCond[175];
    m[186] = run?((((m[65]&~m[122]&m[256])|(~m[65]&m[122]&m[256]))&BiasedRNG[105])|(((m[65]&m[122]&~m[256]))&~BiasedRNG[105])|((m[65]&m[122]&m[256]))):InitCond[176];
    m[187] = run?((((m[73]&~m[123]&m[271])|(~m[73]&m[123]&m[271]))&BiasedRNG[106])|(((m[73]&m[123]&~m[271]))&~BiasedRNG[106])|((m[73]&m[123]&m[271]))):InitCond[177];
    m[188] = run?((((m[81]&~m[124]&m[291])|(~m[81]&m[124]&m[291]))&BiasedRNG[107])|(((m[81]&m[124]&~m[291]))&~BiasedRNG[107])|((m[81]&m[124]&m[291]))):InitCond[178];
    m[189] = run?((((m[89]&~m[125]&m[316])|(~m[89]&m[125]&m[316]))&BiasedRNG[108])|(((m[89]&m[125]&~m[316]))&~BiasedRNG[108])|((m[89]&m[125]&m[316]))):InitCond[179];
    m[190] = run?((((m[97]&~m[126]&m[346])|(~m[97]&m[126]&m[346]))&BiasedRNG[109])|(((m[97]&m[126]&~m[346]))&~BiasedRNG[109])|((m[97]&m[126]&m[346]))):InitCond[180];
    m[191] = run?((((m[105]&~m[127]&m[381])|(~m[105]&m[127]&m[381]))&BiasedRNG[110])|(((m[105]&m[127]&~m[381]))&~BiasedRNG[110])|((m[105]&m[127]&m[381]))):InitCond[181];
    m[192] = run?((((m[50]&~m[128]&m[251])|(~m[50]&m[128]&m[251]))&BiasedRNG[111])|(((m[50]&m[128]&~m[251]))&~BiasedRNG[111])|((m[50]&m[128]&m[251]))):InitCond[182];
    m[193] = run?((((m[58]&~m[129]&m[261])|(~m[58]&m[129]&m[261]))&BiasedRNG[112])|(((m[58]&m[129]&~m[261]))&~BiasedRNG[112])|((m[58]&m[129]&m[261]))):InitCond[183];
    m[194] = run?((((m[66]&~m[130]&m[276])|(~m[66]&m[130]&m[276]))&BiasedRNG[113])|(((m[66]&m[130]&~m[276]))&~BiasedRNG[113])|((m[66]&m[130]&m[276]))):InitCond[184];
    m[195] = run?((((m[74]&~m[131]&m[296])|(~m[74]&m[131]&m[296]))&BiasedRNG[114])|(((m[74]&m[131]&~m[296]))&~BiasedRNG[114])|((m[74]&m[131]&m[296]))):InitCond[185];
    m[196] = run?((((m[82]&~m[132]&m[321])|(~m[82]&m[132]&m[321]))&BiasedRNG[115])|(((m[82]&m[132]&~m[321]))&~BiasedRNG[115])|((m[82]&m[132]&m[321]))):InitCond[186];
    m[197] = run?((((m[90]&~m[133]&m[351])|(~m[90]&m[133]&m[351]))&BiasedRNG[116])|(((m[90]&m[133]&~m[351]))&~BiasedRNG[116])|((m[90]&m[133]&m[351]))):InitCond[187];
    m[198] = run?((((m[98]&~m[134]&m[386])|(~m[98]&m[134]&m[386]))&BiasedRNG[117])|(((m[98]&m[134]&~m[386]))&~BiasedRNG[117])|((m[98]&m[134]&m[386]))):InitCond[188];
    m[199] = run?((((m[106]&~m[135]&m[416])|(~m[106]&m[135]&m[416]))&BiasedRNG[118])|(((m[106]&m[135]&~m[416]))&~BiasedRNG[118])|((m[106]&m[135]&m[416]))):InitCond[189];
    m[200] = run?((((m[51]&~m[136]&m[266])|(~m[51]&m[136]&m[266]))&BiasedRNG[119])|(((m[51]&m[136]&~m[266]))&~BiasedRNG[119])|((m[51]&m[136]&m[266]))):InitCond[190];
    m[201] = run?((((m[59]&~m[137]&m[281])|(~m[59]&m[137]&m[281]))&BiasedRNG[120])|(((m[59]&m[137]&~m[281]))&~BiasedRNG[120])|((m[59]&m[137]&m[281]))):InitCond[191];
    m[202] = run?((((m[67]&~m[138]&m[301])|(~m[67]&m[138]&m[301]))&BiasedRNG[121])|(((m[67]&m[138]&~m[301]))&~BiasedRNG[121])|((m[67]&m[138]&m[301]))):InitCond[192];
    m[203] = run?((((m[75]&~m[139]&m[326])|(~m[75]&m[139]&m[326]))&BiasedRNG[122])|(((m[75]&m[139]&~m[326]))&~BiasedRNG[122])|((m[75]&m[139]&m[326]))):InitCond[193];
    m[204] = run?((((m[83]&~m[140]&m[356])|(~m[83]&m[140]&m[356]))&BiasedRNG[123])|(((m[83]&m[140]&~m[356]))&~BiasedRNG[123])|((m[83]&m[140]&m[356]))):InitCond[194];
    m[205] = run?((((m[91]&~m[141]&m[391])|(~m[91]&m[141]&m[391]))&BiasedRNG[124])|(((m[91]&m[141]&~m[391]))&~BiasedRNG[124])|((m[91]&m[141]&m[391]))):InitCond[195];
    m[206] = run?((((m[99]&~m[142]&m[421])|(~m[99]&m[142]&m[421]))&BiasedRNG[125])|(((m[99]&m[142]&~m[421]))&~BiasedRNG[125])|((m[99]&m[142]&m[421]))):InitCond[196];
    m[207] = run?((((m[107]&~m[143]&m[446])|(~m[107]&m[143]&m[446]))&BiasedRNG[126])|(((m[107]&m[143]&~m[446]))&~BiasedRNG[126])|((m[107]&m[143]&m[446]))):InitCond[197];
    m[208] = run?((((m[52]&~m[144]&m[286])|(~m[52]&m[144]&m[286]))&BiasedRNG[127])|(((m[52]&m[144]&~m[286]))&~BiasedRNG[127])|((m[52]&m[144]&m[286]))):InitCond[198];
    m[209] = run?((((m[60]&~m[145]&m[306])|(~m[60]&m[145]&m[306]))&BiasedRNG[128])|(((m[60]&m[145]&~m[306]))&~BiasedRNG[128])|((m[60]&m[145]&m[306]))):InitCond[199];
    m[210] = run?((((m[68]&~m[146]&m[331])|(~m[68]&m[146]&m[331]))&BiasedRNG[129])|(((m[68]&m[146]&~m[331]))&~BiasedRNG[129])|((m[68]&m[146]&m[331]))):InitCond[200];
    m[211] = run?((((m[76]&~m[147]&m[361])|(~m[76]&m[147]&m[361]))&BiasedRNG[130])|(((m[76]&m[147]&~m[361]))&~BiasedRNG[130])|((m[76]&m[147]&m[361]))):InitCond[201];
    m[212] = run?((((m[84]&~m[148]&m[396])|(~m[84]&m[148]&m[396]))&BiasedRNG[131])|(((m[84]&m[148]&~m[396]))&~BiasedRNG[131])|((m[84]&m[148]&m[396]))):InitCond[202];
    m[213] = run?((((m[92]&~m[149]&m[426])|(~m[92]&m[149]&m[426]))&BiasedRNG[132])|(((m[92]&m[149]&~m[426]))&~BiasedRNG[132])|((m[92]&m[149]&m[426]))):InitCond[203];
    m[214] = run?((((m[100]&~m[150]&m[451])|(~m[100]&m[150]&m[451]))&BiasedRNG[133])|(((m[100]&m[150]&~m[451]))&~BiasedRNG[133])|((m[100]&m[150]&m[451]))):InitCond[204];
    m[215] = run?((((m[108]&~m[151]&m[471])|(~m[108]&m[151]&m[471]))&BiasedRNG[134])|(((m[108]&m[151]&~m[471]))&~BiasedRNG[134])|((m[108]&m[151]&m[471]))):InitCond[205];
    m[216] = run?((((m[53]&~m[152]&m[311])|(~m[53]&m[152]&m[311]))&BiasedRNG[135])|(((m[53]&m[152]&~m[311]))&~BiasedRNG[135])|((m[53]&m[152]&m[311]))):InitCond[206];
    m[217] = run?((((m[61]&~m[153]&m[336])|(~m[61]&m[153]&m[336]))&BiasedRNG[136])|(((m[61]&m[153]&~m[336]))&~BiasedRNG[136])|((m[61]&m[153]&m[336]))):InitCond[207];
    m[218] = run?((((m[69]&~m[154]&m[366])|(~m[69]&m[154]&m[366]))&BiasedRNG[137])|(((m[69]&m[154]&~m[366]))&~BiasedRNG[137])|((m[69]&m[154]&m[366]))):InitCond[208];
    m[219] = run?((((m[77]&~m[155]&m[401])|(~m[77]&m[155]&m[401]))&BiasedRNG[138])|(((m[77]&m[155]&~m[401]))&~BiasedRNG[138])|((m[77]&m[155]&m[401]))):InitCond[209];
    m[220] = run?((((m[85]&~m[156]&m[431])|(~m[85]&m[156]&m[431]))&BiasedRNG[139])|(((m[85]&m[156]&~m[431]))&~BiasedRNG[139])|((m[85]&m[156]&m[431]))):InitCond[210];
    m[221] = run?((((m[93]&~m[157]&m[456])|(~m[93]&m[157]&m[456]))&BiasedRNG[140])|(((m[93]&m[157]&~m[456]))&~BiasedRNG[140])|((m[93]&m[157]&m[456]))):InitCond[211];
    m[222] = run?((((m[101]&~m[158]&m[476])|(~m[101]&m[158]&m[476]))&BiasedRNG[141])|(((m[101]&m[158]&~m[476]))&~BiasedRNG[141])|((m[101]&m[158]&m[476]))):InitCond[212];
    m[223] = run?((((m[109]&~m[159]&m[491])|(~m[109]&m[159]&m[491]))&BiasedRNG[142])|(((m[109]&m[159]&~m[491]))&~BiasedRNG[142])|((m[109]&m[159]&m[491]))):InitCond[213];
    m[224] = run?((((m[54]&~m[160]&m[341])|(~m[54]&m[160]&m[341]))&BiasedRNG[143])|(((m[54]&m[160]&~m[341]))&~BiasedRNG[143])|((m[54]&m[160]&m[341]))):InitCond[214];
    m[225] = run?((((m[62]&~m[161]&m[371])|(~m[62]&m[161]&m[371]))&BiasedRNG[144])|(((m[62]&m[161]&~m[371]))&~BiasedRNG[144])|((m[62]&m[161]&m[371]))):InitCond[215];
    m[226] = run?((((m[70]&~m[162]&m[406])|(~m[70]&m[162]&m[406]))&BiasedRNG[145])|(((m[70]&m[162]&~m[406]))&~BiasedRNG[145])|((m[70]&m[162]&m[406]))):InitCond[216];
    m[227] = run?((((m[78]&~m[163]&m[436])|(~m[78]&m[163]&m[436]))&BiasedRNG[146])|(((m[78]&m[163]&~m[436]))&~BiasedRNG[146])|((m[78]&m[163]&m[436]))):InitCond[217];
    m[228] = run?((((m[86]&~m[164]&m[461])|(~m[86]&m[164]&m[461]))&BiasedRNG[147])|(((m[86]&m[164]&~m[461]))&~BiasedRNG[147])|((m[86]&m[164]&m[461]))):InitCond[218];
    m[229] = run?((((m[94]&~m[165]&m[481])|(~m[94]&m[165]&m[481]))&BiasedRNG[148])|(((m[94]&m[165]&~m[481]))&~BiasedRNG[148])|((m[94]&m[165]&m[481]))):InitCond[219];
    m[230] = run?((((m[102]&~m[166]&m[496])|(~m[102]&m[166]&m[496]))&BiasedRNG[149])|(((m[102]&m[166]&~m[496]))&~BiasedRNG[149])|((m[102]&m[166]&m[496]))):InitCond[220];
    m[231] = run?((((m[110]&~m[167]&m[506])|(~m[110]&m[167]&m[506]))&BiasedRNG[150])|(((m[110]&m[167]&~m[506]))&~BiasedRNG[150])|((m[110]&m[167]&m[506]))):InitCond[221];
    m[232] = run?((((m[55]&~m[168]&m[376])|(~m[55]&m[168]&m[376]))&BiasedRNG[151])|(((m[55]&m[168]&~m[376]))&~BiasedRNG[151])|((m[55]&m[168]&m[376]))):InitCond[222];
    m[233] = run?((((m[63]&~m[169]&m[411])|(~m[63]&m[169]&m[411]))&BiasedRNG[152])|(((m[63]&m[169]&~m[411]))&~BiasedRNG[152])|((m[63]&m[169]&m[411]))):InitCond[223];
    m[234] = run?((((m[71]&~m[170]&m[441])|(~m[71]&m[170]&m[441]))&BiasedRNG[153])|(((m[71]&m[170]&~m[441]))&~BiasedRNG[153])|((m[71]&m[170]&m[441]))):InitCond[224];
    m[235] = run?((((m[79]&~m[171]&m[466])|(~m[79]&m[171]&m[466]))&BiasedRNG[154])|(((m[79]&m[171]&~m[466]))&~BiasedRNG[154])|((m[79]&m[171]&m[466]))):InitCond[225];
    m[236] = run?((((m[87]&~m[172]&m[486])|(~m[87]&m[172]&m[486]))&BiasedRNG[155])|(((m[87]&m[172]&~m[486]))&~BiasedRNG[155])|((m[87]&m[172]&m[486]))):InitCond[226];
    m[237] = run?((((m[95]&~m[173]&m[501])|(~m[95]&m[173]&m[501]))&BiasedRNG[156])|(((m[95]&m[173]&~m[501]))&~BiasedRNG[156])|((m[95]&m[173]&m[501]))):InitCond[227];
    m[238] = run?((((m[103]&~m[174]&m[511])|(~m[103]&m[174]&m[511]))&BiasedRNG[157])|(((m[103]&m[174]&~m[511]))&~BiasedRNG[157])|((m[103]&m[174]&m[511]))):InitCond[228];
    m[239] = run?((((m[111]&~m[175]&m[516])|(~m[111]&m[175]&m[516]))&BiasedRNG[158])|(((m[111]&m[175]&~m[516]))&~BiasedRNG[158])|((m[111]&m[175]&m[516]))):InitCond[229];
    m[247] = run?((((m[244]&~m[245]&~m[246]&~m[248]&~m[249])|(~m[244]&~m[245]&~m[246]&m[248]&~m[249])|(m[244]&m[245]&~m[246]&m[248]&~m[249])|(m[244]&~m[245]&m[246]&m[248]&~m[249])|(~m[244]&m[245]&~m[246]&~m[248]&m[249])|(~m[244]&~m[245]&m[246]&~m[248]&m[249])|(m[244]&m[245]&m[246]&~m[248]&m[249])|(~m[244]&m[245]&m[246]&m[248]&m[249]))&UnbiasedRNG[71])|((m[244]&~m[245]&~m[246]&m[248]&~m[249])|(~m[244]&~m[245]&~m[246]&~m[248]&m[249])|(m[244]&~m[245]&~m[246]&~m[248]&m[249])|(m[244]&m[245]&~m[246]&~m[248]&m[249])|(m[244]&~m[245]&m[246]&~m[248]&m[249])|(~m[244]&~m[245]&~m[246]&m[248]&m[249])|(m[244]&~m[245]&~m[246]&m[248]&m[249])|(~m[244]&m[245]&~m[246]&m[248]&m[249])|(m[244]&m[245]&~m[246]&m[248]&m[249])|(~m[244]&~m[245]&m[246]&m[248]&m[249])|(m[244]&~m[245]&m[246]&m[248]&m[249])|(m[244]&m[245]&m[246]&m[248]&m[249]))):InitCond[230];
    m[257] = run?((((m[249]&~m[255]&~m[256]&~m[258]&~m[259])|(~m[249]&~m[255]&~m[256]&m[258]&~m[259])|(m[249]&m[255]&~m[256]&m[258]&~m[259])|(m[249]&~m[255]&m[256]&m[258]&~m[259])|(~m[249]&m[255]&~m[256]&~m[258]&m[259])|(~m[249]&~m[255]&m[256]&~m[258]&m[259])|(m[249]&m[255]&m[256]&~m[258]&m[259])|(~m[249]&m[255]&m[256]&m[258]&m[259]))&UnbiasedRNG[72])|((m[249]&~m[255]&~m[256]&m[258]&~m[259])|(~m[249]&~m[255]&~m[256]&~m[258]&m[259])|(m[249]&~m[255]&~m[256]&~m[258]&m[259])|(m[249]&m[255]&~m[256]&~m[258]&m[259])|(m[249]&~m[255]&m[256]&~m[258]&m[259])|(~m[249]&~m[255]&~m[256]&m[258]&m[259])|(m[249]&~m[255]&~m[256]&m[258]&m[259])|(~m[249]&m[255]&~m[256]&m[258]&m[259])|(m[249]&m[255]&~m[256]&m[258]&m[259])|(~m[249]&~m[255]&m[256]&m[258]&m[259])|(m[249]&~m[255]&m[256]&m[258]&m[259])|(m[249]&m[255]&m[256]&m[258]&m[259]))):InitCond[231];
    m[262] = run?((((m[254]&~m[260]&~m[261]&~m[263]&~m[264])|(~m[254]&~m[260]&~m[261]&m[263]&~m[264])|(m[254]&m[260]&~m[261]&m[263]&~m[264])|(m[254]&~m[260]&m[261]&m[263]&~m[264])|(~m[254]&m[260]&~m[261]&~m[263]&m[264])|(~m[254]&~m[260]&m[261]&~m[263]&m[264])|(m[254]&m[260]&m[261]&~m[263]&m[264])|(~m[254]&m[260]&m[261]&m[263]&m[264]))&UnbiasedRNG[73])|((m[254]&~m[260]&~m[261]&m[263]&~m[264])|(~m[254]&~m[260]&~m[261]&~m[263]&m[264])|(m[254]&~m[260]&~m[261]&~m[263]&m[264])|(m[254]&m[260]&~m[261]&~m[263]&m[264])|(m[254]&~m[260]&m[261]&~m[263]&m[264])|(~m[254]&~m[260]&~m[261]&m[263]&m[264])|(m[254]&~m[260]&~m[261]&m[263]&m[264])|(~m[254]&m[260]&~m[261]&m[263]&m[264])|(m[254]&m[260]&~m[261]&m[263]&m[264])|(~m[254]&~m[260]&m[261]&m[263]&m[264])|(m[254]&~m[260]&m[261]&m[263]&m[264])|(m[254]&m[260]&m[261]&m[263]&m[264]))):InitCond[232];
    m[272] = run?((((m[259]&~m[270]&~m[271]&~m[273]&~m[274])|(~m[259]&~m[270]&~m[271]&m[273]&~m[274])|(m[259]&m[270]&~m[271]&m[273]&~m[274])|(m[259]&~m[270]&m[271]&m[273]&~m[274])|(~m[259]&m[270]&~m[271]&~m[273]&m[274])|(~m[259]&~m[270]&m[271]&~m[273]&m[274])|(m[259]&m[270]&m[271]&~m[273]&m[274])|(~m[259]&m[270]&m[271]&m[273]&m[274]))&UnbiasedRNG[74])|((m[259]&~m[270]&~m[271]&m[273]&~m[274])|(~m[259]&~m[270]&~m[271]&~m[273]&m[274])|(m[259]&~m[270]&~m[271]&~m[273]&m[274])|(m[259]&m[270]&~m[271]&~m[273]&m[274])|(m[259]&~m[270]&m[271]&~m[273]&m[274])|(~m[259]&~m[270]&~m[271]&m[273]&m[274])|(m[259]&~m[270]&~m[271]&m[273]&m[274])|(~m[259]&m[270]&~m[271]&m[273]&m[274])|(m[259]&m[270]&~m[271]&m[273]&m[274])|(~m[259]&~m[270]&m[271]&m[273]&m[274])|(m[259]&~m[270]&m[271]&m[273]&m[274])|(m[259]&m[270]&m[271]&m[273]&m[274]))):InitCond[233];
    m[277] = run?((((m[264]&~m[275]&~m[276]&~m[278]&~m[279])|(~m[264]&~m[275]&~m[276]&m[278]&~m[279])|(m[264]&m[275]&~m[276]&m[278]&~m[279])|(m[264]&~m[275]&m[276]&m[278]&~m[279])|(~m[264]&m[275]&~m[276]&~m[278]&m[279])|(~m[264]&~m[275]&m[276]&~m[278]&m[279])|(m[264]&m[275]&m[276]&~m[278]&m[279])|(~m[264]&m[275]&m[276]&m[278]&m[279]))&UnbiasedRNG[75])|((m[264]&~m[275]&~m[276]&m[278]&~m[279])|(~m[264]&~m[275]&~m[276]&~m[278]&m[279])|(m[264]&~m[275]&~m[276]&~m[278]&m[279])|(m[264]&m[275]&~m[276]&~m[278]&m[279])|(m[264]&~m[275]&m[276]&~m[278]&m[279])|(~m[264]&~m[275]&~m[276]&m[278]&m[279])|(m[264]&~m[275]&~m[276]&m[278]&m[279])|(~m[264]&m[275]&~m[276]&m[278]&m[279])|(m[264]&m[275]&~m[276]&m[278]&m[279])|(~m[264]&~m[275]&m[276]&m[278]&m[279])|(m[264]&~m[275]&m[276]&m[278]&m[279])|(m[264]&m[275]&m[276]&m[278]&m[279]))):InitCond[234];
    m[282] = run?((((m[269]&~m[280]&~m[281]&~m[283]&~m[284])|(~m[269]&~m[280]&~m[281]&m[283]&~m[284])|(m[269]&m[280]&~m[281]&m[283]&~m[284])|(m[269]&~m[280]&m[281]&m[283]&~m[284])|(~m[269]&m[280]&~m[281]&~m[283]&m[284])|(~m[269]&~m[280]&m[281]&~m[283]&m[284])|(m[269]&m[280]&m[281]&~m[283]&m[284])|(~m[269]&m[280]&m[281]&m[283]&m[284]))&UnbiasedRNG[76])|((m[269]&~m[280]&~m[281]&m[283]&~m[284])|(~m[269]&~m[280]&~m[281]&~m[283]&m[284])|(m[269]&~m[280]&~m[281]&~m[283]&m[284])|(m[269]&m[280]&~m[281]&~m[283]&m[284])|(m[269]&~m[280]&m[281]&~m[283]&m[284])|(~m[269]&~m[280]&~m[281]&m[283]&m[284])|(m[269]&~m[280]&~m[281]&m[283]&m[284])|(~m[269]&m[280]&~m[281]&m[283]&m[284])|(m[269]&m[280]&~m[281]&m[283]&m[284])|(~m[269]&~m[280]&m[281]&m[283]&m[284])|(m[269]&~m[280]&m[281]&m[283]&m[284])|(m[269]&m[280]&m[281]&m[283]&m[284]))):InitCond[235];
    m[292] = run?((((m[274]&~m[290]&~m[291]&~m[293]&~m[294])|(~m[274]&~m[290]&~m[291]&m[293]&~m[294])|(m[274]&m[290]&~m[291]&m[293]&~m[294])|(m[274]&~m[290]&m[291]&m[293]&~m[294])|(~m[274]&m[290]&~m[291]&~m[293]&m[294])|(~m[274]&~m[290]&m[291]&~m[293]&m[294])|(m[274]&m[290]&m[291]&~m[293]&m[294])|(~m[274]&m[290]&m[291]&m[293]&m[294]))&UnbiasedRNG[77])|((m[274]&~m[290]&~m[291]&m[293]&~m[294])|(~m[274]&~m[290]&~m[291]&~m[293]&m[294])|(m[274]&~m[290]&~m[291]&~m[293]&m[294])|(m[274]&m[290]&~m[291]&~m[293]&m[294])|(m[274]&~m[290]&m[291]&~m[293]&m[294])|(~m[274]&~m[290]&~m[291]&m[293]&m[294])|(m[274]&~m[290]&~m[291]&m[293]&m[294])|(~m[274]&m[290]&~m[291]&m[293]&m[294])|(m[274]&m[290]&~m[291]&m[293]&m[294])|(~m[274]&~m[290]&m[291]&m[293]&m[294])|(m[274]&~m[290]&m[291]&m[293]&m[294])|(m[274]&m[290]&m[291]&m[293]&m[294]))):InitCond[236];
    m[297] = run?((((m[279]&~m[295]&~m[296]&~m[298]&~m[299])|(~m[279]&~m[295]&~m[296]&m[298]&~m[299])|(m[279]&m[295]&~m[296]&m[298]&~m[299])|(m[279]&~m[295]&m[296]&m[298]&~m[299])|(~m[279]&m[295]&~m[296]&~m[298]&m[299])|(~m[279]&~m[295]&m[296]&~m[298]&m[299])|(m[279]&m[295]&m[296]&~m[298]&m[299])|(~m[279]&m[295]&m[296]&m[298]&m[299]))&UnbiasedRNG[78])|((m[279]&~m[295]&~m[296]&m[298]&~m[299])|(~m[279]&~m[295]&~m[296]&~m[298]&m[299])|(m[279]&~m[295]&~m[296]&~m[298]&m[299])|(m[279]&m[295]&~m[296]&~m[298]&m[299])|(m[279]&~m[295]&m[296]&~m[298]&m[299])|(~m[279]&~m[295]&~m[296]&m[298]&m[299])|(m[279]&~m[295]&~m[296]&m[298]&m[299])|(~m[279]&m[295]&~m[296]&m[298]&m[299])|(m[279]&m[295]&~m[296]&m[298]&m[299])|(~m[279]&~m[295]&m[296]&m[298]&m[299])|(m[279]&~m[295]&m[296]&m[298]&m[299])|(m[279]&m[295]&m[296]&m[298]&m[299]))):InitCond[237];
    m[302] = run?((((m[284]&~m[300]&~m[301]&~m[303]&~m[304])|(~m[284]&~m[300]&~m[301]&m[303]&~m[304])|(m[284]&m[300]&~m[301]&m[303]&~m[304])|(m[284]&~m[300]&m[301]&m[303]&~m[304])|(~m[284]&m[300]&~m[301]&~m[303]&m[304])|(~m[284]&~m[300]&m[301]&~m[303]&m[304])|(m[284]&m[300]&m[301]&~m[303]&m[304])|(~m[284]&m[300]&m[301]&m[303]&m[304]))&UnbiasedRNG[79])|((m[284]&~m[300]&~m[301]&m[303]&~m[304])|(~m[284]&~m[300]&~m[301]&~m[303]&m[304])|(m[284]&~m[300]&~m[301]&~m[303]&m[304])|(m[284]&m[300]&~m[301]&~m[303]&m[304])|(m[284]&~m[300]&m[301]&~m[303]&m[304])|(~m[284]&~m[300]&~m[301]&m[303]&m[304])|(m[284]&~m[300]&~m[301]&m[303]&m[304])|(~m[284]&m[300]&~m[301]&m[303]&m[304])|(m[284]&m[300]&~m[301]&m[303]&m[304])|(~m[284]&~m[300]&m[301]&m[303]&m[304])|(m[284]&~m[300]&m[301]&m[303]&m[304])|(m[284]&m[300]&m[301]&m[303]&m[304]))):InitCond[238];
    m[307] = run?((((m[289]&~m[305]&~m[306]&~m[308]&~m[309])|(~m[289]&~m[305]&~m[306]&m[308]&~m[309])|(m[289]&m[305]&~m[306]&m[308]&~m[309])|(m[289]&~m[305]&m[306]&m[308]&~m[309])|(~m[289]&m[305]&~m[306]&~m[308]&m[309])|(~m[289]&~m[305]&m[306]&~m[308]&m[309])|(m[289]&m[305]&m[306]&~m[308]&m[309])|(~m[289]&m[305]&m[306]&m[308]&m[309]))&UnbiasedRNG[80])|((m[289]&~m[305]&~m[306]&m[308]&~m[309])|(~m[289]&~m[305]&~m[306]&~m[308]&m[309])|(m[289]&~m[305]&~m[306]&~m[308]&m[309])|(m[289]&m[305]&~m[306]&~m[308]&m[309])|(m[289]&~m[305]&m[306]&~m[308]&m[309])|(~m[289]&~m[305]&~m[306]&m[308]&m[309])|(m[289]&~m[305]&~m[306]&m[308]&m[309])|(~m[289]&m[305]&~m[306]&m[308]&m[309])|(m[289]&m[305]&~m[306]&m[308]&m[309])|(~m[289]&~m[305]&m[306]&m[308]&m[309])|(m[289]&~m[305]&m[306]&m[308]&m[309])|(m[289]&m[305]&m[306]&m[308]&m[309]))):InitCond[239];
    m[317] = run?((((m[294]&~m[315]&~m[316]&~m[318]&~m[319])|(~m[294]&~m[315]&~m[316]&m[318]&~m[319])|(m[294]&m[315]&~m[316]&m[318]&~m[319])|(m[294]&~m[315]&m[316]&m[318]&~m[319])|(~m[294]&m[315]&~m[316]&~m[318]&m[319])|(~m[294]&~m[315]&m[316]&~m[318]&m[319])|(m[294]&m[315]&m[316]&~m[318]&m[319])|(~m[294]&m[315]&m[316]&m[318]&m[319]))&UnbiasedRNG[81])|((m[294]&~m[315]&~m[316]&m[318]&~m[319])|(~m[294]&~m[315]&~m[316]&~m[318]&m[319])|(m[294]&~m[315]&~m[316]&~m[318]&m[319])|(m[294]&m[315]&~m[316]&~m[318]&m[319])|(m[294]&~m[315]&m[316]&~m[318]&m[319])|(~m[294]&~m[315]&~m[316]&m[318]&m[319])|(m[294]&~m[315]&~m[316]&m[318]&m[319])|(~m[294]&m[315]&~m[316]&m[318]&m[319])|(m[294]&m[315]&~m[316]&m[318]&m[319])|(~m[294]&~m[315]&m[316]&m[318]&m[319])|(m[294]&~m[315]&m[316]&m[318]&m[319])|(m[294]&m[315]&m[316]&m[318]&m[319]))):InitCond[240];
    m[322] = run?((((m[299]&~m[320]&~m[321]&~m[323]&~m[324])|(~m[299]&~m[320]&~m[321]&m[323]&~m[324])|(m[299]&m[320]&~m[321]&m[323]&~m[324])|(m[299]&~m[320]&m[321]&m[323]&~m[324])|(~m[299]&m[320]&~m[321]&~m[323]&m[324])|(~m[299]&~m[320]&m[321]&~m[323]&m[324])|(m[299]&m[320]&m[321]&~m[323]&m[324])|(~m[299]&m[320]&m[321]&m[323]&m[324]))&UnbiasedRNG[82])|((m[299]&~m[320]&~m[321]&m[323]&~m[324])|(~m[299]&~m[320]&~m[321]&~m[323]&m[324])|(m[299]&~m[320]&~m[321]&~m[323]&m[324])|(m[299]&m[320]&~m[321]&~m[323]&m[324])|(m[299]&~m[320]&m[321]&~m[323]&m[324])|(~m[299]&~m[320]&~m[321]&m[323]&m[324])|(m[299]&~m[320]&~m[321]&m[323]&m[324])|(~m[299]&m[320]&~m[321]&m[323]&m[324])|(m[299]&m[320]&~m[321]&m[323]&m[324])|(~m[299]&~m[320]&m[321]&m[323]&m[324])|(m[299]&~m[320]&m[321]&m[323]&m[324])|(m[299]&m[320]&m[321]&m[323]&m[324]))):InitCond[241];
    m[327] = run?((((m[304]&~m[325]&~m[326]&~m[328]&~m[329])|(~m[304]&~m[325]&~m[326]&m[328]&~m[329])|(m[304]&m[325]&~m[326]&m[328]&~m[329])|(m[304]&~m[325]&m[326]&m[328]&~m[329])|(~m[304]&m[325]&~m[326]&~m[328]&m[329])|(~m[304]&~m[325]&m[326]&~m[328]&m[329])|(m[304]&m[325]&m[326]&~m[328]&m[329])|(~m[304]&m[325]&m[326]&m[328]&m[329]))&UnbiasedRNG[83])|((m[304]&~m[325]&~m[326]&m[328]&~m[329])|(~m[304]&~m[325]&~m[326]&~m[328]&m[329])|(m[304]&~m[325]&~m[326]&~m[328]&m[329])|(m[304]&m[325]&~m[326]&~m[328]&m[329])|(m[304]&~m[325]&m[326]&~m[328]&m[329])|(~m[304]&~m[325]&~m[326]&m[328]&m[329])|(m[304]&~m[325]&~m[326]&m[328]&m[329])|(~m[304]&m[325]&~m[326]&m[328]&m[329])|(m[304]&m[325]&~m[326]&m[328]&m[329])|(~m[304]&~m[325]&m[326]&m[328]&m[329])|(m[304]&~m[325]&m[326]&m[328]&m[329])|(m[304]&m[325]&m[326]&m[328]&m[329]))):InitCond[242];
    m[332] = run?((((m[309]&~m[330]&~m[331]&~m[333]&~m[334])|(~m[309]&~m[330]&~m[331]&m[333]&~m[334])|(m[309]&m[330]&~m[331]&m[333]&~m[334])|(m[309]&~m[330]&m[331]&m[333]&~m[334])|(~m[309]&m[330]&~m[331]&~m[333]&m[334])|(~m[309]&~m[330]&m[331]&~m[333]&m[334])|(m[309]&m[330]&m[331]&~m[333]&m[334])|(~m[309]&m[330]&m[331]&m[333]&m[334]))&UnbiasedRNG[84])|((m[309]&~m[330]&~m[331]&m[333]&~m[334])|(~m[309]&~m[330]&~m[331]&~m[333]&m[334])|(m[309]&~m[330]&~m[331]&~m[333]&m[334])|(m[309]&m[330]&~m[331]&~m[333]&m[334])|(m[309]&~m[330]&m[331]&~m[333]&m[334])|(~m[309]&~m[330]&~m[331]&m[333]&m[334])|(m[309]&~m[330]&~m[331]&m[333]&m[334])|(~m[309]&m[330]&~m[331]&m[333]&m[334])|(m[309]&m[330]&~m[331]&m[333]&m[334])|(~m[309]&~m[330]&m[331]&m[333]&m[334])|(m[309]&~m[330]&m[331]&m[333]&m[334])|(m[309]&m[330]&m[331]&m[333]&m[334]))):InitCond[243];
    m[337] = run?((((m[314]&~m[335]&~m[336]&~m[338]&~m[339])|(~m[314]&~m[335]&~m[336]&m[338]&~m[339])|(m[314]&m[335]&~m[336]&m[338]&~m[339])|(m[314]&~m[335]&m[336]&m[338]&~m[339])|(~m[314]&m[335]&~m[336]&~m[338]&m[339])|(~m[314]&~m[335]&m[336]&~m[338]&m[339])|(m[314]&m[335]&m[336]&~m[338]&m[339])|(~m[314]&m[335]&m[336]&m[338]&m[339]))&UnbiasedRNG[85])|((m[314]&~m[335]&~m[336]&m[338]&~m[339])|(~m[314]&~m[335]&~m[336]&~m[338]&m[339])|(m[314]&~m[335]&~m[336]&~m[338]&m[339])|(m[314]&m[335]&~m[336]&~m[338]&m[339])|(m[314]&~m[335]&m[336]&~m[338]&m[339])|(~m[314]&~m[335]&~m[336]&m[338]&m[339])|(m[314]&~m[335]&~m[336]&m[338]&m[339])|(~m[314]&m[335]&~m[336]&m[338]&m[339])|(m[314]&m[335]&~m[336]&m[338]&m[339])|(~m[314]&~m[335]&m[336]&m[338]&m[339])|(m[314]&~m[335]&m[336]&m[338]&m[339])|(m[314]&m[335]&m[336]&m[338]&m[339]))):InitCond[244];
    m[347] = run?((((m[319]&~m[345]&~m[346]&~m[348]&~m[349])|(~m[319]&~m[345]&~m[346]&m[348]&~m[349])|(m[319]&m[345]&~m[346]&m[348]&~m[349])|(m[319]&~m[345]&m[346]&m[348]&~m[349])|(~m[319]&m[345]&~m[346]&~m[348]&m[349])|(~m[319]&~m[345]&m[346]&~m[348]&m[349])|(m[319]&m[345]&m[346]&~m[348]&m[349])|(~m[319]&m[345]&m[346]&m[348]&m[349]))&UnbiasedRNG[86])|((m[319]&~m[345]&~m[346]&m[348]&~m[349])|(~m[319]&~m[345]&~m[346]&~m[348]&m[349])|(m[319]&~m[345]&~m[346]&~m[348]&m[349])|(m[319]&m[345]&~m[346]&~m[348]&m[349])|(m[319]&~m[345]&m[346]&~m[348]&m[349])|(~m[319]&~m[345]&~m[346]&m[348]&m[349])|(m[319]&~m[345]&~m[346]&m[348]&m[349])|(~m[319]&m[345]&~m[346]&m[348]&m[349])|(m[319]&m[345]&~m[346]&m[348]&m[349])|(~m[319]&~m[345]&m[346]&m[348]&m[349])|(m[319]&~m[345]&m[346]&m[348]&m[349])|(m[319]&m[345]&m[346]&m[348]&m[349]))):InitCond[245];
    m[352] = run?((((m[324]&~m[350]&~m[351]&~m[353]&~m[354])|(~m[324]&~m[350]&~m[351]&m[353]&~m[354])|(m[324]&m[350]&~m[351]&m[353]&~m[354])|(m[324]&~m[350]&m[351]&m[353]&~m[354])|(~m[324]&m[350]&~m[351]&~m[353]&m[354])|(~m[324]&~m[350]&m[351]&~m[353]&m[354])|(m[324]&m[350]&m[351]&~m[353]&m[354])|(~m[324]&m[350]&m[351]&m[353]&m[354]))&UnbiasedRNG[87])|((m[324]&~m[350]&~m[351]&m[353]&~m[354])|(~m[324]&~m[350]&~m[351]&~m[353]&m[354])|(m[324]&~m[350]&~m[351]&~m[353]&m[354])|(m[324]&m[350]&~m[351]&~m[353]&m[354])|(m[324]&~m[350]&m[351]&~m[353]&m[354])|(~m[324]&~m[350]&~m[351]&m[353]&m[354])|(m[324]&~m[350]&~m[351]&m[353]&m[354])|(~m[324]&m[350]&~m[351]&m[353]&m[354])|(m[324]&m[350]&~m[351]&m[353]&m[354])|(~m[324]&~m[350]&m[351]&m[353]&m[354])|(m[324]&~m[350]&m[351]&m[353]&m[354])|(m[324]&m[350]&m[351]&m[353]&m[354]))):InitCond[246];
    m[357] = run?((((m[329]&~m[355]&~m[356]&~m[358]&~m[359])|(~m[329]&~m[355]&~m[356]&m[358]&~m[359])|(m[329]&m[355]&~m[356]&m[358]&~m[359])|(m[329]&~m[355]&m[356]&m[358]&~m[359])|(~m[329]&m[355]&~m[356]&~m[358]&m[359])|(~m[329]&~m[355]&m[356]&~m[358]&m[359])|(m[329]&m[355]&m[356]&~m[358]&m[359])|(~m[329]&m[355]&m[356]&m[358]&m[359]))&UnbiasedRNG[88])|((m[329]&~m[355]&~m[356]&m[358]&~m[359])|(~m[329]&~m[355]&~m[356]&~m[358]&m[359])|(m[329]&~m[355]&~m[356]&~m[358]&m[359])|(m[329]&m[355]&~m[356]&~m[358]&m[359])|(m[329]&~m[355]&m[356]&~m[358]&m[359])|(~m[329]&~m[355]&~m[356]&m[358]&m[359])|(m[329]&~m[355]&~m[356]&m[358]&m[359])|(~m[329]&m[355]&~m[356]&m[358]&m[359])|(m[329]&m[355]&~m[356]&m[358]&m[359])|(~m[329]&~m[355]&m[356]&m[358]&m[359])|(m[329]&~m[355]&m[356]&m[358]&m[359])|(m[329]&m[355]&m[356]&m[358]&m[359]))):InitCond[247];
    m[362] = run?((((m[334]&~m[360]&~m[361]&~m[363]&~m[364])|(~m[334]&~m[360]&~m[361]&m[363]&~m[364])|(m[334]&m[360]&~m[361]&m[363]&~m[364])|(m[334]&~m[360]&m[361]&m[363]&~m[364])|(~m[334]&m[360]&~m[361]&~m[363]&m[364])|(~m[334]&~m[360]&m[361]&~m[363]&m[364])|(m[334]&m[360]&m[361]&~m[363]&m[364])|(~m[334]&m[360]&m[361]&m[363]&m[364]))&UnbiasedRNG[89])|((m[334]&~m[360]&~m[361]&m[363]&~m[364])|(~m[334]&~m[360]&~m[361]&~m[363]&m[364])|(m[334]&~m[360]&~m[361]&~m[363]&m[364])|(m[334]&m[360]&~m[361]&~m[363]&m[364])|(m[334]&~m[360]&m[361]&~m[363]&m[364])|(~m[334]&~m[360]&~m[361]&m[363]&m[364])|(m[334]&~m[360]&~m[361]&m[363]&m[364])|(~m[334]&m[360]&~m[361]&m[363]&m[364])|(m[334]&m[360]&~m[361]&m[363]&m[364])|(~m[334]&~m[360]&m[361]&m[363]&m[364])|(m[334]&~m[360]&m[361]&m[363]&m[364])|(m[334]&m[360]&m[361]&m[363]&m[364]))):InitCond[248];
    m[367] = run?((((m[339]&~m[365]&~m[366]&~m[368]&~m[369])|(~m[339]&~m[365]&~m[366]&m[368]&~m[369])|(m[339]&m[365]&~m[366]&m[368]&~m[369])|(m[339]&~m[365]&m[366]&m[368]&~m[369])|(~m[339]&m[365]&~m[366]&~m[368]&m[369])|(~m[339]&~m[365]&m[366]&~m[368]&m[369])|(m[339]&m[365]&m[366]&~m[368]&m[369])|(~m[339]&m[365]&m[366]&m[368]&m[369]))&UnbiasedRNG[90])|((m[339]&~m[365]&~m[366]&m[368]&~m[369])|(~m[339]&~m[365]&~m[366]&~m[368]&m[369])|(m[339]&~m[365]&~m[366]&~m[368]&m[369])|(m[339]&m[365]&~m[366]&~m[368]&m[369])|(m[339]&~m[365]&m[366]&~m[368]&m[369])|(~m[339]&~m[365]&~m[366]&m[368]&m[369])|(m[339]&~m[365]&~m[366]&m[368]&m[369])|(~m[339]&m[365]&~m[366]&m[368]&m[369])|(m[339]&m[365]&~m[366]&m[368]&m[369])|(~m[339]&~m[365]&m[366]&m[368]&m[369])|(m[339]&~m[365]&m[366]&m[368]&m[369])|(m[339]&m[365]&m[366]&m[368]&m[369]))):InitCond[249];
    m[372] = run?((((m[344]&~m[370]&~m[371]&~m[373]&~m[374])|(~m[344]&~m[370]&~m[371]&m[373]&~m[374])|(m[344]&m[370]&~m[371]&m[373]&~m[374])|(m[344]&~m[370]&m[371]&m[373]&~m[374])|(~m[344]&m[370]&~m[371]&~m[373]&m[374])|(~m[344]&~m[370]&m[371]&~m[373]&m[374])|(m[344]&m[370]&m[371]&~m[373]&m[374])|(~m[344]&m[370]&m[371]&m[373]&m[374]))&UnbiasedRNG[91])|((m[344]&~m[370]&~m[371]&m[373]&~m[374])|(~m[344]&~m[370]&~m[371]&~m[373]&m[374])|(m[344]&~m[370]&~m[371]&~m[373]&m[374])|(m[344]&m[370]&~m[371]&~m[373]&m[374])|(m[344]&~m[370]&m[371]&~m[373]&m[374])|(~m[344]&~m[370]&~m[371]&m[373]&m[374])|(m[344]&~m[370]&~m[371]&m[373]&m[374])|(~m[344]&m[370]&~m[371]&m[373]&m[374])|(m[344]&m[370]&~m[371]&m[373]&m[374])|(~m[344]&~m[370]&m[371]&m[373]&m[374])|(m[344]&~m[370]&m[371]&m[373]&m[374])|(m[344]&m[370]&m[371]&m[373]&m[374]))):InitCond[250];
    m[382] = run?((((m[349]&~m[380]&~m[381]&~m[383]&~m[384])|(~m[349]&~m[380]&~m[381]&m[383]&~m[384])|(m[349]&m[380]&~m[381]&m[383]&~m[384])|(m[349]&~m[380]&m[381]&m[383]&~m[384])|(~m[349]&m[380]&~m[381]&~m[383]&m[384])|(~m[349]&~m[380]&m[381]&~m[383]&m[384])|(m[349]&m[380]&m[381]&~m[383]&m[384])|(~m[349]&m[380]&m[381]&m[383]&m[384]))&UnbiasedRNG[92])|((m[349]&~m[380]&~m[381]&m[383]&~m[384])|(~m[349]&~m[380]&~m[381]&~m[383]&m[384])|(m[349]&~m[380]&~m[381]&~m[383]&m[384])|(m[349]&m[380]&~m[381]&~m[383]&m[384])|(m[349]&~m[380]&m[381]&~m[383]&m[384])|(~m[349]&~m[380]&~m[381]&m[383]&m[384])|(m[349]&~m[380]&~m[381]&m[383]&m[384])|(~m[349]&m[380]&~m[381]&m[383]&m[384])|(m[349]&m[380]&~m[381]&m[383]&m[384])|(~m[349]&~m[380]&m[381]&m[383]&m[384])|(m[349]&~m[380]&m[381]&m[383]&m[384])|(m[349]&m[380]&m[381]&m[383]&m[384]))):InitCond[251];
    m[387] = run?((((m[354]&~m[385]&~m[386]&~m[388]&~m[389])|(~m[354]&~m[385]&~m[386]&m[388]&~m[389])|(m[354]&m[385]&~m[386]&m[388]&~m[389])|(m[354]&~m[385]&m[386]&m[388]&~m[389])|(~m[354]&m[385]&~m[386]&~m[388]&m[389])|(~m[354]&~m[385]&m[386]&~m[388]&m[389])|(m[354]&m[385]&m[386]&~m[388]&m[389])|(~m[354]&m[385]&m[386]&m[388]&m[389]))&UnbiasedRNG[93])|((m[354]&~m[385]&~m[386]&m[388]&~m[389])|(~m[354]&~m[385]&~m[386]&~m[388]&m[389])|(m[354]&~m[385]&~m[386]&~m[388]&m[389])|(m[354]&m[385]&~m[386]&~m[388]&m[389])|(m[354]&~m[385]&m[386]&~m[388]&m[389])|(~m[354]&~m[385]&~m[386]&m[388]&m[389])|(m[354]&~m[385]&~m[386]&m[388]&m[389])|(~m[354]&m[385]&~m[386]&m[388]&m[389])|(m[354]&m[385]&~m[386]&m[388]&m[389])|(~m[354]&~m[385]&m[386]&m[388]&m[389])|(m[354]&~m[385]&m[386]&m[388]&m[389])|(m[354]&m[385]&m[386]&m[388]&m[389]))):InitCond[252];
    m[392] = run?((((m[359]&~m[390]&~m[391]&~m[393]&~m[394])|(~m[359]&~m[390]&~m[391]&m[393]&~m[394])|(m[359]&m[390]&~m[391]&m[393]&~m[394])|(m[359]&~m[390]&m[391]&m[393]&~m[394])|(~m[359]&m[390]&~m[391]&~m[393]&m[394])|(~m[359]&~m[390]&m[391]&~m[393]&m[394])|(m[359]&m[390]&m[391]&~m[393]&m[394])|(~m[359]&m[390]&m[391]&m[393]&m[394]))&UnbiasedRNG[94])|((m[359]&~m[390]&~m[391]&m[393]&~m[394])|(~m[359]&~m[390]&~m[391]&~m[393]&m[394])|(m[359]&~m[390]&~m[391]&~m[393]&m[394])|(m[359]&m[390]&~m[391]&~m[393]&m[394])|(m[359]&~m[390]&m[391]&~m[393]&m[394])|(~m[359]&~m[390]&~m[391]&m[393]&m[394])|(m[359]&~m[390]&~m[391]&m[393]&m[394])|(~m[359]&m[390]&~m[391]&m[393]&m[394])|(m[359]&m[390]&~m[391]&m[393]&m[394])|(~m[359]&~m[390]&m[391]&m[393]&m[394])|(m[359]&~m[390]&m[391]&m[393]&m[394])|(m[359]&m[390]&m[391]&m[393]&m[394]))):InitCond[253];
    m[397] = run?((((m[364]&~m[395]&~m[396]&~m[398]&~m[399])|(~m[364]&~m[395]&~m[396]&m[398]&~m[399])|(m[364]&m[395]&~m[396]&m[398]&~m[399])|(m[364]&~m[395]&m[396]&m[398]&~m[399])|(~m[364]&m[395]&~m[396]&~m[398]&m[399])|(~m[364]&~m[395]&m[396]&~m[398]&m[399])|(m[364]&m[395]&m[396]&~m[398]&m[399])|(~m[364]&m[395]&m[396]&m[398]&m[399]))&UnbiasedRNG[95])|((m[364]&~m[395]&~m[396]&m[398]&~m[399])|(~m[364]&~m[395]&~m[396]&~m[398]&m[399])|(m[364]&~m[395]&~m[396]&~m[398]&m[399])|(m[364]&m[395]&~m[396]&~m[398]&m[399])|(m[364]&~m[395]&m[396]&~m[398]&m[399])|(~m[364]&~m[395]&~m[396]&m[398]&m[399])|(m[364]&~m[395]&~m[396]&m[398]&m[399])|(~m[364]&m[395]&~m[396]&m[398]&m[399])|(m[364]&m[395]&~m[396]&m[398]&m[399])|(~m[364]&~m[395]&m[396]&m[398]&m[399])|(m[364]&~m[395]&m[396]&m[398]&m[399])|(m[364]&m[395]&m[396]&m[398]&m[399]))):InitCond[254];
    m[402] = run?((((m[369]&~m[400]&~m[401]&~m[403]&~m[404])|(~m[369]&~m[400]&~m[401]&m[403]&~m[404])|(m[369]&m[400]&~m[401]&m[403]&~m[404])|(m[369]&~m[400]&m[401]&m[403]&~m[404])|(~m[369]&m[400]&~m[401]&~m[403]&m[404])|(~m[369]&~m[400]&m[401]&~m[403]&m[404])|(m[369]&m[400]&m[401]&~m[403]&m[404])|(~m[369]&m[400]&m[401]&m[403]&m[404]))&UnbiasedRNG[96])|((m[369]&~m[400]&~m[401]&m[403]&~m[404])|(~m[369]&~m[400]&~m[401]&~m[403]&m[404])|(m[369]&~m[400]&~m[401]&~m[403]&m[404])|(m[369]&m[400]&~m[401]&~m[403]&m[404])|(m[369]&~m[400]&m[401]&~m[403]&m[404])|(~m[369]&~m[400]&~m[401]&m[403]&m[404])|(m[369]&~m[400]&~m[401]&m[403]&m[404])|(~m[369]&m[400]&~m[401]&m[403]&m[404])|(m[369]&m[400]&~m[401]&m[403]&m[404])|(~m[369]&~m[400]&m[401]&m[403]&m[404])|(m[369]&~m[400]&m[401]&m[403]&m[404])|(m[369]&m[400]&m[401]&m[403]&m[404]))):InitCond[255];
    m[407] = run?((((m[374]&~m[405]&~m[406]&~m[408]&~m[409])|(~m[374]&~m[405]&~m[406]&m[408]&~m[409])|(m[374]&m[405]&~m[406]&m[408]&~m[409])|(m[374]&~m[405]&m[406]&m[408]&~m[409])|(~m[374]&m[405]&~m[406]&~m[408]&m[409])|(~m[374]&~m[405]&m[406]&~m[408]&m[409])|(m[374]&m[405]&m[406]&~m[408]&m[409])|(~m[374]&m[405]&m[406]&m[408]&m[409]))&UnbiasedRNG[97])|((m[374]&~m[405]&~m[406]&m[408]&~m[409])|(~m[374]&~m[405]&~m[406]&~m[408]&m[409])|(m[374]&~m[405]&~m[406]&~m[408]&m[409])|(m[374]&m[405]&~m[406]&~m[408]&m[409])|(m[374]&~m[405]&m[406]&~m[408]&m[409])|(~m[374]&~m[405]&~m[406]&m[408]&m[409])|(m[374]&~m[405]&~m[406]&m[408]&m[409])|(~m[374]&m[405]&~m[406]&m[408]&m[409])|(m[374]&m[405]&~m[406]&m[408]&m[409])|(~m[374]&~m[405]&m[406]&m[408]&m[409])|(m[374]&~m[405]&m[406]&m[408]&m[409])|(m[374]&m[405]&m[406]&m[408]&m[409]))):InitCond[256];
    m[412] = run?((((m[379]&~m[410]&~m[411]&~m[413]&~m[414])|(~m[379]&~m[410]&~m[411]&m[413]&~m[414])|(m[379]&m[410]&~m[411]&m[413]&~m[414])|(m[379]&~m[410]&m[411]&m[413]&~m[414])|(~m[379]&m[410]&~m[411]&~m[413]&m[414])|(~m[379]&~m[410]&m[411]&~m[413]&m[414])|(m[379]&m[410]&m[411]&~m[413]&m[414])|(~m[379]&m[410]&m[411]&m[413]&m[414]))&UnbiasedRNG[98])|((m[379]&~m[410]&~m[411]&m[413]&~m[414])|(~m[379]&~m[410]&~m[411]&~m[413]&m[414])|(m[379]&~m[410]&~m[411]&~m[413]&m[414])|(m[379]&m[410]&~m[411]&~m[413]&m[414])|(m[379]&~m[410]&m[411]&~m[413]&m[414])|(~m[379]&~m[410]&~m[411]&m[413]&m[414])|(m[379]&~m[410]&~m[411]&m[413]&m[414])|(~m[379]&m[410]&~m[411]&m[413]&m[414])|(m[379]&m[410]&~m[411]&m[413]&m[414])|(~m[379]&~m[410]&m[411]&m[413]&m[414])|(m[379]&~m[410]&m[411]&m[413]&m[414])|(m[379]&m[410]&m[411]&m[413]&m[414]))):InitCond[257];
    m[417] = run?((((m[389]&~m[415]&~m[416]&~m[418]&~m[419])|(~m[389]&~m[415]&~m[416]&m[418]&~m[419])|(m[389]&m[415]&~m[416]&m[418]&~m[419])|(m[389]&~m[415]&m[416]&m[418]&~m[419])|(~m[389]&m[415]&~m[416]&~m[418]&m[419])|(~m[389]&~m[415]&m[416]&~m[418]&m[419])|(m[389]&m[415]&m[416]&~m[418]&m[419])|(~m[389]&m[415]&m[416]&m[418]&m[419]))&UnbiasedRNG[99])|((m[389]&~m[415]&~m[416]&m[418]&~m[419])|(~m[389]&~m[415]&~m[416]&~m[418]&m[419])|(m[389]&~m[415]&~m[416]&~m[418]&m[419])|(m[389]&m[415]&~m[416]&~m[418]&m[419])|(m[389]&~m[415]&m[416]&~m[418]&m[419])|(~m[389]&~m[415]&~m[416]&m[418]&m[419])|(m[389]&~m[415]&~m[416]&m[418]&m[419])|(~m[389]&m[415]&~m[416]&m[418]&m[419])|(m[389]&m[415]&~m[416]&m[418]&m[419])|(~m[389]&~m[415]&m[416]&m[418]&m[419])|(m[389]&~m[415]&m[416]&m[418]&m[419])|(m[389]&m[415]&m[416]&m[418]&m[419]))):InitCond[258];
    m[422] = run?((((m[394]&~m[420]&~m[421]&~m[423]&~m[424])|(~m[394]&~m[420]&~m[421]&m[423]&~m[424])|(m[394]&m[420]&~m[421]&m[423]&~m[424])|(m[394]&~m[420]&m[421]&m[423]&~m[424])|(~m[394]&m[420]&~m[421]&~m[423]&m[424])|(~m[394]&~m[420]&m[421]&~m[423]&m[424])|(m[394]&m[420]&m[421]&~m[423]&m[424])|(~m[394]&m[420]&m[421]&m[423]&m[424]))&UnbiasedRNG[100])|((m[394]&~m[420]&~m[421]&m[423]&~m[424])|(~m[394]&~m[420]&~m[421]&~m[423]&m[424])|(m[394]&~m[420]&~m[421]&~m[423]&m[424])|(m[394]&m[420]&~m[421]&~m[423]&m[424])|(m[394]&~m[420]&m[421]&~m[423]&m[424])|(~m[394]&~m[420]&~m[421]&m[423]&m[424])|(m[394]&~m[420]&~m[421]&m[423]&m[424])|(~m[394]&m[420]&~m[421]&m[423]&m[424])|(m[394]&m[420]&~m[421]&m[423]&m[424])|(~m[394]&~m[420]&m[421]&m[423]&m[424])|(m[394]&~m[420]&m[421]&m[423]&m[424])|(m[394]&m[420]&m[421]&m[423]&m[424]))):InitCond[259];
    m[427] = run?((((m[399]&~m[425]&~m[426]&~m[428]&~m[429])|(~m[399]&~m[425]&~m[426]&m[428]&~m[429])|(m[399]&m[425]&~m[426]&m[428]&~m[429])|(m[399]&~m[425]&m[426]&m[428]&~m[429])|(~m[399]&m[425]&~m[426]&~m[428]&m[429])|(~m[399]&~m[425]&m[426]&~m[428]&m[429])|(m[399]&m[425]&m[426]&~m[428]&m[429])|(~m[399]&m[425]&m[426]&m[428]&m[429]))&UnbiasedRNG[101])|((m[399]&~m[425]&~m[426]&m[428]&~m[429])|(~m[399]&~m[425]&~m[426]&~m[428]&m[429])|(m[399]&~m[425]&~m[426]&~m[428]&m[429])|(m[399]&m[425]&~m[426]&~m[428]&m[429])|(m[399]&~m[425]&m[426]&~m[428]&m[429])|(~m[399]&~m[425]&~m[426]&m[428]&m[429])|(m[399]&~m[425]&~m[426]&m[428]&m[429])|(~m[399]&m[425]&~m[426]&m[428]&m[429])|(m[399]&m[425]&~m[426]&m[428]&m[429])|(~m[399]&~m[425]&m[426]&m[428]&m[429])|(m[399]&~m[425]&m[426]&m[428]&m[429])|(m[399]&m[425]&m[426]&m[428]&m[429]))):InitCond[260];
    m[432] = run?((((m[404]&~m[430]&~m[431]&~m[433]&~m[434])|(~m[404]&~m[430]&~m[431]&m[433]&~m[434])|(m[404]&m[430]&~m[431]&m[433]&~m[434])|(m[404]&~m[430]&m[431]&m[433]&~m[434])|(~m[404]&m[430]&~m[431]&~m[433]&m[434])|(~m[404]&~m[430]&m[431]&~m[433]&m[434])|(m[404]&m[430]&m[431]&~m[433]&m[434])|(~m[404]&m[430]&m[431]&m[433]&m[434]))&UnbiasedRNG[102])|((m[404]&~m[430]&~m[431]&m[433]&~m[434])|(~m[404]&~m[430]&~m[431]&~m[433]&m[434])|(m[404]&~m[430]&~m[431]&~m[433]&m[434])|(m[404]&m[430]&~m[431]&~m[433]&m[434])|(m[404]&~m[430]&m[431]&~m[433]&m[434])|(~m[404]&~m[430]&~m[431]&m[433]&m[434])|(m[404]&~m[430]&~m[431]&m[433]&m[434])|(~m[404]&m[430]&~m[431]&m[433]&m[434])|(m[404]&m[430]&~m[431]&m[433]&m[434])|(~m[404]&~m[430]&m[431]&m[433]&m[434])|(m[404]&~m[430]&m[431]&m[433]&m[434])|(m[404]&m[430]&m[431]&m[433]&m[434]))):InitCond[261];
    m[437] = run?((((m[409]&~m[435]&~m[436]&~m[438]&~m[439])|(~m[409]&~m[435]&~m[436]&m[438]&~m[439])|(m[409]&m[435]&~m[436]&m[438]&~m[439])|(m[409]&~m[435]&m[436]&m[438]&~m[439])|(~m[409]&m[435]&~m[436]&~m[438]&m[439])|(~m[409]&~m[435]&m[436]&~m[438]&m[439])|(m[409]&m[435]&m[436]&~m[438]&m[439])|(~m[409]&m[435]&m[436]&m[438]&m[439]))&UnbiasedRNG[103])|((m[409]&~m[435]&~m[436]&m[438]&~m[439])|(~m[409]&~m[435]&~m[436]&~m[438]&m[439])|(m[409]&~m[435]&~m[436]&~m[438]&m[439])|(m[409]&m[435]&~m[436]&~m[438]&m[439])|(m[409]&~m[435]&m[436]&~m[438]&m[439])|(~m[409]&~m[435]&~m[436]&m[438]&m[439])|(m[409]&~m[435]&~m[436]&m[438]&m[439])|(~m[409]&m[435]&~m[436]&m[438]&m[439])|(m[409]&m[435]&~m[436]&m[438]&m[439])|(~m[409]&~m[435]&m[436]&m[438]&m[439])|(m[409]&~m[435]&m[436]&m[438]&m[439])|(m[409]&m[435]&m[436]&m[438]&m[439]))):InitCond[262];
    m[442] = run?((((m[414]&~m[440]&~m[441]&~m[443]&~m[444])|(~m[414]&~m[440]&~m[441]&m[443]&~m[444])|(m[414]&m[440]&~m[441]&m[443]&~m[444])|(m[414]&~m[440]&m[441]&m[443]&~m[444])|(~m[414]&m[440]&~m[441]&~m[443]&m[444])|(~m[414]&~m[440]&m[441]&~m[443]&m[444])|(m[414]&m[440]&m[441]&~m[443]&m[444])|(~m[414]&m[440]&m[441]&m[443]&m[444]))&UnbiasedRNG[104])|((m[414]&~m[440]&~m[441]&m[443]&~m[444])|(~m[414]&~m[440]&~m[441]&~m[443]&m[444])|(m[414]&~m[440]&~m[441]&~m[443]&m[444])|(m[414]&m[440]&~m[441]&~m[443]&m[444])|(m[414]&~m[440]&m[441]&~m[443]&m[444])|(~m[414]&~m[440]&~m[441]&m[443]&m[444])|(m[414]&~m[440]&~m[441]&m[443]&m[444])|(~m[414]&m[440]&~m[441]&m[443]&m[444])|(m[414]&m[440]&~m[441]&m[443]&m[444])|(~m[414]&~m[440]&m[441]&m[443]&m[444])|(m[414]&~m[440]&m[441]&m[443]&m[444])|(m[414]&m[440]&m[441]&m[443]&m[444]))):InitCond[263];
    m[447] = run?((((m[424]&~m[445]&~m[446]&~m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&m[448]&~m[449])|(m[424]&m[445]&~m[446]&m[448]&~m[449])|(m[424]&~m[445]&m[446]&m[448]&~m[449])|(~m[424]&m[445]&~m[446]&~m[448]&m[449])|(~m[424]&~m[445]&m[446]&~m[448]&m[449])|(m[424]&m[445]&m[446]&~m[448]&m[449])|(~m[424]&m[445]&m[446]&m[448]&m[449]))&UnbiasedRNG[105])|((m[424]&~m[445]&~m[446]&m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&m[446]&~m[448]&m[449])|(~m[424]&~m[445]&~m[446]&m[448]&m[449])|(m[424]&~m[445]&~m[446]&m[448]&m[449])|(~m[424]&m[445]&~m[446]&m[448]&m[449])|(m[424]&m[445]&~m[446]&m[448]&m[449])|(~m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&m[445]&m[446]&m[448]&m[449]))):InitCond[264];
    m[452] = run?((((m[429]&~m[450]&~m[451]&~m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&m[453]&~m[454])|(m[429]&m[450]&~m[451]&m[453]&~m[454])|(m[429]&~m[450]&m[451]&m[453]&~m[454])|(~m[429]&m[450]&~m[451]&~m[453]&m[454])|(~m[429]&~m[450]&m[451]&~m[453]&m[454])|(m[429]&m[450]&m[451]&~m[453]&m[454])|(~m[429]&m[450]&m[451]&m[453]&m[454]))&UnbiasedRNG[106])|((m[429]&~m[450]&~m[451]&m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&m[451]&~m[453]&m[454])|(~m[429]&~m[450]&~m[451]&m[453]&m[454])|(m[429]&~m[450]&~m[451]&m[453]&m[454])|(~m[429]&m[450]&~m[451]&m[453]&m[454])|(m[429]&m[450]&~m[451]&m[453]&m[454])|(~m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&m[450]&m[451]&m[453]&m[454]))):InitCond[265];
    m[457] = run?((((m[434]&~m[455]&~m[456]&~m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&m[458]&~m[459])|(m[434]&m[455]&~m[456]&m[458]&~m[459])|(m[434]&~m[455]&m[456]&m[458]&~m[459])|(~m[434]&m[455]&~m[456]&~m[458]&m[459])|(~m[434]&~m[455]&m[456]&~m[458]&m[459])|(m[434]&m[455]&m[456]&~m[458]&m[459])|(~m[434]&m[455]&m[456]&m[458]&m[459]))&UnbiasedRNG[107])|((m[434]&~m[455]&~m[456]&m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&m[456]&~m[458]&m[459])|(~m[434]&~m[455]&~m[456]&m[458]&m[459])|(m[434]&~m[455]&~m[456]&m[458]&m[459])|(~m[434]&m[455]&~m[456]&m[458]&m[459])|(m[434]&m[455]&~m[456]&m[458]&m[459])|(~m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&m[455]&m[456]&m[458]&m[459]))):InitCond[266];
    m[462] = run?((((m[439]&~m[460]&~m[461]&~m[463]&~m[464])|(~m[439]&~m[460]&~m[461]&m[463]&~m[464])|(m[439]&m[460]&~m[461]&m[463]&~m[464])|(m[439]&~m[460]&m[461]&m[463]&~m[464])|(~m[439]&m[460]&~m[461]&~m[463]&m[464])|(~m[439]&~m[460]&m[461]&~m[463]&m[464])|(m[439]&m[460]&m[461]&~m[463]&m[464])|(~m[439]&m[460]&m[461]&m[463]&m[464]))&UnbiasedRNG[108])|((m[439]&~m[460]&~m[461]&m[463]&~m[464])|(~m[439]&~m[460]&~m[461]&~m[463]&m[464])|(m[439]&~m[460]&~m[461]&~m[463]&m[464])|(m[439]&m[460]&~m[461]&~m[463]&m[464])|(m[439]&~m[460]&m[461]&~m[463]&m[464])|(~m[439]&~m[460]&~m[461]&m[463]&m[464])|(m[439]&~m[460]&~m[461]&m[463]&m[464])|(~m[439]&m[460]&~m[461]&m[463]&m[464])|(m[439]&m[460]&~m[461]&m[463]&m[464])|(~m[439]&~m[460]&m[461]&m[463]&m[464])|(m[439]&~m[460]&m[461]&m[463]&m[464])|(m[439]&m[460]&m[461]&m[463]&m[464]))):InitCond[267];
    m[467] = run?((((m[444]&~m[465]&~m[466]&~m[468]&~m[469])|(~m[444]&~m[465]&~m[466]&m[468]&~m[469])|(m[444]&m[465]&~m[466]&m[468]&~m[469])|(m[444]&~m[465]&m[466]&m[468]&~m[469])|(~m[444]&m[465]&~m[466]&~m[468]&m[469])|(~m[444]&~m[465]&m[466]&~m[468]&m[469])|(m[444]&m[465]&m[466]&~m[468]&m[469])|(~m[444]&m[465]&m[466]&m[468]&m[469]))&UnbiasedRNG[109])|((m[444]&~m[465]&~m[466]&m[468]&~m[469])|(~m[444]&~m[465]&~m[466]&~m[468]&m[469])|(m[444]&~m[465]&~m[466]&~m[468]&m[469])|(m[444]&m[465]&~m[466]&~m[468]&m[469])|(m[444]&~m[465]&m[466]&~m[468]&m[469])|(~m[444]&~m[465]&~m[466]&m[468]&m[469])|(m[444]&~m[465]&~m[466]&m[468]&m[469])|(~m[444]&m[465]&~m[466]&m[468]&m[469])|(m[444]&m[465]&~m[466]&m[468]&m[469])|(~m[444]&~m[465]&m[466]&m[468]&m[469])|(m[444]&~m[465]&m[466]&m[468]&m[469])|(m[444]&m[465]&m[466]&m[468]&m[469]))):InitCond[268];
    m[472] = run?((((m[454]&~m[470]&~m[471]&~m[473]&~m[474])|(~m[454]&~m[470]&~m[471]&m[473]&~m[474])|(m[454]&m[470]&~m[471]&m[473]&~m[474])|(m[454]&~m[470]&m[471]&m[473]&~m[474])|(~m[454]&m[470]&~m[471]&~m[473]&m[474])|(~m[454]&~m[470]&m[471]&~m[473]&m[474])|(m[454]&m[470]&m[471]&~m[473]&m[474])|(~m[454]&m[470]&m[471]&m[473]&m[474]))&UnbiasedRNG[110])|((m[454]&~m[470]&~m[471]&m[473]&~m[474])|(~m[454]&~m[470]&~m[471]&~m[473]&m[474])|(m[454]&~m[470]&~m[471]&~m[473]&m[474])|(m[454]&m[470]&~m[471]&~m[473]&m[474])|(m[454]&~m[470]&m[471]&~m[473]&m[474])|(~m[454]&~m[470]&~m[471]&m[473]&m[474])|(m[454]&~m[470]&~m[471]&m[473]&m[474])|(~m[454]&m[470]&~m[471]&m[473]&m[474])|(m[454]&m[470]&~m[471]&m[473]&m[474])|(~m[454]&~m[470]&m[471]&m[473]&m[474])|(m[454]&~m[470]&m[471]&m[473]&m[474])|(m[454]&m[470]&m[471]&m[473]&m[474]))):InitCond[269];
    m[477] = run?((((m[459]&~m[475]&~m[476]&~m[478]&~m[479])|(~m[459]&~m[475]&~m[476]&m[478]&~m[479])|(m[459]&m[475]&~m[476]&m[478]&~m[479])|(m[459]&~m[475]&m[476]&m[478]&~m[479])|(~m[459]&m[475]&~m[476]&~m[478]&m[479])|(~m[459]&~m[475]&m[476]&~m[478]&m[479])|(m[459]&m[475]&m[476]&~m[478]&m[479])|(~m[459]&m[475]&m[476]&m[478]&m[479]))&UnbiasedRNG[111])|((m[459]&~m[475]&~m[476]&m[478]&~m[479])|(~m[459]&~m[475]&~m[476]&~m[478]&m[479])|(m[459]&~m[475]&~m[476]&~m[478]&m[479])|(m[459]&m[475]&~m[476]&~m[478]&m[479])|(m[459]&~m[475]&m[476]&~m[478]&m[479])|(~m[459]&~m[475]&~m[476]&m[478]&m[479])|(m[459]&~m[475]&~m[476]&m[478]&m[479])|(~m[459]&m[475]&~m[476]&m[478]&m[479])|(m[459]&m[475]&~m[476]&m[478]&m[479])|(~m[459]&~m[475]&m[476]&m[478]&m[479])|(m[459]&~m[475]&m[476]&m[478]&m[479])|(m[459]&m[475]&m[476]&m[478]&m[479]))):InitCond[270];
    m[482] = run?((((m[464]&~m[480]&~m[481]&~m[483]&~m[484])|(~m[464]&~m[480]&~m[481]&m[483]&~m[484])|(m[464]&m[480]&~m[481]&m[483]&~m[484])|(m[464]&~m[480]&m[481]&m[483]&~m[484])|(~m[464]&m[480]&~m[481]&~m[483]&m[484])|(~m[464]&~m[480]&m[481]&~m[483]&m[484])|(m[464]&m[480]&m[481]&~m[483]&m[484])|(~m[464]&m[480]&m[481]&m[483]&m[484]))&UnbiasedRNG[112])|((m[464]&~m[480]&~m[481]&m[483]&~m[484])|(~m[464]&~m[480]&~m[481]&~m[483]&m[484])|(m[464]&~m[480]&~m[481]&~m[483]&m[484])|(m[464]&m[480]&~m[481]&~m[483]&m[484])|(m[464]&~m[480]&m[481]&~m[483]&m[484])|(~m[464]&~m[480]&~m[481]&m[483]&m[484])|(m[464]&~m[480]&~m[481]&m[483]&m[484])|(~m[464]&m[480]&~m[481]&m[483]&m[484])|(m[464]&m[480]&~m[481]&m[483]&m[484])|(~m[464]&~m[480]&m[481]&m[483]&m[484])|(m[464]&~m[480]&m[481]&m[483]&m[484])|(m[464]&m[480]&m[481]&m[483]&m[484]))):InitCond[271];
    m[487] = run?((((m[469]&~m[485]&~m[486]&~m[488]&~m[489])|(~m[469]&~m[485]&~m[486]&m[488]&~m[489])|(m[469]&m[485]&~m[486]&m[488]&~m[489])|(m[469]&~m[485]&m[486]&m[488]&~m[489])|(~m[469]&m[485]&~m[486]&~m[488]&m[489])|(~m[469]&~m[485]&m[486]&~m[488]&m[489])|(m[469]&m[485]&m[486]&~m[488]&m[489])|(~m[469]&m[485]&m[486]&m[488]&m[489]))&UnbiasedRNG[113])|((m[469]&~m[485]&~m[486]&m[488]&~m[489])|(~m[469]&~m[485]&~m[486]&~m[488]&m[489])|(m[469]&~m[485]&~m[486]&~m[488]&m[489])|(m[469]&m[485]&~m[486]&~m[488]&m[489])|(m[469]&~m[485]&m[486]&~m[488]&m[489])|(~m[469]&~m[485]&~m[486]&m[488]&m[489])|(m[469]&~m[485]&~m[486]&m[488]&m[489])|(~m[469]&m[485]&~m[486]&m[488]&m[489])|(m[469]&m[485]&~m[486]&m[488]&m[489])|(~m[469]&~m[485]&m[486]&m[488]&m[489])|(m[469]&~m[485]&m[486]&m[488]&m[489])|(m[469]&m[485]&m[486]&m[488]&m[489]))):InitCond[272];
    m[492] = run?((((m[479]&~m[490]&~m[491]&~m[493]&~m[494])|(~m[479]&~m[490]&~m[491]&m[493]&~m[494])|(m[479]&m[490]&~m[491]&m[493]&~m[494])|(m[479]&~m[490]&m[491]&m[493]&~m[494])|(~m[479]&m[490]&~m[491]&~m[493]&m[494])|(~m[479]&~m[490]&m[491]&~m[493]&m[494])|(m[479]&m[490]&m[491]&~m[493]&m[494])|(~m[479]&m[490]&m[491]&m[493]&m[494]))&UnbiasedRNG[114])|((m[479]&~m[490]&~m[491]&m[493]&~m[494])|(~m[479]&~m[490]&~m[491]&~m[493]&m[494])|(m[479]&~m[490]&~m[491]&~m[493]&m[494])|(m[479]&m[490]&~m[491]&~m[493]&m[494])|(m[479]&~m[490]&m[491]&~m[493]&m[494])|(~m[479]&~m[490]&~m[491]&m[493]&m[494])|(m[479]&~m[490]&~m[491]&m[493]&m[494])|(~m[479]&m[490]&~m[491]&m[493]&m[494])|(m[479]&m[490]&~m[491]&m[493]&m[494])|(~m[479]&~m[490]&m[491]&m[493]&m[494])|(m[479]&~m[490]&m[491]&m[493]&m[494])|(m[479]&m[490]&m[491]&m[493]&m[494]))):InitCond[273];
    m[497] = run?((((m[484]&~m[495]&~m[496]&~m[498]&~m[499])|(~m[484]&~m[495]&~m[496]&m[498]&~m[499])|(m[484]&m[495]&~m[496]&m[498]&~m[499])|(m[484]&~m[495]&m[496]&m[498]&~m[499])|(~m[484]&m[495]&~m[496]&~m[498]&m[499])|(~m[484]&~m[495]&m[496]&~m[498]&m[499])|(m[484]&m[495]&m[496]&~m[498]&m[499])|(~m[484]&m[495]&m[496]&m[498]&m[499]))&UnbiasedRNG[115])|((m[484]&~m[495]&~m[496]&m[498]&~m[499])|(~m[484]&~m[495]&~m[496]&~m[498]&m[499])|(m[484]&~m[495]&~m[496]&~m[498]&m[499])|(m[484]&m[495]&~m[496]&~m[498]&m[499])|(m[484]&~m[495]&m[496]&~m[498]&m[499])|(~m[484]&~m[495]&~m[496]&m[498]&m[499])|(m[484]&~m[495]&~m[496]&m[498]&m[499])|(~m[484]&m[495]&~m[496]&m[498]&m[499])|(m[484]&m[495]&~m[496]&m[498]&m[499])|(~m[484]&~m[495]&m[496]&m[498]&m[499])|(m[484]&~m[495]&m[496]&m[498]&m[499])|(m[484]&m[495]&m[496]&m[498]&m[499]))):InitCond[274];
    m[502] = run?((((m[489]&~m[500]&~m[501]&~m[503]&~m[504])|(~m[489]&~m[500]&~m[501]&m[503]&~m[504])|(m[489]&m[500]&~m[501]&m[503]&~m[504])|(m[489]&~m[500]&m[501]&m[503]&~m[504])|(~m[489]&m[500]&~m[501]&~m[503]&m[504])|(~m[489]&~m[500]&m[501]&~m[503]&m[504])|(m[489]&m[500]&m[501]&~m[503]&m[504])|(~m[489]&m[500]&m[501]&m[503]&m[504]))&UnbiasedRNG[116])|((m[489]&~m[500]&~m[501]&m[503]&~m[504])|(~m[489]&~m[500]&~m[501]&~m[503]&m[504])|(m[489]&~m[500]&~m[501]&~m[503]&m[504])|(m[489]&m[500]&~m[501]&~m[503]&m[504])|(m[489]&~m[500]&m[501]&~m[503]&m[504])|(~m[489]&~m[500]&~m[501]&m[503]&m[504])|(m[489]&~m[500]&~m[501]&m[503]&m[504])|(~m[489]&m[500]&~m[501]&m[503]&m[504])|(m[489]&m[500]&~m[501]&m[503]&m[504])|(~m[489]&~m[500]&m[501]&m[503]&m[504])|(m[489]&~m[500]&m[501]&m[503]&m[504])|(m[489]&m[500]&m[501]&m[503]&m[504]))):InitCond[275];
    m[507] = run?((((m[499]&~m[505]&~m[506]&~m[508]&~m[509])|(~m[499]&~m[505]&~m[506]&m[508]&~m[509])|(m[499]&m[505]&~m[506]&m[508]&~m[509])|(m[499]&~m[505]&m[506]&m[508]&~m[509])|(~m[499]&m[505]&~m[506]&~m[508]&m[509])|(~m[499]&~m[505]&m[506]&~m[508]&m[509])|(m[499]&m[505]&m[506]&~m[508]&m[509])|(~m[499]&m[505]&m[506]&m[508]&m[509]))&UnbiasedRNG[117])|((m[499]&~m[505]&~m[506]&m[508]&~m[509])|(~m[499]&~m[505]&~m[506]&~m[508]&m[509])|(m[499]&~m[505]&~m[506]&~m[508]&m[509])|(m[499]&m[505]&~m[506]&~m[508]&m[509])|(m[499]&~m[505]&m[506]&~m[508]&m[509])|(~m[499]&~m[505]&~m[506]&m[508]&m[509])|(m[499]&~m[505]&~m[506]&m[508]&m[509])|(~m[499]&m[505]&~m[506]&m[508]&m[509])|(m[499]&m[505]&~m[506]&m[508]&m[509])|(~m[499]&~m[505]&m[506]&m[508]&m[509])|(m[499]&~m[505]&m[506]&m[508]&m[509])|(m[499]&m[505]&m[506]&m[508]&m[509]))):InitCond[276];
    m[512] = run?((((m[504]&~m[510]&~m[511]&~m[513]&~m[514])|(~m[504]&~m[510]&~m[511]&m[513]&~m[514])|(m[504]&m[510]&~m[511]&m[513]&~m[514])|(m[504]&~m[510]&m[511]&m[513]&~m[514])|(~m[504]&m[510]&~m[511]&~m[513]&m[514])|(~m[504]&~m[510]&m[511]&~m[513]&m[514])|(m[504]&m[510]&m[511]&~m[513]&m[514])|(~m[504]&m[510]&m[511]&m[513]&m[514]))&UnbiasedRNG[118])|((m[504]&~m[510]&~m[511]&m[513]&~m[514])|(~m[504]&~m[510]&~m[511]&~m[513]&m[514])|(m[504]&~m[510]&~m[511]&~m[513]&m[514])|(m[504]&m[510]&~m[511]&~m[513]&m[514])|(m[504]&~m[510]&m[511]&~m[513]&m[514])|(~m[504]&~m[510]&~m[511]&m[513]&m[514])|(m[504]&~m[510]&~m[511]&m[513]&m[514])|(~m[504]&m[510]&~m[511]&m[513]&m[514])|(m[504]&m[510]&~m[511]&m[513]&m[514])|(~m[504]&~m[510]&m[511]&m[513]&m[514])|(m[504]&~m[510]&m[511]&m[513]&m[514])|(m[504]&m[510]&m[511]&m[513]&m[514]))):InitCond[277];
    m[517] = run?((((m[514]&~m[515]&~m[516]&~m[518]&~m[519])|(~m[514]&~m[515]&~m[516]&m[518]&~m[519])|(m[514]&m[515]&~m[516]&m[518]&~m[519])|(m[514]&~m[515]&m[516]&m[518]&~m[519])|(~m[514]&m[515]&~m[516]&~m[518]&m[519])|(~m[514]&~m[515]&m[516]&~m[518]&m[519])|(m[514]&m[515]&m[516]&~m[518]&m[519])|(~m[514]&m[515]&m[516]&m[518]&m[519]))&UnbiasedRNG[119])|((m[514]&~m[515]&~m[516]&m[518]&~m[519])|(~m[514]&~m[515]&~m[516]&~m[518]&m[519])|(m[514]&~m[515]&~m[516]&~m[518]&m[519])|(m[514]&m[515]&~m[516]&~m[518]&m[519])|(m[514]&~m[515]&m[516]&~m[518]&m[519])|(~m[514]&~m[515]&~m[516]&m[518]&m[519])|(m[514]&~m[515]&~m[516]&m[518]&m[519])|(~m[514]&m[515]&~m[516]&m[518]&m[519])|(m[514]&m[515]&~m[516]&m[518]&m[519])|(~m[514]&~m[515]&m[516]&m[518]&m[519])|(m[514]&~m[515]&m[516]&m[518]&m[519])|(m[514]&m[515]&m[516]&m[518]&m[519]))):InitCond[278];
end

always @(posedge color2_clk) begin
    m[112] = run?((((~m[32]&~m[48]&~m[176])|(m[32]&m[48]&~m[176]))&BiasedRNG[159])|(((m[32]&~m[48]&~m[176])|(~m[32]&m[48]&m[176]))&~BiasedRNG[159])|((~m[32]&~m[48]&m[176])|(m[32]&~m[48]&m[176])|(m[32]&m[48]&m[176]))):InitCond[279];
    m[113] = run?((((~m[32]&~m[56]&~m[177])|(m[32]&m[56]&~m[177]))&BiasedRNG[160])|(((m[32]&~m[56]&~m[177])|(~m[32]&m[56]&m[177]))&~BiasedRNG[160])|((~m[32]&~m[56]&m[177])|(m[32]&~m[56]&m[177])|(m[32]&m[56]&m[177]))):InitCond[280];
    m[114] = run?((((~m[32]&~m[64]&~m[178])|(m[32]&m[64]&~m[178]))&BiasedRNG[161])|(((m[32]&~m[64]&~m[178])|(~m[32]&m[64]&m[178]))&~BiasedRNG[161])|((~m[32]&~m[64]&m[178])|(m[32]&~m[64]&m[178])|(m[32]&m[64]&m[178]))):InitCond[281];
    m[115] = run?((((~m[32]&~m[72]&~m[179])|(m[32]&m[72]&~m[179]))&BiasedRNG[162])|(((m[32]&~m[72]&~m[179])|(~m[32]&m[72]&m[179]))&~BiasedRNG[162])|((~m[32]&~m[72]&m[179])|(m[32]&~m[72]&m[179])|(m[32]&m[72]&m[179]))):InitCond[282];
    m[116] = run?((((~m[33]&~m[80]&~m[180])|(m[33]&m[80]&~m[180]))&BiasedRNG[163])|(((m[33]&~m[80]&~m[180])|(~m[33]&m[80]&m[180]))&~BiasedRNG[163])|((~m[33]&~m[80]&m[180])|(m[33]&~m[80]&m[180])|(m[33]&m[80]&m[180]))):InitCond[283];
    m[117] = run?((((~m[33]&~m[88]&~m[181])|(m[33]&m[88]&~m[181]))&BiasedRNG[164])|(((m[33]&~m[88]&~m[181])|(~m[33]&m[88]&m[181]))&~BiasedRNG[164])|((~m[33]&~m[88]&m[181])|(m[33]&~m[88]&m[181])|(m[33]&m[88]&m[181]))):InitCond[284];
    m[118] = run?((((~m[33]&~m[96]&~m[182])|(m[33]&m[96]&~m[182]))&BiasedRNG[165])|(((m[33]&~m[96]&~m[182])|(~m[33]&m[96]&m[182]))&~BiasedRNG[165])|((~m[33]&~m[96]&m[182])|(m[33]&~m[96]&m[182])|(m[33]&m[96]&m[182]))):InitCond[285];
    m[119] = run?((((~m[33]&~m[104]&~m[183])|(m[33]&m[104]&~m[183]))&BiasedRNG[166])|(((m[33]&~m[104]&~m[183])|(~m[33]&m[104]&m[183]))&~BiasedRNG[166])|((~m[33]&~m[104]&m[183])|(m[33]&~m[104]&m[183])|(m[33]&m[104]&m[183]))):InitCond[286];
    m[120] = run?((((~m[34]&~m[49]&~m[184])|(m[34]&m[49]&~m[184]))&BiasedRNG[167])|(((m[34]&~m[49]&~m[184])|(~m[34]&m[49]&m[184]))&~BiasedRNG[167])|((~m[34]&~m[49]&m[184])|(m[34]&~m[49]&m[184])|(m[34]&m[49]&m[184]))):InitCond[287];
    m[121] = run?((((~m[34]&~m[57]&~m[185])|(m[34]&m[57]&~m[185]))&BiasedRNG[168])|(((m[34]&~m[57]&~m[185])|(~m[34]&m[57]&m[185]))&~BiasedRNG[168])|((~m[34]&~m[57]&m[185])|(m[34]&~m[57]&m[185])|(m[34]&m[57]&m[185]))):InitCond[288];
    m[122] = run?((((~m[34]&~m[65]&~m[186])|(m[34]&m[65]&~m[186]))&BiasedRNG[169])|(((m[34]&~m[65]&~m[186])|(~m[34]&m[65]&m[186]))&~BiasedRNG[169])|((~m[34]&~m[65]&m[186])|(m[34]&~m[65]&m[186])|(m[34]&m[65]&m[186]))):InitCond[289];
    m[123] = run?((((~m[34]&~m[73]&~m[187])|(m[34]&m[73]&~m[187]))&BiasedRNG[170])|(((m[34]&~m[73]&~m[187])|(~m[34]&m[73]&m[187]))&~BiasedRNG[170])|((~m[34]&~m[73]&m[187])|(m[34]&~m[73]&m[187])|(m[34]&m[73]&m[187]))):InitCond[290];
    m[124] = run?((((~m[35]&~m[81]&~m[188])|(m[35]&m[81]&~m[188]))&BiasedRNG[171])|(((m[35]&~m[81]&~m[188])|(~m[35]&m[81]&m[188]))&~BiasedRNG[171])|((~m[35]&~m[81]&m[188])|(m[35]&~m[81]&m[188])|(m[35]&m[81]&m[188]))):InitCond[291];
    m[125] = run?((((~m[35]&~m[89]&~m[189])|(m[35]&m[89]&~m[189]))&BiasedRNG[172])|(((m[35]&~m[89]&~m[189])|(~m[35]&m[89]&m[189]))&~BiasedRNG[172])|((~m[35]&~m[89]&m[189])|(m[35]&~m[89]&m[189])|(m[35]&m[89]&m[189]))):InitCond[292];
    m[126] = run?((((~m[35]&~m[97]&~m[190])|(m[35]&m[97]&~m[190]))&BiasedRNG[173])|(((m[35]&~m[97]&~m[190])|(~m[35]&m[97]&m[190]))&~BiasedRNG[173])|((~m[35]&~m[97]&m[190])|(m[35]&~m[97]&m[190])|(m[35]&m[97]&m[190]))):InitCond[293];
    m[127] = run?((((~m[35]&~m[105]&~m[191])|(m[35]&m[105]&~m[191]))&BiasedRNG[174])|(((m[35]&~m[105]&~m[191])|(~m[35]&m[105]&m[191]))&~BiasedRNG[174])|((~m[35]&~m[105]&m[191])|(m[35]&~m[105]&m[191])|(m[35]&m[105]&m[191]))):InitCond[294];
    m[128] = run?((((~m[36]&~m[50]&~m[192])|(m[36]&m[50]&~m[192]))&BiasedRNG[175])|(((m[36]&~m[50]&~m[192])|(~m[36]&m[50]&m[192]))&~BiasedRNG[175])|((~m[36]&~m[50]&m[192])|(m[36]&~m[50]&m[192])|(m[36]&m[50]&m[192]))):InitCond[295];
    m[129] = run?((((~m[36]&~m[58]&~m[193])|(m[36]&m[58]&~m[193]))&BiasedRNG[176])|(((m[36]&~m[58]&~m[193])|(~m[36]&m[58]&m[193]))&~BiasedRNG[176])|((~m[36]&~m[58]&m[193])|(m[36]&~m[58]&m[193])|(m[36]&m[58]&m[193]))):InitCond[296];
    m[130] = run?((((~m[36]&~m[66]&~m[194])|(m[36]&m[66]&~m[194]))&BiasedRNG[177])|(((m[36]&~m[66]&~m[194])|(~m[36]&m[66]&m[194]))&~BiasedRNG[177])|((~m[36]&~m[66]&m[194])|(m[36]&~m[66]&m[194])|(m[36]&m[66]&m[194]))):InitCond[297];
    m[131] = run?((((~m[36]&~m[74]&~m[195])|(m[36]&m[74]&~m[195]))&BiasedRNG[178])|(((m[36]&~m[74]&~m[195])|(~m[36]&m[74]&m[195]))&~BiasedRNG[178])|((~m[36]&~m[74]&m[195])|(m[36]&~m[74]&m[195])|(m[36]&m[74]&m[195]))):InitCond[298];
    m[132] = run?((((~m[37]&~m[82]&~m[196])|(m[37]&m[82]&~m[196]))&BiasedRNG[179])|(((m[37]&~m[82]&~m[196])|(~m[37]&m[82]&m[196]))&~BiasedRNG[179])|((~m[37]&~m[82]&m[196])|(m[37]&~m[82]&m[196])|(m[37]&m[82]&m[196]))):InitCond[299];
    m[133] = run?((((~m[37]&~m[90]&~m[197])|(m[37]&m[90]&~m[197]))&BiasedRNG[180])|(((m[37]&~m[90]&~m[197])|(~m[37]&m[90]&m[197]))&~BiasedRNG[180])|((~m[37]&~m[90]&m[197])|(m[37]&~m[90]&m[197])|(m[37]&m[90]&m[197]))):InitCond[300];
    m[134] = run?((((~m[37]&~m[98]&~m[198])|(m[37]&m[98]&~m[198]))&BiasedRNG[181])|(((m[37]&~m[98]&~m[198])|(~m[37]&m[98]&m[198]))&~BiasedRNG[181])|((~m[37]&~m[98]&m[198])|(m[37]&~m[98]&m[198])|(m[37]&m[98]&m[198]))):InitCond[301];
    m[135] = run?((((~m[37]&~m[106]&~m[199])|(m[37]&m[106]&~m[199]))&BiasedRNG[182])|(((m[37]&~m[106]&~m[199])|(~m[37]&m[106]&m[199]))&~BiasedRNG[182])|((~m[37]&~m[106]&m[199])|(m[37]&~m[106]&m[199])|(m[37]&m[106]&m[199]))):InitCond[302];
    m[136] = run?((((~m[38]&~m[51]&~m[200])|(m[38]&m[51]&~m[200]))&BiasedRNG[183])|(((m[38]&~m[51]&~m[200])|(~m[38]&m[51]&m[200]))&~BiasedRNG[183])|((~m[38]&~m[51]&m[200])|(m[38]&~m[51]&m[200])|(m[38]&m[51]&m[200]))):InitCond[303];
    m[137] = run?((((~m[38]&~m[59]&~m[201])|(m[38]&m[59]&~m[201]))&BiasedRNG[184])|(((m[38]&~m[59]&~m[201])|(~m[38]&m[59]&m[201]))&~BiasedRNG[184])|((~m[38]&~m[59]&m[201])|(m[38]&~m[59]&m[201])|(m[38]&m[59]&m[201]))):InitCond[304];
    m[138] = run?((((~m[38]&~m[67]&~m[202])|(m[38]&m[67]&~m[202]))&BiasedRNG[185])|(((m[38]&~m[67]&~m[202])|(~m[38]&m[67]&m[202]))&~BiasedRNG[185])|((~m[38]&~m[67]&m[202])|(m[38]&~m[67]&m[202])|(m[38]&m[67]&m[202]))):InitCond[305];
    m[139] = run?((((~m[38]&~m[75]&~m[203])|(m[38]&m[75]&~m[203]))&BiasedRNG[186])|(((m[38]&~m[75]&~m[203])|(~m[38]&m[75]&m[203]))&~BiasedRNG[186])|((~m[38]&~m[75]&m[203])|(m[38]&~m[75]&m[203])|(m[38]&m[75]&m[203]))):InitCond[306];
    m[140] = run?((((~m[39]&~m[83]&~m[204])|(m[39]&m[83]&~m[204]))&BiasedRNG[187])|(((m[39]&~m[83]&~m[204])|(~m[39]&m[83]&m[204]))&~BiasedRNG[187])|((~m[39]&~m[83]&m[204])|(m[39]&~m[83]&m[204])|(m[39]&m[83]&m[204]))):InitCond[307];
    m[141] = run?((((~m[39]&~m[91]&~m[205])|(m[39]&m[91]&~m[205]))&BiasedRNG[188])|(((m[39]&~m[91]&~m[205])|(~m[39]&m[91]&m[205]))&~BiasedRNG[188])|((~m[39]&~m[91]&m[205])|(m[39]&~m[91]&m[205])|(m[39]&m[91]&m[205]))):InitCond[308];
    m[142] = run?((((~m[39]&~m[99]&~m[206])|(m[39]&m[99]&~m[206]))&BiasedRNG[189])|(((m[39]&~m[99]&~m[206])|(~m[39]&m[99]&m[206]))&~BiasedRNG[189])|((~m[39]&~m[99]&m[206])|(m[39]&~m[99]&m[206])|(m[39]&m[99]&m[206]))):InitCond[309];
    m[143] = run?((((~m[39]&~m[107]&~m[207])|(m[39]&m[107]&~m[207]))&BiasedRNG[190])|(((m[39]&~m[107]&~m[207])|(~m[39]&m[107]&m[207]))&~BiasedRNG[190])|((~m[39]&~m[107]&m[207])|(m[39]&~m[107]&m[207])|(m[39]&m[107]&m[207]))):InitCond[310];
    m[144] = run?((((~m[40]&~m[52]&~m[208])|(m[40]&m[52]&~m[208]))&BiasedRNG[191])|(((m[40]&~m[52]&~m[208])|(~m[40]&m[52]&m[208]))&~BiasedRNG[191])|((~m[40]&~m[52]&m[208])|(m[40]&~m[52]&m[208])|(m[40]&m[52]&m[208]))):InitCond[311];
    m[145] = run?((((~m[40]&~m[60]&~m[209])|(m[40]&m[60]&~m[209]))&BiasedRNG[192])|(((m[40]&~m[60]&~m[209])|(~m[40]&m[60]&m[209]))&~BiasedRNG[192])|((~m[40]&~m[60]&m[209])|(m[40]&~m[60]&m[209])|(m[40]&m[60]&m[209]))):InitCond[312];
    m[146] = run?((((~m[40]&~m[68]&~m[210])|(m[40]&m[68]&~m[210]))&BiasedRNG[193])|(((m[40]&~m[68]&~m[210])|(~m[40]&m[68]&m[210]))&~BiasedRNG[193])|((~m[40]&~m[68]&m[210])|(m[40]&~m[68]&m[210])|(m[40]&m[68]&m[210]))):InitCond[313];
    m[147] = run?((((~m[40]&~m[76]&~m[211])|(m[40]&m[76]&~m[211]))&BiasedRNG[194])|(((m[40]&~m[76]&~m[211])|(~m[40]&m[76]&m[211]))&~BiasedRNG[194])|((~m[40]&~m[76]&m[211])|(m[40]&~m[76]&m[211])|(m[40]&m[76]&m[211]))):InitCond[314];
    m[148] = run?((((~m[41]&~m[84]&~m[212])|(m[41]&m[84]&~m[212]))&BiasedRNG[195])|(((m[41]&~m[84]&~m[212])|(~m[41]&m[84]&m[212]))&~BiasedRNG[195])|((~m[41]&~m[84]&m[212])|(m[41]&~m[84]&m[212])|(m[41]&m[84]&m[212]))):InitCond[315];
    m[149] = run?((((~m[41]&~m[92]&~m[213])|(m[41]&m[92]&~m[213]))&BiasedRNG[196])|(((m[41]&~m[92]&~m[213])|(~m[41]&m[92]&m[213]))&~BiasedRNG[196])|((~m[41]&~m[92]&m[213])|(m[41]&~m[92]&m[213])|(m[41]&m[92]&m[213]))):InitCond[316];
    m[150] = run?((((~m[41]&~m[100]&~m[214])|(m[41]&m[100]&~m[214]))&BiasedRNG[197])|(((m[41]&~m[100]&~m[214])|(~m[41]&m[100]&m[214]))&~BiasedRNG[197])|((~m[41]&~m[100]&m[214])|(m[41]&~m[100]&m[214])|(m[41]&m[100]&m[214]))):InitCond[317];
    m[151] = run?((((~m[41]&~m[108]&~m[215])|(m[41]&m[108]&~m[215]))&BiasedRNG[198])|(((m[41]&~m[108]&~m[215])|(~m[41]&m[108]&m[215]))&~BiasedRNG[198])|((~m[41]&~m[108]&m[215])|(m[41]&~m[108]&m[215])|(m[41]&m[108]&m[215]))):InitCond[318];
    m[152] = run?((((~m[42]&~m[53]&~m[216])|(m[42]&m[53]&~m[216]))&BiasedRNG[199])|(((m[42]&~m[53]&~m[216])|(~m[42]&m[53]&m[216]))&~BiasedRNG[199])|((~m[42]&~m[53]&m[216])|(m[42]&~m[53]&m[216])|(m[42]&m[53]&m[216]))):InitCond[319];
    m[153] = run?((((~m[42]&~m[61]&~m[217])|(m[42]&m[61]&~m[217]))&BiasedRNG[200])|(((m[42]&~m[61]&~m[217])|(~m[42]&m[61]&m[217]))&~BiasedRNG[200])|((~m[42]&~m[61]&m[217])|(m[42]&~m[61]&m[217])|(m[42]&m[61]&m[217]))):InitCond[320];
    m[154] = run?((((~m[42]&~m[69]&~m[218])|(m[42]&m[69]&~m[218]))&BiasedRNG[201])|(((m[42]&~m[69]&~m[218])|(~m[42]&m[69]&m[218]))&~BiasedRNG[201])|((~m[42]&~m[69]&m[218])|(m[42]&~m[69]&m[218])|(m[42]&m[69]&m[218]))):InitCond[321];
    m[155] = run?((((~m[42]&~m[77]&~m[219])|(m[42]&m[77]&~m[219]))&BiasedRNG[202])|(((m[42]&~m[77]&~m[219])|(~m[42]&m[77]&m[219]))&~BiasedRNG[202])|((~m[42]&~m[77]&m[219])|(m[42]&~m[77]&m[219])|(m[42]&m[77]&m[219]))):InitCond[322];
    m[156] = run?((((~m[43]&~m[85]&~m[220])|(m[43]&m[85]&~m[220]))&BiasedRNG[203])|(((m[43]&~m[85]&~m[220])|(~m[43]&m[85]&m[220]))&~BiasedRNG[203])|((~m[43]&~m[85]&m[220])|(m[43]&~m[85]&m[220])|(m[43]&m[85]&m[220]))):InitCond[323];
    m[157] = run?((((~m[43]&~m[93]&~m[221])|(m[43]&m[93]&~m[221]))&BiasedRNG[204])|(((m[43]&~m[93]&~m[221])|(~m[43]&m[93]&m[221]))&~BiasedRNG[204])|((~m[43]&~m[93]&m[221])|(m[43]&~m[93]&m[221])|(m[43]&m[93]&m[221]))):InitCond[324];
    m[158] = run?((((~m[43]&~m[101]&~m[222])|(m[43]&m[101]&~m[222]))&BiasedRNG[205])|(((m[43]&~m[101]&~m[222])|(~m[43]&m[101]&m[222]))&~BiasedRNG[205])|((~m[43]&~m[101]&m[222])|(m[43]&~m[101]&m[222])|(m[43]&m[101]&m[222]))):InitCond[325];
    m[159] = run?((((~m[43]&~m[109]&~m[223])|(m[43]&m[109]&~m[223]))&BiasedRNG[206])|(((m[43]&~m[109]&~m[223])|(~m[43]&m[109]&m[223]))&~BiasedRNG[206])|((~m[43]&~m[109]&m[223])|(m[43]&~m[109]&m[223])|(m[43]&m[109]&m[223]))):InitCond[326];
    m[160] = run?((((~m[44]&~m[54]&~m[224])|(m[44]&m[54]&~m[224]))&BiasedRNG[207])|(((m[44]&~m[54]&~m[224])|(~m[44]&m[54]&m[224]))&~BiasedRNG[207])|((~m[44]&~m[54]&m[224])|(m[44]&~m[54]&m[224])|(m[44]&m[54]&m[224]))):InitCond[327];
    m[161] = run?((((~m[44]&~m[62]&~m[225])|(m[44]&m[62]&~m[225]))&BiasedRNG[208])|(((m[44]&~m[62]&~m[225])|(~m[44]&m[62]&m[225]))&~BiasedRNG[208])|((~m[44]&~m[62]&m[225])|(m[44]&~m[62]&m[225])|(m[44]&m[62]&m[225]))):InitCond[328];
    m[162] = run?((((~m[44]&~m[70]&~m[226])|(m[44]&m[70]&~m[226]))&BiasedRNG[209])|(((m[44]&~m[70]&~m[226])|(~m[44]&m[70]&m[226]))&~BiasedRNG[209])|((~m[44]&~m[70]&m[226])|(m[44]&~m[70]&m[226])|(m[44]&m[70]&m[226]))):InitCond[329];
    m[163] = run?((((~m[44]&~m[78]&~m[227])|(m[44]&m[78]&~m[227]))&BiasedRNG[210])|(((m[44]&~m[78]&~m[227])|(~m[44]&m[78]&m[227]))&~BiasedRNG[210])|((~m[44]&~m[78]&m[227])|(m[44]&~m[78]&m[227])|(m[44]&m[78]&m[227]))):InitCond[330];
    m[164] = run?((((~m[45]&~m[86]&~m[228])|(m[45]&m[86]&~m[228]))&BiasedRNG[211])|(((m[45]&~m[86]&~m[228])|(~m[45]&m[86]&m[228]))&~BiasedRNG[211])|((~m[45]&~m[86]&m[228])|(m[45]&~m[86]&m[228])|(m[45]&m[86]&m[228]))):InitCond[331];
    m[165] = run?((((~m[45]&~m[94]&~m[229])|(m[45]&m[94]&~m[229]))&BiasedRNG[212])|(((m[45]&~m[94]&~m[229])|(~m[45]&m[94]&m[229]))&~BiasedRNG[212])|((~m[45]&~m[94]&m[229])|(m[45]&~m[94]&m[229])|(m[45]&m[94]&m[229]))):InitCond[332];
    m[166] = run?((((~m[45]&~m[102]&~m[230])|(m[45]&m[102]&~m[230]))&BiasedRNG[213])|(((m[45]&~m[102]&~m[230])|(~m[45]&m[102]&m[230]))&~BiasedRNG[213])|((~m[45]&~m[102]&m[230])|(m[45]&~m[102]&m[230])|(m[45]&m[102]&m[230]))):InitCond[333];
    m[167] = run?((((~m[45]&~m[110]&~m[231])|(m[45]&m[110]&~m[231]))&BiasedRNG[214])|(((m[45]&~m[110]&~m[231])|(~m[45]&m[110]&m[231]))&~BiasedRNG[214])|((~m[45]&~m[110]&m[231])|(m[45]&~m[110]&m[231])|(m[45]&m[110]&m[231]))):InitCond[334];
    m[168] = run?((((~m[46]&~m[55]&~m[232])|(m[46]&m[55]&~m[232]))&BiasedRNG[215])|(((m[46]&~m[55]&~m[232])|(~m[46]&m[55]&m[232]))&~BiasedRNG[215])|((~m[46]&~m[55]&m[232])|(m[46]&~m[55]&m[232])|(m[46]&m[55]&m[232]))):InitCond[335];
    m[169] = run?((((~m[46]&~m[63]&~m[233])|(m[46]&m[63]&~m[233]))&BiasedRNG[216])|(((m[46]&~m[63]&~m[233])|(~m[46]&m[63]&m[233]))&~BiasedRNG[216])|((~m[46]&~m[63]&m[233])|(m[46]&~m[63]&m[233])|(m[46]&m[63]&m[233]))):InitCond[336];
    m[170] = run?((((~m[46]&~m[71]&~m[234])|(m[46]&m[71]&~m[234]))&BiasedRNG[217])|(((m[46]&~m[71]&~m[234])|(~m[46]&m[71]&m[234]))&~BiasedRNG[217])|((~m[46]&~m[71]&m[234])|(m[46]&~m[71]&m[234])|(m[46]&m[71]&m[234]))):InitCond[337];
    m[171] = run?((((~m[46]&~m[79]&~m[235])|(m[46]&m[79]&~m[235]))&BiasedRNG[218])|(((m[46]&~m[79]&~m[235])|(~m[46]&m[79]&m[235]))&~BiasedRNG[218])|((~m[46]&~m[79]&m[235])|(m[46]&~m[79]&m[235])|(m[46]&m[79]&m[235]))):InitCond[338];
    m[172] = run?((((~m[47]&~m[87]&~m[236])|(m[47]&m[87]&~m[236]))&BiasedRNG[219])|(((m[47]&~m[87]&~m[236])|(~m[47]&m[87]&m[236]))&~BiasedRNG[219])|((~m[47]&~m[87]&m[236])|(m[47]&~m[87]&m[236])|(m[47]&m[87]&m[236]))):InitCond[339];
    m[173] = run?((((~m[47]&~m[95]&~m[237])|(m[47]&m[95]&~m[237]))&BiasedRNG[220])|(((m[47]&~m[95]&~m[237])|(~m[47]&m[95]&m[237]))&~BiasedRNG[220])|((~m[47]&~m[95]&m[237])|(m[47]&~m[95]&m[237])|(m[47]&m[95]&m[237]))):InitCond[340];
    m[174] = run?((((~m[47]&~m[103]&~m[238])|(m[47]&m[103]&~m[238]))&BiasedRNG[221])|(((m[47]&~m[103]&~m[238])|(~m[47]&m[103]&m[238]))&~BiasedRNG[221])|((~m[47]&~m[103]&m[238])|(m[47]&~m[103]&m[238])|(m[47]&m[103]&m[238]))):InitCond[341];
    m[175] = run?((((~m[47]&~m[111]&~m[239])|(m[47]&m[111]&~m[239]))&BiasedRNG[222])|(((m[47]&~m[111]&~m[239])|(~m[47]&m[111]&m[239]))&~BiasedRNG[222])|((~m[47]&~m[111]&m[239])|(m[47]&~m[111]&m[239])|(m[47]&m[111]&m[239]))):InitCond[342];
    m[241] = run?((((m[184]&~m[240]&~m[242]&~m[243]&~m[244])|(~m[184]&~m[240]&~m[242]&m[243]&~m[244])|(m[184]&m[240]&~m[242]&m[243]&~m[244])|(m[184]&~m[240]&m[242]&m[243]&~m[244])|(~m[184]&m[240]&~m[242]&~m[243]&m[244])|(~m[184]&~m[240]&m[242]&~m[243]&m[244])|(m[184]&m[240]&m[242]&~m[243]&m[244])|(~m[184]&m[240]&m[242]&m[243]&m[244]))&UnbiasedRNG[120])|((m[184]&~m[240]&~m[242]&m[243]&~m[244])|(~m[184]&~m[240]&~m[242]&~m[243]&m[244])|(m[184]&~m[240]&~m[242]&~m[243]&m[244])|(m[184]&m[240]&~m[242]&~m[243]&m[244])|(m[184]&~m[240]&m[242]&~m[243]&m[244])|(~m[184]&~m[240]&~m[242]&m[243]&m[244])|(m[184]&~m[240]&~m[242]&m[243]&m[244])|(~m[184]&m[240]&~m[242]&m[243]&m[244])|(m[184]&m[240]&~m[242]&m[243]&m[244])|(~m[184]&~m[240]&m[242]&m[243]&m[244])|(m[184]&~m[240]&m[242]&m[243]&m[244])|(m[184]&m[240]&m[242]&m[243]&m[244]))):InitCond[343];
    m[246] = run?((((m[185]&~m[245]&~m[247]&~m[248]&~m[249])|(~m[185]&~m[245]&~m[247]&m[248]&~m[249])|(m[185]&m[245]&~m[247]&m[248]&~m[249])|(m[185]&~m[245]&m[247]&m[248]&~m[249])|(~m[185]&m[245]&~m[247]&~m[248]&m[249])|(~m[185]&~m[245]&m[247]&~m[248]&m[249])|(m[185]&m[245]&m[247]&~m[248]&m[249])|(~m[185]&m[245]&m[247]&m[248]&m[249]))&UnbiasedRNG[121])|((m[185]&~m[245]&~m[247]&m[248]&~m[249])|(~m[185]&~m[245]&~m[247]&~m[248]&m[249])|(m[185]&~m[245]&~m[247]&~m[248]&m[249])|(m[185]&m[245]&~m[247]&~m[248]&m[249])|(m[185]&~m[245]&m[247]&~m[248]&m[249])|(~m[185]&~m[245]&~m[247]&m[248]&m[249])|(m[185]&~m[245]&~m[247]&m[248]&m[249])|(~m[185]&m[245]&~m[247]&m[248]&m[249])|(m[185]&m[245]&~m[247]&m[248]&m[249])|(~m[185]&~m[245]&m[247]&m[248]&m[249])|(m[185]&~m[245]&m[247]&m[248]&m[249])|(m[185]&m[245]&m[247]&m[248]&m[249]))):InitCond[344];
    m[251] = run?((((m[192]&~m[250]&~m[252]&~m[253]&~m[254])|(~m[192]&~m[250]&~m[252]&m[253]&~m[254])|(m[192]&m[250]&~m[252]&m[253]&~m[254])|(m[192]&~m[250]&m[252]&m[253]&~m[254])|(~m[192]&m[250]&~m[252]&~m[253]&m[254])|(~m[192]&~m[250]&m[252]&~m[253]&m[254])|(m[192]&m[250]&m[252]&~m[253]&m[254])|(~m[192]&m[250]&m[252]&m[253]&m[254]))&UnbiasedRNG[122])|((m[192]&~m[250]&~m[252]&m[253]&~m[254])|(~m[192]&~m[250]&~m[252]&~m[253]&m[254])|(m[192]&~m[250]&~m[252]&~m[253]&m[254])|(m[192]&m[250]&~m[252]&~m[253]&m[254])|(m[192]&~m[250]&m[252]&~m[253]&m[254])|(~m[192]&~m[250]&~m[252]&m[253]&m[254])|(m[192]&~m[250]&~m[252]&m[253]&m[254])|(~m[192]&m[250]&~m[252]&m[253]&m[254])|(m[192]&m[250]&~m[252]&m[253]&m[254])|(~m[192]&~m[250]&m[252]&m[253]&m[254])|(m[192]&~m[250]&m[252]&m[253]&m[254])|(m[192]&m[250]&m[252]&m[253]&m[254]))):InitCond[345];
    m[256] = run?((((m[186]&~m[255]&~m[257]&~m[258]&~m[259])|(~m[186]&~m[255]&~m[257]&m[258]&~m[259])|(m[186]&m[255]&~m[257]&m[258]&~m[259])|(m[186]&~m[255]&m[257]&m[258]&~m[259])|(~m[186]&m[255]&~m[257]&~m[258]&m[259])|(~m[186]&~m[255]&m[257]&~m[258]&m[259])|(m[186]&m[255]&m[257]&~m[258]&m[259])|(~m[186]&m[255]&m[257]&m[258]&m[259]))&UnbiasedRNG[123])|((m[186]&~m[255]&~m[257]&m[258]&~m[259])|(~m[186]&~m[255]&~m[257]&~m[258]&m[259])|(m[186]&~m[255]&~m[257]&~m[258]&m[259])|(m[186]&m[255]&~m[257]&~m[258]&m[259])|(m[186]&~m[255]&m[257]&~m[258]&m[259])|(~m[186]&~m[255]&~m[257]&m[258]&m[259])|(m[186]&~m[255]&~m[257]&m[258]&m[259])|(~m[186]&m[255]&~m[257]&m[258]&m[259])|(m[186]&m[255]&~m[257]&m[258]&m[259])|(~m[186]&~m[255]&m[257]&m[258]&m[259])|(m[186]&~m[255]&m[257]&m[258]&m[259])|(m[186]&m[255]&m[257]&m[258]&m[259]))):InitCond[346];
    m[261] = run?((((m[193]&~m[260]&~m[262]&~m[263]&~m[264])|(~m[193]&~m[260]&~m[262]&m[263]&~m[264])|(m[193]&m[260]&~m[262]&m[263]&~m[264])|(m[193]&~m[260]&m[262]&m[263]&~m[264])|(~m[193]&m[260]&~m[262]&~m[263]&m[264])|(~m[193]&~m[260]&m[262]&~m[263]&m[264])|(m[193]&m[260]&m[262]&~m[263]&m[264])|(~m[193]&m[260]&m[262]&m[263]&m[264]))&UnbiasedRNG[124])|((m[193]&~m[260]&~m[262]&m[263]&~m[264])|(~m[193]&~m[260]&~m[262]&~m[263]&m[264])|(m[193]&~m[260]&~m[262]&~m[263]&m[264])|(m[193]&m[260]&~m[262]&~m[263]&m[264])|(m[193]&~m[260]&m[262]&~m[263]&m[264])|(~m[193]&~m[260]&~m[262]&m[263]&m[264])|(m[193]&~m[260]&~m[262]&m[263]&m[264])|(~m[193]&m[260]&~m[262]&m[263]&m[264])|(m[193]&m[260]&~m[262]&m[263]&m[264])|(~m[193]&~m[260]&m[262]&m[263]&m[264])|(m[193]&~m[260]&m[262]&m[263]&m[264])|(m[193]&m[260]&m[262]&m[263]&m[264]))):InitCond[347];
    m[266] = run?((((m[200]&~m[265]&~m[267]&~m[268]&~m[269])|(~m[200]&~m[265]&~m[267]&m[268]&~m[269])|(m[200]&m[265]&~m[267]&m[268]&~m[269])|(m[200]&~m[265]&m[267]&m[268]&~m[269])|(~m[200]&m[265]&~m[267]&~m[268]&m[269])|(~m[200]&~m[265]&m[267]&~m[268]&m[269])|(m[200]&m[265]&m[267]&~m[268]&m[269])|(~m[200]&m[265]&m[267]&m[268]&m[269]))&UnbiasedRNG[125])|((m[200]&~m[265]&~m[267]&m[268]&~m[269])|(~m[200]&~m[265]&~m[267]&~m[268]&m[269])|(m[200]&~m[265]&~m[267]&~m[268]&m[269])|(m[200]&m[265]&~m[267]&~m[268]&m[269])|(m[200]&~m[265]&m[267]&~m[268]&m[269])|(~m[200]&~m[265]&~m[267]&m[268]&m[269])|(m[200]&~m[265]&~m[267]&m[268]&m[269])|(~m[200]&m[265]&~m[267]&m[268]&m[269])|(m[200]&m[265]&~m[267]&m[268]&m[269])|(~m[200]&~m[265]&m[267]&m[268]&m[269])|(m[200]&~m[265]&m[267]&m[268]&m[269])|(m[200]&m[265]&m[267]&m[268]&m[269]))):InitCond[348];
    m[271] = run?((((m[187]&~m[270]&~m[272]&~m[273]&~m[274])|(~m[187]&~m[270]&~m[272]&m[273]&~m[274])|(m[187]&m[270]&~m[272]&m[273]&~m[274])|(m[187]&~m[270]&m[272]&m[273]&~m[274])|(~m[187]&m[270]&~m[272]&~m[273]&m[274])|(~m[187]&~m[270]&m[272]&~m[273]&m[274])|(m[187]&m[270]&m[272]&~m[273]&m[274])|(~m[187]&m[270]&m[272]&m[273]&m[274]))&UnbiasedRNG[126])|((m[187]&~m[270]&~m[272]&m[273]&~m[274])|(~m[187]&~m[270]&~m[272]&~m[273]&m[274])|(m[187]&~m[270]&~m[272]&~m[273]&m[274])|(m[187]&m[270]&~m[272]&~m[273]&m[274])|(m[187]&~m[270]&m[272]&~m[273]&m[274])|(~m[187]&~m[270]&~m[272]&m[273]&m[274])|(m[187]&~m[270]&~m[272]&m[273]&m[274])|(~m[187]&m[270]&~m[272]&m[273]&m[274])|(m[187]&m[270]&~m[272]&m[273]&m[274])|(~m[187]&~m[270]&m[272]&m[273]&m[274])|(m[187]&~m[270]&m[272]&m[273]&m[274])|(m[187]&m[270]&m[272]&m[273]&m[274]))):InitCond[349];
    m[276] = run?((((m[194]&~m[275]&~m[277]&~m[278]&~m[279])|(~m[194]&~m[275]&~m[277]&m[278]&~m[279])|(m[194]&m[275]&~m[277]&m[278]&~m[279])|(m[194]&~m[275]&m[277]&m[278]&~m[279])|(~m[194]&m[275]&~m[277]&~m[278]&m[279])|(~m[194]&~m[275]&m[277]&~m[278]&m[279])|(m[194]&m[275]&m[277]&~m[278]&m[279])|(~m[194]&m[275]&m[277]&m[278]&m[279]))&UnbiasedRNG[127])|((m[194]&~m[275]&~m[277]&m[278]&~m[279])|(~m[194]&~m[275]&~m[277]&~m[278]&m[279])|(m[194]&~m[275]&~m[277]&~m[278]&m[279])|(m[194]&m[275]&~m[277]&~m[278]&m[279])|(m[194]&~m[275]&m[277]&~m[278]&m[279])|(~m[194]&~m[275]&~m[277]&m[278]&m[279])|(m[194]&~m[275]&~m[277]&m[278]&m[279])|(~m[194]&m[275]&~m[277]&m[278]&m[279])|(m[194]&m[275]&~m[277]&m[278]&m[279])|(~m[194]&~m[275]&m[277]&m[278]&m[279])|(m[194]&~m[275]&m[277]&m[278]&m[279])|(m[194]&m[275]&m[277]&m[278]&m[279]))):InitCond[350];
    m[281] = run?((((m[201]&~m[280]&~m[282]&~m[283]&~m[284])|(~m[201]&~m[280]&~m[282]&m[283]&~m[284])|(m[201]&m[280]&~m[282]&m[283]&~m[284])|(m[201]&~m[280]&m[282]&m[283]&~m[284])|(~m[201]&m[280]&~m[282]&~m[283]&m[284])|(~m[201]&~m[280]&m[282]&~m[283]&m[284])|(m[201]&m[280]&m[282]&~m[283]&m[284])|(~m[201]&m[280]&m[282]&m[283]&m[284]))&UnbiasedRNG[128])|((m[201]&~m[280]&~m[282]&m[283]&~m[284])|(~m[201]&~m[280]&~m[282]&~m[283]&m[284])|(m[201]&~m[280]&~m[282]&~m[283]&m[284])|(m[201]&m[280]&~m[282]&~m[283]&m[284])|(m[201]&~m[280]&m[282]&~m[283]&m[284])|(~m[201]&~m[280]&~m[282]&m[283]&m[284])|(m[201]&~m[280]&~m[282]&m[283]&m[284])|(~m[201]&m[280]&~m[282]&m[283]&m[284])|(m[201]&m[280]&~m[282]&m[283]&m[284])|(~m[201]&~m[280]&m[282]&m[283]&m[284])|(m[201]&~m[280]&m[282]&m[283]&m[284])|(m[201]&m[280]&m[282]&m[283]&m[284]))):InitCond[351];
    m[286] = run?((((m[208]&~m[285]&~m[287]&~m[288]&~m[289])|(~m[208]&~m[285]&~m[287]&m[288]&~m[289])|(m[208]&m[285]&~m[287]&m[288]&~m[289])|(m[208]&~m[285]&m[287]&m[288]&~m[289])|(~m[208]&m[285]&~m[287]&~m[288]&m[289])|(~m[208]&~m[285]&m[287]&~m[288]&m[289])|(m[208]&m[285]&m[287]&~m[288]&m[289])|(~m[208]&m[285]&m[287]&m[288]&m[289]))&UnbiasedRNG[129])|((m[208]&~m[285]&~m[287]&m[288]&~m[289])|(~m[208]&~m[285]&~m[287]&~m[288]&m[289])|(m[208]&~m[285]&~m[287]&~m[288]&m[289])|(m[208]&m[285]&~m[287]&~m[288]&m[289])|(m[208]&~m[285]&m[287]&~m[288]&m[289])|(~m[208]&~m[285]&~m[287]&m[288]&m[289])|(m[208]&~m[285]&~m[287]&m[288]&m[289])|(~m[208]&m[285]&~m[287]&m[288]&m[289])|(m[208]&m[285]&~m[287]&m[288]&m[289])|(~m[208]&~m[285]&m[287]&m[288]&m[289])|(m[208]&~m[285]&m[287]&m[288]&m[289])|(m[208]&m[285]&m[287]&m[288]&m[289]))):InitCond[352];
    m[291] = run?((((m[188]&~m[290]&~m[292]&~m[293]&~m[294])|(~m[188]&~m[290]&~m[292]&m[293]&~m[294])|(m[188]&m[290]&~m[292]&m[293]&~m[294])|(m[188]&~m[290]&m[292]&m[293]&~m[294])|(~m[188]&m[290]&~m[292]&~m[293]&m[294])|(~m[188]&~m[290]&m[292]&~m[293]&m[294])|(m[188]&m[290]&m[292]&~m[293]&m[294])|(~m[188]&m[290]&m[292]&m[293]&m[294]))&UnbiasedRNG[130])|((m[188]&~m[290]&~m[292]&m[293]&~m[294])|(~m[188]&~m[290]&~m[292]&~m[293]&m[294])|(m[188]&~m[290]&~m[292]&~m[293]&m[294])|(m[188]&m[290]&~m[292]&~m[293]&m[294])|(m[188]&~m[290]&m[292]&~m[293]&m[294])|(~m[188]&~m[290]&~m[292]&m[293]&m[294])|(m[188]&~m[290]&~m[292]&m[293]&m[294])|(~m[188]&m[290]&~m[292]&m[293]&m[294])|(m[188]&m[290]&~m[292]&m[293]&m[294])|(~m[188]&~m[290]&m[292]&m[293]&m[294])|(m[188]&~m[290]&m[292]&m[293]&m[294])|(m[188]&m[290]&m[292]&m[293]&m[294]))):InitCond[353];
    m[296] = run?((((m[195]&~m[295]&~m[297]&~m[298]&~m[299])|(~m[195]&~m[295]&~m[297]&m[298]&~m[299])|(m[195]&m[295]&~m[297]&m[298]&~m[299])|(m[195]&~m[295]&m[297]&m[298]&~m[299])|(~m[195]&m[295]&~m[297]&~m[298]&m[299])|(~m[195]&~m[295]&m[297]&~m[298]&m[299])|(m[195]&m[295]&m[297]&~m[298]&m[299])|(~m[195]&m[295]&m[297]&m[298]&m[299]))&UnbiasedRNG[131])|((m[195]&~m[295]&~m[297]&m[298]&~m[299])|(~m[195]&~m[295]&~m[297]&~m[298]&m[299])|(m[195]&~m[295]&~m[297]&~m[298]&m[299])|(m[195]&m[295]&~m[297]&~m[298]&m[299])|(m[195]&~m[295]&m[297]&~m[298]&m[299])|(~m[195]&~m[295]&~m[297]&m[298]&m[299])|(m[195]&~m[295]&~m[297]&m[298]&m[299])|(~m[195]&m[295]&~m[297]&m[298]&m[299])|(m[195]&m[295]&~m[297]&m[298]&m[299])|(~m[195]&~m[295]&m[297]&m[298]&m[299])|(m[195]&~m[295]&m[297]&m[298]&m[299])|(m[195]&m[295]&m[297]&m[298]&m[299]))):InitCond[354];
    m[301] = run?((((m[202]&~m[300]&~m[302]&~m[303]&~m[304])|(~m[202]&~m[300]&~m[302]&m[303]&~m[304])|(m[202]&m[300]&~m[302]&m[303]&~m[304])|(m[202]&~m[300]&m[302]&m[303]&~m[304])|(~m[202]&m[300]&~m[302]&~m[303]&m[304])|(~m[202]&~m[300]&m[302]&~m[303]&m[304])|(m[202]&m[300]&m[302]&~m[303]&m[304])|(~m[202]&m[300]&m[302]&m[303]&m[304]))&UnbiasedRNG[132])|((m[202]&~m[300]&~m[302]&m[303]&~m[304])|(~m[202]&~m[300]&~m[302]&~m[303]&m[304])|(m[202]&~m[300]&~m[302]&~m[303]&m[304])|(m[202]&m[300]&~m[302]&~m[303]&m[304])|(m[202]&~m[300]&m[302]&~m[303]&m[304])|(~m[202]&~m[300]&~m[302]&m[303]&m[304])|(m[202]&~m[300]&~m[302]&m[303]&m[304])|(~m[202]&m[300]&~m[302]&m[303]&m[304])|(m[202]&m[300]&~m[302]&m[303]&m[304])|(~m[202]&~m[300]&m[302]&m[303]&m[304])|(m[202]&~m[300]&m[302]&m[303]&m[304])|(m[202]&m[300]&m[302]&m[303]&m[304]))):InitCond[355];
    m[306] = run?((((m[209]&~m[305]&~m[307]&~m[308]&~m[309])|(~m[209]&~m[305]&~m[307]&m[308]&~m[309])|(m[209]&m[305]&~m[307]&m[308]&~m[309])|(m[209]&~m[305]&m[307]&m[308]&~m[309])|(~m[209]&m[305]&~m[307]&~m[308]&m[309])|(~m[209]&~m[305]&m[307]&~m[308]&m[309])|(m[209]&m[305]&m[307]&~m[308]&m[309])|(~m[209]&m[305]&m[307]&m[308]&m[309]))&UnbiasedRNG[133])|((m[209]&~m[305]&~m[307]&m[308]&~m[309])|(~m[209]&~m[305]&~m[307]&~m[308]&m[309])|(m[209]&~m[305]&~m[307]&~m[308]&m[309])|(m[209]&m[305]&~m[307]&~m[308]&m[309])|(m[209]&~m[305]&m[307]&~m[308]&m[309])|(~m[209]&~m[305]&~m[307]&m[308]&m[309])|(m[209]&~m[305]&~m[307]&m[308]&m[309])|(~m[209]&m[305]&~m[307]&m[308]&m[309])|(m[209]&m[305]&~m[307]&m[308]&m[309])|(~m[209]&~m[305]&m[307]&m[308]&m[309])|(m[209]&~m[305]&m[307]&m[308]&m[309])|(m[209]&m[305]&m[307]&m[308]&m[309]))):InitCond[356];
    m[311] = run?((((m[216]&~m[310]&~m[312]&~m[313]&~m[314])|(~m[216]&~m[310]&~m[312]&m[313]&~m[314])|(m[216]&m[310]&~m[312]&m[313]&~m[314])|(m[216]&~m[310]&m[312]&m[313]&~m[314])|(~m[216]&m[310]&~m[312]&~m[313]&m[314])|(~m[216]&~m[310]&m[312]&~m[313]&m[314])|(m[216]&m[310]&m[312]&~m[313]&m[314])|(~m[216]&m[310]&m[312]&m[313]&m[314]))&UnbiasedRNG[134])|((m[216]&~m[310]&~m[312]&m[313]&~m[314])|(~m[216]&~m[310]&~m[312]&~m[313]&m[314])|(m[216]&~m[310]&~m[312]&~m[313]&m[314])|(m[216]&m[310]&~m[312]&~m[313]&m[314])|(m[216]&~m[310]&m[312]&~m[313]&m[314])|(~m[216]&~m[310]&~m[312]&m[313]&m[314])|(m[216]&~m[310]&~m[312]&m[313]&m[314])|(~m[216]&m[310]&~m[312]&m[313]&m[314])|(m[216]&m[310]&~m[312]&m[313]&m[314])|(~m[216]&~m[310]&m[312]&m[313]&m[314])|(m[216]&~m[310]&m[312]&m[313]&m[314])|(m[216]&m[310]&m[312]&m[313]&m[314]))):InitCond[357];
    m[316] = run?((((m[189]&~m[315]&~m[317]&~m[318]&~m[319])|(~m[189]&~m[315]&~m[317]&m[318]&~m[319])|(m[189]&m[315]&~m[317]&m[318]&~m[319])|(m[189]&~m[315]&m[317]&m[318]&~m[319])|(~m[189]&m[315]&~m[317]&~m[318]&m[319])|(~m[189]&~m[315]&m[317]&~m[318]&m[319])|(m[189]&m[315]&m[317]&~m[318]&m[319])|(~m[189]&m[315]&m[317]&m[318]&m[319]))&UnbiasedRNG[135])|((m[189]&~m[315]&~m[317]&m[318]&~m[319])|(~m[189]&~m[315]&~m[317]&~m[318]&m[319])|(m[189]&~m[315]&~m[317]&~m[318]&m[319])|(m[189]&m[315]&~m[317]&~m[318]&m[319])|(m[189]&~m[315]&m[317]&~m[318]&m[319])|(~m[189]&~m[315]&~m[317]&m[318]&m[319])|(m[189]&~m[315]&~m[317]&m[318]&m[319])|(~m[189]&m[315]&~m[317]&m[318]&m[319])|(m[189]&m[315]&~m[317]&m[318]&m[319])|(~m[189]&~m[315]&m[317]&m[318]&m[319])|(m[189]&~m[315]&m[317]&m[318]&m[319])|(m[189]&m[315]&m[317]&m[318]&m[319]))):InitCond[358];
    m[321] = run?((((m[196]&~m[320]&~m[322]&~m[323]&~m[324])|(~m[196]&~m[320]&~m[322]&m[323]&~m[324])|(m[196]&m[320]&~m[322]&m[323]&~m[324])|(m[196]&~m[320]&m[322]&m[323]&~m[324])|(~m[196]&m[320]&~m[322]&~m[323]&m[324])|(~m[196]&~m[320]&m[322]&~m[323]&m[324])|(m[196]&m[320]&m[322]&~m[323]&m[324])|(~m[196]&m[320]&m[322]&m[323]&m[324]))&UnbiasedRNG[136])|((m[196]&~m[320]&~m[322]&m[323]&~m[324])|(~m[196]&~m[320]&~m[322]&~m[323]&m[324])|(m[196]&~m[320]&~m[322]&~m[323]&m[324])|(m[196]&m[320]&~m[322]&~m[323]&m[324])|(m[196]&~m[320]&m[322]&~m[323]&m[324])|(~m[196]&~m[320]&~m[322]&m[323]&m[324])|(m[196]&~m[320]&~m[322]&m[323]&m[324])|(~m[196]&m[320]&~m[322]&m[323]&m[324])|(m[196]&m[320]&~m[322]&m[323]&m[324])|(~m[196]&~m[320]&m[322]&m[323]&m[324])|(m[196]&~m[320]&m[322]&m[323]&m[324])|(m[196]&m[320]&m[322]&m[323]&m[324]))):InitCond[359];
    m[326] = run?((((m[203]&~m[325]&~m[327]&~m[328]&~m[329])|(~m[203]&~m[325]&~m[327]&m[328]&~m[329])|(m[203]&m[325]&~m[327]&m[328]&~m[329])|(m[203]&~m[325]&m[327]&m[328]&~m[329])|(~m[203]&m[325]&~m[327]&~m[328]&m[329])|(~m[203]&~m[325]&m[327]&~m[328]&m[329])|(m[203]&m[325]&m[327]&~m[328]&m[329])|(~m[203]&m[325]&m[327]&m[328]&m[329]))&UnbiasedRNG[137])|((m[203]&~m[325]&~m[327]&m[328]&~m[329])|(~m[203]&~m[325]&~m[327]&~m[328]&m[329])|(m[203]&~m[325]&~m[327]&~m[328]&m[329])|(m[203]&m[325]&~m[327]&~m[328]&m[329])|(m[203]&~m[325]&m[327]&~m[328]&m[329])|(~m[203]&~m[325]&~m[327]&m[328]&m[329])|(m[203]&~m[325]&~m[327]&m[328]&m[329])|(~m[203]&m[325]&~m[327]&m[328]&m[329])|(m[203]&m[325]&~m[327]&m[328]&m[329])|(~m[203]&~m[325]&m[327]&m[328]&m[329])|(m[203]&~m[325]&m[327]&m[328]&m[329])|(m[203]&m[325]&m[327]&m[328]&m[329]))):InitCond[360];
    m[331] = run?((((m[210]&~m[330]&~m[332]&~m[333]&~m[334])|(~m[210]&~m[330]&~m[332]&m[333]&~m[334])|(m[210]&m[330]&~m[332]&m[333]&~m[334])|(m[210]&~m[330]&m[332]&m[333]&~m[334])|(~m[210]&m[330]&~m[332]&~m[333]&m[334])|(~m[210]&~m[330]&m[332]&~m[333]&m[334])|(m[210]&m[330]&m[332]&~m[333]&m[334])|(~m[210]&m[330]&m[332]&m[333]&m[334]))&UnbiasedRNG[138])|((m[210]&~m[330]&~m[332]&m[333]&~m[334])|(~m[210]&~m[330]&~m[332]&~m[333]&m[334])|(m[210]&~m[330]&~m[332]&~m[333]&m[334])|(m[210]&m[330]&~m[332]&~m[333]&m[334])|(m[210]&~m[330]&m[332]&~m[333]&m[334])|(~m[210]&~m[330]&~m[332]&m[333]&m[334])|(m[210]&~m[330]&~m[332]&m[333]&m[334])|(~m[210]&m[330]&~m[332]&m[333]&m[334])|(m[210]&m[330]&~m[332]&m[333]&m[334])|(~m[210]&~m[330]&m[332]&m[333]&m[334])|(m[210]&~m[330]&m[332]&m[333]&m[334])|(m[210]&m[330]&m[332]&m[333]&m[334]))):InitCond[361];
    m[336] = run?((((m[217]&~m[335]&~m[337]&~m[338]&~m[339])|(~m[217]&~m[335]&~m[337]&m[338]&~m[339])|(m[217]&m[335]&~m[337]&m[338]&~m[339])|(m[217]&~m[335]&m[337]&m[338]&~m[339])|(~m[217]&m[335]&~m[337]&~m[338]&m[339])|(~m[217]&~m[335]&m[337]&~m[338]&m[339])|(m[217]&m[335]&m[337]&~m[338]&m[339])|(~m[217]&m[335]&m[337]&m[338]&m[339]))&UnbiasedRNG[139])|((m[217]&~m[335]&~m[337]&m[338]&~m[339])|(~m[217]&~m[335]&~m[337]&~m[338]&m[339])|(m[217]&~m[335]&~m[337]&~m[338]&m[339])|(m[217]&m[335]&~m[337]&~m[338]&m[339])|(m[217]&~m[335]&m[337]&~m[338]&m[339])|(~m[217]&~m[335]&~m[337]&m[338]&m[339])|(m[217]&~m[335]&~m[337]&m[338]&m[339])|(~m[217]&m[335]&~m[337]&m[338]&m[339])|(m[217]&m[335]&~m[337]&m[338]&m[339])|(~m[217]&~m[335]&m[337]&m[338]&m[339])|(m[217]&~m[335]&m[337]&m[338]&m[339])|(m[217]&m[335]&m[337]&m[338]&m[339]))):InitCond[362];
    m[341] = run?((((m[224]&~m[340]&~m[342]&~m[343]&~m[344])|(~m[224]&~m[340]&~m[342]&m[343]&~m[344])|(m[224]&m[340]&~m[342]&m[343]&~m[344])|(m[224]&~m[340]&m[342]&m[343]&~m[344])|(~m[224]&m[340]&~m[342]&~m[343]&m[344])|(~m[224]&~m[340]&m[342]&~m[343]&m[344])|(m[224]&m[340]&m[342]&~m[343]&m[344])|(~m[224]&m[340]&m[342]&m[343]&m[344]))&UnbiasedRNG[140])|((m[224]&~m[340]&~m[342]&m[343]&~m[344])|(~m[224]&~m[340]&~m[342]&~m[343]&m[344])|(m[224]&~m[340]&~m[342]&~m[343]&m[344])|(m[224]&m[340]&~m[342]&~m[343]&m[344])|(m[224]&~m[340]&m[342]&~m[343]&m[344])|(~m[224]&~m[340]&~m[342]&m[343]&m[344])|(m[224]&~m[340]&~m[342]&m[343]&m[344])|(~m[224]&m[340]&~m[342]&m[343]&m[344])|(m[224]&m[340]&~m[342]&m[343]&m[344])|(~m[224]&~m[340]&m[342]&m[343]&m[344])|(m[224]&~m[340]&m[342]&m[343]&m[344])|(m[224]&m[340]&m[342]&m[343]&m[344]))):InitCond[363];
    m[346] = run?((((m[190]&~m[345]&~m[347]&~m[348]&~m[349])|(~m[190]&~m[345]&~m[347]&m[348]&~m[349])|(m[190]&m[345]&~m[347]&m[348]&~m[349])|(m[190]&~m[345]&m[347]&m[348]&~m[349])|(~m[190]&m[345]&~m[347]&~m[348]&m[349])|(~m[190]&~m[345]&m[347]&~m[348]&m[349])|(m[190]&m[345]&m[347]&~m[348]&m[349])|(~m[190]&m[345]&m[347]&m[348]&m[349]))&UnbiasedRNG[141])|((m[190]&~m[345]&~m[347]&m[348]&~m[349])|(~m[190]&~m[345]&~m[347]&~m[348]&m[349])|(m[190]&~m[345]&~m[347]&~m[348]&m[349])|(m[190]&m[345]&~m[347]&~m[348]&m[349])|(m[190]&~m[345]&m[347]&~m[348]&m[349])|(~m[190]&~m[345]&~m[347]&m[348]&m[349])|(m[190]&~m[345]&~m[347]&m[348]&m[349])|(~m[190]&m[345]&~m[347]&m[348]&m[349])|(m[190]&m[345]&~m[347]&m[348]&m[349])|(~m[190]&~m[345]&m[347]&m[348]&m[349])|(m[190]&~m[345]&m[347]&m[348]&m[349])|(m[190]&m[345]&m[347]&m[348]&m[349]))):InitCond[364];
    m[351] = run?((((m[197]&~m[350]&~m[352]&~m[353]&~m[354])|(~m[197]&~m[350]&~m[352]&m[353]&~m[354])|(m[197]&m[350]&~m[352]&m[353]&~m[354])|(m[197]&~m[350]&m[352]&m[353]&~m[354])|(~m[197]&m[350]&~m[352]&~m[353]&m[354])|(~m[197]&~m[350]&m[352]&~m[353]&m[354])|(m[197]&m[350]&m[352]&~m[353]&m[354])|(~m[197]&m[350]&m[352]&m[353]&m[354]))&UnbiasedRNG[142])|((m[197]&~m[350]&~m[352]&m[353]&~m[354])|(~m[197]&~m[350]&~m[352]&~m[353]&m[354])|(m[197]&~m[350]&~m[352]&~m[353]&m[354])|(m[197]&m[350]&~m[352]&~m[353]&m[354])|(m[197]&~m[350]&m[352]&~m[353]&m[354])|(~m[197]&~m[350]&~m[352]&m[353]&m[354])|(m[197]&~m[350]&~m[352]&m[353]&m[354])|(~m[197]&m[350]&~m[352]&m[353]&m[354])|(m[197]&m[350]&~m[352]&m[353]&m[354])|(~m[197]&~m[350]&m[352]&m[353]&m[354])|(m[197]&~m[350]&m[352]&m[353]&m[354])|(m[197]&m[350]&m[352]&m[353]&m[354]))):InitCond[365];
    m[356] = run?((((m[204]&~m[355]&~m[357]&~m[358]&~m[359])|(~m[204]&~m[355]&~m[357]&m[358]&~m[359])|(m[204]&m[355]&~m[357]&m[358]&~m[359])|(m[204]&~m[355]&m[357]&m[358]&~m[359])|(~m[204]&m[355]&~m[357]&~m[358]&m[359])|(~m[204]&~m[355]&m[357]&~m[358]&m[359])|(m[204]&m[355]&m[357]&~m[358]&m[359])|(~m[204]&m[355]&m[357]&m[358]&m[359]))&UnbiasedRNG[143])|((m[204]&~m[355]&~m[357]&m[358]&~m[359])|(~m[204]&~m[355]&~m[357]&~m[358]&m[359])|(m[204]&~m[355]&~m[357]&~m[358]&m[359])|(m[204]&m[355]&~m[357]&~m[358]&m[359])|(m[204]&~m[355]&m[357]&~m[358]&m[359])|(~m[204]&~m[355]&~m[357]&m[358]&m[359])|(m[204]&~m[355]&~m[357]&m[358]&m[359])|(~m[204]&m[355]&~m[357]&m[358]&m[359])|(m[204]&m[355]&~m[357]&m[358]&m[359])|(~m[204]&~m[355]&m[357]&m[358]&m[359])|(m[204]&~m[355]&m[357]&m[358]&m[359])|(m[204]&m[355]&m[357]&m[358]&m[359]))):InitCond[366];
    m[361] = run?((((m[211]&~m[360]&~m[362]&~m[363]&~m[364])|(~m[211]&~m[360]&~m[362]&m[363]&~m[364])|(m[211]&m[360]&~m[362]&m[363]&~m[364])|(m[211]&~m[360]&m[362]&m[363]&~m[364])|(~m[211]&m[360]&~m[362]&~m[363]&m[364])|(~m[211]&~m[360]&m[362]&~m[363]&m[364])|(m[211]&m[360]&m[362]&~m[363]&m[364])|(~m[211]&m[360]&m[362]&m[363]&m[364]))&UnbiasedRNG[144])|((m[211]&~m[360]&~m[362]&m[363]&~m[364])|(~m[211]&~m[360]&~m[362]&~m[363]&m[364])|(m[211]&~m[360]&~m[362]&~m[363]&m[364])|(m[211]&m[360]&~m[362]&~m[363]&m[364])|(m[211]&~m[360]&m[362]&~m[363]&m[364])|(~m[211]&~m[360]&~m[362]&m[363]&m[364])|(m[211]&~m[360]&~m[362]&m[363]&m[364])|(~m[211]&m[360]&~m[362]&m[363]&m[364])|(m[211]&m[360]&~m[362]&m[363]&m[364])|(~m[211]&~m[360]&m[362]&m[363]&m[364])|(m[211]&~m[360]&m[362]&m[363]&m[364])|(m[211]&m[360]&m[362]&m[363]&m[364]))):InitCond[367];
    m[366] = run?((((m[218]&~m[365]&~m[367]&~m[368]&~m[369])|(~m[218]&~m[365]&~m[367]&m[368]&~m[369])|(m[218]&m[365]&~m[367]&m[368]&~m[369])|(m[218]&~m[365]&m[367]&m[368]&~m[369])|(~m[218]&m[365]&~m[367]&~m[368]&m[369])|(~m[218]&~m[365]&m[367]&~m[368]&m[369])|(m[218]&m[365]&m[367]&~m[368]&m[369])|(~m[218]&m[365]&m[367]&m[368]&m[369]))&UnbiasedRNG[145])|((m[218]&~m[365]&~m[367]&m[368]&~m[369])|(~m[218]&~m[365]&~m[367]&~m[368]&m[369])|(m[218]&~m[365]&~m[367]&~m[368]&m[369])|(m[218]&m[365]&~m[367]&~m[368]&m[369])|(m[218]&~m[365]&m[367]&~m[368]&m[369])|(~m[218]&~m[365]&~m[367]&m[368]&m[369])|(m[218]&~m[365]&~m[367]&m[368]&m[369])|(~m[218]&m[365]&~m[367]&m[368]&m[369])|(m[218]&m[365]&~m[367]&m[368]&m[369])|(~m[218]&~m[365]&m[367]&m[368]&m[369])|(m[218]&~m[365]&m[367]&m[368]&m[369])|(m[218]&m[365]&m[367]&m[368]&m[369]))):InitCond[368];
    m[371] = run?((((m[225]&~m[370]&~m[372]&~m[373]&~m[374])|(~m[225]&~m[370]&~m[372]&m[373]&~m[374])|(m[225]&m[370]&~m[372]&m[373]&~m[374])|(m[225]&~m[370]&m[372]&m[373]&~m[374])|(~m[225]&m[370]&~m[372]&~m[373]&m[374])|(~m[225]&~m[370]&m[372]&~m[373]&m[374])|(m[225]&m[370]&m[372]&~m[373]&m[374])|(~m[225]&m[370]&m[372]&m[373]&m[374]))&UnbiasedRNG[146])|((m[225]&~m[370]&~m[372]&m[373]&~m[374])|(~m[225]&~m[370]&~m[372]&~m[373]&m[374])|(m[225]&~m[370]&~m[372]&~m[373]&m[374])|(m[225]&m[370]&~m[372]&~m[373]&m[374])|(m[225]&~m[370]&m[372]&~m[373]&m[374])|(~m[225]&~m[370]&~m[372]&m[373]&m[374])|(m[225]&~m[370]&~m[372]&m[373]&m[374])|(~m[225]&m[370]&~m[372]&m[373]&m[374])|(m[225]&m[370]&~m[372]&m[373]&m[374])|(~m[225]&~m[370]&m[372]&m[373]&m[374])|(m[225]&~m[370]&m[372]&m[373]&m[374])|(m[225]&m[370]&m[372]&m[373]&m[374]))):InitCond[369];
    m[376] = run?((((m[232]&~m[375]&~m[377]&~m[378]&~m[379])|(~m[232]&~m[375]&~m[377]&m[378]&~m[379])|(m[232]&m[375]&~m[377]&m[378]&~m[379])|(m[232]&~m[375]&m[377]&m[378]&~m[379])|(~m[232]&m[375]&~m[377]&~m[378]&m[379])|(~m[232]&~m[375]&m[377]&~m[378]&m[379])|(m[232]&m[375]&m[377]&~m[378]&m[379])|(~m[232]&m[375]&m[377]&m[378]&m[379]))&UnbiasedRNG[147])|((m[232]&~m[375]&~m[377]&m[378]&~m[379])|(~m[232]&~m[375]&~m[377]&~m[378]&m[379])|(m[232]&~m[375]&~m[377]&~m[378]&m[379])|(m[232]&m[375]&~m[377]&~m[378]&m[379])|(m[232]&~m[375]&m[377]&~m[378]&m[379])|(~m[232]&~m[375]&~m[377]&m[378]&m[379])|(m[232]&~m[375]&~m[377]&m[378]&m[379])|(~m[232]&m[375]&~m[377]&m[378]&m[379])|(m[232]&m[375]&~m[377]&m[378]&m[379])|(~m[232]&~m[375]&m[377]&m[378]&m[379])|(m[232]&~m[375]&m[377]&m[378]&m[379])|(m[232]&m[375]&m[377]&m[378]&m[379]))):InitCond[370];
    m[381] = run?((((m[191]&~m[380]&~m[382]&~m[383]&~m[384])|(~m[191]&~m[380]&~m[382]&m[383]&~m[384])|(m[191]&m[380]&~m[382]&m[383]&~m[384])|(m[191]&~m[380]&m[382]&m[383]&~m[384])|(~m[191]&m[380]&~m[382]&~m[383]&m[384])|(~m[191]&~m[380]&m[382]&~m[383]&m[384])|(m[191]&m[380]&m[382]&~m[383]&m[384])|(~m[191]&m[380]&m[382]&m[383]&m[384]))&UnbiasedRNG[148])|((m[191]&~m[380]&~m[382]&m[383]&~m[384])|(~m[191]&~m[380]&~m[382]&~m[383]&m[384])|(m[191]&~m[380]&~m[382]&~m[383]&m[384])|(m[191]&m[380]&~m[382]&~m[383]&m[384])|(m[191]&~m[380]&m[382]&~m[383]&m[384])|(~m[191]&~m[380]&~m[382]&m[383]&m[384])|(m[191]&~m[380]&~m[382]&m[383]&m[384])|(~m[191]&m[380]&~m[382]&m[383]&m[384])|(m[191]&m[380]&~m[382]&m[383]&m[384])|(~m[191]&~m[380]&m[382]&m[383]&m[384])|(m[191]&~m[380]&m[382]&m[383]&m[384])|(m[191]&m[380]&m[382]&m[383]&m[384]))):InitCond[371];
    m[386] = run?((((m[198]&~m[385]&~m[387]&~m[388]&~m[389])|(~m[198]&~m[385]&~m[387]&m[388]&~m[389])|(m[198]&m[385]&~m[387]&m[388]&~m[389])|(m[198]&~m[385]&m[387]&m[388]&~m[389])|(~m[198]&m[385]&~m[387]&~m[388]&m[389])|(~m[198]&~m[385]&m[387]&~m[388]&m[389])|(m[198]&m[385]&m[387]&~m[388]&m[389])|(~m[198]&m[385]&m[387]&m[388]&m[389]))&UnbiasedRNG[149])|((m[198]&~m[385]&~m[387]&m[388]&~m[389])|(~m[198]&~m[385]&~m[387]&~m[388]&m[389])|(m[198]&~m[385]&~m[387]&~m[388]&m[389])|(m[198]&m[385]&~m[387]&~m[388]&m[389])|(m[198]&~m[385]&m[387]&~m[388]&m[389])|(~m[198]&~m[385]&~m[387]&m[388]&m[389])|(m[198]&~m[385]&~m[387]&m[388]&m[389])|(~m[198]&m[385]&~m[387]&m[388]&m[389])|(m[198]&m[385]&~m[387]&m[388]&m[389])|(~m[198]&~m[385]&m[387]&m[388]&m[389])|(m[198]&~m[385]&m[387]&m[388]&m[389])|(m[198]&m[385]&m[387]&m[388]&m[389]))):InitCond[372];
    m[391] = run?((((m[205]&~m[390]&~m[392]&~m[393]&~m[394])|(~m[205]&~m[390]&~m[392]&m[393]&~m[394])|(m[205]&m[390]&~m[392]&m[393]&~m[394])|(m[205]&~m[390]&m[392]&m[393]&~m[394])|(~m[205]&m[390]&~m[392]&~m[393]&m[394])|(~m[205]&~m[390]&m[392]&~m[393]&m[394])|(m[205]&m[390]&m[392]&~m[393]&m[394])|(~m[205]&m[390]&m[392]&m[393]&m[394]))&UnbiasedRNG[150])|((m[205]&~m[390]&~m[392]&m[393]&~m[394])|(~m[205]&~m[390]&~m[392]&~m[393]&m[394])|(m[205]&~m[390]&~m[392]&~m[393]&m[394])|(m[205]&m[390]&~m[392]&~m[393]&m[394])|(m[205]&~m[390]&m[392]&~m[393]&m[394])|(~m[205]&~m[390]&~m[392]&m[393]&m[394])|(m[205]&~m[390]&~m[392]&m[393]&m[394])|(~m[205]&m[390]&~m[392]&m[393]&m[394])|(m[205]&m[390]&~m[392]&m[393]&m[394])|(~m[205]&~m[390]&m[392]&m[393]&m[394])|(m[205]&~m[390]&m[392]&m[393]&m[394])|(m[205]&m[390]&m[392]&m[393]&m[394]))):InitCond[373];
    m[396] = run?((((m[212]&~m[395]&~m[397]&~m[398]&~m[399])|(~m[212]&~m[395]&~m[397]&m[398]&~m[399])|(m[212]&m[395]&~m[397]&m[398]&~m[399])|(m[212]&~m[395]&m[397]&m[398]&~m[399])|(~m[212]&m[395]&~m[397]&~m[398]&m[399])|(~m[212]&~m[395]&m[397]&~m[398]&m[399])|(m[212]&m[395]&m[397]&~m[398]&m[399])|(~m[212]&m[395]&m[397]&m[398]&m[399]))&UnbiasedRNG[151])|((m[212]&~m[395]&~m[397]&m[398]&~m[399])|(~m[212]&~m[395]&~m[397]&~m[398]&m[399])|(m[212]&~m[395]&~m[397]&~m[398]&m[399])|(m[212]&m[395]&~m[397]&~m[398]&m[399])|(m[212]&~m[395]&m[397]&~m[398]&m[399])|(~m[212]&~m[395]&~m[397]&m[398]&m[399])|(m[212]&~m[395]&~m[397]&m[398]&m[399])|(~m[212]&m[395]&~m[397]&m[398]&m[399])|(m[212]&m[395]&~m[397]&m[398]&m[399])|(~m[212]&~m[395]&m[397]&m[398]&m[399])|(m[212]&~m[395]&m[397]&m[398]&m[399])|(m[212]&m[395]&m[397]&m[398]&m[399]))):InitCond[374];
    m[401] = run?((((m[219]&~m[400]&~m[402]&~m[403]&~m[404])|(~m[219]&~m[400]&~m[402]&m[403]&~m[404])|(m[219]&m[400]&~m[402]&m[403]&~m[404])|(m[219]&~m[400]&m[402]&m[403]&~m[404])|(~m[219]&m[400]&~m[402]&~m[403]&m[404])|(~m[219]&~m[400]&m[402]&~m[403]&m[404])|(m[219]&m[400]&m[402]&~m[403]&m[404])|(~m[219]&m[400]&m[402]&m[403]&m[404]))&UnbiasedRNG[152])|((m[219]&~m[400]&~m[402]&m[403]&~m[404])|(~m[219]&~m[400]&~m[402]&~m[403]&m[404])|(m[219]&~m[400]&~m[402]&~m[403]&m[404])|(m[219]&m[400]&~m[402]&~m[403]&m[404])|(m[219]&~m[400]&m[402]&~m[403]&m[404])|(~m[219]&~m[400]&~m[402]&m[403]&m[404])|(m[219]&~m[400]&~m[402]&m[403]&m[404])|(~m[219]&m[400]&~m[402]&m[403]&m[404])|(m[219]&m[400]&~m[402]&m[403]&m[404])|(~m[219]&~m[400]&m[402]&m[403]&m[404])|(m[219]&~m[400]&m[402]&m[403]&m[404])|(m[219]&m[400]&m[402]&m[403]&m[404]))):InitCond[375];
    m[406] = run?((((m[226]&~m[405]&~m[407]&~m[408]&~m[409])|(~m[226]&~m[405]&~m[407]&m[408]&~m[409])|(m[226]&m[405]&~m[407]&m[408]&~m[409])|(m[226]&~m[405]&m[407]&m[408]&~m[409])|(~m[226]&m[405]&~m[407]&~m[408]&m[409])|(~m[226]&~m[405]&m[407]&~m[408]&m[409])|(m[226]&m[405]&m[407]&~m[408]&m[409])|(~m[226]&m[405]&m[407]&m[408]&m[409]))&UnbiasedRNG[153])|((m[226]&~m[405]&~m[407]&m[408]&~m[409])|(~m[226]&~m[405]&~m[407]&~m[408]&m[409])|(m[226]&~m[405]&~m[407]&~m[408]&m[409])|(m[226]&m[405]&~m[407]&~m[408]&m[409])|(m[226]&~m[405]&m[407]&~m[408]&m[409])|(~m[226]&~m[405]&~m[407]&m[408]&m[409])|(m[226]&~m[405]&~m[407]&m[408]&m[409])|(~m[226]&m[405]&~m[407]&m[408]&m[409])|(m[226]&m[405]&~m[407]&m[408]&m[409])|(~m[226]&~m[405]&m[407]&m[408]&m[409])|(m[226]&~m[405]&m[407]&m[408]&m[409])|(m[226]&m[405]&m[407]&m[408]&m[409]))):InitCond[376];
    m[411] = run?((((m[233]&~m[410]&~m[412]&~m[413]&~m[414])|(~m[233]&~m[410]&~m[412]&m[413]&~m[414])|(m[233]&m[410]&~m[412]&m[413]&~m[414])|(m[233]&~m[410]&m[412]&m[413]&~m[414])|(~m[233]&m[410]&~m[412]&~m[413]&m[414])|(~m[233]&~m[410]&m[412]&~m[413]&m[414])|(m[233]&m[410]&m[412]&~m[413]&m[414])|(~m[233]&m[410]&m[412]&m[413]&m[414]))&UnbiasedRNG[154])|((m[233]&~m[410]&~m[412]&m[413]&~m[414])|(~m[233]&~m[410]&~m[412]&~m[413]&m[414])|(m[233]&~m[410]&~m[412]&~m[413]&m[414])|(m[233]&m[410]&~m[412]&~m[413]&m[414])|(m[233]&~m[410]&m[412]&~m[413]&m[414])|(~m[233]&~m[410]&~m[412]&m[413]&m[414])|(m[233]&~m[410]&~m[412]&m[413]&m[414])|(~m[233]&m[410]&~m[412]&m[413]&m[414])|(m[233]&m[410]&~m[412]&m[413]&m[414])|(~m[233]&~m[410]&m[412]&m[413]&m[414])|(m[233]&~m[410]&m[412]&m[413]&m[414])|(m[233]&m[410]&m[412]&m[413]&m[414]))):InitCond[377];
    m[416] = run?((((m[199]&~m[415]&~m[417]&~m[418]&~m[419])|(~m[199]&~m[415]&~m[417]&m[418]&~m[419])|(m[199]&m[415]&~m[417]&m[418]&~m[419])|(m[199]&~m[415]&m[417]&m[418]&~m[419])|(~m[199]&m[415]&~m[417]&~m[418]&m[419])|(~m[199]&~m[415]&m[417]&~m[418]&m[419])|(m[199]&m[415]&m[417]&~m[418]&m[419])|(~m[199]&m[415]&m[417]&m[418]&m[419]))&UnbiasedRNG[155])|((m[199]&~m[415]&~m[417]&m[418]&~m[419])|(~m[199]&~m[415]&~m[417]&~m[418]&m[419])|(m[199]&~m[415]&~m[417]&~m[418]&m[419])|(m[199]&m[415]&~m[417]&~m[418]&m[419])|(m[199]&~m[415]&m[417]&~m[418]&m[419])|(~m[199]&~m[415]&~m[417]&m[418]&m[419])|(m[199]&~m[415]&~m[417]&m[418]&m[419])|(~m[199]&m[415]&~m[417]&m[418]&m[419])|(m[199]&m[415]&~m[417]&m[418]&m[419])|(~m[199]&~m[415]&m[417]&m[418]&m[419])|(m[199]&~m[415]&m[417]&m[418]&m[419])|(m[199]&m[415]&m[417]&m[418]&m[419]))):InitCond[378];
    m[421] = run?((((m[206]&~m[420]&~m[422]&~m[423]&~m[424])|(~m[206]&~m[420]&~m[422]&m[423]&~m[424])|(m[206]&m[420]&~m[422]&m[423]&~m[424])|(m[206]&~m[420]&m[422]&m[423]&~m[424])|(~m[206]&m[420]&~m[422]&~m[423]&m[424])|(~m[206]&~m[420]&m[422]&~m[423]&m[424])|(m[206]&m[420]&m[422]&~m[423]&m[424])|(~m[206]&m[420]&m[422]&m[423]&m[424]))&UnbiasedRNG[156])|((m[206]&~m[420]&~m[422]&m[423]&~m[424])|(~m[206]&~m[420]&~m[422]&~m[423]&m[424])|(m[206]&~m[420]&~m[422]&~m[423]&m[424])|(m[206]&m[420]&~m[422]&~m[423]&m[424])|(m[206]&~m[420]&m[422]&~m[423]&m[424])|(~m[206]&~m[420]&~m[422]&m[423]&m[424])|(m[206]&~m[420]&~m[422]&m[423]&m[424])|(~m[206]&m[420]&~m[422]&m[423]&m[424])|(m[206]&m[420]&~m[422]&m[423]&m[424])|(~m[206]&~m[420]&m[422]&m[423]&m[424])|(m[206]&~m[420]&m[422]&m[423]&m[424])|(m[206]&m[420]&m[422]&m[423]&m[424]))):InitCond[379];
    m[426] = run?((((m[213]&~m[425]&~m[427]&~m[428]&~m[429])|(~m[213]&~m[425]&~m[427]&m[428]&~m[429])|(m[213]&m[425]&~m[427]&m[428]&~m[429])|(m[213]&~m[425]&m[427]&m[428]&~m[429])|(~m[213]&m[425]&~m[427]&~m[428]&m[429])|(~m[213]&~m[425]&m[427]&~m[428]&m[429])|(m[213]&m[425]&m[427]&~m[428]&m[429])|(~m[213]&m[425]&m[427]&m[428]&m[429]))&UnbiasedRNG[157])|((m[213]&~m[425]&~m[427]&m[428]&~m[429])|(~m[213]&~m[425]&~m[427]&~m[428]&m[429])|(m[213]&~m[425]&~m[427]&~m[428]&m[429])|(m[213]&m[425]&~m[427]&~m[428]&m[429])|(m[213]&~m[425]&m[427]&~m[428]&m[429])|(~m[213]&~m[425]&~m[427]&m[428]&m[429])|(m[213]&~m[425]&~m[427]&m[428]&m[429])|(~m[213]&m[425]&~m[427]&m[428]&m[429])|(m[213]&m[425]&~m[427]&m[428]&m[429])|(~m[213]&~m[425]&m[427]&m[428]&m[429])|(m[213]&~m[425]&m[427]&m[428]&m[429])|(m[213]&m[425]&m[427]&m[428]&m[429]))):InitCond[380];
    m[431] = run?((((m[220]&~m[430]&~m[432]&~m[433]&~m[434])|(~m[220]&~m[430]&~m[432]&m[433]&~m[434])|(m[220]&m[430]&~m[432]&m[433]&~m[434])|(m[220]&~m[430]&m[432]&m[433]&~m[434])|(~m[220]&m[430]&~m[432]&~m[433]&m[434])|(~m[220]&~m[430]&m[432]&~m[433]&m[434])|(m[220]&m[430]&m[432]&~m[433]&m[434])|(~m[220]&m[430]&m[432]&m[433]&m[434]))&UnbiasedRNG[158])|((m[220]&~m[430]&~m[432]&m[433]&~m[434])|(~m[220]&~m[430]&~m[432]&~m[433]&m[434])|(m[220]&~m[430]&~m[432]&~m[433]&m[434])|(m[220]&m[430]&~m[432]&~m[433]&m[434])|(m[220]&~m[430]&m[432]&~m[433]&m[434])|(~m[220]&~m[430]&~m[432]&m[433]&m[434])|(m[220]&~m[430]&~m[432]&m[433]&m[434])|(~m[220]&m[430]&~m[432]&m[433]&m[434])|(m[220]&m[430]&~m[432]&m[433]&m[434])|(~m[220]&~m[430]&m[432]&m[433]&m[434])|(m[220]&~m[430]&m[432]&m[433]&m[434])|(m[220]&m[430]&m[432]&m[433]&m[434]))):InitCond[381];
    m[436] = run?((((m[227]&~m[435]&~m[437]&~m[438]&~m[439])|(~m[227]&~m[435]&~m[437]&m[438]&~m[439])|(m[227]&m[435]&~m[437]&m[438]&~m[439])|(m[227]&~m[435]&m[437]&m[438]&~m[439])|(~m[227]&m[435]&~m[437]&~m[438]&m[439])|(~m[227]&~m[435]&m[437]&~m[438]&m[439])|(m[227]&m[435]&m[437]&~m[438]&m[439])|(~m[227]&m[435]&m[437]&m[438]&m[439]))&UnbiasedRNG[159])|((m[227]&~m[435]&~m[437]&m[438]&~m[439])|(~m[227]&~m[435]&~m[437]&~m[438]&m[439])|(m[227]&~m[435]&~m[437]&~m[438]&m[439])|(m[227]&m[435]&~m[437]&~m[438]&m[439])|(m[227]&~m[435]&m[437]&~m[438]&m[439])|(~m[227]&~m[435]&~m[437]&m[438]&m[439])|(m[227]&~m[435]&~m[437]&m[438]&m[439])|(~m[227]&m[435]&~m[437]&m[438]&m[439])|(m[227]&m[435]&~m[437]&m[438]&m[439])|(~m[227]&~m[435]&m[437]&m[438]&m[439])|(m[227]&~m[435]&m[437]&m[438]&m[439])|(m[227]&m[435]&m[437]&m[438]&m[439]))):InitCond[382];
    m[441] = run?((((m[234]&~m[440]&~m[442]&~m[443]&~m[444])|(~m[234]&~m[440]&~m[442]&m[443]&~m[444])|(m[234]&m[440]&~m[442]&m[443]&~m[444])|(m[234]&~m[440]&m[442]&m[443]&~m[444])|(~m[234]&m[440]&~m[442]&~m[443]&m[444])|(~m[234]&~m[440]&m[442]&~m[443]&m[444])|(m[234]&m[440]&m[442]&~m[443]&m[444])|(~m[234]&m[440]&m[442]&m[443]&m[444]))&UnbiasedRNG[160])|((m[234]&~m[440]&~m[442]&m[443]&~m[444])|(~m[234]&~m[440]&~m[442]&~m[443]&m[444])|(m[234]&~m[440]&~m[442]&~m[443]&m[444])|(m[234]&m[440]&~m[442]&~m[443]&m[444])|(m[234]&~m[440]&m[442]&~m[443]&m[444])|(~m[234]&~m[440]&~m[442]&m[443]&m[444])|(m[234]&~m[440]&~m[442]&m[443]&m[444])|(~m[234]&m[440]&~m[442]&m[443]&m[444])|(m[234]&m[440]&~m[442]&m[443]&m[444])|(~m[234]&~m[440]&m[442]&m[443]&m[444])|(m[234]&~m[440]&m[442]&m[443]&m[444])|(m[234]&m[440]&m[442]&m[443]&m[444]))):InitCond[383];
    m[446] = run?((((m[207]&~m[445]&~m[447]&~m[448]&~m[449])|(~m[207]&~m[445]&~m[447]&m[448]&~m[449])|(m[207]&m[445]&~m[447]&m[448]&~m[449])|(m[207]&~m[445]&m[447]&m[448]&~m[449])|(~m[207]&m[445]&~m[447]&~m[448]&m[449])|(~m[207]&~m[445]&m[447]&~m[448]&m[449])|(m[207]&m[445]&m[447]&~m[448]&m[449])|(~m[207]&m[445]&m[447]&m[448]&m[449]))&UnbiasedRNG[161])|((m[207]&~m[445]&~m[447]&m[448]&~m[449])|(~m[207]&~m[445]&~m[447]&~m[448]&m[449])|(m[207]&~m[445]&~m[447]&~m[448]&m[449])|(m[207]&m[445]&~m[447]&~m[448]&m[449])|(m[207]&~m[445]&m[447]&~m[448]&m[449])|(~m[207]&~m[445]&~m[447]&m[448]&m[449])|(m[207]&~m[445]&~m[447]&m[448]&m[449])|(~m[207]&m[445]&~m[447]&m[448]&m[449])|(m[207]&m[445]&~m[447]&m[448]&m[449])|(~m[207]&~m[445]&m[447]&m[448]&m[449])|(m[207]&~m[445]&m[447]&m[448]&m[449])|(m[207]&m[445]&m[447]&m[448]&m[449]))):InitCond[384];
    m[451] = run?((((m[214]&~m[450]&~m[452]&~m[453]&~m[454])|(~m[214]&~m[450]&~m[452]&m[453]&~m[454])|(m[214]&m[450]&~m[452]&m[453]&~m[454])|(m[214]&~m[450]&m[452]&m[453]&~m[454])|(~m[214]&m[450]&~m[452]&~m[453]&m[454])|(~m[214]&~m[450]&m[452]&~m[453]&m[454])|(m[214]&m[450]&m[452]&~m[453]&m[454])|(~m[214]&m[450]&m[452]&m[453]&m[454]))&UnbiasedRNG[162])|((m[214]&~m[450]&~m[452]&m[453]&~m[454])|(~m[214]&~m[450]&~m[452]&~m[453]&m[454])|(m[214]&~m[450]&~m[452]&~m[453]&m[454])|(m[214]&m[450]&~m[452]&~m[453]&m[454])|(m[214]&~m[450]&m[452]&~m[453]&m[454])|(~m[214]&~m[450]&~m[452]&m[453]&m[454])|(m[214]&~m[450]&~m[452]&m[453]&m[454])|(~m[214]&m[450]&~m[452]&m[453]&m[454])|(m[214]&m[450]&~m[452]&m[453]&m[454])|(~m[214]&~m[450]&m[452]&m[453]&m[454])|(m[214]&~m[450]&m[452]&m[453]&m[454])|(m[214]&m[450]&m[452]&m[453]&m[454]))):InitCond[385];
    m[456] = run?((((m[221]&~m[455]&~m[457]&~m[458]&~m[459])|(~m[221]&~m[455]&~m[457]&m[458]&~m[459])|(m[221]&m[455]&~m[457]&m[458]&~m[459])|(m[221]&~m[455]&m[457]&m[458]&~m[459])|(~m[221]&m[455]&~m[457]&~m[458]&m[459])|(~m[221]&~m[455]&m[457]&~m[458]&m[459])|(m[221]&m[455]&m[457]&~m[458]&m[459])|(~m[221]&m[455]&m[457]&m[458]&m[459]))&UnbiasedRNG[163])|((m[221]&~m[455]&~m[457]&m[458]&~m[459])|(~m[221]&~m[455]&~m[457]&~m[458]&m[459])|(m[221]&~m[455]&~m[457]&~m[458]&m[459])|(m[221]&m[455]&~m[457]&~m[458]&m[459])|(m[221]&~m[455]&m[457]&~m[458]&m[459])|(~m[221]&~m[455]&~m[457]&m[458]&m[459])|(m[221]&~m[455]&~m[457]&m[458]&m[459])|(~m[221]&m[455]&~m[457]&m[458]&m[459])|(m[221]&m[455]&~m[457]&m[458]&m[459])|(~m[221]&~m[455]&m[457]&m[458]&m[459])|(m[221]&~m[455]&m[457]&m[458]&m[459])|(m[221]&m[455]&m[457]&m[458]&m[459]))):InitCond[386];
    m[461] = run?((((m[228]&~m[460]&~m[462]&~m[463]&~m[464])|(~m[228]&~m[460]&~m[462]&m[463]&~m[464])|(m[228]&m[460]&~m[462]&m[463]&~m[464])|(m[228]&~m[460]&m[462]&m[463]&~m[464])|(~m[228]&m[460]&~m[462]&~m[463]&m[464])|(~m[228]&~m[460]&m[462]&~m[463]&m[464])|(m[228]&m[460]&m[462]&~m[463]&m[464])|(~m[228]&m[460]&m[462]&m[463]&m[464]))&UnbiasedRNG[164])|((m[228]&~m[460]&~m[462]&m[463]&~m[464])|(~m[228]&~m[460]&~m[462]&~m[463]&m[464])|(m[228]&~m[460]&~m[462]&~m[463]&m[464])|(m[228]&m[460]&~m[462]&~m[463]&m[464])|(m[228]&~m[460]&m[462]&~m[463]&m[464])|(~m[228]&~m[460]&~m[462]&m[463]&m[464])|(m[228]&~m[460]&~m[462]&m[463]&m[464])|(~m[228]&m[460]&~m[462]&m[463]&m[464])|(m[228]&m[460]&~m[462]&m[463]&m[464])|(~m[228]&~m[460]&m[462]&m[463]&m[464])|(m[228]&~m[460]&m[462]&m[463]&m[464])|(m[228]&m[460]&m[462]&m[463]&m[464]))):InitCond[387];
    m[466] = run?((((m[235]&~m[465]&~m[467]&~m[468]&~m[469])|(~m[235]&~m[465]&~m[467]&m[468]&~m[469])|(m[235]&m[465]&~m[467]&m[468]&~m[469])|(m[235]&~m[465]&m[467]&m[468]&~m[469])|(~m[235]&m[465]&~m[467]&~m[468]&m[469])|(~m[235]&~m[465]&m[467]&~m[468]&m[469])|(m[235]&m[465]&m[467]&~m[468]&m[469])|(~m[235]&m[465]&m[467]&m[468]&m[469]))&UnbiasedRNG[165])|((m[235]&~m[465]&~m[467]&m[468]&~m[469])|(~m[235]&~m[465]&~m[467]&~m[468]&m[469])|(m[235]&~m[465]&~m[467]&~m[468]&m[469])|(m[235]&m[465]&~m[467]&~m[468]&m[469])|(m[235]&~m[465]&m[467]&~m[468]&m[469])|(~m[235]&~m[465]&~m[467]&m[468]&m[469])|(m[235]&~m[465]&~m[467]&m[468]&m[469])|(~m[235]&m[465]&~m[467]&m[468]&m[469])|(m[235]&m[465]&~m[467]&m[468]&m[469])|(~m[235]&~m[465]&m[467]&m[468]&m[469])|(m[235]&~m[465]&m[467]&m[468]&m[469])|(m[235]&m[465]&m[467]&m[468]&m[469]))):InitCond[388];
    m[471] = run?((((m[215]&~m[470]&~m[472]&~m[473]&~m[474])|(~m[215]&~m[470]&~m[472]&m[473]&~m[474])|(m[215]&m[470]&~m[472]&m[473]&~m[474])|(m[215]&~m[470]&m[472]&m[473]&~m[474])|(~m[215]&m[470]&~m[472]&~m[473]&m[474])|(~m[215]&~m[470]&m[472]&~m[473]&m[474])|(m[215]&m[470]&m[472]&~m[473]&m[474])|(~m[215]&m[470]&m[472]&m[473]&m[474]))&UnbiasedRNG[166])|((m[215]&~m[470]&~m[472]&m[473]&~m[474])|(~m[215]&~m[470]&~m[472]&~m[473]&m[474])|(m[215]&~m[470]&~m[472]&~m[473]&m[474])|(m[215]&m[470]&~m[472]&~m[473]&m[474])|(m[215]&~m[470]&m[472]&~m[473]&m[474])|(~m[215]&~m[470]&~m[472]&m[473]&m[474])|(m[215]&~m[470]&~m[472]&m[473]&m[474])|(~m[215]&m[470]&~m[472]&m[473]&m[474])|(m[215]&m[470]&~m[472]&m[473]&m[474])|(~m[215]&~m[470]&m[472]&m[473]&m[474])|(m[215]&~m[470]&m[472]&m[473]&m[474])|(m[215]&m[470]&m[472]&m[473]&m[474]))):InitCond[389];
    m[476] = run?((((m[222]&~m[475]&~m[477]&~m[478]&~m[479])|(~m[222]&~m[475]&~m[477]&m[478]&~m[479])|(m[222]&m[475]&~m[477]&m[478]&~m[479])|(m[222]&~m[475]&m[477]&m[478]&~m[479])|(~m[222]&m[475]&~m[477]&~m[478]&m[479])|(~m[222]&~m[475]&m[477]&~m[478]&m[479])|(m[222]&m[475]&m[477]&~m[478]&m[479])|(~m[222]&m[475]&m[477]&m[478]&m[479]))&UnbiasedRNG[167])|((m[222]&~m[475]&~m[477]&m[478]&~m[479])|(~m[222]&~m[475]&~m[477]&~m[478]&m[479])|(m[222]&~m[475]&~m[477]&~m[478]&m[479])|(m[222]&m[475]&~m[477]&~m[478]&m[479])|(m[222]&~m[475]&m[477]&~m[478]&m[479])|(~m[222]&~m[475]&~m[477]&m[478]&m[479])|(m[222]&~m[475]&~m[477]&m[478]&m[479])|(~m[222]&m[475]&~m[477]&m[478]&m[479])|(m[222]&m[475]&~m[477]&m[478]&m[479])|(~m[222]&~m[475]&m[477]&m[478]&m[479])|(m[222]&~m[475]&m[477]&m[478]&m[479])|(m[222]&m[475]&m[477]&m[478]&m[479]))):InitCond[390];
    m[481] = run?((((m[229]&~m[480]&~m[482]&~m[483]&~m[484])|(~m[229]&~m[480]&~m[482]&m[483]&~m[484])|(m[229]&m[480]&~m[482]&m[483]&~m[484])|(m[229]&~m[480]&m[482]&m[483]&~m[484])|(~m[229]&m[480]&~m[482]&~m[483]&m[484])|(~m[229]&~m[480]&m[482]&~m[483]&m[484])|(m[229]&m[480]&m[482]&~m[483]&m[484])|(~m[229]&m[480]&m[482]&m[483]&m[484]))&UnbiasedRNG[168])|((m[229]&~m[480]&~m[482]&m[483]&~m[484])|(~m[229]&~m[480]&~m[482]&~m[483]&m[484])|(m[229]&~m[480]&~m[482]&~m[483]&m[484])|(m[229]&m[480]&~m[482]&~m[483]&m[484])|(m[229]&~m[480]&m[482]&~m[483]&m[484])|(~m[229]&~m[480]&~m[482]&m[483]&m[484])|(m[229]&~m[480]&~m[482]&m[483]&m[484])|(~m[229]&m[480]&~m[482]&m[483]&m[484])|(m[229]&m[480]&~m[482]&m[483]&m[484])|(~m[229]&~m[480]&m[482]&m[483]&m[484])|(m[229]&~m[480]&m[482]&m[483]&m[484])|(m[229]&m[480]&m[482]&m[483]&m[484]))):InitCond[391];
    m[486] = run?((((m[236]&~m[485]&~m[487]&~m[488]&~m[489])|(~m[236]&~m[485]&~m[487]&m[488]&~m[489])|(m[236]&m[485]&~m[487]&m[488]&~m[489])|(m[236]&~m[485]&m[487]&m[488]&~m[489])|(~m[236]&m[485]&~m[487]&~m[488]&m[489])|(~m[236]&~m[485]&m[487]&~m[488]&m[489])|(m[236]&m[485]&m[487]&~m[488]&m[489])|(~m[236]&m[485]&m[487]&m[488]&m[489]))&UnbiasedRNG[169])|((m[236]&~m[485]&~m[487]&m[488]&~m[489])|(~m[236]&~m[485]&~m[487]&~m[488]&m[489])|(m[236]&~m[485]&~m[487]&~m[488]&m[489])|(m[236]&m[485]&~m[487]&~m[488]&m[489])|(m[236]&~m[485]&m[487]&~m[488]&m[489])|(~m[236]&~m[485]&~m[487]&m[488]&m[489])|(m[236]&~m[485]&~m[487]&m[488]&m[489])|(~m[236]&m[485]&~m[487]&m[488]&m[489])|(m[236]&m[485]&~m[487]&m[488]&m[489])|(~m[236]&~m[485]&m[487]&m[488]&m[489])|(m[236]&~m[485]&m[487]&m[488]&m[489])|(m[236]&m[485]&m[487]&m[488]&m[489]))):InitCond[392];
    m[491] = run?((((m[223]&~m[490]&~m[492]&~m[493]&~m[494])|(~m[223]&~m[490]&~m[492]&m[493]&~m[494])|(m[223]&m[490]&~m[492]&m[493]&~m[494])|(m[223]&~m[490]&m[492]&m[493]&~m[494])|(~m[223]&m[490]&~m[492]&~m[493]&m[494])|(~m[223]&~m[490]&m[492]&~m[493]&m[494])|(m[223]&m[490]&m[492]&~m[493]&m[494])|(~m[223]&m[490]&m[492]&m[493]&m[494]))&UnbiasedRNG[170])|((m[223]&~m[490]&~m[492]&m[493]&~m[494])|(~m[223]&~m[490]&~m[492]&~m[493]&m[494])|(m[223]&~m[490]&~m[492]&~m[493]&m[494])|(m[223]&m[490]&~m[492]&~m[493]&m[494])|(m[223]&~m[490]&m[492]&~m[493]&m[494])|(~m[223]&~m[490]&~m[492]&m[493]&m[494])|(m[223]&~m[490]&~m[492]&m[493]&m[494])|(~m[223]&m[490]&~m[492]&m[493]&m[494])|(m[223]&m[490]&~m[492]&m[493]&m[494])|(~m[223]&~m[490]&m[492]&m[493]&m[494])|(m[223]&~m[490]&m[492]&m[493]&m[494])|(m[223]&m[490]&m[492]&m[493]&m[494]))):InitCond[393];
    m[496] = run?((((m[230]&~m[495]&~m[497]&~m[498]&~m[499])|(~m[230]&~m[495]&~m[497]&m[498]&~m[499])|(m[230]&m[495]&~m[497]&m[498]&~m[499])|(m[230]&~m[495]&m[497]&m[498]&~m[499])|(~m[230]&m[495]&~m[497]&~m[498]&m[499])|(~m[230]&~m[495]&m[497]&~m[498]&m[499])|(m[230]&m[495]&m[497]&~m[498]&m[499])|(~m[230]&m[495]&m[497]&m[498]&m[499]))&UnbiasedRNG[171])|((m[230]&~m[495]&~m[497]&m[498]&~m[499])|(~m[230]&~m[495]&~m[497]&~m[498]&m[499])|(m[230]&~m[495]&~m[497]&~m[498]&m[499])|(m[230]&m[495]&~m[497]&~m[498]&m[499])|(m[230]&~m[495]&m[497]&~m[498]&m[499])|(~m[230]&~m[495]&~m[497]&m[498]&m[499])|(m[230]&~m[495]&~m[497]&m[498]&m[499])|(~m[230]&m[495]&~m[497]&m[498]&m[499])|(m[230]&m[495]&~m[497]&m[498]&m[499])|(~m[230]&~m[495]&m[497]&m[498]&m[499])|(m[230]&~m[495]&m[497]&m[498]&m[499])|(m[230]&m[495]&m[497]&m[498]&m[499]))):InitCond[394];
    m[501] = run?((((m[237]&~m[500]&~m[502]&~m[503]&~m[504])|(~m[237]&~m[500]&~m[502]&m[503]&~m[504])|(m[237]&m[500]&~m[502]&m[503]&~m[504])|(m[237]&~m[500]&m[502]&m[503]&~m[504])|(~m[237]&m[500]&~m[502]&~m[503]&m[504])|(~m[237]&~m[500]&m[502]&~m[503]&m[504])|(m[237]&m[500]&m[502]&~m[503]&m[504])|(~m[237]&m[500]&m[502]&m[503]&m[504]))&UnbiasedRNG[172])|((m[237]&~m[500]&~m[502]&m[503]&~m[504])|(~m[237]&~m[500]&~m[502]&~m[503]&m[504])|(m[237]&~m[500]&~m[502]&~m[503]&m[504])|(m[237]&m[500]&~m[502]&~m[503]&m[504])|(m[237]&~m[500]&m[502]&~m[503]&m[504])|(~m[237]&~m[500]&~m[502]&m[503]&m[504])|(m[237]&~m[500]&~m[502]&m[503]&m[504])|(~m[237]&m[500]&~m[502]&m[503]&m[504])|(m[237]&m[500]&~m[502]&m[503]&m[504])|(~m[237]&~m[500]&m[502]&m[503]&m[504])|(m[237]&~m[500]&m[502]&m[503]&m[504])|(m[237]&m[500]&m[502]&m[503]&m[504]))):InitCond[395];
    m[506] = run?((((m[231]&~m[505]&~m[507]&~m[508]&~m[509])|(~m[231]&~m[505]&~m[507]&m[508]&~m[509])|(m[231]&m[505]&~m[507]&m[508]&~m[509])|(m[231]&~m[505]&m[507]&m[508]&~m[509])|(~m[231]&m[505]&~m[507]&~m[508]&m[509])|(~m[231]&~m[505]&m[507]&~m[508]&m[509])|(m[231]&m[505]&m[507]&~m[508]&m[509])|(~m[231]&m[505]&m[507]&m[508]&m[509]))&UnbiasedRNG[173])|((m[231]&~m[505]&~m[507]&m[508]&~m[509])|(~m[231]&~m[505]&~m[507]&~m[508]&m[509])|(m[231]&~m[505]&~m[507]&~m[508]&m[509])|(m[231]&m[505]&~m[507]&~m[508]&m[509])|(m[231]&~m[505]&m[507]&~m[508]&m[509])|(~m[231]&~m[505]&~m[507]&m[508]&m[509])|(m[231]&~m[505]&~m[507]&m[508]&m[509])|(~m[231]&m[505]&~m[507]&m[508]&m[509])|(m[231]&m[505]&~m[507]&m[508]&m[509])|(~m[231]&~m[505]&m[507]&m[508]&m[509])|(m[231]&~m[505]&m[507]&m[508]&m[509])|(m[231]&m[505]&m[507]&m[508]&m[509]))):InitCond[396];
    m[511] = run?((((m[238]&~m[510]&~m[512]&~m[513]&~m[514])|(~m[238]&~m[510]&~m[512]&m[513]&~m[514])|(m[238]&m[510]&~m[512]&m[513]&~m[514])|(m[238]&~m[510]&m[512]&m[513]&~m[514])|(~m[238]&m[510]&~m[512]&~m[513]&m[514])|(~m[238]&~m[510]&m[512]&~m[513]&m[514])|(m[238]&m[510]&m[512]&~m[513]&m[514])|(~m[238]&m[510]&m[512]&m[513]&m[514]))&UnbiasedRNG[174])|((m[238]&~m[510]&~m[512]&m[513]&~m[514])|(~m[238]&~m[510]&~m[512]&~m[513]&m[514])|(m[238]&~m[510]&~m[512]&~m[513]&m[514])|(m[238]&m[510]&~m[512]&~m[513]&m[514])|(m[238]&~m[510]&m[512]&~m[513]&m[514])|(~m[238]&~m[510]&~m[512]&m[513]&m[514])|(m[238]&~m[510]&~m[512]&m[513]&m[514])|(~m[238]&m[510]&~m[512]&m[513]&m[514])|(m[238]&m[510]&~m[512]&m[513]&m[514])|(~m[238]&~m[510]&m[512]&m[513]&m[514])|(m[238]&~m[510]&m[512]&m[513]&m[514])|(m[238]&m[510]&m[512]&m[513]&m[514]))):InitCond[397];
    m[516] = run?((((m[239]&~m[515]&~m[517]&~m[518]&~m[519])|(~m[239]&~m[515]&~m[517]&m[518]&~m[519])|(m[239]&m[515]&~m[517]&m[518]&~m[519])|(m[239]&~m[515]&m[517]&m[518]&~m[519])|(~m[239]&m[515]&~m[517]&~m[518]&m[519])|(~m[239]&~m[515]&m[517]&~m[518]&m[519])|(m[239]&m[515]&m[517]&~m[518]&m[519])|(~m[239]&m[515]&m[517]&m[518]&m[519]))&UnbiasedRNG[175])|((m[239]&~m[515]&~m[517]&m[518]&~m[519])|(~m[239]&~m[515]&~m[517]&~m[518]&m[519])|(m[239]&~m[515]&~m[517]&~m[518]&m[519])|(m[239]&m[515]&~m[517]&~m[518]&m[519])|(m[239]&~m[515]&m[517]&~m[518]&m[519])|(~m[239]&~m[515]&~m[517]&m[518]&m[519])|(m[239]&~m[515]&~m[517]&m[518]&m[519])|(~m[239]&m[515]&~m[517]&m[518]&m[519])|(m[239]&m[515]&~m[517]&m[518]&m[519])|(~m[239]&~m[515]&m[517]&m[518]&m[519])|(m[239]&~m[515]&m[517]&m[518]&m[519])|(m[239]&m[515]&m[517]&m[518]&m[519]))):InitCond[398];
end

always @(posedge color3_clk) begin
    m[248] = run?((((m[245]&~m[246]&~m[247]&~m[249]&~m[250])|(~m[245]&m[246]&~m[247]&~m[249]&~m[250])|(~m[245]&~m[246]&m[247]&~m[249]&~m[250])|(m[245]&m[246]&m[247]&m[249]&~m[250])|(~m[245]&~m[246]&~m[247]&~m[249]&m[250])|(m[245]&m[246]&~m[247]&m[249]&m[250])|(m[245]&~m[246]&m[247]&m[249]&m[250])|(~m[245]&m[246]&m[247]&m[249]&m[250]))&UnbiasedRNG[176])|((m[245]&m[246]&~m[247]&~m[249]&~m[250])|(m[245]&~m[246]&m[247]&~m[249]&~m[250])|(~m[245]&m[246]&m[247]&~m[249]&~m[250])|(m[245]&m[246]&m[247]&~m[249]&~m[250])|(m[245]&~m[246]&~m[247]&~m[249]&m[250])|(~m[245]&m[246]&~m[247]&~m[249]&m[250])|(m[245]&m[246]&~m[247]&~m[249]&m[250])|(~m[245]&~m[246]&m[247]&~m[249]&m[250])|(m[245]&~m[246]&m[247]&~m[249]&m[250])|(~m[245]&m[246]&m[247]&~m[249]&m[250])|(m[245]&m[246]&m[247]&~m[249]&m[250])|(m[245]&m[246]&m[247]&m[249]&m[250]))):InitCond[399];
    m[258] = run?((((m[255]&~m[256]&~m[257]&~m[259]&~m[260])|(~m[255]&m[256]&~m[257]&~m[259]&~m[260])|(~m[255]&~m[256]&m[257]&~m[259]&~m[260])|(m[255]&m[256]&m[257]&m[259]&~m[260])|(~m[255]&~m[256]&~m[257]&~m[259]&m[260])|(m[255]&m[256]&~m[257]&m[259]&m[260])|(m[255]&~m[256]&m[257]&m[259]&m[260])|(~m[255]&m[256]&m[257]&m[259]&m[260]))&UnbiasedRNG[177])|((m[255]&m[256]&~m[257]&~m[259]&~m[260])|(m[255]&~m[256]&m[257]&~m[259]&~m[260])|(~m[255]&m[256]&m[257]&~m[259]&~m[260])|(m[255]&m[256]&m[257]&~m[259]&~m[260])|(m[255]&~m[256]&~m[257]&~m[259]&m[260])|(~m[255]&m[256]&~m[257]&~m[259]&m[260])|(m[255]&m[256]&~m[257]&~m[259]&m[260])|(~m[255]&~m[256]&m[257]&~m[259]&m[260])|(m[255]&~m[256]&m[257]&~m[259]&m[260])|(~m[255]&m[256]&m[257]&~m[259]&m[260])|(m[255]&m[256]&m[257]&~m[259]&m[260])|(m[255]&m[256]&m[257]&m[259]&m[260]))):InitCond[400];
    m[263] = run?((((m[260]&~m[261]&~m[262]&~m[264]&~m[265])|(~m[260]&m[261]&~m[262]&~m[264]&~m[265])|(~m[260]&~m[261]&m[262]&~m[264]&~m[265])|(m[260]&m[261]&m[262]&m[264]&~m[265])|(~m[260]&~m[261]&~m[262]&~m[264]&m[265])|(m[260]&m[261]&~m[262]&m[264]&m[265])|(m[260]&~m[261]&m[262]&m[264]&m[265])|(~m[260]&m[261]&m[262]&m[264]&m[265]))&UnbiasedRNG[178])|((m[260]&m[261]&~m[262]&~m[264]&~m[265])|(m[260]&~m[261]&m[262]&~m[264]&~m[265])|(~m[260]&m[261]&m[262]&~m[264]&~m[265])|(m[260]&m[261]&m[262]&~m[264]&~m[265])|(m[260]&~m[261]&~m[262]&~m[264]&m[265])|(~m[260]&m[261]&~m[262]&~m[264]&m[265])|(m[260]&m[261]&~m[262]&~m[264]&m[265])|(~m[260]&~m[261]&m[262]&~m[264]&m[265])|(m[260]&~m[261]&m[262]&~m[264]&m[265])|(~m[260]&m[261]&m[262]&~m[264]&m[265])|(m[260]&m[261]&m[262]&~m[264]&m[265])|(m[260]&m[261]&m[262]&m[264]&m[265]))):InitCond[401];
    m[273] = run?((((m[270]&~m[271]&~m[272]&~m[274]&~m[275])|(~m[270]&m[271]&~m[272]&~m[274]&~m[275])|(~m[270]&~m[271]&m[272]&~m[274]&~m[275])|(m[270]&m[271]&m[272]&m[274]&~m[275])|(~m[270]&~m[271]&~m[272]&~m[274]&m[275])|(m[270]&m[271]&~m[272]&m[274]&m[275])|(m[270]&~m[271]&m[272]&m[274]&m[275])|(~m[270]&m[271]&m[272]&m[274]&m[275]))&UnbiasedRNG[179])|((m[270]&m[271]&~m[272]&~m[274]&~m[275])|(m[270]&~m[271]&m[272]&~m[274]&~m[275])|(~m[270]&m[271]&m[272]&~m[274]&~m[275])|(m[270]&m[271]&m[272]&~m[274]&~m[275])|(m[270]&~m[271]&~m[272]&~m[274]&m[275])|(~m[270]&m[271]&~m[272]&~m[274]&m[275])|(m[270]&m[271]&~m[272]&~m[274]&m[275])|(~m[270]&~m[271]&m[272]&~m[274]&m[275])|(m[270]&~m[271]&m[272]&~m[274]&m[275])|(~m[270]&m[271]&m[272]&~m[274]&m[275])|(m[270]&m[271]&m[272]&~m[274]&m[275])|(m[270]&m[271]&m[272]&m[274]&m[275]))):InitCond[402];
    m[278] = run?((((m[275]&~m[276]&~m[277]&~m[279]&~m[280])|(~m[275]&m[276]&~m[277]&~m[279]&~m[280])|(~m[275]&~m[276]&m[277]&~m[279]&~m[280])|(m[275]&m[276]&m[277]&m[279]&~m[280])|(~m[275]&~m[276]&~m[277]&~m[279]&m[280])|(m[275]&m[276]&~m[277]&m[279]&m[280])|(m[275]&~m[276]&m[277]&m[279]&m[280])|(~m[275]&m[276]&m[277]&m[279]&m[280]))&UnbiasedRNG[180])|((m[275]&m[276]&~m[277]&~m[279]&~m[280])|(m[275]&~m[276]&m[277]&~m[279]&~m[280])|(~m[275]&m[276]&m[277]&~m[279]&~m[280])|(m[275]&m[276]&m[277]&~m[279]&~m[280])|(m[275]&~m[276]&~m[277]&~m[279]&m[280])|(~m[275]&m[276]&~m[277]&~m[279]&m[280])|(m[275]&m[276]&~m[277]&~m[279]&m[280])|(~m[275]&~m[276]&m[277]&~m[279]&m[280])|(m[275]&~m[276]&m[277]&~m[279]&m[280])|(~m[275]&m[276]&m[277]&~m[279]&m[280])|(m[275]&m[276]&m[277]&~m[279]&m[280])|(m[275]&m[276]&m[277]&m[279]&m[280]))):InitCond[403];
    m[283] = run?((((m[280]&~m[281]&~m[282]&~m[284]&~m[285])|(~m[280]&m[281]&~m[282]&~m[284]&~m[285])|(~m[280]&~m[281]&m[282]&~m[284]&~m[285])|(m[280]&m[281]&m[282]&m[284]&~m[285])|(~m[280]&~m[281]&~m[282]&~m[284]&m[285])|(m[280]&m[281]&~m[282]&m[284]&m[285])|(m[280]&~m[281]&m[282]&m[284]&m[285])|(~m[280]&m[281]&m[282]&m[284]&m[285]))&UnbiasedRNG[181])|((m[280]&m[281]&~m[282]&~m[284]&~m[285])|(m[280]&~m[281]&m[282]&~m[284]&~m[285])|(~m[280]&m[281]&m[282]&~m[284]&~m[285])|(m[280]&m[281]&m[282]&~m[284]&~m[285])|(m[280]&~m[281]&~m[282]&~m[284]&m[285])|(~m[280]&m[281]&~m[282]&~m[284]&m[285])|(m[280]&m[281]&~m[282]&~m[284]&m[285])|(~m[280]&~m[281]&m[282]&~m[284]&m[285])|(m[280]&~m[281]&m[282]&~m[284]&m[285])|(~m[280]&m[281]&m[282]&~m[284]&m[285])|(m[280]&m[281]&m[282]&~m[284]&m[285])|(m[280]&m[281]&m[282]&m[284]&m[285]))):InitCond[404];
    m[293] = run?((((m[290]&~m[291]&~m[292]&~m[294]&~m[295])|(~m[290]&m[291]&~m[292]&~m[294]&~m[295])|(~m[290]&~m[291]&m[292]&~m[294]&~m[295])|(m[290]&m[291]&m[292]&m[294]&~m[295])|(~m[290]&~m[291]&~m[292]&~m[294]&m[295])|(m[290]&m[291]&~m[292]&m[294]&m[295])|(m[290]&~m[291]&m[292]&m[294]&m[295])|(~m[290]&m[291]&m[292]&m[294]&m[295]))&UnbiasedRNG[182])|((m[290]&m[291]&~m[292]&~m[294]&~m[295])|(m[290]&~m[291]&m[292]&~m[294]&~m[295])|(~m[290]&m[291]&m[292]&~m[294]&~m[295])|(m[290]&m[291]&m[292]&~m[294]&~m[295])|(m[290]&~m[291]&~m[292]&~m[294]&m[295])|(~m[290]&m[291]&~m[292]&~m[294]&m[295])|(m[290]&m[291]&~m[292]&~m[294]&m[295])|(~m[290]&~m[291]&m[292]&~m[294]&m[295])|(m[290]&~m[291]&m[292]&~m[294]&m[295])|(~m[290]&m[291]&m[292]&~m[294]&m[295])|(m[290]&m[291]&m[292]&~m[294]&m[295])|(m[290]&m[291]&m[292]&m[294]&m[295]))):InitCond[405];
    m[298] = run?((((m[295]&~m[296]&~m[297]&~m[299]&~m[300])|(~m[295]&m[296]&~m[297]&~m[299]&~m[300])|(~m[295]&~m[296]&m[297]&~m[299]&~m[300])|(m[295]&m[296]&m[297]&m[299]&~m[300])|(~m[295]&~m[296]&~m[297]&~m[299]&m[300])|(m[295]&m[296]&~m[297]&m[299]&m[300])|(m[295]&~m[296]&m[297]&m[299]&m[300])|(~m[295]&m[296]&m[297]&m[299]&m[300]))&UnbiasedRNG[183])|((m[295]&m[296]&~m[297]&~m[299]&~m[300])|(m[295]&~m[296]&m[297]&~m[299]&~m[300])|(~m[295]&m[296]&m[297]&~m[299]&~m[300])|(m[295]&m[296]&m[297]&~m[299]&~m[300])|(m[295]&~m[296]&~m[297]&~m[299]&m[300])|(~m[295]&m[296]&~m[297]&~m[299]&m[300])|(m[295]&m[296]&~m[297]&~m[299]&m[300])|(~m[295]&~m[296]&m[297]&~m[299]&m[300])|(m[295]&~m[296]&m[297]&~m[299]&m[300])|(~m[295]&m[296]&m[297]&~m[299]&m[300])|(m[295]&m[296]&m[297]&~m[299]&m[300])|(m[295]&m[296]&m[297]&m[299]&m[300]))):InitCond[406];
    m[303] = run?((((m[300]&~m[301]&~m[302]&~m[304]&~m[305])|(~m[300]&m[301]&~m[302]&~m[304]&~m[305])|(~m[300]&~m[301]&m[302]&~m[304]&~m[305])|(m[300]&m[301]&m[302]&m[304]&~m[305])|(~m[300]&~m[301]&~m[302]&~m[304]&m[305])|(m[300]&m[301]&~m[302]&m[304]&m[305])|(m[300]&~m[301]&m[302]&m[304]&m[305])|(~m[300]&m[301]&m[302]&m[304]&m[305]))&UnbiasedRNG[184])|((m[300]&m[301]&~m[302]&~m[304]&~m[305])|(m[300]&~m[301]&m[302]&~m[304]&~m[305])|(~m[300]&m[301]&m[302]&~m[304]&~m[305])|(m[300]&m[301]&m[302]&~m[304]&~m[305])|(m[300]&~m[301]&~m[302]&~m[304]&m[305])|(~m[300]&m[301]&~m[302]&~m[304]&m[305])|(m[300]&m[301]&~m[302]&~m[304]&m[305])|(~m[300]&~m[301]&m[302]&~m[304]&m[305])|(m[300]&~m[301]&m[302]&~m[304]&m[305])|(~m[300]&m[301]&m[302]&~m[304]&m[305])|(m[300]&m[301]&m[302]&~m[304]&m[305])|(m[300]&m[301]&m[302]&m[304]&m[305]))):InitCond[407];
    m[308] = run?((((m[305]&~m[306]&~m[307]&~m[309]&~m[310])|(~m[305]&m[306]&~m[307]&~m[309]&~m[310])|(~m[305]&~m[306]&m[307]&~m[309]&~m[310])|(m[305]&m[306]&m[307]&m[309]&~m[310])|(~m[305]&~m[306]&~m[307]&~m[309]&m[310])|(m[305]&m[306]&~m[307]&m[309]&m[310])|(m[305]&~m[306]&m[307]&m[309]&m[310])|(~m[305]&m[306]&m[307]&m[309]&m[310]))&UnbiasedRNG[185])|((m[305]&m[306]&~m[307]&~m[309]&~m[310])|(m[305]&~m[306]&m[307]&~m[309]&~m[310])|(~m[305]&m[306]&m[307]&~m[309]&~m[310])|(m[305]&m[306]&m[307]&~m[309]&~m[310])|(m[305]&~m[306]&~m[307]&~m[309]&m[310])|(~m[305]&m[306]&~m[307]&~m[309]&m[310])|(m[305]&m[306]&~m[307]&~m[309]&m[310])|(~m[305]&~m[306]&m[307]&~m[309]&m[310])|(m[305]&~m[306]&m[307]&~m[309]&m[310])|(~m[305]&m[306]&m[307]&~m[309]&m[310])|(m[305]&m[306]&m[307]&~m[309]&m[310])|(m[305]&m[306]&m[307]&m[309]&m[310]))):InitCond[408];
    m[318] = run?((((m[315]&~m[316]&~m[317]&~m[319]&~m[320])|(~m[315]&m[316]&~m[317]&~m[319]&~m[320])|(~m[315]&~m[316]&m[317]&~m[319]&~m[320])|(m[315]&m[316]&m[317]&m[319]&~m[320])|(~m[315]&~m[316]&~m[317]&~m[319]&m[320])|(m[315]&m[316]&~m[317]&m[319]&m[320])|(m[315]&~m[316]&m[317]&m[319]&m[320])|(~m[315]&m[316]&m[317]&m[319]&m[320]))&UnbiasedRNG[186])|((m[315]&m[316]&~m[317]&~m[319]&~m[320])|(m[315]&~m[316]&m[317]&~m[319]&~m[320])|(~m[315]&m[316]&m[317]&~m[319]&~m[320])|(m[315]&m[316]&m[317]&~m[319]&~m[320])|(m[315]&~m[316]&~m[317]&~m[319]&m[320])|(~m[315]&m[316]&~m[317]&~m[319]&m[320])|(m[315]&m[316]&~m[317]&~m[319]&m[320])|(~m[315]&~m[316]&m[317]&~m[319]&m[320])|(m[315]&~m[316]&m[317]&~m[319]&m[320])|(~m[315]&m[316]&m[317]&~m[319]&m[320])|(m[315]&m[316]&m[317]&~m[319]&m[320])|(m[315]&m[316]&m[317]&m[319]&m[320]))):InitCond[409];
    m[323] = run?((((m[320]&~m[321]&~m[322]&~m[324]&~m[325])|(~m[320]&m[321]&~m[322]&~m[324]&~m[325])|(~m[320]&~m[321]&m[322]&~m[324]&~m[325])|(m[320]&m[321]&m[322]&m[324]&~m[325])|(~m[320]&~m[321]&~m[322]&~m[324]&m[325])|(m[320]&m[321]&~m[322]&m[324]&m[325])|(m[320]&~m[321]&m[322]&m[324]&m[325])|(~m[320]&m[321]&m[322]&m[324]&m[325]))&UnbiasedRNG[187])|((m[320]&m[321]&~m[322]&~m[324]&~m[325])|(m[320]&~m[321]&m[322]&~m[324]&~m[325])|(~m[320]&m[321]&m[322]&~m[324]&~m[325])|(m[320]&m[321]&m[322]&~m[324]&~m[325])|(m[320]&~m[321]&~m[322]&~m[324]&m[325])|(~m[320]&m[321]&~m[322]&~m[324]&m[325])|(m[320]&m[321]&~m[322]&~m[324]&m[325])|(~m[320]&~m[321]&m[322]&~m[324]&m[325])|(m[320]&~m[321]&m[322]&~m[324]&m[325])|(~m[320]&m[321]&m[322]&~m[324]&m[325])|(m[320]&m[321]&m[322]&~m[324]&m[325])|(m[320]&m[321]&m[322]&m[324]&m[325]))):InitCond[410];
    m[328] = run?((((m[325]&~m[326]&~m[327]&~m[329]&~m[330])|(~m[325]&m[326]&~m[327]&~m[329]&~m[330])|(~m[325]&~m[326]&m[327]&~m[329]&~m[330])|(m[325]&m[326]&m[327]&m[329]&~m[330])|(~m[325]&~m[326]&~m[327]&~m[329]&m[330])|(m[325]&m[326]&~m[327]&m[329]&m[330])|(m[325]&~m[326]&m[327]&m[329]&m[330])|(~m[325]&m[326]&m[327]&m[329]&m[330]))&UnbiasedRNG[188])|((m[325]&m[326]&~m[327]&~m[329]&~m[330])|(m[325]&~m[326]&m[327]&~m[329]&~m[330])|(~m[325]&m[326]&m[327]&~m[329]&~m[330])|(m[325]&m[326]&m[327]&~m[329]&~m[330])|(m[325]&~m[326]&~m[327]&~m[329]&m[330])|(~m[325]&m[326]&~m[327]&~m[329]&m[330])|(m[325]&m[326]&~m[327]&~m[329]&m[330])|(~m[325]&~m[326]&m[327]&~m[329]&m[330])|(m[325]&~m[326]&m[327]&~m[329]&m[330])|(~m[325]&m[326]&m[327]&~m[329]&m[330])|(m[325]&m[326]&m[327]&~m[329]&m[330])|(m[325]&m[326]&m[327]&m[329]&m[330]))):InitCond[411];
    m[333] = run?((((m[330]&~m[331]&~m[332]&~m[334]&~m[335])|(~m[330]&m[331]&~m[332]&~m[334]&~m[335])|(~m[330]&~m[331]&m[332]&~m[334]&~m[335])|(m[330]&m[331]&m[332]&m[334]&~m[335])|(~m[330]&~m[331]&~m[332]&~m[334]&m[335])|(m[330]&m[331]&~m[332]&m[334]&m[335])|(m[330]&~m[331]&m[332]&m[334]&m[335])|(~m[330]&m[331]&m[332]&m[334]&m[335]))&UnbiasedRNG[189])|((m[330]&m[331]&~m[332]&~m[334]&~m[335])|(m[330]&~m[331]&m[332]&~m[334]&~m[335])|(~m[330]&m[331]&m[332]&~m[334]&~m[335])|(m[330]&m[331]&m[332]&~m[334]&~m[335])|(m[330]&~m[331]&~m[332]&~m[334]&m[335])|(~m[330]&m[331]&~m[332]&~m[334]&m[335])|(m[330]&m[331]&~m[332]&~m[334]&m[335])|(~m[330]&~m[331]&m[332]&~m[334]&m[335])|(m[330]&~m[331]&m[332]&~m[334]&m[335])|(~m[330]&m[331]&m[332]&~m[334]&m[335])|(m[330]&m[331]&m[332]&~m[334]&m[335])|(m[330]&m[331]&m[332]&m[334]&m[335]))):InitCond[412];
    m[338] = run?((((m[335]&~m[336]&~m[337]&~m[339]&~m[340])|(~m[335]&m[336]&~m[337]&~m[339]&~m[340])|(~m[335]&~m[336]&m[337]&~m[339]&~m[340])|(m[335]&m[336]&m[337]&m[339]&~m[340])|(~m[335]&~m[336]&~m[337]&~m[339]&m[340])|(m[335]&m[336]&~m[337]&m[339]&m[340])|(m[335]&~m[336]&m[337]&m[339]&m[340])|(~m[335]&m[336]&m[337]&m[339]&m[340]))&UnbiasedRNG[190])|((m[335]&m[336]&~m[337]&~m[339]&~m[340])|(m[335]&~m[336]&m[337]&~m[339]&~m[340])|(~m[335]&m[336]&m[337]&~m[339]&~m[340])|(m[335]&m[336]&m[337]&~m[339]&~m[340])|(m[335]&~m[336]&~m[337]&~m[339]&m[340])|(~m[335]&m[336]&~m[337]&~m[339]&m[340])|(m[335]&m[336]&~m[337]&~m[339]&m[340])|(~m[335]&~m[336]&m[337]&~m[339]&m[340])|(m[335]&~m[336]&m[337]&~m[339]&m[340])|(~m[335]&m[336]&m[337]&~m[339]&m[340])|(m[335]&m[336]&m[337]&~m[339]&m[340])|(m[335]&m[336]&m[337]&m[339]&m[340]))):InitCond[413];
    m[348] = run?((((m[345]&~m[346]&~m[347]&~m[349]&~m[350])|(~m[345]&m[346]&~m[347]&~m[349]&~m[350])|(~m[345]&~m[346]&m[347]&~m[349]&~m[350])|(m[345]&m[346]&m[347]&m[349]&~m[350])|(~m[345]&~m[346]&~m[347]&~m[349]&m[350])|(m[345]&m[346]&~m[347]&m[349]&m[350])|(m[345]&~m[346]&m[347]&m[349]&m[350])|(~m[345]&m[346]&m[347]&m[349]&m[350]))&UnbiasedRNG[191])|((m[345]&m[346]&~m[347]&~m[349]&~m[350])|(m[345]&~m[346]&m[347]&~m[349]&~m[350])|(~m[345]&m[346]&m[347]&~m[349]&~m[350])|(m[345]&m[346]&m[347]&~m[349]&~m[350])|(m[345]&~m[346]&~m[347]&~m[349]&m[350])|(~m[345]&m[346]&~m[347]&~m[349]&m[350])|(m[345]&m[346]&~m[347]&~m[349]&m[350])|(~m[345]&~m[346]&m[347]&~m[349]&m[350])|(m[345]&~m[346]&m[347]&~m[349]&m[350])|(~m[345]&m[346]&m[347]&~m[349]&m[350])|(m[345]&m[346]&m[347]&~m[349]&m[350])|(m[345]&m[346]&m[347]&m[349]&m[350]))):InitCond[414];
    m[353] = run?((((m[350]&~m[351]&~m[352]&~m[354]&~m[355])|(~m[350]&m[351]&~m[352]&~m[354]&~m[355])|(~m[350]&~m[351]&m[352]&~m[354]&~m[355])|(m[350]&m[351]&m[352]&m[354]&~m[355])|(~m[350]&~m[351]&~m[352]&~m[354]&m[355])|(m[350]&m[351]&~m[352]&m[354]&m[355])|(m[350]&~m[351]&m[352]&m[354]&m[355])|(~m[350]&m[351]&m[352]&m[354]&m[355]))&UnbiasedRNG[192])|((m[350]&m[351]&~m[352]&~m[354]&~m[355])|(m[350]&~m[351]&m[352]&~m[354]&~m[355])|(~m[350]&m[351]&m[352]&~m[354]&~m[355])|(m[350]&m[351]&m[352]&~m[354]&~m[355])|(m[350]&~m[351]&~m[352]&~m[354]&m[355])|(~m[350]&m[351]&~m[352]&~m[354]&m[355])|(m[350]&m[351]&~m[352]&~m[354]&m[355])|(~m[350]&~m[351]&m[352]&~m[354]&m[355])|(m[350]&~m[351]&m[352]&~m[354]&m[355])|(~m[350]&m[351]&m[352]&~m[354]&m[355])|(m[350]&m[351]&m[352]&~m[354]&m[355])|(m[350]&m[351]&m[352]&m[354]&m[355]))):InitCond[415];
    m[358] = run?((((m[355]&~m[356]&~m[357]&~m[359]&~m[360])|(~m[355]&m[356]&~m[357]&~m[359]&~m[360])|(~m[355]&~m[356]&m[357]&~m[359]&~m[360])|(m[355]&m[356]&m[357]&m[359]&~m[360])|(~m[355]&~m[356]&~m[357]&~m[359]&m[360])|(m[355]&m[356]&~m[357]&m[359]&m[360])|(m[355]&~m[356]&m[357]&m[359]&m[360])|(~m[355]&m[356]&m[357]&m[359]&m[360]))&UnbiasedRNG[193])|((m[355]&m[356]&~m[357]&~m[359]&~m[360])|(m[355]&~m[356]&m[357]&~m[359]&~m[360])|(~m[355]&m[356]&m[357]&~m[359]&~m[360])|(m[355]&m[356]&m[357]&~m[359]&~m[360])|(m[355]&~m[356]&~m[357]&~m[359]&m[360])|(~m[355]&m[356]&~m[357]&~m[359]&m[360])|(m[355]&m[356]&~m[357]&~m[359]&m[360])|(~m[355]&~m[356]&m[357]&~m[359]&m[360])|(m[355]&~m[356]&m[357]&~m[359]&m[360])|(~m[355]&m[356]&m[357]&~m[359]&m[360])|(m[355]&m[356]&m[357]&~m[359]&m[360])|(m[355]&m[356]&m[357]&m[359]&m[360]))):InitCond[416];
    m[363] = run?((((m[360]&~m[361]&~m[362]&~m[364]&~m[365])|(~m[360]&m[361]&~m[362]&~m[364]&~m[365])|(~m[360]&~m[361]&m[362]&~m[364]&~m[365])|(m[360]&m[361]&m[362]&m[364]&~m[365])|(~m[360]&~m[361]&~m[362]&~m[364]&m[365])|(m[360]&m[361]&~m[362]&m[364]&m[365])|(m[360]&~m[361]&m[362]&m[364]&m[365])|(~m[360]&m[361]&m[362]&m[364]&m[365]))&UnbiasedRNG[194])|((m[360]&m[361]&~m[362]&~m[364]&~m[365])|(m[360]&~m[361]&m[362]&~m[364]&~m[365])|(~m[360]&m[361]&m[362]&~m[364]&~m[365])|(m[360]&m[361]&m[362]&~m[364]&~m[365])|(m[360]&~m[361]&~m[362]&~m[364]&m[365])|(~m[360]&m[361]&~m[362]&~m[364]&m[365])|(m[360]&m[361]&~m[362]&~m[364]&m[365])|(~m[360]&~m[361]&m[362]&~m[364]&m[365])|(m[360]&~m[361]&m[362]&~m[364]&m[365])|(~m[360]&m[361]&m[362]&~m[364]&m[365])|(m[360]&m[361]&m[362]&~m[364]&m[365])|(m[360]&m[361]&m[362]&m[364]&m[365]))):InitCond[417];
    m[368] = run?((((m[365]&~m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&~m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&m[369]&~m[370])|(~m[365]&~m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&m[369]&m[370])|(m[365]&~m[366]&m[367]&m[369]&m[370])|(~m[365]&m[366]&m[367]&m[369]&m[370]))&UnbiasedRNG[195])|((m[365]&m[366]&~m[367]&~m[369]&~m[370])|(m[365]&~m[366]&m[367]&~m[369]&~m[370])|(~m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&~m[366]&~m[367]&~m[369]&m[370])|(~m[365]&m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&~m[369]&m[370])|(~m[365]&~m[366]&m[367]&~m[369]&m[370])|(m[365]&~m[366]&m[367]&~m[369]&m[370])|(~m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&m[369]&m[370]))):InitCond[418];
    m[373] = run?((((m[370]&~m[371]&~m[372]&~m[374]&~m[375])|(~m[370]&m[371]&~m[372]&~m[374]&~m[375])|(~m[370]&~m[371]&m[372]&~m[374]&~m[375])|(m[370]&m[371]&m[372]&m[374]&~m[375])|(~m[370]&~m[371]&~m[372]&~m[374]&m[375])|(m[370]&m[371]&~m[372]&m[374]&m[375])|(m[370]&~m[371]&m[372]&m[374]&m[375])|(~m[370]&m[371]&m[372]&m[374]&m[375]))&UnbiasedRNG[196])|((m[370]&m[371]&~m[372]&~m[374]&~m[375])|(m[370]&~m[371]&m[372]&~m[374]&~m[375])|(~m[370]&m[371]&m[372]&~m[374]&~m[375])|(m[370]&m[371]&m[372]&~m[374]&~m[375])|(m[370]&~m[371]&~m[372]&~m[374]&m[375])|(~m[370]&m[371]&~m[372]&~m[374]&m[375])|(m[370]&m[371]&~m[372]&~m[374]&m[375])|(~m[370]&~m[371]&m[372]&~m[374]&m[375])|(m[370]&~m[371]&m[372]&~m[374]&m[375])|(~m[370]&m[371]&m[372]&~m[374]&m[375])|(m[370]&m[371]&m[372]&~m[374]&m[375])|(m[370]&m[371]&m[372]&m[374]&m[375]))):InitCond[419];
    m[383] = run?((((m[380]&~m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&~m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&m[384]&~m[385])|(~m[380]&~m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&m[384]&m[385])|(m[380]&~m[381]&m[382]&m[384]&m[385])|(~m[380]&m[381]&m[382]&m[384]&m[385]))&UnbiasedRNG[197])|((m[380]&m[381]&~m[382]&~m[384]&~m[385])|(m[380]&~m[381]&m[382]&~m[384]&~m[385])|(~m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&~m[381]&~m[382]&~m[384]&m[385])|(~m[380]&m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&~m[384]&m[385])|(~m[380]&~m[381]&m[382]&~m[384]&m[385])|(m[380]&~m[381]&m[382]&~m[384]&m[385])|(~m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&m[384]&m[385]))):InitCond[420];
    m[388] = run?((((m[385]&~m[386]&~m[387]&~m[389]&~m[390])|(~m[385]&m[386]&~m[387]&~m[389]&~m[390])|(~m[385]&~m[386]&m[387]&~m[389]&~m[390])|(m[385]&m[386]&m[387]&m[389]&~m[390])|(~m[385]&~m[386]&~m[387]&~m[389]&m[390])|(m[385]&m[386]&~m[387]&m[389]&m[390])|(m[385]&~m[386]&m[387]&m[389]&m[390])|(~m[385]&m[386]&m[387]&m[389]&m[390]))&UnbiasedRNG[198])|((m[385]&m[386]&~m[387]&~m[389]&~m[390])|(m[385]&~m[386]&m[387]&~m[389]&~m[390])|(~m[385]&m[386]&m[387]&~m[389]&~m[390])|(m[385]&m[386]&m[387]&~m[389]&~m[390])|(m[385]&~m[386]&~m[387]&~m[389]&m[390])|(~m[385]&m[386]&~m[387]&~m[389]&m[390])|(m[385]&m[386]&~m[387]&~m[389]&m[390])|(~m[385]&~m[386]&m[387]&~m[389]&m[390])|(m[385]&~m[386]&m[387]&~m[389]&m[390])|(~m[385]&m[386]&m[387]&~m[389]&m[390])|(m[385]&m[386]&m[387]&~m[389]&m[390])|(m[385]&m[386]&m[387]&m[389]&m[390]))):InitCond[421];
    m[393] = run?((((m[390]&~m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&~m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&m[394]&~m[395])|(~m[390]&~m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&m[394]&m[395])|(m[390]&~m[391]&m[392]&m[394]&m[395])|(~m[390]&m[391]&m[392]&m[394]&m[395]))&UnbiasedRNG[199])|((m[390]&m[391]&~m[392]&~m[394]&~m[395])|(m[390]&~m[391]&m[392]&~m[394]&~m[395])|(~m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&~m[391]&~m[392]&~m[394]&m[395])|(~m[390]&m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&~m[394]&m[395])|(~m[390]&~m[391]&m[392]&~m[394]&m[395])|(m[390]&~m[391]&m[392]&~m[394]&m[395])|(~m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&m[394]&m[395]))):InitCond[422];
    m[398] = run?((((m[395]&~m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&~m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&m[399]&~m[400])|(~m[395]&~m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&m[399]&m[400])|(m[395]&~m[396]&m[397]&m[399]&m[400])|(~m[395]&m[396]&m[397]&m[399]&m[400]))&UnbiasedRNG[200])|((m[395]&m[396]&~m[397]&~m[399]&~m[400])|(m[395]&~m[396]&m[397]&~m[399]&~m[400])|(~m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&~m[396]&~m[397]&~m[399]&m[400])|(~m[395]&m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&~m[399]&m[400])|(~m[395]&~m[396]&m[397]&~m[399]&m[400])|(m[395]&~m[396]&m[397]&~m[399]&m[400])|(~m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&m[399]&m[400]))):InitCond[423];
    m[403] = run?((((m[400]&~m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&~m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&m[404]&~m[405])|(~m[400]&~m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&m[404]&m[405])|(m[400]&~m[401]&m[402]&m[404]&m[405])|(~m[400]&m[401]&m[402]&m[404]&m[405]))&UnbiasedRNG[201])|((m[400]&m[401]&~m[402]&~m[404]&~m[405])|(m[400]&~m[401]&m[402]&~m[404]&~m[405])|(~m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&~m[401]&~m[402]&~m[404]&m[405])|(~m[400]&m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&~m[404]&m[405])|(~m[400]&~m[401]&m[402]&~m[404]&m[405])|(m[400]&~m[401]&m[402]&~m[404]&m[405])|(~m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&m[404]&m[405]))):InitCond[424];
    m[408] = run?((((m[405]&~m[406]&~m[407]&~m[409]&~m[410])|(~m[405]&m[406]&~m[407]&~m[409]&~m[410])|(~m[405]&~m[406]&m[407]&~m[409]&~m[410])|(m[405]&m[406]&m[407]&m[409]&~m[410])|(~m[405]&~m[406]&~m[407]&~m[409]&m[410])|(m[405]&m[406]&~m[407]&m[409]&m[410])|(m[405]&~m[406]&m[407]&m[409]&m[410])|(~m[405]&m[406]&m[407]&m[409]&m[410]))&UnbiasedRNG[202])|((m[405]&m[406]&~m[407]&~m[409]&~m[410])|(m[405]&~m[406]&m[407]&~m[409]&~m[410])|(~m[405]&m[406]&m[407]&~m[409]&~m[410])|(m[405]&m[406]&m[407]&~m[409]&~m[410])|(m[405]&~m[406]&~m[407]&~m[409]&m[410])|(~m[405]&m[406]&~m[407]&~m[409]&m[410])|(m[405]&m[406]&~m[407]&~m[409]&m[410])|(~m[405]&~m[406]&m[407]&~m[409]&m[410])|(m[405]&~m[406]&m[407]&~m[409]&m[410])|(~m[405]&m[406]&m[407]&~m[409]&m[410])|(m[405]&m[406]&m[407]&~m[409]&m[410])|(m[405]&m[406]&m[407]&m[409]&m[410]))):InitCond[425];
    m[418] = run?((((m[415]&~m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&~m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&m[419]&~m[420])|(~m[415]&~m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&m[419]&m[420])|(m[415]&~m[416]&m[417]&m[419]&m[420])|(~m[415]&m[416]&m[417]&m[419]&m[420]))&UnbiasedRNG[203])|((m[415]&m[416]&~m[417]&~m[419]&~m[420])|(m[415]&~m[416]&m[417]&~m[419]&~m[420])|(~m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&~m[416]&~m[417]&~m[419]&m[420])|(~m[415]&m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&~m[419]&m[420])|(~m[415]&~m[416]&m[417]&~m[419]&m[420])|(m[415]&~m[416]&m[417]&~m[419]&m[420])|(~m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&m[419]&m[420]))):InitCond[426];
    m[423] = run?((((m[420]&~m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&~m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&m[424]&~m[425])|(~m[420]&~m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&m[424]&m[425])|(m[420]&~m[421]&m[422]&m[424]&m[425])|(~m[420]&m[421]&m[422]&m[424]&m[425]))&UnbiasedRNG[204])|((m[420]&m[421]&~m[422]&~m[424]&~m[425])|(m[420]&~m[421]&m[422]&~m[424]&~m[425])|(~m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&~m[421]&~m[422]&~m[424]&m[425])|(~m[420]&m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&~m[424]&m[425])|(~m[420]&~m[421]&m[422]&~m[424]&m[425])|(m[420]&~m[421]&m[422]&~m[424]&m[425])|(~m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&m[424]&m[425]))):InitCond[427];
    m[428] = run?((((m[425]&~m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&~m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&m[429]&~m[430])|(~m[425]&~m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&m[429]&m[430])|(m[425]&~m[426]&m[427]&m[429]&m[430])|(~m[425]&m[426]&m[427]&m[429]&m[430]))&UnbiasedRNG[205])|((m[425]&m[426]&~m[427]&~m[429]&~m[430])|(m[425]&~m[426]&m[427]&~m[429]&~m[430])|(~m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&~m[426]&~m[427]&~m[429]&m[430])|(~m[425]&m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&~m[429]&m[430])|(~m[425]&~m[426]&m[427]&~m[429]&m[430])|(m[425]&~m[426]&m[427]&~m[429]&m[430])|(~m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&m[429]&m[430]))):InitCond[428];
    m[433] = run?((((m[430]&~m[431]&~m[432]&~m[434]&~m[435])|(~m[430]&m[431]&~m[432]&~m[434]&~m[435])|(~m[430]&~m[431]&m[432]&~m[434]&~m[435])|(m[430]&m[431]&m[432]&m[434]&~m[435])|(~m[430]&~m[431]&~m[432]&~m[434]&m[435])|(m[430]&m[431]&~m[432]&m[434]&m[435])|(m[430]&~m[431]&m[432]&m[434]&m[435])|(~m[430]&m[431]&m[432]&m[434]&m[435]))&UnbiasedRNG[206])|((m[430]&m[431]&~m[432]&~m[434]&~m[435])|(m[430]&~m[431]&m[432]&~m[434]&~m[435])|(~m[430]&m[431]&m[432]&~m[434]&~m[435])|(m[430]&m[431]&m[432]&~m[434]&~m[435])|(m[430]&~m[431]&~m[432]&~m[434]&m[435])|(~m[430]&m[431]&~m[432]&~m[434]&m[435])|(m[430]&m[431]&~m[432]&~m[434]&m[435])|(~m[430]&~m[431]&m[432]&~m[434]&m[435])|(m[430]&~m[431]&m[432]&~m[434]&m[435])|(~m[430]&m[431]&m[432]&~m[434]&m[435])|(m[430]&m[431]&m[432]&~m[434]&m[435])|(m[430]&m[431]&m[432]&m[434]&m[435]))):InitCond[429];
    m[438] = run?((((m[435]&~m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&~m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&m[439]&~m[440])|(~m[435]&~m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&m[439]&m[440])|(m[435]&~m[436]&m[437]&m[439]&m[440])|(~m[435]&m[436]&m[437]&m[439]&m[440]))&UnbiasedRNG[207])|((m[435]&m[436]&~m[437]&~m[439]&~m[440])|(m[435]&~m[436]&m[437]&~m[439]&~m[440])|(~m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&~m[436]&~m[437]&~m[439]&m[440])|(~m[435]&m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&~m[439]&m[440])|(~m[435]&~m[436]&m[437]&~m[439]&m[440])|(m[435]&~m[436]&m[437]&~m[439]&m[440])|(~m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&m[439]&m[440]))):InitCond[430];
    m[448] = run?((((m[445]&~m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&~m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&m[449]&~m[450])|(~m[445]&~m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&m[449]&m[450])|(m[445]&~m[446]&m[447]&m[449]&m[450])|(~m[445]&m[446]&m[447]&m[449]&m[450]))&UnbiasedRNG[208])|((m[445]&m[446]&~m[447]&~m[449]&~m[450])|(m[445]&~m[446]&m[447]&~m[449]&~m[450])|(~m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&~m[446]&~m[447]&~m[449]&m[450])|(~m[445]&m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&~m[449]&m[450])|(~m[445]&~m[446]&m[447]&~m[449]&m[450])|(m[445]&~m[446]&m[447]&~m[449]&m[450])|(~m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&m[449]&m[450]))):InitCond[431];
    m[453] = run?((((m[450]&~m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&~m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&m[454]&~m[455])|(~m[450]&~m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&m[454]&m[455])|(m[450]&~m[451]&m[452]&m[454]&m[455])|(~m[450]&m[451]&m[452]&m[454]&m[455]))&UnbiasedRNG[209])|((m[450]&m[451]&~m[452]&~m[454]&~m[455])|(m[450]&~m[451]&m[452]&~m[454]&~m[455])|(~m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&~m[451]&~m[452]&~m[454]&m[455])|(~m[450]&m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&~m[454]&m[455])|(~m[450]&~m[451]&m[452]&~m[454]&m[455])|(m[450]&~m[451]&m[452]&~m[454]&m[455])|(~m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&m[454]&m[455]))):InitCond[432];
    m[458] = run?((((m[455]&~m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&~m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&m[459]&~m[460])|(~m[455]&~m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&m[459]&m[460])|(m[455]&~m[456]&m[457]&m[459]&m[460])|(~m[455]&m[456]&m[457]&m[459]&m[460]))&UnbiasedRNG[210])|((m[455]&m[456]&~m[457]&~m[459]&~m[460])|(m[455]&~m[456]&m[457]&~m[459]&~m[460])|(~m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&~m[456]&~m[457]&~m[459]&m[460])|(~m[455]&m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&~m[459]&m[460])|(~m[455]&~m[456]&m[457]&~m[459]&m[460])|(m[455]&~m[456]&m[457]&~m[459]&m[460])|(~m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&m[459]&m[460]))):InitCond[433];
    m[463] = run?((((m[460]&~m[461]&~m[462]&~m[464]&~m[465])|(~m[460]&m[461]&~m[462]&~m[464]&~m[465])|(~m[460]&~m[461]&m[462]&~m[464]&~m[465])|(m[460]&m[461]&m[462]&m[464]&~m[465])|(~m[460]&~m[461]&~m[462]&~m[464]&m[465])|(m[460]&m[461]&~m[462]&m[464]&m[465])|(m[460]&~m[461]&m[462]&m[464]&m[465])|(~m[460]&m[461]&m[462]&m[464]&m[465]))&UnbiasedRNG[211])|((m[460]&m[461]&~m[462]&~m[464]&~m[465])|(m[460]&~m[461]&m[462]&~m[464]&~m[465])|(~m[460]&m[461]&m[462]&~m[464]&~m[465])|(m[460]&m[461]&m[462]&~m[464]&~m[465])|(m[460]&~m[461]&~m[462]&~m[464]&m[465])|(~m[460]&m[461]&~m[462]&~m[464]&m[465])|(m[460]&m[461]&~m[462]&~m[464]&m[465])|(~m[460]&~m[461]&m[462]&~m[464]&m[465])|(m[460]&~m[461]&m[462]&~m[464]&m[465])|(~m[460]&m[461]&m[462]&~m[464]&m[465])|(m[460]&m[461]&m[462]&~m[464]&m[465])|(m[460]&m[461]&m[462]&m[464]&m[465]))):InitCond[434];
    m[473] = run?((((m[470]&~m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&~m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&m[474]&~m[475])|(~m[470]&~m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&m[474]&m[475])|(m[470]&~m[471]&m[472]&m[474]&m[475])|(~m[470]&m[471]&m[472]&m[474]&m[475]))&UnbiasedRNG[212])|((m[470]&m[471]&~m[472]&~m[474]&~m[475])|(m[470]&~m[471]&m[472]&~m[474]&~m[475])|(~m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&~m[471]&~m[472]&~m[474]&m[475])|(~m[470]&m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&~m[474]&m[475])|(~m[470]&~m[471]&m[472]&~m[474]&m[475])|(m[470]&~m[471]&m[472]&~m[474]&m[475])|(~m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&m[474]&m[475]))):InitCond[435];
    m[478] = run?((((m[475]&~m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&~m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&m[479]&~m[480])|(~m[475]&~m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&m[479]&m[480])|(m[475]&~m[476]&m[477]&m[479]&m[480])|(~m[475]&m[476]&m[477]&m[479]&m[480]))&UnbiasedRNG[213])|((m[475]&m[476]&~m[477]&~m[479]&~m[480])|(m[475]&~m[476]&m[477]&~m[479]&~m[480])|(~m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&~m[476]&~m[477]&~m[479]&m[480])|(~m[475]&m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&~m[479]&m[480])|(~m[475]&~m[476]&m[477]&~m[479]&m[480])|(m[475]&~m[476]&m[477]&~m[479]&m[480])|(~m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&m[479]&m[480]))):InitCond[436];
    m[483] = run?((((m[480]&~m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&~m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&m[484]&~m[485])|(~m[480]&~m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&m[484]&m[485])|(m[480]&~m[481]&m[482]&m[484]&m[485])|(~m[480]&m[481]&m[482]&m[484]&m[485]))&UnbiasedRNG[214])|((m[480]&m[481]&~m[482]&~m[484]&~m[485])|(m[480]&~m[481]&m[482]&~m[484]&~m[485])|(~m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&~m[481]&~m[482]&~m[484]&m[485])|(~m[480]&m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&~m[484]&m[485])|(~m[480]&~m[481]&m[482]&~m[484]&m[485])|(m[480]&~m[481]&m[482]&~m[484]&m[485])|(~m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&m[484]&m[485]))):InitCond[437];
    m[493] = run?((((m[490]&~m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&~m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&m[494]&~m[495])|(~m[490]&~m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&m[494]&m[495])|(m[490]&~m[491]&m[492]&m[494]&m[495])|(~m[490]&m[491]&m[492]&m[494]&m[495]))&UnbiasedRNG[215])|((m[490]&m[491]&~m[492]&~m[494]&~m[495])|(m[490]&~m[491]&m[492]&~m[494]&~m[495])|(~m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&~m[491]&~m[492]&~m[494]&m[495])|(~m[490]&m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&~m[494]&m[495])|(~m[490]&~m[491]&m[492]&~m[494]&m[495])|(m[490]&~m[491]&m[492]&~m[494]&m[495])|(~m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&m[494]&m[495]))):InitCond[438];
    m[498] = run?((((m[495]&~m[496]&~m[497]&~m[499]&~m[500])|(~m[495]&m[496]&~m[497]&~m[499]&~m[500])|(~m[495]&~m[496]&m[497]&~m[499]&~m[500])|(m[495]&m[496]&m[497]&m[499]&~m[500])|(~m[495]&~m[496]&~m[497]&~m[499]&m[500])|(m[495]&m[496]&~m[497]&m[499]&m[500])|(m[495]&~m[496]&m[497]&m[499]&m[500])|(~m[495]&m[496]&m[497]&m[499]&m[500]))&UnbiasedRNG[216])|((m[495]&m[496]&~m[497]&~m[499]&~m[500])|(m[495]&~m[496]&m[497]&~m[499]&~m[500])|(~m[495]&m[496]&m[497]&~m[499]&~m[500])|(m[495]&m[496]&m[497]&~m[499]&~m[500])|(m[495]&~m[496]&~m[497]&~m[499]&m[500])|(~m[495]&m[496]&~m[497]&~m[499]&m[500])|(m[495]&m[496]&~m[497]&~m[499]&m[500])|(~m[495]&~m[496]&m[497]&~m[499]&m[500])|(m[495]&~m[496]&m[497]&~m[499]&m[500])|(~m[495]&m[496]&m[497]&~m[499]&m[500])|(m[495]&m[496]&m[497]&~m[499]&m[500])|(m[495]&m[496]&m[497]&m[499]&m[500]))):InitCond[439];
    m[508] = run?((((m[505]&~m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&~m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&m[509]&~m[510])|(~m[505]&~m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&m[509]&m[510])|(m[505]&~m[506]&m[507]&m[509]&m[510])|(~m[505]&m[506]&m[507]&m[509]&m[510]))&UnbiasedRNG[217])|((m[505]&m[506]&~m[507]&~m[509]&~m[510])|(m[505]&~m[506]&m[507]&~m[509]&~m[510])|(~m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&~m[506]&~m[507]&~m[509]&m[510])|(~m[505]&m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&~m[509]&m[510])|(~m[505]&~m[506]&m[507]&~m[509]&m[510])|(m[505]&~m[506]&m[507]&~m[509]&m[510])|(~m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&m[509]&m[510]))):InitCond[440];
end

always @(posedge color4_clk) begin
    m[244] = run?((((m[240]&~m[241]&~m[242]&~m[243]&~m[247])|(~m[240]&m[241]&~m[242]&~m[243]&~m[247])|(~m[240]&~m[241]&m[242]&~m[243]&~m[247])|(m[240]&m[241]&~m[242]&m[243]&~m[247])|(m[240]&~m[241]&m[242]&m[243]&~m[247])|(~m[240]&m[241]&m[242]&m[243]&~m[247]))&BiasedRNG[223])|(((m[240]&~m[241]&~m[242]&~m[243]&m[247])|(~m[240]&m[241]&~m[242]&~m[243]&m[247])|(~m[240]&~m[241]&m[242]&~m[243]&m[247])|(m[240]&m[241]&~m[242]&m[243]&m[247])|(m[240]&~m[241]&m[242]&m[243]&m[247])|(~m[240]&m[241]&m[242]&m[243]&m[247]))&~BiasedRNG[223])|((m[240]&m[241]&~m[242]&~m[243]&~m[247])|(m[240]&~m[241]&m[242]&~m[243]&~m[247])|(~m[240]&m[241]&m[242]&~m[243]&~m[247])|(m[240]&m[241]&m[242]&~m[243]&~m[247])|(m[240]&m[241]&m[242]&m[243]&~m[247])|(m[240]&m[241]&~m[242]&~m[243]&m[247])|(m[240]&~m[241]&m[242]&~m[243]&m[247])|(~m[240]&m[241]&m[242]&~m[243]&m[247])|(m[240]&m[241]&m[242]&~m[243]&m[247])|(m[240]&m[241]&m[242]&m[243]&m[247]))):InitCond[441];
    m[249] = run?((((m[245]&~m[246]&~m[247]&~m[248]&~m[257])|(~m[245]&m[246]&~m[247]&~m[248]&~m[257])|(~m[245]&~m[246]&m[247]&~m[248]&~m[257])|(m[245]&m[246]&~m[247]&m[248]&~m[257])|(m[245]&~m[246]&m[247]&m[248]&~m[257])|(~m[245]&m[246]&m[247]&m[248]&~m[257]))&BiasedRNG[224])|(((m[245]&~m[246]&~m[247]&~m[248]&m[257])|(~m[245]&m[246]&~m[247]&~m[248]&m[257])|(~m[245]&~m[246]&m[247]&~m[248]&m[257])|(m[245]&m[246]&~m[247]&m[248]&m[257])|(m[245]&~m[246]&m[247]&m[248]&m[257])|(~m[245]&m[246]&m[247]&m[248]&m[257]))&~BiasedRNG[224])|((m[245]&m[246]&~m[247]&~m[248]&~m[257])|(m[245]&~m[246]&m[247]&~m[248]&~m[257])|(~m[245]&m[246]&m[247]&~m[248]&~m[257])|(m[245]&m[246]&m[247]&~m[248]&~m[257])|(m[245]&m[246]&m[247]&m[248]&~m[257])|(m[245]&m[246]&~m[247]&~m[248]&m[257])|(m[245]&~m[246]&m[247]&~m[248]&m[257])|(~m[245]&m[246]&m[247]&~m[248]&m[257])|(m[245]&m[246]&m[247]&~m[248]&m[257])|(m[245]&m[246]&m[247]&m[248]&m[257]))):InitCond[442];
    m[254] = run?((((m[250]&~m[251]&~m[252]&~m[253]&~m[262])|(~m[250]&m[251]&~m[252]&~m[253]&~m[262])|(~m[250]&~m[251]&m[252]&~m[253]&~m[262])|(m[250]&m[251]&~m[252]&m[253]&~m[262])|(m[250]&~m[251]&m[252]&m[253]&~m[262])|(~m[250]&m[251]&m[252]&m[253]&~m[262]))&BiasedRNG[225])|(((m[250]&~m[251]&~m[252]&~m[253]&m[262])|(~m[250]&m[251]&~m[252]&~m[253]&m[262])|(~m[250]&~m[251]&m[252]&~m[253]&m[262])|(m[250]&m[251]&~m[252]&m[253]&m[262])|(m[250]&~m[251]&m[252]&m[253]&m[262])|(~m[250]&m[251]&m[252]&m[253]&m[262]))&~BiasedRNG[225])|((m[250]&m[251]&~m[252]&~m[253]&~m[262])|(m[250]&~m[251]&m[252]&~m[253]&~m[262])|(~m[250]&m[251]&m[252]&~m[253]&~m[262])|(m[250]&m[251]&m[252]&~m[253]&~m[262])|(m[250]&m[251]&m[252]&m[253]&~m[262])|(m[250]&m[251]&~m[252]&~m[253]&m[262])|(m[250]&~m[251]&m[252]&~m[253]&m[262])|(~m[250]&m[251]&m[252]&~m[253]&m[262])|(m[250]&m[251]&m[252]&~m[253]&m[262])|(m[250]&m[251]&m[252]&m[253]&m[262]))):InitCond[443];
    m[259] = run?((((m[255]&~m[256]&~m[257]&~m[258]&~m[272])|(~m[255]&m[256]&~m[257]&~m[258]&~m[272])|(~m[255]&~m[256]&m[257]&~m[258]&~m[272])|(m[255]&m[256]&~m[257]&m[258]&~m[272])|(m[255]&~m[256]&m[257]&m[258]&~m[272])|(~m[255]&m[256]&m[257]&m[258]&~m[272]))&BiasedRNG[226])|(((m[255]&~m[256]&~m[257]&~m[258]&m[272])|(~m[255]&m[256]&~m[257]&~m[258]&m[272])|(~m[255]&~m[256]&m[257]&~m[258]&m[272])|(m[255]&m[256]&~m[257]&m[258]&m[272])|(m[255]&~m[256]&m[257]&m[258]&m[272])|(~m[255]&m[256]&m[257]&m[258]&m[272]))&~BiasedRNG[226])|((m[255]&m[256]&~m[257]&~m[258]&~m[272])|(m[255]&~m[256]&m[257]&~m[258]&~m[272])|(~m[255]&m[256]&m[257]&~m[258]&~m[272])|(m[255]&m[256]&m[257]&~m[258]&~m[272])|(m[255]&m[256]&m[257]&m[258]&~m[272])|(m[255]&m[256]&~m[257]&~m[258]&m[272])|(m[255]&~m[256]&m[257]&~m[258]&m[272])|(~m[255]&m[256]&m[257]&~m[258]&m[272])|(m[255]&m[256]&m[257]&~m[258]&m[272])|(m[255]&m[256]&m[257]&m[258]&m[272]))):InitCond[444];
    m[264] = run?((((m[260]&~m[261]&~m[262]&~m[263]&~m[277])|(~m[260]&m[261]&~m[262]&~m[263]&~m[277])|(~m[260]&~m[261]&m[262]&~m[263]&~m[277])|(m[260]&m[261]&~m[262]&m[263]&~m[277])|(m[260]&~m[261]&m[262]&m[263]&~m[277])|(~m[260]&m[261]&m[262]&m[263]&~m[277]))&BiasedRNG[227])|(((m[260]&~m[261]&~m[262]&~m[263]&m[277])|(~m[260]&m[261]&~m[262]&~m[263]&m[277])|(~m[260]&~m[261]&m[262]&~m[263]&m[277])|(m[260]&m[261]&~m[262]&m[263]&m[277])|(m[260]&~m[261]&m[262]&m[263]&m[277])|(~m[260]&m[261]&m[262]&m[263]&m[277]))&~BiasedRNG[227])|((m[260]&m[261]&~m[262]&~m[263]&~m[277])|(m[260]&~m[261]&m[262]&~m[263]&~m[277])|(~m[260]&m[261]&m[262]&~m[263]&~m[277])|(m[260]&m[261]&m[262]&~m[263]&~m[277])|(m[260]&m[261]&m[262]&m[263]&~m[277])|(m[260]&m[261]&~m[262]&~m[263]&m[277])|(m[260]&~m[261]&m[262]&~m[263]&m[277])|(~m[260]&m[261]&m[262]&~m[263]&m[277])|(m[260]&m[261]&m[262]&~m[263]&m[277])|(m[260]&m[261]&m[262]&m[263]&m[277]))):InitCond[445];
    m[269] = run?((((m[265]&~m[266]&~m[267]&~m[268]&~m[282])|(~m[265]&m[266]&~m[267]&~m[268]&~m[282])|(~m[265]&~m[266]&m[267]&~m[268]&~m[282])|(m[265]&m[266]&~m[267]&m[268]&~m[282])|(m[265]&~m[266]&m[267]&m[268]&~m[282])|(~m[265]&m[266]&m[267]&m[268]&~m[282]))&BiasedRNG[228])|(((m[265]&~m[266]&~m[267]&~m[268]&m[282])|(~m[265]&m[266]&~m[267]&~m[268]&m[282])|(~m[265]&~m[266]&m[267]&~m[268]&m[282])|(m[265]&m[266]&~m[267]&m[268]&m[282])|(m[265]&~m[266]&m[267]&m[268]&m[282])|(~m[265]&m[266]&m[267]&m[268]&m[282]))&~BiasedRNG[228])|((m[265]&m[266]&~m[267]&~m[268]&~m[282])|(m[265]&~m[266]&m[267]&~m[268]&~m[282])|(~m[265]&m[266]&m[267]&~m[268]&~m[282])|(m[265]&m[266]&m[267]&~m[268]&~m[282])|(m[265]&m[266]&m[267]&m[268]&~m[282])|(m[265]&m[266]&~m[267]&~m[268]&m[282])|(m[265]&~m[266]&m[267]&~m[268]&m[282])|(~m[265]&m[266]&m[267]&~m[268]&m[282])|(m[265]&m[266]&m[267]&~m[268]&m[282])|(m[265]&m[266]&m[267]&m[268]&m[282]))):InitCond[446];
    m[274] = run?((((m[270]&~m[271]&~m[272]&~m[273]&~m[292])|(~m[270]&m[271]&~m[272]&~m[273]&~m[292])|(~m[270]&~m[271]&m[272]&~m[273]&~m[292])|(m[270]&m[271]&~m[272]&m[273]&~m[292])|(m[270]&~m[271]&m[272]&m[273]&~m[292])|(~m[270]&m[271]&m[272]&m[273]&~m[292]))&BiasedRNG[229])|(((m[270]&~m[271]&~m[272]&~m[273]&m[292])|(~m[270]&m[271]&~m[272]&~m[273]&m[292])|(~m[270]&~m[271]&m[272]&~m[273]&m[292])|(m[270]&m[271]&~m[272]&m[273]&m[292])|(m[270]&~m[271]&m[272]&m[273]&m[292])|(~m[270]&m[271]&m[272]&m[273]&m[292]))&~BiasedRNG[229])|((m[270]&m[271]&~m[272]&~m[273]&~m[292])|(m[270]&~m[271]&m[272]&~m[273]&~m[292])|(~m[270]&m[271]&m[272]&~m[273]&~m[292])|(m[270]&m[271]&m[272]&~m[273]&~m[292])|(m[270]&m[271]&m[272]&m[273]&~m[292])|(m[270]&m[271]&~m[272]&~m[273]&m[292])|(m[270]&~m[271]&m[272]&~m[273]&m[292])|(~m[270]&m[271]&m[272]&~m[273]&m[292])|(m[270]&m[271]&m[272]&~m[273]&m[292])|(m[270]&m[271]&m[272]&m[273]&m[292]))):InitCond[447];
    m[279] = run?((((m[275]&~m[276]&~m[277]&~m[278]&~m[297])|(~m[275]&m[276]&~m[277]&~m[278]&~m[297])|(~m[275]&~m[276]&m[277]&~m[278]&~m[297])|(m[275]&m[276]&~m[277]&m[278]&~m[297])|(m[275]&~m[276]&m[277]&m[278]&~m[297])|(~m[275]&m[276]&m[277]&m[278]&~m[297]))&BiasedRNG[230])|(((m[275]&~m[276]&~m[277]&~m[278]&m[297])|(~m[275]&m[276]&~m[277]&~m[278]&m[297])|(~m[275]&~m[276]&m[277]&~m[278]&m[297])|(m[275]&m[276]&~m[277]&m[278]&m[297])|(m[275]&~m[276]&m[277]&m[278]&m[297])|(~m[275]&m[276]&m[277]&m[278]&m[297]))&~BiasedRNG[230])|((m[275]&m[276]&~m[277]&~m[278]&~m[297])|(m[275]&~m[276]&m[277]&~m[278]&~m[297])|(~m[275]&m[276]&m[277]&~m[278]&~m[297])|(m[275]&m[276]&m[277]&~m[278]&~m[297])|(m[275]&m[276]&m[277]&m[278]&~m[297])|(m[275]&m[276]&~m[277]&~m[278]&m[297])|(m[275]&~m[276]&m[277]&~m[278]&m[297])|(~m[275]&m[276]&m[277]&~m[278]&m[297])|(m[275]&m[276]&m[277]&~m[278]&m[297])|(m[275]&m[276]&m[277]&m[278]&m[297]))):InitCond[448];
    m[284] = run?((((m[280]&~m[281]&~m[282]&~m[283]&~m[302])|(~m[280]&m[281]&~m[282]&~m[283]&~m[302])|(~m[280]&~m[281]&m[282]&~m[283]&~m[302])|(m[280]&m[281]&~m[282]&m[283]&~m[302])|(m[280]&~m[281]&m[282]&m[283]&~m[302])|(~m[280]&m[281]&m[282]&m[283]&~m[302]))&BiasedRNG[231])|(((m[280]&~m[281]&~m[282]&~m[283]&m[302])|(~m[280]&m[281]&~m[282]&~m[283]&m[302])|(~m[280]&~m[281]&m[282]&~m[283]&m[302])|(m[280]&m[281]&~m[282]&m[283]&m[302])|(m[280]&~m[281]&m[282]&m[283]&m[302])|(~m[280]&m[281]&m[282]&m[283]&m[302]))&~BiasedRNG[231])|((m[280]&m[281]&~m[282]&~m[283]&~m[302])|(m[280]&~m[281]&m[282]&~m[283]&~m[302])|(~m[280]&m[281]&m[282]&~m[283]&~m[302])|(m[280]&m[281]&m[282]&~m[283]&~m[302])|(m[280]&m[281]&m[282]&m[283]&~m[302])|(m[280]&m[281]&~m[282]&~m[283]&m[302])|(m[280]&~m[281]&m[282]&~m[283]&m[302])|(~m[280]&m[281]&m[282]&~m[283]&m[302])|(m[280]&m[281]&m[282]&~m[283]&m[302])|(m[280]&m[281]&m[282]&m[283]&m[302]))):InitCond[449];
    m[289] = run?((((m[285]&~m[286]&~m[287]&~m[288]&~m[307])|(~m[285]&m[286]&~m[287]&~m[288]&~m[307])|(~m[285]&~m[286]&m[287]&~m[288]&~m[307])|(m[285]&m[286]&~m[287]&m[288]&~m[307])|(m[285]&~m[286]&m[287]&m[288]&~m[307])|(~m[285]&m[286]&m[287]&m[288]&~m[307]))&BiasedRNG[232])|(((m[285]&~m[286]&~m[287]&~m[288]&m[307])|(~m[285]&m[286]&~m[287]&~m[288]&m[307])|(~m[285]&~m[286]&m[287]&~m[288]&m[307])|(m[285]&m[286]&~m[287]&m[288]&m[307])|(m[285]&~m[286]&m[287]&m[288]&m[307])|(~m[285]&m[286]&m[287]&m[288]&m[307]))&~BiasedRNG[232])|((m[285]&m[286]&~m[287]&~m[288]&~m[307])|(m[285]&~m[286]&m[287]&~m[288]&~m[307])|(~m[285]&m[286]&m[287]&~m[288]&~m[307])|(m[285]&m[286]&m[287]&~m[288]&~m[307])|(m[285]&m[286]&m[287]&m[288]&~m[307])|(m[285]&m[286]&~m[287]&~m[288]&m[307])|(m[285]&~m[286]&m[287]&~m[288]&m[307])|(~m[285]&m[286]&m[287]&~m[288]&m[307])|(m[285]&m[286]&m[287]&~m[288]&m[307])|(m[285]&m[286]&m[287]&m[288]&m[307]))):InitCond[450];
    m[294] = run?((((m[290]&~m[291]&~m[292]&~m[293]&~m[317])|(~m[290]&m[291]&~m[292]&~m[293]&~m[317])|(~m[290]&~m[291]&m[292]&~m[293]&~m[317])|(m[290]&m[291]&~m[292]&m[293]&~m[317])|(m[290]&~m[291]&m[292]&m[293]&~m[317])|(~m[290]&m[291]&m[292]&m[293]&~m[317]))&BiasedRNG[233])|(((m[290]&~m[291]&~m[292]&~m[293]&m[317])|(~m[290]&m[291]&~m[292]&~m[293]&m[317])|(~m[290]&~m[291]&m[292]&~m[293]&m[317])|(m[290]&m[291]&~m[292]&m[293]&m[317])|(m[290]&~m[291]&m[292]&m[293]&m[317])|(~m[290]&m[291]&m[292]&m[293]&m[317]))&~BiasedRNG[233])|((m[290]&m[291]&~m[292]&~m[293]&~m[317])|(m[290]&~m[291]&m[292]&~m[293]&~m[317])|(~m[290]&m[291]&m[292]&~m[293]&~m[317])|(m[290]&m[291]&m[292]&~m[293]&~m[317])|(m[290]&m[291]&m[292]&m[293]&~m[317])|(m[290]&m[291]&~m[292]&~m[293]&m[317])|(m[290]&~m[291]&m[292]&~m[293]&m[317])|(~m[290]&m[291]&m[292]&~m[293]&m[317])|(m[290]&m[291]&m[292]&~m[293]&m[317])|(m[290]&m[291]&m[292]&m[293]&m[317]))):InitCond[451];
    m[299] = run?((((m[295]&~m[296]&~m[297]&~m[298]&~m[322])|(~m[295]&m[296]&~m[297]&~m[298]&~m[322])|(~m[295]&~m[296]&m[297]&~m[298]&~m[322])|(m[295]&m[296]&~m[297]&m[298]&~m[322])|(m[295]&~m[296]&m[297]&m[298]&~m[322])|(~m[295]&m[296]&m[297]&m[298]&~m[322]))&BiasedRNG[234])|(((m[295]&~m[296]&~m[297]&~m[298]&m[322])|(~m[295]&m[296]&~m[297]&~m[298]&m[322])|(~m[295]&~m[296]&m[297]&~m[298]&m[322])|(m[295]&m[296]&~m[297]&m[298]&m[322])|(m[295]&~m[296]&m[297]&m[298]&m[322])|(~m[295]&m[296]&m[297]&m[298]&m[322]))&~BiasedRNG[234])|((m[295]&m[296]&~m[297]&~m[298]&~m[322])|(m[295]&~m[296]&m[297]&~m[298]&~m[322])|(~m[295]&m[296]&m[297]&~m[298]&~m[322])|(m[295]&m[296]&m[297]&~m[298]&~m[322])|(m[295]&m[296]&m[297]&m[298]&~m[322])|(m[295]&m[296]&~m[297]&~m[298]&m[322])|(m[295]&~m[296]&m[297]&~m[298]&m[322])|(~m[295]&m[296]&m[297]&~m[298]&m[322])|(m[295]&m[296]&m[297]&~m[298]&m[322])|(m[295]&m[296]&m[297]&m[298]&m[322]))):InitCond[452];
    m[304] = run?((((m[300]&~m[301]&~m[302]&~m[303]&~m[327])|(~m[300]&m[301]&~m[302]&~m[303]&~m[327])|(~m[300]&~m[301]&m[302]&~m[303]&~m[327])|(m[300]&m[301]&~m[302]&m[303]&~m[327])|(m[300]&~m[301]&m[302]&m[303]&~m[327])|(~m[300]&m[301]&m[302]&m[303]&~m[327]))&BiasedRNG[235])|(((m[300]&~m[301]&~m[302]&~m[303]&m[327])|(~m[300]&m[301]&~m[302]&~m[303]&m[327])|(~m[300]&~m[301]&m[302]&~m[303]&m[327])|(m[300]&m[301]&~m[302]&m[303]&m[327])|(m[300]&~m[301]&m[302]&m[303]&m[327])|(~m[300]&m[301]&m[302]&m[303]&m[327]))&~BiasedRNG[235])|((m[300]&m[301]&~m[302]&~m[303]&~m[327])|(m[300]&~m[301]&m[302]&~m[303]&~m[327])|(~m[300]&m[301]&m[302]&~m[303]&~m[327])|(m[300]&m[301]&m[302]&~m[303]&~m[327])|(m[300]&m[301]&m[302]&m[303]&~m[327])|(m[300]&m[301]&~m[302]&~m[303]&m[327])|(m[300]&~m[301]&m[302]&~m[303]&m[327])|(~m[300]&m[301]&m[302]&~m[303]&m[327])|(m[300]&m[301]&m[302]&~m[303]&m[327])|(m[300]&m[301]&m[302]&m[303]&m[327]))):InitCond[453];
    m[309] = run?((((m[305]&~m[306]&~m[307]&~m[308]&~m[332])|(~m[305]&m[306]&~m[307]&~m[308]&~m[332])|(~m[305]&~m[306]&m[307]&~m[308]&~m[332])|(m[305]&m[306]&~m[307]&m[308]&~m[332])|(m[305]&~m[306]&m[307]&m[308]&~m[332])|(~m[305]&m[306]&m[307]&m[308]&~m[332]))&BiasedRNG[236])|(((m[305]&~m[306]&~m[307]&~m[308]&m[332])|(~m[305]&m[306]&~m[307]&~m[308]&m[332])|(~m[305]&~m[306]&m[307]&~m[308]&m[332])|(m[305]&m[306]&~m[307]&m[308]&m[332])|(m[305]&~m[306]&m[307]&m[308]&m[332])|(~m[305]&m[306]&m[307]&m[308]&m[332]))&~BiasedRNG[236])|((m[305]&m[306]&~m[307]&~m[308]&~m[332])|(m[305]&~m[306]&m[307]&~m[308]&~m[332])|(~m[305]&m[306]&m[307]&~m[308]&~m[332])|(m[305]&m[306]&m[307]&~m[308]&~m[332])|(m[305]&m[306]&m[307]&m[308]&~m[332])|(m[305]&m[306]&~m[307]&~m[308]&m[332])|(m[305]&~m[306]&m[307]&~m[308]&m[332])|(~m[305]&m[306]&m[307]&~m[308]&m[332])|(m[305]&m[306]&m[307]&~m[308]&m[332])|(m[305]&m[306]&m[307]&m[308]&m[332]))):InitCond[454];
    m[314] = run?((((m[310]&~m[311]&~m[312]&~m[313]&~m[337])|(~m[310]&m[311]&~m[312]&~m[313]&~m[337])|(~m[310]&~m[311]&m[312]&~m[313]&~m[337])|(m[310]&m[311]&~m[312]&m[313]&~m[337])|(m[310]&~m[311]&m[312]&m[313]&~m[337])|(~m[310]&m[311]&m[312]&m[313]&~m[337]))&BiasedRNG[237])|(((m[310]&~m[311]&~m[312]&~m[313]&m[337])|(~m[310]&m[311]&~m[312]&~m[313]&m[337])|(~m[310]&~m[311]&m[312]&~m[313]&m[337])|(m[310]&m[311]&~m[312]&m[313]&m[337])|(m[310]&~m[311]&m[312]&m[313]&m[337])|(~m[310]&m[311]&m[312]&m[313]&m[337]))&~BiasedRNG[237])|((m[310]&m[311]&~m[312]&~m[313]&~m[337])|(m[310]&~m[311]&m[312]&~m[313]&~m[337])|(~m[310]&m[311]&m[312]&~m[313]&~m[337])|(m[310]&m[311]&m[312]&~m[313]&~m[337])|(m[310]&m[311]&m[312]&m[313]&~m[337])|(m[310]&m[311]&~m[312]&~m[313]&m[337])|(m[310]&~m[311]&m[312]&~m[313]&m[337])|(~m[310]&m[311]&m[312]&~m[313]&m[337])|(m[310]&m[311]&m[312]&~m[313]&m[337])|(m[310]&m[311]&m[312]&m[313]&m[337]))):InitCond[455];
    m[319] = run?((((m[315]&~m[316]&~m[317]&~m[318]&~m[347])|(~m[315]&m[316]&~m[317]&~m[318]&~m[347])|(~m[315]&~m[316]&m[317]&~m[318]&~m[347])|(m[315]&m[316]&~m[317]&m[318]&~m[347])|(m[315]&~m[316]&m[317]&m[318]&~m[347])|(~m[315]&m[316]&m[317]&m[318]&~m[347]))&BiasedRNG[238])|(((m[315]&~m[316]&~m[317]&~m[318]&m[347])|(~m[315]&m[316]&~m[317]&~m[318]&m[347])|(~m[315]&~m[316]&m[317]&~m[318]&m[347])|(m[315]&m[316]&~m[317]&m[318]&m[347])|(m[315]&~m[316]&m[317]&m[318]&m[347])|(~m[315]&m[316]&m[317]&m[318]&m[347]))&~BiasedRNG[238])|((m[315]&m[316]&~m[317]&~m[318]&~m[347])|(m[315]&~m[316]&m[317]&~m[318]&~m[347])|(~m[315]&m[316]&m[317]&~m[318]&~m[347])|(m[315]&m[316]&m[317]&~m[318]&~m[347])|(m[315]&m[316]&m[317]&m[318]&~m[347])|(m[315]&m[316]&~m[317]&~m[318]&m[347])|(m[315]&~m[316]&m[317]&~m[318]&m[347])|(~m[315]&m[316]&m[317]&~m[318]&m[347])|(m[315]&m[316]&m[317]&~m[318]&m[347])|(m[315]&m[316]&m[317]&m[318]&m[347]))):InitCond[456];
    m[324] = run?((((m[320]&~m[321]&~m[322]&~m[323]&~m[352])|(~m[320]&m[321]&~m[322]&~m[323]&~m[352])|(~m[320]&~m[321]&m[322]&~m[323]&~m[352])|(m[320]&m[321]&~m[322]&m[323]&~m[352])|(m[320]&~m[321]&m[322]&m[323]&~m[352])|(~m[320]&m[321]&m[322]&m[323]&~m[352]))&BiasedRNG[239])|(((m[320]&~m[321]&~m[322]&~m[323]&m[352])|(~m[320]&m[321]&~m[322]&~m[323]&m[352])|(~m[320]&~m[321]&m[322]&~m[323]&m[352])|(m[320]&m[321]&~m[322]&m[323]&m[352])|(m[320]&~m[321]&m[322]&m[323]&m[352])|(~m[320]&m[321]&m[322]&m[323]&m[352]))&~BiasedRNG[239])|((m[320]&m[321]&~m[322]&~m[323]&~m[352])|(m[320]&~m[321]&m[322]&~m[323]&~m[352])|(~m[320]&m[321]&m[322]&~m[323]&~m[352])|(m[320]&m[321]&m[322]&~m[323]&~m[352])|(m[320]&m[321]&m[322]&m[323]&~m[352])|(m[320]&m[321]&~m[322]&~m[323]&m[352])|(m[320]&~m[321]&m[322]&~m[323]&m[352])|(~m[320]&m[321]&m[322]&~m[323]&m[352])|(m[320]&m[321]&m[322]&~m[323]&m[352])|(m[320]&m[321]&m[322]&m[323]&m[352]))):InitCond[457];
    m[329] = run?((((m[325]&~m[326]&~m[327]&~m[328]&~m[357])|(~m[325]&m[326]&~m[327]&~m[328]&~m[357])|(~m[325]&~m[326]&m[327]&~m[328]&~m[357])|(m[325]&m[326]&~m[327]&m[328]&~m[357])|(m[325]&~m[326]&m[327]&m[328]&~m[357])|(~m[325]&m[326]&m[327]&m[328]&~m[357]))&BiasedRNG[240])|(((m[325]&~m[326]&~m[327]&~m[328]&m[357])|(~m[325]&m[326]&~m[327]&~m[328]&m[357])|(~m[325]&~m[326]&m[327]&~m[328]&m[357])|(m[325]&m[326]&~m[327]&m[328]&m[357])|(m[325]&~m[326]&m[327]&m[328]&m[357])|(~m[325]&m[326]&m[327]&m[328]&m[357]))&~BiasedRNG[240])|((m[325]&m[326]&~m[327]&~m[328]&~m[357])|(m[325]&~m[326]&m[327]&~m[328]&~m[357])|(~m[325]&m[326]&m[327]&~m[328]&~m[357])|(m[325]&m[326]&m[327]&~m[328]&~m[357])|(m[325]&m[326]&m[327]&m[328]&~m[357])|(m[325]&m[326]&~m[327]&~m[328]&m[357])|(m[325]&~m[326]&m[327]&~m[328]&m[357])|(~m[325]&m[326]&m[327]&~m[328]&m[357])|(m[325]&m[326]&m[327]&~m[328]&m[357])|(m[325]&m[326]&m[327]&m[328]&m[357]))):InitCond[458];
    m[334] = run?((((m[330]&~m[331]&~m[332]&~m[333]&~m[362])|(~m[330]&m[331]&~m[332]&~m[333]&~m[362])|(~m[330]&~m[331]&m[332]&~m[333]&~m[362])|(m[330]&m[331]&~m[332]&m[333]&~m[362])|(m[330]&~m[331]&m[332]&m[333]&~m[362])|(~m[330]&m[331]&m[332]&m[333]&~m[362]))&BiasedRNG[241])|(((m[330]&~m[331]&~m[332]&~m[333]&m[362])|(~m[330]&m[331]&~m[332]&~m[333]&m[362])|(~m[330]&~m[331]&m[332]&~m[333]&m[362])|(m[330]&m[331]&~m[332]&m[333]&m[362])|(m[330]&~m[331]&m[332]&m[333]&m[362])|(~m[330]&m[331]&m[332]&m[333]&m[362]))&~BiasedRNG[241])|((m[330]&m[331]&~m[332]&~m[333]&~m[362])|(m[330]&~m[331]&m[332]&~m[333]&~m[362])|(~m[330]&m[331]&m[332]&~m[333]&~m[362])|(m[330]&m[331]&m[332]&~m[333]&~m[362])|(m[330]&m[331]&m[332]&m[333]&~m[362])|(m[330]&m[331]&~m[332]&~m[333]&m[362])|(m[330]&~m[331]&m[332]&~m[333]&m[362])|(~m[330]&m[331]&m[332]&~m[333]&m[362])|(m[330]&m[331]&m[332]&~m[333]&m[362])|(m[330]&m[331]&m[332]&m[333]&m[362]))):InitCond[459];
    m[339] = run?((((m[335]&~m[336]&~m[337]&~m[338]&~m[367])|(~m[335]&m[336]&~m[337]&~m[338]&~m[367])|(~m[335]&~m[336]&m[337]&~m[338]&~m[367])|(m[335]&m[336]&~m[337]&m[338]&~m[367])|(m[335]&~m[336]&m[337]&m[338]&~m[367])|(~m[335]&m[336]&m[337]&m[338]&~m[367]))&BiasedRNG[242])|(((m[335]&~m[336]&~m[337]&~m[338]&m[367])|(~m[335]&m[336]&~m[337]&~m[338]&m[367])|(~m[335]&~m[336]&m[337]&~m[338]&m[367])|(m[335]&m[336]&~m[337]&m[338]&m[367])|(m[335]&~m[336]&m[337]&m[338]&m[367])|(~m[335]&m[336]&m[337]&m[338]&m[367]))&~BiasedRNG[242])|((m[335]&m[336]&~m[337]&~m[338]&~m[367])|(m[335]&~m[336]&m[337]&~m[338]&~m[367])|(~m[335]&m[336]&m[337]&~m[338]&~m[367])|(m[335]&m[336]&m[337]&~m[338]&~m[367])|(m[335]&m[336]&m[337]&m[338]&~m[367])|(m[335]&m[336]&~m[337]&~m[338]&m[367])|(m[335]&~m[336]&m[337]&~m[338]&m[367])|(~m[335]&m[336]&m[337]&~m[338]&m[367])|(m[335]&m[336]&m[337]&~m[338]&m[367])|(m[335]&m[336]&m[337]&m[338]&m[367]))):InitCond[460];
    m[344] = run?((((m[340]&~m[341]&~m[342]&~m[343]&~m[372])|(~m[340]&m[341]&~m[342]&~m[343]&~m[372])|(~m[340]&~m[341]&m[342]&~m[343]&~m[372])|(m[340]&m[341]&~m[342]&m[343]&~m[372])|(m[340]&~m[341]&m[342]&m[343]&~m[372])|(~m[340]&m[341]&m[342]&m[343]&~m[372]))&BiasedRNG[243])|(((m[340]&~m[341]&~m[342]&~m[343]&m[372])|(~m[340]&m[341]&~m[342]&~m[343]&m[372])|(~m[340]&~m[341]&m[342]&~m[343]&m[372])|(m[340]&m[341]&~m[342]&m[343]&m[372])|(m[340]&~m[341]&m[342]&m[343]&m[372])|(~m[340]&m[341]&m[342]&m[343]&m[372]))&~BiasedRNG[243])|((m[340]&m[341]&~m[342]&~m[343]&~m[372])|(m[340]&~m[341]&m[342]&~m[343]&~m[372])|(~m[340]&m[341]&m[342]&~m[343]&~m[372])|(m[340]&m[341]&m[342]&~m[343]&~m[372])|(m[340]&m[341]&m[342]&m[343]&~m[372])|(m[340]&m[341]&~m[342]&~m[343]&m[372])|(m[340]&~m[341]&m[342]&~m[343]&m[372])|(~m[340]&m[341]&m[342]&~m[343]&m[372])|(m[340]&m[341]&m[342]&~m[343]&m[372])|(m[340]&m[341]&m[342]&m[343]&m[372]))):InitCond[461];
    m[349] = run?((((m[345]&~m[346]&~m[347]&~m[348]&~m[382])|(~m[345]&m[346]&~m[347]&~m[348]&~m[382])|(~m[345]&~m[346]&m[347]&~m[348]&~m[382])|(m[345]&m[346]&~m[347]&m[348]&~m[382])|(m[345]&~m[346]&m[347]&m[348]&~m[382])|(~m[345]&m[346]&m[347]&m[348]&~m[382]))&BiasedRNG[244])|(((m[345]&~m[346]&~m[347]&~m[348]&m[382])|(~m[345]&m[346]&~m[347]&~m[348]&m[382])|(~m[345]&~m[346]&m[347]&~m[348]&m[382])|(m[345]&m[346]&~m[347]&m[348]&m[382])|(m[345]&~m[346]&m[347]&m[348]&m[382])|(~m[345]&m[346]&m[347]&m[348]&m[382]))&~BiasedRNG[244])|((m[345]&m[346]&~m[347]&~m[348]&~m[382])|(m[345]&~m[346]&m[347]&~m[348]&~m[382])|(~m[345]&m[346]&m[347]&~m[348]&~m[382])|(m[345]&m[346]&m[347]&~m[348]&~m[382])|(m[345]&m[346]&m[347]&m[348]&~m[382])|(m[345]&m[346]&~m[347]&~m[348]&m[382])|(m[345]&~m[346]&m[347]&~m[348]&m[382])|(~m[345]&m[346]&m[347]&~m[348]&m[382])|(m[345]&m[346]&m[347]&~m[348]&m[382])|(m[345]&m[346]&m[347]&m[348]&m[382]))):InitCond[462];
    m[354] = run?((((m[350]&~m[351]&~m[352]&~m[353]&~m[387])|(~m[350]&m[351]&~m[352]&~m[353]&~m[387])|(~m[350]&~m[351]&m[352]&~m[353]&~m[387])|(m[350]&m[351]&~m[352]&m[353]&~m[387])|(m[350]&~m[351]&m[352]&m[353]&~m[387])|(~m[350]&m[351]&m[352]&m[353]&~m[387]))&BiasedRNG[245])|(((m[350]&~m[351]&~m[352]&~m[353]&m[387])|(~m[350]&m[351]&~m[352]&~m[353]&m[387])|(~m[350]&~m[351]&m[352]&~m[353]&m[387])|(m[350]&m[351]&~m[352]&m[353]&m[387])|(m[350]&~m[351]&m[352]&m[353]&m[387])|(~m[350]&m[351]&m[352]&m[353]&m[387]))&~BiasedRNG[245])|((m[350]&m[351]&~m[352]&~m[353]&~m[387])|(m[350]&~m[351]&m[352]&~m[353]&~m[387])|(~m[350]&m[351]&m[352]&~m[353]&~m[387])|(m[350]&m[351]&m[352]&~m[353]&~m[387])|(m[350]&m[351]&m[352]&m[353]&~m[387])|(m[350]&m[351]&~m[352]&~m[353]&m[387])|(m[350]&~m[351]&m[352]&~m[353]&m[387])|(~m[350]&m[351]&m[352]&~m[353]&m[387])|(m[350]&m[351]&m[352]&~m[353]&m[387])|(m[350]&m[351]&m[352]&m[353]&m[387]))):InitCond[463];
    m[359] = run?((((m[355]&~m[356]&~m[357]&~m[358]&~m[392])|(~m[355]&m[356]&~m[357]&~m[358]&~m[392])|(~m[355]&~m[356]&m[357]&~m[358]&~m[392])|(m[355]&m[356]&~m[357]&m[358]&~m[392])|(m[355]&~m[356]&m[357]&m[358]&~m[392])|(~m[355]&m[356]&m[357]&m[358]&~m[392]))&BiasedRNG[246])|(((m[355]&~m[356]&~m[357]&~m[358]&m[392])|(~m[355]&m[356]&~m[357]&~m[358]&m[392])|(~m[355]&~m[356]&m[357]&~m[358]&m[392])|(m[355]&m[356]&~m[357]&m[358]&m[392])|(m[355]&~m[356]&m[357]&m[358]&m[392])|(~m[355]&m[356]&m[357]&m[358]&m[392]))&~BiasedRNG[246])|((m[355]&m[356]&~m[357]&~m[358]&~m[392])|(m[355]&~m[356]&m[357]&~m[358]&~m[392])|(~m[355]&m[356]&m[357]&~m[358]&~m[392])|(m[355]&m[356]&m[357]&~m[358]&~m[392])|(m[355]&m[356]&m[357]&m[358]&~m[392])|(m[355]&m[356]&~m[357]&~m[358]&m[392])|(m[355]&~m[356]&m[357]&~m[358]&m[392])|(~m[355]&m[356]&m[357]&~m[358]&m[392])|(m[355]&m[356]&m[357]&~m[358]&m[392])|(m[355]&m[356]&m[357]&m[358]&m[392]))):InitCond[464];
    m[364] = run?((((m[360]&~m[361]&~m[362]&~m[363]&~m[397])|(~m[360]&m[361]&~m[362]&~m[363]&~m[397])|(~m[360]&~m[361]&m[362]&~m[363]&~m[397])|(m[360]&m[361]&~m[362]&m[363]&~m[397])|(m[360]&~m[361]&m[362]&m[363]&~m[397])|(~m[360]&m[361]&m[362]&m[363]&~m[397]))&BiasedRNG[247])|(((m[360]&~m[361]&~m[362]&~m[363]&m[397])|(~m[360]&m[361]&~m[362]&~m[363]&m[397])|(~m[360]&~m[361]&m[362]&~m[363]&m[397])|(m[360]&m[361]&~m[362]&m[363]&m[397])|(m[360]&~m[361]&m[362]&m[363]&m[397])|(~m[360]&m[361]&m[362]&m[363]&m[397]))&~BiasedRNG[247])|((m[360]&m[361]&~m[362]&~m[363]&~m[397])|(m[360]&~m[361]&m[362]&~m[363]&~m[397])|(~m[360]&m[361]&m[362]&~m[363]&~m[397])|(m[360]&m[361]&m[362]&~m[363]&~m[397])|(m[360]&m[361]&m[362]&m[363]&~m[397])|(m[360]&m[361]&~m[362]&~m[363]&m[397])|(m[360]&~m[361]&m[362]&~m[363]&m[397])|(~m[360]&m[361]&m[362]&~m[363]&m[397])|(m[360]&m[361]&m[362]&~m[363]&m[397])|(m[360]&m[361]&m[362]&m[363]&m[397]))):InitCond[465];
    m[369] = run?((((m[365]&~m[366]&~m[367]&~m[368]&~m[402])|(~m[365]&m[366]&~m[367]&~m[368]&~m[402])|(~m[365]&~m[366]&m[367]&~m[368]&~m[402])|(m[365]&m[366]&~m[367]&m[368]&~m[402])|(m[365]&~m[366]&m[367]&m[368]&~m[402])|(~m[365]&m[366]&m[367]&m[368]&~m[402]))&BiasedRNG[248])|(((m[365]&~m[366]&~m[367]&~m[368]&m[402])|(~m[365]&m[366]&~m[367]&~m[368]&m[402])|(~m[365]&~m[366]&m[367]&~m[368]&m[402])|(m[365]&m[366]&~m[367]&m[368]&m[402])|(m[365]&~m[366]&m[367]&m[368]&m[402])|(~m[365]&m[366]&m[367]&m[368]&m[402]))&~BiasedRNG[248])|((m[365]&m[366]&~m[367]&~m[368]&~m[402])|(m[365]&~m[366]&m[367]&~m[368]&~m[402])|(~m[365]&m[366]&m[367]&~m[368]&~m[402])|(m[365]&m[366]&m[367]&~m[368]&~m[402])|(m[365]&m[366]&m[367]&m[368]&~m[402])|(m[365]&m[366]&~m[367]&~m[368]&m[402])|(m[365]&~m[366]&m[367]&~m[368]&m[402])|(~m[365]&m[366]&m[367]&~m[368]&m[402])|(m[365]&m[366]&m[367]&~m[368]&m[402])|(m[365]&m[366]&m[367]&m[368]&m[402]))):InitCond[466];
    m[374] = run?((((m[370]&~m[371]&~m[372]&~m[373]&~m[407])|(~m[370]&m[371]&~m[372]&~m[373]&~m[407])|(~m[370]&~m[371]&m[372]&~m[373]&~m[407])|(m[370]&m[371]&~m[372]&m[373]&~m[407])|(m[370]&~m[371]&m[372]&m[373]&~m[407])|(~m[370]&m[371]&m[372]&m[373]&~m[407]))&BiasedRNG[249])|(((m[370]&~m[371]&~m[372]&~m[373]&m[407])|(~m[370]&m[371]&~m[372]&~m[373]&m[407])|(~m[370]&~m[371]&m[372]&~m[373]&m[407])|(m[370]&m[371]&~m[372]&m[373]&m[407])|(m[370]&~m[371]&m[372]&m[373]&m[407])|(~m[370]&m[371]&m[372]&m[373]&m[407]))&~BiasedRNG[249])|((m[370]&m[371]&~m[372]&~m[373]&~m[407])|(m[370]&~m[371]&m[372]&~m[373]&~m[407])|(~m[370]&m[371]&m[372]&~m[373]&~m[407])|(m[370]&m[371]&m[372]&~m[373]&~m[407])|(m[370]&m[371]&m[372]&m[373]&~m[407])|(m[370]&m[371]&~m[372]&~m[373]&m[407])|(m[370]&~m[371]&m[372]&~m[373]&m[407])|(~m[370]&m[371]&m[372]&~m[373]&m[407])|(m[370]&m[371]&m[372]&~m[373]&m[407])|(m[370]&m[371]&m[372]&m[373]&m[407]))):InitCond[467];
    m[379] = run?((((m[375]&~m[376]&~m[377]&~m[378]&~m[412])|(~m[375]&m[376]&~m[377]&~m[378]&~m[412])|(~m[375]&~m[376]&m[377]&~m[378]&~m[412])|(m[375]&m[376]&~m[377]&m[378]&~m[412])|(m[375]&~m[376]&m[377]&m[378]&~m[412])|(~m[375]&m[376]&m[377]&m[378]&~m[412]))&BiasedRNG[250])|(((m[375]&~m[376]&~m[377]&~m[378]&m[412])|(~m[375]&m[376]&~m[377]&~m[378]&m[412])|(~m[375]&~m[376]&m[377]&~m[378]&m[412])|(m[375]&m[376]&~m[377]&m[378]&m[412])|(m[375]&~m[376]&m[377]&m[378]&m[412])|(~m[375]&m[376]&m[377]&m[378]&m[412]))&~BiasedRNG[250])|((m[375]&m[376]&~m[377]&~m[378]&~m[412])|(m[375]&~m[376]&m[377]&~m[378]&~m[412])|(~m[375]&m[376]&m[377]&~m[378]&~m[412])|(m[375]&m[376]&m[377]&~m[378]&~m[412])|(m[375]&m[376]&m[377]&m[378]&~m[412])|(m[375]&m[376]&~m[377]&~m[378]&m[412])|(m[375]&~m[376]&m[377]&~m[378]&m[412])|(~m[375]&m[376]&m[377]&~m[378]&m[412])|(m[375]&m[376]&m[377]&~m[378]&m[412])|(m[375]&m[376]&m[377]&m[378]&m[412]))):InitCond[468];
    m[384] = run?((((m[380]&~m[381]&~m[382]&~m[383]&~m[415])|(~m[380]&m[381]&~m[382]&~m[383]&~m[415])|(~m[380]&~m[381]&m[382]&~m[383]&~m[415])|(m[380]&m[381]&~m[382]&m[383]&~m[415])|(m[380]&~m[381]&m[382]&m[383]&~m[415])|(~m[380]&m[381]&m[382]&m[383]&~m[415]))&BiasedRNG[251])|(((m[380]&~m[381]&~m[382]&~m[383]&m[415])|(~m[380]&m[381]&~m[382]&~m[383]&m[415])|(~m[380]&~m[381]&m[382]&~m[383]&m[415])|(m[380]&m[381]&~m[382]&m[383]&m[415])|(m[380]&~m[381]&m[382]&m[383]&m[415])|(~m[380]&m[381]&m[382]&m[383]&m[415]))&~BiasedRNG[251])|((m[380]&m[381]&~m[382]&~m[383]&~m[415])|(m[380]&~m[381]&m[382]&~m[383]&~m[415])|(~m[380]&m[381]&m[382]&~m[383]&~m[415])|(m[380]&m[381]&m[382]&~m[383]&~m[415])|(m[380]&m[381]&m[382]&m[383]&~m[415])|(m[380]&m[381]&~m[382]&~m[383]&m[415])|(m[380]&~m[381]&m[382]&~m[383]&m[415])|(~m[380]&m[381]&m[382]&~m[383]&m[415])|(m[380]&m[381]&m[382]&~m[383]&m[415])|(m[380]&m[381]&m[382]&m[383]&m[415]))):InitCond[469];
    m[389] = run?((((m[385]&~m[386]&~m[387]&~m[388]&~m[417])|(~m[385]&m[386]&~m[387]&~m[388]&~m[417])|(~m[385]&~m[386]&m[387]&~m[388]&~m[417])|(m[385]&m[386]&~m[387]&m[388]&~m[417])|(m[385]&~m[386]&m[387]&m[388]&~m[417])|(~m[385]&m[386]&m[387]&m[388]&~m[417]))&BiasedRNG[252])|(((m[385]&~m[386]&~m[387]&~m[388]&m[417])|(~m[385]&m[386]&~m[387]&~m[388]&m[417])|(~m[385]&~m[386]&m[387]&~m[388]&m[417])|(m[385]&m[386]&~m[387]&m[388]&m[417])|(m[385]&~m[386]&m[387]&m[388]&m[417])|(~m[385]&m[386]&m[387]&m[388]&m[417]))&~BiasedRNG[252])|((m[385]&m[386]&~m[387]&~m[388]&~m[417])|(m[385]&~m[386]&m[387]&~m[388]&~m[417])|(~m[385]&m[386]&m[387]&~m[388]&~m[417])|(m[385]&m[386]&m[387]&~m[388]&~m[417])|(m[385]&m[386]&m[387]&m[388]&~m[417])|(m[385]&m[386]&~m[387]&~m[388]&m[417])|(m[385]&~m[386]&m[387]&~m[388]&m[417])|(~m[385]&m[386]&m[387]&~m[388]&m[417])|(m[385]&m[386]&m[387]&~m[388]&m[417])|(m[385]&m[386]&m[387]&m[388]&m[417]))):InitCond[470];
    m[394] = run?((((m[390]&~m[391]&~m[392]&~m[393]&~m[422])|(~m[390]&m[391]&~m[392]&~m[393]&~m[422])|(~m[390]&~m[391]&m[392]&~m[393]&~m[422])|(m[390]&m[391]&~m[392]&m[393]&~m[422])|(m[390]&~m[391]&m[392]&m[393]&~m[422])|(~m[390]&m[391]&m[392]&m[393]&~m[422]))&BiasedRNG[253])|(((m[390]&~m[391]&~m[392]&~m[393]&m[422])|(~m[390]&m[391]&~m[392]&~m[393]&m[422])|(~m[390]&~m[391]&m[392]&~m[393]&m[422])|(m[390]&m[391]&~m[392]&m[393]&m[422])|(m[390]&~m[391]&m[392]&m[393]&m[422])|(~m[390]&m[391]&m[392]&m[393]&m[422]))&~BiasedRNG[253])|((m[390]&m[391]&~m[392]&~m[393]&~m[422])|(m[390]&~m[391]&m[392]&~m[393]&~m[422])|(~m[390]&m[391]&m[392]&~m[393]&~m[422])|(m[390]&m[391]&m[392]&~m[393]&~m[422])|(m[390]&m[391]&m[392]&m[393]&~m[422])|(m[390]&m[391]&~m[392]&~m[393]&m[422])|(m[390]&~m[391]&m[392]&~m[393]&m[422])|(~m[390]&m[391]&m[392]&~m[393]&m[422])|(m[390]&m[391]&m[392]&~m[393]&m[422])|(m[390]&m[391]&m[392]&m[393]&m[422]))):InitCond[471];
    m[399] = run?((((m[395]&~m[396]&~m[397]&~m[398]&~m[427])|(~m[395]&m[396]&~m[397]&~m[398]&~m[427])|(~m[395]&~m[396]&m[397]&~m[398]&~m[427])|(m[395]&m[396]&~m[397]&m[398]&~m[427])|(m[395]&~m[396]&m[397]&m[398]&~m[427])|(~m[395]&m[396]&m[397]&m[398]&~m[427]))&BiasedRNG[254])|(((m[395]&~m[396]&~m[397]&~m[398]&m[427])|(~m[395]&m[396]&~m[397]&~m[398]&m[427])|(~m[395]&~m[396]&m[397]&~m[398]&m[427])|(m[395]&m[396]&~m[397]&m[398]&m[427])|(m[395]&~m[396]&m[397]&m[398]&m[427])|(~m[395]&m[396]&m[397]&m[398]&m[427]))&~BiasedRNG[254])|((m[395]&m[396]&~m[397]&~m[398]&~m[427])|(m[395]&~m[396]&m[397]&~m[398]&~m[427])|(~m[395]&m[396]&m[397]&~m[398]&~m[427])|(m[395]&m[396]&m[397]&~m[398]&~m[427])|(m[395]&m[396]&m[397]&m[398]&~m[427])|(m[395]&m[396]&~m[397]&~m[398]&m[427])|(m[395]&~m[396]&m[397]&~m[398]&m[427])|(~m[395]&m[396]&m[397]&~m[398]&m[427])|(m[395]&m[396]&m[397]&~m[398]&m[427])|(m[395]&m[396]&m[397]&m[398]&m[427]))):InitCond[472];
    m[404] = run?((((m[400]&~m[401]&~m[402]&~m[403]&~m[432])|(~m[400]&m[401]&~m[402]&~m[403]&~m[432])|(~m[400]&~m[401]&m[402]&~m[403]&~m[432])|(m[400]&m[401]&~m[402]&m[403]&~m[432])|(m[400]&~m[401]&m[402]&m[403]&~m[432])|(~m[400]&m[401]&m[402]&m[403]&~m[432]))&BiasedRNG[255])|(((m[400]&~m[401]&~m[402]&~m[403]&m[432])|(~m[400]&m[401]&~m[402]&~m[403]&m[432])|(~m[400]&~m[401]&m[402]&~m[403]&m[432])|(m[400]&m[401]&~m[402]&m[403]&m[432])|(m[400]&~m[401]&m[402]&m[403]&m[432])|(~m[400]&m[401]&m[402]&m[403]&m[432]))&~BiasedRNG[255])|((m[400]&m[401]&~m[402]&~m[403]&~m[432])|(m[400]&~m[401]&m[402]&~m[403]&~m[432])|(~m[400]&m[401]&m[402]&~m[403]&~m[432])|(m[400]&m[401]&m[402]&~m[403]&~m[432])|(m[400]&m[401]&m[402]&m[403]&~m[432])|(m[400]&m[401]&~m[402]&~m[403]&m[432])|(m[400]&~m[401]&m[402]&~m[403]&m[432])|(~m[400]&m[401]&m[402]&~m[403]&m[432])|(m[400]&m[401]&m[402]&~m[403]&m[432])|(m[400]&m[401]&m[402]&m[403]&m[432]))):InitCond[473];
    m[409] = run?((((m[405]&~m[406]&~m[407]&~m[408]&~m[437])|(~m[405]&m[406]&~m[407]&~m[408]&~m[437])|(~m[405]&~m[406]&m[407]&~m[408]&~m[437])|(m[405]&m[406]&~m[407]&m[408]&~m[437])|(m[405]&~m[406]&m[407]&m[408]&~m[437])|(~m[405]&m[406]&m[407]&m[408]&~m[437]))&BiasedRNG[256])|(((m[405]&~m[406]&~m[407]&~m[408]&m[437])|(~m[405]&m[406]&~m[407]&~m[408]&m[437])|(~m[405]&~m[406]&m[407]&~m[408]&m[437])|(m[405]&m[406]&~m[407]&m[408]&m[437])|(m[405]&~m[406]&m[407]&m[408]&m[437])|(~m[405]&m[406]&m[407]&m[408]&m[437]))&~BiasedRNG[256])|((m[405]&m[406]&~m[407]&~m[408]&~m[437])|(m[405]&~m[406]&m[407]&~m[408]&~m[437])|(~m[405]&m[406]&m[407]&~m[408]&~m[437])|(m[405]&m[406]&m[407]&~m[408]&~m[437])|(m[405]&m[406]&m[407]&m[408]&~m[437])|(m[405]&m[406]&~m[407]&~m[408]&m[437])|(m[405]&~m[406]&m[407]&~m[408]&m[437])|(~m[405]&m[406]&m[407]&~m[408]&m[437])|(m[405]&m[406]&m[407]&~m[408]&m[437])|(m[405]&m[406]&m[407]&m[408]&m[437]))):InitCond[474];
    m[414] = run?((((m[410]&~m[411]&~m[412]&~m[413]&~m[442])|(~m[410]&m[411]&~m[412]&~m[413]&~m[442])|(~m[410]&~m[411]&m[412]&~m[413]&~m[442])|(m[410]&m[411]&~m[412]&m[413]&~m[442])|(m[410]&~m[411]&m[412]&m[413]&~m[442])|(~m[410]&m[411]&m[412]&m[413]&~m[442]))&BiasedRNG[257])|(((m[410]&~m[411]&~m[412]&~m[413]&m[442])|(~m[410]&m[411]&~m[412]&~m[413]&m[442])|(~m[410]&~m[411]&m[412]&~m[413]&m[442])|(m[410]&m[411]&~m[412]&m[413]&m[442])|(m[410]&~m[411]&m[412]&m[413]&m[442])|(~m[410]&m[411]&m[412]&m[413]&m[442]))&~BiasedRNG[257])|((m[410]&m[411]&~m[412]&~m[413]&~m[442])|(m[410]&~m[411]&m[412]&~m[413]&~m[442])|(~m[410]&m[411]&m[412]&~m[413]&~m[442])|(m[410]&m[411]&m[412]&~m[413]&~m[442])|(m[410]&m[411]&m[412]&m[413]&~m[442])|(m[410]&m[411]&~m[412]&~m[413]&m[442])|(m[410]&~m[411]&m[412]&~m[413]&m[442])|(~m[410]&m[411]&m[412]&~m[413]&m[442])|(m[410]&m[411]&m[412]&~m[413]&m[442])|(m[410]&m[411]&m[412]&m[413]&m[442]))):InitCond[475];
    m[419] = run?((((m[415]&~m[416]&~m[417]&~m[418]&~m[445])|(~m[415]&m[416]&~m[417]&~m[418]&~m[445])|(~m[415]&~m[416]&m[417]&~m[418]&~m[445])|(m[415]&m[416]&~m[417]&m[418]&~m[445])|(m[415]&~m[416]&m[417]&m[418]&~m[445])|(~m[415]&m[416]&m[417]&m[418]&~m[445]))&BiasedRNG[258])|(((m[415]&~m[416]&~m[417]&~m[418]&m[445])|(~m[415]&m[416]&~m[417]&~m[418]&m[445])|(~m[415]&~m[416]&m[417]&~m[418]&m[445])|(m[415]&m[416]&~m[417]&m[418]&m[445])|(m[415]&~m[416]&m[417]&m[418]&m[445])|(~m[415]&m[416]&m[417]&m[418]&m[445]))&~BiasedRNG[258])|((m[415]&m[416]&~m[417]&~m[418]&~m[445])|(m[415]&~m[416]&m[417]&~m[418]&~m[445])|(~m[415]&m[416]&m[417]&~m[418]&~m[445])|(m[415]&m[416]&m[417]&~m[418]&~m[445])|(m[415]&m[416]&m[417]&m[418]&~m[445])|(m[415]&m[416]&~m[417]&~m[418]&m[445])|(m[415]&~m[416]&m[417]&~m[418]&m[445])|(~m[415]&m[416]&m[417]&~m[418]&m[445])|(m[415]&m[416]&m[417]&~m[418]&m[445])|(m[415]&m[416]&m[417]&m[418]&m[445]))):InitCond[476];
    m[424] = run?((((m[420]&~m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&~m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&~m[422]&m[423]&~m[447])|(m[420]&~m[421]&m[422]&m[423]&~m[447])|(~m[420]&m[421]&m[422]&m[423]&~m[447]))&BiasedRNG[259])|(((m[420]&~m[421]&~m[422]&~m[423]&m[447])|(~m[420]&m[421]&~m[422]&~m[423]&m[447])|(~m[420]&~m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&~m[422]&m[423]&m[447])|(m[420]&~m[421]&m[422]&m[423]&m[447])|(~m[420]&m[421]&m[422]&m[423]&m[447]))&~BiasedRNG[259])|((m[420]&m[421]&~m[422]&~m[423]&~m[447])|(m[420]&~m[421]&m[422]&~m[423]&~m[447])|(~m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&m[423]&~m[447])|(m[420]&m[421]&~m[422]&~m[423]&m[447])|(m[420]&~m[421]&m[422]&~m[423]&m[447])|(~m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&m[423]&m[447]))):InitCond[477];
    m[429] = run?((((m[425]&~m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&~m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&~m[427]&m[428]&~m[452])|(m[425]&~m[426]&m[427]&m[428]&~m[452])|(~m[425]&m[426]&m[427]&m[428]&~m[452]))&BiasedRNG[260])|(((m[425]&~m[426]&~m[427]&~m[428]&m[452])|(~m[425]&m[426]&~m[427]&~m[428]&m[452])|(~m[425]&~m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&~m[427]&m[428]&m[452])|(m[425]&~m[426]&m[427]&m[428]&m[452])|(~m[425]&m[426]&m[427]&m[428]&m[452]))&~BiasedRNG[260])|((m[425]&m[426]&~m[427]&~m[428]&~m[452])|(m[425]&~m[426]&m[427]&~m[428]&~m[452])|(~m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&m[428]&~m[452])|(m[425]&m[426]&~m[427]&~m[428]&m[452])|(m[425]&~m[426]&m[427]&~m[428]&m[452])|(~m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&m[428]&m[452]))):InitCond[478];
    m[434] = run?((((m[430]&~m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&~m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&~m[432]&m[433]&~m[457])|(m[430]&~m[431]&m[432]&m[433]&~m[457])|(~m[430]&m[431]&m[432]&m[433]&~m[457]))&BiasedRNG[261])|(((m[430]&~m[431]&~m[432]&~m[433]&m[457])|(~m[430]&m[431]&~m[432]&~m[433]&m[457])|(~m[430]&~m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&~m[432]&m[433]&m[457])|(m[430]&~m[431]&m[432]&m[433]&m[457])|(~m[430]&m[431]&m[432]&m[433]&m[457]))&~BiasedRNG[261])|((m[430]&m[431]&~m[432]&~m[433]&~m[457])|(m[430]&~m[431]&m[432]&~m[433]&~m[457])|(~m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&m[433]&~m[457])|(m[430]&m[431]&~m[432]&~m[433]&m[457])|(m[430]&~m[431]&m[432]&~m[433]&m[457])|(~m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&m[433]&m[457]))):InitCond[479];
    m[439] = run?((((m[435]&~m[436]&~m[437]&~m[438]&~m[462])|(~m[435]&m[436]&~m[437]&~m[438]&~m[462])|(~m[435]&~m[436]&m[437]&~m[438]&~m[462])|(m[435]&m[436]&~m[437]&m[438]&~m[462])|(m[435]&~m[436]&m[437]&m[438]&~m[462])|(~m[435]&m[436]&m[437]&m[438]&~m[462]))&BiasedRNG[262])|(((m[435]&~m[436]&~m[437]&~m[438]&m[462])|(~m[435]&m[436]&~m[437]&~m[438]&m[462])|(~m[435]&~m[436]&m[437]&~m[438]&m[462])|(m[435]&m[436]&~m[437]&m[438]&m[462])|(m[435]&~m[436]&m[437]&m[438]&m[462])|(~m[435]&m[436]&m[437]&m[438]&m[462]))&~BiasedRNG[262])|((m[435]&m[436]&~m[437]&~m[438]&~m[462])|(m[435]&~m[436]&m[437]&~m[438]&~m[462])|(~m[435]&m[436]&m[437]&~m[438]&~m[462])|(m[435]&m[436]&m[437]&~m[438]&~m[462])|(m[435]&m[436]&m[437]&m[438]&~m[462])|(m[435]&m[436]&~m[437]&~m[438]&m[462])|(m[435]&~m[436]&m[437]&~m[438]&m[462])|(~m[435]&m[436]&m[437]&~m[438]&m[462])|(m[435]&m[436]&m[437]&~m[438]&m[462])|(m[435]&m[436]&m[437]&m[438]&m[462]))):InitCond[480];
    m[444] = run?((((m[440]&~m[441]&~m[442]&~m[443]&~m[467])|(~m[440]&m[441]&~m[442]&~m[443]&~m[467])|(~m[440]&~m[441]&m[442]&~m[443]&~m[467])|(m[440]&m[441]&~m[442]&m[443]&~m[467])|(m[440]&~m[441]&m[442]&m[443]&~m[467])|(~m[440]&m[441]&m[442]&m[443]&~m[467]))&BiasedRNG[263])|(((m[440]&~m[441]&~m[442]&~m[443]&m[467])|(~m[440]&m[441]&~m[442]&~m[443]&m[467])|(~m[440]&~m[441]&m[442]&~m[443]&m[467])|(m[440]&m[441]&~m[442]&m[443]&m[467])|(m[440]&~m[441]&m[442]&m[443]&m[467])|(~m[440]&m[441]&m[442]&m[443]&m[467]))&~BiasedRNG[263])|((m[440]&m[441]&~m[442]&~m[443]&~m[467])|(m[440]&~m[441]&m[442]&~m[443]&~m[467])|(~m[440]&m[441]&m[442]&~m[443]&~m[467])|(m[440]&m[441]&m[442]&~m[443]&~m[467])|(m[440]&m[441]&m[442]&m[443]&~m[467])|(m[440]&m[441]&~m[442]&~m[443]&m[467])|(m[440]&~m[441]&m[442]&~m[443]&m[467])|(~m[440]&m[441]&m[442]&~m[443]&m[467])|(m[440]&m[441]&m[442]&~m[443]&m[467])|(m[440]&m[441]&m[442]&m[443]&m[467]))):InitCond[481];
    m[449] = run?((((m[445]&~m[446]&~m[447]&~m[448]&~m[470])|(~m[445]&m[446]&~m[447]&~m[448]&~m[470])|(~m[445]&~m[446]&m[447]&~m[448]&~m[470])|(m[445]&m[446]&~m[447]&m[448]&~m[470])|(m[445]&~m[446]&m[447]&m[448]&~m[470])|(~m[445]&m[446]&m[447]&m[448]&~m[470]))&BiasedRNG[264])|(((m[445]&~m[446]&~m[447]&~m[448]&m[470])|(~m[445]&m[446]&~m[447]&~m[448]&m[470])|(~m[445]&~m[446]&m[447]&~m[448]&m[470])|(m[445]&m[446]&~m[447]&m[448]&m[470])|(m[445]&~m[446]&m[447]&m[448]&m[470])|(~m[445]&m[446]&m[447]&m[448]&m[470]))&~BiasedRNG[264])|((m[445]&m[446]&~m[447]&~m[448]&~m[470])|(m[445]&~m[446]&m[447]&~m[448]&~m[470])|(~m[445]&m[446]&m[447]&~m[448]&~m[470])|(m[445]&m[446]&m[447]&~m[448]&~m[470])|(m[445]&m[446]&m[447]&m[448]&~m[470])|(m[445]&m[446]&~m[447]&~m[448]&m[470])|(m[445]&~m[446]&m[447]&~m[448]&m[470])|(~m[445]&m[446]&m[447]&~m[448]&m[470])|(m[445]&m[446]&m[447]&~m[448]&m[470])|(m[445]&m[446]&m[447]&m[448]&m[470]))):InitCond[482];
    m[454] = run?((((m[450]&~m[451]&~m[452]&~m[453]&~m[472])|(~m[450]&m[451]&~m[452]&~m[453]&~m[472])|(~m[450]&~m[451]&m[452]&~m[453]&~m[472])|(m[450]&m[451]&~m[452]&m[453]&~m[472])|(m[450]&~m[451]&m[452]&m[453]&~m[472])|(~m[450]&m[451]&m[452]&m[453]&~m[472]))&BiasedRNG[265])|(((m[450]&~m[451]&~m[452]&~m[453]&m[472])|(~m[450]&m[451]&~m[452]&~m[453]&m[472])|(~m[450]&~m[451]&m[452]&~m[453]&m[472])|(m[450]&m[451]&~m[452]&m[453]&m[472])|(m[450]&~m[451]&m[452]&m[453]&m[472])|(~m[450]&m[451]&m[452]&m[453]&m[472]))&~BiasedRNG[265])|((m[450]&m[451]&~m[452]&~m[453]&~m[472])|(m[450]&~m[451]&m[452]&~m[453]&~m[472])|(~m[450]&m[451]&m[452]&~m[453]&~m[472])|(m[450]&m[451]&m[452]&~m[453]&~m[472])|(m[450]&m[451]&m[452]&m[453]&~m[472])|(m[450]&m[451]&~m[452]&~m[453]&m[472])|(m[450]&~m[451]&m[452]&~m[453]&m[472])|(~m[450]&m[451]&m[452]&~m[453]&m[472])|(m[450]&m[451]&m[452]&~m[453]&m[472])|(m[450]&m[451]&m[452]&m[453]&m[472]))):InitCond[483];
    m[459] = run?((((m[455]&~m[456]&~m[457]&~m[458]&~m[477])|(~m[455]&m[456]&~m[457]&~m[458]&~m[477])|(~m[455]&~m[456]&m[457]&~m[458]&~m[477])|(m[455]&m[456]&~m[457]&m[458]&~m[477])|(m[455]&~m[456]&m[457]&m[458]&~m[477])|(~m[455]&m[456]&m[457]&m[458]&~m[477]))&BiasedRNG[266])|(((m[455]&~m[456]&~m[457]&~m[458]&m[477])|(~m[455]&m[456]&~m[457]&~m[458]&m[477])|(~m[455]&~m[456]&m[457]&~m[458]&m[477])|(m[455]&m[456]&~m[457]&m[458]&m[477])|(m[455]&~m[456]&m[457]&m[458]&m[477])|(~m[455]&m[456]&m[457]&m[458]&m[477]))&~BiasedRNG[266])|((m[455]&m[456]&~m[457]&~m[458]&~m[477])|(m[455]&~m[456]&m[457]&~m[458]&~m[477])|(~m[455]&m[456]&m[457]&~m[458]&~m[477])|(m[455]&m[456]&m[457]&~m[458]&~m[477])|(m[455]&m[456]&m[457]&m[458]&~m[477])|(m[455]&m[456]&~m[457]&~m[458]&m[477])|(m[455]&~m[456]&m[457]&~m[458]&m[477])|(~m[455]&m[456]&m[457]&~m[458]&m[477])|(m[455]&m[456]&m[457]&~m[458]&m[477])|(m[455]&m[456]&m[457]&m[458]&m[477]))):InitCond[484];
    m[464] = run?((((m[460]&~m[461]&~m[462]&~m[463]&~m[482])|(~m[460]&m[461]&~m[462]&~m[463]&~m[482])|(~m[460]&~m[461]&m[462]&~m[463]&~m[482])|(m[460]&m[461]&~m[462]&m[463]&~m[482])|(m[460]&~m[461]&m[462]&m[463]&~m[482])|(~m[460]&m[461]&m[462]&m[463]&~m[482]))&BiasedRNG[267])|(((m[460]&~m[461]&~m[462]&~m[463]&m[482])|(~m[460]&m[461]&~m[462]&~m[463]&m[482])|(~m[460]&~m[461]&m[462]&~m[463]&m[482])|(m[460]&m[461]&~m[462]&m[463]&m[482])|(m[460]&~m[461]&m[462]&m[463]&m[482])|(~m[460]&m[461]&m[462]&m[463]&m[482]))&~BiasedRNG[267])|((m[460]&m[461]&~m[462]&~m[463]&~m[482])|(m[460]&~m[461]&m[462]&~m[463]&~m[482])|(~m[460]&m[461]&m[462]&~m[463]&~m[482])|(m[460]&m[461]&m[462]&~m[463]&~m[482])|(m[460]&m[461]&m[462]&m[463]&~m[482])|(m[460]&m[461]&~m[462]&~m[463]&m[482])|(m[460]&~m[461]&m[462]&~m[463]&m[482])|(~m[460]&m[461]&m[462]&~m[463]&m[482])|(m[460]&m[461]&m[462]&~m[463]&m[482])|(m[460]&m[461]&m[462]&m[463]&m[482]))):InitCond[485];
    m[469] = run?((((m[465]&~m[466]&~m[467]&~m[468]&~m[487])|(~m[465]&m[466]&~m[467]&~m[468]&~m[487])|(~m[465]&~m[466]&m[467]&~m[468]&~m[487])|(m[465]&m[466]&~m[467]&m[468]&~m[487])|(m[465]&~m[466]&m[467]&m[468]&~m[487])|(~m[465]&m[466]&m[467]&m[468]&~m[487]))&BiasedRNG[268])|(((m[465]&~m[466]&~m[467]&~m[468]&m[487])|(~m[465]&m[466]&~m[467]&~m[468]&m[487])|(~m[465]&~m[466]&m[467]&~m[468]&m[487])|(m[465]&m[466]&~m[467]&m[468]&m[487])|(m[465]&~m[466]&m[467]&m[468]&m[487])|(~m[465]&m[466]&m[467]&m[468]&m[487]))&~BiasedRNG[268])|((m[465]&m[466]&~m[467]&~m[468]&~m[487])|(m[465]&~m[466]&m[467]&~m[468]&~m[487])|(~m[465]&m[466]&m[467]&~m[468]&~m[487])|(m[465]&m[466]&m[467]&~m[468]&~m[487])|(m[465]&m[466]&m[467]&m[468]&~m[487])|(m[465]&m[466]&~m[467]&~m[468]&m[487])|(m[465]&~m[466]&m[467]&~m[468]&m[487])|(~m[465]&m[466]&m[467]&~m[468]&m[487])|(m[465]&m[466]&m[467]&~m[468]&m[487])|(m[465]&m[466]&m[467]&m[468]&m[487]))):InitCond[486];
    m[474] = run?((((m[470]&~m[471]&~m[472]&~m[473]&~m[490])|(~m[470]&m[471]&~m[472]&~m[473]&~m[490])|(~m[470]&~m[471]&m[472]&~m[473]&~m[490])|(m[470]&m[471]&~m[472]&m[473]&~m[490])|(m[470]&~m[471]&m[472]&m[473]&~m[490])|(~m[470]&m[471]&m[472]&m[473]&~m[490]))&BiasedRNG[269])|(((m[470]&~m[471]&~m[472]&~m[473]&m[490])|(~m[470]&m[471]&~m[472]&~m[473]&m[490])|(~m[470]&~m[471]&m[472]&~m[473]&m[490])|(m[470]&m[471]&~m[472]&m[473]&m[490])|(m[470]&~m[471]&m[472]&m[473]&m[490])|(~m[470]&m[471]&m[472]&m[473]&m[490]))&~BiasedRNG[269])|((m[470]&m[471]&~m[472]&~m[473]&~m[490])|(m[470]&~m[471]&m[472]&~m[473]&~m[490])|(~m[470]&m[471]&m[472]&~m[473]&~m[490])|(m[470]&m[471]&m[472]&~m[473]&~m[490])|(m[470]&m[471]&m[472]&m[473]&~m[490])|(m[470]&m[471]&~m[472]&~m[473]&m[490])|(m[470]&~m[471]&m[472]&~m[473]&m[490])|(~m[470]&m[471]&m[472]&~m[473]&m[490])|(m[470]&m[471]&m[472]&~m[473]&m[490])|(m[470]&m[471]&m[472]&m[473]&m[490]))):InitCond[487];
    m[479] = run?((((m[475]&~m[476]&~m[477]&~m[478]&~m[492])|(~m[475]&m[476]&~m[477]&~m[478]&~m[492])|(~m[475]&~m[476]&m[477]&~m[478]&~m[492])|(m[475]&m[476]&~m[477]&m[478]&~m[492])|(m[475]&~m[476]&m[477]&m[478]&~m[492])|(~m[475]&m[476]&m[477]&m[478]&~m[492]))&BiasedRNG[270])|(((m[475]&~m[476]&~m[477]&~m[478]&m[492])|(~m[475]&m[476]&~m[477]&~m[478]&m[492])|(~m[475]&~m[476]&m[477]&~m[478]&m[492])|(m[475]&m[476]&~m[477]&m[478]&m[492])|(m[475]&~m[476]&m[477]&m[478]&m[492])|(~m[475]&m[476]&m[477]&m[478]&m[492]))&~BiasedRNG[270])|((m[475]&m[476]&~m[477]&~m[478]&~m[492])|(m[475]&~m[476]&m[477]&~m[478]&~m[492])|(~m[475]&m[476]&m[477]&~m[478]&~m[492])|(m[475]&m[476]&m[477]&~m[478]&~m[492])|(m[475]&m[476]&m[477]&m[478]&~m[492])|(m[475]&m[476]&~m[477]&~m[478]&m[492])|(m[475]&~m[476]&m[477]&~m[478]&m[492])|(~m[475]&m[476]&m[477]&~m[478]&m[492])|(m[475]&m[476]&m[477]&~m[478]&m[492])|(m[475]&m[476]&m[477]&m[478]&m[492]))):InitCond[488];
    m[484] = run?((((m[480]&~m[481]&~m[482]&~m[483]&~m[497])|(~m[480]&m[481]&~m[482]&~m[483]&~m[497])|(~m[480]&~m[481]&m[482]&~m[483]&~m[497])|(m[480]&m[481]&~m[482]&m[483]&~m[497])|(m[480]&~m[481]&m[482]&m[483]&~m[497])|(~m[480]&m[481]&m[482]&m[483]&~m[497]))&BiasedRNG[271])|(((m[480]&~m[481]&~m[482]&~m[483]&m[497])|(~m[480]&m[481]&~m[482]&~m[483]&m[497])|(~m[480]&~m[481]&m[482]&~m[483]&m[497])|(m[480]&m[481]&~m[482]&m[483]&m[497])|(m[480]&~m[481]&m[482]&m[483]&m[497])|(~m[480]&m[481]&m[482]&m[483]&m[497]))&~BiasedRNG[271])|((m[480]&m[481]&~m[482]&~m[483]&~m[497])|(m[480]&~m[481]&m[482]&~m[483]&~m[497])|(~m[480]&m[481]&m[482]&~m[483]&~m[497])|(m[480]&m[481]&m[482]&~m[483]&~m[497])|(m[480]&m[481]&m[482]&m[483]&~m[497])|(m[480]&m[481]&~m[482]&~m[483]&m[497])|(m[480]&~m[481]&m[482]&~m[483]&m[497])|(~m[480]&m[481]&m[482]&~m[483]&m[497])|(m[480]&m[481]&m[482]&~m[483]&m[497])|(m[480]&m[481]&m[482]&m[483]&m[497]))):InitCond[489];
    m[489] = run?((((m[485]&~m[486]&~m[487]&~m[488]&~m[502])|(~m[485]&m[486]&~m[487]&~m[488]&~m[502])|(~m[485]&~m[486]&m[487]&~m[488]&~m[502])|(m[485]&m[486]&~m[487]&m[488]&~m[502])|(m[485]&~m[486]&m[487]&m[488]&~m[502])|(~m[485]&m[486]&m[487]&m[488]&~m[502]))&BiasedRNG[272])|(((m[485]&~m[486]&~m[487]&~m[488]&m[502])|(~m[485]&m[486]&~m[487]&~m[488]&m[502])|(~m[485]&~m[486]&m[487]&~m[488]&m[502])|(m[485]&m[486]&~m[487]&m[488]&m[502])|(m[485]&~m[486]&m[487]&m[488]&m[502])|(~m[485]&m[486]&m[487]&m[488]&m[502]))&~BiasedRNG[272])|((m[485]&m[486]&~m[487]&~m[488]&~m[502])|(m[485]&~m[486]&m[487]&~m[488]&~m[502])|(~m[485]&m[486]&m[487]&~m[488]&~m[502])|(m[485]&m[486]&m[487]&~m[488]&~m[502])|(m[485]&m[486]&m[487]&m[488]&~m[502])|(m[485]&m[486]&~m[487]&~m[488]&m[502])|(m[485]&~m[486]&m[487]&~m[488]&m[502])|(~m[485]&m[486]&m[487]&~m[488]&m[502])|(m[485]&m[486]&m[487]&~m[488]&m[502])|(m[485]&m[486]&m[487]&m[488]&m[502]))):InitCond[490];
    m[494] = run?((((m[490]&~m[491]&~m[492]&~m[493]&~m[505])|(~m[490]&m[491]&~m[492]&~m[493]&~m[505])|(~m[490]&~m[491]&m[492]&~m[493]&~m[505])|(m[490]&m[491]&~m[492]&m[493]&~m[505])|(m[490]&~m[491]&m[492]&m[493]&~m[505])|(~m[490]&m[491]&m[492]&m[493]&~m[505]))&BiasedRNG[273])|(((m[490]&~m[491]&~m[492]&~m[493]&m[505])|(~m[490]&m[491]&~m[492]&~m[493]&m[505])|(~m[490]&~m[491]&m[492]&~m[493]&m[505])|(m[490]&m[491]&~m[492]&m[493]&m[505])|(m[490]&~m[491]&m[492]&m[493]&m[505])|(~m[490]&m[491]&m[492]&m[493]&m[505]))&~BiasedRNG[273])|((m[490]&m[491]&~m[492]&~m[493]&~m[505])|(m[490]&~m[491]&m[492]&~m[493]&~m[505])|(~m[490]&m[491]&m[492]&~m[493]&~m[505])|(m[490]&m[491]&m[492]&~m[493]&~m[505])|(m[490]&m[491]&m[492]&m[493]&~m[505])|(m[490]&m[491]&~m[492]&~m[493]&m[505])|(m[490]&~m[491]&m[492]&~m[493]&m[505])|(~m[490]&m[491]&m[492]&~m[493]&m[505])|(m[490]&m[491]&m[492]&~m[493]&m[505])|(m[490]&m[491]&m[492]&m[493]&m[505]))):InitCond[491];
    m[499] = run?((((m[495]&~m[496]&~m[497]&~m[498]&~m[507])|(~m[495]&m[496]&~m[497]&~m[498]&~m[507])|(~m[495]&~m[496]&m[497]&~m[498]&~m[507])|(m[495]&m[496]&~m[497]&m[498]&~m[507])|(m[495]&~m[496]&m[497]&m[498]&~m[507])|(~m[495]&m[496]&m[497]&m[498]&~m[507]))&BiasedRNG[274])|(((m[495]&~m[496]&~m[497]&~m[498]&m[507])|(~m[495]&m[496]&~m[497]&~m[498]&m[507])|(~m[495]&~m[496]&m[497]&~m[498]&m[507])|(m[495]&m[496]&~m[497]&m[498]&m[507])|(m[495]&~m[496]&m[497]&m[498]&m[507])|(~m[495]&m[496]&m[497]&m[498]&m[507]))&~BiasedRNG[274])|((m[495]&m[496]&~m[497]&~m[498]&~m[507])|(m[495]&~m[496]&m[497]&~m[498]&~m[507])|(~m[495]&m[496]&m[497]&~m[498]&~m[507])|(m[495]&m[496]&m[497]&~m[498]&~m[507])|(m[495]&m[496]&m[497]&m[498]&~m[507])|(m[495]&m[496]&~m[497]&~m[498]&m[507])|(m[495]&~m[496]&m[497]&~m[498]&m[507])|(~m[495]&m[496]&m[497]&~m[498]&m[507])|(m[495]&m[496]&m[497]&~m[498]&m[507])|(m[495]&m[496]&m[497]&m[498]&m[507]))):InitCond[492];
    m[504] = run?((((m[500]&~m[501]&~m[502]&~m[503]&~m[512])|(~m[500]&m[501]&~m[502]&~m[503]&~m[512])|(~m[500]&~m[501]&m[502]&~m[503]&~m[512])|(m[500]&m[501]&~m[502]&m[503]&~m[512])|(m[500]&~m[501]&m[502]&m[503]&~m[512])|(~m[500]&m[501]&m[502]&m[503]&~m[512]))&BiasedRNG[275])|(((m[500]&~m[501]&~m[502]&~m[503]&m[512])|(~m[500]&m[501]&~m[502]&~m[503]&m[512])|(~m[500]&~m[501]&m[502]&~m[503]&m[512])|(m[500]&m[501]&~m[502]&m[503]&m[512])|(m[500]&~m[501]&m[502]&m[503]&m[512])|(~m[500]&m[501]&m[502]&m[503]&m[512]))&~BiasedRNG[275])|((m[500]&m[501]&~m[502]&~m[503]&~m[512])|(m[500]&~m[501]&m[502]&~m[503]&~m[512])|(~m[500]&m[501]&m[502]&~m[503]&~m[512])|(m[500]&m[501]&m[502]&~m[503]&~m[512])|(m[500]&m[501]&m[502]&m[503]&~m[512])|(m[500]&m[501]&~m[502]&~m[503]&m[512])|(m[500]&~m[501]&m[502]&~m[503]&m[512])|(~m[500]&m[501]&m[502]&~m[503]&m[512])|(m[500]&m[501]&m[502]&~m[503]&m[512])|(m[500]&m[501]&m[502]&m[503]&m[512]))):InitCond[493];
    m[509] = run?((((m[505]&~m[506]&~m[507]&~m[508]&~m[515])|(~m[505]&m[506]&~m[507]&~m[508]&~m[515])|(~m[505]&~m[506]&m[507]&~m[508]&~m[515])|(m[505]&m[506]&~m[507]&m[508]&~m[515])|(m[505]&~m[506]&m[507]&m[508]&~m[515])|(~m[505]&m[506]&m[507]&m[508]&~m[515]))&BiasedRNG[276])|(((m[505]&~m[506]&~m[507]&~m[508]&m[515])|(~m[505]&m[506]&~m[507]&~m[508]&m[515])|(~m[505]&~m[506]&m[507]&~m[508]&m[515])|(m[505]&m[506]&~m[507]&m[508]&m[515])|(m[505]&~m[506]&m[507]&m[508]&m[515])|(~m[505]&m[506]&m[507]&m[508]&m[515]))&~BiasedRNG[276])|((m[505]&m[506]&~m[507]&~m[508]&~m[515])|(m[505]&~m[506]&m[507]&~m[508]&~m[515])|(~m[505]&m[506]&m[507]&~m[508]&~m[515])|(m[505]&m[506]&m[507]&~m[508]&~m[515])|(m[505]&m[506]&m[507]&m[508]&~m[515])|(m[505]&m[506]&~m[507]&~m[508]&m[515])|(m[505]&~m[506]&m[507]&~m[508]&m[515])|(~m[505]&m[506]&m[507]&~m[508]&m[515])|(m[505]&m[506]&m[507]&~m[508]&m[515])|(m[505]&m[506]&m[507]&m[508]&m[515]))):InitCond[494];
    m[514] = run?((((m[510]&~m[511]&~m[512]&~m[513]&~m[517])|(~m[510]&m[511]&~m[512]&~m[513]&~m[517])|(~m[510]&~m[511]&m[512]&~m[513]&~m[517])|(m[510]&m[511]&~m[512]&m[513]&~m[517])|(m[510]&~m[511]&m[512]&m[513]&~m[517])|(~m[510]&m[511]&m[512]&m[513]&~m[517]))&BiasedRNG[277])|(((m[510]&~m[511]&~m[512]&~m[513]&m[517])|(~m[510]&m[511]&~m[512]&~m[513]&m[517])|(~m[510]&~m[511]&m[512]&~m[513]&m[517])|(m[510]&m[511]&~m[512]&m[513]&m[517])|(m[510]&~m[511]&m[512]&m[513]&m[517])|(~m[510]&m[511]&m[512]&m[513]&m[517]))&~BiasedRNG[277])|((m[510]&m[511]&~m[512]&~m[513]&~m[517])|(m[510]&~m[511]&m[512]&~m[513]&~m[517])|(~m[510]&m[511]&m[512]&~m[513]&~m[517])|(m[510]&m[511]&m[512]&~m[513]&~m[517])|(m[510]&m[511]&m[512]&m[513]&~m[517])|(m[510]&m[511]&~m[512]&~m[513]&m[517])|(m[510]&~m[511]&m[512]&~m[513]&m[517])|(~m[510]&m[511]&m[512]&~m[513]&m[517])|(m[510]&m[511]&m[512]&~m[513]&m[517])|(m[510]&m[511]&m[512]&m[513]&m[517]))):InitCond[495];
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[119]&LFSRcolor0[178]&LFSRcolor0[106]);
    BiasedRNG[1] = (LFSRcolor0[109]&LFSRcolor0[1]&LFSRcolor0[30]);
    BiasedRNG[2] = (LFSRcolor0[180]&LFSRcolor0[195]&LFSRcolor0[37]);
    BiasedRNG[3] = (LFSRcolor0[51]&LFSRcolor0[104]&LFSRcolor0[161]);
    BiasedRNG[4] = (LFSRcolor0[90]&LFSRcolor0[230]&LFSRcolor0[78]);
    BiasedRNG[5] = (LFSRcolor0[247]&LFSRcolor0[203]&LFSRcolor0[163]);
    BiasedRNG[6] = (LFSRcolor0[250]&LFSRcolor0[245]&LFSRcolor0[14]);
    BiasedRNG[7] = (LFSRcolor0[112]&LFSRcolor0[207]&LFSRcolor0[91]);
    BiasedRNG[8] = (LFSRcolor0[93]&LFSRcolor0[130]&LFSRcolor0[113]);
    BiasedRNG[9] = (LFSRcolor0[52]&LFSRcolor0[162]&LFSRcolor0[26]);
    BiasedRNG[10] = (LFSRcolor0[6]&LFSRcolor0[141]&LFSRcolor0[271]);
    BiasedRNG[11] = (LFSRcolor0[80]&LFSRcolor0[160]&LFSRcolor0[40]);
    BiasedRNG[12] = (LFSRcolor0[204]&LFSRcolor0[274]&LFSRcolor0[33]);
    BiasedRNG[13] = (LFSRcolor0[116]&LFSRcolor0[63]&LFSRcolor0[138]);
    BiasedRNG[14] = (LFSRcolor0[122]&LFSRcolor0[202]&LFSRcolor0[210]);
    BiasedRNG[15] = (LFSRcolor0[21]&LFSRcolor0[273]&LFSRcolor0[168]);
    BiasedRNG[16] = (LFSRcolor0[265]&LFSRcolor0[25]&LFSRcolor0[58]);
    BiasedRNG[17] = (LFSRcolor0[166]&LFSRcolor0[244]&LFSRcolor0[86]);
    BiasedRNG[18] = (LFSRcolor0[155]&LFSRcolor0[13]&LFSRcolor0[68]);
    BiasedRNG[19] = (LFSRcolor0[3]&LFSRcolor0[154]&LFSRcolor0[17]);
    BiasedRNG[20] = (LFSRcolor0[231]&LFSRcolor0[65]&LFSRcolor0[146]);
    BiasedRNG[21] = (LFSRcolor0[239]&LFSRcolor0[186]&LFSRcolor0[38]);
    BiasedRNG[22] = (LFSRcolor0[228]&LFSRcolor0[107]&LFSRcolor0[173]);
    BiasedRNG[23] = (LFSRcolor0[187]&LFSRcolor0[272]&LFSRcolor0[246]);
    BiasedRNG[24] = (LFSRcolor0[142]&LFSRcolor0[35]&LFSRcolor0[124]);
    BiasedRNG[25] = (LFSRcolor0[54]&LFSRcolor0[24]&LFSRcolor0[42]);
    BiasedRNG[26] = (LFSRcolor0[192]&LFSRcolor0[46]&LFSRcolor0[132]);
    BiasedRNG[27] = (LFSRcolor0[100]&LFSRcolor0[164]&LFSRcolor0[2]);
    BiasedRNG[28] = (LFSRcolor0[200]&LFSRcolor0[172]&LFSRcolor0[151]);
    BiasedRNG[29] = (LFSRcolor0[19]&LFSRcolor0[12]&LFSRcolor0[236]);
    BiasedRNG[30] = (LFSRcolor0[97]&LFSRcolor0[227]&LFSRcolor0[177]);
    BiasedRNG[31] = (LFSRcolor0[152]&LFSRcolor0[243]&LFSRcolor0[148]);
    BiasedRNG[32] = (LFSRcolor0[118]&LFSRcolor0[34]&LFSRcolor0[85]);
    BiasedRNG[33] = (LFSRcolor0[89]&LFSRcolor0[240]&LFSRcolor0[275]);
    BiasedRNG[34] = (LFSRcolor0[208]&LFSRcolor0[147]&LFSRcolor0[221]);
    BiasedRNG[35] = (LFSRcolor0[223]&LFSRcolor0[175]&LFSRcolor0[182]);
    BiasedRNG[36] = (LFSRcolor0[238]&LFSRcolor0[31]&LFSRcolor0[153]);
    BiasedRNG[37] = (LFSRcolor0[127]&LFSRcolor0[50]&LFSRcolor0[55]);
    BiasedRNG[38] = (LFSRcolor0[115]&LFSRcolor0[196]&LFSRcolor0[249]);
    BiasedRNG[39] = (LFSRcolor0[129]&LFSRcolor0[57]&LFSRcolor0[62]);
    BiasedRNG[40] = (LFSRcolor0[61]&LFSRcolor0[184]&LFSRcolor0[242]);
    BiasedRNG[41] = (LFSRcolor0[111]&LFSRcolor0[235]&LFSRcolor0[20]);
    BiasedRNG[42] = (LFSRcolor0[74]&LFSRcolor0[181]&LFSRcolor0[103]);
    BiasedRNG[43] = (LFSRcolor0[0]&LFSRcolor0[258]&LFSRcolor0[16]);
    BiasedRNG[44] = (LFSRcolor0[27]&LFSRcolor0[135]&LFSRcolor0[139]);
    BiasedRNG[45] = (LFSRcolor0[7]&LFSRcolor0[22]&LFSRcolor0[237]);
    BiasedRNG[46] = (LFSRcolor0[169]&LFSRcolor0[9]&LFSRcolor0[70]);
    BiasedRNG[47] = (LFSRcolor0[264]&LFSRcolor0[18]&LFSRcolor0[226]);
    BiasedRNG[48] = (LFSRcolor0[99]&LFSRcolor0[45]&LFSRcolor0[188]);
    BiasedRNG[49] = (LFSRcolor0[56]&LFSRcolor0[83]&LFSRcolor0[137]);
    BiasedRNG[50] = (LFSRcolor0[266]&LFSRcolor0[205]&LFSRcolor0[157]);
    BiasedRNG[51] = (LFSRcolor0[149]&LFSRcolor0[233]&LFSRcolor0[225]);
    BiasedRNG[52] = (LFSRcolor0[253]&LFSRcolor0[255]&LFSRcolor0[36]);
    BiasedRNG[53] = (LFSRcolor0[79]&LFSRcolor0[201]&LFSRcolor0[260]);
    BiasedRNG[54] = (LFSRcolor0[120]&LFSRcolor0[5]&LFSRcolor0[82]);
    BiasedRNG[55] = (LFSRcolor0[262]&LFSRcolor0[252]&LFSRcolor0[257]);
    BiasedRNG[56] = (LFSRcolor0[259]&LFSRcolor0[32]&LFSRcolor0[193]);
    BiasedRNG[57] = (LFSRcolor0[81]&LFSRcolor0[217]&LFSRcolor0[110]);
    BiasedRNG[58] = (LFSRcolor0[156]&LFSRcolor0[165]&LFSRcolor0[261]);
    BiasedRNG[59] = (LFSRcolor0[263]&LFSRcolor0[96]&LFSRcolor0[114]);
    BiasedRNG[60] = (LFSRcolor0[197]&LFSRcolor0[256]&LFSRcolor0[8]);
    BiasedRNG[61] = (LFSRcolor0[123]&LFSRcolor0[213]&LFSRcolor0[84]);
    BiasedRNG[62] = (LFSRcolor0[176]&LFSRcolor0[140]&LFSRcolor0[194]);
    BiasedRNG[63] = (LFSRcolor0[214]&LFSRcolor0[28]&LFSRcolor0[71]);
    UnbiasedRNG[0] = LFSRcolor0[224];
    UnbiasedRNG[1] = LFSRcolor0[49];
    UnbiasedRNG[2] = LFSRcolor0[128];
    UnbiasedRNG[3] = LFSRcolor0[234];
    UnbiasedRNG[4] = LFSRcolor0[43];
    UnbiasedRNG[5] = LFSRcolor0[183];
    UnbiasedRNG[6] = LFSRcolor0[126];
    UnbiasedRNG[7] = LFSRcolor0[53];
    UnbiasedRNG[8] = LFSRcolor0[198];
    UnbiasedRNG[9] = LFSRcolor0[254];
    UnbiasedRNG[10] = LFSRcolor0[241];
    UnbiasedRNG[11] = LFSRcolor0[145];
    UnbiasedRNG[12] = LFSRcolor0[11];
    UnbiasedRNG[13] = LFSRcolor0[219];
    UnbiasedRNG[14] = LFSRcolor0[76];
    UnbiasedRNG[15] = LFSRcolor0[15];
    UnbiasedRNG[16] = LFSRcolor0[94];
    UnbiasedRNG[17] = LFSRcolor0[267];
    UnbiasedRNG[18] = LFSRcolor0[144];
    UnbiasedRNG[19] = LFSRcolor0[150];
    UnbiasedRNG[20] = LFSRcolor0[77];
    UnbiasedRNG[21] = LFSRcolor0[143];
    UnbiasedRNG[22] = LFSRcolor0[41];
    UnbiasedRNG[23] = LFSRcolor0[44];
    UnbiasedRNG[24] = LFSRcolor0[48];
    UnbiasedRNG[25] = LFSRcolor0[174];
    UnbiasedRNG[26] = LFSRcolor0[220];
    UnbiasedRNG[27] = LFSRcolor0[212];
    UnbiasedRNG[28] = LFSRcolor0[159];
    UnbiasedRNG[29] = LFSRcolor0[218];
    UnbiasedRNG[30] = LFSRcolor0[248];
    UnbiasedRNG[31] = LFSRcolor0[158];
    UnbiasedRNG[32] = LFSRcolor0[270];
    UnbiasedRNG[33] = LFSRcolor0[215];
    UnbiasedRNG[34] = LFSRcolor0[136];
    UnbiasedRNG[35] = LFSRcolor0[108];
    UnbiasedRNG[36] = LFSRcolor0[268];
    UnbiasedRNG[37] = LFSRcolor0[269];
    UnbiasedRNG[38] = LFSRcolor0[47];
    UnbiasedRNG[39] = LFSRcolor0[92];
    UnbiasedRNG[40] = LFSRcolor0[102];
    UnbiasedRNG[41] = LFSRcolor0[134];
    UnbiasedRNG[42] = LFSRcolor0[88];
    UnbiasedRNG[43] = LFSRcolor0[105];
    UnbiasedRNG[44] = LFSRcolor0[170];
    UnbiasedRNG[45] = LFSRcolor0[206];
    UnbiasedRNG[46] = LFSRcolor0[4];
    UnbiasedRNG[47] = LFSRcolor0[73];
    UnbiasedRNG[48] = LFSRcolor0[251];
    UnbiasedRNG[49] = LFSRcolor0[167];
    UnbiasedRNG[50] = LFSRcolor0[98];
    UnbiasedRNG[51] = LFSRcolor0[29];
    UnbiasedRNG[52] = LFSRcolor0[59];
    UnbiasedRNG[53] = LFSRcolor0[95];
    UnbiasedRNG[54] = LFSRcolor0[209];
    UnbiasedRNG[55] = LFSRcolor0[101];
    UnbiasedRNG[56] = LFSRcolor0[232];
    UnbiasedRNG[57] = LFSRcolor0[171];
    UnbiasedRNG[58] = LFSRcolor0[87];
    UnbiasedRNG[59] = LFSRcolor0[23];
    UnbiasedRNG[60] = LFSRcolor0[39];
    UnbiasedRNG[61] = LFSRcolor0[69];
    UnbiasedRNG[62] = LFSRcolor0[64];
    UnbiasedRNG[63] = LFSRcolor0[211];
    UnbiasedRNG[64] = LFSRcolor0[117];
    UnbiasedRNG[65] = LFSRcolor0[189];
    UnbiasedRNG[66] = LFSRcolor0[191];
    UnbiasedRNG[67] = LFSRcolor0[75];
    UnbiasedRNG[68] = LFSRcolor0[67];
    UnbiasedRNG[69] = LFSRcolor0[190];
    UnbiasedRNG[70] = LFSRcolor0[10];
end

always @(posedge color0_clk) begin
    BiasedRNG[64] = (LFSRcolor1[39]&LFSRcolor1[278]&LFSRcolor1[234]);
    BiasedRNG[65] = (LFSRcolor1[165]&LFSRcolor1[320]&LFSRcolor1[152]);
    BiasedRNG[66] = (LFSRcolor1[177]&LFSRcolor1[357]&LFSRcolor1[199]);
    BiasedRNG[67] = (LFSRcolor1[365]&LFSRcolor1[46]&LFSRcolor1[269]);
    BiasedRNG[68] = (LFSRcolor1[105]&LFSRcolor1[142]&LFSRcolor1[158]);
    BiasedRNG[69] = (LFSRcolor1[140]&LFSRcolor1[224]&LFSRcolor1[248]);
    BiasedRNG[70] = (LFSRcolor1[354]&LFSRcolor1[8]&LFSRcolor1[208]);
    BiasedRNG[71] = (LFSRcolor1[350]&LFSRcolor1[3]&LFSRcolor1[103]);
    BiasedRNG[72] = (LFSRcolor1[4]&LFSRcolor1[173]&LFSRcolor1[207]);
    BiasedRNG[73] = (LFSRcolor1[77]&LFSRcolor1[115]&LFSRcolor1[108]);
    BiasedRNG[74] = (LFSRcolor1[112]&LFSRcolor1[306]&LFSRcolor1[213]);
    BiasedRNG[75] = (LFSRcolor1[221]&LFSRcolor1[290]&LFSRcolor1[124]);
    BiasedRNG[76] = (LFSRcolor1[82]&LFSRcolor1[136]&LFSRcolor1[264]);
    BiasedRNG[77] = (LFSRcolor1[318]&LFSRcolor1[49]&LFSRcolor1[229]);
    BiasedRNG[78] = (LFSRcolor1[344]&LFSRcolor1[190]&LFSRcolor1[361]);
    BiasedRNG[79] = (LFSRcolor1[338]&LFSRcolor1[170]&LFSRcolor1[56]);
    BiasedRNG[80] = (LFSRcolor1[200]&LFSRcolor1[174]&LFSRcolor1[113]);
    BiasedRNG[81] = (LFSRcolor1[125]&LFSRcolor1[265]&LFSRcolor1[257]);
    BiasedRNG[82] = (LFSRcolor1[315]&LFSRcolor1[276]&LFSRcolor1[28]);
    BiasedRNG[83] = (LFSRcolor1[88]&LFSRcolor1[246]&LFSRcolor1[24]);
    BiasedRNG[84] = (LFSRcolor1[206]&LFSRcolor1[7]&LFSRcolor1[272]);
    BiasedRNG[85] = (LFSRcolor1[6]&LFSRcolor1[138]&LFSRcolor1[171]);
    BiasedRNG[86] = (LFSRcolor1[220]&LFSRcolor1[331]&LFSRcolor1[346]);
    BiasedRNG[87] = (LFSRcolor1[232]&LFSRcolor1[79]&LFSRcolor1[282]);
    BiasedRNG[88] = (LFSRcolor1[226]&LFSRcolor1[319]&LFSRcolor1[321]);
    BiasedRNG[89] = (LFSRcolor1[367]&LFSRcolor1[355]&LFSRcolor1[145]);
    BiasedRNG[90] = (LFSRcolor1[218]&LFSRcolor1[85]&LFSRcolor1[19]);
    BiasedRNG[91] = (LFSRcolor1[227]&LFSRcolor1[96]&LFSRcolor1[216]);
    BiasedRNG[92] = (LFSRcolor1[256]&LFSRcolor1[341]&LFSRcolor1[308]);
    BiasedRNG[93] = (LFSRcolor1[0]&LFSRcolor1[188]&LFSRcolor1[111]);
    BiasedRNG[94] = (LFSRcolor1[57]&LFSRcolor1[363]&LFSRcolor1[83]);
    BiasedRNG[95] = (LFSRcolor1[304]&LFSRcolor1[243]&LFSRcolor1[134]);
    BiasedRNG[96] = (LFSRcolor1[347]&LFSRcolor1[149]&LFSRcolor1[100]);
    BiasedRNG[97] = (LFSRcolor1[65]&LFSRcolor1[179]&LFSRcolor1[117]);
    BiasedRNG[98] = (LFSRcolor1[62]&LFSRcolor1[102]&LFSRcolor1[84]);
    BiasedRNG[99] = (LFSRcolor1[31]&LFSRcolor1[230]&LFSRcolor1[285]);
    BiasedRNG[100] = (LFSRcolor1[130]&LFSRcolor1[160]&LFSRcolor1[120]);
    BiasedRNG[101] = (LFSRcolor1[237]&LFSRcolor1[40]&LFSRcolor1[240]);
    BiasedRNG[102] = (LFSRcolor1[186]&LFSRcolor1[143]&LFSRcolor1[348]);
    BiasedRNG[103] = (LFSRcolor1[274]&LFSRcolor1[121]&LFSRcolor1[250]);
    BiasedRNG[104] = (LFSRcolor1[157]&LFSRcolor1[148]&LFSRcolor1[135]);
    BiasedRNG[105] = (LFSRcolor1[326]&LFSRcolor1[61]&LFSRcolor1[172]);
    BiasedRNG[106] = (LFSRcolor1[13]&LFSRcolor1[233]&LFSRcolor1[328]);
    BiasedRNG[107] = (LFSRcolor1[50]&LFSRcolor1[260]&LFSRcolor1[296]);
    BiasedRNG[108] = (LFSRcolor1[182]&LFSRcolor1[301]&LFSRcolor1[305]);
    BiasedRNG[109] = (LFSRcolor1[110]&LFSRcolor1[330]&LFSRcolor1[317]);
    BiasedRNG[110] = (LFSRcolor1[2]&LFSRcolor1[231]&LFSRcolor1[68]);
    BiasedRNG[111] = (LFSRcolor1[21]&LFSRcolor1[212]&LFSRcolor1[52]);
    BiasedRNG[112] = (LFSRcolor1[129]&LFSRcolor1[273]&LFSRcolor1[128]);
    BiasedRNG[113] = (LFSRcolor1[154]&LFSRcolor1[176]&LFSRcolor1[195]);
    BiasedRNG[114] = (LFSRcolor1[55]&LFSRcolor1[191]&LFSRcolor1[340]);
    BiasedRNG[115] = (LFSRcolor1[261]&LFSRcolor1[307]&LFSRcolor1[223]);
    BiasedRNG[116] = (LFSRcolor1[364]&LFSRcolor1[187]&LFSRcolor1[298]);
    BiasedRNG[117] = (LFSRcolor1[332]&LFSRcolor1[300]&LFSRcolor1[91]);
    BiasedRNG[118] = (LFSRcolor1[87]&LFSRcolor1[137]&LFSRcolor1[72]);
    BiasedRNG[119] = (LFSRcolor1[169]&LFSRcolor1[325]&LFSRcolor1[342]);
    BiasedRNG[120] = (LFSRcolor1[59]&LFSRcolor1[180]&LFSRcolor1[185]);
    BiasedRNG[121] = (LFSRcolor1[313]&LFSRcolor1[147]&LFSRcolor1[241]);
    BiasedRNG[122] = (LFSRcolor1[41]&LFSRcolor1[255]&LFSRcolor1[242]);
    BiasedRNG[123] = (LFSRcolor1[294]&LFSRcolor1[245]&LFSRcolor1[345]);
    BiasedRNG[124] = (LFSRcolor1[38]&LFSRcolor1[193]&LFSRcolor1[153]);
    BiasedRNG[125] = (LFSRcolor1[201]&LFSRcolor1[132]&LFSRcolor1[109]);
    BiasedRNG[126] = (LFSRcolor1[262]&LFSRcolor1[175]&LFSRcolor1[196]);
    BiasedRNG[127] = (LFSRcolor1[67]&LFSRcolor1[360]&LFSRcolor1[316]);
    BiasedRNG[128] = (LFSRcolor1[51]&LFSRcolor1[215]&LFSRcolor1[17]);
    BiasedRNG[129] = (LFSRcolor1[219]&LFSRcolor1[310]&LFSRcolor1[80]);
    BiasedRNG[130] = (LFSRcolor1[277]&LFSRcolor1[334]&LFSRcolor1[42]);
    BiasedRNG[131] = (LFSRcolor1[312]&LFSRcolor1[178]&LFSRcolor1[209]);
    BiasedRNG[132] = (LFSRcolor1[205]&LFSRcolor1[214]&LFSRcolor1[311]);
    BiasedRNG[133] = (LFSRcolor1[225]&LFSRcolor1[69]&LFSRcolor1[283]);
    BiasedRNG[134] = (LFSRcolor1[329]&LFSRcolor1[18]&LFSRcolor1[295]);
    BiasedRNG[135] = (LFSRcolor1[97]&LFSRcolor1[15]&LFSRcolor1[25]);
    BiasedRNG[136] = (LFSRcolor1[239]&LFSRcolor1[279]&LFSRcolor1[63]);
    BiasedRNG[137] = (LFSRcolor1[75]&LFSRcolor1[189]&LFSRcolor1[90]);
    BiasedRNG[138] = (LFSRcolor1[14]&LFSRcolor1[150]&LFSRcolor1[47]);
    BiasedRNG[139] = (LFSRcolor1[235]&LFSRcolor1[34]&LFSRcolor1[339]);
    BiasedRNG[140] = (LFSRcolor1[45]&LFSRcolor1[118]&LFSRcolor1[131]);
    BiasedRNG[141] = (LFSRcolor1[16]&LFSRcolor1[322]&LFSRcolor1[197]);
    BiasedRNG[142] = (LFSRcolor1[291]&LFSRcolor1[366]&LFSRcolor1[26]);
    BiasedRNG[143] = (LFSRcolor1[106]&LFSRcolor1[114]&LFSRcolor1[133]);
    BiasedRNG[144] = (LFSRcolor1[222]&LFSRcolor1[211]&LFSRcolor1[181]);
    BiasedRNG[145] = (LFSRcolor1[252]&LFSRcolor1[95]&LFSRcolor1[254]);
    BiasedRNG[146] = (LFSRcolor1[98]&LFSRcolor1[309]&LFSRcolor1[119]);
    BiasedRNG[147] = (LFSRcolor1[48]&LFSRcolor1[352]&LFSRcolor1[297]);
    BiasedRNG[148] = (LFSRcolor1[362]&LFSRcolor1[253]&LFSRcolor1[53]);
    BiasedRNG[149] = (LFSRcolor1[64]&LFSRcolor1[198]&LFSRcolor1[122]);
    BiasedRNG[150] = (LFSRcolor1[336]&LFSRcolor1[284]&LFSRcolor1[166]);
    BiasedRNG[151] = (LFSRcolor1[73]&LFSRcolor1[280]&LFSRcolor1[139]);
    BiasedRNG[152] = (LFSRcolor1[271]&LFSRcolor1[20]&LFSRcolor1[356]);
    BiasedRNG[153] = (LFSRcolor1[151]&LFSRcolor1[30]&LFSRcolor1[293]);
    BiasedRNG[154] = (LFSRcolor1[1]&LFSRcolor1[156]&LFSRcolor1[289]);
    BiasedRNG[155] = (LFSRcolor1[244]&LFSRcolor1[33]&LFSRcolor1[35]);
    BiasedRNG[156] = (LFSRcolor1[70]&LFSRcolor1[324]&LFSRcolor1[5]);
    BiasedRNG[157] = (LFSRcolor1[164]&LFSRcolor1[36]&LFSRcolor1[314]);
    BiasedRNG[158] = (LFSRcolor1[351]&LFSRcolor1[268]&LFSRcolor1[92]);
    UnbiasedRNG[71] = LFSRcolor1[204];
    UnbiasedRNG[72] = LFSRcolor1[9];
    UnbiasedRNG[73] = LFSRcolor1[359];
    UnbiasedRNG[74] = LFSRcolor1[168];
    UnbiasedRNG[75] = LFSRcolor1[94];
    UnbiasedRNG[76] = LFSRcolor1[286];
    UnbiasedRNG[77] = LFSRcolor1[81];
    UnbiasedRNG[78] = LFSRcolor1[11];
    UnbiasedRNG[79] = LFSRcolor1[162];
    UnbiasedRNG[80] = LFSRcolor1[270];
    UnbiasedRNG[81] = LFSRcolor1[275];
    UnbiasedRNG[82] = LFSRcolor1[247];
    UnbiasedRNG[83] = LFSRcolor1[66];
    UnbiasedRNG[84] = LFSRcolor1[266];
    UnbiasedRNG[85] = LFSRcolor1[251];
    UnbiasedRNG[86] = LFSRcolor1[184];
    UnbiasedRNG[87] = LFSRcolor1[22];
    UnbiasedRNG[88] = LFSRcolor1[238];
    UnbiasedRNG[89] = LFSRcolor1[101];
    UnbiasedRNG[90] = LFSRcolor1[203];
    UnbiasedRNG[91] = LFSRcolor1[99];
    UnbiasedRNG[92] = LFSRcolor1[144];
    UnbiasedRNG[93] = LFSRcolor1[89];
    UnbiasedRNG[94] = LFSRcolor1[74];
    UnbiasedRNG[95] = LFSRcolor1[86];
    UnbiasedRNG[96] = LFSRcolor1[281];
    UnbiasedRNG[97] = LFSRcolor1[163];
    UnbiasedRNG[98] = LFSRcolor1[202];
    UnbiasedRNG[99] = LFSRcolor1[107];
    UnbiasedRNG[100] = LFSRcolor1[335];
    UnbiasedRNG[101] = LFSRcolor1[349];
    UnbiasedRNG[102] = LFSRcolor1[27];
    UnbiasedRNG[103] = LFSRcolor1[259];
    UnbiasedRNG[104] = LFSRcolor1[217];
    UnbiasedRNG[105] = LFSRcolor1[161];
    UnbiasedRNG[106] = LFSRcolor1[126];
    UnbiasedRNG[107] = LFSRcolor1[127];
    UnbiasedRNG[108] = LFSRcolor1[343];
    UnbiasedRNG[109] = LFSRcolor1[29];
    UnbiasedRNG[110] = LFSRcolor1[333];
    UnbiasedRNG[111] = LFSRcolor1[288];
    UnbiasedRNG[112] = LFSRcolor1[194];
    UnbiasedRNG[113] = LFSRcolor1[302];
    UnbiasedRNG[114] = LFSRcolor1[353];
    UnbiasedRNG[115] = LFSRcolor1[60];
    UnbiasedRNG[116] = LFSRcolor1[299];
    UnbiasedRNG[117] = LFSRcolor1[358];
    UnbiasedRNG[118] = LFSRcolor1[71];
    UnbiasedRNG[119] = LFSRcolor1[159];
end

always @(posedge color1_clk) begin
    BiasedRNG[159] = (LFSRcolor2[253]&LFSRcolor2[274]&LFSRcolor2[122]);
    BiasedRNG[160] = (LFSRcolor2[125]&LFSRcolor2[88]&LFSRcolor2[162]);
    BiasedRNG[161] = (LFSRcolor2[44]&LFSRcolor2[18]&LFSRcolor2[25]);
    BiasedRNG[162] = (LFSRcolor2[260]&LFSRcolor2[42]&LFSRcolor2[198]);
    BiasedRNG[163] = (LFSRcolor2[192]&LFSRcolor2[57]&LFSRcolor2[74]);
    BiasedRNG[164] = (LFSRcolor2[19]&LFSRcolor2[188]&LFSRcolor2[115]);
    BiasedRNG[165] = (LFSRcolor2[136]&LFSRcolor2[254]&LFSRcolor2[222]);
    BiasedRNG[166] = (LFSRcolor2[189]&LFSRcolor2[244]&LFSRcolor2[261]);
    BiasedRNG[167] = (LFSRcolor2[8]&LFSRcolor2[36]&LFSRcolor2[69]);
    BiasedRNG[168] = (LFSRcolor2[13]&LFSRcolor2[181]&LFSRcolor2[6]);
    BiasedRNG[169] = (LFSRcolor2[120]&LFSRcolor2[82]&LFSRcolor2[175]);
    BiasedRNG[170] = (LFSRcolor2[135]&LFSRcolor2[217]&LFSRcolor2[235]);
    BiasedRNG[171] = (LFSRcolor2[216]&LFSRcolor2[171]&LFSRcolor2[102]);
    BiasedRNG[172] = (LFSRcolor2[223]&LFSRcolor2[178]&LFSRcolor2[111]);
    BiasedRNG[173] = (LFSRcolor2[60]&LFSRcolor2[163]&LFSRcolor2[56]);
    BiasedRNG[174] = (LFSRcolor2[170]&LFSRcolor2[154]&LFSRcolor2[240]);
    BiasedRNG[175] = (LFSRcolor2[194]&LFSRcolor2[186]&LFSRcolor2[262]);
    BiasedRNG[176] = (LFSRcolor2[20]&LFSRcolor2[161]&LFSRcolor2[75]);
    BiasedRNG[177] = (LFSRcolor2[251]&LFSRcolor2[221]&LFSRcolor2[73]);
    BiasedRNG[178] = (LFSRcolor2[242]&LFSRcolor2[53]&LFSRcolor2[127]);
    BiasedRNG[179] = (LFSRcolor2[47]&LFSRcolor2[77]&LFSRcolor2[9]);
    BiasedRNG[180] = (LFSRcolor2[7]&LFSRcolor2[72]&LFSRcolor2[264]);
    BiasedRNG[181] = (LFSRcolor2[27]&LFSRcolor2[220]&LFSRcolor2[90]);
    BiasedRNG[182] = (LFSRcolor2[193]&LFSRcolor2[100]&LFSRcolor2[237]);
    BiasedRNG[183] = (LFSRcolor2[184]&LFSRcolor2[201]&LFSRcolor2[55]);
    BiasedRNG[184] = (LFSRcolor2[11]&LFSRcolor2[58]&LFSRcolor2[156]);
    BiasedRNG[185] = (LFSRcolor2[24]&LFSRcolor2[227]&LFSRcolor2[252]);
    BiasedRNG[186] = (LFSRcolor2[139]&LFSRcolor2[267]&LFSRcolor2[144]);
    BiasedRNG[187] = (LFSRcolor2[43]&LFSRcolor2[26]&LFSRcolor2[99]);
    BiasedRNG[188] = (LFSRcolor2[199]&LFSRcolor2[208]&LFSRcolor2[39]);
    BiasedRNG[189] = (LFSRcolor2[79]&LFSRcolor2[12]&LFSRcolor2[113]);
    BiasedRNG[190] = (LFSRcolor2[233]&LFSRcolor2[76]&LFSRcolor2[232]);
    BiasedRNG[191] = (LFSRcolor2[93]&LFSRcolor2[91]&LFSRcolor2[143]);
    BiasedRNG[192] = (LFSRcolor2[95]&LFSRcolor2[152]&LFSRcolor2[225]);
    BiasedRNG[193] = (LFSRcolor2[64]&LFSRcolor2[197]&LFSRcolor2[157]);
    BiasedRNG[194] = (LFSRcolor2[272]&LFSRcolor2[185]&LFSRcolor2[146]);
    BiasedRNG[195] = (LFSRcolor2[23]&LFSRcolor2[248]&LFSRcolor2[176]);
    BiasedRNG[196] = (LFSRcolor2[268]&LFSRcolor2[204]&LFSRcolor2[2]);
    BiasedRNG[197] = (LFSRcolor2[159]&LFSRcolor2[65]&LFSRcolor2[228]);
    BiasedRNG[198] = (LFSRcolor2[249]&LFSRcolor2[123]&LFSRcolor2[104]);
    BiasedRNG[199] = (LFSRcolor2[59]&LFSRcolor2[211]&LFSRcolor2[70]);
    BiasedRNG[200] = (LFSRcolor2[50]&LFSRcolor2[187]&LFSRcolor2[141]);
    BiasedRNG[201] = (LFSRcolor2[195]&LFSRcolor2[66]&LFSRcolor2[138]);
    BiasedRNG[202] = (LFSRcolor2[112]&LFSRcolor2[116]&LFSRcolor2[29]);
    BiasedRNG[203] = (LFSRcolor2[119]&LFSRcolor2[172]&LFSRcolor2[3]);
    BiasedRNG[204] = (LFSRcolor2[103]&LFSRcolor2[212]&LFSRcolor2[63]);
    BiasedRNG[205] = (LFSRcolor2[31]&LFSRcolor2[33]&LFSRcolor2[173]);
    BiasedRNG[206] = (LFSRcolor2[255]&LFSRcolor2[140]&LFSRcolor2[164]);
    BiasedRNG[207] = (LFSRcolor2[202]&LFSRcolor2[54]&LFSRcolor2[247]);
    BiasedRNG[208] = (LFSRcolor2[166]&LFSRcolor2[270]&LFSRcolor2[207]);
    BiasedRNG[209] = (LFSRcolor2[49]&LFSRcolor2[200]&LFSRcolor2[41]);
    BiasedRNG[210] = (LFSRcolor2[14]&LFSRcolor2[86]&LFSRcolor2[196]);
    BiasedRNG[211] = (LFSRcolor2[149]&LFSRcolor2[229]&LFSRcolor2[275]);
    BiasedRNG[212] = (LFSRcolor2[230]&LFSRcolor2[250]&LFSRcolor2[238]);
    BiasedRNG[213] = (LFSRcolor2[61]&LFSRcolor2[94]&LFSRcolor2[206]);
    BiasedRNG[214] = (LFSRcolor2[219]&LFSRcolor2[213]&LFSRcolor2[84]);
    BiasedRNG[215] = (LFSRcolor2[105]&LFSRcolor2[110]&LFSRcolor2[98]);
    BiasedRNG[216] = (LFSRcolor2[205]&LFSRcolor2[259]&LFSRcolor2[231]);
    BiasedRNG[217] = (LFSRcolor2[269]&LFSRcolor2[224]&LFSRcolor2[180]);
    BiasedRNG[218] = (LFSRcolor2[226]&LFSRcolor2[130]&LFSRcolor2[131]);
    BiasedRNG[219] = (LFSRcolor2[133]&LFSRcolor2[215]&LFSRcolor2[256]);
    BiasedRNG[220] = (LFSRcolor2[108]&LFSRcolor2[28]&LFSRcolor2[10]);
    BiasedRNG[221] = (LFSRcolor2[168]&LFSRcolor2[101]&LFSRcolor2[147]);
    BiasedRNG[222] = (LFSRcolor2[241]&LFSRcolor2[78]&LFSRcolor2[32]);
    UnbiasedRNG[120] = LFSRcolor2[97];
    UnbiasedRNG[121] = LFSRcolor2[85];
    UnbiasedRNG[122] = LFSRcolor2[191];
    UnbiasedRNG[123] = LFSRcolor2[174];
    UnbiasedRNG[124] = LFSRcolor2[210];
    UnbiasedRNG[125] = LFSRcolor2[179];
    UnbiasedRNG[126] = LFSRcolor2[37];
    UnbiasedRNG[127] = LFSRcolor2[266];
    UnbiasedRNG[128] = LFSRcolor2[118];
    UnbiasedRNG[129] = LFSRcolor2[81];
    UnbiasedRNG[130] = LFSRcolor2[234];
    UnbiasedRNG[131] = LFSRcolor2[243];
    UnbiasedRNG[132] = LFSRcolor2[126];
    UnbiasedRNG[133] = LFSRcolor2[153];
    UnbiasedRNG[134] = LFSRcolor2[158];
    UnbiasedRNG[135] = LFSRcolor2[35];
    UnbiasedRNG[136] = LFSRcolor2[21];
    UnbiasedRNG[137] = LFSRcolor2[0];
    UnbiasedRNG[138] = LFSRcolor2[257];
    UnbiasedRNG[139] = LFSRcolor2[46];
    UnbiasedRNG[140] = LFSRcolor2[22];
    UnbiasedRNG[141] = LFSRcolor2[263];
    UnbiasedRNG[142] = LFSRcolor2[71];
    UnbiasedRNG[143] = LFSRcolor2[17];
    UnbiasedRNG[144] = LFSRcolor2[15];
    UnbiasedRNG[145] = LFSRcolor2[190];
    UnbiasedRNG[146] = LFSRcolor2[40];
    UnbiasedRNG[147] = LFSRcolor2[148];
    UnbiasedRNG[148] = LFSRcolor2[214];
    UnbiasedRNG[149] = LFSRcolor2[87];
    UnbiasedRNG[150] = LFSRcolor2[236];
    UnbiasedRNG[151] = LFSRcolor2[160];
    UnbiasedRNG[152] = LFSRcolor2[177];
    UnbiasedRNG[153] = LFSRcolor2[265];
    UnbiasedRNG[154] = LFSRcolor2[4];
    UnbiasedRNG[155] = LFSRcolor2[151];
    UnbiasedRNG[156] = LFSRcolor2[182];
    UnbiasedRNG[157] = LFSRcolor2[129];
    UnbiasedRNG[158] = LFSRcolor2[271];
    UnbiasedRNG[159] = LFSRcolor2[1];
    UnbiasedRNG[160] = LFSRcolor2[80];
    UnbiasedRNG[161] = LFSRcolor2[106];
    UnbiasedRNG[162] = LFSRcolor2[165];
    UnbiasedRNG[163] = LFSRcolor2[169];
    UnbiasedRNG[164] = LFSRcolor2[246];
    UnbiasedRNG[165] = LFSRcolor2[5];
    UnbiasedRNG[166] = LFSRcolor2[38];
    UnbiasedRNG[167] = LFSRcolor2[155];
    UnbiasedRNG[168] = LFSRcolor2[16];
    UnbiasedRNG[169] = LFSRcolor2[30];
    UnbiasedRNG[170] = LFSRcolor2[132];
    UnbiasedRNG[171] = LFSRcolor2[45];
    UnbiasedRNG[172] = LFSRcolor2[51];
    UnbiasedRNG[173] = LFSRcolor2[209];
    UnbiasedRNG[174] = LFSRcolor2[150];
    UnbiasedRNG[175] = LFSRcolor2[117];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[176] = LFSRcolor3[18];
    UnbiasedRNG[177] = LFSRcolor3[17];
    UnbiasedRNG[178] = LFSRcolor3[29];
    UnbiasedRNG[179] = LFSRcolor3[11];
    UnbiasedRNG[180] = LFSRcolor3[28];
    UnbiasedRNG[181] = LFSRcolor3[8];
    UnbiasedRNG[182] = LFSRcolor3[2];
    UnbiasedRNG[183] = LFSRcolor3[37];
    UnbiasedRNG[184] = LFSRcolor3[24];
    UnbiasedRNG[185] = LFSRcolor3[45];
    UnbiasedRNG[186] = LFSRcolor3[41];
    UnbiasedRNG[187] = LFSRcolor3[40];
    UnbiasedRNG[188] = LFSRcolor3[5];
    UnbiasedRNG[189] = LFSRcolor3[33];
    UnbiasedRNG[190] = LFSRcolor3[12];
    UnbiasedRNG[191] = LFSRcolor3[9];
    UnbiasedRNG[192] = LFSRcolor3[31];
    UnbiasedRNG[193] = LFSRcolor3[32];
    UnbiasedRNG[194] = LFSRcolor3[20];
    UnbiasedRNG[195] = LFSRcolor3[4];
    UnbiasedRNG[196] = LFSRcolor3[3];
    UnbiasedRNG[197] = LFSRcolor3[25];
    UnbiasedRNG[198] = LFSRcolor3[10];
    UnbiasedRNG[199] = LFSRcolor3[36];
    UnbiasedRNG[200] = LFSRcolor3[30];
    UnbiasedRNG[201] = LFSRcolor3[13];
    UnbiasedRNG[202] = LFSRcolor3[42];
    UnbiasedRNG[203] = LFSRcolor3[0];
    UnbiasedRNG[204] = LFSRcolor3[44];
    UnbiasedRNG[205] = LFSRcolor3[15];
    UnbiasedRNG[206] = LFSRcolor3[19];
    UnbiasedRNG[207] = LFSRcolor3[23];
    UnbiasedRNG[208] = LFSRcolor3[38];
    UnbiasedRNG[209] = LFSRcolor3[26];
    UnbiasedRNG[210] = LFSRcolor3[22];
    UnbiasedRNG[211] = LFSRcolor3[7];
    UnbiasedRNG[212] = LFSRcolor3[27];
    UnbiasedRNG[213] = LFSRcolor3[14];
    UnbiasedRNG[214] = LFSRcolor3[43];
    UnbiasedRNG[215] = LFSRcolor3[6];
    UnbiasedRNG[216] = LFSRcolor3[34];
    UnbiasedRNG[217] = LFSRcolor3[1];
end

always @(posedge color3_clk) begin
    BiasedRNG[223] = (LFSRcolor4[95]&LFSRcolor4[64]&LFSRcolor4[42]);
    BiasedRNG[224] = (LFSRcolor4[174]&LFSRcolor4[76]&LFSRcolor4[74]);
    BiasedRNG[225] = (LFSRcolor4[137]&LFSRcolor4[150]&LFSRcolor4[126]);
    BiasedRNG[226] = (LFSRcolor4[18]&LFSRcolor4[121]&LFSRcolor4[163]);
    BiasedRNG[227] = (LFSRcolor4[130]&LFSRcolor4[52]&LFSRcolor4[106]);
    BiasedRNG[228] = (LFSRcolor4[99]&LFSRcolor4[164]&LFSRcolor4[138]);
    BiasedRNG[229] = (LFSRcolor4[120]&LFSRcolor4[78]&LFSRcolor4[123]);
    BiasedRNG[230] = (LFSRcolor4[41]&LFSRcolor4[131]&LFSRcolor4[118]);
    BiasedRNG[231] = (LFSRcolor4[160]&LFSRcolor4[90]&LFSRcolor4[92]);
    BiasedRNG[232] = (LFSRcolor4[58]&LFSRcolor4[14]&LFSRcolor4[69]);
    BiasedRNG[233] = (LFSRcolor4[107]&LFSRcolor4[141]&LFSRcolor4[45]);
    BiasedRNG[234] = (LFSRcolor4[5]&LFSRcolor4[105]&LFSRcolor4[122]);
    BiasedRNG[235] = (LFSRcolor4[182]&LFSRcolor4[66]&LFSRcolor4[140]);
    BiasedRNG[236] = (LFSRcolor4[148]&LFSRcolor4[23]&LFSRcolor4[104]);
    BiasedRNG[237] = (LFSRcolor4[59]&LFSRcolor4[75]&LFSRcolor4[67]);
    BiasedRNG[238] = (LFSRcolor4[111]&LFSRcolor4[70]&LFSRcolor4[110]);
    BiasedRNG[239] = (LFSRcolor4[93]&LFSRcolor4[54]&LFSRcolor4[39]);
    BiasedRNG[240] = (LFSRcolor4[83]&LFSRcolor4[65]&LFSRcolor4[145]);
    BiasedRNG[241] = (LFSRcolor4[60]&LFSRcolor4[171]&LFSRcolor4[117]);
    BiasedRNG[242] = (LFSRcolor4[27]&LFSRcolor4[155]&LFSRcolor4[119]);
    BiasedRNG[243] = (LFSRcolor4[85]&LFSRcolor4[4]&LFSRcolor4[89]);
    BiasedRNG[244] = (LFSRcolor4[116]&LFSRcolor4[77]&LFSRcolor4[178]);
    BiasedRNG[245] = (LFSRcolor4[167]&LFSRcolor4[48]&LFSRcolor4[32]);
    BiasedRNG[246] = (LFSRcolor4[35]&LFSRcolor4[136]&LFSRcolor4[112]);
    BiasedRNG[247] = (LFSRcolor4[56]&LFSRcolor4[91]&LFSRcolor4[26]);
    BiasedRNG[248] = (LFSRcolor4[180]&LFSRcolor4[169]&LFSRcolor4[47]);
    BiasedRNG[249] = (LFSRcolor4[152]&LFSRcolor4[132]&LFSRcolor4[24]);
    BiasedRNG[250] = (LFSRcolor4[20]&LFSRcolor4[33]&LFSRcolor4[168]);
    BiasedRNG[251] = (LFSRcolor4[175]&LFSRcolor4[149]&LFSRcolor4[133]);
    BiasedRNG[252] = (LFSRcolor4[147]&LFSRcolor4[57]&LFSRcolor4[177]);
    BiasedRNG[253] = (LFSRcolor4[96]&LFSRcolor4[21]&LFSRcolor4[100]);
    BiasedRNG[254] = (LFSRcolor4[159]&LFSRcolor4[43]&LFSRcolor4[25]);
    BiasedRNG[255] = (LFSRcolor4[179]&LFSRcolor4[73]&LFSRcolor4[165]);
    BiasedRNG[256] = (LFSRcolor4[1]&LFSRcolor4[103]&LFSRcolor4[7]);
    BiasedRNG[257] = (LFSRcolor4[8]&LFSRcolor4[71]&LFSRcolor4[55]);
    BiasedRNG[258] = (LFSRcolor4[9]&LFSRcolor4[88]&LFSRcolor4[146]);
    BiasedRNG[259] = (LFSRcolor4[81]&LFSRcolor4[97]&LFSRcolor4[16]);
    BiasedRNG[260] = (LFSRcolor4[30]&LFSRcolor4[166]&LFSRcolor4[17]);
    BiasedRNG[261] = (LFSRcolor4[101]&LFSRcolor4[157]&LFSRcolor4[128]);
    BiasedRNG[262] = (LFSRcolor4[143]&LFSRcolor4[6]&LFSRcolor4[13]);
    BiasedRNG[263] = (LFSRcolor4[156]&LFSRcolor4[79]&LFSRcolor4[109]);
    BiasedRNG[264] = (LFSRcolor4[115]&LFSRcolor4[153]&LFSRcolor4[15]);
    BiasedRNG[265] = (LFSRcolor4[84]&LFSRcolor4[108]&LFSRcolor4[10]);
    BiasedRNG[266] = (LFSRcolor4[68]&LFSRcolor4[154]&LFSRcolor4[144]);
    BiasedRNG[267] = (LFSRcolor4[37]&LFSRcolor4[63]&LFSRcolor4[46]);
    BiasedRNG[268] = (LFSRcolor4[53]&LFSRcolor4[142]&LFSRcolor4[113]);
    BiasedRNG[269] = (LFSRcolor4[0]&LFSRcolor4[61]&LFSRcolor4[176]);
    BiasedRNG[270] = (LFSRcolor4[183]&LFSRcolor4[2]&LFSRcolor4[129]);
    BiasedRNG[271] = (LFSRcolor4[127]&LFSRcolor4[12]&LFSRcolor4[31]);
    BiasedRNG[272] = (LFSRcolor4[181]&LFSRcolor4[28]&LFSRcolor4[114]);
    BiasedRNG[273] = (LFSRcolor4[158]&LFSRcolor4[139]&LFSRcolor4[80]);
    BiasedRNG[274] = (LFSRcolor4[38]&LFSRcolor4[172]&LFSRcolor4[3]);
    BiasedRNG[275] = (LFSRcolor4[86]&LFSRcolor4[50]&LFSRcolor4[161]);
    BiasedRNG[276] = (LFSRcolor4[135]&LFSRcolor4[29]&LFSRcolor4[173]);
    BiasedRNG[277] = (LFSRcolor4[151]&LFSRcolor4[19]&LFSRcolor4[62]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

//Generate the ILA for data collection:
ila_0 ILAinst(.clk(sample_clk),.probe0(run),.probe1(solution_flag),.probe2(failure),.probe3(counter[37:0]));

//Instantiate VIO:
vio_0 VIOinst (.clk(sample_clk),.probe_out0(reset),.probe_out1(solution_set[15:0]));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule