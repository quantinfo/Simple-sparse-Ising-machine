//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [37:0] counter;
initial counter = 38'b0;
reg [11:0] solution;
reg [11:0] solution_check;
wire [11:0] solution_set;
initial solution_check = 12'b110010100001;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
reg [0:263] InitCond;
reg run;
wire [183:0] LFSRcolor0;
wire [183:0] LFSRcolor1;
wire [137:0] LFSRcolor2;
wire [45:0] LFSRcolor3;
wire [91:0] LFSRcolor4;
reg [159:0] BiasedRNG;       //For I=+/-1 cases
reg [103:0] UnbiasedRNG;   //For I=0 cases
reg [0:281] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[96] = 1'b1;
initial m[135] = 1'b0;
initial m[145] = 1'b0;
initial m[160] = 1'b0;
initial m[180] = 1'b0;
initial m[205] = 1'b1;
initial m[230] = 1'b0;
initial m[250] = 1'b1;
initial m[265] = 1'b0;
initial m[275] = 1'b0;
initial m[280] = 1'b1;
initial m[281] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[134] = 1'b0;
initial m[144] = 1'b0;
initial m[159] = 1'b0;
initial m[179] = 1'b0;
initial m[204] = 1'b0;
initial m[207] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
//To control whether the system runs or resets using VIO and counter:
always @(posedge sample_clk) begin
    if (reset) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 12'b0;
        failure = 1'b0;
        solution_check = solution_set;
        m[96] = solution_set[0];
        m[135] = solution_set[1];
        m[145] = solution_set[2];
        m[160] = solution_set[3];
        m[180] = solution_set[4];
        m[205] = solution_set[5];
        m[230] = solution_set[6];
        m[250] = solution_set[7];
        m[265] = solution_set[8];
        m[275] = solution_set[9];
        m[280] = solution_set[10];
        m[281] = solution_set[11];
    end else if (solution_flag) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 12'b0;
        failure = 1'b0;
    end else if (counter < 38'b11111111111111111111111111111111111111) begin
        if (counter == 1) begin
            InitCond[0] = UnbiasedRNG[0];
            InitCond[1] = UnbiasedRNG[1];
            InitCond[2] = UnbiasedRNG[2];
            InitCond[3] = UnbiasedRNG[3];
            InitCond[4] = UnbiasedRNG[4];
            InitCond[5] = UnbiasedRNG[5];
            InitCond[6] = UnbiasedRNG[6];
            InitCond[7] = UnbiasedRNG[7];
            InitCond[8] = UnbiasedRNG[8];
            InitCond[9] = UnbiasedRNG[9];
            InitCond[10] = UnbiasedRNG[10];
            InitCond[11] = UnbiasedRNG[11];
            InitCond[12] = UnbiasedRNG[12];
            InitCond[13] = UnbiasedRNG[13];
            InitCond[14] = UnbiasedRNG[14];
            InitCond[15] = UnbiasedRNG[15];
            InitCond[16] = UnbiasedRNG[16];
            InitCond[17] = UnbiasedRNG[17];
            InitCond[18] = UnbiasedRNG[18];
            InitCond[19] = UnbiasedRNG[19];
            InitCond[20] = UnbiasedRNG[20];
            InitCond[21] = UnbiasedRNG[21];
            InitCond[22] = UnbiasedRNG[22];
            InitCond[23] = UnbiasedRNG[23];
            InitCond[24] = UnbiasedRNG[24];
            InitCond[25] = UnbiasedRNG[25];
            InitCond[26] = UnbiasedRNG[26];
            InitCond[27] = UnbiasedRNG[27];
            InitCond[28] = UnbiasedRNG[28];
            InitCond[29] = UnbiasedRNG[29];
            InitCond[30] = UnbiasedRNG[30];
            InitCond[31] = UnbiasedRNG[31];
            InitCond[32] = UnbiasedRNG[32];
            InitCond[33] = UnbiasedRNG[33];
            InitCond[34] = UnbiasedRNG[34];
            InitCond[35] = UnbiasedRNG[35];
            InitCond[36] = UnbiasedRNG[36];
            InitCond[37] = UnbiasedRNG[37];
            InitCond[38] = UnbiasedRNG[38];
            InitCond[39] = UnbiasedRNG[39];
            InitCond[40] = UnbiasedRNG[40];
            InitCond[41] = UnbiasedRNG[41];
            InitCond[42] = UnbiasedRNG[42];
            InitCond[43] = UnbiasedRNG[43];
            InitCond[44] = UnbiasedRNG[44];
            InitCond[45] = UnbiasedRNG[45];
            InitCond[46] = UnbiasedRNG[46];
            InitCond[47] = UnbiasedRNG[47];
            InitCond[48] = UnbiasedRNG[48];
            InitCond[49] = UnbiasedRNG[49];
            InitCond[50] = UnbiasedRNG[50];
            InitCond[51] = UnbiasedRNG[51];
            InitCond[52] = UnbiasedRNG[52];
            InitCond[53] = UnbiasedRNG[53];
            InitCond[54] = UnbiasedRNG[54];
            InitCond[55] = UnbiasedRNG[55];
            InitCond[56] = UnbiasedRNG[56];
            InitCond[57] = UnbiasedRNG[57];
            InitCond[58] = UnbiasedRNG[58];
            InitCond[59] = UnbiasedRNG[59];
            InitCond[60] = UnbiasedRNG[60];
            InitCond[61] = UnbiasedRNG[61];
            InitCond[62] = UnbiasedRNG[62];
            InitCond[63] = UnbiasedRNG[63];
            InitCond[64] = UnbiasedRNG[64];
            InitCond[65] = UnbiasedRNG[65];
            InitCond[66] = UnbiasedRNG[66];
            InitCond[67] = UnbiasedRNG[67];
            InitCond[68] = UnbiasedRNG[68];
            InitCond[69] = UnbiasedRNG[69];
            InitCond[70] = UnbiasedRNG[70];
            InitCond[71] = UnbiasedRNG[71];
            InitCond[72] = UnbiasedRNG[72];
            InitCond[73] = UnbiasedRNG[73];
            InitCond[74] = UnbiasedRNG[74];
            InitCond[75] = UnbiasedRNG[75];
            InitCond[76] = UnbiasedRNG[76];
            InitCond[77] = UnbiasedRNG[77];
            InitCond[78] = UnbiasedRNG[78];
            InitCond[79] = UnbiasedRNG[79];
            InitCond[80] = UnbiasedRNG[80];
            InitCond[81] = UnbiasedRNG[81];
            InitCond[82] = UnbiasedRNG[82];
            InitCond[83] = UnbiasedRNG[83];
            InitCond[84] = UnbiasedRNG[84];
            InitCond[85] = UnbiasedRNG[85];
            InitCond[86] = UnbiasedRNG[86];
            InitCond[87] = UnbiasedRNG[87];
            InitCond[88] = UnbiasedRNG[88];
            InitCond[89] = UnbiasedRNG[89];
            InitCond[90] = UnbiasedRNG[90];
            InitCond[91] = UnbiasedRNG[91];
            InitCond[92] = UnbiasedRNG[92];
            InitCond[93] = UnbiasedRNG[93];
            InitCond[94] = UnbiasedRNG[94];
            InitCond[95] = UnbiasedRNG[95];
            InitCond[96] = UnbiasedRNG[96];
            InitCond[97] = UnbiasedRNG[97];
            InitCond[98] = UnbiasedRNG[98];
            InitCond[99] = UnbiasedRNG[99];
            InitCond[100] = UnbiasedRNG[100];
            InitCond[101] = UnbiasedRNG[101];
            InitCond[102] = UnbiasedRNG[102];
            InitCond[103] = UnbiasedRNG[103];
        end
        else if (counter == 2) begin
            InitCond[104] = UnbiasedRNG[0];
            InitCond[105] = UnbiasedRNG[1];
            InitCond[106] = UnbiasedRNG[2];
            InitCond[107] = UnbiasedRNG[3];
            InitCond[108] = UnbiasedRNG[4];
            InitCond[109] = UnbiasedRNG[5];
            InitCond[110] = UnbiasedRNG[6];
            InitCond[111] = UnbiasedRNG[7];
            InitCond[112] = UnbiasedRNG[8];
            InitCond[113] = UnbiasedRNG[9];
            InitCond[114] = UnbiasedRNG[10];
            InitCond[115] = UnbiasedRNG[11];
            InitCond[116] = UnbiasedRNG[12];
            InitCond[117] = UnbiasedRNG[13];
            InitCond[118] = UnbiasedRNG[14];
            InitCond[119] = UnbiasedRNG[15];
            InitCond[120] = UnbiasedRNG[16];
            InitCond[121] = UnbiasedRNG[17];
            InitCond[122] = UnbiasedRNG[18];
            InitCond[123] = UnbiasedRNG[19];
            InitCond[124] = UnbiasedRNG[20];
            InitCond[125] = UnbiasedRNG[21];
            InitCond[126] = UnbiasedRNG[22];
            InitCond[127] = UnbiasedRNG[23];
            InitCond[128] = UnbiasedRNG[24];
            InitCond[129] = UnbiasedRNG[25];
            InitCond[130] = UnbiasedRNG[26];
            InitCond[131] = UnbiasedRNG[27];
            InitCond[132] = UnbiasedRNG[28];
            InitCond[133] = UnbiasedRNG[29];
            InitCond[134] = UnbiasedRNG[30];
            InitCond[135] = UnbiasedRNG[31];
            InitCond[136] = UnbiasedRNG[32];
            InitCond[137] = UnbiasedRNG[33];
            InitCond[138] = UnbiasedRNG[34];
            InitCond[139] = UnbiasedRNG[35];
            InitCond[140] = UnbiasedRNG[36];
            InitCond[141] = UnbiasedRNG[37];
            InitCond[142] = UnbiasedRNG[38];
            InitCond[143] = UnbiasedRNG[39];
            InitCond[144] = UnbiasedRNG[40];
            InitCond[145] = UnbiasedRNG[41];
            InitCond[146] = UnbiasedRNG[42];
            InitCond[147] = UnbiasedRNG[43];
            InitCond[148] = UnbiasedRNG[44];
            InitCond[149] = UnbiasedRNG[45];
            InitCond[150] = UnbiasedRNG[46];
            InitCond[151] = UnbiasedRNG[47];
            InitCond[152] = UnbiasedRNG[48];
            InitCond[153] = UnbiasedRNG[49];
            InitCond[154] = UnbiasedRNG[50];
            InitCond[155] = UnbiasedRNG[51];
            InitCond[156] = UnbiasedRNG[52];
            InitCond[157] = UnbiasedRNG[53];
            InitCond[158] = UnbiasedRNG[54];
            InitCond[159] = UnbiasedRNG[55];
            InitCond[160] = UnbiasedRNG[56];
            InitCond[161] = UnbiasedRNG[57];
            InitCond[162] = UnbiasedRNG[58];
            InitCond[163] = UnbiasedRNG[59];
            InitCond[164] = UnbiasedRNG[60];
            InitCond[165] = UnbiasedRNG[61];
            InitCond[166] = UnbiasedRNG[62];
            InitCond[167] = UnbiasedRNG[63];
            InitCond[168] = UnbiasedRNG[64];
            InitCond[169] = UnbiasedRNG[65];
            InitCond[170] = UnbiasedRNG[66];
            InitCond[171] = UnbiasedRNG[67];
            InitCond[172] = UnbiasedRNG[68];
            InitCond[173] = UnbiasedRNG[69];
            InitCond[174] = UnbiasedRNG[70];
            InitCond[175] = UnbiasedRNG[71];
            InitCond[176] = UnbiasedRNG[72];
            InitCond[177] = UnbiasedRNG[73];
            InitCond[178] = UnbiasedRNG[74];
            InitCond[179] = UnbiasedRNG[75];
            InitCond[180] = UnbiasedRNG[76];
            InitCond[181] = UnbiasedRNG[77];
            InitCond[182] = UnbiasedRNG[78];
            InitCond[183] = UnbiasedRNG[79];
            InitCond[184] = UnbiasedRNG[80];
            InitCond[185] = UnbiasedRNG[81];
            InitCond[186] = UnbiasedRNG[82];
            InitCond[187] = UnbiasedRNG[83];
            InitCond[188] = UnbiasedRNG[84];
            InitCond[189] = UnbiasedRNG[85];
            InitCond[190] = UnbiasedRNG[86];
            InitCond[191] = UnbiasedRNG[87];
            InitCond[192] = UnbiasedRNG[88];
            InitCond[193] = UnbiasedRNG[89];
            InitCond[194] = UnbiasedRNG[90];
            InitCond[195] = UnbiasedRNG[91];
            InitCond[196] = UnbiasedRNG[92];
            InitCond[197] = UnbiasedRNG[93];
            InitCond[198] = UnbiasedRNG[94];
            InitCond[199] = UnbiasedRNG[95];
            InitCond[200] = UnbiasedRNG[96];
            InitCond[201] = UnbiasedRNG[97];
            InitCond[202] = UnbiasedRNG[98];
            InitCond[203] = UnbiasedRNG[99];
            InitCond[204] = UnbiasedRNG[100];
            InitCond[205] = UnbiasedRNG[101];
            InitCond[206] = UnbiasedRNG[102];
            InitCond[207] = UnbiasedRNG[103];
        end
        else if (counter == 3) begin
            InitCond[208] = UnbiasedRNG[0];
            InitCond[209] = UnbiasedRNG[1];
            InitCond[210] = UnbiasedRNG[2];
            InitCond[211] = UnbiasedRNG[3];
            InitCond[212] = UnbiasedRNG[4];
            InitCond[213] = UnbiasedRNG[5];
            InitCond[214] = UnbiasedRNG[6];
            InitCond[215] = UnbiasedRNG[7];
            InitCond[216] = UnbiasedRNG[8];
            InitCond[217] = UnbiasedRNG[9];
            InitCond[218] = UnbiasedRNG[10];
            InitCond[219] = UnbiasedRNG[11];
            InitCond[220] = UnbiasedRNG[12];
            InitCond[221] = UnbiasedRNG[13];
            InitCond[222] = UnbiasedRNG[14];
            InitCond[223] = UnbiasedRNG[15];
            InitCond[224] = UnbiasedRNG[16];
            InitCond[225] = UnbiasedRNG[17];
            InitCond[226] = UnbiasedRNG[18];
            InitCond[227] = UnbiasedRNG[19];
            InitCond[228] = UnbiasedRNG[20];
            InitCond[229] = UnbiasedRNG[21];
            InitCond[230] = UnbiasedRNG[22];
            InitCond[231] = UnbiasedRNG[23];
            InitCond[232] = UnbiasedRNG[24];
            InitCond[233] = UnbiasedRNG[25];
            InitCond[234] = UnbiasedRNG[26];
            InitCond[235] = UnbiasedRNG[27];
            InitCond[236] = UnbiasedRNG[28];
            InitCond[237] = UnbiasedRNG[29];
            InitCond[238] = UnbiasedRNG[30];
            InitCond[239] = UnbiasedRNG[31];
            InitCond[240] = UnbiasedRNG[32];
            InitCond[241] = UnbiasedRNG[33];
            InitCond[242] = UnbiasedRNG[34];
            InitCond[243] = UnbiasedRNG[35];
            InitCond[244] = UnbiasedRNG[36];
            InitCond[245] = UnbiasedRNG[37];
            InitCond[246] = UnbiasedRNG[38];
            InitCond[247] = UnbiasedRNG[39];
            InitCond[248] = UnbiasedRNG[40];
            InitCond[249] = UnbiasedRNG[41];
            InitCond[250] = UnbiasedRNG[42];
            InitCond[251] = UnbiasedRNG[43];
            InitCond[252] = UnbiasedRNG[44];
            InitCond[253] = UnbiasedRNG[45];
            InitCond[254] = UnbiasedRNG[46];
            InitCond[255] = UnbiasedRNG[47];
            InitCond[256] = UnbiasedRNG[48];
            InitCond[257] = UnbiasedRNG[49];
            InitCond[258] = UnbiasedRNG[50];
            InitCond[259] = UnbiasedRNG[51];
            InitCond[260] = UnbiasedRNG[52];
            InitCond[261] = UnbiasedRNG[53];
            InitCond[262] = UnbiasedRNG[54];
            InitCond[263] = UnbiasedRNG[55];
        end
        else if (counter==5)
            run = 1'b1;
        counter = counter+38'b1;
        solution = {m[5],m[4],m[3],m[2],m[1],m[0]}*{m[11],m[10],m[9],m[8],m[7],m[6]};
    end else begin 
        counter = 38'b0;
        failure = 1'b1;
        run = 1'b0;
    end
end

//To measure on only the last step using ILA:
always @(negedge sample_clk) begin
    if (solution_flag)
        solution_flag = 1'b0;
    else if ((run & (solution == solution_check)) | failure)
        solution_flag = 1'b1;
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = run?((((m[12]&~m[24]&~m[25])|(~m[12]&m[24]&~m[25])|(~m[12]&~m[24]&m[25]))&BiasedRNG[0])|(((m[12]&m[24]&~m[25])|(m[12]&~m[24]&m[25])|(~m[12]&m[24]&m[25]))&~BiasedRNG[0])|((m[12]&m[24]&m[25]))):InitCond[0];
    m[1] = run?((((m[13]&~m[30]&~m[31])|(~m[13]&m[30]&~m[31])|(~m[13]&~m[30]&m[31]))&BiasedRNG[1])|(((m[13]&m[30]&~m[31])|(m[13]&~m[30]&m[31])|(~m[13]&m[30]&m[31]))&~BiasedRNG[1])|((m[13]&m[30]&m[31]))):InitCond[1];
    m[2] = run?((((m[14]&~m[36]&~m[37])|(~m[14]&m[36]&~m[37])|(~m[14]&~m[36]&m[37]))&BiasedRNG[2])|(((m[14]&m[36]&~m[37])|(m[14]&~m[36]&m[37])|(~m[14]&m[36]&m[37]))&~BiasedRNG[2])|((m[14]&m[36]&m[37]))):InitCond[2];
    m[3] = run?((((m[15]&~m[42]&~m[43])|(~m[15]&m[42]&~m[43])|(~m[15]&~m[42]&m[43]))&BiasedRNG[3])|(((m[15]&m[42]&~m[43])|(m[15]&~m[42]&m[43])|(~m[15]&m[42]&m[43]))&~BiasedRNG[3])|((m[15]&m[42]&m[43]))):InitCond[3];
    m[4] = run?((((m[16]&~m[48]&~m[49])|(~m[16]&m[48]&~m[49])|(~m[16]&~m[48]&m[49]))&BiasedRNG[4])|(((m[16]&m[48]&~m[49])|(m[16]&~m[48]&m[49])|(~m[16]&m[48]&m[49]))&~BiasedRNG[4])|((m[16]&m[48]&m[49]))):InitCond[4];
    m[5] = run?((((m[17]&~m[54]&~m[55])|(~m[17]&m[54]&~m[55])|(~m[17]&~m[54]&m[55]))&BiasedRNG[5])|(((m[17]&m[54]&~m[55])|(m[17]&~m[54]&m[55])|(~m[17]&m[54]&m[55]))&~BiasedRNG[5])|((m[17]&m[54]&m[55]))):InitCond[5];
    m[6] = run?((((m[18]&~m[60]&~m[61])|(~m[18]&m[60]&~m[61])|(~m[18]&~m[60]&m[61]))&BiasedRNG[6])|(((m[18]&m[60]&~m[61])|(m[18]&~m[60]&m[61])|(~m[18]&m[60]&m[61]))&~BiasedRNG[6])|((m[18]&m[60]&m[61]))):InitCond[6];
    m[7] = run?((((m[19]&~m[66]&~m[67])|(~m[19]&m[66]&~m[67])|(~m[19]&~m[66]&m[67]))&BiasedRNG[7])|(((m[19]&m[66]&~m[67])|(m[19]&~m[66]&m[67])|(~m[19]&m[66]&m[67]))&~BiasedRNG[7])|((m[19]&m[66]&m[67]))):InitCond[7];
    m[8] = run?((((m[20]&~m[72]&~m[73])|(~m[20]&m[72]&~m[73])|(~m[20]&~m[72]&m[73]))&BiasedRNG[8])|(((m[20]&m[72]&~m[73])|(m[20]&~m[72]&m[73])|(~m[20]&m[72]&m[73]))&~BiasedRNG[8])|((m[20]&m[72]&m[73]))):InitCond[8];
    m[9] = run?((((m[21]&~m[78]&~m[79])|(~m[21]&m[78]&~m[79])|(~m[21]&~m[78]&m[79]))&BiasedRNG[9])|(((m[21]&m[78]&~m[79])|(m[21]&~m[78]&m[79])|(~m[21]&m[78]&m[79]))&~BiasedRNG[9])|((m[21]&m[78]&m[79]))):InitCond[9];
    m[10] = run?((((m[22]&~m[84]&~m[85])|(~m[22]&m[84]&~m[85])|(~m[22]&~m[84]&m[85]))&BiasedRNG[10])|(((m[22]&m[84]&~m[85])|(m[22]&~m[84]&m[85])|(~m[22]&m[84]&m[85]))&~BiasedRNG[10])|((m[22]&m[84]&m[85]))):InitCond[10];
    m[11] = run?((((m[23]&~m[90]&~m[91])|(~m[23]&m[90]&~m[91])|(~m[23]&~m[90]&m[91]))&BiasedRNG[11])|(((m[23]&m[90]&~m[91])|(m[23]&~m[90]&m[91])|(~m[23]&m[90]&m[91]))&~BiasedRNG[11])|((m[23]&m[90]&m[91]))):InitCond[11];
    m[26] = run?((((~m[12]&~m[72]&~m[108])|(m[12]&m[72]&~m[108]))&BiasedRNG[12])|(((m[12]&~m[72]&~m[108])|(~m[12]&m[72]&m[108]))&~BiasedRNG[12])|((~m[12]&~m[72]&m[108])|(m[12]&~m[72]&m[108])|(m[12]&m[72]&m[108]))):InitCond[12];
    m[27] = run?((((~m[12]&~m[78]&~m[114])|(m[12]&m[78]&~m[114]))&BiasedRNG[13])|(((m[12]&~m[78]&~m[114])|(~m[12]&m[78]&m[114]))&~BiasedRNG[13])|((~m[12]&~m[78]&m[114])|(m[12]&~m[78]&m[114])|(m[12]&m[78]&m[114]))):InitCond[13];
    m[28] = run?((((~m[12]&~m[84]&~m[120])|(m[12]&m[84]&~m[120]))&BiasedRNG[14])|(((m[12]&~m[84]&~m[120])|(~m[12]&m[84]&m[120]))&~BiasedRNG[14])|((~m[12]&~m[84]&m[120])|(m[12]&~m[84]&m[120])|(m[12]&m[84]&m[120]))):InitCond[14];
    m[29] = run?((((~m[12]&~m[90]&~m[126])|(m[12]&m[90]&~m[126]))&BiasedRNG[15])|(((m[12]&~m[90]&~m[126])|(~m[12]&m[90]&m[126]))&~BiasedRNG[15])|((~m[12]&~m[90]&m[126])|(m[12]&~m[90]&m[126])|(m[12]&m[90]&m[126]))):InitCond[15];
    m[32] = run?((((~m[13]&~m[73]&~m[109])|(m[13]&m[73]&~m[109]))&BiasedRNG[16])|(((m[13]&~m[73]&~m[109])|(~m[13]&m[73]&m[109]))&~BiasedRNG[16])|((~m[13]&~m[73]&m[109])|(m[13]&~m[73]&m[109])|(m[13]&m[73]&m[109]))):InitCond[16];
    m[33] = run?((((~m[13]&~m[79]&~m[115])|(m[13]&m[79]&~m[115]))&BiasedRNG[17])|(((m[13]&~m[79]&~m[115])|(~m[13]&m[79]&m[115]))&~BiasedRNG[17])|((~m[13]&~m[79]&m[115])|(m[13]&~m[79]&m[115])|(m[13]&m[79]&m[115]))):InitCond[17];
    m[34] = run?((((~m[13]&~m[85]&~m[121])|(m[13]&m[85]&~m[121]))&BiasedRNG[18])|(((m[13]&~m[85]&~m[121])|(~m[13]&m[85]&m[121]))&~BiasedRNG[18])|((~m[13]&~m[85]&m[121])|(m[13]&~m[85]&m[121])|(m[13]&m[85]&m[121]))):InitCond[18];
    m[35] = run?((((~m[13]&~m[91]&~m[127])|(m[13]&m[91]&~m[127]))&BiasedRNG[19])|(((m[13]&~m[91]&~m[127])|(~m[13]&m[91]&m[127]))&~BiasedRNG[19])|((~m[13]&~m[91]&m[127])|(m[13]&~m[91]&m[127])|(m[13]&m[91]&m[127]))):InitCond[19];
    m[38] = run?((((~m[14]&~m[74]&~m[110])|(m[14]&m[74]&~m[110]))&BiasedRNG[20])|(((m[14]&~m[74]&~m[110])|(~m[14]&m[74]&m[110]))&~BiasedRNG[20])|((~m[14]&~m[74]&m[110])|(m[14]&~m[74]&m[110])|(m[14]&m[74]&m[110]))):InitCond[20];
    m[39] = run?((((~m[14]&~m[80]&~m[116])|(m[14]&m[80]&~m[116]))&BiasedRNG[21])|(((m[14]&~m[80]&~m[116])|(~m[14]&m[80]&m[116]))&~BiasedRNG[21])|((~m[14]&~m[80]&m[116])|(m[14]&~m[80]&m[116])|(m[14]&m[80]&m[116]))):InitCond[21];
    m[40] = run?((((~m[14]&~m[86]&~m[122])|(m[14]&m[86]&~m[122]))&BiasedRNG[22])|(((m[14]&~m[86]&~m[122])|(~m[14]&m[86]&m[122]))&~BiasedRNG[22])|((~m[14]&~m[86]&m[122])|(m[14]&~m[86]&m[122])|(m[14]&m[86]&m[122]))):InitCond[22];
    m[41] = run?((((~m[14]&~m[92]&~m[128])|(m[14]&m[92]&~m[128]))&BiasedRNG[23])|(((m[14]&~m[92]&~m[128])|(~m[14]&m[92]&m[128]))&~BiasedRNG[23])|((~m[14]&~m[92]&m[128])|(m[14]&~m[92]&m[128])|(m[14]&m[92]&m[128]))):InitCond[23];
    m[44] = run?((((~m[15]&~m[75]&~m[111])|(m[15]&m[75]&~m[111]))&BiasedRNG[24])|(((m[15]&~m[75]&~m[111])|(~m[15]&m[75]&m[111]))&~BiasedRNG[24])|((~m[15]&~m[75]&m[111])|(m[15]&~m[75]&m[111])|(m[15]&m[75]&m[111]))):InitCond[24];
    m[45] = run?((((~m[15]&~m[81]&~m[117])|(m[15]&m[81]&~m[117]))&BiasedRNG[25])|(((m[15]&~m[81]&~m[117])|(~m[15]&m[81]&m[117]))&~BiasedRNG[25])|((~m[15]&~m[81]&m[117])|(m[15]&~m[81]&m[117])|(m[15]&m[81]&m[117]))):InitCond[25];
    m[46] = run?((((~m[15]&~m[87]&~m[123])|(m[15]&m[87]&~m[123]))&BiasedRNG[26])|(((m[15]&~m[87]&~m[123])|(~m[15]&m[87]&m[123]))&~BiasedRNG[26])|((~m[15]&~m[87]&m[123])|(m[15]&~m[87]&m[123])|(m[15]&m[87]&m[123]))):InitCond[26];
    m[47] = run?((((~m[15]&~m[93]&~m[129])|(m[15]&m[93]&~m[129]))&BiasedRNG[27])|(((m[15]&~m[93]&~m[129])|(~m[15]&m[93]&m[129]))&~BiasedRNG[27])|((~m[15]&~m[93]&m[129])|(m[15]&~m[93]&m[129])|(m[15]&m[93]&m[129]))):InitCond[27];
    m[50] = run?((((~m[16]&~m[76]&~m[112])|(m[16]&m[76]&~m[112]))&BiasedRNG[28])|(((m[16]&~m[76]&~m[112])|(~m[16]&m[76]&m[112]))&~BiasedRNG[28])|((~m[16]&~m[76]&m[112])|(m[16]&~m[76]&m[112])|(m[16]&m[76]&m[112]))):InitCond[28];
    m[51] = run?((((~m[16]&~m[82]&~m[118])|(m[16]&m[82]&~m[118]))&BiasedRNG[29])|(((m[16]&~m[82]&~m[118])|(~m[16]&m[82]&m[118]))&~BiasedRNG[29])|((~m[16]&~m[82]&m[118])|(m[16]&~m[82]&m[118])|(m[16]&m[82]&m[118]))):InitCond[29];
    m[52] = run?((((~m[16]&~m[88]&~m[124])|(m[16]&m[88]&~m[124]))&BiasedRNG[30])|(((m[16]&~m[88]&~m[124])|(~m[16]&m[88]&m[124]))&~BiasedRNG[30])|((~m[16]&~m[88]&m[124])|(m[16]&~m[88]&m[124])|(m[16]&m[88]&m[124]))):InitCond[30];
    m[53] = run?((((~m[16]&~m[94]&~m[130])|(m[16]&m[94]&~m[130]))&BiasedRNG[31])|(((m[16]&~m[94]&~m[130])|(~m[16]&m[94]&m[130]))&~BiasedRNG[31])|((~m[16]&~m[94]&m[130])|(m[16]&~m[94]&m[130])|(m[16]&m[94]&m[130]))):InitCond[31];
    m[56] = run?((((~m[17]&~m[77]&~m[113])|(m[17]&m[77]&~m[113]))&BiasedRNG[32])|(((m[17]&~m[77]&~m[113])|(~m[17]&m[77]&m[113]))&~BiasedRNG[32])|((~m[17]&~m[77]&m[113])|(m[17]&~m[77]&m[113])|(m[17]&m[77]&m[113]))):InitCond[32];
    m[57] = run?((((~m[17]&~m[83]&~m[119])|(m[17]&m[83]&~m[119]))&BiasedRNG[33])|(((m[17]&~m[83]&~m[119])|(~m[17]&m[83]&m[119]))&~BiasedRNG[33])|((~m[17]&~m[83]&m[119])|(m[17]&~m[83]&m[119])|(m[17]&m[83]&m[119]))):InitCond[33];
    m[58] = run?((((~m[17]&~m[89]&~m[125])|(m[17]&m[89]&~m[125]))&BiasedRNG[34])|(((m[17]&~m[89]&~m[125])|(~m[17]&m[89]&m[125]))&~BiasedRNG[34])|((~m[17]&~m[89]&m[125])|(m[17]&~m[89]&m[125])|(m[17]&m[89]&m[125]))):InitCond[34];
    m[59] = run?((((~m[17]&~m[95]&~m[131])|(m[17]&m[95]&~m[131]))&BiasedRNG[35])|(((m[17]&~m[95]&~m[131])|(~m[17]&m[95]&m[131]))&~BiasedRNG[35])|((~m[17]&~m[95]&m[131])|(m[17]&~m[95]&m[131])|(m[17]&m[95]&m[131]))):InitCond[35];
    m[62] = run?((((~m[18]&~m[36]&~m[98])|(m[18]&m[36]&~m[98]))&BiasedRNG[36])|(((m[18]&~m[36]&~m[98])|(~m[18]&m[36]&m[98]))&~BiasedRNG[36])|((~m[18]&~m[36]&m[98])|(m[18]&~m[36]&m[98])|(m[18]&m[36]&m[98]))):InitCond[36];
    m[63] = run?((((~m[18]&~m[42]&~m[99])|(m[18]&m[42]&~m[99]))&BiasedRNG[37])|(((m[18]&~m[42]&~m[99])|(~m[18]&m[42]&m[99]))&~BiasedRNG[37])|((~m[18]&~m[42]&m[99])|(m[18]&~m[42]&m[99])|(m[18]&m[42]&m[99]))):InitCond[37];
    m[64] = run?((((~m[18]&~m[48]&~m[100])|(m[18]&m[48]&~m[100]))&BiasedRNG[38])|(((m[18]&~m[48]&~m[100])|(~m[18]&m[48]&m[100]))&~BiasedRNG[38])|((~m[18]&~m[48]&m[100])|(m[18]&~m[48]&m[100])|(m[18]&m[48]&m[100]))):InitCond[38];
    m[65] = run?((((~m[18]&~m[54]&~m[101])|(m[18]&m[54]&~m[101]))&BiasedRNG[39])|(((m[18]&~m[54]&~m[101])|(~m[18]&m[54]&m[101]))&~BiasedRNG[39])|((~m[18]&~m[54]&m[101])|(m[18]&~m[54]&m[101])|(m[18]&m[54]&m[101]))):InitCond[39];
    m[68] = run?((((~m[19]&~m[37]&~m[104])|(m[19]&m[37]&~m[104]))&BiasedRNG[40])|(((m[19]&~m[37]&~m[104])|(~m[19]&m[37]&m[104]))&~BiasedRNG[40])|((~m[19]&~m[37]&m[104])|(m[19]&~m[37]&m[104])|(m[19]&m[37]&m[104]))):InitCond[40];
    m[69] = run?((((~m[19]&~m[43]&~m[105])|(m[19]&m[43]&~m[105]))&BiasedRNG[41])|(((m[19]&~m[43]&~m[105])|(~m[19]&m[43]&m[105]))&~BiasedRNG[41])|((~m[19]&~m[43]&m[105])|(m[19]&~m[43]&m[105])|(m[19]&m[43]&m[105]))):InitCond[41];
    m[70] = run?((((~m[19]&~m[49]&~m[106])|(m[19]&m[49]&~m[106]))&BiasedRNG[42])|(((m[19]&~m[49]&~m[106])|(~m[19]&m[49]&m[106]))&~BiasedRNG[42])|((~m[19]&~m[49]&m[106])|(m[19]&~m[49]&m[106])|(m[19]&m[49]&m[106]))):InitCond[42];
    m[71] = run?((((~m[19]&~m[55]&~m[107])|(m[19]&m[55]&~m[107]))&BiasedRNG[43])|(((m[19]&~m[55]&~m[107])|(~m[19]&m[55]&m[107]))&~BiasedRNG[43])|((~m[19]&~m[55]&m[107])|(m[19]&~m[55]&m[107])|(m[19]&m[55]&m[107]))):InitCond[43];
    m[97] = run?((((m[30]&~m[61]&m[132])|(~m[30]&m[61]&m[132]))&BiasedRNG[44])|(((m[30]&m[61]&~m[132]))&~BiasedRNG[44])|((m[30]&m[61]&m[132]))):InitCond[44];
    m[102] = run?((((m[25]&~m[66]&m[133])|(~m[25]&m[66]&m[133]))&BiasedRNG[45])|(((m[25]&m[66]&~m[133]))&~BiasedRNG[45])|((m[25]&m[66]&m[133]))):InitCond[45];
    m[103] = run?((((m[31]&~m[67]&m[138])|(~m[31]&m[67]&m[138]))&BiasedRNG[46])|(((m[31]&m[67]&~m[138]))&~BiasedRNG[46])|((m[31]&m[67]&m[138]))):InitCond[46];
    m[137] = run?((((m[98]&~m[138]&~m[139]&~m[140]&~m[141])|(~m[98]&~m[138]&~m[139]&m[140]&~m[141])|(m[98]&m[138]&~m[139]&m[140]&~m[141])|(m[98]&~m[138]&m[139]&m[140]&~m[141])|(~m[98]&m[138]&~m[139]&~m[140]&m[141])|(~m[98]&~m[138]&m[139]&~m[140]&m[141])|(m[98]&m[138]&m[139]&~m[140]&m[141])|(~m[98]&m[138]&m[139]&m[140]&m[141]))&UnbiasedRNG[0])|((m[98]&~m[138]&~m[139]&m[140]&~m[141])|(~m[98]&~m[138]&~m[139]&~m[140]&m[141])|(m[98]&~m[138]&~m[139]&~m[140]&m[141])|(m[98]&m[138]&~m[139]&~m[140]&m[141])|(m[98]&~m[138]&m[139]&~m[140]&m[141])|(~m[98]&~m[138]&~m[139]&m[140]&m[141])|(m[98]&~m[138]&~m[139]&m[140]&m[141])|(~m[98]&m[138]&~m[139]&m[140]&m[141])|(m[98]&m[138]&~m[139]&m[140]&m[141])|(~m[98]&~m[138]&m[139]&m[140]&m[141])|(m[98]&~m[138]&m[139]&m[140]&m[141])|(m[98]&m[138]&m[139]&m[140]&m[141]))):InitCond[47];
    m[142] = run?((((m[140]&~m[143]&~m[144]&~m[145]&~m[146])|(~m[140]&~m[143]&~m[144]&m[145]&~m[146])|(m[140]&m[143]&~m[144]&m[145]&~m[146])|(m[140]&~m[143]&m[144]&m[145]&~m[146])|(~m[140]&m[143]&~m[144]&~m[145]&m[146])|(~m[140]&~m[143]&m[144]&~m[145]&m[146])|(m[140]&m[143]&m[144]&~m[145]&m[146])|(~m[140]&m[143]&m[144]&m[145]&m[146]))&UnbiasedRNG[1])|((m[140]&~m[143]&~m[144]&m[145]&~m[146])|(~m[140]&~m[143]&~m[144]&~m[145]&m[146])|(m[140]&~m[143]&~m[144]&~m[145]&m[146])|(m[140]&m[143]&~m[144]&~m[145]&m[146])|(m[140]&~m[143]&m[144]&~m[145]&m[146])|(~m[140]&~m[143]&~m[144]&m[145]&m[146])|(m[140]&~m[143]&~m[144]&m[145]&m[146])|(~m[140]&m[143]&~m[144]&m[145]&m[146])|(m[140]&m[143]&~m[144]&m[145]&m[146])|(~m[140]&~m[143]&m[144]&m[145]&m[146])|(m[140]&~m[143]&m[144]&m[145]&m[146])|(m[140]&m[143]&m[144]&m[145]&m[146]))):InitCond[48];
    m[147] = run?((((m[99]&~m[148]&~m[149]&~m[150]&~m[151])|(~m[99]&~m[148]&~m[149]&m[150]&~m[151])|(m[99]&m[148]&~m[149]&m[150]&~m[151])|(m[99]&~m[148]&m[149]&m[150]&~m[151])|(~m[99]&m[148]&~m[149]&~m[150]&m[151])|(~m[99]&~m[148]&m[149]&~m[150]&m[151])|(m[99]&m[148]&m[149]&~m[150]&m[151])|(~m[99]&m[148]&m[149]&m[150]&m[151]))&UnbiasedRNG[2])|((m[99]&~m[148]&~m[149]&m[150]&~m[151])|(~m[99]&~m[148]&~m[149]&~m[150]&m[151])|(m[99]&~m[148]&~m[149]&~m[150]&m[151])|(m[99]&m[148]&~m[149]&~m[150]&m[151])|(m[99]&~m[148]&m[149]&~m[150]&m[151])|(~m[99]&~m[148]&~m[149]&m[150]&m[151])|(m[99]&~m[148]&~m[149]&m[150]&m[151])|(~m[99]&m[148]&~m[149]&m[150]&m[151])|(m[99]&m[148]&~m[149]&m[150]&m[151])|(~m[99]&~m[148]&m[149]&m[150]&m[151])|(m[99]&~m[148]&m[149]&m[150]&m[151])|(m[99]&m[148]&m[149]&m[150]&m[151]))):InitCond[49];
    m[152] = run?((((m[150]&~m[153]&~m[154]&~m[155]&~m[156])|(~m[150]&~m[153]&~m[154]&m[155]&~m[156])|(m[150]&m[153]&~m[154]&m[155]&~m[156])|(m[150]&~m[153]&m[154]&m[155]&~m[156])|(~m[150]&m[153]&~m[154]&~m[155]&m[156])|(~m[150]&~m[153]&m[154]&~m[155]&m[156])|(m[150]&m[153]&m[154]&~m[155]&m[156])|(~m[150]&m[153]&m[154]&m[155]&m[156]))&UnbiasedRNG[3])|((m[150]&~m[153]&~m[154]&m[155]&~m[156])|(~m[150]&~m[153]&~m[154]&~m[155]&m[156])|(m[150]&~m[153]&~m[154]&~m[155]&m[156])|(m[150]&m[153]&~m[154]&~m[155]&m[156])|(m[150]&~m[153]&m[154]&~m[155]&m[156])|(~m[150]&~m[153]&~m[154]&m[155]&m[156])|(m[150]&~m[153]&~m[154]&m[155]&m[156])|(~m[150]&m[153]&~m[154]&m[155]&m[156])|(m[150]&m[153]&~m[154]&m[155]&m[156])|(~m[150]&~m[153]&m[154]&m[155]&m[156])|(m[150]&~m[153]&m[154]&m[155]&m[156])|(m[150]&m[153]&m[154]&m[155]&m[156]))):InitCond[50];
    m[157] = run?((((m[155]&~m[158]&~m[159]&~m[160]&~m[161])|(~m[155]&~m[158]&~m[159]&m[160]&~m[161])|(m[155]&m[158]&~m[159]&m[160]&~m[161])|(m[155]&~m[158]&m[159]&m[160]&~m[161])|(~m[155]&m[158]&~m[159]&~m[160]&m[161])|(~m[155]&~m[158]&m[159]&~m[160]&m[161])|(m[155]&m[158]&m[159]&~m[160]&m[161])|(~m[155]&m[158]&m[159]&m[160]&m[161]))&UnbiasedRNG[4])|((m[155]&~m[158]&~m[159]&m[160]&~m[161])|(~m[155]&~m[158]&~m[159]&~m[160]&m[161])|(m[155]&~m[158]&~m[159]&~m[160]&m[161])|(m[155]&m[158]&~m[159]&~m[160]&m[161])|(m[155]&~m[158]&m[159]&~m[160]&m[161])|(~m[155]&~m[158]&~m[159]&m[160]&m[161])|(m[155]&~m[158]&~m[159]&m[160]&m[161])|(~m[155]&m[158]&~m[159]&m[160]&m[161])|(m[155]&m[158]&~m[159]&m[160]&m[161])|(~m[155]&~m[158]&m[159]&m[160]&m[161])|(m[155]&~m[158]&m[159]&m[160]&m[161])|(m[155]&m[158]&m[159]&m[160]&m[161]))):InitCond[51];
    m[162] = run?((((m[100]&~m[163]&~m[164]&~m[165]&~m[166])|(~m[100]&~m[163]&~m[164]&m[165]&~m[166])|(m[100]&m[163]&~m[164]&m[165]&~m[166])|(m[100]&~m[163]&m[164]&m[165]&~m[166])|(~m[100]&m[163]&~m[164]&~m[165]&m[166])|(~m[100]&~m[163]&m[164]&~m[165]&m[166])|(m[100]&m[163]&m[164]&~m[165]&m[166])|(~m[100]&m[163]&m[164]&m[165]&m[166]))&UnbiasedRNG[5])|((m[100]&~m[163]&~m[164]&m[165]&~m[166])|(~m[100]&~m[163]&~m[164]&~m[165]&m[166])|(m[100]&~m[163]&~m[164]&~m[165]&m[166])|(m[100]&m[163]&~m[164]&~m[165]&m[166])|(m[100]&~m[163]&m[164]&~m[165]&m[166])|(~m[100]&~m[163]&~m[164]&m[165]&m[166])|(m[100]&~m[163]&~m[164]&m[165]&m[166])|(~m[100]&m[163]&~m[164]&m[165]&m[166])|(m[100]&m[163]&~m[164]&m[165]&m[166])|(~m[100]&~m[163]&m[164]&m[165]&m[166])|(m[100]&~m[163]&m[164]&m[165]&m[166])|(m[100]&m[163]&m[164]&m[165]&m[166]))):InitCond[52];
    m[167] = run?((((m[165]&~m[168]&~m[169]&~m[170]&~m[171])|(~m[165]&~m[168]&~m[169]&m[170]&~m[171])|(m[165]&m[168]&~m[169]&m[170]&~m[171])|(m[165]&~m[168]&m[169]&m[170]&~m[171])|(~m[165]&m[168]&~m[169]&~m[170]&m[171])|(~m[165]&~m[168]&m[169]&~m[170]&m[171])|(m[165]&m[168]&m[169]&~m[170]&m[171])|(~m[165]&m[168]&m[169]&m[170]&m[171]))&UnbiasedRNG[6])|((m[165]&~m[168]&~m[169]&m[170]&~m[171])|(~m[165]&~m[168]&~m[169]&~m[170]&m[171])|(m[165]&~m[168]&~m[169]&~m[170]&m[171])|(m[165]&m[168]&~m[169]&~m[170]&m[171])|(m[165]&~m[168]&m[169]&~m[170]&m[171])|(~m[165]&~m[168]&~m[169]&m[170]&m[171])|(m[165]&~m[168]&~m[169]&m[170]&m[171])|(~m[165]&m[168]&~m[169]&m[170]&m[171])|(m[165]&m[168]&~m[169]&m[170]&m[171])|(~m[165]&~m[168]&m[169]&m[170]&m[171])|(m[165]&~m[168]&m[169]&m[170]&m[171])|(m[165]&m[168]&m[169]&m[170]&m[171]))):InitCond[53];
    m[172] = run?((((m[170]&~m[173]&~m[174]&~m[175]&~m[176])|(~m[170]&~m[173]&~m[174]&m[175]&~m[176])|(m[170]&m[173]&~m[174]&m[175]&~m[176])|(m[170]&~m[173]&m[174]&m[175]&~m[176])|(~m[170]&m[173]&~m[174]&~m[175]&m[176])|(~m[170]&~m[173]&m[174]&~m[175]&m[176])|(m[170]&m[173]&m[174]&~m[175]&m[176])|(~m[170]&m[173]&m[174]&m[175]&m[176]))&UnbiasedRNG[7])|((m[170]&~m[173]&~m[174]&m[175]&~m[176])|(~m[170]&~m[173]&~m[174]&~m[175]&m[176])|(m[170]&~m[173]&~m[174]&~m[175]&m[176])|(m[170]&m[173]&~m[174]&~m[175]&m[176])|(m[170]&~m[173]&m[174]&~m[175]&m[176])|(~m[170]&~m[173]&~m[174]&m[175]&m[176])|(m[170]&~m[173]&~m[174]&m[175]&m[176])|(~m[170]&m[173]&~m[174]&m[175]&m[176])|(m[170]&m[173]&~m[174]&m[175]&m[176])|(~m[170]&~m[173]&m[174]&m[175]&m[176])|(m[170]&~m[173]&m[174]&m[175]&m[176])|(m[170]&m[173]&m[174]&m[175]&m[176]))):InitCond[54];
    m[177] = run?((((m[175]&~m[178]&~m[179]&~m[180]&~m[181])|(~m[175]&~m[178]&~m[179]&m[180]&~m[181])|(m[175]&m[178]&~m[179]&m[180]&~m[181])|(m[175]&~m[178]&m[179]&m[180]&~m[181])|(~m[175]&m[178]&~m[179]&~m[180]&m[181])|(~m[175]&~m[178]&m[179]&~m[180]&m[181])|(m[175]&m[178]&m[179]&~m[180]&m[181])|(~m[175]&m[178]&m[179]&m[180]&m[181]))&UnbiasedRNG[8])|((m[175]&~m[178]&~m[179]&m[180]&~m[181])|(~m[175]&~m[178]&~m[179]&~m[180]&m[181])|(m[175]&~m[178]&~m[179]&~m[180]&m[181])|(m[175]&m[178]&~m[179]&~m[180]&m[181])|(m[175]&~m[178]&m[179]&~m[180]&m[181])|(~m[175]&~m[178]&~m[179]&m[180]&m[181])|(m[175]&~m[178]&~m[179]&m[180]&m[181])|(~m[175]&m[178]&~m[179]&m[180]&m[181])|(m[175]&m[178]&~m[179]&m[180]&m[181])|(~m[175]&~m[178]&m[179]&m[180]&m[181])|(m[175]&~m[178]&m[179]&m[180]&m[181])|(m[175]&m[178]&m[179]&m[180]&m[181]))):InitCond[55];
    m[182] = run?((((m[101]&~m[183]&~m[184]&~m[185]&~m[186])|(~m[101]&~m[183]&~m[184]&m[185]&~m[186])|(m[101]&m[183]&~m[184]&m[185]&~m[186])|(m[101]&~m[183]&m[184]&m[185]&~m[186])|(~m[101]&m[183]&~m[184]&~m[185]&m[186])|(~m[101]&~m[183]&m[184]&~m[185]&m[186])|(m[101]&m[183]&m[184]&~m[185]&m[186])|(~m[101]&m[183]&m[184]&m[185]&m[186]))&UnbiasedRNG[9])|((m[101]&~m[183]&~m[184]&m[185]&~m[186])|(~m[101]&~m[183]&~m[184]&~m[185]&m[186])|(m[101]&~m[183]&~m[184]&~m[185]&m[186])|(m[101]&m[183]&~m[184]&~m[185]&m[186])|(m[101]&~m[183]&m[184]&~m[185]&m[186])|(~m[101]&~m[183]&~m[184]&m[185]&m[186])|(m[101]&~m[183]&~m[184]&m[185]&m[186])|(~m[101]&m[183]&~m[184]&m[185]&m[186])|(m[101]&m[183]&~m[184]&m[185]&m[186])|(~m[101]&~m[183]&m[184]&m[185]&m[186])|(m[101]&~m[183]&m[184]&m[185]&m[186])|(m[101]&m[183]&m[184]&m[185]&m[186]))):InitCond[56];
    m[187] = run?((((m[185]&~m[188]&~m[189]&~m[190]&~m[191])|(~m[185]&~m[188]&~m[189]&m[190]&~m[191])|(m[185]&m[188]&~m[189]&m[190]&~m[191])|(m[185]&~m[188]&m[189]&m[190]&~m[191])|(~m[185]&m[188]&~m[189]&~m[190]&m[191])|(~m[185]&~m[188]&m[189]&~m[190]&m[191])|(m[185]&m[188]&m[189]&~m[190]&m[191])|(~m[185]&m[188]&m[189]&m[190]&m[191]))&UnbiasedRNG[10])|((m[185]&~m[188]&~m[189]&m[190]&~m[191])|(~m[185]&~m[188]&~m[189]&~m[190]&m[191])|(m[185]&~m[188]&~m[189]&~m[190]&m[191])|(m[185]&m[188]&~m[189]&~m[190]&m[191])|(m[185]&~m[188]&m[189]&~m[190]&m[191])|(~m[185]&~m[188]&~m[189]&m[190]&m[191])|(m[185]&~m[188]&~m[189]&m[190]&m[191])|(~m[185]&m[188]&~m[189]&m[190]&m[191])|(m[185]&m[188]&~m[189]&m[190]&m[191])|(~m[185]&~m[188]&m[189]&m[190]&m[191])|(m[185]&~m[188]&m[189]&m[190]&m[191])|(m[185]&m[188]&m[189]&m[190]&m[191]))):InitCond[57];
    m[192] = run?((((m[190]&~m[193]&~m[194]&~m[195]&~m[196])|(~m[190]&~m[193]&~m[194]&m[195]&~m[196])|(m[190]&m[193]&~m[194]&m[195]&~m[196])|(m[190]&~m[193]&m[194]&m[195]&~m[196])|(~m[190]&m[193]&~m[194]&~m[195]&m[196])|(~m[190]&~m[193]&m[194]&~m[195]&m[196])|(m[190]&m[193]&m[194]&~m[195]&m[196])|(~m[190]&m[193]&m[194]&m[195]&m[196]))&UnbiasedRNG[11])|((m[190]&~m[193]&~m[194]&m[195]&~m[196])|(~m[190]&~m[193]&~m[194]&~m[195]&m[196])|(m[190]&~m[193]&~m[194]&~m[195]&m[196])|(m[190]&m[193]&~m[194]&~m[195]&m[196])|(m[190]&~m[193]&m[194]&~m[195]&m[196])|(~m[190]&~m[193]&~m[194]&m[195]&m[196])|(m[190]&~m[193]&~m[194]&m[195]&m[196])|(~m[190]&m[193]&~m[194]&m[195]&m[196])|(m[190]&m[193]&~m[194]&m[195]&m[196])|(~m[190]&~m[193]&m[194]&m[195]&m[196])|(m[190]&~m[193]&m[194]&m[195]&m[196])|(m[190]&m[193]&m[194]&m[195]&m[196]))):InitCond[58];
    m[197] = run?((((m[195]&~m[198]&~m[199]&~m[200]&~m[201])|(~m[195]&~m[198]&~m[199]&m[200]&~m[201])|(m[195]&m[198]&~m[199]&m[200]&~m[201])|(m[195]&~m[198]&m[199]&m[200]&~m[201])|(~m[195]&m[198]&~m[199]&~m[200]&m[201])|(~m[195]&~m[198]&m[199]&~m[200]&m[201])|(m[195]&m[198]&m[199]&~m[200]&m[201])|(~m[195]&m[198]&m[199]&m[200]&m[201]))&UnbiasedRNG[12])|((m[195]&~m[198]&~m[199]&m[200]&~m[201])|(~m[195]&~m[198]&~m[199]&~m[200]&m[201])|(m[195]&~m[198]&~m[199]&~m[200]&m[201])|(m[195]&m[198]&~m[199]&~m[200]&m[201])|(m[195]&~m[198]&m[199]&~m[200]&m[201])|(~m[195]&~m[198]&~m[199]&m[200]&m[201])|(m[195]&~m[198]&~m[199]&m[200]&m[201])|(~m[195]&m[198]&~m[199]&m[200]&m[201])|(m[195]&m[198]&~m[199]&m[200]&m[201])|(~m[195]&~m[198]&m[199]&m[200]&m[201])|(m[195]&~m[198]&m[199]&m[200]&m[201])|(m[195]&m[198]&m[199]&m[200]&m[201]))):InitCond[59];
    m[202] = run?((((m[200]&~m[203]&~m[204]&~m[205]&~m[206])|(~m[200]&~m[203]&~m[204]&m[205]&~m[206])|(m[200]&m[203]&~m[204]&m[205]&~m[206])|(m[200]&~m[203]&m[204]&m[205]&~m[206])|(~m[200]&m[203]&~m[204]&~m[205]&m[206])|(~m[200]&~m[203]&m[204]&~m[205]&m[206])|(m[200]&m[203]&m[204]&~m[205]&m[206])|(~m[200]&m[203]&m[204]&m[205]&m[206]))&UnbiasedRNG[13])|((m[200]&~m[203]&~m[204]&m[205]&~m[206])|(~m[200]&~m[203]&~m[204]&~m[205]&m[206])|(m[200]&~m[203]&~m[204]&~m[205]&m[206])|(m[200]&m[203]&~m[204]&~m[205]&m[206])|(m[200]&~m[203]&m[204]&~m[205]&m[206])|(~m[200]&~m[203]&~m[204]&m[205]&m[206])|(m[200]&~m[203]&~m[204]&m[205]&m[206])|(~m[200]&m[203]&~m[204]&m[205]&m[206])|(m[200]&m[203]&~m[204]&m[205]&m[206])|(~m[200]&~m[203]&m[204]&m[205]&m[206])|(m[200]&~m[203]&m[204]&m[205]&m[206])|(m[200]&m[203]&m[204]&m[205]&m[206]))):InitCond[60];
    m[212] = run?((((m[210]&~m[213]&~m[214]&~m[215]&~m[216])|(~m[210]&~m[213]&~m[214]&m[215]&~m[216])|(m[210]&m[213]&~m[214]&m[215]&~m[216])|(m[210]&~m[213]&m[214]&m[215]&~m[216])|(~m[210]&m[213]&~m[214]&~m[215]&m[216])|(~m[210]&~m[213]&m[214]&~m[215]&m[216])|(m[210]&m[213]&m[214]&~m[215]&m[216])|(~m[210]&m[213]&m[214]&m[215]&m[216]))&UnbiasedRNG[14])|((m[210]&~m[213]&~m[214]&m[215]&~m[216])|(~m[210]&~m[213]&~m[214]&~m[215]&m[216])|(m[210]&~m[213]&~m[214]&~m[215]&m[216])|(m[210]&m[213]&~m[214]&~m[215]&m[216])|(m[210]&~m[213]&m[214]&~m[215]&m[216])|(~m[210]&~m[213]&~m[214]&m[215]&m[216])|(m[210]&~m[213]&~m[214]&m[215]&m[216])|(~m[210]&m[213]&~m[214]&m[215]&m[216])|(m[210]&m[213]&~m[214]&m[215]&m[216])|(~m[210]&~m[213]&m[214]&m[215]&m[216])|(m[210]&~m[213]&m[214]&m[215]&m[216])|(m[210]&m[213]&m[214]&m[215]&m[216]))):InitCond[61];
    m[217] = run?((((m[215]&~m[218]&~m[219]&~m[220]&~m[221])|(~m[215]&~m[218]&~m[219]&m[220]&~m[221])|(m[215]&m[218]&~m[219]&m[220]&~m[221])|(m[215]&~m[218]&m[219]&m[220]&~m[221])|(~m[215]&m[218]&~m[219]&~m[220]&m[221])|(~m[215]&~m[218]&m[219]&~m[220]&m[221])|(m[215]&m[218]&m[219]&~m[220]&m[221])|(~m[215]&m[218]&m[219]&m[220]&m[221]))&UnbiasedRNG[15])|((m[215]&~m[218]&~m[219]&m[220]&~m[221])|(~m[215]&~m[218]&~m[219]&~m[220]&m[221])|(m[215]&~m[218]&~m[219]&~m[220]&m[221])|(m[215]&m[218]&~m[219]&~m[220]&m[221])|(m[215]&~m[218]&m[219]&~m[220]&m[221])|(~m[215]&~m[218]&~m[219]&m[220]&m[221])|(m[215]&~m[218]&~m[219]&m[220]&m[221])|(~m[215]&m[218]&~m[219]&m[220]&m[221])|(m[215]&m[218]&~m[219]&m[220]&m[221])|(~m[215]&~m[218]&m[219]&m[220]&m[221])|(m[215]&~m[218]&m[219]&m[220]&m[221])|(m[215]&m[218]&m[219]&m[220]&m[221]))):InitCond[62];
    m[222] = run?((((m[220]&~m[223]&~m[224]&~m[225]&~m[226])|(~m[220]&~m[223]&~m[224]&m[225]&~m[226])|(m[220]&m[223]&~m[224]&m[225]&~m[226])|(m[220]&~m[223]&m[224]&m[225]&~m[226])|(~m[220]&m[223]&~m[224]&~m[225]&m[226])|(~m[220]&~m[223]&m[224]&~m[225]&m[226])|(m[220]&m[223]&m[224]&~m[225]&m[226])|(~m[220]&m[223]&m[224]&m[225]&m[226]))&UnbiasedRNG[16])|((m[220]&~m[223]&~m[224]&m[225]&~m[226])|(~m[220]&~m[223]&~m[224]&~m[225]&m[226])|(m[220]&~m[223]&~m[224]&~m[225]&m[226])|(m[220]&m[223]&~m[224]&~m[225]&m[226])|(m[220]&~m[223]&m[224]&~m[225]&m[226])|(~m[220]&~m[223]&~m[224]&m[225]&m[226])|(m[220]&~m[223]&~m[224]&m[225]&m[226])|(~m[220]&m[223]&~m[224]&m[225]&m[226])|(m[220]&m[223]&~m[224]&m[225]&m[226])|(~m[220]&~m[223]&m[224]&m[225]&m[226])|(m[220]&~m[223]&m[224]&m[225]&m[226])|(m[220]&m[223]&m[224]&m[225]&m[226]))):InitCond[63];
    m[227] = run?((((m[225]&~m[228]&~m[229]&~m[230]&~m[231])|(~m[225]&~m[228]&~m[229]&m[230]&~m[231])|(m[225]&m[228]&~m[229]&m[230]&~m[231])|(m[225]&~m[228]&m[229]&m[230]&~m[231])|(~m[225]&m[228]&~m[229]&~m[230]&m[231])|(~m[225]&~m[228]&m[229]&~m[230]&m[231])|(m[225]&m[228]&m[229]&~m[230]&m[231])|(~m[225]&m[228]&m[229]&m[230]&m[231]))&UnbiasedRNG[17])|((m[225]&~m[228]&~m[229]&m[230]&~m[231])|(~m[225]&~m[228]&~m[229]&~m[230]&m[231])|(m[225]&~m[228]&~m[229]&~m[230]&m[231])|(m[225]&m[228]&~m[229]&~m[230]&m[231])|(m[225]&~m[228]&m[229]&~m[230]&m[231])|(~m[225]&~m[228]&~m[229]&m[230]&m[231])|(m[225]&~m[228]&~m[229]&m[230]&m[231])|(~m[225]&m[228]&~m[229]&m[230]&m[231])|(m[225]&m[228]&~m[229]&m[230]&m[231])|(~m[225]&~m[228]&m[229]&m[230]&m[231])|(m[225]&~m[228]&m[229]&m[230]&m[231])|(m[225]&m[228]&m[229]&m[230]&m[231]))):InitCond[64];
    m[232] = run?((((m[211]&~m[233]&~m[234]&~m[235]&~m[236])|(~m[211]&~m[233]&~m[234]&m[235]&~m[236])|(m[211]&m[233]&~m[234]&m[235]&~m[236])|(m[211]&~m[233]&m[234]&m[235]&~m[236])|(~m[211]&m[233]&~m[234]&~m[235]&m[236])|(~m[211]&~m[233]&m[234]&~m[235]&m[236])|(m[211]&m[233]&m[234]&~m[235]&m[236])|(~m[211]&m[233]&m[234]&m[235]&m[236]))&UnbiasedRNG[18])|((m[211]&~m[233]&~m[234]&m[235]&~m[236])|(~m[211]&~m[233]&~m[234]&~m[235]&m[236])|(m[211]&~m[233]&~m[234]&~m[235]&m[236])|(m[211]&m[233]&~m[234]&~m[235]&m[236])|(m[211]&~m[233]&m[234]&~m[235]&m[236])|(~m[211]&~m[233]&~m[234]&m[235]&m[236])|(m[211]&~m[233]&~m[234]&m[235]&m[236])|(~m[211]&m[233]&~m[234]&m[235]&m[236])|(m[211]&m[233]&~m[234]&m[235]&m[236])|(~m[211]&~m[233]&m[234]&m[235]&m[236])|(m[211]&~m[233]&m[234]&m[235]&m[236])|(m[211]&m[233]&m[234]&m[235]&m[236]))):InitCond[65];
    m[237] = run?((((m[235]&~m[238]&~m[239]&~m[240]&~m[241])|(~m[235]&~m[238]&~m[239]&m[240]&~m[241])|(m[235]&m[238]&~m[239]&m[240]&~m[241])|(m[235]&~m[238]&m[239]&m[240]&~m[241])|(~m[235]&m[238]&~m[239]&~m[240]&m[241])|(~m[235]&~m[238]&m[239]&~m[240]&m[241])|(m[235]&m[238]&m[239]&~m[240]&m[241])|(~m[235]&m[238]&m[239]&m[240]&m[241]))&UnbiasedRNG[19])|((m[235]&~m[238]&~m[239]&m[240]&~m[241])|(~m[235]&~m[238]&~m[239]&~m[240]&m[241])|(m[235]&~m[238]&~m[239]&~m[240]&m[241])|(m[235]&m[238]&~m[239]&~m[240]&m[241])|(m[235]&~m[238]&m[239]&~m[240]&m[241])|(~m[235]&~m[238]&~m[239]&m[240]&m[241])|(m[235]&~m[238]&~m[239]&m[240]&m[241])|(~m[235]&m[238]&~m[239]&m[240]&m[241])|(m[235]&m[238]&~m[239]&m[240]&m[241])|(~m[235]&~m[238]&m[239]&m[240]&m[241])|(m[235]&~m[238]&m[239]&m[240]&m[241])|(m[235]&m[238]&m[239]&m[240]&m[241]))):InitCond[66];
    m[242] = run?((((m[240]&~m[243]&~m[244]&~m[245]&~m[246])|(~m[240]&~m[243]&~m[244]&m[245]&~m[246])|(m[240]&m[243]&~m[244]&m[245]&~m[246])|(m[240]&~m[243]&m[244]&m[245]&~m[246])|(~m[240]&m[243]&~m[244]&~m[245]&m[246])|(~m[240]&~m[243]&m[244]&~m[245]&m[246])|(m[240]&m[243]&m[244]&~m[245]&m[246])|(~m[240]&m[243]&m[244]&m[245]&m[246]))&UnbiasedRNG[20])|((m[240]&~m[243]&~m[244]&m[245]&~m[246])|(~m[240]&~m[243]&~m[244]&~m[245]&m[246])|(m[240]&~m[243]&~m[244]&~m[245]&m[246])|(m[240]&m[243]&~m[244]&~m[245]&m[246])|(m[240]&~m[243]&m[244]&~m[245]&m[246])|(~m[240]&~m[243]&~m[244]&m[245]&m[246])|(m[240]&~m[243]&~m[244]&m[245]&m[246])|(~m[240]&m[243]&~m[244]&m[245]&m[246])|(m[240]&m[243]&~m[244]&m[245]&m[246])|(~m[240]&~m[243]&m[244]&m[245]&m[246])|(m[240]&~m[243]&m[244]&m[245]&m[246])|(m[240]&m[243]&m[244]&m[245]&m[246]))):InitCond[67];
    m[247] = run?((((m[245]&~m[248]&~m[249]&~m[250]&~m[251])|(~m[245]&~m[248]&~m[249]&m[250]&~m[251])|(m[245]&m[248]&~m[249]&m[250]&~m[251])|(m[245]&~m[248]&m[249]&m[250]&~m[251])|(~m[245]&m[248]&~m[249]&~m[250]&m[251])|(~m[245]&~m[248]&m[249]&~m[250]&m[251])|(m[245]&m[248]&m[249]&~m[250]&m[251])|(~m[245]&m[248]&m[249]&m[250]&m[251]))&UnbiasedRNG[21])|((m[245]&~m[248]&~m[249]&m[250]&~m[251])|(~m[245]&~m[248]&~m[249]&~m[250]&m[251])|(m[245]&~m[248]&~m[249]&~m[250]&m[251])|(m[245]&m[248]&~m[249]&~m[250]&m[251])|(m[245]&~m[248]&m[249]&~m[250]&m[251])|(~m[245]&~m[248]&~m[249]&m[250]&m[251])|(m[245]&~m[248]&~m[249]&m[250]&m[251])|(~m[245]&m[248]&~m[249]&m[250]&m[251])|(m[245]&m[248]&~m[249]&m[250]&m[251])|(~m[245]&~m[248]&m[249]&m[250]&m[251])|(m[245]&~m[248]&m[249]&m[250]&m[251])|(m[245]&m[248]&m[249]&m[250]&m[251]))):InitCond[68];
    m[252] = run?((((m[236]&~m[253]&~m[254]&~m[255]&~m[256])|(~m[236]&~m[253]&~m[254]&m[255]&~m[256])|(m[236]&m[253]&~m[254]&m[255]&~m[256])|(m[236]&~m[253]&m[254]&m[255]&~m[256])|(~m[236]&m[253]&~m[254]&~m[255]&m[256])|(~m[236]&~m[253]&m[254]&~m[255]&m[256])|(m[236]&m[253]&m[254]&~m[255]&m[256])|(~m[236]&m[253]&m[254]&m[255]&m[256]))&UnbiasedRNG[22])|((m[236]&~m[253]&~m[254]&m[255]&~m[256])|(~m[236]&~m[253]&~m[254]&~m[255]&m[256])|(m[236]&~m[253]&~m[254]&~m[255]&m[256])|(m[236]&m[253]&~m[254]&~m[255]&m[256])|(m[236]&~m[253]&m[254]&~m[255]&m[256])|(~m[236]&~m[253]&~m[254]&m[255]&m[256])|(m[236]&~m[253]&~m[254]&m[255]&m[256])|(~m[236]&m[253]&~m[254]&m[255]&m[256])|(m[236]&m[253]&~m[254]&m[255]&m[256])|(~m[236]&~m[253]&m[254]&m[255]&m[256])|(m[236]&~m[253]&m[254]&m[255]&m[256])|(m[236]&m[253]&m[254]&m[255]&m[256]))):InitCond[69];
    m[257] = run?((((m[255]&~m[258]&~m[259]&~m[260]&~m[261])|(~m[255]&~m[258]&~m[259]&m[260]&~m[261])|(m[255]&m[258]&~m[259]&m[260]&~m[261])|(m[255]&~m[258]&m[259]&m[260]&~m[261])|(~m[255]&m[258]&~m[259]&~m[260]&m[261])|(~m[255]&~m[258]&m[259]&~m[260]&m[261])|(m[255]&m[258]&m[259]&~m[260]&m[261])|(~m[255]&m[258]&m[259]&m[260]&m[261]))&UnbiasedRNG[23])|((m[255]&~m[258]&~m[259]&m[260]&~m[261])|(~m[255]&~m[258]&~m[259]&~m[260]&m[261])|(m[255]&~m[258]&~m[259]&~m[260]&m[261])|(m[255]&m[258]&~m[259]&~m[260]&m[261])|(m[255]&~m[258]&m[259]&~m[260]&m[261])|(~m[255]&~m[258]&~m[259]&m[260]&m[261])|(m[255]&~m[258]&~m[259]&m[260]&m[261])|(~m[255]&m[258]&~m[259]&m[260]&m[261])|(m[255]&m[258]&~m[259]&m[260]&m[261])|(~m[255]&~m[258]&m[259]&m[260]&m[261])|(m[255]&~m[258]&m[259]&m[260]&m[261])|(m[255]&m[258]&m[259]&m[260]&m[261]))):InitCond[70];
    m[262] = run?((((m[260]&~m[263]&~m[264]&~m[265]&~m[266])|(~m[260]&~m[263]&~m[264]&m[265]&~m[266])|(m[260]&m[263]&~m[264]&m[265]&~m[266])|(m[260]&~m[263]&m[264]&m[265]&~m[266])|(~m[260]&m[263]&~m[264]&~m[265]&m[266])|(~m[260]&~m[263]&m[264]&~m[265]&m[266])|(m[260]&m[263]&m[264]&~m[265]&m[266])|(~m[260]&m[263]&m[264]&m[265]&m[266]))&UnbiasedRNG[24])|((m[260]&~m[263]&~m[264]&m[265]&~m[266])|(~m[260]&~m[263]&~m[264]&~m[265]&m[266])|(m[260]&~m[263]&~m[264]&~m[265]&m[266])|(m[260]&m[263]&~m[264]&~m[265]&m[266])|(m[260]&~m[263]&m[264]&~m[265]&m[266])|(~m[260]&~m[263]&~m[264]&m[265]&m[266])|(m[260]&~m[263]&~m[264]&m[265]&m[266])|(~m[260]&m[263]&~m[264]&m[265]&m[266])|(m[260]&m[263]&~m[264]&m[265]&m[266])|(~m[260]&~m[263]&m[264]&m[265]&m[266])|(m[260]&~m[263]&m[264]&m[265]&m[266])|(m[260]&m[263]&m[264]&m[265]&m[266]))):InitCond[71];
    m[267] = run?((((m[256]&~m[268]&~m[269]&~m[270]&~m[271])|(~m[256]&~m[268]&~m[269]&m[270]&~m[271])|(m[256]&m[268]&~m[269]&m[270]&~m[271])|(m[256]&~m[268]&m[269]&m[270]&~m[271])|(~m[256]&m[268]&~m[269]&~m[270]&m[271])|(~m[256]&~m[268]&m[269]&~m[270]&m[271])|(m[256]&m[268]&m[269]&~m[270]&m[271])|(~m[256]&m[268]&m[269]&m[270]&m[271]))&UnbiasedRNG[25])|((m[256]&~m[268]&~m[269]&m[270]&~m[271])|(~m[256]&~m[268]&~m[269]&~m[270]&m[271])|(m[256]&~m[268]&~m[269]&~m[270]&m[271])|(m[256]&m[268]&~m[269]&~m[270]&m[271])|(m[256]&~m[268]&m[269]&~m[270]&m[271])|(~m[256]&~m[268]&~m[269]&m[270]&m[271])|(m[256]&~m[268]&~m[269]&m[270]&m[271])|(~m[256]&m[268]&~m[269]&m[270]&m[271])|(m[256]&m[268]&~m[269]&m[270]&m[271])|(~m[256]&~m[268]&m[269]&m[270]&m[271])|(m[256]&~m[268]&m[269]&m[270]&m[271])|(m[256]&m[268]&m[269]&m[270]&m[271]))):InitCond[72];
    m[272] = run?((((m[270]&~m[273]&~m[274]&~m[275]&~m[276])|(~m[270]&~m[273]&~m[274]&m[275]&~m[276])|(m[270]&m[273]&~m[274]&m[275]&~m[276])|(m[270]&~m[273]&m[274]&m[275]&~m[276])|(~m[270]&m[273]&~m[274]&~m[275]&m[276])|(~m[270]&~m[273]&m[274]&~m[275]&m[276])|(m[270]&m[273]&m[274]&~m[275]&m[276])|(~m[270]&m[273]&m[274]&m[275]&m[276]))&UnbiasedRNG[26])|((m[270]&~m[273]&~m[274]&m[275]&~m[276])|(~m[270]&~m[273]&~m[274]&~m[275]&m[276])|(m[270]&~m[273]&~m[274]&~m[275]&m[276])|(m[270]&m[273]&~m[274]&~m[275]&m[276])|(m[270]&~m[273]&m[274]&~m[275]&m[276])|(~m[270]&~m[273]&~m[274]&m[275]&m[276])|(m[270]&~m[273]&~m[274]&m[275]&m[276])|(~m[270]&m[273]&~m[274]&m[275]&m[276])|(m[270]&m[273]&~m[274]&m[275]&m[276])|(~m[270]&~m[273]&m[274]&m[275]&m[276])|(m[270]&~m[273]&m[274]&m[275]&m[276])|(m[270]&m[273]&m[274]&m[275]&m[276]))):InitCond[73];
    m[277] = run?((((m[271]&~m[278]&~m[279]&~m[280]&~m[281])|(~m[271]&~m[278]&~m[279]&m[280]&~m[281])|(m[271]&m[278]&~m[279]&m[280]&~m[281])|(m[271]&~m[278]&m[279]&m[280]&~m[281])|(~m[271]&m[278]&~m[279]&~m[280]&m[281])|(~m[271]&~m[278]&m[279]&~m[280]&m[281])|(m[271]&m[278]&m[279]&~m[280]&m[281])|(~m[271]&m[278]&m[279]&m[280]&m[281]))&UnbiasedRNG[27])|((m[271]&~m[278]&~m[279]&m[280]&~m[281])|(~m[271]&~m[278]&~m[279]&~m[280]&m[281])|(m[271]&~m[278]&~m[279]&~m[280]&m[281])|(m[271]&m[278]&~m[279]&~m[280]&m[281])|(m[271]&~m[278]&m[279]&~m[280]&m[281])|(~m[271]&~m[278]&~m[279]&m[280]&m[281])|(m[271]&~m[278]&~m[279]&m[280]&m[281])|(~m[271]&m[278]&~m[279]&m[280]&m[281])|(m[271]&m[278]&~m[279]&m[280]&m[281])|(~m[271]&~m[278]&m[279]&m[280]&m[281])|(m[271]&~m[278]&m[279]&m[280]&m[281])|(m[271]&m[278]&m[279]&m[280]&m[281]))):InitCond[74];
end

always @(posedge color1_clk) begin
    m[12] = run?((((m[0]&m[26]&~m[27]&~m[28]&~m[29])|(m[0]&~m[26]&m[27]&~m[28]&~m[29])|(~m[0]&m[26]&m[27]&~m[28]&~m[29])|(m[0]&~m[26]&~m[27]&m[28]&~m[29])|(~m[0]&m[26]&~m[27]&m[28]&~m[29])|(~m[0]&~m[26]&m[27]&m[28]&~m[29])|(m[0]&~m[26]&~m[27]&~m[28]&m[29])|(~m[0]&m[26]&~m[27]&~m[28]&m[29])|(~m[0]&~m[26]&m[27]&~m[28]&m[29])|(~m[0]&~m[26]&~m[27]&m[28]&m[29]))&BiasedRNG[47])|(((m[0]&m[26]&m[27]&~m[28]&~m[29])|(m[0]&m[26]&~m[27]&m[28]&~m[29])|(m[0]&~m[26]&m[27]&m[28]&~m[29])|(~m[0]&m[26]&m[27]&m[28]&~m[29])|(m[0]&m[26]&~m[27]&~m[28]&m[29])|(m[0]&~m[26]&m[27]&~m[28]&m[29])|(~m[0]&m[26]&m[27]&~m[28]&m[29])|(m[0]&~m[26]&~m[27]&m[28]&m[29])|(~m[0]&m[26]&~m[27]&m[28]&m[29])|(~m[0]&~m[26]&m[27]&m[28]&m[29]))&~BiasedRNG[47])|((m[0]&m[26]&m[27]&m[28]&~m[29])|(m[0]&m[26]&m[27]&~m[28]&m[29])|(m[0]&m[26]&~m[27]&m[28]&m[29])|(m[0]&~m[26]&m[27]&m[28]&m[29])|(~m[0]&m[26]&m[27]&m[28]&m[29])|(m[0]&m[26]&m[27]&m[28]&m[29]))):InitCond[75];
    m[13] = run?((((m[1]&m[32]&~m[33]&~m[34]&~m[35])|(m[1]&~m[32]&m[33]&~m[34]&~m[35])|(~m[1]&m[32]&m[33]&~m[34]&~m[35])|(m[1]&~m[32]&~m[33]&m[34]&~m[35])|(~m[1]&m[32]&~m[33]&m[34]&~m[35])|(~m[1]&~m[32]&m[33]&m[34]&~m[35])|(m[1]&~m[32]&~m[33]&~m[34]&m[35])|(~m[1]&m[32]&~m[33]&~m[34]&m[35])|(~m[1]&~m[32]&m[33]&~m[34]&m[35])|(~m[1]&~m[32]&~m[33]&m[34]&m[35]))&BiasedRNG[48])|(((m[1]&m[32]&m[33]&~m[34]&~m[35])|(m[1]&m[32]&~m[33]&m[34]&~m[35])|(m[1]&~m[32]&m[33]&m[34]&~m[35])|(~m[1]&m[32]&m[33]&m[34]&~m[35])|(m[1]&m[32]&~m[33]&~m[34]&m[35])|(m[1]&~m[32]&m[33]&~m[34]&m[35])|(~m[1]&m[32]&m[33]&~m[34]&m[35])|(m[1]&~m[32]&~m[33]&m[34]&m[35])|(~m[1]&m[32]&~m[33]&m[34]&m[35])|(~m[1]&~m[32]&m[33]&m[34]&m[35]))&~BiasedRNG[48])|((m[1]&m[32]&m[33]&m[34]&~m[35])|(m[1]&m[32]&m[33]&~m[34]&m[35])|(m[1]&m[32]&~m[33]&m[34]&m[35])|(m[1]&~m[32]&m[33]&m[34]&m[35])|(~m[1]&m[32]&m[33]&m[34]&m[35])|(m[1]&m[32]&m[33]&m[34]&m[35]))):InitCond[76];
    m[14] = run?((((m[2]&m[38]&~m[39]&~m[40]&~m[41])|(m[2]&~m[38]&m[39]&~m[40]&~m[41])|(~m[2]&m[38]&m[39]&~m[40]&~m[41])|(m[2]&~m[38]&~m[39]&m[40]&~m[41])|(~m[2]&m[38]&~m[39]&m[40]&~m[41])|(~m[2]&~m[38]&m[39]&m[40]&~m[41])|(m[2]&~m[38]&~m[39]&~m[40]&m[41])|(~m[2]&m[38]&~m[39]&~m[40]&m[41])|(~m[2]&~m[38]&m[39]&~m[40]&m[41])|(~m[2]&~m[38]&~m[39]&m[40]&m[41]))&BiasedRNG[49])|(((m[2]&m[38]&m[39]&~m[40]&~m[41])|(m[2]&m[38]&~m[39]&m[40]&~m[41])|(m[2]&~m[38]&m[39]&m[40]&~m[41])|(~m[2]&m[38]&m[39]&m[40]&~m[41])|(m[2]&m[38]&~m[39]&~m[40]&m[41])|(m[2]&~m[38]&m[39]&~m[40]&m[41])|(~m[2]&m[38]&m[39]&~m[40]&m[41])|(m[2]&~m[38]&~m[39]&m[40]&m[41])|(~m[2]&m[38]&~m[39]&m[40]&m[41])|(~m[2]&~m[38]&m[39]&m[40]&m[41]))&~BiasedRNG[49])|((m[2]&m[38]&m[39]&m[40]&~m[41])|(m[2]&m[38]&m[39]&~m[40]&m[41])|(m[2]&m[38]&~m[39]&m[40]&m[41])|(m[2]&~m[38]&m[39]&m[40]&m[41])|(~m[2]&m[38]&m[39]&m[40]&m[41])|(m[2]&m[38]&m[39]&m[40]&m[41]))):InitCond[77];
    m[15] = run?((((m[3]&m[44]&~m[45]&~m[46]&~m[47])|(m[3]&~m[44]&m[45]&~m[46]&~m[47])|(~m[3]&m[44]&m[45]&~m[46]&~m[47])|(m[3]&~m[44]&~m[45]&m[46]&~m[47])|(~m[3]&m[44]&~m[45]&m[46]&~m[47])|(~m[3]&~m[44]&m[45]&m[46]&~m[47])|(m[3]&~m[44]&~m[45]&~m[46]&m[47])|(~m[3]&m[44]&~m[45]&~m[46]&m[47])|(~m[3]&~m[44]&m[45]&~m[46]&m[47])|(~m[3]&~m[44]&~m[45]&m[46]&m[47]))&BiasedRNG[50])|(((m[3]&m[44]&m[45]&~m[46]&~m[47])|(m[3]&m[44]&~m[45]&m[46]&~m[47])|(m[3]&~m[44]&m[45]&m[46]&~m[47])|(~m[3]&m[44]&m[45]&m[46]&~m[47])|(m[3]&m[44]&~m[45]&~m[46]&m[47])|(m[3]&~m[44]&m[45]&~m[46]&m[47])|(~m[3]&m[44]&m[45]&~m[46]&m[47])|(m[3]&~m[44]&~m[45]&m[46]&m[47])|(~m[3]&m[44]&~m[45]&m[46]&m[47])|(~m[3]&~m[44]&m[45]&m[46]&m[47]))&~BiasedRNG[50])|((m[3]&m[44]&m[45]&m[46]&~m[47])|(m[3]&m[44]&m[45]&~m[46]&m[47])|(m[3]&m[44]&~m[45]&m[46]&m[47])|(m[3]&~m[44]&m[45]&m[46]&m[47])|(~m[3]&m[44]&m[45]&m[46]&m[47])|(m[3]&m[44]&m[45]&m[46]&m[47]))):InitCond[78];
    m[16] = run?((((m[4]&m[50]&~m[51]&~m[52]&~m[53])|(m[4]&~m[50]&m[51]&~m[52]&~m[53])|(~m[4]&m[50]&m[51]&~m[52]&~m[53])|(m[4]&~m[50]&~m[51]&m[52]&~m[53])|(~m[4]&m[50]&~m[51]&m[52]&~m[53])|(~m[4]&~m[50]&m[51]&m[52]&~m[53])|(m[4]&~m[50]&~m[51]&~m[52]&m[53])|(~m[4]&m[50]&~m[51]&~m[52]&m[53])|(~m[4]&~m[50]&m[51]&~m[52]&m[53])|(~m[4]&~m[50]&~m[51]&m[52]&m[53]))&BiasedRNG[51])|(((m[4]&m[50]&m[51]&~m[52]&~m[53])|(m[4]&m[50]&~m[51]&m[52]&~m[53])|(m[4]&~m[50]&m[51]&m[52]&~m[53])|(~m[4]&m[50]&m[51]&m[52]&~m[53])|(m[4]&m[50]&~m[51]&~m[52]&m[53])|(m[4]&~m[50]&m[51]&~m[52]&m[53])|(~m[4]&m[50]&m[51]&~m[52]&m[53])|(m[4]&~m[50]&~m[51]&m[52]&m[53])|(~m[4]&m[50]&~m[51]&m[52]&m[53])|(~m[4]&~m[50]&m[51]&m[52]&m[53]))&~BiasedRNG[51])|((m[4]&m[50]&m[51]&m[52]&~m[53])|(m[4]&m[50]&m[51]&~m[52]&m[53])|(m[4]&m[50]&~m[51]&m[52]&m[53])|(m[4]&~m[50]&m[51]&m[52]&m[53])|(~m[4]&m[50]&m[51]&m[52]&m[53])|(m[4]&m[50]&m[51]&m[52]&m[53]))):InitCond[79];
    m[17] = run?((((m[5]&m[56]&~m[57]&~m[58]&~m[59])|(m[5]&~m[56]&m[57]&~m[58]&~m[59])|(~m[5]&m[56]&m[57]&~m[58]&~m[59])|(m[5]&~m[56]&~m[57]&m[58]&~m[59])|(~m[5]&m[56]&~m[57]&m[58]&~m[59])|(~m[5]&~m[56]&m[57]&m[58]&~m[59])|(m[5]&~m[56]&~m[57]&~m[58]&m[59])|(~m[5]&m[56]&~m[57]&~m[58]&m[59])|(~m[5]&~m[56]&m[57]&~m[58]&m[59])|(~m[5]&~m[56]&~m[57]&m[58]&m[59]))&BiasedRNG[52])|(((m[5]&m[56]&m[57]&~m[58]&~m[59])|(m[5]&m[56]&~m[57]&m[58]&~m[59])|(m[5]&~m[56]&m[57]&m[58]&~m[59])|(~m[5]&m[56]&m[57]&m[58]&~m[59])|(m[5]&m[56]&~m[57]&~m[58]&m[59])|(m[5]&~m[56]&m[57]&~m[58]&m[59])|(~m[5]&m[56]&m[57]&~m[58]&m[59])|(m[5]&~m[56]&~m[57]&m[58]&m[59])|(~m[5]&m[56]&~m[57]&m[58]&m[59])|(~m[5]&~m[56]&m[57]&m[58]&m[59]))&~BiasedRNG[52])|((m[5]&m[56]&m[57]&m[58]&~m[59])|(m[5]&m[56]&m[57]&~m[58]&m[59])|(m[5]&m[56]&~m[57]&m[58]&m[59])|(m[5]&~m[56]&m[57]&m[58]&m[59])|(~m[5]&m[56]&m[57]&m[58]&m[59])|(m[5]&m[56]&m[57]&m[58]&m[59]))):InitCond[80];
    m[18] = run?((((m[6]&m[62]&~m[63]&~m[64]&~m[65])|(m[6]&~m[62]&m[63]&~m[64]&~m[65])|(~m[6]&m[62]&m[63]&~m[64]&~m[65])|(m[6]&~m[62]&~m[63]&m[64]&~m[65])|(~m[6]&m[62]&~m[63]&m[64]&~m[65])|(~m[6]&~m[62]&m[63]&m[64]&~m[65])|(m[6]&~m[62]&~m[63]&~m[64]&m[65])|(~m[6]&m[62]&~m[63]&~m[64]&m[65])|(~m[6]&~m[62]&m[63]&~m[64]&m[65])|(~m[6]&~m[62]&~m[63]&m[64]&m[65]))&BiasedRNG[53])|(((m[6]&m[62]&m[63]&~m[64]&~m[65])|(m[6]&m[62]&~m[63]&m[64]&~m[65])|(m[6]&~m[62]&m[63]&m[64]&~m[65])|(~m[6]&m[62]&m[63]&m[64]&~m[65])|(m[6]&m[62]&~m[63]&~m[64]&m[65])|(m[6]&~m[62]&m[63]&~m[64]&m[65])|(~m[6]&m[62]&m[63]&~m[64]&m[65])|(m[6]&~m[62]&~m[63]&m[64]&m[65])|(~m[6]&m[62]&~m[63]&m[64]&m[65])|(~m[6]&~m[62]&m[63]&m[64]&m[65]))&~BiasedRNG[53])|((m[6]&m[62]&m[63]&m[64]&~m[65])|(m[6]&m[62]&m[63]&~m[64]&m[65])|(m[6]&m[62]&~m[63]&m[64]&m[65])|(m[6]&~m[62]&m[63]&m[64]&m[65])|(~m[6]&m[62]&m[63]&m[64]&m[65])|(m[6]&m[62]&m[63]&m[64]&m[65]))):InitCond[81];
    m[19] = run?((((m[7]&m[68]&~m[69]&~m[70]&~m[71])|(m[7]&~m[68]&m[69]&~m[70]&~m[71])|(~m[7]&m[68]&m[69]&~m[70]&~m[71])|(m[7]&~m[68]&~m[69]&m[70]&~m[71])|(~m[7]&m[68]&~m[69]&m[70]&~m[71])|(~m[7]&~m[68]&m[69]&m[70]&~m[71])|(m[7]&~m[68]&~m[69]&~m[70]&m[71])|(~m[7]&m[68]&~m[69]&~m[70]&m[71])|(~m[7]&~m[68]&m[69]&~m[70]&m[71])|(~m[7]&~m[68]&~m[69]&m[70]&m[71]))&BiasedRNG[54])|(((m[7]&m[68]&m[69]&~m[70]&~m[71])|(m[7]&m[68]&~m[69]&m[70]&~m[71])|(m[7]&~m[68]&m[69]&m[70]&~m[71])|(~m[7]&m[68]&m[69]&m[70]&~m[71])|(m[7]&m[68]&~m[69]&~m[70]&m[71])|(m[7]&~m[68]&m[69]&~m[70]&m[71])|(~m[7]&m[68]&m[69]&~m[70]&m[71])|(m[7]&~m[68]&~m[69]&m[70]&m[71])|(~m[7]&m[68]&~m[69]&m[70]&m[71])|(~m[7]&~m[68]&m[69]&m[70]&m[71]))&~BiasedRNG[54])|((m[7]&m[68]&m[69]&m[70]&~m[71])|(m[7]&m[68]&m[69]&~m[70]&m[71])|(m[7]&m[68]&~m[69]&m[70]&m[71])|(m[7]&~m[68]&m[69]&m[70]&m[71])|(~m[7]&m[68]&m[69]&m[70]&m[71])|(m[7]&m[68]&m[69]&m[70]&m[71]))):InitCond[82];
    m[20] = run?((((m[8]&m[74]&~m[75]&~m[76]&~m[77])|(m[8]&~m[74]&m[75]&~m[76]&~m[77])|(~m[8]&m[74]&m[75]&~m[76]&~m[77])|(m[8]&~m[74]&~m[75]&m[76]&~m[77])|(~m[8]&m[74]&~m[75]&m[76]&~m[77])|(~m[8]&~m[74]&m[75]&m[76]&~m[77])|(m[8]&~m[74]&~m[75]&~m[76]&m[77])|(~m[8]&m[74]&~m[75]&~m[76]&m[77])|(~m[8]&~m[74]&m[75]&~m[76]&m[77])|(~m[8]&~m[74]&~m[75]&m[76]&m[77]))&BiasedRNG[55])|(((m[8]&m[74]&m[75]&~m[76]&~m[77])|(m[8]&m[74]&~m[75]&m[76]&~m[77])|(m[8]&~m[74]&m[75]&m[76]&~m[77])|(~m[8]&m[74]&m[75]&m[76]&~m[77])|(m[8]&m[74]&~m[75]&~m[76]&m[77])|(m[8]&~m[74]&m[75]&~m[76]&m[77])|(~m[8]&m[74]&m[75]&~m[76]&m[77])|(m[8]&~m[74]&~m[75]&m[76]&m[77])|(~m[8]&m[74]&~m[75]&m[76]&m[77])|(~m[8]&~m[74]&m[75]&m[76]&m[77]))&~BiasedRNG[55])|((m[8]&m[74]&m[75]&m[76]&~m[77])|(m[8]&m[74]&m[75]&~m[76]&m[77])|(m[8]&m[74]&~m[75]&m[76]&m[77])|(m[8]&~m[74]&m[75]&m[76]&m[77])|(~m[8]&m[74]&m[75]&m[76]&m[77])|(m[8]&m[74]&m[75]&m[76]&m[77]))):InitCond[83];
    m[21] = run?((((m[9]&m[80]&~m[81]&~m[82]&~m[83])|(m[9]&~m[80]&m[81]&~m[82]&~m[83])|(~m[9]&m[80]&m[81]&~m[82]&~m[83])|(m[9]&~m[80]&~m[81]&m[82]&~m[83])|(~m[9]&m[80]&~m[81]&m[82]&~m[83])|(~m[9]&~m[80]&m[81]&m[82]&~m[83])|(m[9]&~m[80]&~m[81]&~m[82]&m[83])|(~m[9]&m[80]&~m[81]&~m[82]&m[83])|(~m[9]&~m[80]&m[81]&~m[82]&m[83])|(~m[9]&~m[80]&~m[81]&m[82]&m[83]))&BiasedRNG[56])|(((m[9]&m[80]&m[81]&~m[82]&~m[83])|(m[9]&m[80]&~m[81]&m[82]&~m[83])|(m[9]&~m[80]&m[81]&m[82]&~m[83])|(~m[9]&m[80]&m[81]&m[82]&~m[83])|(m[9]&m[80]&~m[81]&~m[82]&m[83])|(m[9]&~m[80]&m[81]&~m[82]&m[83])|(~m[9]&m[80]&m[81]&~m[82]&m[83])|(m[9]&~m[80]&~m[81]&m[82]&m[83])|(~m[9]&m[80]&~m[81]&m[82]&m[83])|(~m[9]&~m[80]&m[81]&m[82]&m[83]))&~BiasedRNG[56])|((m[9]&m[80]&m[81]&m[82]&~m[83])|(m[9]&m[80]&m[81]&~m[82]&m[83])|(m[9]&m[80]&~m[81]&m[82]&m[83])|(m[9]&~m[80]&m[81]&m[82]&m[83])|(~m[9]&m[80]&m[81]&m[82]&m[83])|(m[9]&m[80]&m[81]&m[82]&m[83]))):InitCond[84];
    m[22] = run?((((m[10]&m[86]&~m[87]&~m[88]&~m[89])|(m[10]&~m[86]&m[87]&~m[88]&~m[89])|(~m[10]&m[86]&m[87]&~m[88]&~m[89])|(m[10]&~m[86]&~m[87]&m[88]&~m[89])|(~m[10]&m[86]&~m[87]&m[88]&~m[89])|(~m[10]&~m[86]&m[87]&m[88]&~m[89])|(m[10]&~m[86]&~m[87]&~m[88]&m[89])|(~m[10]&m[86]&~m[87]&~m[88]&m[89])|(~m[10]&~m[86]&m[87]&~m[88]&m[89])|(~m[10]&~m[86]&~m[87]&m[88]&m[89]))&BiasedRNG[57])|(((m[10]&m[86]&m[87]&~m[88]&~m[89])|(m[10]&m[86]&~m[87]&m[88]&~m[89])|(m[10]&~m[86]&m[87]&m[88]&~m[89])|(~m[10]&m[86]&m[87]&m[88]&~m[89])|(m[10]&m[86]&~m[87]&~m[88]&m[89])|(m[10]&~m[86]&m[87]&~m[88]&m[89])|(~m[10]&m[86]&m[87]&~m[88]&m[89])|(m[10]&~m[86]&~m[87]&m[88]&m[89])|(~m[10]&m[86]&~m[87]&m[88]&m[89])|(~m[10]&~m[86]&m[87]&m[88]&m[89]))&~BiasedRNG[57])|((m[10]&m[86]&m[87]&m[88]&~m[89])|(m[10]&m[86]&m[87]&~m[88]&m[89])|(m[10]&m[86]&~m[87]&m[88]&m[89])|(m[10]&~m[86]&m[87]&m[88]&m[89])|(~m[10]&m[86]&m[87]&m[88]&m[89])|(m[10]&m[86]&m[87]&m[88]&m[89]))):InitCond[85];
    m[23] = run?((((m[11]&m[92]&~m[93]&~m[94]&~m[95])|(m[11]&~m[92]&m[93]&~m[94]&~m[95])|(~m[11]&m[92]&m[93]&~m[94]&~m[95])|(m[11]&~m[92]&~m[93]&m[94]&~m[95])|(~m[11]&m[92]&~m[93]&m[94]&~m[95])|(~m[11]&~m[92]&m[93]&m[94]&~m[95])|(m[11]&~m[92]&~m[93]&~m[94]&m[95])|(~m[11]&m[92]&~m[93]&~m[94]&m[95])|(~m[11]&~m[92]&m[93]&~m[94]&m[95])|(~m[11]&~m[92]&~m[93]&m[94]&m[95]))&BiasedRNG[58])|(((m[11]&m[92]&m[93]&~m[94]&~m[95])|(m[11]&m[92]&~m[93]&m[94]&~m[95])|(m[11]&~m[92]&m[93]&m[94]&~m[95])|(~m[11]&m[92]&m[93]&m[94]&~m[95])|(m[11]&m[92]&~m[93]&~m[94]&m[95])|(m[11]&~m[92]&m[93]&~m[94]&m[95])|(~m[11]&m[92]&m[93]&~m[94]&m[95])|(m[11]&~m[92]&~m[93]&m[94]&m[95])|(~m[11]&m[92]&~m[93]&m[94]&m[95])|(~m[11]&~m[92]&m[93]&m[94]&m[95]))&~BiasedRNG[58])|((m[11]&m[92]&m[93]&m[94]&~m[95])|(m[11]&m[92]&m[93]&~m[94]&m[95])|(m[11]&m[92]&~m[93]&m[94]&m[95])|(m[11]&~m[92]&m[93]&m[94]&m[95])|(~m[11]&m[92]&m[93]&m[94]&m[95])|(m[11]&m[92]&m[93]&m[94]&m[95]))):InitCond[86];
    m[24] = run?((((~m[0]&~m[60]&~m[96])|(m[0]&m[60]&~m[96]))&BiasedRNG[59])|(((m[0]&~m[60]&~m[96])|(~m[0]&m[60]&m[96]))&~BiasedRNG[59])|((~m[0]&~m[60]&m[96])|(m[0]&~m[60]&m[96])|(m[0]&m[60]&m[96]))):InitCond[87];
    m[25] = run?((((~m[0]&~m[66]&~m[102])|(m[0]&m[66]&~m[102]))&BiasedRNG[60])|(((m[0]&~m[66]&~m[102])|(~m[0]&m[66]&m[102]))&~BiasedRNG[60])|((~m[0]&~m[66]&m[102])|(m[0]&~m[66]&m[102])|(m[0]&m[66]&m[102]))):InitCond[88];
    m[30] = run?((((~m[1]&~m[61]&~m[97])|(m[1]&m[61]&~m[97]))&BiasedRNG[61])|(((m[1]&~m[61]&~m[97])|(~m[1]&m[61]&m[97]))&~BiasedRNG[61])|((~m[1]&~m[61]&m[97])|(m[1]&~m[61]&m[97])|(m[1]&m[61]&m[97]))):InitCond[89];
    m[31] = run?((((~m[1]&~m[67]&~m[103])|(m[1]&m[67]&~m[103]))&BiasedRNG[62])|(((m[1]&~m[67]&~m[103])|(~m[1]&m[67]&m[103]))&~BiasedRNG[62])|((~m[1]&~m[67]&m[103])|(m[1]&~m[67]&m[103])|(m[1]&m[67]&m[103]))):InitCond[90];
    m[36] = run?((((~m[2]&~m[62]&~m[98])|(m[2]&m[62]&~m[98]))&BiasedRNG[63])|(((m[2]&~m[62]&~m[98])|(~m[2]&m[62]&m[98]))&~BiasedRNG[63])|((~m[2]&~m[62]&m[98])|(m[2]&~m[62]&m[98])|(m[2]&m[62]&m[98]))):InitCond[91];
    m[37] = run?((((~m[2]&~m[68]&~m[104])|(m[2]&m[68]&~m[104]))&BiasedRNG[64])|(((m[2]&~m[68]&~m[104])|(~m[2]&m[68]&m[104]))&~BiasedRNG[64])|((~m[2]&~m[68]&m[104])|(m[2]&~m[68]&m[104])|(m[2]&m[68]&m[104]))):InitCond[92];
    m[42] = run?((((~m[3]&~m[63]&~m[99])|(m[3]&m[63]&~m[99]))&BiasedRNG[65])|(((m[3]&~m[63]&~m[99])|(~m[3]&m[63]&m[99]))&~BiasedRNG[65])|((~m[3]&~m[63]&m[99])|(m[3]&~m[63]&m[99])|(m[3]&m[63]&m[99]))):InitCond[93];
    m[43] = run?((((~m[3]&~m[69]&~m[105])|(m[3]&m[69]&~m[105]))&BiasedRNG[66])|(((m[3]&~m[69]&~m[105])|(~m[3]&m[69]&m[105]))&~BiasedRNG[66])|((~m[3]&~m[69]&m[105])|(m[3]&~m[69]&m[105])|(m[3]&m[69]&m[105]))):InitCond[94];
    m[48] = run?((((~m[4]&~m[64]&~m[100])|(m[4]&m[64]&~m[100]))&BiasedRNG[67])|(((m[4]&~m[64]&~m[100])|(~m[4]&m[64]&m[100]))&~BiasedRNG[67])|((~m[4]&~m[64]&m[100])|(m[4]&~m[64]&m[100])|(m[4]&m[64]&m[100]))):InitCond[95];
    m[49] = run?((((~m[4]&~m[70]&~m[106])|(m[4]&m[70]&~m[106]))&BiasedRNG[68])|(((m[4]&~m[70]&~m[106])|(~m[4]&m[70]&m[106]))&~BiasedRNG[68])|((~m[4]&~m[70]&m[106])|(m[4]&~m[70]&m[106])|(m[4]&m[70]&m[106]))):InitCond[96];
    m[54] = run?((((~m[5]&~m[65]&~m[101])|(m[5]&m[65]&~m[101]))&BiasedRNG[69])|(((m[5]&~m[65]&~m[101])|(~m[5]&m[65]&m[101]))&~BiasedRNG[69])|((~m[5]&~m[65]&m[101])|(m[5]&~m[65]&m[101])|(m[5]&m[65]&m[101]))):InitCond[97];
    m[55] = run?((((~m[5]&~m[71]&~m[107])|(m[5]&m[71]&~m[107]))&BiasedRNG[70])|(((m[5]&~m[71]&~m[107])|(~m[5]&m[71]&m[107]))&~BiasedRNG[70])|((~m[5]&~m[71]&m[107])|(m[5]&~m[71]&m[107])|(m[5]&m[71]&m[107]))):InitCond[98];
    m[72] = run?((((~m[8]&~m[26]&~m[108])|(m[8]&m[26]&~m[108]))&BiasedRNG[71])|(((m[8]&~m[26]&~m[108])|(~m[8]&m[26]&m[108]))&~BiasedRNG[71])|((~m[8]&~m[26]&m[108])|(m[8]&~m[26]&m[108])|(m[8]&m[26]&m[108]))):InitCond[99];
    m[73] = run?((((~m[8]&~m[32]&~m[109])|(m[8]&m[32]&~m[109]))&BiasedRNG[72])|(((m[8]&~m[32]&~m[109])|(~m[8]&m[32]&m[109]))&~BiasedRNG[72])|((~m[8]&~m[32]&m[109])|(m[8]&~m[32]&m[109])|(m[8]&m[32]&m[109]))):InitCond[100];
    m[78] = run?((((~m[9]&~m[27]&~m[114])|(m[9]&m[27]&~m[114]))&BiasedRNG[73])|(((m[9]&~m[27]&~m[114])|(~m[9]&m[27]&m[114]))&~BiasedRNG[73])|((~m[9]&~m[27]&m[114])|(m[9]&~m[27]&m[114])|(m[9]&m[27]&m[114]))):InitCond[101];
    m[79] = run?((((~m[9]&~m[33]&~m[115])|(m[9]&m[33]&~m[115]))&BiasedRNG[74])|(((m[9]&~m[33]&~m[115])|(~m[9]&m[33]&m[115]))&~BiasedRNG[74])|((~m[9]&~m[33]&m[115])|(m[9]&~m[33]&m[115])|(m[9]&m[33]&m[115]))):InitCond[102];
    m[84] = run?((((~m[10]&~m[28]&~m[120])|(m[10]&m[28]&~m[120]))&BiasedRNG[75])|(((m[10]&~m[28]&~m[120])|(~m[10]&m[28]&m[120]))&~BiasedRNG[75])|((~m[10]&~m[28]&m[120])|(m[10]&~m[28]&m[120])|(m[10]&m[28]&m[120]))):InitCond[103];
    m[85] = run?((((~m[10]&~m[34]&~m[121])|(m[10]&m[34]&~m[121]))&BiasedRNG[76])|(((m[10]&~m[34]&~m[121])|(~m[10]&m[34]&m[121]))&~BiasedRNG[76])|((~m[10]&~m[34]&m[121])|(m[10]&~m[34]&m[121])|(m[10]&m[34]&m[121]))):InitCond[104];
    m[90] = run?((((~m[11]&~m[29]&~m[126])|(m[11]&m[29]&~m[126]))&BiasedRNG[77])|(((m[11]&~m[29]&~m[126])|(~m[11]&m[29]&m[126]))&~BiasedRNG[77])|((~m[11]&~m[29]&m[126])|(m[11]&~m[29]&m[126])|(m[11]&m[29]&m[126]))):InitCond[105];
    m[91] = run?((((~m[11]&~m[35]&~m[127])|(m[11]&m[35]&~m[127]))&BiasedRNG[78])|(((m[11]&~m[35]&~m[127])|(~m[11]&m[35]&m[127]))&~BiasedRNG[78])|((~m[11]&~m[35]&m[127])|(m[11]&~m[35]&m[127])|(m[11]&m[35]&m[127]))):InitCond[106];
    m[110] = run?((((m[38]&~m[74]&m[168])|(~m[38]&m[74]&m[168]))&BiasedRNG[79])|(((m[38]&m[74]&~m[168]))&~BiasedRNG[79])|((m[38]&m[74]&m[168]))):InitCond[107];
    m[111] = run?((((m[44]&~m[75]&m[188])|(~m[44]&m[75]&m[188]))&BiasedRNG[80])|(((m[44]&m[75]&~m[188]))&~BiasedRNG[80])|((m[44]&m[75]&m[188]))):InitCond[108];
    m[112] = run?((((m[50]&~m[76]&m[213])|(~m[50]&m[76]&m[213]))&BiasedRNG[81])|(((m[50]&m[76]&~m[213]))&~BiasedRNG[81])|((m[50]&m[76]&m[213]))):InitCond[109];
    m[113] = run?((((m[56]&~m[77]&m[233])|(~m[56]&m[77]&m[233]))&BiasedRNG[82])|(((m[56]&m[77]&~m[233]))&~BiasedRNG[82])|((m[56]&m[77]&m[233]))):InitCond[110];
    m[116] = run?((((m[39]&~m[80]&m[193])|(~m[39]&m[80]&m[193]))&BiasedRNG[83])|(((m[39]&m[80]&~m[193]))&~BiasedRNG[83])|((m[39]&m[80]&m[193]))):InitCond[111];
    m[117] = run?((((m[45]&~m[81]&m[218])|(~m[45]&m[81]&m[218]))&BiasedRNG[84])|(((m[45]&m[81]&~m[218]))&~BiasedRNG[84])|((m[45]&m[81]&m[218]))):InitCond[112];
    m[118] = run?((((m[51]&~m[82]&m[238])|(~m[51]&m[82]&m[238]))&BiasedRNG[85])|(((m[51]&m[82]&~m[238]))&~BiasedRNG[85])|((m[51]&m[82]&m[238]))):InitCond[113];
    m[119] = run?((((m[57]&~m[83]&m[253])|(~m[57]&m[83]&m[253]))&BiasedRNG[86])|(((m[57]&m[83]&~m[253]))&~BiasedRNG[86])|((m[57]&m[83]&m[253]))):InitCond[114];
    m[122] = run?((((m[40]&~m[86]&m[223])|(~m[40]&m[86]&m[223]))&BiasedRNG[87])|(((m[40]&m[86]&~m[223]))&~BiasedRNG[87])|((m[40]&m[86]&m[223]))):InitCond[115];
    m[123] = run?((((m[46]&~m[87]&m[243])|(~m[46]&m[87]&m[243]))&BiasedRNG[88])|(((m[46]&m[87]&~m[243]))&~BiasedRNG[88])|((m[46]&m[87]&m[243]))):InitCond[116];
    m[124] = run?((((m[52]&~m[88]&m[258])|(~m[52]&m[88]&m[258]))&BiasedRNG[89])|(((m[52]&m[88]&~m[258]))&~BiasedRNG[89])|((m[52]&m[88]&m[258]))):InitCond[117];
    m[125] = run?((((m[58]&~m[89]&m[268])|(~m[58]&m[89]&m[268]))&BiasedRNG[90])|(((m[58]&m[89]&~m[268]))&~BiasedRNG[90])|((m[58]&m[89]&m[268]))):InitCond[118];
    m[128] = run?((((m[41]&~m[92]&m[248])|(~m[41]&m[92]&m[248]))&BiasedRNG[91])|(((m[41]&m[92]&~m[248]))&~BiasedRNG[91])|((m[41]&m[92]&m[248]))):InitCond[119];
    m[129] = run?((((m[47]&~m[93]&m[263])|(~m[47]&m[93]&m[263]))&BiasedRNG[92])|(((m[47]&m[93]&~m[263]))&~BiasedRNG[92])|((m[47]&m[93]&m[263]))):InitCond[120];
    m[130] = run?((((m[53]&~m[94]&m[273])|(~m[53]&m[94]&m[273]))&BiasedRNG[93])|(((m[53]&m[94]&~m[273]))&~BiasedRNG[93])|((m[53]&m[94]&m[273]))):InitCond[121];
    m[131] = run?((((m[59]&~m[95]&m[278])|(~m[59]&m[95]&m[278]))&BiasedRNG[94])|(((m[59]&m[95]&~m[278]))&~BiasedRNG[94])|((m[59]&m[95]&m[278]))):InitCond[122];
    m[132] = run?((((m[97]&~m[133]&~m[134]&~m[135]&~m[136])|(~m[97]&~m[133]&~m[134]&m[135]&~m[136])|(m[97]&m[133]&~m[134]&m[135]&~m[136])|(m[97]&~m[133]&m[134]&m[135]&~m[136])|(~m[97]&m[133]&~m[134]&~m[135]&m[136])|(~m[97]&~m[133]&m[134]&~m[135]&m[136])|(m[97]&m[133]&m[134]&~m[135]&m[136])|(~m[97]&m[133]&m[134]&m[135]&m[136]))&UnbiasedRNG[28])|((m[97]&~m[133]&~m[134]&m[135]&~m[136])|(~m[97]&~m[133]&~m[134]&~m[135]&m[136])|(m[97]&~m[133]&~m[134]&~m[135]&m[136])|(m[97]&m[133]&~m[134]&~m[135]&m[136])|(m[97]&~m[133]&m[134]&~m[135]&m[136])|(~m[97]&~m[133]&~m[134]&m[135]&m[136])|(m[97]&~m[133]&~m[134]&m[135]&m[136])|(~m[97]&m[133]&~m[134]&m[135]&m[136])|(m[97]&m[133]&~m[134]&m[135]&m[136])|(~m[97]&~m[133]&m[134]&m[135]&m[136])|(m[97]&~m[133]&m[134]&m[135]&m[136])|(m[97]&m[133]&m[134]&m[135]&m[136]))):InitCond[123];
    m[138] = run?((((m[103]&~m[137]&~m[139]&~m[140]&~m[141])|(~m[103]&~m[137]&~m[139]&m[140]&~m[141])|(m[103]&m[137]&~m[139]&m[140]&~m[141])|(m[103]&~m[137]&m[139]&m[140]&~m[141])|(~m[103]&m[137]&~m[139]&~m[140]&m[141])|(~m[103]&~m[137]&m[139]&~m[140]&m[141])|(m[103]&m[137]&m[139]&~m[140]&m[141])|(~m[103]&m[137]&m[139]&m[140]&m[141]))&UnbiasedRNG[29])|((m[103]&~m[137]&~m[139]&m[140]&~m[141])|(~m[103]&~m[137]&~m[139]&~m[140]&m[141])|(m[103]&~m[137]&~m[139]&~m[140]&m[141])|(m[103]&m[137]&~m[139]&~m[140]&m[141])|(m[103]&~m[137]&m[139]&~m[140]&m[141])|(~m[103]&~m[137]&~m[139]&m[140]&m[141])|(m[103]&~m[137]&~m[139]&m[140]&m[141])|(~m[103]&m[137]&~m[139]&m[140]&m[141])|(m[103]&m[137]&~m[139]&m[140]&m[141])|(~m[103]&~m[137]&m[139]&m[140]&m[141])|(m[103]&~m[137]&m[139]&m[140]&m[141])|(m[103]&m[137]&m[139]&m[140]&m[141]))):InitCond[124];
    m[143] = run?((((m[108]&~m[142]&~m[144]&~m[145]&~m[146])|(~m[108]&~m[142]&~m[144]&m[145]&~m[146])|(m[108]&m[142]&~m[144]&m[145]&~m[146])|(m[108]&~m[142]&m[144]&m[145]&~m[146])|(~m[108]&m[142]&~m[144]&~m[145]&m[146])|(~m[108]&~m[142]&m[144]&~m[145]&m[146])|(m[108]&m[142]&m[144]&~m[145]&m[146])|(~m[108]&m[142]&m[144]&m[145]&m[146]))&UnbiasedRNG[30])|((m[108]&~m[142]&~m[144]&m[145]&~m[146])|(~m[108]&~m[142]&~m[144]&~m[145]&m[146])|(m[108]&~m[142]&~m[144]&~m[145]&m[146])|(m[108]&m[142]&~m[144]&~m[145]&m[146])|(m[108]&~m[142]&m[144]&~m[145]&m[146])|(~m[108]&~m[142]&~m[144]&m[145]&m[146])|(m[108]&~m[142]&~m[144]&m[145]&m[146])|(~m[108]&m[142]&~m[144]&m[145]&m[146])|(m[108]&m[142]&~m[144]&m[145]&m[146])|(~m[108]&~m[142]&m[144]&m[145]&m[146])|(m[108]&~m[142]&m[144]&m[145]&m[146])|(m[108]&m[142]&m[144]&m[145]&m[146]))):InitCond[125];
    m[148] = run?((((m[104]&~m[147]&~m[149]&~m[150]&~m[151])|(~m[104]&~m[147]&~m[149]&m[150]&~m[151])|(m[104]&m[147]&~m[149]&m[150]&~m[151])|(m[104]&~m[147]&m[149]&m[150]&~m[151])|(~m[104]&m[147]&~m[149]&~m[150]&m[151])|(~m[104]&~m[147]&m[149]&~m[150]&m[151])|(m[104]&m[147]&m[149]&~m[150]&m[151])|(~m[104]&m[147]&m[149]&m[150]&m[151]))&UnbiasedRNG[31])|((m[104]&~m[147]&~m[149]&m[150]&~m[151])|(~m[104]&~m[147]&~m[149]&~m[150]&m[151])|(m[104]&~m[147]&~m[149]&~m[150]&m[151])|(m[104]&m[147]&~m[149]&~m[150]&m[151])|(m[104]&~m[147]&m[149]&~m[150]&m[151])|(~m[104]&~m[147]&~m[149]&m[150]&m[151])|(m[104]&~m[147]&~m[149]&m[150]&m[151])|(~m[104]&m[147]&~m[149]&m[150]&m[151])|(m[104]&m[147]&~m[149]&m[150]&m[151])|(~m[104]&~m[147]&m[149]&m[150]&m[151])|(m[104]&~m[147]&m[149]&m[150]&m[151])|(m[104]&m[147]&m[149]&m[150]&m[151]))):InitCond[126];
    m[153] = run?((((m[109]&~m[152]&~m[154]&~m[155]&~m[156])|(~m[109]&~m[152]&~m[154]&m[155]&~m[156])|(m[109]&m[152]&~m[154]&m[155]&~m[156])|(m[109]&~m[152]&m[154]&m[155]&~m[156])|(~m[109]&m[152]&~m[154]&~m[155]&m[156])|(~m[109]&~m[152]&m[154]&~m[155]&m[156])|(m[109]&m[152]&m[154]&~m[155]&m[156])|(~m[109]&m[152]&m[154]&m[155]&m[156]))&UnbiasedRNG[32])|((m[109]&~m[152]&~m[154]&m[155]&~m[156])|(~m[109]&~m[152]&~m[154]&~m[155]&m[156])|(m[109]&~m[152]&~m[154]&~m[155]&m[156])|(m[109]&m[152]&~m[154]&~m[155]&m[156])|(m[109]&~m[152]&m[154]&~m[155]&m[156])|(~m[109]&~m[152]&~m[154]&m[155]&m[156])|(m[109]&~m[152]&~m[154]&m[155]&m[156])|(~m[109]&m[152]&~m[154]&m[155]&m[156])|(m[109]&m[152]&~m[154]&m[155]&m[156])|(~m[109]&~m[152]&m[154]&m[155]&m[156])|(m[109]&~m[152]&m[154]&m[155]&m[156])|(m[109]&m[152]&m[154]&m[155]&m[156]))):InitCond[127];
    m[158] = run?((((m[114]&~m[157]&~m[159]&~m[160]&~m[161])|(~m[114]&~m[157]&~m[159]&m[160]&~m[161])|(m[114]&m[157]&~m[159]&m[160]&~m[161])|(m[114]&~m[157]&m[159]&m[160]&~m[161])|(~m[114]&m[157]&~m[159]&~m[160]&m[161])|(~m[114]&~m[157]&m[159]&~m[160]&m[161])|(m[114]&m[157]&m[159]&~m[160]&m[161])|(~m[114]&m[157]&m[159]&m[160]&m[161]))&UnbiasedRNG[33])|((m[114]&~m[157]&~m[159]&m[160]&~m[161])|(~m[114]&~m[157]&~m[159]&~m[160]&m[161])|(m[114]&~m[157]&~m[159]&~m[160]&m[161])|(m[114]&m[157]&~m[159]&~m[160]&m[161])|(m[114]&~m[157]&m[159]&~m[160]&m[161])|(~m[114]&~m[157]&~m[159]&m[160]&m[161])|(m[114]&~m[157]&~m[159]&m[160]&m[161])|(~m[114]&m[157]&~m[159]&m[160]&m[161])|(m[114]&m[157]&~m[159]&m[160]&m[161])|(~m[114]&~m[157]&m[159]&m[160]&m[161])|(m[114]&~m[157]&m[159]&m[160]&m[161])|(m[114]&m[157]&m[159]&m[160]&m[161]))):InitCond[128];
    m[163] = run?((((m[105]&~m[162]&~m[164]&~m[165]&~m[166])|(~m[105]&~m[162]&~m[164]&m[165]&~m[166])|(m[105]&m[162]&~m[164]&m[165]&~m[166])|(m[105]&~m[162]&m[164]&m[165]&~m[166])|(~m[105]&m[162]&~m[164]&~m[165]&m[166])|(~m[105]&~m[162]&m[164]&~m[165]&m[166])|(m[105]&m[162]&m[164]&~m[165]&m[166])|(~m[105]&m[162]&m[164]&m[165]&m[166]))&UnbiasedRNG[34])|((m[105]&~m[162]&~m[164]&m[165]&~m[166])|(~m[105]&~m[162]&~m[164]&~m[165]&m[166])|(m[105]&~m[162]&~m[164]&~m[165]&m[166])|(m[105]&m[162]&~m[164]&~m[165]&m[166])|(m[105]&~m[162]&m[164]&~m[165]&m[166])|(~m[105]&~m[162]&~m[164]&m[165]&m[166])|(m[105]&~m[162]&~m[164]&m[165]&m[166])|(~m[105]&m[162]&~m[164]&m[165]&m[166])|(m[105]&m[162]&~m[164]&m[165]&m[166])|(~m[105]&~m[162]&m[164]&m[165]&m[166])|(m[105]&~m[162]&m[164]&m[165]&m[166])|(m[105]&m[162]&m[164]&m[165]&m[166]))):InitCond[129];
    m[169] = run?((((m[156]&~m[167]&~m[168]&~m[170]&~m[171])|(~m[156]&~m[167]&~m[168]&m[170]&~m[171])|(m[156]&m[167]&~m[168]&m[170]&~m[171])|(m[156]&~m[167]&m[168]&m[170]&~m[171])|(~m[156]&m[167]&~m[168]&~m[170]&m[171])|(~m[156]&~m[167]&m[168]&~m[170]&m[171])|(m[156]&m[167]&m[168]&~m[170]&m[171])|(~m[156]&m[167]&m[168]&m[170]&m[171]))&UnbiasedRNG[35])|((m[156]&~m[167]&~m[168]&m[170]&~m[171])|(~m[156]&~m[167]&~m[168]&~m[170]&m[171])|(m[156]&~m[167]&~m[168]&~m[170]&m[171])|(m[156]&m[167]&~m[168]&~m[170]&m[171])|(m[156]&~m[167]&m[168]&~m[170]&m[171])|(~m[156]&~m[167]&~m[168]&m[170]&m[171])|(m[156]&~m[167]&~m[168]&m[170]&m[171])|(~m[156]&m[167]&~m[168]&m[170]&m[171])|(m[156]&m[167]&~m[168]&m[170]&m[171])|(~m[156]&~m[167]&m[168]&m[170]&m[171])|(m[156]&~m[167]&m[168]&m[170]&m[171])|(m[156]&m[167]&m[168]&m[170]&m[171]))):InitCond[130];
    m[173] = run?((((m[115]&~m[172]&~m[174]&~m[175]&~m[176])|(~m[115]&~m[172]&~m[174]&m[175]&~m[176])|(m[115]&m[172]&~m[174]&m[175]&~m[176])|(m[115]&~m[172]&m[174]&m[175]&~m[176])|(~m[115]&m[172]&~m[174]&~m[175]&m[176])|(~m[115]&~m[172]&m[174]&~m[175]&m[176])|(m[115]&m[172]&m[174]&~m[175]&m[176])|(~m[115]&m[172]&m[174]&m[175]&m[176]))&UnbiasedRNG[36])|((m[115]&~m[172]&~m[174]&m[175]&~m[176])|(~m[115]&~m[172]&~m[174]&~m[175]&m[176])|(m[115]&~m[172]&~m[174]&~m[175]&m[176])|(m[115]&m[172]&~m[174]&~m[175]&m[176])|(m[115]&~m[172]&m[174]&~m[175]&m[176])|(~m[115]&~m[172]&~m[174]&m[175]&m[176])|(m[115]&~m[172]&~m[174]&m[175]&m[176])|(~m[115]&m[172]&~m[174]&m[175]&m[176])|(m[115]&m[172]&~m[174]&m[175]&m[176])|(~m[115]&~m[172]&m[174]&m[175]&m[176])|(m[115]&~m[172]&m[174]&m[175]&m[176])|(m[115]&m[172]&m[174]&m[175]&m[176]))):InitCond[131];
    m[178] = run?((((m[120]&~m[177]&~m[179]&~m[180]&~m[181])|(~m[120]&~m[177]&~m[179]&m[180]&~m[181])|(m[120]&m[177]&~m[179]&m[180]&~m[181])|(m[120]&~m[177]&m[179]&m[180]&~m[181])|(~m[120]&m[177]&~m[179]&~m[180]&m[181])|(~m[120]&~m[177]&m[179]&~m[180]&m[181])|(m[120]&m[177]&m[179]&~m[180]&m[181])|(~m[120]&m[177]&m[179]&m[180]&m[181]))&UnbiasedRNG[37])|((m[120]&~m[177]&~m[179]&m[180]&~m[181])|(~m[120]&~m[177]&~m[179]&~m[180]&m[181])|(m[120]&~m[177]&~m[179]&~m[180]&m[181])|(m[120]&m[177]&~m[179]&~m[180]&m[181])|(m[120]&~m[177]&m[179]&~m[180]&m[181])|(~m[120]&~m[177]&~m[179]&m[180]&m[181])|(m[120]&~m[177]&~m[179]&m[180]&m[181])|(~m[120]&m[177]&~m[179]&m[180]&m[181])|(m[120]&m[177]&~m[179]&m[180]&m[181])|(~m[120]&~m[177]&m[179]&m[180]&m[181])|(m[120]&~m[177]&m[179]&m[180]&m[181])|(m[120]&m[177]&m[179]&m[180]&m[181]))):InitCond[132];
    m[183] = run?((((m[106]&~m[182]&~m[184]&~m[185]&~m[186])|(~m[106]&~m[182]&~m[184]&m[185]&~m[186])|(m[106]&m[182]&~m[184]&m[185]&~m[186])|(m[106]&~m[182]&m[184]&m[185]&~m[186])|(~m[106]&m[182]&~m[184]&~m[185]&m[186])|(~m[106]&~m[182]&m[184]&~m[185]&m[186])|(m[106]&m[182]&m[184]&~m[185]&m[186])|(~m[106]&m[182]&m[184]&m[185]&m[186]))&UnbiasedRNG[38])|((m[106]&~m[182]&~m[184]&m[185]&~m[186])|(~m[106]&~m[182]&~m[184]&~m[185]&m[186])|(m[106]&~m[182]&~m[184]&~m[185]&m[186])|(m[106]&m[182]&~m[184]&~m[185]&m[186])|(m[106]&~m[182]&m[184]&~m[185]&m[186])|(~m[106]&~m[182]&~m[184]&m[185]&m[186])|(m[106]&~m[182]&~m[184]&m[185]&m[186])|(~m[106]&m[182]&~m[184]&m[185]&m[186])|(m[106]&m[182]&~m[184]&m[185]&m[186])|(~m[106]&~m[182]&m[184]&m[185]&m[186])|(m[106]&~m[182]&m[184]&m[185]&m[186])|(m[106]&m[182]&m[184]&m[185]&m[186]))):InitCond[133];
    m[189] = run?((((m[171]&~m[187]&~m[188]&~m[190]&~m[191])|(~m[171]&~m[187]&~m[188]&m[190]&~m[191])|(m[171]&m[187]&~m[188]&m[190]&~m[191])|(m[171]&~m[187]&m[188]&m[190]&~m[191])|(~m[171]&m[187]&~m[188]&~m[190]&m[191])|(~m[171]&~m[187]&m[188]&~m[190]&m[191])|(m[171]&m[187]&m[188]&~m[190]&m[191])|(~m[171]&m[187]&m[188]&m[190]&m[191]))&UnbiasedRNG[39])|((m[171]&~m[187]&~m[188]&m[190]&~m[191])|(~m[171]&~m[187]&~m[188]&~m[190]&m[191])|(m[171]&~m[187]&~m[188]&~m[190]&m[191])|(m[171]&m[187]&~m[188]&~m[190]&m[191])|(m[171]&~m[187]&m[188]&~m[190]&m[191])|(~m[171]&~m[187]&~m[188]&m[190]&m[191])|(m[171]&~m[187]&~m[188]&m[190]&m[191])|(~m[171]&m[187]&~m[188]&m[190]&m[191])|(m[171]&m[187]&~m[188]&m[190]&m[191])|(~m[171]&~m[187]&m[188]&m[190]&m[191])|(m[171]&~m[187]&m[188]&m[190]&m[191])|(m[171]&m[187]&m[188]&m[190]&m[191]))):InitCond[134];
    m[194] = run?((((m[176]&~m[192]&~m[193]&~m[195]&~m[196])|(~m[176]&~m[192]&~m[193]&m[195]&~m[196])|(m[176]&m[192]&~m[193]&m[195]&~m[196])|(m[176]&~m[192]&m[193]&m[195]&~m[196])|(~m[176]&m[192]&~m[193]&~m[195]&m[196])|(~m[176]&~m[192]&m[193]&~m[195]&m[196])|(m[176]&m[192]&m[193]&~m[195]&m[196])|(~m[176]&m[192]&m[193]&m[195]&m[196]))&UnbiasedRNG[40])|((m[176]&~m[192]&~m[193]&m[195]&~m[196])|(~m[176]&~m[192]&~m[193]&~m[195]&m[196])|(m[176]&~m[192]&~m[193]&~m[195]&m[196])|(m[176]&m[192]&~m[193]&~m[195]&m[196])|(m[176]&~m[192]&m[193]&~m[195]&m[196])|(~m[176]&~m[192]&~m[193]&m[195]&m[196])|(m[176]&~m[192]&~m[193]&m[195]&m[196])|(~m[176]&m[192]&~m[193]&m[195]&m[196])|(m[176]&m[192]&~m[193]&m[195]&m[196])|(~m[176]&~m[192]&m[193]&m[195]&m[196])|(m[176]&~m[192]&m[193]&m[195]&m[196])|(m[176]&m[192]&m[193]&m[195]&m[196]))):InitCond[135];
    m[198] = run?((((m[121]&~m[197]&~m[199]&~m[200]&~m[201])|(~m[121]&~m[197]&~m[199]&m[200]&~m[201])|(m[121]&m[197]&~m[199]&m[200]&~m[201])|(m[121]&~m[197]&m[199]&m[200]&~m[201])|(~m[121]&m[197]&~m[199]&~m[200]&m[201])|(~m[121]&~m[197]&m[199]&~m[200]&m[201])|(m[121]&m[197]&m[199]&~m[200]&m[201])|(~m[121]&m[197]&m[199]&m[200]&m[201]))&UnbiasedRNG[41])|((m[121]&~m[197]&~m[199]&m[200]&~m[201])|(~m[121]&~m[197]&~m[199]&~m[200]&m[201])|(m[121]&~m[197]&~m[199]&~m[200]&m[201])|(m[121]&m[197]&~m[199]&~m[200]&m[201])|(m[121]&~m[197]&m[199]&~m[200]&m[201])|(~m[121]&~m[197]&~m[199]&m[200]&m[201])|(m[121]&~m[197]&~m[199]&m[200]&m[201])|(~m[121]&m[197]&~m[199]&m[200]&m[201])|(m[121]&m[197]&~m[199]&m[200]&m[201])|(~m[121]&~m[197]&m[199]&m[200]&m[201])|(m[121]&~m[197]&m[199]&m[200]&m[201])|(m[121]&m[197]&m[199]&m[200]&m[201]))):InitCond[136];
    m[203] = run?((((m[126]&~m[202]&~m[204]&~m[205]&~m[206])|(~m[126]&~m[202]&~m[204]&m[205]&~m[206])|(m[126]&m[202]&~m[204]&m[205]&~m[206])|(m[126]&~m[202]&m[204]&m[205]&~m[206])|(~m[126]&m[202]&~m[204]&~m[205]&m[206])|(~m[126]&~m[202]&m[204]&~m[205]&m[206])|(m[126]&m[202]&m[204]&~m[205]&m[206])|(~m[126]&m[202]&m[204]&m[205]&m[206]))&UnbiasedRNG[42])|((m[126]&~m[202]&~m[204]&m[205]&~m[206])|(~m[126]&~m[202]&~m[204]&~m[205]&m[206])|(m[126]&~m[202]&~m[204]&~m[205]&m[206])|(m[126]&m[202]&~m[204]&~m[205]&m[206])|(m[126]&~m[202]&m[204]&~m[205]&m[206])|(~m[126]&~m[202]&~m[204]&m[205]&m[206])|(m[126]&~m[202]&~m[204]&m[205]&m[206])|(~m[126]&m[202]&~m[204]&m[205]&m[206])|(m[126]&m[202]&~m[204]&m[205]&m[206])|(~m[126]&~m[202]&m[204]&m[205]&m[206])|(m[126]&~m[202]&m[204]&m[205]&m[206])|(m[126]&m[202]&m[204]&m[205]&m[206]))):InitCond[137];
    m[208] = run?((((m[107]&~m[207]&~m[209]&~m[210]&~m[211])|(~m[107]&~m[207]&~m[209]&m[210]&~m[211])|(m[107]&m[207]&~m[209]&m[210]&~m[211])|(m[107]&~m[207]&m[209]&m[210]&~m[211])|(~m[107]&m[207]&~m[209]&~m[210]&m[211])|(~m[107]&~m[207]&m[209]&~m[210]&m[211])|(m[107]&m[207]&m[209]&~m[210]&m[211])|(~m[107]&m[207]&m[209]&m[210]&m[211]))&UnbiasedRNG[43])|((m[107]&~m[207]&~m[209]&m[210]&~m[211])|(~m[107]&~m[207]&~m[209]&~m[210]&m[211])|(m[107]&~m[207]&~m[209]&~m[210]&m[211])|(m[107]&m[207]&~m[209]&~m[210]&m[211])|(m[107]&~m[207]&m[209]&~m[210]&m[211])|(~m[107]&~m[207]&~m[209]&m[210]&m[211])|(m[107]&~m[207]&~m[209]&m[210]&m[211])|(~m[107]&m[207]&~m[209]&m[210]&m[211])|(m[107]&m[207]&~m[209]&m[210]&m[211])|(~m[107]&~m[207]&m[209]&m[210]&m[211])|(m[107]&~m[207]&m[209]&m[210]&m[211])|(m[107]&m[207]&m[209]&m[210]&m[211]))):InitCond[138];
    m[214] = run?((((m[191]&~m[212]&~m[213]&~m[215]&~m[216])|(~m[191]&~m[212]&~m[213]&m[215]&~m[216])|(m[191]&m[212]&~m[213]&m[215]&~m[216])|(m[191]&~m[212]&m[213]&m[215]&~m[216])|(~m[191]&m[212]&~m[213]&~m[215]&m[216])|(~m[191]&~m[212]&m[213]&~m[215]&m[216])|(m[191]&m[212]&m[213]&~m[215]&m[216])|(~m[191]&m[212]&m[213]&m[215]&m[216]))&UnbiasedRNG[44])|((m[191]&~m[212]&~m[213]&m[215]&~m[216])|(~m[191]&~m[212]&~m[213]&~m[215]&m[216])|(m[191]&~m[212]&~m[213]&~m[215]&m[216])|(m[191]&m[212]&~m[213]&~m[215]&m[216])|(m[191]&~m[212]&m[213]&~m[215]&m[216])|(~m[191]&~m[212]&~m[213]&m[215]&m[216])|(m[191]&~m[212]&~m[213]&m[215]&m[216])|(~m[191]&m[212]&~m[213]&m[215]&m[216])|(m[191]&m[212]&~m[213]&m[215]&m[216])|(~m[191]&~m[212]&m[213]&m[215]&m[216])|(m[191]&~m[212]&m[213]&m[215]&m[216])|(m[191]&m[212]&m[213]&m[215]&m[216]))):InitCond[139];
    m[219] = run?((((m[196]&~m[217]&~m[218]&~m[220]&~m[221])|(~m[196]&~m[217]&~m[218]&m[220]&~m[221])|(m[196]&m[217]&~m[218]&m[220]&~m[221])|(m[196]&~m[217]&m[218]&m[220]&~m[221])|(~m[196]&m[217]&~m[218]&~m[220]&m[221])|(~m[196]&~m[217]&m[218]&~m[220]&m[221])|(m[196]&m[217]&m[218]&~m[220]&m[221])|(~m[196]&m[217]&m[218]&m[220]&m[221]))&UnbiasedRNG[45])|((m[196]&~m[217]&~m[218]&m[220]&~m[221])|(~m[196]&~m[217]&~m[218]&~m[220]&m[221])|(m[196]&~m[217]&~m[218]&~m[220]&m[221])|(m[196]&m[217]&~m[218]&~m[220]&m[221])|(m[196]&~m[217]&m[218]&~m[220]&m[221])|(~m[196]&~m[217]&~m[218]&m[220]&m[221])|(m[196]&~m[217]&~m[218]&m[220]&m[221])|(~m[196]&m[217]&~m[218]&m[220]&m[221])|(m[196]&m[217]&~m[218]&m[220]&m[221])|(~m[196]&~m[217]&m[218]&m[220]&m[221])|(m[196]&~m[217]&m[218]&m[220]&m[221])|(m[196]&m[217]&m[218]&m[220]&m[221]))):InitCond[140];
    m[224] = run?((((m[201]&~m[222]&~m[223]&~m[225]&~m[226])|(~m[201]&~m[222]&~m[223]&m[225]&~m[226])|(m[201]&m[222]&~m[223]&m[225]&~m[226])|(m[201]&~m[222]&m[223]&m[225]&~m[226])|(~m[201]&m[222]&~m[223]&~m[225]&m[226])|(~m[201]&~m[222]&m[223]&~m[225]&m[226])|(m[201]&m[222]&m[223]&~m[225]&m[226])|(~m[201]&m[222]&m[223]&m[225]&m[226]))&UnbiasedRNG[46])|((m[201]&~m[222]&~m[223]&m[225]&~m[226])|(~m[201]&~m[222]&~m[223]&~m[225]&m[226])|(m[201]&~m[222]&~m[223]&~m[225]&m[226])|(m[201]&m[222]&~m[223]&~m[225]&m[226])|(m[201]&~m[222]&m[223]&~m[225]&m[226])|(~m[201]&~m[222]&~m[223]&m[225]&m[226])|(m[201]&~m[222]&~m[223]&m[225]&m[226])|(~m[201]&m[222]&~m[223]&m[225]&m[226])|(m[201]&m[222]&~m[223]&m[225]&m[226])|(~m[201]&~m[222]&m[223]&m[225]&m[226])|(m[201]&~m[222]&m[223]&m[225]&m[226])|(m[201]&m[222]&m[223]&m[225]&m[226]))):InitCond[141];
    m[228] = run?((((m[127]&~m[227]&~m[229]&~m[230]&~m[231])|(~m[127]&~m[227]&~m[229]&m[230]&~m[231])|(m[127]&m[227]&~m[229]&m[230]&~m[231])|(m[127]&~m[227]&m[229]&m[230]&~m[231])|(~m[127]&m[227]&~m[229]&~m[230]&m[231])|(~m[127]&~m[227]&m[229]&~m[230]&m[231])|(m[127]&m[227]&m[229]&~m[230]&m[231])|(~m[127]&m[227]&m[229]&m[230]&m[231]))&UnbiasedRNG[47])|((m[127]&~m[227]&~m[229]&m[230]&~m[231])|(~m[127]&~m[227]&~m[229]&~m[230]&m[231])|(m[127]&~m[227]&~m[229]&~m[230]&m[231])|(m[127]&m[227]&~m[229]&~m[230]&m[231])|(m[127]&~m[227]&m[229]&~m[230]&m[231])|(~m[127]&~m[227]&~m[229]&m[230]&m[231])|(m[127]&~m[227]&~m[229]&m[230]&m[231])|(~m[127]&m[227]&~m[229]&m[230]&m[231])|(m[127]&m[227]&~m[229]&m[230]&m[231])|(~m[127]&~m[227]&m[229]&m[230]&m[231])|(m[127]&~m[227]&m[229]&m[230]&m[231])|(m[127]&m[227]&m[229]&m[230]&m[231]))):InitCond[142];
    m[234] = run?((((m[216]&~m[232]&~m[233]&~m[235]&~m[236])|(~m[216]&~m[232]&~m[233]&m[235]&~m[236])|(m[216]&m[232]&~m[233]&m[235]&~m[236])|(m[216]&~m[232]&m[233]&m[235]&~m[236])|(~m[216]&m[232]&~m[233]&~m[235]&m[236])|(~m[216]&~m[232]&m[233]&~m[235]&m[236])|(m[216]&m[232]&m[233]&~m[235]&m[236])|(~m[216]&m[232]&m[233]&m[235]&m[236]))&UnbiasedRNG[48])|((m[216]&~m[232]&~m[233]&m[235]&~m[236])|(~m[216]&~m[232]&~m[233]&~m[235]&m[236])|(m[216]&~m[232]&~m[233]&~m[235]&m[236])|(m[216]&m[232]&~m[233]&~m[235]&m[236])|(m[216]&~m[232]&m[233]&~m[235]&m[236])|(~m[216]&~m[232]&~m[233]&m[235]&m[236])|(m[216]&~m[232]&~m[233]&m[235]&m[236])|(~m[216]&m[232]&~m[233]&m[235]&m[236])|(m[216]&m[232]&~m[233]&m[235]&m[236])|(~m[216]&~m[232]&m[233]&m[235]&m[236])|(m[216]&~m[232]&m[233]&m[235]&m[236])|(m[216]&m[232]&m[233]&m[235]&m[236]))):InitCond[143];
    m[239] = run?((((m[221]&~m[237]&~m[238]&~m[240]&~m[241])|(~m[221]&~m[237]&~m[238]&m[240]&~m[241])|(m[221]&m[237]&~m[238]&m[240]&~m[241])|(m[221]&~m[237]&m[238]&m[240]&~m[241])|(~m[221]&m[237]&~m[238]&~m[240]&m[241])|(~m[221]&~m[237]&m[238]&~m[240]&m[241])|(m[221]&m[237]&m[238]&~m[240]&m[241])|(~m[221]&m[237]&m[238]&m[240]&m[241]))&UnbiasedRNG[49])|((m[221]&~m[237]&~m[238]&m[240]&~m[241])|(~m[221]&~m[237]&~m[238]&~m[240]&m[241])|(m[221]&~m[237]&~m[238]&~m[240]&m[241])|(m[221]&m[237]&~m[238]&~m[240]&m[241])|(m[221]&~m[237]&m[238]&~m[240]&m[241])|(~m[221]&~m[237]&~m[238]&m[240]&m[241])|(m[221]&~m[237]&~m[238]&m[240]&m[241])|(~m[221]&m[237]&~m[238]&m[240]&m[241])|(m[221]&m[237]&~m[238]&m[240]&m[241])|(~m[221]&~m[237]&m[238]&m[240]&m[241])|(m[221]&~m[237]&m[238]&m[240]&m[241])|(m[221]&m[237]&m[238]&m[240]&m[241]))):InitCond[144];
    m[244] = run?((((m[226]&~m[242]&~m[243]&~m[245]&~m[246])|(~m[226]&~m[242]&~m[243]&m[245]&~m[246])|(m[226]&m[242]&~m[243]&m[245]&~m[246])|(m[226]&~m[242]&m[243]&m[245]&~m[246])|(~m[226]&m[242]&~m[243]&~m[245]&m[246])|(~m[226]&~m[242]&m[243]&~m[245]&m[246])|(m[226]&m[242]&m[243]&~m[245]&m[246])|(~m[226]&m[242]&m[243]&m[245]&m[246]))&UnbiasedRNG[50])|((m[226]&~m[242]&~m[243]&m[245]&~m[246])|(~m[226]&~m[242]&~m[243]&~m[245]&m[246])|(m[226]&~m[242]&~m[243]&~m[245]&m[246])|(m[226]&m[242]&~m[243]&~m[245]&m[246])|(m[226]&~m[242]&m[243]&~m[245]&m[246])|(~m[226]&~m[242]&~m[243]&m[245]&m[246])|(m[226]&~m[242]&~m[243]&m[245]&m[246])|(~m[226]&m[242]&~m[243]&m[245]&m[246])|(m[226]&m[242]&~m[243]&m[245]&m[246])|(~m[226]&~m[242]&m[243]&m[245]&m[246])|(m[226]&~m[242]&m[243]&m[245]&m[246])|(m[226]&m[242]&m[243]&m[245]&m[246]))):InitCond[145];
    m[249] = run?((((m[231]&~m[247]&~m[248]&~m[250]&~m[251])|(~m[231]&~m[247]&~m[248]&m[250]&~m[251])|(m[231]&m[247]&~m[248]&m[250]&~m[251])|(m[231]&~m[247]&m[248]&m[250]&~m[251])|(~m[231]&m[247]&~m[248]&~m[250]&m[251])|(~m[231]&~m[247]&m[248]&~m[250]&m[251])|(m[231]&m[247]&m[248]&~m[250]&m[251])|(~m[231]&m[247]&m[248]&m[250]&m[251]))&UnbiasedRNG[51])|((m[231]&~m[247]&~m[248]&m[250]&~m[251])|(~m[231]&~m[247]&~m[248]&~m[250]&m[251])|(m[231]&~m[247]&~m[248]&~m[250]&m[251])|(m[231]&m[247]&~m[248]&~m[250]&m[251])|(m[231]&~m[247]&m[248]&~m[250]&m[251])|(~m[231]&~m[247]&~m[248]&m[250]&m[251])|(m[231]&~m[247]&~m[248]&m[250]&m[251])|(~m[231]&m[247]&~m[248]&m[250]&m[251])|(m[231]&m[247]&~m[248]&m[250]&m[251])|(~m[231]&~m[247]&m[248]&m[250]&m[251])|(m[231]&~m[247]&m[248]&m[250]&m[251])|(m[231]&m[247]&m[248]&m[250]&m[251]))):InitCond[146];
    m[254] = run?((((m[241]&~m[252]&~m[253]&~m[255]&~m[256])|(~m[241]&~m[252]&~m[253]&m[255]&~m[256])|(m[241]&m[252]&~m[253]&m[255]&~m[256])|(m[241]&~m[252]&m[253]&m[255]&~m[256])|(~m[241]&m[252]&~m[253]&~m[255]&m[256])|(~m[241]&~m[252]&m[253]&~m[255]&m[256])|(m[241]&m[252]&m[253]&~m[255]&m[256])|(~m[241]&m[252]&m[253]&m[255]&m[256]))&UnbiasedRNG[52])|((m[241]&~m[252]&~m[253]&m[255]&~m[256])|(~m[241]&~m[252]&~m[253]&~m[255]&m[256])|(m[241]&~m[252]&~m[253]&~m[255]&m[256])|(m[241]&m[252]&~m[253]&~m[255]&m[256])|(m[241]&~m[252]&m[253]&~m[255]&m[256])|(~m[241]&~m[252]&~m[253]&m[255]&m[256])|(m[241]&~m[252]&~m[253]&m[255]&m[256])|(~m[241]&m[252]&~m[253]&m[255]&m[256])|(m[241]&m[252]&~m[253]&m[255]&m[256])|(~m[241]&~m[252]&m[253]&m[255]&m[256])|(m[241]&~m[252]&m[253]&m[255]&m[256])|(m[241]&m[252]&m[253]&m[255]&m[256]))):InitCond[147];
    m[259] = run?((((m[246]&~m[257]&~m[258]&~m[260]&~m[261])|(~m[246]&~m[257]&~m[258]&m[260]&~m[261])|(m[246]&m[257]&~m[258]&m[260]&~m[261])|(m[246]&~m[257]&m[258]&m[260]&~m[261])|(~m[246]&m[257]&~m[258]&~m[260]&m[261])|(~m[246]&~m[257]&m[258]&~m[260]&m[261])|(m[246]&m[257]&m[258]&~m[260]&m[261])|(~m[246]&m[257]&m[258]&m[260]&m[261]))&UnbiasedRNG[53])|((m[246]&~m[257]&~m[258]&m[260]&~m[261])|(~m[246]&~m[257]&~m[258]&~m[260]&m[261])|(m[246]&~m[257]&~m[258]&~m[260]&m[261])|(m[246]&m[257]&~m[258]&~m[260]&m[261])|(m[246]&~m[257]&m[258]&~m[260]&m[261])|(~m[246]&~m[257]&~m[258]&m[260]&m[261])|(m[246]&~m[257]&~m[258]&m[260]&m[261])|(~m[246]&m[257]&~m[258]&m[260]&m[261])|(m[246]&m[257]&~m[258]&m[260]&m[261])|(~m[246]&~m[257]&m[258]&m[260]&m[261])|(m[246]&~m[257]&m[258]&m[260]&m[261])|(m[246]&m[257]&m[258]&m[260]&m[261]))):InitCond[148];
    m[264] = run?((((m[251]&~m[262]&~m[263]&~m[265]&~m[266])|(~m[251]&~m[262]&~m[263]&m[265]&~m[266])|(m[251]&m[262]&~m[263]&m[265]&~m[266])|(m[251]&~m[262]&m[263]&m[265]&~m[266])|(~m[251]&m[262]&~m[263]&~m[265]&m[266])|(~m[251]&~m[262]&m[263]&~m[265]&m[266])|(m[251]&m[262]&m[263]&~m[265]&m[266])|(~m[251]&m[262]&m[263]&m[265]&m[266]))&UnbiasedRNG[54])|((m[251]&~m[262]&~m[263]&m[265]&~m[266])|(~m[251]&~m[262]&~m[263]&~m[265]&m[266])|(m[251]&~m[262]&~m[263]&~m[265]&m[266])|(m[251]&m[262]&~m[263]&~m[265]&m[266])|(m[251]&~m[262]&m[263]&~m[265]&m[266])|(~m[251]&~m[262]&~m[263]&m[265]&m[266])|(m[251]&~m[262]&~m[263]&m[265]&m[266])|(~m[251]&m[262]&~m[263]&m[265]&m[266])|(m[251]&m[262]&~m[263]&m[265]&m[266])|(~m[251]&~m[262]&m[263]&m[265]&m[266])|(m[251]&~m[262]&m[263]&m[265]&m[266])|(m[251]&m[262]&m[263]&m[265]&m[266]))):InitCond[149];
    m[269] = run?((((m[261]&~m[267]&~m[268]&~m[270]&~m[271])|(~m[261]&~m[267]&~m[268]&m[270]&~m[271])|(m[261]&m[267]&~m[268]&m[270]&~m[271])|(m[261]&~m[267]&m[268]&m[270]&~m[271])|(~m[261]&m[267]&~m[268]&~m[270]&m[271])|(~m[261]&~m[267]&m[268]&~m[270]&m[271])|(m[261]&m[267]&m[268]&~m[270]&m[271])|(~m[261]&m[267]&m[268]&m[270]&m[271]))&UnbiasedRNG[55])|((m[261]&~m[267]&~m[268]&m[270]&~m[271])|(~m[261]&~m[267]&~m[268]&~m[270]&m[271])|(m[261]&~m[267]&~m[268]&~m[270]&m[271])|(m[261]&m[267]&~m[268]&~m[270]&m[271])|(m[261]&~m[267]&m[268]&~m[270]&m[271])|(~m[261]&~m[267]&~m[268]&m[270]&m[271])|(m[261]&~m[267]&~m[268]&m[270]&m[271])|(~m[261]&m[267]&~m[268]&m[270]&m[271])|(m[261]&m[267]&~m[268]&m[270]&m[271])|(~m[261]&~m[267]&m[268]&m[270]&m[271])|(m[261]&~m[267]&m[268]&m[270]&m[271])|(m[261]&m[267]&m[268]&m[270]&m[271]))):InitCond[150];
    m[274] = run?((((m[266]&~m[272]&~m[273]&~m[275]&~m[276])|(~m[266]&~m[272]&~m[273]&m[275]&~m[276])|(m[266]&m[272]&~m[273]&m[275]&~m[276])|(m[266]&~m[272]&m[273]&m[275]&~m[276])|(~m[266]&m[272]&~m[273]&~m[275]&m[276])|(~m[266]&~m[272]&m[273]&~m[275]&m[276])|(m[266]&m[272]&m[273]&~m[275]&m[276])|(~m[266]&m[272]&m[273]&m[275]&m[276]))&UnbiasedRNG[56])|((m[266]&~m[272]&~m[273]&m[275]&~m[276])|(~m[266]&~m[272]&~m[273]&~m[275]&m[276])|(m[266]&~m[272]&~m[273]&~m[275]&m[276])|(m[266]&m[272]&~m[273]&~m[275]&m[276])|(m[266]&~m[272]&m[273]&~m[275]&m[276])|(~m[266]&~m[272]&~m[273]&m[275]&m[276])|(m[266]&~m[272]&~m[273]&m[275]&m[276])|(~m[266]&m[272]&~m[273]&m[275]&m[276])|(m[266]&m[272]&~m[273]&m[275]&m[276])|(~m[266]&~m[272]&m[273]&m[275]&m[276])|(m[266]&~m[272]&m[273]&m[275]&m[276])|(m[266]&m[272]&m[273]&m[275]&m[276]))):InitCond[151];
    m[279] = run?((((m[276]&~m[277]&~m[278]&~m[280]&~m[281])|(~m[276]&~m[277]&~m[278]&m[280]&~m[281])|(m[276]&m[277]&~m[278]&m[280]&~m[281])|(m[276]&~m[277]&m[278]&m[280]&~m[281])|(~m[276]&m[277]&~m[278]&~m[280]&m[281])|(~m[276]&~m[277]&m[278]&~m[280]&m[281])|(m[276]&m[277]&m[278]&~m[280]&m[281])|(~m[276]&m[277]&m[278]&m[280]&m[281]))&UnbiasedRNG[57])|((m[276]&~m[277]&~m[278]&m[280]&~m[281])|(~m[276]&~m[277]&~m[278]&~m[280]&m[281])|(m[276]&~m[277]&~m[278]&~m[280]&m[281])|(m[276]&m[277]&~m[278]&~m[280]&m[281])|(m[276]&~m[277]&m[278]&~m[280]&m[281])|(~m[276]&~m[277]&~m[278]&m[280]&m[281])|(m[276]&~m[277]&~m[278]&m[280]&m[281])|(~m[276]&m[277]&~m[278]&m[280]&m[281])|(m[276]&m[277]&~m[278]&m[280]&m[281])|(~m[276]&~m[277]&m[278]&m[280]&m[281])|(m[276]&~m[277]&m[278]&m[280]&m[281])|(m[276]&m[277]&m[278]&m[280]&m[281]))):InitCond[152];
end

always @(posedge color2_clk) begin
    m[60] = run?((((~m[6]&~m[24]&~m[96])|(m[6]&m[24]&~m[96]))&BiasedRNG[95])|(((m[6]&~m[24]&~m[96])|(~m[6]&m[24]&m[96]))&~BiasedRNG[95])|((~m[6]&~m[24]&m[96])|(m[6]&~m[24]&m[96])|(m[6]&m[24]&m[96]))):InitCond[153];
    m[61] = run?((((~m[6]&~m[30]&~m[97])|(m[6]&m[30]&~m[97]))&BiasedRNG[96])|(((m[6]&~m[30]&~m[97])|(~m[6]&m[30]&m[97]))&~BiasedRNG[96])|((~m[6]&~m[30]&m[97])|(m[6]&~m[30]&m[97])|(m[6]&m[30]&m[97]))):InitCond[154];
    m[66] = run?((((~m[7]&~m[25]&~m[102])|(m[7]&m[25]&~m[102]))&BiasedRNG[97])|(((m[7]&~m[25]&~m[102])|(~m[7]&m[25]&m[102]))&~BiasedRNG[97])|((~m[7]&~m[25]&m[102])|(m[7]&~m[25]&m[102])|(m[7]&m[25]&m[102]))):InitCond[155];
    m[67] = run?((((~m[7]&~m[31]&~m[103])|(m[7]&m[31]&~m[103]))&BiasedRNG[98])|(((m[7]&~m[31]&~m[103])|(~m[7]&m[31]&m[103]))&~BiasedRNG[98])|((~m[7]&~m[31]&m[103])|(m[7]&~m[31]&m[103])|(m[7]&m[31]&m[103]))):InitCond[156];
    m[74] = run?((((~m[20]&~m[38]&~m[110])|(m[20]&m[38]&~m[110]))&BiasedRNG[99])|(((m[20]&~m[38]&~m[110])|(~m[20]&m[38]&m[110]))&~BiasedRNG[99])|((~m[20]&~m[38]&m[110])|(m[20]&~m[38]&m[110])|(m[20]&m[38]&m[110]))):InitCond[157];
    m[75] = run?((((~m[20]&~m[44]&~m[111])|(m[20]&m[44]&~m[111]))&BiasedRNG[100])|(((m[20]&~m[44]&~m[111])|(~m[20]&m[44]&m[111]))&~BiasedRNG[100])|((~m[20]&~m[44]&m[111])|(m[20]&~m[44]&m[111])|(m[20]&m[44]&m[111]))):InitCond[158];
    m[76] = run?((((~m[20]&~m[50]&~m[112])|(m[20]&m[50]&~m[112]))&BiasedRNG[101])|(((m[20]&~m[50]&~m[112])|(~m[20]&m[50]&m[112]))&~BiasedRNG[101])|((~m[20]&~m[50]&m[112])|(m[20]&~m[50]&m[112])|(m[20]&m[50]&m[112]))):InitCond[159];
    m[77] = run?((((~m[20]&~m[56]&~m[113])|(m[20]&m[56]&~m[113]))&BiasedRNG[102])|(((m[20]&~m[56]&~m[113])|(~m[20]&m[56]&m[113]))&~BiasedRNG[102])|((~m[20]&~m[56]&m[113])|(m[20]&~m[56]&m[113])|(m[20]&m[56]&m[113]))):InitCond[160];
    m[80] = run?((((~m[21]&~m[39]&~m[116])|(m[21]&m[39]&~m[116]))&BiasedRNG[103])|(((m[21]&~m[39]&~m[116])|(~m[21]&m[39]&m[116]))&~BiasedRNG[103])|((~m[21]&~m[39]&m[116])|(m[21]&~m[39]&m[116])|(m[21]&m[39]&m[116]))):InitCond[161];
    m[81] = run?((((~m[21]&~m[45]&~m[117])|(m[21]&m[45]&~m[117]))&BiasedRNG[104])|(((m[21]&~m[45]&~m[117])|(~m[21]&m[45]&m[117]))&~BiasedRNG[104])|((~m[21]&~m[45]&m[117])|(m[21]&~m[45]&m[117])|(m[21]&m[45]&m[117]))):InitCond[162];
    m[82] = run?((((~m[21]&~m[51]&~m[118])|(m[21]&m[51]&~m[118]))&BiasedRNG[105])|(((m[21]&~m[51]&~m[118])|(~m[21]&m[51]&m[118]))&~BiasedRNG[105])|((~m[21]&~m[51]&m[118])|(m[21]&~m[51]&m[118])|(m[21]&m[51]&m[118]))):InitCond[163];
    m[83] = run?((((~m[21]&~m[57]&~m[119])|(m[21]&m[57]&~m[119]))&BiasedRNG[106])|(((m[21]&~m[57]&~m[119])|(~m[21]&m[57]&m[119]))&~BiasedRNG[106])|((~m[21]&~m[57]&m[119])|(m[21]&~m[57]&m[119])|(m[21]&m[57]&m[119]))):InitCond[164];
    m[86] = run?((((~m[22]&~m[40]&~m[122])|(m[22]&m[40]&~m[122]))&BiasedRNG[107])|(((m[22]&~m[40]&~m[122])|(~m[22]&m[40]&m[122]))&~BiasedRNG[107])|((~m[22]&~m[40]&m[122])|(m[22]&~m[40]&m[122])|(m[22]&m[40]&m[122]))):InitCond[165];
    m[87] = run?((((~m[22]&~m[46]&~m[123])|(m[22]&m[46]&~m[123]))&BiasedRNG[108])|(((m[22]&~m[46]&~m[123])|(~m[22]&m[46]&m[123]))&~BiasedRNG[108])|((~m[22]&~m[46]&m[123])|(m[22]&~m[46]&m[123])|(m[22]&m[46]&m[123]))):InitCond[166];
    m[88] = run?((((~m[22]&~m[52]&~m[124])|(m[22]&m[52]&~m[124]))&BiasedRNG[109])|(((m[22]&~m[52]&~m[124])|(~m[22]&m[52]&m[124]))&~BiasedRNG[109])|((~m[22]&~m[52]&m[124])|(m[22]&~m[52]&m[124])|(m[22]&m[52]&m[124]))):InitCond[167];
    m[89] = run?((((~m[22]&~m[58]&~m[125])|(m[22]&m[58]&~m[125]))&BiasedRNG[110])|(((m[22]&~m[58]&~m[125])|(~m[22]&m[58]&m[125]))&~BiasedRNG[110])|((~m[22]&~m[58]&m[125])|(m[22]&~m[58]&m[125])|(m[22]&m[58]&m[125]))):InitCond[168];
    m[92] = run?((((~m[23]&~m[41]&~m[128])|(m[23]&m[41]&~m[128]))&BiasedRNG[111])|(((m[23]&~m[41]&~m[128])|(~m[23]&m[41]&m[128]))&~BiasedRNG[111])|((~m[23]&~m[41]&m[128])|(m[23]&~m[41]&m[128])|(m[23]&m[41]&m[128]))):InitCond[169];
    m[93] = run?((((~m[23]&~m[47]&~m[129])|(m[23]&m[47]&~m[129]))&BiasedRNG[112])|(((m[23]&~m[47]&~m[129])|(~m[23]&m[47]&m[129]))&~BiasedRNG[112])|((~m[23]&~m[47]&m[129])|(m[23]&~m[47]&m[129])|(m[23]&m[47]&m[129]))):InitCond[170];
    m[94] = run?((((~m[23]&~m[53]&~m[130])|(m[23]&m[53]&~m[130]))&BiasedRNG[113])|(((m[23]&~m[53]&~m[130])|(~m[23]&m[53]&m[130]))&~BiasedRNG[113])|((~m[23]&~m[53]&m[130])|(m[23]&~m[53]&m[130])|(m[23]&m[53]&m[130]))):InitCond[171];
    m[95] = run?((((~m[23]&~m[59]&~m[131])|(m[23]&m[59]&~m[131]))&BiasedRNG[114])|(((m[23]&~m[59]&~m[131])|(~m[23]&m[59]&m[131]))&~BiasedRNG[114])|((~m[23]&~m[59]&m[131])|(m[23]&~m[59]&m[131])|(m[23]&m[59]&m[131]))):InitCond[172];
    m[98] = run?((((m[36]&~m[62]&m[137])|(~m[36]&m[62]&m[137]))&BiasedRNG[115])|(((m[36]&m[62]&~m[137]))&~BiasedRNG[115])|((m[36]&m[62]&m[137]))):InitCond[173];
    m[99] = run?((((m[42]&~m[63]&m[147])|(~m[42]&m[63]&m[147]))&BiasedRNG[116])|(((m[42]&m[63]&~m[147]))&~BiasedRNG[116])|((m[42]&m[63]&m[147]))):InitCond[174];
    m[100] = run?((((m[48]&~m[64]&m[162])|(~m[48]&m[64]&m[162]))&BiasedRNG[117])|(((m[48]&m[64]&~m[162]))&~BiasedRNG[117])|((m[48]&m[64]&m[162]))):InitCond[175];
    m[101] = run?((((m[54]&~m[65]&m[182])|(~m[54]&m[65]&m[182]))&BiasedRNG[118])|(((m[54]&m[65]&~m[182]))&~BiasedRNG[118])|((m[54]&m[65]&m[182]))):InitCond[176];
    m[104] = run?((((m[37]&~m[68]&m[148])|(~m[37]&m[68]&m[148]))&BiasedRNG[119])|(((m[37]&m[68]&~m[148]))&~BiasedRNG[119])|((m[37]&m[68]&m[148]))):InitCond[177];
    m[105] = run?((((m[43]&~m[69]&m[163])|(~m[43]&m[69]&m[163]))&BiasedRNG[120])|(((m[43]&m[69]&~m[163]))&~BiasedRNG[120])|((m[43]&m[69]&m[163]))):InitCond[178];
    m[106] = run?((((m[49]&~m[70]&m[183])|(~m[49]&m[70]&m[183]))&BiasedRNG[121])|(((m[49]&m[70]&~m[183]))&~BiasedRNG[121])|((m[49]&m[70]&m[183]))):InitCond[179];
    m[107] = run?((((m[55]&~m[71]&m[208])|(~m[55]&m[71]&m[208]))&BiasedRNG[122])|(((m[55]&m[71]&~m[208]))&~BiasedRNG[122])|((m[55]&m[71]&m[208]))):InitCond[180];
    m[108] = run?((((m[26]&~m[72]&m[143])|(~m[26]&m[72]&m[143]))&BiasedRNG[123])|(((m[26]&m[72]&~m[143]))&~BiasedRNG[123])|((m[26]&m[72]&m[143]))):InitCond[181];
    m[109] = run?((((m[32]&~m[73]&m[153])|(~m[32]&m[73]&m[153]))&BiasedRNG[124])|(((m[32]&m[73]&~m[153]))&~BiasedRNG[124])|((m[32]&m[73]&m[153]))):InitCond[182];
    m[114] = run?((((m[27]&~m[78]&m[158])|(~m[27]&m[78]&m[158]))&BiasedRNG[125])|(((m[27]&m[78]&~m[158]))&~BiasedRNG[125])|((m[27]&m[78]&m[158]))):InitCond[183];
    m[115] = run?((((m[33]&~m[79]&m[173])|(~m[33]&m[79]&m[173]))&BiasedRNG[126])|(((m[33]&m[79]&~m[173]))&~BiasedRNG[126])|((m[33]&m[79]&m[173]))):InitCond[184];
    m[120] = run?((((m[28]&~m[84]&m[178])|(~m[28]&m[84]&m[178]))&BiasedRNG[127])|(((m[28]&m[84]&~m[178]))&~BiasedRNG[127])|((m[28]&m[84]&m[178]))):InitCond[185];
    m[121] = run?((((m[34]&~m[85]&m[198])|(~m[34]&m[85]&m[198]))&BiasedRNG[128])|(((m[34]&m[85]&~m[198]))&~BiasedRNG[128])|((m[34]&m[85]&m[198]))):InitCond[186];
    m[126] = run?((((m[29]&~m[90]&m[203])|(~m[29]&m[90]&m[203]))&BiasedRNG[129])|(((m[29]&m[90]&~m[203]))&~BiasedRNG[129])|((m[29]&m[90]&m[203]))):InitCond[187];
    m[127] = run?((((m[35]&~m[91]&m[228])|(~m[35]&m[91]&m[228]))&BiasedRNG[130])|(((m[35]&m[91]&~m[228]))&~BiasedRNG[130])|((m[35]&m[91]&m[228]))):InitCond[188];
    m[133] = run?((((m[102]&~m[132]&~m[134]&~m[135]&~m[136])|(~m[102]&~m[132]&~m[134]&m[135]&~m[136])|(m[102]&m[132]&~m[134]&m[135]&~m[136])|(m[102]&~m[132]&m[134]&m[135]&~m[136])|(~m[102]&m[132]&~m[134]&~m[135]&m[136])|(~m[102]&~m[132]&m[134]&~m[135]&m[136])|(m[102]&m[132]&m[134]&~m[135]&m[136])|(~m[102]&m[132]&m[134]&m[135]&m[136]))&UnbiasedRNG[58])|((m[102]&~m[132]&~m[134]&m[135]&~m[136])|(~m[102]&~m[132]&~m[134]&~m[135]&m[136])|(m[102]&~m[132]&~m[134]&~m[135]&m[136])|(m[102]&m[132]&~m[134]&~m[135]&m[136])|(m[102]&~m[132]&m[134]&~m[135]&m[136])|(~m[102]&~m[132]&~m[134]&m[135]&m[136])|(m[102]&~m[132]&~m[134]&m[135]&m[136])|(~m[102]&m[132]&~m[134]&m[135]&m[136])|(m[102]&m[132]&~m[134]&m[135]&m[136])|(~m[102]&~m[132]&m[134]&m[135]&m[136])|(m[102]&~m[132]&m[134]&m[135]&m[136])|(m[102]&m[132]&m[134]&m[135]&m[136]))):InitCond[189];
    m[139] = run?((((m[136]&~m[137]&~m[138]&~m[140]&~m[141])|(~m[136]&~m[137]&~m[138]&m[140]&~m[141])|(m[136]&m[137]&~m[138]&m[140]&~m[141])|(m[136]&~m[137]&m[138]&m[140]&~m[141])|(~m[136]&m[137]&~m[138]&~m[140]&m[141])|(~m[136]&~m[137]&m[138]&~m[140]&m[141])|(m[136]&m[137]&m[138]&~m[140]&m[141])|(~m[136]&m[137]&m[138]&m[140]&m[141]))&UnbiasedRNG[59])|((m[136]&~m[137]&~m[138]&m[140]&~m[141])|(~m[136]&~m[137]&~m[138]&~m[140]&m[141])|(m[136]&~m[137]&~m[138]&~m[140]&m[141])|(m[136]&m[137]&~m[138]&~m[140]&m[141])|(m[136]&~m[137]&m[138]&~m[140]&m[141])|(~m[136]&~m[137]&~m[138]&m[140]&m[141])|(m[136]&~m[137]&~m[138]&m[140]&m[141])|(~m[136]&m[137]&~m[138]&m[140]&m[141])|(m[136]&m[137]&~m[138]&m[140]&m[141])|(~m[136]&~m[137]&m[138]&m[140]&m[141])|(m[136]&~m[137]&m[138]&m[140]&m[141])|(m[136]&m[137]&m[138]&m[140]&m[141]))):InitCond[190];
    m[149] = run?((((m[141]&~m[147]&~m[148]&~m[150]&~m[151])|(~m[141]&~m[147]&~m[148]&m[150]&~m[151])|(m[141]&m[147]&~m[148]&m[150]&~m[151])|(m[141]&~m[147]&m[148]&m[150]&~m[151])|(~m[141]&m[147]&~m[148]&~m[150]&m[151])|(~m[141]&~m[147]&m[148]&~m[150]&m[151])|(m[141]&m[147]&m[148]&~m[150]&m[151])|(~m[141]&m[147]&m[148]&m[150]&m[151]))&UnbiasedRNG[60])|((m[141]&~m[147]&~m[148]&m[150]&~m[151])|(~m[141]&~m[147]&~m[148]&~m[150]&m[151])|(m[141]&~m[147]&~m[148]&~m[150]&m[151])|(m[141]&m[147]&~m[148]&~m[150]&m[151])|(m[141]&~m[147]&m[148]&~m[150]&m[151])|(~m[141]&~m[147]&~m[148]&m[150]&m[151])|(m[141]&~m[147]&~m[148]&m[150]&m[151])|(~m[141]&m[147]&~m[148]&m[150]&m[151])|(m[141]&m[147]&~m[148]&m[150]&m[151])|(~m[141]&~m[147]&m[148]&m[150]&m[151])|(m[141]&~m[147]&m[148]&m[150]&m[151])|(m[141]&m[147]&m[148]&m[150]&m[151]))):InitCond[191];
    m[154] = run?((((m[146]&~m[152]&~m[153]&~m[155]&~m[156])|(~m[146]&~m[152]&~m[153]&m[155]&~m[156])|(m[146]&m[152]&~m[153]&m[155]&~m[156])|(m[146]&~m[152]&m[153]&m[155]&~m[156])|(~m[146]&m[152]&~m[153]&~m[155]&m[156])|(~m[146]&~m[152]&m[153]&~m[155]&m[156])|(m[146]&m[152]&m[153]&~m[155]&m[156])|(~m[146]&m[152]&m[153]&m[155]&m[156]))&UnbiasedRNG[61])|((m[146]&~m[152]&~m[153]&m[155]&~m[156])|(~m[146]&~m[152]&~m[153]&~m[155]&m[156])|(m[146]&~m[152]&~m[153]&~m[155]&m[156])|(m[146]&m[152]&~m[153]&~m[155]&m[156])|(m[146]&~m[152]&m[153]&~m[155]&m[156])|(~m[146]&~m[152]&~m[153]&m[155]&m[156])|(m[146]&~m[152]&~m[153]&m[155]&m[156])|(~m[146]&m[152]&~m[153]&m[155]&m[156])|(m[146]&m[152]&~m[153]&m[155]&m[156])|(~m[146]&~m[152]&m[153]&m[155]&m[156])|(m[146]&~m[152]&m[153]&m[155]&m[156])|(m[146]&m[152]&m[153]&m[155]&m[156]))):InitCond[192];
    m[164] = run?((((m[151]&~m[162]&~m[163]&~m[165]&~m[166])|(~m[151]&~m[162]&~m[163]&m[165]&~m[166])|(m[151]&m[162]&~m[163]&m[165]&~m[166])|(m[151]&~m[162]&m[163]&m[165]&~m[166])|(~m[151]&m[162]&~m[163]&~m[165]&m[166])|(~m[151]&~m[162]&m[163]&~m[165]&m[166])|(m[151]&m[162]&m[163]&~m[165]&m[166])|(~m[151]&m[162]&m[163]&m[165]&m[166]))&UnbiasedRNG[62])|((m[151]&~m[162]&~m[163]&m[165]&~m[166])|(~m[151]&~m[162]&~m[163]&~m[165]&m[166])|(m[151]&~m[162]&~m[163]&~m[165]&m[166])|(m[151]&m[162]&~m[163]&~m[165]&m[166])|(m[151]&~m[162]&m[163]&~m[165]&m[166])|(~m[151]&~m[162]&~m[163]&m[165]&m[166])|(m[151]&~m[162]&~m[163]&m[165]&m[166])|(~m[151]&m[162]&~m[163]&m[165]&m[166])|(m[151]&m[162]&~m[163]&m[165]&m[166])|(~m[151]&~m[162]&m[163]&m[165]&m[166])|(m[151]&~m[162]&m[163]&m[165]&m[166])|(m[151]&m[162]&m[163]&m[165]&m[166]))):InitCond[193];
    m[168] = run?((((m[110]&~m[167]&~m[169]&~m[170]&~m[171])|(~m[110]&~m[167]&~m[169]&m[170]&~m[171])|(m[110]&m[167]&~m[169]&m[170]&~m[171])|(m[110]&~m[167]&m[169]&m[170]&~m[171])|(~m[110]&m[167]&~m[169]&~m[170]&m[171])|(~m[110]&~m[167]&m[169]&~m[170]&m[171])|(m[110]&m[167]&m[169]&~m[170]&m[171])|(~m[110]&m[167]&m[169]&m[170]&m[171]))&UnbiasedRNG[63])|((m[110]&~m[167]&~m[169]&m[170]&~m[171])|(~m[110]&~m[167]&~m[169]&~m[170]&m[171])|(m[110]&~m[167]&~m[169]&~m[170]&m[171])|(m[110]&m[167]&~m[169]&~m[170]&m[171])|(m[110]&~m[167]&m[169]&~m[170]&m[171])|(~m[110]&~m[167]&~m[169]&m[170]&m[171])|(m[110]&~m[167]&~m[169]&m[170]&m[171])|(~m[110]&m[167]&~m[169]&m[170]&m[171])|(m[110]&m[167]&~m[169]&m[170]&m[171])|(~m[110]&~m[167]&m[169]&m[170]&m[171])|(m[110]&~m[167]&m[169]&m[170]&m[171])|(m[110]&m[167]&m[169]&m[170]&m[171]))):InitCond[194];
    m[174] = run?((((m[161]&~m[172]&~m[173]&~m[175]&~m[176])|(~m[161]&~m[172]&~m[173]&m[175]&~m[176])|(m[161]&m[172]&~m[173]&m[175]&~m[176])|(m[161]&~m[172]&m[173]&m[175]&~m[176])|(~m[161]&m[172]&~m[173]&~m[175]&m[176])|(~m[161]&~m[172]&m[173]&~m[175]&m[176])|(m[161]&m[172]&m[173]&~m[175]&m[176])|(~m[161]&m[172]&m[173]&m[175]&m[176]))&UnbiasedRNG[64])|((m[161]&~m[172]&~m[173]&m[175]&~m[176])|(~m[161]&~m[172]&~m[173]&~m[175]&m[176])|(m[161]&~m[172]&~m[173]&~m[175]&m[176])|(m[161]&m[172]&~m[173]&~m[175]&m[176])|(m[161]&~m[172]&m[173]&~m[175]&m[176])|(~m[161]&~m[172]&~m[173]&m[175]&m[176])|(m[161]&~m[172]&~m[173]&m[175]&m[176])|(~m[161]&m[172]&~m[173]&m[175]&m[176])|(m[161]&m[172]&~m[173]&m[175]&m[176])|(~m[161]&~m[172]&m[173]&m[175]&m[176])|(m[161]&~m[172]&m[173]&m[175]&m[176])|(m[161]&m[172]&m[173]&m[175]&m[176]))):InitCond[195];
    m[184] = run?((((m[166]&~m[182]&~m[183]&~m[185]&~m[186])|(~m[166]&~m[182]&~m[183]&m[185]&~m[186])|(m[166]&m[182]&~m[183]&m[185]&~m[186])|(m[166]&~m[182]&m[183]&m[185]&~m[186])|(~m[166]&m[182]&~m[183]&~m[185]&m[186])|(~m[166]&~m[182]&m[183]&~m[185]&m[186])|(m[166]&m[182]&m[183]&~m[185]&m[186])|(~m[166]&m[182]&m[183]&m[185]&m[186]))&UnbiasedRNG[65])|((m[166]&~m[182]&~m[183]&m[185]&~m[186])|(~m[166]&~m[182]&~m[183]&~m[185]&m[186])|(m[166]&~m[182]&~m[183]&~m[185]&m[186])|(m[166]&m[182]&~m[183]&~m[185]&m[186])|(m[166]&~m[182]&m[183]&~m[185]&m[186])|(~m[166]&~m[182]&~m[183]&m[185]&m[186])|(m[166]&~m[182]&~m[183]&m[185]&m[186])|(~m[166]&m[182]&~m[183]&m[185]&m[186])|(m[166]&m[182]&~m[183]&m[185]&m[186])|(~m[166]&~m[182]&m[183]&m[185]&m[186])|(m[166]&~m[182]&m[183]&m[185]&m[186])|(m[166]&m[182]&m[183]&m[185]&m[186]))):InitCond[196];
    m[188] = run?((((m[111]&~m[187]&~m[189]&~m[190]&~m[191])|(~m[111]&~m[187]&~m[189]&m[190]&~m[191])|(m[111]&m[187]&~m[189]&m[190]&~m[191])|(m[111]&~m[187]&m[189]&m[190]&~m[191])|(~m[111]&m[187]&~m[189]&~m[190]&m[191])|(~m[111]&~m[187]&m[189]&~m[190]&m[191])|(m[111]&m[187]&m[189]&~m[190]&m[191])|(~m[111]&m[187]&m[189]&m[190]&m[191]))&UnbiasedRNG[66])|((m[111]&~m[187]&~m[189]&m[190]&~m[191])|(~m[111]&~m[187]&~m[189]&~m[190]&m[191])|(m[111]&~m[187]&~m[189]&~m[190]&m[191])|(m[111]&m[187]&~m[189]&~m[190]&m[191])|(m[111]&~m[187]&m[189]&~m[190]&m[191])|(~m[111]&~m[187]&~m[189]&m[190]&m[191])|(m[111]&~m[187]&~m[189]&m[190]&m[191])|(~m[111]&m[187]&~m[189]&m[190]&m[191])|(m[111]&m[187]&~m[189]&m[190]&m[191])|(~m[111]&~m[187]&m[189]&m[190]&m[191])|(m[111]&~m[187]&m[189]&m[190]&m[191])|(m[111]&m[187]&m[189]&m[190]&m[191]))):InitCond[197];
    m[193] = run?((((m[116]&~m[192]&~m[194]&~m[195]&~m[196])|(~m[116]&~m[192]&~m[194]&m[195]&~m[196])|(m[116]&m[192]&~m[194]&m[195]&~m[196])|(m[116]&~m[192]&m[194]&m[195]&~m[196])|(~m[116]&m[192]&~m[194]&~m[195]&m[196])|(~m[116]&~m[192]&m[194]&~m[195]&m[196])|(m[116]&m[192]&m[194]&~m[195]&m[196])|(~m[116]&m[192]&m[194]&m[195]&m[196]))&UnbiasedRNG[67])|((m[116]&~m[192]&~m[194]&m[195]&~m[196])|(~m[116]&~m[192]&~m[194]&~m[195]&m[196])|(m[116]&~m[192]&~m[194]&~m[195]&m[196])|(m[116]&m[192]&~m[194]&~m[195]&m[196])|(m[116]&~m[192]&m[194]&~m[195]&m[196])|(~m[116]&~m[192]&~m[194]&m[195]&m[196])|(m[116]&~m[192]&~m[194]&m[195]&m[196])|(~m[116]&m[192]&~m[194]&m[195]&m[196])|(m[116]&m[192]&~m[194]&m[195]&m[196])|(~m[116]&~m[192]&m[194]&m[195]&m[196])|(m[116]&~m[192]&m[194]&m[195]&m[196])|(m[116]&m[192]&m[194]&m[195]&m[196]))):InitCond[198];
    m[199] = run?((((m[181]&~m[197]&~m[198]&~m[200]&~m[201])|(~m[181]&~m[197]&~m[198]&m[200]&~m[201])|(m[181]&m[197]&~m[198]&m[200]&~m[201])|(m[181]&~m[197]&m[198]&m[200]&~m[201])|(~m[181]&m[197]&~m[198]&~m[200]&m[201])|(~m[181]&~m[197]&m[198]&~m[200]&m[201])|(m[181]&m[197]&m[198]&~m[200]&m[201])|(~m[181]&m[197]&m[198]&m[200]&m[201]))&UnbiasedRNG[68])|((m[181]&~m[197]&~m[198]&m[200]&~m[201])|(~m[181]&~m[197]&~m[198]&~m[200]&m[201])|(m[181]&~m[197]&~m[198]&~m[200]&m[201])|(m[181]&m[197]&~m[198]&~m[200]&m[201])|(m[181]&~m[197]&m[198]&~m[200]&m[201])|(~m[181]&~m[197]&~m[198]&m[200]&m[201])|(m[181]&~m[197]&~m[198]&m[200]&m[201])|(~m[181]&m[197]&~m[198]&m[200]&m[201])|(m[181]&m[197]&~m[198]&m[200]&m[201])|(~m[181]&~m[197]&m[198]&m[200]&m[201])|(m[181]&~m[197]&m[198]&m[200]&m[201])|(m[181]&m[197]&m[198]&m[200]&m[201]))):InitCond[199];
    m[209] = run?((((m[186]&~m[207]&~m[208]&~m[210]&~m[211])|(~m[186]&~m[207]&~m[208]&m[210]&~m[211])|(m[186]&m[207]&~m[208]&m[210]&~m[211])|(m[186]&~m[207]&m[208]&m[210]&~m[211])|(~m[186]&m[207]&~m[208]&~m[210]&m[211])|(~m[186]&~m[207]&m[208]&~m[210]&m[211])|(m[186]&m[207]&m[208]&~m[210]&m[211])|(~m[186]&m[207]&m[208]&m[210]&m[211]))&UnbiasedRNG[69])|((m[186]&~m[207]&~m[208]&m[210]&~m[211])|(~m[186]&~m[207]&~m[208]&~m[210]&m[211])|(m[186]&~m[207]&~m[208]&~m[210]&m[211])|(m[186]&m[207]&~m[208]&~m[210]&m[211])|(m[186]&~m[207]&m[208]&~m[210]&m[211])|(~m[186]&~m[207]&~m[208]&m[210]&m[211])|(m[186]&~m[207]&~m[208]&m[210]&m[211])|(~m[186]&m[207]&~m[208]&m[210]&m[211])|(m[186]&m[207]&~m[208]&m[210]&m[211])|(~m[186]&~m[207]&m[208]&m[210]&m[211])|(m[186]&~m[207]&m[208]&m[210]&m[211])|(m[186]&m[207]&m[208]&m[210]&m[211]))):InitCond[200];
    m[213] = run?((((m[112]&~m[212]&~m[214]&~m[215]&~m[216])|(~m[112]&~m[212]&~m[214]&m[215]&~m[216])|(m[112]&m[212]&~m[214]&m[215]&~m[216])|(m[112]&~m[212]&m[214]&m[215]&~m[216])|(~m[112]&m[212]&~m[214]&~m[215]&m[216])|(~m[112]&~m[212]&m[214]&~m[215]&m[216])|(m[112]&m[212]&m[214]&~m[215]&m[216])|(~m[112]&m[212]&m[214]&m[215]&m[216]))&UnbiasedRNG[70])|((m[112]&~m[212]&~m[214]&m[215]&~m[216])|(~m[112]&~m[212]&~m[214]&~m[215]&m[216])|(m[112]&~m[212]&~m[214]&~m[215]&m[216])|(m[112]&m[212]&~m[214]&~m[215]&m[216])|(m[112]&~m[212]&m[214]&~m[215]&m[216])|(~m[112]&~m[212]&~m[214]&m[215]&m[216])|(m[112]&~m[212]&~m[214]&m[215]&m[216])|(~m[112]&m[212]&~m[214]&m[215]&m[216])|(m[112]&m[212]&~m[214]&m[215]&m[216])|(~m[112]&~m[212]&m[214]&m[215]&m[216])|(m[112]&~m[212]&m[214]&m[215]&m[216])|(m[112]&m[212]&m[214]&m[215]&m[216]))):InitCond[201];
    m[218] = run?((((m[117]&~m[217]&~m[219]&~m[220]&~m[221])|(~m[117]&~m[217]&~m[219]&m[220]&~m[221])|(m[117]&m[217]&~m[219]&m[220]&~m[221])|(m[117]&~m[217]&m[219]&m[220]&~m[221])|(~m[117]&m[217]&~m[219]&~m[220]&m[221])|(~m[117]&~m[217]&m[219]&~m[220]&m[221])|(m[117]&m[217]&m[219]&~m[220]&m[221])|(~m[117]&m[217]&m[219]&m[220]&m[221]))&UnbiasedRNG[71])|((m[117]&~m[217]&~m[219]&m[220]&~m[221])|(~m[117]&~m[217]&~m[219]&~m[220]&m[221])|(m[117]&~m[217]&~m[219]&~m[220]&m[221])|(m[117]&m[217]&~m[219]&~m[220]&m[221])|(m[117]&~m[217]&m[219]&~m[220]&m[221])|(~m[117]&~m[217]&~m[219]&m[220]&m[221])|(m[117]&~m[217]&~m[219]&m[220]&m[221])|(~m[117]&m[217]&~m[219]&m[220]&m[221])|(m[117]&m[217]&~m[219]&m[220]&m[221])|(~m[117]&~m[217]&m[219]&m[220]&m[221])|(m[117]&~m[217]&m[219]&m[220]&m[221])|(m[117]&m[217]&m[219]&m[220]&m[221]))):InitCond[202];
    m[223] = run?((((m[122]&~m[222]&~m[224]&~m[225]&~m[226])|(~m[122]&~m[222]&~m[224]&m[225]&~m[226])|(m[122]&m[222]&~m[224]&m[225]&~m[226])|(m[122]&~m[222]&m[224]&m[225]&~m[226])|(~m[122]&m[222]&~m[224]&~m[225]&m[226])|(~m[122]&~m[222]&m[224]&~m[225]&m[226])|(m[122]&m[222]&m[224]&~m[225]&m[226])|(~m[122]&m[222]&m[224]&m[225]&m[226]))&UnbiasedRNG[72])|((m[122]&~m[222]&~m[224]&m[225]&~m[226])|(~m[122]&~m[222]&~m[224]&~m[225]&m[226])|(m[122]&~m[222]&~m[224]&~m[225]&m[226])|(m[122]&m[222]&~m[224]&~m[225]&m[226])|(m[122]&~m[222]&m[224]&~m[225]&m[226])|(~m[122]&~m[222]&~m[224]&m[225]&m[226])|(m[122]&~m[222]&~m[224]&m[225]&m[226])|(~m[122]&m[222]&~m[224]&m[225]&m[226])|(m[122]&m[222]&~m[224]&m[225]&m[226])|(~m[122]&~m[222]&m[224]&m[225]&m[226])|(m[122]&~m[222]&m[224]&m[225]&m[226])|(m[122]&m[222]&m[224]&m[225]&m[226]))):InitCond[203];
    m[229] = run?((((m[206]&~m[227]&~m[228]&~m[230]&~m[231])|(~m[206]&~m[227]&~m[228]&m[230]&~m[231])|(m[206]&m[227]&~m[228]&m[230]&~m[231])|(m[206]&~m[227]&m[228]&m[230]&~m[231])|(~m[206]&m[227]&~m[228]&~m[230]&m[231])|(~m[206]&~m[227]&m[228]&~m[230]&m[231])|(m[206]&m[227]&m[228]&~m[230]&m[231])|(~m[206]&m[227]&m[228]&m[230]&m[231]))&UnbiasedRNG[73])|((m[206]&~m[227]&~m[228]&m[230]&~m[231])|(~m[206]&~m[227]&~m[228]&~m[230]&m[231])|(m[206]&~m[227]&~m[228]&~m[230]&m[231])|(m[206]&m[227]&~m[228]&~m[230]&m[231])|(m[206]&~m[227]&m[228]&~m[230]&m[231])|(~m[206]&~m[227]&~m[228]&m[230]&m[231])|(m[206]&~m[227]&~m[228]&m[230]&m[231])|(~m[206]&m[227]&~m[228]&m[230]&m[231])|(m[206]&m[227]&~m[228]&m[230]&m[231])|(~m[206]&~m[227]&m[228]&m[230]&m[231])|(m[206]&~m[227]&m[228]&m[230]&m[231])|(m[206]&m[227]&m[228]&m[230]&m[231]))):InitCond[204];
    m[233] = run?((((m[113]&~m[232]&~m[234]&~m[235]&~m[236])|(~m[113]&~m[232]&~m[234]&m[235]&~m[236])|(m[113]&m[232]&~m[234]&m[235]&~m[236])|(m[113]&~m[232]&m[234]&m[235]&~m[236])|(~m[113]&m[232]&~m[234]&~m[235]&m[236])|(~m[113]&~m[232]&m[234]&~m[235]&m[236])|(m[113]&m[232]&m[234]&~m[235]&m[236])|(~m[113]&m[232]&m[234]&m[235]&m[236]))&UnbiasedRNG[74])|((m[113]&~m[232]&~m[234]&m[235]&~m[236])|(~m[113]&~m[232]&~m[234]&~m[235]&m[236])|(m[113]&~m[232]&~m[234]&~m[235]&m[236])|(m[113]&m[232]&~m[234]&~m[235]&m[236])|(m[113]&~m[232]&m[234]&~m[235]&m[236])|(~m[113]&~m[232]&~m[234]&m[235]&m[236])|(m[113]&~m[232]&~m[234]&m[235]&m[236])|(~m[113]&m[232]&~m[234]&m[235]&m[236])|(m[113]&m[232]&~m[234]&m[235]&m[236])|(~m[113]&~m[232]&m[234]&m[235]&m[236])|(m[113]&~m[232]&m[234]&m[235]&m[236])|(m[113]&m[232]&m[234]&m[235]&m[236]))):InitCond[205];
    m[238] = run?((((m[118]&~m[237]&~m[239]&~m[240]&~m[241])|(~m[118]&~m[237]&~m[239]&m[240]&~m[241])|(m[118]&m[237]&~m[239]&m[240]&~m[241])|(m[118]&~m[237]&m[239]&m[240]&~m[241])|(~m[118]&m[237]&~m[239]&~m[240]&m[241])|(~m[118]&~m[237]&m[239]&~m[240]&m[241])|(m[118]&m[237]&m[239]&~m[240]&m[241])|(~m[118]&m[237]&m[239]&m[240]&m[241]))&UnbiasedRNG[75])|((m[118]&~m[237]&~m[239]&m[240]&~m[241])|(~m[118]&~m[237]&~m[239]&~m[240]&m[241])|(m[118]&~m[237]&~m[239]&~m[240]&m[241])|(m[118]&m[237]&~m[239]&~m[240]&m[241])|(m[118]&~m[237]&m[239]&~m[240]&m[241])|(~m[118]&~m[237]&~m[239]&m[240]&m[241])|(m[118]&~m[237]&~m[239]&m[240]&m[241])|(~m[118]&m[237]&~m[239]&m[240]&m[241])|(m[118]&m[237]&~m[239]&m[240]&m[241])|(~m[118]&~m[237]&m[239]&m[240]&m[241])|(m[118]&~m[237]&m[239]&m[240]&m[241])|(m[118]&m[237]&m[239]&m[240]&m[241]))):InitCond[206];
    m[243] = run?((((m[123]&~m[242]&~m[244]&~m[245]&~m[246])|(~m[123]&~m[242]&~m[244]&m[245]&~m[246])|(m[123]&m[242]&~m[244]&m[245]&~m[246])|(m[123]&~m[242]&m[244]&m[245]&~m[246])|(~m[123]&m[242]&~m[244]&~m[245]&m[246])|(~m[123]&~m[242]&m[244]&~m[245]&m[246])|(m[123]&m[242]&m[244]&~m[245]&m[246])|(~m[123]&m[242]&m[244]&m[245]&m[246]))&UnbiasedRNG[76])|((m[123]&~m[242]&~m[244]&m[245]&~m[246])|(~m[123]&~m[242]&~m[244]&~m[245]&m[246])|(m[123]&~m[242]&~m[244]&~m[245]&m[246])|(m[123]&m[242]&~m[244]&~m[245]&m[246])|(m[123]&~m[242]&m[244]&~m[245]&m[246])|(~m[123]&~m[242]&~m[244]&m[245]&m[246])|(m[123]&~m[242]&~m[244]&m[245]&m[246])|(~m[123]&m[242]&~m[244]&m[245]&m[246])|(m[123]&m[242]&~m[244]&m[245]&m[246])|(~m[123]&~m[242]&m[244]&m[245]&m[246])|(m[123]&~m[242]&m[244]&m[245]&m[246])|(m[123]&m[242]&m[244]&m[245]&m[246]))):InitCond[207];
    m[248] = run?((((m[128]&~m[247]&~m[249]&~m[250]&~m[251])|(~m[128]&~m[247]&~m[249]&m[250]&~m[251])|(m[128]&m[247]&~m[249]&m[250]&~m[251])|(m[128]&~m[247]&m[249]&m[250]&~m[251])|(~m[128]&m[247]&~m[249]&~m[250]&m[251])|(~m[128]&~m[247]&m[249]&~m[250]&m[251])|(m[128]&m[247]&m[249]&~m[250]&m[251])|(~m[128]&m[247]&m[249]&m[250]&m[251]))&UnbiasedRNG[77])|((m[128]&~m[247]&~m[249]&m[250]&~m[251])|(~m[128]&~m[247]&~m[249]&~m[250]&m[251])|(m[128]&~m[247]&~m[249]&~m[250]&m[251])|(m[128]&m[247]&~m[249]&~m[250]&m[251])|(m[128]&~m[247]&m[249]&~m[250]&m[251])|(~m[128]&~m[247]&~m[249]&m[250]&m[251])|(m[128]&~m[247]&~m[249]&m[250]&m[251])|(~m[128]&m[247]&~m[249]&m[250]&m[251])|(m[128]&m[247]&~m[249]&m[250]&m[251])|(~m[128]&~m[247]&m[249]&m[250]&m[251])|(m[128]&~m[247]&m[249]&m[250]&m[251])|(m[128]&m[247]&m[249]&m[250]&m[251]))):InitCond[208];
    m[253] = run?((((m[119]&~m[252]&~m[254]&~m[255]&~m[256])|(~m[119]&~m[252]&~m[254]&m[255]&~m[256])|(m[119]&m[252]&~m[254]&m[255]&~m[256])|(m[119]&~m[252]&m[254]&m[255]&~m[256])|(~m[119]&m[252]&~m[254]&~m[255]&m[256])|(~m[119]&~m[252]&m[254]&~m[255]&m[256])|(m[119]&m[252]&m[254]&~m[255]&m[256])|(~m[119]&m[252]&m[254]&m[255]&m[256]))&UnbiasedRNG[78])|((m[119]&~m[252]&~m[254]&m[255]&~m[256])|(~m[119]&~m[252]&~m[254]&~m[255]&m[256])|(m[119]&~m[252]&~m[254]&~m[255]&m[256])|(m[119]&m[252]&~m[254]&~m[255]&m[256])|(m[119]&~m[252]&m[254]&~m[255]&m[256])|(~m[119]&~m[252]&~m[254]&m[255]&m[256])|(m[119]&~m[252]&~m[254]&m[255]&m[256])|(~m[119]&m[252]&~m[254]&m[255]&m[256])|(m[119]&m[252]&~m[254]&m[255]&m[256])|(~m[119]&~m[252]&m[254]&m[255]&m[256])|(m[119]&~m[252]&m[254]&m[255]&m[256])|(m[119]&m[252]&m[254]&m[255]&m[256]))):InitCond[209];
    m[258] = run?((((m[124]&~m[257]&~m[259]&~m[260]&~m[261])|(~m[124]&~m[257]&~m[259]&m[260]&~m[261])|(m[124]&m[257]&~m[259]&m[260]&~m[261])|(m[124]&~m[257]&m[259]&m[260]&~m[261])|(~m[124]&m[257]&~m[259]&~m[260]&m[261])|(~m[124]&~m[257]&m[259]&~m[260]&m[261])|(m[124]&m[257]&m[259]&~m[260]&m[261])|(~m[124]&m[257]&m[259]&m[260]&m[261]))&UnbiasedRNG[79])|((m[124]&~m[257]&~m[259]&m[260]&~m[261])|(~m[124]&~m[257]&~m[259]&~m[260]&m[261])|(m[124]&~m[257]&~m[259]&~m[260]&m[261])|(m[124]&m[257]&~m[259]&~m[260]&m[261])|(m[124]&~m[257]&m[259]&~m[260]&m[261])|(~m[124]&~m[257]&~m[259]&m[260]&m[261])|(m[124]&~m[257]&~m[259]&m[260]&m[261])|(~m[124]&m[257]&~m[259]&m[260]&m[261])|(m[124]&m[257]&~m[259]&m[260]&m[261])|(~m[124]&~m[257]&m[259]&m[260]&m[261])|(m[124]&~m[257]&m[259]&m[260]&m[261])|(m[124]&m[257]&m[259]&m[260]&m[261]))):InitCond[210];
    m[263] = run?((((m[129]&~m[262]&~m[264]&~m[265]&~m[266])|(~m[129]&~m[262]&~m[264]&m[265]&~m[266])|(m[129]&m[262]&~m[264]&m[265]&~m[266])|(m[129]&~m[262]&m[264]&m[265]&~m[266])|(~m[129]&m[262]&~m[264]&~m[265]&m[266])|(~m[129]&~m[262]&m[264]&~m[265]&m[266])|(m[129]&m[262]&m[264]&~m[265]&m[266])|(~m[129]&m[262]&m[264]&m[265]&m[266]))&UnbiasedRNG[80])|((m[129]&~m[262]&~m[264]&m[265]&~m[266])|(~m[129]&~m[262]&~m[264]&~m[265]&m[266])|(m[129]&~m[262]&~m[264]&~m[265]&m[266])|(m[129]&m[262]&~m[264]&~m[265]&m[266])|(m[129]&~m[262]&m[264]&~m[265]&m[266])|(~m[129]&~m[262]&~m[264]&m[265]&m[266])|(m[129]&~m[262]&~m[264]&m[265]&m[266])|(~m[129]&m[262]&~m[264]&m[265]&m[266])|(m[129]&m[262]&~m[264]&m[265]&m[266])|(~m[129]&~m[262]&m[264]&m[265]&m[266])|(m[129]&~m[262]&m[264]&m[265]&m[266])|(m[129]&m[262]&m[264]&m[265]&m[266]))):InitCond[211];
    m[268] = run?((((m[125]&~m[267]&~m[269]&~m[270]&~m[271])|(~m[125]&~m[267]&~m[269]&m[270]&~m[271])|(m[125]&m[267]&~m[269]&m[270]&~m[271])|(m[125]&~m[267]&m[269]&m[270]&~m[271])|(~m[125]&m[267]&~m[269]&~m[270]&m[271])|(~m[125]&~m[267]&m[269]&~m[270]&m[271])|(m[125]&m[267]&m[269]&~m[270]&m[271])|(~m[125]&m[267]&m[269]&m[270]&m[271]))&UnbiasedRNG[81])|((m[125]&~m[267]&~m[269]&m[270]&~m[271])|(~m[125]&~m[267]&~m[269]&~m[270]&m[271])|(m[125]&~m[267]&~m[269]&~m[270]&m[271])|(m[125]&m[267]&~m[269]&~m[270]&m[271])|(m[125]&~m[267]&m[269]&~m[270]&m[271])|(~m[125]&~m[267]&~m[269]&m[270]&m[271])|(m[125]&~m[267]&~m[269]&m[270]&m[271])|(~m[125]&m[267]&~m[269]&m[270]&m[271])|(m[125]&m[267]&~m[269]&m[270]&m[271])|(~m[125]&~m[267]&m[269]&m[270]&m[271])|(m[125]&~m[267]&m[269]&m[270]&m[271])|(m[125]&m[267]&m[269]&m[270]&m[271]))):InitCond[212];
    m[273] = run?((((m[130]&~m[272]&~m[274]&~m[275]&~m[276])|(~m[130]&~m[272]&~m[274]&m[275]&~m[276])|(m[130]&m[272]&~m[274]&m[275]&~m[276])|(m[130]&~m[272]&m[274]&m[275]&~m[276])|(~m[130]&m[272]&~m[274]&~m[275]&m[276])|(~m[130]&~m[272]&m[274]&~m[275]&m[276])|(m[130]&m[272]&m[274]&~m[275]&m[276])|(~m[130]&m[272]&m[274]&m[275]&m[276]))&UnbiasedRNG[82])|((m[130]&~m[272]&~m[274]&m[275]&~m[276])|(~m[130]&~m[272]&~m[274]&~m[275]&m[276])|(m[130]&~m[272]&~m[274]&~m[275]&m[276])|(m[130]&m[272]&~m[274]&~m[275]&m[276])|(m[130]&~m[272]&m[274]&~m[275]&m[276])|(~m[130]&~m[272]&~m[274]&m[275]&m[276])|(m[130]&~m[272]&~m[274]&m[275]&m[276])|(~m[130]&m[272]&~m[274]&m[275]&m[276])|(m[130]&m[272]&~m[274]&m[275]&m[276])|(~m[130]&~m[272]&m[274]&m[275]&m[276])|(m[130]&~m[272]&m[274]&m[275]&m[276])|(m[130]&m[272]&m[274]&m[275]&m[276]))):InitCond[213];
    m[278] = run?((((m[131]&~m[277]&~m[279]&~m[280]&~m[281])|(~m[131]&~m[277]&~m[279]&m[280]&~m[281])|(m[131]&m[277]&~m[279]&m[280]&~m[281])|(m[131]&~m[277]&m[279]&m[280]&~m[281])|(~m[131]&m[277]&~m[279]&~m[280]&m[281])|(~m[131]&~m[277]&m[279]&~m[280]&m[281])|(m[131]&m[277]&m[279]&~m[280]&m[281])|(~m[131]&m[277]&m[279]&m[280]&m[281]))&UnbiasedRNG[83])|((m[131]&~m[277]&~m[279]&m[280]&~m[281])|(~m[131]&~m[277]&~m[279]&~m[280]&m[281])|(m[131]&~m[277]&~m[279]&~m[280]&m[281])|(m[131]&m[277]&~m[279]&~m[280]&m[281])|(m[131]&~m[277]&m[279]&~m[280]&m[281])|(~m[131]&~m[277]&~m[279]&m[280]&m[281])|(m[131]&~m[277]&~m[279]&m[280]&m[281])|(~m[131]&m[277]&~m[279]&m[280]&m[281])|(m[131]&m[277]&~m[279]&m[280]&m[281])|(~m[131]&~m[277]&m[279]&m[280]&m[281])|(m[131]&~m[277]&m[279]&m[280]&m[281])|(m[131]&m[277]&m[279]&m[280]&m[281]))):InitCond[214];
end

always @(posedge color3_clk) begin
    m[140] = run?((((m[137]&~m[138]&~m[139]&~m[141]&~m[142])|(~m[137]&m[138]&~m[139]&~m[141]&~m[142])|(~m[137]&~m[138]&m[139]&~m[141]&~m[142])|(m[137]&m[138]&m[139]&m[141]&~m[142])|(~m[137]&~m[138]&~m[139]&~m[141]&m[142])|(m[137]&m[138]&~m[139]&m[141]&m[142])|(m[137]&~m[138]&m[139]&m[141]&m[142])|(~m[137]&m[138]&m[139]&m[141]&m[142]))&UnbiasedRNG[84])|((m[137]&m[138]&~m[139]&~m[141]&~m[142])|(m[137]&~m[138]&m[139]&~m[141]&~m[142])|(~m[137]&m[138]&m[139]&~m[141]&~m[142])|(m[137]&m[138]&m[139]&~m[141]&~m[142])|(m[137]&~m[138]&~m[139]&~m[141]&m[142])|(~m[137]&m[138]&~m[139]&~m[141]&m[142])|(m[137]&m[138]&~m[139]&~m[141]&m[142])|(~m[137]&~m[138]&m[139]&~m[141]&m[142])|(m[137]&~m[138]&m[139]&~m[141]&m[142])|(~m[137]&m[138]&m[139]&~m[141]&m[142])|(m[137]&m[138]&m[139]&~m[141]&m[142])|(m[137]&m[138]&m[139]&m[141]&m[142]))):InitCond[215];
    m[150] = run?((((m[147]&~m[148]&~m[149]&~m[151]&~m[152])|(~m[147]&m[148]&~m[149]&~m[151]&~m[152])|(~m[147]&~m[148]&m[149]&~m[151]&~m[152])|(m[147]&m[148]&m[149]&m[151]&~m[152])|(~m[147]&~m[148]&~m[149]&~m[151]&m[152])|(m[147]&m[148]&~m[149]&m[151]&m[152])|(m[147]&~m[148]&m[149]&m[151]&m[152])|(~m[147]&m[148]&m[149]&m[151]&m[152]))&UnbiasedRNG[85])|((m[147]&m[148]&~m[149]&~m[151]&~m[152])|(m[147]&~m[148]&m[149]&~m[151]&~m[152])|(~m[147]&m[148]&m[149]&~m[151]&~m[152])|(m[147]&m[148]&m[149]&~m[151]&~m[152])|(m[147]&~m[148]&~m[149]&~m[151]&m[152])|(~m[147]&m[148]&~m[149]&~m[151]&m[152])|(m[147]&m[148]&~m[149]&~m[151]&m[152])|(~m[147]&~m[148]&m[149]&~m[151]&m[152])|(m[147]&~m[148]&m[149]&~m[151]&m[152])|(~m[147]&m[148]&m[149]&~m[151]&m[152])|(m[147]&m[148]&m[149]&~m[151]&m[152])|(m[147]&m[148]&m[149]&m[151]&m[152]))):InitCond[216];
    m[155] = run?((((m[152]&~m[153]&~m[154]&~m[156]&~m[157])|(~m[152]&m[153]&~m[154]&~m[156]&~m[157])|(~m[152]&~m[153]&m[154]&~m[156]&~m[157])|(m[152]&m[153]&m[154]&m[156]&~m[157])|(~m[152]&~m[153]&~m[154]&~m[156]&m[157])|(m[152]&m[153]&~m[154]&m[156]&m[157])|(m[152]&~m[153]&m[154]&m[156]&m[157])|(~m[152]&m[153]&m[154]&m[156]&m[157]))&UnbiasedRNG[86])|((m[152]&m[153]&~m[154]&~m[156]&~m[157])|(m[152]&~m[153]&m[154]&~m[156]&~m[157])|(~m[152]&m[153]&m[154]&~m[156]&~m[157])|(m[152]&m[153]&m[154]&~m[156]&~m[157])|(m[152]&~m[153]&~m[154]&~m[156]&m[157])|(~m[152]&m[153]&~m[154]&~m[156]&m[157])|(m[152]&m[153]&~m[154]&~m[156]&m[157])|(~m[152]&~m[153]&m[154]&~m[156]&m[157])|(m[152]&~m[153]&m[154]&~m[156]&m[157])|(~m[152]&m[153]&m[154]&~m[156]&m[157])|(m[152]&m[153]&m[154]&~m[156]&m[157])|(m[152]&m[153]&m[154]&m[156]&m[157]))):InitCond[217];
    m[165] = run?((((m[162]&~m[163]&~m[164]&~m[166]&~m[167])|(~m[162]&m[163]&~m[164]&~m[166]&~m[167])|(~m[162]&~m[163]&m[164]&~m[166]&~m[167])|(m[162]&m[163]&m[164]&m[166]&~m[167])|(~m[162]&~m[163]&~m[164]&~m[166]&m[167])|(m[162]&m[163]&~m[164]&m[166]&m[167])|(m[162]&~m[163]&m[164]&m[166]&m[167])|(~m[162]&m[163]&m[164]&m[166]&m[167]))&UnbiasedRNG[87])|((m[162]&m[163]&~m[164]&~m[166]&~m[167])|(m[162]&~m[163]&m[164]&~m[166]&~m[167])|(~m[162]&m[163]&m[164]&~m[166]&~m[167])|(m[162]&m[163]&m[164]&~m[166]&~m[167])|(m[162]&~m[163]&~m[164]&~m[166]&m[167])|(~m[162]&m[163]&~m[164]&~m[166]&m[167])|(m[162]&m[163]&~m[164]&~m[166]&m[167])|(~m[162]&~m[163]&m[164]&~m[166]&m[167])|(m[162]&~m[163]&m[164]&~m[166]&m[167])|(~m[162]&m[163]&m[164]&~m[166]&m[167])|(m[162]&m[163]&m[164]&~m[166]&m[167])|(m[162]&m[163]&m[164]&m[166]&m[167]))):InitCond[218];
    m[170] = run?((((m[167]&~m[168]&~m[169]&~m[171]&~m[172])|(~m[167]&m[168]&~m[169]&~m[171]&~m[172])|(~m[167]&~m[168]&m[169]&~m[171]&~m[172])|(m[167]&m[168]&m[169]&m[171]&~m[172])|(~m[167]&~m[168]&~m[169]&~m[171]&m[172])|(m[167]&m[168]&~m[169]&m[171]&m[172])|(m[167]&~m[168]&m[169]&m[171]&m[172])|(~m[167]&m[168]&m[169]&m[171]&m[172]))&UnbiasedRNG[88])|((m[167]&m[168]&~m[169]&~m[171]&~m[172])|(m[167]&~m[168]&m[169]&~m[171]&~m[172])|(~m[167]&m[168]&m[169]&~m[171]&~m[172])|(m[167]&m[168]&m[169]&~m[171]&~m[172])|(m[167]&~m[168]&~m[169]&~m[171]&m[172])|(~m[167]&m[168]&~m[169]&~m[171]&m[172])|(m[167]&m[168]&~m[169]&~m[171]&m[172])|(~m[167]&~m[168]&m[169]&~m[171]&m[172])|(m[167]&~m[168]&m[169]&~m[171]&m[172])|(~m[167]&m[168]&m[169]&~m[171]&m[172])|(m[167]&m[168]&m[169]&~m[171]&m[172])|(m[167]&m[168]&m[169]&m[171]&m[172]))):InitCond[219];
    m[175] = run?((((m[172]&~m[173]&~m[174]&~m[176]&~m[177])|(~m[172]&m[173]&~m[174]&~m[176]&~m[177])|(~m[172]&~m[173]&m[174]&~m[176]&~m[177])|(m[172]&m[173]&m[174]&m[176]&~m[177])|(~m[172]&~m[173]&~m[174]&~m[176]&m[177])|(m[172]&m[173]&~m[174]&m[176]&m[177])|(m[172]&~m[173]&m[174]&m[176]&m[177])|(~m[172]&m[173]&m[174]&m[176]&m[177]))&UnbiasedRNG[89])|((m[172]&m[173]&~m[174]&~m[176]&~m[177])|(m[172]&~m[173]&m[174]&~m[176]&~m[177])|(~m[172]&m[173]&m[174]&~m[176]&~m[177])|(m[172]&m[173]&m[174]&~m[176]&~m[177])|(m[172]&~m[173]&~m[174]&~m[176]&m[177])|(~m[172]&m[173]&~m[174]&~m[176]&m[177])|(m[172]&m[173]&~m[174]&~m[176]&m[177])|(~m[172]&~m[173]&m[174]&~m[176]&m[177])|(m[172]&~m[173]&m[174]&~m[176]&m[177])|(~m[172]&m[173]&m[174]&~m[176]&m[177])|(m[172]&m[173]&m[174]&~m[176]&m[177])|(m[172]&m[173]&m[174]&m[176]&m[177]))):InitCond[220];
    m[185] = run?((((m[182]&~m[183]&~m[184]&~m[186]&~m[187])|(~m[182]&m[183]&~m[184]&~m[186]&~m[187])|(~m[182]&~m[183]&m[184]&~m[186]&~m[187])|(m[182]&m[183]&m[184]&m[186]&~m[187])|(~m[182]&~m[183]&~m[184]&~m[186]&m[187])|(m[182]&m[183]&~m[184]&m[186]&m[187])|(m[182]&~m[183]&m[184]&m[186]&m[187])|(~m[182]&m[183]&m[184]&m[186]&m[187]))&UnbiasedRNG[90])|((m[182]&m[183]&~m[184]&~m[186]&~m[187])|(m[182]&~m[183]&m[184]&~m[186]&~m[187])|(~m[182]&m[183]&m[184]&~m[186]&~m[187])|(m[182]&m[183]&m[184]&~m[186]&~m[187])|(m[182]&~m[183]&~m[184]&~m[186]&m[187])|(~m[182]&m[183]&~m[184]&~m[186]&m[187])|(m[182]&m[183]&~m[184]&~m[186]&m[187])|(~m[182]&~m[183]&m[184]&~m[186]&m[187])|(m[182]&~m[183]&m[184]&~m[186]&m[187])|(~m[182]&m[183]&m[184]&~m[186]&m[187])|(m[182]&m[183]&m[184]&~m[186]&m[187])|(m[182]&m[183]&m[184]&m[186]&m[187]))):InitCond[221];
    m[190] = run?((((m[187]&~m[188]&~m[189]&~m[191]&~m[192])|(~m[187]&m[188]&~m[189]&~m[191]&~m[192])|(~m[187]&~m[188]&m[189]&~m[191]&~m[192])|(m[187]&m[188]&m[189]&m[191]&~m[192])|(~m[187]&~m[188]&~m[189]&~m[191]&m[192])|(m[187]&m[188]&~m[189]&m[191]&m[192])|(m[187]&~m[188]&m[189]&m[191]&m[192])|(~m[187]&m[188]&m[189]&m[191]&m[192]))&UnbiasedRNG[91])|((m[187]&m[188]&~m[189]&~m[191]&~m[192])|(m[187]&~m[188]&m[189]&~m[191]&~m[192])|(~m[187]&m[188]&m[189]&~m[191]&~m[192])|(m[187]&m[188]&m[189]&~m[191]&~m[192])|(m[187]&~m[188]&~m[189]&~m[191]&m[192])|(~m[187]&m[188]&~m[189]&~m[191]&m[192])|(m[187]&m[188]&~m[189]&~m[191]&m[192])|(~m[187]&~m[188]&m[189]&~m[191]&m[192])|(m[187]&~m[188]&m[189]&~m[191]&m[192])|(~m[187]&m[188]&m[189]&~m[191]&m[192])|(m[187]&m[188]&m[189]&~m[191]&m[192])|(m[187]&m[188]&m[189]&m[191]&m[192]))):InitCond[222];
    m[195] = run?((((m[192]&~m[193]&~m[194]&~m[196]&~m[197])|(~m[192]&m[193]&~m[194]&~m[196]&~m[197])|(~m[192]&~m[193]&m[194]&~m[196]&~m[197])|(m[192]&m[193]&m[194]&m[196]&~m[197])|(~m[192]&~m[193]&~m[194]&~m[196]&m[197])|(m[192]&m[193]&~m[194]&m[196]&m[197])|(m[192]&~m[193]&m[194]&m[196]&m[197])|(~m[192]&m[193]&m[194]&m[196]&m[197]))&UnbiasedRNG[92])|((m[192]&m[193]&~m[194]&~m[196]&~m[197])|(m[192]&~m[193]&m[194]&~m[196]&~m[197])|(~m[192]&m[193]&m[194]&~m[196]&~m[197])|(m[192]&m[193]&m[194]&~m[196]&~m[197])|(m[192]&~m[193]&~m[194]&~m[196]&m[197])|(~m[192]&m[193]&~m[194]&~m[196]&m[197])|(m[192]&m[193]&~m[194]&~m[196]&m[197])|(~m[192]&~m[193]&m[194]&~m[196]&m[197])|(m[192]&~m[193]&m[194]&~m[196]&m[197])|(~m[192]&m[193]&m[194]&~m[196]&m[197])|(m[192]&m[193]&m[194]&~m[196]&m[197])|(m[192]&m[193]&m[194]&m[196]&m[197]))):InitCond[223];
    m[200] = run?((((m[197]&~m[198]&~m[199]&~m[201]&~m[202])|(~m[197]&m[198]&~m[199]&~m[201]&~m[202])|(~m[197]&~m[198]&m[199]&~m[201]&~m[202])|(m[197]&m[198]&m[199]&m[201]&~m[202])|(~m[197]&~m[198]&~m[199]&~m[201]&m[202])|(m[197]&m[198]&~m[199]&m[201]&m[202])|(m[197]&~m[198]&m[199]&m[201]&m[202])|(~m[197]&m[198]&m[199]&m[201]&m[202]))&UnbiasedRNG[93])|((m[197]&m[198]&~m[199]&~m[201]&~m[202])|(m[197]&~m[198]&m[199]&~m[201]&~m[202])|(~m[197]&m[198]&m[199]&~m[201]&~m[202])|(m[197]&m[198]&m[199]&~m[201]&~m[202])|(m[197]&~m[198]&~m[199]&~m[201]&m[202])|(~m[197]&m[198]&~m[199]&~m[201]&m[202])|(m[197]&m[198]&~m[199]&~m[201]&m[202])|(~m[197]&~m[198]&m[199]&~m[201]&m[202])|(m[197]&~m[198]&m[199]&~m[201]&m[202])|(~m[197]&m[198]&m[199]&~m[201]&m[202])|(m[197]&m[198]&m[199]&~m[201]&m[202])|(m[197]&m[198]&m[199]&m[201]&m[202]))):InitCond[224];
    m[210] = run?((((m[207]&~m[208]&~m[209]&~m[211]&~m[212])|(~m[207]&m[208]&~m[209]&~m[211]&~m[212])|(~m[207]&~m[208]&m[209]&~m[211]&~m[212])|(m[207]&m[208]&m[209]&m[211]&~m[212])|(~m[207]&~m[208]&~m[209]&~m[211]&m[212])|(m[207]&m[208]&~m[209]&m[211]&m[212])|(m[207]&~m[208]&m[209]&m[211]&m[212])|(~m[207]&m[208]&m[209]&m[211]&m[212]))&UnbiasedRNG[94])|((m[207]&m[208]&~m[209]&~m[211]&~m[212])|(m[207]&~m[208]&m[209]&~m[211]&~m[212])|(~m[207]&m[208]&m[209]&~m[211]&~m[212])|(m[207]&m[208]&m[209]&~m[211]&~m[212])|(m[207]&~m[208]&~m[209]&~m[211]&m[212])|(~m[207]&m[208]&~m[209]&~m[211]&m[212])|(m[207]&m[208]&~m[209]&~m[211]&m[212])|(~m[207]&~m[208]&m[209]&~m[211]&m[212])|(m[207]&~m[208]&m[209]&~m[211]&m[212])|(~m[207]&m[208]&m[209]&~m[211]&m[212])|(m[207]&m[208]&m[209]&~m[211]&m[212])|(m[207]&m[208]&m[209]&m[211]&m[212]))):InitCond[225];
    m[215] = run?((((m[212]&~m[213]&~m[214]&~m[216]&~m[217])|(~m[212]&m[213]&~m[214]&~m[216]&~m[217])|(~m[212]&~m[213]&m[214]&~m[216]&~m[217])|(m[212]&m[213]&m[214]&m[216]&~m[217])|(~m[212]&~m[213]&~m[214]&~m[216]&m[217])|(m[212]&m[213]&~m[214]&m[216]&m[217])|(m[212]&~m[213]&m[214]&m[216]&m[217])|(~m[212]&m[213]&m[214]&m[216]&m[217]))&UnbiasedRNG[95])|((m[212]&m[213]&~m[214]&~m[216]&~m[217])|(m[212]&~m[213]&m[214]&~m[216]&~m[217])|(~m[212]&m[213]&m[214]&~m[216]&~m[217])|(m[212]&m[213]&m[214]&~m[216]&~m[217])|(m[212]&~m[213]&~m[214]&~m[216]&m[217])|(~m[212]&m[213]&~m[214]&~m[216]&m[217])|(m[212]&m[213]&~m[214]&~m[216]&m[217])|(~m[212]&~m[213]&m[214]&~m[216]&m[217])|(m[212]&~m[213]&m[214]&~m[216]&m[217])|(~m[212]&m[213]&m[214]&~m[216]&m[217])|(m[212]&m[213]&m[214]&~m[216]&m[217])|(m[212]&m[213]&m[214]&m[216]&m[217]))):InitCond[226];
    m[220] = run?((((m[217]&~m[218]&~m[219]&~m[221]&~m[222])|(~m[217]&m[218]&~m[219]&~m[221]&~m[222])|(~m[217]&~m[218]&m[219]&~m[221]&~m[222])|(m[217]&m[218]&m[219]&m[221]&~m[222])|(~m[217]&~m[218]&~m[219]&~m[221]&m[222])|(m[217]&m[218]&~m[219]&m[221]&m[222])|(m[217]&~m[218]&m[219]&m[221]&m[222])|(~m[217]&m[218]&m[219]&m[221]&m[222]))&UnbiasedRNG[96])|((m[217]&m[218]&~m[219]&~m[221]&~m[222])|(m[217]&~m[218]&m[219]&~m[221]&~m[222])|(~m[217]&m[218]&m[219]&~m[221]&~m[222])|(m[217]&m[218]&m[219]&~m[221]&~m[222])|(m[217]&~m[218]&~m[219]&~m[221]&m[222])|(~m[217]&m[218]&~m[219]&~m[221]&m[222])|(m[217]&m[218]&~m[219]&~m[221]&m[222])|(~m[217]&~m[218]&m[219]&~m[221]&m[222])|(m[217]&~m[218]&m[219]&~m[221]&m[222])|(~m[217]&m[218]&m[219]&~m[221]&m[222])|(m[217]&m[218]&m[219]&~m[221]&m[222])|(m[217]&m[218]&m[219]&m[221]&m[222]))):InitCond[227];
    m[225] = run?((((m[222]&~m[223]&~m[224]&~m[226]&~m[227])|(~m[222]&m[223]&~m[224]&~m[226]&~m[227])|(~m[222]&~m[223]&m[224]&~m[226]&~m[227])|(m[222]&m[223]&m[224]&m[226]&~m[227])|(~m[222]&~m[223]&~m[224]&~m[226]&m[227])|(m[222]&m[223]&~m[224]&m[226]&m[227])|(m[222]&~m[223]&m[224]&m[226]&m[227])|(~m[222]&m[223]&m[224]&m[226]&m[227]))&UnbiasedRNG[97])|((m[222]&m[223]&~m[224]&~m[226]&~m[227])|(m[222]&~m[223]&m[224]&~m[226]&~m[227])|(~m[222]&m[223]&m[224]&~m[226]&~m[227])|(m[222]&m[223]&m[224]&~m[226]&~m[227])|(m[222]&~m[223]&~m[224]&~m[226]&m[227])|(~m[222]&m[223]&~m[224]&~m[226]&m[227])|(m[222]&m[223]&~m[224]&~m[226]&m[227])|(~m[222]&~m[223]&m[224]&~m[226]&m[227])|(m[222]&~m[223]&m[224]&~m[226]&m[227])|(~m[222]&m[223]&m[224]&~m[226]&m[227])|(m[222]&m[223]&m[224]&~m[226]&m[227])|(m[222]&m[223]&m[224]&m[226]&m[227]))):InitCond[228];
    m[235] = run?((((m[232]&~m[233]&~m[234]&~m[236]&~m[237])|(~m[232]&m[233]&~m[234]&~m[236]&~m[237])|(~m[232]&~m[233]&m[234]&~m[236]&~m[237])|(m[232]&m[233]&m[234]&m[236]&~m[237])|(~m[232]&~m[233]&~m[234]&~m[236]&m[237])|(m[232]&m[233]&~m[234]&m[236]&m[237])|(m[232]&~m[233]&m[234]&m[236]&m[237])|(~m[232]&m[233]&m[234]&m[236]&m[237]))&UnbiasedRNG[98])|((m[232]&m[233]&~m[234]&~m[236]&~m[237])|(m[232]&~m[233]&m[234]&~m[236]&~m[237])|(~m[232]&m[233]&m[234]&~m[236]&~m[237])|(m[232]&m[233]&m[234]&~m[236]&~m[237])|(m[232]&~m[233]&~m[234]&~m[236]&m[237])|(~m[232]&m[233]&~m[234]&~m[236]&m[237])|(m[232]&m[233]&~m[234]&~m[236]&m[237])|(~m[232]&~m[233]&m[234]&~m[236]&m[237])|(m[232]&~m[233]&m[234]&~m[236]&m[237])|(~m[232]&m[233]&m[234]&~m[236]&m[237])|(m[232]&m[233]&m[234]&~m[236]&m[237])|(m[232]&m[233]&m[234]&m[236]&m[237]))):InitCond[229];
    m[240] = run?((((m[237]&~m[238]&~m[239]&~m[241]&~m[242])|(~m[237]&m[238]&~m[239]&~m[241]&~m[242])|(~m[237]&~m[238]&m[239]&~m[241]&~m[242])|(m[237]&m[238]&m[239]&m[241]&~m[242])|(~m[237]&~m[238]&~m[239]&~m[241]&m[242])|(m[237]&m[238]&~m[239]&m[241]&m[242])|(m[237]&~m[238]&m[239]&m[241]&m[242])|(~m[237]&m[238]&m[239]&m[241]&m[242]))&UnbiasedRNG[99])|((m[237]&m[238]&~m[239]&~m[241]&~m[242])|(m[237]&~m[238]&m[239]&~m[241]&~m[242])|(~m[237]&m[238]&m[239]&~m[241]&~m[242])|(m[237]&m[238]&m[239]&~m[241]&~m[242])|(m[237]&~m[238]&~m[239]&~m[241]&m[242])|(~m[237]&m[238]&~m[239]&~m[241]&m[242])|(m[237]&m[238]&~m[239]&~m[241]&m[242])|(~m[237]&~m[238]&m[239]&~m[241]&m[242])|(m[237]&~m[238]&m[239]&~m[241]&m[242])|(~m[237]&m[238]&m[239]&~m[241]&m[242])|(m[237]&m[238]&m[239]&~m[241]&m[242])|(m[237]&m[238]&m[239]&m[241]&m[242]))):InitCond[230];
    m[245] = run?((((m[242]&~m[243]&~m[244]&~m[246]&~m[247])|(~m[242]&m[243]&~m[244]&~m[246]&~m[247])|(~m[242]&~m[243]&m[244]&~m[246]&~m[247])|(m[242]&m[243]&m[244]&m[246]&~m[247])|(~m[242]&~m[243]&~m[244]&~m[246]&m[247])|(m[242]&m[243]&~m[244]&m[246]&m[247])|(m[242]&~m[243]&m[244]&m[246]&m[247])|(~m[242]&m[243]&m[244]&m[246]&m[247]))&UnbiasedRNG[100])|((m[242]&m[243]&~m[244]&~m[246]&~m[247])|(m[242]&~m[243]&m[244]&~m[246]&~m[247])|(~m[242]&m[243]&m[244]&~m[246]&~m[247])|(m[242]&m[243]&m[244]&~m[246]&~m[247])|(m[242]&~m[243]&~m[244]&~m[246]&m[247])|(~m[242]&m[243]&~m[244]&~m[246]&m[247])|(m[242]&m[243]&~m[244]&~m[246]&m[247])|(~m[242]&~m[243]&m[244]&~m[246]&m[247])|(m[242]&~m[243]&m[244]&~m[246]&m[247])|(~m[242]&m[243]&m[244]&~m[246]&m[247])|(m[242]&m[243]&m[244]&~m[246]&m[247])|(m[242]&m[243]&m[244]&m[246]&m[247]))):InitCond[231];
    m[255] = run?((((m[252]&~m[253]&~m[254]&~m[256]&~m[257])|(~m[252]&m[253]&~m[254]&~m[256]&~m[257])|(~m[252]&~m[253]&m[254]&~m[256]&~m[257])|(m[252]&m[253]&m[254]&m[256]&~m[257])|(~m[252]&~m[253]&~m[254]&~m[256]&m[257])|(m[252]&m[253]&~m[254]&m[256]&m[257])|(m[252]&~m[253]&m[254]&m[256]&m[257])|(~m[252]&m[253]&m[254]&m[256]&m[257]))&UnbiasedRNG[101])|((m[252]&m[253]&~m[254]&~m[256]&~m[257])|(m[252]&~m[253]&m[254]&~m[256]&~m[257])|(~m[252]&m[253]&m[254]&~m[256]&~m[257])|(m[252]&m[253]&m[254]&~m[256]&~m[257])|(m[252]&~m[253]&~m[254]&~m[256]&m[257])|(~m[252]&m[253]&~m[254]&~m[256]&m[257])|(m[252]&m[253]&~m[254]&~m[256]&m[257])|(~m[252]&~m[253]&m[254]&~m[256]&m[257])|(m[252]&~m[253]&m[254]&~m[256]&m[257])|(~m[252]&m[253]&m[254]&~m[256]&m[257])|(m[252]&m[253]&m[254]&~m[256]&m[257])|(m[252]&m[253]&m[254]&m[256]&m[257]))):InitCond[232];
    m[260] = run?((((m[257]&~m[258]&~m[259]&~m[261]&~m[262])|(~m[257]&m[258]&~m[259]&~m[261]&~m[262])|(~m[257]&~m[258]&m[259]&~m[261]&~m[262])|(m[257]&m[258]&m[259]&m[261]&~m[262])|(~m[257]&~m[258]&~m[259]&~m[261]&m[262])|(m[257]&m[258]&~m[259]&m[261]&m[262])|(m[257]&~m[258]&m[259]&m[261]&m[262])|(~m[257]&m[258]&m[259]&m[261]&m[262]))&UnbiasedRNG[102])|((m[257]&m[258]&~m[259]&~m[261]&~m[262])|(m[257]&~m[258]&m[259]&~m[261]&~m[262])|(~m[257]&m[258]&m[259]&~m[261]&~m[262])|(m[257]&m[258]&m[259]&~m[261]&~m[262])|(m[257]&~m[258]&~m[259]&~m[261]&m[262])|(~m[257]&m[258]&~m[259]&~m[261]&m[262])|(m[257]&m[258]&~m[259]&~m[261]&m[262])|(~m[257]&~m[258]&m[259]&~m[261]&m[262])|(m[257]&~m[258]&m[259]&~m[261]&m[262])|(~m[257]&m[258]&m[259]&~m[261]&m[262])|(m[257]&m[258]&m[259]&~m[261]&m[262])|(m[257]&m[258]&m[259]&m[261]&m[262]))):InitCond[233];
    m[270] = run?((((m[267]&~m[268]&~m[269]&~m[271]&~m[272])|(~m[267]&m[268]&~m[269]&~m[271]&~m[272])|(~m[267]&~m[268]&m[269]&~m[271]&~m[272])|(m[267]&m[268]&m[269]&m[271]&~m[272])|(~m[267]&~m[268]&~m[269]&~m[271]&m[272])|(m[267]&m[268]&~m[269]&m[271]&m[272])|(m[267]&~m[268]&m[269]&m[271]&m[272])|(~m[267]&m[268]&m[269]&m[271]&m[272]))&UnbiasedRNG[103])|((m[267]&m[268]&~m[269]&~m[271]&~m[272])|(m[267]&~m[268]&m[269]&~m[271]&~m[272])|(~m[267]&m[268]&m[269]&~m[271]&~m[272])|(m[267]&m[268]&m[269]&~m[271]&~m[272])|(m[267]&~m[268]&~m[269]&~m[271]&m[272])|(~m[267]&m[268]&~m[269]&~m[271]&m[272])|(m[267]&m[268]&~m[269]&~m[271]&m[272])|(~m[267]&~m[268]&m[269]&~m[271]&m[272])|(m[267]&~m[268]&m[269]&~m[271]&m[272])|(~m[267]&m[268]&m[269]&~m[271]&m[272])|(m[267]&m[268]&m[269]&~m[271]&m[272])|(m[267]&m[268]&m[269]&m[271]&m[272]))):InitCond[234];
end

always @(posedge color4_clk) begin
    m[136] = run?((((m[132]&~m[133]&~m[134]&~m[135]&~m[139])|(~m[132]&m[133]&~m[134]&~m[135]&~m[139])|(~m[132]&~m[133]&m[134]&~m[135]&~m[139])|(m[132]&m[133]&~m[134]&m[135]&~m[139])|(m[132]&~m[133]&m[134]&m[135]&~m[139])|(~m[132]&m[133]&m[134]&m[135]&~m[139]))&BiasedRNG[131])|(((m[132]&~m[133]&~m[134]&~m[135]&m[139])|(~m[132]&m[133]&~m[134]&~m[135]&m[139])|(~m[132]&~m[133]&m[134]&~m[135]&m[139])|(m[132]&m[133]&~m[134]&m[135]&m[139])|(m[132]&~m[133]&m[134]&m[135]&m[139])|(~m[132]&m[133]&m[134]&m[135]&m[139]))&~BiasedRNG[131])|((m[132]&m[133]&~m[134]&~m[135]&~m[139])|(m[132]&~m[133]&m[134]&~m[135]&~m[139])|(~m[132]&m[133]&m[134]&~m[135]&~m[139])|(m[132]&m[133]&m[134]&~m[135]&~m[139])|(m[132]&m[133]&m[134]&m[135]&~m[139])|(m[132]&m[133]&~m[134]&~m[135]&m[139])|(m[132]&~m[133]&m[134]&~m[135]&m[139])|(~m[132]&m[133]&m[134]&~m[135]&m[139])|(m[132]&m[133]&m[134]&~m[135]&m[139])|(m[132]&m[133]&m[134]&m[135]&m[139]))):InitCond[235];
    m[141] = run?((((m[137]&~m[138]&~m[139]&~m[140]&~m[149])|(~m[137]&m[138]&~m[139]&~m[140]&~m[149])|(~m[137]&~m[138]&m[139]&~m[140]&~m[149])|(m[137]&m[138]&~m[139]&m[140]&~m[149])|(m[137]&~m[138]&m[139]&m[140]&~m[149])|(~m[137]&m[138]&m[139]&m[140]&~m[149]))&BiasedRNG[132])|(((m[137]&~m[138]&~m[139]&~m[140]&m[149])|(~m[137]&m[138]&~m[139]&~m[140]&m[149])|(~m[137]&~m[138]&m[139]&~m[140]&m[149])|(m[137]&m[138]&~m[139]&m[140]&m[149])|(m[137]&~m[138]&m[139]&m[140]&m[149])|(~m[137]&m[138]&m[139]&m[140]&m[149]))&~BiasedRNG[132])|((m[137]&m[138]&~m[139]&~m[140]&~m[149])|(m[137]&~m[138]&m[139]&~m[140]&~m[149])|(~m[137]&m[138]&m[139]&~m[140]&~m[149])|(m[137]&m[138]&m[139]&~m[140]&~m[149])|(m[137]&m[138]&m[139]&m[140]&~m[149])|(m[137]&m[138]&~m[139]&~m[140]&m[149])|(m[137]&~m[138]&m[139]&~m[140]&m[149])|(~m[137]&m[138]&m[139]&~m[140]&m[149])|(m[137]&m[138]&m[139]&~m[140]&m[149])|(m[137]&m[138]&m[139]&m[140]&m[149]))):InitCond[236];
    m[146] = run?((((m[142]&~m[143]&~m[144]&~m[145]&~m[154])|(~m[142]&m[143]&~m[144]&~m[145]&~m[154])|(~m[142]&~m[143]&m[144]&~m[145]&~m[154])|(m[142]&m[143]&~m[144]&m[145]&~m[154])|(m[142]&~m[143]&m[144]&m[145]&~m[154])|(~m[142]&m[143]&m[144]&m[145]&~m[154]))&BiasedRNG[133])|(((m[142]&~m[143]&~m[144]&~m[145]&m[154])|(~m[142]&m[143]&~m[144]&~m[145]&m[154])|(~m[142]&~m[143]&m[144]&~m[145]&m[154])|(m[142]&m[143]&~m[144]&m[145]&m[154])|(m[142]&~m[143]&m[144]&m[145]&m[154])|(~m[142]&m[143]&m[144]&m[145]&m[154]))&~BiasedRNG[133])|((m[142]&m[143]&~m[144]&~m[145]&~m[154])|(m[142]&~m[143]&m[144]&~m[145]&~m[154])|(~m[142]&m[143]&m[144]&~m[145]&~m[154])|(m[142]&m[143]&m[144]&~m[145]&~m[154])|(m[142]&m[143]&m[144]&m[145]&~m[154])|(m[142]&m[143]&~m[144]&~m[145]&m[154])|(m[142]&~m[143]&m[144]&~m[145]&m[154])|(~m[142]&m[143]&m[144]&~m[145]&m[154])|(m[142]&m[143]&m[144]&~m[145]&m[154])|(m[142]&m[143]&m[144]&m[145]&m[154]))):InitCond[237];
    m[151] = run?((((m[147]&~m[148]&~m[149]&~m[150]&~m[164])|(~m[147]&m[148]&~m[149]&~m[150]&~m[164])|(~m[147]&~m[148]&m[149]&~m[150]&~m[164])|(m[147]&m[148]&~m[149]&m[150]&~m[164])|(m[147]&~m[148]&m[149]&m[150]&~m[164])|(~m[147]&m[148]&m[149]&m[150]&~m[164]))&BiasedRNG[134])|(((m[147]&~m[148]&~m[149]&~m[150]&m[164])|(~m[147]&m[148]&~m[149]&~m[150]&m[164])|(~m[147]&~m[148]&m[149]&~m[150]&m[164])|(m[147]&m[148]&~m[149]&m[150]&m[164])|(m[147]&~m[148]&m[149]&m[150]&m[164])|(~m[147]&m[148]&m[149]&m[150]&m[164]))&~BiasedRNG[134])|((m[147]&m[148]&~m[149]&~m[150]&~m[164])|(m[147]&~m[148]&m[149]&~m[150]&~m[164])|(~m[147]&m[148]&m[149]&~m[150]&~m[164])|(m[147]&m[148]&m[149]&~m[150]&~m[164])|(m[147]&m[148]&m[149]&m[150]&~m[164])|(m[147]&m[148]&~m[149]&~m[150]&m[164])|(m[147]&~m[148]&m[149]&~m[150]&m[164])|(~m[147]&m[148]&m[149]&~m[150]&m[164])|(m[147]&m[148]&m[149]&~m[150]&m[164])|(m[147]&m[148]&m[149]&m[150]&m[164]))):InitCond[238];
    m[156] = run?((((m[152]&~m[153]&~m[154]&~m[155]&~m[169])|(~m[152]&m[153]&~m[154]&~m[155]&~m[169])|(~m[152]&~m[153]&m[154]&~m[155]&~m[169])|(m[152]&m[153]&~m[154]&m[155]&~m[169])|(m[152]&~m[153]&m[154]&m[155]&~m[169])|(~m[152]&m[153]&m[154]&m[155]&~m[169]))&BiasedRNG[135])|(((m[152]&~m[153]&~m[154]&~m[155]&m[169])|(~m[152]&m[153]&~m[154]&~m[155]&m[169])|(~m[152]&~m[153]&m[154]&~m[155]&m[169])|(m[152]&m[153]&~m[154]&m[155]&m[169])|(m[152]&~m[153]&m[154]&m[155]&m[169])|(~m[152]&m[153]&m[154]&m[155]&m[169]))&~BiasedRNG[135])|((m[152]&m[153]&~m[154]&~m[155]&~m[169])|(m[152]&~m[153]&m[154]&~m[155]&~m[169])|(~m[152]&m[153]&m[154]&~m[155]&~m[169])|(m[152]&m[153]&m[154]&~m[155]&~m[169])|(m[152]&m[153]&m[154]&m[155]&~m[169])|(m[152]&m[153]&~m[154]&~m[155]&m[169])|(m[152]&~m[153]&m[154]&~m[155]&m[169])|(~m[152]&m[153]&m[154]&~m[155]&m[169])|(m[152]&m[153]&m[154]&~m[155]&m[169])|(m[152]&m[153]&m[154]&m[155]&m[169]))):InitCond[239];
    m[161] = run?((((m[157]&~m[158]&~m[159]&~m[160]&~m[174])|(~m[157]&m[158]&~m[159]&~m[160]&~m[174])|(~m[157]&~m[158]&m[159]&~m[160]&~m[174])|(m[157]&m[158]&~m[159]&m[160]&~m[174])|(m[157]&~m[158]&m[159]&m[160]&~m[174])|(~m[157]&m[158]&m[159]&m[160]&~m[174]))&BiasedRNG[136])|(((m[157]&~m[158]&~m[159]&~m[160]&m[174])|(~m[157]&m[158]&~m[159]&~m[160]&m[174])|(~m[157]&~m[158]&m[159]&~m[160]&m[174])|(m[157]&m[158]&~m[159]&m[160]&m[174])|(m[157]&~m[158]&m[159]&m[160]&m[174])|(~m[157]&m[158]&m[159]&m[160]&m[174]))&~BiasedRNG[136])|((m[157]&m[158]&~m[159]&~m[160]&~m[174])|(m[157]&~m[158]&m[159]&~m[160]&~m[174])|(~m[157]&m[158]&m[159]&~m[160]&~m[174])|(m[157]&m[158]&m[159]&~m[160]&~m[174])|(m[157]&m[158]&m[159]&m[160]&~m[174])|(m[157]&m[158]&~m[159]&~m[160]&m[174])|(m[157]&~m[158]&m[159]&~m[160]&m[174])|(~m[157]&m[158]&m[159]&~m[160]&m[174])|(m[157]&m[158]&m[159]&~m[160]&m[174])|(m[157]&m[158]&m[159]&m[160]&m[174]))):InitCond[240];
    m[166] = run?((((m[162]&~m[163]&~m[164]&~m[165]&~m[184])|(~m[162]&m[163]&~m[164]&~m[165]&~m[184])|(~m[162]&~m[163]&m[164]&~m[165]&~m[184])|(m[162]&m[163]&~m[164]&m[165]&~m[184])|(m[162]&~m[163]&m[164]&m[165]&~m[184])|(~m[162]&m[163]&m[164]&m[165]&~m[184]))&BiasedRNG[137])|(((m[162]&~m[163]&~m[164]&~m[165]&m[184])|(~m[162]&m[163]&~m[164]&~m[165]&m[184])|(~m[162]&~m[163]&m[164]&~m[165]&m[184])|(m[162]&m[163]&~m[164]&m[165]&m[184])|(m[162]&~m[163]&m[164]&m[165]&m[184])|(~m[162]&m[163]&m[164]&m[165]&m[184]))&~BiasedRNG[137])|((m[162]&m[163]&~m[164]&~m[165]&~m[184])|(m[162]&~m[163]&m[164]&~m[165]&~m[184])|(~m[162]&m[163]&m[164]&~m[165]&~m[184])|(m[162]&m[163]&m[164]&~m[165]&~m[184])|(m[162]&m[163]&m[164]&m[165]&~m[184])|(m[162]&m[163]&~m[164]&~m[165]&m[184])|(m[162]&~m[163]&m[164]&~m[165]&m[184])|(~m[162]&m[163]&m[164]&~m[165]&m[184])|(m[162]&m[163]&m[164]&~m[165]&m[184])|(m[162]&m[163]&m[164]&m[165]&m[184]))):InitCond[241];
    m[171] = run?((((m[167]&~m[168]&~m[169]&~m[170]&~m[189])|(~m[167]&m[168]&~m[169]&~m[170]&~m[189])|(~m[167]&~m[168]&m[169]&~m[170]&~m[189])|(m[167]&m[168]&~m[169]&m[170]&~m[189])|(m[167]&~m[168]&m[169]&m[170]&~m[189])|(~m[167]&m[168]&m[169]&m[170]&~m[189]))&BiasedRNG[138])|(((m[167]&~m[168]&~m[169]&~m[170]&m[189])|(~m[167]&m[168]&~m[169]&~m[170]&m[189])|(~m[167]&~m[168]&m[169]&~m[170]&m[189])|(m[167]&m[168]&~m[169]&m[170]&m[189])|(m[167]&~m[168]&m[169]&m[170]&m[189])|(~m[167]&m[168]&m[169]&m[170]&m[189]))&~BiasedRNG[138])|((m[167]&m[168]&~m[169]&~m[170]&~m[189])|(m[167]&~m[168]&m[169]&~m[170]&~m[189])|(~m[167]&m[168]&m[169]&~m[170]&~m[189])|(m[167]&m[168]&m[169]&~m[170]&~m[189])|(m[167]&m[168]&m[169]&m[170]&~m[189])|(m[167]&m[168]&~m[169]&~m[170]&m[189])|(m[167]&~m[168]&m[169]&~m[170]&m[189])|(~m[167]&m[168]&m[169]&~m[170]&m[189])|(m[167]&m[168]&m[169]&~m[170]&m[189])|(m[167]&m[168]&m[169]&m[170]&m[189]))):InitCond[242];
    m[176] = run?((((m[172]&~m[173]&~m[174]&~m[175]&~m[194])|(~m[172]&m[173]&~m[174]&~m[175]&~m[194])|(~m[172]&~m[173]&m[174]&~m[175]&~m[194])|(m[172]&m[173]&~m[174]&m[175]&~m[194])|(m[172]&~m[173]&m[174]&m[175]&~m[194])|(~m[172]&m[173]&m[174]&m[175]&~m[194]))&BiasedRNG[139])|(((m[172]&~m[173]&~m[174]&~m[175]&m[194])|(~m[172]&m[173]&~m[174]&~m[175]&m[194])|(~m[172]&~m[173]&m[174]&~m[175]&m[194])|(m[172]&m[173]&~m[174]&m[175]&m[194])|(m[172]&~m[173]&m[174]&m[175]&m[194])|(~m[172]&m[173]&m[174]&m[175]&m[194]))&~BiasedRNG[139])|((m[172]&m[173]&~m[174]&~m[175]&~m[194])|(m[172]&~m[173]&m[174]&~m[175]&~m[194])|(~m[172]&m[173]&m[174]&~m[175]&~m[194])|(m[172]&m[173]&m[174]&~m[175]&~m[194])|(m[172]&m[173]&m[174]&m[175]&~m[194])|(m[172]&m[173]&~m[174]&~m[175]&m[194])|(m[172]&~m[173]&m[174]&~m[175]&m[194])|(~m[172]&m[173]&m[174]&~m[175]&m[194])|(m[172]&m[173]&m[174]&~m[175]&m[194])|(m[172]&m[173]&m[174]&m[175]&m[194]))):InitCond[243];
    m[181] = run?((((m[177]&~m[178]&~m[179]&~m[180]&~m[199])|(~m[177]&m[178]&~m[179]&~m[180]&~m[199])|(~m[177]&~m[178]&m[179]&~m[180]&~m[199])|(m[177]&m[178]&~m[179]&m[180]&~m[199])|(m[177]&~m[178]&m[179]&m[180]&~m[199])|(~m[177]&m[178]&m[179]&m[180]&~m[199]))&BiasedRNG[140])|(((m[177]&~m[178]&~m[179]&~m[180]&m[199])|(~m[177]&m[178]&~m[179]&~m[180]&m[199])|(~m[177]&~m[178]&m[179]&~m[180]&m[199])|(m[177]&m[178]&~m[179]&m[180]&m[199])|(m[177]&~m[178]&m[179]&m[180]&m[199])|(~m[177]&m[178]&m[179]&m[180]&m[199]))&~BiasedRNG[140])|((m[177]&m[178]&~m[179]&~m[180]&~m[199])|(m[177]&~m[178]&m[179]&~m[180]&~m[199])|(~m[177]&m[178]&m[179]&~m[180]&~m[199])|(m[177]&m[178]&m[179]&~m[180]&~m[199])|(m[177]&m[178]&m[179]&m[180]&~m[199])|(m[177]&m[178]&~m[179]&~m[180]&m[199])|(m[177]&~m[178]&m[179]&~m[180]&m[199])|(~m[177]&m[178]&m[179]&~m[180]&m[199])|(m[177]&m[178]&m[179]&~m[180]&m[199])|(m[177]&m[178]&m[179]&m[180]&m[199]))):InitCond[244];
    m[186] = run?((((m[182]&~m[183]&~m[184]&~m[185]&~m[209])|(~m[182]&m[183]&~m[184]&~m[185]&~m[209])|(~m[182]&~m[183]&m[184]&~m[185]&~m[209])|(m[182]&m[183]&~m[184]&m[185]&~m[209])|(m[182]&~m[183]&m[184]&m[185]&~m[209])|(~m[182]&m[183]&m[184]&m[185]&~m[209]))&BiasedRNG[141])|(((m[182]&~m[183]&~m[184]&~m[185]&m[209])|(~m[182]&m[183]&~m[184]&~m[185]&m[209])|(~m[182]&~m[183]&m[184]&~m[185]&m[209])|(m[182]&m[183]&~m[184]&m[185]&m[209])|(m[182]&~m[183]&m[184]&m[185]&m[209])|(~m[182]&m[183]&m[184]&m[185]&m[209]))&~BiasedRNG[141])|((m[182]&m[183]&~m[184]&~m[185]&~m[209])|(m[182]&~m[183]&m[184]&~m[185]&~m[209])|(~m[182]&m[183]&m[184]&~m[185]&~m[209])|(m[182]&m[183]&m[184]&~m[185]&~m[209])|(m[182]&m[183]&m[184]&m[185]&~m[209])|(m[182]&m[183]&~m[184]&~m[185]&m[209])|(m[182]&~m[183]&m[184]&~m[185]&m[209])|(~m[182]&m[183]&m[184]&~m[185]&m[209])|(m[182]&m[183]&m[184]&~m[185]&m[209])|(m[182]&m[183]&m[184]&m[185]&m[209]))):InitCond[245];
    m[191] = run?((((m[187]&~m[188]&~m[189]&~m[190]&~m[214])|(~m[187]&m[188]&~m[189]&~m[190]&~m[214])|(~m[187]&~m[188]&m[189]&~m[190]&~m[214])|(m[187]&m[188]&~m[189]&m[190]&~m[214])|(m[187]&~m[188]&m[189]&m[190]&~m[214])|(~m[187]&m[188]&m[189]&m[190]&~m[214]))&BiasedRNG[142])|(((m[187]&~m[188]&~m[189]&~m[190]&m[214])|(~m[187]&m[188]&~m[189]&~m[190]&m[214])|(~m[187]&~m[188]&m[189]&~m[190]&m[214])|(m[187]&m[188]&~m[189]&m[190]&m[214])|(m[187]&~m[188]&m[189]&m[190]&m[214])|(~m[187]&m[188]&m[189]&m[190]&m[214]))&~BiasedRNG[142])|((m[187]&m[188]&~m[189]&~m[190]&~m[214])|(m[187]&~m[188]&m[189]&~m[190]&~m[214])|(~m[187]&m[188]&m[189]&~m[190]&~m[214])|(m[187]&m[188]&m[189]&~m[190]&~m[214])|(m[187]&m[188]&m[189]&m[190]&~m[214])|(m[187]&m[188]&~m[189]&~m[190]&m[214])|(m[187]&~m[188]&m[189]&~m[190]&m[214])|(~m[187]&m[188]&m[189]&~m[190]&m[214])|(m[187]&m[188]&m[189]&~m[190]&m[214])|(m[187]&m[188]&m[189]&m[190]&m[214]))):InitCond[246];
    m[196] = run?((((m[192]&~m[193]&~m[194]&~m[195]&~m[219])|(~m[192]&m[193]&~m[194]&~m[195]&~m[219])|(~m[192]&~m[193]&m[194]&~m[195]&~m[219])|(m[192]&m[193]&~m[194]&m[195]&~m[219])|(m[192]&~m[193]&m[194]&m[195]&~m[219])|(~m[192]&m[193]&m[194]&m[195]&~m[219]))&BiasedRNG[143])|(((m[192]&~m[193]&~m[194]&~m[195]&m[219])|(~m[192]&m[193]&~m[194]&~m[195]&m[219])|(~m[192]&~m[193]&m[194]&~m[195]&m[219])|(m[192]&m[193]&~m[194]&m[195]&m[219])|(m[192]&~m[193]&m[194]&m[195]&m[219])|(~m[192]&m[193]&m[194]&m[195]&m[219]))&~BiasedRNG[143])|((m[192]&m[193]&~m[194]&~m[195]&~m[219])|(m[192]&~m[193]&m[194]&~m[195]&~m[219])|(~m[192]&m[193]&m[194]&~m[195]&~m[219])|(m[192]&m[193]&m[194]&~m[195]&~m[219])|(m[192]&m[193]&m[194]&m[195]&~m[219])|(m[192]&m[193]&~m[194]&~m[195]&m[219])|(m[192]&~m[193]&m[194]&~m[195]&m[219])|(~m[192]&m[193]&m[194]&~m[195]&m[219])|(m[192]&m[193]&m[194]&~m[195]&m[219])|(m[192]&m[193]&m[194]&m[195]&m[219]))):InitCond[247];
    m[201] = run?((((m[197]&~m[198]&~m[199]&~m[200]&~m[224])|(~m[197]&m[198]&~m[199]&~m[200]&~m[224])|(~m[197]&~m[198]&m[199]&~m[200]&~m[224])|(m[197]&m[198]&~m[199]&m[200]&~m[224])|(m[197]&~m[198]&m[199]&m[200]&~m[224])|(~m[197]&m[198]&m[199]&m[200]&~m[224]))&BiasedRNG[144])|(((m[197]&~m[198]&~m[199]&~m[200]&m[224])|(~m[197]&m[198]&~m[199]&~m[200]&m[224])|(~m[197]&~m[198]&m[199]&~m[200]&m[224])|(m[197]&m[198]&~m[199]&m[200]&m[224])|(m[197]&~m[198]&m[199]&m[200]&m[224])|(~m[197]&m[198]&m[199]&m[200]&m[224]))&~BiasedRNG[144])|((m[197]&m[198]&~m[199]&~m[200]&~m[224])|(m[197]&~m[198]&m[199]&~m[200]&~m[224])|(~m[197]&m[198]&m[199]&~m[200]&~m[224])|(m[197]&m[198]&m[199]&~m[200]&~m[224])|(m[197]&m[198]&m[199]&m[200]&~m[224])|(m[197]&m[198]&~m[199]&~m[200]&m[224])|(m[197]&~m[198]&m[199]&~m[200]&m[224])|(~m[197]&m[198]&m[199]&~m[200]&m[224])|(m[197]&m[198]&m[199]&~m[200]&m[224])|(m[197]&m[198]&m[199]&m[200]&m[224]))):InitCond[248];
    m[206] = run?((((m[202]&~m[203]&~m[204]&~m[205]&~m[229])|(~m[202]&m[203]&~m[204]&~m[205]&~m[229])|(~m[202]&~m[203]&m[204]&~m[205]&~m[229])|(m[202]&m[203]&~m[204]&m[205]&~m[229])|(m[202]&~m[203]&m[204]&m[205]&~m[229])|(~m[202]&m[203]&m[204]&m[205]&~m[229]))&BiasedRNG[145])|(((m[202]&~m[203]&~m[204]&~m[205]&m[229])|(~m[202]&m[203]&~m[204]&~m[205]&m[229])|(~m[202]&~m[203]&m[204]&~m[205]&m[229])|(m[202]&m[203]&~m[204]&m[205]&m[229])|(m[202]&~m[203]&m[204]&m[205]&m[229])|(~m[202]&m[203]&m[204]&m[205]&m[229]))&~BiasedRNG[145])|((m[202]&m[203]&~m[204]&~m[205]&~m[229])|(m[202]&~m[203]&m[204]&~m[205]&~m[229])|(~m[202]&m[203]&m[204]&~m[205]&~m[229])|(m[202]&m[203]&m[204]&~m[205]&~m[229])|(m[202]&m[203]&m[204]&m[205]&~m[229])|(m[202]&m[203]&~m[204]&~m[205]&m[229])|(m[202]&~m[203]&m[204]&~m[205]&m[229])|(~m[202]&m[203]&m[204]&~m[205]&m[229])|(m[202]&m[203]&m[204]&~m[205]&m[229])|(m[202]&m[203]&m[204]&m[205]&m[229]))):InitCond[249];
    m[211] = run?((((m[207]&~m[208]&~m[209]&~m[210]&~m[232])|(~m[207]&m[208]&~m[209]&~m[210]&~m[232])|(~m[207]&~m[208]&m[209]&~m[210]&~m[232])|(m[207]&m[208]&~m[209]&m[210]&~m[232])|(m[207]&~m[208]&m[209]&m[210]&~m[232])|(~m[207]&m[208]&m[209]&m[210]&~m[232]))&BiasedRNG[146])|(((m[207]&~m[208]&~m[209]&~m[210]&m[232])|(~m[207]&m[208]&~m[209]&~m[210]&m[232])|(~m[207]&~m[208]&m[209]&~m[210]&m[232])|(m[207]&m[208]&~m[209]&m[210]&m[232])|(m[207]&~m[208]&m[209]&m[210]&m[232])|(~m[207]&m[208]&m[209]&m[210]&m[232]))&~BiasedRNG[146])|((m[207]&m[208]&~m[209]&~m[210]&~m[232])|(m[207]&~m[208]&m[209]&~m[210]&~m[232])|(~m[207]&m[208]&m[209]&~m[210]&~m[232])|(m[207]&m[208]&m[209]&~m[210]&~m[232])|(m[207]&m[208]&m[209]&m[210]&~m[232])|(m[207]&m[208]&~m[209]&~m[210]&m[232])|(m[207]&~m[208]&m[209]&~m[210]&m[232])|(~m[207]&m[208]&m[209]&~m[210]&m[232])|(m[207]&m[208]&m[209]&~m[210]&m[232])|(m[207]&m[208]&m[209]&m[210]&m[232]))):InitCond[250];
    m[216] = run?((((m[212]&~m[213]&~m[214]&~m[215]&~m[234])|(~m[212]&m[213]&~m[214]&~m[215]&~m[234])|(~m[212]&~m[213]&m[214]&~m[215]&~m[234])|(m[212]&m[213]&~m[214]&m[215]&~m[234])|(m[212]&~m[213]&m[214]&m[215]&~m[234])|(~m[212]&m[213]&m[214]&m[215]&~m[234]))&BiasedRNG[147])|(((m[212]&~m[213]&~m[214]&~m[215]&m[234])|(~m[212]&m[213]&~m[214]&~m[215]&m[234])|(~m[212]&~m[213]&m[214]&~m[215]&m[234])|(m[212]&m[213]&~m[214]&m[215]&m[234])|(m[212]&~m[213]&m[214]&m[215]&m[234])|(~m[212]&m[213]&m[214]&m[215]&m[234]))&~BiasedRNG[147])|((m[212]&m[213]&~m[214]&~m[215]&~m[234])|(m[212]&~m[213]&m[214]&~m[215]&~m[234])|(~m[212]&m[213]&m[214]&~m[215]&~m[234])|(m[212]&m[213]&m[214]&~m[215]&~m[234])|(m[212]&m[213]&m[214]&m[215]&~m[234])|(m[212]&m[213]&~m[214]&~m[215]&m[234])|(m[212]&~m[213]&m[214]&~m[215]&m[234])|(~m[212]&m[213]&m[214]&~m[215]&m[234])|(m[212]&m[213]&m[214]&~m[215]&m[234])|(m[212]&m[213]&m[214]&m[215]&m[234]))):InitCond[251];
    m[221] = run?((((m[217]&~m[218]&~m[219]&~m[220]&~m[239])|(~m[217]&m[218]&~m[219]&~m[220]&~m[239])|(~m[217]&~m[218]&m[219]&~m[220]&~m[239])|(m[217]&m[218]&~m[219]&m[220]&~m[239])|(m[217]&~m[218]&m[219]&m[220]&~m[239])|(~m[217]&m[218]&m[219]&m[220]&~m[239]))&BiasedRNG[148])|(((m[217]&~m[218]&~m[219]&~m[220]&m[239])|(~m[217]&m[218]&~m[219]&~m[220]&m[239])|(~m[217]&~m[218]&m[219]&~m[220]&m[239])|(m[217]&m[218]&~m[219]&m[220]&m[239])|(m[217]&~m[218]&m[219]&m[220]&m[239])|(~m[217]&m[218]&m[219]&m[220]&m[239]))&~BiasedRNG[148])|((m[217]&m[218]&~m[219]&~m[220]&~m[239])|(m[217]&~m[218]&m[219]&~m[220]&~m[239])|(~m[217]&m[218]&m[219]&~m[220]&~m[239])|(m[217]&m[218]&m[219]&~m[220]&~m[239])|(m[217]&m[218]&m[219]&m[220]&~m[239])|(m[217]&m[218]&~m[219]&~m[220]&m[239])|(m[217]&~m[218]&m[219]&~m[220]&m[239])|(~m[217]&m[218]&m[219]&~m[220]&m[239])|(m[217]&m[218]&m[219]&~m[220]&m[239])|(m[217]&m[218]&m[219]&m[220]&m[239]))):InitCond[252];
    m[226] = run?((((m[222]&~m[223]&~m[224]&~m[225]&~m[244])|(~m[222]&m[223]&~m[224]&~m[225]&~m[244])|(~m[222]&~m[223]&m[224]&~m[225]&~m[244])|(m[222]&m[223]&~m[224]&m[225]&~m[244])|(m[222]&~m[223]&m[224]&m[225]&~m[244])|(~m[222]&m[223]&m[224]&m[225]&~m[244]))&BiasedRNG[149])|(((m[222]&~m[223]&~m[224]&~m[225]&m[244])|(~m[222]&m[223]&~m[224]&~m[225]&m[244])|(~m[222]&~m[223]&m[224]&~m[225]&m[244])|(m[222]&m[223]&~m[224]&m[225]&m[244])|(m[222]&~m[223]&m[224]&m[225]&m[244])|(~m[222]&m[223]&m[224]&m[225]&m[244]))&~BiasedRNG[149])|((m[222]&m[223]&~m[224]&~m[225]&~m[244])|(m[222]&~m[223]&m[224]&~m[225]&~m[244])|(~m[222]&m[223]&m[224]&~m[225]&~m[244])|(m[222]&m[223]&m[224]&~m[225]&~m[244])|(m[222]&m[223]&m[224]&m[225]&~m[244])|(m[222]&m[223]&~m[224]&~m[225]&m[244])|(m[222]&~m[223]&m[224]&~m[225]&m[244])|(~m[222]&m[223]&m[224]&~m[225]&m[244])|(m[222]&m[223]&m[224]&~m[225]&m[244])|(m[222]&m[223]&m[224]&m[225]&m[244]))):InitCond[253];
    m[231] = run?((((m[227]&~m[228]&~m[229]&~m[230]&~m[249])|(~m[227]&m[228]&~m[229]&~m[230]&~m[249])|(~m[227]&~m[228]&m[229]&~m[230]&~m[249])|(m[227]&m[228]&~m[229]&m[230]&~m[249])|(m[227]&~m[228]&m[229]&m[230]&~m[249])|(~m[227]&m[228]&m[229]&m[230]&~m[249]))&BiasedRNG[150])|(((m[227]&~m[228]&~m[229]&~m[230]&m[249])|(~m[227]&m[228]&~m[229]&~m[230]&m[249])|(~m[227]&~m[228]&m[229]&~m[230]&m[249])|(m[227]&m[228]&~m[229]&m[230]&m[249])|(m[227]&~m[228]&m[229]&m[230]&m[249])|(~m[227]&m[228]&m[229]&m[230]&m[249]))&~BiasedRNG[150])|((m[227]&m[228]&~m[229]&~m[230]&~m[249])|(m[227]&~m[228]&m[229]&~m[230]&~m[249])|(~m[227]&m[228]&m[229]&~m[230]&~m[249])|(m[227]&m[228]&m[229]&~m[230]&~m[249])|(m[227]&m[228]&m[229]&m[230]&~m[249])|(m[227]&m[228]&~m[229]&~m[230]&m[249])|(m[227]&~m[228]&m[229]&~m[230]&m[249])|(~m[227]&m[228]&m[229]&~m[230]&m[249])|(m[227]&m[228]&m[229]&~m[230]&m[249])|(m[227]&m[228]&m[229]&m[230]&m[249]))):InitCond[254];
    m[236] = run?((((m[232]&~m[233]&~m[234]&~m[235]&~m[252])|(~m[232]&m[233]&~m[234]&~m[235]&~m[252])|(~m[232]&~m[233]&m[234]&~m[235]&~m[252])|(m[232]&m[233]&~m[234]&m[235]&~m[252])|(m[232]&~m[233]&m[234]&m[235]&~m[252])|(~m[232]&m[233]&m[234]&m[235]&~m[252]))&BiasedRNG[151])|(((m[232]&~m[233]&~m[234]&~m[235]&m[252])|(~m[232]&m[233]&~m[234]&~m[235]&m[252])|(~m[232]&~m[233]&m[234]&~m[235]&m[252])|(m[232]&m[233]&~m[234]&m[235]&m[252])|(m[232]&~m[233]&m[234]&m[235]&m[252])|(~m[232]&m[233]&m[234]&m[235]&m[252]))&~BiasedRNG[151])|((m[232]&m[233]&~m[234]&~m[235]&~m[252])|(m[232]&~m[233]&m[234]&~m[235]&~m[252])|(~m[232]&m[233]&m[234]&~m[235]&~m[252])|(m[232]&m[233]&m[234]&~m[235]&~m[252])|(m[232]&m[233]&m[234]&m[235]&~m[252])|(m[232]&m[233]&~m[234]&~m[235]&m[252])|(m[232]&~m[233]&m[234]&~m[235]&m[252])|(~m[232]&m[233]&m[234]&~m[235]&m[252])|(m[232]&m[233]&m[234]&~m[235]&m[252])|(m[232]&m[233]&m[234]&m[235]&m[252]))):InitCond[255];
    m[241] = run?((((m[237]&~m[238]&~m[239]&~m[240]&~m[254])|(~m[237]&m[238]&~m[239]&~m[240]&~m[254])|(~m[237]&~m[238]&m[239]&~m[240]&~m[254])|(m[237]&m[238]&~m[239]&m[240]&~m[254])|(m[237]&~m[238]&m[239]&m[240]&~m[254])|(~m[237]&m[238]&m[239]&m[240]&~m[254]))&BiasedRNG[152])|(((m[237]&~m[238]&~m[239]&~m[240]&m[254])|(~m[237]&m[238]&~m[239]&~m[240]&m[254])|(~m[237]&~m[238]&m[239]&~m[240]&m[254])|(m[237]&m[238]&~m[239]&m[240]&m[254])|(m[237]&~m[238]&m[239]&m[240]&m[254])|(~m[237]&m[238]&m[239]&m[240]&m[254]))&~BiasedRNG[152])|((m[237]&m[238]&~m[239]&~m[240]&~m[254])|(m[237]&~m[238]&m[239]&~m[240]&~m[254])|(~m[237]&m[238]&m[239]&~m[240]&~m[254])|(m[237]&m[238]&m[239]&~m[240]&~m[254])|(m[237]&m[238]&m[239]&m[240]&~m[254])|(m[237]&m[238]&~m[239]&~m[240]&m[254])|(m[237]&~m[238]&m[239]&~m[240]&m[254])|(~m[237]&m[238]&m[239]&~m[240]&m[254])|(m[237]&m[238]&m[239]&~m[240]&m[254])|(m[237]&m[238]&m[239]&m[240]&m[254]))):InitCond[256];
    m[246] = run?((((m[242]&~m[243]&~m[244]&~m[245]&~m[259])|(~m[242]&m[243]&~m[244]&~m[245]&~m[259])|(~m[242]&~m[243]&m[244]&~m[245]&~m[259])|(m[242]&m[243]&~m[244]&m[245]&~m[259])|(m[242]&~m[243]&m[244]&m[245]&~m[259])|(~m[242]&m[243]&m[244]&m[245]&~m[259]))&BiasedRNG[153])|(((m[242]&~m[243]&~m[244]&~m[245]&m[259])|(~m[242]&m[243]&~m[244]&~m[245]&m[259])|(~m[242]&~m[243]&m[244]&~m[245]&m[259])|(m[242]&m[243]&~m[244]&m[245]&m[259])|(m[242]&~m[243]&m[244]&m[245]&m[259])|(~m[242]&m[243]&m[244]&m[245]&m[259]))&~BiasedRNG[153])|((m[242]&m[243]&~m[244]&~m[245]&~m[259])|(m[242]&~m[243]&m[244]&~m[245]&~m[259])|(~m[242]&m[243]&m[244]&~m[245]&~m[259])|(m[242]&m[243]&m[244]&~m[245]&~m[259])|(m[242]&m[243]&m[244]&m[245]&~m[259])|(m[242]&m[243]&~m[244]&~m[245]&m[259])|(m[242]&~m[243]&m[244]&~m[245]&m[259])|(~m[242]&m[243]&m[244]&~m[245]&m[259])|(m[242]&m[243]&m[244]&~m[245]&m[259])|(m[242]&m[243]&m[244]&m[245]&m[259]))):InitCond[257];
    m[251] = run?((((m[247]&~m[248]&~m[249]&~m[250]&~m[264])|(~m[247]&m[248]&~m[249]&~m[250]&~m[264])|(~m[247]&~m[248]&m[249]&~m[250]&~m[264])|(m[247]&m[248]&~m[249]&m[250]&~m[264])|(m[247]&~m[248]&m[249]&m[250]&~m[264])|(~m[247]&m[248]&m[249]&m[250]&~m[264]))&BiasedRNG[154])|(((m[247]&~m[248]&~m[249]&~m[250]&m[264])|(~m[247]&m[248]&~m[249]&~m[250]&m[264])|(~m[247]&~m[248]&m[249]&~m[250]&m[264])|(m[247]&m[248]&~m[249]&m[250]&m[264])|(m[247]&~m[248]&m[249]&m[250]&m[264])|(~m[247]&m[248]&m[249]&m[250]&m[264]))&~BiasedRNG[154])|((m[247]&m[248]&~m[249]&~m[250]&~m[264])|(m[247]&~m[248]&m[249]&~m[250]&~m[264])|(~m[247]&m[248]&m[249]&~m[250]&~m[264])|(m[247]&m[248]&m[249]&~m[250]&~m[264])|(m[247]&m[248]&m[249]&m[250]&~m[264])|(m[247]&m[248]&~m[249]&~m[250]&m[264])|(m[247]&~m[248]&m[249]&~m[250]&m[264])|(~m[247]&m[248]&m[249]&~m[250]&m[264])|(m[247]&m[248]&m[249]&~m[250]&m[264])|(m[247]&m[248]&m[249]&m[250]&m[264]))):InitCond[258];
    m[256] = run?((((m[252]&~m[253]&~m[254]&~m[255]&~m[267])|(~m[252]&m[253]&~m[254]&~m[255]&~m[267])|(~m[252]&~m[253]&m[254]&~m[255]&~m[267])|(m[252]&m[253]&~m[254]&m[255]&~m[267])|(m[252]&~m[253]&m[254]&m[255]&~m[267])|(~m[252]&m[253]&m[254]&m[255]&~m[267]))&BiasedRNG[155])|(((m[252]&~m[253]&~m[254]&~m[255]&m[267])|(~m[252]&m[253]&~m[254]&~m[255]&m[267])|(~m[252]&~m[253]&m[254]&~m[255]&m[267])|(m[252]&m[253]&~m[254]&m[255]&m[267])|(m[252]&~m[253]&m[254]&m[255]&m[267])|(~m[252]&m[253]&m[254]&m[255]&m[267]))&~BiasedRNG[155])|((m[252]&m[253]&~m[254]&~m[255]&~m[267])|(m[252]&~m[253]&m[254]&~m[255]&~m[267])|(~m[252]&m[253]&m[254]&~m[255]&~m[267])|(m[252]&m[253]&m[254]&~m[255]&~m[267])|(m[252]&m[253]&m[254]&m[255]&~m[267])|(m[252]&m[253]&~m[254]&~m[255]&m[267])|(m[252]&~m[253]&m[254]&~m[255]&m[267])|(~m[252]&m[253]&m[254]&~m[255]&m[267])|(m[252]&m[253]&m[254]&~m[255]&m[267])|(m[252]&m[253]&m[254]&m[255]&m[267]))):InitCond[259];
    m[261] = run?((((m[257]&~m[258]&~m[259]&~m[260]&~m[269])|(~m[257]&m[258]&~m[259]&~m[260]&~m[269])|(~m[257]&~m[258]&m[259]&~m[260]&~m[269])|(m[257]&m[258]&~m[259]&m[260]&~m[269])|(m[257]&~m[258]&m[259]&m[260]&~m[269])|(~m[257]&m[258]&m[259]&m[260]&~m[269]))&BiasedRNG[156])|(((m[257]&~m[258]&~m[259]&~m[260]&m[269])|(~m[257]&m[258]&~m[259]&~m[260]&m[269])|(~m[257]&~m[258]&m[259]&~m[260]&m[269])|(m[257]&m[258]&~m[259]&m[260]&m[269])|(m[257]&~m[258]&m[259]&m[260]&m[269])|(~m[257]&m[258]&m[259]&m[260]&m[269]))&~BiasedRNG[156])|((m[257]&m[258]&~m[259]&~m[260]&~m[269])|(m[257]&~m[258]&m[259]&~m[260]&~m[269])|(~m[257]&m[258]&m[259]&~m[260]&~m[269])|(m[257]&m[258]&m[259]&~m[260]&~m[269])|(m[257]&m[258]&m[259]&m[260]&~m[269])|(m[257]&m[258]&~m[259]&~m[260]&m[269])|(m[257]&~m[258]&m[259]&~m[260]&m[269])|(~m[257]&m[258]&m[259]&~m[260]&m[269])|(m[257]&m[258]&m[259]&~m[260]&m[269])|(m[257]&m[258]&m[259]&m[260]&m[269]))):InitCond[260];
    m[266] = run?((((m[262]&~m[263]&~m[264]&~m[265]&~m[274])|(~m[262]&m[263]&~m[264]&~m[265]&~m[274])|(~m[262]&~m[263]&m[264]&~m[265]&~m[274])|(m[262]&m[263]&~m[264]&m[265]&~m[274])|(m[262]&~m[263]&m[264]&m[265]&~m[274])|(~m[262]&m[263]&m[264]&m[265]&~m[274]))&BiasedRNG[157])|(((m[262]&~m[263]&~m[264]&~m[265]&m[274])|(~m[262]&m[263]&~m[264]&~m[265]&m[274])|(~m[262]&~m[263]&m[264]&~m[265]&m[274])|(m[262]&m[263]&~m[264]&m[265]&m[274])|(m[262]&~m[263]&m[264]&m[265]&m[274])|(~m[262]&m[263]&m[264]&m[265]&m[274]))&~BiasedRNG[157])|((m[262]&m[263]&~m[264]&~m[265]&~m[274])|(m[262]&~m[263]&m[264]&~m[265]&~m[274])|(~m[262]&m[263]&m[264]&~m[265]&~m[274])|(m[262]&m[263]&m[264]&~m[265]&~m[274])|(m[262]&m[263]&m[264]&m[265]&~m[274])|(m[262]&m[263]&~m[264]&~m[265]&m[274])|(m[262]&~m[263]&m[264]&~m[265]&m[274])|(~m[262]&m[263]&m[264]&~m[265]&m[274])|(m[262]&m[263]&m[264]&~m[265]&m[274])|(m[262]&m[263]&m[264]&m[265]&m[274]))):InitCond[261];
    m[271] = run?((((m[267]&~m[268]&~m[269]&~m[270]&~m[277])|(~m[267]&m[268]&~m[269]&~m[270]&~m[277])|(~m[267]&~m[268]&m[269]&~m[270]&~m[277])|(m[267]&m[268]&~m[269]&m[270]&~m[277])|(m[267]&~m[268]&m[269]&m[270]&~m[277])|(~m[267]&m[268]&m[269]&m[270]&~m[277]))&BiasedRNG[158])|(((m[267]&~m[268]&~m[269]&~m[270]&m[277])|(~m[267]&m[268]&~m[269]&~m[270]&m[277])|(~m[267]&~m[268]&m[269]&~m[270]&m[277])|(m[267]&m[268]&~m[269]&m[270]&m[277])|(m[267]&~m[268]&m[269]&m[270]&m[277])|(~m[267]&m[268]&m[269]&m[270]&m[277]))&~BiasedRNG[158])|((m[267]&m[268]&~m[269]&~m[270]&~m[277])|(m[267]&~m[268]&m[269]&~m[270]&~m[277])|(~m[267]&m[268]&m[269]&~m[270]&~m[277])|(m[267]&m[268]&m[269]&~m[270]&~m[277])|(m[267]&m[268]&m[269]&m[270]&~m[277])|(m[267]&m[268]&~m[269]&~m[270]&m[277])|(m[267]&~m[268]&m[269]&~m[270]&m[277])|(~m[267]&m[268]&m[269]&~m[270]&m[277])|(m[267]&m[268]&m[269]&~m[270]&m[277])|(m[267]&m[268]&m[269]&m[270]&m[277]))):InitCond[262];
    m[276] = run?((((m[272]&~m[273]&~m[274]&~m[275]&~m[279])|(~m[272]&m[273]&~m[274]&~m[275]&~m[279])|(~m[272]&~m[273]&m[274]&~m[275]&~m[279])|(m[272]&m[273]&~m[274]&m[275]&~m[279])|(m[272]&~m[273]&m[274]&m[275]&~m[279])|(~m[272]&m[273]&m[274]&m[275]&~m[279]))&BiasedRNG[159])|(((m[272]&~m[273]&~m[274]&~m[275]&m[279])|(~m[272]&m[273]&~m[274]&~m[275]&m[279])|(~m[272]&~m[273]&m[274]&~m[275]&m[279])|(m[272]&m[273]&~m[274]&m[275]&m[279])|(m[272]&~m[273]&m[274]&m[275]&m[279])|(~m[272]&m[273]&m[274]&m[275]&m[279]))&~BiasedRNG[159])|((m[272]&m[273]&~m[274]&~m[275]&~m[279])|(m[272]&~m[273]&m[274]&~m[275]&~m[279])|(~m[272]&m[273]&m[274]&~m[275]&~m[279])|(m[272]&m[273]&m[274]&~m[275]&~m[279])|(m[272]&m[273]&m[274]&m[275]&~m[279])|(m[272]&m[273]&~m[274]&~m[275]&m[279])|(m[272]&~m[273]&m[274]&~m[275]&m[279])|(~m[272]&m[273]&m[274]&~m[275]&m[279])|(m[272]&m[273]&m[274]&~m[275]&m[279])|(m[272]&m[273]&m[274]&m[275]&m[279]))):InitCond[263];
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[53]&LFSRcolor0[100]&LFSRcolor0[77]);
    BiasedRNG[1] = (LFSRcolor0[31]&LFSRcolor0[122]&LFSRcolor0[166]);
    BiasedRNG[2] = (LFSRcolor0[155]&LFSRcolor0[99]&LFSRcolor0[149]);
    BiasedRNG[3] = (LFSRcolor0[164]&LFSRcolor0[38]&LFSRcolor0[57]);
    BiasedRNG[4] = (LFSRcolor0[124]&LFSRcolor0[109]&LFSRcolor0[64]);
    BiasedRNG[5] = (LFSRcolor0[24]&LFSRcolor0[0]&LFSRcolor0[146]);
    BiasedRNG[6] = (LFSRcolor0[28]&LFSRcolor0[2]&LFSRcolor0[44]);
    BiasedRNG[7] = (LFSRcolor0[18]&LFSRcolor0[13]&LFSRcolor0[39]);
    BiasedRNG[8] = (LFSRcolor0[62]&LFSRcolor0[79]&LFSRcolor0[95]);
    BiasedRNG[9] = (LFSRcolor0[176]&LFSRcolor0[97]&LFSRcolor0[129]);
    BiasedRNG[10] = (LFSRcolor0[86]&LFSRcolor0[16]&LFSRcolor0[119]);
    BiasedRNG[11] = (LFSRcolor0[171]&LFSRcolor0[51]&LFSRcolor0[96]);
    BiasedRNG[12] = (LFSRcolor0[85]&LFSRcolor0[174]&LFSRcolor0[118]);
    BiasedRNG[13] = (LFSRcolor0[66]&LFSRcolor0[65]&LFSRcolor0[144]);
    BiasedRNG[14] = (LFSRcolor0[89]&LFSRcolor0[87]&LFSRcolor0[145]);
    BiasedRNG[15] = (LFSRcolor0[121]&LFSRcolor0[148]&LFSRcolor0[158]);
    BiasedRNG[16] = (LFSRcolor0[17]&LFSRcolor0[167]&LFSRcolor0[91]);
    BiasedRNG[17] = (LFSRcolor0[134]&LFSRcolor0[59]&LFSRcolor0[54]);
    BiasedRNG[18] = (LFSRcolor0[177]&LFSRcolor0[151]&LFSRcolor0[1]);
    BiasedRNG[19] = (LFSRcolor0[6]&LFSRcolor0[47]&LFSRcolor0[94]);
    BiasedRNG[20] = (LFSRcolor0[180]&LFSRcolor0[142]&LFSRcolor0[169]);
    BiasedRNG[21] = (LFSRcolor0[36]&LFSRcolor0[74]&LFSRcolor0[9]);
    BiasedRNG[22] = (LFSRcolor0[153]&LFSRcolor0[114]&LFSRcolor0[12]);
    BiasedRNG[23] = (LFSRcolor0[7]&LFSRcolor0[123]&LFSRcolor0[73]);
    BiasedRNG[24] = (LFSRcolor0[20]&LFSRcolor0[137]&LFSRcolor0[108]);
    BiasedRNG[25] = (LFSRcolor0[19]&LFSRcolor0[175]&LFSRcolor0[162]);
    BiasedRNG[26] = (LFSRcolor0[130]&LFSRcolor0[93]&LFSRcolor0[15]);
    BiasedRNG[27] = (LFSRcolor0[56]&LFSRcolor0[181]&LFSRcolor0[140]);
    BiasedRNG[28] = (LFSRcolor0[112]&LFSRcolor0[34]&LFSRcolor0[23]);
    BiasedRNG[29] = (LFSRcolor0[107]&LFSRcolor0[90]&LFSRcolor0[159]);
    BiasedRNG[30] = (LFSRcolor0[165]&LFSRcolor0[22]&LFSRcolor0[37]);
    BiasedRNG[31] = (LFSRcolor0[69]&LFSRcolor0[29]&LFSRcolor0[21]);
    BiasedRNG[32] = (LFSRcolor0[43]&LFSRcolor0[150]&LFSRcolor0[32]);
    BiasedRNG[33] = (LFSRcolor0[116]&LFSRcolor0[179]&LFSRcolor0[52]);
    BiasedRNG[34] = (LFSRcolor0[117]&LFSRcolor0[42]&LFSRcolor0[84]);
    BiasedRNG[35] = (LFSRcolor0[128]&LFSRcolor0[50]&LFSRcolor0[156]);
    BiasedRNG[36] = (LFSRcolor0[133]&LFSRcolor0[183]&LFSRcolor0[81]);
    BiasedRNG[37] = (LFSRcolor0[143]&LFSRcolor0[168]&LFSRcolor0[8]);
    BiasedRNG[38] = (LFSRcolor0[136]&LFSRcolor0[14]&LFSRcolor0[40]);
    BiasedRNG[39] = (LFSRcolor0[70]&LFSRcolor0[49]&LFSRcolor0[141]);
    BiasedRNG[40] = (LFSRcolor0[76]&LFSRcolor0[63]&LFSRcolor0[178]);
    BiasedRNG[41] = (LFSRcolor0[106]&LFSRcolor0[83]&LFSRcolor0[5]);
    BiasedRNG[42] = (LFSRcolor0[135]&LFSRcolor0[82]&LFSRcolor0[48]);
    BiasedRNG[43] = (LFSRcolor0[26]&LFSRcolor0[46]&LFSRcolor0[152]);
    BiasedRNG[44] = (LFSRcolor0[161]&LFSRcolor0[25]&LFSRcolor0[67]);
    BiasedRNG[45] = (LFSRcolor0[173]&LFSRcolor0[92]&LFSRcolor0[103]);
    BiasedRNG[46] = (LFSRcolor0[102]&LFSRcolor0[68]&LFSRcolor0[147]);
    UnbiasedRNG[0] = LFSRcolor0[110];
    UnbiasedRNG[1] = LFSRcolor0[75];
    UnbiasedRNG[2] = LFSRcolor0[60];
    UnbiasedRNG[3] = LFSRcolor0[71];
    UnbiasedRNG[4] = LFSRcolor0[55];
    UnbiasedRNG[5] = LFSRcolor0[126];
    UnbiasedRNG[6] = LFSRcolor0[154];
    UnbiasedRNG[7] = LFSRcolor0[138];
    UnbiasedRNG[8] = LFSRcolor0[125];
    UnbiasedRNG[9] = LFSRcolor0[78];
    UnbiasedRNG[10] = LFSRcolor0[113];
    UnbiasedRNG[11] = LFSRcolor0[88];
    UnbiasedRNG[12] = LFSRcolor0[163];
    UnbiasedRNG[13] = LFSRcolor0[170];
    UnbiasedRNG[14] = LFSRcolor0[61];
    UnbiasedRNG[15] = LFSRcolor0[80];
    UnbiasedRNG[16] = LFSRcolor0[41];
    UnbiasedRNG[17] = LFSRcolor0[104];
    UnbiasedRNG[18] = LFSRcolor0[160];
    UnbiasedRNG[19] = LFSRcolor0[30];
    UnbiasedRNG[20] = LFSRcolor0[139];
    UnbiasedRNG[21] = LFSRcolor0[4];
    UnbiasedRNG[22] = LFSRcolor0[115];
    UnbiasedRNG[23] = LFSRcolor0[120];
    UnbiasedRNG[24] = LFSRcolor0[132];
    UnbiasedRNG[25] = LFSRcolor0[33];
    UnbiasedRNG[26] = LFSRcolor0[101];
    UnbiasedRNG[27] = LFSRcolor0[35];
end

always @(posedge color0_clk) begin
    BiasedRNG[47] = (LFSRcolor1[57]&LFSRcolor1[175]&LFSRcolor1[169]);
    BiasedRNG[48] = (LFSRcolor1[51]&LFSRcolor1[29]&LFSRcolor1[134]);
    BiasedRNG[49] = (LFSRcolor1[11]&LFSRcolor1[91]&LFSRcolor1[126]);
    BiasedRNG[50] = (LFSRcolor1[77]&LFSRcolor1[162]&LFSRcolor1[96]);
    BiasedRNG[51] = (LFSRcolor1[94]&LFSRcolor1[40]&LFSRcolor1[36]);
    BiasedRNG[52] = (LFSRcolor1[171]&LFSRcolor1[173]&LFSRcolor1[54]);
    BiasedRNG[53] = (LFSRcolor1[178]&LFSRcolor1[61]&LFSRcolor1[37]);
    BiasedRNG[54] = (LFSRcolor1[22]&LFSRcolor1[70]&LFSRcolor1[118]);
    BiasedRNG[55] = (LFSRcolor1[147]&LFSRcolor1[4]&LFSRcolor1[155]);
    BiasedRNG[56] = (LFSRcolor1[139]&LFSRcolor1[127]&LFSRcolor1[13]);
    BiasedRNG[57] = (LFSRcolor1[90]&LFSRcolor1[35]&LFSRcolor1[14]);
    BiasedRNG[58] = (LFSRcolor1[59]&LFSRcolor1[164]&LFSRcolor1[69]);
    BiasedRNG[59] = (LFSRcolor1[8]&LFSRcolor1[177]&LFSRcolor1[6]);
    BiasedRNG[60] = (LFSRcolor1[2]&LFSRcolor1[83]&LFSRcolor1[64]);
    BiasedRNG[61] = (LFSRcolor1[50]&LFSRcolor1[161]&LFSRcolor1[103]);
    BiasedRNG[62] = (LFSRcolor1[21]&LFSRcolor1[117]&LFSRcolor1[56]);
    BiasedRNG[63] = (LFSRcolor1[128]&LFSRcolor1[158]&LFSRcolor1[25]);
    BiasedRNG[64] = (LFSRcolor1[144]&LFSRcolor1[67]&LFSRcolor1[47]);
    BiasedRNG[65] = (LFSRcolor1[154]&LFSRcolor1[81]&LFSRcolor1[148]);
    BiasedRNG[66] = (LFSRcolor1[10]&LFSRcolor1[108]&LFSRcolor1[100]);
    BiasedRNG[67] = (LFSRcolor1[182]&LFSRcolor1[105]&LFSRcolor1[19]);
    BiasedRNG[68] = (LFSRcolor1[152]&LFSRcolor1[42]&LFSRcolor1[73]);
    BiasedRNG[69] = (LFSRcolor1[1]&LFSRcolor1[104]&LFSRcolor1[39]);
    BiasedRNG[70] = (LFSRcolor1[16]&LFSRcolor1[23]&LFSRcolor1[60]);
    BiasedRNG[71] = (LFSRcolor1[181]&LFSRcolor1[107]&LFSRcolor1[99]);
    BiasedRNG[72] = (LFSRcolor1[122]&LFSRcolor1[75]&LFSRcolor1[18]);
    BiasedRNG[73] = (LFSRcolor1[157]&LFSRcolor1[183]&LFSRcolor1[102]);
    BiasedRNG[74] = (LFSRcolor1[111]&LFSRcolor1[113]&LFSRcolor1[110]);
    BiasedRNG[75] = (LFSRcolor1[31]&LFSRcolor1[115]&LFSRcolor1[132]);
    BiasedRNG[76] = (LFSRcolor1[120]&LFSRcolor1[78]&LFSRcolor1[153]);
    BiasedRNG[77] = (LFSRcolor1[145]&LFSRcolor1[20]&LFSRcolor1[130]);
    BiasedRNG[78] = (LFSRcolor1[84]&LFSRcolor1[3]&LFSRcolor1[176]);
    BiasedRNG[79] = (LFSRcolor1[66]&LFSRcolor1[46]&LFSRcolor1[41]);
    BiasedRNG[80] = (LFSRcolor1[112]&LFSRcolor1[44]&LFSRcolor1[12]);
    BiasedRNG[81] = (LFSRcolor1[30]&LFSRcolor1[0]&LFSRcolor1[72]);
    BiasedRNG[82] = (LFSRcolor1[15]&LFSRcolor1[160]&LFSRcolor1[168]);
    BiasedRNG[83] = (LFSRcolor1[86]&LFSRcolor1[33]&LFSRcolor1[45]);
    BiasedRNG[84] = (LFSRcolor1[124]&LFSRcolor1[74]&LFSRcolor1[7]);
    BiasedRNG[85] = (LFSRcolor1[136]&LFSRcolor1[135]&LFSRcolor1[48]);
    BiasedRNG[86] = (LFSRcolor1[9]&LFSRcolor1[76]&LFSRcolor1[82]);
    BiasedRNG[87] = (LFSRcolor1[172]&LFSRcolor1[71]&LFSRcolor1[55]);
    BiasedRNG[88] = (LFSRcolor1[123]&LFSRcolor1[97]&LFSRcolor1[165]);
    BiasedRNG[89] = (LFSRcolor1[79]&LFSRcolor1[80]&LFSRcolor1[166]);
    BiasedRNG[90] = (LFSRcolor1[119]&LFSRcolor1[142]&LFSRcolor1[34]);
    BiasedRNG[91] = (LFSRcolor1[93]&LFSRcolor1[106]&LFSRcolor1[65]);
    BiasedRNG[92] = (LFSRcolor1[125]&LFSRcolor1[174]&LFSRcolor1[26]);
    BiasedRNG[93] = (LFSRcolor1[121]&LFSRcolor1[133]&LFSRcolor1[137]);
    BiasedRNG[94] = (LFSRcolor1[49]&LFSRcolor1[88]&LFSRcolor1[156]);
    UnbiasedRNG[28] = LFSRcolor1[146];
    UnbiasedRNG[29] = LFSRcolor1[28];
    UnbiasedRNG[30] = LFSRcolor1[62];
    UnbiasedRNG[31] = LFSRcolor1[138];
    UnbiasedRNG[32] = LFSRcolor1[98];
    UnbiasedRNG[33] = LFSRcolor1[131];
    UnbiasedRNG[34] = LFSRcolor1[151];
    UnbiasedRNG[35] = LFSRcolor1[179];
    UnbiasedRNG[36] = LFSRcolor1[141];
    UnbiasedRNG[37] = LFSRcolor1[63];
    UnbiasedRNG[38] = LFSRcolor1[163];
    UnbiasedRNG[39] = LFSRcolor1[52];
    UnbiasedRNG[40] = LFSRcolor1[87];
    UnbiasedRNG[41] = LFSRcolor1[27];
    UnbiasedRNG[42] = LFSRcolor1[140];
    UnbiasedRNG[43] = LFSRcolor1[43];
    UnbiasedRNG[44] = LFSRcolor1[149];
    UnbiasedRNG[45] = LFSRcolor1[109];
    UnbiasedRNG[46] = LFSRcolor1[85];
    UnbiasedRNG[47] = LFSRcolor1[150];
    UnbiasedRNG[48] = LFSRcolor1[129];
    UnbiasedRNG[49] = LFSRcolor1[5];
    UnbiasedRNG[50] = LFSRcolor1[101];
    UnbiasedRNG[51] = LFSRcolor1[92];
    UnbiasedRNG[52] = LFSRcolor1[143];
    UnbiasedRNG[53] = LFSRcolor1[180];
    UnbiasedRNG[54] = LFSRcolor1[32];
    UnbiasedRNG[55] = LFSRcolor1[89];
    UnbiasedRNG[56] = LFSRcolor1[24];
    UnbiasedRNG[57] = LFSRcolor1[53];
end

always @(posedge color1_clk) begin
    BiasedRNG[95] = (LFSRcolor2[9]&LFSRcolor2[1]&LFSRcolor2[94]);
    BiasedRNG[96] = (LFSRcolor2[41]&LFSRcolor2[83]&LFSRcolor2[95]);
    BiasedRNG[97] = (LFSRcolor2[36]&LFSRcolor2[126]&LFSRcolor2[74]);
    BiasedRNG[98] = (LFSRcolor2[19]&LFSRcolor2[4]&LFSRcolor2[28]);
    BiasedRNG[99] = (LFSRcolor2[7]&LFSRcolor2[99]&LFSRcolor2[63]);
    BiasedRNG[100] = (LFSRcolor2[130]&LFSRcolor2[116]&LFSRcolor2[109]);
    BiasedRNG[101] = (LFSRcolor2[73]&LFSRcolor2[21]&LFSRcolor2[33]);
    BiasedRNG[102] = (LFSRcolor2[128]&LFSRcolor2[65]&LFSRcolor2[86]);
    BiasedRNG[103] = (LFSRcolor2[88]&LFSRcolor2[31]&LFSRcolor2[105]);
    BiasedRNG[104] = (LFSRcolor2[110]&LFSRcolor2[11]&LFSRcolor2[111]);
    BiasedRNG[105] = (LFSRcolor2[10]&LFSRcolor2[75]&LFSRcolor2[72]);
    BiasedRNG[106] = (LFSRcolor2[49]&LFSRcolor2[107]&LFSRcolor2[119]);
    BiasedRNG[107] = (LFSRcolor2[46]&LFSRcolor2[3]&LFSRcolor2[61]);
    BiasedRNG[108] = (LFSRcolor2[79]&LFSRcolor2[92]&LFSRcolor2[16]);
    BiasedRNG[109] = (LFSRcolor2[122]&LFSRcolor2[52]&LFSRcolor2[114]);
    BiasedRNG[110] = (LFSRcolor2[90]&LFSRcolor2[124]&LFSRcolor2[91]);
    BiasedRNG[111] = (LFSRcolor2[97]&LFSRcolor2[101]&LFSRcolor2[106]);
    BiasedRNG[112] = (LFSRcolor2[78]&LFSRcolor2[121]&LFSRcolor2[18]);
    BiasedRNG[113] = (LFSRcolor2[70]&LFSRcolor2[51]&LFSRcolor2[30]);
    BiasedRNG[114] = (LFSRcolor2[56]&LFSRcolor2[117]&LFSRcolor2[71]);
    BiasedRNG[115] = (LFSRcolor2[131]&LFSRcolor2[15]&LFSRcolor2[134]);
    BiasedRNG[116] = (LFSRcolor2[43]&LFSRcolor2[34]&LFSRcolor2[50]);
    BiasedRNG[117] = (LFSRcolor2[53]&LFSRcolor2[32]&LFSRcolor2[98]);
    BiasedRNG[118] = (LFSRcolor2[26]&LFSRcolor2[64]&LFSRcolor2[84]);
    BiasedRNG[119] = (LFSRcolor2[0]&LFSRcolor2[57]&LFSRcolor2[81]);
    BiasedRNG[120] = (LFSRcolor2[42]&LFSRcolor2[59]&LFSRcolor2[47]);
    BiasedRNG[121] = (LFSRcolor2[108]&LFSRcolor2[60]&LFSRcolor2[100]);
    BiasedRNG[122] = (LFSRcolor2[102]&LFSRcolor2[38]&LFSRcolor2[104]);
    BiasedRNG[123] = (LFSRcolor2[129]&LFSRcolor2[103]&LFSRcolor2[76]);
    BiasedRNG[124] = (LFSRcolor2[6]&LFSRcolor2[22]&LFSRcolor2[55]);
    BiasedRNG[125] = (LFSRcolor2[115]&LFSRcolor2[54]&LFSRcolor2[85]);
    BiasedRNG[126] = (LFSRcolor2[24]&LFSRcolor2[87]&LFSRcolor2[44]);
    BiasedRNG[127] = (LFSRcolor2[25]&LFSRcolor2[45]&LFSRcolor2[20]);
    BiasedRNG[128] = (LFSRcolor2[93]&LFSRcolor2[8]&LFSRcolor2[5]);
    BiasedRNG[129] = (LFSRcolor2[120]&LFSRcolor2[69]&LFSRcolor2[35]);
    BiasedRNG[130] = (LFSRcolor2[40]&LFSRcolor2[89]&LFSRcolor2[2]);
    UnbiasedRNG[58] = LFSRcolor2[29];
    UnbiasedRNG[59] = LFSRcolor2[58];
    UnbiasedRNG[60] = LFSRcolor2[113];
    UnbiasedRNG[61] = LFSRcolor2[132];
    UnbiasedRNG[62] = LFSRcolor2[48];
    UnbiasedRNG[63] = LFSRcolor2[13];
    UnbiasedRNG[64] = LFSRcolor2[80];
    UnbiasedRNG[65] = LFSRcolor2[14];
    UnbiasedRNG[66] = LFSRcolor2[68];
    UnbiasedRNG[67] = LFSRcolor2[137];
    UnbiasedRNG[68] = LFSRcolor2[135];
    UnbiasedRNG[69] = LFSRcolor2[62];
    UnbiasedRNG[70] = LFSRcolor2[66];
    UnbiasedRNG[71] = LFSRcolor2[12];
    UnbiasedRNG[72] = LFSRcolor2[118];
    UnbiasedRNG[73] = LFSRcolor2[67];
    UnbiasedRNG[74] = LFSRcolor2[37];
    UnbiasedRNG[75] = LFSRcolor2[82];
    UnbiasedRNG[76] = LFSRcolor2[136];
    UnbiasedRNG[77] = LFSRcolor2[77];
    UnbiasedRNG[78] = LFSRcolor2[127];
    UnbiasedRNG[79] = LFSRcolor2[96];
    UnbiasedRNG[80] = LFSRcolor2[112];
    UnbiasedRNG[81] = LFSRcolor2[125];
    UnbiasedRNG[82] = LFSRcolor2[27];
    UnbiasedRNG[83] = LFSRcolor2[23];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[84] = LFSRcolor3[30];
    UnbiasedRNG[85] = LFSRcolor3[44];
    UnbiasedRNG[86] = LFSRcolor3[14];
    UnbiasedRNG[87] = LFSRcolor3[8];
    UnbiasedRNG[88] = LFSRcolor3[26];
    UnbiasedRNG[89] = LFSRcolor3[45];
    UnbiasedRNG[90] = LFSRcolor3[1];
    UnbiasedRNG[91] = LFSRcolor3[37];
    UnbiasedRNG[92] = LFSRcolor3[22];
    UnbiasedRNG[93] = LFSRcolor3[24];
    UnbiasedRNG[94] = LFSRcolor3[34];
    UnbiasedRNG[95] = LFSRcolor3[42];
    UnbiasedRNG[96] = LFSRcolor3[28];
    UnbiasedRNG[97] = LFSRcolor3[40];
    UnbiasedRNG[98] = LFSRcolor3[16];
    UnbiasedRNG[99] = LFSRcolor3[32];
    UnbiasedRNG[100] = LFSRcolor3[7];
    UnbiasedRNG[101] = LFSRcolor3[20];
    UnbiasedRNG[102] = LFSRcolor3[13];
    UnbiasedRNG[103] = LFSRcolor3[15];
end

always @(posedge color3_clk) begin
    BiasedRNG[131] = (LFSRcolor4[89]&LFSRcolor4[3]&LFSRcolor4[13]);
    BiasedRNG[132] = (LFSRcolor4[8]&LFSRcolor4[83]&LFSRcolor4[17]);
    BiasedRNG[133] = (LFSRcolor4[37]&LFSRcolor4[79]&LFSRcolor4[10]);
    BiasedRNG[134] = (LFSRcolor4[28]&LFSRcolor4[66]&LFSRcolor4[44]);
    BiasedRNG[135] = (LFSRcolor4[51]&LFSRcolor4[76]&LFSRcolor4[63]);
    BiasedRNG[136] = (LFSRcolor4[42]&LFSRcolor4[20]&LFSRcolor4[72]);
    BiasedRNG[137] = (LFSRcolor4[77]&LFSRcolor4[55]&LFSRcolor4[88]);
    BiasedRNG[138] = (LFSRcolor4[47]&LFSRcolor4[41]&LFSRcolor4[56]);
    BiasedRNG[139] = (LFSRcolor4[18]&LFSRcolor4[85]&LFSRcolor4[15]);
    BiasedRNG[140] = (LFSRcolor4[86]&LFSRcolor4[62]&LFSRcolor4[75]);
    BiasedRNG[141] = (LFSRcolor4[38]&LFSRcolor4[60]&LFSRcolor4[70]);
    BiasedRNG[142] = (LFSRcolor4[49]&LFSRcolor4[58]&LFSRcolor4[34]);
    BiasedRNG[143] = (LFSRcolor4[7]&LFSRcolor4[16]&LFSRcolor4[26]);
    BiasedRNG[144] = (LFSRcolor4[90]&LFSRcolor4[53]&LFSRcolor4[30]);
    BiasedRNG[145] = (LFSRcolor4[61]&LFSRcolor4[91]&LFSRcolor4[52]);
    BiasedRNG[146] = (LFSRcolor4[6]&LFSRcolor4[80]&LFSRcolor4[46]);
    BiasedRNG[147] = (LFSRcolor4[32]&LFSRcolor4[35]&LFSRcolor4[40]);
    BiasedRNG[148] = (LFSRcolor4[69]&LFSRcolor4[71]&LFSRcolor4[65]);
    BiasedRNG[149] = (LFSRcolor4[36]&LFSRcolor4[14]&LFSRcolor4[39]);
    BiasedRNG[150] = (LFSRcolor4[57]&LFSRcolor4[0]&LFSRcolor4[59]);
    BiasedRNG[151] = (LFSRcolor4[27]&LFSRcolor4[2]&LFSRcolor4[4]);
    BiasedRNG[152] = (LFSRcolor4[84]&LFSRcolor4[74]&LFSRcolor4[5]);
    BiasedRNG[153] = (LFSRcolor4[43]&LFSRcolor4[23]&LFSRcolor4[21]);
    BiasedRNG[154] = (LFSRcolor4[24]&LFSRcolor4[1]&LFSRcolor4[22]);
    BiasedRNG[155] = (LFSRcolor4[68]&LFSRcolor4[45]&LFSRcolor4[48]);
    BiasedRNG[156] = (LFSRcolor4[78]&LFSRcolor4[19]&LFSRcolor4[67]);
    BiasedRNG[157] = (LFSRcolor4[73]&LFSRcolor4[33]&LFSRcolor4[29]);
    BiasedRNG[158] = (LFSRcolor4[50]&LFSRcolor4[31]&LFSRcolor4[12]);
    BiasedRNG[159] = (LFSRcolor4[11]&LFSRcolor4[82]&LFSRcolor4[9]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

//Generate the ILA for data collection:
ila_0 ILAinst(.clk(sample_clk),.probe0(run),.probe1(solution_flag),.probe2(failure),.probe3(counter[37:0]));

//Instantiate VIO:
vio_0 VIOinst (.clk(sample_clk),.probe_out0(reset),.probe_out1(solution_set[11:0]));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule