//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [5:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [91:0] LFSRcolor0;
wire [45:0] LFSRcolor1;
wire [45:0] LFSRcolor2;
wire [45:0] LFSRcolor3;
wire [45:0] LFSRcolor4;
reg [36:0] BiasedRNG;       //For I=+/-1 cases
reg [16:0] UnbiasedRNG;   //For I=0 cases
reg [0:62] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[24] = 1'b0;
initial m[36] = 1'b1;
initial m[46] = 1'b0;
initial m[56] = 1'b1;
initial m[61] = 1'b0;
initial m[62] = 1'b0;

//Initialize the PBits clamped to zero:
initial m[35] = 1'b0;
initial m[45] = 1'b0;
initial m[48] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 0;
initial m[1] = 1;
initial m[2] = 0;
initial m[3] = 0;
initial m[4] = 0;
initial m[5] = 0;
initial m[6] = 0;
initial m[7] = 1;
initial m[8] = 1;
initial m[9] = 0;
initial m[10] = 0;
initial m[11] = 1;
initial m[12] = 1;
initial m[13] = 0;
initial m[14] = 0;
initial m[15] = 0;
initial m[16] = 0;
initial m[17] = 1;
initial m[18] = 1;
initial m[19] = 0;
initial m[20] = 0;
initial m[21] = 1;
initial m[22] = 1;
initial m[23] = 1;
initial m[25] = 1;
initial m[26] = 0;
initial m[27] = 0;
initial m[28] = 0;
initial m[29] = 1;
initial m[30] = 1;
initial m[31] = 0;
initial m[32] = 1;
initial m[33] = 0;
initial m[34] = 1;
initial m[37] = 0;
initial m[38] = 0;
initial m[39] = 1;
initial m[40] = 1;
initial m[41] = 0;
initial m[42] = 0;
initial m[43] = 1;
initial m[44] = 1;
initial m[47] = 1;
initial m[49] = 1;
initial m[50] = 1;
initial m[51] = 0;
initial m[52] = 1;
initial m[53] = 1;
initial m[54] = 1;
initial m[55] = 1;
initial m[57] = 1;
initial m[58] = 1;
initial m[59] = 0;
initial m[60] = 0;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[2],m[1],m[0]}*{m[5],m[4],m[3]};
end

always @(negedge sample_clk) begin
    if (solution == 6'b001010)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[6]&~m[7]&~m[8])|(~m[6]&m[7]&~m[8])|(~m[6]&~m[7]&m[8]))&BiasedRNG[0])|(((m[6]&m[7]&~m[8])|(m[6]&~m[7]&m[8])|(~m[6]&m[7]&m[8]))&~BiasedRNG[0])|((m[6]&m[7]&m[8]));
    m[1] = (((m[9]&~m[10]&~m[11])|(~m[9]&m[10]&~m[11])|(~m[9]&~m[10]&m[11]))&BiasedRNG[1])|(((m[9]&m[10]&~m[11])|(m[9]&~m[10]&m[11])|(~m[9]&m[10]&m[11]))&~BiasedRNG[1])|((m[9]&m[10]&m[11]));
    m[2] = (((m[12]&~m[13]&~m[14])|(~m[12]&m[13]&~m[14])|(~m[12]&~m[13]&m[14]))&BiasedRNG[2])|(((m[12]&m[13]&~m[14])|(m[12]&~m[13]&m[14])|(~m[12]&m[13]&m[14]))&~BiasedRNG[2])|((m[12]&m[13]&m[14]));
    m[3] = (((m[15]&~m[16]&~m[17])|(~m[15]&m[16]&~m[17])|(~m[15]&~m[16]&m[17]))&BiasedRNG[3])|(((m[15]&m[16]&~m[17])|(m[15]&~m[16]&m[17])|(~m[15]&m[16]&m[17]))&~BiasedRNG[3])|((m[15]&m[16]&m[17]));
    m[4] = (((m[18]&~m[19]&~m[20])|(~m[18]&m[19]&~m[20])|(~m[18]&~m[19]&m[20]))&BiasedRNG[4])|(((m[18]&m[19]&~m[20])|(m[18]&~m[19]&m[20])|(~m[18]&m[19]&m[20]))&~BiasedRNG[4])|((m[18]&m[19]&m[20]));
    m[5] = (((m[21]&~m[22]&~m[23])|(~m[21]&m[22]&~m[23])|(~m[21]&~m[22]&m[23]))&BiasedRNG[5])|(((m[21]&m[22]&~m[23])|(m[21]&~m[22]&m[23])|(~m[21]&m[22]&m[23]))&~BiasedRNG[5])|((m[21]&m[22]&m[23]));
    m[25] = (((m[9]&~m[16]&m[33])|(~m[9]&m[16]&m[33]))&BiasedRNG[6])|(((m[9]&m[16]&~m[33]))&~BiasedRNG[6])|((m[9]&m[16]&m[33]));
    m[26] = (((m[12]&~m[17]&m[38])|(~m[12]&m[17]&m[38]))&BiasedRNG[7])|(((m[12]&m[17]&~m[38]))&~BiasedRNG[7])|((m[12]&m[17]&m[38]));
    m[27] = (((m[7]&~m[18]&m[34])|(~m[7]&m[18]&m[34]))&BiasedRNG[8])|(((m[7]&m[18]&~m[34]))&~BiasedRNG[8])|((m[7]&m[18]&m[34]));
    m[28] = (((m[10]&~m[19]&m[39])|(~m[10]&m[19]&m[39]))&BiasedRNG[9])|(((m[10]&m[19]&~m[39]))&~BiasedRNG[9])|((m[10]&m[19]&m[39]));
    m[29] = (((m[13]&~m[20]&m[49])|(~m[13]&m[20]&m[49]))&BiasedRNG[10])|(((m[13]&m[20]&~m[49]))&~BiasedRNG[10])|((m[13]&m[20]&m[49]));
    m[30] = (((m[8]&~m[21]&m[44])|(~m[8]&m[21]&m[44]))&BiasedRNG[11])|(((m[8]&m[21]&~m[44]))&~BiasedRNG[11])|((m[8]&m[21]&m[44]));
    m[31] = (((m[11]&~m[22]&m[54])|(~m[11]&m[22]&m[54]))&BiasedRNG[12])|(((m[11]&m[22]&~m[54]))&~BiasedRNG[12])|((m[11]&m[22]&m[54]));
    m[32] = (((m[14]&~m[23]&m[59])|(~m[14]&m[23]&m[59]))&BiasedRNG[13])|(((m[14]&m[23]&~m[59]))&~BiasedRNG[13])|((m[14]&m[23]&m[59]));
    m[40] = (((m[37]&~m[38]&~m[39]&~m[41]&~m[42])|(~m[37]&~m[38]&~m[39]&m[41]&~m[42])|(m[37]&m[38]&~m[39]&m[41]&~m[42])|(m[37]&~m[38]&m[39]&m[41]&~m[42])|(~m[37]&m[38]&~m[39]&~m[41]&m[42])|(~m[37]&~m[38]&m[39]&~m[41]&m[42])|(m[37]&m[38]&m[39]&~m[41]&m[42])|(~m[37]&m[38]&m[39]&m[41]&m[42]))&UnbiasedRNG[0])|((m[37]&~m[38]&~m[39]&m[41]&~m[42])|(~m[37]&~m[38]&~m[39]&~m[41]&m[42])|(m[37]&~m[38]&~m[39]&~m[41]&m[42])|(m[37]&m[38]&~m[39]&~m[41]&m[42])|(m[37]&~m[38]&m[39]&~m[41]&m[42])|(~m[37]&~m[38]&~m[39]&m[41]&m[42])|(m[37]&~m[38]&~m[39]&m[41]&m[42])|(~m[37]&m[38]&~m[39]&m[41]&m[42])|(m[37]&m[38]&~m[39]&m[41]&m[42])|(~m[37]&~m[38]&m[39]&m[41]&m[42])|(m[37]&~m[38]&m[39]&m[41]&m[42])|(m[37]&m[38]&m[39]&m[41]&m[42]));
    m[43] = (((m[41]&~m[44]&~m[45]&~m[46]&~m[47])|(~m[41]&~m[44]&~m[45]&m[46]&~m[47])|(m[41]&m[44]&~m[45]&m[46]&~m[47])|(m[41]&~m[44]&m[45]&m[46]&~m[47])|(~m[41]&m[44]&~m[45]&~m[46]&m[47])|(~m[41]&~m[44]&m[45]&~m[46]&m[47])|(m[41]&m[44]&m[45]&~m[46]&m[47])|(~m[41]&m[44]&m[45]&m[46]&m[47]))&UnbiasedRNG[1])|((m[41]&~m[44]&~m[45]&m[46]&~m[47])|(~m[41]&~m[44]&~m[45]&~m[46]&m[47])|(m[41]&~m[44]&~m[45]&~m[46]&m[47])|(m[41]&m[44]&~m[45]&~m[46]&m[47])|(m[41]&~m[44]&m[45]&~m[46]&m[47])|(~m[41]&~m[44]&~m[45]&m[46]&m[47])|(m[41]&~m[44]&~m[45]&m[46]&m[47])|(~m[41]&m[44]&~m[45]&m[46]&m[47])|(m[41]&m[44]&~m[45]&m[46]&m[47])|(~m[41]&~m[44]&m[45]&m[46]&m[47])|(m[41]&~m[44]&m[45]&m[46]&m[47])|(m[41]&m[44]&m[45]&m[46]&m[47]));
    m[53] = (((m[51]&~m[54]&~m[55]&~m[56]&~m[57])|(~m[51]&~m[54]&~m[55]&m[56]&~m[57])|(m[51]&m[54]&~m[55]&m[56]&~m[57])|(m[51]&~m[54]&m[55]&m[56]&~m[57])|(~m[51]&m[54]&~m[55]&~m[56]&m[57])|(~m[51]&~m[54]&m[55]&~m[56]&m[57])|(m[51]&m[54]&m[55]&~m[56]&m[57])|(~m[51]&m[54]&m[55]&m[56]&m[57]))&UnbiasedRNG[2])|((m[51]&~m[54]&~m[55]&m[56]&~m[57])|(~m[51]&~m[54]&~m[55]&~m[56]&m[57])|(m[51]&~m[54]&~m[55]&~m[56]&m[57])|(m[51]&m[54]&~m[55]&~m[56]&m[57])|(m[51]&~m[54]&m[55]&~m[56]&m[57])|(~m[51]&~m[54]&~m[55]&m[56]&m[57])|(m[51]&~m[54]&~m[55]&m[56]&m[57])|(~m[51]&m[54]&~m[55]&m[56]&m[57])|(m[51]&m[54]&~m[55]&m[56]&m[57])|(~m[51]&~m[54]&m[55]&m[56]&m[57])|(m[51]&~m[54]&m[55]&m[56]&m[57])|(m[51]&m[54]&m[55]&m[56]&m[57]));
    m[58] = (((m[52]&~m[59]&~m[60]&~m[61]&~m[62])|(~m[52]&~m[59]&~m[60]&m[61]&~m[62])|(m[52]&m[59]&~m[60]&m[61]&~m[62])|(m[52]&~m[59]&m[60]&m[61]&~m[62])|(~m[52]&m[59]&~m[60]&~m[61]&m[62])|(~m[52]&~m[59]&m[60]&~m[61]&m[62])|(m[52]&m[59]&m[60]&~m[61]&m[62])|(~m[52]&m[59]&m[60]&m[61]&m[62]))&UnbiasedRNG[3])|((m[52]&~m[59]&~m[60]&m[61]&~m[62])|(~m[52]&~m[59]&~m[60]&~m[61]&m[62])|(m[52]&~m[59]&~m[60]&~m[61]&m[62])|(m[52]&m[59]&~m[60]&~m[61]&m[62])|(m[52]&~m[59]&m[60]&~m[61]&m[62])|(~m[52]&~m[59]&~m[60]&m[61]&m[62])|(m[52]&~m[59]&~m[60]&m[61]&m[62])|(~m[52]&m[59]&~m[60]&m[61]&m[62])|(m[52]&m[59]&~m[60]&m[61]&m[62])|(~m[52]&~m[59]&m[60]&m[61]&m[62])|(m[52]&~m[59]&m[60]&m[61]&m[62])|(m[52]&m[59]&m[60]&m[61]&m[62]));
end

always @(posedge color1_clk) begin
    m[6] = (((~m[0]&~m[15]&~m[24])|(m[0]&m[15]&~m[24]))&BiasedRNG[14])|(((m[0]&~m[15]&~m[24])|(~m[0]&m[15]&m[24]))&~BiasedRNG[14])|((~m[0]&~m[15]&m[24])|(m[0]&~m[15]&m[24])|(m[0]&m[15]&m[24]));
    m[7] = (((~m[0]&~m[18]&~m[27])|(m[0]&m[18]&~m[27]))&BiasedRNG[15])|(((m[0]&~m[18]&~m[27])|(~m[0]&m[18]&m[27]))&~BiasedRNG[15])|((~m[0]&~m[18]&m[27])|(m[0]&~m[18]&m[27])|(m[0]&m[18]&m[27]));
    m[8] = (((~m[0]&~m[21]&~m[30])|(m[0]&m[21]&~m[30]))&BiasedRNG[16])|(((m[0]&~m[21]&~m[30])|(~m[0]&m[21]&m[30]))&~BiasedRNG[16])|((~m[0]&~m[21]&m[30])|(m[0]&~m[21]&m[30])|(m[0]&m[21]&m[30]));
    m[9] = (((~m[1]&~m[16]&~m[25])|(m[1]&m[16]&~m[25]))&BiasedRNG[17])|(((m[1]&~m[16]&~m[25])|(~m[1]&m[16]&m[25]))&~BiasedRNG[17])|((~m[1]&~m[16]&m[25])|(m[1]&~m[16]&m[25])|(m[1]&m[16]&m[25]));
    m[10] = (((~m[1]&~m[19]&~m[28])|(m[1]&m[19]&~m[28]))&BiasedRNG[18])|(((m[1]&~m[19]&~m[28])|(~m[1]&m[19]&m[28]))&~BiasedRNG[18])|((~m[1]&~m[19]&m[28])|(m[1]&~m[19]&m[28])|(m[1]&m[19]&m[28]));
    m[11] = (((~m[1]&~m[22]&~m[31])|(m[1]&m[22]&~m[31]))&BiasedRNG[19])|(((m[1]&~m[22]&~m[31])|(~m[1]&m[22]&m[31]))&~BiasedRNG[19])|((~m[1]&~m[22]&m[31])|(m[1]&~m[22]&m[31])|(m[1]&m[22]&m[31]));
    m[12] = (((~m[2]&~m[17]&~m[26])|(m[2]&m[17]&~m[26]))&BiasedRNG[20])|(((m[2]&~m[17]&~m[26])|(~m[2]&m[17]&m[26]))&~BiasedRNG[20])|((~m[2]&~m[17]&m[26])|(m[2]&~m[17]&m[26])|(m[2]&m[17]&m[26]));
    m[13] = (((~m[2]&~m[20]&~m[29])|(m[2]&m[20]&~m[29]))&BiasedRNG[21])|(((m[2]&~m[20]&~m[29])|(~m[2]&m[20]&m[29]))&~BiasedRNG[21])|((~m[2]&~m[20]&m[29])|(m[2]&~m[20]&m[29])|(m[2]&m[20]&m[29]));
    m[14] = (((~m[2]&~m[23]&~m[32])|(m[2]&m[23]&~m[32]))&BiasedRNG[22])|(((m[2]&~m[23]&~m[32])|(~m[2]&m[23]&m[32]))&~BiasedRNG[22])|((~m[2]&~m[23]&m[32])|(m[2]&~m[23]&m[32])|(m[2]&m[23]&m[32]));
    m[33] = (((m[25]&~m[34]&~m[35]&~m[36]&~m[37])|(~m[25]&~m[34]&~m[35]&m[36]&~m[37])|(m[25]&m[34]&~m[35]&m[36]&~m[37])|(m[25]&~m[34]&m[35]&m[36]&~m[37])|(~m[25]&m[34]&~m[35]&~m[36]&m[37])|(~m[25]&~m[34]&m[35]&~m[36]&m[37])|(m[25]&m[34]&m[35]&~m[36]&m[37])|(~m[25]&m[34]&m[35]&m[36]&m[37]))&UnbiasedRNG[4])|((m[25]&~m[34]&~m[35]&m[36]&~m[37])|(~m[25]&~m[34]&~m[35]&~m[36]&m[37])|(m[25]&~m[34]&~m[35]&~m[36]&m[37])|(m[25]&m[34]&~m[35]&~m[36]&m[37])|(m[25]&~m[34]&m[35]&~m[36]&m[37])|(~m[25]&~m[34]&~m[35]&m[36]&m[37])|(m[25]&~m[34]&~m[35]&m[36]&m[37])|(~m[25]&m[34]&~m[35]&m[36]&m[37])|(m[25]&m[34]&~m[35]&m[36]&m[37])|(~m[25]&~m[34]&m[35]&m[36]&m[37])|(m[25]&~m[34]&m[35]&m[36]&m[37])|(m[25]&m[34]&m[35]&m[36]&m[37]));
    m[38] = (((m[26]&~m[39]&~m[40]&~m[41]&~m[42])|(~m[26]&~m[39]&~m[40]&m[41]&~m[42])|(m[26]&m[39]&~m[40]&m[41]&~m[42])|(m[26]&~m[39]&m[40]&m[41]&~m[42])|(~m[26]&m[39]&~m[40]&~m[41]&m[42])|(~m[26]&~m[39]&m[40]&~m[41]&m[42])|(m[26]&m[39]&m[40]&~m[41]&m[42])|(~m[26]&m[39]&m[40]&m[41]&m[42]))&UnbiasedRNG[5])|((m[26]&~m[39]&~m[40]&m[41]&~m[42])|(~m[26]&~m[39]&~m[40]&~m[41]&m[42])|(m[26]&~m[39]&~m[40]&~m[41]&m[42])|(m[26]&m[39]&~m[40]&~m[41]&m[42])|(m[26]&~m[39]&m[40]&~m[41]&m[42])|(~m[26]&~m[39]&~m[40]&m[41]&m[42])|(m[26]&~m[39]&~m[40]&m[41]&m[42])|(~m[26]&m[39]&~m[40]&m[41]&m[42])|(m[26]&m[39]&~m[40]&m[41]&m[42])|(~m[26]&~m[39]&m[40]&m[41]&m[42])|(m[26]&~m[39]&m[40]&m[41]&m[42])|(m[26]&m[39]&m[40]&m[41]&m[42]));
    m[44] = (((m[30]&~m[43]&~m[45]&~m[46]&~m[47])|(~m[30]&~m[43]&~m[45]&m[46]&~m[47])|(m[30]&m[43]&~m[45]&m[46]&~m[47])|(m[30]&~m[43]&m[45]&m[46]&~m[47])|(~m[30]&m[43]&~m[45]&~m[46]&m[47])|(~m[30]&~m[43]&m[45]&~m[46]&m[47])|(m[30]&m[43]&m[45]&~m[46]&m[47])|(~m[30]&m[43]&m[45]&m[46]&m[47]))&UnbiasedRNG[6])|((m[30]&~m[43]&~m[45]&m[46]&~m[47])|(~m[30]&~m[43]&~m[45]&~m[46]&m[47])|(m[30]&~m[43]&~m[45]&~m[46]&m[47])|(m[30]&m[43]&~m[45]&~m[46]&m[47])|(m[30]&~m[43]&m[45]&~m[46]&m[47])|(~m[30]&~m[43]&~m[45]&m[46]&m[47])|(m[30]&~m[43]&~m[45]&m[46]&m[47])|(~m[30]&m[43]&~m[45]&m[46]&m[47])|(m[30]&m[43]&~m[45]&m[46]&m[47])|(~m[30]&~m[43]&m[45]&m[46]&m[47])|(m[30]&~m[43]&m[45]&m[46]&m[47])|(m[30]&m[43]&m[45]&m[46]&m[47]));
    m[49] = (((m[29]&~m[48]&~m[50]&~m[51]&~m[52])|(~m[29]&~m[48]&~m[50]&m[51]&~m[52])|(m[29]&m[48]&~m[50]&m[51]&~m[52])|(m[29]&~m[48]&m[50]&m[51]&~m[52])|(~m[29]&m[48]&~m[50]&~m[51]&m[52])|(~m[29]&~m[48]&m[50]&~m[51]&m[52])|(m[29]&m[48]&m[50]&~m[51]&m[52])|(~m[29]&m[48]&m[50]&m[51]&m[52]))&UnbiasedRNG[7])|((m[29]&~m[48]&~m[50]&m[51]&~m[52])|(~m[29]&~m[48]&~m[50]&~m[51]&m[52])|(m[29]&~m[48]&~m[50]&~m[51]&m[52])|(m[29]&m[48]&~m[50]&~m[51]&m[52])|(m[29]&~m[48]&m[50]&~m[51]&m[52])|(~m[29]&~m[48]&~m[50]&m[51]&m[52])|(m[29]&~m[48]&~m[50]&m[51]&m[52])|(~m[29]&m[48]&~m[50]&m[51]&m[52])|(m[29]&m[48]&~m[50]&m[51]&m[52])|(~m[29]&~m[48]&m[50]&m[51]&m[52])|(m[29]&~m[48]&m[50]&m[51]&m[52])|(m[29]&m[48]&m[50]&m[51]&m[52]));
    m[54] = (((m[31]&~m[53]&~m[55]&~m[56]&~m[57])|(~m[31]&~m[53]&~m[55]&m[56]&~m[57])|(m[31]&m[53]&~m[55]&m[56]&~m[57])|(m[31]&~m[53]&m[55]&m[56]&~m[57])|(~m[31]&m[53]&~m[55]&~m[56]&m[57])|(~m[31]&~m[53]&m[55]&~m[56]&m[57])|(m[31]&m[53]&m[55]&~m[56]&m[57])|(~m[31]&m[53]&m[55]&m[56]&m[57]))&UnbiasedRNG[8])|((m[31]&~m[53]&~m[55]&m[56]&~m[57])|(~m[31]&~m[53]&~m[55]&~m[56]&m[57])|(m[31]&~m[53]&~m[55]&~m[56]&m[57])|(m[31]&m[53]&~m[55]&~m[56]&m[57])|(m[31]&~m[53]&m[55]&~m[56]&m[57])|(~m[31]&~m[53]&~m[55]&m[56]&m[57])|(m[31]&~m[53]&~m[55]&m[56]&m[57])|(~m[31]&m[53]&~m[55]&m[56]&m[57])|(m[31]&m[53]&~m[55]&m[56]&m[57])|(~m[31]&~m[53]&m[55]&m[56]&m[57])|(m[31]&~m[53]&m[55]&m[56]&m[57])|(m[31]&m[53]&m[55]&m[56]&m[57]));
    m[59] = (((m[32]&~m[58]&~m[60]&~m[61]&~m[62])|(~m[32]&~m[58]&~m[60]&m[61]&~m[62])|(m[32]&m[58]&~m[60]&m[61]&~m[62])|(m[32]&~m[58]&m[60]&m[61]&~m[62])|(~m[32]&m[58]&~m[60]&~m[61]&m[62])|(~m[32]&~m[58]&m[60]&~m[61]&m[62])|(m[32]&m[58]&m[60]&~m[61]&m[62])|(~m[32]&m[58]&m[60]&m[61]&m[62]))&UnbiasedRNG[9])|((m[32]&~m[58]&~m[60]&m[61]&~m[62])|(~m[32]&~m[58]&~m[60]&~m[61]&m[62])|(m[32]&~m[58]&~m[60]&~m[61]&m[62])|(m[32]&m[58]&~m[60]&~m[61]&m[62])|(m[32]&~m[58]&m[60]&~m[61]&m[62])|(~m[32]&~m[58]&~m[60]&m[61]&m[62])|(m[32]&~m[58]&~m[60]&m[61]&m[62])|(~m[32]&m[58]&~m[60]&m[61]&m[62])|(m[32]&m[58]&~m[60]&m[61]&m[62])|(~m[32]&~m[58]&m[60]&m[61]&m[62])|(m[32]&~m[58]&m[60]&m[61]&m[62])|(m[32]&m[58]&m[60]&m[61]&m[62]));
end

always @(posedge color2_clk) begin
    m[15] = (((~m[3]&~m[6]&~m[24])|(m[3]&m[6]&~m[24]))&BiasedRNG[23])|(((m[3]&~m[6]&~m[24])|(~m[3]&m[6]&m[24]))&~BiasedRNG[23])|((~m[3]&~m[6]&m[24])|(m[3]&~m[6]&m[24])|(m[3]&m[6]&m[24]));
    m[16] = (((~m[3]&~m[9]&~m[25])|(m[3]&m[9]&~m[25]))&BiasedRNG[24])|(((m[3]&~m[9]&~m[25])|(~m[3]&m[9]&m[25]))&~BiasedRNG[24])|((~m[3]&~m[9]&m[25])|(m[3]&~m[9]&m[25])|(m[3]&m[9]&m[25]));
    m[17] = (((~m[3]&~m[12]&~m[26])|(m[3]&m[12]&~m[26]))&BiasedRNG[25])|(((m[3]&~m[12]&~m[26])|(~m[3]&m[12]&m[26]))&~BiasedRNG[25])|((~m[3]&~m[12]&m[26])|(m[3]&~m[12]&m[26])|(m[3]&m[12]&m[26]));
    m[18] = (((~m[4]&~m[7]&~m[27])|(m[4]&m[7]&~m[27]))&BiasedRNG[26])|(((m[4]&~m[7]&~m[27])|(~m[4]&m[7]&m[27]))&~BiasedRNG[26])|((~m[4]&~m[7]&m[27])|(m[4]&~m[7]&m[27])|(m[4]&m[7]&m[27]));
    m[19] = (((~m[4]&~m[10]&~m[28])|(m[4]&m[10]&~m[28]))&BiasedRNG[27])|(((m[4]&~m[10]&~m[28])|(~m[4]&m[10]&m[28]))&~BiasedRNG[27])|((~m[4]&~m[10]&m[28])|(m[4]&~m[10]&m[28])|(m[4]&m[10]&m[28]));
    m[20] = (((~m[4]&~m[13]&~m[29])|(m[4]&m[13]&~m[29]))&BiasedRNG[28])|(((m[4]&~m[13]&~m[29])|(~m[4]&m[13]&m[29]))&~BiasedRNG[28])|((~m[4]&~m[13]&m[29])|(m[4]&~m[13]&m[29])|(m[4]&m[13]&m[29]));
    m[21] = (((~m[5]&~m[8]&~m[30])|(m[5]&m[8]&~m[30]))&BiasedRNG[29])|(((m[5]&~m[8]&~m[30])|(~m[5]&m[8]&m[30]))&~BiasedRNG[29])|((~m[5]&~m[8]&m[30])|(m[5]&~m[8]&m[30])|(m[5]&m[8]&m[30]));
    m[22] = (((~m[5]&~m[11]&~m[31])|(m[5]&m[11]&~m[31]))&BiasedRNG[30])|(((m[5]&~m[11]&~m[31])|(~m[5]&m[11]&m[31]))&~BiasedRNG[30])|((~m[5]&~m[11]&m[31])|(m[5]&~m[11]&m[31])|(m[5]&m[11]&m[31]));
    m[23] = (((~m[5]&~m[14]&~m[32])|(m[5]&m[14]&~m[32]))&BiasedRNG[31])|(((m[5]&~m[14]&~m[32])|(~m[5]&m[14]&m[32]))&~BiasedRNG[31])|((~m[5]&~m[14]&m[32])|(m[5]&~m[14]&m[32])|(m[5]&m[14]&m[32]));
    m[34] = (((m[27]&~m[33]&~m[35]&~m[36]&~m[37])|(~m[27]&~m[33]&~m[35]&m[36]&~m[37])|(m[27]&m[33]&~m[35]&m[36]&~m[37])|(m[27]&~m[33]&m[35]&m[36]&~m[37])|(~m[27]&m[33]&~m[35]&~m[36]&m[37])|(~m[27]&~m[33]&m[35]&~m[36]&m[37])|(m[27]&m[33]&m[35]&~m[36]&m[37])|(~m[27]&m[33]&m[35]&m[36]&m[37]))&UnbiasedRNG[10])|((m[27]&~m[33]&~m[35]&m[36]&~m[37])|(~m[27]&~m[33]&~m[35]&~m[36]&m[37])|(m[27]&~m[33]&~m[35]&~m[36]&m[37])|(m[27]&m[33]&~m[35]&~m[36]&m[37])|(m[27]&~m[33]&m[35]&~m[36]&m[37])|(~m[27]&~m[33]&~m[35]&m[36]&m[37])|(m[27]&~m[33]&~m[35]&m[36]&m[37])|(~m[27]&m[33]&~m[35]&m[36]&m[37])|(m[27]&m[33]&~m[35]&m[36]&m[37])|(~m[27]&~m[33]&m[35]&m[36]&m[37])|(m[27]&~m[33]&m[35]&m[36]&m[37])|(m[27]&m[33]&m[35]&m[36]&m[37]));
    m[39] = (((m[28]&~m[38]&~m[40]&~m[41]&~m[42])|(~m[28]&~m[38]&~m[40]&m[41]&~m[42])|(m[28]&m[38]&~m[40]&m[41]&~m[42])|(m[28]&~m[38]&m[40]&m[41]&~m[42])|(~m[28]&m[38]&~m[40]&~m[41]&m[42])|(~m[28]&~m[38]&m[40]&~m[41]&m[42])|(m[28]&m[38]&m[40]&~m[41]&m[42])|(~m[28]&m[38]&m[40]&m[41]&m[42]))&UnbiasedRNG[11])|((m[28]&~m[38]&~m[40]&m[41]&~m[42])|(~m[28]&~m[38]&~m[40]&~m[41]&m[42])|(m[28]&~m[38]&~m[40]&~m[41]&m[42])|(m[28]&m[38]&~m[40]&~m[41]&m[42])|(m[28]&~m[38]&m[40]&~m[41]&m[42])|(~m[28]&~m[38]&~m[40]&m[41]&m[42])|(m[28]&~m[38]&~m[40]&m[41]&m[42])|(~m[28]&m[38]&~m[40]&m[41]&m[42])|(m[28]&m[38]&~m[40]&m[41]&m[42])|(~m[28]&~m[38]&m[40]&m[41]&m[42])|(m[28]&~m[38]&m[40]&m[41]&m[42])|(m[28]&m[38]&m[40]&m[41]&m[42]));
    m[50] = (((m[42]&~m[48]&~m[49]&~m[51]&~m[52])|(~m[42]&~m[48]&~m[49]&m[51]&~m[52])|(m[42]&m[48]&~m[49]&m[51]&~m[52])|(m[42]&~m[48]&m[49]&m[51]&~m[52])|(~m[42]&m[48]&~m[49]&~m[51]&m[52])|(~m[42]&~m[48]&m[49]&~m[51]&m[52])|(m[42]&m[48]&m[49]&~m[51]&m[52])|(~m[42]&m[48]&m[49]&m[51]&m[52]))&UnbiasedRNG[12])|((m[42]&~m[48]&~m[49]&m[51]&~m[52])|(~m[42]&~m[48]&~m[49]&~m[51]&m[52])|(m[42]&~m[48]&~m[49]&~m[51]&m[52])|(m[42]&m[48]&~m[49]&~m[51]&m[52])|(m[42]&~m[48]&m[49]&~m[51]&m[52])|(~m[42]&~m[48]&~m[49]&m[51]&m[52])|(m[42]&~m[48]&~m[49]&m[51]&m[52])|(~m[42]&m[48]&~m[49]&m[51]&m[52])|(m[42]&m[48]&~m[49]&m[51]&m[52])|(~m[42]&~m[48]&m[49]&m[51]&m[52])|(m[42]&~m[48]&m[49]&m[51]&m[52])|(m[42]&m[48]&m[49]&m[51]&m[52]));
    m[55] = (((m[47]&~m[53]&~m[54]&~m[56]&~m[57])|(~m[47]&~m[53]&~m[54]&m[56]&~m[57])|(m[47]&m[53]&~m[54]&m[56]&~m[57])|(m[47]&~m[53]&m[54]&m[56]&~m[57])|(~m[47]&m[53]&~m[54]&~m[56]&m[57])|(~m[47]&~m[53]&m[54]&~m[56]&m[57])|(m[47]&m[53]&m[54]&~m[56]&m[57])|(~m[47]&m[53]&m[54]&m[56]&m[57]))&UnbiasedRNG[13])|((m[47]&~m[53]&~m[54]&m[56]&~m[57])|(~m[47]&~m[53]&~m[54]&~m[56]&m[57])|(m[47]&~m[53]&~m[54]&~m[56]&m[57])|(m[47]&m[53]&~m[54]&~m[56]&m[57])|(m[47]&~m[53]&m[54]&~m[56]&m[57])|(~m[47]&~m[53]&~m[54]&m[56]&m[57])|(m[47]&~m[53]&~m[54]&m[56]&m[57])|(~m[47]&m[53]&~m[54]&m[56]&m[57])|(m[47]&m[53]&~m[54]&m[56]&m[57])|(~m[47]&~m[53]&m[54]&m[56]&m[57])|(m[47]&~m[53]&m[54]&m[56]&m[57])|(m[47]&m[53]&m[54]&m[56]&m[57]));
    m[60] = (((m[57]&~m[58]&~m[59]&~m[61]&~m[62])|(~m[57]&~m[58]&~m[59]&m[61]&~m[62])|(m[57]&m[58]&~m[59]&m[61]&~m[62])|(m[57]&~m[58]&m[59]&m[61]&~m[62])|(~m[57]&m[58]&~m[59]&~m[61]&m[62])|(~m[57]&~m[58]&m[59]&~m[61]&m[62])|(m[57]&m[58]&m[59]&~m[61]&m[62])|(~m[57]&m[58]&m[59]&m[61]&m[62]))&UnbiasedRNG[14])|((m[57]&~m[58]&~m[59]&m[61]&~m[62])|(~m[57]&~m[58]&~m[59]&~m[61]&m[62])|(m[57]&~m[58]&~m[59]&~m[61]&m[62])|(m[57]&m[58]&~m[59]&~m[61]&m[62])|(m[57]&~m[58]&m[59]&~m[61]&m[62])|(~m[57]&~m[58]&~m[59]&m[61]&m[62])|(m[57]&~m[58]&~m[59]&m[61]&m[62])|(~m[57]&m[58]&~m[59]&m[61]&m[62])|(m[57]&m[58]&~m[59]&m[61]&m[62])|(~m[57]&~m[58]&m[59]&m[61]&m[62])|(m[57]&~m[58]&m[59]&m[61]&m[62])|(m[57]&m[58]&m[59]&m[61]&m[62]));
end

always @(posedge color3_clk) begin
    m[41] = (((m[38]&~m[39]&~m[40]&~m[42]&~m[43])|(~m[38]&m[39]&~m[40]&~m[42]&~m[43])|(~m[38]&~m[39]&m[40]&~m[42]&~m[43])|(m[38]&m[39]&m[40]&m[42]&~m[43])|(~m[38]&~m[39]&~m[40]&~m[42]&m[43])|(m[38]&m[39]&~m[40]&m[42]&m[43])|(m[38]&~m[39]&m[40]&m[42]&m[43])|(~m[38]&m[39]&m[40]&m[42]&m[43]))&UnbiasedRNG[15])|((m[38]&m[39]&~m[40]&~m[42]&~m[43])|(m[38]&~m[39]&m[40]&~m[42]&~m[43])|(~m[38]&m[39]&m[40]&~m[42]&~m[43])|(m[38]&m[39]&m[40]&~m[42]&~m[43])|(m[38]&~m[39]&~m[40]&~m[42]&m[43])|(~m[38]&m[39]&~m[40]&~m[42]&m[43])|(m[38]&m[39]&~m[40]&~m[42]&m[43])|(~m[38]&~m[39]&m[40]&~m[42]&m[43])|(m[38]&~m[39]&m[40]&~m[42]&m[43])|(~m[38]&m[39]&m[40]&~m[42]&m[43])|(m[38]&m[39]&m[40]&~m[42]&m[43])|(m[38]&m[39]&m[40]&m[42]&m[43]));
    m[51] = (((m[48]&~m[49]&~m[50]&~m[52]&~m[53])|(~m[48]&m[49]&~m[50]&~m[52]&~m[53])|(~m[48]&~m[49]&m[50]&~m[52]&~m[53])|(m[48]&m[49]&m[50]&m[52]&~m[53])|(~m[48]&~m[49]&~m[50]&~m[52]&m[53])|(m[48]&m[49]&~m[50]&m[52]&m[53])|(m[48]&~m[49]&m[50]&m[52]&m[53])|(~m[48]&m[49]&m[50]&m[52]&m[53]))&UnbiasedRNG[16])|((m[48]&m[49]&~m[50]&~m[52]&~m[53])|(m[48]&~m[49]&m[50]&~m[52]&~m[53])|(~m[48]&m[49]&m[50]&~m[52]&~m[53])|(m[48]&m[49]&m[50]&~m[52]&~m[53])|(m[48]&~m[49]&~m[50]&~m[52]&m[53])|(~m[48]&m[49]&~m[50]&~m[52]&m[53])|(m[48]&m[49]&~m[50]&~m[52]&m[53])|(~m[48]&~m[49]&m[50]&~m[52]&m[53])|(m[48]&~m[49]&m[50]&~m[52]&m[53])|(~m[48]&m[49]&m[50]&~m[52]&m[53])|(m[48]&m[49]&m[50]&~m[52]&m[53])|(m[48]&m[49]&m[50]&m[52]&m[53]));
end

always @(posedge color4_clk) begin
    m[37] = (((m[33]&~m[34]&~m[35]&~m[36]&~m[40])|(~m[33]&m[34]&~m[35]&~m[36]&~m[40])|(~m[33]&~m[34]&m[35]&~m[36]&~m[40])|(m[33]&m[34]&~m[35]&m[36]&~m[40])|(m[33]&~m[34]&m[35]&m[36]&~m[40])|(~m[33]&m[34]&m[35]&m[36]&~m[40]))&BiasedRNG[32])|(((m[33]&~m[34]&~m[35]&~m[36]&m[40])|(~m[33]&m[34]&~m[35]&~m[36]&m[40])|(~m[33]&~m[34]&m[35]&~m[36]&m[40])|(m[33]&m[34]&~m[35]&m[36]&m[40])|(m[33]&~m[34]&m[35]&m[36]&m[40])|(~m[33]&m[34]&m[35]&m[36]&m[40]))&~BiasedRNG[32])|((m[33]&m[34]&~m[35]&~m[36]&~m[40])|(m[33]&~m[34]&m[35]&~m[36]&~m[40])|(~m[33]&m[34]&m[35]&~m[36]&~m[40])|(m[33]&m[34]&m[35]&~m[36]&~m[40])|(m[33]&m[34]&m[35]&m[36]&~m[40])|(m[33]&m[34]&~m[35]&~m[36]&m[40])|(m[33]&~m[34]&m[35]&~m[36]&m[40])|(~m[33]&m[34]&m[35]&~m[36]&m[40])|(m[33]&m[34]&m[35]&~m[36]&m[40])|(m[33]&m[34]&m[35]&m[36]&m[40]));
    m[42] = (((m[38]&~m[39]&~m[40]&~m[41]&~m[50])|(~m[38]&m[39]&~m[40]&~m[41]&~m[50])|(~m[38]&~m[39]&m[40]&~m[41]&~m[50])|(m[38]&m[39]&~m[40]&m[41]&~m[50])|(m[38]&~m[39]&m[40]&m[41]&~m[50])|(~m[38]&m[39]&m[40]&m[41]&~m[50]))&BiasedRNG[33])|(((m[38]&~m[39]&~m[40]&~m[41]&m[50])|(~m[38]&m[39]&~m[40]&~m[41]&m[50])|(~m[38]&~m[39]&m[40]&~m[41]&m[50])|(m[38]&m[39]&~m[40]&m[41]&m[50])|(m[38]&~m[39]&m[40]&m[41]&m[50])|(~m[38]&m[39]&m[40]&m[41]&m[50]))&~BiasedRNG[33])|((m[38]&m[39]&~m[40]&~m[41]&~m[50])|(m[38]&~m[39]&m[40]&~m[41]&~m[50])|(~m[38]&m[39]&m[40]&~m[41]&~m[50])|(m[38]&m[39]&m[40]&~m[41]&~m[50])|(m[38]&m[39]&m[40]&m[41]&~m[50])|(m[38]&m[39]&~m[40]&~m[41]&m[50])|(m[38]&~m[39]&m[40]&~m[41]&m[50])|(~m[38]&m[39]&m[40]&~m[41]&m[50])|(m[38]&m[39]&m[40]&~m[41]&m[50])|(m[38]&m[39]&m[40]&m[41]&m[50]));
    m[47] = (((m[43]&~m[44]&~m[45]&~m[46]&~m[55])|(~m[43]&m[44]&~m[45]&~m[46]&~m[55])|(~m[43]&~m[44]&m[45]&~m[46]&~m[55])|(m[43]&m[44]&~m[45]&m[46]&~m[55])|(m[43]&~m[44]&m[45]&m[46]&~m[55])|(~m[43]&m[44]&m[45]&m[46]&~m[55]))&BiasedRNG[34])|(((m[43]&~m[44]&~m[45]&~m[46]&m[55])|(~m[43]&m[44]&~m[45]&~m[46]&m[55])|(~m[43]&~m[44]&m[45]&~m[46]&m[55])|(m[43]&m[44]&~m[45]&m[46]&m[55])|(m[43]&~m[44]&m[45]&m[46]&m[55])|(~m[43]&m[44]&m[45]&m[46]&m[55]))&~BiasedRNG[34])|((m[43]&m[44]&~m[45]&~m[46]&~m[55])|(m[43]&~m[44]&m[45]&~m[46]&~m[55])|(~m[43]&m[44]&m[45]&~m[46]&~m[55])|(m[43]&m[44]&m[45]&~m[46]&~m[55])|(m[43]&m[44]&m[45]&m[46]&~m[55])|(m[43]&m[44]&~m[45]&~m[46]&m[55])|(m[43]&~m[44]&m[45]&~m[46]&m[55])|(~m[43]&m[44]&m[45]&~m[46]&m[55])|(m[43]&m[44]&m[45]&~m[46]&m[55])|(m[43]&m[44]&m[45]&m[46]&m[55]));
    m[52] = (((m[48]&~m[49]&~m[50]&~m[51]&~m[58])|(~m[48]&m[49]&~m[50]&~m[51]&~m[58])|(~m[48]&~m[49]&m[50]&~m[51]&~m[58])|(m[48]&m[49]&~m[50]&m[51]&~m[58])|(m[48]&~m[49]&m[50]&m[51]&~m[58])|(~m[48]&m[49]&m[50]&m[51]&~m[58]))&BiasedRNG[35])|(((m[48]&~m[49]&~m[50]&~m[51]&m[58])|(~m[48]&m[49]&~m[50]&~m[51]&m[58])|(~m[48]&~m[49]&m[50]&~m[51]&m[58])|(m[48]&m[49]&~m[50]&m[51]&m[58])|(m[48]&~m[49]&m[50]&m[51]&m[58])|(~m[48]&m[49]&m[50]&m[51]&m[58]))&~BiasedRNG[35])|((m[48]&m[49]&~m[50]&~m[51]&~m[58])|(m[48]&~m[49]&m[50]&~m[51]&~m[58])|(~m[48]&m[49]&m[50]&~m[51]&~m[58])|(m[48]&m[49]&m[50]&~m[51]&~m[58])|(m[48]&m[49]&m[50]&m[51]&~m[58])|(m[48]&m[49]&~m[50]&~m[51]&m[58])|(m[48]&~m[49]&m[50]&~m[51]&m[58])|(~m[48]&m[49]&m[50]&~m[51]&m[58])|(m[48]&m[49]&m[50]&~m[51]&m[58])|(m[48]&m[49]&m[50]&m[51]&m[58]));
    m[57] = (((m[53]&~m[54]&~m[55]&~m[56]&~m[60])|(~m[53]&m[54]&~m[55]&~m[56]&~m[60])|(~m[53]&~m[54]&m[55]&~m[56]&~m[60])|(m[53]&m[54]&~m[55]&m[56]&~m[60])|(m[53]&~m[54]&m[55]&m[56]&~m[60])|(~m[53]&m[54]&m[55]&m[56]&~m[60]))&BiasedRNG[36])|(((m[53]&~m[54]&~m[55]&~m[56]&m[60])|(~m[53]&m[54]&~m[55]&~m[56]&m[60])|(~m[53]&~m[54]&m[55]&~m[56]&m[60])|(m[53]&m[54]&~m[55]&m[56]&m[60])|(m[53]&~m[54]&m[55]&m[56]&m[60])|(~m[53]&m[54]&m[55]&m[56]&m[60]))&~BiasedRNG[36])|((m[53]&m[54]&~m[55]&~m[56]&~m[60])|(m[53]&~m[54]&m[55]&~m[56]&~m[60])|(~m[53]&m[54]&m[55]&~m[56]&~m[60])|(m[53]&m[54]&m[55]&~m[56]&~m[60])|(m[53]&m[54]&m[55]&m[56]&~m[60])|(m[53]&m[54]&~m[55]&~m[56]&m[60])|(m[53]&~m[54]&m[55]&~m[56]&m[60])|(~m[53]&m[54]&m[55]&~m[56]&m[60])|(m[53]&m[54]&m[55]&~m[56]&m[60])|(m[53]&m[54]&m[55]&m[56]&m[60]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[70]&LFSRcolor0[40]&LFSRcolor0[6]&LFSRcolor0[19]);
    BiasedRNG[1] = (LFSRcolor0[52]&LFSRcolor0[8]&LFSRcolor0[76]&LFSRcolor0[77]);
    BiasedRNG[2] = (LFSRcolor0[27]&LFSRcolor0[59]&LFSRcolor0[69]&LFSRcolor0[64]);
    BiasedRNG[3] = (LFSRcolor0[65]&LFSRcolor0[26]&LFSRcolor0[62]&LFSRcolor0[82]);
    BiasedRNG[4] = (LFSRcolor0[83]&LFSRcolor0[10]&LFSRcolor0[13]&LFSRcolor0[1]);
    BiasedRNG[5] = (LFSRcolor0[25]&LFSRcolor0[0]&LFSRcolor0[28]&LFSRcolor0[89]);
    BiasedRNG[6] = (LFSRcolor0[86]&LFSRcolor0[47]&LFSRcolor0[20]&LFSRcolor0[75]);
    BiasedRNG[7] = (LFSRcolor0[33]&LFSRcolor0[9]&LFSRcolor0[39]&LFSRcolor0[90]);
    BiasedRNG[8] = (LFSRcolor0[71]&LFSRcolor0[84]&LFSRcolor0[21]&LFSRcolor0[51]);
    BiasedRNG[9] = (LFSRcolor0[66]&LFSRcolor0[73]&LFSRcolor0[85]&LFSRcolor0[12]);
    BiasedRNG[10] = (LFSRcolor0[87]&LFSRcolor0[41]&LFSRcolor0[46]&LFSRcolor0[4]);
    BiasedRNG[11] = (LFSRcolor0[68]&LFSRcolor0[16]&LFSRcolor0[79]&LFSRcolor0[53]);
    BiasedRNG[12] = (LFSRcolor0[29]&LFSRcolor0[57]&LFSRcolor0[58]&LFSRcolor0[17]);
    BiasedRNG[13] = (LFSRcolor0[81]&LFSRcolor0[32]&LFSRcolor0[45]&LFSRcolor0[67]);
    UnbiasedRNG[0] = LFSRcolor0[15];
    UnbiasedRNG[1] = LFSRcolor0[5];
    UnbiasedRNG[2] = LFSRcolor0[63];
    UnbiasedRNG[3] = LFSRcolor0[74];
end

always @(posedge color0_clk) begin
    BiasedRNG[14] = (LFSRcolor1[13]&LFSRcolor1[28]&LFSRcolor1[44]&LFSRcolor1[32]);
    BiasedRNG[15] = (LFSRcolor1[42]&LFSRcolor1[10]&LFSRcolor1[15]&LFSRcolor1[27]);
    BiasedRNG[16] = (LFSRcolor1[8]&LFSRcolor1[19]&LFSRcolor1[11]&LFSRcolor1[23]);
    BiasedRNG[17] = (LFSRcolor1[7]&LFSRcolor1[40]&LFSRcolor1[41]&LFSRcolor1[4]);
    BiasedRNG[18] = (LFSRcolor1[31]&LFSRcolor1[24]&LFSRcolor1[2]&LFSRcolor1[22]);
    BiasedRNG[19] = (LFSRcolor1[17]&LFSRcolor1[35]&LFSRcolor1[37]&LFSRcolor1[5]);
    BiasedRNG[20] = (LFSRcolor1[29]&LFSRcolor1[38]&LFSRcolor1[30]&LFSRcolor1[33]);
    BiasedRNG[21] = (LFSRcolor1[43]&LFSRcolor1[1]&LFSRcolor1[21]&LFSRcolor1[20]);
    BiasedRNG[22] = (LFSRcolor1[26]&LFSRcolor1[34]&LFSRcolor1[45]&LFSRcolor1[9]);
    UnbiasedRNG[4] = LFSRcolor1[12];
    UnbiasedRNG[5] = LFSRcolor1[3];
    UnbiasedRNG[6] = LFSRcolor1[25];
    UnbiasedRNG[7] = LFSRcolor1[39];
    UnbiasedRNG[8] = LFSRcolor1[16];
    UnbiasedRNG[9] = LFSRcolor1[0];
end

always @(posedge color1_clk) begin
    BiasedRNG[23] = (LFSRcolor2[23]&LFSRcolor2[15]&LFSRcolor2[0]&LFSRcolor2[20]);
    BiasedRNG[24] = (LFSRcolor2[16]&LFSRcolor2[37]&LFSRcolor2[9]&LFSRcolor2[6]);
    BiasedRNG[25] = (LFSRcolor2[25]&LFSRcolor2[29]&LFSRcolor2[3]&LFSRcolor2[14]);
    BiasedRNG[26] = (LFSRcolor2[8]&LFSRcolor2[28]&LFSRcolor2[21]&LFSRcolor2[24]);
    BiasedRNG[27] = (LFSRcolor2[18]&LFSRcolor2[38]&LFSRcolor2[43]&LFSRcolor2[5]);
    BiasedRNG[28] = (LFSRcolor2[2]&LFSRcolor2[35]&LFSRcolor2[34]&LFSRcolor2[32]);
    BiasedRNG[29] = (LFSRcolor2[26]&LFSRcolor2[11]&LFSRcolor2[13]&LFSRcolor2[40]);
    BiasedRNG[30] = (LFSRcolor2[44]&LFSRcolor2[17]&LFSRcolor2[12]&LFSRcolor2[30]);
    BiasedRNG[31] = (LFSRcolor2[10]&LFSRcolor2[4]&LFSRcolor2[42]&LFSRcolor2[45]);
    UnbiasedRNG[10] = LFSRcolor2[19];
    UnbiasedRNG[11] = LFSRcolor2[31];
    UnbiasedRNG[12] = LFSRcolor2[41];
    UnbiasedRNG[13] = LFSRcolor2[22];
    UnbiasedRNG[14] = LFSRcolor2[27];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[15] = LFSRcolor3[11];
    UnbiasedRNG[16] = LFSRcolor3[1];
end

always @(posedge color3_clk) begin
    BiasedRNG[32] = (LFSRcolor4[28]&LFSRcolor4[34]&LFSRcolor4[0]&LFSRcolor4[43]);
    BiasedRNG[33] = (LFSRcolor4[12]&LFSRcolor4[45]&LFSRcolor4[39]&LFSRcolor4[13]);
    BiasedRNG[34] = (LFSRcolor4[11]&LFSRcolor4[21]&LFSRcolor4[6]&LFSRcolor4[36]);
    BiasedRNG[35] = (LFSRcolor4[33]&LFSRcolor4[8]&LFSRcolor4[41]&LFSRcolor4[16]);
    BiasedRNG[36] = (LFSRcolor4[40]&LFSRcolor4[4]&LFSRcolor4[22]&LFSRcolor4[29]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule