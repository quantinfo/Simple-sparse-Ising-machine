//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [19:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [505:0] LFSRcolor0;
wire [689:0] LFSRcolor1;
wire [505:0] LFSRcolor2;
wire [91:0] LFSRcolor3;
wire [367:0] LFSRcolor4;
reg [427:0] BiasedRNG;       //For I=+/-1 cases
reg [351:0] UnbiasedRNG;   //For I=0 cases
reg [0:809] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[260] = 1'b1;
initial m[363] = 1'b1;
initial m[373] = 1'b1;
initial m[388] = 1'b1;
initial m[408] = 1'b0;
initial m[433] = 1'b1;
initial m[463] = 1'b1;
initial m[498] = 1'b1;
initial m[538] = 1'b1;
initial m[583] = 1'b0;
initial m[628] = 1'b0;
initial m[668] = 1'b0;
initial m[703] = 1'b0;
initial m[733] = 1'b0;
initial m[758] = 1'b1;
initial m[778] = 1'b0;
initial m[793] = 1'b1;
initial m[803] = 1'b1;
initial m[808] = 1'b1;
initial m[809] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[362] = 1'b0;
initial m[372] = 1'b0;
initial m[387] = 1'b0;
initial m[407] = 1'b0;
initial m[432] = 1'b0;
initial m[462] = 1'b0;
initial m[497] = 1'b0;
initial m[537] = 1'b0;
initial m[582] = 1'b0;
initial m[585] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 0;
initial m[1] = 0;
initial m[2] = 1;
initial m[3] = 1;
initial m[4] = 0;
initial m[5] = 0;
initial m[6] = 1;
initial m[7] = 0;
initial m[8] = 0;
initial m[9] = 0;
initial m[10] = 0;
initial m[11] = 1;
initial m[12] = 0;
initial m[13] = 0;
initial m[14] = 0;
initial m[15] = 1;
initial m[16] = 0;
initial m[17] = 0;
initial m[18] = 1;
initial m[19] = 1;
initial m[20] = 1;
initial m[21] = 1;
initial m[22] = 0;
initial m[23] = 0;
initial m[24] = 1;
initial m[25] = 1;
initial m[26] = 1;
initial m[27] = 0;
initial m[28] = 1;
initial m[29] = 0;
initial m[30] = 1;
initial m[31] = 1;
initial m[32] = 1;
initial m[33] = 1;
initial m[34] = 0;
initial m[35] = 1;
initial m[36] = 1;
initial m[37] = 1;
initial m[38] = 1;
initial m[39] = 1;
initial m[40] = 0;
initial m[41] = 0;
initial m[42] = 0;
initial m[43] = 1;
initial m[44] = 1;
initial m[45] = 0;
initial m[46] = 0;
initial m[47] = 1;
initial m[48] = 0;
initial m[49] = 1;
initial m[50] = 0;
initial m[51] = 0;
initial m[52] = 0;
initial m[53] = 1;
initial m[54] = 1;
initial m[55] = 0;
initial m[56] = 1;
initial m[57] = 0;
initial m[58] = 0;
initial m[59] = 0;
initial m[60] = 0;
initial m[61] = 0;
initial m[62] = 0;
initial m[63] = 1;
initial m[64] = 0;
initial m[65] = 1;
initial m[66] = 0;
initial m[67] = 1;
initial m[68] = 0;
initial m[69] = 0;
initial m[70] = 1;
initial m[71] = 0;
initial m[72] = 0;
initial m[73] = 0;
initial m[74] = 0;
initial m[75] = 1;
initial m[76] = 0;
initial m[77] = 0;
initial m[78] = 0;
initial m[79] = 0;
initial m[80] = 1;
initial m[81] = 0;
initial m[82] = 1;
initial m[83] = 1;
initial m[84] = 0;
initial m[85] = 1;
initial m[86] = 1;
initial m[87] = 0;
initial m[88] = 0;
initial m[89] = 1;
initial m[90] = 1;
initial m[91] = 0;
initial m[92] = 1;
initial m[93] = 1;
initial m[94] = 1;
initial m[95] = 0;
initial m[96] = 0;
initial m[97] = 1;
initial m[98] = 1;
initial m[99] = 0;
initial m[100] = 1;
initial m[101] = 0;
initial m[102] = 0;
initial m[103] = 1;
initial m[104] = 0;
initial m[105] = 0;
initial m[106] = 1;
initial m[107] = 1;
initial m[108] = 0;
initial m[109] = 0;
initial m[110] = 1;
initial m[111] = 0;
initial m[112] = 1;
initial m[113] = 0;
initial m[114] = 1;
initial m[115] = 1;
initial m[116] = 1;
initial m[117] = 0;
initial m[118] = 1;
initial m[119] = 0;
initial m[120] = 1;
initial m[121] = 0;
initial m[122] = 0;
initial m[123] = 1;
initial m[124] = 0;
initial m[125] = 1;
initial m[126] = 1;
initial m[127] = 1;
initial m[128] = 1;
initial m[129] = 1;
initial m[130] = 1;
initial m[131] = 1;
initial m[132] = 1;
initial m[133] = 0;
initial m[134] = 0;
initial m[135] = 0;
initial m[136] = 0;
initial m[137] = 0;
initial m[138] = 1;
initial m[139] = 0;
initial m[140] = 0;
initial m[141] = 1;
initial m[142] = 1;
initial m[143] = 1;
initial m[144] = 1;
initial m[145] = 0;
initial m[146] = 0;
initial m[147] = 0;
initial m[148] = 0;
initial m[149] = 1;
initial m[150] = 0;
initial m[151] = 1;
initial m[152] = 0;
initial m[153] = 0;
initial m[154] = 1;
initial m[155] = 0;
initial m[156] = 0;
initial m[157] = 0;
initial m[158] = 0;
initial m[159] = 1;
initial m[160] = 1;
initial m[161] = 0;
initial m[162] = 0;
initial m[163] = 0;
initial m[164] = 1;
initial m[165] = 0;
initial m[166] = 1;
initial m[167] = 1;
initial m[168] = 0;
initial m[169] = 0;
initial m[170] = 0;
initial m[171] = 0;
initial m[172] = 0;
initial m[173] = 0;
initial m[174] = 1;
initial m[175] = 1;
initial m[176] = 1;
initial m[177] = 1;
initial m[178] = 1;
initial m[179] = 0;
initial m[180] = 1;
initial m[181] = 0;
initial m[182] = 1;
initial m[183] = 1;
initial m[184] = 0;
initial m[185] = 0;
initial m[186] = 1;
initial m[187] = 1;
initial m[188] = 1;
initial m[189] = 0;
initial m[190] = 1;
initial m[191] = 0;
initial m[192] = 0;
initial m[193] = 1;
initial m[194] = 1;
initial m[195] = 1;
initial m[196] = 1;
initial m[197] = 1;
initial m[198] = 0;
initial m[199] = 0;
initial m[200] = 1;
initial m[201] = 1;
initial m[202] = 0;
initial m[203] = 1;
initial m[204] = 1;
initial m[205] = 1;
initial m[206] = 0;
initial m[207] = 0;
initial m[208] = 0;
initial m[209] = 0;
initial m[210] = 0;
initial m[211] = 0;
initial m[212] = 0;
initial m[213] = 1;
initial m[214] = 0;
initial m[215] = 0;
initial m[216] = 0;
initial m[217] = 0;
initial m[218] = 1;
initial m[219] = 0;
initial m[220] = 1;
initial m[221] = 1;
initial m[222] = 0;
initial m[223] = 0;
initial m[224] = 1;
initial m[225] = 1;
initial m[226] = 1;
initial m[227] = 1;
initial m[228] = 1;
initial m[229] = 0;
initial m[230] = 1;
initial m[231] = 0;
initial m[232] = 1;
initial m[233] = 0;
initial m[234] = 1;
initial m[235] = 1;
initial m[236] = 1;
initial m[237] = 0;
initial m[238] = 1;
initial m[239] = 0;
initial m[240] = 0;
initial m[241] = 0;
initial m[242] = 1;
initial m[243] = 1;
initial m[244] = 0;
initial m[245] = 0;
initial m[246] = 0;
initial m[247] = 0;
initial m[248] = 1;
initial m[249] = 1;
initial m[250] = 0;
initial m[251] = 0;
initial m[252] = 0;
initial m[253] = 1;
initial m[254] = 0;
initial m[255] = 1;
initial m[256] = 1;
initial m[257] = 0;
initial m[258] = 0;
initial m[259] = 1;
initial m[261] = 0;
initial m[262] = 0;
initial m[263] = 1;
initial m[264] = 1;
initial m[265] = 1;
initial m[266] = 0;
initial m[267] = 0;
initial m[268] = 1;
initial m[269] = 0;
initial m[270] = 0;
initial m[271] = 1;
initial m[272] = 0;
initial m[273] = 1;
initial m[274] = 1;
initial m[275] = 0;
initial m[276] = 0;
initial m[277] = 1;
initial m[278] = 1;
initial m[279] = 0;
initial m[280] = 1;
initial m[281] = 0;
initial m[282] = 1;
initial m[283] = 0;
initial m[284] = 0;
initial m[285] = 0;
initial m[286] = 0;
initial m[287] = 1;
initial m[288] = 1;
initial m[289] = 0;
initial m[290] = 0;
initial m[291] = 0;
initial m[292] = 1;
initial m[293] = 0;
initial m[294] = 0;
initial m[295] = 0;
initial m[296] = 0;
initial m[297] = 0;
initial m[298] = 1;
initial m[299] = 0;
initial m[300] = 1;
initial m[301] = 1;
initial m[302] = 0;
initial m[303] = 1;
initial m[304] = 0;
initial m[305] = 1;
initial m[306] = 1;
initial m[307] = 0;
initial m[308] = 1;
initial m[309] = 0;
initial m[310] = 0;
initial m[311] = 0;
initial m[312] = 1;
initial m[313] = 0;
initial m[314] = 0;
initial m[315] = 0;
initial m[316] = 0;
initial m[317] = 1;
initial m[318] = 1;
initial m[319] = 0;
initial m[320] = 1;
initial m[321] = 0;
initial m[322] = 1;
initial m[323] = 0;
initial m[324] = 1;
initial m[325] = 1;
initial m[326] = 1;
initial m[327] = 1;
initial m[328] = 1;
initial m[329] = 1;
initial m[330] = 0;
initial m[331] = 0;
initial m[332] = 0;
initial m[333] = 0;
initial m[334] = 0;
initial m[335] = 1;
initial m[336] = 0;
initial m[337] = 0;
initial m[338] = 1;
initial m[339] = 0;
initial m[340] = 1;
initial m[341] = 0;
initial m[342] = 0;
initial m[343] = 0;
initial m[344] = 1;
initial m[345] = 1;
initial m[346] = 0;
initial m[347] = 0;
initial m[348] = 0;
initial m[349] = 1;
initial m[350] = 1;
initial m[351] = 0;
initial m[352] = 0;
initial m[353] = 1;
initial m[354] = 1;
initial m[355] = 1;
initial m[356] = 0;
initial m[357] = 1;
initial m[358] = 1;
initial m[359] = 0;
initial m[360] = 1;
initial m[361] = 0;
initial m[364] = 1;
initial m[365] = 1;
initial m[366] = 0;
initial m[367] = 1;
initial m[368] = 0;
initial m[369] = 0;
initial m[370] = 1;
initial m[371] = 0;
initial m[374] = 1;
initial m[375] = 1;
initial m[376] = 1;
initial m[377] = 0;
initial m[378] = 1;
initial m[379] = 1;
initial m[380] = 1;
initial m[381] = 1;
initial m[382] = 0;
initial m[383] = 1;
initial m[384] = 0;
initial m[385] = 1;
initial m[386] = 1;
initial m[389] = 0;
initial m[390] = 0;
initial m[391] = 1;
initial m[392] = 0;
initial m[393] = 0;
initial m[394] = 0;
initial m[395] = 0;
initial m[396] = 1;
initial m[397] = 1;
initial m[398] = 1;
initial m[399] = 1;
initial m[400] = 0;
initial m[401] = 0;
initial m[402] = 0;
initial m[403] = 0;
initial m[404] = 0;
initial m[405] = 1;
initial m[406] = 0;
initial m[409] = 0;
initial m[410] = 1;
initial m[411] = 1;
initial m[412] = 1;
initial m[413] = 1;
initial m[414] = 0;
initial m[415] = 0;
initial m[416] = 1;
initial m[417] = 0;
initial m[418] = 1;
initial m[419] = 0;
initial m[420] = 0;
initial m[421] = 1;
initial m[422] = 0;
initial m[423] = 0;
initial m[424] = 1;
initial m[425] = 1;
initial m[426] = 0;
initial m[427] = 0;
initial m[428] = 1;
initial m[429] = 0;
initial m[430] = 0;
initial m[431] = 0;
initial m[434] = 1;
initial m[435] = 0;
initial m[436] = 1;
initial m[437] = 1;
initial m[438] = 0;
initial m[439] = 1;
initial m[440] = 1;
initial m[441] = 1;
initial m[442] = 1;
initial m[443] = 1;
initial m[444] = 1;
initial m[445] = 0;
initial m[446] = 0;
initial m[447] = 0;
initial m[448] = 0;
initial m[449] = 0;
initial m[450] = 0;
initial m[451] = 0;
initial m[452] = 0;
initial m[453] = 1;
initial m[454] = 1;
initial m[455] = 0;
initial m[456] = 0;
initial m[457] = 1;
initial m[458] = 1;
initial m[459] = 0;
initial m[460] = 1;
initial m[461] = 1;
initial m[464] = 1;
initial m[465] = 1;
initial m[466] = 0;
initial m[467] = 0;
initial m[468] = 0;
initial m[469] = 0;
initial m[470] = 1;
initial m[471] = 0;
initial m[472] = 0;
initial m[473] = 1;
initial m[474] = 1;
initial m[475] = 0;
initial m[476] = 0;
initial m[477] = 1;
initial m[478] = 0;
initial m[479] = 1;
initial m[480] = 1;
initial m[481] = 0;
initial m[482] = 1;
initial m[483] = 0;
initial m[484] = 0;
initial m[485] = 1;
initial m[486] = 0;
initial m[487] = 0;
initial m[488] = 1;
initial m[489] = 1;
initial m[490] = 1;
initial m[491] = 0;
initial m[492] = 0;
initial m[493] = 1;
initial m[494] = 0;
initial m[495] = 0;
initial m[496] = 1;
initial m[499] = 1;
initial m[500] = 1;
initial m[501] = 0;
initial m[502] = 1;
initial m[503] = 1;
initial m[504] = 1;
initial m[505] = 0;
initial m[506] = 0;
initial m[507] = 0;
initial m[508] = 0;
initial m[509] = 0;
initial m[510] = 0;
initial m[511] = 1;
initial m[512] = 1;
initial m[513] = 1;
initial m[514] = 0;
initial m[515] = 1;
initial m[516] = 1;
initial m[517] = 1;
initial m[518] = 1;
initial m[519] = 1;
initial m[520] = 1;
initial m[521] = 1;
initial m[522] = 1;
initial m[523] = 1;
initial m[524] = 0;
initial m[525] = 0;
initial m[526] = 1;
initial m[527] = 0;
initial m[528] = 1;
initial m[529] = 0;
initial m[530] = 0;
initial m[531] = 0;
initial m[532] = 0;
initial m[533] = 0;
initial m[534] = 0;
initial m[535] = 1;
initial m[536] = 1;
initial m[539] = 1;
initial m[540] = 0;
initial m[541] = 0;
initial m[542] = 1;
initial m[543] = 1;
initial m[544] = 1;
initial m[545] = 1;
initial m[546] = 1;
initial m[547] = 0;
initial m[548] = 0;
initial m[549] = 1;
initial m[550] = 1;
initial m[551] = 0;
initial m[552] = 0;
initial m[553] = 0;
initial m[554] = 0;
initial m[555] = 0;
initial m[556] = 1;
initial m[557] = 0;
initial m[558] = 0;
initial m[559] = 1;
initial m[560] = 0;
initial m[561] = 0;
initial m[562] = 0;
initial m[563] = 0;
initial m[564] = 0;
initial m[565] = 0;
initial m[566] = 1;
initial m[567] = 0;
initial m[568] = 1;
initial m[569] = 1;
initial m[570] = 1;
initial m[571] = 0;
initial m[572] = 0;
initial m[573] = 1;
initial m[574] = 1;
initial m[575] = 1;
initial m[576] = 1;
initial m[577] = 1;
initial m[578] = 0;
initial m[579] = 1;
initial m[580] = 1;
initial m[581] = 1;
initial m[584] = 1;
initial m[586] = 1;
initial m[587] = 0;
initial m[588] = 0;
initial m[589] = 0;
initial m[590] = 0;
initial m[591] = 1;
initial m[592] = 0;
initial m[593] = 1;
initial m[594] = 1;
initial m[595] = 1;
initial m[596] = 0;
initial m[597] = 1;
initial m[598] = 0;
initial m[599] = 1;
initial m[600] = 0;
initial m[601] = 1;
initial m[602] = 0;
initial m[603] = 1;
initial m[604] = 1;
initial m[605] = 1;
initial m[606] = 1;
initial m[607] = 1;
initial m[608] = 1;
initial m[609] = 0;
initial m[610] = 1;
initial m[611] = 0;
initial m[612] = 1;
initial m[613] = 0;
initial m[614] = 1;
initial m[615] = 0;
initial m[616] = 0;
initial m[617] = 0;
initial m[618] = 1;
initial m[619] = 1;
initial m[620] = 0;
initial m[621] = 1;
initial m[622] = 1;
initial m[623] = 0;
initial m[624] = 1;
initial m[625] = 0;
initial m[626] = 0;
initial m[627] = 0;
initial m[629] = 1;
initial m[630] = 1;
initial m[631] = 0;
initial m[632] = 1;
initial m[633] = 1;
initial m[634] = 1;
initial m[635] = 0;
initial m[636] = 0;
initial m[637] = 1;
initial m[638] = 1;
initial m[639] = 1;
initial m[640] = 0;
initial m[641] = 1;
initial m[642] = 1;
initial m[643] = 1;
initial m[644] = 1;
initial m[645] = 1;
initial m[646] = 1;
initial m[647] = 0;
initial m[648] = 1;
initial m[649] = 1;
initial m[650] = 0;
initial m[651] = 1;
initial m[652] = 1;
initial m[653] = 1;
initial m[654] = 0;
initial m[655] = 0;
initial m[656] = 0;
initial m[657] = 1;
initial m[658] = 1;
initial m[659] = 1;
initial m[660] = 1;
initial m[661] = 1;
initial m[662] = 1;
initial m[663] = 0;
initial m[664] = 1;
initial m[665] = 1;
initial m[666] = 0;
initial m[667] = 1;
initial m[669] = 1;
initial m[670] = 1;
initial m[671] = 0;
initial m[672] = 0;
initial m[673] = 1;
initial m[674] = 1;
initial m[675] = 1;
initial m[676] = 1;
initial m[677] = 0;
initial m[678] = 1;
initial m[679] = 0;
initial m[680] = 1;
initial m[681] = 1;
initial m[682] = 1;
initial m[683] = 1;
initial m[684] = 0;
initial m[685] = 0;
initial m[686] = 0;
initial m[687] = 0;
initial m[688] = 0;
initial m[689] = 0;
initial m[690] = 1;
initial m[691] = 1;
initial m[692] = 0;
initial m[693] = 1;
initial m[694] = 1;
initial m[695] = 1;
initial m[696] = 1;
initial m[697] = 1;
initial m[698] = 0;
initial m[699] = 0;
initial m[700] = 0;
initial m[701] = 0;
initial m[702] = 1;
initial m[704] = 1;
initial m[705] = 1;
initial m[706] = 1;
initial m[707] = 1;
initial m[708] = 0;
initial m[709] = 0;
initial m[710] = 0;
initial m[711] = 1;
initial m[712] = 1;
initial m[713] = 1;
initial m[714] = 0;
initial m[715] = 0;
initial m[716] = 0;
initial m[717] = 0;
initial m[718] = 1;
initial m[719] = 1;
initial m[720] = 1;
initial m[721] = 0;
initial m[722] = 1;
initial m[723] = 0;
initial m[724] = 1;
initial m[725] = 0;
initial m[726] = 1;
initial m[727] = 0;
initial m[728] = 0;
initial m[729] = 1;
initial m[730] = 1;
initial m[731] = 0;
initial m[732] = 1;
initial m[734] = 1;
initial m[735] = 1;
initial m[736] = 0;
initial m[737] = 1;
initial m[738] = 0;
initial m[739] = 0;
initial m[740] = 0;
initial m[741] = 0;
initial m[742] = 0;
initial m[743] = 0;
initial m[744] = 0;
initial m[745] = 1;
initial m[746] = 1;
initial m[747] = 1;
initial m[748] = 0;
initial m[749] = 0;
initial m[750] = 0;
initial m[751] = 1;
initial m[752] = 1;
initial m[753] = 1;
initial m[754] = 0;
initial m[755] = 1;
initial m[756] = 0;
initial m[757] = 1;
initial m[759] = 1;
initial m[760] = 1;
initial m[761] = 0;
initial m[762] = 0;
initial m[763] = 1;
initial m[764] = 1;
initial m[765] = 0;
initial m[766] = 0;
initial m[767] = 1;
initial m[768] = 0;
initial m[769] = 0;
initial m[770] = 1;
initial m[771] = 1;
initial m[772] = 0;
initial m[773] = 1;
initial m[774] = 1;
initial m[775] = 0;
initial m[776] = 0;
initial m[777] = 1;
initial m[779] = 0;
initial m[780] = 1;
initial m[781] = 1;
initial m[782] = 1;
initial m[783] = 0;
initial m[784] = 1;
initial m[785] = 1;
initial m[786] = 0;
initial m[787] = 0;
initial m[788] = 0;
initial m[789] = 1;
initial m[790] = 0;
initial m[791] = 1;
initial m[792] = 1;
initial m[794] = 1;
initial m[795] = 0;
initial m[796] = 0;
initial m[797] = 1;
initial m[798] = 0;
initial m[799] = 0;
initial m[800] = 1;
initial m[801] = 0;
initial m[802] = 0;
initial m[804] = 1;
initial m[805] = 1;
initial m[806] = 0;
initial m[807] = 0;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[19],m[18],m[17],m[16],m[15],m[14],m[13],m[12],m[11],m[10]};
end

always @(negedge sample_clk) begin
    if (solution == 20'b11110100000111101111)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[20]&m[21]&~m[60]&~m[61])|(m[20]&~m[21]&m[60]&~m[61])|(~m[20]&m[21]&m[60]&~m[61])|(m[20]&~m[21]&~m[60]&m[61])|(~m[20]&m[21]&~m[60]&m[61])|(~m[20]&~m[21]&m[60]&m[61]))&UnbiasedRNG[0])|((m[20]&m[21]&m[60]&~m[61])|(m[20]&m[21]&~m[60]&m[61])|(m[20]&~m[21]&m[60]&m[61])|(~m[20]&m[21]&m[60]&m[61])|(m[20]&m[21]&m[60]&m[61]));
    m[1] = (((m[22]&m[23]&~m[70]&~m[71])|(m[22]&~m[23]&m[70]&~m[71])|(~m[22]&m[23]&m[70]&~m[71])|(m[22]&~m[23]&~m[70]&m[71])|(~m[22]&m[23]&~m[70]&m[71])|(~m[22]&~m[23]&m[70]&m[71]))&UnbiasedRNG[1])|((m[22]&m[23]&m[70]&~m[71])|(m[22]&m[23]&~m[70]&m[71])|(m[22]&~m[23]&m[70]&m[71])|(~m[22]&m[23]&m[70]&m[71])|(m[22]&m[23]&m[70]&m[71]));
    m[2] = (((m[24]&m[25]&~m[80]&~m[81])|(m[24]&~m[25]&m[80]&~m[81])|(~m[24]&m[25]&m[80]&~m[81])|(m[24]&~m[25]&~m[80]&m[81])|(~m[24]&m[25]&~m[80]&m[81])|(~m[24]&~m[25]&m[80]&m[81]))&UnbiasedRNG[2])|((m[24]&m[25]&m[80]&~m[81])|(m[24]&m[25]&~m[80]&m[81])|(m[24]&~m[25]&m[80]&m[81])|(~m[24]&m[25]&m[80]&m[81])|(m[24]&m[25]&m[80]&m[81]));
    m[3] = (((m[26]&m[27]&~m[90]&~m[91])|(m[26]&~m[27]&m[90]&~m[91])|(~m[26]&m[27]&m[90]&~m[91])|(m[26]&~m[27]&~m[90]&m[91])|(~m[26]&m[27]&~m[90]&m[91])|(~m[26]&~m[27]&m[90]&m[91]))&UnbiasedRNG[3])|((m[26]&m[27]&m[90]&~m[91])|(m[26]&m[27]&~m[90]&m[91])|(m[26]&~m[27]&m[90]&m[91])|(~m[26]&m[27]&m[90]&m[91])|(m[26]&m[27]&m[90]&m[91]));
    m[4] = (((m[28]&m[29]&~m[100]&~m[101])|(m[28]&~m[29]&m[100]&~m[101])|(~m[28]&m[29]&m[100]&~m[101])|(m[28]&~m[29]&~m[100]&m[101])|(~m[28]&m[29]&~m[100]&m[101])|(~m[28]&~m[29]&m[100]&m[101]))&UnbiasedRNG[4])|((m[28]&m[29]&m[100]&~m[101])|(m[28]&m[29]&~m[100]&m[101])|(m[28]&~m[29]&m[100]&m[101])|(~m[28]&m[29]&m[100]&m[101])|(m[28]&m[29]&m[100]&m[101]));
    m[5] = (((m[30]&m[31]&~m[110]&~m[111])|(m[30]&~m[31]&m[110]&~m[111])|(~m[30]&m[31]&m[110]&~m[111])|(m[30]&~m[31]&~m[110]&m[111])|(~m[30]&m[31]&~m[110]&m[111])|(~m[30]&~m[31]&m[110]&m[111]))&UnbiasedRNG[5])|((m[30]&m[31]&m[110]&~m[111])|(m[30]&m[31]&~m[110]&m[111])|(m[30]&~m[31]&m[110]&m[111])|(~m[30]&m[31]&m[110]&m[111])|(m[30]&m[31]&m[110]&m[111]));
    m[6] = (((m[32]&m[33]&~m[120]&~m[121])|(m[32]&~m[33]&m[120]&~m[121])|(~m[32]&m[33]&m[120]&~m[121])|(m[32]&~m[33]&~m[120]&m[121])|(~m[32]&m[33]&~m[120]&m[121])|(~m[32]&~m[33]&m[120]&m[121]))&UnbiasedRNG[6])|((m[32]&m[33]&m[120]&~m[121])|(m[32]&m[33]&~m[120]&m[121])|(m[32]&~m[33]&m[120]&m[121])|(~m[32]&m[33]&m[120]&m[121])|(m[32]&m[33]&m[120]&m[121]));
    m[7] = (((m[34]&m[35]&~m[130]&~m[131])|(m[34]&~m[35]&m[130]&~m[131])|(~m[34]&m[35]&m[130]&~m[131])|(m[34]&~m[35]&~m[130]&m[131])|(~m[34]&m[35]&~m[130]&m[131])|(~m[34]&~m[35]&m[130]&m[131]))&UnbiasedRNG[7])|((m[34]&m[35]&m[130]&~m[131])|(m[34]&m[35]&~m[130]&m[131])|(m[34]&~m[35]&m[130]&m[131])|(~m[34]&m[35]&m[130]&m[131])|(m[34]&m[35]&m[130]&m[131]));
    m[8] = (((m[36]&m[37]&~m[140]&~m[141])|(m[36]&~m[37]&m[140]&~m[141])|(~m[36]&m[37]&m[140]&~m[141])|(m[36]&~m[37]&~m[140]&m[141])|(~m[36]&m[37]&~m[140]&m[141])|(~m[36]&~m[37]&m[140]&m[141]))&UnbiasedRNG[8])|((m[36]&m[37]&m[140]&~m[141])|(m[36]&m[37]&~m[140]&m[141])|(m[36]&~m[37]&m[140]&m[141])|(~m[36]&m[37]&m[140]&m[141])|(m[36]&m[37]&m[140]&m[141]));
    m[9] = (((m[38]&m[39]&~m[150]&~m[151])|(m[38]&~m[39]&m[150]&~m[151])|(~m[38]&m[39]&m[150]&~m[151])|(m[38]&~m[39]&~m[150]&m[151])|(~m[38]&m[39]&~m[150]&m[151])|(~m[38]&~m[39]&m[150]&m[151]))&UnbiasedRNG[9])|((m[38]&m[39]&m[150]&~m[151])|(m[38]&m[39]&~m[150]&m[151])|(m[38]&~m[39]&m[150]&m[151])|(~m[38]&m[39]&m[150]&m[151])|(m[38]&m[39]&m[150]&m[151]));
    m[10] = (((m[40]&m[41]&~m[160]&~m[161])|(m[40]&~m[41]&m[160]&~m[161])|(~m[40]&m[41]&m[160]&~m[161])|(m[40]&~m[41]&~m[160]&m[161])|(~m[40]&m[41]&~m[160]&m[161])|(~m[40]&~m[41]&m[160]&m[161]))&UnbiasedRNG[10])|((m[40]&m[41]&m[160]&~m[161])|(m[40]&m[41]&~m[160]&m[161])|(m[40]&~m[41]&m[160]&m[161])|(~m[40]&m[41]&m[160]&m[161])|(m[40]&m[41]&m[160]&m[161]));
    m[11] = (((m[42]&m[43]&~m[170]&~m[171])|(m[42]&~m[43]&m[170]&~m[171])|(~m[42]&m[43]&m[170]&~m[171])|(m[42]&~m[43]&~m[170]&m[171])|(~m[42]&m[43]&~m[170]&m[171])|(~m[42]&~m[43]&m[170]&m[171]))&UnbiasedRNG[11])|((m[42]&m[43]&m[170]&~m[171])|(m[42]&m[43]&~m[170]&m[171])|(m[42]&~m[43]&m[170]&m[171])|(~m[42]&m[43]&m[170]&m[171])|(m[42]&m[43]&m[170]&m[171]));
    m[12] = (((m[44]&m[45]&~m[180]&~m[181])|(m[44]&~m[45]&m[180]&~m[181])|(~m[44]&m[45]&m[180]&~m[181])|(m[44]&~m[45]&~m[180]&m[181])|(~m[44]&m[45]&~m[180]&m[181])|(~m[44]&~m[45]&m[180]&m[181]))&UnbiasedRNG[12])|((m[44]&m[45]&m[180]&~m[181])|(m[44]&m[45]&~m[180]&m[181])|(m[44]&~m[45]&m[180]&m[181])|(~m[44]&m[45]&m[180]&m[181])|(m[44]&m[45]&m[180]&m[181]));
    m[13] = (((m[46]&m[47]&~m[190]&~m[191])|(m[46]&~m[47]&m[190]&~m[191])|(~m[46]&m[47]&m[190]&~m[191])|(m[46]&~m[47]&~m[190]&m[191])|(~m[46]&m[47]&~m[190]&m[191])|(~m[46]&~m[47]&m[190]&m[191]))&UnbiasedRNG[13])|((m[46]&m[47]&m[190]&~m[191])|(m[46]&m[47]&~m[190]&m[191])|(m[46]&~m[47]&m[190]&m[191])|(~m[46]&m[47]&m[190]&m[191])|(m[46]&m[47]&m[190]&m[191]));
    m[14] = (((m[48]&m[49]&~m[200]&~m[201])|(m[48]&~m[49]&m[200]&~m[201])|(~m[48]&m[49]&m[200]&~m[201])|(m[48]&~m[49]&~m[200]&m[201])|(~m[48]&m[49]&~m[200]&m[201])|(~m[48]&~m[49]&m[200]&m[201]))&UnbiasedRNG[14])|((m[48]&m[49]&m[200]&~m[201])|(m[48]&m[49]&~m[200]&m[201])|(m[48]&~m[49]&m[200]&m[201])|(~m[48]&m[49]&m[200]&m[201])|(m[48]&m[49]&m[200]&m[201]));
    m[15] = (((m[50]&m[51]&~m[210]&~m[211])|(m[50]&~m[51]&m[210]&~m[211])|(~m[50]&m[51]&m[210]&~m[211])|(m[50]&~m[51]&~m[210]&m[211])|(~m[50]&m[51]&~m[210]&m[211])|(~m[50]&~m[51]&m[210]&m[211]))&UnbiasedRNG[15])|((m[50]&m[51]&m[210]&~m[211])|(m[50]&m[51]&~m[210]&m[211])|(m[50]&~m[51]&m[210]&m[211])|(~m[50]&m[51]&m[210]&m[211])|(m[50]&m[51]&m[210]&m[211]));
    m[16] = (((m[52]&m[53]&~m[220]&~m[221])|(m[52]&~m[53]&m[220]&~m[221])|(~m[52]&m[53]&m[220]&~m[221])|(m[52]&~m[53]&~m[220]&m[221])|(~m[52]&m[53]&~m[220]&m[221])|(~m[52]&~m[53]&m[220]&m[221]))&UnbiasedRNG[16])|((m[52]&m[53]&m[220]&~m[221])|(m[52]&m[53]&~m[220]&m[221])|(m[52]&~m[53]&m[220]&m[221])|(~m[52]&m[53]&m[220]&m[221])|(m[52]&m[53]&m[220]&m[221]));
    m[17] = (((m[54]&m[55]&~m[230]&~m[231])|(m[54]&~m[55]&m[230]&~m[231])|(~m[54]&m[55]&m[230]&~m[231])|(m[54]&~m[55]&~m[230]&m[231])|(~m[54]&m[55]&~m[230]&m[231])|(~m[54]&~m[55]&m[230]&m[231]))&UnbiasedRNG[17])|((m[54]&m[55]&m[230]&~m[231])|(m[54]&m[55]&~m[230]&m[231])|(m[54]&~m[55]&m[230]&m[231])|(~m[54]&m[55]&m[230]&m[231])|(m[54]&m[55]&m[230]&m[231]));
    m[18] = (((m[56]&m[57]&~m[240]&~m[241])|(m[56]&~m[57]&m[240]&~m[241])|(~m[56]&m[57]&m[240]&~m[241])|(m[56]&~m[57]&~m[240]&m[241])|(~m[56]&m[57]&~m[240]&m[241])|(~m[56]&~m[57]&m[240]&m[241]))&UnbiasedRNG[18])|((m[56]&m[57]&m[240]&~m[241])|(m[56]&m[57]&~m[240]&m[241])|(m[56]&~m[57]&m[240]&m[241])|(~m[56]&m[57]&m[240]&m[241])|(m[56]&m[57]&m[240]&m[241]));
    m[19] = (((m[58]&m[59]&~m[250]&~m[251])|(m[58]&~m[59]&m[250]&~m[251])|(~m[58]&m[59]&m[250]&~m[251])|(m[58]&~m[59]&~m[250]&m[251])|(~m[58]&m[59]&~m[250]&m[251])|(~m[58]&~m[59]&m[250]&m[251]))&UnbiasedRNG[19])|((m[58]&m[59]&m[250]&~m[251])|(m[58]&m[59]&~m[250]&m[251])|(m[58]&~m[59]&m[250]&m[251])|(~m[58]&m[59]&m[250]&m[251])|(m[58]&m[59]&m[250]&m[251]));
    m[62] = (((~m[20]&~m[180]&~m[280])|(m[20]&m[180]&~m[280]))&BiasedRNG[0])|(((m[20]&~m[180]&~m[280])|(~m[20]&m[180]&m[280]))&~BiasedRNG[0])|((~m[20]&~m[180]&m[280])|(m[20]&~m[180]&m[280])|(m[20]&m[180]&m[280]));
    m[63] = (((~m[20]&~m[190]&~m[290])|(m[20]&m[190]&~m[290]))&BiasedRNG[1])|(((m[20]&~m[190]&~m[290])|(~m[20]&m[190]&m[290]))&~BiasedRNG[1])|((~m[20]&~m[190]&m[290])|(m[20]&~m[190]&m[290])|(m[20]&m[190]&m[290]));
    m[64] = (((~m[20]&~m[200]&~m[300])|(m[20]&m[200]&~m[300]))&BiasedRNG[2])|(((m[20]&~m[200]&~m[300])|(~m[20]&m[200]&m[300]))&~BiasedRNG[2])|((~m[20]&~m[200]&m[300])|(m[20]&~m[200]&m[300])|(m[20]&m[200]&m[300]));
    m[65] = (((~m[20]&~m[210]&~m[310])|(m[20]&m[210]&~m[310]))&BiasedRNG[3])|(((m[20]&~m[210]&~m[310])|(~m[20]&m[210]&m[310]))&~BiasedRNG[3])|((~m[20]&~m[210]&m[310])|(m[20]&~m[210]&m[310])|(m[20]&m[210]&m[310]));
    m[66] = (((~m[21]&~m[220]&~m[320])|(m[21]&m[220]&~m[320]))&BiasedRNG[4])|(((m[21]&~m[220]&~m[320])|(~m[21]&m[220]&m[320]))&~BiasedRNG[4])|((~m[21]&~m[220]&m[320])|(m[21]&~m[220]&m[320])|(m[21]&m[220]&m[320]));
    m[67] = (((~m[21]&~m[230]&~m[330])|(m[21]&m[230]&~m[330]))&BiasedRNG[5])|(((m[21]&~m[230]&~m[330])|(~m[21]&m[230]&m[330]))&~BiasedRNG[5])|((~m[21]&~m[230]&m[330])|(m[21]&~m[230]&m[330])|(m[21]&m[230]&m[330]));
    m[68] = (((~m[21]&~m[240]&~m[340])|(m[21]&m[240]&~m[340]))&BiasedRNG[6])|(((m[21]&~m[240]&~m[340])|(~m[21]&m[240]&m[340]))&~BiasedRNG[6])|((~m[21]&~m[240]&m[340])|(m[21]&~m[240]&m[340])|(m[21]&m[240]&m[340]));
    m[69] = (((~m[21]&~m[250]&~m[350])|(m[21]&m[250]&~m[350]))&BiasedRNG[7])|(((m[21]&~m[250]&~m[350])|(~m[21]&m[250]&m[350]))&~BiasedRNG[7])|((~m[21]&~m[250]&m[350])|(m[21]&~m[250]&m[350])|(m[21]&m[250]&m[350]));
    m[72] = (((~m[22]&~m[181]&~m[281])|(m[22]&m[181]&~m[281]))&BiasedRNG[8])|(((m[22]&~m[181]&~m[281])|(~m[22]&m[181]&m[281]))&~BiasedRNG[8])|((~m[22]&~m[181]&m[281])|(m[22]&~m[181]&m[281])|(m[22]&m[181]&m[281]));
    m[73] = (((~m[22]&~m[191]&~m[291])|(m[22]&m[191]&~m[291]))&BiasedRNG[9])|(((m[22]&~m[191]&~m[291])|(~m[22]&m[191]&m[291]))&~BiasedRNG[9])|((~m[22]&~m[191]&m[291])|(m[22]&~m[191]&m[291])|(m[22]&m[191]&m[291]));
    m[74] = (((~m[22]&~m[201]&~m[301])|(m[22]&m[201]&~m[301]))&BiasedRNG[10])|(((m[22]&~m[201]&~m[301])|(~m[22]&m[201]&m[301]))&~BiasedRNG[10])|((~m[22]&~m[201]&m[301])|(m[22]&~m[201]&m[301])|(m[22]&m[201]&m[301]));
    m[75] = (((~m[22]&~m[211]&~m[311])|(m[22]&m[211]&~m[311]))&BiasedRNG[11])|(((m[22]&~m[211]&~m[311])|(~m[22]&m[211]&m[311]))&~BiasedRNG[11])|((~m[22]&~m[211]&m[311])|(m[22]&~m[211]&m[311])|(m[22]&m[211]&m[311]));
    m[76] = (((~m[23]&~m[221]&~m[321])|(m[23]&m[221]&~m[321]))&BiasedRNG[12])|(((m[23]&~m[221]&~m[321])|(~m[23]&m[221]&m[321]))&~BiasedRNG[12])|((~m[23]&~m[221]&m[321])|(m[23]&~m[221]&m[321])|(m[23]&m[221]&m[321]));
    m[77] = (((~m[23]&~m[231]&~m[331])|(m[23]&m[231]&~m[331]))&BiasedRNG[13])|(((m[23]&~m[231]&~m[331])|(~m[23]&m[231]&m[331]))&~BiasedRNG[13])|((~m[23]&~m[231]&m[331])|(m[23]&~m[231]&m[331])|(m[23]&m[231]&m[331]));
    m[78] = (((~m[23]&~m[241]&~m[341])|(m[23]&m[241]&~m[341]))&BiasedRNG[14])|(((m[23]&~m[241]&~m[341])|(~m[23]&m[241]&m[341]))&~BiasedRNG[14])|((~m[23]&~m[241]&m[341])|(m[23]&~m[241]&m[341])|(m[23]&m[241]&m[341]));
    m[79] = (((~m[23]&~m[251]&~m[351])|(m[23]&m[251]&~m[351]))&BiasedRNG[15])|(((m[23]&~m[251]&~m[351])|(~m[23]&m[251]&m[351]))&~BiasedRNG[15])|((~m[23]&~m[251]&m[351])|(m[23]&~m[251]&m[351])|(m[23]&m[251]&m[351]));
    m[82] = (((~m[24]&~m[182]&~m[282])|(m[24]&m[182]&~m[282]))&BiasedRNG[16])|(((m[24]&~m[182]&~m[282])|(~m[24]&m[182]&m[282]))&~BiasedRNG[16])|((~m[24]&~m[182]&m[282])|(m[24]&~m[182]&m[282])|(m[24]&m[182]&m[282]));
    m[83] = (((~m[24]&~m[192]&~m[292])|(m[24]&m[192]&~m[292]))&BiasedRNG[17])|(((m[24]&~m[192]&~m[292])|(~m[24]&m[192]&m[292]))&~BiasedRNG[17])|((~m[24]&~m[192]&m[292])|(m[24]&~m[192]&m[292])|(m[24]&m[192]&m[292]));
    m[84] = (((~m[24]&~m[202]&~m[302])|(m[24]&m[202]&~m[302]))&BiasedRNG[18])|(((m[24]&~m[202]&~m[302])|(~m[24]&m[202]&m[302]))&~BiasedRNG[18])|((~m[24]&~m[202]&m[302])|(m[24]&~m[202]&m[302])|(m[24]&m[202]&m[302]));
    m[85] = (((~m[24]&~m[212]&~m[312])|(m[24]&m[212]&~m[312]))&BiasedRNG[19])|(((m[24]&~m[212]&~m[312])|(~m[24]&m[212]&m[312]))&~BiasedRNG[19])|((~m[24]&~m[212]&m[312])|(m[24]&~m[212]&m[312])|(m[24]&m[212]&m[312]));
    m[86] = (((~m[25]&~m[222]&~m[322])|(m[25]&m[222]&~m[322]))&BiasedRNG[20])|(((m[25]&~m[222]&~m[322])|(~m[25]&m[222]&m[322]))&~BiasedRNG[20])|((~m[25]&~m[222]&m[322])|(m[25]&~m[222]&m[322])|(m[25]&m[222]&m[322]));
    m[87] = (((~m[25]&~m[232]&~m[332])|(m[25]&m[232]&~m[332]))&BiasedRNG[21])|(((m[25]&~m[232]&~m[332])|(~m[25]&m[232]&m[332]))&~BiasedRNG[21])|((~m[25]&~m[232]&m[332])|(m[25]&~m[232]&m[332])|(m[25]&m[232]&m[332]));
    m[88] = (((~m[25]&~m[242]&~m[342])|(m[25]&m[242]&~m[342]))&BiasedRNG[22])|(((m[25]&~m[242]&~m[342])|(~m[25]&m[242]&m[342]))&~BiasedRNG[22])|((~m[25]&~m[242]&m[342])|(m[25]&~m[242]&m[342])|(m[25]&m[242]&m[342]));
    m[89] = (((~m[25]&~m[252]&~m[352])|(m[25]&m[252]&~m[352]))&BiasedRNG[23])|(((m[25]&~m[252]&~m[352])|(~m[25]&m[252]&m[352]))&~BiasedRNG[23])|((~m[25]&~m[252]&m[352])|(m[25]&~m[252]&m[352])|(m[25]&m[252]&m[352]));
    m[92] = (((~m[26]&~m[183]&~m[283])|(m[26]&m[183]&~m[283]))&BiasedRNG[24])|(((m[26]&~m[183]&~m[283])|(~m[26]&m[183]&m[283]))&~BiasedRNG[24])|((~m[26]&~m[183]&m[283])|(m[26]&~m[183]&m[283])|(m[26]&m[183]&m[283]));
    m[93] = (((~m[26]&~m[193]&~m[293])|(m[26]&m[193]&~m[293]))&BiasedRNG[25])|(((m[26]&~m[193]&~m[293])|(~m[26]&m[193]&m[293]))&~BiasedRNG[25])|((~m[26]&~m[193]&m[293])|(m[26]&~m[193]&m[293])|(m[26]&m[193]&m[293]));
    m[94] = (((~m[26]&~m[203]&~m[303])|(m[26]&m[203]&~m[303]))&BiasedRNG[26])|(((m[26]&~m[203]&~m[303])|(~m[26]&m[203]&m[303]))&~BiasedRNG[26])|((~m[26]&~m[203]&m[303])|(m[26]&~m[203]&m[303])|(m[26]&m[203]&m[303]));
    m[95] = (((~m[26]&~m[213]&~m[313])|(m[26]&m[213]&~m[313]))&BiasedRNG[27])|(((m[26]&~m[213]&~m[313])|(~m[26]&m[213]&m[313]))&~BiasedRNG[27])|((~m[26]&~m[213]&m[313])|(m[26]&~m[213]&m[313])|(m[26]&m[213]&m[313]));
    m[96] = (((~m[27]&~m[223]&~m[323])|(m[27]&m[223]&~m[323]))&BiasedRNG[28])|(((m[27]&~m[223]&~m[323])|(~m[27]&m[223]&m[323]))&~BiasedRNG[28])|((~m[27]&~m[223]&m[323])|(m[27]&~m[223]&m[323])|(m[27]&m[223]&m[323]));
    m[97] = (((~m[27]&~m[233]&~m[333])|(m[27]&m[233]&~m[333]))&BiasedRNG[29])|(((m[27]&~m[233]&~m[333])|(~m[27]&m[233]&m[333]))&~BiasedRNG[29])|((~m[27]&~m[233]&m[333])|(m[27]&~m[233]&m[333])|(m[27]&m[233]&m[333]));
    m[98] = (((~m[27]&~m[243]&~m[343])|(m[27]&m[243]&~m[343]))&BiasedRNG[30])|(((m[27]&~m[243]&~m[343])|(~m[27]&m[243]&m[343]))&~BiasedRNG[30])|((~m[27]&~m[243]&m[343])|(m[27]&~m[243]&m[343])|(m[27]&m[243]&m[343]));
    m[99] = (((~m[27]&~m[253]&~m[353])|(m[27]&m[253]&~m[353]))&BiasedRNG[31])|(((m[27]&~m[253]&~m[353])|(~m[27]&m[253]&m[353]))&~BiasedRNG[31])|((~m[27]&~m[253]&m[353])|(m[27]&~m[253]&m[353])|(m[27]&m[253]&m[353]));
    m[102] = (((~m[28]&~m[184]&~m[284])|(m[28]&m[184]&~m[284]))&BiasedRNG[32])|(((m[28]&~m[184]&~m[284])|(~m[28]&m[184]&m[284]))&~BiasedRNG[32])|((~m[28]&~m[184]&m[284])|(m[28]&~m[184]&m[284])|(m[28]&m[184]&m[284]));
    m[103] = (((~m[28]&~m[194]&~m[294])|(m[28]&m[194]&~m[294]))&BiasedRNG[33])|(((m[28]&~m[194]&~m[294])|(~m[28]&m[194]&m[294]))&~BiasedRNG[33])|((~m[28]&~m[194]&m[294])|(m[28]&~m[194]&m[294])|(m[28]&m[194]&m[294]));
    m[104] = (((~m[28]&~m[204]&~m[304])|(m[28]&m[204]&~m[304]))&BiasedRNG[34])|(((m[28]&~m[204]&~m[304])|(~m[28]&m[204]&m[304]))&~BiasedRNG[34])|((~m[28]&~m[204]&m[304])|(m[28]&~m[204]&m[304])|(m[28]&m[204]&m[304]));
    m[105] = (((~m[28]&~m[214]&~m[314])|(m[28]&m[214]&~m[314]))&BiasedRNG[35])|(((m[28]&~m[214]&~m[314])|(~m[28]&m[214]&m[314]))&~BiasedRNG[35])|((~m[28]&~m[214]&m[314])|(m[28]&~m[214]&m[314])|(m[28]&m[214]&m[314]));
    m[106] = (((~m[29]&~m[224]&~m[324])|(m[29]&m[224]&~m[324]))&BiasedRNG[36])|(((m[29]&~m[224]&~m[324])|(~m[29]&m[224]&m[324]))&~BiasedRNG[36])|((~m[29]&~m[224]&m[324])|(m[29]&~m[224]&m[324])|(m[29]&m[224]&m[324]));
    m[107] = (((~m[29]&~m[234]&~m[334])|(m[29]&m[234]&~m[334]))&BiasedRNG[37])|(((m[29]&~m[234]&~m[334])|(~m[29]&m[234]&m[334]))&~BiasedRNG[37])|((~m[29]&~m[234]&m[334])|(m[29]&~m[234]&m[334])|(m[29]&m[234]&m[334]));
    m[108] = (((~m[29]&~m[244]&~m[344])|(m[29]&m[244]&~m[344]))&BiasedRNG[38])|(((m[29]&~m[244]&~m[344])|(~m[29]&m[244]&m[344]))&~BiasedRNG[38])|((~m[29]&~m[244]&m[344])|(m[29]&~m[244]&m[344])|(m[29]&m[244]&m[344]));
    m[109] = (((~m[29]&~m[254]&~m[354])|(m[29]&m[254]&~m[354]))&BiasedRNG[39])|(((m[29]&~m[254]&~m[354])|(~m[29]&m[254]&m[354]))&~BiasedRNG[39])|((~m[29]&~m[254]&m[354])|(m[29]&~m[254]&m[354])|(m[29]&m[254]&m[354]));
    m[112] = (((~m[30]&~m[185]&~m[285])|(m[30]&m[185]&~m[285]))&BiasedRNG[40])|(((m[30]&~m[185]&~m[285])|(~m[30]&m[185]&m[285]))&~BiasedRNG[40])|((~m[30]&~m[185]&m[285])|(m[30]&~m[185]&m[285])|(m[30]&m[185]&m[285]));
    m[113] = (((~m[30]&~m[195]&~m[295])|(m[30]&m[195]&~m[295]))&BiasedRNG[41])|(((m[30]&~m[195]&~m[295])|(~m[30]&m[195]&m[295]))&~BiasedRNG[41])|((~m[30]&~m[195]&m[295])|(m[30]&~m[195]&m[295])|(m[30]&m[195]&m[295]));
    m[114] = (((~m[30]&~m[205]&~m[305])|(m[30]&m[205]&~m[305]))&BiasedRNG[42])|(((m[30]&~m[205]&~m[305])|(~m[30]&m[205]&m[305]))&~BiasedRNG[42])|((~m[30]&~m[205]&m[305])|(m[30]&~m[205]&m[305])|(m[30]&m[205]&m[305]));
    m[115] = (((~m[30]&~m[215]&~m[315])|(m[30]&m[215]&~m[315]))&BiasedRNG[43])|(((m[30]&~m[215]&~m[315])|(~m[30]&m[215]&m[315]))&~BiasedRNG[43])|((~m[30]&~m[215]&m[315])|(m[30]&~m[215]&m[315])|(m[30]&m[215]&m[315]));
    m[116] = (((~m[31]&~m[225]&~m[325])|(m[31]&m[225]&~m[325]))&BiasedRNG[44])|(((m[31]&~m[225]&~m[325])|(~m[31]&m[225]&m[325]))&~BiasedRNG[44])|((~m[31]&~m[225]&m[325])|(m[31]&~m[225]&m[325])|(m[31]&m[225]&m[325]));
    m[117] = (((~m[31]&~m[235]&~m[335])|(m[31]&m[235]&~m[335]))&BiasedRNG[45])|(((m[31]&~m[235]&~m[335])|(~m[31]&m[235]&m[335]))&~BiasedRNG[45])|((~m[31]&~m[235]&m[335])|(m[31]&~m[235]&m[335])|(m[31]&m[235]&m[335]));
    m[118] = (((~m[31]&~m[245]&~m[345])|(m[31]&m[245]&~m[345]))&BiasedRNG[46])|(((m[31]&~m[245]&~m[345])|(~m[31]&m[245]&m[345]))&~BiasedRNG[46])|((~m[31]&~m[245]&m[345])|(m[31]&~m[245]&m[345])|(m[31]&m[245]&m[345]));
    m[119] = (((~m[31]&~m[255]&~m[355])|(m[31]&m[255]&~m[355]))&BiasedRNG[47])|(((m[31]&~m[255]&~m[355])|(~m[31]&m[255]&m[355]))&~BiasedRNG[47])|((~m[31]&~m[255]&m[355])|(m[31]&~m[255]&m[355])|(m[31]&m[255]&m[355]));
    m[122] = (((~m[32]&~m[186]&~m[286])|(m[32]&m[186]&~m[286]))&BiasedRNG[48])|(((m[32]&~m[186]&~m[286])|(~m[32]&m[186]&m[286]))&~BiasedRNG[48])|((~m[32]&~m[186]&m[286])|(m[32]&~m[186]&m[286])|(m[32]&m[186]&m[286]));
    m[123] = (((~m[32]&~m[196]&~m[296])|(m[32]&m[196]&~m[296]))&BiasedRNG[49])|(((m[32]&~m[196]&~m[296])|(~m[32]&m[196]&m[296]))&~BiasedRNG[49])|((~m[32]&~m[196]&m[296])|(m[32]&~m[196]&m[296])|(m[32]&m[196]&m[296]));
    m[124] = (((~m[32]&~m[206]&~m[306])|(m[32]&m[206]&~m[306]))&BiasedRNG[50])|(((m[32]&~m[206]&~m[306])|(~m[32]&m[206]&m[306]))&~BiasedRNG[50])|((~m[32]&~m[206]&m[306])|(m[32]&~m[206]&m[306])|(m[32]&m[206]&m[306]));
    m[125] = (((~m[32]&~m[216]&~m[316])|(m[32]&m[216]&~m[316]))&BiasedRNG[51])|(((m[32]&~m[216]&~m[316])|(~m[32]&m[216]&m[316]))&~BiasedRNG[51])|((~m[32]&~m[216]&m[316])|(m[32]&~m[216]&m[316])|(m[32]&m[216]&m[316]));
    m[126] = (((~m[33]&~m[226]&~m[326])|(m[33]&m[226]&~m[326]))&BiasedRNG[52])|(((m[33]&~m[226]&~m[326])|(~m[33]&m[226]&m[326]))&~BiasedRNG[52])|((~m[33]&~m[226]&m[326])|(m[33]&~m[226]&m[326])|(m[33]&m[226]&m[326]));
    m[127] = (((~m[33]&~m[236]&~m[336])|(m[33]&m[236]&~m[336]))&BiasedRNG[53])|(((m[33]&~m[236]&~m[336])|(~m[33]&m[236]&m[336]))&~BiasedRNG[53])|((~m[33]&~m[236]&m[336])|(m[33]&~m[236]&m[336])|(m[33]&m[236]&m[336]));
    m[128] = (((~m[33]&~m[246]&~m[346])|(m[33]&m[246]&~m[346]))&BiasedRNG[54])|(((m[33]&~m[246]&~m[346])|(~m[33]&m[246]&m[346]))&~BiasedRNG[54])|((~m[33]&~m[246]&m[346])|(m[33]&~m[246]&m[346])|(m[33]&m[246]&m[346]));
    m[129] = (((~m[33]&~m[256]&~m[356])|(m[33]&m[256]&~m[356]))&BiasedRNG[55])|(((m[33]&~m[256]&~m[356])|(~m[33]&m[256]&m[356]))&~BiasedRNG[55])|((~m[33]&~m[256]&m[356])|(m[33]&~m[256]&m[356])|(m[33]&m[256]&m[356]));
    m[132] = (((~m[34]&~m[187]&~m[287])|(m[34]&m[187]&~m[287]))&BiasedRNG[56])|(((m[34]&~m[187]&~m[287])|(~m[34]&m[187]&m[287]))&~BiasedRNG[56])|((~m[34]&~m[187]&m[287])|(m[34]&~m[187]&m[287])|(m[34]&m[187]&m[287]));
    m[133] = (((~m[34]&~m[197]&~m[297])|(m[34]&m[197]&~m[297]))&BiasedRNG[57])|(((m[34]&~m[197]&~m[297])|(~m[34]&m[197]&m[297]))&~BiasedRNG[57])|((~m[34]&~m[197]&m[297])|(m[34]&~m[197]&m[297])|(m[34]&m[197]&m[297]));
    m[134] = (((~m[34]&~m[207]&~m[307])|(m[34]&m[207]&~m[307]))&BiasedRNG[58])|(((m[34]&~m[207]&~m[307])|(~m[34]&m[207]&m[307]))&~BiasedRNG[58])|((~m[34]&~m[207]&m[307])|(m[34]&~m[207]&m[307])|(m[34]&m[207]&m[307]));
    m[135] = (((~m[34]&~m[217]&~m[317])|(m[34]&m[217]&~m[317]))&BiasedRNG[59])|(((m[34]&~m[217]&~m[317])|(~m[34]&m[217]&m[317]))&~BiasedRNG[59])|((~m[34]&~m[217]&m[317])|(m[34]&~m[217]&m[317])|(m[34]&m[217]&m[317]));
    m[136] = (((~m[35]&~m[227]&~m[327])|(m[35]&m[227]&~m[327]))&BiasedRNG[60])|(((m[35]&~m[227]&~m[327])|(~m[35]&m[227]&m[327]))&~BiasedRNG[60])|((~m[35]&~m[227]&m[327])|(m[35]&~m[227]&m[327])|(m[35]&m[227]&m[327]));
    m[137] = (((~m[35]&~m[237]&~m[337])|(m[35]&m[237]&~m[337]))&BiasedRNG[61])|(((m[35]&~m[237]&~m[337])|(~m[35]&m[237]&m[337]))&~BiasedRNG[61])|((~m[35]&~m[237]&m[337])|(m[35]&~m[237]&m[337])|(m[35]&m[237]&m[337]));
    m[138] = (((~m[35]&~m[247]&~m[347])|(m[35]&m[247]&~m[347]))&BiasedRNG[62])|(((m[35]&~m[247]&~m[347])|(~m[35]&m[247]&m[347]))&~BiasedRNG[62])|((~m[35]&~m[247]&m[347])|(m[35]&~m[247]&m[347])|(m[35]&m[247]&m[347]));
    m[139] = (((~m[35]&~m[257]&~m[357])|(m[35]&m[257]&~m[357]))&BiasedRNG[63])|(((m[35]&~m[257]&~m[357])|(~m[35]&m[257]&m[357]))&~BiasedRNG[63])|((~m[35]&~m[257]&m[357])|(m[35]&~m[257]&m[357])|(m[35]&m[257]&m[357]));
    m[142] = (((~m[36]&~m[188]&~m[288])|(m[36]&m[188]&~m[288]))&BiasedRNG[64])|(((m[36]&~m[188]&~m[288])|(~m[36]&m[188]&m[288]))&~BiasedRNG[64])|((~m[36]&~m[188]&m[288])|(m[36]&~m[188]&m[288])|(m[36]&m[188]&m[288]));
    m[143] = (((~m[36]&~m[198]&~m[298])|(m[36]&m[198]&~m[298]))&BiasedRNG[65])|(((m[36]&~m[198]&~m[298])|(~m[36]&m[198]&m[298]))&~BiasedRNG[65])|((~m[36]&~m[198]&m[298])|(m[36]&~m[198]&m[298])|(m[36]&m[198]&m[298]));
    m[144] = (((~m[36]&~m[208]&~m[308])|(m[36]&m[208]&~m[308]))&BiasedRNG[66])|(((m[36]&~m[208]&~m[308])|(~m[36]&m[208]&m[308]))&~BiasedRNG[66])|((~m[36]&~m[208]&m[308])|(m[36]&~m[208]&m[308])|(m[36]&m[208]&m[308]));
    m[145] = (((~m[36]&~m[218]&~m[318])|(m[36]&m[218]&~m[318]))&BiasedRNG[67])|(((m[36]&~m[218]&~m[318])|(~m[36]&m[218]&m[318]))&~BiasedRNG[67])|((~m[36]&~m[218]&m[318])|(m[36]&~m[218]&m[318])|(m[36]&m[218]&m[318]));
    m[146] = (((~m[37]&~m[228]&~m[328])|(m[37]&m[228]&~m[328]))&BiasedRNG[68])|(((m[37]&~m[228]&~m[328])|(~m[37]&m[228]&m[328]))&~BiasedRNG[68])|((~m[37]&~m[228]&m[328])|(m[37]&~m[228]&m[328])|(m[37]&m[228]&m[328]));
    m[147] = (((~m[37]&~m[238]&~m[338])|(m[37]&m[238]&~m[338]))&BiasedRNG[69])|(((m[37]&~m[238]&~m[338])|(~m[37]&m[238]&m[338]))&~BiasedRNG[69])|((~m[37]&~m[238]&m[338])|(m[37]&~m[238]&m[338])|(m[37]&m[238]&m[338]));
    m[148] = (((~m[37]&~m[248]&~m[348])|(m[37]&m[248]&~m[348]))&BiasedRNG[70])|(((m[37]&~m[248]&~m[348])|(~m[37]&m[248]&m[348]))&~BiasedRNG[70])|((~m[37]&~m[248]&m[348])|(m[37]&~m[248]&m[348])|(m[37]&m[248]&m[348]));
    m[149] = (((~m[37]&~m[258]&~m[358])|(m[37]&m[258]&~m[358]))&BiasedRNG[71])|(((m[37]&~m[258]&~m[358])|(~m[37]&m[258]&m[358]))&~BiasedRNG[71])|((~m[37]&~m[258]&m[358])|(m[37]&~m[258]&m[358])|(m[37]&m[258]&m[358]));
    m[152] = (((~m[38]&~m[189]&~m[289])|(m[38]&m[189]&~m[289]))&BiasedRNG[72])|(((m[38]&~m[189]&~m[289])|(~m[38]&m[189]&m[289]))&~BiasedRNG[72])|((~m[38]&~m[189]&m[289])|(m[38]&~m[189]&m[289])|(m[38]&m[189]&m[289]));
    m[153] = (((~m[38]&~m[199]&~m[299])|(m[38]&m[199]&~m[299]))&BiasedRNG[73])|(((m[38]&~m[199]&~m[299])|(~m[38]&m[199]&m[299]))&~BiasedRNG[73])|((~m[38]&~m[199]&m[299])|(m[38]&~m[199]&m[299])|(m[38]&m[199]&m[299]));
    m[154] = (((~m[38]&~m[209]&~m[309])|(m[38]&m[209]&~m[309]))&BiasedRNG[74])|(((m[38]&~m[209]&~m[309])|(~m[38]&m[209]&m[309]))&~BiasedRNG[74])|((~m[38]&~m[209]&m[309])|(m[38]&~m[209]&m[309])|(m[38]&m[209]&m[309]));
    m[155] = (((~m[38]&~m[219]&~m[319])|(m[38]&m[219]&~m[319]))&BiasedRNG[75])|(((m[38]&~m[219]&~m[319])|(~m[38]&m[219]&m[319]))&~BiasedRNG[75])|((~m[38]&~m[219]&m[319])|(m[38]&~m[219]&m[319])|(m[38]&m[219]&m[319]));
    m[156] = (((~m[39]&~m[229]&~m[329])|(m[39]&m[229]&~m[329]))&BiasedRNG[76])|(((m[39]&~m[229]&~m[329])|(~m[39]&m[229]&m[329]))&~BiasedRNG[76])|((~m[39]&~m[229]&m[329])|(m[39]&~m[229]&m[329])|(m[39]&m[229]&m[329]));
    m[157] = (((~m[39]&~m[239]&~m[339])|(m[39]&m[239]&~m[339]))&BiasedRNG[77])|(((m[39]&~m[239]&~m[339])|(~m[39]&m[239]&m[339]))&~BiasedRNG[77])|((~m[39]&~m[239]&m[339])|(m[39]&~m[239]&m[339])|(m[39]&m[239]&m[339]));
    m[158] = (((~m[39]&~m[249]&~m[349])|(m[39]&m[249]&~m[349]))&BiasedRNG[78])|(((m[39]&~m[249]&~m[349])|(~m[39]&m[249]&m[349]))&~BiasedRNG[78])|((~m[39]&~m[249]&m[349])|(m[39]&~m[249]&m[349])|(m[39]&m[249]&m[349]));
    m[159] = (((~m[39]&~m[259]&~m[359])|(m[39]&m[259]&~m[359]))&BiasedRNG[79])|(((m[39]&~m[259]&~m[359])|(~m[39]&m[259]&m[359]))&~BiasedRNG[79])|((~m[39]&~m[259]&m[359])|(m[39]&~m[259]&m[359])|(m[39]&m[259]&m[359]));
    m[162] = (((~m[40]&~m[80]&~m[262])|(m[40]&m[80]&~m[262]))&BiasedRNG[80])|(((m[40]&~m[80]&~m[262])|(~m[40]&m[80]&m[262]))&~BiasedRNG[80])|((~m[40]&~m[80]&m[262])|(m[40]&~m[80]&m[262])|(m[40]&m[80]&m[262]));
    m[163] = (((~m[40]&~m[90]&~m[263])|(m[40]&m[90]&~m[263]))&BiasedRNG[81])|(((m[40]&~m[90]&~m[263])|(~m[40]&m[90]&m[263]))&~BiasedRNG[81])|((~m[40]&~m[90]&m[263])|(m[40]&~m[90]&m[263])|(m[40]&m[90]&m[263]));
    m[164] = (((~m[40]&~m[100]&~m[264])|(m[40]&m[100]&~m[264]))&BiasedRNG[82])|(((m[40]&~m[100]&~m[264])|(~m[40]&m[100]&m[264]))&~BiasedRNG[82])|((~m[40]&~m[100]&m[264])|(m[40]&~m[100]&m[264])|(m[40]&m[100]&m[264]));
    m[165] = (((~m[40]&~m[110]&~m[265])|(m[40]&m[110]&~m[265]))&BiasedRNG[83])|(((m[40]&~m[110]&~m[265])|(~m[40]&m[110]&m[265]))&~BiasedRNG[83])|((~m[40]&~m[110]&m[265])|(m[40]&~m[110]&m[265])|(m[40]&m[110]&m[265]));
    m[166] = (((~m[41]&~m[120]&~m[266])|(m[41]&m[120]&~m[266]))&BiasedRNG[84])|(((m[41]&~m[120]&~m[266])|(~m[41]&m[120]&m[266]))&~BiasedRNG[84])|((~m[41]&~m[120]&m[266])|(m[41]&~m[120]&m[266])|(m[41]&m[120]&m[266]));
    m[167] = (((~m[41]&~m[130]&~m[267])|(m[41]&m[130]&~m[267]))&BiasedRNG[85])|(((m[41]&~m[130]&~m[267])|(~m[41]&m[130]&m[267]))&~BiasedRNG[85])|((~m[41]&~m[130]&m[267])|(m[41]&~m[130]&m[267])|(m[41]&m[130]&m[267]));
    m[168] = (((~m[41]&~m[140]&~m[268])|(m[41]&m[140]&~m[268]))&BiasedRNG[86])|(((m[41]&~m[140]&~m[268])|(~m[41]&m[140]&m[268]))&~BiasedRNG[86])|((~m[41]&~m[140]&m[268])|(m[41]&~m[140]&m[268])|(m[41]&m[140]&m[268]));
    m[169] = (((~m[41]&~m[150]&~m[269])|(m[41]&m[150]&~m[269]))&BiasedRNG[87])|(((m[41]&~m[150]&~m[269])|(~m[41]&m[150]&m[269]))&~BiasedRNG[87])|((~m[41]&~m[150]&m[269])|(m[41]&~m[150]&m[269])|(m[41]&m[150]&m[269]));
    m[172] = (((~m[42]&~m[81]&~m[272])|(m[42]&m[81]&~m[272]))&BiasedRNG[88])|(((m[42]&~m[81]&~m[272])|(~m[42]&m[81]&m[272]))&~BiasedRNG[88])|((~m[42]&~m[81]&m[272])|(m[42]&~m[81]&m[272])|(m[42]&m[81]&m[272]));
    m[173] = (((~m[42]&~m[91]&~m[273])|(m[42]&m[91]&~m[273]))&BiasedRNG[89])|(((m[42]&~m[91]&~m[273])|(~m[42]&m[91]&m[273]))&~BiasedRNG[89])|((~m[42]&~m[91]&m[273])|(m[42]&~m[91]&m[273])|(m[42]&m[91]&m[273]));
    m[174] = (((~m[42]&~m[101]&~m[274])|(m[42]&m[101]&~m[274]))&BiasedRNG[90])|(((m[42]&~m[101]&~m[274])|(~m[42]&m[101]&m[274]))&~BiasedRNG[90])|((~m[42]&~m[101]&m[274])|(m[42]&~m[101]&m[274])|(m[42]&m[101]&m[274]));
    m[175] = (((~m[42]&~m[111]&~m[275])|(m[42]&m[111]&~m[275]))&BiasedRNG[91])|(((m[42]&~m[111]&~m[275])|(~m[42]&m[111]&m[275]))&~BiasedRNG[91])|((~m[42]&~m[111]&m[275])|(m[42]&~m[111]&m[275])|(m[42]&m[111]&m[275]));
    m[176] = (((~m[43]&~m[121]&~m[276])|(m[43]&m[121]&~m[276]))&BiasedRNG[92])|(((m[43]&~m[121]&~m[276])|(~m[43]&m[121]&m[276]))&~BiasedRNG[92])|((~m[43]&~m[121]&m[276])|(m[43]&~m[121]&m[276])|(m[43]&m[121]&m[276]));
    m[177] = (((~m[43]&~m[131]&~m[277])|(m[43]&m[131]&~m[277]))&BiasedRNG[93])|(((m[43]&~m[131]&~m[277])|(~m[43]&m[131]&m[277]))&~BiasedRNG[93])|((~m[43]&~m[131]&m[277])|(m[43]&~m[131]&m[277])|(m[43]&m[131]&m[277]));
    m[178] = (((~m[43]&~m[141]&~m[278])|(m[43]&m[141]&~m[278]))&BiasedRNG[94])|(((m[43]&~m[141]&~m[278])|(~m[43]&m[141]&m[278]))&~BiasedRNG[94])|((~m[43]&~m[141]&m[278])|(m[43]&~m[141]&m[278])|(m[43]&m[141]&m[278]));
    m[179] = (((~m[43]&~m[151]&~m[279])|(m[43]&m[151]&~m[279]))&BiasedRNG[95])|(((m[43]&~m[151]&~m[279])|(~m[43]&m[151]&m[279]))&~BiasedRNG[95])|((~m[43]&~m[151]&m[279])|(m[43]&~m[151]&m[279])|(m[43]&m[151]&m[279]));
    m[261] = (((m[70]&~m[161]&m[360])|(~m[70]&m[161]&m[360]))&BiasedRNG[96])|(((m[70]&m[161]&~m[360]))&~BiasedRNG[96])|((m[70]&m[161]&m[360]));
    m[270] = (((m[61]&~m[170]&m[361])|(~m[61]&m[170]&m[361]))&BiasedRNG[97])|(((m[61]&m[170]&~m[361]))&~BiasedRNG[97])|((m[61]&m[170]&m[361]));
    m[271] = (((m[71]&~m[171]&m[366])|(~m[71]&m[171]&m[366]))&BiasedRNG[98])|(((m[71]&m[171]&~m[366]))&~BiasedRNG[98])|((m[71]&m[171]&m[366]));
    m[365] = (((m[262]&~m[366]&~m[367]&~m[368]&~m[369])|(~m[262]&~m[366]&~m[367]&m[368]&~m[369])|(m[262]&m[366]&~m[367]&m[368]&~m[369])|(m[262]&~m[366]&m[367]&m[368]&~m[369])|(~m[262]&m[366]&~m[367]&~m[368]&m[369])|(~m[262]&~m[366]&m[367]&~m[368]&m[369])|(m[262]&m[366]&m[367]&~m[368]&m[369])|(~m[262]&m[366]&m[367]&m[368]&m[369]))&UnbiasedRNG[20])|((m[262]&~m[366]&~m[367]&m[368]&~m[369])|(~m[262]&~m[366]&~m[367]&~m[368]&m[369])|(m[262]&~m[366]&~m[367]&~m[368]&m[369])|(m[262]&m[366]&~m[367]&~m[368]&m[369])|(m[262]&~m[366]&m[367]&~m[368]&m[369])|(~m[262]&~m[366]&~m[367]&m[368]&m[369])|(m[262]&~m[366]&~m[367]&m[368]&m[369])|(~m[262]&m[366]&~m[367]&m[368]&m[369])|(m[262]&m[366]&~m[367]&m[368]&m[369])|(~m[262]&~m[366]&m[367]&m[368]&m[369])|(m[262]&~m[366]&m[367]&m[368]&m[369])|(m[262]&m[366]&m[367]&m[368]&m[369]));
    m[370] = (((m[368]&~m[371]&~m[372]&~m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&m[373]&~m[374])|(m[368]&m[371]&~m[372]&m[373]&~m[374])|(m[368]&~m[371]&m[372]&m[373]&~m[374])|(~m[368]&m[371]&~m[372]&~m[373]&m[374])|(~m[368]&~m[371]&m[372]&~m[373]&m[374])|(m[368]&m[371]&m[372]&~m[373]&m[374])|(~m[368]&m[371]&m[372]&m[373]&m[374]))&UnbiasedRNG[21])|((m[368]&~m[371]&~m[372]&m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&m[372]&~m[373]&m[374])|(~m[368]&~m[371]&~m[372]&m[373]&m[374])|(m[368]&~m[371]&~m[372]&m[373]&m[374])|(~m[368]&m[371]&~m[372]&m[373]&m[374])|(m[368]&m[371]&~m[372]&m[373]&m[374])|(~m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&m[371]&m[372]&m[373]&m[374]));
    m[375] = (((m[263]&~m[376]&~m[377]&~m[378]&~m[379])|(~m[263]&~m[376]&~m[377]&m[378]&~m[379])|(m[263]&m[376]&~m[377]&m[378]&~m[379])|(m[263]&~m[376]&m[377]&m[378]&~m[379])|(~m[263]&m[376]&~m[377]&~m[378]&m[379])|(~m[263]&~m[376]&m[377]&~m[378]&m[379])|(m[263]&m[376]&m[377]&~m[378]&m[379])|(~m[263]&m[376]&m[377]&m[378]&m[379]))&UnbiasedRNG[22])|((m[263]&~m[376]&~m[377]&m[378]&~m[379])|(~m[263]&~m[376]&~m[377]&~m[378]&m[379])|(m[263]&~m[376]&~m[377]&~m[378]&m[379])|(m[263]&m[376]&~m[377]&~m[378]&m[379])|(m[263]&~m[376]&m[377]&~m[378]&m[379])|(~m[263]&~m[376]&~m[377]&m[378]&m[379])|(m[263]&~m[376]&~m[377]&m[378]&m[379])|(~m[263]&m[376]&~m[377]&m[378]&m[379])|(m[263]&m[376]&~m[377]&m[378]&m[379])|(~m[263]&~m[376]&m[377]&m[378]&m[379])|(m[263]&~m[376]&m[377]&m[378]&m[379])|(m[263]&m[376]&m[377]&m[378]&m[379]));
    m[380] = (((m[378]&~m[381]&~m[382]&~m[383]&~m[384])|(~m[378]&~m[381]&~m[382]&m[383]&~m[384])|(m[378]&m[381]&~m[382]&m[383]&~m[384])|(m[378]&~m[381]&m[382]&m[383]&~m[384])|(~m[378]&m[381]&~m[382]&~m[383]&m[384])|(~m[378]&~m[381]&m[382]&~m[383]&m[384])|(m[378]&m[381]&m[382]&~m[383]&m[384])|(~m[378]&m[381]&m[382]&m[383]&m[384]))&UnbiasedRNG[23])|((m[378]&~m[381]&~m[382]&m[383]&~m[384])|(~m[378]&~m[381]&~m[382]&~m[383]&m[384])|(m[378]&~m[381]&~m[382]&~m[383]&m[384])|(m[378]&m[381]&~m[382]&~m[383]&m[384])|(m[378]&~m[381]&m[382]&~m[383]&m[384])|(~m[378]&~m[381]&~m[382]&m[383]&m[384])|(m[378]&~m[381]&~m[382]&m[383]&m[384])|(~m[378]&m[381]&~m[382]&m[383]&m[384])|(m[378]&m[381]&~m[382]&m[383]&m[384])|(~m[378]&~m[381]&m[382]&m[383]&m[384])|(m[378]&~m[381]&m[382]&m[383]&m[384])|(m[378]&m[381]&m[382]&m[383]&m[384]));
    m[385] = (((m[383]&~m[386]&~m[387]&~m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&m[388]&~m[389])|(m[383]&m[386]&~m[387]&m[388]&~m[389])|(m[383]&~m[386]&m[387]&m[388]&~m[389])|(~m[383]&m[386]&~m[387]&~m[388]&m[389])|(~m[383]&~m[386]&m[387]&~m[388]&m[389])|(m[383]&m[386]&m[387]&~m[388]&m[389])|(~m[383]&m[386]&m[387]&m[388]&m[389]))&UnbiasedRNG[24])|((m[383]&~m[386]&~m[387]&m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&m[387]&~m[388]&m[389])|(~m[383]&~m[386]&~m[387]&m[388]&m[389])|(m[383]&~m[386]&~m[387]&m[388]&m[389])|(~m[383]&m[386]&~m[387]&m[388]&m[389])|(m[383]&m[386]&~m[387]&m[388]&m[389])|(~m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&m[386]&m[387]&m[388]&m[389]));
    m[390] = (((m[264]&~m[391]&~m[392]&~m[393]&~m[394])|(~m[264]&~m[391]&~m[392]&m[393]&~m[394])|(m[264]&m[391]&~m[392]&m[393]&~m[394])|(m[264]&~m[391]&m[392]&m[393]&~m[394])|(~m[264]&m[391]&~m[392]&~m[393]&m[394])|(~m[264]&~m[391]&m[392]&~m[393]&m[394])|(m[264]&m[391]&m[392]&~m[393]&m[394])|(~m[264]&m[391]&m[392]&m[393]&m[394]))&UnbiasedRNG[25])|((m[264]&~m[391]&~m[392]&m[393]&~m[394])|(~m[264]&~m[391]&~m[392]&~m[393]&m[394])|(m[264]&~m[391]&~m[392]&~m[393]&m[394])|(m[264]&m[391]&~m[392]&~m[393]&m[394])|(m[264]&~m[391]&m[392]&~m[393]&m[394])|(~m[264]&~m[391]&~m[392]&m[393]&m[394])|(m[264]&~m[391]&~m[392]&m[393]&m[394])|(~m[264]&m[391]&~m[392]&m[393]&m[394])|(m[264]&m[391]&~m[392]&m[393]&m[394])|(~m[264]&~m[391]&m[392]&m[393]&m[394])|(m[264]&~m[391]&m[392]&m[393]&m[394])|(m[264]&m[391]&m[392]&m[393]&m[394]));
    m[395] = (((m[393]&~m[396]&~m[397]&~m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&m[398]&~m[399])|(m[393]&m[396]&~m[397]&m[398]&~m[399])|(m[393]&~m[396]&m[397]&m[398]&~m[399])|(~m[393]&m[396]&~m[397]&~m[398]&m[399])|(~m[393]&~m[396]&m[397]&~m[398]&m[399])|(m[393]&m[396]&m[397]&~m[398]&m[399])|(~m[393]&m[396]&m[397]&m[398]&m[399]))&UnbiasedRNG[26])|((m[393]&~m[396]&~m[397]&m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&m[397]&~m[398]&m[399])|(~m[393]&~m[396]&~m[397]&m[398]&m[399])|(m[393]&~m[396]&~m[397]&m[398]&m[399])|(~m[393]&m[396]&~m[397]&m[398]&m[399])|(m[393]&m[396]&~m[397]&m[398]&m[399])|(~m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&m[396]&m[397]&m[398]&m[399]));
    m[400] = (((m[398]&~m[401]&~m[402]&~m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&m[403]&~m[404])|(m[398]&m[401]&~m[402]&m[403]&~m[404])|(m[398]&~m[401]&m[402]&m[403]&~m[404])|(~m[398]&m[401]&~m[402]&~m[403]&m[404])|(~m[398]&~m[401]&m[402]&~m[403]&m[404])|(m[398]&m[401]&m[402]&~m[403]&m[404])|(~m[398]&m[401]&m[402]&m[403]&m[404]))&UnbiasedRNG[27])|((m[398]&~m[401]&~m[402]&m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&m[402]&~m[403]&m[404])|(~m[398]&~m[401]&~m[402]&m[403]&m[404])|(m[398]&~m[401]&~m[402]&m[403]&m[404])|(~m[398]&m[401]&~m[402]&m[403]&m[404])|(m[398]&m[401]&~m[402]&m[403]&m[404])|(~m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&m[401]&m[402]&m[403]&m[404]));
    m[405] = (((m[403]&~m[406]&~m[407]&~m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&m[408]&~m[409])|(m[403]&m[406]&~m[407]&m[408]&~m[409])|(m[403]&~m[406]&m[407]&m[408]&~m[409])|(~m[403]&m[406]&~m[407]&~m[408]&m[409])|(~m[403]&~m[406]&m[407]&~m[408]&m[409])|(m[403]&m[406]&m[407]&~m[408]&m[409])|(~m[403]&m[406]&m[407]&m[408]&m[409]))&UnbiasedRNG[28])|((m[403]&~m[406]&~m[407]&m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&m[407]&~m[408]&m[409])|(~m[403]&~m[406]&~m[407]&m[408]&m[409])|(m[403]&~m[406]&~m[407]&m[408]&m[409])|(~m[403]&m[406]&~m[407]&m[408]&m[409])|(m[403]&m[406]&~m[407]&m[408]&m[409])|(~m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&m[406]&m[407]&m[408]&m[409]));
    m[410] = (((m[265]&~m[411]&~m[412]&~m[413]&~m[414])|(~m[265]&~m[411]&~m[412]&m[413]&~m[414])|(m[265]&m[411]&~m[412]&m[413]&~m[414])|(m[265]&~m[411]&m[412]&m[413]&~m[414])|(~m[265]&m[411]&~m[412]&~m[413]&m[414])|(~m[265]&~m[411]&m[412]&~m[413]&m[414])|(m[265]&m[411]&m[412]&~m[413]&m[414])|(~m[265]&m[411]&m[412]&m[413]&m[414]))&UnbiasedRNG[29])|((m[265]&~m[411]&~m[412]&m[413]&~m[414])|(~m[265]&~m[411]&~m[412]&~m[413]&m[414])|(m[265]&~m[411]&~m[412]&~m[413]&m[414])|(m[265]&m[411]&~m[412]&~m[413]&m[414])|(m[265]&~m[411]&m[412]&~m[413]&m[414])|(~m[265]&~m[411]&~m[412]&m[413]&m[414])|(m[265]&~m[411]&~m[412]&m[413]&m[414])|(~m[265]&m[411]&~m[412]&m[413]&m[414])|(m[265]&m[411]&~m[412]&m[413]&m[414])|(~m[265]&~m[411]&m[412]&m[413]&m[414])|(m[265]&~m[411]&m[412]&m[413]&m[414])|(m[265]&m[411]&m[412]&m[413]&m[414]));
    m[415] = (((m[413]&~m[416]&~m[417]&~m[418]&~m[419])|(~m[413]&~m[416]&~m[417]&m[418]&~m[419])|(m[413]&m[416]&~m[417]&m[418]&~m[419])|(m[413]&~m[416]&m[417]&m[418]&~m[419])|(~m[413]&m[416]&~m[417]&~m[418]&m[419])|(~m[413]&~m[416]&m[417]&~m[418]&m[419])|(m[413]&m[416]&m[417]&~m[418]&m[419])|(~m[413]&m[416]&m[417]&m[418]&m[419]))&UnbiasedRNG[30])|((m[413]&~m[416]&~m[417]&m[418]&~m[419])|(~m[413]&~m[416]&~m[417]&~m[418]&m[419])|(m[413]&~m[416]&~m[417]&~m[418]&m[419])|(m[413]&m[416]&~m[417]&~m[418]&m[419])|(m[413]&~m[416]&m[417]&~m[418]&m[419])|(~m[413]&~m[416]&~m[417]&m[418]&m[419])|(m[413]&~m[416]&~m[417]&m[418]&m[419])|(~m[413]&m[416]&~m[417]&m[418]&m[419])|(m[413]&m[416]&~m[417]&m[418]&m[419])|(~m[413]&~m[416]&m[417]&m[418]&m[419])|(m[413]&~m[416]&m[417]&m[418]&m[419])|(m[413]&m[416]&m[417]&m[418]&m[419]));
    m[420] = (((m[418]&~m[421]&~m[422]&~m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&m[423]&~m[424])|(m[418]&m[421]&~m[422]&m[423]&~m[424])|(m[418]&~m[421]&m[422]&m[423]&~m[424])|(~m[418]&m[421]&~m[422]&~m[423]&m[424])|(~m[418]&~m[421]&m[422]&~m[423]&m[424])|(m[418]&m[421]&m[422]&~m[423]&m[424])|(~m[418]&m[421]&m[422]&m[423]&m[424]))&UnbiasedRNG[31])|((m[418]&~m[421]&~m[422]&m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&m[422]&~m[423]&m[424])|(~m[418]&~m[421]&~m[422]&m[423]&m[424])|(m[418]&~m[421]&~m[422]&m[423]&m[424])|(~m[418]&m[421]&~m[422]&m[423]&m[424])|(m[418]&m[421]&~m[422]&m[423]&m[424])|(~m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&m[421]&m[422]&m[423]&m[424]));
    m[425] = (((m[423]&~m[426]&~m[427]&~m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&m[428]&~m[429])|(m[423]&m[426]&~m[427]&m[428]&~m[429])|(m[423]&~m[426]&m[427]&m[428]&~m[429])|(~m[423]&m[426]&~m[427]&~m[428]&m[429])|(~m[423]&~m[426]&m[427]&~m[428]&m[429])|(m[423]&m[426]&m[427]&~m[428]&m[429])|(~m[423]&m[426]&m[427]&m[428]&m[429]))&UnbiasedRNG[32])|((m[423]&~m[426]&~m[427]&m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&m[427]&~m[428]&m[429])|(~m[423]&~m[426]&~m[427]&m[428]&m[429])|(m[423]&~m[426]&~m[427]&m[428]&m[429])|(~m[423]&m[426]&~m[427]&m[428]&m[429])|(m[423]&m[426]&~m[427]&m[428]&m[429])|(~m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&m[426]&m[427]&m[428]&m[429]));
    m[430] = (((m[428]&~m[431]&~m[432]&~m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&m[433]&~m[434])|(m[428]&m[431]&~m[432]&m[433]&~m[434])|(m[428]&~m[431]&m[432]&m[433]&~m[434])|(~m[428]&m[431]&~m[432]&~m[433]&m[434])|(~m[428]&~m[431]&m[432]&~m[433]&m[434])|(m[428]&m[431]&m[432]&~m[433]&m[434])|(~m[428]&m[431]&m[432]&m[433]&m[434]))&UnbiasedRNG[33])|((m[428]&~m[431]&~m[432]&m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&m[432]&~m[433]&m[434])|(~m[428]&~m[431]&~m[432]&m[433]&m[434])|(m[428]&~m[431]&~m[432]&m[433]&m[434])|(~m[428]&m[431]&~m[432]&m[433]&m[434])|(m[428]&m[431]&~m[432]&m[433]&m[434])|(~m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&m[431]&m[432]&m[433]&m[434]));
    m[435] = (((m[266]&~m[436]&~m[437]&~m[438]&~m[439])|(~m[266]&~m[436]&~m[437]&m[438]&~m[439])|(m[266]&m[436]&~m[437]&m[438]&~m[439])|(m[266]&~m[436]&m[437]&m[438]&~m[439])|(~m[266]&m[436]&~m[437]&~m[438]&m[439])|(~m[266]&~m[436]&m[437]&~m[438]&m[439])|(m[266]&m[436]&m[437]&~m[438]&m[439])|(~m[266]&m[436]&m[437]&m[438]&m[439]))&UnbiasedRNG[34])|((m[266]&~m[436]&~m[437]&m[438]&~m[439])|(~m[266]&~m[436]&~m[437]&~m[438]&m[439])|(m[266]&~m[436]&~m[437]&~m[438]&m[439])|(m[266]&m[436]&~m[437]&~m[438]&m[439])|(m[266]&~m[436]&m[437]&~m[438]&m[439])|(~m[266]&~m[436]&~m[437]&m[438]&m[439])|(m[266]&~m[436]&~m[437]&m[438]&m[439])|(~m[266]&m[436]&~m[437]&m[438]&m[439])|(m[266]&m[436]&~m[437]&m[438]&m[439])|(~m[266]&~m[436]&m[437]&m[438]&m[439])|(m[266]&~m[436]&m[437]&m[438]&m[439])|(m[266]&m[436]&m[437]&m[438]&m[439]));
    m[440] = (((m[438]&~m[441]&~m[442]&~m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&m[443]&~m[444])|(m[438]&m[441]&~m[442]&m[443]&~m[444])|(m[438]&~m[441]&m[442]&m[443]&~m[444])|(~m[438]&m[441]&~m[442]&~m[443]&m[444])|(~m[438]&~m[441]&m[442]&~m[443]&m[444])|(m[438]&m[441]&m[442]&~m[443]&m[444])|(~m[438]&m[441]&m[442]&m[443]&m[444]))&UnbiasedRNG[35])|((m[438]&~m[441]&~m[442]&m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&m[442]&~m[443]&m[444])|(~m[438]&~m[441]&~m[442]&m[443]&m[444])|(m[438]&~m[441]&~m[442]&m[443]&m[444])|(~m[438]&m[441]&~m[442]&m[443]&m[444])|(m[438]&m[441]&~m[442]&m[443]&m[444])|(~m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&m[441]&m[442]&m[443]&m[444]));
    m[445] = (((m[443]&~m[446]&~m[447]&~m[448]&~m[449])|(~m[443]&~m[446]&~m[447]&m[448]&~m[449])|(m[443]&m[446]&~m[447]&m[448]&~m[449])|(m[443]&~m[446]&m[447]&m[448]&~m[449])|(~m[443]&m[446]&~m[447]&~m[448]&m[449])|(~m[443]&~m[446]&m[447]&~m[448]&m[449])|(m[443]&m[446]&m[447]&~m[448]&m[449])|(~m[443]&m[446]&m[447]&m[448]&m[449]))&UnbiasedRNG[36])|((m[443]&~m[446]&~m[447]&m[448]&~m[449])|(~m[443]&~m[446]&~m[447]&~m[448]&m[449])|(m[443]&~m[446]&~m[447]&~m[448]&m[449])|(m[443]&m[446]&~m[447]&~m[448]&m[449])|(m[443]&~m[446]&m[447]&~m[448]&m[449])|(~m[443]&~m[446]&~m[447]&m[448]&m[449])|(m[443]&~m[446]&~m[447]&m[448]&m[449])|(~m[443]&m[446]&~m[447]&m[448]&m[449])|(m[443]&m[446]&~m[447]&m[448]&m[449])|(~m[443]&~m[446]&m[447]&m[448]&m[449])|(m[443]&~m[446]&m[447]&m[448]&m[449])|(m[443]&m[446]&m[447]&m[448]&m[449]));
    m[450] = (((m[448]&~m[451]&~m[452]&~m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&m[453]&~m[454])|(m[448]&m[451]&~m[452]&m[453]&~m[454])|(m[448]&~m[451]&m[452]&m[453]&~m[454])|(~m[448]&m[451]&~m[452]&~m[453]&m[454])|(~m[448]&~m[451]&m[452]&~m[453]&m[454])|(m[448]&m[451]&m[452]&~m[453]&m[454])|(~m[448]&m[451]&m[452]&m[453]&m[454]))&UnbiasedRNG[37])|((m[448]&~m[451]&~m[452]&m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&m[452]&~m[453]&m[454])|(~m[448]&~m[451]&~m[452]&m[453]&m[454])|(m[448]&~m[451]&~m[452]&m[453]&m[454])|(~m[448]&m[451]&~m[452]&m[453]&m[454])|(m[448]&m[451]&~m[452]&m[453]&m[454])|(~m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&m[451]&m[452]&m[453]&m[454]));
    m[455] = (((m[453]&~m[456]&~m[457]&~m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&m[458]&~m[459])|(m[453]&m[456]&~m[457]&m[458]&~m[459])|(m[453]&~m[456]&m[457]&m[458]&~m[459])|(~m[453]&m[456]&~m[457]&~m[458]&m[459])|(~m[453]&~m[456]&m[457]&~m[458]&m[459])|(m[453]&m[456]&m[457]&~m[458]&m[459])|(~m[453]&m[456]&m[457]&m[458]&m[459]))&UnbiasedRNG[38])|((m[453]&~m[456]&~m[457]&m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&m[457]&~m[458]&m[459])|(~m[453]&~m[456]&~m[457]&m[458]&m[459])|(m[453]&~m[456]&~m[457]&m[458]&m[459])|(~m[453]&m[456]&~m[457]&m[458]&m[459])|(m[453]&m[456]&~m[457]&m[458]&m[459])|(~m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&m[456]&m[457]&m[458]&m[459]));
    m[460] = (((m[458]&~m[461]&~m[462]&~m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&m[463]&~m[464])|(m[458]&m[461]&~m[462]&m[463]&~m[464])|(m[458]&~m[461]&m[462]&m[463]&~m[464])|(~m[458]&m[461]&~m[462]&~m[463]&m[464])|(~m[458]&~m[461]&m[462]&~m[463]&m[464])|(m[458]&m[461]&m[462]&~m[463]&m[464])|(~m[458]&m[461]&m[462]&m[463]&m[464]))&UnbiasedRNG[39])|((m[458]&~m[461]&~m[462]&m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&m[462]&~m[463]&m[464])|(~m[458]&~m[461]&~m[462]&m[463]&m[464])|(m[458]&~m[461]&~m[462]&m[463]&m[464])|(~m[458]&m[461]&~m[462]&m[463]&m[464])|(m[458]&m[461]&~m[462]&m[463]&m[464])|(~m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&m[461]&m[462]&m[463]&m[464]));
    m[465] = (((m[267]&~m[466]&~m[467]&~m[468]&~m[469])|(~m[267]&~m[466]&~m[467]&m[468]&~m[469])|(m[267]&m[466]&~m[467]&m[468]&~m[469])|(m[267]&~m[466]&m[467]&m[468]&~m[469])|(~m[267]&m[466]&~m[467]&~m[468]&m[469])|(~m[267]&~m[466]&m[467]&~m[468]&m[469])|(m[267]&m[466]&m[467]&~m[468]&m[469])|(~m[267]&m[466]&m[467]&m[468]&m[469]))&UnbiasedRNG[40])|((m[267]&~m[466]&~m[467]&m[468]&~m[469])|(~m[267]&~m[466]&~m[467]&~m[468]&m[469])|(m[267]&~m[466]&~m[467]&~m[468]&m[469])|(m[267]&m[466]&~m[467]&~m[468]&m[469])|(m[267]&~m[466]&m[467]&~m[468]&m[469])|(~m[267]&~m[466]&~m[467]&m[468]&m[469])|(m[267]&~m[466]&~m[467]&m[468]&m[469])|(~m[267]&m[466]&~m[467]&m[468]&m[469])|(m[267]&m[466]&~m[467]&m[468]&m[469])|(~m[267]&~m[466]&m[467]&m[468]&m[469])|(m[267]&~m[466]&m[467]&m[468]&m[469])|(m[267]&m[466]&m[467]&m[468]&m[469]));
    m[470] = (((m[468]&~m[471]&~m[472]&~m[473]&~m[474])|(~m[468]&~m[471]&~m[472]&m[473]&~m[474])|(m[468]&m[471]&~m[472]&m[473]&~m[474])|(m[468]&~m[471]&m[472]&m[473]&~m[474])|(~m[468]&m[471]&~m[472]&~m[473]&m[474])|(~m[468]&~m[471]&m[472]&~m[473]&m[474])|(m[468]&m[471]&m[472]&~m[473]&m[474])|(~m[468]&m[471]&m[472]&m[473]&m[474]))&UnbiasedRNG[41])|((m[468]&~m[471]&~m[472]&m[473]&~m[474])|(~m[468]&~m[471]&~m[472]&~m[473]&m[474])|(m[468]&~m[471]&~m[472]&~m[473]&m[474])|(m[468]&m[471]&~m[472]&~m[473]&m[474])|(m[468]&~m[471]&m[472]&~m[473]&m[474])|(~m[468]&~m[471]&~m[472]&m[473]&m[474])|(m[468]&~m[471]&~m[472]&m[473]&m[474])|(~m[468]&m[471]&~m[472]&m[473]&m[474])|(m[468]&m[471]&~m[472]&m[473]&m[474])|(~m[468]&~m[471]&m[472]&m[473]&m[474])|(m[468]&~m[471]&m[472]&m[473]&m[474])|(m[468]&m[471]&m[472]&m[473]&m[474]));
    m[475] = (((m[473]&~m[476]&~m[477]&~m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&m[478]&~m[479])|(m[473]&m[476]&~m[477]&m[478]&~m[479])|(m[473]&~m[476]&m[477]&m[478]&~m[479])|(~m[473]&m[476]&~m[477]&~m[478]&m[479])|(~m[473]&~m[476]&m[477]&~m[478]&m[479])|(m[473]&m[476]&m[477]&~m[478]&m[479])|(~m[473]&m[476]&m[477]&m[478]&m[479]))&UnbiasedRNG[42])|((m[473]&~m[476]&~m[477]&m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&m[477]&~m[478]&m[479])|(~m[473]&~m[476]&~m[477]&m[478]&m[479])|(m[473]&~m[476]&~m[477]&m[478]&m[479])|(~m[473]&m[476]&~m[477]&m[478]&m[479])|(m[473]&m[476]&~m[477]&m[478]&m[479])|(~m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&m[476]&m[477]&m[478]&m[479]));
    m[480] = (((m[478]&~m[481]&~m[482]&~m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&m[483]&~m[484])|(m[478]&m[481]&~m[482]&m[483]&~m[484])|(m[478]&~m[481]&m[482]&m[483]&~m[484])|(~m[478]&m[481]&~m[482]&~m[483]&m[484])|(~m[478]&~m[481]&m[482]&~m[483]&m[484])|(m[478]&m[481]&m[482]&~m[483]&m[484])|(~m[478]&m[481]&m[482]&m[483]&m[484]))&UnbiasedRNG[43])|((m[478]&~m[481]&~m[482]&m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&m[482]&~m[483]&m[484])|(~m[478]&~m[481]&~m[482]&m[483]&m[484])|(m[478]&~m[481]&~m[482]&m[483]&m[484])|(~m[478]&m[481]&~m[482]&m[483]&m[484])|(m[478]&m[481]&~m[482]&m[483]&m[484])|(~m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&m[481]&m[482]&m[483]&m[484]));
    m[485] = (((m[483]&~m[486]&~m[487]&~m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&m[488]&~m[489])|(m[483]&m[486]&~m[487]&m[488]&~m[489])|(m[483]&~m[486]&m[487]&m[488]&~m[489])|(~m[483]&m[486]&~m[487]&~m[488]&m[489])|(~m[483]&~m[486]&m[487]&~m[488]&m[489])|(m[483]&m[486]&m[487]&~m[488]&m[489])|(~m[483]&m[486]&m[487]&m[488]&m[489]))&UnbiasedRNG[44])|((m[483]&~m[486]&~m[487]&m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&m[487]&~m[488]&m[489])|(~m[483]&~m[486]&~m[487]&m[488]&m[489])|(m[483]&~m[486]&~m[487]&m[488]&m[489])|(~m[483]&m[486]&~m[487]&m[488]&m[489])|(m[483]&m[486]&~m[487]&m[488]&m[489])|(~m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&m[486]&m[487]&m[488]&m[489]));
    m[490] = (((m[488]&~m[491]&~m[492]&~m[493]&~m[494])|(~m[488]&~m[491]&~m[492]&m[493]&~m[494])|(m[488]&m[491]&~m[492]&m[493]&~m[494])|(m[488]&~m[491]&m[492]&m[493]&~m[494])|(~m[488]&m[491]&~m[492]&~m[493]&m[494])|(~m[488]&~m[491]&m[492]&~m[493]&m[494])|(m[488]&m[491]&m[492]&~m[493]&m[494])|(~m[488]&m[491]&m[492]&m[493]&m[494]))&UnbiasedRNG[45])|((m[488]&~m[491]&~m[492]&m[493]&~m[494])|(~m[488]&~m[491]&~m[492]&~m[493]&m[494])|(m[488]&~m[491]&~m[492]&~m[493]&m[494])|(m[488]&m[491]&~m[492]&~m[493]&m[494])|(m[488]&~m[491]&m[492]&~m[493]&m[494])|(~m[488]&~m[491]&~m[492]&m[493]&m[494])|(m[488]&~m[491]&~m[492]&m[493]&m[494])|(~m[488]&m[491]&~m[492]&m[493]&m[494])|(m[488]&m[491]&~m[492]&m[493]&m[494])|(~m[488]&~m[491]&m[492]&m[493]&m[494])|(m[488]&~m[491]&m[492]&m[493]&m[494])|(m[488]&m[491]&m[492]&m[493]&m[494]));
    m[495] = (((m[493]&~m[496]&~m[497]&~m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&m[498]&~m[499])|(m[493]&m[496]&~m[497]&m[498]&~m[499])|(m[493]&~m[496]&m[497]&m[498]&~m[499])|(~m[493]&m[496]&~m[497]&~m[498]&m[499])|(~m[493]&~m[496]&m[497]&~m[498]&m[499])|(m[493]&m[496]&m[497]&~m[498]&m[499])|(~m[493]&m[496]&m[497]&m[498]&m[499]))&UnbiasedRNG[46])|((m[493]&~m[496]&~m[497]&m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&m[497]&~m[498]&m[499])|(~m[493]&~m[496]&~m[497]&m[498]&m[499])|(m[493]&~m[496]&~m[497]&m[498]&m[499])|(~m[493]&m[496]&~m[497]&m[498]&m[499])|(m[493]&m[496]&~m[497]&m[498]&m[499])|(~m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&m[496]&m[497]&m[498]&m[499]));
    m[500] = (((m[268]&~m[501]&~m[502]&~m[503]&~m[504])|(~m[268]&~m[501]&~m[502]&m[503]&~m[504])|(m[268]&m[501]&~m[502]&m[503]&~m[504])|(m[268]&~m[501]&m[502]&m[503]&~m[504])|(~m[268]&m[501]&~m[502]&~m[503]&m[504])|(~m[268]&~m[501]&m[502]&~m[503]&m[504])|(m[268]&m[501]&m[502]&~m[503]&m[504])|(~m[268]&m[501]&m[502]&m[503]&m[504]))&UnbiasedRNG[47])|((m[268]&~m[501]&~m[502]&m[503]&~m[504])|(~m[268]&~m[501]&~m[502]&~m[503]&m[504])|(m[268]&~m[501]&~m[502]&~m[503]&m[504])|(m[268]&m[501]&~m[502]&~m[503]&m[504])|(m[268]&~m[501]&m[502]&~m[503]&m[504])|(~m[268]&~m[501]&~m[502]&m[503]&m[504])|(m[268]&~m[501]&~m[502]&m[503]&m[504])|(~m[268]&m[501]&~m[502]&m[503]&m[504])|(m[268]&m[501]&~m[502]&m[503]&m[504])|(~m[268]&~m[501]&m[502]&m[503]&m[504])|(m[268]&~m[501]&m[502]&m[503]&m[504])|(m[268]&m[501]&m[502]&m[503]&m[504]));
    m[505] = (((m[503]&~m[506]&~m[507]&~m[508]&~m[509])|(~m[503]&~m[506]&~m[507]&m[508]&~m[509])|(m[503]&m[506]&~m[507]&m[508]&~m[509])|(m[503]&~m[506]&m[507]&m[508]&~m[509])|(~m[503]&m[506]&~m[507]&~m[508]&m[509])|(~m[503]&~m[506]&m[507]&~m[508]&m[509])|(m[503]&m[506]&m[507]&~m[508]&m[509])|(~m[503]&m[506]&m[507]&m[508]&m[509]))&UnbiasedRNG[48])|((m[503]&~m[506]&~m[507]&m[508]&~m[509])|(~m[503]&~m[506]&~m[507]&~m[508]&m[509])|(m[503]&~m[506]&~m[507]&~m[508]&m[509])|(m[503]&m[506]&~m[507]&~m[508]&m[509])|(m[503]&~m[506]&m[507]&~m[508]&m[509])|(~m[503]&~m[506]&~m[507]&m[508]&m[509])|(m[503]&~m[506]&~m[507]&m[508]&m[509])|(~m[503]&m[506]&~m[507]&m[508]&m[509])|(m[503]&m[506]&~m[507]&m[508]&m[509])|(~m[503]&~m[506]&m[507]&m[508]&m[509])|(m[503]&~m[506]&m[507]&m[508]&m[509])|(m[503]&m[506]&m[507]&m[508]&m[509]));
    m[510] = (((m[508]&~m[511]&~m[512]&~m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&m[513]&~m[514])|(m[508]&m[511]&~m[512]&m[513]&~m[514])|(m[508]&~m[511]&m[512]&m[513]&~m[514])|(~m[508]&m[511]&~m[512]&~m[513]&m[514])|(~m[508]&~m[511]&m[512]&~m[513]&m[514])|(m[508]&m[511]&m[512]&~m[513]&m[514])|(~m[508]&m[511]&m[512]&m[513]&m[514]))&UnbiasedRNG[49])|((m[508]&~m[511]&~m[512]&m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&m[512]&~m[513]&m[514])|(~m[508]&~m[511]&~m[512]&m[513]&m[514])|(m[508]&~m[511]&~m[512]&m[513]&m[514])|(~m[508]&m[511]&~m[512]&m[513]&m[514])|(m[508]&m[511]&~m[512]&m[513]&m[514])|(~m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&m[511]&m[512]&m[513]&m[514]));
    m[515] = (((m[513]&~m[516]&~m[517]&~m[518]&~m[519])|(~m[513]&~m[516]&~m[517]&m[518]&~m[519])|(m[513]&m[516]&~m[517]&m[518]&~m[519])|(m[513]&~m[516]&m[517]&m[518]&~m[519])|(~m[513]&m[516]&~m[517]&~m[518]&m[519])|(~m[513]&~m[516]&m[517]&~m[518]&m[519])|(m[513]&m[516]&m[517]&~m[518]&m[519])|(~m[513]&m[516]&m[517]&m[518]&m[519]))&UnbiasedRNG[50])|((m[513]&~m[516]&~m[517]&m[518]&~m[519])|(~m[513]&~m[516]&~m[517]&~m[518]&m[519])|(m[513]&~m[516]&~m[517]&~m[518]&m[519])|(m[513]&m[516]&~m[517]&~m[518]&m[519])|(m[513]&~m[516]&m[517]&~m[518]&m[519])|(~m[513]&~m[516]&~m[517]&m[518]&m[519])|(m[513]&~m[516]&~m[517]&m[518]&m[519])|(~m[513]&m[516]&~m[517]&m[518]&m[519])|(m[513]&m[516]&~m[517]&m[518]&m[519])|(~m[513]&~m[516]&m[517]&m[518]&m[519])|(m[513]&~m[516]&m[517]&m[518]&m[519])|(m[513]&m[516]&m[517]&m[518]&m[519]));
    m[520] = (((m[518]&~m[521]&~m[522]&~m[523]&~m[524])|(~m[518]&~m[521]&~m[522]&m[523]&~m[524])|(m[518]&m[521]&~m[522]&m[523]&~m[524])|(m[518]&~m[521]&m[522]&m[523]&~m[524])|(~m[518]&m[521]&~m[522]&~m[523]&m[524])|(~m[518]&~m[521]&m[522]&~m[523]&m[524])|(m[518]&m[521]&m[522]&~m[523]&m[524])|(~m[518]&m[521]&m[522]&m[523]&m[524]))&UnbiasedRNG[51])|((m[518]&~m[521]&~m[522]&m[523]&~m[524])|(~m[518]&~m[521]&~m[522]&~m[523]&m[524])|(m[518]&~m[521]&~m[522]&~m[523]&m[524])|(m[518]&m[521]&~m[522]&~m[523]&m[524])|(m[518]&~m[521]&m[522]&~m[523]&m[524])|(~m[518]&~m[521]&~m[522]&m[523]&m[524])|(m[518]&~m[521]&~m[522]&m[523]&m[524])|(~m[518]&m[521]&~m[522]&m[523]&m[524])|(m[518]&m[521]&~m[522]&m[523]&m[524])|(~m[518]&~m[521]&m[522]&m[523]&m[524])|(m[518]&~m[521]&m[522]&m[523]&m[524])|(m[518]&m[521]&m[522]&m[523]&m[524]));
    m[525] = (((m[523]&~m[526]&~m[527]&~m[528]&~m[529])|(~m[523]&~m[526]&~m[527]&m[528]&~m[529])|(m[523]&m[526]&~m[527]&m[528]&~m[529])|(m[523]&~m[526]&m[527]&m[528]&~m[529])|(~m[523]&m[526]&~m[527]&~m[528]&m[529])|(~m[523]&~m[526]&m[527]&~m[528]&m[529])|(m[523]&m[526]&m[527]&~m[528]&m[529])|(~m[523]&m[526]&m[527]&m[528]&m[529]))&UnbiasedRNG[52])|((m[523]&~m[526]&~m[527]&m[528]&~m[529])|(~m[523]&~m[526]&~m[527]&~m[528]&m[529])|(m[523]&~m[526]&~m[527]&~m[528]&m[529])|(m[523]&m[526]&~m[527]&~m[528]&m[529])|(m[523]&~m[526]&m[527]&~m[528]&m[529])|(~m[523]&~m[526]&~m[527]&m[528]&m[529])|(m[523]&~m[526]&~m[527]&m[528]&m[529])|(~m[523]&m[526]&~m[527]&m[528]&m[529])|(m[523]&m[526]&~m[527]&m[528]&m[529])|(~m[523]&~m[526]&m[527]&m[528]&m[529])|(m[523]&~m[526]&m[527]&m[528]&m[529])|(m[523]&m[526]&m[527]&m[528]&m[529]));
    m[530] = (((m[528]&~m[531]&~m[532]&~m[533]&~m[534])|(~m[528]&~m[531]&~m[532]&m[533]&~m[534])|(m[528]&m[531]&~m[532]&m[533]&~m[534])|(m[528]&~m[531]&m[532]&m[533]&~m[534])|(~m[528]&m[531]&~m[532]&~m[533]&m[534])|(~m[528]&~m[531]&m[532]&~m[533]&m[534])|(m[528]&m[531]&m[532]&~m[533]&m[534])|(~m[528]&m[531]&m[532]&m[533]&m[534]))&UnbiasedRNG[53])|((m[528]&~m[531]&~m[532]&m[533]&~m[534])|(~m[528]&~m[531]&~m[532]&~m[533]&m[534])|(m[528]&~m[531]&~m[532]&~m[533]&m[534])|(m[528]&m[531]&~m[532]&~m[533]&m[534])|(m[528]&~m[531]&m[532]&~m[533]&m[534])|(~m[528]&~m[531]&~m[532]&m[533]&m[534])|(m[528]&~m[531]&~m[532]&m[533]&m[534])|(~m[528]&m[531]&~m[532]&m[533]&m[534])|(m[528]&m[531]&~m[532]&m[533]&m[534])|(~m[528]&~m[531]&m[532]&m[533]&m[534])|(m[528]&~m[531]&m[532]&m[533]&m[534])|(m[528]&m[531]&m[532]&m[533]&m[534]));
    m[535] = (((m[533]&~m[536]&~m[537]&~m[538]&~m[539])|(~m[533]&~m[536]&~m[537]&m[538]&~m[539])|(m[533]&m[536]&~m[537]&m[538]&~m[539])|(m[533]&~m[536]&m[537]&m[538]&~m[539])|(~m[533]&m[536]&~m[537]&~m[538]&m[539])|(~m[533]&~m[536]&m[537]&~m[538]&m[539])|(m[533]&m[536]&m[537]&~m[538]&m[539])|(~m[533]&m[536]&m[537]&m[538]&m[539]))&UnbiasedRNG[54])|((m[533]&~m[536]&~m[537]&m[538]&~m[539])|(~m[533]&~m[536]&~m[537]&~m[538]&m[539])|(m[533]&~m[536]&~m[537]&~m[538]&m[539])|(m[533]&m[536]&~m[537]&~m[538]&m[539])|(m[533]&~m[536]&m[537]&~m[538]&m[539])|(~m[533]&~m[536]&~m[537]&m[538]&m[539])|(m[533]&~m[536]&~m[537]&m[538]&m[539])|(~m[533]&m[536]&~m[537]&m[538]&m[539])|(m[533]&m[536]&~m[537]&m[538]&m[539])|(~m[533]&~m[536]&m[537]&m[538]&m[539])|(m[533]&~m[536]&m[537]&m[538]&m[539])|(m[533]&m[536]&m[537]&m[538]&m[539]));
    m[540] = (((m[269]&~m[541]&~m[542]&~m[543]&~m[544])|(~m[269]&~m[541]&~m[542]&m[543]&~m[544])|(m[269]&m[541]&~m[542]&m[543]&~m[544])|(m[269]&~m[541]&m[542]&m[543]&~m[544])|(~m[269]&m[541]&~m[542]&~m[543]&m[544])|(~m[269]&~m[541]&m[542]&~m[543]&m[544])|(m[269]&m[541]&m[542]&~m[543]&m[544])|(~m[269]&m[541]&m[542]&m[543]&m[544]))&UnbiasedRNG[55])|((m[269]&~m[541]&~m[542]&m[543]&~m[544])|(~m[269]&~m[541]&~m[542]&~m[543]&m[544])|(m[269]&~m[541]&~m[542]&~m[543]&m[544])|(m[269]&m[541]&~m[542]&~m[543]&m[544])|(m[269]&~m[541]&m[542]&~m[543]&m[544])|(~m[269]&~m[541]&~m[542]&m[543]&m[544])|(m[269]&~m[541]&~m[542]&m[543]&m[544])|(~m[269]&m[541]&~m[542]&m[543]&m[544])|(m[269]&m[541]&~m[542]&m[543]&m[544])|(~m[269]&~m[541]&m[542]&m[543]&m[544])|(m[269]&~m[541]&m[542]&m[543]&m[544])|(m[269]&m[541]&m[542]&m[543]&m[544]));
    m[545] = (((m[543]&~m[546]&~m[547]&~m[548]&~m[549])|(~m[543]&~m[546]&~m[547]&m[548]&~m[549])|(m[543]&m[546]&~m[547]&m[548]&~m[549])|(m[543]&~m[546]&m[547]&m[548]&~m[549])|(~m[543]&m[546]&~m[547]&~m[548]&m[549])|(~m[543]&~m[546]&m[547]&~m[548]&m[549])|(m[543]&m[546]&m[547]&~m[548]&m[549])|(~m[543]&m[546]&m[547]&m[548]&m[549]))&UnbiasedRNG[56])|((m[543]&~m[546]&~m[547]&m[548]&~m[549])|(~m[543]&~m[546]&~m[547]&~m[548]&m[549])|(m[543]&~m[546]&~m[547]&~m[548]&m[549])|(m[543]&m[546]&~m[547]&~m[548]&m[549])|(m[543]&~m[546]&m[547]&~m[548]&m[549])|(~m[543]&~m[546]&~m[547]&m[548]&m[549])|(m[543]&~m[546]&~m[547]&m[548]&m[549])|(~m[543]&m[546]&~m[547]&m[548]&m[549])|(m[543]&m[546]&~m[547]&m[548]&m[549])|(~m[543]&~m[546]&m[547]&m[548]&m[549])|(m[543]&~m[546]&m[547]&m[548]&m[549])|(m[543]&m[546]&m[547]&m[548]&m[549]));
    m[550] = (((m[548]&~m[551]&~m[552]&~m[553]&~m[554])|(~m[548]&~m[551]&~m[552]&m[553]&~m[554])|(m[548]&m[551]&~m[552]&m[553]&~m[554])|(m[548]&~m[551]&m[552]&m[553]&~m[554])|(~m[548]&m[551]&~m[552]&~m[553]&m[554])|(~m[548]&~m[551]&m[552]&~m[553]&m[554])|(m[548]&m[551]&m[552]&~m[553]&m[554])|(~m[548]&m[551]&m[552]&m[553]&m[554]))&UnbiasedRNG[57])|((m[548]&~m[551]&~m[552]&m[553]&~m[554])|(~m[548]&~m[551]&~m[552]&~m[553]&m[554])|(m[548]&~m[551]&~m[552]&~m[553]&m[554])|(m[548]&m[551]&~m[552]&~m[553]&m[554])|(m[548]&~m[551]&m[552]&~m[553]&m[554])|(~m[548]&~m[551]&~m[552]&m[553]&m[554])|(m[548]&~m[551]&~m[552]&m[553]&m[554])|(~m[548]&m[551]&~m[552]&m[553]&m[554])|(m[548]&m[551]&~m[552]&m[553]&m[554])|(~m[548]&~m[551]&m[552]&m[553]&m[554])|(m[548]&~m[551]&m[552]&m[553]&m[554])|(m[548]&m[551]&m[552]&m[553]&m[554]));
    m[555] = (((m[553]&~m[556]&~m[557]&~m[558]&~m[559])|(~m[553]&~m[556]&~m[557]&m[558]&~m[559])|(m[553]&m[556]&~m[557]&m[558]&~m[559])|(m[553]&~m[556]&m[557]&m[558]&~m[559])|(~m[553]&m[556]&~m[557]&~m[558]&m[559])|(~m[553]&~m[556]&m[557]&~m[558]&m[559])|(m[553]&m[556]&m[557]&~m[558]&m[559])|(~m[553]&m[556]&m[557]&m[558]&m[559]))&UnbiasedRNG[58])|((m[553]&~m[556]&~m[557]&m[558]&~m[559])|(~m[553]&~m[556]&~m[557]&~m[558]&m[559])|(m[553]&~m[556]&~m[557]&~m[558]&m[559])|(m[553]&m[556]&~m[557]&~m[558]&m[559])|(m[553]&~m[556]&m[557]&~m[558]&m[559])|(~m[553]&~m[556]&~m[557]&m[558]&m[559])|(m[553]&~m[556]&~m[557]&m[558]&m[559])|(~m[553]&m[556]&~m[557]&m[558]&m[559])|(m[553]&m[556]&~m[557]&m[558]&m[559])|(~m[553]&~m[556]&m[557]&m[558]&m[559])|(m[553]&~m[556]&m[557]&m[558]&m[559])|(m[553]&m[556]&m[557]&m[558]&m[559]));
    m[560] = (((m[558]&~m[561]&~m[562]&~m[563]&~m[564])|(~m[558]&~m[561]&~m[562]&m[563]&~m[564])|(m[558]&m[561]&~m[562]&m[563]&~m[564])|(m[558]&~m[561]&m[562]&m[563]&~m[564])|(~m[558]&m[561]&~m[562]&~m[563]&m[564])|(~m[558]&~m[561]&m[562]&~m[563]&m[564])|(m[558]&m[561]&m[562]&~m[563]&m[564])|(~m[558]&m[561]&m[562]&m[563]&m[564]))&UnbiasedRNG[59])|((m[558]&~m[561]&~m[562]&m[563]&~m[564])|(~m[558]&~m[561]&~m[562]&~m[563]&m[564])|(m[558]&~m[561]&~m[562]&~m[563]&m[564])|(m[558]&m[561]&~m[562]&~m[563]&m[564])|(m[558]&~m[561]&m[562]&~m[563]&m[564])|(~m[558]&~m[561]&~m[562]&m[563]&m[564])|(m[558]&~m[561]&~m[562]&m[563]&m[564])|(~m[558]&m[561]&~m[562]&m[563]&m[564])|(m[558]&m[561]&~m[562]&m[563]&m[564])|(~m[558]&~m[561]&m[562]&m[563]&m[564])|(m[558]&~m[561]&m[562]&m[563]&m[564])|(m[558]&m[561]&m[562]&m[563]&m[564]));
    m[565] = (((m[563]&~m[566]&~m[567]&~m[568]&~m[569])|(~m[563]&~m[566]&~m[567]&m[568]&~m[569])|(m[563]&m[566]&~m[567]&m[568]&~m[569])|(m[563]&~m[566]&m[567]&m[568]&~m[569])|(~m[563]&m[566]&~m[567]&~m[568]&m[569])|(~m[563]&~m[566]&m[567]&~m[568]&m[569])|(m[563]&m[566]&m[567]&~m[568]&m[569])|(~m[563]&m[566]&m[567]&m[568]&m[569]))&UnbiasedRNG[60])|((m[563]&~m[566]&~m[567]&m[568]&~m[569])|(~m[563]&~m[566]&~m[567]&~m[568]&m[569])|(m[563]&~m[566]&~m[567]&~m[568]&m[569])|(m[563]&m[566]&~m[567]&~m[568]&m[569])|(m[563]&~m[566]&m[567]&~m[568]&m[569])|(~m[563]&~m[566]&~m[567]&m[568]&m[569])|(m[563]&~m[566]&~m[567]&m[568]&m[569])|(~m[563]&m[566]&~m[567]&m[568]&m[569])|(m[563]&m[566]&~m[567]&m[568]&m[569])|(~m[563]&~m[566]&m[567]&m[568]&m[569])|(m[563]&~m[566]&m[567]&m[568]&m[569])|(m[563]&m[566]&m[567]&m[568]&m[569]));
    m[570] = (((m[568]&~m[571]&~m[572]&~m[573]&~m[574])|(~m[568]&~m[571]&~m[572]&m[573]&~m[574])|(m[568]&m[571]&~m[572]&m[573]&~m[574])|(m[568]&~m[571]&m[572]&m[573]&~m[574])|(~m[568]&m[571]&~m[572]&~m[573]&m[574])|(~m[568]&~m[571]&m[572]&~m[573]&m[574])|(m[568]&m[571]&m[572]&~m[573]&m[574])|(~m[568]&m[571]&m[572]&m[573]&m[574]))&UnbiasedRNG[61])|((m[568]&~m[571]&~m[572]&m[573]&~m[574])|(~m[568]&~m[571]&~m[572]&~m[573]&m[574])|(m[568]&~m[571]&~m[572]&~m[573]&m[574])|(m[568]&m[571]&~m[572]&~m[573]&m[574])|(m[568]&~m[571]&m[572]&~m[573]&m[574])|(~m[568]&~m[571]&~m[572]&m[573]&m[574])|(m[568]&~m[571]&~m[572]&m[573]&m[574])|(~m[568]&m[571]&~m[572]&m[573]&m[574])|(m[568]&m[571]&~m[572]&m[573]&m[574])|(~m[568]&~m[571]&m[572]&m[573]&m[574])|(m[568]&~m[571]&m[572]&m[573]&m[574])|(m[568]&m[571]&m[572]&m[573]&m[574]));
    m[575] = (((m[573]&~m[576]&~m[577]&~m[578]&~m[579])|(~m[573]&~m[576]&~m[577]&m[578]&~m[579])|(m[573]&m[576]&~m[577]&m[578]&~m[579])|(m[573]&~m[576]&m[577]&m[578]&~m[579])|(~m[573]&m[576]&~m[577]&~m[578]&m[579])|(~m[573]&~m[576]&m[577]&~m[578]&m[579])|(m[573]&m[576]&m[577]&~m[578]&m[579])|(~m[573]&m[576]&m[577]&m[578]&m[579]))&UnbiasedRNG[62])|((m[573]&~m[576]&~m[577]&m[578]&~m[579])|(~m[573]&~m[576]&~m[577]&~m[578]&m[579])|(m[573]&~m[576]&~m[577]&~m[578]&m[579])|(m[573]&m[576]&~m[577]&~m[578]&m[579])|(m[573]&~m[576]&m[577]&~m[578]&m[579])|(~m[573]&~m[576]&~m[577]&m[578]&m[579])|(m[573]&~m[576]&~m[577]&m[578]&m[579])|(~m[573]&m[576]&~m[577]&m[578]&m[579])|(m[573]&m[576]&~m[577]&m[578]&m[579])|(~m[573]&~m[576]&m[577]&m[578]&m[579])|(m[573]&~m[576]&m[577]&m[578]&m[579])|(m[573]&m[576]&m[577]&m[578]&m[579]));
    m[580] = (((m[578]&~m[581]&~m[582]&~m[583]&~m[584])|(~m[578]&~m[581]&~m[582]&m[583]&~m[584])|(m[578]&m[581]&~m[582]&m[583]&~m[584])|(m[578]&~m[581]&m[582]&m[583]&~m[584])|(~m[578]&m[581]&~m[582]&~m[583]&m[584])|(~m[578]&~m[581]&m[582]&~m[583]&m[584])|(m[578]&m[581]&m[582]&~m[583]&m[584])|(~m[578]&m[581]&m[582]&m[583]&m[584]))&UnbiasedRNG[63])|((m[578]&~m[581]&~m[582]&m[583]&~m[584])|(~m[578]&~m[581]&~m[582]&~m[583]&m[584])|(m[578]&~m[581]&~m[582]&~m[583]&m[584])|(m[578]&m[581]&~m[582]&~m[583]&m[584])|(m[578]&~m[581]&m[582]&~m[583]&m[584])|(~m[578]&~m[581]&~m[582]&m[583]&m[584])|(m[578]&~m[581]&~m[582]&m[583]&m[584])|(~m[578]&m[581]&~m[582]&m[583]&m[584])|(m[578]&m[581]&~m[582]&m[583]&m[584])|(~m[578]&~m[581]&m[582]&m[583]&m[584])|(m[578]&~m[581]&m[582]&m[583]&m[584])|(m[578]&m[581]&m[582]&m[583]&m[584]));
    m[590] = (((m[588]&~m[591]&~m[592]&~m[593]&~m[594])|(~m[588]&~m[591]&~m[592]&m[593]&~m[594])|(m[588]&m[591]&~m[592]&m[593]&~m[594])|(m[588]&~m[591]&m[592]&m[593]&~m[594])|(~m[588]&m[591]&~m[592]&~m[593]&m[594])|(~m[588]&~m[591]&m[592]&~m[593]&m[594])|(m[588]&m[591]&m[592]&~m[593]&m[594])|(~m[588]&m[591]&m[592]&m[593]&m[594]))&UnbiasedRNG[64])|((m[588]&~m[591]&~m[592]&m[593]&~m[594])|(~m[588]&~m[591]&~m[592]&~m[593]&m[594])|(m[588]&~m[591]&~m[592]&~m[593]&m[594])|(m[588]&m[591]&~m[592]&~m[593]&m[594])|(m[588]&~m[591]&m[592]&~m[593]&m[594])|(~m[588]&~m[591]&~m[592]&m[593]&m[594])|(m[588]&~m[591]&~m[592]&m[593]&m[594])|(~m[588]&m[591]&~m[592]&m[593]&m[594])|(m[588]&m[591]&~m[592]&m[593]&m[594])|(~m[588]&~m[591]&m[592]&m[593]&m[594])|(m[588]&~m[591]&m[592]&m[593]&m[594])|(m[588]&m[591]&m[592]&m[593]&m[594]));
    m[595] = (((m[593]&~m[596]&~m[597]&~m[598]&~m[599])|(~m[593]&~m[596]&~m[597]&m[598]&~m[599])|(m[593]&m[596]&~m[597]&m[598]&~m[599])|(m[593]&~m[596]&m[597]&m[598]&~m[599])|(~m[593]&m[596]&~m[597]&~m[598]&m[599])|(~m[593]&~m[596]&m[597]&~m[598]&m[599])|(m[593]&m[596]&m[597]&~m[598]&m[599])|(~m[593]&m[596]&m[597]&m[598]&m[599]))&UnbiasedRNG[65])|((m[593]&~m[596]&~m[597]&m[598]&~m[599])|(~m[593]&~m[596]&~m[597]&~m[598]&m[599])|(m[593]&~m[596]&~m[597]&~m[598]&m[599])|(m[593]&m[596]&~m[597]&~m[598]&m[599])|(m[593]&~m[596]&m[597]&~m[598]&m[599])|(~m[593]&~m[596]&~m[597]&m[598]&m[599])|(m[593]&~m[596]&~m[597]&m[598]&m[599])|(~m[593]&m[596]&~m[597]&m[598]&m[599])|(m[593]&m[596]&~m[597]&m[598]&m[599])|(~m[593]&~m[596]&m[597]&m[598]&m[599])|(m[593]&~m[596]&m[597]&m[598]&m[599])|(m[593]&m[596]&m[597]&m[598]&m[599]));
    m[600] = (((m[598]&~m[601]&~m[602]&~m[603]&~m[604])|(~m[598]&~m[601]&~m[602]&m[603]&~m[604])|(m[598]&m[601]&~m[602]&m[603]&~m[604])|(m[598]&~m[601]&m[602]&m[603]&~m[604])|(~m[598]&m[601]&~m[602]&~m[603]&m[604])|(~m[598]&~m[601]&m[602]&~m[603]&m[604])|(m[598]&m[601]&m[602]&~m[603]&m[604])|(~m[598]&m[601]&m[602]&m[603]&m[604]))&UnbiasedRNG[66])|((m[598]&~m[601]&~m[602]&m[603]&~m[604])|(~m[598]&~m[601]&~m[602]&~m[603]&m[604])|(m[598]&~m[601]&~m[602]&~m[603]&m[604])|(m[598]&m[601]&~m[602]&~m[603]&m[604])|(m[598]&~m[601]&m[602]&~m[603]&m[604])|(~m[598]&~m[601]&~m[602]&m[603]&m[604])|(m[598]&~m[601]&~m[602]&m[603]&m[604])|(~m[598]&m[601]&~m[602]&m[603]&m[604])|(m[598]&m[601]&~m[602]&m[603]&m[604])|(~m[598]&~m[601]&m[602]&m[603]&m[604])|(m[598]&~m[601]&m[602]&m[603]&m[604])|(m[598]&m[601]&m[602]&m[603]&m[604]));
    m[605] = (((m[603]&~m[606]&~m[607]&~m[608]&~m[609])|(~m[603]&~m[606]&~m[607]&m[608]&~m[609])|(m[603]&m[606]&~m[607]&m[608]&~m[609])|(m[603]&~m[606]&m[607]&m[608]&~m[609])|(~m[603]&m[606]&~m[607]&~m[608]&m[609])|(~m[603]&~m[606]&m[607]&~m[608]&m[609])|(m[603]&m[606]&m[607]&~m[608]&m[609])|(~m[603]&m[606]&m[607]&m[608]&m[609]))&UnbiasedRNG[67])|((m[603]&~m[606]&~m[607]&m[608]&~m[609])|(~m[603]&~m[606]&~m[607]&~m[608]&m[609])|(m[603]&~m[606]&~m[607]&~m[608]&m[609])|(m[603]&m[606]&~m[607]&~m[608]&m[609])|(m[603]&~m[606]&m[607]&~m[608]&m[609])|(~m[603]&~m[606]&~m[607]&m[608]&m[609])|(m[603]&~m[606]&~m[607]&m[608]&m[609])|(~m[603]&m[606]&~m[607]&m[608]&m[609])|(m[603]&m[606]&~m[607]&m[608]&m[609])|(~m[603]&~m[606]&m[607]&m[608]&m[609])|(m[603]&~m[606]&m[607]&m[608]&m[609])|(m[603]&m[606]&m[607]&m[608]&m[609]));
    m[610] = (((m[608]&~m[611]&~m[612]&~m[613]&~m[614])|(~m[608]&~m[611]&~m[612]&m[613]&~m[614])|(m[608]&m[611]&~m[612]&m[613]&~m[614])|(m[608]&~m[611]&m[612]&m[613]&~m[614])|(~m[608]&m[611]&~m[612]&~m[613]&m[614])|(~m[608]&~m[611]&m[612]&~m[613]&m[614])|(m[608]&m[611]&m[612]&~m[613]&m[614])|(~m[608]&m[611]&m[612]&m[613]&m[614]))&UnbiasedRNG[68])|((m[608]&~m[611]&~m[612]&m[613]&~m[614])|(~m[608]&~m[611]&~m[612]&~m[613]&m[614])|(m[608]&~m[611]&~m[612]&~m[613]&m[614])|(m[608]&m[611]&~m[612]&~m[613]&m[614])|(m[608]&~m[611]&m[612]&~m[613]&m[614])|(~m[608]&~m[611]&~m[612]&m[613]&m[614])|(m[608]&~m[611]&~m[612]&m[613]&m[614])|(~m[608]&m[611]&~m[612]&m[613]&m[614])|(m[608]&m[611]&~m[612]&m[613]&m[614])|(~m[608]&~m[611]&m[612]&m[613]&m[614])|(m[608]&~m[611]&m[612]&m[613]&m[614])|(m[608]&m[611]&m[612]&m[613]&m[614]));
    m[615] = (((m[613]&~m[616]&~m[617]&~m[618]&~m[619])|(~m[613]&~m[616]&~m[617]&m[618]&~m[619])|(m[613]&m[616]&~m[617]&m[618]&~m[619])|(m[613]&~m[616]&m[617]&m[618]&~m[619])|(~m[613]&m[616]&~m[617]&~m[618]&m[619])|(~m[613]&~m[616]&m[617]&~m[618]&m[619])|(m[613]&m[616]&m[617]&~m[618]&m[619])|(~m[613]&m[616]&m[617]&m[618]&m[619]))&UnbiasedRNG[69])|((m[613]&~m[616]&~m[617]&m[618]&~m[619])|(~m[613]&~m[616]&~m[617]&~m[618]&m[619])|(m[613]&~m[616]&~m[617]&~m[618]&m[619])|(m[613]&m[616]&~m[617]&~m[618]&m[619])|(m[613]&~m[616]&m[617]&~m[618]&m[619])|(~m[613]&~m[616]&~m[617]&m[618]&m[619])|(m[613]&~m[616]&~m[617]&m[618]&m[619])|(~m[613]&m[616]&~m[617]&m[618]&m[619])|(m[613]&m[616]&~m[617]&m[618]&m[619])|(~m[613]&~m[616]&m[617]&m[618]&m[619])|(m[613]&~m[616]&m[617]&m[618]&m[619])|(m[613]&m[616]&m[617]&m[618]&m[619]));
    m[620] = (((m[618]&~m[621]&~m[622]&~m[623]&~m[624])|(~m[618]&~m[621]&~m[622]&m[623]&~m[624])|(m[618]&m[621]&~m[622]&m[623]&~m[624])|(m[618]&~m[621]&m[622]&m[623]&~m[624])|(~m[618]&m[621]&~m[622]&~m[623]&m[624])|(~m[618]&~m[621]&m[622]&~m[623]&m[624])|(m[618]&m[621]&m[622]&~m[623]&m[624])|(~m[618]&m[621]&m[622]&m[623]&m[624]))&UnbiasedRNG[70])|((m[618]&~m[621]&~m[622]&m[623]&~m[624])|(~m[618]&~m[621]&~m[622]&~m[623]&m[624])|(m[618]&~m[621]&~m[622]&~m[623]&m[624])|(m[618]&m[621]&~m[622]&~m[623]&m[624])|(m[618]&~m[621]&m[622]&~m[623]&m[624])|(~m[618]&~m[621]&~m[622]&m[623]&m[624])|(m[618]&~m[621]&~m[622]&m[623]&m[624])|(~m[618]&m[621]&~m[622]&m[623]&m[624])|(m[618]&m[621]&~m[622]&m[623]&m[624])|(~m[618]&~m[621]&m[622]&m[623]&m[624])|(m[618]&~m[621]&m[622]&m[623]&m[624])|(m[618]&m[621]&m[622]&m[623]&m[624]));
    m[625] = (((m[623]&~m[626]&~m[627]&~m[628]&~m[629])|(~m[623]&~m[626]&~m[627]&m[628]&~m[629])|(m[623]&m[626]&~m[627]&m[628]&~m[629])|(m[623]&~m[626]&m[627]&m[628]&~m[629])|(~m[623]&m[626]&~m[627]&~m[628]&m[629])|(~m[623]&~m[626]&m[627]&~m[628]&m[629])|(m[623]&m[626]&m[627]&~m[628]&m[629])|(~m[623]&m[626]&m[627]&m[628]&m[629]))&UnbiasedRNG[71])|((m[623]&~m[626]&~m[627]&m[628]&~m[629])|(~m[623]&~m[626]&~m[627]&~m[628]&m[629])|(m[623]&~m[626]&~m[627]&~m[628]&m[629])|(m[623]&m[626]&~m[627]&~m[628]&m[629])|(m[623]&~m[626]&m[627]&~m[628]&m[629])|(~m[623]&~m[626]&~m[627]&m[628]&m[629])|(m[623]&~m[626]&~m[627]&m[628]&m[629])|(~m[623]&m[626]&~m[627]&m[628]&m[629])|(m[623]&m[626]&~m[627]&m[628]&m[629])|(~m[623]&~m[626]&m[627]&m[628]&m[629])|(m[623]&~m[626]&m[627]&m[628]&m[629])|(m[623]&m[626]&m[627]&m[628]&m[629]));
    m[630] = (((m[589]&~m[631]&~m[632]&~m[633]&~m[634])|(~m[589]&~m[631]&~m[632]&m[633]&~m[634])|(m[589]&m[631]&~m[632]&m[633]&~m[634])|(m[589]&~m[631]&m[632]&m[633]&~m[634])|(~m[589]&m[631]&~m[632]&~m[633]&m[634])|(~m[589]&~m[631]&m[632]&~m[633]&m[634])|(m[589]&m[631]&m[632]&~m[633]&m[634])|(~m[589]&m[631]&m[632]&m[633]&m[634]))&UnbiasedRNG[72])|((m[589]&~m[631]&~m[632]&m[633]&~m[634])|(~m[589]&~m[631]&~m[632]&~m[633]&m[634])|(m[589]&~m[631]&~m[632]&~m[633]&m[634])|(m[589]&m[631]&~m[632]&~m[633]&m[634])|(m[589]&~m[631]&m[632]&~m[633]&m[634])|(~m[589]&~m[631]&~m[632]&m[633]&m[634])|(m[589]&~m[631]&~m[632]&m[633]&m[634])|(~m[589]&m[631]&~m[632]&m[633]&m[634])|(m[589]&m[631]&~m[632]&m[633]&m[634])|(~m[589]&~m[631]&m[632]&m[633]&m[634])|(m[589]&~m[631]&m[632]&m[633]&m[634])|(m[589]&m[631]&m[632]&m[633]&m[634]));
    m[635] = (((m[633]&~m[636]&~m[637]&~m[638]&~m[639])|(~m[633]&~m[636]&~m[637]&m[638]&~m[639])|(m[633]&m[636]&~m[637]&m[638]&~m[639])|(m[633]&~m[636]&m[637]&m[638]&~m[639])|(~m[633]&m[636]&~m[637]&~m[638]&m[639])|(~m[633]&~m[636]&m[637]&~m[638]&m[639])|(m[633]&m[636]&m[637]&~m[638]&m[639])|(~m[633]&m[636]&m[637]&m[638]&m[639]))&UnbiasedRNG[73])|((m[633]&~m[636]&~m[637]&m[638]&~m[639])|(~m[633]&~m[636]&~m[637]&~m[638]&m[639])|(m[633]&~m[636]&~m[637]&~m[638]&m[639])|(m[633]&m[636]&~m[637]&~m[638]&m[639])|(m[633]&~m[636]&m[637]&~m[638]&m[639])|(~m[633]&~m[636]&~m[637]&m[638]&m[639])|(m[633]&~m[636]&~m[637]&m[638]&m[639])|(~m[633]&m[636]&~m[637]&m[638]&m[639])|(m[633]&m[636]&~m[637]&m[638]&m[639])|(~m[633]&~m[636]&m[637]&m[638]&m[639])|(m[633]&~m[636]&m[637]&m[638]&m[639])|(m[633]&m[636]&m[637]&m[638]&m[639]));
    m[640] = (((m[638]&~m[641]&~m[642]&~m[643]&~m[644])|(~m[638]&~m[641]&~m[642]&m[643]&~m[644])|(m[638]&m[641]&~m[642]&m[643]&~m[644])|(m[638]&~m[641]&m[642]&m[643]&~m[644])|(~m[638]&m[641]&~m[642]&~m[643]&m[644])|(~m[638]&~m[641]&m[642]&~m[643]&m[644])|(m[638]&m[641]&m[642]&~m[643]&m[644])|(~m[638]&m[641]&m[642]&m[643]&m[644]))&UnbiasedRNG[74])|((m[638]&~m[641]&~m[642]&m[643]&~m[644])|(~m[638]&~m[641]&~m[642]&~m[643]&m[644])|(m[638]&~m[641]&~m[642]&~m[643]&m[644])|(m[638]&m[641]&~m[642]&~m[643]&m[644])|(m[638]&~m[641]&m[642]&~m[643]&m[644])|(~m[638]&~m[641]&~m[642]&m[643]&m[644])|(m[638]&~m[641]&~m[642]&m[643]&m[644])|(~m[638]&m[641]&~m[642]&m[643]&m[644])|(m[638]&m[641]&~m[642]&m[643]&m[644])|(~m[638]&~m[641]&m[642]&m[643]&m[644])|(m[638]&~m[641]&m[642]&m[643]&m[644])|(m[638]&m[641]&m[642]&m[643]&m[644]));
    m[645] = (((m[643]&~m[646]&~m[647]&~m[648]&~m[649])|(~m[643]&~m[646]&~m[647]&m[648]&~m[649])|(m[643]&m[646]&~m[647]&m[648]&~m[649])|(m[643]&~m[646]&m[647]&m[648]&~m[649])|(~m[643]&m[646]&~m[647]&~m[648]&m[649])|(~m[643]&~m[646]&m[647]&~m[648]&m[649])|(m[643]&m[646]&m[647]&~m[648]&m[649])|(~m[643]&m[646]&m[647]&m[648]&m[649]))&UnbiasedRNG[75])|((m[643]&~m[646]&~m[647]&m[648]&~m[649])|(~m[643]&~m[646]&~m[647]&~m[648]&m[649])|(m[643]&~m[646]&~m[647]&~m[648]&m[649])|(m[643]&m[646]&~m[647]&~m[648]&m[649])|(m[643]&~m[646]&m[647]&~m[648]&m[649])|(~m[643]&~m[646]&~m[647]&m[648]&m[649])|(m[643]&~m[646]&~m[647]&m[648]&m[649])|(~m[643]&m[646]&~m[647]&m[648]&m[649])|(m[643]&m[646]&~m[647]&m[648]&m[649])|(~m[643]&~m[646]&m[647]&m[648]&m[649])|(m[643]&~m[646]&m[647]&m[648]&m[649])|(m[643]&m[646]&m[647]&m[648]&m[649]));
    m[650] = (((m[648]&~m[651]&~m[652]&~m[653]&~m[654])|(~m[648]&~m[651]&~m[652]&m[653]&~m[654])|(m[648]&m[651]&~m[652]&m[653]&~m[654])|(m[648]&~m[651]&m[652]&m[653]&~m[654])|(~m[648]&m[651]&~m[652]&~m[653]&m[654])|(~m[648]&~m[651]&m[652]&~m[653]&m[654])|(m[648]&m[651]&m[652]&~m[653]&m[654])|(~m[648]&m[651]&m[652]&m[653]&m[654]))&UnbiasedRNG[76])|((m[648]&~m[651]&~m[652]&m[653]&~m[654])|(~m[648]&~m[651]&~m[652]&~m[653]&m[654])|(m[648]&~m[651]&~m[652]&~m[653]&m[654])|(m[648]&m[651]&~m[652]&~m[653]&m[654])|(m[648]&~m[651]&m[652]&~m[653]&m[654])|(~m[648]&~m[651]&~m[652]&m[653]&m[654])|(m[648]&~m[651]&~m[652]&m[653]&m[654])|(~m[648]&m[651]&~m[652]&m[653]&m[654])|(m[648]&m[651]&~m[652]&m[653]&m[654])|(~m[648]&~m[651]&m[652]&m[653]&m[654])|(m[648]&~m[651]&m[652]&m[653]&m[654])|(m[648]&m[651]&m[652]&m[653]&m[654]));
    m[655] = (((m[653]&~m[656]&~m[657]&~m[658]&~m[659])|(~m[653]&~m[656]&~m[657]&m[658]&~m[659])|(m[653]&m[656]&~m[657]&m[658]&~m[659])|(m[653]&~m[656]&m[657]&m[658]&~m[659])|(~m[653]&m[656]&~m[657]&~m[658]&m[659])|(~m[653]&~m[656]&m[657]&~m[658]&m[659])|(m[653]&m[656]&m[657]&~m[658]&m[659])|(~m[653]&m[656]&m[657]&m[658]&m[659]))&UnbiasedRNG[77])|((m[653]&~m[656]&~m[657]&m[658]&~m[659])|(~m[653]&~m[656]&~m[657]&~m[658]&m[659])|(m[653]&~m[656]&~m[657]&~m[658]&m[659])|(m[653]&m[656]&~m[657]&~m[658]&m[659])|(m[653]&~m[656]&m[657]&~m[658]&m[659])|(~m[653]&~m[656]&~m[657]&m[658]&m[659])|(m[653]&~m[656]&~m[657]&m[658]&m[659])|(~m[653]&m[656]&~m[657]&m[658]&m[659])|(m[653]&m[656]&~m[657]&m[658]&m[659])|(~m[653]&~m[656]&m[657]&m[658]&m[659])|(m[653]&~m[656]&m[657]&m[658]&m[659])|(m[653]&m[656]&m[657]&m[658]&m[659]));
    m[660] = (((m[658]&~m[661]&~m[662]&~m[663]&~m[664])|(~m[658]&~m[661]&~m[662]&m[663]&~m[664])|(m[658]&m[661]&~m[662]&m[663]&~m[664])|(m[658]&~m[661]&m[662]&m[663]&~m[664])|(~m[658]&m[661]&~m[662]&~m[663]&m[664])|(~m[658]&~m[661]&m[662]&~m[663]&m[664])|(m[658]&m[661]&m[662]&~m[663]&m[664])|(~m[658]&m[661]&m[662]&m[663]&m[664]))&UnbiasedRNG[78])|((m[658]&~m[661]&~m[662]&m[663]&~m[664])|(~m[658]&~m[661]&~m[662]&~m[663]&m[664])|(m[658]&~m[661]&~m[662]&~m[663]&m[664])|(m[658]&m[661]&~m[662]&~m[663]&m[664])|(m[658]&~m[661]&m[662]&~m[663]&m[664])|(~m[658]&~m[661]&~m[662]&m[663]&m[664])|(m[658]&~m[661]&~m[662]&m[663]&m[664])|(~m[658]&m[661]&~m[662]&m[663]&m[664])|(m[658]&m[661]&~m[662]&m[663]&m[664])|(~m[658]&~m[661]&m[662]&m[663]&m[664])|(m[658]&~m[661]&m[662]&m[663]&m[664])|(m[658]&m[661]&m[662]&m[663]&m[664]));
    m[665] = (((m[663]&~m[666]&~m[667]&~m[668]&~m[669])|(~m[663]&~m[666]&~m[667]&m[668]&~m[669])|(m[663]&m[666]&~m[667]&m[668]&~m[669])|(m[663]&~m[666]&m[667]&m[668]&~m[669])|(~m[663]&m[666]&~m[667]&~m[668]&m[669])|(~m[663]&~m[666]&m[667]&~m[668]&m[669])|(m[663]&m[666]&m[667]&~m[668]&m[669])|(~m[663]&m[666]&m[667]&m[668]&m[669]))&UnbiasedRNG[79])|((m[663]&~m[666]&~m[667]&m[668]&~m[669])|(~m[663]&~m[666]&~m[667]&~m[668]&m[669])|(m[663]&~m[666]&~m[667]&~m[668]&m[669])|(m[663]&m[666]&~m[667]&~m[668]&m[669])|(m[663]&~m[666]&m[667]&~m[668]&m[669])|(~m[663]&~m[666]&~m[667]&m[668]&m[669])|(m[663]&~m[666]&~m[667]&m[668]&m[669])|(~m[663]&m[666]&~m[667]&m[668]&m[669])|(m[663]&m[666]&~m[667]&m[668]&m[669])|(~m[663]&~m[666]&m[667]&m[668]&m[669])|(m[663]&~m[666]&m[667]&m[668]&m[669])|(m[663]&m[666]&m[667]&m[668]&m[669]));
    m[670] = (((m[634]&~m[671]&~m[672]&~m[673]&~m[674])|(~m[634]&~m[671]&~m[672]&m[673]&~m[674])|(m[634]&m[671]&~m[672]&m[673]&~m[674])|(m[634]&~m[671]&m[672]&m[673]&~m[674])|(~m[634]&m[671]&~m[672]&~m[673]&m[674])|(~m[634]&~m[671]&m[672]&~m[673]&m[674])|(m[634]&m[671]&m[672]&~m[673]&m[674])|(~m[634]&m[671]&m[672]&m[673]&m[674]))&UnbiasedRNG[80])|((m[634]&~m[671]&~m[672]&m[673]&~m[674])|(~m[634]&~m[671]&~m[672]&~m[673]&m[674])|(m[634]&~m[671]&~m[672]&~m[673]&m[674])|(m[634]&m[671]&~m[672]&~m[673]&m[674])|(m[634]&~m[671]&m[672]&~m[673]&m[674])|(~m[634]&~m[671]&~m[672]&m[673]&m[674])|(m[634]&~m[671]&~m[672]&m[673]&m[674])|(~m[634]&m[671]&~m[672]&m[673]&m[674])|(m[634]&m[671]&~m[672]&m[673]&m[674])|(~m[634]&~m[671]&m[672]&m[673]&m[674])|(m[634]&~m[671]&m[672]&m[673]&m[674])|(m[634]&m[671]&m[672]&m[673]&m[674]));
    m[675] = (((m[673]&~m[676]&~m[677]&~m[678]&~m[679])|(~m[673]&~m[676]&~m[677]&m[678]&~m[679])|(m[673]&m[676]&~m[677]&m[678]&~m[679])|(m[673]&~m[676]&m[677]&m[678]&~m[679])|(~m[673]&m[676]&~m[677]&~m[678]&m[679])|(~m[673]&~m[676]&m[677]&~m[678]&m[679])|(m[673]&m[676]&m[677]&~m[678]&m[679])|(~m[673]&m[676]&m[677]&m[678]&m[679]))&UnbiasedRNG[81])|((m[673]&~m[676]&~m[677]&m[678]&~m[679])|(~m[673]&~m[676]&~m[677]&~m[678]&m[679])|(m[673]&~m[676]&~m[677]&~m[678]&m[679])|(m[673]&m[676]&~m[677]&~m[678]&m[679])|(m[673]&~m[676]&m[677]&~m[678]&m[679])|(~m[673]&~m[676]&~m[677]&m[678]&m[679])|(m[673]&~m[676]&~m[677]&m[678]&m[679])|(~m[673]&m[676]&~m[677]&m[678]&m[679])|(m[673]&m[676]&~m[677]&m[678]&m[679])|(~m[673]&~m[676]&m[677]&m[678]&m[679])|(m[673]&~m[676]&m[677]&m[678]&m[679])|(m[673]&m[676]&m[677]&m[678]&m[679]));
    m[680] = (((m[678]&~m[681]&~m[682]&~m[683]&~m[684])|(~m[678]&~m[681]&~m[682]&m[683]&~m[684])|(m[678]&m[681]&~m[682]&m[683]&~m[684])|(m[678]&~m[681]&m[682]&m[683]&~m[684])|(~m[678]&m[681]&~m[682]&~m[683]&m[684])|(~m[678]&~m[681]&m[682]&~m[683]&m[684])|(m[678]&m[681]&m[682]&~m[683]&m[684])|(~m[678]&m[681]&m[682]&m[683]&m[684]))&UnbiasedRNG[82])|((m[678]&~m[681]&~m[682]&m[683]&~m[684])|(~m[678]&~m[681]&~m[682]&~m[683]&m[684])|(m[678]&~m[681]&~m[682]&~m[683]&m[684])|(m[678]&m[681]&~m[682]&~m[683]&m[684])|(m[678]&~m[681]&m[682]&~m[683]&m[684])|(~m[678]&~m[681]&~m[682]&m[683]&m[684])|(m[678]&~m[681]&~m[682]&m[683]&m[684])|(~m[678]&m[681]&~m[682]&m[683]&m[684])|(m[678]&m[681]&~m[682]&m[683]&m[684])|(~m[678]&~m[681]&m[682]&m[683]&m[684])|(m[678]&~m[681]&m[682]&m[683]&m[684])|(m[678]&m[681]&m[682]&m[683]&m[684]));
    m[685] = (((m[683]&~m[686]&~m[687]&~m[688]&~m[689])|(~m[683]&~m[686]&~m[687]&m[688]&~m[689])|(m[683]&m[686]&~m[687]&m[688]&~m[689])|(m[683]&~m[686]&m[687]&m[688]&~m[689])|(~m[683]&m[686]&~m[687]&~m[688]&m[689])|(~m[683]&~m[686]&m[687]&~m[688]&m[689])|(m[683]&m[686]&m[687]&~m[688]&m[689])|(~m[683]&m[686]&m[687]&m[688]&m[689]))&UnbiasedRNG[83])|((m[683]&~m[686]&~m[687]&m[688]&~m[689])|(~m[683]&~m[686]&~m[687]&~m[688]&m[689])|(m[683]&~m[686]&~m[687]&~m[688]&m[689])|(m[683]&m[686]&~m[687]&~m[688]&m[689])|(m[683]&~m[686]&m[687]&~m[688]&m[689])|(~m[683]&~m[686]&~m[687]&m[688]&m[689])|(m[683]&~m[686]&~m[687]&m[688]&m[689])|(~m[683]&m[686]&~m[687]&m[688]&m[689])|(m[683]&m[686]&~m[687]&m[688]&m[689])|(~m[683]&~m[686]&m[687]&m[688]&m[689])|(m[683]&~m[686]&m[687]&m[688]&m[689])|(m[683]&m[686]&m[687]&m[688]&m[689]));
    m[690] = (((m[688]&~m[691]&~m[692]&~m[693]&~m[694])|(~m[688]&~m[691]&~m[692]&m[693]&~m[694])|(m[688]&m[691]&~m[692]&m[693]&~m[694])|(m[688]&~m[691]&m[692]&m[693]&~m[694])|(~m[688]&m[691]&~m[692]&~m[693]&m[694])|(~m[688]&~m[691]&m[692]&~m[693]&m[694])|(m[688]&m[691]&m[692]&~m[693]&m[694])|(~m[688]&m[691]&m[692]&m[693]&m[694]))&UnbiasedRNG[84])|((m[688]&~m[691]&~m[692]&m[693]&~m[694])|(~m[688]&~m[691]&~m[692]&~m[693]&m[694])|(m[688]&~m[691]&~m[692]&~m[693]&m[694])|(m[688]&m[691]&~m[692]&~m[693]&m[694])|(m[688]&~m[691]&m[692]&~m[693]&m[694])|(~m[688]&~m[691]&~m[692]&m[693]&m[694])|(m[688]&~m[691]&~m[692]&m[693]&m[694])|(~m[688]&m[691]&~m[692]&m[693]&m[694])|(m[688]&m[691]&~m[692]&m[693]&m[694])|(~m[688]&~m[691]&m[692]&m[693]&m[694])|(m[688]&~m[691]&m[692]&m[693]&m[694])|(m[688]&m[691]&m[692]&m[693]&m[694]));
    m[695] = (((m[693]&~m[696]&~m[697]&~m[698]&~m[699])|(~m[693]&~m[696]&~m[697]&m[698]&~m[699])|(m[693]&m[696]&~m[697]&m[698]&~m[699])|(m[693]&~m[696]&m[697]&m[698]&~m[699])|(~m[693]&m[696]&~m[697]&~m[698]&m[699])|(~m[693]&~m[696]&m[697]&~m[698]&m[699])|(m[693]&m[696]&m[697]&~m[698]&m[699])|(~m[693]&m[696]&m[697]&m[698]&m[699]))&UnbiasedRNG[85])|((m[693]&~m[696]&~m[697]&m[698]&~m[699])|(~m[693]&~m[696]&~m[697]&~m[698]&m[699])|(m[693]&~m[696]&~m[697]&~m[698]&m[699])|(m[693]&m[696]&~m[697]&~m[698]&m[699])|(m[693]&~m[696]&m[697]&~m[698]&m[699])|(~m[693]&~m[696]&~m[697]&m[698]&m[699])|(m[693]&~m[696]&~m[697]&m[698]&m[699])|(~m[693]&m[696]&~m[697]&m[698]&m[699])|(m[693]&m[696]&~m[697]&m[698]&m[699])|(~m[693]&~m[696]&m[697]&m[698]&m[699])|(m[693]&~m[696]&m[697]&m[698]&m[699])|(m[693]&m[696]&m[697]&m[698]&m[699]));
    m[700] = (((m[698]&~m[701]&~m[702]&~m[703]&~m[704])|(~m[698]&~m[701]&~m[702]&m[703]&~m[704])|(m[698]&m[701]&~m[702]&m[703]&~m[704])|(m[698]&~m[701]&m[702]&m[703]&~m[704])|(~m[698]&m[701]&~m[702]&~m[703]&m[704])|(~m[698]&~m[701]&m[702]&~m[703]&m[704])|(m[698]&m[701]&m[702]&~m[703]&m[704])|(~m[698]&m[701]&m[702]&m[703]&m[704]))&UnbiasedRNG[86])|((m[698]&~m[701]&~m[702]&m[703]&~m[704])|(~m[698]&~m[701]&~m[702]&~m[703]&m[704])|(m[698]&~m[701]&~m[702]&~m[703]&m[704])|(m[698]&m[701]&~m[702]&~m[703]&m[704])|(m[698]&~m[701]&m[702]&~m[703]&m[704])|(~m[698]&~m[701]&~m[702]&m[703]&m[704])|(m[698]&~m[701]&~m[702]&m[703]&m[704])|(~m[698]&m[701]&~m[702]&m[703]&m[704])|(m[698]&m[701]&~m[702]&m[703]&m[704])|(~m[698]&~m[701]&m[702]&m[703]&m[704])|(m[698]&~m[701]&m[702]&m[703]&m[704])|(m[698]&m[701]&m[702]&m[703]&m[704]));
    m[705] = (((m[674]&~m[706]&~m[707]&~m[708]&~m[709])|(~m[674]&~m[706]&~m[707]&m[708]&~m[709])|(m[674]&m[706]&~m[707]&m[708]&~m[709])|(m[674]&~m[706]&m[707]&m[708]&~m[709])|(~m[674]&m[706]&~m[707]&~m[708]&m[709])|(~m[674]&~m[706]&m[707]&~m[708]&m[709])|(m[674]&m[706]&m[707]&~m[708]&m[709])|(~m[674]&m[706]&m[707]&m[708]&m[709]))&UnbiasedRNG[87])|((m[674]&~m[706]&~m[707]&m[708]&~m[709])|(~m[674]&~m[706]&~m[707]&~m[708]&m[709])|(m[674]&~m[706]&~m[707]&~m[708]&m[709])|(m[674]&m[706]&~m[707]&~m[708]&m[709])|(m[674]&~m[706]&m[707]&~m[708]&m[709])|(~m[674]&~m[706]&~m[707]&m[708]&m[709])|(m[674]&~m[706]&~m[707]&m[708]&m[709])|(~m[674]&m[706]&~m[707]&m[708]&m[709])|(m[674]&m[706]&~m[707]&m[708]&m[709])|(~m[674]&~m[706]&m[707]&m[708]&m[709])|(m[674]&~m[706]&m[707]&m[708]&m[709])|(m[674]&m[706]&m[707]&m[708]&m[709]));
    m[710] = (((m[708]&~m[711]&~m[712]&~m[713]&~m[714])|(~m[708]&~m[711]&~m[712]&m[713]&~m[714])|(m[708]&m[711]&~m[712]&m[713]&~m[714])|(m[708]&~m[711]&m[712]&m[713]&~m[714])|(~m[708]&m[711]&~m[712]&~m[713]&m[714])|(~m[708]&~m[711]&m[712]&~m[713]&m[714])|(m[708]&m[711]&m[712]&~m[713]&m[714])|(~m[708]&m[711]&m[712]&m[713]&m[714]))&UnbiasedRNG[88])|((m[708]&~m[711]&~m[712]&m[713]&~m[714])|(~m[708]&~m[711]&~m[712]&~m[713]&m[714])|(m[708]&~m[711]&~m[712]&~m[713]&m[714])|(m[708]&m[711]&~m[712]&~m[713]&m[714])|(m[708]&~m[711]&m[712]&~m[713]&m[714])|(~m[708]&~m[711]&~m[712]&m[713]&m[714])|(m[708]&~m[711]&~m[712]&m[713]&m[714])|(~m[708]&m[711]&~m[712]&m[713]&m[714])|(m[708]&m[711]&~m[712]&m[713]&m[714])|(~m[708]&~m[711]&m[712]&m[713]&m[714])|(m[708]&~m[711]&m[712]&m[713]&m[714])|(m[708]&m[711]&m[712]&m[713]&m[714]));
    m[715] = (((m[713]&~m[716]&~m[717]&~m[718]&~m[719])|(~m[713]&~m[716]&~m[717]&m[718]&~m[719])|(m[713]&m[716]&~m[717]&m[718]&~m[719])|(m[713]&~m[716]&m[717]&m[718]&~m[719])|(~m[713]&m[716]&~m[717]&~m[718]&m[719])|(~m[713]&~m[716]&m[717]&~m[718]&m[719])|(m[713]&m[716]&m[717]&~m[718]&m[719])|(~m[713]&m[716]&m[717]&m[718]&m[719]))&UnbiasedRNG[89])|((m[713]&~m[716]&~m[717]&m[718]&~m[719])|(~m[713]&~m[716]&~m[717]&~m[718]&m[719])|(m[713]&~m[716]&~m[717]&~m[718]&m[719])|(m[713]&m[716]&~m[717]&~m[718]&m[719])|(m[713]&~m[716]&m[717]&~m[718]&m[719])|(~m[713]&~m[716]&~m[717]&m[718]&m[719])|(m[713]&~m[716]&~m[717]&m[718]&m[719])|(~m[713]&m[716]&~m[717]&m[718]&m[719])|(m[713]&m[716]&~m[717]&m[718]&m[719])|(~m[713]&~m[716]&m[717]&m[718]&m[719])|(m[713]&~m[716]&m[717]&m[718]&m[719])|(m[713]&m[716]&m[717]&m[718]&m[719]));
    m[720] = (((m[718]&~m[721]&~m[722]&~m[723]&~m[724])|(~m[718]&~m[721]&~m[722]&m[723]&~m[724])|(m[718]&m[721]&~m[722]&m[723]&~m[724])|(m[718]&~m[721]&m[722]&m[723]&~m[724])|(~m[718]&m[721]&~m[722]&~m[723]&m[724])|(~m[718]&~m[721]&m[722]&~m[723]&m[724])|(m[718]&m[721]&m[722]&~m[723]&m[724])|(~m[718]&m[721]&m[722]&m[723]&m[724]))&UnbiasedRNG[90])|((m[718]&~m[721]&~m[722]&m[723]&~m[724])|(~m[718]&~m[721]&~m[722]&~m[723]&m[724])|(m[718]&~m[721]&~m[722]&~m[723]&m[724])|(m[718]&m[721]&~m[722]&~m[723]&m[724])|(m[718]&~m[721]&m[722]&~m[723]&m[724])|(~m[718]&~m[721]&~m[722]&m[723]&m[724])|(m[718]&~m[721]&~m[722]&m[723]&m[724])|(~m[718]&m[721]&~m[722]&m[723]&m[724])|(m[718]&m[721]&~m[722]&m[723]&m[724])|(~m[718]&~m[721]&m[722]&m[723]&m[724])|(m[718]&~m[721]&m[722]&m[723]&m[724])|(m[718]&m[721]&m[722]&m[723]&m[724]));
    m[725] = (((m[723]&~m[726]&~m[727]&~m[728]&~m[729])|(~m[723]&~m[726]&~m[727]&m[728]&~m[729])|(m[723]&m[726]&~m[727]&m[728]&~m[729])|(m[723]&~m[726]&m[727]&m[728]&~m[729])|(~m[723]&m[726]&~m[727]&~m[728]&m[729])|(~m[723]&~m[726]&m[727]&~m[728]&m[729])|(m[723]&m[726]&m[727]&~m[728]&m[729])|(~m[723]&m[726]&m[727]&m[728]&m[729]))&UnbiasedRNG[91])|((m[723]&~m[726]&~m[727]&m[728]&~m[729])|(~m[723]&~m[726]&~m[727]&~m[728]&m[729])|(m[723]&~m[726]&~m[727]&~m[728]&m[729])|(m[723]&m[726]&~m[727]&~m[728]&m[729])|(m[723]&~m[726]&m[727]&~m[728]&m[729])|(~m[723]&~m[726]&~m[727]&m[728]&m[729])|(m[723]&~m[726]&~m[727]&m[728]&m[729])|(~m[723]&m[726]&~m[727]&m[728]&m[729])|(m[723]&m[726]&~m[727]&m[728]&m[729])|(~m[723]&~m[726]&m[727]&m[728]&m[729])|(m[723]&~m[726]&m[727]&m[728]&m[729])|(m[723]&m[726]&m[727]&m[728]&m[729]));
    m[730] = (((m[728]&~m[731]&~m[732]&~m[733]&~m[734])|(~m[728]&~m[731]&~m[732]&m[733]&~m[734])|(m[728]&m[731]&~m[732]&m[733]&~m[734])|(m[728]&~m[731]&m[732]&m[733]&~m[734])|(~m[728]&m[731]&~m[732]&~m[733]&m[734])|(~m[728]&~m[731]&m[732]&~m[733]&m[734])|(m[728]&m[731]&m[732]&~m[733]&m[734])|(~m[728]&m[731]&m[732]&m[733]&m[734]))&UnbiasedRNG[92])|((m[728]&~m[731]&~m[732]&m[733]&~m[734])|(~m[728]&~m[731]&~m[732]&~m[733]&m[734])|(m[728]&~m[731]&~m[732]&~m[733]&m[734])|(m[728]&m[731]&~m[732]&~m[733]&m[734])|(m[728]&~m[731]&m[732]&~m[733]&m[734])|(~m[728]&~m[731]&~m[732]&m[733]&m[734])|(m[728]&~m[731]&~m[732]&m[733]&m[734])|(~m[728]&m[731]&~m[732]&m[733]&m[734])|(m[728]&m[731]&~m[732]&m[733]&m[734])|(~m[728]&~m[731]&m[732]&m[733]&m[734])|(m[728]&~m[731]&m[732]&m[733]&m[734])|(m[728]&m[731]&m[732]&m[733]&m[734]));
    m[735] = (((m[709]&~m[736]&~m[737]&~m[738]&~m[739])|(~m[709]&~m[736]&~m[737]&m[738]&~m[739])|(m[709]&m[736]&~m[737]&m[738]&~m[739])|(m[709]&~m[736]&m[737]&m[738]&~m[739])|(~m[709]&m[736]&~m[737]&~m[738]&m[739])|(~m[709]&~m[736]&m[737]&~m[738]&m[739])|(m[709]&m[736]&m[737]&~m[738]&m[739])|(~m[709]&m[736]&m[737]&m[738]&m[739]))&UnbiasedRNG[93])|((m[709]&~m[736]&~m[737]&m[738]&~m[739])|(~m[709]&~m[736]&~m[737]&~m[738]&m[739])|(m[709]&~m[736]&~m[737]&~m[738]&m[739])|(m[709]&m[736]&~m[737]&~m[738]&m[739])|(m[709]&~m[736]&m[737]&~m[738]&m[739])|(~m[709]&~m[736]&~m[737]&m[738]&m[739])|(m[709]&~m[736]&~m[737]&m[738]&m[739])|(~m[709]&m[736]&~m[737]&m[738]&m[739])|(m[709]&m[736]&~m[737]&m[738]&m[739])|(~m[709]&~m[736]&m[737]&m[738]&m[739])|(m[709]&~m[736]&m[737]&m[738]&m[739])|(m[709]&m[736]&m[737]&m[738]&m[739]));
    m[740] = (((m[738]&~m[741]&~m[742]&~m[743]&~m[744])|(~m[738]&~m[741]&~m[742]&m[743]&~m[744])|(m[738]&m[741]&~m[742]&m[743]&~m[744])|(m[738]&~m[741]&m[742]&m[743]&~m[744])|(~m[738]&m[741]&~m[742]&~m[743]&m[744])|(~m[738]&~m[741]&m[742]&~m[743]&m[744])|(m[738]&m[741]&m[742]&~m[743]&m[744])|(~m[738]&m[741]&m[742]&m[743]&m[744]))&UnbiasedRNG[94])|((m[738]&~m[741]&~m[742]&m[743]&~m[744])|(~m[738]&~m[741]&~m[742]&~m[743]&m[744])|(m[738]&~m[741]&~m[742]&~m[743]&m[744])|(m[738]&m[741]&~m[742]&~m[743]&m[744])|(m[738]&~m[741]&m[742]&~m[743]&m[744])|(~m[738]&~m[741]&~m[742]&m[743]&m[744])|(m[738]&~m[741]&~m[742]&m[743]&m[744])|(~m[738]&m[741]&~m[742]&m[743]&m[744])|(m[738]&m[741]&~m[742]&m[743]&m[744])|(~m[738]&~m[741]&m[742]&m[743]&m[744])|(m[738]&~m[741]&m[742]&m[743]&m[744])|(m[738]&m[741]&m[742]&m[743]&m[744]));
    m[745] = (((m[743]&~m[746]&~m[747]&~m[748]&~m[749])|(~m[743]&~m[746]&~m[747]&m[748]&~m[749])|(m[743]&m[746]&~m[747]&m[748]&~m[749])|(m[743]&~m[746]&m[747]&m[748]&~m[749])|(~m[743]&m[746]&~m[747]&~m[748]&m[749])|(~m[743]&~m[746]&m[747]&~m[748]&m[749])|(m[743]&m[746]&m[747]&~m[748]&m[749])|(~m[743]&m[746]&m[747]&m[748]&m[749]))&UnbiasedRNG[95])|((m[743]&~m[746]&~m[747]&m[748]&~m[749])|(~m[743]&~m[746]&~m[747]&~m[748]&m[749])|(m[743]&~m[746]&~m[747]&~m[748]&m[749])|(m[743]&m[746]&~m[747]&~m[748]&m[749])|(m[743]&~m[746]&m[747]&~m[748]&m[749])|(~m[743]&~m[746]&~m[747]&m[748]&m[749])|(m[743]&~m[746]&~m[747]&m[748]&m[749])|(~m[743]&m[746]&~m[747]&m[748]&m[749])|(m[743]&m[746]&~m[747]&m[748]&m[749])|(~m[743]&~m[746]&m[747]&m[748]&m[749])|(m[743]&~m[746]&m[747]&m[748]&m[749])|(m[743]&m[746]&m[747]&m[748]&m[749]));
    m[750] = (((m[748]&~m[751]&~m[752]&~m[753]&~m[754])|(~m[748]&~m[751]&~m[752]&m[753]&~m[754])|(m[748]&m[751]&~m[752]&m[753]&~m[754])|(m[748]&~m[751]&m[752]&m[753]&~m[754])|(~m[748]&m[751]&~m[752]&~m[753]&m[754])|(~m[748]&~m[751]&m[752]&~m[753]&m[754])|(m[748]&m[751]&m[752]&~m[753]&m[754])|(~m[748]&m[751]&m[752]&m[753]&m[754]))&UnbiasedRNG[96])|((m[748]&~m[751]&~m[752]&m[753]&~m[754])|(~m[748]&~m[751]&~m[752]&~m[753]&m[754])|(m[748]&~m[751]&~m[752]&~m[753]&m[754])|(m[748]&m[751]&~m[752]&~m[753]&m[754])|(m[748]&~m[751]&m[752]&~m[753]&m[754])|(~m[748]&~m[751]&~m[752]&m[753]&m[754])|(m[748]&~m[751]&~m[752]&m[753]&m[754])|(~m[748]&m[751]&~m[752]&m[753]&m[754])|(m[748]&m[751]&~m[752]&m[753]&m[754])|(~m[748]&~m[751]&m[752]&m[753]&m[754])|(m[748]&~m[751]&m[752]&m[753]&m[754])|(m[748]&m[751]&m[752]&m[753]&m[754]));
    m[755] = (((m[753]&~m[756]&~m[757]&~m[758]&~m[759])|(~m[753]&~m[756]&~m[757]&m[758]&~m[759])|(m[753]&m[756]&~m[757]&m[758]&~m[759])|(m[753]&~m[756]&m[757]&m[758]&~m[759])|(~m[753]&m[756]&~m[757]&~m[758]&m[759])|(~m[753]&~m[756]&m[757]&~m[758]&m[759])|(m[753]&m[756]&m[757]&~m[758]&m[759])|(~m[753]&m[756]&m[757]&m[758]&m[759]))&UnbiasedRNG[97])|((m[753]&~m[756]&~m[757]&m[758]&~m[759])|(~m[753]&~m[756]&~m[757]&~m[758]&m[759])|(m[753]&~m[756]&~m[757]&~m[758]&m[759])|(m[753]&m[756]&~m[757]&~m[758]&m[759])|(m[753]&~m[756]&m[757]&~m[758]&m[759])|(~m[753]&~m[756]&~m[757]&m[758]&m[759])|(m[753]&~m[756]&~m[757]&m[758]&m[759])|(~m[753]&m[756]&~m[757]&m[758]&m[759])|(m[753]&m[756]&~m[757]&m[758]&m[759])|(~m[753]&~m[756]&m[757]&m[758]&m[759])|(m[753]&~m[756]&m[757]&m[758]&m[759])|(m[753]&m[756]&m[757]&m[758]&m[759]));
    m[760] = (((m[739]&~m[761]&~m[762]&~m[763]&~m[764])|(~m[739]&~m[761]&~m[762]&m[763]&~m[764])|(m[739]&m[761]&~m[762]&m[763]&~m[764])|(m[739]&~m[761]&m[762]&m[763]&~m[764])|(~m[739]&m[761]&~m[762]&~m[763]&m[764])|(~m[739]&~m[761]&m[762]&~m[763]&m[764])|(m[739]&m[761]&m[762]&~m[763]&m[764])|(~m[739]&m[761]&m[762]&m[763]&m[764]))&UnbiasedRNG[98])|((m[739]&~m[761]&~m[762]&m[763]&~m[764])|(~m[739]&~m[761]&~m[762]&~m[763]&m[764])|(m[739]&~m[761]&~m[762]&~m[763]&m[764])|(m[739]&m[761]&~m[762]&~m[763]&m[764])|(m[739]&~m[761]&m[762]&~m[763]&m[764])|(~m[739]&~m[761]&~m[762]&m[763]&m[764])|(m[739]&~m[761]&~m[762]&m[763]&m[764])|(~m[739]&m[761]&~m[762]&m[763]&m[764])|(m[739]&m[761]&~m[762]&m[763]&m[764])|(~m[739]&~m[761]&m[762]&m[763]&m[764])|(m[739]&~m[761]&m[762]&m[763]&m[764])|(m[739]&m[761]&m[762]&m[763]&m[764]));
    m[765] = (((m[763]&~m[766]&~m[767]&~m[768]&~m[769])|(~m[763]&~m[766]&~m[767]&m[768]&~m[769])|(m[763]&m[766]&~m[767]&m[768]&~m[769])|(m[763]&~m[766]&m[767]&m[768]&~m[769])|(~m[763]&m[766]&~m[767]&~m[768]&m[769])|(~m[763]&~m[766]&m[767]&~m[768]&m[769])|(m[763]&m[766]&m[767]&~m[768]&m[769])|(~m[763]&m[766]&m[767]&m[768]&m[769]))&UnbiasedRNG[99])|((m[763]&~m[766]&~m[767]&m[768]&~m[769])|(~m[763]&~m[766]&~m[767]&~m[768]&m[769])|(m[763]&~m[766]&~m[767]&~m[768]&m[769])|(m[763]&m[766]&~m[767]&~m[768]&m[769])|(m[763]&~m[766]&m[767]&~m[768]&m[769])|(~m[763]&~m[766]&~m[767]&m[768]&m[769])|(m[763]&~m[766]&~m[767]&m[768]&m[769])|(~m[763]&m[766]&~m[767]&m[768]&m[769])|(m[763]&m[766]&~m[767]&m[768]&m[769])|(~m[763]&~m[766]&m[767]&m[768]&m[769])|(m[763]&~m[766]&m[767]&m[768]&m[769])|(m[763]&m[766]&m[767]&m[768]&m[769]));
    m[770] = (((m[768]&~m[771]&~m[772]&~m[773]&~m[774])|(~m[768]&~m[771]&~m[772]&m[773]&~m[774])|(m[768]&m[771]&~m[772]&m[773]&~m[774])|(m[768]&~m[771]&m[772]&m[773]&~m[774])|(~m[768]&m[771]&~m[772]&~m[773]&m[774])|(~m[768]&~m[771]&m[772]&~m[773]&m[774])|(m[768]&m[771]&m[772]&~m[773]&m[774])|(~m[768]&m[771]&m[772]&m[773]&m[774]))&UnbiasedRNG[100])|((m[768]&~m[771]&~m[772]&m[773]&~m[774])|(~m[768]&~m[771]&~m[772]&~m[773]&m[774])|(m[768]&~m[771]&~m[772]&~m[773]&m[774])|(m[768]&m[771]&~m[772]&~m[773]&m[774])|(m[768]&~m[771]&m[772]&~m[773]&m[774])|(~m[768]&~m[771]&~m[772]&m[773]&m[774])|(m[768]&~m[771]&~m[772]&m[773]&m[774])|(~m[768]&m[771]&~m[772]&m[773]&m[774])|(m[768]&m[771]&~m[772]&m[773]&m[774])|(~m[768]&~m[771]&m[772]&m[773]&m[774])|(m[768]&~m[771]&m[772]&m[773]&m[774])|(m[768]&m[771]&m[772]&m[773]&m[774]));
    m[775] = (((m[773]&~m[776]&~m[777]&~m[778]&~m[779])|(~m[773]&~m[776]&~m[777]&m[778]&~m[779])|(m[773]&m[776]&~m[777]&m[778]&~m[779])|(m[773]&~m[776]&m[777]&m[778]&~m[779])|(~m[773]&m[776]&~m[777]&~m[778]&m[779])|(~m[773]&~m[776]&m[777]&~m[778]&m[779])|(m[773]&m[776]&m[777]&~m[778]&m[779])|(~m[773]&m[776]&m[777]&m[778]&m[779]))&UnbiasedRNG[101])|((m[773]&~m[776]&~m[777]&m[778]&~m[779])|(~m[773]&~m[776]&~m[777]&~m[778]&m[779])|(m[773]&~m[776]&~m[777]&~m[778]&m[779])|(m[773]&m[776]&~m[777]&~m[778]&m[779])|(m[773]&~m[776]&m[777]&~m[778]&m[779])|(~m[773]&~m[776]&~m[777]&m[778]&m[779])|(m[773]&~m[776]&~m[777]&m[778]&m[779])|(~m[773]&m[776]&~m[777]&m[778]&m[779])|(m[773]&m[776]&~m[777]&m[778]&m[779])|(~m[773]&~m[776]&m[777]&m[778]&m[779])|(m[773]&~m[776]&m[777]&m[778]&m[779])|(m[773]&m[776]&m[777]&m[778]&m[779]));
    m[780] = (((m[764]&~m[781]&~m[782]&~m[783]&~m[784])|(~m[764]&~m[781]&~m[782]&m[783]&~m[784])|(m[764]&m[781]&~m[782]&m[783]&~m[784])|(m[764]&~m[781]&m[782]&m[783]&~m[784])|(~m[764]&m[781]&~m[782]&~m[783]&m[784])|(~m[764]&~m[781]&m[782]&~m[783]&m[784])|(m[764]&m[781]&m[782]&~m[783]&m[784])|(~m[764]&m[781]&m[782]&m[783]&m[784]))&UnbiasedRNG[102])|((m[764]&~m[781]&~m[782]&m[783]&~m[784])|(~m[764]&~m[781]&~m[782]&~m[783]&m[784])|(m[764]&~m[781]&~m[782]&~m[783]&m[784])|(m[764]&m[781]&~m[782]&~m[783]&m[784])|(m[764]&~m[781]&m[782]&~m[783]&m[784])|(~m[764]&~m[781]&~m[782]&m[783]&m[784])|(m[764]&~m[781]&~m[782]&m[783]&m[784])|(~m[764]&m[781]&~m[782]&m[783]&m[784])|(m[764]&m[781]&~m[782]&m[783]&m[784])|(~m[764]&~m[781]&m[782]&m[783]&m[784])|(m[764]&~m[781]&m[782]&m[783]&m[784])|(m[764]&m[781]&m[782]&m[783]&m[784]));
    m[785] = (((m[783]&~m[786]&~m[787]&~m[788]&~m[789])|(~m[783]&~m[786]&~m[787]&m[788]&~m[789])|(m[783]&m[786]&~m[787]&m[788]&~m[789])|(m[783]&~m[786]&m[787]&m[788]&~m[789])|(~m[783]&m[786]&~m[787]&~m[788]&m[789])|(~m[783]&~m[786]&m[787]&~m[788]&m[789])|(m[783]&m[786]&m[787]&~m[788]&m[789])|(~m[783]&m[786]&m[787]&m[788]&m[789]))&UnbiasedRNG[103])|((m[783]&~m[786]&~m[787]&m[788]&~m[789])|(~m[783]&~m[786]&~m[787]&~m[788]&m[789])|(m[783]&~m[786]&~m[787]&~m[788]&m[789])|(m[783]&m[786]&~m[787]&~m[788]&m[789])|(m[783]&~m[786]&m[787]&~m[788]&m[789])|(~m[783]&~m[786]&~m[787]&m[788]&m[789])|(m[783]&~m[786]&~m[787]&m[788]&m[789])|(~m[783]&m[786]&~m[787]&m[788]&m[789])|(m[783]&m[786]&~m[787]&m[788]&m[789])|(~m[783]&~m[786]&m[787]&m[788]&m[789])|(m[783]&~m[786]&m[787]&m[788]&m[789])|(m[783]&m[786]&m[787]&m[788]&m[789]));
    m[790] = (((m[788]&~m[791]&~m[792]&~m[793]&~m[794])|(~m[788]&~m[791]&~m[792]&m[793]&~m[794])|(m[788]&m[791]&~m[792]&m[793]&~m[794])|(m[788]&~m[791]&m[792]&m[793]&~m[794])|(~m[788]&m[791]&~m[792]&~m[793]&m[794])|(~m[788]&~m[791]&m[792]&~m[793]&m[794])|(m[788]&m[791]&m[792]&~m[793]&m[794])|(~m[788]&m[791]&m[792]&m[793]&m[794]))&UnbiasedRNG[104])|((m[788]&~m[791]&~m[792]&m[793]&~m[794])|(~m[788]&~m[791]&~m[792]&~m[793]&m[794])|(m[788]&~m[791]&~m[792]&~m[793]&m[794])|(m[788]&m[791]&~m[792]&~m[793]&m[794])|(m[788]&~m[791]&m[792]&~m[793]&m[794])|(~m[788]&~m[791]&~m[792]&m[793]&m[794])|(m[788]&~m[791]&~m[792]&m[793]&m[794])|(~m[788]&m[791]&~m[792]&m[793]&m[794])|(m[788]&m[791]&~m[792]&m[793]&m[794])|(~m[788]&~m[791]&m[792]&m[793]&m[794])|(m[788]&~m[791]&m[792]&m[793]&m[794])|(m[788]&m[791]&m[792]&m[793]&m[794]));
    m[795] = (((m[784]&~m[796]&~m[797]&~m[798]&~m[799])|(~m[784]&~m[796]&~m[797]&m[798]&~m[799])|(m[784]&m[796]&~m[797]&m[798]&~m[799])|(m[784]&~m[796]&m[797]&m[798]&~m[799])|(~m[784]&m[796]&~m[797]&~m[798]&m[799])|(~m[784]&~m[796]&m[797]&~m[798]&m[799])|(m[784]&m[796]&m[797]&~m[798]&m[799])|(~m[784]&m[796]&m[797]&m[798]&m[799]))&UnbiasedRNG[105])|((m[784]&~m[796]&~m[797]&m[798]&~m[799])|(~m[784]&~m[796]&~m[797]&~m[798]&m[799])|(m[784]&~m[796]&~m[797]&~m[798]&m[799])|(m[784]&m[796]&~m[797]&~m[798]&m[799])|(m[784]&~m[796]&m[797]&~m[798]&m[799])|(~m[784]&~m[796]&~m[797]&m[798]&m[799])|(m[784]&~m[796]&~m[797]&m[798]&m[799])|(~m[784]&m[796]&~m[797]&m[798]&m[799])|(m[784]&m[796]&~m[797]&m[798]&m[799])|(~m[784]&~m[796]&m[797]&m[798]&m[799])|(m[784]&~m[796]&m[797]&m[798]&m[799])|(m[784]&m[796]&m[797]&m[798]&m[799]));
    m[800] = (((m[798]&~m[801]&~m[802]&~m[803]&~m[804])|(~m[798]&~m[801]&~m[802]&m[803]&~m[804])|(m[798]&m[801]&~m[802]&m[803]&~m[804])|(m[798]&~m[801]&m[802]&m[803]&~m[804])|(~m[798]&m[801]&~m[802]&~m[803]&m[804])|(~m[798]&~m[801]&m[802]&~m[803]&m[804])|(m[798]&m[801]&m[802]&~m[803]&m[804])|(~m[798]&m[801]&m[802]&m[803]&m[804]))&UnbiasedRNG[106])|((m[798]&~m[801]&~m[802]&m[803]&~m[804])|(~m[798]&~m[801]&~m[802]&~m[803]&m[804])|(m[798]&~m[801]&~m[802]&~m[803]&m[804])|(m[798]&m[801]&~m[802]&~m[803]&m[804])|(m[798]&~m[801]&m[802]&~m[803]&m[804])|(~m[798]&~m[801]&~m[802]&m[803]&m[804])|(m[798]&~m[801]&~m[802]&m[803]&m[804])|(~m[798]&m[801]&~m[802]&m[803]&m[804])|(m[798]&m[801]&~m[802]&m[803]&m[804])|(~m[798]&~m[801]&m[802]&m[803]&m[804])|(m[798]&~m[801]&m[802]&m[803]&m[804])|(m[798]&m[801]&m[802]&m[803]&m[804]));
    m[805] = (((m[799]&~m[806]&~m[807]&~m[808]&~m[809])|(~m[799]&~m[806]&~m[807]&m[808]&~m[809])|(m[799]&m[806]&~m[807]&m[808]&~m[809])|(m[799]&~m[806]&m[807]&m[808]&~m[809])|(~m[799]&m[806]&~m[807]&~m[808]&m[809])|(~m[799]&~m[806]&m[807]&~m[808]&m[809])|(m[799]&m[806]&m[807]&~m[808]&m[809])|(~m[799]&m[806]&m[807]&m[808]&m[809]))&UnbiasedRNG[107])|((m[799]&~m[806]&~m[807]&m[808]&~m[809])|(~m[799]&~m[806]&~m[807]&~m[808]&m[809])|(m[799]&~m[806]&~m[807]&~m[808]&m[809])|(m[799]&m[806]&~m[807]&~m[808]&m[809])|(m[799]&~m[806]&m[807]&~m[808]&m[809])|(~m[799]&~m[806]&~m[807]&m[808]&m[809])|(m[799]&~m[806]&~m[807]&m[808]&m[809])|(~m[799]&m[806]&~m[807]&m[808]&m[809])|(m[799]&m[806]&~m[807]&m[808]&m[809])|(~m[799]&~m[806]&m[807]&m[808]&m[809])|(m[799]&~m[806]&m[807]&m[808]&m[809])|(m[799]&m[806]&m[807]&m[808]&m[809]));
end

always @(posedge color1_clk) begin
    m[20] = (((m[0]&m[62]&~m[63]&~m[64]&~m[65])|(m[0]&~m[62]&m[63]&~m[64]&~m[65])|(~m[0]&m[62]&m[63]&~m[64]&~m[65])|(m[0]&~m[62]&~m[63]&m[64]&~m[65])|(~m[0]&m[62]&~m[63]&m[64]&~m[65])|(~m[0]&~m[62]&m[63]&m[64]&~m[65])|(m[0]&~m[62]&~m[63]&~m[64]&m[65])|(~m[0]&m[62]&~m[63]&~m[64]&m[65])|(~m[0]&~m[62]&m[63]&~m[64]&m[65])|(~m[0]&~m[62]&~m[63]&m[64]&m[65]))&BiasedRNG[99])|(((m[0]&m[62]&m[63]&~m[64]&~m[65])|(m[0]&m[62]&~m[63]&m[64]&~m[65])|(m[0]&~m[62]&m[63]&m[64]&~m[65])|(~m[0]&m[62]&m[63]&m[64]&~m[65])|(m[0]&m[62]&~m[63]&~m[64]&m[65])|(m[0]&~m[62]&m[63]&~m[64]&m[65])|(~m[0]&m[62]&m[63]&~m[64]&m[65])|(m[0]&~m[62]&~m[63]&m[64]&m[65])|(~m[0]&m[62]&~m[63]&m[64]&m[65])|(~m[0]&~m[62]&m[63]&m[64]&m[65]))&~BiasedRNG[99])|((m[0]&m[62]&m[63]&m[64]&~m[65])|(m[0]&m[62]&m[63]&~m[64]&m[65])|(m[0]&m[62]&~m[63]&m[64]&m[65])|(m[0]&~m[62]&m[63]&m[64]&m[65])|(~m[0]&m[62]&m[63]&m[64]&m[65])|(m[0]&m[62]&m[63]&m[64]&m[65]));
    m[21] = (((m[0]&m[66]&~m[67]&~m[68]&~m[69])|(m[0]&~m[66]&m[67]&~m[68]&~m[69])|(~m[0]&m[66]&m[67]&~m[68]&~m[69])|(m[0]&~m[66]&~m[67]&m[68]&~m[69])|(~m[0]&m[66]&~m[67]&m[68]&~m[69])|(~m[0]&~m[66]&m[67]&m[68]&~m[69])|(m[0]&~m[66]&~m[67]&~m[68]&m[69])|(~m[0]&m[66]&~m[67]&~m[68]&m[69])|(~m[0]&~m[66]&m[67]&~m[68]&m[69])|(~m[0]&~m[66]&~m[67]&m[68]&m[69]))&BiasedRNG[100])|(((m[0]&m[66]&m[67]&~m[68]&~m[69])|(m[0]&m[66]&~m[67]&m[68]&~m[69])|(m[0]&~m[66]&m[67]&m[68]&~m[69])|(~m[0]&m[66]&m[67]&m[68]&~m[69])|(m[0]&m[66]&~m[67]&~m[68]&m[69])|(m[0]&~m[66]&m[67]&~m[68]&m[69])|(~m[0]&m[66]&m[67]&~m[68]&m[69])|(m[0]&~m[66]&~m[67]&m[68]&m[69])|(~m[0]&m[66]&~m[67]&m[68]&m[69])|(~m[0]&~m[66]&m[67]&m[68]&m[69]))&~BiasedRNG[100])|((m[0]&m[66]&m[67]&m[68]&~m[69])|(m[0]&m[66]&m[67]&~m[68]&m[69])|(m[0]&m[66]&~m[67]&m[68]&m[69])|(m[0]&~m[66]&m[67]&m[68]&m[69])|(~m[0]&m[66]&m[67]&m[68]&m[69])|(m[0]&m[66]&m[67]&m[68]&m[69]));
    m[22] = (((m[1]&m[72]&~m[73]&~m[74]&~m[75])|(m[1]&~m[72]&m[73]&~m[74]&~m[75])|(~m[1]&m[72]&m[73]&~m[74]&~m[75])|(m[1]&~m[72]&~m[73]&m[74]&~m[75])|(~m[1]&m[72]&~m[73]&m[74]&~m[75])|(~m[1]&~m[72]&m[73]&m[74]&~m[75])|(m[1]&~m[72]&~m[73]&~m[74]&m[75])|(~m[1]&m[72]&~m[73]&~m[74]&m[75])|(~m[1]&~m[72]&m[73]&~m[74]&m[75])|(~m[1]&~m[72]&~m[73]&m[74]&m[75]))&BiasedRNG[101])|(((m[1]&m[72]&m[73]&~m[74]&~m[75])|(m[1]&m[72]&~m[73]&m[74]&~m[75])|(m[1]&~m[72]&m[73]&m[74]&~m[75])|(~m[1]&m[72]&m[73]&m[74]&~m[75])|(m[1]&m[72]&~m[73]&~m[74]&m[75])|(m[1]&~m[72]&m[73]&~m[74]&m[75])|(~m[1]&m[72]&m[73]&~m[74]&m[75])|(m[1]&~m[72]&~m[73]&m[74]&m[75])|(~m[1]&m[72]&~m[73]&m[74]&m[75])|(~m[1]&~m[72]&m[73]&m[74]&m[75]))&~BiasedRNG[101])|((m[1]&m[72]&m[73]&m[74]&~m[75])|(m[1]&m[72]&m[73]&~m[74]&m[75])|(m[1]&m[72]&~m[73]&m[74]&m[75])|(m[1]&~m[72]&m[73]&m[74]&m[75])|(~m[1]&m[72]&m[73]&m[74]&m[75])|(m[1]&m[72]&m[73]&m[74]&m[75]));
    m[23] = (((m[1]&m[76]&~m[77]&~m[78]&~m[79])|(m[1]&~m[76]&m[77]&~m[78]&~m[79])|(~m[1]&m[76]&m[77]&~m[78]&~m[79])|(m[1]&~m[76]&~m[77]&m[78]&~m[79])|(~m[1]&m[76]&~m[77]&m[78]&~m[79])|(~m[1]&~m[76]&m[77]&m[78]&~m[79])|(m[1]&~m[76]&~m[77]&~m[78]&m[79])|(~m[1]&m[76]&~m[77]&~m[78]&m[79])|(~m[1]&~m[76]&m[77]&~m[78]&m[79])|(~m[1]&~m[76]&~m[77]&m[78]&m[79]))&BiasedRNG[102])|(((m[1]&m[76]&m[77]&~m[78]&~m[79])|(m[1]&m[76]&~m[77]&m[78]&~m[79])|(m[1]&~m[76]&m[77]&m[78]&~m[79])|(~m[1]&m[76]&m[77]&m[78]&~m[79])|(m[1]&m[76]&~m[77]&~m[78]&m[79])|(m[1]&~m[76]&m[77]&~m[78]&m[79])|(~m[1]&m[76]&m[77]&~m[78]&m[79])|(m[1]&~m[76]&~m[77]&m[78]&m[79])|(~m[1]&m[76]&~m[77]&m[78]&m[79])|(~m[1]&~m[76]&m[77]&m[78]&m[79]))&~BiasedRNG[102])|((m[1]&m[76]&m[77]&m[78]&~m[79])|(m[1]&m[76]&m[77]&~m[78]&m[79])|(m[1]&m[76]&~m[77]&m[78]&m[79])|(m[1]&~m[76]&m[77]&m[78]&m[79])|(~m[1]&m[76]&m[77]&m[78]&m[79])|(m[1]&m[76]&m[77]&m[78]&m[79]));
    m[24] = (((m[2]&m[82]&~m[83]&~m[84]&~m[85])|(m[2]&~m[82]&m[83]&~m[84]&~m[85])|(~m[2]&m[82]&m[83]&~m[84]&~m[85])|(m[2]&~m[82]&~m[83]&m[84]&~m[85])|(~m[2]&m[82]&~m[83]&m[84]&~m[85])|(~m[2]&~m[82]&m[83]&m[84]&~m[85])|(m[2]&~m[82]&~m[83]&~m[84]&m[85])|(~m[2]&m[82]&~m[83]&~m[84]&m[85])|(~m[2]&~m[82]&m[83]&~m[84]&m[85])|(~m[2]&~m[82]&~m[83]&m[84]&m[85]))&BiasedRNG[103])|(((m[2]&m[82]&m[83]&~m[84]&~m[85])|(m[2]&m[82]&~m[83]&m[84]&~m[85])|(m[2]&~m[82]&m[83]&m[84]&~m[85])|(~m[2]&m[82]&m[83]&m[84]&~m[85])|(m[2]&m[82]&~m[83]&~m[84]&m[85])|(m[2]&~m[82]&m[83]&~m[84]&m[85])|(~m[2]&m[82]&m[83]&~m[84]&m[85])|(m[2]&~m[82]&~m[83]&m[84]&m[85])|(~m[2]&m[82]&~m[83]&m[84]&m[85])|(~m[2]&~m[82]&m[83]&m[84]&m[85]))&~BiasedRNG[103])|((m[2]&m[82]&m[83]&m[84]&~m[85])|(m[2]&m[82]&m[83]&~m[84]&m[85])|(m[2]&m[82]&~m[83]&m[84]&m[85])|(m[2]&~m[82]&m[83]&m[84]&m[85])|(~m[2]&m[82]&m[83]&m[84]&m[85])|(m[2]&m[82]&m[83]&m[84]&m[85]));
    m[25] = (((m[2]&m[86]&~m[87]&~m[88]&~m[89])|(m[2]&~m[86]&m[87]&~m[88]&~m[89])|(~m[2]&m[86]&m[87]&~m[88]&~m[89])|(m[2]&~m[86]&~m[87]&m[88]&~m[89])|(~m[2]&m[86]&~m[87]&m[88]&~m[89])|(~m[2]&~m[86]&m[87]&m[88]&~m[89])|(m[2]&~m[86]&~m[87]&~m[88]&m[89])|(~m[2]&m[86]&~m[87]&~m[88]&m[89])|(~m[2]&~m[86]&m[87]&~m[88]&m[89])|(~m[2]&~m[86]&~m[87]&m[88]&m[89]))&BiasedRNG[104])|(((m[2]&m[86]&m[87]&~m[88]&~m[89])|(m[2]&m[86]&~m[87]&m[88]&~m[89])|(m[2]&~m[86]&m[87]&m[88]&~m[89])|(~m[2]&m[86]&m[87]&m[88]&~m[89])|(m[2]&m[86]&~m[87]&~m[88]&m[89])|(m[2]&~m[86]&m[87]&~m[88]&m[89])|(~m[2]&m[86]&m[87]&~m[88]&m[89])|(m[2]&~m[86]&~m[87]&m[88]&m[89])|(~m[2]&m[86]&~m[87]&m[88]&m[89])|(~m[2]&~m[86]&m[87]&m[88]&m[89]))&~BiasedRNG[104])|((m[2]&m[86]&m[87]&m[88]&~m[89])|(m[2]&m[86]&m[87]&~m[88]&m[89])|(m[2]&m[86]&~m[87]&m[88]&m[89])|(m[2]&~m[86]&m[87]&m[88]&m[89])|(~m[2]&m[86]&m[87]&m[88]&m[89])|(m[2]&m[86]&m[87]&m[88]&m[89]));
    m[26] = (((m[3]&m[92]&~m[93]&~m[94]&~m[95])|(m[3]&~m[92]&m[93]&~m[94]&~m[95])|(~m[3]&m[92]&m[93]&~m[94]&~m[95])|(m[3]&~m[92]&~m[93]&m[94]&~m[95])|(~m[3]&m[92]&~m[93]&m[94]&~m[95])|(~m[3]&~m[92]&m[93]&m[94]&~m[95])|(m[3]&~m[92]&~m[93]&~m[94]&m[95])|(~m[3]&m[92]&~m[93]&~m[94]&m[95])|(~m[3]&~m[92]&m[93]&~m[94]&m[95])|(~m[3]&~m[92]&~m[93]&m[94]&m[95]))&BiasedRNG[105])|(((m[3]&m[92]&m[93]&~m[94]&~m[95])|(m[3]&m[92]&~m[93]&m[94]&~m[95])|(m[3]&~m[92]&m[93]&m[94]&~m[95])|(~m[3]&m[92]&m[93]&m[94]&~m[95])|(m[3]&m[92]&~m[93]&~m[94]&m[95])|(m[3]&~m[92]&m[93]&~m[94]&m[95])|(~m[3]&m[92]&m[93]&~m[94]&m[95])|(m[3]&~m[92]&~m[93]&m[94]&m[95])|(~m[3]&m[92]&~m[93]&m[94]&m[95])|(~m[3]&~m[92]&m[93]&m[94]&m[95]))&~BiasedRNG[105])|((m[3]&m[92]&m[93]&m[94]&~m[95])|(m[3]&m[92]&m[93]&~m[94]&m[95])|(m[3]&m[92]&~m[93]&m[94]&m[95])|(m[3]&~m[92]&m[93]&m[94]&m[95])|(~m[3]&m[92]&m[93]&m[94]&m[95])|(m[3]&m[92]&m[93]&m[94]&m[95]));
    m[27] = (((m[3]&m[96]&~m[97]&~m[98]&~m[99])|(m[3]&~m[96]&m[97]&~m[98]&~m[99])|(~m[3]&m[96]&m[97]&~m[98]&~m[99])|(m[3]&~m[96]&~m[97]&m[98]&~m[99])|(~m[3]&m[96]&~m[97]&m[98]&~m[99])|(~m[3]&~m[96]&m[97]&m[98]&~m[99])|(m[3]&~m[96]&~m[97]&~m[98]&m[99])|(~m[3]&m[96]&~m[97]&~m[98]&m[99])|(~m[3]&~m[96]&m[97]&~m[98]&m[99])|(~m[3]&~m[96]&~m[97]&m[98]&m[99]))&BiasedRNG[106])|(((m[3]&m[96]&m[97]&~m[98]&~m[99])|(m[3]&m[96]&~m[97]&m[98]&~m[99])|(m[3]&~m[96]&m[97]&m[98]&~m[99])|(~m[3]&m[96]&m[97]&m[98]&~m[99])|(m[3]&m[96]&~m[97]&~m[98]&m[99])|(m[3]&~m[96]&m[97]&~m[98]&m[99])|(~m[3]&m[96]&m[97]&~m[98]&m[99])|(m[3]&~m[96]&~m[97]&m[98]&m[99])|(~m[3]&m[96]&~m[97]&m[98]&m[99])|(~m[3]&~m[96]&m[97]&m[98]&m[99]))&~BiasedRNG[106])|((m[3]&m[96]&m[97]&m[98]&~m[99])|(m[3]&m[96]&m[97]&~m[98]&m[99])|(m[3]&m[96]&~m[97]&m[98]&m[99])|(m[3]&~m[96]&m[97]&m[98]&m[99])|(~m[3]&m[96]&m[97]&m[98]&m[99])|(m[3]&m[96]&m[97]&m[98]&m[99]));
    m[28] = (((m[4]&m[102]&~m[103]&~m[104]&~m[105])|(m[4]&~m[102]&m[103]&~m[104]&~m[105])|(~m[4]&m[102]&m[103]&~m[104]&~m[105])|(m[4]&~m[102]&~m[103]&m[104]&~m[105])|(~m[4]&m[102]&~m[103]&m[104]&~m[105])|(~m[4]&~m[102]&m[103]&m[104]&~m[105])|(m[4]&~m[102]&~m[103]&~m[104]&m[105])|(~m[4]&m[102]&~m[103]&~m[104]&m[105])|(~m[4]&~m[102]&m[103]&~m[104]&m[105])|(~m[4]&~m[102]&~m[103]&m[104]&m[105]))&BiasedRNG[107])|(((m[4]&m[102]&m[103]&~m[104]&~m[105])|(m[4]&m[102]&~m[103]&m[104]&~m[105])|(m[4]&~m[102]&m[103]&m[104]&~m[105])|(~m[4]&m[102]&m[103]&m[104]&~m[105])|(m[4]&m[102]&~m[103]&~m[104]&m[105])|(m[4]&~m[102]&m[103]&~m[104]&m[105])|(~m[4]&m[102]&m[103]&~m[104]&m[105])|(m[4]&~m[102]&~m[103]&m[104]&m[105])|(~m[4]&m[102]&~m[103]&m[104]&m[105])|(~m[4]&~m[102]&m[103]&m[104]&m[105]))&~BiasedRNG[107])|((m[4]&m[102]&m[103]&m[104]&~m[105])|(m[4]&m[102]&m[103]&~m[104]&m[105])|(m[4]&m[102]&~m[103]&m[104]&m[105])|(m[4]&~m[102]&m[103]&m[104]&m[105])|(~m[4]&m[102]&m[103]&m[104]&m[105])|(m[4]&m[102]&m[103]&m[104]&m[105]));
    m[29] = (((m[4]&m[106]&~m[107]&~m[108]&~m[109])|(m[4]&~m[106]&m[107]&~m[108]&~m[109])|(~m[4]&m[106]&m[107]&~m[108]&~m[109])|(m[4]&~m[106]&~m[107]&m[108]&~m[109])|(~m[4]&m[106]&~m[107]&m[108]&~m[109])|(~m[4]&~m[106]&m[107]&m[108]&~m[109])|(m[4]&~m[106]&~m[107]&~m[108]&m[109])|(~m[4]&m[106]&~m[107]&~m[108]&m[109])|(~m[4]&~m[106]&m[107]&~m[108]&m[109])|(~m[4]&~m[106]&~m[107]&m[108]&m[109]))&BiasedRNG[108])|(((m[4]&m[106]&m[107]&~m[108]&~m[109])|(m[4]&m[106]&~m[107]&m[108]&~m[109])|(m[4]&~m[106]&m[107]&m[108]&~m[109])|(~m[4]&m[106]&m[107]&m[108]&~m[109])|(m[4]&m[106]&~m[107]&~m[108]&m[109])|(m[4]&~m[106]&m[107]&~m[108]&m[109])|(~m[4]&m[106]&m[107]&~m[108]&m[109])|(m[4]&~m[106]&~m[107]&m[108]&m[109])|(~m[4]&m[106]&~m[107]&m[108]&m[109])|(~m[4]&~m[106]&m[107]&m[108]&m[109]))&~BiasedRNG[108])|((m[4]&m[106]&m[107]&m[108]&~m[109])|(m[4]&m[106]&m[107]&~m[108]&m[109])|(m[4]&m[106]&~m[107]&m[108]&m[109])|(m[4]&~m[106]&m[107]&m[108]&m[109])|(~m[4]&m[106]&m[107]&m[108]&m[109])|(m[4]&m[106]&m[107]&m[108]&m[109]));
    m[30] = (((m[5]&m[112]&~m[113]&~m[114]&~m[115])|(m[5]&~m[112]&m[113]&~m[114]&~m[115])|(~m[5]&m[112]&m[113]&~m[114]&~m[115])|(m[5]&~m[112]&~m[113]&m[114]&~m[115])|(~m[5]&m[112]&~m[113]&m[114]&~m[115])|(~m[5]&~m[112]&m[113]&m[114]&~m[115])|(m[5]&~m[112]&~m[113]&~m[114]&m[115])|(~m[5]&m[112]&~m[113]&~m[114]&m[115])|(~m[5]&~m[112]&m[113]&~m[114]&m[115])|(~m[5]&~m[112]&~m[113]&m[114]&m[115]))&BiasedRNG[109])|(((m[5]&m[112]&m[113]&~m[114]&~m[115])|(m[5]&m[112]&~m[113]&m[114]&~m[115])|(m[5]&~m[112]&m[113]&m[114]&~m[115])|(~m[5]&m[112]&m[113]&m[114]&~m[115])|(m[5]&m[112]&~m[113]&~m[114]&m[115])|(m[5]&~m[112]&m[113]&~m[114]&m[115])|(~m[5]&m[112]&m[113]&~m[114]&m[115])|(m[5]&~m[112]&~m[113]&m[114]&m[115])|(~m[5]&m[112]&~m[113]&m[114]&m[115])|(~m[5]&~m[112]&m[113]&m[114]&m[115]))&~BiasedRNG[109])|((m[5]&m[112]&m[113]&m[114]&~m[115])|(m[5]&m[112]&m[113]&~m[114]&m[115])|(m[5]&m[112]&~m[113]&m[114]&m[115])|(m[5]&~m[112]&m[113]&m[114]&m[115])|(~m[5]&m[112]&m[113]&m[114]&m[115])|(m[5]&m[112]&m[113]&m[114]&m[115]));
    m[31] = (((m[5]&m[116]&~m[117]&~m[118]&~m[119])|(m[5]&~m[116]&m[117]&~m[118]&~m[119])|(~m[5]&m[116]&m[117]&~m[118]&~m[119])|(m[5]&~m[116]&~m[117]&m[118]&~m[119])|(~m[5]&m[116]&~m[117]&m[118]&~m[119])|(~m[5]&~m[116]&m[117]&m[118]&~m[119])|(m[5]&~m[116]&~m[117]&~m[118]&m[119])|(~m[5]&m[116]&~m[117]&~m[118]&m[119])|(~m[5]&~m[116]&m[117]&~m[118]&m[119])|(~m[5]&~m[116]&~m[117]&m[118]&m[119]))&BiasedRNG[110])|(((m[5]&m[116]&m[117]&~m[118]&~m[119])|(m[5]&m[116]&~m[117]&m[118]&~m[119])|(m[5]&~m[116]&m[117]&m[118]&~m[119])|(~m[5]&m[116]&m[117]&m[118]&~m[119])|(m[5]&m[116]&~m[117]&~m[118]&m[119])|(m[5]&~m[116]&m[117]&~m[118]&m[119])|(~m[5]&m[116]&m[117]&~m[118]&m[119])|(m[5]&~m[116]&~m[117]&m[118]&m[119])|(~m[5]&m[116]&~m[117]&m[118]&m[119])|(~m[5]&~m[116]&m[117]&m[118]&m[119]))&~BiasedRNG[110])|((m[5]&m[116]&m[117]&m[118]&~m[119])|(m[5]&m[116]&m[117]&~m[118]&m[119])|(m[5]&m[116]&~m[117]&m[118]&m[119])|(m[5]&~m[116]&m[117]&m[118]&m[119])|(~m[5]&m[116]&m[117]&m[118]&m[119])|(m[5]&m[116]&m[117]&m[118]&m[119]));
    m[32] = (((m[6]&m[122]&~m[123]&~m[124]&~m[125])|(m[6]&~m[122]&m[123]&~m[124]&~m[125])|(~m[6]&m[122]&m[123]&~m[124]&~m[125])|(m[6]&~m[122]&~m[123]&m[124]&~m[125])|(~m[6]&m[122]&~m[123]&m[124]&~m[125])|(~m[6]&~m[122]&m[123]&m[124]&~m[125])|(m[6]&~m[122]&~m[123]&~m[124]&m[125])|(~m[6]&m[122]&~m[123]&~m[124]&m[125])|(~m[6]&~m[122]&m[123]&~m[124]&m[125])|(~m[6]&~m[122]&~m[123]&m[124]&m[125]))&BiasedRNG[111])|(((m[6]&m[122]&m[123]&~m[124]&~m[125])|(m[6]&m[122]&~m[123]&m[124]&~m[125])|(m[6]&~m[122]&m[123]&m[124]&~m[125])|(~m[6]&m[122]&m[123]&m[124]&~m[125])|(m[6]&m[122]&~m[123]&~m[124]&m[125])|(m[6]&~m[122]&m[123]&~m[124]&m[125])|(~m[6]&m[122]&m[123]&~m[124]&m[125])|(m[6]&~m[122]&~m[123]&m[124]&m[125])|(~m[6]&m[122]&~m[123]&m[124]&m[125])|(~m[6]&~m[122]&m[123]&m[124]&m[125]))&~BiasedRNG[111])|((m[6]&m[122]&m[123]&m[124]&~m[125])|(m[6]&m[122]&m[123]&~m[124]&m[125])|(m[6]&m[122]&~m[123]&m[124]&m[125])|(m[6]&~m[122]&m[123]&m[124]&m[125])|(~m[6]&m[122]&m[123]&m[124]&m[125])|(m[6]&m[122]&m[123]&m[124]&m[125]));
    m[33] = (((m[6]&m[126]&~m[127]&~m[128]&~m[129])|(m[6]&~m[126]&m[127]&~m[128]&~m[129])|(~m[6]&m[126]&m[127]&~m[128]&~m[129])|(m[6]&~m[126]&~m[127]&m[128]&~m[129])|(~m[6]&m[126]&~m[127]&m[128]&~m[129])|(~m[6]&~m[126]&m[127]&m[128]&~m[129])|(m[6]&~m[126]&~m[127]&~m[128]&m[129])|(~m[6]&m[126]&~m[127]&~m[128]&m[129])|(~m[6]&~m[126]&m[127]&~m[128]&m[129])|(~m[6]&~m[126]&~m[127]&m[128]&m[129]))&BiasedRNG[112])|(((m[6]&m[126]&m[127]&~m[128]&~m[129])|(m[6]&m[126]&~m[127]&m[128]&~m[129])|(m[6]&~m[126]&m[127]&m[128]&~m[129])|(~m[6]&m[126]&m[127]&m[128]&~m[129])|(m[6]&m[126]&~m[127]&~m[128]&m[129])|(m[6]&~m[126]&m[127]&~m[128]&m[129])|(~m[6]&m[126]&m[127]&~m[128]&m[129])|(m[6]&~m[126]&~m[127]&m[128]&m[129])|(~m[6]&m[126]&~m[127]&m[128]&m[129])|(~m[6]&~m[126]&m[127]&m[128]&m[129]))&~BiasedRNG[112])|((m[6]&m[126]&m[127]&m[128]&~m[129])|(m[6]&m[126]&m[127]&~m[128]&m[129])|(m[6]&m[126]&~m[127]&m[128]&m[129])|(m[6]&~m[126]&m[127]&m[128]&m[129])|(~m[6]&m[126]&m[127]&m[128]&m[129])|(m[6]&m[126]&m[127]&m[128]&m[129]));
    m[34] = (((m[7]&m[132]&~m[133]&~m[134]&~m[135])|(m[7]&~m[132]&m[133]&~m[134]&~m[135])|(~m[7]&m[132]&m[133]&~m[134]&~m[135])|(m[7]&~m[132]&~m[133]&m[134]&~m[135])|(~m[7]&m[132]&~m[133]&m[134]&~m[135])|(~m[7]&~m[132]&m[133]&m[134]&~m[135])|(m[7]&~m[132]&~m[133]&~m[134]&m[135])|(~m[7]&m[132]&~m[133]&~m[134]&m[135])|(~m[7]&~m[132]&m[133]&~m[134]&m[135])|(~m[7]&~m[132]&~m[133]&m[134]&m[135]))&BiasedRNG[113])|(((m[7]&m[132]&m[133]&~m[134]&~m[135])|(m[7]&m[132]&~m[133]&m[134]&~m[135])|(m[7]&~m[132]&m[133]&m[134]&~m[135])|(~m[7]&m[132]&m[133]&m[134]&~m[135])|(m[7]&m[132]&~m[133]&~m[134]&m[135])|(m[7]&~m[132]&m[133]&~m[134]&m[135])|(~m[7]&m[132]&m[133]&~m[134]&m[135])|(m[7]&~m[132]&~m[133]&m[134]&m[135])|(~m[7]&m[132]&~m[133]&m[134]&m[135])|(~m[7]&~m[132]&m[133]&m[134]&m[135]))&~BiasedRNG[113])|((m[7]&m[132]&m[133]&m[134]&~m[135])|(m[7]&m[132]&m[133]&~m[134]&m[135])|(m[7]&m[132]&~m[133]&m[134]&m[135])|(m[7]&~m[132]&m[133]&m[134]&m[135])|(~m[7]&m[132]&m[133]&m[134]&m[135])|(m[7]&m[132]&m[133]&m[134]&m[135]));
    m[35] = (((m[7]&m[136]&~m[137]&~m[138]&~m[139])|(m[7]&~m[136]&m[137]&~m[138]&~m[139])|(~m[7]&m[136]&m[137]&~m[138]&~m[139])|(m[7]&~m[136]&~m[137]&m[138]&~m[139])|(~m[7]&m[136]&~m[137]&m[138]&~m[139])|(~m[7]&~m[136]&m[137]&m[138]&~m[139])|(m[7]&~m[136]&~m[137]&~m[138]&m[139])|(~m[7]&m[136]&~m[137]&~m[138]&m[139])|(~m[7]&~m[136]&m[137]&~m[138]&m[139])|(~m[7]&~m[136]&~m[137]&m[138]&m[139]))&BiasedRNG[114])|(((m[7]&m[136]&m[137]&~m[138]&~m[139])|(m[7]&m[136]&~m[137]&m[138]&~m[139])|(m[7]&~m[136]&m[137]&m[138]&~m[139])|(~m[7]&m[136]&m[137]&m[138]&~m[139])|(m[7]&m[136]&~m[137]&~m[138]&m[139])|(m[7]&~m[136]&m[137]&~m[138]&m[139])|(~m[7]&m[136]&m[137]&~m[138]&m[139])|(m[7]&~m[136]&~m[137]&m[138]&m[139])|(~m[7]&m[136]&~m[137]&m[138]&m[139])|(~m[7]&~m[136]&m[137]&m[138]&m[139]))&~BiasedRNG[114])|((m[7]&m[136]&m[137]&m[138]&~m[139])|(m[7]&m[136]&m[137]&~m[138]&m[139])|(m[7]&m[136]&~m[137]&m[138]&m[139])|(m[7]&~m[136]&m[137]&m[138]&m[139])|(~m[7]&m[136]&m[137]&m[138]&m[139])|(m[7]&m[136]&m[137]&m[138]&m[139]));
    m[36] = (((m[8]&m[142]&~m[143]&~m[144]&~m[145])|(m[8]&~m[142]&m[143]&~m[144]&~m[145])|(~m[8]&m[142]&m[143]&~m[144]&~m[145])|(m[8]&~m[142]&~m[143]&m[144]&~m[145])|(~m[8]&m[142]&~m[143]&m[144]&~m[145])|(~m[8]&~m[142]&m[143]&m[144]&~m[145])|(m[8]&~m[142]&~m[143]&~m[144]&m[145])|(~m[8]&m[142]&~m[143]&~m[144]&m[145])|(~m[8]&~m[142]&m[143]&~m[144]&m[145])|(~m[8]&~m[142]&~m[143]&m[144]&m[145]))&BiasedRNG[115])|(((m[8]&m[142]&m[143]&~m[144]&~m[145])|(m[8]&m[142]&~m[143]&m[144]&~m[145])|(m[8]&~m[142]&m[143]&m[144]&~m[145])|(~m[8]&m[142]&m[143]&m[144]&~m[145])|(m[8]&m[142]&~m[143]&~m[144]&m[145])|(m[8]&~m[142]&m[143]&~m[144]&m[145])|(~m[8]&m[142]&m[143]&~m[144]&m[145])|(m[8]&~m[142]&~m[143]&m[144]&m[145])|(~m[8]&m[142]&~m[143]&m[144]&m[145])|(~m[8]&~m[142]&m[143]&m[144]&m[145]))&~BiasedRNG[115])|((m[8]&m[142]&m[143]&m[144]&~m[145])|(m[8]&m[142]&m[143]&~m[144]&m[145])|(m[8]&m[142]&~m[143]&m[144]&m[145])|(m[8]&~m[142]&m[143]&m[144]&m[145])|(~m[8]&m[142]&m[143]&m[144]&m[145])|(m[8]&m[142]&m[143]&m[144]&m[145]));
    m[37] = (((m[8]&m[146]&~m[147]&~m[148]&~m[149])|(m[8]&~m[146]&m[147]&~m[148]&~m[149])|(~m[8]&m[146]&m[147]&~m[148]&~m[149])|(m[8]&~m[146]&~m[147]&m[148]&~m[149])|(~m[8]&m[146]&~m[147]&m[148]&~m[149])|(~m[8]&~m[146]&m[147]&m[148]&~m[149])|(m[8]&~m[146]&~m[147]&~m[148]&m[149])|(~m[8]&m[146]&~m[147]&~m[148]&m[149])|(~m[8]&~m[146]&m[147]&~m[148]&m[149])|(~m[8]&~m[146]&~m[147]&m[148]&m[149]))&BiasedRNG[116])|(((m[8]&m[146]&m[147]&~m[148]&~m[149])|(m[8]&m[146]&~m[147]&m[148]&~m[149])|(m[8]&~m[146]&m[147]&m[148]&~m[149])|(~m[8]&m[146]&m[147]&m[148]&~m[149])|(m[8]&m[146]&~m[147]&~m[148]&m[149])|(m[8]&~m[146]&m[147]&~m[148]&m[149])|(~m[8]&m[146]&m[147]&~m[148]&m[149])|(m[8]&~m[146]&~m[147]&m[148]&m[149])|(~m[8]&m[146]&~m[147]&m[148]&m[149])|(~m[8]&~m[146]&m[147]&m[148]&m[149]))&~BiasedRNG[116])|((m[8]&m[146]&m[147]&m[148]&~m[149])|(m[8]&m[146]&m[147]&~m[148]&m[149])|(m[8]&m[146]&~m[147]&m[148]&m[149])|(m[8]&~m[146]&m[147]&m[148]&m[149])|(~m[8]&m[146]&m[147]&m[148]&m[149])|(m[8]&m[146]&m[147]&m[148]&m[149]));
    m[38] = (((m[9]&m[152]&~m[153]&~m[154]&~m[155])|(m[9]&~m[152]&m[153]&~m[154]&~m[155])|(~m[9]&m[152]&m[153]&~m[154]&~m[155])|(m[9]&~m[152]&~m[153]&m[154]&~m[155])|(~m[9]&m[152]&~m[153]&m[154]&~m[155])|(~m[9]&~m[152]&m[153]&m[154]&~m[155])|(m[9]&~m[152]&~m[153]&~m[154]&m[155])|(~m[9]&m[152]&~m[153]&~m[154]&m[155])|(~m[9]&~m[152]&m[153]&~m[154]&m[155])|(~m[9]&~m[152]&~m[153]&m[154]&m[155]))&BiasedRNG[117])|(((m[9]&m[152]&m[153]&~m[154]&~m[155])|(m[9]&m[152]&~m[153]&m[154]&~m[155])|(m[9]&~m[152]&m[153]&m[154]&~m[155])|(~m[9]&m[152]&m[153]&m[154]&~m[155])|(m[9]&m[152]&~m[153]&~m[154]&m[155])|(m[9]&~m[152]&m[153]&~m[154]&m[155])|(~m[9]&m[152]&m[153]&~m[154]&m[155])|(m[9]&~m[152]&~m[153]&m[154]&m[155])|(~m[9]&m[152]&~m[153]&m[154]&m[155])|(~m[9]&~m[152]&m[153]&m[154]&m[155]))&~BiasedRNG[117])|((m[9]&m[152]&m[153]&m[154]&~m[155])|(m[9]&m[152]&m[153]&~m[154]&m[155])|(m[9]&m[152]&~m[153]&m[154]&m[155])|(m[9]&~m[152]&m[153]&m[154]&m[155])|(~m[9]&m[152]&m[153]&m[154]&m[155])|(m[9]&m[152]&m[153]&m[154]&m[155]));
    m[39] = (((m[9]&m[156]&~m[157]&~m[158]&~m[159])|(m[9]&~m[156]&m[157]&~m[158]&~m[159])|(~m[9]&m[156]&m[157]&~m[158]&~m[159])|(m[9]&~m[156]&~m[157]&m[158]&~m[159])|(~m[9]&m[156]&~m[157]&m[158]&~m[159])|(~m[9]&~m[156]&m[157]&m[158]&~m[159])|(m[9]&~m[156]&~m[157]&~m[158]&m[159])|(~m[9]&m[156]&~m[157]&~m[158]&m[159])|(~m[9]&~m[156]&m[157]&~m[158]&m[159])|(~m[9]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[118])|(((m[9]&m[156]&m[157]&~m[158]&~m[159])|(m[9]&m[156]&~m[157]&m[158]&~m[159])|(m[9]&~m[156]&m[157]&m[158]&~m[159])|(~m[9]&m[156]&m[157]&m[158]&~m[159])|(m[9]&m[156]&~m[157]&~m[158]&m[159])|(m[9]&~m[156]&m[157]&~m[158]&m[159])|(~m[9]&m[156]&m[157]&~m[158]&m[159])|(m[9]&~m[156]&~m[157]&m[158]&m[159])|(~m[9]&m[156]&~m[157]&m[158]&m[159])|(~m[9]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[118])|((m[9]&m[156]&m[157]&m[158]&~m[159])|(m[9]&m[156]&m[157]&~m[158]&m[159])|(m[9]&m[156]&~m[157]&m[158]&m[159])|(m[9]&~m[156]&m[157]&m[158]&m[159])|(~m[9]&m[156]&m[157]&m[158]&m[159])|(m[9]&m[156]&m[157]&m[158]&m[159]));
    m[40] = (((m[10]&m[162]&~m[163]&~m[164]&~m[165])|(m[10]&~m[162]&m[163]&~m[164]&~m[165])|(~m[10]&m[162]&m[163]&~m[164]&~m[165])|(m[10]&~m[162]&~m[163]&m[164]&~m[165])|(~m[10]&m[162]&~m[163]&m[164]&~m[165])|(~m[10]&~m[162]&m[163]&m[164]&~m[165])|(m[10]&~m[162]&~m[163]&~m[164]&m[165])|(~m[10]&m[162]&~m[163]&~m[164]&m[165])|(~m[10]&~m[162]&m[163]&~m[164]&m[165])|(~m[10]&~m[162]&~m[163]&m[164]&m[165]))&BiasedRNG[119])|(((m[10]&m[162]&m[163]&~m[164]&~m[165])|(m[10]&m[162]&~m[163]&m[164]&~m[165])|(m[10]&~m[162]&m[163]&m[164]&~m[165])|(~m[10]&m[162]&m[163]&m[164]&~m[165])|(m[10]&m[162]&~m[163]&~m[164]&m[165])|(m[10]&~m[162]&m[163]&~m[164]&m[165])|(~m[10]&m[162]&m[163]&~m[164]&m[165])|(m[10]&~m[162]&~m[163]&m[164]&m[165])|(~m[10]&m[162]&~m[163]&m[164]&m[165])|(~m[10]&~m[162]&m[163]&m[164]&m[165]))&~BiasedRNG[119])|((m[10]&m[162]&m[163]&m[164]&~m[165])|(m[10]&m[162]&m[163]&~m[164]&m[165])|(m[10]&m[162]&~m[163]&m[164]&m[165])|(m[10]&~m[162]&m[163]&m[164]&m[165])|(~m[10]&m[162]&m[163]&m[164]&m[165])|(m[10]&m[162]&m[163]&m[164]&m[165]));
    m[41] = (((m[10]&m[166]&~m[167]&~m[168]&~m[169])|(m[10]&~m[166]&m[167]&~m[168]&~m[169])|(~m[10]&m[166]&m[167]&~m[168]&~m[169])|(m[10]&~m[166]&~m[167]&m[168]&~m[169])|(~m[10]&m[166]&~m[167]&m[168]&~m[169])|(~m[10]&~m[166]&m[167]&m[168]&~m[169])|(m[10]&~m[166]&~m[167]&~m[168]&m[169])|(~m[10]&m[166]&~m[167]&~m[168]&m[169])|(~m[10]&~m[166]&m[167]&~m[168]&m[169])|(~m[10]&~m[166]&~m[167]&m[168]&m[169]))&BiasedRNG[120])|(((m[10]&m[166]&m[167]&~m[168]&~m[169])|(m[10]&m[166]&~m[167]&m[168]&~m[169])|(m[10]&~m[166]&m[167]&m[168]&~m[169])|(~m[10]&m[166]&m[167]&m[168]&~m[169])|(m[10]&m[166]&~m[167]&~m[168]&m[169])|(m[10]&~m[166]&m[167]&~m[168]&m[169])|(~m[10]&m[166]&m[167]&~m[168]&m[169])|(m[10]&~m[166]&~m[167]&m[168]&m[169])|(~m[10]&m[166]&~m[167]&m[168]&m[169])|(~m[10]&~m[166]&m[167]&m[168]&m[169]))&~BiasedRNG[120])|((m[10]&m[166]&m[167]&m[168]&~m[169])|(m[10]&m[166]&m[167]&~m[168]&m[169])|(m[10]&m[166]&~m[167]&m[168]&m[169])|(m[10]&~m[166]&m[167]&m[168]&m[169])|(~m[10]&m[166]&m[167]&m[168]&m[169])|(m[10]&m[166]&m[167]&m[168]&m[169]));
    m[42] = (((m[11]&m[172]&~m[173]&~m[174]&~m[175])|(m[11]&~m[172]&m[173]&~m[174]&~m[175])|(~m[11]&m[172]&m[173]&~m[174]&~m[175])|(m[11]&~m[172]&~m[173]&m[174]&~m[175])|(~m[11]&m[172]&~m[173]&m[174]&~m[175])|(~m[11]&~m[172]&m[173]&m[174]&~m[175])|(m[11]&~m[172]&~m[173]&~m[174]&m[175])|(~m[11]&m[172]&~m[173]&~m[174]&m[175])|(~m[11]&~m[172]&m[173]&~m[174]&m[175])|(~m[11]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[121])|(((m[11]&m[172]&m[173]&~m[174]&~m[175])|(m[11]&m[172]&~m[173]&m[174]&~m[175])|(m[11]&~m[172]&m[173]&m[174]&~m[175])|(~m[11]&m[172]&m[173]&m[174]&~m[175])|(m[11]&m[172]&~m[173]&~m[174]&m[175])|(m[11]&~m[172]&m[173]&~m[174]&m[175])|(~m[11]&m[172]&m[173]&~m[174]&m[175])|(m[11]&~m[172]&~m[173]&m[174]&m[175])|(~m[11]&m[172]&~m[173]&m[174]&m[175])|(~m[11]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[121])|((m[11]&m[172]&m[173]&m[174]&~m[175])|(m[11]&m[172]&m[173]&~m[174]&m[175])|(m[11]&m[172]&~m[173]&m[174]&m[175])|(m[11]&~m[172]&m[173]&m[174]&m[175])|(~m[11]&m[172]&m[173]&m[174]&m[175])|(m[11]&m[172]&m[173]&m[174]&m[175]));
    m[43] = (((m[11]&m[176]&~m[177]&~m[178]&~m[179])|(m[11]&~m[176]&m[177]&~m[178]&~m[179])|(~m[11]&m[176]&m[177]&~m[178]&~m[179])|(m[11]&~m[176]&~m[177]&m[178]&~m[179])|(~m[11]&m[176]&~m[177]&m[178]&~m[179])|(~m[11]&~m[176]&m[177]&m[178]&~m[179])|(m[11]&~m[176]&~m[177]&~m[178]&m[179])|(~m[11]&m[176]&~m[177]&~m[178]&m[179])|(~m[11]&~m[176]&m[177]&~m[178]&m[179])|(~m[11]&~m[176]&~m[177]&m[178]&m[179]))&BiasedRNG[122])|(((m[11]&m[176]&m[177]&~m[178]&~m[179])|(m[11]&m[176]&~m[177]&m[178]&~m[179])|(m[11]&~m[176]&m[177]&m[178]&~m[179])|(~m[11]&m[176]&m[177]&m[178]&~m[179])|(m[11]&m[176]&~m[177]&~m[178]&m[179])|(m[11]&~m[176]&m[177]&~m[178]&m[179])|(~m[11]&m[176]&m[177]&~m[178]&m[179])|(m[11]&~m[176]&~m[177]&m[178]&m[179])|(~m[11]&m[176]&~m[177]&m[178]&m[179])|(~m[11]&~m[176]&m[177]&m[178]&m[179]))&~BiasedRNG[122])|((m[11]&m[176]&m[177]&m[178]&~m[179])|(m[11]&m[176]&m[177]&~m[178]&m[179])|(m[11]&m[176]&~m[177]&m[178]&m[179])|(m[11]&~m[176]&m[177]&m[178]&m[179])|(~m[11]&m[176]&m[177]&m[178]&m[179])|(m[11]&m[176]&m[177]&m[178]&m[179]));
    m[44] = (((m[12]&m[182]&~m[183]&~m[184]&~m[185])|(m[12]&~m[182]&m[183]&~m[184]&~m[185])|(~m[12]&m[182]&m[183]&~m[184]&~m[185])|(m[12]&~m[182]&~m[183]&m[184]&~m[185])|(~m[12]&m[182]&~m[183]&m[184]&~m[185])|(~m[12]&~m[182]&m[183]&m[184]&~m[185])|(m[12]&~m[182]&~m[183]&~m[184]&m[185])|(~m[12]&m[182]&~m[183]&~m[184]&m[185])|(~m[12]&~m[182]&m[183]&~m[184]&m[185])|(~m[12]&~m[182]&~m[183]&m[184]&m[185]))&BiasedRNG[123])|(((m[12]&m[182]&m[183]&~m[184]&~m[185])|(m[12]&m[182]&~m[183]&m[184]&~m[185])|(m[12]&~m[182]&m[183]&m[184]&~m[185])|(~m[12]&m[182]&m[183]&m[184]&~m[185])|(m[12]&m[182]&~m[183]&~m[184]&m[185])|(m[12]&~m[182]&m[183]&~m[184]&m[185])|(~m[12]&m[182]&m[183]&~m[184]&m[185])|(m[12]&~m[182]&~m[183]&m[184]&m[185])|(~m[12]&m[182]&~m[183]&m[184]&m[185])|(~m[12]&~m[182]&m[183]&m[184]&m[185]))&~BiasedRNG[123])|((m[12]&m[182]&m[183]&m[184]&~m[185])|(m[12]&m[182]&m[183]&~m[184]&m[185])|(m[12]&m[182]&~m[183]&m[184]&m[185])|(m[12]&~m[182]&m[183]&m[184]&m[185])|(~m[12]&m[182]&m[183]&m[184]&m[185])|(m[12]&m[182]&m[183]&m[184]&m[185]));
    m[45] = (((m[12]&m[186]&~m[187]&~m[188]&~m[189])|(m[12]&~m[186]&m[187]&~m[188]&~m[189])|(~m[12]&m[186]&m[187]&~m[188]&~m[189])|(m[12]&~m[186]&~m[187]&m[188]&~m[189])|(~m[12]&m[186]&~m[187]&m[188]&~m[189])|(~m[12]&~m[186]&m[187]&m[188]&~m[189])|(m[12]&~m[186]&~m[187]&~m[188]&m[189])|(~m[12]&m[186]&~m[187]&~m[188]&m[189])|(~m[12]&~m[186]&m[187]&~m[188]&m[189])|(~m[12]&~m[186]&~m[187]&m[188]&m[189]))&BiasedRNG[124])|(((m[12]&m[186]&m[187]&~m[188]&~m[189])|(m[12]&m[186]&~m[187]&m[188]&~m[189])|(m[12]&~m[186]&m[187]&m[188]&~m[189])|(~m[12]&m[186]&m[187]&m[188]&~m[189])|(m[12]&m[186]&~m[187]&~m[188]&m[189])|(m[12]&~m[186]&m[187]&~m[188]&m[189])|(~m[12]&m[186]&m[187]&~m[188]&m[189])|(m[12]&~m[186]&~m[187]&m[188]&m[189])|(~m[12]&m[186]&~m[187]&m[188]&m[189])|(~m[12]&~m[186]&m[187]&m[188]&m[189]))&~BiasedRNG[124])|((m[12]&m[186]&m[187]&m[188]&~m[189])|(m[12]&m[186]&m[187]&~m[188]&m[189])|(m[12]&m[186]&~m[187]&m[188]&m[189])|(m[12]&~m[186]&m[187]&m[188]&m[189])|(~m[12]&m[186]&m[187]&m[188]&m[189])|(m[12]&m[186]&m[187]&m[188]&m[189]));
    m[46] = (((m[13]&m[192]&~m[193]&~m[194]&~m[195])|(m[13]&~m[192]&m[193]&~m[194]&~m[195])|(~m[13]&m[192]&m[193]&~m[194]&~m[195])|(m[13]&~m[192]&~m[193]&m[194]&~m[195])|(~m[13]&m[192]&~m[193]&m[194]&~m[195])|(~m[13]&~m[192]&m[193]&m[194]&~m[195])|(m[13]&~m[192]&~m[193]&~m[194]&m[195])|(~m[13]&m[192]&~m[193]&~m[194]&m[195])|(~m[13]&~m[192]&m[193]&~m[194]&m[195])|(~m[13]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[125])|(((m[13]&m[192]&m[193]&~m[194]&~m[195])|(m[13]&m[192]&~m[193]&m[194]&~m[195])|(m[13]&~m[192]&m[193]&m[194]&~m[195])|(~m[13]&m[192]&m[193]&m[194]&~m[195])|(m[13]&m[192]&~m[193]&~m[194]&m[195])|(m[13]&~m[192]&m[193]&~m[194]&m[195])|(~m[13]&m[192]&m[193]&~m[194]&m[195])|(m[13]&~m[192]&~m[193]&m[194]&m[195])|(~m[13]&m[192]&~m[193]&m[194]&m[195])|(~m[13]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[125])|((m[13]&m[192]&m[193]&m[194]&~m[195])|(m[13]&m[192]&m[193]&~m[194]&m[195])|(m[13]&m[192]&~m[193]&m[194]&m[195])|(m[13]&~m[192]&m[193]&m[194]&m[195])|(~m[13]&m[192]&m[193]&m[194]&m[195])|(m[13]&m[192]&m[193]&m[194]&m[195]));
    m[47] = (((m[13]&m[196]&~m[197]&~m[198]&~m[199])|(m[13]&~m[196]&m[197]&~m[198]&~m[199])|(~m[13]&m[196]&m[197]&~m[198]&~m[199])|(m[13]&~m[196]&~m[197]&m[198]&~m[199])|(~m[13]&m[196]&~m[197]&m[198]&~m[199])|(~m[13]&~m[196]&m[197]&m[198]&~m[199])|(m[13]&~m[196]&~m[197]&~m[198]&m[199])|(~m[13]&m[196]&~m[197]&~m[198]&m[199])|(~m[13]&~m[196]&m[197]&~m[198]&m[199])|(~m[13]&~m[196]&~m[197]&m[198]&m[199]))&BiasedRNG[126])|(((m[13]&m[196]&m[197]&~m[198]&~m[199])|(m[13]&m[196]&~m[197]&m[198]&~m[199])|(m[13]&~m[196]&m[197]&m[198]&~m[199])|(~m[13]&m[196]&m[197]&m[198]&~m[199])|(m[13]&m[196]&~m[197]&~m[198]&m[199])|(m[13]&~m[196]&m[197]&~m[198]&m[199])|(~m[13]&m[196]&m[197]&~m[198]&m[199])|(m[13]&~m[196]&~m[197]&m[198]&m[199])|(~m[13]&m[196]&~m[197]&m[198]&m[199])|(~m[13]&~m[196]&m[197]&m[198]&m[199]))&~BiasedRNG[126])|((m[13]&m[196]&m[197]&m[198]&~m[199])|(m[13]&m[196]&m[197]&~m[198]&m[199])|(m[13]&m[196]&~m[197]&m[198]&m[199])|(m[13]&~m[196]&m[197]&m[198]&m[199])|(~m[13]&m[196]&m[197]&m[198]&m[199])|(m[13]&m[196]&m[197]&m[198]&m[199]));
    m[48] = (((m[14]&m[202]&~m[203]&~m[204]&~m[205])|(m[14]&~m[202]&m[203]&~m[204]&~m[205])|(~m[14]&m[202]&m[203]&~m[204]&~m[205])|(m[14]&~m[202]&~m[203]&m[204]&~m[205])|(~m[14]&m[202]&~m[203]&m[204]&~m[205])|(~m[14]&~m[202]&m[203]&m[204]&~m[205])|(m[14]&~m[202]&~m[203]&~m[204]&m[205])|(~m[14]&m[202]&~m[203]&~m[204]&m[205])|(~m[14]&~m[202]&m[203]&~m[204]&m[205])|(~m[14]&~m[202]&~m[203]&m[204]&m[205]))&BiasedRNG[127])|(((m[14]&m[202]&m[203]&~m[204]&~m[205])|(m[14]&m[202]&~m[203]&m[204]&~m[205])|(m[14]&~m[202]&m[203]&m[204]&~m[205])|(~m[14]&m[202]&m[203]&m[204]&~m[205])|(m[14]&m[202]&~m[203]&~m[204]&m[205])|(m[14]&~m[202]&m[203]&~m[204]&m[205])|(~m[14]&m[202]&m[203]&~m[204]&m[205])|(m[14]&~m[202]&~m[203]&m[204]&m[205])|(~m[14]&m[202]&~m[203]&m[204]&m[205])|(~m[14]&~m[202]&m[203]&m[204]&m[205]))&~BiasedRNG[127])|((m[14]&m[202]&m[203]&m[204]&~m[205])|(m[14]&m[202]&m[203]&~m[204]&m[205])|(m[14]&m[202]&~m[203]&m[204]&m[205])|(m[14]&~m[202]&m[203]&m[204]&m[205])|(~m[14]&m[202]&m[203]&m[204]&m[205])|(m[14]&m[202]&m[203]&m[204]&m[205]));
    m[49] = (((m[14]&m[206]&~m[207]&~m[208]&~m[209])|(m[14]&~m[206]&m[207]&~m[208]&~m[209])|(~m[14]&m[206]&m[207]&~m[208]&~m[209])|(m[14]&~m[206]&~m[207]&m[208]&~m[209])|(~m[14]&m[206]&~m[207]&m[208]&~m[209])|(~m[14]&~m[206]&m[207]&m[208]&~m[209])|(m[14]&~m[206]&~m[207]&~m[208]&m[209])|(~m[14]&m[206]&~m[207]&~m[208]&m[209])|(~m[14]&~m[206]&m[207]&~m[208]&m[209])|(~m[14]&~m[206]&~m[207]&m[208]&m[209]))&BiasedRNG[128])|(((m[14]&m[206]&m[207]&~m[208]&~m[209])|(m[14]&m[206]&~m[207]&m[208]&~m[209])|(m[14]&~m[206]&m[207]&m[208]&~m[209])|(~m[14]&m[206]&m[207]&m[208]&~m[209])|(m[14]&m[206]&~m[207]&~m[208]&m[209])|(m[14]&~m[206]&m[207]&~m[208]&m[209])|(~m[14]&m[206]&m[207]&~m[208]&m[209])|(m[14]&~m[206]&~m[207]&m[208]&m[209])|(~m[14]&m[206]&~m[207]&m[208]&m[209])|(~m[14]&~m[206]&m[207]&m[208]&m[209]))&~BiasedRNG[128])|((m[14]&m[206]&m[207]&m[208]&~m[209])|(m[14]&m[206]&m[207]&~m[208]&m[209])|(m[14]&m[206]&~m[207]&m[208]&m[209])|(m[14]&~m[206]&m[207]&m[208]&m[209])|(~m[14]&m[206]&m[207]&m[208]&m[209])|(m[14]&m[206]&m[207]&m[208]&m[209]));
    m[50] = (((m[15]&m[212]&~m[213]&~m[214]&~m[215])|(m[15]&~m[212]&m[213]&~m[214]&~m[215])|(~m[15]&m[212]&m[213]&~m[214]&~m[215])|(m[15]&~m[212]&~m[213]&m[214]&~m[215])|(~m[15]&m[212]&~m[213]&m[214]&~m[215])|(~m[15]&~m[212]&m[213]&m[214]&~m[215])|(m[15]&~m[212]&~m[213]&~m[214]&m[215])|(~m[15]&m[212]&~m[213]&~m[214]&m[215])|(~m[15]&~m[212]&m[213]&~m[214]&m[215])|(~m[15]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[129])|(((m[15]&m[212]&m[213]&~m[214]&~m[215])|(m[15]&m[212]&~m[213]&m[214]&~m[215])|(m[15]&~m[212]&m[213]&m[214]&~m[215])|(~m[15]&m[212]&m[213]&m[214]&~m[215])|(m[15]&m[212]&~m[213]&~m[214]&m[215])|(m[15]&~m[212]&m[213]&~m[214]&m[215])|(~m[15]&m[212]&m[213]&~m[214]&m[215])|(m[15]&~m[212]&~m[213]&m[214]&m[215])|(~m[15]&m[212]&~m[213]&m[214]&m[215])|(~m[15]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[129])|((m[15]&m[212]&m[213]&m[214]&~m[215])|(m[15]&m[212]&m[213]&~m[214]&m[215])|(m[15]&m[212]&~m[213]&m[214]&m[215])|(m[15]&~m[212]&m[213]&m[214]&m[215])|(~m[15]&m[212]&m[213]&m[214]&m[215])|(m[15]&m[212]&m[213]&m[214]&m[215]));
    m[51] = (((m[15]&m[216]&~m[217]&~m[218]&~m[219])|(m[15]&~m[216]&m[217]&~m[218]&~m[219])|(~m[15]&m[216]&m[217]&~m[218]&~m[219])|(m[15]&~m[216]&~m[217]&m[218]&~m[219])|(~m[15]&m[216]&~m[217]&m[218]&~m[219])|(~m[15]&~m[216]&m[217]&m[218]&~m[219])|(m[15]&~m[216]&~m[217]&~m[218]&m[219])|(~m[15]&m[216]&~m[217]&~m[218]&m[219])|(~m[15]&~m[216]&m[217]&~m[218]&m[219])|(~m[15]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[130])|(((m[15]&m[216]&m[217]&~m[218]&~m[219])|(m[15]&m[216]&~m[217]&m[218]&~m[219])|(m[15]&~m[216]&m[217]&m[218]&~m[219])|(~m[15]&m[216]&m[217]&m[218]&~m[219])|(m[15]&m[216]&~m[217]&~m[218]&m[219])|(m[15]&~m[216]&m[217]&~m[218]&m[219])|(~m[15]&m[216]&m[217]&~m[218]&m[219])|(m[15]&~m[216]&~m[217]&m[218]&m[219])|(~m[15]&m[216]&~m[217]&m[218]&m[219])|(~m[15]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[130])|((m[15]&m[216]&m[217]&m[218]&~m[219])|(m[15]&m[216]&m[217]&~m[218]&m[219])|(m[15]&m[216]&~m[217]&m[218]&m[219])|(m[15]&~m[216]&m[217]&m[218]&m[219])|(~m[15]&m[216]&m[217]&m[218]&m[219])|(m[15]&m[216]&m[217]&m[218]&m[219]));
    m[52] = (((m[16]&m[222]&~m[223]&~m[224]&~m[225])|(m[16]&~m[222]&m[223]&~m[224]&~m[225])|(~m[16]&m[222]&m[223]&~m[224]&~m[225])|(m[16]&~m[222]&~m[223]&m[224]&~m[225])|(~m[16]&m[222]&~m[223]&m[224]&~m[225])|(~m[16]&~m[222]&m[223]&m[224]&~m[225])|(m[16]&~m[222]&~m[223]&~m[224]&m[225])|(~m[16]&m[222]&~m[223]&~m[224]&m[225])|(~m[16]&~m[222]&m[223]&~m[224]&m[225])|(~m[16]&~m[222]&~m[223]&m[224]&m[225]))&BiasedRNG[131])|(((m[16]&m[222]&m[223]&~m[224]&~m[225])|(m[16]&m[222]&~m[223]&m[224]&~m[225])|(m[16]&~m[222]&m[223]&m[224]&~m[225])|(~m[16]&m[222]&m[223]&m[224]&~m[225])|(m[16]&m[222]&~m[223]&~m[224]&m[225])|(m[16]&~m[222]&m[223]&~m[224]&m[225])|(~m[16]&m[222]&m[223]&~m[224]&m[225])|(m[16]&~m[222]&~m[223]&m[224]&m[225])|(~m[16]&m[222]&~m[223]&m[224]&m[225])|(~m[16]&~m[222]&m[223]&m[224]&m[225]))&~BiasedRNG[131])|((m[16]&m[222]&m[223]&m[224]&~m[225])|(m[16]&m[222]&m[223]&~m[224]&m[225])|(m[16]&m[222]&~m[223]&m[224]&m[225])|(m[16]&~m[222]&m[223]&m[224]&m[225])|(~m[16]&m[222]&m[223]&m[224]&m[225])|(m[16]&m[222]&m[223]&m[224]&m[225]));
    m[53] = (((m[16]&m[226]&~m[227]&~m[228]&~m[229])|(m[16]&~m[226]&m[227]&~m[228]&~m[229])|(~m[16]&m[226]&m[227]&~m[228]&~m[229])|(m[16]&~m[226]&~m[227]&m[228]&~m[229])|(~m[16]&m[226]&~m[227]&m[228]&~m[229])|(~m[16]&~m[226]&m[227]&m[228]&~m[229])|(m[16]&~m[226]&~m[227]&~m[228]&m[229])|(~m[16]&m[226]&~m[227]&~m[228]&m[229])|(~m[16]&~m[226]&m[227]&~m[228]&m[229])|(~m[16]&~m[226]&~m[227]&m[228]&m[229]))&BiasedRNG[132])|(((m[16]&m[226]&m[227]&~m[228]&~m[229])|(m[16]&m[226]&~m[227]&m[228]&~m[229])|(m[16]&~m[226]&m[227]&m[228]&~m[229])|(~m[16]&m[226]&m[227]&m[228]&~m[229])|(m[16]&m[226]&~m[227]&~m[228]&m[229])|(m[16]&~m[226]&m[227]&~m[228]&m[229])|(~m[16]&m[226]&m[227]&~m[228]&m[229])|(m[16]&~m[226]&~m[227]&m[228]&m[229])|(~m[16]&m[226]&~m[227]&m[228]&m[229])|(~m[16]&~m[226]&m[227]&m[228]&m[229]))&~BiasedRNG[132])|((m[16]&m[226]&m[227]&m[228]&~m[229])|(m[16]&m[226]&m[227]&~m[228]&m[229])|(m[16]&m[226]&~m[227]&m[228]&m[229])|(m[16]&~m[226]&m[227]&m[228]&m[229])|(~m[16]&m[226]&m[227]&m[228]&m[229])|(m[16]&m[226]&m[227]&m[228]&m[229]));
    m[54] = (((m[17]&m[232]&~m[233]&~m[234]&~m[235])|(m[17]&~m[232]&m[233]&~m[234]&~m[235])|(~m[17]&m[232]&m[233]&~m[234]&~m[235])|(m[17]&~m[232]&~m[233]&m[234]&~m[235])|(~m[17]&m[232]&~m[233]&m[234]&~m[235])|(~m[17]&~m[232]&m[233]&m[234]&~m[235])|(m[17]&~m[232]&~m[233]&~m[234]&m[235])|(~m[17]&m[232]&~m[233]&~m[234]&m[235])|(~m[17]&~m[232]&m[233]&~m[234]&m[235])|(~m[17]&~m[232]&~m[233]&m[234]&m[235]))&BiasedRNG[133])|(((m[17]&m[232]&m[233]&~m[234]&~m[235])|(m[17]&m[232]&~m[233]&m[234]&~m[235])|(m[17]&~m[232]&m[233]&m[234]&~m[235])|(~m[17]&m[232]&m[233]&m[234]&~m[235])|(m[17]&m[232]&~m[233]&~m[234]&m[235])|(m[17]&~m[232]&m[233]&~m[234]&m[235])|(~m[17]&m[232]&m[233]&~m[234]&m[235])|(m[17]&~m[232]&~m[233]&m[234]&m[235])|(~m[17]&m[232]&~m[233]&m[234]&m[235])|(~m[17]&~m[232]&m[233]&m[234]&m[235]))&~BiasedRNG[133])|((m[17]&m[232]&m[233]&m[234]&~m[235])|(m[17]&m[232]&m[233]&~m[234]&m[235])|(m[17]&m[232]&~m[233]&m[234]&m[235])|(m[17]&~m[232]&m[233]&m[234]&m[235])|(~m[17]&m[232]&m[233]&m[234]&m[235])|(m[17]&m[232]&m[233]&m[234]&m[235]));
    m[55] = (((m[17]&m[236]&~m[237]&~m[238]&~m[239])|(m[17]&~m[236]&m[237]&~m[238]&~m[239])|(~m[17]&m[236]&m[237]&~m[238]&~m[239])|(m[17]&~m[236]&~m[237]&m[238]&~m[239])|(~m[17]&m[236]&~m[237]&m[238]&~m[239])|(~m[17]&~m[236]&m[237]&m[238]&~m[239])|(m[17]&~m[236]&~m[237]&~m[238]&m[239])|(~m[17]&m[236]&~m[237]&~m[238]&m[239])|(~m[17]&~m[236]&m[237]&~m[238]&m[239])|(~m[17]&~m[236]&~m[237]&m[238]&m[239]))&BiasedRNG[134])|(((m[17]&m[236]&m[237]&~m[238]&~m[239])|(m[17]&m[236]&~m[237]&m[238]&~m[239])|(m[17]&~m[236]&m[237]&m[238]&~m[239])|(~m[17]&m[236]&m[237]&m[238]&~m[239])|(m[17]&m[236]&~m[237]&~m[238]&m[239])|(m[17]&~m[236]&m[237]&~m[238]&m[239])|(~m[17]&m[236]&m[237]&~m[238]&m[239])|(m[17]&~m[236]&~m[237]&m[238]&m[239])|(~m[17]&m[236]&~m[237]&m[238]&m[239])|(~m[17]&~m[236]&m[237]&m[238]&m[239]))&~BiasedRNG[134])|((m[17]&m[236]&m[237]&m[238]&~m[239])|(m[17]&m[236]&m[237]&~m[238]&m[239])|(m[17]&m[236]&~m[237]&m[238]&m[239])|(m[17]&~m[236]&m[237]&m[238]&m[239])|(~m[17]&m[236]&m[237]&m[238]&m[239])|(m[17]&m[236]&m[237]&m[238]&m[239]));
    m[56] = (((m[18]&m[242]&~m[243]&~m[244]&~m[245])|(m[18]&~m[242]&m[243]&~m[244]&~m[245])|(~m[18]&m[242]&m[243]&~m[244]&~m[245])|(m[18]&~m[242]&~m[243]&m[244]&~m[245])|(~m[18]&m[242]&~m[243]&m[244]&~m[245])|(~m[18]&~m[242]&m[243]&m[244]&~m[245])|(m[18]&~m[242]&~m[243]&~m[244]&m[245])|(~m[18]&m[242]&~m[243]&~m[244]&m[245])|(~m[18]&~m[242]&m[243]&~m[244]&m[245])|(~m[18]&~m[242]&~m[243]&m[244]&m[245]))&BiasedRNG[135])|(((m[18]&m[242]&m[243]&~m[244]&~m[245])|(m[18]&m[242]&~m[243]&m[244]&~m[245])|(m[18]&~m[242]&m[243]&m[244]&~m[245])|(~m[18]&m[242]&m[243]&m[244]&~m[245])|(m[18]&m[242]&~m[243]&~m[244]&m[245])|(m[18]&~m[242]&m[243]&~m[244]&m[245])|(~m[18]&m[242]&m[243]&~m[244]&m[245])|(m[18]&~m[242]&~m[243]&m[244]&m[245])|(~m[18]&m[242]&~m[243]&m[244]&m[245])|(~m[18]&~m[242]&m[243]&m[244]&m[245]))&~BiasedRNG[135])|((m[18]&m[242]&m[243]&m[244]&~m[245])|(m[18]&m[242]&m[243]&~m[244]&m[245])|(m[18]&m[242]&~m[243]&m[244]&m[245])|(m[18]&~m[242]&m[243]&m[244]&m[245])|(~m[18]&m[242]&m[243]&m[244]&m[245])|(m[18]&m[242]&m[243]&m[244]&m[245]));
    m[57] = (((m[18]&m[246]&~m[247]&~m[248]&~m[249])|(m[18]&~m[246]&m[247]&~m[248]&~m[249])|(~m[18]&m[246]&m[247]&~m[248]&~m[249])|(m[18]&~m[246]&~m[247]&m[248]&~m[249])|(~m[18]&m[246]&~m[247]&m[248]&~m[249])|(~m[18]&~m[246]&m[247]&m[248]&~m[249])|(m[18]&~m[246]&~m[247]&~m[248]&m[249])|(~m[18]&m[246]&~m[247]&~m[248]&m[249])|(~m[18]&~m[246]&m[247]&~m[248]&m[249])|(~m[18]&~m[246]&~m[247]&m[248]&m[249]))&BiasedRNG[136])|(((m[18]&m[246]&m[247]&~m[248]&~m[249])|(m[18]&m[246]&~m[247]&m[248]&~m[249])|(m[18]&~m[246]&m[247]&m[248]&~m[249])|(~m[18]&m[246]&m[247]&m[248]&~m[249])|(m[18]&m[246]&~m[247]&~m[248]&m[249])|(m[18]&~m[246]&m[247]&~m[248]&m[249])|(~m[18]&m[246]&m[247]&~m[248]&m[249])|(m[18]&~m[246]&~m[247]&m[248]&m[249])|(~m[18]&m[246]&~m[247]&m[248]&m[249])|(~m[18]&~m[246]&m[247]&m[248]&m[249]))&~BiasedRNG[136])|((m[18]&m[246]&m[247]&m[248]&~m[249])|(m[18]&m[246]&m[247]&~m[248]&m[249])|(m[18]&m[246]&~m[247]&m[248]&m[249])|(m[18]&~m[246]&m[247]&m[248]&m[249])|(~m[18]&m[246]&m[247]&m[248]&m[249])|(m[18]&m[246]&m[247]&m[248]&m[249]));
    m[58] = (((m[19]&m[252]&~m[253]&~m[254]&~m[255])|(m[19]&~m[252]&m[253]&~m[254]&~m[255])|(~m[19]&m[252]&m[253]&~m[254]&~m[255])|(m[19]&~m[252]&~m[253]&m[254]&~m[255])|(~m[19]&m[252]&~m[253]&m[254]&~m[255])|(~m[19]&~m[252]&m[253]&m[254]&~m[255])|(m[19]&~m[252]&~m[253]&~m[254]&m[255])|(~m[19]&m[252]&~m[253]&~m[254]&m[255])|(~m[19]&~m[252]&m[253]&~m[254]&m[255])|(~m[19]&~m[252]&~m[253]&m[254]&m[255]))&BiasedRNG[137])|(((m[19]&m[252]&m[253]&~m[254]&~m[255])|(m[19]&m[252]&~m[253]&m[254]&~m[255])|(m[19]&~m[252]&m[253]&m[254]&~m[255])|(~m[19]&m[252]&m[253]&m[254]&~m[255])|(m[19]&m[252]&~m[253]&~m[254]&m[255])|(m[19]&~m[252]&m[253]&~m[254]&m[255])|(~m[19]&m[252]&m[253]&~m[254]&m[255])|(m[19]&~m[252]&~m[253]&m[254]&m[255])|(~m[19]&m[252]&~m[253]&m[254]&m[255])|(~m[19]&~m[252]&m[253]&m[254]&m[255]))&~BiasedRNG[137])|((m[19]&m[252]&m[253]&m[254]&~m[255])|(m[19]&m[252]&m[253]&~m[254]&m[255])|(m[19]&m[252]&~m[253]&m[254]&m[255])|(m[19]&~m[252]&m[253]&m[254]&m[255])|(~m[19]&m[252]&m[253]&m[254]&m[255])|(m[19]&m[252]&m[253]&m[254]&m[255]));
    m[59] = (((m[19]&m[256]&~m[257]&~m[258]&~m[259])|(m[19]&~m[256]&m[257]&~m[258]&~m[259])|(~m[19]&m[256]&m[257]&~m[258]&~m[259])|(m[19]&~m[256]&~m[257]&m[258]&~m[259])|(~m[19]&m[256]&~m[257]&m[258]&~m[259])|(~m[19]&~m[256]&m[257]&m[258]&~m[259])|(m[19]&~m[256]&~m[257]&~m[258]&m[259])|(~m[19]&m[256]&~m[257]&~m[258]&m[259])|(~m[19]&~m[256]&m[257]&~m[258]&m[259])|(~m[19]&~m[256]&~m[257]&m[258]&m[259]))&BiasedRNG[138])|(((m[19]&m[256]&m[257]&~m[258]&~m[259])|(m[19]&m[256]&~m[257]&m[258]&~m[259])|(m[19]&~m[256]&m[257]&m[258]&~m[259])|(~m[19]&m[256]&m[257]&m[258]&~m[259])|(m[19]&m[256]&~m[257]&~m[258]&m[259])|(m[19]&~m[256]&m[257]&~m[258]&m[259])|(~m[19]&m[256]&m[257]&~m[258]&m[259])|(m[19]&~m[256]&~m[257]&m[258]&m[259])|(~m[19]&m[256]&~m[257]&m[258]&m[259])|(~m[19]&~m[256]&m[257]&m[258]&m[259]))&~BiasedRNG[138])|((m[19]&m[256]&m[257]&m[258]&~m[259])|(m[19]&m[256]&m[257]&~m[258]&m[259])|(m[19]&m[256]&~m[257]&m[258]&m[259])|(m[19]&~m[256]&m[257]&m[258]&m[259])|(~m[19]&m[256]&m[257]&m[258]&m[259])|(m[19]&m[256]&m[257]&m[258]&m[259]));
    m[60] = (((~m[0]&~m[160]&~m[260])|(m[0]&m[160]&~m[260]))&BiasedRNG[139])|(((m[0]&~m[160]&~m[260])|(~m[0]&m[160]&m[260]))&~BiasedRNG[139])|((~m[0]&~m[160]&m[260])|(m[0]&~m[160]&m[260])|(m[0]&m[160]&m[260]));
    m[61] = (((~m[0]&~m[170]&~m[270])|(m[0]&m[170]&~m[270]))&BiasedRNG[140])|(((m[0]&~m[170]&~m[270])|(~m[0]&m[170]&m[270]))&~BiasedRNG[140])|((~m[0]&~m[170]&m[270])|(m[0]&~m[170]&m[270])|(m[0]&m[170]&m[270]));
    m[70] = (((~m[1]&~m[161]&~m[261])|(m[1]&m[161]&~m[261]))&BiasedRNG[141])|(((m[1]&~m[161]&~m[261])|(~m[1]&m[161]&m[261]))&~BiasedRNG[141])|((~m[1]&~m[161]&m[261])|(m[1]&~m[161]&m[261])|(m[1]&m[161]&m[261]));
    m[71] = (((~m[1]&~m[171]&~m[271])|(m[1]&m[171]&~m[271]))&BiasedRNG[142])|(((m[1]&~m[171]&~m[271])|(~m[1]&m[171]&m[271]))&~BiasedRNG[142])|((~m[1]&~m[171]&m[271])|(m[1]&~m[171]&m[271])|(m[1]&m[171]&m[271]));
    m[80] = (((~m[2]&~m[162]&~m[262])|(m[2]&m[162]&~m[262]))&BiasedRNG[143])|(((m[2]&~m[162]&~m[262])|(~m[2]&m[162]&m[262]))&~BiasedRNG[143])|((~m[2]&~m[162]&m[262])|(m[2]&~m[162]&m[262])|(m[2]&m[162]&m[262]));
    m[81] = (((~m[2]&~m[172]&~m[272])|(m[2]&m[172]&~m[272]))&BiasedRNG[144])|(((m[2]&~m[172]&~m[272])|(~m[2]&m[172]&m[272]))&~BiasedRNG[144])|((~m[2]&~m[172]&m[272])|(m[2]&~m[172]&m[272])|(m[2]&m[172]&m[272]));
    m[90] = (((~m[3]&~m[163]&~m[263])|(m[3]&m[163]&~m[263]))&BiasedRNG[145])|(((m[3]&~m[163]&~m[263])|(~m[3]&m[163]&m[263]))&~BiasedRNG[145])|((~m[3]&~m[163]&m[263])|(m[3]&~m[163]&m[263])|(m[3]&m[163]&m[263]));
    m[91] = (((~m[3]&~m[173]&~m[273])|(m[3]&m[173]&~m[273]))&BiasedRNG[146])|(((m[3]&~m[173]&~m[273])|(~m[3]&m[173]&m[273]))&~BiasedRNG[146])|((~m[3]&~m[173]&m[273])|(m[3]&~m[173]&m[273])|(m[3]&m[173]&m[273]));
    m[100] = (((~m[4]&~m[164]&~m[264])|(m[4]&m[164]&~m[264]))&BiasedRNG[147])|(((m[4]&~m[164]&~m[264])|(~m[4]&m[164]&m[264]))&~BiasedRNG[147])|((~m[4]&~m[164]&m[264])|(m[4]&~m[164]&m[264])|(m[4]&m[164]&m[264]));
    m[101] = (((~m[4]&~m[174]&~m[274])|(m[4]&m[174]&~m[274]))&BiasedRNG[148])|(((m[4]&~m[174]&~m[274])|(~m[4]&m[174]&m[274]))&~BiasedRNG[148])|((~m[4]&~m[174]&m[274])|(m[4]&~m[174]&m[274])|(m[4]&m[174]&m[274]));
    m[110] = (((~m[5]&~m[165]&~m[265])|(m[5]&m[165]&~m[265]))&BiasedRNG[149])|(((m[5]&~m[165]&~m[265])|(~m[5]&m[165]&m[265]))&~BiasedRNG[149])|((~m[5]&~m[165]&m[265])|(m[5]&~m[165]&m[265])|(m[5]&m[165]&m[265]));
    m[111] = (((~m[5]&~m[175]&~m[275])|(m[5]&m[175]&~m[275]))&BiasedRNG[150])|(((m[5]&~m[175]&~m[275])|(~m[5]&m[175]&m[275]))&~BiasedRNG[150])|((~m[5]&~m[175]&m[275])|(m[5]&~m[175]&m[275])|(m[5]&m[175]&m[275]));
    m[120] = (((~m[6]&~m[166]&~m[266])|(m[6]&m[166]&~m[266]))&BiasedRNG[151])|(((m[6]&~m[166]&~m[266])|(~m[6]&m[166]&m[266]))&~BiasedRNG[151])|((~m[6]&~m[166]&m[266])|(m[6]&~m[166]&m[266])|(m[6]&m[166]&m[266]));
    m[121] = (((~m[6]&~m[176]&~m[276])|(m[6]&m[176]&~m[276]))&BiasedRNG[152])|(((m[6]&~m[176]&~m[276])|(~m[6]&m[176]&m[276]))&~BiasedRNG[152])|((~m[6]&~m[176]&m[276])|(m[6]&~m[176]&m[276])|(m[6]&m[176]&m[276]));
    m[130] = (((~m[7]&~m[167]&~m[267])|(m[7]&m[167]&~m[267]))&BiasedRNG[153])|(((m[7]&~m[167]&~m[267])|(~m[7]&m[167]&m[267]))&~BiasedRNG[153])|((~m[7]&~m[167]&m[267])|(m[7]&~m[167]&m[267])|(m[7]&m[167]&m[267]));
    m[131] = (((~m[7]&~m[177]&~m[277])|(m[7]&m[177]&~m[277]))&BiasedRNG[154])|(((m[7]&~m[177]&~m[277])|(~m[7]&m[177]&m[277]))&~BiasedRNG[154])|((~m[7]&~m[177]&m[277])|(m[7]&~m[177]&m[277])|(m[7]&m[177]&m[277]));
    m[140] = (((~m[8]&~m[168]&~m[268])|(m[8]&m[168]&~m[268]))&BiasedRNG[155])|(((m[8]&~m[168]&~m[268])|(~m[8]&m[168]&m[268]))&~BiasedRNG[155])|((~m[8]&~m[168]&m[268])|(m[8]&~m[168]&m[268])|(m[8]&m[168]&m[268]));
    m[141] = (((~m[8]&~m[178]&~m[278])|(m[8]&m[178]&~m[278]))&BiasedRNG[156])|(((m[8]&~m[178]&~m[278])|(~m[8]&m[178]&m[278]))&~BiasedRNG[156])|((~m[8]&~m[178]&m[278])|(m[8]&~m[178]&m[278])|(m[8]&m[178]&m[278]));
    m[150] = (((~m[9]&~m[169]&~m[269])|(m[9]&m[169]&~m[269]))&BiasedRNG[157])|(((m[9]&~m[169]&~m[269])|(~m[9]&m[169]&m[269]))&~BiasedRNG[157])|((~m[9]&~m[169]&m[269])|(m[9]&~m[169]&m[269])|(m[9]&m[169]&m[269]));
    m[151] = (((~m[9]&~m[179]&~m[279])|(m[9]&m[179]&~m[279]))&BiasedRNG[158])|(((m[9]&~m[179]&~m[279])|(~m[9]&m[179]&m[279]))&~BiasedRNG[158])|((~m[9]&~m[179]&m[279])|(m[9]&~m[179]&m[279])|(m[9]&m[179]&m[279]));
    m[180] = (((~m[12]&~m[62]&~m[280])|(m[12]&m[62]&~m[280]))&BiasedRNG[159])|(((m[12]&~m[62]&~m[280])|(~m[12]&m[62]&m[280]))&~BiasedRNG[159])|((~m[12]&~m[62]&m[280])|(m[12]&~m[62]&m[280])|(m[12]&m[62]&m[280]));
    m[181] = (((~m[12]&~m[72]&~m[281])|(m[12]&m[72]&~m[281]))&BiasedRNG[160])|(((m[12]&~m[72]&~m[281])|(~m[12]&m[72]&m[281]))&~BiasedRNG[160])|((~m[12]&~m[72]&m[281])|(m[12]&~m[72]&m[281])|(m[12]&m[72]&m[281]));
    m[190] = (((~m[13]&~m[63]&~m[290])|(m[13]&m[63]&~m[290]))&BiasedRNG[161])|(((m[13]&~m[63]&~m[290])|(~m[13]&m[63]&m[290]))&~BiasedRNG[161])|((~m[13]&~m[63]&m[290])|(m[13]&~m[63]&m[290])|(m[13]&m[63]&m[290]));
    m[191] = (((~m[13]&~m[73]&~m[291])|(m[13]&m[73]&~m[291]))&BiasedRNG[162])|(((m[13]&~m[73]&~m[291])|(~m[13]&m[73]&m[291]))&~BiasedRNG[162])|((~m[13]&~m[73]&m[291])|(m[13]&~m[73]&m[291])|(m[13]&m[73]&m[291]));
    m[200] = (((~m[14]&~m[64]&~m[300])|(m[14]&m[64]&~m[300]))&BiasedRNG[163])|(((m[14]&~m[64]&~m[300])|(~m[14]&m[64]&m[300]))&~BiasedRNG[163])|((~m[14]&~m[64]&m[300])|(m[14]&~m[64]&m[300])|(m[14]&m[64]&m[300]));
    m[201] = (((~m[14]&~m[74]&~m[301])|(m[14]&m[74]&~m[301]))&BiasedRNG[164])|(((m[14]&~m[74]&~m[301])|(~m[14]&m[74]&m[301]))&~BiasedRNG[164])|((~m[14]&~m[74]&m[301])|(m[14]&~m[74]&m[301])|(m[14]&m[74]&m[301]));
    m[210] = (((~m[15]&~m[65]&~m[310])|(m[15]&m[65]&~m[310]))&BiasedRNG[165])|(((m[15]&~m[65]&~m[310])|(~m[15]&m[65]&m[310]))&~BiasedRNG[165])|((~m[15]&~m[65]&m[310])|(m[15]&~m[65]&m[310])|(m[15]&m[65]&m[310]));
    m[211] = (((~m[15]&~m[75]&~m[311])|(m[15]&m[75]&~m[311]))&BiasedRNG[166])|(((m[15]&~m[75]&~m[311])|(~m[15]&m[75]&m[311]))&~BiasedRNG[166])|((~m[15]&~m[75]&m[311])|(m[15]&~m[75]&m[311])|(m[15]&m[75]&m[311]));
    m[220] = (((~m[16]&~m[66]&~m[320])|(m[16]&m[66]&~m[320]))&BiasedRNG[167])|(((m[16]&~m[66]&~m[320])|(~m[16]&m[66]&m[320]))&~BiasedRNG[167])|((~m[16]&~m[66]&m[320])|(m[16]&~m[66]&m[320])|(m[16]&m[66]&m[320]));
    m[221] = (((~m[16]&~m[76]&~m[321])|(m[16]&m[76]&~m[321]))&BiasedRNG[168])|(((m[16]&~m[76]&~m[321])|(~m[16]&m[76]&m[321]))&~BiasedRNG[168])|((~m[16]&~m[76]&m[321])|(m[16]&~m[76]&m[321])|(m[16]&m[76]&m[321]));
    m[230] = (((~m[17]&~m[67]&~m[330])|(m[17]&m[67]&~m[330]))&BiasedRNG[169])|(((m[17]&~m[67]&~m[330])|(~m[17]&m[67]&m[330]))&~BiasedRNG[169])|((~m[17]&~m[67]&m[330])|(m[17]&~m[67]&m[330])|(m[17]&m[67]&m[330]));
    m[231] = (((~m[17]&~m[77]&~m[331])|(m[17]&m[77]&~m[331]))&BiasedRNG[170])|(((m[17]&~m[77]&~m[331])|(~m[17]&m[77]&m[331]))&~BiasedRNG[170])|((~m[17]&~m[77]&m[331])|(m[17]&~m[77]&m[331])|(m[17]&m[77]&m[331]));
    m[240] = (((~m[18]&~m[68]&~m[340])|(m[18]&m[68]&~m[340]))&BiasedRNG[171])|(((m[18]&~m[68]&~m[340])|(~m[18]&m[68]&m[340]))&~BiasedRNG[171])|((~m[18]&~m[68]&m[340])|(m[18]&~m[68]&m[340])|(m[18]&m[68]&m[340]));
    m[241] = (((~m[18]&~m[78]&~m[341])|(m[18]&m[78]&~m[341]))&BiasedRNG[172])|(((m[18]&~m[78]&~m[341])|(~m[18]&m[78]&m[341]))&~BiasedRNG[172])|((~m[18]&~m[78]&m[341])|(m[18]&~m[78]&m[341])|(m[18]&m[78]&m[341]));
    m[250] = (((~m[19]&~m[69]&~m[350])|(m[19]&m[69]&~m[350]))&BiasedRNG[173])|(((m[19]&~m[69]&~m[350])|(~m[19]&m[69]&m[350]))&~BiasedRNG[173])|((~m[19]&~m[69]&m[350])|(m[19]&~m[69]&m[350])|(m[19]&m[69]&m[350]));
    m[251] = (((~m[19]&~m[79]&~m[351])|(m[19]&m[79]&~m[351]))&BiasedRNG[174])|(((m[19]&~m[79]&~m[351])|(~m[19]&m[79]&m[351]))&~BiasedRNG[174])|((~m[19]&~m[79]&m[351])|(m[19]&~m[79]&m[351])|(m[19]&m[79]&m[351]));
    m[282] = (((m[82]&~m[182]&m[396])|(~m[82]&m[182]&m[396]))&BiasedRNG[175])|(((m[82]&m[182]&~m[396]))&~BiasedRNG[175])|((m[82]&m[182]&m[396]));
    m[283] = (((m[92]&~m[183]&m[416])|(~m[92]&m[183]&m[416]))&BiasedRNG[176])|(((m[92]&m[183]&~m[416]))&~BiasedRNG[176])|((m[92]&m[183]&m[416]));
    m[284] = (((m[102]&~m[184]&m[441])|(~m[102]&m[184]&m[441]))&BiasedRNG[177])|(((m[102]&m[184]&~m[441]))&~BiasedRNG[177])|((m[102]&m[184]&m[441]));
    m[285] = (((m[112]&~m[185]&m[471])|(~m[112]&m[185]&m[471]))&BiasedRNG[178])|(((m[112]&m[185]&~m[471]))&~BiasedRNG[178])|((m[112]&m[185]&m[471]));
    m[286] = (((m[122]&~m[186]&m[506])|(~m[122]&m[186]&m[506]))&BiasedRNG[179])|(((m[122]&m[186]&~m[506]))&~BiasedRNG[179])|((m[122]&m[186]&m[506]));
    m[287] = (((m[132]&~m[187]&m[546])|(~m[132]&m[187]&m[546]))&BiasedRNG[180])|(((m[132]&m[187]&~m[546]))&~BiasedRNG[180])|((m[132]&m[187]&m[546]));
    m[288] = (((m[142]&~m[188]&m[591])|(~m[142]&m[188]&m[591]))&BiasedRNG[181])|(((m[142]&m[188]&~m[591]))&~BiasedRNG[181])|((m[142]&m[188]&m[591]));
    m[289] = (((m[152]&~m[189]&m[631])|(~m[152]&m[189]&m[631]))&BiasedRNG[182])|(((m[152]&m[189]&~m[631]))&~BiasedRNG[182])|((m[152]&m[189]&m[631]));
    m[292] = (((m[83]&~m[192]&m[421])|(~m[83]&m[192]&m[421]))&BiasedRNG[183])|(((m[83]&m[192]&~m[421]))&~BiasedRNG[183])|((m[83]&m[192]&m[421]));
    m[293] = (((m[93]&~m[193]&m[446])|(~m[93]&m[193]&m[446]))&BiasedRNG[184])|(((m[93]&m[193]&~m[446]))&~BiasedRNG[184])|((m[93]&m[193]&m[446]));
    m[294] = (((m[103]&~m[194]&m[476])|(~m[103]&m[194]&m[476]))&BiasedRNG[185])|(((m[103]&m[194]&~m[476]))&~BiasedRNG[185])|((m[103]&m[194]&m[476]));
    m[295] = (((m[113]&~m[195]&m[511])|(~m[113]&m[195]&m[511]))&BiasedRNG[186])|(((m[113]&m[195]&~m[511]))&~BiasedRNG[186])|((m[113]&m[195]&m[511]));
    m[296] = (((m[123]&~m[196]&m[551])|(~m[123]&m[196]&m[551]))&BiasedRNG[187])|(((m[123]&m[196]&~m[551]))&~BiasedRNG[187])|((m[123]&m[196]&m[551]));
    m[297] = (((m[133]&~m[197]&m[596])|(~m[133]&m[197]&m[596]))&BiasedRNG[188])|(((m[133]&m[197]&~m[596]))&~BiasedRNG[188])|((m[133]&m[197]&m[596]));
    m[298] = (((m[143]&~m[198]&m[636])|(~m[143]&m[198]&m[636]))&BiasedRNG[189])|(((m[143]&m[198]&~m[636]))&~BiasedRNG[189])|((m[143]&m[198]&m[636]));
    m[299] = (((m[153]&~m[199]&m[671])|(~m[153]&m[199]&m[671]))&BiasedRNG[190])|(((m[153]&m[199]&~m[671]))&~BiasedRNG[190])|((m[153]&m[199]&m[671]));
    m[302] = (((m[84]&~m[202]&m[451])|(~m[84]&m[202]&m[451]))&BiasedRNG[191])|(((m[84]&m[202]&~m[451]))&~BiasedRNG[191])|((m[84]&m[202]&m[451]));
    m[303] = (((m[94]&~m[203]&m[481])|(~m[94]&m[203]&m[481]))&BiasedRNG[192])|(((m[94]&m[203]&~m[481]))&~BiasedRNG[192])|((m[94]&m[203]&m[481]));
    m[304] = (((m[104]&~m[204]&m[516])|(~m[104]&m[204]&m[516]))&BiasedRNG[193])|(((m[104]&m[204]&~m[516]))&~BiasedRNG[193])|((m[104]&m[204]&m[516]));
    m[305] = (((m[114]&~m[205]&m[556])|(~m[114]&m[205]&m[556]))&BiasedRNG[194])|(((m[114]&m[205]&~m[556]))&~BiasedRNG[194])|((m[114]&m[205]&m[556]));
    m[306] = (((m[124]&~m[206]&m[601])|(~m[124]&m[206]&m[601]))&BiasedRNG[195])|(((m[124]&m[206]&~m[601]))&~BiasedRNG[195])|((m[124]&m[206]&m[601]));
    m[307] = (((m[134]&~m[207]&m[641])|(~m[134]&m[207]&m[641]))&BiasedRNG[196])|(((m[134]&m[207]&~m[641]))&~BiasedRNG[196])|((m[134]&m[207]&m[641]));
    m[308] = (((m[144]&~m[208]&m[676])|(~m[144]&m[208]&m[676]))&BiasedRNG[197])|(((m[144]&m[208]&~m[676]))&~BiasedRNG[197])|((m[144]&m[208]&m[676]));
    m[309] = (((m[154]&~m[209]&m[706])|(~m[154]&m[209]&m[706]))&BiasedRNG[198])|(((m[154]&m[209]&~m[706]))&~BiasedRNG[198])|((m[154]&m[209]&m[706]));
    m[312] = (((m[85]&~m[212]&m[486])|(~m[85]&m[212]&m[486]))&BiasedRNG[199])|(((m[85]&m[212]&~m[486]))&~BiasedRNG[199])|((m[85]&m[212]&m[486]));
    m[313] = (((m[95]&~m[213]&m[521])|(~m[95]&m[213]&m[521]))&BiasedRNG[200])|(((m[95]&m[213]&~m[521]))&~BiasedRNG[200])|((m[95]&m[213]&m[521]));
    m[314] = (((m[105]&~m[214]&m[561])|(~m[105]&m[214]&m[561]))&BiasedRNG[201])|(((m[105]&m[214]&~m[561]))&~BiasedRNG[201])|((m[105]&m[214]&m[561]));
    m[315] = (((m[115]&~m[215]&m[606])|(~m[115]&m[215]&m[606]))&BiasedRNG[202])|(((m[115]&m[215]&~m[606]))&~BiasedRNG[202])|((m[115]&m[215]&m[606]));
    m[316] = (((m[125]&~m[216]&m[646])|(~m[125]&m[216]&m[646]))&BiasedRNG[203])|(((m[125]&m[216]&~m[646]))&~BiasedRNG[203])|((m[125]&m[216]&m[646]));
    m[317] = (((m[135]&~m[217]&m[681])|(~m[135]&m[217]&m[681]))&BiasedRNG[204])|(((m[135]&m[217]&~m[681]))&~BiasedRNG[204])|((m[135]&m[217]&m[681]));
    m[318] = (((m[145]&~m[218]&m[711])|(~m[145]&m[218]&m[711]))&BiasedRNG[205])|(((m[145]&m[218]&~m[711]))&~BiasedRNG[205])|((m[145]&m[218]&m[711]));
    m[319] = (((m[155]&~m[219]&m[736])|(~m[155]&m[219]&m[736]))&BiasedRNG[206])|(((m[155]&m[219]&~m[736]))&~BiasedRNG[206])|((m[155]&m[219]&m[736]));
    m[322] = (((m[86]&~m[222]&m[526])|(~m[86]&m[222]&m[526]))&BiasedRNG[207])|(((m[86]&m[222]&~m[526]))&~BiasedRNG[207])|((m[86]&m[222]&m[526]));
    m[323] = (((m[96]&~m[223]&m[566])|(~m[96]&m[223]&m[566]))&BiasedRNG[208])|(((m[96]&m[223]&~m[566]))&~BiasedRNG[208])|((m[96]&m[223]&m[566]));
    m[324] = (((m[106]&~m[224]&m[611])|(~m[106]&m[224]&m[611]))&BiasedRNG[209])|(((m[106]&m[224]&~m[611]))&~BiasedRNG[209])|((m[106]&m[224]&m[611]));
    m[325] = (((m[116]&~m[225]&m[651])|(~m[116]&m[225]&m[651]))&BiasedRNG[210])|(((m[116]&m[225]&~m[651]))&~BiasedRNG[210])|((m[116]&m[225]&m[651]));
    m[326] = (((m[126]&~m[226]&m[686])|(~m[126]&m[226]&m[686]))&BiasedRNG[211])|(((m[126]&m[226]&~m[686]))&~BiasedRNG[211])|((m[126]&m[226]&m[686]));
    m[327] = (((m[136]&~m[227]&m[716])|(~m[136]&m[227]&m[716]))&BiasedRNG[212])|(((m[136]&m[227]&~m[716]))&~BiasedRNG[212])|((m[136]&m[227]&m[716]));
    m[328] = (((m[146]&~m[228]&m[741])|(~m[146]&m[228]&m[741]))&BiasedRNG[213])|(((m[146]&m[228]&~m[741]))&~BiasedRNG[213])|((m[146]&m[228]&m[741]));
    m[329] = (((m[156]&~m[229]&m[761])|(~m[156]&m[229]&m[761]))&BiasedRNG[214])|(((m[156]&m[229]&~m[761]))&~BiasedRNG[214])|((m[156]&m[229]&m[761]));
    m[332] = (((m[87]&~m[232]&m[571])|(~m[87]&m[232]&m[571]))&BiasedRNG[215])|(((m[87]&m[232]&~m[571]))&~BiasedRNG[215])|((m[87]&m[232]&m[571]));
    m[333] = (((m[97]&~m[233]&m[616])|(~m[97]&m[233]&m[616]))&BiasedRNG[216])|(((m[97]&m[233]&~m[616]))&~BiasedRNG[216])|((m[97]&m[233]&m[616]));
    m[334] = (((m[107]&~m[234]&m[656])|(~m[107]&m[234]&m[656]))&BiasedRNG[217])|(((m[107]&m[234]&~m[656]))&~BiasedRNG[217])|((m[107]&m[234]&m[656]));
    m[335] = (((m[117]&~m[235]&m[691])|(~m[117]&m[235]&m[691]))&BiasedRNG[218])|(((m[117]&m[235]&~m[691]))&~BiasedRNG[218])|((m[117]&m[235]&m[691]));
    m[336] = (((m[127]&~m[236]&m[721])|(~m[127]&m[236]&m[721]))&BiasedRNG[219])|(((m[127]&m[236]&~m[721]))&~BiasedRNG[219])|((m[127]&m[236]&m[721]));
    m[337] = (((m[137]&~m[237]&m[746])|(~m[137]&m[237]&m[746]))&BiasedRNG[220])|(((m[137]&m[237]&~m[746]))&~BiasedRNG[220])|((m[137]&m[237]&m[746]));
    m[338] = (((m[147]&~m[238]&m[766])|(~m[147]&m[238]&m[766]))&BiasedRNG[221])|(((m[147]&m[238]&~m[766]))&~BiasedRNG[221])|((m[147]&m[238]&m[766]));
    m[339] = (((m[157]&~m[239]&m[781])|(~m[157]&m[239]&m[781]))&BiasedRNG[222])|(((m[157]&m[239]&~m[781]))&~BiasedRNG[222])|((m[157]&m[239]&m[781]));
    m[342] = (((m[88]&~m[242]&m[621])|(~m[88]&m[242]&m[621]))&BiasedRNG[223])|(((m[88]&m[242]&~m[621]))&~BiasedRNG[223])|((m[88]&m[242]&m[621]));
    m[343] = (((m[98]&~m[243]&m[661])|(~m[98]&m[243]&m[661]))&BiasedRNG[224])|(((m[98]&m[243]&~m[661]))&~BiasedRNG[224])|((m[98]&m[243]&m[661]));
    m[344] = (((m[108]&~m[244]&m[696])|(~m[108]&m[244]&m[696]))&BiasedRNG[225])|(((m[108]&m[244]&~m[696]))&~BiasedRNG[225])|((m[108]&m[244]&m[696]));
    m[345] = (((m[118]&~m[245]&m[726])|(~m[118]&m[245]&m[726]))&BiasedRNG[226])|(((m[118]&m[245]&~m[726]))&~BiasedRNG[226])|((m[118]&m[245]&m[726]));
    m[346] = (((m[128]&~m[246]&m[751])|(~m[128]&m[246]&m[751]))&BiasedRNG[227])|(((m[128]&m[246]&~m[751]))&~BiasedRNG[227])|((m[128]&m[246]&m[751]));
    m[347] = (((m[138]&~m[247]&m[771])|(~m[138]&m[247]&m[771]))&BiasedRNG[228])|(((m[138]&m[247]&~m[771]))&~BiasedRNG[228])|((m[138]&m[247]&m[771]));
    m[348] = (((m[148]&~m[248]&m[786])|(~m[148]&m[248]&m[786]))&BiasedRNG[229])|(((m[148]&m[248]&~m[786]))&~BiasedRNG[229])|((m[148]&m[248]&m[786]));
    m[349] = (((m[158]&~m[249]&m[796])|(~m[158]&m[249]&m[796]))&BiasedRNG[230])|(((m[158]&m[249]&~m[796]))&~BiasedRNG[230])|((m[158]&m[249]&m[796]));
    m[352] = (((m[89]&~m[252]&m[666])|(~m[89]&m[252]&m[666]))&BiasedRNG[231])|(((m[89]&m[252]&~m[666]))&~BiasedRNG[231])|((m[89]&m[252]&m[666]));
    m[353] = (((m[99]&~m[253]&m[701])|(~m[99]&m[253]&m[701]))&BiasedRNG[232])|(((m[99]&m[253]&~m[701]))&~BiasedRNG[232])|((m[99]&m[253]&m[701]));
    m[354] = (((m[109]&~m[254]&m[731])|(~m[109]&m[254]&m[731]))&BiasedRNG[233])|(((m[109]&m[254]&~m[731]))&~BiasedRNG[233])|((m[109]&m[254]&m[731]));
    m[355] = (((m[119]&~m[255]&m[756])|(~m[119]&m[255]&m[756]))&BiasedRNG[234])|(((m[119]&m[255]&~m[756]))&~BiasedRNG[234])|((m[119]&m[255]&m[756]));
    m[356] = (((m[129]&~m[256]&m[776])|(~m[129]&m[256]&m[776]))&BiasedRNG[235])|(((m[129]&m[256]&~m[776]))&~BiasedRNG[235])|((m[129]&m[256]&m[776]));
    m[357] = (((m[139]&~m[257]&m[791])|(~m[139]&m[257]&m[791]))&BiasedRNG[236])|(((m[139]&m[257]&~m[791]))&~BiasedRNG[236])|((m[139]&m[257]&m[791]));
    m[358] = (((m[149]&~m[258]&m[801])|(~m[149]&m[258]&m[801]))&BiasedRNG[237])|(((m[149]&m[258]&~m[801]))&~BiasedRNG[237])|((m[149]&m[258]&m[801]));
    m[359] = (((m[159]&~m[259]&m[806])|(~m[159]&m[259]&m[806]))&BiasedRNG[238])|(((m[159]&m[259]&~m[806]))&~BiasedRNG[238])|((m[159]&m[259]&m[806]));
    m[360] = (((m[261]&~m[361]&~m[362]&~m[363]&~m[364])|(~m[261]&~m[361]&~m[362]&m[363]&~m[364])|(m[261]&m[361]&~m[362]&m[363]&~m[364])|(m[261]&~m[361]&m[362]&m[363]&~m[364])|(~m[261]&m[361]&~m[362]&~m[363]&m[364])|(~m[261]&~m[361]&m[362]&~m[363]&m[364])|(m[261]&m[361]&m[362]&~m[363]&m[364])|(~m[261]&m[361]&m[362]&m[363]&m[364]))&UnbiasedRNG[108])|((m[261]&~m[361]&~m[362]&m[363]&~m[364])|(~m[261]&~m[361]&~m[362]&~m[363]&m[364])|(m[261]&~m[361]&~m[362]&~m[363]&m[364])|(m[261]&m[361]&~m[362]&~m[363]&m[364])|(m[261]&~m[361]&m[362]&~m[363]&m[364])|(~m[261]&~m[361]&~m[362]&m[363]&m[364])|(m[261]&~m[361]&~m[362]&m[363]&m[364])|(~m[261]&m[361]&~m[362]&m[363]&m[364])|(m[261]&m[361]&~m[362]&m[363]&m[364])|(~m[261]&~m[361]&m[362]&m[363]&m[364])|(m[261]&~m[361]&m[362]&m[363]&m[364])|(m[261]&m[361]&m[362]&m[363]&m[364]));
    m[366] = (((m[271]&~m[365]&~m[367]&~m[368]&~m[369])|(~m[271]&~m[365]&~m[367]&m[368]&~m[369])|(m[271]&m[365]&~m[367]&m[368]&~m[369])|(m[271]&~m[365]&m[367]&m[368]&~m[369])|(~m[271]&m[365]&~m[367]&~m[368]&m[369])|(~m[271]&~m[365]&m[367]&~m[368]&m[369])|(m[271]&m[365]&m[367]&~m[368]&m[369])|(~m[271]&m[365]&m[367]&m[368]&m[369]))&UnbiasedRNG[109])|((m[271]&~m[365]&~m[367]&m[368]&~m[369])|(~m[271]&~m[365]&~m[367]&~m[368]&m[369])|(m[271]&~m[365]&~m[367]&~m[368]&m[369])|(m[271]&m[365]&~m[367]&~m[368]&m[369])|(m[271]&~m[365]&m[367]&~m[368]&m[369])|(~m[271]&~m[365]&~m[367]&m[368]&m[369])|(m[271]&~m[365]&~m[367]&m[368]&m[369])|(~m[271]&m[365]&~m[367]&m[368]&m[369])|(m[271]&m[365]&~m[367]&m[368]&m[369])|(~m[271]&~m[365]&m[367]&m[368]&m[369])|(m[271]&~m[365]&m[367]&m[368]&m[369])|(m[271]&m[365]&m[367]&m[368]&m[369]));
    m[371] = (((m[280]&~m[370]&~m[372]&~m[373]&~m[374])|(~m[280]&~m[370]&~m[372]&m[373]&~m[374])|(m[280]&m[370]&~m[372]&m[373]&~m[374])|(m[280]&~m[370]&m[372]&m[373]&~m[374])|(~m[280]&m[370]&~m[372]&~m[373]&m[374])|(~m[280]&~m[370]&m[372]&~m[373]&m[374])|(m[280]&m[370]&m[372]&~m[373]&m[374])|(~m[280]&m[370]&m[372]&m[373]&m[374]))&UnbiasedRNG[110])|((m[280]&~m[370]&~m[372]&m[373]&~m[374])|(~m[280]&~m[370]&~m[372]&~m[373]&m[374])|(m[280]&~m[370]&~m[372]&~m[373]&m[374])|(m[280]&m[370]&~m[372]&~m[373]&m[374])|(m[280]&~m[370]&m[372]&~m[373]&m[374])|(~m[280]&~m[370]&~m[372]&m[373]&m[374])|(m[280]&~m[370]&~m[372]&m[373]&m[374])|(~m[280]&m[370]&~m[372]&m[373]&m[374])|(m[280]&m[370]&~m[372]&m[373]&m[374])|(~m[280]&~m[370]&m[372]&m[373]&m[374])|(m[280]&~m[370]&m[372]&m[373]&m[374])|(m[280]&m[370]&m[372]&m[373]&m[374]));
    m[376] = (((m[272]&~m[375]&~m[377]&~m[378]&~m[379])|(~m[272]&~m[375]&~m[377]&m[378]&~m[379])|(m[272]&m[375]&~m[377]&m[378]&~m[379])|(m[272]&~m[375]&m[377]&m[378]&~m[379])|(~m[272]&m[375]&~m[377]&~m[378]&m[379])|(~m[272]&~m[375]&m[377]&~m[378]&m[379])|(m[272]&m[375]&m[377]&~m[378]&m[379])|(~m[272]&m[375]&m[377]&m[378]&m[379]))&UnbiasedRNG[111])|((m[272]&~m[375]&~m[377]&m[378]&~m[379])|(~m[272]&~m[375]&~m[377]&~m[378]&m[379])|(m[272]&~m[375]&~m[377]&~m[378]&m[379])|(m[272]&m[375]&~m[377]&~m[378]&m[379])|(m[272]&~m[375]&m[377]&~m[378]&m[379])|(~m[272]&~m[375]&~m[377]&m[378]&m[379])|(m[272]&~m[375]&~m[377]&m[378]&m[379])|(~m[272]&m[375]&~m[377]&m[378]&m[379])|(m[272]&m[375]&~m[377]&m[378]&m[379])|(~m[272]&~m[375]&m[377]&m[378]&m[379])|(m[272]&~m[375]&m[377]&m[378]&m[379])|(m[272]&m[375]&m[377]&m[378]&m[379]));
    m[381] = (((m[281]&~m[380]&~m[382]&~m[383]&~m[384])|(~m[281]&~m[380]&~m[382]&m[383]&~m[384])|(m[281]&m[380]&~m[382]&m[383]&~m[384])|(m[281]&~m[380]&m[382]&m[383]&~m[384])|(~m[281]&m[380]&~m[382]&~m[383]&m[384])|(~m[281]&~m[380]&m[382]&~m[383]&m[384])|(m[281]&m[380]&m[382]&~m[383]&m[384])|(~m[281]&m[380]&m[382]&m[383]&m[384]))&UnbiasedRNG[112])|((m[281]&~m[380]&~m[382]&m[383]&~m[384])|(~m[281]&~m[380]&~m[382]&~m[383]&m[384])|(m[281]&~m[380]&~m[382]&~m[383]&m[384])|(m[281]&m[380]&~m[382]&~m[383]&m[384])|(m[281]&~m[380]&m[382]&~m[383]&m[384])|(~m[281]&~m[380]&~m[382]&m[383]&m[384])|(m[281]&~m[380]&~m[382]&m[383]&m[384])|(~m[281]&m[380]&~m[382]&m[383]&m[384])|(m[281]&m[380]&~m[382]&m[383]&m[384])|(~m[281]&~m[380]&m[382]&m[383]&m[384])|(m[281]&~m[380]&m[382]&m[383]&m[384])|(m[281]&m[380]&m[382]&m[383]&m[384]));
    m[386] = (((m[290]&~m[385]&~m[387]&~m[388]&~m[389])|(~m[290]&~m[385]&~m[387]&m[388]&~m[389])|(m[290]&m[385]&~m[387]&m[388]&~m[389])|(m[290]&~m[385]&m[387]&m[388]&~m[389])|(~m[290]&m[385]&~m[387]&~m[388]&m[389])|(~m[290]&~m[385]&m[387]&~m[388]&m[389])|(m[290]&m[385]&m[387]&~m[388]&m[389])|(~m[290]&m[385]&m[387]&m[388]&m[389]))&UnbiasedRNG[113])|((m[290]&~m[385]&~m[387]&m[388]&~m[389])|(~m[290]&~m[385]&~m[387]&~m[388]&m[389])|(m[290]&~m[385]&~m[387]&~m[388]&m[389])|(m[290]&m[385]&~m[387]&~m[388]&m[389])|(m[290]&~m[385]&m[387]&~m[388]&m[389])|(~m[290]&~m[385]&~m[387]&m[388]&m[389])|(m[290]&~m[385]&~m[387]&m[388]&m[389])|(~m[290]&m[385]&~m[387]&m[388]&m[389])|(m[290]&m[385]&~m[387]&m[388]&m[389])|(~m[290]&~m[385]&m[387]&m[388]&m[389])|(m[290]&~m[385]&m[387]&m[388]&m[389])|(m[290]&m[385]&m[387]&m[388]&m[389]));
    m[391] = (((m[273]&~m[390]&~m[392]&~m[393]&~m[394])|(~m[273]&~m[390]&~m[392]&m[393]&~m[394])|(m[273]&m[390]&~m[392]&m[393]&~m[394])|(m[273]&~m[390]&m[392]&m[393]&~m[394])|(~m[273]&m[390]&~m[392]&~m[393]&m[394])|(~m[273]&~m[390]&m[392]&~m[393]&m[394])|(m[273]&m[390]&m[392]&~m[393]&m[394])|(~m[273]&m[390]&m[392]&m[393]&m[394]))&UnbiasedRNG[114])|((m[273]&~m[390]&~m[392]&m[393]&~m[394])|(~m[273]&~m[390]&~m[392]&~m[393]&m[394])|(m[273]&~m[390]&~m[392]&~m[393]&m[394])|(m[273]&m[390]&~m[392]&~m[393]&m[394])|(m[273]&~m[390]&m[392]&~m[393]&m[394])|(~m[273]&~m[390]&~m[392]&m[393]&m[394])|(m[273]&~m[390]&~m[392]&m[393]&m[394])|(~m[273]&m[390]&~m[392]&m[393]&m[394])|(m[273]&m[390]&~m[392]&m[393]&m[394])|(~m[273]&~m[390]&m[392]&m[393]&m[394])|(m[273]&~m[390]&m[392]&m[393]&m[394])|(m[273]&m[390]&m[392]&m[393]&m[394]));
    m[397] = (((m[384]&~m[395]&~m[396]&~m[398]&~m[399])|(~m[384]&~m[395]&~m[396]&m[398]&~m[399])|(m[384]&m[395]&~m[396]&m[398]&~m[399])|(m[384]&~m[395]&m[396]&m[398]&~m[399])|(~m[384]&m[395]&~m[396]&~m[398]&m[399])|(~m[384]&~m[395]&m[396]&~m[398]&m[399])|(m[384]&m[395]&m[396]&~m[398]&m[399])|(~m[384]&m[395]&m[396]&m[398]&m[399]))&UnbiasedRNG[115])|((m[384]&~m[395]&~m[396]&m[398]&~m[399])|(~m[384]&~m[395]&~m[396]&~m[398]&m[399])|(m[384]&~m[395]&~m[396]&~m[398]&m[399])|(m[384]&m[395]&~m[396]&~m[398]&m[399])|(m[384]&~m[395]&m[396]&~m[398]&m[399])|(~m[384]&~m[395]&~m[396]&m[398]&m[399])|(m[384]&~m[395]&~m[396]&m[398]&m[399])|(~m[384]&m[395]&~m[396]&m[398]&m[399])|(m[384]&m[395]&~m[396]&m[398]&m[399])|(~m[384]&~m[395]&m[396]&m[398]&m[399])|(m[384]&~m[395]&m[396]&m[398]&m[399])|(m[384]&m[395]&m[396]&m[398]&m[399]));
    m[401] = (((m[291]&~m[400]&~m[402]&~m[403]&~m[404])|(~m[291]&~m[400]&~m[402]&m[403]&~m[404])|(m[291]&m[400]&~m[402]&m[403]&~m[404])|(m[291]&~m[400]&m[402]&m[403]&~m[404])|(~m[291]&m[400]&~m[402]&~m[403]&m[404])|(~m[291]&~m[400]&m[402]&~m[403]&m[404])|(m[291]&m[400]&m[402]&~m[403]&m[404])|(~m[291]&m[400]&m[402]&m[403]&m[404]))&UnbiasedRNG[116])|((m[291]&~m[400]&~m[402]&m[403]&~m[404])|(~m[291]&~m[400]&~m[402]&~m[403]&m[404])|(m[291]&~m[400]&~m[402]&~m[403]&m[404])|(m[291]&m[400]&~m[402]&~m[403]&m[404])|(m[291]&~m[400]&m[402]&~m[403]&m[404])|(~m[291]&~m[400]&~m[402]&m[403]&m[404])|(m[291]&~m[400]&~m[402]&m[403]&m[404])|(~m[291]&m[400]&~m[402]&m[403]&m[404])|(m[291]&m[400]&~m[402]&m[403]&m[404])|(~m[291]&~m[400]&m[402]&m[403]&m[404])|(m[291]&~m[400]&m[402]&m[403]&m[404])|(m[291]&m[400]&m[402]&m[403]&m[404]));
    m[406] = (((m[300]&~m[405]&~m[407]&~m[408]&~m[409])|(~m[300]&~m[405]&~m[407]&m[408]&~m[409])|(m[300]&m[405]&~m[407]&m[408]&~m[409])|(m[300]&~m[405]&m[407]&m[408]&~m[409])|(~m[300]&m[405]&~m[407]&~m[408]&m[409])|(~m[300]&~m[405]&m[407]&~m[408]&m[409])|(m[300]&m[405]&m[407]&~m[408]&m[409])|(~m[300]&m[405]&m[407]&m[408]&m[409]))&UnbiasedRNG[117])|((m[300]&~m[405]&~m[407]&m[408]&~m[409])|(~m[300]&~m[405]&~m[407]&~m[408]&m[409])|(m[300]&~m[405]&~m[407]&~m[408]&m[409])|(m[300]&m[405]&~m[407]&~m[408]&m[409])|(m[300]&~m[405]&m[407]&~m[408]&m[409])|(~m[300]&~m[405]&~m[407]&m[408]&m[409])|(m[300]&~m[405]&~m[407]&m[408]&m[409])|(~m[300]&m[405]&~m[407]&m[408]&m[409])|(m[300]&m[405]&~m[407]&m[408]&m[409])|(~m[300]&~m[405]&m[407]&m[408]&m[409])|(m[300]&~m[405]&m[407]&m[408]&m[409])|(m[300]&m[405]&m[407]&m[408]&m[409]));
    m[411] = (((m[274]&~m[410]&~m[412]&~m[413]&~m[414])|(~m[274]&~m[410]&~m[412]&m[413]&~m[414])|(m[274]&m[410]&~m[412]&m[413]&~m[414])|(m[274]&~m[410]&m[412]&m[413]&~m[414])|(~m[274]&m[410]&~m[412]&~m[413]&m[414])|(~m[274]&~m[410]&m[412]&~m[413]&m[414])|(m[274]&m[410]&m[412]&~m[413]&m[414])|(~m[274]&m[410]&m[412]&m[413]&m[414]))&UnbiasedRNG[118])|((m[274]&~m[410]&~m[412]&m[413]&~m[414])|(~m[274]&~m[410]&~m[412]&~m[413]&m[414])|(m[274]&~m[410]&~m[412]&~m[413]&m[414])|(m[274]&m[410]&~m[412]&~m[413]&m[414])|(m[274]&~m[410]&m[412]&~m[413]&m[414])|(~m[274]&~m[410]&~m[412]&m[413]&m[414])|(m[274]&~m[410]&~m[412]&m[413]&m[414])|(~m[274]&m[410]&~m[412]&m[413]&m[414])|(m[274]&m[410]&~m[412]&m[413]&m[414])|(~m[274]&~m[410]&m[412]&m[413]&m[414])|(m[274]&~m[410]&m[412]&m[413]&m[414])|(m[274]&m[410]&m[412]&m[413]&m[414]));
    m[417] = (((m[399]&~m[415]&~m[416]&~m[418]&~m[419])|(~m[399]&~m[415]&~m[416]&m[418]&~m[419])|(m[399]&m[415]&~m[416]&m[418]&~m[419])|(m[399]&~m[415]&m[416]&m[418]&~m[419])|(~m[399]&m[415]&~m[416]&~m[418]&m[419])|(~m[399]&~m[415]&m[416]&~m[418]&m[419])|(m[399]&m[415]&m[416]&~m[418]&m[419])|(~m[399]&m[415]&m[416]&m[418]&m[419]))&UnbiasedRNG[119])|((m[399]&~m[415]&~m[416]&m[418]&~m[419])|(~m[399]&~m[415]&~m[416]&~m[418]&m[419])|(m[399]&~m[415]&~m[416]&~m[418]&m[419])|(m[399]&m[415]&~m[416]&~m[418]&m[419])|(m[399]&~m[415]&m[416]&~m[418]&m[419])|(~m[399]&~m[415]&~m[416]&m[418]&m[419])|(m[399]&~m[415]&~m[416]&m[418]&m[419])|(~m[399]&m[415]&~m[416]&m[418]&m[419])|(m[399]&m[415]&~m[416]&m[418]&m[419])|(~m[399]&~m[415]&m[416]&m[418]&m[419])|(m[399]&~m[415]&m[416]&m[418]&m[419])|(m[399]&m[415]&m[416]&m[418]&m[419]));
    m[422] = (((m[404]&~m[420]&~m[421]&~m[423]&~m[424])|(~m[404]&~m[420]&~m[421]&m[423]&~m[424])|(m[404]&m[420]&~m[421]&m[423]&~m[424])|(m[404]&~m[420]&m[421]&m[423]&~m[424])|(~m[404]&m[420]&~m[421]&~m[423]&m[424])|(~m[404]&~m[420]&m[421]&~m[423]&m[424])|(m[404]&m[420]&m[421]&~m[423]&m[424])|(~m[404]&m[420]&m[421]&m[423]&m[424]))&UnbiasedRNG[120])|((m[404]&~m[420]&~m[421]&m[423]&~m[424])|(~m[404]&~m[420]&~m[421]&~m[423]&m[424])|(m[404]&~m[420]&~m[421]&~m[423]&m[424])|(m[404]&m[420]&~m[421]&~m[423]&m[424])|(m[404]&~m[420]&m[421]&~m[423]&m[424])|(~m[404]&~m[420]&~m[421]&m[423]&m[424])|(m[404]&~m[420]&~m[421]&m[423]&m[424])|(~m[404]&m[420]&~m[421]&m[423]&m[424])|(m[404]&m[420]&~m[421]&m[423]&m[424])|(~m[404]&~m[420]&m[421]&m[423]&m[424])|(m[404]&~m[420]&m[421]&m[423]&m[424])|(m[404]&m[420]&m[421]&m[423]&m[424]));
    m[426] = (((m[301]&~m[425]&~m[427]&~m[428]&~m[429])|(~m[301]&~m[425]&~m[427]&m[428]&~m[429])|(m[301]&m[425]&~m[427]&m[428]&~m[429])|(m[301]&~m[425]&m[427]&m[428]&~m[429])|(~m[301]&m[425]&~m[427]&~m[428]&m[429])|(~m[301]&~m[425]&m[427]&~m[428]&m[429])|(m[301]&m[425]&m[427]&~m[428]&m[429])|(~m[301]&m[425]&m[427]&m[428]&m[429]))&UnbiasedRNG[121])|((m[301]&~m[425]&~m[427]&m[428]&~m[429])|(~m[301]&~m[425]&~m[427]&~m[428]&m[429])|(m[301]&~m[425]&~m[427]&~m[428]&m[429])|(m[301]&m[425]&~m[427]&~m[428]&m[429])|(m[301]&~m[425]&m[427]&~m[428]&m[429])|(~m[301]&~m[425]&~m[427]&m[428]&m[429])|(m[301]&~m[425]&~m[427]&m[428]&m[429])|(~m[301]&m[425]&~m[427]&m[428]&m[429])|(m[301]&m[425]&~m[427]&m[428]&m[429])|(~m[301]&~m[425]&m[427]&m[428]&m[429])|(m[301]&~m[425]&m[427]&m[428]&m[429])|(m[301]&m[425]&m[427]&m[428]&m[429]));
    m[431] = (((m[310]&~m[430]&~m[432]&~m[433]&~m[434])|(~m[310]&~m[430]&~m[432]&m[433]&~m[434])|(m[310]&m[430]&~m[432]&m[433]&~m[434])|(m[310]&~m[430]&m[432]&m[433]&~m[434])|(~m[310]&m[430]&~m[432]&~m[433]&m[434])|(~m[310]&~m[430]&m[432]&~m[433]&m[434])|(m[310]&m[430]&m[432]&~m[433]&m[434])|(~m[310]&m[430]&m[432]&m[433]&m[434]))&UnbiasedRNG[122])|((m[310]&~m[430]&~m[432]&m[433]&~m[434])|(~m[310]&~m[430]&~m[432]&~m[433]&m[434])|(m[310]&~m[430]&~m[432]&~m[433]&m[434])|(m[310]&m[430]&~m[432]&~m[433]&m[434])|(m[310]&~m[430]&m[432]&~m[433]&m[434])|(~m[310]&~m[430]&~m[432]&m[433]&m[434])|(m[310]&~m[430]&~m[432]&m[433]&m[434])|(~m[310]&m[430]&~m[432]&m[433]&m[434])|(m[310]&m[430]&~m[432]&m[433]&m[434])|(~m[310]&~m[430]&m[432]&m[433]&m[434])|(m[310]&~m[430]&m[432]&m[433]&m[434])|(m[310]&m[430]&m[432]&m[433]&m[434]));
    m[436] = (((m[275]&~m[435]&~m[437]&~m[438]&~m[439])|(~m[275]&~m[435]&~m[437]&m[438]&~m[439])|(m[275]&m[435]&~m[437]&m[438]&~m[439])|(m[275]&~m[435]&m[437]&m[438]&~m[439])|(~m[275]&m[435]&~m[437]&~m[438]&m[439])|(~m[275]&~m[435]&m[437]&~m[438]&m[439])|(m[275]&m[435]&m[437]&~m[438]&m[439])|(~m[275]&m[435]&m[437]&m[438]&m[439]))&UnbiasedRNG[123])|((m[275]&~m[435]&~m[437]&m[438]&~m[439])|(~m[275]&~m[435]&~m[437]&~m[438]&m[439])|(m[275]&~m[435]&~m[437]&~m[438]&m[439])|(m[275]&m[435]&~m[437]&~m[438]&m[439])|(m[275]&~m[435]&m[437]&~m[438]&m[439])|(~m[275]&~m[435]&~m[437]&m[438]&m[439])|(m[275]&~m[435]&~m[437]&m[438]&m[439])|(~m[275]&m[435]&~m[437]&m[438]&m[439])|(m[275]&m[435]&~m[437]&m[438]&m[439])|(~m[275]&~m[435]&m[437]&m[438]&m[439])|(m[275]&~m[435]&m[437]&m[438]&m[439])|(m[275]&m[435]&m[437]&m[438]&m[439]));
    m[442] = (((m[419]&~m[440]&~m[441]&~m[443]&~m[444])|(~m[419]&~m[440]&~m[441]&m[443]&~m[444])|(m[419]&m[440]&~m[441]&m[443]&~m[444])|(m[419]&~m[440]&m[441]&m[443]&~m[444])|(~m[419]&m[440]&~m[441]&~m[443]&m[444])|(~m[419]&~m[440]&m[441]&~m[443]&m[444])|(m[419]&m[440]&m[441]&~m[443]&m[444])|(~m[419]&m[440]&m[441]&m[443]&m[444]))&UnbiasedRNG[124])|((m[419]&~m[440]&~m[441]&m[443]&~m[444])|(~m[419]&~m[440]&~m[441]&~m[443]&m[444])|(m[419]&~m[440]&~m[441]&~m[443]&m[444])|(m[419]&m[440]&~m[441]&~m[443]&m[444])|(m[419]&~m[440]&m[441]&~m[443]&m[444])|(~m[419]&~m[440]&~m[441]&m[443]&m[444])|(m[419]&~m[440]&~m[441]&m[443]&m[444])|(~m[419]&m[440]&~m[441]&m[443]&m[444])|(m[419]&m[440]&~m[441]&m[443]&m[444])|(~m[419]&~m[440]&m[441]&m[443]&m[444])|(m[419]&~m[440]&m[441]&m[443]&m[444])|(m[419]&m[440]&m[441]&m[443]&m[444]));
    m[447] = (((m[424]&~m[445]&~m[446]&~m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&m[448]&~m[449])|(m[424]&m[445]&~m[446]&m[448]&~m[449])|(m[424]&~m[445]&m[446]&m[448]&~m[449])|(~m[424]&m[445]&~m[446]&~m[448]&m[449])|(~m[424]&~m[445]&m[446]&~m[448]&m[449])|(m[424]&m[445]&m[446]&~m[448]&m[449])|(~m[424]&m[445]&m[446]&m[448]&m[449]))&UnbiasedRNG[125])|((m[424]&~m[445]&~m[446]&m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&m[446]&~m[448]&m[449])|(~m[424]&~m[445]&~m[446]&m[448]&m[449])|(m[424]&~m[445]&~m[446]&m[448]&m[449])|(~m[424]&m[445]&~m[446]&m[448]&m[449])|(m[424]&m[445]&~m[446]&m[448]&m[449])|(~m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&m[445]&m[446]&m[448]&m[449]));
    m[452] = (((m[429]&~m[450]&~m[451]&~m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&m[453]&~m[454])|(m[429]&m[450]&~m[451]&m[453]&~m[454])|(m[429]&~m[450]&m[451]&m[453]&~m[454])|(~m[429]&m[450]&~m[451]&~m[453]&m[454])|(~m[429]&~m[450]&m[451]&~m[453]&m[454])|(m[429]&m[450]&m[451]&~m[453]&m[454])|(~m[429]&m[450]&m[451]&m[453]&m[454]))&UnbiasedRNG[126])|((m[429]&~m[450]&~m[451]&m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&m[451]&~m[453]&m[454])|(~m[429]&~m[450]&~m[451]&m[453]&m[454])|(m[429]&~m[450]&~m[451]&m[453]&m[454])|(~m[429]&m[450]&~m[451]&m[453]&m[454])|(m[429]&m[450]&~m[451]&m[453]&m[454])|(~m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&m[450]&m[451]&m[453]&m[454]));
    m[456] = (((m[311]&~m[455]&~m[457]&~m[458]&~m[459])|(~m[311]&~m[455]&~m[457]&m[458]&~m[459])|(m[311]&m[455]&~m[457]&m[458]&~m[459])|(m[311]&~m[455]&m[457]&m[458]&~m[459])|(~m[311]&m[455]&~m[457]&~m[458]&m[459])|(~m[311]&~m[455]&m[457]&~m[458]&m[459])|(m[311]&m[455]&m[457]&~m[458]&m[459])|(~m[311]&m[455]&m[457]&m[458]&m[459]))&UnbiasedRNG[127])|((m[311]&~m[455]&~m[457]&m[458]&~m[459])|(~m[311]&~m[455]&~m[457]&~m[458]&m[459])|(m[311]&~m[455]&~m[457]&~m[458]&m[459])|(m[311]&m[455]&~m[457]&~m[458]&m[459])|(m[311]&~m[455]&m[457]&~m[458]&m[459])|(~m[311]&~m[455]&~m[457]&m[458]&m[459])|(m[311]&~m[455]&~m[457]&m[458]&m[459])|(~m[311]&m[455]&~m[457]&m[458]&m[459])|(m[311]&m[455]&~m[457]&m[458]&m[459])|(~m[311]&~m[455]&m[457]&m[458]&m[459])|(m[311]&~m[455]&m[457]&m[458]&m[459])|(m[311]&m[455]&m[457]&m[458]&m[459]));
    m[461] = (((m[320]&~m[460]&~m[462]&~m[463]&~m[464])|(~m[320]&~m[460]&~m[462]&m[463]&~m[464])|(m[320]&m[460]&~m[462]&m[463]&~m[464])|(m[320]&~m[460]&m[462]&m[463]&~m[464])|(~m[320]&m[460]&~m[462]&~m[463]&m[464])|(~m[320]&~m[460]&m[462]&~m[463]&m[464])|(m[320]&m[460]&m[462]&~m[463]&m[464])|(~m[320]&m[460]&m[462]&m[463]&m[464]))&UnbiasedRNG[128])|((m[320]&~m[460]&~m[462]&m[463]&~m[464])|(~m[320]&~m[460]&~m[462]&~m[463]&m[464])|(m[320]&~m[460]&~m[462]&~m[463]&m[464])|(m[320]&m[460]&~m[462]&~m[463]&m[464])|(m[320]&~m[460]&m[462]&~m[463]&m[464])|(~m[320]&~m[460]&~m[462]&m[463]&m[464])|(m[320]&~m[460]&~m[462]&m[463]&m[464])|(~m[320]&m[460]&~m[462]&m[463]&m[464])|(m[320]&m[460]&~m[462]&m[463]&m[464])|(~m[320]&~m[460]&m[462]&m[463]&m[464])|(m[320]&~m[460]&m[462]&m[463]&m[464])|(m[320]&m[460]&m[462]&m[463]&m[464]));
    m[466] = (((m[276]&~m[465]&~m[467]&~m[468]&~m[469])|(~m[276]&~m[465]&~m[467]&m[468]&~m[469])|(m[276]&m[465]&~m[467]&m[468]&~m[469])|(m[276]&~m[465]&m[467]&m[468]&~m[469])|(~m[276]&m[465]&~m[467]&~m[468]&m[469])|(~m[276]&~m[465]&m[467]&~m[468]&m[469])|(m[276]&m[465]&m[467]&~m[468]&m[469])|(~m[276]&m[465]&m[467]&m[468]&m[469]))&UnbiasedRNG[129])|((m[276]&~m[465]&~m[467]&m[468]&~m[469])|(~m[276]&~m[465]&~m[467]&~m[468]&m[469])|(m[276]&~m[465]&~m[467]&~m[468]&m[469])|(m[276]&m[465]&~m[467]&~m[468]&m[469])|(m[276]&~m[465]&m[467]&~m[468]&m[469])|(~m[276]&~m[465]&~m[467]&m[468]&m[469])|(m[276]&~m[465]&~m[467]&m[468]&m[469])|(~m[276]&m[465]&~m[467]&m[468]&m[469])|(m[276]&m[465]&~m[467]&m[468]&m[469])|(~m[276]&~m[465]&m[467]&m[468]&m[469])|(m[276]&~m[465]&m[467]&m[468]&m[469])|(m[276]&m[465]&m[467]&m[468]&m[469]));
    m[472] = (((m[444]&~m[470]&~m[471]&~m[473]&~m[474])|(~m[444]&~m[470]&~m[471]&m[473]&~m[474])|(m[444]&m[470]&~m[471]&m[473]&~m[474])|(m[444]&~m[470]&m[471]&m[473]&~m[474])|(~m[444]&m[470]&~m[471]&~m[473]&m[474])|(~m[444]&~m[470]&m[471]&~m[473]&m[474])|(m[444]&m[470]&m[471]&~m[473]&m[474])|(~m[444]&m[470]&m[471]&m[473]&m[474]))&UnbiasedRNG[130])|((m[444]&~m[470]&~m[471]&m[473]&~m[474])|(~m[444]&~m[470]&~m[471]&~m[473]&m[474])|(m[444]&~m[470]&~m[471]&~m[473]&m[474])|(m[444]&m[470]&~m[471]&~m[473]&m[474])|(m[444]&~m[470]&m[471]&~m[473]&m[474])|(~m[444]&~m[470]&~m[471]&m[473]&m[474])|(m[444]&~m[470]&~m[471]&m[473]&m[474])|(~m[444]&m[470]&~m[471]&m[473]&m[474])|(m[444]&m[470]&~m[471]&m[473]&m[474])|(~m[444]&~m[470]&m[471]&m[473]&m[474])|(m[444]&~m[470]&m[471]&m[473]&m[474])|(m[444]&m[470]&m[471]&m[473]&m[474]));
    m[477] = (((m[449]&~m[475]&~m[476]&~m[478]&~m[479])|(~m[449]&~m[475]&~m[476]&m[478]&~m[479])|(m[449]&m[475]&~m[476]&m[478]&~m[479])|(m[449]&~m[475]&m[476]&m[478]&~m[479])|(~m[449]&m[475]&~m[476]&~m[478]&m[479])|(~m[449]&~m[475]&m[476]&~m[478]&m[479])|(m[449]&m[475]&m[476]&~m[478]&m[479])|(~m[449]&m[475]&m[476]&m[478]&m[479]))&UnbiasedRNG[131])|((m[449]&~m[475]&~m[476]&m[478]&~m[479])|(~m[449]&~m[475]&~m[476]&~m[478]&m[479])|(m[449]&~m[475]&~m[476]&~m[478]&m[479])|(m[449]&m[475]&~m[476]&~m[478]&m[479])|(m[449]&~m[475]&m[476]&~m[478]&m[479])|(~m[449]&~m[475]&~m[476]&m[478]&m[479])|(m[449]&~m[475]&~m[476]&m[478]&m[479])|(~m[449]&m[475]&~m[476]&m[478]&m[479])|(m[449]&m[475]&~m[476]&m[478]&m[479])|(~m[449]&~m[475]&m[476]&m[478]&m[479])|(m[449]&~m[475]&m[476]&m[478]&m[479])|(m[449]&m[475]&m[476]&m[478]&m[479]));
    m[482] = (((m[454]&~m[480]&~m[481]&~m[483]&~m[484])|(~m[454]&~m[480]&~m[481]&m[483]&~m[484])|(m[454]&m[480]&~m[481]&m[483]&~m[484])|(m[454]&~m[480]&m[481]&m[483]&~m[484])|(~m[454]&m[480]&~m[481]&~m[483]&m[484])|(~m[454]&~m[480]&m[481]&~m[483]&m[484])|(m[454]&m[480]&m[481]&~m[483]&m[484])|(~m[454]&m[480]&m[481]&m[483]&m[484]))&UnbiasedRNG[132])|((m[454]&~m[480]&~m[481]&m[483]&~m[484])|(~m[454]&~m[480]&~m[481]&~m[483]&m[484])|(m[454]&~m[480]&~m[481]&~m[483]&m[484])|(m[454]&m[480]&~m[481]&~m[483]&m[484])|(m[454]&~m[480]&m[481]&~m[483]&m[484])|(~m[454]&~m[480]&~m[481]&m[483]&m[484])|(m[454]&~m[480]&~m[481]&m[483]&m[484])|(~m[454]&m[480]&~m[481]&m[483]&m[484])|(m[454]&m[480]&~m[481]&m[483]&m[484])|(~m[454]&~m[480]&m[481]&m[483]&m[484])|(m[454]&~m[480]&m[481]&m[483]&m[484])|(m[454]&m[480]&m[481]&m[483]&m[484]));
    m[487] = (((m[459]&~m[485]&~m[486]&~m[488]&~m[489])|(~m[459]&~m[485]&~m[486]&m[488]&~m[489])|(m[459]&m[485]&~m[486]&m[488]&~m[489])|(m[459]&~m[485]&m[486]&m[488]&~m[489])|(~m[459]&m[485]&~m[486]&~m[488]&m[489])|(~m[459]&~m[485]&m[486]&~m[488]&m[489])|(m[459]&m[485]&m[486]&~m[488]&m[489])|(~m[459]&m[485]&m[486]&m[488]&m[489]))&UnbiasedRNG[133])|((m[459]&~m[485]&~m[486]&m[488]&~m[489])|(~m[459]&~m[485]&~m[486]&~m[488]&m[489])|(m[459]&~m[485]&~m[486]&~m[488]&m[489])|(m[459]&m[485]&~m[486]&~m[488]&m[489])|(m[459]&~m[485]&m[486]&~m[488]&m[489])|(~m[459]&~m[485]&~m[486]&m[488]&m[489])|(m[459]&~m[485]&~m[486]&m[488]&m[489])|(~m[459]&m[485]&~m[486]&m[488]&m[489])|(m[459]&m[485]&~m[486]&m[488]&m[489])|(~m[459]&~m[485]&m[486]&m[488]&m[489])|(m[459]&~m[485]&m[486]&m[488]&m[489])|(m[459]&m[485]&m[486]&m[488]&m[489]));
    m[491] = (((m[321]&~m[490]&~m[492]&~m[493]&~m[494])|(~m[321]&~m[490]&~m[492]&m[493]&~m[494])|(m[321]&m[490]&~m[492]&m[493]&~m[494])|(m[321]&~m[490]&m[492]&m[493]&~m[494])|(~m[321]&m[490]&~m[492]&~m[493]&m[494])|(~m[321]&~m[490]&m[492]&~m[493]&m[494])|(m[321]&m[490]&m[492]&~m[493]&m[494])|(~m[321]&m[490]&m[492]&m[493]&m[494]))&UnbiasedRNG[134])|((m[321]&~m[490]&~m[492]&m[493]&~m[494])|(~m[321]&~m[490]&~m[492]&~m[493]&m[494])|(m[321]&~m[490]&~m[492]&~m[493]&m[494])|(m[321]&m[490]&~m[492]&~m[493]&m[494])|(m[321]&~m[490]&m[492]&~m[493]&m[494])|(~m[321]&~m[490]&~m[492]&m[493]&m[494])|(m[321]&~m[490]&~m[492]&m[493]&m[494])|(~m[321]&m[490]&~m[492]&m[493]&m[494])|(m[321]&m[490]&~m[492]&m[493]&m[494])|(~m[321]&~m[490]&m[492]&m[493]&m[494])|(m[321]&~m[490]&m[492]&m[493]&m[494])|(m[321]&m[490]&m[492]&m[493]&m[494]));
    m[496] = (((m[330]&~m[495]&~m[497]&~m[498]&~m[499])|(~m[330]&~m[495]&~m[497]&m[498]&~m[499])|(m[330]&m[495]&~m[497]&m[498]&~m[499])|(m[330]&~m[495]&m[497]&m[498]&~m[499])|(~m[330]&m[495]&~m[497]&~m[498]&m[499])|(~m[330]&~m[495]&m[497]&~m[498]&m[499])|(m[330]&m[495]&m[497]&~m[498]&m[499])|(~m[330]&m[495]&m[497]&m[498]&m[499]))&UnbiasedRNG[135])|((m[330]&~m[495]&~m[497]&m[498]&~m[499])|(~m[330]&~m[495]&~m[497]&~m[498]&m[499])|(m[330]&~m[495]&~m[497]&~m[498]&m[499])|(m[330]&m[495]&~m[497]&~m[498]&m[499])|(m[330]&~m[495]&m[497]&~m[498]&m[499])|(~m[330]&~m[495]&~m[497]&m[498]&m[499])|(m[330]&~m[495]&~m[497]&m[498]&m[499])|(~m[330]&m[495]&~m[497]&m[498]&m[499])|(m[330]&m[495]&~m[497]&m[498]&m[499])|(~m[330]&~m[495]&m[497]&m[498]&m[499])|(m[330]&~m[495]&m[497]&m[498]&m[499])|(m[330]&m[495]&m[497]&m[498]&m[499]));
    m[501] = (((m[277]&~m[500]&~m[502]&~m[503]&~m[504])|(~m[277]&~m[500]&~m[502]&m[503]&~m[504])|(m[277]&m[500]&~m[502]&m[503]&~m[504])|(m[277]&~m[500]&m[502]&m[503]&~m[504])|(~m[277]&m[500]&~m[502]&~m[503]&m[504])|(~m[277]&~m[500]&m[502]&~m[503]&m[504])|(m[277]&m[500]&m[502]&~m[503]&m[504])|(~m[277]&m[500]&m[502]&m[503]&m[504]))&UnbiasedRNG[136])|((m[277]&~m[500]&~m[502]&m[503]&~m[504])|(~m[277]&~m[500]&~m[502]&~m[503]&m[504])|(m[277]&~m[500]&~m[502]&~m[503]&m[504])|(m[277]&m[500]&~m[502]&~m[503]&m[504])|(m[277]&~m[500]&m[502]&~m[503]&m[504])|(~m[277]&~m[500]&~m[502]&m[503]&m[504])|(m[277]&~m[500]&~m[502]&m[503]&m[504])|(~m[277]&m[500]&~m[502]&m[503]&m[504])|(m[277]&m[500]&~m[502]&m[503]&m[504])|(~m[277]&~m[500]&m[502]&m[503]&m[504])|(m[277]&~m[500]&m[502]&m[503]&m[504])|(m[277]&m[500]&m[502]&m[503]&m[504]));
    m[507] = (((m[474]&~m[505]&~m[506]&~m[508]&~m[509])|(~m[474]&~m[505]&~m[506]&m[508]&~m[509])|(m[474]&m[505]&~m[506]&m[508]&~m[509])|(m[474]&~m[505]&m[506]&m[508]&~m[509])|(~m[474]&m[505]&~m[506]&~m[508]&m[509])|(~m[474]&~m[505]&m[506]&~m[508]&m[509])|(m[474]&m[505]&m[506]&~m[508]&m[509])|(~m[474]&m[505]&m[506]&m[508]&m[509]))&UnbiasedRNG[137])|((m[474]&~m[505]&~m[506]&m[508]&~m[509])|(~m[474]&~m[505]&~m[506]&~m[508]&m[509])|(m[474]&~m[505]&~m[506]&~m[508]&m[509])|(m[474]&m[505]&~m[506]&~m[508]&m[509])|(m[474]&~m[505]&m[506]&~m[508]&m[509])|(~m[474]&~m[505]&~m[506]&m[508]&m[509])|(m[474]&~m[505]&~m[506]&m[508]&m[509])|(~m[474]&m[505]&~m[506]&m[508]&m[509])|(m[474]&m[505]&~m[506]&m[508]&m[509])|(~m[474]&~m[505]&m[506]&m[508]&m[509])|(m[474]&~m[505]&m[506]&m[508]&m[509])|(m[474]&m[505]&m[506]&m[508]&m[509]));
    m[512] = (((m[479]&~m[510]&~m[511]&~m[513]&~m[514])|(~m[479]&~m[510]&~m[511]&m[513]&~m[514])|(m[479]&m[510]&~m[511]&m[513]&~m[514])|(m[479]&~m[510]&m[511]&m[513]&~m[514])|(~m[479]&m[510]&~m[511]&~m[513]&m[514])|(~m[479]&~m[510]&m[511]&~m[513]&m[514])|(m[479]&m[510]&m[511]&~m[513]&m[514])|(~m[479]&m[510]&m[511]&m[513]&m[514]))&UnbiasedRNG[138])|((m[479]&~m[510]&~m[511]&m[513]&~m[514])|(~m[479]&~m[510]&~m[511]&~m[513]&m[514])|(m[479]&~m[510]&~m[511]&~m[513]&m[514])|(m[479]&m[510]&~m[511]&~m[513]&m[514])|(m[479]&~m[510]&m[511]&~m[513]&m[514])|(~m[479]&~m[510]&~m[511]&m[513]&m[514])|(m[479]&~m[510]&~m[511]&m[513]&m[514])|(~m[479]&m[510]&~m[511]&m[513]&m[514])|(m[479]&m[510]&~m[511]&m[513]&m[514])|(~m[479]&~m[510]&m[511]&m[513]&m[514])|(m[479]&~m[510]&m[511]&m[513]&m[514])|(m[479]&m[510]&m[511]&m[513]&m[514]));
    m[517] = (((m[484]&~m[515]&~m[516]&~m[518]&~m[519])|(~m[484]&~m[515]&~m[516]&m[518]&~m[519])|(m[484]&m[515]&~m[516]&m[518]&~m[519])|(m[484]&~m[515]&m[516]&m[518]&~m[519])|(~m[484]&m[515]&~m[516]&~m[518]&m[519])|(~m[484]&~m[515]&m[516]&~m[518]&m[519])|(m[484]&m[515]&m[516]&~m[518]&m[519])|(~m[484]&m[515]&m[516]&m[518]&m[519]))&UnbiasedRNG[139])|((m[484]&~m[515]&~m[516]&m[518]&~m[519])|(~m[484]&~m[515]&~m[516]&~m[518]&m[519])|(m[484]&~m[515]&~m[516]&~m[518]&m[519])|(m[484]&m[515]&~m[516]&~m[518]&m[519])|(m[484]&~m[515]&m[516]&~m[518]&m[519])|(~m[484]&~m[515]&~m[516]&m[518]&m[519])|(m[484]&~m[515]&~m[516]&m[518]&m[519])|(~m[484]&m[515]&~m[516]&m[518]&m[519])|(m[484]&m[515]&~m[516]&m[518]&m[519])|(~m[484]&~m[515]&m[516]&m[518]&m[519])|(m[484]&~m[515]&m[516]&m[518]&m[519])|(m[484]&m[515]&m[516]&m[518]&m[519]));
    m[522] = (((m[489]&~m[520]&~m[521]&~m[523]&~m[524])|(~m[489]&~m[520]&~m[521]&m[523]&~m[524])|(m[489]&m[520]&~m[521]&m[523]&~m[524])|(m[489]&~m[520]&m[521]&m[523]&~m[524])|(~m[489]&m[520]&~m[521]&~m[523]&m[524])|(~m[489]&~m[520]&m[521]&~m[523]&m[524])|(m[489]&m[520]&m[521]&~m[523]&m[524])|(~m[489]&m[520]&m[521]&m[523]&m[524]))&UnbiasedRNG[140])|((m[489]&~m[520]&~m[521]&m[523]&~m[524])|(~m[489]&~m[520]&~m[521]&~m[523]&m[524])|(m[489]&~m[520]&~m[521]&~m[523]&m[524])|(m[489]&m[520]&~m[521]&~m[523]&m[524])|(m[489]&~m[520]&m[521]&~m[523]&m[524])|(~m[489]&~m[520]&~m[521]&m[523]&m[524])|(m[489]&~m[520]&~m[521]&m[523]&m[524])|(~m[489]&m[520]&~m[521]&m[523]&m[524])|(m[489]&m[520]&~m[521]&m[523]&m[524])|(~m[489]&~m[520]&m[521]&m[523]&m[524])|(m[489]&~m[520]&m[521]&m[523]&m[524])|(m[489]&m[520]&m[521]&m[523]&m[524]));
    m[527] = (((m[494]&~m[525]&~m[526]&~m[528]&~m[529])|(~m[494]&~m[525]&~m[526]&m[528]&~m[529])|(m[494]&m[525]&~m[526]&m[528]&~m[529])|(m[494]&~m[525]&m[526]&m[528]&~m[529])|(~m[494]&m[525]&~m[526]&~m[528]&m[529])|(~m[494]&~m[525]&m[526]&~m[528]&m[529])|(m[494]&m[525]&m[526]&~m[528]&m[529])|(~m[494]&m[525]&m[526]&m[528]&m[529]))&UnbiasedRNG[141])|((m[494]&~m[525]&~m[526]&m[528]&~m[529])|(~m[494]&~m[525]&~m[526]&~m[528]&m[529])|(m[494]&~m[525]&~m[526]&~m[528]&m[529])|(m[494]&m[525]&~m[526]&~m[528]&m[529])|(m[494]&~m[525]&m[526]&~m[528]&m[529])|(~m[494]&~m[525]&~m[526]&m[528]&m[529])|(m[494]&~m[525]&~m[526]&m[528]&m[529])|(~m[494]&m[525]&~m[526]&m[528]&m[529])|(m[494]&m[525]&~m[526]&m[528]&m[529])|(~m[494]&~m[525]&m[526]&m[528]&m[529])|(m[494]&~m[525]&m[526]&m[528]&m[529])|(m[494]&m[525]&m[526]&m[528]&m[529]));
    m[531] = (((m[331]&~m[530]&~m[532]&~m[533]&~m[534])|(~m[331]&~m[530]&~m[532]&m[533]&~m[534])|(m[331]&m[530]&~m[532]&m[533]&~m[534])|(m[331]&~m[530]&m[532]&m[533]&~m[534])|(~m[331]&m[530]&~m[532]&~m[533]&m[534])|(~m[331]&~m[530]&m[532]&~m[533]&m[534])|(m[331]&m[530]&m[532]&~m[533]&m[534])|(~m[331]&m[530]&m[532]&m[533]&m[534]))&UnbiasedRNG[142])|((m[331]&~m[530]&~m[532]&m[533]&~m[534])|(~m[331]&~m[530]&~m[532]&~m[533]&m[534])|(m[331]&~m[530]&~m[532]&~m[533]&m[534])|(m[331]&m[530]&~m[532]&~m[533]&m[534])|(m[331]&~m[530]&m[532]&~m[533]&m[534])|(~m[331]&~m[530]&~m[532]&m[533]&m[534])|(m[331]&~m[530]&~m[532]&m[533]&m[534])|(~m[331]&m[530]&~m[532]&m[533]&m[534])|(m[331]&m[530]&~m[532]&m[533]&m[534])|(~m[331]&~m[530]&m[532]&m[533]&m[534])|(m[331]&~m[530]&m[532]&m[533]&m[534])|(m[331]&m[530]&m[532]&m[533]&m[534]));
    m[536] = (((m[340]&~m[535]&~m[537]&~m[538]&~m[539])|(~m[340]&~m[535]&~m[537]&m[538]&~m[539])|(m[340]&m[535]&~m[537]&m[538]&~m[539])|(m[340]&~m[535]&m[537]&m[538]&~m[539])|(~m[340]&m[535]&~m[537]&~m[538]&m[539])|(~m[340]&~m[535]&m[537]&~m[538]&m[539])|(m[340]&m[535]&m[537]&~m[538]&m[539])|(~m[340]&m[535]&m[537]&m[538]&m[539]))&UnbiasedRNG[143])|((m[340]&~m[535]&~m[537]&m[538]&~m[539])|(~m[340]&~m[535]&~m[537]&~m[538]&m[539])|(m[340]&~m[535]&~m[537]&~m[538]&m[539])|(m[340]&m[535]&~m[537]&~m[538]&m[539])|(m[340]&~m[535]&m[537]&~m[538]&m[539])|(~m[340]&~m[535]&~m[537]&m[538]&m[539])|(m[340]&~m[535]&~m[537]&m[538]&m[539])|(~m[340]&m[535]&~m[537]&m[538]&m[539])|(m[340]&m[535]&~m[537]&m[538]&m[539])|(~m[340]&~m[535]&m[537]&m[538]&m[539])|(m[340]&~m[535]&m[537]&m[538]&m[539])|(m[340]&m[535]&m[537]&m[538]&m[539]));
    m[541] = (((m[278]&~m[540]&~m[542]&~m[543]&~m[544])|(~m[278]&~m[540]&~m[542]&m[543]&~m[544])|(m[278]&m[540]&~m[542]&m[543]&~m[544])|(m[278]&~m[540]&m[542]&m[543]&~m[544])|(~m[278]&m[540]&~m[542]&~m[543]&m[544])|(~m[278]&~m[540]&m[542]&~m[543]&m[544])|(m[278]&m[540]&m[542]&~m[543]&m[544])|(~m[278]&m[540]&m[542]&m[543]&m[544]))&UnbiasedRNG[144])|((m[278]&~m[540]&~m[542]&m[543]&~m[544])|(~m[278]&~m[540]&~m[542]&~m[543]&m[544])|(m[278]&~m[540]&~m[542]&~m[543]&m[544])|(m[278]&m[540]&~m[542]&~m[543]&m[544])|(m[278]&~m[540]&m[542]&~m[543]&m[544])|(~m[278]&~m[540]&~m[542]&m[543]&m[544])|(m[278]&~m[540]&~m[542]&m[543]&m[544])|(~m[278]&m[540]&~m[542]&m[543]&m[544])|(m[278]&m[540]&~m[542]&m[543]&m[544])|(~m[278]&~m[540]&m[542]&m[543]&m[544])|(m[278]&~m[540]&m[542]&m[543]&m[544])|(m[278]&m[540]&m[542]&m[543]&m[544]));
    m[547] = (((m[509]&~m[545]&~m[546]&~m[548]&~m[549])|(~m[509]&~m[545]&~m[546]&m[548]&~m[549])|(m[509]&m[545]&~m[546]&m[548]&~m[549])|(m[509]&~m[545]&m[546]&m[548]&~m[549])|(~m[509]&m[545]&~m[546]&~m[548]&m[549])|(~m[509]&~m[545]&m[546]&~m[548]&m[549])|(m[509]&m[545]&m[546]&~m[548]&m[549])|(~m[509]&m[545]&m[546]&m[548]&m[549]))&UnbiasedRNG[145])|((m[509]&~m[545]&~m[546]&m[548]&~m[549])|(~m[509]&~m[545]&~m[546]&~m[548]&m[549])|(m[509]&~m[545]&~m[546]&~m[548]&m[549])|(m[509]&m[545]&~m[546]&~m[548]&m[549])|(m[509]&~m[545]&m[546]&~m[548]&m[549])|(~m[509]&~m[545]&~m[546]&m[548]&m[549])|(m[509]&~m[545]&~m[546]&m[548]&m[549])|(~m[509]&m[545]&~m[546]&m[548]&m[549])|(m[509]&m[545]&~m[546]&m[548]&m[549])|(~m[509]&~m[545]&m[546]&m[548]&m[549])|(m[509]&~m[545]&m[546]&m[548]&m[549])|(m[509]&m[545]&m[546]&m[548]&m[549]));
    m[552] = (((m[514]&~m[550]&~m[551]&~m[553]&~m[554])|(~m[514]&~m[550]&~m[551]&m[553]&~m[554])|(m[514]&m[550]&~m[551]&m[553]&~m[554])|(m[514]&~m[550]&m[551]&m[553]&~m[554])|(~m[514]&m[550]&~m[551]&~m[553]&m[554])|(~m[514]&~m[550]&m[551]&~m[553]&m[554])|(m[514]&m[550]&m[551]&~m[553]&m[554])|(~m[514]&m[550]&m[551]&m[553]&m[554]))&UnbiasedRNG[146])|((m[514]&~m[550]&~m[551]&m[553]&~m[554])|(~m[514]&~m[550]&~m[551]&~m[553]&m[554])|(m[514]&~m[550]&~m[551]&~m[553]&m[554])|(m[514]&m[550]&~m[551]&~m[553]&m[554])|(m[514]&~m[550]&m[551]&~m[553]&m[554])|(~m[514]&~m[550]&~m[551]&m[553]&m[554])|(m[514]&~m[550]&~m[551]&m[553]&m[554])|(~m[514]&m[550]&~m[551]&m[553]&m[554])|(m[514]&m[550]&~m[551]&m[553]&m[554])|(~m[514]&~m[550]&m[551]&m[553]&m[554])|(m[514]&~m[550]&m[551]&m[553]&m[554])|(m[514]&m[550]&m[551]&m[553]&m[554]));
    m[557] = (((m[519]&~m[555]&~m[556]&~m[558]&~m[559])|(~m[519]&~m[555]&~m[556]&m[558]&~m[559])|(m[519]&m[555]&~m[556]&m[558]&~m[559])|(m[519]&~m[555]&m[556]&m[558]&~m[559])|(~m[519]&m[555]&~m[556]&~m[558]&m[559])|(~m[519]&~m[555]&m[556]&~m[558]&m[559])|(m[519]&m[555]&m[556]&~m[558]&m[559])|(~m[519]&m[555]&m[556]&m[558]&m[559]))&UnbiasedRNG[147])|((m[519]&~m[555]&~m[556]&m[558]&~m[559])|(~m[519]&~m[555]&~m[556]&~m[558]&m[559])|(m[519]&~m[555]&~m[556]&~m[558]&m[559])|(m[519]&m[555]&~m[556]&~m[558]&m[559])|(m[519]&~m[555]&m[556]&~m[558]&m[559])|(~m[519]&~m[555]&~m[556]&m[558]&m[559])|(m[519]&~m[555]&~m[556]&m[558]&m[559])|(~m[519]&m[555]&~m[556]&m[558]&m[559])|(m[519]&m[555]&~m[556]&m[558]&m[559])|(~m[519]&~m[555]&m[556]&m[558]&m[559])|(m[519]&~m[555]&m[556]&m[558]&m[559])|(m[519]&m[555]&m[556]&m[558]&m[559]));
    m[562] = (((m[524]&~m[560]&~m[561]&~m[563]&~m[564])|(~m[524]&~m[560]&~m[561]&m[563]&~m[564])|(m[524]&m[560]&~m[561]&m[563]&~m[564])|(m[524]&~m[560]&m[561]&m[563]&~m[564])|(~m[524]&m[560]&~m[561]&~m[563]&m[564])|(~m[524]&~m[560]&m[561]&~m[563]&m[564])|(m[524]&m[560]&m[561]&~m[563]&m[564])|(~m[524]&m[560]&m[561]&m[563]&m[564]))&UnbiasedRNG[148])|((m[524]&~m[560]&~m[561]&m[563]&~m[564])|(~m[524]&~m[560]&~m[561]&~m[563]&m[564])|(m[524]&~m[560]&~m[561]&~m[563]&m[564])|(m[524]&m[560]&~m[561]&~m[563]&m[564])|(m[524]&~m[560]&m[561]&~m[563]&m[564])|(~m[524]&~m[560]&~m[561]&m[563]&m[564])|(m[524]&~m[560]&~m[561]&m[563]&m[564])|(~m[524]&m[560]&~m[561]&m[563]&m[564])|(m[524]&m[560]&~m[561]&m[563]&m[564])|(~m[524]&~m[560]&m[561]&m[563]&m[564])|(m[524]&~m[560]&m[561]&m[563]&m[564])|(m[524]&m[560]&m[561]&m[563]&m[564]));
    m[567] = (((m[529]&~m[565]&~m[566]&~m[568]&~m[569])|(~m[529]&~m[565]&~m[566]&m[568]&~m[569])|(m[529]&m[565]&~m[566]&m[568]&~m[569])|(m[529]&~m[565]&m[566]&m[568]&~m[569])|(~m[529]&m[565]&~m[566]&~m[568]&m[569])|(~m[529]&~m[565]&m[566]&~m[568]&m[569])|(m[529]&m[565]&m[566]&~m[568]&m[569])|(~m[529]&m[565]&m[566]&m[568]&m[569]))&UnbiasedRNG[149])|((m[529]&~m[565]&~m[566]&m[568]&~m[569])|(~m[529]&~m[565]&~m[566]&~m[568]&m[569])|(m[529]&~m[565]&~m[566]&~m[568]&m[569])|(m[529]&m[565]&~m[566]&~m[568]&m[569])|(m[529]&~m[565]&m[566]&~m[568]&m[569])|(~m[529]&~m[565]&~m[566]&m[568]&m[569])|(m[529]&~m[565]&~m[566]&m[568]&m[569])|(~m[529]&m[565]&~m[566]&m[568]&m[569])|(m[529]&m[565]&~m[566]&m[568]&m[569])|(~m[529]&~m[565]&m[566]&m[568]&m[569])|(m[529]&~m[565]&m[566]&m[568]&m[569])|(m[529]&m[565]&m[566]&m[568]&m[569]));
    m[572] = (((m[534]&~m[570]&~m[571]&~m[573]&~m[574])|(~m[534]&~m[570]&~m[571]&m[573]&~m[574])|(m[534]&m[570]&~m[571]&m[573]&~m[574])|(m[534]&~m[570]&m[571]&m[573]&~m[574])|(~m[534]&m[570]&~m[571]&~m[573]&m[574])|(~m[534]&~m[570]&m[571]&~m[573]&m[574])|(m[534]&m[570]&m[571]&~m[573]&m[574])|(~m[534]&m[570]&m[571]&m[573]&m[574]))&UnbiasedRNG[150])|((m[534]&~m[570]&~m[571]&m[573]&~m[574])|(~m[534]&~m[570]&~m[571]&~m[573]&m[574])|(m[534]&~m[570]&~m[571]&~m[573]&m[574])|(m[534]&m[570]&~m[571]&~m[573]&m[574])|(m[534]&~m[570]&m[571]&~m[573]&m[574])|(~m[534]&~m[570]&~m[571]&m[573]&m[574])|(m[534]&~m[570]&~m[571]&m[573]&m[574])|(~m[534]&m[570]&~m[571]&m[573]&m[574])|(m[534]&m[570]&~m[571]&m[573]&m[574])|(~m[534]&~m[570]&m[571]&m[573]&m[574])|(m[534]&~m[570]&m[571]&m[573]&m[574])|(m[534]&m[570]&m[571]&m[573]&m[574]));
    m[576] = (((m[341]&~m[575]&~m[577]&~m[578]&~m[579])|(~m[341]&~m[575]&~m[577]&m[578]&~m[579])|(m[341]&m[575]&~m[577]&m[578]&~m[579])|(m[341]&~m[575]&m[577]&m[578]&~m[579])|(~m[341]&m[575]&~m[577]&~m[578]&m[579])|(~m[341]&~m[575]&m[577]&~m[578]&m[579])|(m[341]&m[575]&m[577]&~m[578]&m[579])|(~m[341]&m[575]&m[577]&m[578]&m[579]))&UnbiasedRNG[151])|((m[341]&~m[575]&~m[577]&m[578]&~m[579])|(~m[341]&~m[575]&~m[577]&~m[578]&m[579])|(m[341]&~m[575]&~m[577]&~m[578]&m[579])|(m[341]&m[575]&~m[577]&~m[578]&m[579])|(m[341]&~m[575]&m[577]&~m[578]&m[579])|(~m[341]&~m[575]&~m[577]&m[578]&m[579])|(m[341]&~m[575]&~m[577]&m[578]&m[579])|(~m[341]&m[575]&~m[577]&m[578]&m[579])|(m[341]&m[575]&~m[577]&m[578]&m[579])|(~m[341]&~m[575]&m[577]&m[578]&m[579])|(m[341]&~m[575]&m[577]&m[578]&m[579])|(m[341]&m[575]&m[577]&m[578]&m[579]));
    m[581] = (((m[350]&~m[580]&~m[582]&~m[583]&~m[584])|(~m[350]&~m[580]&~m[582]&m[583]&~m[584])|(m[350]&m[580]&~m[582]&m[583]&~m[584])|(m[350]&~m[580]&m[582]&m[583]&~m[584])|(~m[350]&m[580]&~m[582]&~m[583]&m[584])|(~m[350]&~m[580]&m[582]&~m[583]&m[584])|(m[350]&m[580]&m[582]&~m[583]&m[584])|(~m[350]&m[580]&m[582]&m[583]&m[584]))&UnbiasedRNG[152])|((m[350]&~m[580]&~m[582]&m[583]&~m[584])|(~m[350]&~m[580]&~m[582]&~m[583]&m[584])|(m[350]&~m[580]&~m[582]&~m[583]&m[584])|(m[350]&m[580]&~m[582]&~m[583]&m[584])|(m[350]&~m[580]&m[582]&~m[583]&m[584])|(~m[350]&~m[580]&~m[582]&m[583]&m[584])|(m[350]&~m[580]&~m[582]&m[583]&m[584])|(~m[350]&m[580]&~m[582]&m[583]&m[584])|(m[350]&m[580]&~m[582]&m[583]&m[584])|(~m[350]&~m[580]&m[582]&m[583]&m[584])|(m[350]&~m[580]&m[582]&m[583]&m[584])|(m[350]&m[580]&m[582]&m[583]&m[584]));
    m[586] = (((m[279]&~m[585]&~m[587]&~m[588]&~m[589])|(~m[279]&~m[585]&~m[587]&m[588]&~m[589])|(m[279]&m[585]&~m[587]&m[588]&~m[589])|(m[279]&~m[585]&m[587]&m[588]&~m[589])|(~m[279]&m[585]&~m[587]&~m[588]&m[589])|(~m[279]&~m[585]&m[587]&~m[588]&m[589])|(m[279]&m[585]&m[587]&~m[588]&m[589])|(~m[279]&m[585]&m[587]&m[588]&m[589]))&UnbiasedRNG[153])|((m[279]&~m[585]&~m[587]&m[588]&~m[589])|(~m[279]&~m[585]&~m[587]&~m[588]&m[589])|(m[279]&~m[585]&~m[587]&~m[588]&m[589])|(m[279]&m[585]&~m[587]&~m[588]&m[589])|(m[279]&~m[585]&m[587]&~m[588]&m[589])|(~m[279]&~m[585]&~m[587]&m[588]&m[589])|(m[279]&~m[585]&~m[587]&m[588]&m[589])|(~m[279]&m[585]&~m[587]&m[588]&m[589])|(m[279]&m[585]&~m[587]&m[588]&m[589])|(~m[279]&~m[585]&m[587]&m[588]&m[589])|(m[279]&~m[585]&m[587]&m[588]&m[589])|(m[279]&m[585]&m[587]&m[588]&m[589]));
    m[592] = (((m[549]&~m[590]&~m[591]&~m[593]&~m[594])|(~m[549]&~m[590]&~m[591]&m[593]&~m[594])|(m[549]&m[590]&~m[591]&m[593]&~m[594])|(m[549]&~m[590]&m[591]&m[593]&~m[594])|(~m[549]&m[590]&~m[591]&~m[593]&m[594])|(~m[549]&~m[590]&m[591]&~m[593]&m[594])|(m[549]&m[590]&m[591]&~m[593]&m[594])|(~m[549]&m[590]&m[591]&m[593]&m[594]))&UnbiasedRNG[154])|((m[549]&~m[590]&~m[591]&m[593]&~m[594])|(~m[549]&~m[590]&~m[591]&~m[593]&m[594])|(m[549]&~m[590]&~m[591]&~m[593]&m[594])|(m[549]&m[590]&~m[591]&~m[593]&m[594])|(m[549]&~m[590]&m[591]&~m[593]&m[594])|(~m[549]&~m[590]&~m[591]&m[593]&m[594])|(m[549]&~m[590]&~m[591]&m[593]&m[594])|(~m[549]&m[590]&~m[591]&m[593]&m[594])|(m[549]&m[590]&~m[591]&m[593]&m[594])|(~m[549]&~m[590]&m[591]&m[593]&m[594])|(m[549]&~m[590]&m[591]&m[593]&m[594])|(m[549]&m[590]&m[591]&m[593]&m[594]));
    m[597] = (((m[554]&~m[595]&~m[596]&~m[598]&~m[599])|(~m[554]&~m[595]&~m[596]&m[598]&~m[599])|(m[554]&m[595]&~m[596]&m[598]&~m[599])|(m[554]&~m[595]&m[596]&m[598]&~m[599])|(~m[554]&m[595]&~m[596]&~m[598]&m[599])|(~m[554]&~m[595]&m[596]&~m[598]&m[599])|(m[554]&m[595]&m[596]&~m[598]&m[599])|(~m[554]&m[595]&m[596]&m[598]&m[599]))&UnbiasedRNG[155])|((m[554]&~m[595]&~m[596]&m[598]&~m[599])|(~m[554]&~m[595]&~m[596]&~m[598]&m[599])|(m[554]&~m[595]&~m[596]&~m[598]&m[599])|(m[554]&m[595]&~m[596]&~m[598]&m[599])|(m[554]&~m[595]&m[596]&~m[598]&m[599])|(~m[554]&~m[595]&~m[596]&m[598]&m[599])|(m[554]&~m[595]&~m[596]&m[598]&m[599])|(~m[554]&m[595]&~m[596]&m[598]&m[599])|(m[554]&m[595]&~m[596]&m[598]&m[599])|(~m[554]&~m[595]&m[596]&m[598]&m[599])|(m[554]&~m[595]&m[596]&m[598]&m[599])|(m[554]&m[595]&m[596]&m[598]&m[599]));
    m[602] = (((m[559]&~m[600]&~m[601]&~m[603]&~m[604])|(~m[559]&~m[600]&~m[601]&m[603]&~m[604])|(m[559]&m[600]&~m[601]&m[603]&~m[604])|(m[559]&~m[600]&m[601]&m[603]&~m[604])|(~m[559]&m[600]&~m[601]&~m[603]&m[604])|(~m[559]&~m[600]&m[601]&~m[603]&m[604])|(m[559]&m[600]&m[601]&~m[603]&m[604])|(~m[559]&m[600]&m[601]&m[603]&m[604]))&UnbiasedRNG[156])|((m[559]&~m[600]&~m[601]&m[603]&~m[604])|(~m[559]&~m[600]&~m[601]&~m[603]&m[604])|(m[559]&~m[600]&~m[601]&~m[603]&m[604])|(m[559]&m[600]&~m[601]&~m[603]&m[604])|(m[559]&~m[600]&m[601]&~m[603]&m[604])|(~m[559]&~m[600]&~m[601]&m[603]&m[604])|(m[559]&~m[600]&~m[601]&m[603]&m[604])|(~m[559]&m[600]&~m[601]&m[603]&m[604])|(m[559]&m[600]&~m[601]&m[603]&m[604])|(~m[559]&~m[600]&m[601]&m[603]&m[604])|(m[559]&~m[600]&m[601]&m[603]&m[604])|(m[559]&m[600]&m[601]&m[603]&m[604]));
    m[607] = (((m[564]&~m[605]&~m[606]&~m[608]&~m[609])|(~m[564]&~m[605]&~m[606]&m[608]&~m[609])|(m[564]&m[605]&~m[606]&m[608]&~m[609])|(m[564]&~m[605]&m[606]&m[608]&~m[609])|(~m[564]&m[605]&~m[606]&~m[608]&m[609])|(~m[564]&~m[605]&m[606]&~m[608]&m[609])|(m[564]&m[605]&m[606]&~m[608]&m[609])|(~m[564]&m[605]&m[606]&m[608]&m[609]))&UnbiasedRNG[157])|((m[564]&~m[605]&~m[606]&m[608]&~m[609])|(~m[564]&~m[605]&~m[606]&~m[608]&m[609])|(m[564]&~m[605]&~m[606]&~m[608]&m[609])|(m[564]&m[605]&~m[606]&~m[608]&m[609])|(m[564]&~m[605]&m[606]&~m[608]&m[609])|(~m[564]&~m[605]&~m[606]&m[608]&m[609])|(m[564]&~m[605]&~m[606]&m[608]&m[609])|(~m[564]&m[605]&~m[606]&m[608]&m[609])|(m[564]&m[605]&~m[606]&m[608]&m[609])|(~m[564]&~m[605]&m[606]&m[608]&m[609])|(m[564]&~m[605]&m[606]&m[608]&m[609])|(m[564]&m[605]&m[606]&m[608]&m[609]));
    m[612] = (((m[569]&~m[610]&~m[611]&~m[613]&~m[614])|(~m[569]&~m[610]&~m[611]&m[613]&~m[614])|(m[569]&m[610]&~m[611]&m[613]&~m[614])|(m[569]&~m[610]&m[611]&m[613]&~m[614])|(~m[569]&m[610]&~m[611]&~m[613]&m[614])|(~m[569]&~m[610]&m[611]&~m[613]&m[614])|(m[569]&m[610]&m[611]&~m[613]&m[614])|(~m[569]&m[610]&m[611]&m[613]&m[614]))&UnbiasedRNG[158])|((m[569]&~m[610]&~m[611]&m[613]&~m[614])|(~m[569]&~m[610]&~m[611]&~m[613]&m[614])|(m[569]&~m[610]&~m[611]&~m[613]&m[614])|(m[569]&m[610]&~m[611]&~m[613]&m[614])|(m[569]&~m[610]&m[611]&~m[613]&m[614])|(~m[569]&~m[610]&~m[611]&m[613]&m[614])|(m[569]&~m[610]&~m[611]&m[613]&m[614])|(~m[569]&m[610]&~m[611]&m[613]&m[614])|(m[569]&m[610]&~m[611]&m[613]&m[614])|(~m[569]&~m[610]&m[611]&m[613]&m[614])|(m[569]&~m[610]&m[611]&m[613]&m[614])|(m[569]&m[610]&m[611]&m[613]&m[614]));
    m[617] = (((m[574]&~m[615]&~m[616]&~m[618]&~m[619])|(~m[574]&~m[615]&~m[616]&m[618]&~m[619])|(m[574]&m[615]&~m[616]&m[618]&~m[619])|(m[574]&~m[615]&m[616]&m[618]&~m[619])|(~m[574]&m[615]&~m[616]&~m[618]&m[619])|(~m[574]&~m[615]&m[616]&~m[618]&m[619])|(m[574]&m[615]&m[616]&~m[618]&m[619])|(~m[574]&m[615]&m[616]&m[618]&m[619]))&UnbiasedRNG[159])|((m[574]&~m[615]&~m[616]&m[618]&~m[619])|(~m[574]&~m[615]&~m[616]&~m[618]&m[619])|(m[574]&~m[615]&~m[616]&~m[618]&m[619])|(m[574]&m[615]&~m[616]&~m[618]&m[619])|(m[574]&~m[615]&m[616]&~m[618]&m[619])|(~m[574]&~m[615]&~m[616]&m[618]&m[619])|(m[574]&~m[615]&~m[616]&m[618]&m[619])|(~m[574]&m[615]&~m[616]&m[618]&m[619])|(m[574]&m[615]&~m[616]&m[618]&m[619])|(~m[574]&~m[615]&m[616]&m[618]&m[619])|(m[574]&~m[615]&m[616]&m[618]&m[619])|(m[574]&m[615]&m[616]&m[618]&m[619]));
    m[622] = (((m[579]&~m[620]&~m[621]&~m[623]&~m[624])|(~m[579]&~m[620]&~m[621]&m[623]&~m[624])|(m[579]&m[620]&~m[621]&m[623]&~m[624])|(m[579]&~m[620]&m[621]&m[623]&~m[624])|(~m[579]&m[620]&~m[621]&~m[623]&m[624])|(~m[579]&~m[620]&m[621]&~m[623]&m[624])|(m[579]&m[620]&m[621]&~m[623]&m[624])|(~m[579]&m[620]&m[621]&m[623]&m[624]))&UnbiasedRNG[160])|((m[579]&~m[620]&~m[621]&m[623]&~m[624])|(~m[579]&~m[620]&~m[621]&~m[623]&m[624])|(m[579]&~m[620]&~m[621]&~m[623]&m[624])|(m[579]&m[620]&~m[621]&~m[623]&m[624])|(m[579]&~m[620]&m[621]&~m[623]&m[624])|(~m[579]&~m[620]&~m[621]&m[623]&m[624])|(m[579]&~m[620]&~m[621]&m[623]&m[624])|(~m[579]&m[620]&~m[621]&m[623]&m[624])|(m[579]&m[620]&~m[621]&m[623]&m[624])|(~m[579]&~m[620]&m[621]&m[623]&m[624])|(m[579]&~m[620]&m[621]&m[623]&m[624])|(m[579]&m[620]&m[621]&m[623]&m[624]));
    m[626] = (((m[351]&~m[625]&~m[627]&~m[628]&~m[629])|(~m[351]&~m[625]&~m[627]&m[628]&~m[629])|(m[351]&m[625]&~m[627]&m[628]&~m[629])|(m[351]&~m[625]&m[627]&m[628]&~m[629])|(~m[351]&m[625]&~m[627]&~m[628]&m[629])|(~m[351]&~m[625]&m[627]&~m[628]&m[629])|(m[351]&m[625]&m[627]&~m[628]&m[629])|(~m[351]&m[625]&m[627]&m[628]&m[629]))&UnbiasedRNG[161])|((m[351]&~m[625]&~m[627]&m[628]&~m[629])|(~m[351]&~m[625]&~m[627]&~m[628]&m[629])|(m[351]&~m[625]&~m[627]&~m[628]&m[629])|(m[351]&m[625]&~m[627]&~m[628]&m[629])|(m[351]&~m[625]&m[627]&~m[628]&m[629])|(~m[351]&~m[625]&~m[627]&m[628]&m[629])|(m[351]&~m[625]&~m[627]&m[628]&m[629])|(~m[351]&m[625]&~m[627]&m[628]&m[629])|(m[351]&m[625]&~m[627]&m[628]&m[629])|(~m[351]&~m[625]&m[627]&m[628]&m[629])|(m[351]&~m[625]&m[627]&m[628]&m[629])|(m[351]&m[625]&m[627]&m[628]&m[629]));
    m[632] = (((m[594]&~m[630]&~m[631]&~m[633]&~m[634])|(~m[594]&~m[630]&~m[631]&m[633]&~m[634])|(m[594]&m[630]&~m[631]&m[633]&~m[634])|(m[594]&~m[630]&m[631]&m[633]&~m[634])|(~m[594]&m[630]&~m[631]&~m[633]&m[634])|(~m[594]&~m[630]&m[631]&~m[633]&m[634])|(m[594]&m[630]&m[631]&~m[633]&m[634])|(~m[594]&m[630]&m[631]&m[633]&m[634]))&UnbiasedRNG[162])|((m[594]&~m[630]&~m[631]&m[633]&~m[634])|(~m[594]&~m[630]&~m[631]&~m[633]&m[634])|(m[594]&~m[630]&~m[631]&~m[633]&m[634])|(m[594]&m[630]&~m[631]&~m[633]&m[634])|(m[594]&~m[630]&m[631]&~m[633]&m[634])|(~m[594]&~m[630]&~m[631]&m[633]&m[634])|(m[594]&~m[630]&~m[631]&m[633]&m[634])|(~m[594]&m[630]&~m[631]&m[633]&m[634])|(m[594]&m[630]&~m[631]&m[633]&m[634])|(~m[594]&~m[630]&m[631]&m[633]&m[634])|(m[594]&~m[630]&m[631]&m[633]&m[634])|(m[594]&m[630]&m[631]&m[633]&m[634]));
    m[637] = (((m[599]&~m[635]&~m[636]&~m[638]&~m[639])|(~m[599]&~m[635]&~m[636]&m[638]&~m[639])|(m[599]&m[635]&~m[636]&m[638]&~m[639])|(m[599]&~m[635]&m[636]&m[638]&~m[639])|(~m[599]&m[635]&~m[636]&~m[638]&m[639])|(~m[599]&~m[635]&m[636]&~m[638]&m[639])|(m[599]&m[635]&m[636]&~m[638]&m[639])|(~m[599]&m[635]&m[636]&m[638]&m[639]))&UnbiasedRNG[163])|((m[599]&~m[635]&~m[636]&m[638]&~m[639])|(~m[599]&~m[635]&~m[636]&~m[638]&m[639])|(m[599]&~m[635]&~m[636]&~m[638]&m[639])|(m[599]&m[635]&~m[636]&~m[638]&m[639])|(m[599]&~m[635]&m[636]&~m[638]&m[639])|(~m[599]&~m[635]&~m[636]&m[638]&m[639])|(m[599]&~m[635]&~m[636]&m[638]&m[639])|(~m[599]&m[635]&~m[636]&m[638]&m[639])|(m[599]&m[635]&~m[636]&m[638]&m[639])|(~m[599]&~m[635]&m[636]&m[638]&m[639])|(m[599]&~m[635]&m[636]&m[638]&m[639])|(m[599]&m[635]&m[636]&m[638]&m[639]));
    m[642] = (((m[604]&~m[640]&~m[641]&~m[643]&~m[644])|(~m[604]&~m[640]&~m[641]&m[643]&~m[644])|(m[604]&m[640]&~m[641]&m[643]&~m[644])|(m[604]&~m[640]&m[641]&m[643]&~m[644])|(~m[604]&m[640]&~m[641]&~m[643]&m[644])|(~m[604]&~m[640]&m[641]&~m[643]&m[644])|(m[604]&m[640]&m[641]&~m[643]&m[644])|(~m[604]&m[640]&m[641]&m[643]&m[644]))&UnbiasedRNG[164])|((m[604]&~m[640]&~m[641]&m[643]&~m[644])|(~m[604]&~m[640]&~m[641]&~m[643]&m[644])|(m[604]&~m[640]&~m[641]&~m[643]&m[644])|(m[604]&m[640]&~m[641]&~m[643]&m[644])|(m[604]&~m[640]&m[641]&~m[643]&m[644])|(~m[604]&~m[640]&~m[641]&m[643]&m[644])|(m[604]&~m[640]&~m[641]&m[643]&m[644])|(~m[604]&m[640]&~m[641]&m[643]&m[644])|(m[604]&m[640]&~m[641]&m[643]&m[644])|(~m[604]&~m[640]&m[641]&m[643]&m[644])|(m[604]&~m[640]&m[641]&m[643]&m[644])|(m[604]&m[640]&m[641]&m[643]&m[644]));
    m[647] = (((m[609]&~m[645]&~m[646]&~m[648]&~m[649])|(~m[609]&~m[645]&~m[646]&m[648]&~m[649])|(m[609]&m[645]&~m[646]&m[648]&~m[649])|(m[609]&~m[645]&m[646]&m[648]&~m[649])|(~m[609]&m[645]&~m[646]&~m[648]&m[649])|(~m[609]&~m[645]&m[646]&~m[648]&m[649])|(m[609]&m[645]&m[646]&~m[648]&m[649])|(~m[609]&m[645]&m[646]&m[648]&m[649]))&UnbiasedRNG[165])|((m[609]&~m[645]&~m[646]&m[648]&~m[649])|(~m[609]&~m[645]&~m[646]&~m[648]&m[649])|(m[609]&~m[645]&~m[646]&~m[648]&m[649])|(m[609]&m[645]&~m[646]&~m[648]&m[649])|(m[609]&~m[645]&m[646]&~m[648]&m[649])|(~m[609]&~m[645]&~m[646]&m[648]&m[649])|(m[609]&~m[645]&~m[646]&m[648]&m[649])|(~m[609]&m[645]&~m[646]&m[648]&m[649])|(m[609]&m[645]&~m[646]&m[648]&m[649])|(~m[609]&~m[645]&m[646]&m[648]&m[649])|(m[609]&~m[645]&m[646]&m[648]&m[649])|(m[609]&m[645]&m[646]&m[648]&m[649]));
    m[652] = (((m[614]&~m[650]&~m[651]&~m[653]&~m[654])|(~m[614]&~m[650]&~m[651]&m[653]&~m[654])|(m[614]&m[650]&~m[651]&m[653]&~m[654])|(m[614]&~m[650]&m[651]&m[653]&~m[654])|(~m[614]&m[650]&~m[651]&~m[653]&m[654])|(~m[614]&~m[650]&m[651]&~m[653]&m[654])|(m[614]&m[650]&m[651]&~m[653]&m[654])|(~m[614]&m[650]&m[651]&m[653]&m[654]))&UnbiasedRNG[166])|((m[614]&~m[650]&~m[651]&m[653]&~m[654])|(~m[614]&~m[650]&~m[651]&~m[653]&m[654])|(m[614]&~m[650]&~m[651]&~m[653]&m[654])|(m[614]&m[650]&~m[651]&~m[653]&m[654])|(m[614]&~m[650]&m[651]&~m[653]&m[654])|(~m[614]&~m[650]&~m[651]&m[653]&m[654])|(m[614]&~m[650]&~m[651]&m[653]&m[654])|(~m[614]&m[650]&~m[651]&m[653]&m[654])|(m[614]&m[650]&~m[651]&m[653]&m[654])|(~m[614]&~m[650]&m[651]&m[653]&m[654])|(m[614]&~m[650]&m[651]&m[653]&m[654])|(m[614]&m[650]&m[651]&m[653]&m[654]));
    m[657] = (((m[619]&~m[655]&~m[656]&~m[658]&~m[659])|(~m[619]&~m[655]&~m[656]&m[658]&~m[659])|(m[619]&m[655]&~m[656]&m[658]&~m[659])|(m[619]&~m[655]&m[656]&m[658]&~m[659])|(~m[619]&m[655]&~m[656]&~m[658]&m[659])|(~m[619]&~m[655]&m[656]&~m[658]&m[659])|(m[619]&m[655]&m[656]&~m[658]&m[659])|(~m[619]&m[655]&m[656]&m[658]&m[659]))&UnbiasedRNG[167])|((m[619]&~m[655]&~m[656]&m[658]&~m[659])|(~m[619]&~m[655]&~m[656]&~m[658]&m[659])|(m[619]&~m[655]&~m[656]&~m[658]&m[659])|(m[619]&m[655]&~m[656]&~m[658]&m[659])|(m[619]&~m[655]&m[656]&~m[658]&m[659])|(~m[619]&~m[655]&~m[656]&m[658]&m[659])|(m[619]&~m[655]&~m[656]&m[658]&m[659])|(~m[619]&m[655]&~m[656]&m[658]&m[659])|(m[619]&m[655]&~m[656]&m[658]&m[659])|(~m[619]&~m[655]&m[656]&m[658]&m[659])|(m[619]&~m[655]&m[656]&m[658]&m[659])|(m[619]&m[655]&m[656]&m[658]&m[659]));
    m[662] = (((m[624]&~m[660]&~m[661]&~m[663]&~m[664])|(~m[624]&~m[660]&~m[661]&m[663]&~m[664])|(m[624]&m[660]&~m[661]&m[663]&~m[664])|(m[624]&~m[660]&m[661]&m[663]&~m[664])|(~m[624]&m[660]&~m[661]&~m[663]&m[664])|(~m[624]&~m[660]&m[661]&~m[663]&m[664])|(m[624]&m[660]&m[661]&~m[663]&m[664])|(~m[624]&m[660]&m[661]&m[663]&m[664]))&UnbiasedRNG[168])|((m[624]&~m[660]&~m[661]&m[663]&~m[664])|(~m[624]&~m[660]&~m[661]&~m[663]&m[664])|(m[624]&~m[660]&~m[661]&~m[663]&m[664])|(m[624]&m[660]&~m[661]&~m[663]&m[664])|(m[624]&~m[660]&m[661]&~m[663]&m[664])|(~m[624]&~m[660]&~m[661]&m[663]&m[664])|(m[624]&~m[660]&~m[661]&m[663]&m[664])|(~m[624]&m[660]&~m[661]&m[663]&m[664])|(m[624]&m[660]&~m[661]&m[663]&m[664])|(~m[624]&~m[660]&m[661]&m[663]&m[664])|(m[624]&~m[660]&m[661]&m[663]&m[664])|(m[624]&m[660]&m[661]&m[663]&m[664]));
    m[667] = (((m[629]&~m[665]&~m[666]&~m[668]&~m[669])|(~m[629]&~m[665]&~m[666]&m[668]&~m[669])|(m[629]&m[665]&~m[666]&m[668]&~m[669])|(m[629]&~m[665]&m[666]&m[668]&~m[669])|(~m[629]&m[665]&~m[666]&~m[668]&m[669])|(~m[629]&~m[665]&m[666]&~m[668]&m[669])|(m[629]&m[665]&m[666]&~m[668]&m[669])|(~m[629]&m[665]&m[666]&m[668]&m[669]))&UnbiasedRNG[169])|((m[629]&~m[665]&~m[666]&m[668]&~m[669])|(~m[629]&~m[665]&~m[666]&~m[668]&m[669])|(m[629]&~m[665]&~m[666]&~m[668]&m[669])|(m[629]&m[665]&~m[666]&~m[668]&m[669])|(m[629]&~m[665]&m[666]&~m[668]&m[669])|(~m[629]&~m[665]&~m[666]&m[668]&m[669])|(m[629]&~m[665]&~m[666]&m[668]&m[669])|(~m[629]&m[665]&~m[666]&m[668]&m[669])|(m[629]&m[665]&~m[666]&m[668]&m[669])|(~m[629]&~m[665]&m[666]&m[668]&m[669])|(m[629]&~m[665]&m[666]&m[668]&m[669])|(m[629]&m[665]&m[666]&m[668]&m[669]));
    m[672] = (((m[639]&~m[670]&~m[671]&~m[673]&~m[674])|(~m[639]&~m[670]&~m[671]&m[673]&~m[674])|(m[639]&m[670]&~m[671]&m[673]&~m[674])|(m[639]&~m[670]&m[671]&m[673]&~m[674])|(~m[639]&m[670]&~m[671]&~m[673]&m[674])|(~m[639]&~m[670]&m[671]&~m[673]&m[674])|(m[639]&m[670]&m[671]&~m[673]&m[674])|(~m[639]&m[670]&m[671]&m[673]&m[674]))&UnbiasedRNG[170])|((m[639]&~m[670]&~m[671]&m[673]&~m[674])|(~m[639]&~m[670]&~m[671]&~m[673]&m[674])|(m[639]&~m[670]&~m[671]&~m[673]&m[674])|(m[639]&m[670]&~m[671]&~m[673]&m[674])|(m[639]&~m[670]&m[671]&~m[673]&m[674])|(~m[639]&~m[670]&~m[671]&m[673]&m[674])|(m[639]&~m[670]&~m[671]&m[673]&m[674])|(~m[639]&m[670]&~m[671]&m[673]&m[674])|(m[639]&m[670]&~m[671]&m[673]&m[674])|(~m[639]&~m[670]&m[671]&m[673]&m[674])|(m[639]&~m[670]&m[671]&m[673]&m[674])|(m[639]&m[670]&m[671]&m[673]&m[674]));
    m[677] = (((m[644]&~m[675]&~m[676]&~m[678]&~m[679])|(~m[644]&~m[675]&~m[676]&m[678]&~m[679])|(m[644]&m[675]&~m[676]&m[678]&~m[679])|(m[644]&~m[675]&m[676]&m[678]&~m[679])|(~m[644]&m[675]&~m[676]&~m[678]&m[679])|(~m[644]&~m[675]&m[676]&~m[678]&m[679])|(m[644]&m[675]&m[676]&~m[678]&m[679])|(~m[644]&m[675]&m[676]&m[678]&m[679]))&UnbiasedRNG[171])|((m[644]&~m[675]&~m[676]&m[678]&~m[679])|(~m[644]&~m[675]&~m[676]&~m[678]&m[679])|(m[644]&~m[675]&~m[676]&~m[678]&m[679])|(m[644]&m[675]&~m[676]&~m[678]&m[679])|(m[644]&~m[675]&m[676]&~m[678]&m[679])|(~m[644]&~m[675]&~m[676]&m[678]&m[679])|(m[644]&~m[675]&~m[676]&m[678]&m[679])|(~m[644]&m[675]&~m[676]&m[678]&m[679])|(m[644]&m[675]&~m[676]&m[678]&m[679])|(~m[644]&~m[675]&m[676]&m[678]&m[679])|(m[644]&~m[675]&m[676]&m[678]&m[679])|(m[644]&m[675]&m[676]&m[678]&m[679]));
    m[682] = (((m[649]&~m[680]&~m[681]&~m[683]&~m[684])|(~m[649]&~m[680]&~m[681]&m[683]&~m[684])|(m[649]&m[680]&~m[681]&m[683]&~m[684])|(m[649]&~m[680]&m[681]&m[683]&~m[684])|(~m[649]&m[680]&~m[681]&~m[683]&m[684])|(~m[649]&~m[680]&m[681]&~m[683]&m[684])|(m[649]&m[680]&m[681]&~m[683]&m[684])|(~m[649]&m[680]&m[681]&m[683]&m[684]))&UnbiasedRNG[172])|((m[649]&~m[680]&~m[681]&m[683]&~m[684])|(~m[649]&~m[680]&~m[681]&~m[683]&m[684])|(m[649]&~m[680]&~m[681]&~m[683]&m[684])|(m[649]&m[680]&~m[681]&~m[683]&m[684])|(m[649]&~m[680]&m[681]&~m[683]&m[684])|(~m[649]&~m[680]&~m[681]&m[683]&m[684])|(m[649]&~m[680]&~m[681]&m[683]&m[684])|(~m[649]&m[680]&~m[681]&m[683]&m[684])|(m[649]&m[680]&~m[681]&m[683]&m[684])|(~m[649]&~m[680]&m[681]&m[683]&m[684])|(m[649]&~m[680]&m[681]&m[683]&m[684])|(m[649]&m[680]&m[681]&m[683]&m[684]));
    m[687] = (((m[654]&~m[685]&~m[686]&~m[688]&~m[689])|(~m[654]&~m[685]&~m[686]&m[688]&~m[689])|(m[654]&m[685]&~m[686]&m[688]&~m[689])|(m[654]&~m[685]&m[686]&m[688]&~m[689])|(~m[654]&m[685]&~m[686]&~m[688]&m[689])|(~m[654]&~m[685]&m[686]&~m[688]&m[689])|(m[654]&m[685]&m[686]&~m[688]&m[689])|(~m[654]&m[685]&m[686]&m[688]&m[689]))&UnbiasedRNG[173])|((m[654]&~m[685]&~m[686]&m[688]&~m[689])|(~m[654]&~m[685]&~m[686]&~m[688]&m[689])|(m[654]&~m[685]&~m[686]&~m[688]&m[689])|(m[654]&m[685]&~m[686]&~m[688]&m[689])|(m[654]&~m[685]&m[686]&~m[688]&m[689])|(~m[654]&~m[685]&~m[686]&m[688]&m[689])|(m[654]&~m[685]&~m[686]&m[688]&m[689])|(~m[654]&m[685]&~m[686]&m[688]&m[689])|(m[654]&m[685]&~m[686]&m[688]&m[689])|(~m[654]&~m[685]&m[686]&m[688]&m[689])|(m[654]&~m[685]&m[686]&m[688]&m[689])|(m[654]&m[685]&m[686]&m[688]&m[689]));
    m[692] = (((m[659]&~m[690]&~m[691]&~m[693]&~m[694])|(~m[659]&~m[690]&~m[691]&m[693]&~m[694])|(m[659]&m[690]&~m[691]&m[693]&~m[694])|(m[659]&~m[690]&m[691]&m[693]&~m[694])|(~m[659]&m[690]&~m[691]&~m[693]&m[694])|(~m[659]&~m[690]&m[691]&~m[693]&m[694])|(m[659]&m[690]&m[691]&~m[693]&m[694])|(~m[659]&m[690]&m[691]&m[693]&m[694]))&UnbiasedRNG[174])|((m[659]&~m[690]&~m[691]&m[693]&~m[694])|(~m[659]&~m[690]&~m[691]&~m[693]&m[694])|(m[659]&~m[690]&~m[691]&~m[693]&m[694])|(m[659]&m[690]&~m[691]&~m[693]&m[694])|(m[659]&~m[690]&m[691]&~m[693]&m[694])|(~m[659]&~m[690]&~m[691]&m[693]&m[694])|(m[659]&~m[690]&~m[691]&m[693]&m[694])|(~m[659]&m[690]&~m[691]&m[693]&m[694])|(m[659]&m[690]&~m[691]&m[693]&m[694])|(~m[659]&~m[690]&m[691]&m[693]&m[694])|(m[659]&~m[690]&m[691]&m[693]&m[694])|(m[659]&m[690]&m[691]&m[693]&m[694]));
    m[697] = (((m[664]&~m[695]&~m[696]&~m[698]&~m[699])|(~m[664]&~m[695]&~m[696]&m[698]&~m[699])|(m[664]&m[695]&~m[696]&m[698]&~m[699])|(m[664]&~m[695]&m[696]&m[698]&~m[699])|(~m[664]&m[695]&~m[696]&~m[698]&m[699])|(~m[664]&~m[695]&m[696]&~m[698]&m[699])|(m[664]&m[695]&m[696]&~m[698]&m[699])|(~m[664]&m[695]&m[696]&m[698]&m[699]))&UnbiasedRNG[175])|((m[664]&~m[695]&~m[696]&m[698]&~m[699])|(~m[664]&~m[695]&~m[696]&~m[698]&m[699])|(m[664]&~m[695]&~m[696]&~m[698]&m[699])|(m[664]&m[695]&~m[696]&~m[698]&m[699])|(m[664]&~m[695]&m[696]&~m[698]&m[699])|(~m[664]&~m[695]&~m[696]&m[698]&m[699])|(m[664]&~m[695]&~m[696]&m[698]&m[699])|(~m[664]&m[695]&~m[696]&m[698]&m[699])|(m[664]&m[695]&~m[696]&m[698]&m[699])|(~m[664]&~m[695]&m[696]&m[698]&m[699])|(m[664]&~m[695]&m[696]&m[698]&m[699])|(m[664]&m[695]&m[696]&m[698]&m[699]));
    m[702] = (((m[669]&~m[700]&~m[701]&~m[703]&~m[704])|(~m[669]&~m[700]&~m[701]&m[703]&~m[704])|(m[669]&m[700]&~m[701]&m[703]&~m[704])|(m[669]&~m[700]&m[701]&m[703]&~m[704])|(~m[669]&m[700]&~m[701]&~m[703]&m[704])|(~m[669]&~m[700]&m[701]&~m[703]&m[704])|(m[669]&m[700]&m[701]&~m[703]&m[704])|(~m[669]&m[700]&m[701]&m[703]&m[704]))&UnbiasedRNG[176])|((m[669]&~m[700]&~m[701]&m[703]&~m[704])|(~m[669]&~m[700]&~m[701]&~m[703]&m[704])|(m[669]&~m[700]&~m[701]&~m[703]&m[704])|(m[669]&m[700]&~m[701]&~m[703]&m[704])|(m[669]&~m[700]&m[701]&~m[703]&m[704])|(~m[669]&~m[700]&~m[701]&m[703]&m[704])|(m[669]&~m[700]&~m[701]&m[703]&m[704])|(~m[669]&m[700]&~m[701]&m[703]&m[704])|(m[669]&m[700]&~m[701]&m[703]&m[704])|(~m[669]&~m[700]&m[701]&m[703]&m[704])|(m[669]&~m[700]&m[701]&m[703]&m[704])|(m[669]&m[700]&m[701]&m[703]&m[704]));
    m[707] = (((m[679]&~m[705]&~m[706]&~m[708]&~m[709])|(~m[679]&~m[705]&~m[706]&m[708]&~m[709])|(m[679]&m[705]&~m[706]&m[708]&~m[709])|(m[679]&~m[705]&m[706]&m[708]&~m[709])|(~m[679]&m[705]&~m[706]&~m[708]&m[709])|(~m[679]&~m[705]&m[706]&~m[708]&m[709])|(m[679]&m[705]&m[706]&~m[708]&m[709])|(~m[679]&m[705]&m[706]&m[708]&m[709]))&UnbiasedRNG[177])|((m[679]&~m[705]&~m[706]&m[708]&~m[709])|(~m[679]&~m[705]&~m[706]&~m[708]&m[709])|(m[679]&~m[705]&~m[706]&~m[708]&m[709])|(m[679]&m[705]&~m[706]&~m[708]&m[709])|(m[679]&~m[705]&m[706]&~m[708]&m[709])|(~m[679]&~m[705]&~m[706]&m[708]&m[709])|(m[679]&~m[705]&~m[706]&m[708]&m[709])|(~m[679]&m[705]&~m[706]&m[708]&m[709])|(m[679]&m[705]&~m[706]&m[708]&m[709])|(~m[679]&~m[705]&m[706]&m[708]&m[709])|(m[679]&~m[705]&m[706]&m[708]&m[709])|(m[679]&m[705]&m[706]&m[708]&m[709]));
    m[712] = (((m[684]&~m[710]&~m[711]&~m[713]&~m[714])|(~m[684]&~m[710]&~m[711]&m[713]&~m[714])|(m[684]&m[710]&~m[711]&m[713]&~m[714])|(m[684]&~m[710]&m[711]&m[713]&~m[714])|(~m[684]&m[710]&~m[711]&~m[713]&m[714])|(~m[684]&~m[710]&m[711]&~m[713]&m[714])|(m[684]&m[710]&m[711]&~m[713]&m[714])|(~m[684]&m[710]&m[711]&m[713]&m[714]))&UnbiasedRNG[178])|((m[684]&~m[710]&~m[711]&m[713]&~m[714])|(~m[684]&~m[710]&~m[711]&~m[713]&m[714])|(m[684]&~m[710]&~m[711]&~m[713]&m[714])|(m[684]&m[710]&~m[711]&~m[713]&m[714])|(m[684]&~m[710]&m[711]&~m[713]&m[714])|(~m[684]&~m[710]&~m[711]&m[713]&m[714])|(m[684]&~m[710]&~m[711]&m[713]&m[714])|(~m[684]&m[710]&~m[711]&m[713]&m[714])|(m[684]&m[710]&~m[711]&m[713]&m[714])|(~m[684]&~m[710]&m[711]&m[713]&m[714])|(m[684]&~m[710]&m[711]&m[713]&m[714])|(m[684]&m[710]&m[711]&m[713]&m[714]));
    m[717] = (((m[689]&~m[715]&~m[716]&~m[718]&~m[719])|(~m[689]&~m[715]&~m[716]&m[718]&~m[719])|(m[689]&m[715]&~m[716]&m[718]&~m[719])|(m[689]&~m[715]&m[716]&m[718]&~m[719])|(~m[689]&m[715]&~m[716]&~m[718]&m[719])|(~m[689]&~m[715]&m[716]&~m[718]&m[719])|(m[689]&m[715]&m[716]&~m[718]&m[719])|(~m[689]&m[715]&m[716]&m[718]&m[719]))&UnbiasedRNG[179])|((m[689]&~m[715]&~m[716]&m[718]&~m[719])|(~m[689]&~m[715]&~m[716]&~m[718]&m[719])|(m[689]&~m[715]&~m[716]&~m[718]&m[719])|(m[689]&m[715]&~m[716]&~m[718]&m[719])|(m[689]&~m[715]&m[716]&~m[718]&m[719])|(~m[689]&~m[715]&~m[716]&m[718]&m[719])|(m[689]&~m[715]&~m[716]&m[718]&m[719])|(~m[689]&m[715]&~m[716]&m[718]&m[719])|(m[689]&m[715]&~m[716]&m[718]&m[719])|(~m[689]&~m[715]&m[716]&m[718]&m[719])|(m[689]&~m[715]&m[716]&m[718]&m[719])|(m[689]&m[715]&m[716]&m[718]&m[719]));
    m[722] = (((m[694]&~m[720]&~m[721]&~m[723]&~m[724])|(~m[694]&~m[720]&~m[721]&m[723]&~m[724])|(m[694]&m[720]&~m[721]&m[723]&~m[724])|(m[694]&~m[720]&m[721]&m[723]&~m[724])|(~m[694]&m[720]&~m[721]&~m[723]&m[724])|(~m[694]&~m[720]&m[721]&~m[723]&m[724])|(m[694]&m[720]&m[721]&~m[723]&m[724])|(~m[694]&m[720]&m[721]&m[723]&m[724]))&UnbiasedRNG[180])|((m[694]&~m[720]&~m[721]&m[723]&~m[724])|(~m[694]&~m[720]&~m[721]&~m[723]&m[724])|(m[694]&~m[720]&~m[721]&~m[723]&m[724])|(m[694]&m[720]&~m[721]&~m[723]&m[724])|(m[694]&~m[720]&m[721]&~m[723]&m[724])|(~m[694]&~m[720]&~m[721]&m[723]&m[724])|(m[694]&~m[720]&~m[721]&m[723]&m[724])|(~m[694]&m[720]&~m[721]&m[723]&m[724])|(m[694]&m[720]&~m[721]&m[723]&m[724])|(~m[694]&~m[720]&m[721]&m[723]&m[724])|(m[694]&~m[720]&m[721]&m[723]&m[724])|(m[694]&m[720]&m[721]&m[723]&m[724]));
    m[727] = (((m[699]&~m[725]&~m[726]&~m[728]&~m[729])|(~m[699]&~m[725]&~m[726]&m[728]&~m[729])|(m[699]&m[725]&~m[726]&m[728]&~m[729])|(m[699]&~m[725]&m[726]&m[728]&~m[729])|(~m[699]&m[725]&~m[726]&~m[728]&m[729])|(~m[699]&~m[725]&m[726]&~m[728]&m[729])|(m[699]&m[725]&m[726]&~m[728]&m[729])|(~m[699]&m[725]&m[726]&m[728]&m[729]))&UnbiasedRNG[181])|((m[699]&~m[725]&~m[726]&m[728]&~m[729])|(~m[699]&~m[725]&~m[726]&~m[728]&m[729])|(m[699]&~m[725]&~m[726]&~m[728]&m[729])|(m[699]&m[725]&~m[726]&~m[728]&m[729])|(m[699]&~m[725]&m[726]&~m[728]&m[729])|(~m[699]&~m[725]&~m[726]&m[728]&m[729])|(m[699]&~m[725]&~m[726]&m[728]&m[729])|(~m[699]&m[725]&~m[726]&m[728]&m[729])|(m[699]&m[725]&~m[726]&m[728]&m[729])|(~m[699]&~m[725]&m[726]&m[728]&m[729])|(m[699]&~m[725]&m[726]&m[728]&m[729])|(m[699]&m[725]&m[726]&m[728]&m[729]));
    m[732] = (((m[704]&~m[730]&~m[731]&~m[733]&~m[734])|(~m[704]&~m[730]&~m[731]&m[733]&~m[734])|(m[704]&m[730]&~m[731]&m[733]&~m[734])|(m[704]&~m[730]&m[731]&m[733]&~m[734])|(~m[704]&m[730]&~m[731]&~m[733]&m[734])|(~m[704]&~m[730]&m[731]&~m[733]&m[734])|(m[704]&m[730]&m[731]&~m[733]&m[734])|(~m[704]&m[730]&m[731]&m[733]&m[734]))&UnbiasedRNG[182])|((m[704]&~m[730]&~m[731]&m[733]&~m[734])|(~m[704]&~m[730]&~m[731]&~m[733]&m[734])|(m[704]&~m[730]&~m[731]&~m[733]&m[734])|(m[704]&m[730]&~m[731]&~m[733]&m[734])|(m[704]&~m[730]&m[731]&~m[733]&m[734])|(~m[704]&~m[730]&~m[731]&m[733]&m[734])|(m[704]&~m[730]&~m[731]&m[733]&m[734])|(~m[704]&m[730]&~m[731]&m[733]&m[734])|(m[704]&m[730]&~m[731]&m[733]&m[734])|(~m[704]&~m[730]&m[731]&m[733]&m[734])|(m[704]&~m[730]&m[731]&m[733]&m[734])|(m[704]&m[730]&m[731]&m[733]&m[734]));
    m[737] = (((m[714]&~m[735]&~m[736]&~m[738]&~m[739])|(~m[714]&~m[735]&~m[736]&m[738]&~m[739])|(m[714]&m[735]&~m[736]&m[738]&~m[739])|(m[714]&~m[735]&m[736]&m[738]&~m[739])|(~m[714]&m[735]&~m[736]&~m[738]&m[739])|(~m[714]&~m[735]&m[736]&~m[738]&m[739])|(m[714]&m[735]&m[736]&~m[738]&m[739])|(~m[714]&m[735]&m[736]&m[738]&m[739]))&UnbiasedRNG[183])|((m[714]&~m[735]&~m[736]&m[738]&~m[739])|(~m[714]&~m[735]&~m[736]&~m[738]&m[739])|(m[714]&~m[735]&~m[736]&~m[738]&m[739])|(m[714]&m[735]&~m[736]&~m[738]&m[739])|(m[714]&~m[735]&m[736]&~m[738]&m[739])|(~m[714]&~m[735]&~m[736]&m[738]&m[739])|(m[714]&~m[735]&~m[736]&m[738]&m[739])|(~m[714]&m[735]&~m[736]&m[738]&m[739])|(m[714]&m[735]&~m[736]&m[738]&m[739])|(~m[714]&~m[735]&m[736]&m[738]&m[739])|(m[714]&~m[735]&m[736]&m[738]&m[739])|(m[714]&m[735]&m[736]&m[738]&m[739]));
    m[742] = (((m[719]&~m[740]&~m[741]&~m[743]&~m[744])|(~m[719]&~m[740]&~m[741]&m[743]&~m[744])|(m[719]&m[740]&~m[741]&m[743]&~m[744])|(m[719]&~m[740]&m[741]&m[743]&~m[744])|(~m[719]&m[740]&~m[741]&~m[743]&m[744])|(~m[719]&~m[740]&m[741]&~m[743]&m[744])|(m[719]&m[740]&m[741]&~m[743]&m[744])|(~m[719]&m[740]&m[741]&m[743]&m[744]))&UnbiasedRNG[184])|((m[719]&~m[740]&~m[741]&m[743]&~m[744])|(~m[719]&~m[740]&~m[741]&~m[743]&m[744])|(m[719]&~m[740]&~m[741]&~m[743]&m[744])|(m[719]&m[740]&~m[741]&~m[743]&m[744])|(m[719]&~m[740]&m[741]&~m[743]&m[744])|(~m[719]&~m[740]&~m[741]&m[743]&m[744])|(m[719]&~m[740]&~m[741]&m[743]&m[744])|(~m[719]&m[740]&~m[741]&m[743]&m[744])|(m[719]&m[740]&~m[741]&m[743]&m[744])|(~m[719]&~m[740]&m[741]&m[743]&m[744])|(m[719]&~m[740]&m[741]&m[743]&m[744])|(m[719]&m[740]&m[741]&m[743]&m[744]));
    m[747] = (((m[724]&~m[745]&~m[746]&~m[748]&~m[749])|(~m[724]&~m[745]&~m[746]&m[748]&~m[749])|(m[724]&m[745]&~m[746]&m[748]&~m[749])|(m[724]&~m[745]&m[746]&m[748]&~m[749])|(~m[724]&m[745]&~m[746]&~m[748]&m[749])|(~m[724]&~m[745]&m[746]&~m[748]&m[749])|(m[724]&m[745]&m[746]&~m[748]&m[749])|(~m[724]&m[745]&m[746]&m[748]&m[749]))&UnbiasedRNG[185])|((m[724]&~m[745]&~m[746]&m[748]&~m[749])|(~m[724]&~m[745]&~m[746]&~m[748]&m[749])|(m[724]&~m[745]&~m[746]&~m[748]&m[749])|(m[724]&m[745]&~m[746]&~m[748]&m[749])|(m[724]&~m[745]&m[746]&~m[748]&m[749])|(~m[724]&~m[745]&~m[746]&m[748]&m[749])|(m[724]&~m[745]&~m[746]&m[748]&m[749])|(~m[724]&m[745]&~m[746]&m[748]&m[749])|(m[724]&m[745]&~m[746]&m[748]&m[749])|(~m[724]&~m[745]&m[746]&m[748]&m[749])|(m[724]&~m[745]&m[746]&m[748]&m[749])|(m[724]&m[745]&m[746]&m[748]&m[749]));
    m[752] = (((m[729]&~m[750]&~m[751]&~m[753]&~m[754])|(~m[729]&~m[750]&~m[751]&m[753]&~m[754])|(m[729]&m[750]&~m[751]&m[753]&~m[754])|(m[729]&~m[750]&m[751]&m[753]&~m[754])|(~m[729]&m[750]&~m[751]&~m[753]&m[754])|(~m[729]&~m[750]&m[751]&~m[753]&m[754])|(m[729]&m[750]&m[751]&~m[753]&m[754])|(~m[729]&m[750]&m[751]&m[753]&m[754]))&UnbiasedRNG[186])|((m[729]&~m[750]&~m[751]&m[753]&~m[754])|(~m[729]&~m[750]&~m[751]&~m[753]&m[754])|(m[729]&~m[750]&~m[751]&~m[753]&m[754])|(m[729]&m[750]&~m[751]&~m[753]&m[754])|(m[729]&~m[750]&m[751]&~m[753]&m[754])|(~m[729]&~m[750]&~m[751]&m[753]&m[754])|(m[729]&~m[750]&~m[751]&m[753]&m[754])|(~m[729]&m[750]&~m[751]&m[753]&m[754])|(m[729]&m[750]&~m[751]&m[753]&m[754])|(~m[729]&~m[750]&m[751]&m[753]&m[754])|(m[729]&~m[750]&m[751]&m[753]&m[754])|(m[729]&m[750]&m[751]&m[753]&m[754]));
    m[757] = (((m[734]&~m[755]&~m[756]&~m[758]&~m[759])|(~m[734]&~m[755]&~m[756]&m[758]&~m[759])|(m[734]&m[755]&~m[756]&m[758]&~m[759])|(m[734]&~m[755]&m[756]&m[758]&~m[759])|(~m[734]&m[755]&~m[756]&~m[758]&m[759])|(~m[734]&~m[755]&m[756]&~m[758]&m[759])|(m[734]&m[755]&m[756]&~m[758]&m[759])|(~m[734]&m[755]&m[756]&m[758]&m[759]))&UnbiasedRNG[187])|((m[734]&~m[755]&~m[756]&m[758]&~m[759])|(~m[734]&~m[755]&~m[756]&~m[758]&m[759])|(m[734]&~m[755]&~m[756]&~m[758]&m[759])|(m[734]&m[755]&~m[756]&~m[758]&m[759])|(m[734]&~m[755]&m[756]&~m[758]&m[759])|(~m[734]&~m[755]&~m[756]&m[758]&m[759])|(m[734]&~m[755]&~m[756]&m[758]&m[759])|(~m[734]&m[755]&~m[756]&m[758]&m[759])|(m[734]&m[755]&~m[756]&m[758]&m[759])|(~m[734]&~m[755]&m[756]&m[758]&m[759])|(m[734]&~m[755]&m[756]&m[758]&m[759])|(m[734]&m[755]&m[756]&m[758]&m[759]));
    m[762] = (((m[744]&~m[760]&~m[761]&~m[763]&~m[764])|(~m[744]&~m[760]&~m[761]&m[763]&~m[764])|(m[744]&m[760]&~m[761]&m[763]&~m[764])|(m[744]&~m[760]&m[761]&m[763]&~m[764])|(~m[744]&m[760]&~m[761]&~m[763]&m[764])|(~m[744]&~m[760]&m[761]&~m[763]&m[764])|(m[744]&m[760]&m[761]&~m[763]&m[764])|(~m[744]&m[760]&m[761]&m[763]&m[764]))&UnbiasedRNG[188])|((m[744]&~m[760]&~m[761]&m[763]&~m[764])|(~m[744]&~m[760]&~m[761]&~m[763]&m[764])|(m[744]&~m[760]&~m[761]&~m[763]&m[764])|(m[744]&m[760]&~m[761]&~m[763]&m[764])|(m[744]&~m[760]&m[761]&~m[763]&m[764])|(~m[744]&~m[760]&~m[761]&m[763]&m[764])|(m[744]&~m[760]&~m[761]&m[763]&m[764])|(~m[744]&m[760]&~m[761]&m[763]&m[764])|(m[744]&m[760]&~m[761]&m[763]&m[764])|(~m[744]&~m[760]&m[761]&m[763]&m[764])|(m[744]&~m[760]&m[761]&m[763]&m[764])|(m[744]&m[760]&m[761]&m[763]&m[764]));
    m[767] = (((m[749]&~m[765]&~m[766]&~m[768]&~m[769])|(~m[749]&~m[765]&~m[766]&m[768]&~m[769])|(m[749]&m[765]&~m[766]&m[768]&~m[769])|(m[749]&~m[765]&m[766]&m[768]&~m[769])|(~m[749]&m[765]&~m[766]&~m[768]&m[769])|(~m[749]&~m[765]&m[766]&~m[768]&m[769])|(m[749]&m[765]&m[766]&~m[768]&m[769])|(~m[749]&m[765]&m[766]&m[768]&m[769]))&UnbiasedRNG[189])|((m[749]&~m[765]&~m[766]&m[768]&~m[769])|(~m[749]&~m[765]&~m[766]&~m[768]&m[769])|(m[749]&~m[765]&~m[766]&~m[768]&m[769])|(m[749]&m[765]&~m[766]&~m[768]&m[769])|(m[749]&~m[765]&m[766]&~m[768]&m[769])|(~m[749]&~m[765]&~m[766]&m[768]&m[769])|(m[749]&~m[765]&~m[766]&m[768]&m[769])|(~m[749]&m[765]&~m[766]&m[768]&m[769])|(m[749]&m[765]&~m[766]&m[768]&m[769])|(~m[749]&~m[765]&m[766]&m[768]&m[769])|(m[749]&~m[765]&m[766]&m[768]&m[769])|(m[749]&m[765]&m[766]&m[768]&m[769]));
    m[772] = (((m[754]&~m[770]&~m[771]&~m[773]&~m[774])|(~m[754]&~m[770]&~m[771]&m[773]&~m[774])|(m[754]&m[770]&~m[771]&m[773]&~m[774])|(m[754]&~m[770]&m[771]&m[773]&~m[774])|(~m[754]&m[770]&~m[771]&~m[773]&m[774])|(~m[754]&~m[770]&m[771]&~m[773]&m[774])|(m[754]&m[770]&m[771]&~m[773]&m[774])|(~m[754]&m[770]&m[771]&m[773]&m[774]))&UnbiasedRNG[190])|((m[754]&~m[770]&~m[771]&m[773]&~m[774])|(~m[754]&~m[770]&~m[771]&~m[773]&m[774])|(m[754]&~m[770]&~m[771]&~m[773]&m[774])|(m[754]&m[770]&~m[771]&~m[773]&m[774])|(m[754]&~m[770]&m[771]&~m[773]&m[774])|(~m[754]&~m[770]&~m[771]&m[773]&m[774])|(m[754]&~m[770]&~m[771]&m[773]&m[774])|(~m[754]&m[770]&~m[771]&m[773]&m[774])|(m[754]&m[770]&~m[771]&m[773]&m[774])|(~m[754]&~m[770]&m[771]&m[773]&m[774])|(m[754]&~m[770]&m[771]&m[773]&m[774])|(m[754]&m[770]&m[771]&m[773]&m[774]));
    m[777] = (((m[759]&~m[775]&~m[776]&~m[778]&~m[779])|(~m[759]&~m[775]&~m[776]&m[778]&~m[779])|(m[759]&m[775]&~m[776]&m[778]&~m[779])|(m[759]&~m[775]&m[776]&m[778]&~m[779])|(~m[759]&m[775]&~m[776]&~m[778]&m[779])|(~m[759]&~m[775]&m[776]&~m[778]&m[779])|(m[759]&m[775]&m[776]&~m[778]&m[779])|(~m[759]&m[775]&m[776]&m[778]&m[779]))&UnbiasedRNG[191])|((m[759]&~m[775]&~m[776]&m[778]&~m[779])|(~m[759]&~m[775]&~m[776]&~m[778]&m[779])|(m[759]&~m[775]&~m[776]&~m[778]&m[779])|(m[759]&m[775]&~m[776]&~m[778]&m[779])|(m[759]&~m[775]&m[776]&~m[778]&m[779])|(~m[759]&~m[775]&~m[776]&m[778]&m[779])|(m[759]&~m[775]&~m[776]&m[778]&m[779])|(~m[759]&m[775]&~m[776]&m[778]&m[779])|(m[759]&m[775]&~m[776]&m[778]&m[779])|(~m[759]&~m[775]&m[776]&m[778]&m[779])|(m[759]&~m[775]&m[776]&m[778]&m[779])|(m[759]&m[775]&m[776]&m[778]&m[779]));
    m[782] = (((m[769]&~m[780]&~m[781]&~m[783]&~m[784])|(~m[769]&~m[780]&~m[781]&m[783]&~m[784])|(m[769]&m[780]&~m[781]&m[783]&~m[784])|(m[769]&~m[780]&m[781]&m[783]&~m[784])|(~m[769]&m[780]&~m[781]&~m[783]&m[784])|(~m[769]&~m[780]&m[781]&~m[783]&m[784])|(m[769]&m[780]&m[781]&~m[783]&m[784])|(~m[769]&m[780]&m[781]&m[783]&m[784]))&UnbiasedRNG[192])|((m[769]&~m[780]&~m[781]&m[783]&~m[784])|(~m[769]&~m[780]&~m[781]&~m[783]&m[784])|(m[769]&~m[780]&~m[781]&~m[783]&m[784])|(m[769]&m[780]&~m[781]&~m[783]&m[784])|(m[769]&~m[780]&m[781]&~m[783]&m[784])|(~m[769]&~m[780]&~m[781]&m[783]&m[784])|(m[769]&~m[780]&~m[781]&m[783]&m[784])|(~m[769]&m[780]&~m[781]&m[783]&m[784])|(m[769]&m[780]&~m[781]&m[783]&m[784])|(~m[769]&~m[780]&m[781]&m[783]&m[784])|(m[769]&~m[780]&m[781]&m[783]&m[784])|(m[769]&m[780]&m[781]&m[783]&m[784]));
    m[787] = (((m[774]&~m[785]&~m[786]&~m[788]&~m[789])|(~m[774]&~m[785]&~m[786]&m[788]&~m[789])|(m[774]&m[785]&~m[786]&m[788]&~m[789])|(m[774]&~m[785]&m[786]&m[788]&~m[789])|(~m[774]&m[785]&~m[786]&~m[788]&m[789])|(~m[774]&~m[785]&m[786]&~m[788]&m[789])|(m[774]&m[785]&m[786]&~m[788]&m[789])|(~m[774]&m[785]&m[786]&m[788]&m[789]))&UnbiasedRNG[193])|((m[774]&~m[785]&~m[786]&m[788]&~m[789])|(~m[774]&~m[785]&~m[786]&~m[788]&m[789])|(m[774]&~m[785]&~m[786]&~m[788]&m[789])|(m[774]&m[785]&~m[786]&~m[788]&m[789])|(m[774]&~m[785]&m[786]&~m[788]&m[789])|(~m[774]&~m[785]&~m[786]&m[788]&m[789])|(m[774]&~m[785]&~m[786]&m[788]&m[789])|(~m[774]&m[785]&~m[786]&m[788]&m[789])|(m[774]&m[785]&~m[786]&m[788]&m[789])|(~m[774]&~m[785]&m[786]&m[788]&m[789])|(m[774]&~m[785]&m[786]&m[788]&m[789])|(m[774]&m[785]&m[786]&m[788]&m[789]));
    m[792] = (((m[779]&~m[790]&~m[791]&~m[793]&~m[794])|(~m[779]&~m[790]&~m[791]&m[793]&~m[794])|(m[779]&m[790]&~m[791]&m[793]&~m[794])|(m[779]&~m[790]&m[791]&m[793]&~m[794])|(~m[779]&m[790]&~m[791]&~m[793]&m[794])|(~m[779]&~m[790]&m[791]&~m[793]&m[794])|(m[779]&m[790]&m[791]&~m[793]&m[794])|(~m[779]&m[790]&m[791]&m[793]&m[794]))&UnbiasedRNG[194])|((m[779]&~m[790]&~m[791]&m[793]&~m[794])|(~m[779]&~m[790]&~m[791]&~m[793]&m[794])|(m[779]&~m[790]&~m[791]&~m[793]&m[794])|(m[779]&m[790]&~m[791]&~m[793]&m[794])|(m[779]&~m[790]&m[791]&~m[793]&m[794])|(~m[779]&~m[790]&~m[791]&m[793]&m[794])|(m[779]&~m[790]&~m[791]&m[793]&m[794])|(~m[779]&m[790]&~m[791]&m[793]&m[794])|(m[779]&m[790]&~m[791]&m[793]&m[794])|(~m[779]&~m[790]&m[791]&m[793]&m[794])|(m[779]&~m[790]&m[791]&m[793]&m[794])|(m[779]&m[790]&m[791]&m[793]&m[794]));
    m[797] = (((m[789]&~m[795]&~m[796]&~m[798]&~m[799])|(~m[789]&~m[795]&~m[796]&m[798]&~m[799])|(m[789]&m[795]&~m[796]&m[798]&~m[799])|(m[789]&~m[795]&m[796]&m[798]&~m[799])|(~m[789]&m[795]&~m[796]&~m[798]&m[799])|(~m[789]&~m[795]&m[796]&~m[798]&m[799])|(m[789]&m[795]&m[796]&~m[798]&m[799])|(~m[789]&m[795]&m[796]&m[798]&m[799]))&UnbiasedRNG[195])|((m[789]&~m[795]&~m[796]&m[798]&~m[799])|(~m[789]&~m[795]&~m[796]&~m[798]&m[799])|(m[789]&~m[795]&~m[796]&~m[798]&m[799])|(m[789]&m[795]&~m[796]&~m[798]&m[799])|(m[789]&~m[795]&m[796]&~m[798]&m[799])|(~m[789]&~m[795]&~m[796]&m[798]&m[799])|(m[789]&~m[795]&~m[796]&m[798]&m[799])|(~m[789]&m[795]&~m[796]&m[798]&m[799])|(m[789]&m[795]&~m[796]&m[798]&m[799])|(~m[789]&~m[795]&m[796]&m[798]&m[799])|(m[789]&~m[795]&m[796]&m[798]&m[799])|(m[789]&m[795]&m[796]&m[798]&m[799]));
    m[802] = (((m[794]&~m[800]&~m[801]&~m[803]&~m[804])|(~m[794]&~m[800]&~m[801]&m[803]&~m[804])|(m[794]&m[800]&~m[801]&m[803]&~m[804])|(m[794]&~m[800]&m[801]&m[803]&~m[804])|(~m[794]&m[800]&~m[801]&~m[803]&m[804])|(~m[794]&~m[800]&m[801]&~m[803]&m[804])|(m[794]&m[800]&m[801]&~m[803]&m[804])|(~m[794]&m[800]&m[801]&m[803]&m[804]))&UnbiasedRNG[196])|((m[794]&~m[800]&~m[801]&m[803]&~m[804])|(~m[794]&~m[800]&~m[801]&~m[803]&m[804])|(m[794]&~m[800]&~m[801]&~m[803]&m[804])|(m[794]&m[800]&~m[801]&~m[803]&m[804])|(m[794]&~m[800]&m[801]&~m[803]&m[804])|(~m[794]&~m[800]&~m[801]&m[803]&m[804])|(m[794]&~m[800]&~m[801]&m[803]&m[804])|(~m[794]&m[800]&~m[801]&m[803]&m[804])|(m[794]&m[800]&~m[801]&m[803]&m[804])|(~m[794]&~m[800]&m[801]&m[803]&m[804])|(m[794]&~m[800]&m[801]&m[803]&m[804])|(m[794]&m[800]&m[801]&m[803]&m[804]));
    m[807] = (((m[804]&~m[805]&~m[806]&~m[808]&~m[809])|(~m[804]&~m[805]&~m[806]&m[808]&~m[809])|(m[804]&m[805]&~m[806]&m[808]&~m[809])|(m[804]&~m[805]&m[806]&m[808]&~m[809])|(~m[804]&m[805]&~m[806]&~m[808]&m[809])|(~m[804]&~m[805]&m[806]&~m[808]&m[809])|(m[804]&m[805]&m[806]&~m[808]&m[809])|(~m[804]&m[805]&m[806]&m[808]&m[809]))&UnbiasedRNG[197])|((m[804]&~m[805]&~m[806]&m[808]&~m[809])|(~m[804]&~m[805]&~m[806]&~m[808]&m[809])|(m[804]&~m[805]&~m[806]&~m[808]&m[809])|(m[804]&m[805]&~m[806]&~m[808]&m[809])|(m[804]&~m[805]&m[806]&~m[808]&m[809])|(~m[804]&~m[805]&~m[806]&m[808]&m[809])|(m[804]&~m[805]&~m[806]&m[808]&m[809])|(~m[804]&m[805]&~m[806]&m[808]&m[809])|(m[804]&m[805]&~m[806]&m[808]&m[809])|(~m[804]&~m[805]&m[806]&m[808]&m[809])|(m[804]&~m[805]&m[806]&m[808]&m[809])|(m[804]&m[805]&m[806]&m[808]&m[809]));
end

always @(posedge color2_clk) begin
    m[160] = (((~m[10]&~m[60]&~m[260])|(m[10]&m[60]&~m[260]))&BiasedRNG[239])|(((m[10]&~m[60]&~m[260])|(~m[10]&m[60]&m[260]))&~BiasedRNG[239])|((~m[10]&~m[60]&m[260])|(m[10]&~m[60]&m[260])|(m[10]&m[60]&m[260]));
    m[161] = (((~m[10]&~m[70]&~m[261])|(m[10]&m[70]&~m[261]))&BiasedRNG[240])|(((m[10]&~m[70]&~m[261])|(~m[10]&m[70]&m[261]))&~BiasedRNG[240])|((~m[10]&~m[70]&m[261])|(m[10]&~m[70]&m[261])|(m[10]&m[70]&m[261]));
    m[170] = (((~m[11]&~m[61]&~m[270])|(m[11]&m[61]&~m[270]))&BiasedRNG[241])|(((m[11]&~m[61]&~m[270])|(~m[11]&m[61]&m[270]))&~BiasedRNG[241])|((~m[11]&~m[61]&m[270])|(m[11]&~m[61]&m[270])|(m[11]&m[61]&m[270]));
    m[171] = (((~m[11]&~m[71]&~m[271])|(m[11]&m[71]&~m[271]))&BiasedRNG[242])|(((m[11]&~m[71]&~m[271])|(~m[11]&m[71]&m[271]))&~BiasedRNG[242])|((~m[11]&~m[71]&m[271])|(m[11]&~m[71]&m[271])|(m[11]&m[71]&m[271]));
    m[182] = (((~m[44]&~m[82]&~m[282])|(m[44]&m[82]&~m[282]))&BiasedRNG[243])|(((m[44]&~m[82]&~m[282])|(~m[44]&m[82]&m[282]))&~BiasedRNG[243])|((~m[44]&~m[82]&m[282])|(m[44]&~m[82]&m[282])|(m[44]&m[82]&m[282]));
    m[183] = (((~m[44]&~m[92]&~m[283])|(m[44]&m[92]&~m[283]))&BiasedRNG[244])|(((m[44]&~m[92]&~m[283])|(~m[44]&m[92]&m[283]))&~BiasedRNG[244])|((~m[44]&~m[92]&m[283])|(m[44]&~m[92]&m[283])|(m[44]&m[92]&m[283]));
    m[184] = (((~m[44]&~m[102]&~m[284])|(m[44]&m[102]&~m[284]))&BiasedRNG[245])|(((m[44]&~m[102]&~m[284])|(~m[44]&m[102]&m[284]))&~BiasedRNG[245])|((~m[44]&~m[102]&m[284])|(m[44]&~m[102]&m[284])|(m[44]&m[102]&m[284]));
    m[185] = (((~m[44]&~m[112]&~m[285])|(m[44]&m[112]&~m[285]))&BiasedRNG[246])|(((m[44]&~m[112]&~m[285])|(~m[44]&m[112]&m[285]))&~BiasedRNG[246])|((~m[44]&~m[112]&m[285])|(m[44]&~m[112]&m[285])|(m[44]&m[112]&m[285]));
    m[186] = (((~m[45]&~m[122]&~m[286])|(m[45]&m[122]&~m[286]))&BiasedRNG[247])|(((m[45]&~m[122]&~m[286])|(~m[45]&m[122]&m[286]))&~BiasedRNG[247])|((~m[45]&~m[122]&m[286])|(m[45]&~m[122]&m[286])|(m[45]&m[122]&m[286]));
    m[187] = (((~m[45]&~m[132]&~m[287])|(m[45]&m[132]&~m[287]))&BiasedRNG[248])|(((m[45]&~m[132]&~m[287])|(~m[45]&m[132]&m[287]))&~BiasedRNG[248])|((~m[45]&~m[132]&m[287])|(m[45]&~m[132]&m[287])|(m[45]&m[132]&m[287]));
    m[188] = (((~m[45]&~m[142]&~m[288])|(m[45]&m[142]&~m[288]))&BiasedRNG[249])|(((m[45]&~m[142]&~m[288])|(~m[45]&m[142]&m[288]))&~BiasedRNG[249])|((~m[45]&~m[142]&m[288])|(m[45]&~m[142]&m[288])|(m[45]&m[142]&m[288]));
    m[189] = (((~m[45]&~m[152]&~m[289])|(m[45]&m[152]&~m[289]))&BiasedRNG[250])|(((m[45]&~m[152]&~m[289])|(~m[45]&m[152]&m[289]))&~BiasedRNG[250])|((~m[45]&~m[152]&m[289])|(m[45]&~m[152]&m[289])|(m[45]&m[152]&m[289]));
    m[192] = (((~m[46]&~m[83]&~m[292])|(m[46]&m[83]&~m[292]))&BiasedRNG[251])|(((m[46]&~m[83]&~m[292])|(~m[46]&m[83]&m[292]))&~BiasedRNG[251])|((~m[46]&~m[83]&m[292])|(m[46]&~m[83]&m[292])|(m[46]&m[83]&m[292]));
    m[193] = (((~m[46]&~m[93]&~m[293])|(m[46]&m[93]&~m[293]))&BiasedRNG[252])|(((m[46]&~m[93]&~m[293])|(~m[46]&m[93]&m[293]))&~BiasedRNG[252])|((~m[46]&~m[93]&m[293])|(m[46]&~m[93]&m[293])|(m[46]&m[93]&m[293]));
    m[194] = (((~m[46]&~m[103]&~m[294])|(m[46]&m[103]&~m[294]))&BiasedRNG[253])|(((m[46]&~m[103]&~m[294])|(~m[46]&m[103]&m[294]))&~BiasedRNG[253])|((~m[46]&~m[103]&m[294])|(m[46]&~m[103]&m[294])|(m[46]&m[103]&m[294]));
    m[195] = (((~m[46]&~m[113]&~m[295])|(m[46]&m[113]&~m[295]))&BiasedRNG[254])|(((m[46]&~m[113]&~m[295])|(~m[46]&m[113]&m[295]))&~BiasedRNG[254])|((~m[46]&~m[113]&m[295])|(m[46]&~m[113]&m[295])|(m[46]&m[113]&m[295]));
    m[196] = (((~m[47]&~m[123]&~m[296])|(m[47]&m[123]&~m[296]))&BiasedRNG[255])|(((m[47]&~m[123]&~m[296])|(~m[47]&m[123]&m[296]))&~BiasedRNG[255])|((~m[47]&~m[123]&m[296])|(m[47]&~m[123]&m[296])|(m[47]&m[123]&m[296]));
    m[197] = (((~m[47]&~m[133]&~m[297])|(m[47]&m[133]&~m[297]))&BiasedRNG[256])|(((m[47]&~m[133]&~m[297])|(~m[47]&m[133]&m[297]))&~BiasedRNG[256])|((~m[47]&~m[133]&m[297])|(m[47]&~m[133]&m[297])|(m[47]&m[133]&m[297]));
    m[198] = (((~m[47]&~m[143]&~m[298])|(m[47]&m[143]&~m[298]))&BiasedRNG[257])|(((m[47]&~m[143]&~m[298])|(~m[47]&m[143]&m[298]))&~BiasedRNG[257])|((~m[47]&~m[143]&m[298])|(m[47]&~m[143]&m[298])|(m[47]&m[143]&m[298]));
    m[199] = (((~m[47]&~m[153]&~m[299])|(m[47]&m[153]&~m[299]))&BiasedRNG[258])|(((m[47]&~m[153]&~m[299])|(~m[47]&m[153]&m[299]))&~BiasedRNG[258])|((~m[47]&~m[153]&m[299])|(m[47]&~m[153]&m[299])|(m[47]&m[153]&m[299]));
    m[202] = (((~m[48]&~m[84]&~m[302])|(m[48]&m[84]&~m[302]))&BiasedRNG[259])|(((m[48]&~m[84]&~m[302])|(~m[48]&m[84]&m[302]))&~BiasedRNG[259])|((~m[48]&~m[84]&m[302])|(m[48]&~m[84]&m[302])|(m[48]&m[84]&m[302]));
    m[203] = (((~m[48]&~m[94]&~m[303])|(m[48]&m[94]&~m[303]))&BiasedRNG[260])|(((m[48]&~m[94]&~m[303])|(~m[48]&m[94]&m[303]))&~BiasedRNG[260])|((~m[48]&~m[94]&m[303])|(m[48]&~m[94]&m[303])|(m[48]&m[94]&m[303]));
    m[204] = (((~m[48]&~m[104]&~m[304])|(m[48]&m[104]&~m[304]))&BiasedRNG[261])|(((m[48]&~m[104]&~m[304])|(~m[48]&m[104]&m[304]))&~BiasedRNG[261])|((~m[48]&~m[104]&m[304])|(m[48]&~m[104]&m[304])|(m[48]&m[104]&m[304]));
    m[205] = (((~m[48]&~m[114]&~m[305])|(m[48]&m[114]&~m[305]))&BiasedRNG[262])|(((m[48]&~m[114]&~m[305])|(~m[48]&m[114]&m[305]))&~BiasedRNG[262])|((~m[48]&~m[114]&m[305])|(m[48]&~m[114]&m[305])|(m[48]&m[114]&m[305]));
    m[206] = (((~m[49]&~m[124]&~m[306])|(m[49]&m[124]&~m[306]))&BiasedRNG[263])|(((m[49]&~m[124]&~m[306])|(~m[49]&m[124]&m[306]))&~BiasedRNG[263])|((~m[49]&~m[124]&m[306])|(m[49]&~m[124]&m[306])|(m[49]&m[124]&m[306]));
    m[207] = (((~m[49]&~m[134]&~m[307])|(m[49]&m[134]&~m[307]))&BiasedRNG[264])|(((m[49]&~m[134]&~m[307])|(~m[49]&m[134]&m[307]))&~BiasedRNG[264])|((~m[49]&~m[134]&m[307])|(m[49]&~m[134]&m[307])|(m[49]&m[134]&m[307]));
    m[208] = (((~m[49]&~m[144]&~m[308])|(m[49]&m[144]&~m[308]))&BiasedRNG[265])|(((m[49]&~m[144]&~m[308])|(~m[49]&m[144]&m[308]))&~BiasedRNG[265])|((~m[49]&~m[144]&m[308])|(m[49]&~m[144]&m[308])|(m[49]&m[144]&m[308]));
    m[209] = (((~m[49]&~m[154]&~m[309])|(m[49]&m[154]&~m[309]))&BiasedRNG[266])|(((m[49]&~m[154]&~m[309])|(~m[49]&m[154]&m[309]))&~BiasedRNG[266])|((~m[49]&~m[154]&m[309])|(m[49]&~m[154]&m[309])|(m[49]&m[154]&m[309]));
    m[212] = (((~m[50]&~m[85]&~m[312])|(m[50]&m[85]&~m[312]))&BiasedRNG[267])|(((m[50]&~m[85]&~m[312])|(~m[50]&m[85]&m[312]))&~BiasedRNG[267])|((~m[50]&~m[85]&m[312])|(m[50]&~m[85]&m[312])|(m[50]&m[85]&m[312]));
    m[213] = (((~m[50]&~m[95]&~m[313])|(m[50]&m[95]&~m[313]))&BiasedRNG[268])|(((m[50]&~m[95]&~m[313])|(~m[50]&m[95]&m[313]))&~BiasedRNG[268])|((~m[50]&~m[95]&m[313])|(m[50]&~m[95]&m[313])|(m[50]&m[95]&m[313]));
    m[214] = (((~m[50]&~m[105]&~m[314])|(m[50]&m[105]&~m[314]))&BiasedRNG[269])|(((m[50]&~m[105]&~m[314])|(~m[50]&m[105]&m[314]))&~BiasedRNG[269])|((~m[50]&~m[105]&m[314])|(m[50]&~m[105]&m[314])|(m[50]&m[105]&m[314]));
    m[215] = (((~m[50]&~m[115]&~m[315])|(m[50]&m[115]&~m[315]))&BiasedRNG[270])|(((m[50]&~m[115]&~m[315])|(~m[50]&m[115]&m[315]))&~BiasedRNG[270])|((~m[50]&~m[115]&m[315])|(m[50]&~m[115]&m[315])|(m[50]&m[115]&m[315]));
    m[216] = (((~m[51]&~m[125]&~m[316])|(m[51]&m[125]&~m[316]))&BiasedRNG[271])|(((m[51]&~m[125]&~m[316])|(~m[51]&m[125]&m[316]))&~BiasedRNG[271])|((~m[51]&~m[125]&m[316])|(m[51]&~m[125]&m[316])|(m[51]&m[125]&m[316]));
    m[217] = (((~m[51]&~m[135]&~m[317])|(m[51]&m[135]&~m[317]))&BiasedRNG[272])|(((m[51]&~m[135]&~m[317])|(~m[51]&m[135]&m[317]))&~BiasedRNG[272])|((~m[51]&~m[135]&m[317])|(m[51]&~m[135]&m[317])|(m[51]&m[135]&m[317]));
    m[218] = (((~m[51]&~m[145]&~m[318])|(m[51]&m[145]&~m[318]))&BiasedRNG[273])|(((m[51]&~m[145]&~m[318])|(~m[51]&m[145]&m[318]))&~BiasedRNG[273])|((~m[51]&~m[145]&m[318])|(m[51]&~m[145]&m[318])|(m[51]&m[145]&m[318]));
    m[219] = (((~m[51]&~m[155]&~m[319])|(m[51]&m[155]&~m[319]))&BiasedRNG[274])|(((m[51]&~m[155]&~m[319])|(~m[51]&m[155]&m[319]))&~BiasedRNG[274])|((~m[51]&~m[155]&m[319])|(m[51]&~m[155]&m[319])|(m[51]&m[155]&m[319]));
    m[222] = (((~m[52]&~m[86]&~m[322])|(m[52]&m[86]&~m[322]))&BiasedRNG[275])|(((m[52]&~m[86]&~m[322])|(~m[52]&m[86]&m[322]))&~BiasedRNG[275])|((~m[52]&~m[86]&m[322])|(m[52]&~m[86]&m[322])|(m[52]&m[86]&m[322]));
    m[223] = (((~m[52]&~m[96]&~m[323])|(m[52]&m[96]&~m[323]))&BiasedRNG[276])|(((m[52]&~m[96]&~m[323])|(~m[52]&m[96]&m[323]))&~BiasedRNG[276])|((~m[52]&~m[96]&m[323])|(m[52]&~m[96]&m[323])|(m[52]&m[96]&m[323]));
    m[224] = (((~m[52]&~m[106]&~m[324])|(m[52]&m[106]&~m[324]))&BiasedRNG[277])|(((m[52]&~m[106]&~m[324])|(~m[52]&m[106]&m[324]))&~BiasedRNG[277])|((~m[52]&~m[106]&m[324])|(m[52]&~m[106]&m[324])|(m[52]&m[106]&m[324]));
    m[225] = (((~m[52]&~m[116]&~m[325])|(m[52]&m[116]&~m[325]))&BiasedRNG[278])|(((m[52]&~m[116]&~m[325])|(~m[52]&m[116]&m[325]))&~BiasedRNG[278])|((~m[52]&~m[116]&m[325])|(m[52]&~m[116]&m[325])|(m[52]&m[116]&m[325]));
    m[226] = (((~m[53]&~m[126]&~m[326])|(m[53]&m[126]&~m[326]))&BiasedRNG[279])|(((m[53]&~m[126]&~m[326])|(~m[53]&m[126]&m[326]))&~BiasedRNG[279])|((~m[53]&~m[126]&m[326])|(m[53]&~m[126]&m[326])|(m[53]&m[126]&m[326]));
    m[227] = (((~m[53]&~m[136]&~m[327])|(m[53]&m[136]&~m[327]))&BiasedRNG[280])|(((m[53]&~m[136]&~m[327])|(~m[53]&m[136]&m[327]))&~BiasedRNG[280])|((~m[53]&~m[136]&m[327])|(m[53]&~m[136]&m[327])|(m[53]&m[136]&m[327]));
    m[228] = (((~m[53]&~m[146]&~m[328])|(m[53]&m[146]&~m[328]))&BiasedRNG[281])|(((m[53]&~m[146]&~m[328])|(~m[53]&m[146]&m[328]))&~BiasedRNG[281])|((~m[53]&~m[146]&m[328])|(m[53]&~m[146]&m[328])|(m[53]&m[146]&m[328]));
    m[229] = (((~m[53]&~m[156]&~m[329])|(m[53]&m[156]&~m[329]))&BiasedRNG[282])|(((m[53]&~m[156]&~m[329])|(~m[53]&m[156]&m[329]))&~BiasedRNG[282])|((~m[53]&~m[156]&m[329])|(m[53]&~m[156]&m[329])|(m[53]&m[156]&m[329]));
    m[232] = (((~m[54]&~m[87]&~m[332])|(m[54]&m[87]&~m[332]))&BiasedRNG[283])|(((m[54]&~m[87]&~m[332])|(~m[54]&m[87]&m[332]))&~BiasedRNG[283])|((~m[54]&~m[87]&m[332])|(m[54]&~m[87]&m[332])|(m[54]&m[87]&m[332]));
    m[233] = (((~m[54]&~m[97]&~m[333])|(m[54]&m[97]&~m[333]))&BiasedRNG[284])|(((m[54]&~m[97]&~m[333])|(~m[54]&m[97]&m[333]))&~BiasedRNG[284])|((~m[54]&~m[97]&m[333])|(m[54]&~m[97]&m[333])|(m[54]&m[97]&m[333]));
    m[234] = (((~m[54]&~m[107]&~m[334])|(m[54]&m[107]&~m[334]))&BiasedRNG[285])|(((m[54]&~m[107]&~m[334])|(~m[54]&m[107]&m[334]))&~BiasedRNG[285])|((~m[54]&~m[107]&m[334])|(m[54]&~m[107]&m[334])|(m[54]&m[107]&m[334]));
    m[235] = (((~m[54]&~m[117]&~m[335])|(m[54]&m[117]&~m[335]))&BiasedRNG[286])|(((m[54]&~m[117]&~m[335])|(~m[54]&m[117]&m[335]))&~BiasedRNG[286])|((~m[54]&~m[117]&m[335])|(m[54]&~m[117]&m[335])|(m[54]&m[117]&m[335]));
    m[236] = (((~m[55]&~m[127]&~m[336])|(m[55]&m[127]&~m[336]))&BiasedRNG[287])|(((m[55]&~m[127]&~m[336])|(~m[55]&m[127]&m[336]))&~BiasedRNG[287])|((~m[55]&~m[127]&m[336])|(m[55]&~m[127]&m[336])|(m[55]&m[127]&m[336]));
    m[237] = (((~m[55]&~m[137]&~m[337])|(m[55]&m[137]&~m[337]))&BiasedRNG[288])|(((m[55]&~m[137]&~m[337])|(~m[55]&m[137]&m[337]))&~BiasedRNG[288])|((~m[55]&~m[137]&m[337])|(m[55]&~m[137]&m[337])|(m[55]&m[137]&m[337]));
    m[238] = (((~m[55]&~m[147]&~m[338])|(m[55]&m[147]&~m[338]))&BiasedRNG[289])|(((m[55]&~m[147]&~m[338])|(~m[55]&m[147]&m[338]))&~BiasedRNG[289])|((~m[55]&~m[147]&m[338])|(m[55]&~m[147]&m[338])|(m[55]&m[147]&m[338]));
    m[239] = (((~m[55]&~m[157]&~m[339])|(m[55]&m[157]&~m[339]))&BiasedRNG[290])|(((m[55]&~m[157]&~m[339])|(~m[55]&m[157]&m[339]))&~BiasedRNG[290])|((~m[55]&~m[157]&m[339])|(m[55]&~m[157]&m[339])|(m[55]&m[157]&m[339]));
    m[242] = (((~m[56]&~m[88]&~m[342])|(m[56]&m[88]&~m[342]))&BiasedRNG[291])|(((m[56]&~m[88]&~m[342])|(~m[56]&m[88]&m[342]))&~BiasedRNG[291])|((~m[56]&~m[88]&m[342])|(m[56]&~m[88]&m[342])|(m[56]&m[88]&m[342]));
    m[243] = (((~m[56]&~m[98]&~m[343])|(m[56]&m[98]&~m[343]))&BiasedRNG[292])|(((m[56]&~m[98]&~m[343])|(~m[56]&m[98]&m[343]))&~BiasedRNG[292])|((~m[56]&~m[98]&m[343])|(m[56]&~m[98]&m[343])|(m[56]&m[98]&m[343]));
    m[244] = (((~m[56]&~m[108]&~m[344])|(m[56]&m[108]&~m[344]))&BiasedRNG[293])|(((m[56]&~m[108]&~m[344])|(~m[56]&m[108]&m[344]))&~BiasedRNG[293])|((~m[56]&~m[108]&m[344])|(m[56]&~m[108]&m[344])|(m[56]&m[108]&m[344]));
    m[245] = (((~m[56]&~m[118]&~m[345])|(m[56]&m[118]&~m[345]))&BiasedRNG[294])|(((m[56]&~m[118]&~m[345])|(~m[56]&m[118]&m[345]))&~BiasedRNG[294])|((~m[56]&~m[118]&m[345])|(m[56]&~m[118]&m[345])|(m[56]&m[118]&m[345]));
    m[246] = (((~m[57]&~m[128]&~m[346])|(m[57]&m[128]&~m[346]))&BiasedRNG[295])|(((m[57]&~m[128]&~m[346])|(~m[57]&m[128]&m[346]))&~BiasedRNG[295])|((~m[57]&~m[128]&m[346])|(m[57]&~m[128]&m[346])|(m[57]&m[128]&m[346]));
    m[247] = (((~m[57]&~m[138]&~m[347])|(m[57]&m[138]&~m[347]))&BiasedRNG[296])|(((m[57]&~m[138]&~m[347])|(~m[57]&m[138]&m[347]))&~BiasedRNG[296])|((~m[57]&~m[138]&m[347])|(m[57]&~m[138]&m[347])|(m[57]&m[138]&m[347]));
    m[248] = (((~m[57]&~m[148]&~m[348])|(m[57]&m[148]&~m[348]))&BiasedRNG[297])|(((m[57]&~m[148]&~m[348])|(~m[57]&m[148]&m[348]))&~BiasedRNG[297])|((~m[57]&~m[148]&m[348])|(m[57]&~m[148]&m[348])|(m[57]&m[148]&m[348]));
    m[249] = (((~m[57]&~m[158]&~m[349])|(m[57]&m[158]&~m[349]))&BiasedRNG[298])|(((m[57]&~m[158]&~m[349])|(~m[57]&m[158]&m[349]))&~BiasedRNG[298])|((~m[57]&~m[158]&m[349])|(m[57]&~m[158]&m[349])|(m[57]&m[158]&m[349]));
    m[252] = (((~m[58]&~m[89]&~m[352])|(m[58]&m[89]&~m[352]))&BiasedRNG[299])|(((m[58]&~m[89]&~m[352])|(~m[58]&m[89]&m[352]))&~BiasedRNG[299])|((~m[58]&~m[89]&m[352])|(m[58]&~m[89]&m[352])|(m[58]&m[89]&m[352]));
    m[253] = (((~m[58]&~m[99]&~m[353])|(m[58]&m[99]&~m[353]))&BiasedRNG[300])|(((m[58]&~m[99]&~m[353])|(~m[58]&m[99]&m[353]))&~BiasedRNG[300])|((~m[58]&~m[99]&m[353])|(m[58]&~m[99]&m[353])|(m[58]&m[99]&m[353]));
    m[254] = (((~m[58]&~m[109]&~m[354])|(m[58]&m[109]&~m[354]))&BiasedRNG[301])|(((m[58]&~m[109]&~m[354])|(~m[58]&m[109]&m[354]))&~BiasedRNG[301])|((~m[58]&~m[109]&m[354])|(m[58]&~m[109]&m[354])|(m[58]&m[109]&m[354]));
    m[255] = (((~m[58]&~m[119]&~m[355])|(m[58]&m[119]&~m[355]))&BiasedRNG[302])|(((m[58]&~m[119]&~m[355])|(~m[58]&m[119]&m[355]))&~BiasedRNG[302])|((~m[58]&~m[119]&m[355])|(m[58]&~m[119]&m[355])|(m[58]&m[119]&m[355]));
    m[256] = (((~m[59]&~m[129]&~m[356])|(m[59]&m[129]&~m[356]))&BiasedRNG[303])|(((m[59]&~m[129]&~m[356])|(~m[59]&m[129]&m[356]))&~BiasedRNG[303])|((~m[59]&~m[129]&m[356])|(m[59]&~m[129]&m[356])|(m[59]&m[129]&m[356]));
    m[257] = (((~m[59]&~m[139]&~m[357])|(m[59]&m[139]&~m[357]))&BiasedRNG[304])|(((m[59]&~m[139]&~m[357])|(~m[59]&m[139]&m[357]))&~BiasedRNG[304])|((~m[59]&~m[139]&m[357])|(m[59]&~m[139]&m[357])|(m[59]&m[139]&m[357]));
    m[258] = (((~m[59]&~m[149]&~m[358])|(m[59]&m[149]&~m[358]))&BiasedRNG[305])|(((m[59]&~m[149]&~m[358])|(~m[59]&m[149]&m[358]))&~BiasedRNG[305])|((~m[59]&~m[149]&m[358])|(m[59]&~m[149]&m[358])|(m[59]&m[149]&m[358]));
    m[259] = (((~m[59]&~m[159]&~m[359])|(m[59]&m[159]&~m[359]))&BiasedRNG[306])|(((m[59]&~m[159]&~m[359])|(~m[59]&m[159]&m[359]))&~BiasedRNG[306])|((~m[59]&~m[159]&m[359])|(m[59]&~m[159]&m[359])|(m[59]&m[159]&m[359]));
    m[262] = (((m[80]&~m[162]&m[365])|(~m[80]&m[162]&m[365]))&BiasedRNG[307])|(((m[80]&m[162]&~m[365]))&~BiasedRNG[307])|((m[80]&m[162]&m[365]));
    m[263] = (((m[90]&~m[163]&m[375])|(~m[90]&m[163]&m[375]))&BiasedRNG[308])|(((m[90]&m[163]&~m[375]))&~BiasedRNG[308])|((m[90]&m[163]&m[375]));
    m[264] = (((m[100]&~m[164]&m[390])|(~m[100]&m[164]&m[390]))&BiasedRNG[309])|(((m[100]&m[164]&~m[390]))&~BiasedRNG[309])|((m[100]&m[164]&m[390]));
    m[265] = (((m[110]&~m[165]&m[410])|(~m[110]&m[165]&m[410]))&BiasedRNG[310])|(((m[110]&m[165]&~m[410]))&~BiasedRNG[310])|((m[110]&m[165]&m[410]));
    m[266] = (((m[120]&~m[166]&m[435])|(~m[120]&m[166]&m[435]))&BiasedRNG[311])|(((m[120]&m[166]&~m[435]))&~BiasedRNG[311])|((m[120]&m[166]&m[435]));
    m[267] = (((m[130]&~m[167]&m[465])|(~m[130]&m[167]&m[465]))&BiasedRNG[312])|(((m[130]&m[167]&~m[465]))&~BiasedRNG[312])|((m[130]&m[167]&m[465]));
    m[268] = (((m[140]&~m[168]&m[500])|(~m[140]&m[168]&m[500]))&BiasedRNG[313])|(((m[140]&m[168]&~m[500]))&~BiasedRNG[313])|((m[140]&m[168]&m[500]));
    m[269] = (((m[150]&~m[169]&m[540])|(~m[150]&m[169]&m[540]))&BiasedRNG[314])|(((m[150]&m[169]&~m[540]))&~BiasedRNG[314])|((m[150]&m[169]&m[540]));
    m[272] = (((m[81]&~m[172]&m[376])|(~m[81]&m[172]&m[376]))&BiasedRNG[315])|(((m[81]&m[172]&~m[376]))&~BiasedRNG[315])|((m[81]&m[172]&m[376]));
    m[273] = (((m[91]&~m[173]&m[391])|(~m[91]&m[173]&m[391]))&BiasedRNG[316])|(((m[91]&m[173]&~m[391]))&~BiasedRNG[316])|((m[91]&m[173]&m[391]));
    m[274] = (((m[101]&~m[174]&m[411])|(~m[101]&m[174]&m[411]))&BiasedRNG[317])|(((m[101]&m[174]&~m[411]))&~BiasedRNG[317])|((m[101]&m[174]&m[411]));
    m[275] = (((m[111]&~m[175]&m[436])|(~m[111]&m[175]&m[436]))&BiasedRNG[318])|(((m[111]&m[175]&~m[436]))&~BiasedRNG[318])|((m[111]&m[175]&m[436]));
    m[276] = (((m[121]&~m[176]&m[466])|(~m[121]&m[176]&m[466]))&BiasedRNG[319])|(((m[121]&m[176]&~m[466]))&~BiasedRNG[319])|((m[121]&m[176]&m[466]));
    m[277] = (((m[131]&~m[177]&m[501])|(~m[131]&m[177]&m[501]))&BiasedRNG[320])|(((m[131]&m[177]&~m[501]))&~BiasedRNG[320])|((m[131]&m[177]&m[501]));
    m[278] = (((m[141]&~m[178]&m[541])|(~m[141]&m[178]&m[541]))&BiasedRNG[321])|(((m[141]&m[178]&~m[541]))&~BiasedRNG[321])|((m[141]&m[178]&m[541]));
    m[279] = (((m[151]&~m[179]&m[586])|(~m[151]&m[179]&m[586]))&BiasedRNG[322])|(((m[151]&m[179]&~m[586]))&~BiasedRNG[322])|((m[151]&m[179]&m[586]));
    m[280] = (((m[62]&~m[180]&m[371])|(~m[62]&m[180]&m[371]))&BiasedRNG[323])|(((m[62]&m[180]&~m[371]))&~BiasedRNG[323])|((m[62]&m[180]&m[371]));
    m[281] = (((m[72]&~m[181]&m[381])|(~m[72]&m[181]&m[381]))&BiasedRNG[324])|(((m[72]&m[181]&~m[381]))&~BiasedRNG[324])|((m[72]&m[181]&m[381]));
    m[290] = (((m[63]&~m[190]&m[386])|(~m[63]&m[190]&m[386]))&BiasedRNG[325])|(((m[63]&m[190]&~m[386]))&~BiasedRNG[325])|((m[63]&m[190]&m[386]));
    m[291] = (((m[73]&~m[191]&m[401])|(~m[73]&m[191]&m[401]))&BiasedRNG[326])|(((m[73]&m[191]&~m[401]))&~BiasedRNG[326])|((m[73]&m[191]&m[401]));
    m[300] = (((m[64]&~m[200]&m[406])|(~m[64]&m[200]&m[406]))&BiasedRNG[327])|(((m[64]&m[200]&~m[406]))&~BiasedRNG[327])|((m[64]&m[200]&m[406]));
    m[301] = (((m[74]&~m[201]&m[426])|(~m[74]&m[201]&m[426]))&BiasedRNG[328])|(((m[74]&m[201]&~m[426]))&~BiasedRNG[328])|((m[74]&m[201]&m[426]));
    m[310] = (((m[65]&~m[210]&m[431])|(~m[65]&m[210]&m[431]))&BiasedRNG[329])|(((m[65]&m[210]&~m[431]))&~BiasedRNG[329])|((m[65]&m[210]&m[431]));
    m[311] = (((m[75]&~m[211]&m[456])|(~m[75]&m[211]&m[456]))&BiasedRNG[330])|(((m[75]&m[211]&~m[456]))&~BiasedRNG[330])|((m[75]&m[211]&m[456]));
    m[320] = (((m[66]&~m[220]&m[461])|(~m[66]&m[220]&m[461]))&BiasedRNG[331])|(((m[66]&m[220]&~m[461]))&~BiasedRNG[331])|((m[66]&m[220]&m[461]));
    m[321] = (((m[76]&~m[221]&m[491])|(~m[76]&m[221]&m[491]))&BiasedRNG[332])|(((m[76]&m[221]&~m[491]))&~BiasedRNG[332])|((m[76]&m[221]&m[491]));
    m[330] = (((m[67]&~m[230]&m[496])|(~m[67]&m[230]&m[496]))&BiasedRNG[333])|(((m[67]&m[230]&~m[496]))&~BiasedRNG[333])|((m[67]&m[230]&m[496]));
    m[331] = (((m[77]&~m[231]&m[531])|(~m[77]&m[231]&m[531]))&BiasedRNG[334])|(((m[77]&m[231]&~m[531]))&~BiasedRNG[334])|((m[77]&m[231]&m[531]));
    m[340] = (((m[68]&~m[240]&m[536])|(~m[68]&m[240]&m[536]))&BiasedRNG[335])|(((m[68]&m[240]&~m[536]))&~BiasedRNG[335])|((m[68]&m[240]&m[536]));
    m[341] = (((m[78]&~m[241]&m[576])|(~m[78]&m[241]&m[576]))&BiasedRNG[336])|(((m[78]&m[241]&~m[576]))&~BiasedRNG[336])|((m[78]&m[241]&m[576]));
    m[350] = (((m[69]&~m[250]&m[581])|(~m[69]&m[250]&m[581]))&BiasedRNG[337])|(((m[69]&m[250]&~m[581]))&~BiasedRNG[337])|((m[69]&m[250]&m[581]));
    m[351] = (((m[79]&~m[251]&m[626])|(~m[79]&m[251]&m[626]))&BiasedRNG[338])|(((m[79]&m[251]&~m[626]))&~BiasedRNG[338])|((m[79]&m[251]&m[626]));
    m[361] = (((m[270]&~m[360]&~m[362]&~m[363]&~m[364])|(~m[270]&~m[360]&~m[362]&m[363]&~m[364])|(m[270]&m[360]&~m[362]&m[363]&~m[364])|(m[270]&~m[360]&m[362]&m[363]&~m[364])|(~m[270]&m[360]&~m[362]&~m[363]&m[364])|(~m[270]&~m[360]&m[362]&~m[363]&m[364])|(m[270]&m[360]&m[362]&~m[363]&m[364])|(~m[270]&m[360]&m[362]&m[363]&m[364]))&UnbiasedRNG[198])|((m[270]&~m[360]&~m[362]&m[363]&~m[364])|(~m[270]&~m[360]&~m[362]&~m[363]&m[364])|(m[270]&~m[360]&~m[362]&~m[363]&m[364])|(m[270]&m[360]&~m[362]&~m[363]&m[364])|(m[270]&~m[360]&m[362]&~m[363]&m[364])|(~m[270]&~m[360]&~m[362]&m[363]&m[364])|(m[270]&~m[360]&~m[362]&m[363]&m[364])|(~m[270]&m[360]&~m[362]&m[363]&m[364])|(m[270]&m[360]&~m[362]&m[363]&m[364])|(~m[270]&~m[360]&m[362]&m[363]&m[364])|(m[270]&~m[360]&m[362]&m[363]&m[364])|(m[270]&m[360]&m[362]&m[363]&m[364]));
    m[367] = (((m[364]&~m[365]&~m[366]&~m[368]&~m[369])|(~m[364]&~m[365]&~m[366]&m[368]&~m[369])|(m[364]&m[365]&~m[366]&m[368]&~m[369])|(m[364]&~m[365]&m[366]&m[368]&~m[369])|(~m[364]&m[365]&~m[366]&~m[368]&m[369])|(~m[364]&~m[365]&m[366]&~m[368]&m[369])|(m[364]&m[365]&m[366]&~m[368]&m[369])|(~m[364]&m[365]&m[366]&m[368]&m[369]))&UnbiasedRNG[199])|((m[364]&~m[365]&~m[366]&m[368]&~m[369])|(~m[364]&~m[365]&~m[366]&~m[368]&m[369])|(m[364]&~m[365]&~m[366]&~m[368]&m[369])|(m[364]&m[365]&~m[366]&~m[368]&m[369])|(m[364]&~m[365]&m[366]&~m[368]&m[369])|(~m[364]&~m[365]&~m[366]&m[368]&m[369])|(m[364]&~m[365]&~m[366]&m[368]&m[369])|(~m[364]&m[365]&~m[366]&m[368]&m[369])|(m[364]&m[365]&~m[366]&m[368]&m[369])|(~m[364]&~m[365]&m[366]&m[368]&m[369])|(m[364]&~m[365]&m[366]&m[368]&m[369])|(m[364]&m[365]&m[366]&m[368]&m[369]));
    m[377] = (((m[369]&~m[375]&~m[376]&~m[378]&~m[379])|(~m[369]&~m[375]&~m[376]&m[378]&~m[379])|(m[369]&m[375]&~m[376]&m[378]&~m[379])|(m[369]&~m[375]&m[376]&m[378]&~m[379])|(~m[369]&m[375]&~m[376]&~m[378]&m[379])|(~m[369]&~m[375]&m[376]&~m[378]&m[379])|(m[369]&m[375]&m[376]&~m[378]&m[379])|(~m[369]&m[375]&m[376]&m[378]&m[379]))&UnbiasedRNG[200])|((m[369]&~m[375]&~m[376]&m[378]&~m[379])|(~m[369]&~m[375]&~m[376]&~m[378]&m[379])|(m[369]&~m[375]&~m[376]&~m[378]&m[379])|(m[369]&m[375]&~m[376]&~m[378]&m[379])|(m[369]&~m[375]&m[376]&~m[378]&m[379])|(~m[369]&~m[375]&~m[376]&m[378]&m[379])|(m[369]&~m[375]&~m[376]&m[378]&m[379])|(~m[369]&m[375]&~m[376]&m[378]&m[379])|(m[369]&m[375]&~m[376]&m[378]&m[379])|(~m[369]&~m[375]&m[376]&m[378]&m[379])|(m[369]&~m[375]&m[376]&m[378]&m[379])|(m[369]&m[375]&m[376]&m[378]&m[379]));
    m[382] = (((m[374]&~m[380]&~m[381]&~m[383]&~m[384])|(~m[374]&~m[380]&~m[381]&m[383]&~m[384])|(m[374]&m[380]&~m[381]&m[383]&~m[384])|(m[374]&~m[380]&m[381]&m[383]&~m[384])|(~m[374]&m[380]&~m[381]&~m[383]&m[384])|(~m[374]&~m[380]&m[381]&~m[383]&m[384])|(m[374]&m[380]&m[381]&~m[383]&m[384])|(~m[374]&m[380]&m[381]&m[383]&m[384]))&UnbiasedRNG[201])|((m[374]&~m[380]&~m[381]&m[383]&~m[384])|(~m[374]&~m[380]&~m[381]&~m[383]&m[384])|(m[374]&~m[380]&~m[381]&~m[383]&m[384])|(m[374]&m[380]&~m[381]&~m[383]&m[384])|(m[374]&~m[380]&m[381]&~m[383]&m[384])|(~m[374]&~m[380]&~m[381]&m[383]&m[384])|(m[374]&~m[380]&~m[381]&m[383]&m[384])|(~m[374]&m[380]&~m[381]&m[383]&m[384])|(m[374]&m[380]&~m[381]&m[383]&m[384])|(~m[374]&~m[380]&m[381]&m[383]&m[384])|(m[374]&~m[380]&m[381]&m[383]&m[384])|(m[374]&m[380]&m[381]&m[383]&m[384]));
    m[392] = (((m[379]&~m[390]&~m[391]&~m[393]&~m[394])|(~m[379]&~m[390]&~m[391]&m[393]&~m[394])|(m[379]&m[390]&~m[391]&m[393]&~m[394])|(m[379]&~m[390]&m[391]&m[393]&~m[394])|(~m[379]&m[390]&~m[391]&~m[393]&m[394])|(~m[379]&~m[390]&m[391]&~m[393]&m[394])|(m[379]&m[390]&m[391]&~m[393]&m[394])|(~m[379]&m[390]&m[391]&m[393]&m[394]))&UnbiasedRNG[202])|((m[379]&~m[390]&~m[391]&m[393]&~m[394])|(~m[379]&~m[390]&~m[391]&~m[393]&m[394])|(m[379]&~m[390]&~m[391]&~m[393]&m[394])|(m[379]&m[390]&~m[391]&~m[393]&m[394])|(m[379]&~m[390]&m[391]&~m[393]&m[394])|(~m[379]&~m[390]&~m[391]&m[393]&m[394])|(m[379]&~m[390]&~m[391]&m[393]&m[394])|(~m[379]&m[390]&~m[391]&m[393]&m[394])|(m[379]&m[390]&~m[391]&m[393]&m[394])|(~m[379]&~m[390]&m[391]&m[393]&m[394])|(m[379]&~m[390]&m[391]&m[393]&m[394])|(m[379]&m[390]&m[391]&m[393]&m[394]));
    m[396] = (((m[282]&~m[395]&~m[397]&~m[398]&~m[399])|(~m[282]&~m[395]&~m[397]&m[398]&~m[399])|(m[282]&m[395]&~m[397]&m[398]&~m[399])|(m[282]&~m[395]&m[397]&m[398]&~m[399])|(~m[282]&m[395]&~m[397]&~m[398]&m[399])|(~m[282]&~m[395]&m[397]&~m[398]&m[399])|(m[282]&m[395]&m[397]&~m[398]&m[399])|(~m[282]&m[395]&m[397]&m[398]&m[399]))&UnbiasedRNG[203])|((m[282]&~m[395]&~m[397]&m[398]&~m[399])|(~m[282]&~m[395]&~m[397]&~m[398]&m[399])|(m[282]&~m[395]&~m[397]&~m[398]&m[399])|(m[282]&m[395]&~m[397]&~m[398]&m[399])|(m[282]&~m[395]&m[397]&~m[398]&m[399])|(~m[282]&~m[395]&~m[397]&m[398]&m[399])|(m[282]&~m[395]&~m[397]&m[398]&m[399])|(~m[282]&m[395]&~m[397]&m[398]&m[399])|(m[282]&m[395]&~m[397]&m[398]&m[399])|(~m[282]&~m[395]&m[397]&m[398]&m[399])|(m[282]&~m[395]&m[397]&m[398]&m[399])|(m[282]&m[395]&m[397]&m[398]&m[399]));
    m[402] = (((m[389]&~m[400]&~m[401]&~m[403]&~m[404])|(~m[389]&~m[400]&~m[401]&m[403]&~m[404])|(m[389]&m[400]&~m[401]&m[403]&~m[404])|(m[389]&~m[400]&m[401]&m[403]&~m[404])|(~m[389]&m[400]&~m[401]&~m[403]&m[404])|(~m[389]&~m[400]&m[401]&~m[403]&m[404])|(m[389]&m[400]&m[401]&~m[403]&m[404])|(~m[389]&m[400]&m[401]&m[403]&m[404]))&UnbiasedRNG[204])|((m[389]&~m[400]&~m[401]&m[403]&~m[404])|(~m[389]&~m[400]&~m[401]&~m[403]&m[404])|(m[389]&~m[400]&~m[401]&~m[403]&m[404])|(m[389]&m[400]&~m[401]&~m[403]&m[404])|(m[389]&~m[400]&m[401]&~m[403]&m[404])|(~m[389]&~m[400]&~m[401]&m[403]&m[404])|(m[389]&~m[400]&~m[401]&m[403]&m[404])|(~m[389]&m[400]&~m[401]&m[403]&m[404])|(m[389]&m[400]&~m[401]&m[403]&m[404])|(~m[389]&~m[400]&m[401]&m[403]&m[404])|(m[389]&~m[400]&m[401]&m[403]&m[404])|(m[389]&m[400]&m[401]&m[403]&m[404]));
    m[412] = (((m[394]&~m[410]&~m[411]&~m[413]&~m[414])|(~m[394]&~m[410]&~m[411]&m[413]&~m[414])|(m[394]&m[410]&~m[411]&m[413]&~m[414])|(m[394]&~m[410]&m[411]&m[413]&~m[414])|(~m[394]&m[410]&~m[411]&~m[413]&m[414])|(~m[394]&~m[410]&m[411]&~m[413]&m[414])|(m[394]&m[410]&m[411]&~m[413]&m[414])|(~m[394]&m[410]&m[411]&m[413]&m[414]))&UnbiasedRNG[205])|((m[394]&~m[410]&~m[411]&m[413]&~m[414])|(~m[394]&~m[410]&~m[411]&~m[413]&m[414])|(m[394]&~m[410]&~m[411]&~m[413]&m[414])|(m[394]&m[410]&~m[411]&~m[413]&m[414])|(m[394]&~m[410]&m[411]&~m[413]&m[414])|(~m[394]&~m[410]&~m[411]&m[413]&m[414])|(m[394]&~m[410]&~m[411]&m[413]&m[414])|(~m[394]&m[410]&~m[411]&m[413]&m[414])|(m[394]&m[410]&~m[411]&m[413]&m[414])|(~m[394]&~m[410]&m[411]&m[413]&m[414])|(m[394]&~m[410]&m[411]&m[413]&m[414])|(m[394]&m[410]&m[411]&m[413]&m[414]));
    m[416] = (((m[283]&~m[415]&~m[417]&~m[418]&~m[419])|(~m[283]&~m[415]&~m[417]&m[418]&~m[419])|(m[283]&m[415]&~m[417]&m[418]&~m[419])|(m[283]&~m[415]&m[417]&m[418]&~m[419])|(~m[283]&m[415]&~m[417]&~m[418]&m[419])|(~m[283]&~m[415]&m[417]&~m[418]&m[419])|(m[283]&m[415]&m[417]&~m[418]&m[419])|(~m[283]&m[415]&m[417]&m[418]&m[419]))&UnbiasedRNG[206])|((m[283]&~m[415]&~m[417]&m[418]&~m[419])|(~m[283]&~m[415]&~m[417]&~m[418]&m[419])|(m[283]&~m[415]&~m[417]&~m[418]&m[419])|(m[283]&m[415]&~m[417]&~m[418]&m[419])|(m[283]&~m[415]&m[417]&~m[418]&m[419])|(~m[283]&~m[415]&~m[417]&m[418]&m[419])|(m[283]&~m[415]&~m[417]&m[418]&m[419])|(~m[283]&m[415]&~m[417]&m[418]&m[419])|(m[283]&m[415]&~m[417]&m[418]&m[419])|(~m[283]&~m[415]&m[417]&m[418]&m[419])|(m[283]&~m[415]&m[417]&m[418]&m[419])|(m[283]&m[415]&m[417]&m[418]&m[419]));
    m[421] = (((m[292]&~m[420]&~m[422]&~m[423]&~m[424])|(~m[292]&~m[420]&~m[422]&m[423]&~m[424])|(m[292]&m[420]&~m[422]&m[423]&~m[424])|(m[292]&~m[420]&m[422]&m[423]&~m[424])|(~m[292]&m[420]&~m[422]&~m[423]&m[424])|(~m[292]&~m[420]&m[422]&~m[423]&m[424])|(m[292]&m[420]&m[422]&~m[423]&m[424])|(~m[292]&m[420]&m[422]&m[423]&m[424]))&UnbiasedRNG[207])|((m[292]&~m[420]&~m[422]&m[423]&~m[424])|(~m[292]&~m[420]&~m[422]&~m[423]&m[424])|(m[292]&~m[420]&~m[422]&~m[423]&m[424])|(m[292]&m[420]&~m[422]&~m[423]&m[424])|(m[292]&~m[420]&m[422]&~m[423]&m[424])|(~m[292]&~m[420]&~m[422]&m[423]&m[424])|(m[292]&~m[420]&~m[422]&m[423]&m[424])|(~m[292]&m[420]&~m[422]&m[423]&m[424])|(m[292]&m[420]&~m[422]&m[423]&m[424])|(~m[292]&~m[420]&m[422]&m[423]&m[424])|(m[292]&~m[420]&m[422]&m[423]&m[424])|(m[292]&m[420]&m[422]&m[423]&m[424]));
    m[427] = (((m[409]&~m[425]&~m[426]&~m[428]&~m[429])|(~m[409]&~m[425]&~m[426]&m[428]&~m[429])|(m[409]&m[425]&~m[426]&m[428]&~m[429])|(m[409]&~m[425]&m[426]&m[428]&~m[429])|(~m[409]&m[425]&~m[426]&~m[428]&m[429])|(~m[409]&~m[425]&m[426]&~m[428]&m[429])|(m[409]&m[425]&m[426]&~m[428]&m[429])|(~m[409]&m[425]&m[426]&m[428]&m[429]))&UnbiasedRNG[208])|((m[409]&~m[425]&~m[426]&m[428]&~m[429])|(~m[409]&~m[425]&~m[426]&~m[428]&m[429])|(m[409]&~m[425]&~m[426]&~m[428]&m[429])|(m[409]&m[425]&~m[426]&~m[428]&m[429])|(m[409]&~m[425]&m[426]&~m[428]&m[429])|(~m[409]&~m[425]&~m[426]&m[428]&m[429])|(m[409]&~m[425]&~m[426]&m[428]&m[429])|(~m[409]&m[425]&~m[426]&m[428]&m[429])|(m[409]&m[425]&~m[426]&m[428]&m[429])|(~m[409]&~m[425]&m[426]&m[428]&m[429])|(m[409]&~m[425]&m[426]&m[428]&m[429])|(m[409]&m[425]&m[426]&m[428]&m[429]));
    m[437] = (((m[414]&~m[435]&~m[436]&~m[438]&~m[439])|(~m[414]&~m[435]&~m[436]&m[438]&~m[439])|(m[414]&m[435]&~m[436]&m[438]&~m[439])|(m[414]&~m[435]&m[436]&m[438]&~m[439])|(~m[414]&m[435]&~m[436]&~m[438]&m[439])|(~m[414]&~m[435]&m[436]&~m[438]&m[439])|(m[414]&m[435]&m[436]&~m[438]&m[439])|(~m[414]&m[435]&m[436]&m[438]&m[439]))&UnbiasedRNG[209])|((m[414]&~m[435]&~m[436]&m[438]&~m[439])|(~m[414]&~m[435]&~m[436]&~m[438]&m[439])|(m[414]&~m[435]&~m[436]&~m[438]&m[439])|(m[414]&m[435]&~m[436]&~m[438]&m[439])|(m[414]&~m[435]&m[436]&~m[438]&m[439])|(~m[414]&~m[435]&~m[436]&m[438]&m[439])|(m[414]&~m[435]&~m[436]&m[438]&m[439])|(~m[414]&m[435]&~m[436]&m[438]&m[439])|(m[414]&m[435]&~m[436]&m[438]&m[439])|(~m[414]&~m[435]&m[436]&m[438]&m[439])|(m[414]&~m[435]&m[436]&m[438]&m[439])|(m[414]&m[435]&m[436]&m[438]&m[439]));
    m[441] = (((m[284]&~m[440]&~m[442]&~m[443]&~m[444])|(~m[284]&~m[440]&~m[442]&m[443]&~m[444])|(m[284]&m[440]&~m[442]&m[443]&~m[444])|(m[284]&~m[440]&m[442]&m[443]&~m[444])|(~m[284]&m[440]&~m[442]&~m[443]&m[444])|(~m[284]&~m[440]&m[442]&~m[443]&m[444])|(m[284]&m[440]&m[442]&~m[443]&m[444])|(~m[284]&m[440]&m[442]&m[443]&m[444]))&UnbiasedRNG[210])|((m[284]&~m[440]&~m[442]&m[443]&~m[444])|(~m[284]&~m[440]&~m[442]&~m[443]&m[444])|(m[284]&~m[440]&~m[442]&~m[443]&m[444])|(m[284]&m[440]&~m[442]&~m[443]&m[444])|(m[284]&~m[440]&m[442]&~m[443]&m[444])|(~m[284]&~m[440]&~m[442]&m[443]&m[444])|(m[284]&~m[440]&~m[442]&m[443]&m[444])|(~m[284]&m[440]&~m[442]&m[443]&m[444])|(m[284]&m[440]&~m[442]&m[443]&m[444])|(~m[284]&~m[440]&m[442]&m[443]&m[444])|(m[284]&~m[440]&m[442]&m[443]&m[444])|(m[284]&m[440]&m[442]&m[443]&m[444]));
    m[446] = (((m[293]&~m[445]&~m[447]&~m[448]&~m[449])|(~m[293]&~m[445]&~m[447]&m[448]&~m[449])|(m[293]&m[445]&~m[447]&m[448]&~m[449])|(m[293]&~m[445]&m[447]&m[448]&~m[449])|(~m[293]&m[445]&~m[447]&~m[448]&m[449])|(~m[293]&~m[445]&m[447]&~m[448]&m[449])|(m[293]&m[445]&m[447]&~m[448]&m[449])|(~m[293]&m[445]&m[447]&m[448]&m[449]))&UnbiasedRNG[211])|((m[293]&~m[445]&~m[447]&m[448]&~m[449])|(~m[293]&~m[445]&~m[447]&~m[448]&m[449])|(m[293]&~m[445]&~m[447]&~m[448]&m[449])|(m[293]&m[445]&~m[447]&~m[448]&m[449])|(m[293]&~m[445]&m[447]&~m[448]&m[449])|(~m[293]&~m[445]&~m[447]&m[448]&m[449])|(m[293]&~m[445]&~m[447]&m[448]&m[449])|(~m[293]&m[445]&~m[447]&m[448]&m[449])|(m[293]&m[445]&~m[447]&m[448]&m[449])|(~m[293]&~m[445]&m[447]&m[448]&m[449])|(m[293]&~m[445]&m[447]&m[448]&m[449])|(m[293]&m[445]&m[447]&m[448]&m[449]));
    m[451] = (((m[302]&~m[450]&~m[452]&~m[453]&~m[454])|(~m[302]&~m[450]&~m[452]&m[453]&~m[454])|(m[302]&m[450]&~m[452]&m[453]&~m[454])|(m[302]&~m[450]&m[452]&m[453]&~m[454])|(~m[302]&m[450]&~m[452]&~m[453]&m[454])|(~m[302]&~m[450]&m[452]&~m[453]&m[454])|(m[302]&m[450]&m[452]&~m[453]&m[454])|(~m[302]&m[450]&m[452]&m[453]&m[454]))&UnbiasedRNG[212])|((m[302]&~m[450]&~m[452]&m[453]&~m[454])|(~m[302]&~m[450]&~m[452]&~m[453]&m[454])|(m[302]&~m[450]&~m[452]&~m[453]&m[454])|(m[302]&m[450]&~m[452]&~m[453]&m[454])|(m[302]&~m[450]&m[452]&~m[453]&m[454])|(~m[302]&~m[450]&~m[452]&m[453]&m[454])|(m[302]&~m[450]&~m[452]&m[453]&m[454])|(~m[302]&m[450]&~m[452]&m[453]&m[454])|(m[302]&m[450]&~m[452]&m[453]&m[454])|(~m[302]&~m[450]&m[452]&m[453]&m[454])|(m[302]&~m[450]&m[452]&m[453]&m[454])|(m[302]&m[450]&m[452]&m[453]&m[454]));
    m[457] = (((m[434]&~m[455]&~m[456]&~m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&m[458]&~m[459])|(m[434]&m[455]&~m[456]&m[458]&~m[459])|(m[434]&~m[455]&m[456]&m[458]&~m[459])|(~m[434]&m[455]&~m[456]&~m[458]&m[459])|(~m[434]&~m[455]&m[456]&~m[458]&m[459])|(m[434]&m[455]&m[456]&~m[458]&m[459])|(~m[434]&m[455]&m[456]&m[458]&m[459]))&UnbiasedRNG[213])|((m[434]&~m[455]&~m[456]&m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&m[456]&~m[458]&m[459])|(~m[434]&~m[455]&~m[456]&m[458]&m[459])|(m[434]&~m[455]&~m[456]&m[458]&m[459])|(~m[434]&m[455]&~m[456]&m[458]&m[459])|(m[434]&m[455]&~m[456]&m[458]&m[459])|(~m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&m[455]&m[456]&m[458]&m[459]));
    m[467] = (((m[439]&~m[465]&~m[466]&~m[468]&~m[469])|(~m[439]&~m[465]&~m[466]&m[468]&~m[469])|(m[439]&m[465]&~m[466]&m[468]&~m[469])|(m[439]&~m[465]&m[466]&m[468]&~m[469])|(~m[439]&m[465]&~m[466]&~m[468]&m[469])|(~m[439]&~m[465]&m[466]&~m[468]&m[469])|(m[439]&m[465]&m[466]&~m[468]&m[469])|(~m[439]&m[465]&m[466]&m[468]&m[469]))&UnbiasedRNG[214])|((m[439]&~m[465]&~m[466]&m[468]&~m[469])|(~m[439]&~m[465]&~m[466]&~m[468]&m[469])|(m[439]&~m[465]&~m[466]&~m[468]&m[469])|(m[439]&m[465]&~m[466]&~m[468]&m[469])|(m[439]&~m[465]&m[466]&~m[468]&m[469])|(~m[439]&~m[465]&~m[466]&m[468]&m[469])|(m[439]&~m[465]&~m[466]&m[468]&m[469])|(~m[439]&m[465]&~m[466]&m[468]&m[469])|(m[439]&m[465]&~m[466]&m[468]&m[469])|(~m[439]&~m[465]&m[466]&m[468]&m[469])|(m[439]&~m[465]&m[466]&m[468]&m[469])|(m[439]&m[465]&m[466]&m[468]&m[469]));
    m[471] = (((m[285]&~m[470]&~m[472]&~m[473]&~m[474])|(~m[285]&~m[470]&~m[472]&m[473]&~m[474])|(m[285]&m[470]&~m[472]&m[473]&~m[474])|(m[285]&~m[470]&m[472]&m[473]&~m[474])|(~m[285]&m[470]&~m[472]&~m[473]&m[474])|(~m[285]&~m[470]&m[472]&~m[473]&m[474])|(m[285]&m[470]&m[472]&~m[473]&m[474])|(~m[285]&m[470]&m[472]&m[473]&m[474]))&UnbiasedRNG[215])|((m[285]&~m[470]&~m[472]&m[473]&~m[474])|(~m[285]&~m[470]&~m[472]&~m[473]&m[474])|(m[285]&~m[470]&~m[472]&~m[473]&m[474])|(m[285]&m[470]&~m[472]&~m[473]&m[474])|(m[285]&~m[470]&m[472]&~m[473]&m[474])|(~m[285]&~m[470]&~m[472]&m[473]&m[474])|(m[285]&~m[470]&~m[472]&m[473]&m[474])|(~m[285]&m[470]&~m[472]&m[473]&m[474])|(m[285]&m[470]&~m[472]&m[473]&m[474])|(~m[285]&~m[470]&m[472]&m[473]&m[474])|(m[285]&~m[470]&m[472]&m[473]&m[474])|(m[285]&m[470]&m[472]&m[473]&m[474]));
    m[476] = (((m[294]&~m[475]&~m[477]&~m[478]&~m[479])|(~m[294]&~m[475]&~m[477]&m[478]&~m[479])|(m[294]&m[475]&~m[477]&m[478]&~m[479])|(m[294]&~m[475]&m[477]&m[478]&~m[479])|(~m[294]&m[475]&~m[477]&~m[478]&m[479])|(~m[294]&~m[475]&m[477]&~m[478]&m[479])|(m[294]&m[475]&m[477]&~m[478]&m[479])|(~m[294]&m[475]&m[477]&m[478]&m[479]))&UnbiasedRNG[216])|((m[294]&~m[475]&~m[477]&m[478]&~m[479])|(~m[294]&~m[475]&~m[477]&~m[478]&m[479])|(m[294]&~m[475]&~m[477]&~m[478]&m[479])|(m[294]&m[475]&~m[477]&~m[478]&m[479])|(m[294]&~m[475]&m[477]&~m[478]&m[479])|(~m[294]&~m[475]&~m[477]&m[478]&m[479])|(m[294]&~m[475]&~m[477]&m[478]&m[479])|(~m[294]&m[475]&~m[477]&m[478]&m[479])|(m[294]&m[475]&~m[477]&m[478]&m[479])|(~m[294]&~m[475]&m[477]&m[478]&m[479])|(m[294]&~m[475]&m[477]&m[478]&m[479])|(m[294]&m[475]&m[477]&m[478]&m[479]));
    m[481] = (((m[303]&~m[480]&~m[482]&~m[483]&~m[484])|(~m[303]&~m[480]&~m[482]&m[483]&~m[484])|(m[303]&m[480]&~m[482]&m[483]&~m[484])|(m[303]&~m[480]&m[482]&m[483]&~m[484])|(~m[303]&m[480]&~m[482]&~m[483]&m[484])|(~m[303]&~m[480]&m[482]&~m[483]&m[484])|(m[303]&m[480]&m[482]&~m[483]&m[484])|(~m[303]&m[480]&m[482]&m[483]&m[484]))&UnbiasedRNG[217])|((m[303]&~m[480]&~m[482]&m[483]&~m[484])|(~m[303]&~m[480]&~m[482]&~m[483]&m[484])|(m[303]&~m[480]&~m[482]&~m[483]&m[484])|(m[303]&m[480]&~m[482]&~m[483]&m[484])|(m[303]&~m[480]&m[482]&~m[483]&m[484])|(~m[303]&~m[480]&~m[482]&m[483]&m[484])|(m[303]&~m[480]&~m[482]&m[483]&m[484])|(~m[303]&m[480]&~m[482]&m[483]&m[484])|(m[303]&m[480]&~m[482]&m[483]&m[484])|(~m[303]&~m[480]&m[482]&m[483]&m[484])|(m[303]&~m[480]&m[482]&m[483]&m[484])|(m[303]&m[480]&m[482]&m[483]&m[484]));
    m[486] = (((m[312]&~m[485]&~m[487]&~m[488]&~m[489])|(~m[312]&~m[485]&~m[487]&m[488]&~m[489])|(m[312]&m[485]&~m[487]&m[488]&~m[489])|(m[312]&~m[485]&m[487]&m[488]&~m[489])|(~m[312]&m[485]&~m[487]&~m[488]&m[489])|(~m[312]&~m[485]&m[487]&~m[488]&m[489])|(m[312]&m[485]&m[487]&~m[488]&m[489])|(~m[312]&m[485]&m[487]&m[488]&m[489]))&UnbiasedRNG[218])|((m[312]&~m[485]&~m[487]&m[488]&~m[489])|(~m[312]&~m[485]&~m[487]&~m[488]&m[489])|(m[312]&~m[485]&~m[487]&~m[488]&m[489])|(m[312]&m[485]&~m[487]&~m[488]&m[489])|(m[312]&~m[485]&m[487]&~m[488]&m[489])|(~m[312]&~m[485]&~m[487]&m[488]&m[489])|(m[312]&~m[485]&~m[487]&m[488]&m[489])|(~m[312]&m[485]&~m[487]&m[488]&m[489])|(m[312]&m[485]&~m[487]&m[488]&m[489])|(~m[312]&~m[485]&m[487]&m[488]&m[489])|(m[312]&~m[485]&m[487]&m[488]&m[489])|(m[312]&m[485]&m[487]&m[488]&m[489]));
    m[492] = (((m[464]&~m[490]&~m[491]&~m[493]&~m[494])|(~m[464]&~m[490]&~m[491]&m[493]&~m[494])|(m[464]&m[490]&~m[491]&m[493]&~m[494])|(m[464]&~m[490]&m[491]&m[493]&~m[494])|(~m[464]&m[490]&~m[491]&~m[493]&m[494])|(~m[464]&~m[490]&m[491]&~m[493]&m[494])|(m[464]&m[490]&m[491]&~m[493]&m[494])|(~m[464]&m[490]&m[491]&m[493]&m[494]))&UnbiasedRNG[219])|((m[464]&~m[490]&~m[491]&m[493]&~m[494])|(~m[464]&~m[490]&~m[491]&~m[493]&m[494])|(m[464]&~m[490]&~m[491]&~m[493]&m[494])|(m[464]&m[490]&~m[491]&~m[493]&m[494])|(m[464]&~m[490]&m[491]&~m[493]&m[494])|(~m[464]&~m[490]&~m[491]&m[493]&m[494])|(m[464]&~m[490]&~m[491]&m[493]&m[494])|(~m[464]&m[490]&~m[491]&m[493]&m[494])|(m[464]&m[490]&~m[491]&m[493]&m[494])|(~m[464]&~m[490]&m[491]&m[493]&m[494])|(m[464]&~m[490]&m[491]&m[493]&m[494])|(m[464]&m[490]&m[491]&m[493]&m[494]));
    m[502] = (((m[469]&~m[500]&~m[501]&~m[503]&~m[504])|(~m[469]&~m[500]&~m[501]&m[503]&~m[504])|(m[469]&m[500]&~m[501]&m[503]&~m[504])|(m[469]&~m[500]&m[501]&m[503]&~m[504])|(~m[469]&m[500]&~m[501]&~m[503]&m[504])|(~m[469]&~m[500]&m[501]&~m[503]&m[504])|(m[469]&m[500]&m[501]&~m[503]&m[504])|(~m[469]&m[500]&m[501]&m[503]&m[504]))&UnbiasedRNG[220])|((m[469]&~m[500]&~m[501]&m[503]&~m[504])|(~m[469]&~m[500]&~m[501]&~m[503]&m[504])|(m[469]&~m[500]&~m[501]&~m[503]&m[504])|(m[469]&m[500]&~m[501]&~m[503]&m[504])|(m[469]&~m[500]&m[501]&~m[503]&m[504])|(~m[469]&~m[500]&~m[501]&m[503]&m[504])|(m[469]&~m[500]&~m[501]&m[503]&m[504])|(~m[469]&m[500]&~m[501]&m[503]&m[504])|(m[469]&m[500]&~m[501]&m[503]&m[504])|(~m[469]&~m[500]&m[501]&m[503]&m[504])|(m[469]&~m[500]&m[501]&m[503]&m[504])|(m[469]&m[500]&m[501]&m[503]&m[504]));
    m[506] = (((m[286]&~m[505]&~m[507]&~m[508]&~m[509])|(~m[286]&~m[505]&~m[507]&m[508]&~m[509])|(m[286]&m[505]&~m[507]&m[508]&~m[509])|(m[286]&~m[505]&m[507]&m[508]&~m[509])|(~m[286]&m[505]&~m[507]&~m[508]&m[509])|(~m[286]&~m[505]&m[507]&~m[508]&m[509])|(m[286]&m[505]&m[507]&~m[508]&m[509])|(~m[286]&m[505]&m[507]&m[508]&m[509]))&UnbiasedRNG[221])|((m[286]&~m[505]&~m[507]&m[508]&~m[509])|(~m[286]&~m[505]&~m[507]&~m[508]&m[509])|(m[286]&~m[505]&~m[507]&~m[508]&m[509])|(m[286]&m[505]&~m[507]&~m[508]&m[509])|(m[286]&~m[505]&m[507]&~m[508]&m[509])|(~m[286]&~m[505]&~m[507]&m[508]&m[509])|(m[286]&~m[505]&~m[507]&m[508]&m[509])|(~m[286]&m[505]&~m[507]&m[508]&m[509])|(m[286]&m[505]&~m[507]&m[508]&m[509])|(~m[286]&~m[505]&m[507]&m[508]&m[509])|(m[286]&~m[505]&m[507]&m[508]&m[509])|(m[286]&m[505]&m[507]&m[508]&m[509]));
    m[511] = (((m[295]&~m[510]&~m[512]&~m[513]&~m[514])|(~m[295]&~m[510]&~m[512]&m[513]&~m[514])|(m[295]&m[510]&~m[512]&m[513]&~m[514])|(m[295]&~m[510]&m[512]&m[513]&~m[514])|(~m[295]&m[510]&~m[512]&~m[513]&m[514])|(~m[295]&~m[510]&m[512]&~m[513]&m[514])|(m[295]&m[510]&m[512]&~m[513]&m[514])|(~m[295]&m[510]&m[512]&m[513]&m[514]))&UnbiasedRNG[222])|((m[295]&~m[510]&~m[512]&m[513]&~m[514])|(~m[295]&~m[510]&~m[512]&~m[513]&m[514])|(m[295]&~m[510]&~m[512]&~m[513]&m[514])|(m[295]&m[510]&~m[512]&~m[513]&m[514])|(m[295]&~m[510]&m[512]&~m[513]&m[514])|(~m[295]&~m[510]&~m[512]&m[513]&m[514])|(m[295]&~m[510]&~m[512]&m[513]&m[514])|(~m[295]&m[510]&~m[512]&m[513]&m[514])|(m[295]&m[510]&~m[512]&m[513]&m[514])|(~m[295]&~m[510]&m[512]&m[513]&m[514])|(m[295]&~m[510]&m[512]&m[513]&m[514])|(m[295]&m[510]&m[512]&m[513]&m[514]));
    m[516] = (((m[304]&~m[515]&~m[517]&~m[518]&~m[519])|(~m[304]&~m[515]&~m[517]&m[518]&~m[519])|(m[304]&m[515]&~m[517]&m[518]&~m[519])|(m[304]&~m[515]&m[517]&m[518]&~m[519])|(~m[304]&m[515]&~m[517]&~m[518]&m[519])|(~m[304]&~m[515]&m[517]&~m[518]&m[519])|(m[304]&m[515]&m[517]&~m[518]&m[519])|(~m[304]&m[515]&m[517]&m[518]&m[519]))&UnbiasedRNG[223])|((m[304]&~m[515]&~m[517]&m[518]&~m[519])|(~m[304]&~m[515]&~m[517]&~m[518]&m[519])|(m[304]&~m[515]&~m[517]&~m[518]&m[519])|(m[304]&m[515]&~m[517]&~m[518]&m[519])|(m[304]&~m[515]&m[517]&~m[518]&m[519])|(~m[304]&~m[515]&~m[517]&m[518]&m[519])|(m[304]&~m[515]&~m[517]&m[518]&m[519])|(~m[304]&m[515]&~m[517]&m[518]&m[519])|(m[304]&m[515]&~m[517]&m[518]&m[519])|(~m[304]&~m[515]&m[517]&m[518]&m[519])|(m[304]&~m[515]&m[517]&m[518]&m[519])|(m[304]&m[515]&m[517]&m[518]&m[519]));
    m[521] = (((m[313]&~m[520]&~m[522]&~m[523]&~m[524])|(~m[313]&~m[520]&~m[522]&m[523]&~m[524])|(m[313]&m[520]&~m[522]&m[523]&~m[524])|(m[313]&~m[520]&m[522]&m[523]&~m[524])|(~m[313]&m[520]&~m[522]&~m[523]&m[524])|(~m[313]&~m[520]&m[522]&~m[523]&m[524])|(m[313]&m[520]&m[522]&~m[523]&m[524])|(~m[313]&m[520]&m[522]&m[523]&m[524]))&UnbiasedRNG[224])|((m[313]&~m[520]&~m[522]&m[523]&~m[524])|(~m[313]&~m[520]&~m[522]&~m[523]&m[524])|(m[313]&~m[520]&~m[522]&~m[523]&m[524])|(m[313]&m[520]&~m[522]&~m[523]&m[524])|(m[313]&~m[520]&m[522]&~m[523]&m[524])|(~m[313]&~m[520]&~m[522]&m[523]&m[524])|(m[313]&~m[520]&~m[522]&m[523]&m[524])|(~m[313]&m[520]&~m[522]&m[523]&m[524])|(m[313]&m[520]&~m[522]&m[523]&m[524])|(~m[313]&~m[520]&m[522]&m[523]&m[524])|(m[313]&~m[520]&m[522]&m[523]&m[524])|(m[313]&m[520]&m[522]&m[523]&m[524]));
    m[526] = (((m[322]&~m[525]&~m[527]&~m[528]&~m[529])|(~m[322]&~m[525]&~m[527]&m[528]&~m[529])|(m[322]&m[525]&~m[527]&m[528]&~m[529])|(m[322]&~m[525]&m[527]&m[528]&~m[529])|(~m[322]&m[525]&~m[527]&~m[528]&m[529])|(~m[322]&~m[525]&m[527]&~m[528]&m[529])|(m[322]&m[525]&m[527]&~m[528]&m[529])|(~m[322]&m[525]&m[527]&m[528]&m[529]))&UnbiasedRNG[225])|((m[322]&~m[525]&~m[527]&m[528]&~m[529])|(~m[322]&~m[525]&~m[527]&~m[528]&m[529])|(m[322]&~m[525]&~m[527]&~m[528]&m[529])|(m[322]&m[525]&~m[527]&~m[528]&m[529])|(m[322]&~m[525]&m[527]&~m[528]&m[529])|(~m[322]&~m[525]&~m[527]&m[528]&m[529])|(m[322]&~m[525]&~m[527]&m[528]&m[529])|(~m[322]&m[525]&~m[527]&m[528]&m[529])|(m[322]&m[525]&~m[527]&m[528]&m[529])|(~m[322]&~m[525]&m[527]&m[528]&m[529])|(m[322]&~m[525]&m[527]&m[528]&m[529])|(m[322]&m[525]&m[527]&m[528]&m[529]));
    m[532] = (((m[499]&~m[530]&~m[531]&~m[533]&~m[534])|(~m[499]&~m[530]&~m[531]&m[533]&~m[534])|(m[499]&m[530]&~m[531]&m[533]&~m[534])|(m[499]&~m[530]&m[531]&m[533]&~m[534])|(~m[499]&m[530]&~m[531]&~m[533]&m[534])|(~m[499]&~m[530]&m[531]&~m[533]&m[534])|(m[499]&m[530]&m[531]&~m[533]&m[534])|(~m[499]&m[530]&m[531]&m[533]&m[534]))&UnbiasedRNG[226])|((m[499]&~m[530]&~m[531]&m[533]&~m[534])|(~m[499]&~m[530]&~m[531]&~m[533]&m[534])|(m[499]&~m[530]&~m[531]&~m[533]&m[534])|(m[499]&m[530]&~m[531]&~m[533]&m[534])|(m[499]&~m[530]&m[531]&~m[533]&m[534])|(~m[499]&~m[530]&~m[531]&m[533]&m[534])|(m[499]&~m[530]&~m[531]&m[533]&m[534])|(~m[499]&m[530]&~m[531]&m[533]&m[534])|(m[499]&m[530]&~m[531]&m[533]&m[534])|(~m[499]&~m[530]&m[531]&m[533]&m[534])|(m[499]&~m[530]&m[531]&m[533]&m[534])|(m[499]&m[530]&m[531]&m[533]&m[534]));
    m[542] = (((m[504]&~m[540]&~m[541]&~m[543]&~m[544])|(~m[504]&~m[540]&~m[541]&m[543]&~m[544])|(m[504]&m[540]&~m[541]&m[543]&~m[544])|(m[504]&~m[540]&m[541]&m[543]&~m[544])|(~m[504]&m[540]&~m[541]&~m[543]&m[544])|(~m[504]&~m[540]&m[541]&~m[543]&m[544])|(m[504]&m[540]&m[541]&~m[543]&m[544])|(~m[504]&m[540]&m[541]&m[543]&m[544]))&UnbiasedRNG[227])|((m[504]&~m[540]&~m[541]&m[543]&~m[544])|(~m[504]&~m[540]&~m[541]&~m[543]&m[544])|(m[504]&~m[540]&~m[541]&~m[543]&m[544])|(m[504]&m[540]&~m[541]&~m[543]&m[544])|(m[504]&~m[540]&m[541]&~m[543]&m[544])|(~m[504]&~m[540]&~m[541]&m[543]&m[544])|(m[504]&~m[540]&~m[541]&m[543]&m[544])|(~m[504]&m[540]&~m[541]&m[543]&m[544])|(m[504]&m[540]&~m[541]&m[543]&m[544])|(~m[504]&~m[540]&m[541]&m[543]&m[544])|(m[504]&~m[540]&m[541]&m[543]&m[544])|(m[504]&m[540]&m[541]&m[543]&m[544]));
    m[546] = (((m[287]&~m[545]&~m[547]&~m[548]&~m[549])|(~m[287]&~m[545]&~m[547]&m[548]&~m[549])|(m[287]&m[545]&~m[547]&m[548]&~m[549])|(m[287]&~m[545]&m[547]&m[548]&~m[549])|(~m[287]&m[545]&~m[547]&~m[548]&m[549])|(~m[287]&~m[545]&m[547]&~m[548]&m[549])|(m[287]&m[545]&m[547]&~m[548]&m[549])|(~m[287]&m[545]&m[547]&m[548]&m[549]))&UnbiasedRNG[228])|((m[287]&~m[545]&~m[547]&m[548]&~m[549])|(~m[287]&~m[545]&~m[547]&~m[548]&m[549])|(m[287]&~m[545]&~m[547]&~m[548]&m[549])|(m[287]&m[545]&~m[547]&~m[548]&m[549])|(m[287]&~m[545]&m[547]&~m[548]&m[549])|(~m[287]&~m[545]&~m[547]&m[548]&m[549])|(m[287]&~m[545]&~m[547]&m[548]&m[549])|(~m[287]&m[545]&~m[547]&m[548]&m[549])|(m[287]&m[545]&~m[547]&m[548]&m[549])|(~m[287]&~m[545]&m[547]&m[548]&m[549])|(m[287]&~m[545]&m[547]&m[548]&m[549])|(m[287]&m[545]&m[547]&m[548]&m[549]));
    m[551] = (((m[296]&~m[550]&~m[552]&~m[553]&~m[554])|(~m[296]&~m[550]&~m[552]&m[553]&~m[554])|(m[296]&m[550]&~m[552]&m[553]&~m[554])|(m[296]&~m[550]&m[552]&m[553]&~m[554])|(~m[296]&m[550]&~m[552]&~m[553]&m[554])|(~m[296]&~m[550]&m[552]&~m[553]&m[554])|(m[296]&m[550]&m[552]&~m[553]&m[554])|(~m[296]&m[550]&m[552]&m[553]&m[554]))&UnbiasedRNG[229])|((m[296]&~m[550]&~m[552]&m[553]&~m[554])|(~m[296]&~m[550]&~m[552]&~m[553]&m[554])|(m[296]&~m[550]&~m[552]&~m[553]&m[554])|(m[296]&m[550]&~m[552]&~m[553]&m[554])|(m[296]&~m[550]&m[552]&~m[553]&m[554])|(~m[296]&~m[550]&~m[552]&m[553]&m[554])|(m[296]&~m[550]&~m[552]&m[553]&m[554])|(~m[296]&m[550]&~m[552]&m[553]&m[554])|(m[296]&m[550]&~m[552]&m[553]&m[554])|(~m[296]&~m[550]&m[552]&m[553]&m[554])|(m[296]&~m[550]&m[552]&m[553]&m[554])|(m[296]&m[550]&m[552]&m[553]&m[554]));
    m[556] = (((m[305]&~m[555]&~m[557]&~m[558]&~m[559])|(~m[305]&~m[555]&~m[557]&m[558]&~m[559])|(m[305]&m[555]&~m[557]&m[558]&~m[559])|(m[305]&~m[555]&m[557]&m[558]&~m[559])|(~m[305]&m[555]&~m[557]&~m[558]&m[559])|(~m[305]&~m[555]&m[557]&~m[558]&m[559])|(m[305]&m[555]&m[557]&~m[558]&m[559])|(~m[305]&m[555]&m[557]&m[558]&m[559]))&UnbiasedRNG[230])|((m[305]&~m[555]&~m[557]&m[558]&~m[559])|(~m[305]&~m[555]&~m[557]&~m[558]&m[559])|(m[305]&~m[555]&~m[557]&~m[558]&m[559])|(m[305]&m[555]&~m[557]&~m[558]&m[559])|(m[305]&~m[555]&m[557]&~m[558]&m[559])|(~m[305]&~m[555]&~m[557]&m[558]&m[559])|(m[305]&~m[555]&~m[557]&m[558]&m[559])|(~m[305]&m[555]&~m[557]&m[558]&m[559])|(m[305]&m[555]&~m[557]&m[558]&m[559])|(~m[305]&~m[555]&m[557]&m[558]&m[559])|(m[305]&~m[555]&m[557]&m[558]&m[559])|(m[305]&m[555]&m[557]&m[558]&m[559]));
    m[561] = (((m[314]&~m[560]&~m[562]&~m[563]&~m[564])|(~m[314]&~m[560]&~m[562]&m[563]&~m[564])|(m[314]&m[560]&~m[562]&m[563]&~m[564])|(m[314]&~m[560]&m[562]&m[563]&~m[564])|(~m[314]&m[560]&~m[562]&~m[563]&m[564])|(~m[314]&~m[560]&m[562]&~m[563]&m[564])|(m[314]&m[560]&m[562]&~m[563]&m[564])|(~m[314]&m[560]&m[562]&m[563]&m[564]))&UnbiasedRNG[231])|((m[314]&~m[560]&~m[562]&m[563]&~m[564])|(~m[314]&~m[560]&~m[562]&~m[563]&m[564])|(m[314]&~m[560]&~m[562]&~m[563]&m[564])|(m[314]&m[560]&~m[562]&~m[563]&m[564])|(m[314]&~m[560]&m[562]&~m[563]&m[564])|(~m[314]&~m[560]&~m[562]&m[563]&m[564])|(m[314]&~m[560]&~m[562]&m[563]&m[564])|(~m[314]&m[560]&~m[562]&m[563]&m[564])|(m[314]&m[560]&~m[562]&m[563]&m[564])|(~m[314]&~m[560]&m[562]&m[563]&m[564])|(m[314]&~m[560]&m[562]&m[563]&m[564])|(m[314]&m[560]&m[562]&m[563]&m[564]));
    m[566] = (((m[323]&~m[565]&~m[567]&~m[568]&~m[569])|(~m[323]&~m[565]&~m[567]&m[568]&~m[569])|(m[323]&m[565]&~m[567]&m[568]&~m[569])|(m[323]&~m[565]&m[567]&m[568]&~m[569])|(~m[323]&m[565]&~m[567]&~m[568]&m[569])|(~m[323]&~m[565]&m[567]&~m[568]&m[569])|(m[323]&m[565]&m[567]&~m[568]&m[569])|(~m[323]&m[565]&m[567]&m[568]&m[569]))&UnbiasedRNG[232])|((m[323]&~m[565]&~m[567]&m[568]&~m[569])|(~m[323]&~m[565]&~m[567]&~m[568]&m[569])|(m[323]&~m[565]&~m[567]&~m[568]&m[569])|(m[323]&m[565]&~m[567]&~m[568]&m[569])|(m[323]&~m[565]&m[567]&~m[568]&m[569])|(~m[323]&~m[565]&~m[567]&m[568]&m[569])|(m[323]&~m[565]&~m[567]&m[568]&m[569])|(~m[323]&m[565]&~m[567]&m[568]&m[569])|(m[323]&m[565]&~m[567]&m[568]&m[569])|(~m[323]&~m[565]&m[567]&m[568]&m[569])|(m[323]&~m[565]&m[567]&m[568]&m[569])|(m[323]&m[565]&m[567]&m[568]&m[569]));
    m[571] = (((m[332]&~m[570]&~m[572]&~m[573]&~m[574])|(~m[332]&~m[570]&~m[572]&m[573]&~m[574])|(m[332]&m[570]&~m[572]&m[573]&~m[574])|(m[332]&~m[570]&m[572]&m[573]&~m[574])|(~m[332]&m[570]&~m[572]&~m[573]&m[574])|(~m[332]&~m[570]&m[572]&~m[573]&m[574])|(m[332]&m[570]&m[572]&~m[573]&m[574])|(~m[332]&m[570]&m[572]&m[573]&m[574]))&UnbiasedRNG[233])|((m[332]&~m[570]&~m[572]&m[573]&~m[574])|(~m[332]&~m[570]&~m[572]&~m[573]&m[574])|(m[332]&~m[570]&~m[572]&~m[573]&m[574])|(m[332]&m[570]&~m[572]&~m[573]&m[574])|(m[332]&~m[570]&m[572]&~m[573]&m[574])|(~m[332]&~m[570]&~m[572]&m[573]&m[574])|(m[332]&~m[570]&~m[572]&m[573]&m[574])|(~m[332]&m[570]&~m[572]&m[573]&m[574])|(m[332]&m[570]&~m[572]&m[573]&m[574])|(~m[332]&~m[570]&m[572]&m[573]&m[574])|(m[332]&~m[570]&m[572]&m[573]&m[574])|(m[332]&m[570]&m[572]&m[573]&m[574]));
    m[577] = (((m[539]&~m[575]&~m[576]&~m[578]&~m[579])|(~m[539]&~m[575]&~m[576]&m[578]&~m[579])|(m[539]&m[575]&~m[576]&m[578]&~m[579])|(m[539]&~m[575]&m[576]&m[578]&~m[579])|(~m[539]&m[575]&~m[576]&~m[578]&m[579])|(~m[539]&~m[575]&m[576]&~m[578]&m[579])|(m[539]&m[575]&m[576]&~m[578]&m[579])|(~m[539]&m[575]&m[576]&m[578]&m[579]))&UnbiasedRNG[234])|((m[539]&~m[575]&~m[576]&m[578]&~m[579])|(~m[539]&~m[575]&~m[576]&~m[578]&m[579])|(m[539]&~m[575]&~m[576]&~m[578]&m[579])|(m[539]&m[575]&~m[576]&~m[578]&m[579])|(m[539]&~m[575]&m[576]&~m[578]&m[579])|(~m[539]&~m[575]&~m[576]&m[578]&m[579])|(m[539]&~m[575]&~m[576]&m[578]&m[579])|(~m[539]&m[575]&~m[576]&m[578]&m[579])|(m[539]&m[575]&~m[576]&m[578]&m[579])|(~m[539]&~m[575]&m[576]&m[578]&m[579])|(m[539]&~m[575]&m[576]&m[578]&m[579])|(m[539]&m[575]&m[576]&m[578]&m[579]));
    m[587] = (((m[544]&~m[585]&~m[586]&~m[588]&~m[589])|(~m[544]&~m[585]&~m[586]&m[588]&~m[589])|(m[544]&m[585]&~m[586]&m[588]&~m[589])|(m[544]&~m[585]&m[586]&m[588]&~m[589])|(~m[544]&m[585]&~m[586]&~m[588]&m[589])|(~m[544]&~m[585]&m[586]&~m[588]&m[589])|(m[544]&m[585]&m[586]&~m[588]&m[589])|(~m[544]&m[585]&m[586]&m[588]&m[589]))&UnbiasedRNG[235])|((m[544]&~m[585]&~m[586]&m[588]&~m[589])|(~m[544]&~m[585]&~m[586]&~m[588]&m[589])|(m[544]&~m[585]&~m[586]&~m[588]&m[589])|(m[544]&m[585]&~m[586]&~m[588]&m[589])|(m[544]&~m[585]&m[586]&~m[588]&m[589])|(~m[544]&~m[585]&~m[586]&m[588]&m[589])|(m[544]&~m[585]&~m[586]&m[588]&m[589])|(~m[544]&m[585]&~m[586]&m[588]&m[589])|(m[544]&m[585]&~m[586]&m[588]&m[589])|(~m[544]&~m[585]&m[586]&m[588]&m[589])|(m[544]&~m[585]&m[586]&m[588]&m[589])|(m[544]&m[585]&m[586]&m[588]&m[589]));
    m[591] = (((m[288]&~m[590]&~m[592]&~m[593]&~m[594])|(~m[288]&~m[590]&~m[592]&m[593]&~m[594])|(m[288]&m[590]&~m[592]&m[593]&~m[594])|(m[288]&~m[590]&m[592]&m[593]&~m[594])|(~m[288]&m[590]&~m[592]&~m[593]&m[594])|(~m[288]&~m[590]&m[592]&~m[593]&m[594])|(m[288]&m[590]&m[592]&~m[593]&m[594])|(~m[288]&m[590]&m[592]&m[593]&m[594]))&UnbiasedRNG[236])|((m[288]&~m[590]&~m[592]&m[593]&~m[594])|(~m[288]&~m[590]&~m[592]&~m[593]&m[594])|(m[288]&~m[590]&~m[592]&~m[593]&m[594])|(m[288]&m[590]&~m[592]&~m[593]&m[594])|(m[288]&~m[590]&m[592]&~m[593]&m[594])|(~m[288]&~m[590]&~m[592]&m[593]&m[594])|(m[288]&~m[590]&~m[592]&m[593]&m[594])|(~m[288]&m[590]&~m[592]&m[593]&m[594])|(m[288]&m[590]&~m[592]&m[593]&m[594])|(~m[288]&~m[590]&m[592]&m[593]&m[594])|(m[288]&~m[590]&m[592]&m[593]&m[594])|(m[288]&m[590]&m[592]&m[593]&m[594]));
    m[596] = (((m[297]&~m[595]&~m[597]&~m[598]&~m[599])|(~m[297]&~m[595]&~m[597]&m[598]&~m[599])|(m[297]&m[595]&~m[597]&m[598]&~m[599])|(m[297]&~m[595]&m[597]&m[598]&~m[599])|(~m[297]&m[595]&~m[597]&~m[598]&m[599])|(~m[297]&~m[595]&m[597]&~m[598]&m[599])|(m[297]&m[595]&m[597]&~m[598]&m[599])|(~m[297]&m[595]&m[597]&m[598]&m[599]))&UnbiasedRNG[237])|((m[297]&~m[595]&~m[597]&m[598]&~m[599])|(~m[297]&~m[595]&~m[597]&~m[598]&m[599])|(m[297]&~m[595]&~m[597]&~m[598]&m[599])|(m[297]&m[595]&~m[597]&~m[598]&m[599])|(m[297]&~m[595]&m[597]&~m[598]&m[599])|(~m[297]&~m[595]&~m[597]&m[598]&m[599])|(m[297]&~m[595]&~m[597]&m[598]&m[599])|(~m[297]&m[595]&~m[597]&m[598]&m[599])|(m[297]&m[595]&~m[597]&m[598]&m[599])|(~m[297]&~m[595]&m[597]&m[598]&m[599])|(m[297]&~m[595]&m[597]&m[598]&m[599])|(m[297]&m[595]&m[597]&m[598]&m[599]));
    m[601] = (((m[306]&~m[600]&~m[602]&~m[603]&~m[604])|(~m[306]&~m[600]&~m[602]&m[603]&~m[604])|(m[306]&m[600]&~m[602]&m[603]&~m[604])|(m[306]&~m[600]&m[602]&m[603]&~m[604])|(~m[306]&m[600]&~m[602]&~m[603]&m[604])|(~m[306]&~m[600]&m[602]&~m[603]&m[604])|(m[306]&m[600]&m[602]&~m[603]&m[604])|(~m[306]&m[600]&m[602]&m[603]&m[604]))&UnbiasedRNG[238])|((m[306]&~m[600]&~m[602]&m[603]&~m[604])|(~m[306]&~m[600]&~m[602]&~m[603]&m[604])|(m[306]&~m[600]&~m[602]&~m[603]&m[604])|(m[306]&m[600]&~m[602]&~m[603]&m[604])|(m[306]&~m[600]&m[602]&~m[603]&m[604])|(~m[306]&~m[600]&~m[602]&m[603]&m[604])|(m[306]&~m[600]&~m[602]&m[603]&m[604])|(~m[306]&m[600]&~m[602]&m[603]&m[604])|(m[306]&m[600]&~m[602]&m[603]&m[604])|(~m[306]&~m[600]&m[602]&m[603]&m[604])|(m[306]&~m[600]&m[602]&m[603]&m[604])|(m[306]&m[600]&m[602]&m[603]&m[604]));
    m[606] = (((m[315]&~m[605]&~m[607]&~m[608]&~m[609])|(~m[315]&~m[605]&~m[607]&m[608]&~m[609])|(m[315]&m[605]&~m[607]&m[608]&~m[609])|(m[315]&~m[605]&m[607]&m[608]&~m[609])|(~m[315]&m[605]&~m[607]&~m[608]&m[609])|(~m[315]&~m[605]&m[607]&~m[608]&m[609])|(m[315]&m[605]&m[607]&~m[608]&m[609])|(~m[315]&m[605]&m[607]&m[608]&m[609]))&UnbiasedRNG[239])|((m[315]&~m[605]&~m[607]&m[608]&~m[609])|(~m[315]&~m[605]&~m[607]&~m[608]&m[609])|(m[315]&~m[605]&~m[607]&~m[608]&m[609])|(m[315]&m[605]&~m[607]&~m[608]&m[609])|(m[315]&~m[605]&m[607]&~m[608]&m[609])|(~m[315]&~m[605]&~m[607]&m[608]&m[609])|(m[315]&~m[605]&~m[607]&m[608]&m[609])|(~m[315]&m[605]&~m[607]&m[608]&m[609])|(m[315]&m[605]&~m[607]&m[608]&m[609])|(~m[315]&~m[605]&m[607]&m[608]&m[609])|(m[315]&~m[605]&m[607]&m[608]&m[609])|(m[315]&m[605]&m[607]&m[608]&m[609]));
    m[611] = (((m[324]&~m[610]&~m[612]&~m[613]&~m[614])|(~m[324]&~m[610]&~m[612]&m[613]&~m[614])|(m[324]&m[610]&~m[612]&m[613]&~m[614])|(m[324]&~m[610]&m[612]&m[613]&~m[614])|(~m[324]&m[610]&~m[612]&~m[613]&m[614])|(~m[324]&~m[610]&m[612]&~m[613]&m[614])|(m[324]&m[610]&m[612]&~m[613]&m[614])|(~m[324]&m[610]&m[612]&m[613]&m[614]))&UnbiasedRNG[240])|((m[324]&~m[610]&~m[612]&m[613]&~m[614])|(~m[324]&~m[610]&~m[612]&~m[613]&m[614])|(m[324]&~m[610]&~m[612]&~m[613]&m[614])|(m[324]&m[610]&~m[612]&~m[613]&m[614])|(m[324]&~m[610]&m[612]&~m[613]&m[614])|(~m[324]&~m[610]&~m[612]&m[613]&m[614])|(m[324]&~m[610]&~m[612]&m[613]&m[614])|(~m[324]&m[610]&~m[612]&m[613]&m[614])|(m[324]&m[610]&~m[612]&m[613]&m[614])|(~m[324]&~m[610]&m[612]&m[613]&m[614])|(m[324]&~m[610]&m[612]&m[613]&m[614])|(m[324]&m[610]&m[612]&m[613]&m[614]));
    m[616] = (((m[333]&~m[615]&~m[617]&~m[618]&~m[619])|(~m[333]&~m[615]&~m[617]&m[618]&~m[619])|(m[333]&m[615]&~m[617]&m[618]&~m[619])|(m[333]&~m[615]&m[617]&m[618]&~m[619])|(~m[333]&m[615]&~m[617]&~m[618]&m[619])|(~m[333]&~m[615]&m[617]&~m[618]&m[619])|(m[333]&m[615]&m[617]&~m[618]&m[619])|(~m[333]&m[615]&m[617]&m[618]&m[619]))&UnbiasedRNG[241])|((m[333]&~m[615]&~m[617]&m[618]&~m[619])|(~m[333]&~m[615]&~m[617]&~m[618]&m[619])|(m[333]&~m[615]&~m[617]&~m[618]&m[619])|(m[333]&m[615]&~m[617]&~m[618]&m[619])|(m[333]&~m[615]&m[617]&~m[618]&m[619])|(~m[333]&~m[615]&~m[617]&m[618]&m[619])|(m[333]&~m[615]&~m[617]&m[618]&m[619])|(~m[333]&m[615]&~m[617]&m[618]&m[619])|(m[333]&m[615]&~m[617]&m[618]&m[619])|(~m[333]&~m[615]&m[617]&m[618]&m[619])|(m[333]&~m[615]&m[617]&m[618]&m[619])|(m[333]&m[615]&m[617]&m[618]&m[619]));
    m[621] = (((m[342]&~m[620]&~m[622]&~m[623]&~m[624])|(~m[342]&~m[620]&~m[622]&m[623]&~m[624])|(m[342]&m[620]&~m[622]&m[623]&~m[624])|(m[342]&~m[620]&m[622]&m[623]&~m[624])|(~m[342]&m[620]&~m[622]&~m[623]&m[624])|(~m[342]&~m[620]&m[622]&~m[623]&m[624])|(m[342]&m[620]&m[622]&~m[623]&m[624])|(~m[342]&m[620]&m[622]&m[623]&m[624]))&UnbiasedRNG[242])|((m[342]&~m[620]&~m[622]&m[623]&~m[624])|(~m[342]&~m[620]&~m[622]&~m[623]&m[624])|(m[342]&~m[620]&~m[622]&~m[623]&m[624])|(m[342]&m[620]&~m[622]&~m[623]&m[624])|(m[342]&~m[620]&m[622]&~m[623]&m[624])|(~m[342]&~m[620]&~m[622]&m[623]&m[624])|(m[342]&~m[620]&~m[622]&m[623]&m[624])|(~m[342]&m[620]&~m[622]&m[623]&m[624])|(m[342]&m[620]&~m[622]&m[623]&m[624])|(~m[342]&~m[620]&m[622]&m[623]&m[624])|(m[342]&~m[620]&m[622]&m[623]&m[624])|(m[342]&m[620]&m[622]&m[623]&m[624]));
    m[627] = (((m[584]&~m[625]&~m[626]&~m[628]&~m[629])|(~m[584]&~m[625]&~m[626]&m[628]&~m[629])|(m[584]&m[625]&~m[626]&m[628]&~m[629])|(m[584]&~m[625]&m[626]&m[628]&~m[629])|(~m[584]&m[625]&~m[626]&~m[628]&m[629])|(~m[584]&~m[625]&m[626]&~m[628]&m[629])|(m[584]&m[625]&m[626]&~m[628]&m[629])|(~m[584]&m[625]&m[626]&m[628]&m[629]))&UnbiasedRNG[243])|((m[584]&~m[625]&~m[626]&m[628]&~m[629])|(~m[584]&~m[625]&~m[626]&~m[628]&m[629])|(m[584]&~m[625]&~m[626]&~m[628]&m[629])|(m[584]&m[625]&~m[626]&~m[628]&m[629])|(m[584]&~m[625]&m[626]&~m[628]&m[629])|(~m[584]&~m[625]&~m[626]&m[628]&m[629])|(m[584]&~m[625]&~m[626]&m[628]&m[629])|(~m[584]&m[625]&~m[626]&m[628]&m[629])|(m[584]&m[625]&~m[626]&m[628]&m[629])|(~m[584]&~m[625]&m[626]&m[628]&m[629])|(m[584]&~m[625]&m[626]&m[628]&m[629])|(m[584]&m[625]&m[626]&m[628]&m[629]));
    m[631] = (((m[289]&~m[630]&~m[632]&~m[633]&~m[634])|(~m[289]&~m[630]&~m[632]&m[633]&~m[634])|(m[289]&m[630]&~m[632]&m[633]&~m[634])|(m[289]&~m[630]&m[632]&m[633]&~m[634])|(~m[289]&m[630]&~m[632]&~m[633]&m[634])|(~m[289]&~m[630]&m[632]&~m[633]&m[634])|(m[289]&m[630]&m[632]&~m[633]&m[634])|(~m[289]&m[630]&m[632]&m[633]&m[634]))&UnbiasedRNG[244])|((m[289]&~m[630]&~m[632]&m[633]&~m[634])|(~m[289]&~m[630]&~m[632]&~m[633]&m[634])|(m[289]&~m[630]&~m[632]&~m[633]&m[634])|(m[289]&m[630]&~m[632]&~m[633]&m[634])|(m[289]&~m[630]&m[632]&~m[633]&m[634])|(~m[289]&~m[630]&~m[632]&m[633]&m[634])|(m[289]&~m[630]&~m[632]&m[633]&m[634])|(~m[289]&m[630]&~m[632]&m[633]&m[634])|(m[289]&m[630]&~m[632]&m[633]&m[634])|(~m[289]&~m[630]&m[632]&m[633]&m[634])|(m[289]&~m[630]&m[632]&m[633]&m[634])|(m[289]&m[630]&m[632]&m[633]&m[634]));
    m[636] = (((m[298]&~m[635]&~m[637]&~m[638]&~m[639])|(~m[298]&~m[635]&~m[637]&m[638]&~m[639])|(m[298]&m[635]&~m[637]&m[638]&~m[639])|(m[298]&~m[635]&m[637]&m[638]&~m[639])|(~m[298]&m[635]&~m[637]&~m[638]&m[639])|(~m[298]&~m[635]&m[637]&~m[638]&m[639])|(m[298]&m[635]&m[637]&~m[638]&m[639])|(~m[298]&m[635]&m[637]&m[638]&m[639]))&UnbiasedRNG[245])|((m[298]&~m[635]&~m[637]&m[638]&~m[639])|(~m[298]&~m[635]&~m[637]&~m[638]&m[639])|(m[298]&~m[635]&~m[637]&~m[638]&m[639])|(m[298]&m[635]&~m[637]&~m[638]&m[639])|(m[298]&~m[635]&m[637]&~m[638]&m[639])|(~m[298]&~m[635]&~m[637]&m[638]&m[639])|(m[298]&~m[635]&~m[637]&m[638]&m[639])|(~m[298]&m[635]&~m[637]&m[638]&m[639])|(m[298]&m[635]&~m[637]&m[638]&m[639])|(~m[298]&~m[635]&m[637]&m[638]&m[639])|(m[298]&~m[635]&m[637]&m[638]&m[639])|(m[298]&m[635]&m[637]&m[638]&m[639]));
    m[641] = (((m[307]&~m[640]&~m[642]&~m[643]&~m[644])|(~m[307]&~m[640]&~m[642]&m[643]&~m[644])|(m[307]&m[640]&~m[642]&m[643]&~m[644])|(m[307]&~m[640]&m[642]&m[643]&~m[644])|(~m[307]&m[640]&~m[642]&~m[643]&m[644])|(~m[307]&~m[640]&m[642]&~m[643]&m[644])|(m[307]&m[640]&m[642]&~m[643]&m[644])|(~m[307]&m[640]&m[642]&m[643]&m[644]))&UnbiasedRNG[246])|((m[307]&~m[640]&~m[642]&m[643]&~m[644])|(~m[307]&~m[640]&~m[642]&~m[643]&m[644])|(m[307]&~m[640]&~m[642]&~m[643]&m[644])|(m[307]&m[640]&~m[642]&~m[643]&m[644])|(m[307]&~m[640]&m[642]&~m[643]&m[644])|(~m[307]&~m[640]&~m[642]&m[643]&m[644])|(m[307]&~m[640]&~m[642]&m[643]&m[644])|(~m[307]&m[640]&~m[642]&m[643]&m[644])|(m[307]&m[640]&~m[642]&m[643]&m[644])|(~m[307]&~m[640]&m[642]&m[643]&m[644])|(m[307]&~m[640]&m[642]&m[643]&m[644])|(m[307]&m[640]&m[642]&m[643]&m[644]));
    m[646] = (((m[316]&~m[645]&~m[647]&~m[648]&~m[649])|(~m[316]&~m[645]&~m[647]&m[648]&~m[649])|(m[316]&m[645]&~m[647]&m[648]&~m[649])|(m[316]&~m[645]&m[647]&m[648]&~m[649])|(~m[316]&m[645]&~m[647]&~m[648]&m[649])|(~m[316]&~m[645]&m[647]&~m[648]&m[649])|(m[316]&m[645]&m[647]&~m[648]&m[649])|(~m[316]&m[645]&m[647]&m[648]&m[649]))&UnbiasedRNG[247])|((m[316]&~m[645]&~m[647]&m[648]&~m[649])|(~m[316]&~m[645]&~m[647]&~m[648]&m[649])|(m[316]&~m[645]&~m[647]&~m[648]&m[649])|(m[316]&m[645]&~m[647]&~m[648]&m[649])|(m[316]&~m[645]&m[647]&~m[648]&m[649])|(~m[316]&~m[645]&~m[647]&m[648]&m[649])|(m[316]&~m[645]&~m[647]&m[648]&m[649])|(~m[316]&m[645]&~m[647]&m[648]&m[649])|(m[316]&m[645]&~m[647]&m[648]&m[649])|(~m[316]&~m[645]&m[647]&m[648]&m[649])|(m[316]&~m[645]&m[647]&m[648]&m[649])|(m[316]&m[645]&m[647]&m[648]&m[649]));
    m[651] = (((m[325]&~m[650]&~m[652]&~m[653]&~m[654])|(~m[325]&~m[650]&~m[652]&m[653]&~m[654])|(m[325]&m[650]&~m[652]&m[653]&~m[654])|(m[325]&~m[650]&m[652]&m[653]&~m[654])|(~m[325]&m[650]&~m[652]&~m[653]&m[654])|(~m[325]&~m[650]&m[652]&~m[653]&m[654])|(m[325]&m[650]&m[652]&~m[653]&m[654])|(~m[325]&m[650]&m[652]&m[653]&m[654]))&UnbiasedRNG[248])|((m[325]&~m[650]&~m[652]&m[653]&~m[654])|(~m[325]&~m[650]&~m[652]&~m[653]&m[654])|(m[325]&~m[650]&~m[652]&~m[653]&m[654])|(m[325]&m[650]&~m[652]&~m[653]&m[654])|(m[325]&~m[650]&m[652]&~m[653]&m[654])|(~m[325]&~m[650]&~m[652]&m[653]&m[654])|(m[325]&~m[650]&~m[652]&m[653]&m[654])|(~m[325]&m[650]&~m[652]&m[653]&m[654])|(m[325]&m[650]&~m[652]&m[653]&m[654])|(~m[325]&~m[650]&m[652]&m[653]&m[654])|(m[325]&~m[650]&m[652]&m[653]&m[654])|(m[325]&m[650]&m[652]&m[653]&m[654]));
    m[656] = (((m[334]&~m[655]&~m[657]&~m[658]&~m[659])|(~m[334]&~m[655]&~m[657]&m[658]&~m[659])|(m[334]&m[655]&~m[657]&m[658]&~m[659])|(m[334]&~m[655]&m[657]&m[658]&~m[659])|(~m[334]&m[655]&~m[657]&~m[658]&m[659])|(~m[334]&~m[655]&m[657]&~m[658]&m[659])|(m[334]&m[655]&m[657]&~m[658]&m[659])|(~m[334]&m[655]&m[657]&m[658]&m[659]))&UnbiasedRNG[249])|((m[334]&~m[655]&~m[657]&m[658]&~m[659])|(~m[334]&~m[655]&~m[657]&~m[658]&m[659])|(m[334]&~m[655]&~m[657]&~m[658]&m[659])|(m[334]&m[655]&~m[657]&~m[658]&m[659])|(m[334]&~m[655]&m[657]&~m[658]&m[659])|(~m[334]&~m[655]&~m[657]&m[658]&m[659])|(m[334]&~m[655]&~m[657]&m[658]&m[659])|(~m[334]&m[655]&~m[657]&m[658]&m[659])|(m[334]&m[655]&~m[657]&m[658]&m[659])|(~m[334]&~m[655]&m[657]&m[658]&m[659])|(m[334]&~m[655]&m[657]&m[658]&m[659])|(m[334]&m[655]&m[657]&m[658]&m[659]));
    m[661] = (((m[343]&~m[660]&~m[662]&~m[663]&~m[664])|(~m[343]&~m[660]&~m[662]&m[663]&~m[664])|(m[343]&m[660]&~m[662]&m[663]&~m[664])|(m[343]&~m[660]&m[662]&m[663]&~m[664])|(~m[343]&m[660]&~m[662]&~m[663]&m[664])|(~m[343]&~m[660]&m[662]&~m[663]&m[664])|(m[343]&m[660]&m[662]&~m[663]&m[664])|(~m[343]&m[660]&m[662]&m[663]&m[664]))&UnbiasedRNG[250])|((m[343]&~m[660]&~m[662]&m[663]&~m[664])|(~m[343]&~m[660]&~m[662]&~m[663]&m[664])|(m[343]&~m[660]&~m[662]&~m[663]&m[664])|(m[343]&m[660]&~m[662]&~m[663]&m[664])|(m[343]&~m[660]&m[662]&~m[663]&m[664])|(~m[343]&~m[660]&~m[662]&m[663]&m[664])|(m[343]&~m[660]&~m[662]&m[663]&m[664])|(~m[343]&m[660]&~m[662]&m[663]&m[664])|(m[343]&m[660]&~m[662]&m[663]&m[664])|(~m[343]&~m[660]&m[662]&m[663]&m[664])|(m[343]&~m[660]&m[662]&m[663]&m[664])|(m[343]&m[660]&m[662]&m[663]&m[664]));
    m[666] = (((m[352]&~m[665]&~m[667]&~m[668]&~m[669])|(~m[352]&~m[665]&~m[667]&m[668]&~m[669])|(m[352]&m[665]&~m[667]&m[668]&~m[669])|(m[352]&~m[665]&m[667]&m[668]&~m[669])|(~m[352]&m[665]&~m[667]&~m[668]&m[669])|(~m[352]&~m[665]&m[667]&~m[668]&m[669])|(m[352]&m[665]&m[667]&~m[668]&m[669])|(~m[352]&m[665]&m[667]&m[668]&m[669]))&UnbiasedRNG[251])|((m[352]&~m[665]&~m[667]&m[668]&~m[669])|(~m[352]&~m[665]&~m[667]&~m[668]&m[669])|(m[352]&~m[665]&~m[667]&~m[668]&m[669])|(m[352]&m[665]&~m[667]&~m[668]&m[669])|(m[352]&~m[665]&m[667]&~m[668]&m[669])|(~m[352]&~m[665]&~m[667]&m[668]&m[669])|(m[352]&~m[665]&~m[667]&m[668]&m[669])|(~m[352]&m[665]&~m[667]&m[668]&m[669])|(m[352]&m[665]&~m[667]&m[668]&m[669])|(~m[352]&~m[665]&m[667]&m[668]&m[669])|(m[352]&~m[665]&m[667]&m[668]&m[669])|(m[352]&m[665]&m[667]&m[668]&m[669]));
    m[671] = (((m[299]&~m[670]&~m[672]&~m[673]&~m[674])|(~m[299]&~m[670]&~m[672]&m[673]&~m[674])|(m[299]&m[670]&~m[672]&m[673]&~m[674])|(m[299]&~m[670]&m[672]&m[673]&~m[674])|(~m[299]&m[670]&~m[672]&~m[673]&m[674])|(~m[299]&~m[670]&m[672]&~m[673]&m[674])|(m[299]&m[670]&m[672]&~m[673]&m[674])|(~m[299]&m[670]&m[672]&m[673]&m[674]))&UnbiasedRNG[252])|((m[299]&~m[670]&~m[672]&m[673]&~m[674])|(~m[299]&~m[670]&~m[672]&~m[673]&m[674])|(m[299]&~m[670]&~m[672]&~m[673]&m[674])|(m[299]&m[670]&~m[672]&~m[673]&m[674])|(m[299]&~m[670]&m[672]&~m[673]&m[674])|(~m[299]&~m[670]&~m[672]&m[673]&m[674])|(m[299]&~m[670]&~m[672]&m[673]&m[674])|(~m[299]&m[670]&~m[672]&m[673]&m[674])|(m[299]&m[670]&~m[672]&m[673]&m[674])|(~m[299]&~m[670]&m[672]&m[673]&m[674])|(m[299]&~m[670]&m[672]&m[673]&m[674])|(m[299]&m[670]&m[672]&m[673]&m[674]));
    m[676] = (((m[308]&~m[675]&~m[677]&~m[678]&~m[679])|(~m[308]&~m[675]&~m[677]&m[678]&~m[679])|(m[308]&m[675]&~m[677]&m[678]&~m[679])|(m[308]&~m[675]&m[677]&m[678]&~m[679])|(~m[308]&m[675]&~m[677]&~m[678]&m[679])|(~m[308]&~m[675]&m[677]&~m[678]&m[679])|(m[308]&m[675]&m[677]&~m[678]&m[679])|(~m[308]&m[675]&m[677]&m[678]&m[679]))&UnbiasedRNG[253])|((m[308]&~m[675]&~m[677]&m[678]&~m[679])|(~m[308]&~m[675]&~m[677]&~m[678]&m[679])|(m[308]&~m[675]&~m[677]&~m[678]&m[679])|(m[308]&m[675]&~m[677]&~m[678]&m[679])|(m[308]&~m[675]&m[677]&~m[678]&m[679])|(~m[308]&~m[675]&~m[677]&m[678]&m[679])|(m[308]&~m[675]&~m[677]&m[678]&m[679])|(~m[308]&m[675]&~m[677]&m[678]&m[679])|(m[308]&m[675]&~m[677]&m[678]&m[679])|(~m[308]&~m[675]&m[677]&m[678]&m[679])|(m[308]&~m[675]&m[677]&m[678]&m[679])|(m[308]&m[675]&m[677]&m[678]&m[679]));
    m[681] = (((m[317]&~m[680]&~m[682]&~m[683]&~m[684])|(~m[317]&~m[680]&~m[682]&m[683]&~m[684])|(m[317]&m[680]&~m[682]&m[683]&~m[684])|(m[317]&~m[680]&m[682]&m[683]&~m[684])|(~m[317]&m[680]&~m[682]&~m[683]&m[684])|(~m[317]&~m[680]&m[682]&~m[683]&m[684])|(m[317]&m[680]&m[682]&~m[683]&m[684])|(~m[317]&m[680]&m[682]&m[683]&m[684]))&UnbiasedRNG[254])|((m[317]&~m[680]&~m[682]&m[683]&~m[684])|(~m[317]&~m[680]&~m[682]&~m[683]&m[684])|(m[317]&~m[680]&~m[682]&~m[683]&m[684])|(m[317]&m[680]&~m[682]&~m[683]&m[684])|(m[317]&~m[680]&m[682]&~m[683]&m[684])|(~m[317]&~m[680]&~m[682]&m[683]&m[684])|(m[317]&~m[680]&~m[682]&m[683]&m[684])|(~m[317]&m[680]&~m[682]&m[683]&m[684])|(m[317]&m[680]&~m[682]&m[683]&m[684])|(~m[317]&~m[680]&m[682]&m[683]&m[684])|(m[317]&~m[680]&m[682]&m[683]&m[684])|(m[317]&m[680]&m[682]&m[683]&m[684]));
    m[686] = (((m[326]&~m[685]&~m[687]&~m[688]&~m[689])|(~m[326]&~m[685]&~m[687]&m[688]&~m[689])|(m[326]&m[685]&~m[687]&m[688]&~m[689])|(m[326]&~m[685]&m[687]&m[688]&~m[689])|(~m[326]&m[685]&~m[687]&~m[688]&m[689])|(~m[326]&~m[685]&m[687]&~m[688]&m[689])|(m[326]&m[685]&m[687]&~m[688]&m[689])|(~m[326]&m[685]&m[687]&m[688]&m[689]))&UnbiasedRNG[255])|((m[326]&~m[685]&~m[687]&m[688]&~m[689])|(~m[326]&~m[685]&~m[687]&~m[688]&m[689])|(m[326]&~m[685]&~m[687]&~m[688]&m[689])|(m[326]&m[685]&~m[687]&~m[688]&m[689])|(m[326]&~m[685]&m[687]&~m[688]&m[689])|(~m[326]&~m[685]&~m[687]&m[688]&m[689])|(m[326]&~m[685]&~m[687]&m[688]&m[689])|(~m[326]&m[685]&~m[687]&m[688]&m[689])|(m[326]&m[685]&~m[687]&m[688]&m[689])|(~m[326]&~m[685]&m[687]&m[688]&m[689])|(m[326]&~m[685]&m[687]&m[688]&m[689])|(m[326]&m[685]&m[687]&m[688]&m[689]));
    m[691] = (((m[335]&~m[690]&~m[692]&~m[693]&~m[694])|(~m[335]&~m[690]&~m[692]&m[693]&~m[694])|(m[335]&m[690]&~m[692]&m[693]&~m[694])|(m[335]&~m[690]&m[692]&m[693]&~m[694])|(~m[335]&m[690]&~m[692]&~m[693]&m[694])|(~m[335]&~m[690]&m[692]&~m[693]&m[694])|(m[335]&m[690]&m[692]&~m[693]&m[694])|(~m[335]&m[690]&m[692]&m[693]&m[694]))&UnbiasedRNG[256])|((m[335]&~m[690]&~m[692]&m[693]&~m[694])|(~m[335]&~m[690]&~m[692]&~m[693]&m[694])|(m[335]&~m[690]&~m[692]&~m[693]&m[694])|(m[335]&m[690]&~m[692]&~m[693]&m[694])|(m[335]&~m[690]&m[692]&~m[693]&m[694])|(~m[335]&~m[690]&~m[692]&m[693]&m[694])|(m[335]&~m[690]&~m[692]&m[693]&m[694])|(~m[335]&m[690]&~m[692]&m[693]&m[694])|(m[335]&m[690]&~m[692]&m[693]&m[694])|(~m[335]&~m[690]&m[692]&m[693]&m[694])|(m[335]&~m[690]&m[692]&m[693]&m[694])|(m[335]&m[690]&m[692]&m[693]&m[694]));
    m[696] = (((m[344]&~m[695]&~m[697]&~m[698]&~m[699])|(~m[344]&~m[695]&~m[697]&m[698]&~m[699])|(m[344]&m[695]&~m[697]&m[698]&~m[699])|(m[344]&~m[695]&m[697]&m[698]&~m[699])|(~m[344]&m[695]&~m[697]&~m[698]&m[699])|(~m[344]&~m[695]&m[697]&~m[698]&m[699])|(m[344]&m[695]&m[697]&~m[698]&m[699])|(~m[344]&m[695]&m[697]&m[698]&m[699]))&UnbiasedRNG[257])|((m[344]&~m[695]&~m[697]&m[698]&~m[699])|(~m[344]&~m[695]&~m[697]&~m[698]&m[699])|(m[344]&~m[695]&~m[697]&~m[698]&m[699])|(m[344]&m[695]&~m[697]&~m[698]&m[699])|(m[344]&~m[695]&m[697]&~m[698]&m[699])|(~m[344]&~m[695]&~m[697]&m[698]&m[699])|(m[344]&~m[695]&~m[697]&m[698]&m[699])|(~m[344]&m[695]&~m[697]&m[698]&m[699])|(m[344]&m[695]&~m[697]&m[698]&m[699])|(~m[344]&~m[695]&m[697]&m[698]&m[699])|(m[344]&~m[695]&m[697]&m[698]&m[699])|(m[344]&m[695]&m[697]&m[698]&m[699]));
    m[701] = (((m[353]&~m[700]&~m[702]&~m[703]&~m[704])|(~m[353]&~m[700]&~m[702]&m[703]&~m[704])|(m[353]&m[700]&~m[702]&m[703]&~m[704])|(m[353]&~m[700]&m[702]&m[703]&~m[704])|(~m[353]&m[700]&~m[702]&~m[703]&m[704])|(~m[353]&~m[700]&m[702]&~m[703]&m[704])|(m[353]&m[700]&m[702]&~m[703]&m[704])|(~m[353]&m[700]&m[702]&m[703]&m[704]))&UnbiasedRNG[258])|((m[353]&~m[700]&~m[702]&m[703]&~m[704])|(~m[353]&~m[700]&~m[702]&~m[703]&m[704])|(m[353]&~m[700]&~m[702]&~m[703]&m[704])|(m[353]&m[700]&~m[702]&~m[703]&m[704])|(m[353]&~m[700]&m[702]&~m[703]&m[704])|(~m[353]&~m[700]&~m[702]&m[703]&m[704])|(m[353]&~m[700]&~m[702]&m[703]&m[704])|(~m[353]&m[700]&~m[702]&m[703]&m[704])|(m[353]&m[700]&~m[702]&m[703]&m[704])|(~m[353]&~m[700]&m[702]&m[703]&m[704])|(m[353]&~m[700]&m[702]&m[703]&m[704])|(m[353]&m[700]&m[702]&m[703]&m[704]));
    m[706] = (((m[309]&~m[705]&~m[707]&~m[708]&~m[709])|(~m[309]&~m[705]&~m[707]&m[708]&~m[709])|(m[309]&m[705]&~m[707]&m[708]&~m[709])|(m[309]&~m[705]&m[707]&m[708]&~m[709])|(~m[309]&m[705]&~m[707]&~m[708]&m[709])|(~m[309]&~m[705]&m[707]&~m[708]&m[709])|(m[309]&m[705]&m[707]&~m[708]&m[709])|(~m[309]&m[705]&m[707]&m[708]&m[709]))&UnbiasedRNG[259])|((m[309]&~m[705]&~m[707]&m[708]&~m[709])|(~m[309]&~m[705]&~m[707]&~m[708]&m[709])|(m[309]&~m[705]&~m[707]&~m[708]&m[709])|(m[309]&m[705]&~m[707]&~m[708]&m[709])|(m[309]&~m[705]&m[707]&~m[708]&m[709])|(~m[309]&~m[705]&~m[707]&m[708]&m[709])|(m[309]&~m[705]&~m[707]&m[708]&m[709])|(~m[309]&m[705]&~m[707]&m[708]&m[709])|(m[309]&m[705]&~m[707]&m[708]&m[709])|(~m[309]&~m[705]&m[707]&m[708]&m[709])|(m[309]&~m[705]&m[707]&m[708]&m[709])|(m[309]&m[705]&m[707]&m[708]&m[709]));
    m[711] = (((m[318]&~m[710]&~m[712]&~m[713]&~m[714])|(~m[318]&~m[710]&~m[712]&m[713]&~m[714])|(m[318]&m[710]&~m[712]&m[713]&~m[714])|(m[318]&~m[710]&m[712]&m[713]&~m[714])|(~m[318]&m[710]&~m[712]&~m[713]&m[714])|(~m[318]&~m[710]&m[712]&~m[713]&m[714])|(m[318]&m[710]&m[712]&~m[713]&m[714])|(~m[318]&m[710]&m[712]&m[713]&m[714]))&UnbiasedRNG[260])|((m[318]&~m[710]&~m[712]&m[713]&~m[714])|(~m[318]&~m[710]&~m[712]&~m[713]&m[714])|(m[318]&~m[710]&~m[712]&~m[713]&m[714])|(m[318]&m[710]&~m[712]&~m[713]&m[714])|(m[318]&~m[710]&m[712]&~m[713]&m[714])|(~m[318]&~m[710]&~m[712]&m[713]&m[714])|(m[318]&~m[710]&~m[712]&m[713]&m[714])|(~m[318]&m[710]&~m[712]&m[713]&m[714])|(m[318]&m[710]&~m[712]&m[713]&m[714])|(~m[318]&~m[710]&m[712]&m[713]&m[714])|(m[318]&~m[710]&m[712]&m[713]&m[714])|(m[318]&m[710]&m[712]&m[713]&m[714]));
    m[716] = (((m[327]&~m[715]&~m[717]&~m[718]&~m[719])|(~m[327]&~m[715]&~m[717]&m[718]&~m[719])|(m[327]&m[715]&~m[717]&m[718]&~m[719])|(m[327]&~m[715]&m[717]&m[718]&~m[719])|(~m[327]&m[715]&~m[717]&~m[718]&m[719])|(~m[327]&~m[715]&m[717]&~m[718]&m[719])|(m[327]&m[715]&m[717]&~m[718]&m[719])|(~m[327]&m[715]&m[717]&m[718]&m[719]))&UnbiasedRNG[261])|((m[327]&~m[715]&~m[717]&m[718]&~m[719])|(~m[327]&~m[715]&~m[717]&~m[718]&m[719])|(m[327]&~m[715]&~m[717]&~m[718]&m[719])|(m[327]&m[715]&~m[717]&~m[718]&m[719])|(m[327]&~m[715]&m[717]&~m[718]&m[719])|(~m[327]&~m[715]&~m[717]&m[718]&m[719])|(m[327]&~m[715]&~m[717]&m[718]&m[719])|(~m[327]&m[715]&~m[717]&m[718]&m[719])|(m[327]&m[715]&~m[717]&m[718]&m[719])|(~m[327]&~m[715]&m[717]&m[718]&m[719])|(m[327]&~m[715]&m[717]&m[718]&m[719])|(m[327]&m[715]&m[717]&m[718]&m[719]));
    m[721] = (((m[336]&~m[720]&~m[722]&~m[723]&~m[724])|(~m[336]&~m[720]&~m[722]&m[723]&~m[724])|(m[336]&m[720]&~m[722]&m[723]&~m[724])|(m[336]&~m[720]&m[722]&m[723]&~m[724])|(~m[336]&m[720]&~m[722]&~m[723]&m[724])|(~m[336]&~m[720]&m[722]&~m[723]&m[724])|(m[336]&m[720]&m[722]&~m[723]&m[724])|(~m[336]&m[720]&m[722]&m[723]&m[724]))&UnbiasedRNG[262])|((m[336]&~m[720]&~m[722]&m[723]&~m[724])|(~m[336]&~m[720]&~m[722]&~m[723]&m[724])|(m[336]&~m[720]&~m[722]&~m[723]&m[724])|(m[336]&m[720]&~m[722]&~m[723]&m[724])|(m[336]&~m[720]&m[722]&~m[723]&m[724])|(~m[336]&~m[720]&~m[722]&m[723]&m[724])|(m[336]&~m[720]&~m[722]&m[723]&m[724])|(~m[336]&m[720]&~m[722]&m[723]&m[724])|(m[336]&m[720]&~m[722]&m[723]&m[724])|(~m[336]&~m[720]&m[722]&m[723]&m[724])|(m[336]&~m[720]&m[722]&m[723]&m[724])|(m[336]&m[720]&m[722]&m[723]&m[724]));
    m[726] = (((m[345]&~m[725]&~m[727]&~m[728]&~m[729])|(~m[345]&~m[725]&~m[727]&m[728]&~m[729])|(m[345]&m[725]&~m[727]&m[728]&~m[729])|(m[345]&~m[725]&m[727]&m[728]&~m[729])|(~m[345]&m[725]&~m[727]&~m[728]&m[729])|(~m[345]&~m[725]&m[727]&~m[728]&m[729])|(m[345]&m[725]&m[727]&~m[728]&m[729])|(~m[345]&m[725]&m[727]&m[728]&m[729]))&UnbiasedRNG[263])|((m[345]&~m[725]&~m[727]&m[728]&~m[729])|(~m[345]&~m[725]&~m[727]&~m[728]&m[729])|(m[345]&~m[725]&~m[727]&~m[728]&m[729])|(m[345]&m[725]&~m[727]&~m[728]&m[729])|(m[345]&~m[725]&m[727]&~m[728]&m[729])|(~m[345]&~m[725]&~m[727]&m[728]&m[729])|(m[345]&~m[725]&~m[727]&m[728]&m[729])|(~m[345]&m[725]&~m[727]&m[728]&m[729])|(m[345]&m[725]&~m[727]&m[728]&m[729])|(~m[345]&~m[725]&m[727]&m[728]&m[729])|(m[345]&~m[725]&m[727]&m[728]&m[729])|(m[345]&m[725]&m[727]&m[728]&m[729]));
    m[731] = (((m[354]&~m[730]&~m[732]&~m[733]&~m[734])|(~m[354]&~m[730]&~m[732]&m[733]&~m[734])|(m[354]&m[730]&~m[732]&m[733]&~m[734])|(m[354]&~m[730]&m[732]&m[733]&~m[734])|(~m[354]&m[730]&~m[732]&~m[733]&m[734])|(~m[354]&~m[730]&m[732]&~m[733]&m[734])|(m[354]&m[730]&m[732]&~m[733]&m[734])|(~m[354]&m[730]&m[732]&m[733]&m[734]))&UnbiasedRNG[264])|((m[354]&~m[730]&~m[732]&m[733]&~m[734])|(~m[354]&~m[730]&~m[732]&~m[733]&m[734])|(m[354]&~m[730]&~m[732]&~m[733]&m[734])|(m[354]&m[730]&~m[732]&~m[733]&m[734])|(m[354]&~m[730]&m[732]&~m[733]&m[734])|(~m[354]&~m[730]&~m[732]&m[733]&m[734])|(m[354]&~m[730]&~m[732]&m[733]&m[734])|(~m[354]&m[730]&~m[732]&m[733]&m[734])|(m[354]&m[730]&~m[732]&m[733]&m[734])|(~m[354]&~m[730]&m[732]&m[733]&m[734])|(m[354]&~m[730]&m[732]&m[733]&m[734])|(m[354]&m[730]&m[732]&m[733]&m[734]));
    m[736] = (((m[319]&~m[735]&~m[737]&~m[738]&~m[739])|(~m[319]&~m[735]&~m[737]&m[738]&~m[739])|(m[319]&m[735]&~m[737]&m[738]&~m[739])|(m[319]&~m[735]&m[737]&m[738]&~m[739])|(~m[319]&m[735]&~m[737]&~m[738]&m[739])|(~m[319]&~m[735]&m[737]&~m[738]&m[739])|(m[319]&m[735]&m[737]&~m[738]&m[739])|(~m[319]&m[735]&m[737]&m[738]&m[739]))&UnbiasedRNG[265])|((m[319]&~m[735]&~m[737]&m[738]&~m[739])|(~m[319]&~m[735]&~m[737]&~m[738]&m[739])|(m[319]&~m[735]&~m[737]&~m[738]&m[739])|(m[319]&m[735]&~m[737]&~m[738]&m[739])|(m[319]&~m[735]&m[737]&~m[738]&m[739])|(~m[319]&~m[735]&~m[737]&m[738]&m[739])|(m[319]&~m[735]&~m[737]&m[738]&m[739])|(~m[319]&m[735]&~m[737]&m[738]&m[739])|(m[319]&m[735]&~m[737]&m[738]&m[739])|(~m[319]&~m[735]&m[737]&m[738]&m[739])|(m[319]&~m[735]&m[737]&m[738]&m[739])|(m[319]&m[735]&m[737]&m[738]&m[739]));
    m[741] = (((m[328]&~m[740]&~m[742]&~m[743]&~m[744])|(~m[328]&~m[740]&~m[742]&m[743]&~m[744])|(m[328]&m[740]&~m[742]&m[743]&~m[744])|(m[328]&~m[740]&m[742]&m[743]&~m[744])|(~m[328]&m[740]&~m[742]&~m[743]&m[744])|(~m[328]&~m[740]&m[742]&~m[743]&m[744])|(m[328]&m[740]&m[742]&~m[743]&m[744])|(~m[328]&m[740]&m[742]&m[743]&m[744]))&UnbiasedRNG[266])|((m[328]&~m[740]&~m[742]&m[743]&~m[744])|(~m[328]&~m[740]&~m[742]&~m[743]&m[744])|(m[328]&~m[740]&~m[742]&~m[743]&m[744])|(m[328]&m[740]&~m[742]&~m[743]&m[744])|(m[328]&~m[740]&m[742]&~m[743]&m[744])|(~m[328]&~m[740]&~m[742]&m[743]&m[744])|(m[328]&~m[740]&~m[742]&m[743]&m[744])|(~m[328]&m[740]&~m[742]&m[743]&m[744])|(m[328]&m[740]&~m[742]&m[743]&m[744])|(~m[328]&~m[740]&m[742]&m[743]&m[744])|(m[328]&~m[740]&m[742]&m[743]&m[744])|(m[328]&m[740]&m[742]&m[743]&m[744]));
    m[746] = (((m[337]&~m[745]&~m[747]&~m[748]&~m[749])|(~m[337]&~m[745]&~m[747]&m[748]&~m[749])|(m[337]&m[745]&~m[747]&m[748]&~m[749])|(m[337]&~m[745]&m[747]&m[748]&~m[749])|(~m[337]&m[745]&~m[747]&~m[748]&m[749])|(~m[337]&~m[745]&m[747]&~m[748]&m[749])|(m[337]&m[745]&m[747]&~m[748]&m[749])|(~m[337]&m[745]&m[747]&m[748]&m[749]))&UnbiasedRNG[267])|((m[337]&~m[745]&~m[747]&m[748]&~m[749])|(~m[337]&~m[745]&~m[747]&~m[748]&m[749])|(m[337]&~m[745]&~m[747]&~m[748]&m[749])|(m[337]&m[745]&~m[747]&~m[748]&m[749])|(m[337]&~m[745]&m[747]&~m[748]&m[749])|(~m[337]&~m[745]&~m[747]&m[748]&m[749])|(m[337]&~m[745]&~m[747]&m[748]&m[749])|(~m[337]&m[745]&~m[747]&m[748]&m[749])|(m[337]&m[745]&~m[747]&m[748]&m[749])|(~m[337]&~m[745]&m[747]&m[748]&m[749])|(m[337]&~m[745]&m[747]&m[748]&m[749])|(m[337]&m[745]&m[747]&m[748]&m[749]));
    m[751] = (((m[346]&~m[750]&~m[752]&~m[753]&~m[754])|(~m[346]&~m[750]&~m[752]&m[753]&~m[754])|(m[346]&m[750]&~m[752]&m[753]&~m[754])|(m[346]&~m[750]&m[752]&m[753]&~m[754])|(~m[346]&m[750]&~m[752]&~m[753]&m[754])|(~m[346]&~m[750]&m[752]&~m[753]&m[754])|(m[346]&m[750]&m[752]&~m[753]&m[754])|(~m[346]&m[750]&m[752]&m[753]&m[754]))&UnbiasedRNG[268])|((m[346]&~m[750]&~m[752]&m[753]&~m[754])|(~m[346]&~m[750]&~m[752]&~m[753]&m[754])|(m[346]&~m[750]&~m[752]&~m[753]&m[754])|(m[346]&m[750]&~m[752]&~m[753]&m[754])|(m[346]&~m[750]&m[752]&~m[753]&m[754])|(~m[346]&~m[750]&~m[752]&m[753]&m[754])|(m[346]&~m[750]&~m[752]&m[753]&m[754])|(~m[346]&m[750]&~m[752]&m[753]&m[754])|(m[346]&m[750]&~m[752]&m[753]&m[754])|(~m[346]&~m[750]&m[752]&m[753]&m[754])|(m[346]&~m[750]&m[752]&m[753]&m[754])|(m[346]&m[750]&m[752]&m[753]&m[754]));
    m[756] = (((m[355]&~m[755]&~m[757]&~m[758]&~m[759])|(~m[355]&~m[755]&~m[757]&m[758]&~m[759])|(m[355]&m[755]&~m[757]&m[758]&~m[759])|(m[355]&~m[755]&m[757]&m[758]&~m[759])|(~m[355]&m[755]&~m[757]&~m[758]&m[759])|(~m[355]&~m[755]&m[757]&~m[758]&m[759])|(m[355]&m[755]&m[757]&~m[758]&m[759])|(~m[355]&m[755]&m[757]&m[758]&m[759]))&UnbiasedRNG[269])|((m[355]&~m[755]&~m[757]&m[758]&~m[759])|(~m[355]&~m[755]&~m[757]&~m[758]&m[759])|(m[355]&~m[755]&~m[757]&~m[758]&m[759])|(m[355]&m[755]&~m[757]&~m[758]&m[759])|(m[355]&~m[755]&m[757]&~m[758]&m[759])|(~m[355]&~m[755]&~m[757]&m[758]&m[759])|(m[355]&~m[755]&~m[757]&m[758]&m[759])|(~m[355]&m[755]&~m[757]&m[758]&m[759])|(m[355]&m[755]&~m[757]&m[758]&m[759])|(~m[355]&~m[755]&m[757]&m[758]&m[759])|(m[355]&~m[755]&m[757]&m[758]&m[759])|(m[355]&m[755]&m[757]&m[758]&m[759]));
    m[761] = (((m[329]&~m[760]&~m[762]&~m[763]&~m[764])|(~m[329]&~m[760]&~m[762]&m[763]&~m[764])|(m[329]&m[760]&~m[762]&m[763]&~m[764])|(m[329]&~m[760]&m[762]&m[763]&~m[764])|(~m[329]&m[760]&~m[762]&~m[763]&m[764])|(~m[329]&~m[760]&m[762]&~m[763]&m[764])|(m[329]&m[760]&m[762]&~m[763]&m[764])|(~m[329]&m[760]&m[762]&m[763]&m[764]))&UnbiasedRNG[270])|((m[329]&~m[760]&~m[762]&m[763]&~m[764])|(~m[329]&~m[760]&~m[762]&~m[763]&m[764])|(m[329]&~m[760]&~m[762]&~m[763]&m[764])|(m[329]&m[760]&~m[762]&~m[763]&m[764])|(m[329]&~m[760]&m[762]&~m[763]&m[764])|(~m[329]&~m[760]&~m[762]&m[763]&m[764])|(m[329]&~m[760]&~m[762]&m[763]&m[764])|(~m[329]&m[760]&~m[762]&m[763]&m[764])|(m[329]&m[760]&~m[762]&m[763]&m[764])|(~m[329]&~m[760]&m[762]&m[763]&m[764])|(m[329]&~m[760]&m[762]&m[763]&m[764])|(m[329]&m[760]&m[762]&m[763]&m[764]));
    m[766] = (((m[338]&~m[765]&~m[767]&~m[768]&~m[769])|(~m[338]&~m[765]&~m[767]&m[768]&~m[769])|(m[338]&m[765]&~m[767]&m[768]&~m[769])|(m[338]&~m[765]&m[767]&m[768]&~m[769])|(~m[338]&m[765]&~m[767]&~m[768]&m[769])|(~m[338]&~m[765]&m[767]&~m[768]&m[769])|(m[338]&m[765]&m[767]&~m[768]&m[769])|(~m[338]&m[765]&m[767]&m[768]&m[769]))&UnbiasedRNG[271])|((m[338]&~m[765]&~m[767]&m[768]&~m[769])|(~m[338]&~m[765]&~m[767]&~m[768]&m[769])|(m[338]&~m[765]&~m[767]&~m[768]&m[769])|(m[338]&m[765]&~m[767]&~m[768]&m[769])|(m[338]&~m[765]&m[767]&~m[768]&m[769])|(~m[338]&~m[765]&~m[767]&m[768]&m[769])|(m[338]&~m[765]&~m[767]&m[768]&m[769])|(~m[338]&m[765]&~m[767]&m[768]&m[769])|(m[338]&m[765]&~m[767]&m[768]&m[769])|(~m[338]&~m[765]&m[767]&m[768]&m[769])|(m[338]&~m[765]&m[767]&m[768]&m[769])|(m[338]&m[765]&m[767]&m[768]&m[769]));
    m[771] = (((m[347]&~m[770]&~m[772]&~m[773]&~m[774])|(~m[347]&~m[770]&~m[772]&m[773]&~m[774])|(m[347]&m[770]&~m[772]&m[773]&~m[774])|(m[347]&~m[770]&m[772]&m[773]&~m[774])|(~m[347]&m[770]&~m[772]&~m[773]&m[774])|(~m[347]&~m[770]&m[772]&~m[773]&m[774])|(m[347]&m[770]&m[772]&~m[773]&m[774])|(~m[347]&m[770]&m[772]&m[773]&m[774]))&UnbiasedRNG[272])|((m[347]&~m[770]&~m[772]&m[773]&~m[774])|(~m[347]&~m[770]&~m[772]&~m[773]&m[774])|(m[347]&~m[770]&~m[772]&~m[773]&m[774])|(m[347]&m[770]&~m[772]&~m[773]&m[774])|(m[347]&~m[770]&m[772]&~m[773]&m[774])|(~m[347]&~m[770]&~m[772]&m[773]&m[774])|(m[347]&~m[770]&~m[772]&m[773]&m[774])|(~m[347]&m[770]&~m[772]&m[773]&m[774])|(m[347]&m[770]&~m[772]&m[773]&m[774])|(~m[347]&~m[770]&m[772]&m[773]&m[774])|(m[347]&~m[770]&m[772]&m[773]&m[774])|(m[347]&m[770]&m[772]&m[773]&m[774]));
    m[776] = (((m[356]&~m[775]&~m[777]&~m[778]&~m[779])|(~m[356]&~m[775]&~m[777]&m[778]&~m[779])|(m[356]&m[775]&~m[777]&m[778]&~m[779])|(m[356]&~m[775]&m[777]&m[778]&~m[779])|(~m[356]&m[775]&~m[777]&~m[778]&m[779])|(~m[356]&~m[775]&m[777]&~m[778]&m[779])|(m[356]&m[775]&m[777]&~m[778]&m[779])|(~m[356]&m[775]&m[777]&m[778]&m[779]))&UnbiasedRNG[273])|((m[356]&~m[775]&~m[777]&m[778]&~m[779])|(~m[356]&~m[775]&~m[777]&~m[778]&m[779])|(m[356]&~m[775]&~m[777]&~m[778]&m[779])|(m[356]&m[775]&~m[777]&~m[778]&m[779])|(m[356]&~m[775]&m[777]&~m[778]&m[779])|(~m[356]&~m[775]&~m[777]&m[778]&m[779])|(m[356]&~m[775]&~m[777]&m[778]&m[779])|(~m[356]&m[775]&~m[777]&m[778]&m[779])|(m[356]&m[775]&~m[777]&m[778]&m[779])|(~m[356]&~m[775]&m[777]&m[778]&m[779])|(m[356]&~m[775]&m[777]&m[778]&m[779])|(m[356]&m[775]&m[777]&m[778]&m[779]));
    m[781] = (((m[339]&~m[780]&~m[782]&~m[783]&~m[784])|(~m[339]&~m[780]&~m[782]&m[783]&~m[784])|(m[339]&m[780]&~m[782]&m[783]&~m[784])|(m[339]&~m[780]&m[782]&m[783]&~m[784])|(~m[339]&m[780]&~m[782]&~m[783]&m[784])|(~m[339]&~m[780]&m[782]&~m[783]&m[784])|(m[339]&m[780]&m[782]&~m[783]&m[784])|(~m[339]&m[780]&m[782]&m[783]&m[784]))&UnbiasedRNG[274])|((m[339]&~m[780]&~m[782]&m[783]&~m[784])|(~m[339]&~m[780]&~m[782]&~m[783]&m[784])|(m[339]&~m[780]&~m[782]&~m[783]&m[784])|(m[339]&m[780]&~m[782]&~m[783]&m[784])|(m[339]&~m[780]&m[782]&~m[783]&m[784])|(~m[339]&~m[780]&~m[782]&m[783]&m[784])|(m[339]&~m[780]&~m[782]&m[783]&m[784])|(~m[339]&m[780]&~m[782]&m[783]&m[784])|(m[339]&m[780]&~m[782]&m[783]&m[784])|(~m[339]&~m[780]&m[782]&m[783]&m[784])|(m[339]&~m[780]&m[782]&m[783]&m[784])|(m[339]&m[780]&m[782]&m[783]&m[784]));
    m[786] = (((m[348]&~m[785]&~m[787]&~m[788]&~m[789])|(~m[348]&~m[785]&~m[787]&m[788]&~m[789])|(m[348]&m[785]&~m[787]&m[788]&~m[789])|(m[348]&~m[785]&m[787]&m[788]&~m[789])|(~m[348]&m[785]&~m[787]&~m[788]&m[789])|(~m[348]&~m[785]&m[787]&~m[788]&m[789])|(m[348]&m[785]&m[787]&~m[788]&m[789])|(~m[348]&m[785]&m[787]&m[788]&m[789]))&UnbiasedRNG[275])|((m[348]&~m[785]&~m[787]&m[788]&~m[789])|(~m[348]&~m[785]&~m[787]&~m[788]&m[789])|(m[348]&~m[785]&~m[787]&~m[788]&m[789])|(m[348]&m[785]&~m[787]&~m[788]&m[789])|(m[348]&~m[785]&m[787]&~m[788]&m[789])|(~m[348]&~m[785]&~m[787]&m[788]&m[789])|(m[348]&~m[785]&~m[787]&m[788]&m[789])|(~m[348]&m[785]&~m[787]&m[788]&m[789])|(m[348]&m[785]&~m[787]&m[788]&m[789])|(~m[348]&~m[785]&m[787]&m[788]&m[789])|(m[348]&~m[785]&m[787]&m[788]&m[789])|(m[348]&m[785]&m[787]&m[788]&m[789]));
    m[791] = (((m[357]&~m[790]&~m[792]&~m[793]&~m[794])|(~m[357]&~m[790]&~m[792]&m[793]&~m[794])|(m[357]&m[790]&~m[792]&m[793]&~m[794])|(m[357]&~m[790]&m[792]&m[793]&~m[794])|(~m[357]&m[790]&~m[792]&~m[793]&m[794])|(~m[357]&~m[790]&m[792]&~m[793]&m[794])|(m[357]&m[790]&m[792]&~m[793]&m[794])|(~m[357]&m[790]&m[792]&m[793]&m[794]))&UnbiasedRNG[276])|((m[357]&~m[790]&~m[792]&m[793]&~m[794])|(~m[357]&~m[790]&~m[792]&~m[793]&m[794])|(m[357]&~m[790]&~m[792]&~m[793]&m[794])|(m[357]&m[790]&~m[792]&~m[793]&m[794])|(m[357]&~m[790]&m[792]&~m[793]&m[794])|(~m[357]&~m[790]&~m[792]&m[793]&m[794])|(m[357]&~m[790]&~m[792]&m[793]&m[794])|(~m[357]&m[790]&~m[792]&m[793]&m[794])|(m[357]&m[790]&~m[792]&m[793]&m[794])|(~m[357]&~m[790]&m[792]&m[793]&m[794])|(m[357]&~m[790]&m[792]&m[793]&m[794])|(m[357]&m[790]&m[792]&m[793]&m[794]));
    m[796] = (((m[349]&~m[795]&~m[797]&~m[798]&~m[799])|(~m[349]&~m[795]&~m[797]&m[798]&~m[799])|(m[349]&m[795]&~m[797]&m[798]&~m[799])|(m[349]&~m[795]&m[797]&m[798]&~m[799])|(~m[349]&m[795]&~m[797]&~m[798]&m[799])|(~m[349]&~m[795]&m[797]&~m[798]&m[799])|(m[349]&m[795]&m[797]&~m[798]&m[799])|(~m[349]&m[795]&m[797]&m[798]&m[799]))&UnbiasedRNG[277])|((m[349]&~m[795]&~m[797]&m[798]&~m[799])|(~m[349]&~m[795]&~m[797]&~m[798]&m[799])|(m[349]&~m[795]&~m[797]&~m[798]&m[799])|(m[349]&m[795]&~m[797]&~m[798]&m[799])|(m[349]&~m[795]&m[797]&~m[798]&m[799])|(~m[349]&~m[795]&~m[797]&m[798]&m[799])|(m[349]&~m[795]&~m[797]&m[798]&m[799])|(~m[349]&m[795]&~m[797]&m[798]&m[799])|(m[349]&m[795]&~m[797]&m[798]&m[799])|(~m[349]&~m[795]&m[797]&m[798]&m[799])|(m[349]&~m[795]&m[797]&m[798]&m[799])|(m[349]&m[795]&m[797]&m[798]&m[799]));
    m[801] = (((m[358]&~m[800]&~m[802]&~m[803]&~m[804])|(~m[358]&~m[800]&~m[802]&m[803]&~m[804])|(m[358]&m[800]&~m[802]&m[803]&~m[804])|(m[358]&~m[800]&m[802]&m[803]&~m[804])|(~m[358]&m[800]&~m[802]&~m[803]&m[804])|(~m[358]&~m[800]&m[802]&~m[803]&m[804])|(m[358]&m[800]&m[802]&~m[803]&m[804])|(~m[358]&m[800]&m[802]&m[803]&m[804]))&UnbiasedRNG[278])|((m[358]&~m[800]&~m[802]&m[803]&~m[804])|(~m[358]&~m[800]&~m[802]&~m[803]&m[804])|(m[358]&~m[800]&~m[802]&~m[803]&m[804])|(m[358]&m[800]&~m[802]&~m[803]&m[804])|(m[358]&~m[800]&m[802]&~m[803]&m[804])|(~m[358]&~m[800]&~m[802]&m[803]&m[804])|(m[358]&~m[800]&~m[802]&m[803]&m[804])|(~m[358]&m[800]&~m[802]&m[803]&m[804])|(m[358]&m[800]&~m[802]&m[803]&m[804])|(~m[358]&~m[800]&m[802]&m[803]&m[804])|(m[358]&~m[800]&m[802]&m[803]&m[804])|(m[358]&m[800]&m[802]&m[803]&m[804]));
    m[806] = (((m[359]&~m[805]&~m[807]&~m[808]&~m[809])|(~m[359]&~m[805]&~m[807]&m[808]&~m[809])|(m[359]&m[805]&~m[807]&m[808]&~m[809])|(m[359]&~m[805]&m[807]&m[808]&~m[809])|(~m[359]&m[805]&~m[807]&~m[808]&m[809])|(~m[359]&~m[805]&m[807]&~m[808]&m[809])|(m[359]&m[805]&m[807]&~m[808]&m[809])|(~m[359]&m[805]&m[807]&m[808]&m[809]))&UnbiasedRNG[279])|((m[359]&~m[805]&~m[807]&m[808]&~m[809])|(~m[359]&~m[805]&~m[807]&~m[808]&m[809])|(m[359]&~m[805]&~m[807]&~m[808]&m[809])|(m[359]&m[805]&~m[807]&~m[808]&m[809])|(m[359]&~m[805]&m[807]&~m[808]&m[809])|(~m[359]&~m[805]&~m[807]&m[808]&m[809])|(m[359]&~m[805]&~m[807]&m[808]&m[809])|(~m[359]&m[805]&~m[807]&m[808]&m[809])|(m[359]&m[805]&~m[807]&m[808]&m[809])|(~m[359]&~m[805]&m[807]&m[808]&m[809])|(m[359]&~m[805]&m[807]&m[808]&m[809])|(m[359]&m[805]&m[807]&m[808]&m[809]));
end

always @(posedge color3_clk) begin
    m[368] = (((m[365]&~m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&~m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&m[369]&~m[370])|(~m[365]&~m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&m[369]&m[370])|(m[365]&~m[366]&m[367]&m[369]&m[370])|(~m[365]&m[366]&m[367]&m[369]&m[370]))&UnbiasedRNG[280])|((m[365]&m[366]&~m[367]&~m[369]&~m[370])|(m[365]&~m[366]&m[367]&~m[369]&~m[370])|(~m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&~m[366]&~m[367]&~m[369]&m[370])|(~m[365]&m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&~m[369]&m[370])|(~m[365]&~m[366]&m[367]&~m[369]&m[370])|(m[365]&~m[366]&m[367]&~m[369]&m[370])|(~m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&m[369]&m[370]));
    m[378] = (((m[375]&~m[376]&~m[377]&~m[379]&~m[380])|(~m[375]&m[376]&~m[377]&~m[379]&~m[380])|(~m[375]&~m[376]&m[377]&~m[379]&~m[380])|(m[375]&m[376]&m[377]&m[379]&~m[380])|(~m[375]&~m[376]&~m[377]&~m[379]&m[380])|(m[375]&m[376]&~m[377]&m[379]&m[380])|(m[375]&~m[376]&m[377]&m[379]&m[380])|(~m[375]&m[376]&m[377]&m[379]&m[380]))&UnbiasedRNG[281])|((m[375]&m[376]&~m[377]&~m[379]&~m[380])|(m[375]&~m[376]&m[377]&~m[379]&~m[380])|(~m[375]&m[376]&m[377]&~m[379]&~m[380])|(m[375]&m[376]&m[377]&~m[379]&~m[380])|(m[375]&~m[376]&~m[377]&~m[379]&m[380])|(~m[375]&m[376]&~m[377]&~m[379]&m[380])|(m[375]&m[376]&~m[377]&~m[379]&m[380])|(~m[375]&~m[376]&m[377]&~m[379]&m[380])|(m[375]&~m[376]&m[377]&~m[379]&m[380])|(~m[375]&m[376]&m[377]&~m[379]&m[380])|(m[375]&m[376]&m[377]&~m[379]&m[380])|(m[375]&m[376]&m[377]&m[379]&m[380]));
    m[383] = (((m[380]&~m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&~m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&m[384]&~m[385])|(~m[380]&~m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&m[384]&m[385])|(m[380]&~m[381]&m[382]&m[384]&m[385])|(~m[380]&m[381]&m[382]&m[384]&m[385]))&UnbiasedRNG[282])|((m[380]&m[381]&~m[382]&~m[384]&~m[385])|(m[380]&~m[381]&m[382]&~m[384]&~m[385])|(~m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&~m[381]&~m[382]&~m[384]&m[385])|(~m[380]&m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&~m[384]&m[385])|(~m[380]&~m[381]&m[382]&~m[384]&m[385])|(m[380]&~m[381]&m[382]&~m[384]&m[385])|(~m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&m[384]&m[385]));
    m[393] = (((m[390]&~m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&~m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&m[394]&~m[395])|(~m[390]&~m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&m[394]&m[395])|(m[390]&~m[391]&m[392]&m[394]&m[395])|(~m[390]&m[391]&m[392]&m[394]&m[395]))&UnbiasedRNG[283])|((m[390]&m[391]&~m[392]&~m[394]&~m[395])|(m[390]&~m[391]&m[392]&~m[394]&~m[395])|(~m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&~m[391]&~m[392]&~m[394]&m[395])|(~m[390]&m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&~m[394]&m[395])|(~m[390]&~m[391]&m[392]&~m[394]&m[395])|(m[390]&~m[391]&m[392]&~m[394]&m[395])|(~m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&m[394]&m[395]));
    m[398] = (((m[395]&~m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&~m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&m[399]&~m[400])|(~m[395]&~m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&m[399]&m[400])|(m[395]&~m[396]&m[397]&m[399]&m[400])|(~m[395]&m[396]&m[397]&m[399]&m[400]))&UnbiasedRNG[284])|((m[395]&m[396]&~m[397]&~m[399]&~m[400])|(m[395]&~m[396]&m[397]&~m[399]&~m[400])|(~m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&~m[396]&~m[397]&~m[399]&m[400])|(~m[395]&m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&~m[399]&m[400])|(~m[395]&~m[396]&m[397]&~m[399]&m[400])|(m[395]&~m[396]&m[397]&~m[399]&m[400])|(~m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&m[399]&m[400]));
    m[403] = (((m[400]&~m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&~m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&m[404]&~m[405])|(~m[400]&~m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&m[404]&m[405])|(m[400]&~m[401]&m[402]&m[404]&m[405])|(~m[400]&m[401]&m[402]&m[404]&m[405]))&UnbiasedRNG[285])|((m[400]&m[401]&~m[402]&~m[404]&~m[405])|(m[400]&~m[401]&m[402]&~m[404]&~m[405])|(~m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&~m[401]&~m[402]&~m[404]&m[405])|(~m[400]&m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&~m[404]&m[405])|(~m[400]&~m[401]&m[402]&~m[404]&m[405])|(m[400]&~m[401]&m[402]&~m[404]&m[405])|(~m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&m[404]&m[405]));
    m[413] = (((m[410]&~m[411]&~m[412]&~m[414]&~m[415])|(~m[410]&m[411]&~m[412]&~m[414]&~m[415])|(~m[410]&~m[411]&m[412]&~m[414]&~m[415])|(m[410]&m[411]&m[412]&m[414]&~m[415])|(~m[410]&~m[411]&~m[412]&~m[414]&m[415])|(m[410]&m[411]&~m[412]&m[414]&m[415])|(m[410]&~m[411]&m[412]&m[414]&m[415])|(~m[410]&m[411]&m[412]&m[414]&m[415]))&UnbiasedRNG[286])|((m[410]&m[411]&~m[412]&~m[414]&~m[415])|(m[410]&~m[411]&m[412]&~m[414]&~m[415])|(~m[410]&m[411]&m[412]&~m[414]&~m[415])|(m[410]&m[411]&m[412]&~m[414]&~m[415])|(m[410]&~m[411]&~m[412]&~m[414]&m[415])|(~m[410]&m[411]&~m[412]&~m[414]&m[415])|(m[410]&m[411]&~m[412]&~m[414]&m[415])|(~m[410]&~m[411]&m[412]&~m[414]&m[415])|(m[410]&~m[411]&m[412]&~m[414]&m[415])|(~m[410]&m[411]&m[412]&~m[414]&m[415])|(m[410]&m[411]&m[412]&~m[414]&m[415])|(m[410]&m[411]&m[412]&m[414]&m[415]));
    m[418] = (((m[415]&~m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&~m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&m[419]&~m[420])|(~m[415]&~m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&m[419]&m[420])|(m[415]&~m[416]&m[417]&m[419]&m[420])|(~m[415]&m[416]&m[417]&m[419]&m[420]))&UnbiasedRNG[287])|((m[415]&m[416]&~m[417]&~m[419]&~m[420])|(m[415]&~m[416]&m[417]&~m[419]&~m[420])|(~m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&~m[416]&~m[417]&~m[419]&m[420])|(~m[415]&m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&~m[419]&m[420])|(~m[415]&~m[416]&m[417]&~m[419]&m[420])|(m[415]&~m[416]&m[417]&~m[419]&m[420])|(~m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&m[419]&m[420]));
    m[423] = (((m[420]&~m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&~m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&m[424]&~m[425])|(~m[420]&~m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&m[424]&m[425])|(m[420]&~m[421]&m[422]&m[424]&m[425])|(~m[420]&m[421]&m[422]&m[424]&m[425]))&UnbiasedRNG[288])|((m[420]&m[421]&~m[422]&~m[424]&~m[425])|(m[420]&~m[421]&m[422]&~m[424]&~m[425])|(~m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&~m[421]&~m[422]&~m[424]&m[425])|(~m[420]&m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&~m[424]&m[425])|(~m[420]&~m[421]&m[422]&~m[424]&m[425])|(m[420]&~m[421]&m[422]&~m[424]&m[425])|(~m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&m[424]&m[425]));
    m[428] = (((m[425]&~m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&~m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&m[429]&~m[430])|(~m[425]&~m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&m[429]&m[430])|(m[425]&~m[426]&m[427]&m[429]&m[430])|(~m[425]&m[426]&m[427]&m[429]&m[430]))&UnbiasedRNG[289])|((m[425]&m[426]&~m[427]&~m[429]&~m[430])|(m[425]&~m[426]&m[427]&~m[429]&~m[430])|(~m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&~m[426]&~m[427]&~m[429]&m[430])|(~m[425]&m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&~m[429]&m[430])|(~m[425]&~m[426]&m[427]&~m[429]&m[430])|(m[425]&~m[426]&m[427]&~m[429]&m[430])|(~m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&m[429]&m[430]));
    m[438] = (((m[435]&~m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&~m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&m[439]&~m[440])|(~m[435]&~m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&m[439]&m[440])|(m[435]&~m[436]&m[437]&m[439]&m[440])|(~m[435]&m[436]&m[437]&m[439]&m[440]))&UnbiasedRNG[290])|((m[435]&m[436]&~m[437]&~m[439]&~m[440])|(m[435]&~m[436]&m[437]&~m[439]&~m[440])|(~m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&~m[436]&~m[437]&~m[439]&m[440])|(~m[435]&m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&~m[439]&m[440])|(~m[435]&~m[436]&m[437]&~m[439]&m[440])|(m[435]&~m[436]&m[437]&~m[439]&m[440])|(~m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&m[439]&m[440]));
    m[443] = (((m[440]&~m[441]&~m[442]&~m[444]&~m[445])|(~m[440]&m[441]&~m[442]&~m[444]&~m[445])|(~m[440]&~m[441]&m[442]&~m[444]&~m[445])|(m[440]&m[441]&m[442]&m[444]&~m[445])|(~m[440]&~m[441]&~m[442]&~m[444]&m[445])|(m[440]&m[441]&~m[442]&m[444]&m[445])|(m[440]&~m[441]&m[442]&m[444]&m[445])|(~m[440]&m[441]&m[442]&m[444]&m[445]))&UnbiasedRNG[291])|((m[440]&m[441]&~m[442]&~m[444]&~m[445])|(m[440]&~m[441]&m[442]&~m[444]&~m[445])|(~m[440]&m[441]&m[442]&~m[444]&~m[445])|(m[440]&m[441]&m[442]&~m[444]&~m[445])|(m[440]&~m[441]&~m[442]&~m[444]&m[445])|(~m[440]&m[441]&~m[442]&~m[444]&m[445])|(m[440]&m[441]&~m[442]&~m[444]&m[445])|(~m[440]&~m[441]&m[442]&~m[444]&m[445])|(m[440]&~m[441]&m[442]&~m[444]&m[445])|(~m[440]&m[441]&m[442]&~m[444]&m[445])|(m[440]&m[441]&m[442]&~m[444]&m[445])|(m[440]&m[441]&m[442]&m[444]&m[445]));
    m[448] = (((m[445]&~m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&~m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&m[449]&~m[450])|(~m[445]&~m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&m[449]&m[450])|(m[445]&~m[446]&m[447]&m[449]&m[450])|(~m[445]&m[446]&m[447]&m[449]&m[450]))&UnbiasedRNG[292])|((m[445]&m[446]&~m[447]&~m[449]&~m[450])|(m[445]&~m[446]&m[447]&~m[449]&~m[450])|(~m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&~m[446]&~m[447]&~m[449]&m[450])|(~m[445]&m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&~m[449]&m[450])|(~m[445]&~m[446]&m[447]&~m[449]&m[450])|(m[445]&~m[446]&m[447]&~m[449]&m[450])|(~m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&m[449]&m[450]));
    m[453] = (((m[450]&~m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&~m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&m[454]&~m[455])|(~m[450]&~m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&m[454]&m[455])|(m[450]&~m[451]&m[452]&m[454]&m[455])|(~m[450]&m[451]&m[452]&m[454]&m[455]))&UnbiasedRNG[293])|((m[450]&m[451]&~m[452]&~m[454]&~m[455])|(m[450]&~m[451]&m[452]&~m[454]&~m[455])|(~m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&~m[451]&~m[452]&~m[454]&m[455])|(~m[450]&m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&~m[454]&m[455])|(~m[450]&~m[451]&m[452]&~m[454]&m[455])|(m[450]&~m[451]&m[452]&~m[454]&m[455])|(~m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&m[454]&m[455]));
    m[458] = (((m[455]&~m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&~m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&m[459]&~m[460])|(~m[455]&~m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&m[459]&m[460])|(m[455]&~m[456]&m[457]&m[459]&m[460])|(~m[455]&m[456]&m[457]&m[459]&m[460]))&UnbiasedRNG[294])|((m[455]&m[456]&~m[457]&~m[459]&~m[460])|(m[455]&~m[456]&m[457]&~m[459]&~m[460])|(~m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&~m[456]&~m[457]&~m[459]&m[460])|(~m[455]&m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&~m[459]&m[460])|(~m[455]&~m[456]&m[457]&~m[459]&m[460])|(m[455]&~m[456]&m[457]&~m[459]&m[460])|(~m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&m[459]&m[460]));
    m[468] = (((m[465]&~m[466]&~m[467]&~m[469]&~m[470])|(~m[465]&m[466]&~m[467]&~m[469]&~m[470])|(~m[465]&~m[466]&m[467]&~m[469]&~m[470])|(m[465]&m[466]&m[467]&m[469]&~m[470])|(~m[465]&~m[466]&~m[467]&~m[469]&m[470])|(m[465]&m[466]&~m[467]&m[469]&m[470])|(m[465]&~m[466]&m[467]&m[469]&m[470])|(~m[465]&m[466]&m[467]&m[469]&m[470]))&UnbiasedRNG[295])|((m[465]&m[466]&~m[467]&~m[469]&~m[470])|(m[465]&~m[466]&m[467]&~m[469]&~m[470])|(~m[465]&m[466]&m[467]&~m[469]&~m[470])|(m[465]&m[466]&m[467]&~m[469]&~m[470])|(m[465]&~m[466]&~m[467]&~m[469]&m[470])|(~m[465]&m[466]&~m[467]&~m[469]&m[470])|(m[465]&m[466]&~m[467]&~m[469]&m[470])|(~m[465]&~m[466]&m[467]&~m[469]&m[470])|(m[465]&~m[466]&m[467]&~m[469]&m[470])|(~m[465]&m[466]&m[467]&~m[469]&m[470])|(m[465]&m[466]&m[467]&~m[469]&m[470])|(m[465]&m[466]&m[467]&m[469]&m[470]));
    m[473] = (((m[470]&~m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&~m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&m[474]&~m[475])|(~m[470]&~m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&m[474]&m[475])|(m[470]&~m[471]&m[472]&m[474]&m[475])|(~m[470]&m[471]&m[472]&m[474]&m[475]))&UnbiasedRNG[296])|((m[470]&m[471]&~m[472]&~m[474]&~m[475])|(m[470]&~m[471]&m[472]&~m[474]&~m[475])|(~m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&~m[471]&~m[472]&~m[474]&m[475])|(~m[470]&m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&~m[474]&m[475])|(~m[470]&~m[471]&m[472]&~m[474]&m[475])|(m[470]&~m[471]&m[472]&~m[474]&m[475])|(~m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&m[474]&m[475]));
    m[478] = (((m[475]&~m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&~m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&m[479]&~m[480])|(~m[475]&~m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&m[479]&m[480])|(m[475]&~m[476]&m[477]&m[479]&m[480])|(~m[475]&m[476]&m[477]&m[479]&m[480]))&UnbiasedRNG[297])|((m[475]&m[476]&~m[477]&~m[479]&~m[480])|(m[475]&~m[476]&m[477]&~m[479]&~m[480])|(~m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&~m[476]&~m[477]&~m[479]&m[480])|(~m[475]&m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&~m[479]&m[480])|(~m[475]&~m[476]&m[477]&~m[479]&m[480])|(m[475]&~m[476]&m[477]&~m[479]&m[480])|(~m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&m[479]&m[480]));
    m[483] = (((m[480]&~m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&~m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&m[484]&~m[485])|(~m[480]&~m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&m[484]&m[485])|(m[480]&~m[481]&m[482]&m[484]&m[485])|(~m[480]&m[481]&m[482]&m[484]&m[485]))&UnbiasedRNG[298])|((m[480]&m[481]&~m[482]&~m[484]&~m[485])|(m[480]&~m[481]&m[482]&~m[484]&~m[485])|(~m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&~m[481]&~m[482]&~m[484]&m[485])|(~m[480]&m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&~m[484]&m[485])|(~m[480]&~m[481]&m[482]&~m[484]&m[485])|(m[480]&~m[481]&m[482]&~m[484]&m[485])|(~m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&m[484]&m[485]));
    m[488] = (((m[485]&~m[486]&~m[487]&~m[489]&~m[490])|(~m[485]&m[486]&~m[487]&~m[489]&~m[490])|(~m[485]&~m[486]&m[487]&~m[489]&~m[490])|(m[485]&m[486]&m[487]&m[489]&~m[490])|(~m[485]&~m[486]&~m[487]&~m[489]&m[490])|(m[485]&m[486]&~m[487]&m[489]&m[490])|(m[485]&~m[486]&m[487]&m[489]&m[490])|(~m[485]&m[486]&m[487]&m[489]&m[490]))&UnbiasedRNG[299])|((m[485]&m[486]&~m[487]&~m[489]&~m[490])|(m[485]&~m[486]&m[487]&~m[489]&~m[490])|(~m[485]&m[486]&m[487]&~m[489]&~m[490])|(m[485]&m[486]&m[487]&~m[489]&~m[490])|(m[485]&~m[486]&~m[487]&~m[489]&m[490])|(~m[485]&m[486]&~m[487]&~m[489]&m[490])|(m[485]&m[486]&~m[487]&~m[489]&m[490])|(~m[485]&~m[486]&m[487]&~m[489]&m[490])|(m[485]&~m[486]&m[487]&~m[489]&m[490])|(~m[485]&m[486]&m[487]&~m[489]&m[490])|(m[485]&m[486]&m[487]&~m[489]&m[490])|(m[485]&m[486]&m[487]&m[489]&m[490]));
    m[493] = (((m[490]&~m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&~m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&m[494]&~m[495])|(~m[490]&~m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&m[494]&m[495])|(m[490]&~m[491]&m[492]&m[494]&m[495])|(~m[490]&m[491]&m[492]&m[494]&m[495]))&UnbiasedRNG[300])|((m[490]&m[491]&~m[492]&~m[494]&~m[495])|(m[490]&~m[491]&m[492]&~m[494]&~m[495])|(~m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&~m[491]&~m[492]&~m[494]&m[495])|(~m[490]&m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&~m[494]&m[495])|(~m[490]&~m[491]&m[492]&~m[494]&m[495])|(m[490]&~m[491]&m[492]&~m[494]&m[495])|(~m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&m[494]&m[495]));
    m[503] = (((m[500]&~m[501]&~m[502]&~m[504]&~m[505])|(~m[500]&m[501]&~m[502]&~m[504]&~m[505])|(~m[500]&~m[501]&m[502]&~m[504]&~m[505])|(m[500]&m[501]&m[502]&m[504]&~m[505])|(~m[500]&~m[501]&~m[502]&~m[504]&m[505])|(m[500]&m[501]&~m[502]&m[504]&m[505])|(m[500]&~m[501]&m[502]&m[504]&m[505])|(~m[500]&m[501]&m[502]&m[504]&m[505]))&UnbiasedRNG[301])|((m[500]&m[501]&~m[502]&~m[504]&~m[505])|(m[500]&~m[501]&m[502]&~m[504]&~m[505])|(~m[500]&m[501]&m[502]&~m[504]&~m[505])|(m[500]&m[501]&m[502]&~m[504]&~m[505])|(m[500]&~m[501]&~m[502]&~m[504]&m[505])|(~m[500]&m[501]&~m[502]&~m[504]&m[505])|(m[500]&m[501]&~m[502]&~m[504]&m[505])|(~m[500]&~m[501]&m[502]&~m[504]&m[505])|(m[500]&~m[501]&m[502]&~m[504]&m[505])|(~m[500]&m[501]&m[502]&~m[504]&m[505])|(m[500]&m[501]&m[502]&~m[504]&m[505])|(m[500]&m[501]&m[502]&m[504]&m[505]));
    m[508] = (((m[505]&~m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&~m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&m[509]&~m[510])|(~m[505]&~m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&m[509]&m[510])|(m[505]&~m[506]&m[507]&m[509]&m[510])|(~m[505]&m[506]&m[507]&m[509]&m[510]))&UnbiasedRNG[302])|((m[505]&m[506]&~m[507]&~m[509]&~m[510])|(m[505]&~m[506]&m[507]&~m[509]&~m[510])|(~m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&~m[506]&~m[507]&~m[509]&m[510])|(~m[505]&m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&~m[509]&m[510])|(~m[505]&~m[506]&m[507]&~m[509]&m[510])|(m[505]&~m[506]&m[507]&~m[509]&m[510])|(~m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&m[509]&m[510]));
    m[513] = (((m[510]&~m[511]&~m[512]&~m[514]&~m[515])|(~m[510]&m[511]&~m[512]&~m[514]&~m[515])|(~m[510]&~m[511]&m[512]&~m[514]&~m[515])|(m[510]&m[511]&m[512]&m[514]&~m[515])|(~m[510]&~m[511]&~m[512]&~m[514]&m[515])|(m[510]&m[511]&~m[512]&m[514]&m[515])|(m[510]&~m[511]&m[512]&m[514]&m[515])|(~m[510]&m[511]&m[512]&m[514]&m[515]))&UnbiasedRNG[303])|((m[510]&m[511]&~m[512]&~m[514]&~m[515])|(m[510]&~m[511]&m[512]&~m[514]&~m[515])|(~m[510]&m[511]&m[512]&~m[514]&~m[515])|(m[510]&m[511]&m[512]&~m[514]&~m[515])|(m[510]&~m[511]&~m[512]&~m[514]&m[515])|(~m[510]&m[511]&~m[512]&~m[514]&m[515])|(m[510]&m[511]&~m[512]&~m[514]&m[515])|(~m[510]&~m[511]&m[512]&~m[514]&m[515])|(m[510]&~m[511]&m[512]&~m[514]&m[515])|(~m[510]&m[511]&m[512]&~m[514]&m[515])|(m[510]&m[511]&m[512]&~m[514]&m[515])|(m[510]&m[511]&m[512]&m[514]&m[515]));
    m[518] = (((m[515]&~m[516]&~m[517]&~m[519]&~m[520])|(~m[515]&m[516]&~m[517]&~m[519]&~m[520])|(~m[515]&~m[516]&m[517]&~m[519]&~m[520])|(m[515]&m[516]&m[517]&m[519]&~m[520])|(~m[515]&~m[516]&~m[517]&~m[519]&m[520])|(m[515]&m[516]&~m[517]&m[519]&m[520])|(m[515]&~m[516]&m[517]&m[519]&m[520])|(~m[515]&m[516]&m[517]&m[519]&m[520]))&UnbiasedRNG[304])|((m[515]&m[516]&~m[517]&~m[519]&~m[520])|(m[515]&~m[516]&m[517]&~m[519]&~m[520])|(~m[515]&m[516]&m[517]&~m[519]&~m[520])|(m[515]&m[516]&m[517]&~m[519]&~m[520])|(m[515]&~m[516]&~m[517]&~m[519]&m[520])|(~m[515]&m[516]&~m[517]&~m[519]&m[520])|(m[515]&m[516]&~m[517]&~m[519]&m[520])|(~m[515]&~m[516]&m[517]&~m[519]&m[520])|(m[515]&~m[516]&m[517]&~m[519]&m[520])|(~m[515]&m[516]&m[517]&~m[519]&m[520])|(m[515]&m[516]&m[517]&~m[519]&m[520])|(m[515]&m[516]&m[517]&m[519]&m[520]));
    m[523] = (((m[520]&~m[521]&~m[522]&~m[524]&~m[525])|(~m[520]&m[521]&~m[522]&~m[524]&~m[525])|(~m[520]&~m[521]&m[522]&~m[524]&~m[525])|(m[520]&m[521]&m[522]&m[524]&~m[525])|(~m[520]&~m[521]&~m[522]&~m[524]&m[525])|(m[520]&m[521]&~m[522]&m[524]&m[525])|(m[520]&~m[521]&m[522]&m[524]&m[525])|(~m[520]&m[521]&m[522]&m[524]&m[525]))&UnbiasedRNG[305])|((m[520]&m[521]&~m[522]&~m[524]&~m[525])|(m[520]&~m[521]&m[522]&~m[524]&~m[525])|(~m[520]&m[521]&m[522]&~m[524]&~m[525])|(m[520]&m[521]&m[522]&~m[524]&~m[525])|(m[520]&~m[521]&~m[522]&~m[524]&m[525])|(~m[520]&m[521]&~m[522]&~m[524]&m[525])|(m[520]&m[521]&~m[522]&~m[524]&m[525])|(~m[520]&~m[521]&m[522]&~m[524]&m[525])|(m[520]&~m[521]&m[522]&~m[524]&m[525])|(~m[520]&m[521]&m[522]&~m[524]&m[525])|(m[520]&m[521]&m[522]&~m[524]&m[525])|(m[520]&m[521]&m[522]&m[524]&m[525]));
    m[528] = (((m[525]&~m[526]&~m[527]&~m[529]&~m[530])|(~m[525]&m[526]&~m[527]&~m[529]&~m[530])|(~m[525]&~m[526]&m[527]&~m[529]&~m[530])|(m[525]&m[526]&m[527]&m[529]&~m[530])|(~m[525]&~m[526]&~m[527]&~m[529]&m[530])|(m[525]&m[526]&~m[527]&m[529]&m[530])|(m[525]&~m[526]&m[527]&m[529]&m[530])|(~m[525]&m[526]&m[527]&m[529]&m[530]))&UnbiasedRNG[306])|((m[525]&m[526]&~m[527]&~m[529]&~m[530])|(m[525]&~m[526]&m[527]&~m[529]&~m[530])|(~m[525]&m[526]&m[527]&~m[529]&~m[530])|(m[525]&m[526]&m[527]&~m[529]&~m[530])|(m[525]&~m[526]&~m[527]&~m[529]&m[530])|(~m[525]&m[526]&~m[527]&~m[529]&m[530])|(m[525]&m[526]&~m[527]&~m[529]&m[530])|(~m[525]&~m[526]&m[527]&~m[529]&m[530])|(m[525]&~m[526]&m[527]&~m[529]&m[530])|(~m[525]&m[526]&m[527]&~m[529]&m[530])|(m[525]&m[526]&m[527]&~m[529]&m[530])|(m[525]&m[526]&m[527]&m[529]&m[530]));
    m[533] = (((m[530]&~m[531]&~m[532]&~m[534]&~m[535])|(~m[530]&m[531]&~m[532]&~m[534]&~m[535])|(~m[530]&~m[531]&m[532]&~m[534]&~m[535])|(m[530]&m[531]&m[532]&m[534]&~m[535])|(~m[530]&~m[531]&~m[532]&~m[534]&m[535])|(m[530]&m[531]&~m[532]&m[534]&m[535])|(m[530]&~m[531]&m[532]&m[534]&m[535])|(~m[530]&m[531]&m[532]&m[534]&m[535]))&UnbiasedRNG[307])|((m[530]&m[531]&~m[532]&~m[534]&~m[535])|(m[530]&~m[531]&m[532]&~m[534]&~m[535])|(~m[530]&m[531]&m[532]&~m[534]&~m[535])|(m[530]&m[531]&m[532]&~m[534]&~m[535])|(m[530]&~m[531]&~m[532]&~m[534]&m[535])|(~m[530]&m[531]&~m[532]&~m[534]&m[535])|(m[530]&m[531]&~m[532]&~m[534]&m[535])|(~m[530]&~m[531]&m[532]&~m[534]&m[535])|(m[530]&~m[531]&m[532]&~m[534]&m[535])|(~m[530]&m[531]&m[532]&~m[534]&m[535])|(m[530]&m[531]&m[532]&~m[534]&m[535])|(m[530]&m[531]&m[532]&m[534]&m[535]));
    m[543] = (((m[540]&~m[541]&~m[542]&~m[544]&~m[545])|(~m[540]&m[541]&~m[542]&~m[544]&~m[545])|(~m[540]&~m[541]&m[542]&~m[544]&~m[545])|(m[540]&m[541]&m[542]&m[544]&~m[545])|(~m[540]&~m[541]&~m[542]&~m[544]&m[545])|(m[540]&m[541]&~m[542]&m[544]&m[545])|(m[540]&~m[541]&m[542]&m[544]&m[545])|(~m[540]&m[541]&m[542]&m[544]&m[545]))&UnbiasedRNG[308])|((m[540]&m[541]&~m[542]&~m[544]&~m[545])|(m[540]&~m[541]&m[542]&~m[544]&~m[545])|(~m[540]&m[541]&m[542]&~m[544]&~m[545])|(m[540]&m[541]&m[542]&~m[544]&~m[545])|(m[540]&~m[541]&~m[542]&~m[544]&m[545])|(~m[540]&m[541]&~m[542]&~m[544]&m[545])|(m[540]&m[541]&~m[542]&~m[544]&m[545])|(~m[540]&~m[541]&m[542]&~m[544]&m[545])|(m[540]&~m[541]&m[542]&~m[544]&m[545])|(~m[540]&m[541]&m[542]&~m[544]&m[545])|(m[540]&m[541]&m[542]&~m[544]&m[545])|(m[540]&m[541]&m[542]&m[544]&m[545]));
    m[548] = (((m[545]&~m[546]&~m[547]&~m[549]&~m[550])|(~m[545]&m[546]&~m[547]&~m[549]&~m[550])|(~m[545]&~m[546]&m[547]&~m[549]&~m[550])|(m[545]&m[546]&m[547]&m[549]&~m[550])|(~m[545]&~m[546]&~m[547]&~m[549]&m[550])|(m[545]&m[546]&~m[547]&m[549]&m[550])|(m[545]&~m[546]&m[547]&m[549]&m[550])|(~m[545]&m[546]&m[547]&m[549]&m[550]))&UnbiasedRNG[309])|((m[545]&m[546]&~m[547]&~m[549]&~m[550])|(m[545]&~m[546]&m[547]&~m[549]&~m[550])|(~m[545]&m[546]&m[547]&~m[549]&~m[550])|(m[545]&m[546]&m[547]&~m[549]&~m[550])|(m[545]&~m[546]&~m[547]&~m[549]&m[550])|(~m[545]&m[546]&~m[547]&~m[549]&m[550])|(m[545]&m[546]&~m[547]&~m[549]&m[550])|(~m[545]&~m[546]&m[547]&~m[549]&m[550])|(m[545]&~m[546]&m[547]&~m[549]&m[550])|(~m[545]&m[546]&m[547]&~m[549]&m[550])|(m[545]&m[546]&m[547]&~m[549]&m[550])|(m[545]&m[546]&m[547]&m[549]&m[550]));
    m[553] = (((m[550]&~m[551]&~m[552]&~m[554]&~m[555])|(~m[550]&m[551]&~m[552]&~m[554]&~m[555])|(~m[550]&~m[551]&m[552]&~m[554]&~m[555])|(m[550]&m[551]&m[552]&m[554]&~m[555])|(~m[550]&~m[551]&~m[552]&~m[554]&m[555])|(m[550]&m[551]&~m[552]&m[554]&m[555])|(m[550]&~m[551]&m[552]&m[554]&m[555])|(~m[550]&m[551]&m[552]&m[554]&m[555]))&UnbiasedRNG[310])|((m[550]&m[551]&~m[552]&~m[554]&~m[555])|(m[550]&~m[551]&m[552]&~m[554]&~m[555])|(~m[550]&m[551]&m[552]&~m[554]&~m[555])|(m[550]&m[551]&m[552]&~m[554]&~m[555])|(m[550]&~m[551]&~m[552]&~m[554]&m[555])|(~m[550]&m[551]&~m[552]&~m[554]&m[555])|(m[550]&m[551]&~m[552]&~m[554]&m[555])|(~m[550]&~m[551]&m[552]&~m[554]&m[555])|(m[550]&~m[551]&m[552]&~m[554]&m[555])|(~m[550]&m[551]&m[552]&~m[554]&m[555])|(m[550]&m[551]&m[552]&~m[554]&m[555])|(m[550]&m[551]&m[552]&m[554]&m[555]));
    m[558] = (((m[555]&~m[556]&~m[557]&~m[559]&~m[560])|(~m[555]&m[556]&~m[557]&~m[559]&~m[560])|(~m[555]&~m[556]&m[557]&~m[559]&~m[560])|(m[555]&m[556]&m[557]&m[559]&~m[560])|(~m[555]&~m[556]&~m[557]&~m[559]&m[560])|(m[555]&m[556]&~m[557]&m[559]&m[560])|(m[555]&~m[556]&m[557]&m[559]&m[560])|(~m[555]&m[556]&m[557]&m[559]&m[560]))&UnbiasedRNG[311])|((m[555]&m[556]&~m[557]&~m[559]&~m[560])|(m[555]&~m[556]&m[557]&~m[559]&~m[560])|(~m[555]&m[556]&m[557]&~m[559]&~m[560])|(m[555]&m[556]&m[557]&~m[559]&~m[560])|(m[555]&~m[556]&~m[557]&~m[559]&m[560])|(~m[555]&m[556]&~m[557]&~m[559]&m[560])|(m[555]&m[556]&~m[557]&~m[559]&m[560])|(~m[555]&~m[556]&m[557]&~m[559]&m[560])|(m[555]&~m[556]&m[557]&~m[559]&m[560])|(~m[555]&m[556]&m[557]&~m[559]&m[560])|(m[555]&m[556]&m[557]&~m[559]&m[560])|(m[555]&m[556]&m[557]&m[559]&m[560]));
    m[563] = (((m[560]&~m[561]&~m[562]&~m[564]&~m[565])|(~m[560]&m[561]&~m[562]&~m[564]&~m[565])|(~m[560]&~m[561]&m[562]&~m[564]&~m[565])|(m[560]&m[561]&m[562]&m[564]&~m[565])|(~m[560]&~m[561]&~m[562]&~m[564]&m[565])|(m[560]&m[561]&~m[562]&m[564]&m[565])|(m[560]&~m[561]&m[562]&m[564]&m[565])|(~m[560]&m[561]&m[562]&m[564]&m[565]))&UnbiasedRNG[312])|((m[560]&m[561]&~m[562]&~m[564]&~m[565])|(m[560]&~m[561]&m[562]&~m[564]&~m[565])|(~m[560]&m[561]&m[562]&~m[564]&~m[565])|(m[560]&m[561]&m[562]&~m[564]&~m[565])|(m[560]&~m[561]&~m[562]&~m[564]&m[565])|(~m[560]&m[561]&~m[562]&~m[564]&m[565])|(m[560]&m[561]&~m[562]&~m[564]&m[565])|(~m[560]&~m[561]&m[562]&~m[564]&m[565])|(m[560]&~m[561]&m[562]&~m[564]&m[565])|(~m[560]&m[561]&m[562]&~m[564]&m[565])|(m[560]&m[561]&m[562]&~m[564]&m[565])|(m[560]&m[561]&m[562]&m[564]&m[565]));
    m[568] = (((m[565]&~m[566]&~m[567]&~m[569]&~m[570])|(~m[565]&m[566]&~m[567]&~m[569]&~m[570])|(~m[565]&~m[566]&m[567]&~m[569]&~m[570])|(m[565]&m[566]&m[567]&m[569]&~m[570])|(~m[565]&~m[566]&~m[567]&~m[569]&m[570])|(m[565]&m[566]&~m[567]&m[569]&m[570])|(m[565]&~m[566]&m[567]&m[569]&m[570])|(~m[565]&m[566]&m[567]&m[569]&m[570]))&UnbiasedRNG[313])|((m[565]&m[566]&~m[567]&~m[569]&~m[570])|(m[565]&~m[566]&m[567]&~m[569]&~m[570])|(~m[565]&m[566]&m[567]&~m[569]&~m[570])|(m[565]&m[566]&m[567]&~m[569]&~m[570])|(m[565]&~m[566]&~m[567]&~m[569]&m[570])|(~m[565]&m[566]&~m[567]&~m[569]&m[570])|(m[565]&m[566]&~m[567]&~m[569]&m[570])|(~m[565]&~m[566]&m[567]&~m[569]&m[570])|(m[565]&~m[566]&m[567]&~m[569]&m[570])|(~m[565]&m[566]&m[567]&~m[569]&m[570])|(m[565]&m[566]&m[567]&~m[569]&m[570])|(m[565]&m[566]&m[567]&m[569]&m[570]));
    m[573] = (((m[570]&~m[571]&~m[572]&~m[574]&~m[575])|(~m[570]&m[571]&~m[572]&~m[574]&~m[575])|(~m[570]&~m[571]&m[572]&~m[574]&~m[575])|(m[570]&m[571]&m[572]&m[574]&~m[575])|(~m[570]&~m[571]&~m[572]&~m[574]&m[575])|(m[570]&m[571]&~m[572]&m[574]&m[575])|(m[570]&~m[571]&m[572]&m[574]&m[575])|(~m[570]&m[571]&m[572]&m[574]&m[575]))&UnbiasedRNG[314])|((m[570]&m[571]&~m[572]&~m[574]&~m[575])|(m[570]&~m[571]&m[572]&~m[574]&~m[575])|(~m[570]&m[571]&m[572]&~m[574]&~m[575])|(m[570]&m[571]&m[572]&~m[574]&~m[575])|(m[570]&~m[571]&~m[572]&~m[574]&m[575])|(~m[570]&m[571]&~m[572]&~m[574]&m[575])|(m[570]&m[571]&~m[572]&~m[574]&m[575])|(~m[570]&~m[571]&m[572]&~m[574]&m[575])|(m[570]&~m[571]&m[572]&~m[574]&m[575])|(~m[570]&m[571]&m[572]&~m[574]&m[575])|(m[570]&m[571]&m[572]&~m[574]&m[575])|(m[570]&m[571]&m[572]&m[574]&m[575]));
    m[578] = (((m[575]&~m[576]&~m[577]&~m[579]&~m[580])|(~m[575]&m[576]&~m[577]&~m[579]&~m[580])|(~m[575]&~m[576]&m[577]&~m[579]&~m[580])|(m[575]&m[576]&m[577]&m[579]&~m[580])|(~m[575]&~m[576]&~m[577]&~m[579]&m[580])|(m[575]&m[576]&~m[577]&m[579]&m[580])|(m[575]&~m[576]&m[577]&m[579]&m[580])|(~m[575]&m[576]&m[577]&m[579]&m[580]))&UnbiasedRNG[315])|((m[575]&m[576]&~m[577]&~m[579]&~m[580])|(m[575]&~m[576]&m[577]&~m[579]&~m[580])|(~m[575]&m[576]&m[577]&~m[579]&~m[580])|(m[575]&m[576]&m[577]&~m[579]&~m[580])|(m[575]&~m[576]&~m[577]&~m[579]&m[580])|(~m[575]&m[576]&~m[577]&~m[579]&m[580])|(m[575]&m[576]&~m[577]&~m[579]&m[580])|(~m[575]&~m[576]&m[577]&~m[579]&m[580])|(m[575]&~m[576]&m[577]&~m[579]&m[580])|(~m[575]&m[576]&m[577]&~m[579]&m[580])|(m[575]&m[576]&m[577]&~m[579]&m[580])|(m[575]&m[576]&m[577]&m[579]&m[580]));
    m[588] = (((m[585]&~m[586]&~m[587]&~m[589]&~m[590])|(~m[585]&m[586]&~m[587]&~m[589]&~m[590])|(~m[585]&~m[586]&m[587]&~m[589]&~m[590])|(m[585]&m[586]&m[587]&m[589]&~m[590])|(~m[585]&~m[586]&~m[587]&~m[589]&m[590])|(m[585]&m[586]&~m[587]&m[589]&m[590])|(m[585]&~m[586]&m[587]&m[589]&m[590])|(~m[585]&m[586]&m[587]&m[589]&m[590]))&UnbiasedRNG[316])|((m[585]&m[586]&~m[587]&~m[589]&~m[590])|(m[585]&~m[586]&m[587]&~m[589]&~m[590])|(~m[585]&m[586]&m[587]&~m[589]&~m[590])|(m[585]&m[586]&m[587]&~m[589]&~m[590])|(m[585]&~m[586]&~m[587]&~m[589]&m[590])|(~m[585]&m[586]&~m[587]&~m[589]&m[590])|(m[585]&m[586]&~m[587]&~m[589]&m[590])|(~m[585]&~m[586]&m[587]&~m[589]&m[590])|(m[585]&~m[586]&m[587]&~m[589]&m[590])|(~m[585]&m[586]&m[587]&~m[589]&m[590])|(m[585]&m[586]&m[587]&~m[589]&m[590])|(m[585]&m[586]&m[587]&m[589]&m[590]));
    m[593] = (((m[590]&~m[591]&~m[592]&~m[594]&~m[595])|(~m[590]&m[591]&~m[592]&~m[594]&~m[595])|(~m[590]&~m[591]&m[592]&~m[594]&~m[595])|(m[590]&m[591]&m[592]&m[594]&~m[595])|(~m[590]&~m[591]&~m[592]&~m[594]&m[595])|(m[590]&m[591]&~m[592]&m[594]&m[595])|(m[590]&~m[591]&m[592]&m[594]&m[595])|(~m[590]&m[591]&m[592]&m[594]&m[595]))&UnbiasedRNG[317])|((m[590]&m[591]&~m[592]&~m[594]&~m[595])|(m[590]&~m[591]&m[592]&~m[594]&~m[595])|(~m[590]&m[591]&m[592]&~m[594]&~m[595])|(m[590]&m[591]&m[592]&~m[594]&~m[595])|(m[590]&~m[591]&~m[592]&~m[594]&m[595])|(~m[590]&m[591]&~m[592]&~m[594]&m[595])|(m[590]&m[591]&~m[592]&~m[594]&m[595])|(~m[590]&~m[591]&m[592]&~m[594]&m[595])|(m[590]&~m[591]&m[592]&~m[594]&m[595])|(~m[590]&m[591]&m[592]&~m[594]&m[595])|(m[590]&m[591]&m[592]&~m[594]&m[595])|(m[590]&m[591]&m[592]&m[594]&m[595]));
    m[598] = (((m[595]&~m[596]&~m[597]&~m[599]&~m[600])|(~m[595]&m[596]&~m[597]&~m[599]&~m[600])|(~m[595]&~m[596]&m[597]&~m[599]&~m[600])|(m[595]&m[596]&m[597]&m[599]&~m[600])|(~m[595]&~m[596]&~m[597]&~m[599]&m[600])|(m[595]&m[596]&~m[597]&m[599]&m[600])|(m[595]&~m[596]&m[597]&m[599]&m[600])|(~m[595]&m[596]&m[597]&m[599]&m[600]))&UnbiasedRNG[318])|((m[595]&m[596]&~m[597]&~m[599]&~m[600])|(m[595]&~m[596]&m[597]&~m[599]&~m[600])|(~m[595]&m[596]&m[597]&~m[599]&~m[600])|(m[595]&m[596]&m[597]&~m[599]&~m[600])|(m[595]&~m[596]&~m[597]&~m[599]&m[600])|(~m[595]&m[596]&~m[597]&~m[599]&m[600])|(m[595]&m[596]&~m[597]&~m[599]&m[600])|(~m[595]&~m[596]&m[597]&~m[599]&m[600])|(m[595]&~m[596]&m[597]&~m[599]&m[600])|(~m[595]&m[596]&m[597]&~m[599]&m[600])|(m[595]&m[596]&m[597]&~m[599]&m[600])|(m[595]&m[596]&m[597]&m[599]&m[600]));
    m[603] = (((m[600]&~m[601]&~m[602]&~m[604]&~m[605])|(~m[600]&m[601]&~m[602]&~m[604]&~m[605])|(~m[600]&~m[601]&m[602]&~m[604]&~m[605])|(m[600]&m[601]&m[602]&m[604]&~m[605])|(~m[600]&~m[601]&~m[602]&~m[604]&m[605])|(m[600]&m[601]&~m[602]&m[604]&m[605])|(m[600]&~m[601]&m[602]&m[604]&m[605])|(~m[600]&m[601]&m[602]&m[604]&m[605]))&UnbiasedRNG[319])|((m[600]&m[601]&~m[602]&~m[604]&~m[605])|(m[600]&~m[601]&m[602]&~m[604]&~m[605])|(~m[600]&m[601]&m[602]&~m[604]&~m[605])|(m[600]&m[601]&m[602]&~m[604]&~m[605])|(m[600]&~m[601]&~m[602]&~m[604]&m[605])|(~m[600]&m[601]&~m[602]&~m[604]&m[605])|(m[600]&m[601]&~m[602]&~m[604]&m[605])|(~m[600]&~m[601]&m[602]&~m[604]&m[605])|(m[600]&~m[601]&m[602]&~m[604]&m[605])|(~m[600]&m[601]&m[602]&~m[604]&m[605])|(m[600]&m[601]&m[602]&~m[604]&m[605])|(m[600]&m[601]&m[602]&m[604]&m[605]));
    m[608] = (((m[605]&~m[606]&~m[607]&~m[609]&~m[610])|(~m[605]&m[606]&~m[607]&~m[609]&~m[610])|(~m[605]&~m[606]&m[607]&~m[609]&~m[610])|(m[605]&m[606]&m[607]&m[609]&~m[610])|(~m[605]&~m[606]&~m[607]&~m[609]&m[610])|(m[605]&m[606]&~m[607]&m[609]&m[610])|(m[605]&~m[606]&m[607]&m[609]&m[610])|(~m[605]&m[606]&m[607]&m[609]&m[610]))&UnbiasedRNG[320])|((m[605]&m[606]&~m[607]&~m[609]&~m[610])|(m[605]&~m[606]&m[607]&~m[609]&~m[610])|(~m[605]&m[606]&m[607]&~m[609]&~m[610])|(m[605]&m[606]&m[607]&~m[609]&~m[610])|(m[605]&~m[606]&~m[607]&~m[609]&m[610])|(~m[605]&m[606]&~m[607]&~m[609]&m[610])|(m[605]&m[606]&~m[607]&~m[609]&m[610])|(~m[605]&~m[606]&m[607]&~m[609]&m[610])|(m[605]&~m[606]&m[607]&~m[609]&m[610])|(~m[605]&m[606]&m[607]&~m[609]&m[610])|(m[605]&m[606]&m[607]&~m[609]&m[610])|(m[605]&m[606]&m[607]&m[609]&m[610]));
    m[613] = (((m[610]&~m[611]&~m[612]&~m[614]&~m[615])|(~m[610]&m[611]&~m[612]&~m[614]&~m[615])|(~m[610]&~m[611]&m[612]&~m[614]&~m[615])|(m[610]&m[611]&m[612]&m[614]&~m[615])|(~m[610]&~m[611]&~m[612]&~m[614]&m[615])|(m[610]&m[611]&~m[612]&m[614]&m[615])|(m[610]&~m[611]&m[612]&m[614]&m[615])|(~m[610]&m[611]&m[612]&m[614]&m[615]))&UnbiasedRNG[321])|((m[610]&m[611]&~m[612]&~m[614]&~m[615])|(m[610]&~m[611]&m[612]&~m[614]&~m[615])|(~m[610]&m[611]&m[612]&~m[614]&~m[615])|(m[610]&m[611]&m[612]&~m[614]&~m[615])|(m[610]&~m[611]&~m[612]&~m[614]&m[615])|(~m[610]&m[611]&~m[612]&~m[614]&m[615])|(m[610]&m[611]&~m[612]&~m[614]&m[615])|(~m[610]&~m[611]&m[612]&~m[614]&m[615])|(m[610]&~m[611]&m[612]&~m[614]&m[615])|(~m[610]&m[611]&m[612]&~m[614]&m[615])|(m[610]&m[611]&m[612]&~m[614]&m[615])|(m[610]&m[611]&m[612]&m[614]&m[615]));
    m[618] = (((m[615]&~m[616]&~m[617]&~m[619]&~m[620])|(~m[615]&m[616]&~m[617]&~m[619]&~m[620])|(~m[615]&~m[616]&m[617]&~m[619]&~m[620])|(m[615]&m[616]&m[617]&m[619]&~m[620])|(~m[615]&~m[616]&~m[617]&~m[619]&m[620])|(m[615]&m[616]&~m[617]&m[619]&m[620])|(m[615]&~m[616]&m[617]&m[619]&m[620])|(~m[615]&m[616]&m[617]&m[619]&m[620]))&UnbiasedRNG[322])|((m[615]&m[616]&~m[617]&~m[619]&~m[620])|(m[615]&~m[616]&m[617]&~m[619]&~m[620])|(~m[615]&m[616]&m[617]&~m[619]&~m[620])|(m[615]&m[616]&m[617]&~m[619]&~m[620])|(m[615]&~m[616]&~m[617]&~m[619]&m[620])|(~m[615]&m[616]&~m[617]&~m[619]&m[620])|(m[615]&m[616]&~m[617]&~m[619]&m[620])|(~m[615]&~m[616]&m[617]&~m[619]&m[620])|(m[615]&~m[616]&m[617]&~m[619]&m[620])|(~m[615]&m[616]&m[617]&~m[619]&m[620])|(m[615]&m[616]&m[617]&~m[619]&m[620])|(m[615]&m[616]&m[617]&m[619]&m[620]));
    m[623] = (((m[620]&~m[621]&~m[622]&~m[624]&~m[625])|(~m[620]&m[621]&~m[622]&~m[624]&~m[625])|(~m[620]&~m[621]&m[622]&~m[624]&~m[625])|(m[620]&m[621]&m[622]&m[624]&~m[625])|(~m[620]&~m[621]&~m[622]&~m[624]&m[625])|(m[620]&m[621]&~m[622]&m[624]&m[625])|(m[620]&~m[621]&m[622]&m[624]&m[625])|(~m[620]&m[621]&m[622]&m[624]&m[625]))&UnbiasedRNG[323])|((m[620]&m[621]&~m[622]&~m[624]&~m[625])|(m[620]&~m[621]&m[622]&~m[624]&~m[625])|(~m[620]&m[621]&m[622]&~m[624]&~m[625])|(m[620]&m[621]&m[622]&~m[624]&~m[625])|(m[620]&~m[621]&~m[622]&~m[624]&m[625])|(~m[620]&m[621]&~m[622]&~m[624]&m[625])|(m[620]&m[621]&~m[622]&~m[624]&m[625])|(~m[620]&~m[621]&m[622]&~m[624]&m[625])|(m[620]&~m[621]&m[622]&~m[624]&m[625])|(~m[620]&m[621]&m[622]&~m[624]&m[625])|(m[620]&m[621]&m[622]&~m[624]&m[625])|(m[620]&m[621]&m[622]&m[624]&m[625]));
    m[633] = (((m[630]&~m[631]&~m[632]&~m[634]&~m[635])|(~m[630]&m[631]&~m[632]&~m[634]&~m[635])|(~m[630]&~m[631]&m[632]&~m[634]&~m[635])|(m[630]&m[631]&m[632]&m[634]&~m[635])|(~m[630]&~m[631]&~m[632]&~m[634]&m[635])|(m[630]&m[631]&~m[632]&m[634]&m[635])|(m[630]&~m[631]&m[632]&m[634]&m[635])|(~m[630]&m[631]&m[632]&m[634]&m[635]))&UnbiasedRNG[324])|((m[630]&m[631]&~m[632]&~m[634]&~m[635])|(m[630]&~m[631]&m[632]&~m[634]&~m[635])|(~m[630]&m[631]&m[632]&~m[634]&~m[635])|(m[630]&m[631]&m[632]&~m[634]&~m[635])|(m[630]&~m[631]&~m[632]&~m[634]&m[635])|(~m[630]&m[631]&~m[632]&~m[634]&m[635])|(m[630]&m[631]&~m[632]&~m[634]&m[635])|(~m[630]&~m[631]&m[632]&~m[634]&m[635])|(m[630]&~m[631]&m[632]&~m[634]&m[635])|(~m[630]&m[631]&m[632]&~m[634]&m[635])|(m[630]&m[631]&m[632]&~m[634]&m[635])|(m[630]&m[631]&m[632]&m[634]&m[635]));
    m[638] = (((m[635]&~m[636]&~m[637]&~m[639]&~m[640])|(~m[635]&m[636]&~m[637]&~m[639]&~m[640])|(~m[635]&~m[636]&m[637]&~m[639]&~m[640])|(m[635]&m[636]&m[637]&m[639]&~m[640])|(~m[635]&~m[636]&~m[637]&~m[639]&m[640])|(m[635]&m[636]&~m[637]&m[639]&m[640])|(m[635]&~m[636]&m[637]&m[639]&m[640])|(~m[635]&m[636]&m[637]&m[639]&m[640]))&UnbiasedRNG[325])|((m[635]&m[636]&~m[637]&~m[639]&~m[640])|(m[635]&~m[636]&m[637]&~m[639]&~m[640])|(~m[635]&m[636]&m[637]&~m[639]&~m[640])|(m[635]&m[636]&m[637]&~m[639]&~m[640])|(m[635]&~m[636]&~m[637]&~m[639]&m[640])|(~m[635]&m[636]&~m[637]&~m[639]&m[640])|(m[635]&m[636]&~m[637]&~m[639]&m[640])|(~m[635]&~m[636]&m[637]&~m[639]&m[640])|(m[635]&~m[636]&m[637]&~m[639]&m[640])|(~m[635]&m[636]&m[637]&~m[639]&m[640])|(m[635]&m[636]&m[637]&~m[639]&m[640])|(m[635]&m[636]&m[637]&m[639]&m[640]));
    m[643] = (((m[640]&~m[641]&~m[642]&~m[644]&~m[645])|(~m[640]&m[641]&~m[642]&~m[644]&~m[645])|(~m[640]&~m[641]&m[642]&~m[644]&~m[645])|(m[640]&m[641]&m[642]&m[644]&~m[645])|(~m[640]&~m[641]&~m[642]&~m[644]&m[645])|(m[640]&m[641]&~m[642]&m[644]&m[645])|(m[640]&~m[641]&m[642]&m[644]&m[645])|(~m[640]&m[641]&m[642]&m[644]&m[645]))&UnbiasedRNG[326])|((m[640]&m[641]&~m[642]&~m[644]&~m[645])|(m[640]&~m[641]&m[642]&~m[644]&~m[645])|(~m[640]&m[641]&m[642]&~m[644]&~m[645])|(m[640]&m[641]&m[642]&~m[644]&~m[645])|(m[640]&~m[641]&~m[642]&~m[644]&m[645])|(~m[640]&m[641]&~m[642]&~m[644]&m[645])|(m[640]&m[641]&~m[642]&~m[644]&m[645])|(~m[640]&~m[641]&m[642]&~m[644]&m[645])|(m[640]&~m[641]&m[642]&~m[644]&m[645])|(~m[640]&m[641]&m[642]&~m[644]&m[645])|(m[640]&m[641]&m[642]&~m[644]&m[645])|(m[640]&m[641]&m[642]&m[644]&m[645]));
    m[648] = (((m[645]&~m[646]&~m[647]&~m[649]&~m[650])|(~m[645]&m[646]&~m[647]&~m[649]&~m[650])|(~m[645]&~m[646]&m[647]&~m[649]&~m[650])|(m[645]&m[646]&m[647]&m[649]&~m[650])|(~m[645]&~m[646]&~m[647]&~m[649]&m[650])|(m[645]&m[646]&~m[647]&m[649]&m[650])|(m[645]&~m[646]&m[647]&m[649]&m[650])|(~m[645]&m[646]&m[647]&m[649]&m[650]))&UnbiasedRNG[327])|((m[645]&m[646]&~m[647]&~m[649]&~m[650])|(m[645]&~m[646]&m[647]&~m[649]&~m[650])|(~m[645]&m[646]&m[647]&~m[649]&~m[650])|(m[645]&m[646]&m[647]&~m[649]&~m[650])|(m[645]&~m[646]&~m[647]&~m[649]&m[650])|(~m[645]&m[646]&~m[647]&~m[649]&m[650])|(m[645]&m[646]&~m[647]&~m[649]&m[650])|(~m[645]&~m[646]&m[647]&~m[649]&m[650])|(m[645]&~m[646]&m[647]&~m[649]&m[650])|(~m[645]&m[646]&m[647]&~m[649]&m[650])|(m[645]&m[646]&m[647]&~m[649]&m[650])|(m[645]&m[646]&m[647]&m[649]&m[650]));
    m[653] = (((m[650]&~m[651]&~m[652]&~m[654]&~m[655])|(~m[650]&m[651]&~m[652]&~m[654]&~m[655])|(~m[650]&~m[651]&m[652]&~m[654]&~m[655])|(m[650]&m[651]&m[652]&m[654]&~m[655])|(~m[650]&~m[651]&~m[652]&~m[654]&m[655])|(m[650]&m[651]&~m[652]&m[654]&m[655])|(m[650]&~m[651]&m[652]&m[654]&m[655])|(~m[650]&m[651]&m[652]&m[654]&m[655]))&UnbiasedRNG[328])|((m[650]&m[651]&~m[652]&~m[654]&~m[655])|(m[650]&~m[651]&m[652]&~m[654]&~m[655])|(~m[650]&m[651]&m[652]&~m[654]&~m[655])|(m[650]&m[651]&m[652]&~m[654]&~m[655])|(m[650]&~m[651]&~m[652]&~m[654]&m[655])|(~m[650]&m[651]&~m[652]&~m[654]&m[655])|(m[650]&m[651]&~m[652]&~m[654]&m[655])|(~m[650]&~m[651]&m[652]&~m[654]&m[655])|(m[650]&~m[651]&m[652]&~m[654]&m[655])|(~m[650]&m[651]&m[652]&~m[654]&m[655])|(m[650]&m[651]&m[652]&~m[654]&m[655])|(m[650]&m[651]&m[652]&m[654]&m[655]));
    m[658] = (((m[655]&~m[656]&~m[657]&~m[659]&~m[660])|(~m[655]&m[656]&~m[657]&~m[659]&~m[660])|(~m[655]&~m[656]&m[657]&~m[659]&~m[660])|(m[655]&m[656]&m[657]&m[659]&~m[660])|(~m[655]&~m[656]&~m[657]&~m[659]&m[660])|(m[655]&m[656]&~m[657]&m[659]&m[660])|(m[655]&~m[656]&m[657]&m[659]&m[660])|(~m[655]&m[656]&m[657]&m[659]&m[660]))&UnbiasedRNG[329])|((m[655]&m[656]&~m[657]&~m[659]&~m[660])|(m[655]&~m[656]&m[657]&~m[659]&~m[660])|(~m[655]&m[656]&m[657]&~m[659]&~m[660])|(m[655]&m[656]&m[657]&~m[659]&~m[660])|(m[655]&~m[656]&~m[657]&~m[659]&m[660])|(~m[655]&m[656]&~m[657]&~m[659]&m[660])|(m[655]&m[656]&~m[657]&~m[659]&m[660])|(~m[655]&~m[656]&m[657]&~m[659]&m[660])|(m[655]&~m[656]&m[657]&~m[659]&m[660])|(~m[655]&m[656]&m[657]&~m[659]&m[660])|(m[655]&m[656]&m[657]&~m[659]&m[660])|(m[655]&m[656]&m[657]&m[659]&m[660]));
    m[663] = (((m[660]&~m[661]&~m[662]&~m[664]&~m[665])|(~m[660]&m[661]&~m[662]&~m[664]&~m[665])|(~m[660]&~m[661]&m[662]&~m[664]&~m[665])|(m[660]&m[661]&m[662]&m[664]&~m[665])|(~m[660]&~m[661]&~m[662]&~m[664]&m[665])|(m[660]&m[661]&~m[662]&m[664]&m[665])|(m[660]&~m[661]&m[662]&m[664]&m[665])|(~m[660]&m[661]&m[662]&m[664]&m[665]))&UnbiasedRNG[330])|((m[660]&m[661]&~m[662]&~m[664]&~m[665])|(m[660]&~m[661]&m[662]&~m[664]&~m[665])|(~m[660]&m[661]&m[662]&~m[664]&~m[665])|(m[660]&m[661]&m[662]&~m[664]&~m[665])|(m[660]&~m[661]&~m[662]&~m[664]&m[665])|(~m[660]&m[661]&~m[662]&~m[664]&m[665])|(m[660]&m[661]&~m[662]&~m[664]&m[665])|(~m[660]&~m[661]&m[662]&~m[664]&m[665])|(m[660]&~m[661]&m[662]&~m[664]&m[665])|(~m[660]&m[661]&m[662]&~m[664]&m[665])|(m[660]&m[661]&m[662]&~m[664]&m[665])|(m[660]&m[661]&m[662]&m[664]&m[665]));
    m[673] = (((m[670]&~m[671]&~m[672]&~m[674]&~m[675])|(~m[670]&m[671]&~m[672]&~m[674]&~m[675])|(~m[670]&~m[671]&m[672]&~m[674]&~m[675])|(m[670]&m[671]&m[672]&m[674]&~m[675])|(~m[670]&~m[671]&~m[672]&~m[674]&m[675])|(m[670]&m[671]&~m[672]&m[674]&m[675])|(m[670]&~m[671]&m[672]&m[674]&m[675])|(~m[670]&m[671]&m[672]&m[674]&m[675]))&UnbiasedRNG[331])|((m[670]&m[671]&~m[672]&~m[674]&~m[675])|(m[670]&~m[671]&m[672]&~m[674]&~m[675])|(~m[670]&m[671]&m[672]&~m[674]&~m[675])|(m[670]&m[671]&m[672]&~m[674]&~m[675])|(m[670]&~m[671]&~m[672]&~m[674]&m[675])|(~m[670]&m[671]&~m[672]&~m[674]&m[675])|(m[670]&m[671]&~m[672]&~m[674]&m[675])|(~m[670]&~m[671]&m[672]&~m[674]&m[675])|(m[670]&~m[671]&m[672]&~m[674]&m[675])|(~m[670]&m[671]&m[672]&~m[674]&m[675])|(m[670]&m[671]&m[672]&~m[674]&m[675])|(m[670]&m[671]&m[672]&m[674]&m[675]));
    m[678] = (((m[675]&~m[676]&~m[677]&~m[679]&~m[680])|(~m[675]&m[676]&~m[677]&~m[679]&~m[680])|(~m[675]&~m[676]&m[677]&~m[679]&~m[680])|(m[675]&m[676]&m[677]&m[679]&~m[680])|(~m[675]&~m[676]&~m[677]&~m[679]&m[680])|(m[675]&m[676]&~m[677]&m[679]&m[680])|(m[675]&~m[676]&m[677]&m[679]&m[680])|(~m[675]&m[676]&m[677]&m[679]&m[680]))&UnbiasedRNG[332])|((m[675]&m[676]&~m[677]&~m[679]&~m[680])|(m[675]&~m[676]&m[677]&~m[679]&~m[680])|(~m[675]&m[676]&m[677]&~m[679]&~m[680])|(m[675]&m[676]&m[677]&~m[679]&~m[680])|(m[675]&~m[676]&~m[677]&~m[679]&m[680])|(~m[675]&m[676]&~m[677]&~m[679]&m[680])|(m[675]&m[676]&~m[677]&~m[679]&m[680])|(~m[675]&~m[676]&m[677]&~m[679]&m[680])|(m[675]&~m[676]&m[677]&~m[679]&m[680])|(~m[675]&m[676]&m[677]&~m[679]&m[680])|(m[675]&m[676]&m[677]&~m[679]&m[680])|(m[675]&m[676]&m[677]&m[679]&m[680]));
    m[683] = (((m[680]&~m[681]&~m[682]&~m[684]&~m[685])|(~m[680]&m[681]&~m[682]&~m[684]&~m[685])|(~m[680]&~m[681]&m[682]&~m[684]&~m[685])|(m[680]&m[681]&m[682]&m[684]&~m[685])|(~m[680]&~m[681]&~m[682]&~m[684]&m[685])|(m[680]&m[681]&~m[682]&m[684]&m[685])|(m[680]&~m[681]&m[682]&m[684]&m[685])|(~m[680]&m[681]&m[682]&m[684]&m[685]))&UnbiasedRNG[333])|((m[680]&m[681]&~m[682]&~m[684]&~m[685])|(m[680]&~m[681]&m[682]&~m[684]&~m[685])|(~m[680]&m[681]&m[682]&~m[684]&~m[685])|(m[680]&m[681]&m[682]&~m[684]&~m[685])|(m[680]&~m[681]&~m[682]&~m[684]&m[685])|(~m[680]&m[681]&~m[682]&~m[684]&m[685])|(m[680]&m[681]&~m[682]&~m[684]&m[685])|(~m[680]&~m[681]&m[682]&~m[684]&m[685])|(m[680]&~m[681]&m[682]&~m[684]&m[685])|(~m[680]&m[681]&m[682]&~m[684]&m[685])|(m[680]&m[681]&m[682]&~m[684]&m[685])|(m[680]&m[681]&m[682]&m[684]&m[685]));
    m[688] = (((m[685]&~m[686]&~m[687]&~m[689]&~m[690])|(~m[685]&m[686]&~m[687]&~m[689]&~m[690])|(~m[685]&~m[686]&m[687]&~m[689]&~m[690])|(m[685]&m[686]&m[687]&m[689]&~m[690])|(~m[685]&~m[686]&~m[687]&~m[689]&m[690])|(m[685]&m[686]&~m[687]&m[689]&m[690])|(m[685]&~m[686]&m[687]&m[689]&m[690])|(~m[685]&m[686]&m[687]&m[689]&m[690]))&UnbiasedRNG[334])|((m[685]&m[686]&~m[687]&~m[689]&~m[690])|(m[685]&~m[686]&m[687]&~m[689]&~m[690])|(~m[685]&m[686]&m[687]&~m[689]&~m[690])|(m[685]&m[686]&m[687]&~m[689]&~m[690])|(m[685]&~m[686]&~m[687]&~m[689]&m[690])|(~m[685]&m[686]&~m[687]&~m[689]&m[690])|(m[685]&m[686]&~m[687]&~m[689]&m[690])|(~m[685]&~m[686]&m[687]&~m[689]&m[690])|(m[685]&~m[686]&m[687]&~m[689]&m[690])|(~m[685]&m[686]&m[687]&~m[689]&m[690])|(m[685]&m[686]&m[687]&~m[689]&m[690])|(m[685]&m[686]&m[687]&m[689]&m[690]));
    m[693] = (((m[690]&~m[691]&~m[692]&~m[694]&~m[695])|(~m[690]&m[691]&~m[692]&~m[694]&~m[695])|(~m[690]&~m[691]&m[692]&~m[694]&~m[695])|(m[690]&m[691]&m[692]&m[694]&~m[695])|(~m[690]&~m[691]&~m[692]&~m[694]&m[695])|(m[690]&m[691]&~m[692]&m[694]&m[695])|(m[690]&~m[691]&m[692]&m[694]&m[695])|(~m[690]&m[691]&m[692]&m[694]&m[695]))&UnbiasedRNG[335])|((m[690]&m[691]&~m[692]&~m[694]&~m[695])|(m[690]&~m[691]&m[692]&~m[694]&~m[695])|(~m[690]&m[691]&m[692]&~m[694]&~m[695])|(m[690]&m[691]&m[692]&~m[694]&~m[695])|(m[690]&~m[691]&~m[692]&~m[694]&m[695])|(~m[690]&m[691]&~m[692]&~m[694]&m[695])|(m[690]&m[691]&~m[692]&~m[694]&m[695])|(~m[690]&~m[691]&m[692]&~m[694]&m[695])|(m[690]&~m[691]&m[692]&~m[694]&m[695])|(~m[690]&m[691]&m[692]&~m[694]&m[695])|(m[690]&m[691]&m[692]&~m[694]&m[695])|(m[690]&m[691]&m[692]&m[694]&m[695]));
    m[698] = (((m[695]&~m[696]&~m[697]&~m[699]&~m[700])|(~m[695]&m[696]&~m[697]&~m[699]&~m[700])|(~m[695]&~m[696]&m[697]&~m[699]&~m[700])|(m[695]&m[696]&m[697]&m[699]&~m[700])|(~m[695]&~m[696]&~m[697]&~m[699]&m[700])|(m[695]&m[696]&~m[697]&m[699]&m[700])|(m[695]&~m[696]&m[697]&m[699]&m[700])|(~m[695]&m[696]&m[697]&m[699]&m[700]))&UnbiasedRNG[336])|((m[695]&m[696]&~m[697]&~m[699]&~m[700])|(m[695]&~m[696]&m[697]&~m[699]&~m[700])|(~m[695]&m[696]&m[697]&~m[699]&~m[700])|(m[695]&m[696]&m[697]&~m[699]&~m[700])|(m[695]&~m[696]&~m[697]&~m[699]&m[700])|(~m[695]&m[696]&~m[697]&~m[699]&m[700])|(m[695]&m[696]&~m[697]&~m[699]&m[700])|(~m[695]&~m[696]&m[697]&~m[699]&m[700])|(m[695]&~m[696]&m[697]&~m[699]&m[700])|(~m[695]&m[696]&m[697]&~m[699]&m[700])|(m[695]&m[696]&m[697]&~m[699]&m[700])|(m[695]&m[696]&m[697]&m[699]&m[700]));
    m[708] = (((m[705]&~m[706]&~m[707]&~m[709]&~m[710])|(~m[705]&m[706]&~m[707]&~m[709]&~m[710])|(~m[705]&~m[706]&m[707]&~m[709]&~m[710])|(m[705]&m[706]&m[707]&m[709]&~m[710])|(~m[705]&~m[706]&~m[707]&~m[709]&m[710])|(m[705]&m[706]&~m[707]&m[709]&m[710])|(m[705]&~m[706]&m[707]&m[709]&m[710])|(~m[705]&m[706]&m[707]&m[709]&m[710]))&UnbiasedRNG[337])|((m[705]&m[706]&~m[707]&~m[709]&~m[710])|(m[705]&~m[706]&m[707]&~m[709]&~m[710])|(~m[705]&m[706]&m[707]&~m[709]&~m[710])|(m[705]&m[706]&m[707]&~m[709]&~m[710])|(m[705]&~m[706]&~m[707]&~m[709]&m[710])|(~m[705]&m[706]&~m[707]&~m[709]&m[710])|(m[705]&m[706]&~m[707]&~m[709]&m[710])|(~m[705]&~m[706]&m[707]&~m[709]&m[710])|(m[705]&~m[706]&m[707]&~m[709]&m[710])|(~m[705]&m[706]&m[707]&~m[709]&m[710])|(m[705]&m[706]&m[707]&~m[709]&m[710])|(m[705]&m[706]&m[707]&m[709]&m[710]));
    m[713] = (((m[710]&~m[711]&~m[712]&~m[714]&~m[715])|(~m[710]&m[711]&~m[712]&~m[714]&~m[715])|(~m[710]&~m[711]&m[712]&~m[714]&~m[715])|(m[710]&m[711]&m[712]&m[714]&~m[715])|(~m[710]&~m[711]&~m[712]&~m[714]&m[715])|(m[710]&m[711]&~m[712]&m[714]&m[715])|(m[710]&~m[711]&m[712]&m[714]&m[715])|(~m[710]&m[711]&m[712]&m[714]&m[715]))&UnbiasedRNG[338])|((m[710]&m[711]&~m[712]&~m[714]&~m[715])|(m[710]&~m[711]&m[712]&~m[714]&~m[715])|(~m[710]&m[711]&m[712]&~m[714]&~m[715])|(m[710]&m[711]&m[712]&~m[714]&~m[715])|(m[710]&~m[711]&~m[712]&~m[714]&m[715])|(~m[710]&m[711]&~m[712]&~m[714]&m[715])|(m[710]&m[711]&~m[712]&~m[714]&m[715])|(~m[710]&~m[711]&m[712]&~m[714]&m[715])|(m[710]&~m[711]&m[712]&~m[714]&m[715])|(~m[710]&m[711]&m[712]&~m[714]&m[715])|(m[710]&m[711]&m[712]&~m[714]&m[715])|(m[710]&m[711]&m[712]&m[714]&m[715]));
    m[718] = (((m[715]&~m[716]&~m[717]&~m[719]&~m[720])|(~m[715]&m[716]&~m[717]&~m[719]&~m[720])|(~m[715]&~m[716]&m[717]&~m[719]&~m[720])|(m[715]&m[716]&m[717]&m[719]&~m[720])|(~m[715]&~m[716]&~m[717]&~m[719]&m[720])|(m[715]&m[716]&~m[717]&m[719]&m[720])|(m[715]&~m[716]&m[717]&m[719]&m[720])|(~m[715]&m[716]&m[717]&m[719]&m[720]))&UnbiasedRNG[339])|((m[715]&m[716]&~m[717]&~m[719]&~m[720])|(m[715]&~m[716]&m[717]&~m[719]&~m[720])|(~m[715]&m[716]&m[717]&~m[719]&~m[720])|(m[715]&m[716]&m[717]&~m[719]&~m[720])|(m[715]&~m[716]&~m[717]&~m[719]&m[720])|(~m[715]&m[716]&~m[717]&~m[719]&m[720])|(m[715]&m[716]&~m[717]&~m[719]&m[720])|(~m[715]&~m[716]&m[717]&~m[719]&m[720])|(m[715]&~m[716]&m[717]&~m[719]&m[720])|(~m[715]&m[716]&m[717]&~m[719]&m[720])|(m[715]&m[716]&m[717]&~m[719]&m[720])|(m[715]&m[716]&m[717]&m[719]&m[720]));
    m[723] = (((m[720]&~m[721]&~m[722]&~m[724]&~m[725])|(~m[720]&m[721]&~m[722]&~m[724]&~m[725])|(~m[720]&~m[721]&m[722]&~m[724]&~m[725])|(m[720]&m[721]&m[722]&m[724]&~m[725])|(~m[720]&~m[721]&~m[722]&~m[724]&m[725])|(m[720]&m[721]&~m[722]&m[724]&m[725])|(m[720]&~m[721]&m[722]&m[724]&m[725])|(~m[720]&m[721]&m[722]&m[724]&m[725]))&UnbiasedRNG[340])|((m[720]&m[721]&~m[722]&~m[724]&~m[725])|(m[720]&~m[721]&m[722]&~m[724]&~m[725])|(~m[720]&m[721]&m[722]&~m[724]&~m[725])|(m[720]&m[721]&m[722]&~m[724]&~m[725])|(m[720]&~m[721]&~m[722]&~m[724]&m[725])|(~m[720]&m[721]&~m[722]&~m[724]&m[725])|(m[720]&m[721]&~m[722]&~m[724]&m[725])|(~m[720]&~m[721]&m[722]&~m[724]&m[725])|(m[720]&~m[721]&m[722]&~m[724]&m[725])|(~m[720]&m[721]&m[722]&~m[724]&m[725])|(m[720]&m[721]&m[722]&~m[724]&m[725])|(m[720]&m[721]&m[722]&m[724]&m[725]));
    m[728] = (((m[725]&~m[726]&~m[727]&~m[729]&~m[730])|(~m[725]&m[726]&~m[727]&~m[729]&~m[730])|(~m[725]&~m[726]&m[727]&~m[729]&~m[730])|(m[725]&m[726]&m[727]&m[729]&~m[730])|(~m[725]&~m[726]&~m[727]&~m[729]&m[730])|(m[725]&m[726]&~m[727]&m[729]&m[730])|(m[725]&~m[726]&m[727]&m[729]&m[730])|(~m[725]&m[726]&m[727]&m[729]&m[730]))&UnbiasedRNG[341])|((m[725]&m[726]&~m[727]&~m[729]&~m[730])|(m[725]&~m[726]&m[727]&~m[729]&~m[730])|(~m[725]&m[726]&m[727]&~m[729]&~m[730])|(m[725]&m[726]&m[727]&~m[729]&~m[730])|(m[725]&~m[726]&~m[727]&~m[729]&m[730])|(~m[725]&m[726]&~m[727]&~m[729]&m[730])|(m[725]&m[726]&~m[727]&~m[729]&m[730])|(~m[725]&~m[726]&m[727]&~m[729]&m[730])|(m[725]&~m[726]&m[727]&~m[729]&m[730])|(~m[725]&m[726]&m[727]&~m[729]&m[730])|(m[725]&m[726]&m[727]&~m[729]&m[730])|(m[725]&m[726]&m[727]&m[729]&m[730]));
    m[738] = (((m[735]&~m[736]&~m[737]&~m[739]&~m[740])|(~m[735]&m[736]&~m[737]&~m[739]&~m[740])|(~m[735]&~m[736]&m[737]&~m[739]&~m[740])|(m[735]&m[736]&m[737]&m[739]&~m[740])|(~m[735]&~m[736]&~m[737]&~m[739]&m[740])|(m[735]&m[736]&~m[737]&m[739]&m[740])|(m[735]&~m[736]&m[737]&m[739]&m[740])|(~m[735]&m[736]&m[737]&m[739]&m[740]))&UnbiasedRNG[342])|((m[735]&m[736]&~m[737]&~m[739]&~m[740])|(m[735]&~m[736]&m[737]&~m[739]&~m[740])|(~m[735]&m[736]&m[737]&~m[739]&~m[740])|(m[735]&m[736]&m[737]&~m[739]&~m[740])|(m[735]&~m[736]&~m[737]&~m[739]&m[740])|(~m[735]&m[736]&~m[737]&~m[739]&m[740])|(m[735]&m[736]&~m[737]&~m[739]&m[740])|(~m[735]&~m[736]&m[737]&~m[739]&m[740])|(m[735]&~m[736]&m[737]&~m[739]&m[740])|(~m[735]&m[736]&m[737]&~m[739]&m[740])|(m[735]&m[736]&m[737]&~m[739]&m[740])|(m[735]&m[736]&m[737]&m[739]&m[740]));
    m[743] = (((m[740]&~m[741]&~m[742]&~m[744]&~m[745])|(~m[740]&m[741]&~m[742]&~m[744]&~m[745])|(~m[740]&~m[741]&m[742]&~m[744]&~m[745])|(m[740]&m[741]&m[742]&m[744]&~m[745])|(~m[740]&~m[741]&~m[742]&~m[744]&m[745])|(m[740]&m[741]&~m[742]&m[744]&m[745])|(m[740]&~m[741]&m[742]&m[744]&m[745])|(~m[740]&m[741]&m[742]&m[744]&m[745]))&UnbiasedRNG[343])|((m[740]&m[741]&~m[742]&~m[744]&~m[745])|(m[740]&~m[741]&m[742]&~m[744]&~m[745])|(~m[740]&m[741]&m[742]&~m[744]&~m[745])|(m[740]&m[741]&m[742]&~m[744]&~m[745])|(m[740]&~m[741]&~m[742]&~m[744]&m[745])|(~m[740]&m[741]&~m[742]&~m[744]&m[745])|(m[740]&m[741]&~m[742]&~m[744]&m[745])|(~m[740]&~m[741]&m[742]&~m[744]&m[745])|(m[740]&~m[741]&m[742]&~m[744]&m[745])|(~m[740]&m[741]&m[742]&~m[744]&m[745])|(m[740]&m[741]&m[742]&~m[744]&m[745])|(m[740]&m[741]&m[742]&m[744]&m[745]));
    m[748] = (((m[745]&~m[746]&~m[747]&~m[749]&~m[750])|(~m[745]&m[746]&~m[747]&~m[749]&~m[750])|(~m[745]&~m[746]&m[747]&~m[749]&~m[750])|(m[745]&m[746]&m[747]&m[749]&~m[750])|(~m[745]&~m[746]&~m[747]&~m[749]&m[750])|(m[745]&m[746]&~m[747]&m[749]&m[750])|(m[745]&~m[746]&m[747]&m[749]&m[750])|(~m[745]&m[746]&m[747]&m[749]&m[750]))&UnbiasedRNG[344])|((m[745]&m[746]&~m[747]&~m[749]&~m[750])|(m[745]&~m[746]&m[747]&~m[749]&~m[750])|(~m[745]&m[746]&m[747]&~m[749]&~m[750])|(m[745]&m[746]&m[747]&~m[749]&~m[750])|(m[745]&~m[746]&~m[747]&~m[749]&m[750])|(~m[745]&m[746]&~m[747]&~m[749]&m[750])|(m[745]&m[746]&~m[747]&~m[749]&m[750])|(~m[745]&~m[746]&m[747]&~m[749]&m[750])|(m[745]&~m[746]&m[747]&~m[749]&m[750])|(~m[745]&m[746]&m[747]&~m[749]&m[750])|(m[745]&m[746]&m[747]&~m[749]&m[750])|(m[745]&m[746]&m[747]&m[749]&m[750]));
    m[753] = (((m[750]&~m[751]&~m[752]&~m[754]&~m[755])|(~m[750]&m[751]&~m[752]&~m[754]&~m[755])|(~m[750]&~m[751]&m[752]&~m[754]&~m[755])|(m[750]&m[751]&m[752]&m[754]&~m[755])|(~m[750]&~m[751]&~m[752]&~m[754]&m[755])|(m[750]&m[751]&~m[752]&m[754]&m[755])|(m[750]&~m[751]&m[752]&m[754]&m[755])|(~m[750]&m[751]&m[752]&m[754]&m[755]))&UnbiasedRNG[345])|((m[750]&m[751]&~m[752]&~m[754]&~m[755])|(m[750]&~m[751]&m[752]&~m[754]&~m[755])|(~m[750]&m[751]&m[752]&~m[754]&~m[755])|(m[750]&m[751]&m[752]&~m[754]&~m[755])|(m[750]&~m[751]&~m[752]&~m[754]&m[755])|(~m[750]&m[751]&~m[752]&~m[754]&m[755])|(m[750]&m[751]&~m[752]&~m[754]&m[755])|(~m[750]&~m[751]&m[752]&~m[754]&m[755])|(m[750]&~m[751]&m[752]&~m[754]&m[755])|(~m[750]&m[751]&m[752]&~m[754]&m[755])|(m[750]&m[751]&m[752]&~m[754]&m[755])|(m[750]&m[751]&m[752]&m[754]&m[755]));
    m[763] = (((m[760]&~m[761]&~m[762]&~m[764]&~m[765])|(~m[760]&m[761]&~m[762]&~m[764]&~m[765])|(~m[760]&~m[761]&m[762]&~m[764]&~m[765])|(m[760]&m[761]&m[762]&m[764]&~m[765])|(~m[760]&~m[761]&~m[762]&~m[764]&m[765])|(m[760]&m[761]&~m[762]&m[764]&m[765])|(m[760]&~m[761]&m[762]&m[764]&m[765])|(~m[760]&m[761]&m[762]&m[764]&m[765]))&UnbiasedRNG[346])|((m[760]&m[761]&~m[762]&~m[764]&~m[765])|(m[760]&~m[761]&m[762]&~m[764]&~m[765])|(~m[760]&m[761]&m[762]&~m[764]&~m[765])|(m[760]&m[761]&m[762]&~m[764]&~m[765])|(m[760]&~m[761]&~m[762]&~m[764]&m[765])|(~m[760]&m[761]&~m[762]&~m[764]&m[765])|(m[760]&m[761]&~m[762]&~m[764]&m[765])|(~m[760]&~m[761]&m[762]&~m[764]&m[765])|(m[760]&~m[761]&m[762]&~m[764]&m[765])|(~m[760]&m[761]&m[762]&~m[764]&m[765])|(m[760]&m[761]&m[762]&~m[764]&m[765])|(m[760]&m[761]&m[762]&m[764]&m[765]));
    m[768] = (((m[765]&~m[766]&~m[767]&~m[769]&~m[770])|(~m[765]&m[766]&~m[767]&~m[769]&~m[770])|(~m[765]&~m[766]&m[767]&~m[769]&~m[770])|(m[765]&m[766]&m[767]&m[769]&~m[770])|(~m[765]&~m[766]&~m[767]&~m[769]&m[770])|(m[765]&m[766]&~m[767]&m[769]&m[770])|(m[765]&~m[766]&m[767]&m[769]&m[770])|(~m[765]&m[766]&m[767]&m[769]&m[770]))&UnbiasedRNG[347])|((m[765]&m[766]&~m[767]&~m[769]&~m[770])|(m[765]&~m[766]&m[767]&~m[769]&~m[770])|(~m[765]&m[766]&m[767]&~m[769]&~m[770])|(m[765]&m[766]&m[767]&~m[769]&~m[770])|(m[765]&~m[766]&~m[767]&~m[769]&m[770])|(~m[765]&m[766]&~m[767]&~m[769]&m[770])|(m[765]&m[766]&~m[767]&~m[769]&m[770])|(~m[765]&~m[766]&m[767]&~m[769]&m[770])|(m[765]&~m[766]&m[767]&~m[769]&m[770])|(~m[765]&m[766]&m[767]&~m[769]&m[770])|(m[765]&m[766]&m[767]&~m[769]&m[770])|(m[765]&m[766]&m[767]&m[769]&m[770]));
    m[773] = (((m[770]&~m[771]&~m[772]&~m[774]&~m[775])|(~m[770]&m[771]&~m[772]&~m[774]&~m[775])|(~m[770]&~m[771]&m[772]&~m[774]&~m[775])|(m[770]&m[771]&m[772]&m[774]&~m[775])|(~m[770]&~m[771]&~m[772]&~m[774]&m[775])|(m[770]&m[771]&~m[772]&m[774]&m[775])|(m[770]&~m[771]&m[772]&m[774]&m[775])|(~m[770]&m[771]&m[772]&m[774]&m[775]))&UnbiasedRNG[348])|((m[770]&m[771]&~m[772]&~m[774]&~m[775])|(m[770]&~m[771]&m[772]&~m[774]&~m[775])|(~m[770]&m[771]&m[772]&~m[774]&~m[775])|(m[770]&m[771]&m[772]&~m[774]&~m[775])|(m[770]&~m[771]&~m[772]&~m[774]&m[775])|(~m[770]&m[771]&~m[772]&~m[774]&m[775])|(m[770]&m[771]&~m[772]&~m[774]&m[775])|(~m[770]&~m[771]&m[772]&~m[774]&m[775])|(m[770]&~m[771]&m[772]&~m[774]&m[775])|(~m[770]&m[771]&m[772]&~m[774]&m[775])|(m[770]&m[771]&m[772]&~m[774]&m[775])|(m[770]&m[771]&m[772]&m[774]&m[775]));
    m[783] = (((m[780]&~m[781]&~m[782]&~m[784]&~m[785])|(~m[780]&m[781]&~m[782]&~m[784]&~m[785])|(~m[780]&~m[781]&m[782]&~m[784]&~m[785])|(m[780]&m[781]&m[782]&m[784]&~m[785])|(~m[780]&~m[781]&~m[782]&~m[784]&m[785])|(m[780]&m[781]&~m[782]&m[784]&m[785])|(m[780]&~m[781]&m[782]&m[784]&m[785])|(~m[780]&m[781]&m[782]&m[784]&m[785]))&UnbiasedRNG[349])|((m[780]&m[781]&~m[782]&~m[784]&~m[785])|(m[780]&~m[781]&m[782]&~m[784]&~m[785])|(~m[780]&m[781]&m[782]&~m[784]&~m[785])|(m[780]&m[781]&m[782]&~m[784]&~m[785])|(m[780]&~m[781]&~m[782]&~m[784]&m[785])|(~m[780]&m[781]&~m[782]&~m[784]&m[785])|(m[780]&m[781]&~m[782]&~m[784]&m[785])|(~m[780]&~m[781]&m[782]&~m[784]&m[785])|(m[780]&~m[781]&m[782]&~m[784]&m[785])|(~m[780]&m[781]&m[782]&~m[784]&m[785])|(m[780]&m[781]&m[782]&~m[784]&m[785])|(m[780]&m[781]&m[782]&m[784]&m[785]));
    m[788] = (((m[785]&~m[786]&~m[787]&~m[789]&~m[790])|(~m[785]&m[786]&~m[787]&~m[789]&~m[790])|(~m[785]&~m[786]&m[787]&~m[789]&~m[790])|(m[785]&m[786]&m[787]&m[789]&~m[790])|(~m[785]&~m[786]&~m[787]&~m[789]&m[790])|(m[785]&m[786]&~m[787]&m[789]&m[790])|(m[785]&~m[786]&m[787]&m[789]&m[790])|(~m[785]&m[786]&m[787]&m[789]&m[790]))&UnbiasedRNG[350])|((m[785]&m[786]&~m[787]&~m[789]&~m[790])|(m[785]&~m[786]&m[787]&~m[789]&~m[790])|(~m[785]&m[786]&m[787]&~m[789]&~m[790])|(m[785]&m[786]&m[787]&~m[789]&~m[790])|(m[785]&~m[786]&~m[787]&~m[789]&m[790])|(~m[785]&m[786]&~m[787]&~m[789]&m[790])|(m[785]&m[786]&~m[787]&~m[789]&m[790])|(~m[785]&~m[786]&m[787]&~m[789]&m[790])|(m[785]&~m[786]&m[787]&~m[789]&m[790])|(~m[785]&m[786]&m[787]&~m[789]&m[790])|(m[785]&m[786]&m[787]&~m[789]&m[790])|(m[785]&m[786]&m[787]&m[789]&m[790]));
    m[798] = (((m[795]&~m[796]&~m[797]&~m[799]&~m[800])|(~m[795]&m[796]&~m[797]&~m[799]&~m[800])|(~m[795]&~m[796]&m[797]&~m[799]&~m[800])|(m[795]&m[796]&m[797]&m[799]&~m[800])|(~m[795]&~m[796]&~m[797]&~m[799]&m[800])|(m[795]&m[796]&~m[797]&m[799]&m[800])|(m[795]&~m[796]&m[797]&m[799]&m[800])|(~m[795]&m[796]&m[797]&m[799]&m[800]))&UnbiasedRNG[351])|((m[795]&m[796]&~m[797]&~m[799]&~m[800])|(m[795]&~m[796]&m[797]&~m[799]&~m[800])|(~m[795]&m[796]&m[797]&~m[799]&~m[800])|(m[795]&m[796]&m[797]&~m[799]&~m[800])|(m[795]&~m[796]&~m[797]&~m[799]&m[800])|(~m[795]&m[796]&~m[797]&~m[799]&m[800])|(m[795]&m[796]&~m[797]&~m[799]&m[800])|(~m[795]&~m[796]&m[797]&~m[799]&m[800])|(m[795]&~m[796]&m[797]&~m[799]&m[800])|(~m[795]&m[796]&m[797]&~m[799]&m[800])|(m[795]&m[796]&m[797]&~m[799]&m[800])|(m[795]&m[796]&m[797]&m[799]&m[800]));
end

always @(posedge color4_clk) begin
    m[364] = (((m[360]&~m[361]&~m[362]&~m[363]&~m[367])|(~m[360]&m[361]&~m[362]&~m[363]&~m[367])|(~m[360]&~m[361]&m[362]&~m[363]&~m[367])|(m[360]&m[361]&~m[362]&m[363]&~m[367])|(m[360]&~m[361]&m[362]&m[363]&~m[367])|(~m[360]&m[361]&m[362]&m[363]&~m[367]))&BiasedRNG[339])|(((m[360]&~m[361]&~m[362]&~m[363]&m[367])|(~m[360]&m[361]&~m[362]&~m[363]&m[367])|(~m[360]&~m[361]&m[362]&~m[363]&m[367])|(m[360]&m[361]&~m[362]&m[363]&m[367])|(m[360]&~m[361]&m[362]&m[363]&m[367])|(~m[360]&m[361]&m[362]&m[363]&m[367]))&~BiasedRNG[339])|((m[360]&m[361]&~m[362]&~m[363]&~m[367])|(m[360]&~m[361]&m[362]&~m[363]&~m[367])|(~m[360]&m[361]&m[362]&~m[363]&~m[367])|(m[360]&m[361]&m[362]&~m[363]&~m[367])|(m[360]&m[361]&m[362]&m[363]&~m[367])|(m[360]&m[361]&~m[362]&~m[363]&m[367])|(m[360]&~m[361]&m[362]&~m[363]&m[367])|(~m[360]&m[361]&m[362]&~m[363]&m[367])|(m[360]&m[361]&m[362]&~m[363]&m[367])|(m[360]&m[361]&m[362]&m[363]&m[367]));
    m[369] = (((m[365]&~m[366]&~m[367]&~m[368]&~m[377])|(~m[365]&m[366]&~m[367]&~m[368]&~m[377])|(~m[365]&~m[366]&m[367]&~m[368]&~m[377])|(m[365]&m[366]&~m[367]&m[368]&~m[377])|(m[365]&~m[366]&m[367]&m[368]&~m[377])|(~m[365]&m[366]&m[367]&m[368]&~m[377]))&BiasedRNG[340])|(((m[365]&~m[366]&~m[367]&~m[368]&m[377])|(~m[365]&m[366]&~m[367]&~m[368]&m[377])|(~m[365]&~m[366]&m[367]&~m[368]&m[377])|(m[365]&m[366]&~m[367]&m[368]&m[377])|(m[365]&~m[366]&m[367]&m[368]&m[377])|(~m[365]&m[366]&m[367]&m[368]&m[377]))&~BiasedRNG[340])|((m[365]&m[366]&~m[367]&~m[368]&~m[377])|(m[365]&~m[366]&m[367]&~m[368]&~m[377])|(~m[365]&m[366]&m[367]&~m[368]&~m[377])|(m[365]&m[366]&m[367]&~m[368]&~m[377])|(m[365]&m[366]&m[367]&m[368]&~m[377])|(m[365]&m[366]&~m[367]&~m[368]&m[377])|(m[365]&~m[366]&m[367]&~m[368]&m[377])|(~m[365]&m[366]&m[367]&~m[368]&m[377])|(m[365]&m[366]&m[367]&~m[368]&m[377])|(m[365]&m[366]&m[367]&m[368]&m[377]));
    m[374] = (((m[370]&~m[371]&~m[372]&~m[373]&~m[382])|(~m[370]&m[371]&~m[372]&~m[373]&~m[382])|(~m[370]&~m[371]&m[372]&~m[373]&~m[382])|(m[370]&m[371]&~m[372]&m[373]&~m[382])|(m[370]&~m[371]&m[372]&m[373]&~m[382])|(~m[370]&m[371]&m[372]&m[373]&~m[382]))&BiasedRNG[341])|(((m[370]&~m[371]&~m[372]&~m[373]&m[382])|(~m[370]&m[371]&~m[372]&~m[373]&m[382])|(~m[370]&~m[371]&m[372]&~m[373]&m[382])|(m[370]&m[371]&~m[372]&m[373]&m[382])|(m[370]&~m[371]&m[372]&m[373]&m[382])|(~m[370]&m[371]&m[372]&m[373]&m[382]))&~BiasedRNG[341])|((m[370]&m[371]&~m[372]&~m[373]&~m[382])|(m[370]&~m[371]&m[372]&~m[373]&~m[382])|(~m[370]&m[371]&m[372]&~m[373]&~m[382])|(m[370]&m[371]&m[372]&~m[373]&~m[382])|(m[370]&m[371]&m[372]&m[373]&~m[382])|(m[370]&m[371]&~m[372]&~m[373]&m[382])|(m[370]&~m[371]&m[372]&~m[373]&m[382])|(~m[370]&m[371]&m[372]&~m[373]&m[382])|(m[370]&m[371]&m[372]&~m[373]&m[382])|(m[370]&m[371]&m[372]&m[373]&m[382]));
    m[379] = (((m[375]&~m[376]&~m[377]&~m[378]&~m[392])|(~m[375]&m[376]&~m[377]&~m[378]&~m[392])|(~m[375]&~m[376]&m[377]&~m[378]&~m[392])|(m[375]&m[376]&~m[377]&m[378]&~m[392])|(m[375]&~m[376]&m[377]&m[378]&~m[392])|(~m[375]&m[376]&m[377]&m[378]&~m[392]))&BiasedRNG[342])|(((m[375]&~m[376]&~m[377]&~m[378]&m[392])|(~m[375]&m[376]&~m[377]&~m[378]&m[392])|(~m[375]&~m[376]&m[377]&~m[378]&m[392])|(m[375]&m[376]&~m[377]&m[378]&m[392])|(m[375]&~m[376]&m[377]&m[378]&m[392])|(~m[375]&m[376]&m[377]&m[378]&m[392]))&~BiasedRNG[342])|((m[375]&m[376]&~m[377]&~m[378]&~m[392])|(m[375]&~m[376]&m[377]&~m[378]&~m[392])|(~m[375]&m[376]&m[377]&~m[378]&~m[392])|(m[375]&m[376]&m[377]&~m[378]&~m[392])|(m[375]&m[376]&m[377]&m[378]&~m[392])|(m[375]&m[376]&~m[377]&~m[378]&m[392])|(m[375]&~m[376]&m[377]&~m[378]&m[392])|(~m[375]&m[376]&m[377]&~m[378]&m[392])|(m[375]&m[376]&m[377]&~m[378]&m[392])|(m[375]&m[376]&m[377]&m[378]&m[392]));
    m[384] = (((m[380]&~m[381]&~m[382]&~m[383]&~m[397])|(~m[380]&m[381]&~m[382]&~m[383]&~m[397])|(~m[380]&~m[381]&m[382]&~m[383]&~m[397])|(m[380]&m[381]&~m[382]&m[383]&~m[397])|(m[380]&~m[381]&m[382]&m[383]&~m[397])|(~m[380]&m[381]&m[382]&m[383]&~m[397]))&BiasedRNG[343])|(((m[380]&~m[381]&~m[382]&~m[383]&m[397])|(~m[380]&m[381]&~m[382]&~m[383]&m[397])|(~m[380]&~m[381]&m[382]&~m[383]&m[397])|(m[380]&m[381]&~m[382]&m[383]&m[397])|(m[380]&~m[381]&m[382]&m[383]&m[397])|(~m[380]&m[381]&m[382]&m[383]&m[397]))&~BiasedRNG[343])|((m[380]&m[381]&~m[382]&~m[383]&~m[397])|(m[380]&~m[381]&m[382]&~m[383]&~m[397])|(~m[380]&m[381]&m[382]&~m[383]&~m[397])|(m[380]&m[381]&m[382]&~m[383]&~m[397])|(m[380]&m[381]&m[382]&m[383]&~m[397])|(m[380]&m[381]&~m[382]&~m[383]&m[397])|(m[380]&~m[381]&m[382]&~m[383]&m[397])|(~m[380]&m[381]&m[382]&~m[383]&m[397])|(m[380]&m[381]&m[382]&~m[383]&m[397])|(m[380]&m[381]&m[382]&m[383]&m[397]));
    m[389] = (((m[385]&~m[386]&~m[387]&~m[388]&~m[402])|(~m[385]&m[386]&~m[387]&~m[388]&~m[402])|(~m[385]&~m[386]&m[387]&~m[388]&~m[402])|(m[385]&m[386]&~m[387]&m[388]&~m[402])|(m[385]&~m[386]&m[387]&m[388]&~m[402])|(~m[385]&m[386]&m[387]&m[388]&~m[402]))&BiasedRNG[344])|(((m[385]&~m[386]&~m[387]&~m[388]&m[402])|(~m[385]&m[386]&~m[387]&~m[388]&m[402])|(~m[385]&~m[386]&m[387]&~m[388]&m[402])|(m[385]&m[386]&~m[387]&m[388]&m[402])|(m[385]&~m[386]&m[387]&m[388]&m[402])|(~m[385]&m[386]&m[387]&m[388]&m[402]))&~BiasedRNG[344])|((m[385]&m[386]&~m[387]&~m[388]&~m[402])|(m[385]&~m[386]&m[387]&~m[388]&~m[402])|(~m[385]&m[386]&m[387]&~m[388]&~m[402])|(m[385]&m[386]&m[387]&~m[388]&~m[402])|(m[385]&m[386]&m[387]&m[388]&~m[402])|(m[385]&m[386]&~m[387]&~m[388]&m[402])|(m[385]&~m[386]&m[387]&~m[388]&m[402])|(~m[385]&m[386]&m[387]&~m[388]&m[402])|(m[385]&m[386]&m[387]&~m[388]&m[402])|(m[385]&m[386]&m[387]&m[388]&m[402]));
    m[394] = (((m[390]&~m[391]&~m[392]&~m[393]&~m[412])|(~m[390]&m[391]&~m[392]&~m[393]&~m[412])|(~m[390]&~m[391]&m[392]&~m[393]&~m[412])|(m[390]&m[391]&~m[392]&m[393]&~m[412])|(m[390]&~m[391]&m[392]&m[393]&~m[412])|(~m[390]&m[391]&m[392]&m[393]&~m[412]))&BiasedRNG[345])|(((m[390]&~m[391]&~m[392]&~m[393]&m[412])|(~m[390]&m[391]&~m[392]&~m[393]&m[412])|(~m[390]&~m[391]&m[392]&~m[393]&m[412])|(m[390]&m[391]&~m[392]&m[393]&m[412])|(m[390]&~m[391]&m[392]&m[393]&m[412])|(~m[390]&m[391]&m[392]&m[393]&m[412]))&~BiasedRNG[345])|((m[390]&m[391]&~m[392]&~m[393]&~m[412])|(m[390]&~m[391]&m[392]&~m[393]&~m[412])|(~m[390]&m[391]&m[392]&~m[393]&~m[412])|(m[390]&m[391]&m[392]&~m[393]&~m[412])|(m[390]&m[391]&m[392]&m[393]&~m[412])|(m[390]&m[391]&~m[392]&~m[393]&m[412])|(m[390]&~m[391]&m[392]&~m[393]&m[412])|(~m[390]&m[391]&m[392]&~m[393]&m[412])|(m[390]&m[391]&m[392]&~m[393]&m[412])|(m[390]&m[391]&m[392]&m[393]&m[412]));
    m[399] = (((m[395]&~m[396]&~m[397]&~m[398]&~m[417])|(~m[395]&m[396]&~m[397]&~m[398]&~m[417])|(~m[395]&~m[396]&m[397]&~m[398]&~m[417])|(m[395]&m[396]&~m[397]&m[398]&~m[417])|(m[395]&~m[396]&m[397]&m[398]&~m[417])|(~m[395]&m[396]&m[397]&m[398]&~m[417]))&BiasedRNG[346])|(((m[395]&~m[396]&~m[397]&~m[398]&m[417])|(~m[395]&m[396]&~m[397]&~m[398]&m[417])|(~m[395]&~m[396]&m[397]&~m[398]&m[417])|(m[395]&m[396]&~m[397]&m[398]&m[417])|(m[395]&~m[396]&m[397]&m[398]&m[417])|(~m[395]&m[396]&m[397]&m[398]&m[417]))&~BiasedRNG[346])|((m[395]&m[396]&~m[397]&~m[398]&~m[417])|(m[395]&~m[396]&m[397]&~m[398]&~m[417])|(~m[395]&m[396]&m[397]&~m[398]&~m[417])|(m[395]&m[396]&m[397]&~m[398]&~m[417])|(m[395]&m[396]&m[397]&m[398]&~m[417])|(m[395]&m[396]&~m[397]&~m[398]&m[417])|(m[395]&~m[396]&m[397]&~m[398]&m[417])|(~m[395]&m[396]&m[397]&~m[398]&m[417])|(m[395]&m[396]&m[397]&~m[398]&m[417])|(m[395]&m[396]&m[397]&m[398]&m[417]));
    m[404] = (((m[400]&~m[401]&~m[402]&~m[403]&~m[422])|(~m[400]&m[401]&~m[402]&~m[403]&~m[422])|(~m[400]&~m[401]&m[402]&~m[403]&~m[422])|(m[400]&m[401]&~m[402]&m[403]&~m[422])|(m[400]&~m[401]&m[402]&m[403]&~m[422])|(~m[400]&m[401]&m[402]&m[403]&~m[422]))&BiasedRNG[347])|(((m[400]&~m[401]&~m[402]&~m[403]&m[422])|(~m[400]&m[401]&~m[402]&~m[403]&m[422])|(~m[400]&~m[401]&m[402]&~m[403]&m[422])|(m[400]&m[401]&~m[402]&m[403]&m[422])|(m[400]&~m[401]&m[402]&m[403]&m[422])|(~m[400]&m[401]&m[402]&m[403]&m[422]))&~BiasedRNG[347])|((m[400]&m[401]&~m[402]&~m[403]&~m[422])|(m[400]&~m[401]&m[402]&~m[403]&~m[422])|(~m[400]&m[401]&m[402]&~m[403]&~m[422])|(m[400]&m[401]&m[402]&~m[403]&~m[422])|(m[400]&m[401]&m[402]&m[403]&~m[422])|(m[400]&m[401]&~m[402]&~m[403]&m[422])|(m[400]&~m[401]&m[402]&~m[403]&m[422])|(~m[400]&m[401]&m[402]&~m[403]&m[422])|(m[400]&m[401]&m[402]&~m[403]&m[422])|(m[400]&m[401]&m[402]&m[403]&m[422]));
    m[409] = (((m[405]&~m[406]&~m[407]&~m[408]&~m[427])|(~m[405]&m[406]&~m[407]&~m[408]&~m[427])|(~m[405]&~m[406]&m[407]&~m[408]&~m[427])|(m[405]&m[406]&~m[407]&m[408]&~m[427])|(m[405]&~m[406]&m[407]&m[408]&~m[427])|(~m[405]&m[406]&m[407]&m[408]&~m[427]))&BiasedRNG[348])|(((m[405]&~m[406]&~m[407]&~m[408]&m[427])|(~m[405]&m[406]&~m[407]&~m[408]&m[427])|(~m[405]&~m[406]&m[407]&~m[408]&m[427])|(m[405]&m[406]&~m[407]&m[408]&m[427])|(m[405]&~m[406]&m[407]&m[408]&m[427])|(~m[405]&m[406]&m[407]&m[408]&m[427]))&~BiasedRNG[348])|((m[405]&m[406]&~m[407]&~m[408]&~m[427])|(m[405]&~m[406]&m[407]&~m[408]&~m[427])|(~m[405]&m[406]&m[407]&~m[408]&~m[427])|(m[405]&m[406]&m[407]&~m[408]&~m[427])|(m[405]&m[406]&m[407]&m[408]&~m[427])|(m[405]&m[406]&~m[407]&~m[408]&m[427])|(m[405]&~m[406]&m[407]&~m[408]&m[427])|(~m[405]&m[406]&m[407]&~m[408]&m[427])|(m[405]&m[406]&m[407]&~m[408]&m[427])|(m[405]&m[406]&m[407]&m[408]&m[427]));
    m[414] = (((m[410]&~m[411]&~m[412]&~m[413]&~m[437])|(~m[410]&m[411]&~m[412]&~m[413]&~m[437])|(~m[410]&~m[411]&m[412]&~m[413]&~m[437])|(m[410]&m[411]&~m[412]&m[413]&~m[437])|(m[410]&~m[411]&m[412]&m[413]&~m[437])|(~m[410]&m[411]&m[412]&m[413]&~m[437]))&BiasedRNG[349])|(((m[410]&~m[411]&~m[412]&~m[413]&m[437])|(~m[410]&m[411]&~m[412]&~m[413]&m[437])|(~m[410]&~m[411]&m[412]&~m[413]&m[437])|(m[410]&m[411]&~m[412]&m[413]&m[437])|(m[410]&~m[411]&m[412]&m[413]&m[437])|(~m[410]&m[411]&m[412]&m[413]&m[437]))&~BiasedRNG[349])|((m[410]&m[411]&~m[412]&~m[413]&~m[437])|(m[410]&~m[411]&m[412]&~m[413]&~m[437])|(~m[410]&m[411]&m[412]&~m[413]&~m[437])|(m[410]&m[411]&m[412]&~m[413]&~m[437])|(m[410]&m[411]&m[412]&m[413]&~m[437])|(m[410]&m[411]&~m[412]&~m[413]&m[437])|(m[410]&~m[411]&m[412]&~m[413]&m[437])|(~m[410]&m[411]&m[412]&~m[413]&m[437])|(m[410]&m[411]&m[412]&~m[413]&m[437])|(m[410]&m[411]&m[412]&m[413]&m[437]));
    m[419] = (((m[415]&~m[416]&~m[417]&~m[418]&~m[442])|(~m[415]&m[416]&~m[417]&~m[418]&~m[442])|(~m[415]&~m[416]&m[417]&~m[418]&~m[442])|(m[415]&m[416]&~m[417]&m[418]&~m[442])|(m[415]&~m[416]&m[417]&m[418]&~m[442])|(~m[415]&m[416]&m[417]&m[418]&~m[442]))&BiasedRNG[350])|(((m[415]&~m[416]&~m[417]&~m[418]&m[442])|(~m[415]&m[416]&~m[417]&~m[418]&m[442])|(~m[415]&~m[416]&m[417]&~m[418]&m[442])|(m[415]&m[416]&~m[417]&m[418]&m[442])|(m[415]&~m[416]&m[417]&m[418]&m[442])|(~m[415]&m[416]&m[417]&m[418]&m[442]))&~BiasedRNG[350])|((m[415]&m[416]&~m[417]&~m[418]&~m[442])|(m[415]&~m[416]&m[417]&~m[418]&~m[442])|(~m[415]&m[416]&m[417]&~m[418]&~m[442])|(m[415]&m[416]&m[417]&~m[418]&~m[442])|(m[415]&m[416]&m[417]&m[418]&~m[442])|(m[415]&m[416]&~m[417]&~m[418]&m[442])|(m[415]&~m[416]&m[417]&~m[418]&m[442])|(~m[415]&m[416]&m[417]&~m[418]&m[442])|(m[415]&m[416]&m[417]&~m[418]&m[442])|(m[415]&m[416]&m[417]&m[418]&m[442]));
    m[424] = (((m[420]&~m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&~m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&~m[422]&m[423]&~m[447])|(m[420]&~m[421]&m[422]&m[423]&~m[447])|(~m[420]&m[421]&m[422]&m[423]&~m[447]))&BiasedRNG[351])|(((m[420]&~m[421]&~m[422]&~m[423]&m[447])|(~m[420]&m[421]&~m[422]&~m[423]&m[447])|(~m[420]&~m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&~m[422]&m[423]&m[447])|(m[420]&~m[421]&m[422]&m[423]&m[447])|(~m[420]&m[421]&m[422]&m[423]&m[447]))&~BiasedRNG[351])|((m[420]&m[421]&~m[422]&~m[423]&~m[447])|(m[420]&~m[421]&m[422]&~m[423]&~m[447])|(~m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&m[423]&~m[447])|(m[420]&m[421]&~m[422]&~m[423]&m[447])|(m[420]&~m[421]&m[422]&~m[423]&m[447])|(~m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&m[423]&m[447]));
    m[429] = (((m[425]&~m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&~m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&~m[427]&m[428]&~m[452])|(m[425]&~m[426]&m[427]&m[428]&~m[452])|(~m[425]&m[426]&m[427]&m[428]&~m[452]))&BiasedRNG[352])|(((m[425]&~m[426]&~m[427]&~m[428]&m[452])|(~m[425]&m[426]&~m[427]&~m[428]&m[452])|(~m[425]&~m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&~m[427]&m[428]&m[452])|(m[425]&~m[426]&m[427]&m[428]&m[452])|(~m[425]&m[426]&m[427]&m[428]&m[452]))&~BiasedRNG[352])|((m[425]&m[426]&~m[427]&~m[428]&~m[452])|(m[425]&~m[426]&m[427]&~m[428]&~m[452])|(~m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&m[428]&~m[452])|(m[425]&m[426]&~m[427]&~m[428]&m[452])|(m[425]&~m[426]&m[427]&~m[428]&m[452])|(~m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&m[428]&m[452]));
    m[434] = (((m[430]&~m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&~m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&~m[432]&m[433]&~m[457])|(m[430]&~m[431]&m[432]&m[433]&~m[457])|(~m[430]&m[431]&m[432]&m[433]&~m[457]))&BiasedRNG[353])|(((m[430]&~m[431]&~m[432]&~m[433]&m[457])|(~m[430]&m[431]&~m[432]&~m[433]&m[457])|(~m[430]&~m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&~m[432]&m[433]&m[457])|(m[430]&~m[431]&m[432]&m[433]&m[457])|(~m[430]&m[431]&m[432]&m[433]&m[457]))&~BiasedRNG[353])|((m[430]&m[431]&~m[432]&~m[433]&~m[457])|(m[430]&~m[431]&m[432]&~m[433]&~m[457])|(~m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&m[433]&~m[457])|(m[430]&m[431]&~m[432]&~m[433]&m[457])|(m[430]&~m[431]&m[432]&~m[433]&m[457])|(~m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&m[433]&m[457]));
    m[439] = (((m[435]&~m[436]&~m[437]&~m[438]&~m[467])|(~m[435]&m[436]&~m[437]&~m[438]&~m[467])|(~m[435]&~m[436]&m[437]&~m[438]&~m[467])|(m[435]&m[436]&~m[437]&m[438]&~m[467])|(m[435]&~m[436]&m[437]&m[438]&~m[467])|(~m[435]&m[436]&m[437]&m[438]&~m[467]))&BiasedRNG[354])|(((m[435]&~m[436]&~m[437]&~m[438]&m[467])|(~m[435]&m[436]&~m[437]&~m[438]&m[467])|(~m[435]&~m[436]&m[437]&~m[438]&m[467])|(m[435]&m[436]&~m[437]&m[438]&m[467])|(m[435]&~m[436]&m[437]&m[438]&m[467])|(~m[435]&m[436]&m[437]&m[438]&m[467]))&~BiasedRNG[354])|((m[435]&m[436]&~m[437]&~m[438]&~m[467])|(m[435]&~m[436]&m[437]&~m[438]&~m[467])|(~m[435]&m[436]&m[437]&~m[438]&~m[467])|(m[435]&m[436]&m[437]&~m[438]&~m[467])|(m[435]&m[436]&m[437]&m[438]&~m[467])|(m[435]&m[436]&~m[437]&~m[438]&m[467])|(m[435]&~m[436]&m[437]&~m[438]&m[467])|(~m[435]&m[436]&m[437]&~m[438]&m[467])|(m[435]&m[436]&m[437]&~m[438]&m[467])|(m[435]&m[436]&m[437]&m[438]&m[467]));
    m[444] = (((m[440]&~m[441]&~m[442]&~m[443]&~m[472])|(~m[440]&m[441]&~m[442]&~m[443]&~m[472])|(~m[440]&~m[441]&m[442]&~m[443]&~m[472])|(m[440]&m[441]&~m[442]&m[443]&~m[472])|(m[440]&~m[441]&m[442]&m[443]&~m[472])|(~m[440]&m[441]&m[442]&m[443]&~m[472]))&BiasedRNG[355])|(((m[440]&~m[441]&~m[442]&~m[443]&m[472])|(~m[440]&m[441]&~m[442]&~m[443]&m[472])|(~m[440]&~m[441]&m[442]&~m[443]&m[472])|(m[440]&m[441]&~m[442]&m[443]&m[472])|(m[440]&~m[441]&m[442]&m[443]&m[472])|(~m[440]&m[441]&m[442]&m[443]&m[472]))&~BiasedRNG[355])|((m[440]&m[441]&~m[442]&~m[443]&~m[472])|(m[440]&~m[441]&m[442]&~m[443]&~m[472])|(~m[440]&m[441]&m[442]&~m[443]&~m[472])|(m[440]&m[441]&m[442]&~m[443]&~m[472])|(m[440]&m[441]&m[442]&m[443]&~m[472])|(m[440]&m[441]&~m[442]&~m[443]&m[472])|(m[440]&~m[441]&m[442]&~m[443]&m[472])|(~m[440]&m[441]&m[442]&~m[443]&m[472])|(m[440]&m[441]&m[442]&~m[443]&m[472])|(m[440]&m[441]&m[442]&m[443]&m[472]));
    m[449] = (((m[445]&~m[446]&~m[447]&~m[448]&~m[477])|(~m[445]&m[446]&~m[447]&~m[448]&~m[477])|(~m[445]&~m[446]&m[447]&~m[448]&~m[477])|(m[445]&m[446]&~m[447]&m[448]&~m[477])|(m[445]&~m[446]&m[447]&m[448]&~m[477])|(~m[445]&m[446]&m[447]&m[448]&~m[477]))&BiasedRNG[356])|(((m[445]&~m[446]&~m[447]&~m[448]&m[477])|(~m[445]&m[446]&~m[447]&~m[448]&m[477])|(~m[445]&~m[446]&m[447]&~m[448]&m[477])|(m[445]&m[446]&~m[447]&m[448]&m[477])|(m[445]&~m[446]&m[447]&m[448]&m[477])|(~m[445]&m[446]&m[447]&m[448]&m[477]))&~BiasedRNG[356])|((m[445]&m[446]&~m[447]&~m[448]&~m[477])|(m[445]&~m[446]&m[447]&~m[448]&~m[477])|(~m[445]&m[446]&m[447]&~m[448]&~m[477])|(m[445]&m[446]&m[447]&~m[448]&~m[477])|(m[445]&m[446]&m[447]&m[448]&~m[477])|(m[445]&m[446]&~m[447]&~m[448]&m[477])|(m[445]&~m[446]&m[447]&~m[448]&m[477])|(~m[445]&m[446]&m[447]&~m[448]&m[477])|(m[445]&m[446]&m[447]&~m[448]&m[477])|(m[445]&m[446]&m[447]&m[448]&m[477]));
    m[454] = (((m[450]&~m[451]&~m[452]&~m[453]&~m[482])|(~m[450]&m[451]&~m[452]&~m[453]&~m[482])|(~m[450]&~m[451]&m[452]&~m[453]&~m[482])|(m[450]&m[451]&~m[452]&m[453]&~m[482])|(m[450]&~m[451]&m[452]&m[453]&~m[482])|(~m[450]&m[451]&m[452]&m[453]&~m[482]))&BiasedRNG[357])|(((m[450]&~m[451]&~m[452]&~m[453]&m[482])|(~m[450]&m[451]&~m[452]&~m[453]&m[482])|(~m[450]&~m[451]&m[452]&~m[453]&m[482])|(m[450]&m[451]&~m[452]&m[453]&m[482])|(m[450]&~m[451]&m[452]&m[453]&m[482])|(~m[450]&m[451]&m[452]&m[453]&m[482]))&~BiasedRNG[357])|((m[450]&m[451]&~m[452]&~m[453]&~m[482])|(m[450]&~m[451]&m[452]&~m[453]&~m[482])|(~m[450]&m[451]&m[452]&~m[453]&~m[482])|(m[450]&m[451]&m[452]&~m[453]&~m[482])|(m[450]&m[451]&m[452]&m[453]&~m[482])|(m[450]&m[451]&~m[452]&~m[453]&m[482])|(m[450]&~m[451]&m[452]&~m[453]&m[482])|(~m[450]&m[451]&m[452]&~m[453]&m[482])|(m[450]&m[451]&m[452]&~m[453]&m[482])|(m[450]&m[451]&m[452]&m[453]&m[482]));
    m[459] = (((m[455]&~m[456]&~m[457]&~m[458]&~m[487])|(~m[455]&m[456]&~m[457]&~m[458]&~m[487])|(~m[455]&~m[456]&m[457]&~m[458]&~m[487])|(m[455]&m[456]&~m[457]&m[458]&~m[487])|(m[455]&~m[456]&m[457]&m[458]&~m[487])|(~m[455]&m[456]&m[457]&m[458]&~m[487]))&BiasedRNG[358])|(((m[455]&~m[456]&~m[457]&~m[458]&m[487])|(~m[455]&m[456]&~m[457]&~m[458]&m[487])|(~m[455]&~m[456]&m[457]&~m[458]&m[487])|(m[455]&m[456]&~m[457]&m[458]&m[487])|(m[455]&~m[456]&m[457]&m[458]&m[487])|(~m[455]&m[456]&m[457]&m[458]&m[487]))&~BiasedRNG[358])|((m[455]&m[456]&~m[457]&~m[458]&~m[487])|(m[455]&~m[456]&m[457]&~m[458]&~m[487])|(~m[455]&m[456]&m[457]&~m[458]&~m[487])|(m[455]&m[456]&m[457]&~m[458]&~m[487])|(m[455]&m[456]&m[457]&m[458]&~m[487])|(m[455]&m[456]&~m[457]&~m[458]&m[487])|(m[455]&~m[456]&m[457]&~m[458]&m[487])|(~m[455]&m[456]&m[457]&~m[458]&m[487])|(m[455]&m[456]&m[457]&~m[458]&m[487])|(m[455]&m[456]&m[457]&m[458]&m[487]));
    m[464] = (((m[460]&~m[461]&~m[462]&~m[463]&~m[492])|(~m[460]&m[461]&~m[462]&~m[463]&~m[492])|(~m[460]&~m[461]&m[462]&~m[463]&~m[492])|(m[460]&m[461]&~m[462]&m[463]&~m[492])|(m[460]&~m[461]&m[462]&m[463]&~m[492])|(~m[460]&m[461]&m[462]&m[463]&~m[492]))&BiasedRNG[359])|(((m[460]&~m[461]&~m[462]&~m[463]&m[492])|(~m[460]&m[461]&~m[462]&~m[463]&m[492])|(~m[460]&~m[461]&m[462]&~m[463]&m[492])|(m[460]&m[461]&~m[462]&m[463]&m[492])|(m[460]&~m[461]&m[462]&m[463]&m[492])|(~m[460]&m[461]&m[462]&m[463]&m[492]))&~BiasedRNG[359])|((m[460]&m[461]&~m[462]&~m[463]&~m[492])|(m[460]&~m[461]&m[462]&~m[463]&~m[492])|(~m[460]&m[461]&m[462]&~m[463]&~m[492])|(m[460]&m[461]&m[462]&~m[463]&~m[492])|(m[460]&m[461]&m[462]&m[463]&~m[492])|(m[460]&m[461]&~m[462]&~m[463]&m[492])|(m[460]&~m[461]&m[462]&~m[463]&m[492])|(~m[460]&m[461]&m[462]&~m[463]&m[492])|(m[460]&m[461]&m[462]&~m[463]&m[492])|(m[460]&m[461]&m[462]&m[463]&m[492]));
    m[469] = (((m[465]&~m[466]&~m[467]&~m[468]&~m[502])|(~m[465]&m[466]&~m[467]&~m[468]&~m[502])|(~m[465]&~m[466]&m[467]&~m[468]&~m[502])|(m[465]&m[466]&~m[467]&m[468]&~m[502])|(m[465]&~m[466]&m[467]&m[468]&~m[502])|(~m[465]&m[466]&m[467]&m[468]&~m[502]))&BiasedRNG[360])|(((m[465]&~m[466]&~m[467]&~m[468]&m[502])|(~m[465]&m[466]&~m[467]&~m[468]&m[502])|(~m[465]&~m[466]&m[467]&~m[468]&m[502])|(m[465]&m[466]&~m[467]&m[468]&m[502])|(m[465]&~m[466]&m[467]&m[468]&m[502])|(~m[465]&m[466]&m[467]&m[468]&m[502]))&~BiasedRNG[360])|((m[465]&m[466]&~m[467]&~m[468]&~m[502])|(m[465]&~m[466]&m[467]&~m[468]&~m[502])|(~m[465]&m[466]&m[467]&~m[468]&~m[502])|(m[465]&m[466]&m[467]&~m[468]&~m[502])|(m[465]&m[466]&m[467]&m[468]&~m[502])|(m[465]&m[466]&~m[467]&~m[468]&m[502])|(m[465]&~m[466]&m[467]&~m[468]&m[502])|(~m[465]&m[466]&m[467]&~m[468]&m[502])|(m[465]&m[466]&m[467]&~m[468]&m[502])|(m[465]&m[466]&m[467]&m[468]&m[502]));
    m[474] = (((m[470]&~m[471]&~m[472]&~m[473]&~m[507])|(~m[470]&m[471]&~m[472]&~m[473]&~m[507])|(~m[470]&~m[471]&m[472]&~m[473]&~m[507])|(m[470]&m[471]&~m[472]&m[473]&~m[507])|(m[470]&~m[471]&m[472]&m[473]&~m[507])|(~m[470]&m[471]&m[472]&m[473]&~m[507]))&BiasedRNG[361])|(((m[470]&~m[471]&~m[472]&~m[473]&m[507])|(~m[470]&m[471]&~m[472]&~m[473]&m[507])|(~m[470]&~m[471]&m[472]&~m[473]&m[507])|(m[470]&m[471]&~m[472]&m[473]&m[507])|(m[470]&~m[471]&m[472]&m[473]&m[507])|(~m[470]&m[471]&m[472]&m[473]&m[507]))&~BiasedRNG[361])|((m[470]&m[471]&~m[472]&~m[473]&~m[507])|(m[470]&~m[471]&m[472]&~m[473]&~m[507])|(~m[470]&m[471]&m[472]&~m[473]&~m[507])|(m[470]&m[471]&m[472]&~m[473]&~m[507])|(m[470]&m[471]&m[472]&m[473]&~m[507])|(m[470]&m[471]&~m[472]&~m[473]&m[507])|(m[470]&~m[471]&m[472]&~m[473]&m[507])|(~m[470]&m[471]&m[472]&~m[473]&m[507])|(m[470]&m[471]&m[472]&~m[473]&m[507])|(m[470]&m[471]&m[472]&m[473]&m[507]));
    m[479] = (((m[475]&~m[476]&~m[477]&~m[478]&~m[512])|(~m[475]&m[476]&~m[477]&~m[478]&~m[512])|(~m[475]&~m[476]&m[477]&~m[478]&~m[512])|(m[475]&m[476]&~m[477]&m[478]&~m[512])|(m[475]&~m[476]&m[477]&m[478]&~m[512])|(~m[475]&m[476]&m[477]&m[478]&~m[512]))&BiasedRNG[362])|(((m[475]&~m[476]&~m[477]&~m[478]&m[512])|(~m[475]&m[476]&~m[477]&~m[478]&m[512])|(~m[475]&~m[476]&m[477]&~m[478]&m[512])|(m[475]&m[476]&~m[477]&m[478]&m[512])|(m[475]&~m[476]&m[477]&m[478]&m[512])|(~m[475]&m[476]&m[477]&m[478]&m[512]))&~BiasedRNG[362])|((m[475]&m[476]&~m[477]&~m[478]&~m[512])|(m[475]&~m[476]&m[477]&~m[478]&~m[512])|(~m[475]&m[476]&m[477]&~m[478]&~m[512])|(m[475]&m[476]&m[477]&~m[478]&~m[512])|(m[475]&m[476]&m[477]&m[478]&~m[512])|(m[475]&m[476]&~m[477]&~m[478]&m[512])|(m[475]&~m[476]&m[477]&~m[478]&m[512])|(~m[475]&m[476]&m[477]&~m[478]&m[512])|(m[475]&m[476]&m[477]&~m[478]&m[512])|(m[475]&m[476]&m[477]&m[478]&m[512]));
    m[484] = (((m[480]&~m[481]&~m[482]&~m[483]&~m[517])|(~m[480]&m[481]&~m[482]&~m[483]&~m[517])|(~m[480]&~m[481]&m[482]&~m[483]&~m[517])|(m[480]&m[481]&~m[482]&m[483]&~m[517])|(m[480]&~m[481]&m[482]&m[483]&~m[517])|(~m[480]&m[481]&m[482]&m[483]&~m[517]))&BiasedRNG[363])|(((m[480]&~m[481]&~m[482]&~m[483]&m[517])|(~m[480]&m[481]&~m[482]&~m[483]&m[517])|(~m[480]&~m[481]&m[482]&~m[483]&m[517])|(m[480]&m[481]&~m[482]&m[483]&m[517])|(m[480]&~m[481]&m[482]&m[483]&m[517])|(~m[480]&m[481]&m[482]&m[483]&m[517]))&~BiasedRNG[363])|((m[480]&m[481]&~m[482]&~m[483]&~m[517])|(m[480]&~m[481]&m[482]&~m[483]&~m[517])|(~m[480]&m[481]&m[482]&~m[483]&~m[517])|(m[480]&m[481]&m[482]&~m[483]&~m[517])|(m[480]&m[481]&m[482]&m[483]&~m[517])|(m[480]&m[481]&~m[482]&~m[483]&m[517])|(m[480]&~m[481]&m[482]&~m[483]&m[517])|(~m[480]&m[481]&m[482]&~m[483]&m[517])|(m[480]&m[481]&m[482]&~m[483]&m[517])|(m[480]&m[481]&m[482]&m[483]&m[517]));
    m[489] = (((m[485]&~m[486]&~m[487]&~m[488]&~m[522])|(~m[485]&m[486]&~m[487]&~m[488]&~m[522])|(~m[485]&~m[486]&m[487]&~m[488]&~m[522])|(m[485]&m[486]&~m[487]&m[488]&~m[522])|(m[485]&~m[486]&m[487]&m[488]&~m[522])|(~m[485]&m[486]&m[487]&m[488]&~m[522]))&BiasedRNG[364])|(((m[485]&~m[486]&~m[487]&~m[488]&m[522])|(~m[485]&m[486]&~m[487]&~m[488]&m[522])|(~m[485]&~m[486]&m[487]&~m[488]&m[522])|(m[485]&m[486]&~m[487]&m[488]&m[522])|(m[485]&~m[486]&m[487]&m[488]&m[522])|(~m[485]&m[486]&m[487]&m[488]&m[522]))&~BiasedRNG[364])|((m[485]&m[486]&~m[487]&~m[488]&~m[522])|(m[485]&~m[486]&m[487]&~m[488]&~m[522])|(~m[485]&m[486]&m[487]&~m[488]&~m[522])|(m[485]&m[486]&m[487]&~m[488]&~m[522])|(m[485]&m[486]&m[487]&m[488]&~m[522])|(m[485]&m[486]&~m[487]&~m[488]&m[522])|(m[485]&~m[486]&m[487]&~m[488]&m[522])|(~m[485]&m[486]&m[487]&~m[488]&m[522])|(m[485]&m[486]&m[487]&~m[488]&m[522])|(m[485]&m[486]&m[487]&m[488]&m[522]));
    m[494] = (((m[490]&~m[491]&~m[492]&~m[493]&~m[527])|(~m[490]&m[491]&~m[492]&~m[493]&~m[527])|(~m[490]&~m[491]&m[492]&~m[493]&~m[527])|(m[490]&m[491]&~m[492]&m[493]&~m[527])|(m[490]&~m[491]&m[492]&m[493]&~m[527])|(~m[490]&m[491]&m[492]&m[493]&~m[527]))&BiasedRNG[365])|(((m[490]&~m[491]&~m[492]&~m[493]&m[527])|(~m[490]&m[491]&~m[492]&~m[493]&m[527])|(~m[490]&~m[491]&m[492]&~m[493]&m[527])|(m[490]&m[491]&~m[492]&m[493]&m[527])|(m[490]&~m[491]&m[492]&m[493]&m[527])|(~m[490]&m[491]&m[492]&m[493]&m[527]))&~BiasedRNG[365])|((m[490]&m[491]&~m[492]&~m[493]&~m[527])|(m[490]&~m[491]&m[492]&~m[493]&~m[527])|(~m[490]&m[491]&m[492]&~m[493]&~m[527])|(m[490]&m[491]&m[492]&~m[493]&~m[527])|(m[490]&m[491]&m[492]&m[493]&~m[527])|(m[490]&m[491]&~m[492]&~m[493]&m[527])|(m[490]&~m[491]&m[492]&~m[493]&m[527])|(~m[490]&m[491]&m[492]&~m[493]&m[527])|(m[490]&m[491]&m[492]&~m[493]&m[527])|(m[490]&m[491]&m[492]&m[493]&m[527]));
    m[499] = (((m[495]&~m[496]&~m[497]&~m[498]&~m[532])|(~m[495]&m[496]&~m[497]&~m[498]&~m[532])|(~m[495]&~m[496]&m[497]&~m[498]&~m[532])|(m[495]&m[496]&~m[497]&m[498]&~m[532])|(m[495]&~m[496]&m[497]&m[498]&~m[532])|(~m[495]&m[496]&m[497]&m[498]&~m[532]))&BiasedRNG[366])|(((m[495]&~m[496]&~m[497]&~m[498]&m[532])|(~m[495]&m[496]&~m[497]&~m[498]&m[532])|(~m[495]&~m[496]&m[497]&~m[498]&m[532])|(m[495]&m[496]&~m[497]&m[498]&m[532])|(m[495]&~m[496]&m[497]&m[498]&m[532])|(~m[495]&m[496]&m[497]&m[498]&m[532]))&~BiasedRNG[366])|((m[495]&m[496]&~m[497]&~m[498]&~m[532])|(m[495]&~m[496]&m[497]&~m[498]&~m[532])|(~m[495]&m[496]&m[497]&~m[498]&~m[532])|(m[495]&m[496]&m[497]&~m[498]&~m[532])|(m[495]&m[496]&m[497]&m[498]&~m[532])|(m[495]&m[496]&~m[497]&~m[498]&m[532])|(m[495]&~m[496]&m[497]&~m[498]&m[532])|(~m[495]&m[496]&m[497]&~m[498]&m[532])|(m[495]&m[496]&m[497]&~m[498]&m[532])|(m[495]&m[496]&m[497]&m[498]&m[532]));
    m[504] = (((m[500]&~m[501]&~m[502]&~m[503]&~m[542])|(~m[500]&m[501]&~m[502]&~m[503]&~m[542])|(~m[500]&~m[501]&m[502]&~m[503]&~m[542])|(m[500]&m[501]&~m[502]&m[503]&~m[542])|(m[500]&~m[501]&m[502]&m[503]&~m[542])|(~m[500]&m[501]&m[502]&m[503]&~m[542]))&BiasedRNG[367])|(((m[500]&~m[501]&~m[502]&~m[503]&m[542])|(~m[500]&m[501]&~m[502]&~m[503]&m[542])|(~m[500]&~m[501]&m[502]&~m[503]&m[542])|(m[500]&m[501]&~m[502]&m[503]&m[542])|(m[500]&~m[501]&m[502]&m[503]&m[542])|(~m[500]&m[501]&m[502]&m[503]&m[542]))&~BiasedRNG[367])|((m[500]&m[501]&~m[502]&~m[503]&~m[542])|(m[500]&~m[501]&m[502]&~m[503]&~m[542])|(~m[500]&m[501]&m[502]&~m[503]&~m[542])|(m[500]&m[501]&m[502]&~m[503]&~m[542])|(m[500]&m[501]&m[502]&m[503]&~m[542])|(m[500]&m[501]&~m[502]&~m[503]&m[542])|(m[500]&~m[501]&m[502]&~m[503]&m[542])|(~m[500]&m[501]&m[502]&~m[503]&m[542])|(m[500]&m[501]&m[502]&~m[503]&m[542])|(m[500]&m[501]&m[502]&m[503]&m[542]));
    m[509] = (((m[505]&~m[506]&~m[507]&~m[508]&~m[547])|(~m[505]&m[506]&~m[507]&~m[508]&~m[547])|(~m[505]&~m[506]&m[507]&~m[508]&~m[547])|(m[505]&m[506]&~m[507]&m[508]&~m[547])|(m[505]&~m[506]&m[507]&m[508]&~m[547])|(~m[505]&m[506]&m[507]&m[508]&~m[547]))&BiasedRNG[368])|(((m[505]&~m[506]&~m[507]&~m[508]&m[547])|(~m[505]&m[506]&~m[507]&~m[508]&m[547])|(~m[505]&~m[506]&m[507]&~m[508]&m[547])|(m[505]&m[506]&~m[507]&m[508]&m[547])|(m[505]&~m[506]&m[507]&m[508]&m[547])|(~m[505]&m[506]&m[507]&m[508]&m[547]))&~BiasedRNG[368])|((m[505]&m[506]&~m[507]&~m[508]&~m[547])|(m[505]&~m[506]&m[507]&~m[508]&~m[547])|(~m[505]&m[506]&m[507]&~m[508]&~m[547])|(m[505]&m[506]&m[507]&~m[508]&~m[547])|(m[505]&m[506]&m[507]&m[508]&~m[547])|(m[505]&m[506]&~m[507]&~m[508]&m[547])|(m[505]&~m[506]&m[507]&~m[508]&m[547])|(~m[505]&m[506]&m[507]&~m[508]&m[547])|(m[505]&m[506]&m[507]&~m[508]&m[547])|(m[505]&m[506]&m[507]&m[508]&m[547]));
    m[514] = (((m[510]&~m[511]&~m[512]&~m[513]&~m[552])|(~m[510]&m[511]&~m[512]&~m[513]&~m[552])|(~m[510]&~m[511]&m[512]&~m[513]&~m[552])|(m[510]&m[511]&~m[512]&m[513]&~m[552])|(m[510]&~m[511]&m[512]&m[513]&~m[552])|(~m[510]&m[511]&m[512]&m[513]&~m[552]))&BiasedRNG[369])|(((m[510]&~m[511]&~m[512]&~m[513]&m[552])|(~m[510]&m[511]&~m[512]&~m[513]&m[552])|(~m[510]&~m[511]&m[512]&~m[513]&m[552])|(m[510]&m[511]&~m[512]&m[513]&m[552])|(m[510]&~m[511]&m[512]&m[513]&m[552])|(~m[510]&m[511]&m[512]&m[513]&m[552]))&~BiasedRNG[369])|((m[510]&m[511]&~m[512]&~m[513]&~m[552])|(m[510]&~m[511]&m[512]&~m[513]&~m[552])|(~m[510]&m[511]&m[512]&~m[513]&~m[552])|(m[510]&m[511]&m[512]&~m[513]&~m[552])|(m[510]&m[511]&m[512]&m[513]&~m[552])|(m[510]&m[511]&~m[512]&~m[513]&m[552])|(m[510]&~m[511]&m[512]&~m[513]&m[552])|(~m[510]&m[511]&m[512]&~m[513]&m[552])|(m[510]&m[511]&m[512]&~m[513]&m[552])|(m[510]&m[511]&m[512]&m[513]&m[552]));
    m[519] = (((m[515]&~m[516]&~m[517]&~m[518]&~m[557])|(~m[515]&m[516]&~m[517]&~m[518]&~m[557])|(~m[515]&~m[516]&m[517]&~m[518]&~m[557])|(m[515]&m[516]&~m[517]&m[518]&~m[557])|(m[515]&~m[516]&m[517]&m[518]&~m[557])|(~m[515]&m[516]&m[517]&m[518]&~m[557]))&BiasedRNG[370])|(((m[515]&~m[516]&~m[517]&~m[518]&m[557])|(~m[515]&m[516]&~m[517]&~m[518]&m[557])|(~m[515]&~m[516]&m[517]&~m[518]&m[557])|(m[515]&m[516]&~m[517]&m[518]&m[557])|(m[515]&~m[516]&m[517]&m[518]&m[557])|(~m[515]&m[516]&m[517]&m[518]&m[557]))&~BiasedRNG[370])|((m[515]&m[516]&~m[517]&~m[518]&~m[557])|(m[515]&~m[516]&m[517]&~m[518]&~m[557])|(~m[515]&m[516]&m[517]&~m[518]&~m[557])|(m[515]&m[516]&m[517]&~m[518]&~m[557])|(m[515]&m[516]&m[517]&m[518]&~m[557])|(m[515]&m[516]&~m[517]&~m[518]&m[557])|(m[515]&~m[516]&m[517]&~m[518]&m[557])|(~m[515]&m[516]&m[517]&~m[518]&m[557])|(m[515]&m[516]&m[517]&~m[518]&m[557])|(m[515]&m[516]&m[517]&m[518]&m[557]));
    m[524] = (((m[520]&~m[521]&~m[522]&~m[523]&~m[562])|(~m[520]&m[521]&~m[522]&~m[523]&~m[562])|(~m[520]&~m[521]&m[522]&~m[523]&~m[562])|(m[520]&m[521]&~m[522]&m[523]&~m[562])|(m[520]&~m[521]&m[522]&m[523]&~m[562])|(~m[520]&m[521]&m[522]&m[523]&~m[562]))&BiasedRNG[371])|(((m[520]&~m[521]&~m[522]&~m[523]&m[562])|(~m[520]&m[521]&~m[522]&~m[523]&m[562])|(~m[520]&~m[521]&m[522]&~m[523]&m[562])|(m[520]&m[521]&~m[522]&m[523]&m[562])|(m[520]&~m[521]&m[522]&m[523]&m[562])|(~m[520]&m[521]&m[522]&m[523]&m[562]))&~BiasedRNG[371])|((m[520]&m[521]&~m[522]&~m[523]&~m[562])|(m[520]&~m[521]&m[522]&~m[523]&~m[562])|(~m[520]&m[521]&m[522]&~m[523]&~m[562])|(m[520]&m[521]&m[522]&~m[523]&~m[562])|(m[520]&m[521]&m[522]&m[523]&~m[562])|(m[520]&m[521]&~m[522]&~m[523]&m[562])|(m[520]&~m[521]&m[522]&~m[523]&m[562])|(~m[520]&m[521]&m[522]&~m[523]&m[562])|(m[520]&m[521]&m[522]&~m[523]&m[562])|(m[520]&m[521]&m[522]&m[523]&m[562]));
    m[529] = (((m[525]&~m[526]&~m[527]&~m[528]&~m[567])|(~m[525]&m[526]&~m[527]&~m[528]&~m[567])|(~m[525]&~m[526]&m[527]&~m[528]&~m[567])|(m[525]&m[526]&~m[527]&m[528]&~m[567])|(m[525]&~m[526]&m[527]&m[528]&~m[567])|(~m[525]&m[526]&m[527]&m[528]&~m[567]))&BiasedRNG[372])|(((m[525]&~m[526]&~m[527]&~m[528]&m[567])|(~m[525]&m[526]&~m[527]&~m[528]&m[567])|(~m[525]&~m[526]&m[527]&~m[528]&m[567])|(m[525]&m[526]&~m[527]&m[528]&m[567])|(m[525]&~m[526]&m[527]&m[528]&m[567])|(~m[525]&m[526]&m[527]&m[528]&m[567]))&~BiasedRNG[372])|((m[525]&m[526]&~m[527]&~m[528]&~m[567])|(m[525]&~m[526]&m[527]&~m[528]&~m[567])|(~m[525]&m[526]&m[527]&~m[528]&~m[567])|(m[525]&m[526]&m[527]&~m[528]&~m[567])|(m[525]&m[526]&m[527]&m[528]&~m[567])|(m[525]&m[526]&~m[527]&~m[528]&m[567])|(m[525]&~m[526]&m[527]&~m[528]&m[567])|(~m[525]&m[526]&m[527]&~m[528]&m[567])|(m[525]&m[526]&m[527]&~m[528]&m[567])|(m[525]&m[526]&m[527]&m[528]&m[567]));
    m[534] = (((m[530]&~m[531]&~m[532]&~m[533]&~m[572])|(~m[530]&m[531]&~m[532]&~m[533]&~m[572])|(~m[530]&~m[531]&m[532]&~m[533]&~m[572])|(m[530]&m[531]&~m[532]&m[533]&~m[572])|(m[530]&~m[531]&m[532]&m[533]&~m[572])|(~m[530]&m[531]&m[532]&m[533]&~m[572]))&BiasedRNG[373])|(((m[530]&~m[531]&~m[532]&~m[533]&m[572])|(~m[530]&m[531]&~m[532]&~m[533]&m[572])|(~m[530]&~m[531]&m[532]&~m[533]&m[572])|(m[530]&m[531]&~m[532]&m[533]&m[572])|(m[530]&~m[531]&m[532]&m[533]&m[572])|(~m[530]&m[531]&m[532]&m[533]&m[572]))&~BiasedRNG[373])|((m[530]&m[531]&~m[532]&~m[533]&~m[572])|(m[530]&~m[531]&m[532]&~m[533]&~m[572])|(~m[530]&m[531]&m[532]&~m[533]&~m[572])|(m[530]&m[531]&m[532]&~m[533]&~m[572])|(m[530]&m[531]&m[532]&m[533]&~m[572])|(m[530]&m[531]&~m[532]&~m[533]&m[572])|(m[530]&~m[531]&m[532]&~m[533]&m[572])|(~m[530]&m[531]&m[532]&~m[533]&m[572])|(m[530]&m[531]&m[532]&~m[533]&m[572])|(m[530]&m[531]&m[532]&m[533]&m[572]));
    m[539] = (((m[535]&~m[536]&~m[537]&~m[538]&~m[577])|(~m[535]&m[536]&~m[537]&~m[538]&~m[577])|(~m[535]&~m[536]&m[537]&~m[538]&~m[577])|(m[535]&m[536]&~m[537]&m[538]&~m[577])|(m[535]&~m[536]&m[537]&m[538]&~m[577])|(~m[535]&m[536]&m[537]&m[538]&~m[577]))&BiasedRNG[374])|(((m[535]&~m[536]&~m[537]&~m[538]&m[577])|(~m[535]&m[536]&~m[537]&~m[538]&m[577])|(~m[535]&~m[536]&m[537]&~m[538]&m[577])|(m[535]&m[536]&~m[537]&m[538]&m[577])|(m[535]&~m[536]&m[537]&m[538]&m[577])|(~m[535]&m[536]&m[537]&m[538]&m[577]))&~BiasedRNG[374])|((m[535]&m[536]&~m[537]&~m[538]&~m[577])|(m[535]&~m[536]&m[537]&~m[538]&~m[577])|(~m[535]&m[536]&m[537]&~m[538]&~m[577])|(m[535]&m[536]&m[537]&~m[538]&~m[577])|(m[535]&m[536]&m[537]&m[538]&~m[577])|(m[535]&m[536]&~m[537]&~m[538]&m[577])|(m[535]&~m[536]&m[537]&~m[538]&m[577])|(~m[535]&m[536]&m[537]&~m[538]&m[577])|(m[535]&m[536]&m[537]&~m[538]&m[577])|(m[535]&m[536]&m[537]&m[538]&m[577]));
    m[544] = (((m[540]&~m[541]&~m[542]&~m[543]&~m[587])|(~m[540]&m[541]&~m[542]&~m[543]&~m[587])|(~m[540]&~m[541]&m[542]&~m[543]&~m[587])|(m[540]&m[541]&~m[542]&m[543]&~m[587])|(m[540]&~m[541]&m[542]&m[543]&~m[587])|(~m[540]&m[541]&m[542]&m[543]&~m[587]))&BiasedRNG[375])|(((m[540]&~m[541]&~m[542]&~m[543]&m[587])|(~m[540]&m[541]&~m[542]&~m[543]&m[587])|(~m[540]&~m[541]&m[542]&~m[543]&m[587])|(m[540]&m[541]&~m[542]&m[543]&m[587])|(m[540]&~m[541]&m[542]&m[543]&m[587])|(~m[540]&m[541]&m[542]&m[543]&m[587]))&~BiasedRNG[375])|((m[540]&m[541]&~m[542]&~m[543]&~m[587])|(m[540]&~m[541]&m[542]&~m[543]&~m[587])|(~m[540]&m[541]&m[542]&~m[543]&~m[587])|(m[540]&m[541]&m[542]&~m[543]&~m[587])|(m[540]&m[541]&m[542]&m[543]&~m[587])|(m[540]&m[541]&~m[542]&~m[543]&m[587])|(m[540]&~m[541]&m[542]&~m[543]&m[587])|(~m[540]&m[541]&m[542]&~m[543]&m[587])|(m[540]&m[541]&m[542]&~m[543]&m[587])|(m[540]&m[541]&m[542]&m[543]&m[587]));
    m[549] = (((m[545]&~m[546]&~m[547]&~m[548]&~m[592])|(~m[545]&m[546]&~m[547]&~m[548]&~m[592])|(~m[545]&~m[546]&m[547]&~m[548]&~m[592])|(m[545]&m[546]&~m[547]&m[548]&~m[592])|(m[545]&~m[546]&m[547]&m[548]&~m[592])|(~m[545]&m[546]&m[547]&m[548]&~m[592]))&BiasedRNG[376])|(((m[545]&~m[546]&~m[547]&~m[548]&m[592])|(~m[545]&m[546]&~m[547]&~m[548]&m[592])|(~m[545]&~m[546]&m[547]&~m[548]&m[592])|(m[545]&m[546]&~m[547]&m[548]&m[592])|(m[545]&~m[546]&m[547]&m[548]&m[592])|(~m[545]&m[546]&m[547]&m[548]&m[592]))&~BiasedRNG[376])|((m[545]&m[546]&~m[547]&~m[548]&~m[592])|(m[545]&~m[546]&m[547]&~m[548]&~m[592])|(~m[545]&m[546]&m[547]&~m[548]&~m[592])|(m[545]&m[546]&m[547]&~m[548]&~m[592])|(m[545]&m[546]&m[547]&m[548]&~m[592])|(m[545]&m[546]&~m[547]&~m[548]&m[592])|(m[545]&~m[546]&m[547]&~m[548]&m[592])|(~m[545]&m[546]&m[547]&~m[548]&m[592])|(m[545]&m[546]&m[547]&~m[548]&m[592])|(m[545]&m[546]&m[547]&m[548]&m[592]));
    m[554] = (((m[550]&~m[551]&~m[552]&~m[553]&~m[597])|(~m[550]&m[551]&~m[552]&~m[553]&~m[597])|(~m[550]&~m[551]&m[552]&~m[553]&~m[597])|(m[550]&m[551]&~m[552]&m[553]&~m[597])|(m[550]&~m[551]&m[552]&m[553]&~m[597])|(~m[550]&m[551]&m[552]&m[553]&~m[597]))&BiasedRNG[377])|(((m[550]&~m[551]&~m[552]&~m[553]&m[597])|(~m[550]&m[551]&~m[552]&~m[553]&m[597])|(~m[550]&~m[551]&m[552]&~m[553]&m[597])|(m[550]&m[551]&~m[552]&m[553]&m[597])|(m[550]&~m[551]&m[552]&m[553]&m[597])|(~m[550]&m[551]&m[552]&m[553]&m[597]))&~BiasedRNG[377])|((m[550]&m[551]&~m[552]&~m[553]&~m[597])|(m[550]&~m[551]&m[552]&~m[553]&~m[597])|(~m[550]&m[551]&m[552]&~m[553]&~m[597])|(m[550]&m[551]&m[552]&~m[553]&~m[597])|(m[550]&m[551]&m[552]&m[553]&~m[597])|(m[550]&m[551]&~m[552]&~m[553]&m[597])|(m[550]&~m[551]&m[552]&~m[553]&m[597])|(~m[550]&m[551]&m[552]&~m[553]&m[597])|(m[550]&m[551]&m[552]&~m[553]&m[597])|(m[550]&m[551]&m[552]&m[553]&m[597]));
    m[559] = (((m[555]&~m[556]&~m[557]&~m[558]&~m[602])|(~m[555]&m[556]&~m[557]&~m[558]&~m[602])|(~m[555]&~m[556]&m[557]&~m[558]&~m[602])|(m[555]&m[556]&~m[557]&m[558]&~m[602])|(m[555]&~m[556]&m[557]&m[558]&~m[602])|(~m[555]&m[556]&m[557]&m[558]&~m[602]))&BiasedRNG[378])|(((m[555]&~m[556]&~m[557]&~m[558]&m[602])|(~m[555]&m[556]&~m[557]&~m[558]&m[602])|(~m[555]&~m[556]&m[557]&~m[558]&m[602])|(m[555]&m[556]&~m[557]&m[558]&m[602])|(m[555]&~m[556]&m[557]&m[558]&m[602])|(~m[555]&m[556]&m[557]&m[558]&m[602]))&~BiasedRNG[378])|((m[555]&m[556]&~m[557]&~m[558]&~m[602])|(m[555]&~m[556]&m[557]&~m[558]&~m[602])|(~m[555]&m[556]&m[557]&~m[558]&~m[602])|(m[555]&m[556]&m[557]&~m[558]&~m[602])|(m[555]&m[556]&m[557]&m[558]&~m[602])|(m[555]&m[556]&~m[557]&~m[558]&m[602])|(m[555]&~m[556]&m[557]&~m[558]&m[602])|(~m[555]&m[556]&m[557]&~m[558]&m[602])|(m[555]&m[556]&m[557]&~m[558]&m[602])|(m[555]&m[556]&m[557]&m[558]&m[602]));
    m[564] = (((m[560]&~m[561]&~m[562]&~m[563]&~m[607])|(~m[560]&m[561]&~m[562]&~m[563]&~m[607])|(~m[560]&~m[561]&m[562]&~m[563]&~m[607])|(m[560]&m[561]&~m[562]&m[563]&~m[607])|(m[560]&~m[561]&m[562]&m[563]&~m[607])|(~m[560]&m[561]&m[562]&m[563]&~m[607]))&BiasedRNG[379])|(((m[560]&~m[561]&~m[562]&~m[563]&m[607])|(~m[560]&m[561]&~m[562]&~m[563]&m[607])|(~m[560]&~m[561]&m[562]&~m[563]&m[607])|(m[560]&m[561]&~m[562]&m[563]&m[607])|(m[560]&~m[561]&m[562]&m[563]&m[607])|(~m[560]&m[561]&m[562]&m[563]&m[607]))&~BiasedRNG[379])|((m[560]&m[561]&~m[562]&~m[563]&~m[607])|(m[560]&~m[561]&m[562]&~m[563]&~m[607])|(~m[560]&m[561]&m[562]&~m[563]&~m[607])|(m[560]&m[561]&m[562]&~m[563]&~m[607])|(m[560]&m[561]&m[562]&m[563]&~m[607])|(m[560]&m[561]&~m[562]&~m[563]&m[607])|(m[560]&~m[561]&m[562]&~m[563]&m[607])|(~m[560]&m[561]&m[562]&~m[563]&m[607])|(m[560]&m[561]&m[562]&~m[563]&m[607])|(m[560]&m[561]&m[562]&m[563]&m[607]));
    m[569] = (((m[565]&~m[566]&~m[567]&~m[568]&~m[612])|(~m[565]&m[566]&~m[567]&~m[568]&~m[612])|(~m[565]&~m[566]&m[567]&~m[568]&~m[612])|(m[565]&m[566]&~m[567]&m[568]&~m[612])|(m[565]&~m[566]&m[567]&m[568]&~m[612])|(~m[565]&m[566]&m[567]&m[568]&~m[612]))&BiasedRNG[380])|(((m[565]&~m[566]&~m[567]&~m[568]&m[612])|(~m[565]&m[566]&~m[567]&~m[568]&m[612])|(~m[565]&~m[566]&m[567]&~m[568]&m[612])|(m[565]&m[566]&~m[567]&m[568]&m[612])|(m[565]&~m[566]&m[567]&m[568]&m[612])|(~m[565]&m[566]&m[567]&m[568]&m[612]))&~BiasedRNG[380])|((m[565]&m[566]&~m[567]&~m[568]&~m[612])|(m[565]&~m[566]&m[567]&~m[568]&~m[612])|(~m[565]&m[566]&m[567]&~m[568]&~m[612])|(m[565]&m[566]&m[567]&~m[568]&~m[612])|(m[565]&m[566]&m[567]&m[568]&~m[612])|(m[565]&m[566]&~m[567]&~m[568]&m[612])|(m[565]&~m[566]&m[567]&~m[568]&m[612])|(~m[565]&m[566]&m[567]&~m[568]&m[612])|(m[565]&m[566]&m[567]&~m[568]&m[612])|(m[565]&m[566]&m[567]&m[568]&m[612]));
    m[574] = (((m[570]&~m[571]&~m[572]&~m[573]&~m[617])|(~m[570]&m[571]&~m[572]&~m[573]&~m[617])|(~m[570]&~m[571]&m[572]&~m[573]&~m[617])|(m[570]&m[571]&~m[572]&m[573]&~m[617])|(m[570]&~m[571]&m[572]&m[573]&~m[617])|(~m[570]&m[571]&m[572]&m[573]&~m[617]))&BiasedRNG[381])|(((m[570]&~m[571]&~m[572]&~m[573]&m[617])|(~m[570]&m[571]&~m[572]&~m[573]&m[617])|(~m[570]&~m[571]&m[572]&~m[573]&m[617])|(m[570]&m[571]&~m[572]&m[573]&m[617])|(m[570]&~m[571]&m[572]&m[573]&m[617])|(~m[570]&m[571]&m[572]&m[573]&m[617]))&~BiasedRNG[381])|((m[570]&m[571]&~m[572]&~m[573]&~m[617])|(m[570]&~m[571]&m[572]&~m[573]&~m[617])|(~m[570]&m[571]&m[572]&~m[573]&~m[617])|(m[570]&m[571]&m[572]&~m[573]&~m[617])|(m[570]&m[571]&m[572]&m[573]&~m[617])|(m[570]&m[571]&~m[572]&~m[573]&m[617])|(m[570]&~m[571]&m[572]&~m[573]&m[617])|(~m[570]&m[571]&m[572]&~m[573]&m[617])|(m[570]&m[571]&m[572]&~m[573]&m[617])|(m[570]&m[571]&m[572]&m[573]&m[617]));
    m[579] = (((m[575]&~m[576]&~m[577]&~m[578]&~m[622])|(~m[575]&m[576]&~m[577]&~m[578]&~m[622])|(~m[575]&~m[576]&m[577]&~m[578]&~m[622])|(m[575]&m[576]&~m[577]&m[578]&~m[622])|(m[575]&~m[576]&m[577]&m[578]&~m[622])|(~m[575]&m[576]&m[577]&m[578]&~m[622]))&BiasedRNG[382])|(((m[575]&~m[576]&~m[577]&~m[578]&m[622])|(~m[575]&m[576]&~m[577]&~m[578]&m[622])|(~m[575]&~m[576]&m[577]&~m[578]&m[622])|(m[575]&m[576]&~m[577]&m[578]&m[622])|(m[575]&~m[576]&m[577]&m[578]&m[622])|(~m[575]&m[576]&m[577]&m[578]&m[622]))&~BiasedRNG[382])|((m[575]&m[576]&~m[577]&~m[578]&~m[622])|(m[575]&~m[576]&m[577]&~m[578]&~m[622])|(~m[575]&m[576]&m[577]&~m[578]&~m[622])|(m[575]&m[576]&m[577]&~m[578]&~m[622])|(m[575]&m[576]&m[577]&m[578]&~m[622])|(m[575]&m[576]&~m[577]&~m[578]&m[622])|(m[575]&~m[576]&m[577]&~m[578]&m[622])|(~m[575]&m[576]&m[577]&~m[578]&m[622])|(m[575]&m[576]&m[577]&~m[578]&m[622])|(m[575]&m[576]&m[577]&m[578]&m[622]));
    m[584] = (((m[580]&~m[581]&~m[582]&~m[583]&~m[627])|(~m[580]&m[581]&~m[582]&~m[583]&~m[627])|(~m[580]&~m[581]&m[582]&~m[583]&~m[627])|(m[580]&m[581]&~m[582]&m[583]&~m[627])|(m[580]&~m[581]&m[582]&m[583]&~m[627])|(~m[580]&m[581]&m[582]&m[583]&~m[627]))&BiasedRNG[383])|(((m[580]&~m[581]&~m[582]&~m[583]&m[627])|(~m[580]&m[581]&~m[582]&~m[583]&m[627])|(~m[580]&~m[581]&m[582]&~m[583]&m[627])|(m[580]&m[581]&~m[582]&m[583]&m[627])|(m[580]&~m[581]&m[582]&m[583]&m[627])|(~m[580]&m[581]&m[582]&m[583]&m[627]))&~BiasedRNG[383])|((m[580]&m[581]&~m[582]&~m[583]&~m[627])|(m[580]&~m[581]&m[582]&~m[583]&~m[627])|(~m[580]&m[581]&m[582]&~m[583]&~m[627])|(m[580]&m[581]&m[582]&~m[583]&~m[627])|(m[580]&m[581]&m[582]&m[583]&~m[627])|(m[580]&m[581]&~m[582]&~m[583]&m[627])|(m[580]&~m[581]&m[582]&~m[583]&m[627])|(~m[580]&m[581]&m[582]&~m[583]&m[627])|(m[580]&m[581]&m[582]&~m[583]&m[627])|(m[580]&m[581]&m[582]&m[583]&m[627]));
    m[589] = (((m[585]&~m[586]&~m[587]&~m[588]&~m[630])|(~m[585]&m[586]&~m[587]&~m[588]&~m[630])|(~m[585]&~m[586]&m[587]&~m[588]&~m[630])|(m[585]&m[586]&~m[587]&m[588]&~m[630])|(m[585]&~m[586]&m[587]&m[588]&~m[630])|(~m[585]&m[586]&m[587]&m[588]&~m[630]))&BiasedRNG[384])|(((m[585]&~m[586]&~m[587]&~m[588]&m[630])|(~m[585]&m[586]&~m[587]&~m[588]&m[630])|(~m[585]&~m[586]&m[587]&~m[588]&m[630])|(m[585]&m[586]&~m[587]&m[588]&m[630])|(m[585]&~m[586]&m[587]&m[588]&m[630])|(~m[585]&m[586]&m[587]&m[588]&m[630]))&~BiasedRNG[384])|((m[585]&m[586]&~m[587]&~m[588]&~m[630])|(m[585]&~m[586]&m[587]&~m[588]&~m[630])|(~m[585]&m[586]&m[587]&~m[588]&~m[630])|(m[585]&m[586]&m[587]&~m[588]&~m[630])|(m[585]&m[586]&m[587]&m[588]&~m[630])|(m[585]&m[586]&~m[587]&~m[588]&m[630])|(m[585]&~m[586]&m[587]&~m[588]&m[630])|(~m[585]&m[586]&m[587]&~m[588]&m[630])|(m[585]&m[586]&m[587]&~m[588]&m[630])|(m[585]&m[586]&m[587]&m[588]&m[630]));
    m[594] = (((m[590]&~m[591]&~m[592]&~m[593]&~m[632])|(~m[590]&m[591]&~m[592]&~m[593]&~m[632])|(~m[590]&~m[591]&m[592]&~m[593]&~m[632])|(m[590]&m[591]&~m[592]&m[593]&~m[632])|(m[590]&~m[591]&m[592]&m[593]&~m[632])|(~m[590]&m[591]&m[592]&m[593]&~m[632]))&BiasedRNG[385])|(((m[590]&~m[591]&~m[592]&~m[593]&m[632])|(~m[590]&m[591]&~m[592]&~m[593]&m[632])|(~m[590]&~m[591]&m[592]&~m[593]&m[632])|(m[590]&m[591]&~m[592]&m[593]&m[632])|(m[590]&~m[591]&m[592]&m[593]&m[632])|(~m[590]&m[591]&m[592]&m[593]&m[632]))&~BiasedRNG[385])|((m[590]&m[591]&~m[592]&~m[593]&~m[632])|(m[590]&~m[591]&m[592]&~m[593]&~m[632])|(~m[590]&m[591]&m[592]&~m[593]&~m[632])|(m[590]&m[591]&m[592]&~m[593]&~m[632])|(m[590]&m[591]&m[592]&m[593]&~m[632])|(m[590]&m[591]&~m[592]&~m[593]&m[632])|(m[590]&~m[591]&m[592]&~m[593]&m[632])|(~m[590]&m[591]&m[592]&~m[593]&m[632])|(m[590]&m[591]&m[592]&~m[593]&m[632])|(m[590]&m[591]&m[592]&m[593]&m[632]));
    m[599] = (((m[595]&~m[596]&~m[597]&~m[598]&~m[637])|(~m[595]&m[596]&~m[597]&~m[598]&~m[637])|(~m[595]&~m[596]&m[597]&~m[598]&~m[637])|(m[595]&m[596]&~m[597]&m[598]&~m[637])|(m[595]&~m[596]&m[597]&m[598]&~m[637])|(~m[595]&m[596]&m[597]&m[598]&~m[637]))&BiasedRNG[386])|(((m[595]&~m[596]&~m[597]&~m[598]&m[637])|(~m[595]&m[596]&~m[597]&~m[598]&m[637])|(~m[595]&~m[596]&m[597]&~m[598]&m[637])|(m[595]&m[596]&~m[597]&m[598]&m[637])|(m[595]&~m[596]&m[597]&m[598]&m[637])|(~m[595]&m[596]&m[597]&m[598]&m[637]))&~BiasedRNG[386])|((m[595]&m[596]&~m[597]&~m[598]&~m[637])|(m[595]&~m[596]&m[597]&~m[598]&~m[637])|(~m[595]&m[596]&m[597]&~m[598]&~m[637])|(m[595]&m[596]&m[597]&~m[598]&~m[637])|(m[595]&m[596]&m[597]&m[598]&~m[637])|(m[595]&m[596]&~m[597]&~m[598]&m[637])|(m[595]&~m[596]&m[597]&~m[598]&m[637])|(~m[595]&m[596]&m[597]&~m[598]&m[637])|(m[595]&m[596]&m[597]&~m[598]&m[637])|(m[595]&m[596]&m[597]&m[598]&m[637]));
    m[604] = (((m[600]&~m[601]&~m[602]&~m[603]&~m[642])|(~m[600]&m[601]&~m[602]&~m[603]&~m[642])|(~m[600]&~m[601]&m[602]&~m[603]&~m[642])|(m[600]&m[601]&~m[602]&m[603]&~m[642])|(m[600]&~m[601]&m[602]&m[603]&~m[642])|(~m[600]&m[601]&m[602]&m[603]&~m[642]))&BiasedRNG[387])|(((m[600]&~m[601]&~m[602]&~m[603]&m[642])|(~m[600]&m[601]&~m[602]&~m[603]&m[642])|(~m[600]&~m[601]&m[602]&~m[603]&m[642])|(m[600]&m[601]&~m[602]&m[603]&m[642])|(m[600]&~m[601]&m[602]&m[603]&m[642])|(~m[600]&m[601]&m[602]&m[603]&m[642]))&~BiasedRNG[387])|((m[600]&m[601]&~m[602]&~m[603]&~m[642])|(m[600]&~m[601]&m[602]&~m[603]&~m[642])|(~m[600]&m[601]&m[602]&~m[603]&~m[642])|(m[600]&m[601]&m[602]&~m[603]&~m[642])|(m[600]&m[601]&m[602]&m[603]&~m[642])|(m[600]&m[601]&~m[602]&~m[603]&m[642])|(m[600]&~m[601]&m[602]&~m[603]&m[642])|(~m[600]&m[601]&m[602]&~m[603]&m[642])|(m[600]&m[601]&m[602]&~m[603]&m[642])|(m[600]&m[601]&m[602]&m[603]&m[642]));
    m[609] = (((m[605]&~m[606]&~m[607]&~m[608]&~m[647])|(~m[605]&m[606]&~m[607]&~m[608]&~m[647])|(~m[605]&~m[606]&m[607]&~m[608]&~m[647])|(m[605]&m[606]&~m[607]&m[608]&~m[647])|(m[605]&~m[606]&m[607]&m[608]&~m[647])|(~m[605]&m[606]&m[607]&m[608]&~m[647]))&BiasedRNG[388])|(((m[605]&~m[606]&~m[607]&~m[608]&m[647])|(~m[605]&m[606]&~m[607]&~m[608]&m[647])|(~m[605]&~m[606]&m[607]&~m[608]&m[647])|(m[605]&m[606]&~m[607]&m[608]&m[647])|(m[605]&~m[606]&m[607]&m[608]&m[647])|(~m[605]&m[606]&m[607]&m[608]&m[647]))&~BiasedRNG[388])|((m[605]&m[606]&~m[607]&~m[608]&~m[647])|(m[605]&~m[606]&m[607]&~m[608]&~m[647])|(~m[605]&m[606]&m[607]&~m[608]&~m[647])|(m[605]&m[606]&m[607]&~m[608]&~m[647])|(m[605]&m[606]&m[607]&m[608]&~m[647])|(m[605]&m[606]&~m[607]&~m[608]&m[647])|(m[605]&~m[606]&m[607]&~m[608]&m[647])|(~m[605]&m[606]&m[607]&~m[608]&m[647])|(m[605]&m[606]&m[607]&~m[608]&m[647])|(m[605]&m[606]&m[607]&m[608]&m[647]));
    m[614] = (((m[610]&~m[611]&~m[612]&~m[613]&~m[652])|(~m[610]&m[611]&~m[612]&~m[613]&~m[652])|(~m[610]&~m[611]&m[612]&~m[613]&~m[652])|(m[610]&m[611]&~m[612]&m[613]&~m[652])|(m[610]&~m[611]&m[612]&m[613]&~m[652])|(~m[610]&m[611]&m[612]&m[613]&~m[652]))&BiasedRNG[389])|(((m[610]&~m[611]&~m[612]&~m[613]&m[652])|(~m[610]&m[611]&~m[612]&~m[613]&m[652])|(~m[610]&~m[611]&m[612]&~m[613]&m[652])|(m[610]&m[611]&~m[612]&m[613]&m[652])|(m[610]&~m[611]&m[612]&m[613]&m[652])|(~m[610]&m[611]&m[612]&m[613]&m[652]))&~BiasedRNG[389])|((m[610]&m[611]&~m[612]&~m[613]&~m[652])|(m[610]&~m[611]&m[612]&~m[613]&~m[652])|(~m[610]&m[611]&m[612]&~m[613]&~m[652])|(m[610]&m[611]&m[612]&~m[613]&~m[652])|(m[610]&m[611]&m[612]&m[613]&~m[652])|(m[610]&m[611]&~m[612]&~m[613]&m[652])|(m[610]&~m[611]&m[612]&~m[613]&m[652])|(~m[610]&m[611]&m[612]&~m[613]&m[652])|(m[610]&m[611]&m[612]&~m[613]&m[652])|(m[610]&m[611]&m[612]&m[613]&m[652]));
    m[619] = (((m[615]&~m[616]&~m[617]&~m[618]&~m[657])|(~m[615]&m[616]&~m[617]&~m[618]&~m[657])|(~m[615]&~m[616]&m[617]&~m[618]&~m[657])|(m[615]&m[616]&~m[617]&m[618]&~m[657])|(m[615]&~m[616]&m[617]&m[618]&~m[657])|(~m[615]&m[616]&m[617]&m[618]&~m[657]))&BiasedRNG[390])|(((m[615]&~m[616]&~m[617]&~m[618]&m[657])|(~m[615]&m[616]&~m[617]&~m[618]&m[657])|(~m[615]&~m[616]&m[617]&~m[618]&m[657])|(m[615]&m[616]&~m[617]&m[618]&m[657])|(m[615]&~m[616]&m[617]&m[618]&m[657])|(~m[615]&m[616]&m[617]&m[618]&m[657]))&~BiasedRNG[390])|((m[615]&m[616]&~m[617]&~m[618]&~m[657])|(m[615]&~m[616]&m[617]&~m[618]&~m[657])|(~m[615]&m[616]&m[617]&~m[618]&~m[657])|(m[615]&m[616]&m[617]&~m[618]&~m[657])|(m[615]&m[616]&m[617]&m[618]&~m[657])|(m[615]&m[616]&~m[617]&~m[618]&m[657])|(m[615]&~m[616]&m[617]&~m[618]&m[657])|(~m[615]&m[616]&m[617]&~m[618]&m[657])|(m[615]&m[616]&m[617]&~m[618]&m[657])|(m[615]&m[616]&m[617]&m[618]&m[657]));
    m[624] = (((m[620]&~m[621]&~m[622]&~m[623]&~m[662])|(~m[620]&m[621]&~m[622]&~m[623]&~m[662])|(~m[620]&~m[621]&m[622]&~m[623]&~m[662])|(m[620]&m[621]&~m[622]&m[623]&~m[662])|(m[620]&~m[621]&m[622]&m[623]&~m[662])|(~m[620]&m[621]&m[622]&m[623]&~m[662]))&BiasedRNG[391])|(((m[620]&~m[621]&~m[622]&~m[623]&m[662])|(~m[620]&m[621]&~m[622]&~m[623]&m[662])|(~m[620]&~m[621]&m[622]&~m[623]&m[662])|(m[620]&m[621]&~m[622]&m[623]&m[662])|(m[620]&~m[621]&m[622]&m[623]&m[662])|(~m[620]&m[621]&m[622]&m[623]&m[662]))&~BiasedRNG[391])|((m[620]&m[621]&~m[622]&~m[623]&~m[662])|(m[620]&~m[621]&m[622]&~m[623]&~m[662])|(~m[620]&m[621]&m[622]&~m[623]&~m[662])|(m[620]&m[621]&m[622]&~m[623]&~m[662])|(m[620]&m[621]&m[622]&m[623]&~m[662])|(m[620]&m[621]&~m[622]&~m[623]&m[662])|(m[620]&~m[621]&m[622]&~m[623]&m[662])|(~m[620]&m[621]&m[622]&~m[623]&m[662])|(m[620]&m[621]&m[622]&~m[623]&m[662])|(m[620]&m[621]&m[622]&m[623]&m[662]));
    m[629] = (((m[625]&~m[626]&~m[627]&~m[628]&~m[667])|(~m[625]&m[626]&~m[627]&~m[628]&~m[667])|(~m[625]&~m[626]&m[627]&~m[628]&~m[667])|(m[625]&m[626]&~m[627]&m[628]&~m[667])|(m[625]&~m[626]&m[627]&m[628]&~m[667])|(~m[625]&m[626]&m[627]&m[628]&~m[667]))&BiasedRNG[392])|(((m[625]&~m[626]&~m[627]&~m[628]&m[667])|(~m[625]&m[626]&~m[627]&~m[628]&m[667])|(~m[625]&~m[626]&m[627]&~m[628]&m[667])|(m[625]&m[626]&~m[627]&m[628]&m[667])|(m[625]&~m[626]&m[627]&m[628]&m[667])|(~m[625]&m[626]&m[627]&m[628]&m[667]))&~BiasedRNG[392])|((m[625]&m[626]&~m[627]&~m[628]&~m[667])|(m[625]&~m[626]&m[627]&~m[628]&~m[667])|(~m[625]&m[626]&m[627]&~m[628]&~m[667])|(m[625]&m[626]&m[627]&~m[628]&~m[667])|(m[625]&m[626]&m[627]&m[628]&~m[667])|(m[625]&m[626]&~m[627]&~m[628]&m[667])|(m[625]&~m[626]&m[627]&~m[628]&m[667])|(~m[625]&m[626]&m[627]&~m[628]&m[667])|(m[625]&m[626]&m[627]&~m[628]&m[667])|(m[625]&m[626]&m[627]&m[628]&m[667]));
    m[634] = (((m[630]&~m[631]&~m[632]&~m[633]&~m[670])|(~m[630]&m[631]&~m[632]&~m[633]&~m[670])|(~m[630]&~m[631]&m[632]&~m[633]&~m[670])|(m[630]&m[631]&~m[632]&m[633]&~m[670])|(m[630]&~m[631]&m[632]&m[633]&~m[670])|(~m[630]&m[631]&m[632]&m[633]&~m[670]))&BiasedRNG[393])|(((m[630]&~m[631]&~m[632]&~m[633]&m[670])|(~m[630]&m[631]&~m[632]&~m[633]&m[670])|(~m[630]&~m[631]&m[632]&~m[633]&m[670])|(m[630]&m[631]&~m[632]&m[633]&m[670])|(m[630]&~m[631]&m[632]&m[633]&m[670])|(~m[630]&m[631]&m[632]&m[633]&m[670]))&~BiasedRNG[393])|((m[630]&m[631]&~m[632]&~m[633]&~m[670])|(m[630]&~m[631]&m[632]&~m[633]&~m[670])|(~m[630]&m[631]&m[632]&~m[633]&~m[670])|(m[630]&m[631]&m[632]&~m[633]&~m[670])|(m[630]&m[631]&m[632]&m[633]&~m[670])|(m[630]&m[631]&~m[632]&~m[633]&m[670])|(m[630]&~m[631]&m[632]&~m[633]&m[670])|(~m[630]&m[631]&m[632]&~m[633]&m[670])|(m[630]&m[631]&m[632]&~m[633]&m[670])|(m[630]&m[631]&m[632]&m[633]&m[670]));
    m[639] = (((m[635]&~m[636]&~m[637]&~m[638]&~m[672])|(~m[635]&m[636]&~m[637]&~m[638]&~m[672])|(~m[635]&~m[636]&m[637]&~m[638]&~m[672])|(m[635]&m[636]&~m[637]&m[638]&~m[672])|(m[635]&~m[636]&m[637]&m[638]&~m[672])|(~m[635]&m[636]&m[637]&m[638]&~m[672]))&BiasedRNG[394])|(((m[635]&~m[636]&~m[637]&~m[638]&m[672])|(~m[635]&m[636]&~m[637]&~m[638]&m[672])|(~m[635]&~m[636]&m[637]&~m[638]&m[672])|(m[635]&m[636]&~m[637]&m[638]&m[672])|(m[635]&~m[636]&m[637]&m[638]&m[672])|(~m[635]&m[636]&m[637]&m[638]&m[672]))&~BiasedRNG[394])|((m[635]&m[636]&~m[637]&~m[638]&~m[672])|(m[635]&~m[636]&m[637]&~m[638]&~m[672])|(~m[635]&m[636]&m[637]&~m[638]&~m[672])|(m[635]&m[636]&m[637]&~m[638]&~m[672])|(m[635]&m[636]&m[637]&m[638]&~m[672])|(m[635]&m[636]&~m[637]&~m[638]&m[672])|(m[635]&~m[636]&m[637]&~m[638]&m[672])|(~m[635]&m[636]&m[637]&~m[638]&m[672])|(m[635]&m[636]&m[637]&~m[638]&m[672])|(m[635]&m[636]&m[637]&m[638]&m[672]));
    m[644] = (((m[640]&~m[641]&~m[642]&~m[643]&~m[677])|(~m[640]&m[641]&~m[642]&~m[643]&~m[677])|(~m[640]&~m[641]&m[642]&~m[643]&~m[677])|(m[640]&m[641]&~m[642]&m[643]&~m[677])|(m[640]&~m[641]&m[642]&m[643]&~m[677])|(~m[640]&m[641]&m[642]&m[643]&~m[677]))&BiasedRNG[395])|(((m[640]&~m[641]&~m[642]&~m[643]&m[677])|(~m[640]&m[641]&~m[642]&~m[643]&m[677])|(~m[640]&~m[641]&m[642]&~m[643]&m[677])|(m[640]&m[641]&~m[642]&m[643]&m[677])|(m[640]&~m[641]&m[642]&m[643]&m[677])|(~m[640]&m[641]&m[642]&m[643]&m[677]))&~BiasedRNG[395])|((m[640]&m[641]&~m[642]&~m[643]&~m[677])|(m[640]&~m[641]&m[642]&~m[643]&~m[677])|(~m[640]&m[641]&m[642]&~m[643]&~m[677])|(m[640]&m[641]&m[642]&~m[643]&~m[677])|(m[640]&m[641]&m[642]&m[643]&~m[677])|(m[640]&m[641]&~m[642]&~m[643]&m[677])|(m[640]&~m[641]&m[642]&~m[643]&m[677])|(~m[640]&m[641]&m[642]&~m[643]&m[677])|(m[640]&m[641]&m[642]&~m[643]&m[677])|(m[640]&m[641]&m[642]&m[643]&m[677]));
    m[649] = (((m[645]&~m[646]&~m[647]&~m[648]&~m[682])|(~m[645]&m[646]&~m[647]&~m[648]&~m[682])|(~m[645]&~m[646]&m[647]&~m[648]&~m[682])|(m[645]&m[646]&~m[647]&m[648]&~m[682])|(m[645]&~m[646]&m[647]&m[648]&~m[682])|(~m[645]&m[646]&m[647]&m[648]&~m[682]))&BiasedRNG[396])|(((m[645]&~m[646]&~m[647]&~m[648]&m[682])|(~m[645]&m[646]&~m[647]&~m[648]&m[682])|(~m[645]&~m[646]&m[647]&~m[648]&m[682])|(m[645]&m[646]&~m[647]&m[648]&m[682])|(m[645]&~m[646]&m[647]&m[648]&m[682])|(~m[645]&m[646]&m[647]&m[648]&m[682]))&~BiasedRNG[396])|((m[645]&m[646]&~m[647]&~m[648]&~m[682])|(m[645]&~m[646]&m[647]&~m[648]&~m[682])|(~m[645]&m[646]&m[647]&~m[648]&~m[682])|(m[645]&m[646]&m[647]&~m[648]&~m[682])|(m[645]&m[646]&m[647]&m[648]&~m[682])|(m[645]&m[646]&~m[647]&~m[648]&m[682])|(m[645]&~m[646]&m[647]&~m[648]&m[682])|(~m[645]&m[646]&m[647]&~m[648]&m[682])|(m[645]&m[646]&m[647]&~m[648]&m[682])|(m[645]&m[646]&m[647]&m[648]&m[682]));
    m[654] = (((m[650]&~m[651]&~m[652]&~m[653]&~m[687])|(~m[650]&m[651]&~m[652]&~m[653]&~m[687])|(~m[650]&~m[651]&m[652]&~m[653]&~m[687])|(m[650]&m[651]&~m[652]&m[653]&~m[687])|(m[650]&~m[651]&m[652]&m[653]&~m[687])|(~m[650]&m[651]&m[652]&m[653]&~m[687]))&BiasedRNG[397])|(((m[650]&~m[651]&~m[652]&~m[653]&m[687])|(~m[650]&m[651]&~m[652]&~m[653]&m[687])|(~m[650]&~m[651]&m[652]&~m[653]&m[687])|(m[650]&m[651]&~m[652]&m[653]&m[687])|(m[650]&~m[651]&m[652]&m[653]&m[687])|(~m[650]&m[651]&m[652]&m[653]&m[687]))&~BiasedRNG[397])|((m[650]&m[651]&~m[652]&~m[653]&~m[687])|(m[650]&~m[651]&m[652]&~m[653]&~m[687])|(~m[650]&m[651]&m[652]&~m[653]&~m[687])|(m[650]&m[651]&m[652]&~m[653]&~m[687])|(m[650]&m[651]&m[652]&m[653]&~m[687])|(m[650]&m[651]&~m[652]&~m[653]&m[687])|(m[650]&~m[651]&m[652]&~m[653]&m[687])|(~m[650]&m[651]&m[652]&~m[653]&m[687])|(m[650]&m[651]&m[652]&~m[653]&m[687])|(m[650]&m[651]&m[652]&m[653]&m[687]));
    m[659] = (((m[655]&~m[656]&~m[657]&~m[658]&~m[692])|(~m[655]&m[656]&~m[657]&~m[658]&~m[692])|(~m[655]&~m[656]&m[657]&~m[658]&~m[692])|(m[655]&m[656]&~m[657]&m[658]&~m[692])|(m[655]&~m[656]&m[657]&m[658]&~m[692])|(~m[655]&m[656]&m[657]&m[658]&~m[692]))&BiasedRNG[398])|(((m[655]&~m[656]&~m[657]&~m[658]&m[692])|(~m[655]&m[656]&~m[657]&~m[658]&m[692])|(~m[655]&~m[656]&m[657]&~m[658]&m[692])|(m[655]&m[656]&~m[657]&m[658]&m[692])|(m[655]&~m[656]&m[657]&m[658]&m[692])|(~m[655]&m[656]&m[657]&m[658]&m[692]))&~BiasedRNG[398])|((m[655]&m[656]&~m[657]&~m[658]&~m[692])|(m[655]&~m[656]&m[657]&~m[658]&~m[692])|(~m[655]&m[656]&m[657]&~m[658]&~m[692])|(m[655]&m[656]&m[657]&~m[658]&~m[692])|(m[655]&m[656]&m[657]&m[658]&~m[692])|(m[655]&m[656]&~m[657]&~m[658]&m[692])|(m[655]&~m[656]&m[657]&~m[658]&m[692])|(~m[655]&m[656]&m[657]&~m[658]&m[692])|(m[655]&m[656]&m[657]&~m[658]&m[692])|(m[655]&m[656]&m[657]&m[658]&m[692]));
    m[664] = (((m[660]&~m[661]&~m[662]&~m[663]&~m[697])|(~m[660]&m[661]&~m[662]&~m[663]&~m[697])|(~m[660]&~m[661]&m[662]&~m[663]&~m[697])|(m[660]&m[661]&~m[662]&m[663]&~m[697])|(m[660]&~m[661]&m[662]&m[663]&~m[697])|(~m[660]&m[661]&m[662]&m[663]&~m[697]))&BiasedRNG[399])|(((m[660]&~m[661]&~m[662]&~m[663]&m[697])|(~m[660]&m[661]&~m[662]&~m[663]&m[697])|(~m[660]&~m[661]&m[662]&~m[663]&m[697])|(m[660]&m[661]&~m[662]&m[663]&m[697])|(m[660]&~m[661]&m[662]&m[663]&m[697])|(~m[660]&m[661]&m[662]&m[663]&m[697]))&~BiasedRNG[399])|((m[660]&m[661]&~m[662]&~m[663]&~m[697])|(m[660]&~m[661]&m[662]&~m[663]&~m[697])|(~m[660]&m[661]&m[662]&~m[663]&~m[697])|(m[660]&m[661]&m[662]&~m[663]&~m[697])|(m[660]&m[661]&m[662]&m[663]&~m[697])|(m[660]&m[661]&~m[662]&~m[663]&m[697])|(m[660]&~m[661]&m[662]&~m[663]&m[697])|(~m[660]&m[661]&m[662]&~m[663]&m[697])|(m[660]&m[661]&m[662]&~m[663]&m[697])|(m[660]&m[661]&m[662]&m[663]&m[697]));
    m[669] = (((m[665]&~m[666]&~m[667]&~m[668]&~m[702])|(~m[665]&m[666]&~m[667]&~m[668]&~m[702])|(~m[665]&~m[666]&m[667]&~m[668]&~m[702])|(m[665]&m[666]&~m[667]&m[668]&~m[702])|(m[665]&~m[666]&m[667]&m[668]&~m[702])|(~m[665]&m[666]&m[667]&m[668]&~m[702]))&BiasedRNG[400])|(((m[665]&~m[666]&~m[667]&~m[668]&m[702])|(~m[665]&m[666]&~m[667]&~m[668]&m[702])|(~m[665]&~m[666]&m[667]&~m[668]&m[702])|(m[665]&m[666]&~m[667]&m[668]&m[702])|(m[665]&~m[666]&m[667]&m[668]&m[702])|(~m[665]&m[666]&m[667]&m[668]&m[702]))&~BiasedRNG[400])|((m[665]&m[666]&~m[667]&~m[668]&~m[702])|(m[665]&~m[666]&m[667]&~m[668]&~m[702])|(~m[665]&m[666]&m[667]&~m[668]&~m[702])|(m[665]&m[666]&m[667]&~m[668]&~m[702])|(m[665]&m[666]&m[667]&m[668]&~m[702])|(m[665]&m[666]&~m[667]&~m[668]&m[702])|(m[665]&~m[666]&m[667]&~m[668]&m[702])|(~m[665]&m[666]&m[667]&~m[668]&m[702])|(m[665]&m[666]&m[667]&~m[668]&m[702])|(m[665]&m[666]&m[667]&m[668]&m[702]));
    m[674] = (((m[670]&~m[671]&~m[672]&~m[673]&~m[705])|(~m[670]&m[671]&~m[672]&~m[673]&~m[705])|(~m[670]&~m[671]&m[672]&~m[673]&~m[705])|(m[670]&m[671]&~m[672]&m[673]&~m[705])|(m[670]&~m[671]&m[672]&m[673]&~m[705])|(~m[670]&m[671]&m[672]&m[673]&~m[705]))&BiasedRNG[401])|(((m[670]&~m[671]&~m[672]&~m[673]&m[705])|(~m[670]&m[671]&~m[672]&~m[673]&m[705])|(~m[670]&~m[671]&m[672]&~m[673]&m[705])|(m[670]&m[671]&~m[672]&m[673]&m[705])|(m[670]&~m[671]&m[672]&m[673]&m[705])|(~m[670]&m[671]&m[672]&m[673]&m[705]))&~BiasedRNG[401])|((m[670]&m[671]&~m[672]&~m[673]&~m[705])|(m[670]&~m[671]&m[672]&~m[673]&~m[705])|(~m[670]&m[671]&m[672]&~m[673]&~m[705])|(m[670]&m[671]&m[672]&~m[673]&~m[705])|(m[670]&m[671]&m[672]&m[673]&~m[705])|(m[670]&m[671]&~m[672]&~m[673]&m[705])|(m[670]&~m[671]&m[672]&~m[673]&m[705])|(~m[670]&m[671]&m[672]&~m[673]&m[705])|(m[670]&m[671]&m[672]&~m[673]&m[705])|(m[670]&m[671]&m[672]&m[673]&m[705]));
    m[679] = (((m[675]&~m[676]&~m[677]&~m[678]&~m[707])|(~m[675]&m[676]&~m[677]&~m[678]&~m[707])|(~m[675]&~m[676]&m[677]&~m[678]&~m[707])|(m[675]&m[676]&~m[677]&m[678]&~m[707])|(m[675]&~m[676]&m[677]&m[678]&~m[707])|(~m[675]&m[676]&m[677]&m[678]&~m[707]))&BiasedRNG[402])|(((m[675]&~m[676]&~m[677]&~m[678]&m[707])|(~m[675]&m[676]&~m[677]&~m[678]&m[707])|(~m[675]&~m[676]&m[677]&~m[678]&m[707])|(m[675]&m[676]&~m[677]&m[678]&m[707])|(m[675]&~m[676]&m[677]&m[678]&m[707])|(~m[675]&m[676]&m[677]&m[678]&m[707]))&~BiasedRNG[402])|((m[675]&m[676]&~m[677]&~m[678]&~m[707])|(m[675]&~m[676]&m[677]&~m[678]&~m[707])|(~m[675]&m[676]&m[677]&~m[678]&~m[707])|(m[675]&m[676]&m[677]&~m[678]&~m[707])|(m[675]&m[676]&m[677]&m[678]&~m[707])|(m[675]&m[676]&~m[677]&~m[678]&m[707])|(m[675]&~m[676]&m[677]&~m[678]&m[707])|(~m[675]&m[676]&m[677]&~m[678]&m[707])|(m[675]&m[676]&m[677]&~m[678]&m[707])|(m[675]&m[676]&m[677]&m[678]&m[707]));
    m[684] = (((m[680]&~m[681]&~m[682]&~m[683]&~m[712])|(~m[680]&m[681]&~m[682]&~m[683]&~m[712])|(~m[680]&~m[681]&m[682]&~m[683]&~m[712])|(m[680]&m[681]&~m[682]&m[683]&~m[712])|(m[680]&~m[681]&m[682]&m[683]&~m[712])|(~m[680]&m[681]&m[682]&m[683]&~m[712]))&BiasedRNG[403])|(((m[680]&~m[681]&~m[682]&~m[683]&m[712])|(~m[680]&m[681]&~m[682]&~m[683]&m[712])|(~m[680]&~m[681]&m[682]&~m[683]&m[712])|(m[680]&m[681]&~m[682]&m[683]&m[712])|(m[680]&~m[681]&m[682]&m[683]&m[712])|(~m[680]&m[681]&m[682]&m[683]&m[712]))&~BiasedRNG[403])|((m[680]&m[681]&~m[682]&~m[683]&~m[712])|(m[680]&~m[681]&m[682]&~m[683]&~m[712])|(~m[680]&m[681]&m[682]&~m[683]&~m[712])|(m[680]&m[681]&m[682]&~m[683]&~m[712])|(m[680]&m[681]&m[682]&m[683]&~m[712])|(m[680]&m[681]&~m[682]&~m[683]&m[712])|(m[680]&~m[681]&m[682]&~m[683]&m[712])|(~m[680]&m[681]&m[682]&~m[683]&m[712])|(m[680]&m[681]&m[682]&~m[683]&m[712])|(m[680]&m[681]&m[682]&m[683]&m[712]));
    m[689] = (((m[685]&~m[686]&~m[687]&~m[688]&~m[717])|(~m[685]&m[686]&~m[687]&~m[688]&~m[717])|(~m[685]&~m[686]&m[687]&~m[688]&~m[717])|(m[685]&m[686]&~m[687]&m[688]&~m[717])|(m[685]&~m[686]&m[687]&m[688]&~m[717])|(~m[685]&m[686]&m[687]&m[688]&~m[717]))&BiasedRNG[404])|(((m[685]&~m[686]&~m[687]&~m[688]&m[717])|(~m[685]&m[686]&~m[687]&~m[688]&m[717])|(~m[685]&~m[686]&m[687]&~m[688]&m[717])|(m[685]&m[686]&~m[687]&m[688]&m[717])|(m[685]&~m[686]&m[687]&m[688]&m[717])|(~m[685]&m[686]&m[687]&m[688]&m[717]))&~BiasedRNG[404])|((m[685]&m[686]&~m[687]&~m[688]&~m[717])|(m[685]&~m[686]&m[687]&~m[688]&~m[717])|(~m[685]&m[686]&m[687]&~m[688]&~m[717])|(m[685]&m[686]&m[687]&~m[688]&~m[717])|(m[685]&m[686]&m[687]&m[688]&~m[717])|(m[685]&m[686]&~m[687]&~m[688]&m[717])|(m[685]&~m[686]&m[687]&~m[688]&m[717])|(~m[685]&m[686]&m[687]&~m[688]&m[717])|(m[685]&m[686]&m[687]&~m[688]&m[717])|(m[685]&m[686]&m[687]&m[688]&m[717]));
    m[694] = (((m[690]&~m[691]&~m[692]&~m[693]&~m[722])|(~m[690]&m[691]&~m[692]&~m[693]&~m[722])|(~m[690]&~m[691]&m[692]&~m[693]&~m[722])|(m[690]&m[691]&~m[692]&m[693]&~m[722])|(m[690]&~m[691]&m[692]&m[693]&~m[722])|(~m[690]&m[691]&m[692]&m[693]&~m[722]))&BiasedRNG[405])|(((m[690]&~m[691]&~m[692]&~m[693]&m[722])|(~m[690]&m[691]&~m[692]&~m[693]&m[722])|(~m[690]&~m[691]&m[692]&~m[693]&m[722])|(m[690]&m[691]&~m[692]&m[693]&m[722])|(m[690]&~m[691]&m[692]&m[693]&m[722])|(~m[690]&m[691]&m[692]&m[693]&m[722]))&~BiasedRNG[405])|((m[690]&m[691]&~m[692]&~m[693]&~m[722])|(m[690]&~m[691]&m[692]&~m[693]&~m[722])|(~m[690]&m[691]&m[692]&~m[693]&~m[722])|(m[690]&m[691]&m[692]&~m[693]&~m[722])|(m[690]&m[691]&m[692]&m[693]&~m[722])|(m[690]&m[691]&~m[692]&~m[693]&m[722])|(m[690]&~m[691]&m[692]&~m[693]&m[722])|(~m[690]&m[691]&m[692]&~m[693]&m[722])|(m[690]&m[691]&m[692]&~m[693]&m[722])|(m[690]&m[691]&m[692]&m[693]&m[722]));
    m[699] = (((m[695]&~m[696]&~m[697]&~m[698]&~m[727])|(~m[695]&m[696]&~m[697]&~m[698]&~m[727])|(~m[695]&~m[696]&m[697]&~m[698]&~m[727])|(m[695]&m[696]&~m[697]&m[698]&~m[727])|(m[695]&~m[696]&m[697]&m[698]&~m[727])|(~m[695]&m[696]&m[697]&m[698]&~m[727]))&BiasedRNG[406])|(((m[695]&~m[696]&~m[697]&~m[698]&m[727])|(~m[695]&m[696]&~m[697]&~m[698]&m[727])|(~m[695]&~m[696]&m[697]&~m[698]&m[727])|(m[695]&m[696]&~m[697]&m[698]&m[727])|(m[695]&~m[696]&m[697]&m[698]&m[727])|(~m[695]&m[696]&m[697]&m[698]&m[727]))&~BiasedRNG[406])|((m[695]&m[696]&~m[697]&~m[698]&~m[727])|(m[695]&~m[696]&m[697]&~m[698]&~m[727])|(~m[695]&m[696]&m[697]&~m[698]&~m[727])|(m[695]&m[696]&m[697]&~m[698]&~m[727])|(m[695]&m[696]&m[697]&m[698]&~m[727])|(m[695]&m[696]&~m[697]&~m[698]&m[727])|(m[695]&~m[696]&m[697]&~m[698]&m[727])|(~m[695]&m[696]&m[697]&~m[698]&m[727])|(m[695]&m[696]&m[697]&~m[698]&m[727])|(m[695]&m[696]&m[697]&m[698]&m[727]));
    m[704] = (((m[700]&~m[701]&~m[702]&~m[703]&~m[732])|(~m[700]&m[701]&~m[702]&~m[703]&~m[732])|(~m[700]&~m[701]&m[702]&~m[703]&~m[732])|(m[700]&m[701]&~m[702]&m[703]&~m[732])|(m[700]&~m[701]&m[702]&m[703]&~m[732])|(~m[700]&m[701]&m[702]&m[703]&~m[732]))&BiasedRNG[407])|(((m[700]&~m[701]&~m[702]&~m[703]&m[732])|(~m[700]&m[701]&~m[702]&~m[703]&m[732])|(~m[700]&~m[701]&m[702]&~m[703]&m[732])|(m[700]&m[701]&~m[702]&m[703]&m[732])|(m[700]&~m[701]&m[702]&m[703]&m[732])|(~m[700]&m[701]&m[702]&m[703]&m[732]))&~BiasedRNG[407])|((m[700]&m[701]&~m[702]&~m[703]&~m[732])|(m[700]&~m[701]&m[702]&~m[703]&~m[732])|(~m[700]&m[701]&m[702]&~m[703]&~m[732])|(m[700]&m[701]&m[702]&~m[703]&~m[732])|(m[700]&m[701]&m[702]&m[703]&~m[732])|(m[700]&m[701]&~m[702]&~m[703]&m[732])|(m[700]&~m[701]&m[702]&~m[703]&m[732])|(~m[700]&m[701]&m[702]&~m[703]&m[732])|(m[700]&m[701]&m[702]&~m[703]&m[732])|(m[700]&m[701]&m[702]&m[703]&m[732]));
    m[709] = (((m[705]&~m[706]&~m[707]&~m[708]&~m[735])|(~m[705]&m[706]&~m[707]&~m[708]&~m[735])|(~m[705]&~m[706]&m[707]&~m[708]&~m[735])|(m[705]&m[706]&~m[707]&m[708]&~m[735])|(m[705]&~m[706]&m[707]&m[708]&~m[735])|(~m[705]&m[706]&m[707]&m[708]&~m[735]))&BiasedRNG[408])|(((m[705]&~m[706]&~m[707]&~m[708]&m[735])|(~m[705]&m[706]&~m[707]&~m[708]&m[735])|(~m[705]&~m[706]&m[707]&~m[708]&m[735])|(m[705]&m[706]&~m[707]&m[708]&m[735])|(m[705]&~m[706]&m[707]&m[708]&m[735])|(~m[705]&m[706]&m[707]&m[708]&m[735]))&~BiasedRNG[408])|((m[705]&m[706]&~m[707]&~m[708]&~m[735])|(m[705]&~m[706]&m[707]&~m[708]&~m[735])|(~m[705]&m[706]&m[707]&~m[708]&~m[735])|(m[705]&m[706]&m[707]&~m[708]&~m[735])|(m[705]&m[706]&m[707]&m[708]&~m[735])|(m[705]&m[706]&~m[707]&~m[708]&m[735])|(m[705]&~m[706]&m[707]&~m[708]&m[735])|(~m[705]&m[706]&m[707]&~m[708]&m[735])|(m[705]&m[706]&m[707]&~m[708]&m[735])|(m[705]&m[706]&m[707]&m[708]&m[735]));
    m[714] = (((m[710]&~m[711]&~m[712]&~m[713]&~m[737])|(~m[710]&m[711]&~m[712]&~m[713]&~m[737])|(~m[710]&~m[711]&m[712]&~m[713]&~m[737])|(m[710]&m[711]&~m[712]&m[713]&~m[737])|(m[710]&~m[711]&m[712]&m[713]&~m[737])|(~m[710]&m[711]&m[712]&m[713]&~m[737]))&BiasedRNG[409])|(((m[710]&~m[711]&~m[712]&~m[713]&m[737])|(~m[710]&m[711]&~m[712]&~m[713]&m[737])|(~m[710]&~m[711]&m[712]&~m[713]&m[737])|(m[710]&m[711]&~m[712]&m[713]&m[737])|(m[710]&~m[711]&m[712]&m[713]&m[737])|(~m[710]&m[711]&m[712]&m[713]&m[737]))&~BiasedRNG[409])|((m[710]&m[711]&~m[712]&~m[713]&~m[737])|(m[710]&~m[711]&m[712]&~m[713]&~m[737])|(~m[710]&m[711]&m[712]&~m[713]&~m[737])|(m[710]&m[711]&m[712]&~m[713]&~m[737])|(m[710]&m[711]&m[712]&m[713]&~m[737])|(m[710]&m[711]&~m[712]&~m[713]&m[737])|(m[710]&~m[711]&m[712]&~m[713]&m[737])|(~m[710]&m[711]&m[712]&~m[713]&m[737])|(m[710]&m[711]&m[712]&~m[713]&m[737])|(m[710]&m[711]&m[712]&m[713]&m[737]));
    m[719] = (((m[715]&~m[716]&~m[717]&~m[718]&~m[742])|(~m[715]&m[716]&~m[717]&~m[718]&~m[742])|(~m[715]&~m[716]&m[717]&~m[718]&~m[742])|(m[715]&m[716]&~m[717]&m[718]&~m[742])|(m[715]&~m[716]&m[717]&m[718]&~m[742])|(~m[715]&m[716]&m[717]&m[718]&~m[742]))&BiasedRNG[410])|(((m[715]&~m[716]&~m[717]&~m[718]&m[742])|(~m[715]&m[716]&~m[717]&~m[718]&m[742])|(~m[715]&~m[716]&m[717]&~m[718]&m[742])|(m[715]&m[716]&~m[717]&m[718]&m[742])|(m[715]&~m[716]&m[717]&m[718]&m[742])|(~m[715]&m[716]&m[717]&m[718]&m[742]))&~BiasedRNG[410])|((m[715]&m[716]&~m[717]&~m[718]&~m[742])|(m[715]&~m[716]&m[717]&~m[718]&~m[742])|(~m[715]&m[716]&m[717]&~m[718]&~m[742])|(m[715]&m[716]&m[717]&~m[718]&~m[742])|(m[715]&m[716]&m[717]&m[718]&~m[742])|(m[715]&m[716]&~m[717]&~m[718]&m[742])|(m[715]&~m[716]&m[717]&~m[718]&m[742])|(~m[715]&m[716]&m[717]&~m[718]&m[742])|(m[715]&m[716]&m[717]&~m[718]&m[742])|(m[715]&m[716]&m[717]&m[718]&m[742]));
    m[724] = (((m[720]&~m[721]&~m[722]&~m[723]&~m[747])|(~m[720]&m[721]&~m[722]&~m[723]&~m[747])|(~m[720]&~m[721]&m[722]&~m[723]&~m[747])|(m[720]&m[721]&~m[722]&m[723]&~m[747])|(m[720]&~m[721]&m[722]&m[723]&~m[747])|(~m[720]&m[721]&m[722]&m[723]&~m[747]))&BiasedRNG[411])|(((m[720]&~m[721]&~m[722]&~m[723]&m[747])|(~m[720]&m[721]&~m[722]&~m[723]&m[747])|(~m[720]&~m[721]&m[722]&~m[723]&m[747])|(m[720]&m[721]&~m[722]&m[723]&m[747])|(m[720]&~m[721]&m[722]&m[723]&m[747])|(~m[720]&m[721]&m[722]&m[723]&m[747]))&~BiasedRNG[411])|((m[720]&m[721]&~m[722]&~m[723]&~m[747])|(m[720]&~m[721]&m[722]&~m[723]&~m[747])|(~m[720]&m[721]&m[722]&~m[723]&~m[747])|(m[720]&m[721]&m[722]&~m[723]&~m[747])|(m[720]&m[721]&m[722]&m[723]&~m[747])|(m[720]&m[721]&~m[722]&~m[723]&m[747])|(m[720]&~m[721]&m[722]&~m[723]&m[747])|(~m[720]&m[721]&m[722]&~m[723]&m[747])|(m[720]&m[721]&m[722]&~m[723]&m[747])|(m[720]&m[721]&m[722]&m[723]&m[747]));
    m[729] = (((m[725]&~m[726]&~m[727]&~m[728]&~m[752])|(~m[725]&m[726]&~m[727]&~m[728]&~m[752])|(~m[725]&~m[726]&m[727]&~m[728]&~m[752])|(m[725]&m[726]&~m[727]&m[728]&~m[752])|(m[725]&~m[726]&m[727]&m[728]&~m[752])|(~m[725]&m[726]&m[727]&m[728]&~m[752]))&BiasedRNG[412])|(((m[725]&~m[726]&~m[727]&~m[728]&m[752])|(~m[725]&m[726]&~m[727]&~m[728]&m[752])|(~m[725]&~m[726]&m[727]&~m[728]&m[752])|(m[725]&m[726]&~m[727]&m[728]&m[752])|(m[725]&~m[726]&m[727]&m[728]&m[752])|(~m[725]&m[726]&m[727]&m[728]&m[752]))&~BiasedRNG[412])|((m[725]&m[726]&~m[727]&~m[728]&~m[752])|(m[725]&~m[726]&m[727]&~m[728]&~m[752])|(~m[725]&m[726]&m[727]&~m[728]&~m[752])|(m[725]&m[726]&m[727]&~m[728]&~m[752])|(m[725]&m[726]&m[727]&m[728]&~m[752])|(m[725]&m[726]&~m[727]&~m[728]&m[752])|(m[725]&~m[726]&m[727]&~m[728]&m[752])|(~m[725]&m[726]&m[727]&~m[728]&m[752])|(m[725]&m[726]&m[727]&~m[728]&m[752])|(m[725]&m[726]&m[727]&m[728]&m[752]));
    m[734] = (((m[730]&~m[731]&~m[732]&~m[733]&~m[757])|(~m[730]&m[731]&~m[732]&~m[733]&~m[757])|(~m[730]&~m[731]&m[732]&~m[733]&~m[757])|(m[730]&m[731]&~m[732]&m[733]&~m[757])|(m[730]&~m[731]&m[732]&m[733]&~m[757])|(~m[730]&m[731]&m[732]&m[733]&~m[757]))&BiasedRNG[413])|(((m[730]&~m[731]&~m[732]&~m[733]&m[757])|(~m[730]&m[731]&~m[732]&~m[733]&m[757])|(~m[730]&~m[731]&m[732]&~m[733]&m[757])|(m[730]&m[731]&~m[732]&m[733]&m[757])|(m[730]&~m[731]&m[732]&m[733]&m[757])|(~m[730]&m[731]&m[732]&m[733]&m[757]))&~BiasedRNG[413])|((m[730]&m[731]&~m[732]&~m[733]&~m[757])|(m[730]&~m[731]&m[732]&~m[733]&~m[757])|(~m[730]&m[731]&m[732]&~m[733]&~m[757])|(m[730]&m[731]&m[732]&~m[733]&~m[757])|(m[730]&m[731]&m[732]&m[733]&~m[757])|(m[730]&m[731]&~m[732]&~m[733]&m[757])|(m[730]&~m[731]&m[732]&~m[733]&m[757])|(~m[730]&m[731]&m[732]&~m[733]&m[757])|(m[730]&m[731]&m[732]&~m[733]&m[757])|(m[730]&m[731]&m[732]&m[733]&m[757]));
    m[739] = (((m[735]&~m[736]&~m[737]&~m[738]&~m[760])|(~m[735]&m[736]&~m[737]&~m[738]&~m[760])|(~m[735]&~m[736]&m[737]&~m[738]&~m[760])|(m[735]&m[736]&~m[737]&m[738]&~m[760])|(m[735]&~m[736]&m[737]&m[738]&~m[760])|(~m[735]&m[736]&m[737]&m[738]&~m[760]))&BiasedRNG[414])|(((m[735]&~m[736]&~m[737]&~m[738]&m[760])|(~m[735]&m[736]&~m[737]&~m[738]&m[760])|(~m[735]&~m[736]&m[737]&~m[738]&m[760])|(m[735]&m[736]&~m[737]&m[738]&m[760])|(m[735]&~m[736]&m[737]&m[738]&m[760])|(~m[735]&m[736]&m[737]&m[738]&m[760]))&~BiasedRNG[414])|((m[735]&m[736]&~m[737]&~m[738]&~m[760])|(m[735]&~m[736]&m[737]&~m[738]&~m[760])|(~m[735]&m[736]&m[737]&~m[738]&~m[760])|(m[735]&m[736]&m[737]&~m[738]&~m[760])|(m[735]&m[736]&m[737]&m[738]&~m[760])|(m[735]&m[736]&~m[737]&~m[738]&m[760])|(m[735]&~m[736]&m[737]&~m[738]&m[760])|(~m[735]&m[736]&m[737]&~m[738]&m[760])|(m[735]&m[736]&m[737]&~m[738]&m[760])|(m[735]&m[736]&m[737]&m[738]&m[760]));
    m[744] = (((m[740]&~m[741]&~m[742]&~m[743]&~m[762])|(~m[740]&m[741]&~m[742]&~m[743]&~m[762])|(~m[740]&~m[741]&m[742]&~m[743]&~m[762])|(m[740]&m[741]&~m[742]&m[743]&~m[762])|(m[740]&~m[741]&m[742]&m[743]&~m[762])|(~m[740]&m[741]&m[742]&m[743]&~m[762]))&BiasedRNG[415])|(((m[740]&~m[741]&~m[742]&~m[743]&m[762])|(~m[740]&m[741]&~m[742]&~m[743]&m[762])|(~m[740]&~m[741]&m[742]&~m[743]&m[762])|(m[740]&m[741]&~m[742]&m[743]&m[762])|(m[740]&~m[741]&m[742]&m[743]&m[762])|(~m[740]&m[741]&m[742]&m[743]&m[762]))&~BiasedRNG[415])|((m[740]&m[741]&~m[742]&~m[743]&~m[762])|(m[740]&~m[741]&m[742]&~m[743]&~m[762])|(~m[740]&m[741]&m[742]&~m[743]&~m[762])|(m[740]&m[741]&m[742]&~m[743]&~m[762])|(m[740]&m[741]&m[742]&m[743]&~m[762])|(m[740]&m[741]&~m[742]&~m[743]&m[762])|(m[740]&~m[741]&m[742]&~m[743]&m[762])|(~m[740]&m[741]&m[742]&~m[743]&m[762])|(m[740]&m[741]&m[742]&~m[743]&m[762])|(m[740]&m[741]&m[742]&m[743]&m[762]));
    m[749] = (((m[745]&~m[746]&~m[747]&~m[748]&~m[767])|(~m[745]&m[746]&~m[747]&~m[748]&~m[767])|(~m[745]&~m[746]&m[747]&~m[748]&~m[767])|(m[745]&m[746]&~m[747]&m[748]&~m[767])|(m[745]&~m[746]&m[747]&m[748]&~m[767])|(~m[745]&m[746]&m[747]&m[748]&~m[767]))&BiasedRNG[416])|(((m[745]&~m[746]&~m[747]&~m[748]&m[767])|(~m[745]&m[746]&~m[747]&~m[748]&m[767])|(~m[745]&~m[746]&m[747]&~m[748]&m[767])|(m[745]&m[746]&~m[747]&m[748]&m[767])|(m[745]&~m[746]&m[747]&m[748]&m[767])|(~m[745]&m[746]&m[747]&m[748]&m[767]))&~BiasedRNG[416])|((m[745]&m[746]&~m[747]&~m[748]&~m[767])|(m[745]&~m[746]&m[747]&~m[748]&~m[767])|(~m[745]&m[746]&m[747]&~m[748]&~m[767])|(m[745]&m[746]&m[747]&~m[748]&~m[767])|(m[745]&m[746]&m[747]&m[748]&~m[767])|(m[745]&m[746]&~m[747]&~m[748]&m[767])|(m[745]&~m[746]&m[747]&~m[748]&m[767])|(~m[745]&m[746]&m[747]&~m[748]&m[767])|(m[745]&m[746]&m[747]&~m[748]&m[767])|(m[745]&m[746]&m[747]&m[748]&m[767]));
    m[754] = (((m[750]&~m[751]&~m[752]&~m[753]&~m[772])|(~m[750]&m[751]&~m[752]&~m[753]&~m[772])|(~m[750]&~m[751]&m[752]&~m[753]&~m[772])|(m[750]&m[751]&~m[752]&m[753]&~m[772])|(m[750]&~m[751]&m[752]&m[753]&~m[772])|(~m[750]&m[751]&m[752]&m[753]&~m[772]))&BiasedRNG[417])|(((m[750]&~m[751]&~m[752]&~m[753]&m[772])|(~m[750]&m[751]&~m[752]&~m[753]&m[772])|(~m[750]&~m[751]&m[752]&~m[753]&m[772])|(m[750]&m[751]&~m[752]&m[753]&m[772])|(m[750]&~m[751]&m[752]&m[753]&m[772])|(~m[750]&m[751]&m[752]&m[753]&m[772]))&~BiasedRNG[417])|((m[750]&m[751]&~m[752]&~m[753]&~m[772])|(m[750]&~m[751]&m[752]&~m[753]&~m[772])|(~m[750]&m[751]&m[752]&~m[753]&~m[772])|(m[750]&m[751]&m[752]&~m[753]&~m[772])|(m[750]&m[751]&m[752]&m[753]&~m[772])|(m[750]&m[751]&~m[752]&~m[753]&m[772])|(m[750]&~m[751]&m[752]&~m[753]&m[772])|(~m[750]&m[751]&m[752]&~m[753]&m[772])|(m[750]&m[751]&m[752]&~m[753]&m[772])|(m[750]&m[751]&m[752]&m[753]&m[772]));
    m[759] = (((m[755]&~m[756]&~m[757]&~m[758]&~m[777])|(~m[755]&m[756]&~m[757]&~m[758]&~m[777])|(~m[755]&~m[756]&m[757]&~m[758]&~m[777])|(m[755]&m[756]&~m[757]&m[758]&~m[777])|(m[755]&~m[756]&m[757]&m[758]&~m[777])|(~m[755]&m[756]&m[757]&m[758]&~m[777]))&BiasedRNG[418])|(((m[755]&~m[756]&~m[757]&~m[758]&m[777])|(~m[755]&m[756]&~m[757]&~m[758]&m[777])|(~m[755]&~m[756]&m[757]&~m[758]&m[777])|(m[755]&m[756]&~m[757]&m[758]&m[777])|(m[755]&~m[756]&m[757]&m[758]&m[777])|(~m[755]&m[756]&m[757]&m[758]&m[777]))&~BiasedRNG[418])|((m[755]&m[756]&~m[757]&~m[758]&~m[777])|(m[755]&~m[756]&m[757]&~m[758]&~m[777])|(~m[755]&m[756]&m[757]&~m[758]&~m[777])|(m[755]&m[756]&m[757]&~m[758]&~m[777])|(m[755]&m[756]&m[757]&m[758]&~m[777])|(m[755]&m[756]&~m[757]&~m[758]&m[777])|(m[755]&~m[756]&m[757]&~m[758]&m[777])|(~m[755]&m[756]&m[757]&~m[758]&m[777])|(m[755]&m[756]&m[757]&~m[758]&m[777])|(m[755]&m[756]&m[757]&m[758]&m[777]));
    m[764] = (((m[760]&~m[761]&~m[762]&~m[763]&~m[780])|(~m[760]&m[761]&~m[762]&~m[763]&~m[780])|(~m[760]&~m[761]&m[762]&~m[763]&~m[780])|(m[760]&m[761]&~m[762]&m[763]&~m[780])|(m[760]&~m[761]&m[762]&m[763]&~m[780])|(~m[760]&m[761]&m[762]&m[763]&~m[780]))&BiasedRNG[419])|(((m[760]&~m[761]&~m[762]&~m[763]&m[780])|(~m[760]&m[761]&~m[762]&~m[763]&m[780])|(~m[760]&~m[761]&m[762]&~m[763]&m[780])|(m[760]&m[761]&~m[762]&m[763]&m[780])|(m[760]&~m[761]&m[762]&m[763]&m[780])|(~m[760]&m[761]&m[762]&m[763]&m[780]))&~BiasedRNG[419])|((m[760]&m[761]&~m[762]&~m[763]&~m[780])|(m[760]&~m[761]&m[762]&~m[763]&~m[780])|(~m[760]&m[761]&m[762]&~m[763]&~m[780])|(m[760]&m[761]&m[762]&~m[763]&~m[780])|(m[760]&m[761]&m[762]&m[763]&~m[780])|(m[760]&m[761]&~m[762]&~m[763]&m[780])|(m[760]&~m[761]&m[762]&~m[763]&m[780])|(~m[760]&m[761]&m[762]&~m[763]&m[780])|(m[760]&m[761]&m[762]&~m[763]&m[780])|(m[760]&m[761]&m[762]&m[763]&m[780]));
    m[769] = (((m[765]&~m[766]&~m[767]&~m[768]&~m[782])|(~m[765]&m[766]&~m[767]&~m[768]&~m[782])|(~m[765]&~m[766]&m[767]&~m[768]&~m[782])|(m[765]&m[766]&~m[767]&m[768]&~m[782])|(m[765]&~m[766]&m[767]&m[768]&~m[782])|(~m[765]&m[766]&m[767]&m[768]&~m[782]))&BiasedRNG[420])|(((m[765]&~m[766]&~m[767]&~m[768]&m[782])|(~m[765]&m[766]&~m[767]&~m[768]&m[782])|(~m[765]&~m[766]&m[767]&~m[768]&m[782])|(m[765]&m[766]&~m[767]&m[768]&m[782])|(m[765]&~m[766]&m[767]&m[768]&m[782])|(~m[765]&m[766]&m[767]&m[768]&m[782]))&~BiasedRNG[420])|((m[765]&m[766]&~m[767]&~m[768]&~m[782])|(m[765]&~m[766]&m[767]&~m[768]&~m[782])|(~m[765]&m[766]&m[767]&~m[768]&~m[782])|(m[765]&m[766]&m[767]&~m[768]&~m[782])|(m[765]&m[766]&m[767]&m[768]&~m[782])|(m[765]&m[766]&~m[767]&~m[768]&m[782])|(m[765]&~m[766]&m[767]&~m[768]&m[782])|(~m[765]&m[766]&m[767]&~m[768]&m[782])|(m[765]&m[766]&m[767]&~m[768]&m[782])|(m[765]&m[766]&m[767]&m[768]&m[782]));
    m[774] = (((m[770]&~m[771]&~m[772]&~m[773]&~m[787])|(~m[770]&m[771]&~m[772]&~m[773]&~m[787])|(~m[770]&~m[771]&m[772]&~m[773]&~m[787])|(m[770]&m[771]&~m[772]&m[773]&~m[787])|(m[770]&~m[771]&m[772]&m[773]&~m[787])|(~m[770]&m[771]&m[772]&m[773]&~m[787]))&BiasedRNG[421])|(((m[770]&~m[771]&~m[772]&~m[773]&m[787])|(~m[770]&m[771]&~m[772]&~m[773]&m[787])|(~m[770]&~m[771]&m[772]&~m[773]&m[787])|(m[770]&m[771]&~m[772]&m[773]&m[787])|(m[770]&~m[771]&m[772]&m[773]&m[787])|(~m[770]&m[771]&m[772]&m[773]&m[787]))&~BiasedRNG[421])|((m[770]&m[771]&~m[772]&~m[773]&~m[787])|(m[770]&~m[771]&m[772]&~m[773]&~m[787])|(~m[770]&m[771]&m[772]&~m[773]&~m[787])|(m[770]&m[771]&m[772]&~m[773]&~m[787])|(m[770]&m[771]&m[772]&m[773]&~m[787])|(m[770]&m[771]&~m[772]&~m[773]&m[787])|(m[770]&~m[771]&m[772]&~m[773]&m[787])|(~m[770]&m[771]&m[772]&~m[773]&m[787])|(m[770]&m[771]&m[772]&~m[773]&m[787])|(m[770]&m[771]&m[772]&m[773]&m[787]));
    m[779] = (((m[775]&~m[776]&~m[777]&~m[778]&~m[792])|(~m[775]&m[776]&~m[777]&~m[778]&~m[792])|(~m[775]&~m[776]&m[777]&~m[778]&~m[792])|(m[775]&m[776]&~m[777]&m[778]&~m[792])|(m[775]&~m[776]&m[777]&m[778]&~m[792])|(~m[775]&m[776]&m[777]&m[778]&~m[792]))&BiasedRNG[422])|(((m[775]&~m[776]&~m[777]&~m[778]&m[792])|(~m[775]&m[776]&~m[777]&~m[778]&m[792])|(~m[775]&~m[776]&m[777]&~m[778]&m[792])|(m[775]&m[776]&~m[777]&m[778]&m[792])|(m[775]&~m[776]&m[777]&m[778]&m[792])|(~m[775]&m[776]&m[777]&m[778]&m[792]))&~BiasedRNG[422])|((m[775]&m[776]&~m[777]&~m[778]&~m[792])|(m[775]&~m[776]&m[777]&~m[778]&~m[792])|(~m[775]&m[776]&m[777]&~m[778]&~m[792])|(m[775]&m[776]&m[777]&~m[778]&~m[792])|(m[775]&m[776]&m[777]&m[778]&~m[792])|(m[775]&m[776]&~m[777]&~m[778]&m[792])|(m[775]&~m[776]&m[777]&~m[778]&m[792])|(~m[775]&m[776]&m[777]&~m[778]&m[792])|(m[775]&m[776]&m[777]&~m[778]&m[792])|(m[775]&m[776]&m[777]&m[778]&m[792]));
    m[784] = (((m[780]&~m[781]&~m[782]&~m[783]&~m[795])|(~m[780]&m[781]&~m[782]&~m[783]&~m[795])|(~m[780]&~m[781]&m[782]&~m[783]&~m[795])|(m[780]&m[781]&~m[782]&m[783]&~m[795])|(m[780]&~m[781]&m[782]&m[783]&~m[795])|(~m[780]&m[781]&m[782]&m[783]&~m[795]))&BiasedRNG[423])|(((m[780]&~m[781]&~m[782]&~m[783]&m[795])|(~m[780]&m[781]&~m[782]&~m[783]&m[795])|(~m[780]&~m[781]&m[782]&~m[783]&m[795])|(m[780]&m[781]&~m[782]&m[783]&m[795])|(m[780]&~m[781]&m[782]&m[783]&m[795])|(~m[780]&m[781]&m[782]&m[783]&m[795]))&~BiasedRNG[423])|((m[780]&m[781]&~m[782]&~m[783]&~m[795])|(m[780]&~m[781]&m[782]&~m[783]&~m[795])|(~m[780]&m[781]&m[782]&~m[783]&~m[795])|(m[780]&m[781]&m[782]&~m[783]&~m[795])|(m[780]&m[781]&m[782]&m[783]&~m[795])|(m[780]&m[781]&~m[782]&~m[783]&m[795])|(m[780]&~m[781]&m[782]&~m[783]&m[795])|(~m[780]&m[781]&m[782]&~m[783]&m[795])|(m[780]&m[781]&m[782]&~m[783]&m[795])|(m[780]&m[781]&m[782]&m[783]&m[795]));
    m[789] = (((m[785]&~m[786]&~m[787]&~m[788]&~m[797])|(~m[785]&m[786]&~m[787]&~m[788]&~m[797])|(~m[785]&~m[786]&m[787]&~m[788]&~m[797])|(m[785]&m[786]&~m[787]&m[788]&~m[797])|(m[785]&~m[786]&m[787]&m[788]&~m[797])|(~m[785]&m[786]&m[787]&m[788]&~m[797]))&BiasedRNG[424])|(((m[785]&~m[786]&~m[787]&~m[788]&m[797])|(~m[785]&m[786]&~m[787]&~m[788]&m[797])|(~m[785]&~m[786]&m[787]&~m[788]&m[797])|(m[785]&m[786]&~m[787]&m[788]&m[797])|(m[785]&~m[786]&m[787]&m[788]&m[797])|(~m[785]&m[786]&m[787]&m[788]&m[797]))&~BiasedRNG[424])|((m[785]&m[786]&~m[787]&~m[788]&~m[797])|(m[785]&~m[786]&m[787]&~m[788]&~m[797])|(~m[785]&m[786]&m[787]&~m[788]&~m[797])|(m[785]&m[786]&m[787]&~m[788]&~m[797])|(m[785]&m[786]&m[787]&m[788]&~m[797])|(m[785]&m[786]&~m[787]&~m[788]&m[797])|(m[785]&~m[786]&m[787]&~m[788]&m[797])|(~m[785]&m[786]&m[787]&~m[788]&m[797])|(m[785]&m[786]&m[787]&~m[788]&m[797])|(m[785]&m[786]&m[787]&m[788]&m[797]));
    m[794] = (((m[790]&~m[791]&~m[792]&~m[793]&~m[802])|(~m[790]&m[791]&~m[792]&~m[793]&~m[802])|(~m[790]&~m[791]&m[792]&~m[793]&~m[802])|(m[790]&m[791]&~m[792]&m[793]&~m[802])|(m[790]&~m[791]&m[792]&m[793]&~m[802])|(~m[790]&m[791]&m[792]&m[793]&~m[802]))&BiasedRNG[425])|(((m[790]&~m[791]&~m[792]&~m[793]&m[802])|(~m[790]&m[791]&~m[792]&~m[793]&m[802])|(~m[790]&~m[791]&m[792]&~m[793]&m[802])|(m[790]&m[791]&~m[792]&m[793]&m[802])|(m[790]&~m[791]&m[792]&m[793]&m[802])|(~m[790]&m[791]&m[792]&m[793]&m[802]))&~BiasedRNG[425])|((m[790]&m[791]&~m[792]&~m[793]&~m[802])|(m[790]&~m[791]&m[792]&~m[793]&~m[802])|(~m[790]&m[791]&m[792]&~m[793]&~m[802])|(m[790]&m[791]&m[792]&~m[793]&~m[802])|(m[790]&m[791]&m[792]&m[793]&~m[802])|(m[790]&m[791]&~m[792]&~m[793]&m[802])|(m[790]&~m[791]&m[792]&~m[793]&m[802])|(~m[790]&m[791]&m[792]&~m[793]&m[802])|(m[790]&m[791]&m[792]&~m[793]&m[802])|(m[790]&m[791]&m[792]&m[793]&m[802]));
    m[799] = (((m[795]&~m[796]&~m[797]&~m[798]&~m[805])|(~m[795]&m[796]&~m[797]&~m[798]&~m[805])|(~m[795]&~m[796]&m[797]&~m[798]&~m[805])|(m[795]&m[796]&~m[797]&m[798]&~m[805])|(m[795]&~m[796]&m[797]&m[798]&~m[805])|(~m[795]&m[796]&m[797]&m[798]&~m[805]))&BiasedRNG[426])|(((m[795]&~m[796]&~m[797]&~m[798]&m[805])|(~m[795]&m[796]&~m[797]&~m[798]&m[805])|(~m[795]&~m[796]&m[797]&~m[798]&m[805])|(m[795]&m[796]&~m[797]&m[798]&m[805])|(m[795]&~m[796]&m[797]&m[798]&m[805])|(~m[795]&m[796]&m[797]&m[798]&m[805]))&~BiasedRNG[426])|((m[795]&m[796]&~m[797]&~m[798]&~m[805])|(m[795]&~m[796]&m[797]&~m[798]&~m[805])|(~m[795]&m[796]&m[797]&~m[798]&~m[805])|(m[795]&m[796]&m[797]&~m[798]&~m[805])|(m[795]&m[796]&m[797]&m[798]&~m[805])|(m[795]&m[796]&~m[797]&~m[798]&m[805])|(m[795]&~m[796]&m[797]&~m[798]&m[805])|(~m[795]&m[796]&m[797]&~m[798]&m[805])|(m[795]&m[796]&m[797]&~m[798]&m[805])|(m[795]&m[796]&m[797]&m[798]&m[805]));
    m[804] = (((m[800]&~m[801]&~m[802]&~m[803]&~m[807])|(~m[800]&m[801]&~m[802]&~m[803]&~m[807])|(~m[800]&~m[801]&m[802]&~m[803]&~m[807])|(m[800]&m[801]&~m[802]&m[803]&~m[807])|(m[800]&~m[801]&m[802]&m[803]&~m[807])|(~m[800]&m[801]&m[802]&m[803]&~m[807]))&BiasedRNG[427])|(((m[800]&~m[801]&~m[802]&~m[803]&m[807])|(~m[800]&m[801]&~m[802]&~m[803]&m[807])|(~m[800]&~m[801]&m[802]&~m[803]&m[807])|(m[800]&m[801]&~m[802]&m[803]&m[807])|(m[800]&~m[801]&m[802]&m[803]&m[807])|(~m[800]&m[801]&m[802]&m[803]&m[807]))&~BiasedRNG[427])|((m[800]&m[801]&~m[802]&~m[803]&~m[807])|(m[800]&~m[801]&m[802]&~m[803]&~m[807])|(~m[800]&m[801]&m[802]&~m[803]&~m[807])|(m[800]&m[801]&m[802]&~m[803]&~m[807])|(m[800]&m[801]&m[802]&m[803]&~m[807])|(m[800]&m[801]&~m[802]&~m[803]&m[807])|(m[800]&~m[801]&m[802]&~m[803]&m[807])|(~m[800]&m[801]&m[802]&~m[803]&m[807])|(m[800]&m[801]&m[802]&~m[803]&m[807])|(m[800]&m[801]&m[802]&m[803]&m[807]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[334]&LFSRcolor0[146]&LFSRcolor0[42]&LFSRcolor0[430]);
    BiasedRNG[1] = (LFSRcolor0[351]&LFSRcolor0[137]&LFSRcolor0[495]&LFSRcolor0[236]);
    BiasedRNG[2] = (LFSRcolor0[237]&LFSRcolor0[381]&LFSRcolor0[101]&LFSRcolor0[480]);
    BiasedRNG[3] = (LFSRcolor0[33]&LFSRcolor0[419]&LFSRcolor0[192]&LFSRcolor0[281]);
    BiasedRNG[4] = (LFSRcolor0[428]&LFSRcolor0[261]&LFSRcolor0[246]&LFSRcolor0[216]);
    BiasedRNG[5] = (LFSRcolor0[394]&LFSRcolor0[51]&LFSRcolor0[313]&LFSRcolor0[404]);
    BiasedRNG[6] = (LFSRcolor0[355]&LFSRcolor0[40]&LFSRcolor0[443]&LFSRcolor0[364]);
    BiasedRNG[7] = (LFSRcolor0[366]&LFSRcolor0[331]&LFSRcolor0[504]&LFSRcolor0[176]);
    BiasedRNG[8] = (LFSRcolor0[466]&LFSRcolor0[361]&LFSRcolor0[385]&LFSRcolor0[124]);
    BiasedRNG[9] = (LFSRcolor0[57]&LFSRcolor0[106]&LFSRcolor0[327]&LFSRcolor0[110]);
    BiasedRNG[10] = (LFSRcolor0[362]&LFSRcolor0[104]&LFSRcolor0[178]&LFSRcolor0[482]);
    BiasedRNG[11] = (LFSRcolor0[312]&LFSRcolor0[69]&LFSRcolor0[147]&LFSRcolor0[84]);
    BiasedRNG[12] = (LFSRcolor0[314]&LFSRcolor0[191]&LFSRcolor0[303]&LFSRcolor0[341]);
    BiasedRNG[13] = (LFSRcolor0[67]&LFSRcolor0[14]&LFSRcolor0[53]&LFSRcolor0[299]);
    BiasedRNG[14] = (LFSRcolor0[289]&LFSRcolor0[166]&LFSRcolor0[224]&LFSRcolor0[348]);
    BiasedRNG[15] = (LFSRcolor0[474]&LFSRcolor0[210]&LFSRcolor0[123]&LFSRcolor0[417]);
    BiasedRNG[16] = (LFSRcolor0[204]&LFSRcolor0[347]&LFSRcolor0[52]&LFSRcolor0[268]);
    BiasedRNG[17] = (LFSRcolor0[481]&LFSRcolor0[346]&LFSRcolor0[456]&LFSRcolor0[477]);
    BiasedRNG[18] = (LFSRcolor0[354]&LFSRcolor0[20]&LFSRcolor0[95]&LFSRcolor0[134]);
    BiasedRNG[19] = (LFSRcolor0[196]&LFSRcolor0[251]&LFSRcolor0[308]&LFSRcolor0[189]);
    BiasedRNG[20] = (LFSRcolor0[399]&LFSRcolor0[382]&LFSRcolor0[181]&LFSRcolor0[490]);
    BiasedRNG[21] = (LFSRcolor0[10]&LFSRcolor0[212]&LFSRcolor0[55]&LFSRcolor0[56]);
    BiasedRNG[22] = (LFSRcolor0[76]&LFSRcolor0[22]&LFSRcolor0[185]&LFSRcolor0[441]);
    BiasedRNG[23] = (LFSRcolor0[409]&LFSRcolor0[398]&LFSRcolor0[282]&LFSRcolor0[335]);
    BiasedRNG[24] = (LFSRcolor0[72]&LFSRcolor0[2]&LFSRcolor0[68]&LFSRcolor0[454]);
    BiasedRNG[25] = (LFSRcolor0[140]&LFSRcolor0[375]&LFSRcolor0[345]&LFSRcolor0[78]);
    BiasedRNG[26] = (LFSRcolor0[437]&LFSRcolor0[183]&LFSRcolor0[242]&LFSRcolor0[152]);
    BiasedRNG[27] = (LFSRcolor0[301]&LFSRcolor0[431]&LFSRcolor0[460]&LFSRcolor0[370]);
    BiasedRNG[28] = (LFSRcolor0[328]&LFSRcolor0[330]&LFSRcolor0[38]&LFSRcolor0[108]);
    BiasedRNG[29] = (LFSRcolor0[115]&LFSRcolor0[378]&LFSRcolor0[352]&LFSRcolor0[471]);
    BiasedRNG[30] = (LFSRcolor0[203]&LFSRcolor0[159]&LFSRcolor0[12]&LFSRcolor0[422]);
    BiasedRNG[31] = (LFSRcolor0[438]&LFSRcolor0[219]&LFSRcolor0[119]&LFSRcolor0[318]);
    BiasedRNG[32] = (LFSRcolor0[424]&LFSRcolor0[35]&LFSRcolor0[85]&LFSRcolor0[49]);
    BiasedRNG[33] = (LFSRcolor0[505]&LFSRcolor0[86]&LFSRcolor0[358]&LFSRcolor0[410]);
    BiasedRNG[34] = (LFSRcolor0[129]&LFSRcolor0[118]&LFSRcolor0[151]&LFSRcolor0[426]);
    BiasedRNG[35] = (LFSRcolor0[93]&LFSRcolor0[70]&LFSRcolor0[28]&LFSRcolor0[80]);
    BiasedRNG[36] = (LFSRcolor0[179]&LFSRcolor0[421]&LFSRcolor0[102]&LFSRcolor0[451]);
    BiasedRNG[37] = (LFSRcolor0[50]&LFSRcolor0[464]&LFSRcolor0[150]&LFSRcolor0[325]);
    BiasedRNG[38] = (LFSRcolor0[255]&LFSRcolor0[478]&LFSRcolor0[66]&LFSRcolor0[31]);
    BiasedRNG[39] = (LFSRcolor0[180]&LFSRcolor0[208]&LFSRcolor0[463]&LFSRcolor0[500]);
    BiasedRNG[40] = (LFSRcolor0[472]&LFSRcolor0[408]&LFSRcolor0[266]&LFSRcolor0[493]);
    BiasedRNG[41] = (LFSRcolor0[243]&LFSRcolor0[496]&LFSRcolor0[186]&LFSRcolor0[158]);
    BiasedRNG[42] = (LFSRcolor0[218]&LFSRcolor0[25]&LFSRcolor0[233]&LFSRcolor0[267]);
    BiasedRNG[43] = (LFSRcolor0[486]&LFSRcolor0[135]&LFSRcolor0[376]&LFSRcolor0[46]);
    BiasedRNG[44] = (LFSRcolor0[254]&LFSRcolor0[143]&LFSRcolor0[332]&LFSRcolor0[407]);
    BiasedRNG[45] = (LFSRcolor0[112]&LFSRcolor0[81]&LFSRcolor0[316]&LFSRcolor0[4]);
    BiasedRNG[46] = (LFSRcolor0[156]&LFSRcolor0[0]&LFSRcolor0[247]&LFSRcolor0[5]);
    BiasedRNG[47] = (LFSRcolor0[194]&LFSRcolor0[436]&LFSRcolor0[479]&LFSRcolor0[402]);
    BiasedRNG[48] = (LFSRcolor0[214]&LFSRcolor0[414]&LFSRcolor0[343]&LFSRcolor0[356]);
    BiasedRNG[49] = (LFSRcolor0[207]&LFSRcolor0[241]&LFSRcolor0[349]&LFSRcolor0[400]);
    BiasedRNG[50] = (LFSRcolor0[295]&LFSRcolor0[461]&LFSRcolor0[256]&LFSRcolor0[162]);
    BiasedRNG[51] = (LFSRcolor0[59]&LFSRcolor0[326]&LFSRcolor0[206]&LFSRcolor0[427]);
    BiasedRNG[52] = (LFSRcolor0[485]&LFSRcolor0[82]&LFSRcolor0[36]&LFSRcolor0[447]);
    BiasedRNG[53] = (LFSRcolor0[369]&LFSRcolor0[322]&LFSRcolor0[293]&LFSRcolor0[501]);
    BiasedRNG[54] = (LFSRcolor0[449]&LFSRcolor0[97]&LFSRcolor0[100]&LFSRcolor0[231]);
    BiasedRNG[55] = (LFSRcolor0[125]&LFSRcolor0[163]&LFSRcolor0[468]&LFSRcolor0[154]);
    BiasedRNG[56] = (LFSRcolor0[155]&LFSRcolor0[445]&LFSRcolor0[309]&LFSRcolor0[277]);
    BiasedRNG[57] = (LFSRcolor0[333]&LFSRcolor0[201]&LFSRcolor0[274]&LFSRcolor0[244]);
    BiasedRNG[58] = (LFSRcolor0[337]&LFSRcolor0[499]&LFSRcolor0[418]&LFSRcolor0[77]);
    BiasedRNG[59] = (LFSRcolor0[232]&LFSRcolor0[103]&LFSRcolor0[287]&LFSRcolor0[462]);
    BiasedRNG[60] = (LFSRcolor0[306]&LFSRcolor0[258]&LFSRcolor0[126]&LFSRcolor0[9]);
    BiasedRNG[61] = (LFSRcolor0[265]&LFSRcolor0[429]&LFSRcolor0[222]&LFSRcolor0[483]);
    BiasedRNG[62] = (LFSRcolor0[305]&LFSRcolor0[395]&LFSRcolor0[223]&LFSRcolor0[453]);
    BiasedRNG[63] = (LFSRcolor0[131]&LFSRcolor0[448]&LFSRcolor0[283]&LFSRcolor0[74]);
    BiasedRNG[64] = (LFSRcolor0[13]&LFSRcolor0[109]&LFSRcolor0[220]&LFSRcolor0[240]);
    BiasedRNG[65] = (LFSRcolor0[434]&LFSRcolor0[487]&LFSRcolor0[75]&LFSRcolor0[433]);
    BiasedRNG[66] = (LFSRcolor0[113]&LFSRcolor0[23]&LFSRcolor0[439]&LFSRcolor0[465]);
    BiasedRNG[67] = (LFSRcolor0[171]&LFSRcolor0[492]&LFSRcolor0[21]&LFSRcolor0[190]);
    BiasedRNG[68] = (LFSRcolor0[489]&LFSRcolor0[435]&LFSRcolor0[167]&LFSRcolor0[459]);
    BiasedRNG[69] = (LFSRcolor0[248]&LFSRcolor0[397]&LFSRcolor0[368]&LFSRcolor0[172]);
    BiasedRNG[70] = (LFSRcolor0[209]&LFSRcolor0[357]&LFSRcolor0[217]&LFSRcolor0[195]);
    BiasedRNG[71] = (LFSRcolor0[132]&LFSRcolor0[275]&LFSRcolor0[188]&LFSRcolor0[469]);
    BiasedRNG[72] = (LFSRcolor0[286]&LFSRcolor0[116]&LFSRcolor0[403]&LFSRcolor0[360]);
    BiasedRNG[73] = (LFSRcolor0[169]&LFSRcolor0[300]&LFSRcolor0[7]&LFSRcolor0[494]);
    BiasedRNG[74] = (LFSRcolor0[442]&LFSRcolor0[392]&LFSRcolor0[393]&LFSRcolor0[262]);
    BiasedRNG[75] = (LFSRcolor0[396]&LFSRcolor0[372]&LFSRcolor0[73]&LFSRcolor0[197]);
    BiasedRNG[76] = (LFSRcolor0[446]&LFSRcolor0[359]&LFSRcolor0[65]&LFSRcolor0[484]);
    BiasedRNG[77] = (LFSRcolor0[229]&LFSRcolor0[27]&LFSRcolor0[401]&LFSRcolor0[39]);
    BiasedRNG[78] = (LFSRcolor0[455]&LFSRcolor0[473]&LFSRcolor0[142]&LFSRcolor0[18]);
    BiasedRNG[79] = (LFSRcolor0[470]&LFSRcolor0[211]&LFSRcolor0[226]&LFSRcolor0[319]);
    BiasedRNG[80] = (LFSRcolor0[141]&LFSRcolor0[32]&LFSRcolor0[285]&LFSRcolor0[122]);
    BiasedRNG[81] = (LFSRcolor0[34]&LFSRcolor0[245]&LFSRcolor0[444]&LFSRcolor0[260]);
    BiasedRNG[82] = (LFSRcolor0[149]&LFSRcolor0[114]&LFSRcolor0[383]&LFSRcolor0[450]);
    BiasedRNG[83] = (LFSRcolor0[89]&LFSRcolor0[193]&LFSRcolor0[175]&LFSRcolor0[177]);
    BiasedRNG[84] = (LFSRcolor0[228]&LFSRcolor0[457]&LFSRcolor0[88]&LFSRcolor0[41]);
    BiasedRNG[85] = (LFSRcolor0[145]&LFSRcolor0[297]&LFSRcolor0[160]&LFSRcolor0[491]);
    BiasedRNG[86] = (LFSRcolor0[111]&LFSRcolor0[272]&LFSRcolor0[234]&LFSRcolor0[227]);
    BiasedRNG[87] = (LFSRcolor0[153]&LFSRcolor0[161]&LFSRcolor0[54]&LFSRcolor0[284]);
    BiasedRNG[88] = (LFSRcolor0[276]&LFSRcolor0[288]&LFSRcolor0[249]&LFSRcolor0[415]);
    BiasedRNG[89] = (LFSRcolor0[182]&LFSRcolor0[8]&LFSRcolor0[329]&LFSRcolor0[202]);
    BiasedRNG[90] = (LFSRcolor0[165]&LFSRcolor0[384]&LFSRcolor0[379]&LFSRcolor0[270]);
    BiasedRNG[91] = (LFSRcolor0[259]&LFSRcolor0[336]&LFSRcolor0[290]&LFSRcolor0[502]);
    BiasedRNG[92] = (LFSRcolor0[1]&LFSRcolor0[307]&LFSRcolor0[174]&LFSRcolor0[339]);
    BiasedRNG[93] = (LFSRcolor0[79]&LFSRcolor0[47]&LFSRcolor0[377]&LFSRcolor0[105]);
    BiasedRNG[94] = (LFSRcolor0[117]&LFSRcolor0[371]&LFSRcolor0[16]&LFSRcolor0[315]);
    BiasedRNG[95] = (LFSRcolor0[37]&LFSRcolor0[298]&LFSRcolor0[389]&LFSRcolor0[127]);
    BiasedRNG[96] = (LFSRcolor0[238]&LFSRcolor0[83]&LFSRcolor0[304]&LFSRcolor0[411]);
    BiasedRNG[97] = (LFSRcolor0[253]&LFSRcolor0[252]&LFSRcolor0[107]&LFSRcolor0[416]);
    BiasedRNG[98] = (LFSRcolor0[94]&LFSRcolor0[296]&LFSRcolor0[440]&LFSRcolor0[387]);
    UnbiasedRNG[0] = LFSRcolor0[452];
    UnbiasedRNG[1] = LFSRcolor0[432];
    UnbiasedRNG[2] = LFSRcolor0[488];
    UnbiasedRNG[3] = LFSRcolor0[235];
    UnbiasedRNG[4] = LFSRcolor0[310];
    UnbiasedRNG[5] = LFSRcolor0[92];
    UnbiasedRNG[6] = LFSRcolor0[230];
    UnbiasedRNG[7] = LFSRcolor0[367];
    UnbiasedRNG[8] = LFSRcolor0[60];
    UnbiasedRNG[9] = LFSRcolor0[302];
    UnbiasedRNG[10] = LFSRcolor0[391];
    UnbiasedRNG[11] = LFSRcolor0[321];
    UnbiasedRNG[12] = LFSRcolor0[264];
    UnbiasedRNG[13] = LFSRcolor0[133];
    UnbiasedRNG[14] = LFSRcolor0[374];
    UnbiasedRNG[15] = LFSRcolor0[64];
    UnbiasedRNG[16] = LFSRcolor0[200];
    UnbiasedRNG[17] = LFSRcolor0[353];
    UnbiasedRNG[18] = LFSRcolor0[338];
    UnbiasedRNG[19] = LFSRcolor0[320];
    UnbiasedRNG[20] = LFSRcolor0[498];
    UnbiasedRNG[21] = LFSRcolor0[386];
    UnbiasedRNG[22] = LFSRcolor0[342];
    UnbiasedRNG[23] = LFSRcolor0[187];
    UnbiasedRNG[24] = LFSRcolor0[273];
    UnbiasedRNG[25] = LFSRcolor0[213];
    UnbiasedRNG[26] = LFSRcolor0[323];
    UnbiasedRNG[27] = LFSRcolor0[373];
    UnbiasedRNG[28] = LFSRcolor0[29];
    UnbiasedRNG[29] = LFSRcolor0[239];
    UnbiasedRNG[30] = LFSRcolor0[221];
    UnbiasedRNG[31] = LFSRcolor0[170];
    UnbiasedRNG[32] = LFSRcolor0[120];
    UnbiasedRNG[33] = LFSRcolor0[91];
    UnbiasedRNG[34] = LFSRcolor0[365];
    UnbiasedRNG[35] = LFSRcolor0[15];
    UnbiasedRNG[36] = LFSRcolor0[263];
    UnbiasedRNG[37] = LFSRcolor0[291];
    UnbiasedRNG[38] = LFSRcolor0[350];
    UnbiasedRNG[39] = LFSRcolor0[48];
    UnbiasedRNG[40] = LFSRcolor0[58];
    UnbiasedRNG[41] = LFSRcolor0[215];
    UnbiasedRNG[42] = LFSRcolor0[497];
    UnbiasedRNG[43] = LFSRcolor0[458];
    UnbiasedRNG[44] = LFSRcolor0[63];
    UnbiasedRNG[45] = LFSRcolor0[205];
    UnbiasedRNG[46] = LFSRcolor0[62];
    UnbiasedRNG[47] = LFSRcolor0[24];
    UnbiasedRNG[48] = LFSRcolor0[71];
    UnbiasedRNG[49] = LFSRcolor0[423];
    UnbiasedRNG[50] = LFSRcolor0[11];
    UnbiasedRNG[51] = LFSRcolor0[280];
    UnbiasedRNG[52] = LFSRcolor0[87];
    UnbiasedRNG[53] = LFSRcolor0[405];
    UnbiasedRNG[54] = LFSRcolor0[199];
    UnbiasedRNG[55] = LFSRcolor0[121];
    UnbiasedRNG[56] = LFSRcolor0[44];
    UnbiasedRNG[57] = LFSRcolor0[96];
    UnbiasedRNG[58] = LFSRcolor0[6];
    UnbiasedRNG[59] = LFSRcolor0[19];
    UnbiasedRNG[60] = LFSRcolor0[61];
    UnbiasedRNG[61] = LFSRcolor0[406];
    UnbiasedRNG[62] = LFSRcolor0[311];
    UnbiasedRNG[63] = LFSRcolor0[340];
    UnbiasedRNG[64] = LFSRcolor0[294];
    UnbiasedRNG[65] = LFSRcolor0[17];
    UnbiasedRNG[66] = LFSRcolor0[138];
    UnbiasedRNG[67] = LFSRcolor0[198];
    UnbiasedRNG[68] = LFSRcolor0[45];
    UnbiasedRNG[69] = LFSRcolor0[130];
    UnbiasedRNG[70] = LFSRcolor0[412];
    UnbiasedRNG[71] = LFSRcolor0[269];
    UnbiasedRNG[72] = LFSRcolor0[388];
    UnbiasedRNG[73] = LFSRcolor0[26];
    UnbiasedRNG[74] = LFSRcolor0[257];
    UnbiasedRNG[75] = LFSRcolor0[271];
    UnbiasedRNG[76] = LFSRcolor0[98];
    UnbiasedRNG[77] = LFSRcolor0[317];
    UnbiasedRNG[78] = LFSRcolor0[164];
    UnbiasedRNG[79] = LFSRcolor0[128];
    UnbiasedRNG[80] = LFSRcolor0[278];
    UnbiasedRNG[81] = LFSRcolor0[475];
    UnbiasedRNG[82] = LFSRcolor0[380];
    UnbiasedRNG[83] = LFSRcolor0[139];
    UnbiasedRNG[84] = LFSRcolor0[250];
    UnbiasedRNG[85] = LFSRcolor0[99];
    UnbiasedRNG[86] = LFSRcolor0[90];
    UnbiasedRNG[87] = LFSRcolor0[168];
    UnbiasedRNG[88] = LFSRcolor0[344];
    UnbiasedRNG[89] = LFSRcolor0[413];
    UnbiasedRNG[90] = LFSRcolor0[148];
    UnbiasedRNG[91] = LFSRcolor0[157];
    UnbiasedRNG[92] = LFSRcolor0[503];
    UnbiasedRNG[93] = LFSRcolor0[225];
    UnbiasedRNG[94] = LFSRcolor0[30];
    UnbiasedRNG[95] = LFSRcolor0[292];
    UnbiasedRNG[96] = LFSRcolor0[173];
    UnbiasedRNG[97] = LFSRcolor0[3];
    UnbiasedRNG[98] = LFSRcolor0[476];
    UnbiasedRNG[99] = LFSRcolor0[324];
    UnbiasedRNG[100] = LFSRcolor0[363];
    UnbiasedRNG[101] = LFSRcolor0[43];
    UnbiasedRNG[102] = LFSRcolor0[425];
    UnbiasedRNG[103] = LFSRcolor0[390];
    UnbiasedRNG[104] = LFSRcolor0[467];
    UnbiasedRNG[105] = LFSRcolor0[136];
    UnbiasedRNG[106] = LFSRcolor0[184];
    UnbiasedRNG[107] = LFSRcolor0[279];
end

always @(posedge color0_clk) begin
    BiasedRNG[99] = (LFSRcolor1[100]&LFSRcolor1[290]&LFSRcolor1[159]&LFSRcolor1[509]);
    BiasedRNG[100] = (LFSRcolor1[445]&LFSRcolor1[658]&LFSRcolor1[676]&LFSRcolor1[377]);
    BiasedRNG[101] = (LFSRcolor1[197]&LFSRcolor1[283]&LFSRcolor1[556]&LFSRcolor1[75]);
    BiasedRNG[102] = (LFSRcolor1[624]&LFSRcolor1[396]&LFSRcolor1[476]&LFSRcolor1[183]);
    BiasedRNG[103] = (LFSRcolor1[298]&LFSRcolor1[54]&LFSRcolor1[558]&LFSRcolor1[160]);
    BiasedRNG[104] = (LFSRcolor1[69]&LFSRcolor1[122]&LFSRcolor1[343]&LFSRcolor1[516]);
    BiasedRNG[105] = (LFSRcolor1[572]&LFSRcolor1[524]&LFSRcolor1[99]&LFSRcolor1[567]);
    BiasedRNG[106] = (LFSRcolor1[352]&LFSRcolor1[346]&LFSRcolor1[469]&LFSRcolor1[460]);
    BiasedRNG[107] = (LFSRcolor1[218]&LFSRcolor1[432]&LFSRcolor1[398]&LFSRcolor1[673]);
    BiasedRNG[108] = (LFSRcolor1[680]&LFSRcolor1[647]&LFSRcolor1[430]&LFSRcolor1[78]);
    BiasedRNG[109] = (LFSRcolor1[301]&LFSRcolor1[161]&LFSRcolor1[230]&LFSRcolor1[621]);
    BiasedRNG[110] = (LFSRcolor1[313]&LFSRcolor1[220]&LFSRcolor1[274]&LFSRcolor1[141]);
    BiasedRNG[111] = (LFSRcolor1[258]&LFSRcolor1[402]&LFSRcolor1[29]&LFSRcolor1[522]);
    BiasedRNG[112] = (LFSRcolor1[131]&LFSRcolor1[137]&LFSRcolor1[547]&LFSRcolor1[265]);
    BiasedRNG[113] = (LFSRcolor1[563]&LFSRcolor1[488]&LFSRcolor1[399]&LFSRcolor1[344]);
    BiasedRNG[114] = (LFSRcolor1[410]&LFSRcolor1[454]&LFSRcolor1[41]&LFSRcolor1[404]);
    BiasedRNG[115] = (LFSRcolor1[413]&LFSRcolor1[32]&LFSRcolor1[307]&LFSRcolor1[580]);
    BiasedRNG[116] = (LFSRcolor1[130]&LFSRcolor1[392]&LFSRcolor1[142]&LFSRcolor1[611]);
    BiasedRNG[117] = (LFSRcolor1[403]&LFSRcolor1[236]&LFSRcolor1[644]&LFSRcolor1[280]);
    BiasedRNG[118] = (LFSRcolor1[257]&LFSRcolor1[121]&LFSRcolor1[273]&LFSRcolor1[35]);
    BiasedRNG[119] = (LFSRcolor1[291]&LFSRcolor1[199]&LFSRcolor1[610]&LFSRcolor1[634]);
    BiasedRNG[120] = (LFSRcolor1[355]&LFSRcolor1[528]&LFSRcolor1[617]&LFSRcolor1[151]);
    BiasedRNG[121] = (LFSRcolor1[115]&LFSRcolor1[478]&LFSRcolor1[44]&LFSRcolor1[95]);
    BiasedRNG[122] = (LFSRcolor1[143]&LFSRcolor1[597]&LFSRcolor1[105]&LFSRcolor1[521]);
    BiasedRNG[123] = (LFSRcolor1[209]&LFSRcolor1[508]&LFSRcolor1[416]&LFSRcolor1[0]);
    BiasedRNG[124] = (LFSRcolor1[670]&LFSRcolor1[217]&LFSRcolor1[112]&LFSRcolor1[571]);
    BiasedRNG[125] = (LFSRcolor1[144]&LFSRcolor1[546]&LFSRcolor1[592]&LFSRcolor1[61]);
    BiasedRNG[126] = (LFSRcolor1[52]&LFSRcolor1[153]&LFSRcolor1[196]&LFSRcolor1[287]);
    BiasedRNG[127] = (LFSRcolor1[165]&LFSRcolor1[233]&LFSRcolor1[574]&LFSRcolor1[684]);
    BiasedRNG[128] = (LFSRcolor1[83]&LFSRcolor1[45]&LFSRcolor1[340]&LFSRcolor1[663]);
    BiasedRNG[129] = (LFSRcolor1[420]&LFSRcolor1[300]&LFSRcolor1[470]&LFSRcolor1[188]);
    BiasedRNG[130] = (LFSRcolor1[13]&LFSRcolor1[285]&LFSRcolor1[455]&LFSRcolor1[408]);
    BiasedRNG[131] = (LFSRcolor1[182]&LFSRcolor1[207]&LFSRcolor1[92]&LFSRcolor1[314]);
    BiasedRNG[132] = (LFSRcolor1[356]&LFSRcolor1[638]&LFSRcolor1[615]&LFSRcolor1[405]);
    BiasedRNG[133] = (LFSRcolor1[4]&LFSRcolor1[664]&LFSRcolor1[630]&LFSRcolor1[324]);
    BiasedRNG[134] = (LFSRcolor1[466]&LFSRcolor1[249]&LFSRcolor1[375]&LFSRcolor1[279]);
    BiasedRNG[135] = (LFSRcolor1[406]&LFSRcolor1[322]&LFSRcolor1[337]&LFSRcolor1[24]);
    BiasedRNG[136] = (LFSRcolor1[662]&LFSRcolor1[85]&LFSRcolor1[120]&LFSRcolor1[349]);
    BiasedRNG[137] = (LFSRcolor1[614]&LFSRcolor1[93]&LFSRcolor1[351]&LFSRcolor1[175]);
    BiasedRNG[138] = (LFSRcolor1[682]&LFSRcolor1[170]&LFSRcolor1[168]&LFSRcolor1[498]);
    BiasedRNG[139] = (LFSRcolor1[421]&LFSRcolor1[28]&LFSRcolor1[319]&LFSRcolor1[483]);
    BiasedRNG[140] = (LFSRcolor1[181]&LFSRcolor1[654]&LFSRcolor1[501]&LFSRcolor1[221]);
    BiasedRNG[141] = (LFSRcolor1[540]&LFSRcolor1[502]&LFSRcolor1[672]&LFSRcolor1[553]);
    BiasedRNG[142] = (LFSRcolor1[79]&LFSRcolor1[335]&LFSRcolor1[472]&LFSRcolor1[62]);
    BiasedRNG[143] = (LFSRcolor1[240]&LFSRcolor1[627]&LFSRcolor1[312]&LFSRcolor1[613]);
    BiasedRNG[144] = (LFSRcolor1[499]&LFSRcolor1[232]&LFSRcolor1[200]&LFSRcolor1[669]);
    BiasedRNG[145] = (LFSRcolor1[140]&LFSRcolor1[158]&LFSRcolor1[560]&LFSRcolor1[526]);
    BiasedRNG[146] = (LFSRcolor1[594]&LFSRcolor1[222]&LFSRcolor1[417]&LFSRcolor1[46]);
    BiasedRNG[147] = (LFSRcolor1[330]&LFSRcolor1[619]&LFSRcolor1[18]&LFSRcolor1[110]);
    BiasedRNG[148] = (LFSRcolor1[511]&LFSRcolor1[250]&LFSRcolor1[510]&LFSRcolor1[451]);
    BiasedRNG[149] = (LFSRcolor1[150]&LFSRcolor1[534]&LFSRcolor1[618]&LFSRcolor1[135]);
    BiasedRNG[150] = (LFSRcolor1[419]&LFSRcolor1[38]&LFSRcolor1[433]&LFSRcolor1[1]);
    BiasedRNG[151] = (LFSRcolor1[91]&LFSRcolor1[30]&LFSRcolor1[271]&LFSRcolor1[177]);
    BiasedRNG[152] = (LFSRcolor1[166]&LFSRcolor1[70]&LFSRcolor1[114]&LFSRcolor1[519]);
    BiasedRNG[153] = (LFSRcolor1[124]&LFSRcolor1[174]&LFSRcolor1[385]&LFSRcolor1[389]);
    BiasedRNG[154] = (LFSRcolor1[667]&LFSRcolor1[51]&LFSRcolor1[195]&LFSRcolor1[34]);
    BiasedRNG[155] = (LFSRcolor1[237]&LFSRcolor1[23]&LFSRcolor1[643]&LFSRcolor1[357]);
    BiasedRNG[156] = (LFSRcolor1[651]&LFSRcolor1[681]&LFSRcolor1[383]&LFSRcolor1[436]);
    BiasedRNG[157] = (LFSRcolor1[639]&LFSRcolor1[163]&LFSRcolor1[395]&LFSRcolor1[123]);
    BiasedRNG[158] = (LFSRcolor1[292]&LFSRcolor1[390]&LFSRcolor1[2]&LFSRcolor1[480]);
    BiasedRNG[159] = (LFSRcolor1[561]&LFSRcolor1[369]&LFSRcolor1[525]&LFSRcolor1[129]);
    BiasedRNG[160] = (LFSRcolor1[342]&LFSRcolor1[668]&LFSRcolor1[213]&LFSRcolor1[164]);
    BiasedRNG[161] = (LFSRcolor1[254]&LFSRcolor1[677]&LFSRcolor1[660]&LFSRcolor1[284]);
    BiasedRNG[162] = (LFSRcolor1[328]&LFSRcolor1[500]&LFSRcolor1[350]&LFSRcolor1[514]);
    BiasedRNG[163] = (LFSRcolor1[457]&LFSRcolor1[481]&LFSRcolor1[479]&LFSRcolor1[552]);
    BiasedRNG[164] = (LFSRcolor1[428]&LFSRcolor1[202]&LFSRcolor1[309]&LFSRcolor1[311]);
    BiasedRNG[165] = (LFSRcolor1[583]&LFSRcolor1[261]&LFSRcolor1[299]&LFSRcolor1[441]);
    BiasedRNG[166] = (LFSRcolor1[53]&LFSRcolor1[575]&LFSRcolor1[600]&LFSRcolor1[189]);
    BiasedRNG[167] = (LFSRcolor1[507]&LFSRcolor1[225]&LFSRcolor1[191]&LFSRcolor1[497]);
    BiasedRNG[168] = (LFSRcolor1[465]&LFSRcolor1[259]&LFSRcolor1[224]&LFSRcolor1[327]);
    BiasedRNG[169] = (LFSRcolor1[642]&LFSRcolor1[527]&LFSRcolor1[513]&LFSRcolor1[591]);
    BiasedRNG[170] = (LFSRcolor1[512]&LFSRcolor1[192]&LFSRcolor1[94]&LFSRcolor1[623]);
    BiasedRNG[171] = (LFSRcolor1[305]&LFSRcolor1[674]&LFSRcolor1[133]&LFSRcolor1[71]);
    BiasedRNG[172] = (LFSRcolor1[208]&LFSRcolor1[109]&LFSRcolor1[76]&LFSRcolor1[461]);
    BiasedRNG[173] = (LFSRcolor1[629]&LFSRcolor1[485]&LFSRcolor1[56]&LFSRcolor1[474]);
    BiasedRNG[174] = (LFSRcolor1[446]&LFSRcolor1[506]&LFSRcolor1[523]&LFSRcolor1[103]);
    BiasedRNG[175] = (LFSRcolor1[228]&LFSRcolor1[173]&LFSRcolor1[223]&LFSRcolor1[184]);
    BiasedRNG[176] = (LFSRcolor1[176]&LFSRcolor1[172]&LFSRcolor1[666]&LFSRcolor1[559]);
    BiasedRNG[177] = (LFSRcolor1[190]&LFSRcolor1[277]&LFSRcolor1[243]&LFSRcolor1[288]);
    BiasedRNG[178] = (LFSRcolor1[65]&LFSRcolor1[341]&LFSRcolor1[3]&LFSRcolor1[411]);
    BiasedRNG[179] = (LFSRcolor1[382]&LFSRcolor1[136]&LFSRcolor1[657]&LFSRcolor1[550]);
    BiasedRNG[180] = (LFSRcolor1[459]&LFSRcolor1[391]&LFSRcolor1[366]&LFSRcolor1[517]);
    BiasedRNG[181] = (LFSRcolor1[582]&LFSRcolor1[424]&LFSRcolor1[543]&LFSRcolor1[248]);
    BiasedRNG[182] = (LFSRcolor1[687]&LFSRcolor1[247]&LFSRcolor1[293]&LFSRcolor1[678]);
    BiasedRNG[183] = (LFSRcolor1[449]&LFSRcolor1[631]&LFSRcolor1[57]&LFSRcolor1[400]);
    BiasedRNG[184] = (LFSRcolor1[648]&LFSRcolor1[671]&LFSRcolor1[187]&LFSRcolor1[204]);
    BiasedRNG[185] = (LFSRcolor1[439]&LFSRcolor1[31]&LFSRcolor1[67]&LFSRcolor1[588]);
    BiasedRNG[186] = (LFSRcolor1[206]&LFSRcolor1[365]&LFSRcolor1[77]&LFSRcolor1[412]);
    BiasedRNG[187] = (LFSRcolor1[484]&LFSRcolor1[440]&LFSRcolor1[198]&LFSRcolor1[318]);
    BiasedRNG[188] = (LFSRcolor1[531]&LFSRcolor1[268]&LFSRcolor1[68]&LFSRcolor1[242]);
    BiasedRNG[189] = (LFSRcolor1[275]&LFSRcolor1[152]&LFSRcolor1[434]&LFSRcolor1[40]);
    BiasedRNG[190] = (LFSRcolor1[303]&LFSRcolor1[444]&LFSRcolor1[650]&LFSRcolor1[134]);
    BiasedRNG[191] = (LFSRcolor1[423]&LFSRcolor1[431]&LFSRcolor1[589]&LFSRcolor1[463]);
    BiasedRNG[192] = (LFSRcolor1[329]&LFSRcolor1[452]&LFSRcolor1[486]&LFSRcolor1[376]);
    BiasedRNG[193] = (LFSRcolor1[443]&LFSRcolor1[96]&LFSRcolor1[127]&LFSRcolor1[6]);
    BiasedRNG[194] = (LFSRcolor1[148]&LFSRcolor1[584]&LFSRcolor1[450]&LFSRcolor1[491]);
    BiasedRNG[195] = (LFSRcolor1[495]&LFSRcolor1[276]&LFSRcolor1[425]&LFSRcolor1[108]);
    BiasedRNG[196] = (LFSRcolor1[39]&LFSRcolor1[427]&LFSRcolor1[214]&LFSRcolor1[162]);
    BiasedRNG[197] = (LFSRcolor1[33]&LFSRcolor1[603]&LFSRcolor1[448]&LFSRcolor1[255]);
    BiasedRNG[198] = (LFSRcolor1[387]&LFSRcolor1[458]&LFSRcolor1[656]&LFSRcolor1[167]);
    BiasedRNG[199] = (LFSRcolor1[178]&LFSRcolor1[551]&LFSRcolor1[80]&LFSRcolor1[585]);
    BiasedRNG[200] = (LFSRcolor1[74]&LFSRcolor1[542]&LFSRcolor1[55]&LFSRcolor1[505]);
    BiasedRNG[201] = (LFSRcolor1[641]&LFSRcolor1[633]&LFSRcolor1[106]&LFSRcolor1[212]);
    BiasedRNG[202] = (LFSRcolor1[201]&LFSRcolor1[326]&LFSRcolor1[227]&LFSRcolor1[438]);
    BiasedRNG[203] = (LFSRcolor1[679]&LFSRcolor1[216]&LFSRcolor1[437]&LFSRcolor1[659]);
    BiasedRNG[204] = (LFSRcolor1[64]&LFSRcolor1[622]&LFSRcolor1[590]&LFSRcolor1[688]);
    BiasedRNG[205] = (LFSRcolor1[596]&LFSRcolor1[598]&LFSRcolor1[665]&LFSRcolor1[347]);
    BiasedRNG[206] = (LFSRcolor1[87]&LFSRcolor1[566]&LFSRcolor1[116]&LFSRcolor1[607]);
    BiasedRNG[207] = (LFSRcolor1[415]&LFSRcolor1[211]&LFSRcolor1[296]&LFSRcolor1[267]);
    BiasedRNG[208] = (LFSRcolor1[601]&LFSRcolor1[145]&LFSRcolor1[636]&LFSRcolor1[331]);
    BiasedRNG[209] = (LFSRcolor1[626]&LFSRcolor1[98]&LFSRcolor1[102]&LFSRcolor1[386]);
    BiasedRNG[210] = (LFSRcolor1[37]&LFSRcolor1[367]&LFSRcolor1[215]&LFSRcolor1[378]);
    BiasedRNG[211] = (LFSRcolor1[180]&LFSRcolor1[147]&LFSRcolor1[599]&LFSRcolor1[294]);
    BiasedRNG[212] = (LFSRcolor1[7]&LFSRcolor1[333]&LFSRcolor1[418]&LFSRcolor1[14]);
    BiasedRNG[213] = (LFSRcolor1[538]&LFSRcolor1[549]&LFSRcolor1[602]&LFSRcolor1[157]);
    BiasedRNG[214] = (LFSRcolor1[520]&LFSRcolor1[568]&LFSRcolor1[640]&LFSRcolor1[235]);
    BiasedRNG[215] = (LFSRcolor1[464]&LFSRcolor1[646]&LFSRcolor1[686]&LFSRcolor1[82]);
    BiasedRNG[216] = (LFSRcolor1[493]&LFSRcolor1[297]&LFSRcolor1[245]&LFSRcolor1[22]);
    BiasedRNG[217] = (LFSRcolor1[154]&LFSRcolor1[169]&LFSRcolor1[555]&LFSRcolor1[17]);
    BiasedRNG[218] = (LFSRcolor1[477]&LFSRcolor1[231]&LFSRcolor1[306]&LFSRcolor1[655]);
    BiasedRNG[219] = (LFSRcolor1[244]&LFSRcolor1[88]&LFSRcolor1[260]&LFSRcolor1[20]);
    BiasedRNG[220] = (LFSRcolor1[338]&LFSRcolor1[364]&LFSRcolor1[194]&LFSRcolor1[15]);
    BiasedRNG[221] = (LFSRcolor1[628]&LFSRcolor1[471]&LFSRcolor1[320]&LFSRcolor1[595]);
    BiasedRNG[222] = (LFSRcolor1[394]&LFSRcolor1[117]&LFSRcolor1[252]&LFSRcolor1[332]);
    BiasedRNG[223] = (LFSRcolor1[593]&LFSRcolor1[146]&LFSRcolor1[58]&LFSRcolor1[570]);
    BiasedRNG[224] = (LFSRcolor1[573]&LFSRcolor1[354]&LFSRcolor1[132]&LFSRcolor1[9]);
    BiasedRNG[225] = (LFSRcolor1[19]&LFSRcolor1[462]&LFSRcolor1[345]&LFSRcolor1[128]);
    BiasedRNG[226] = (LFSRcolor1[609]&LFSRcolor1[565]&LFSRcolor1[42]&LFSRcolor1[577]);
    BiasedRNG[227] = (LFSRcolor1[689]&LFSRcolor1[564]&LFSRcolor1[372]&LFSRcolor1[84]);
    BiasedRNG[228] = (LFSRcolor1[429]&LFSRcolor1[185]&LFSRcolor1[388]&LFSRcolor1[66]);
    BiasedRNG[229] = (LFSRcolor1[89]&LFSRcolor1[149]&LFSRcolor1[155]&LFSRcolor1[48]);
    BiasedRNG[230] = (LFSRcolor1[359]&LFSRcolor1[490]&LFSRcolor1[407]&LFSRcolor1[264]);
    BiasedRNG[231] = (LFSRcolor1[535]&LFSRcolor1[496]&LFSRcolor1[569]&LFSRcolor1[652]);
    BiasedRNG[232] = (LFSRcolor1[219]&LFSRcolor1[308]&LFSRcolor1[373]&LFSRcolor1[304]);
    BiasedRNG[233] = (LFSRcolor1[579]&LFSRcolor1[60]&LFSRcolor1[515]&LFSRcolor1[138]);
    BiasedRNG[234] = (LFSRcolor1[683]&LFSRcolor1[539]&LFSRcolor1[381]&LFSRcolor1[310]);
    BiasedRNG[235] = (LFSRcolor1[336]&LFSRcolor1[363]&LFSRcolor1[282]&LFSRcolor1[435]);
    BiasedRNG[236] = (LFSRcolor1[545]&LFSRcolor1[179]&LFSRcolor1[637]&LFSRcolor1[101]);
    BiasedRNG[237] = (LFSRcolor1[530]&LFSRcolor1[21]&LFSRcolor1[118]&LFSRcolor1[453]);
    BiasedRNG[238] = (LFSRcolor1[548]&LFSRcolor1[27]&LFSRcolor1[47]&LFSRcolor1[649]);
    UnbiasedRNG[108] = LFSRcolor1[63];
    UnbiasedRNG[109] = LFSRcolor1[518];
    UnbiasedRNG[110] = LFSRcolor1[467];
    UnbiasedRNG[111] = LFSRcolor1[239];
    UnbiasedRNG[112] = LFSRcolor1[353];
    UnbiasedRNG[113] = LFSRcolor1[653];
    UnbiasedRNG[114] = LFSRcolor1[186];
    UnbiasedRNG[115] = LFSRcolor1[104];
    UnbiasedRNG[116] = LFSRcolor1[156];
    UnbiasedRNG[117] = LFSRcolor1[302];
    UnbiasedRNG[118] = LFSRcolor1[632];
    UnbiasedRNG[119] = LFSRcolor1[97];
    UnbiasedRNG[120] = LFSRcolor1[10];
    UnbiasedRNG[121] = LFSRcolor1[12];
    UnbiasedRNG[122] = LFSRcolor1[5];
    UnbiasedRNG[123] = LFSRcolor1[612];
    UnbiasedRNG[124] = LFSRcolor1[397];
    UnbiasedRNG[125] = LFSRcolor1[73];
    UnbiasedRNG[126] = LFSRcolor1[380];
    UnbiasedRNG[127] = LFSRcolor1[358];
    UnbiasedRNG[128] = LFSRcolor1[625];
    UnbiasedRNG[129] = LFSRcolor1[339];
    UnbiasedRNG[130] = LFSRcolor1[368];
    UnbiasedRNG[131] = LFSRcolor1[504];
    UnbiasedRNG[132] = LFSRcolor1[468];
    UnbiasedRNG[133] = LFSRcolor1[475];
    UnbiasedRNG[134] = LFSRcolor1[323];
    UnbiasedRNG[135] = LFSRcolor1[272];
    UnbiasedRNG[136] = LFSRcolor1[473];
    UnbiasedRNG[137] = LFSRcolor1[263];
    UnbiasedRNG[138] = LFSRcolor1[489];
    UnbiasedRNG[139] = LFSRcolor1[256];
    UnbiasedRNG[140] = LFSRcolor1[26];
    UnbiasedRNG[141] = LFSRcolor1[270];
    UnbiasedRNG[142] = LFSRcolor1[25];
    UnbiasedRNG[143] = LFSRcolor1[409];
    UnbiasedRNG[144] = LFSRcolor1[374];
    UnbiasedRNG[145] = LFSRcolor1[295];
    UnbiasedRNG[146] = LFSRcolor1[334];
    UnbiasedRNG[147] = LFSRcolor1[246];
    UnbiasedRNG[148] = LFSRcolor1[262];
    UnbiasedRNG[149] = LFSRcolor1[616];
    UnbiasedRNG[150] = LFSRcolor1[370];
    UnbiasedRNG[151] = LFSRcolor1[675];
    UnbiasedRNG[152] = LFSRcolor1[205];
    UnbiasedRNG[153] = LFSRcolor1[266];
    UnbiasedRNG[154] = LFSRcolor1[321];
    UnbiasedRNG[155] = LFSRcolor1[532];
    UnbiasedRNG[156] = LFSRcolor1[50];
    UnbiasedRNG[157] = LFSRcolor1[456];
    UnbiasedRNG[158] = LFSRcolor1[393];
    UnbiasedRNG[159] = LFSRcolor1[494];
    UnbiasedRNG[160] = LFSRcolor1[315];
    UnbiasedRNG[161] = LFSRcolor1[503];
    UnbiasedRNG[162] = LFSRcolor1[487];
    UnbiasedRNG[163] = LFSRcolor1[43];
    UnbiasedRNG[164] = LFSRcolor1[587];
    UnbiasedRNG[165] = LFSRcolor1[8];
    UnbiasedRNG[166] = LFSRcolor1[360];
    UnbiasedRNG[167] = LFSRcolor1[111];
    UnbiasedRNG[168] = LFSRcolor1[49];
    UnbiasedRNG[169] = LFSRcolor1[139];
    UnbiasedRNG[170] = LFSRcolor1[269];
    UnbiasedRNG[171] = LFSRcolor1[562];
    UnbiasedRNG[172] = LFSRcolor1[605];
    UnbiasedRNG[173] = LFSRcolor1[226];
    UnbiasedRNG[174] = LFSRcolor1[362];
    UnbiasedRNG[175] = LFSRcolor1[586];
    UnbiasedRNG[176] = LFSRcolor1[361];
    UnbiasedRNG[177] = LFSRcolor1[171];
    UnbiasedRNG[178] = LFSRcolor1[113];
    UnbiasedRNG[179] = LFSRcolor1[581];
    UnbiasedRNG[180] = LFSRcolor1[442];
    UnbiasedRNG[181] = LFSRcolor1[554];
    UnbiasedRNG[182] = LFSRcolor1[125];
    UnbiasedRNG[183] = LFSRcolor1[529];
    UnbiasedRNG[184] = LFSRcolor1[422];
    UnbiasedRNG[185] = LFSRcolor1[119];
    UnbiasedRNG[186] = LFSRcolor1[541];
    UnbiasedRNG[187] = LFSRcolor1[241];
    UnbiasedRNG[188] = LFSRcolor1[86];
    UnbiasedRNG[189] = LFSRcolor1[203];
    UnbiasedRNG[190] = LFSRcolor1[317];
    UnbiasedRNG[191] = LFSRcolor1[620];
    UnbiasedRNG[192] = LFSRcolor1[325];
    UnbiasedRNG[193] = LFSRcolor1[544];
    UnbiasedRNG[194] = LFSRcolor1[253];
    UnbiasedRNG[195] = LFSRcolor1[371];
    UnbiasedRNG[196] = LFSRcolor1[193];
    UnbiasedRNG[197] = LFSRcolor1[278];
end

always @(posedge color1_clk) begin
    BiasedRNG[239] = (LFSRcolor2[205]&LFSRcolor2[176]&LFSRcolor2[98]&LFSRcolor2[484]);
    BiasedRNG[240] = (LFSRcolor2[21]&LFSRcolor2[299]&LFSRcolor2[101]&LFSRcolor2[273]);
    BiasedRNG[241] = (LFSRcolor2[425]&LFSRcolor2[191]&LFSRcolor2[323]&LFSRcolor2[173]);
    BiasedRNG[242] = (LFSRcolor2[417]&LFSRcolor2[436]&LFSRcolor2[306]&LFSRcolor2[268]);
    BiasedRNG[243] = (LFSRcolor2[289]&LFSRcolor2[316]&LFSRcolor2[263]&LFSRcolor2[125]);
    BiasedRNG[244] = (LFSRcolor2[73]&LFSRcolor2[386]&LFSRcolor2[457]&LFSRcolor2[19]);
    BiasedRNG[245] = (LFSRcolor2[395]&LFSRcolor2[91]&LFSRcolor2[385]&LFSRcolor2[317]);
    BiasedRNG[246] = (LFSRcolor2[459]&LFSRcolor2[275]&LFSRcolor2[85]&LFSRcolor2[96]);
    BiasedRNG[247] = (LFSRcolor2[295]&LFSRcolor2[234]&LFSRcolor2[81]&LFSRcolor2[461]);
    BiasedRNG[248] = (LFSRcolor2[237]&LFSRcolor2[118]&LFSRcolor2[164]&LFSRcolor2[387]);
    BiasedRNG[249] = (LFSRcolor2[207]&LFSRcolor2[65]&LFSRcolor2[190]&LFSRcolor2[121]);
    BiasedRNG[250] = (LFSRcolor2[45]&LFSRcolor2[402]&LFSRcolor2[262]&LFSRcolor2[475]);
    BiasedRNG[251] = (LFSRcolor2[272]&LFSRcolor2[351]&LFSRcolor2[203]&LFSRcolor2[498]);
    BiasedRNG[252] = (LFSRcolor2[418]&LFSRcolor2[119]&LFSRcolor2[162]&LFSRcolor2[408]);
    BiasedRNG[253] = (LFSRcolor2[84]&LFSRcolor2[233]&LFSRcolor2[242]&LFSRcolor2[146]);
    BiasedRNG[254] = (LFSRcolor2[77]&LFSRcolor2[446]&LFSRcolor2[482]&LFSRcolor2[56]);
    BiasedRNG[255] = (LFSRcolor2[94]&LFSRcolor2[60]&LFSRcolor2[269]&LFSRcolor2[251]);
    BiasedRNG[256] = (LFSRcolor2[93]&LFSRcolor2[326]&LFSRcolor2[296]&LFSRcolor2[297]);
    BiasedRNG[257] = (LFSRcolor2[80]&LFSRcolor2[224]&LFSRcolor2[490]&LFSRcolor2[122]);
    BiasedRNG[258] = (LFSRcolor2[375]&LFSRcolor2[79]&LFSRcolor2[491]&LFSRcolor2[312]);
    BiasedRNG[259] = (LFSRcolor2[472]&LFSRcolor2[32]&LFSRcolor2[305]&LFSRcolor2[152]);
    BiasedRNG[260] = (LFSRcolor2[384]&LFSRcolor2[424]&LFSRcolor2[329]&LFSRcolor2[324]);
    BiasedRNG[261] = (LFSRcolor2[249]&LFSRcolor2[478]&LFSRcolor2[336]&LFSRcolor2[499]);
    BiasedRNG[262] = (LFSRcolor2[398]&LFSRcolor2[357]&LFSRcolor2[467]&LFSRcolor2[143]);
    BiasedRNG[263] = (LFSRcolor2[24]&LFSRcolor2[133]&LFSRcolor2[487]&LFSRcolor2[279]);
    BiasedRNG[264] = (LFSRcolor2[136]&LFSRcolor2[53]&LFSRcolor2[213]&LFSRcolor2[181]);
    BiasedRNG[265] = (LFSRcolor2[481]&LFSRcolor2[288]&LFSRcolor2[62]&LFSRcolor2[209]);
    BiasedRNG[266] = (LFSRcolor2[328]&LFSRcolor2[350]&LFSRcolor2[453]&LFSRcolor2[72]);
    BiasedRNG[267] = (LFSRcolor2[206]&LFSRcolor2[41]&LFSRcolor2[103]&LFSRcolor2[155]);
    BiasedRNG[268] = (LFSRcolor2[108]&LFSRcolor2[260]&LFSRcolor2[367]&LFSRcolor2[455]);
    BiasedRNG[269] = (LFSRcolor2[413]&LFSRcolor2[4]&LFSRcolor2[473]&LFSRcolor2[157]);
    BiasedRNG[270] = (LFSRcolor2[75]&LFSRcolor2[2]&LFSRcolor2[180]&LFSRcolor2[495]);
    BiasedRNG[271] = (LFSRcolor2[381]&LFSRcolor2[248]&LFSRcolor2[348]&LFSRcolor2[13]);
    BiasedRNG[272] = (LFSRcolor2[124]&LFSRcolor2[74]&LFSRcolor2[252]&LFSRcolor2[410]);
    BiasedRNG[273] = (LFSRcolor2[369]&LFSRcolor2[466]&LFSRcolor2[458]&LFSRcolor2[244]);
    BiasedRNG[274] = (LFSRcolor2[280]&LFSRcolor2[285]&LFSRcolor2[439]&LFSRcolor2[30]);
    BiasedRNG[275] = (LFSRcolor2[138]&LFSRcolor2[265]&LFSRcolor2[390]&LFSRcolor2[378]);
    BiasedRNG[276] = (LFSRcolor2[304]&LFSRcolor2[188]&LFSRcolor2[366]&LFSRcolor2[212]);
    BiasedRNG[277] = (LFSRcolor2[435]&LFSRcolor2[476]&LFSRcolor2[214]&LFSRcolor2[36]);
    BiasedRNG[278] = (LFSRcolor2[179]&LFSRcolor2[309]&LFSRcolor2[396]&LFSRcolor2[493]);
    BiasedRNG[279] = (LFSRcolor2[428]&LFSRcolor2[447]&LFSRcolor2[241]&LFSRcolor2[35]);
    BiasedRNG[280] = (LFSRcolor2[308]&LFSRcolor2[204]&LFSRcolor2[58]&LFSRcolor2[99]);
    BiasedRNG[281] = (LFSRcolor2[379]&LFSRcolor2[255]&LFSRcolor2[216]&LFSRcolor2[440]);
    BiasedRNG[282] = (LFSRcolor2[175]&LFSRcolor2[86]&LFSRcolor2[442]&LFSRcolor2[327]);
    BiasedRNG[283] = (LFSRcolor2[197]&LFSRcolor2[352]&LFSRcolor2[76]&LFSRcolor2[353]);
    BiasedRNG[284] = (LFSRcolor2[18]&LFSRcolor2[392]&LFSRcolor2[330]&LFSRcolor2[344]);
    BiasedRNG[285] = (LFSRcolor2[92]&LFSRcolor2[131]&LFSRcolor2[465]&LFSRcolor2[360]);
    BiasedRNG[286] = (LFSRcolor2[189]&LFSRcolor2[356]&LFSRcolor2[321]&LFSRcolor2[169]);
    BiasedRNG[287] = (LFSRcolor2[20]&LFSRcolor2[500]&LFSRcolor2[391]&LFSRcolor2[257]);
    BiasedRNG[288] = (LFSRcolor2[127]&LFSRcolor2[167]&LFSRcolor2[82]&LFSRcolor2[40]);
    BiasedRNG[289] = (LFSRcolor2[339]&LFSRcolor2[239]&LFSRcolor2[54]&LFSRcolor2[355]);
    BiasedRNG[290] = (LFSRcolor2[470]&LFSRcolor2[303]&LFSRcolor2[198]&LFSRcolor2[208]);
    BiasedRNG[291] = (LFSRcolor2[423]&LFSRcolor2[120]&LFSRcolor2[345]&LFSRcolor2[300]);
    BiasedRNG[292] = (LFSRcolor2[219]&LFSRcolor2[178]&LFSRcolor2[6]&LFSRcolor2[388]);
    BiasedRNG[293] = (LFSRcolor2[416]&LFSRcolor2[16]&LFSRcolor2[480]&LFSRcolor2[55]);
    BiasedRNG[294] = (LFSRcolor2[14]&LFSRcolor2[38]&LFSRcolor2[114]&LFSRcolor2[128]);
    BiasedRNG[295] = (LFSRcolor2[404]&LFSRcolor2[39]&LFSRcolor2[148]&LFSRcolor2[415]);
    BiasedRNG[296] = (LFSRcolor2[26]&LFSRcolor2[444]&LFSRcolor2[111]&LFSRcolor2[405]);
    BiasedRNG[297] = (LFSRcolor2[374]&LFSRcolor2[46]&LFSRcolor2[170]&LFSRcolor2[411]);
    BiasedRNG[298] = (LFSRcolor2[130]&LFSRcolor2[474]&LFSRcolor2[50]&LFSRcolor2[420]);
    BiasedRNG[299] = (LFSRcolor2[311]&LFSRcolor2[104]&LFSRcolor2[380]&LFSRcolor2[347]);
    BiasedRNG[300] = (LFSRcolor2[215]&LFSRcolor2[302]&LFSRcolor2[200]&LFSRcolor2[292]);
    BiasedRNG[301] = (LFSRcolor2[401]&LFSRcolor2[168]&LFSRcolor2[245]&LFSRcolor2[290]);
    BiasedRNG[302] = (LFSRcolor2[494]&LFSRcolor2[293]&LFSRcolor2[281]&LFSRcolor2[365]);
    BiasedRNG[303] = (LFSRcolor2[477]&LFSRcolor2[322]&LFSRcolor2[438]&LFSRcolor2[483]);
    BiasedRNG[304] = (LFSRcolor2[9]&LFSRcolor2[485]&LFSRcolor2[318]&LFSRcolor2[464]);
    BiasedRNG[305] = (LFSRcolor2[505]&LFSRcolor2[61]&LFSRcolor2[147]&LFSRcolor2[112]);
    BiasedRNG[306] = (LFSRcolor2[373]&LFSRcolor2[319]&LFSRcolor2[228]&LFSRcolor2[132]);
    BiasedRNG[307] = (LFSRcolor2[441]&LFSRcolor2[109]&LFSRcolor2[23]&LFSRcolor2[48]);
    BiasedRNG[308] = (LFSRcolor2[240]&LFSRcolor2[445]&LFSRcolor2[502]&LFSRcolor2[399]);
    BiasedRNG[309] = (LFSRcolor2[8]&LFSRcolor2[186]&LFSRcolor2[140]&LFSRcolor2[195]);
    BiasedRNG[310] = (LFSRcolor2[42]&LFSRcolor2[78]&LFSRcolor2[354]&LFSRcolor2[346]);
    BiasedRNG[311] = (LFSRcolor2[194]&LFSRcolor2[340]&LFSRcolor2[450]&LFSRcolor2[256]);
    BiasedRNG[312] = (LFSRcolor2[421]&LFSRcolor2[412]&LFSRcolor2[64]&LFSRcolor2[49]);
    BiasedRNG[313] = (LFSRcolor2[258]&LFSRcolor2[426]&LFSRcolor2[407]&LFSRcolor2[433]);
    BiasedRNG[314] = (LFSRcolor2[503]&LFSRcolor2[282]&LFSRcolor2[468]&LFSRcolor2[57]);
    BiasedRNG[315] = (LFSRcolor2[271]&LFSRcolor2[221]&LFSRcolor2[479]&LFSRcolor2[51]);
    BiasedRNG[316] = (LFSRcolor2[70]&LFSRcolor2[422]&LFSRcolor2[363]&LFSRcolor2[63]);
    BiasedRNG[317] = (LFSRcolor2[371]&LFSRcolor2[161]&LFSRcolor2[202]&LFSRcolor2[432]);
    BiasedRNG[318] = (LFSRcolor2[211]&LFSRcolor2[7]&LFSRcolor2[12]&LFSRcolor2[67]);
    BiasedRNG[319] = (LFSRcolor2[307]&LFSRcolor2[199]&LFSRcolor2[222]&LFSRcolor2[287]);
    BiasedRNG[320] = (LFSRcolor2[238]&LFSRcolor2[460]&LFSRcolor2[246]&LFSRcolor2[449]);
    BiasedRNG[321] = (LFSRcolor2[105]&LFSRcolor2[158]&LFSRcolor2[462]&LFSRcolor2[486]);
    BiasedRNG[322] = (LFSRcolor2[504]&LFSRcolor2[431]&LFSRcolor2[492]&LFSRcolor2[171]);
    BiasedRNG[323] = (LFSRcolor2[141]&LFSRcolor2[452]&LFSRcolor2[337]&LFSRcolor2[274]);
    BiasedRNG[324] = (LFSRcolor2[427]&LFSRcolor2[437]&LFSRcolor2[389]&LFSRcolor2[144]);
    BiasedRNG[325] = (LFSRcolor2[10]&LFSRcolor2[187]&LFSRcolor2[87]&LFSRcolor2[134]);
    BiasedRNG[326] = (LFSRcolor2[196]&LFSRcolor2[451]&LFSRcolor2[333]&LFSRcolor2[116]);
    BiasedRNG[327] = (LFSRcolor2[47]&LFSRcolor2[5]&LFSRcolor2[135]&LFSRcolor2[361]);
    BiasedRNG[328] = (LFSRcolor2[342]&LFSRcolor2[66]&LFSRcolor2[469]&LFSRcolor2[69]);
    BiasedRNG[329] = (LFSRcolor2[123]&LFSRcolor2[429]&LFSRcolor2[313]&LFSRcolor2[362]);
    BiasedRNG[330] = (LFSRcolor2[151]&LFSRcolor2[149]&LFSRcolor2[95]&LFSRcolor2[294]);
    BiasedRNG[331] = (LFSRcolor2[115]&LFSRcolor2[253]&LFSRcolor2[225]&LFSRcolor2[254]);
    BiasedRNG[332] = (LFSRcolor2[90]&LFSRcolor2[247]&LFSRcolor2[117]&LFSRcolor2[27]);
    BiasedRNG[333] = (LFSRcolor2[184]&LFSRcolor2[193]&LFSRcolor2[400]&LFSRcolor2[335]);
    BiasedRNG[334] = (LFSRcolor2[250]&LFSRcolor2[310]&LFSRcolor2[377]&LFSRcolor2[154]);
    BiasedRNG[335] = (LFSRcolor2[232]&LFSRcolor2[266]&LFSRcolor2[113]&LFSRcolor2[43]);
    BiasedRNG[336] = (LFSRcolor2[267]&LFSRcolor2[226]&LFSRcolor2[372]&LFSRcolor2[160]);
    BiasedRNG[337] = (LFSRcolor2[22]&LFSRcolor2[278]&LFSRcolor2[150]&LFSRcolor2[358]);
    BiasedRNG[338] = (LFSRcolor2[145]&LFSRcolor2[172]&LFSRcolor2[236]&LFSRcolor2[331]);
    UnbiasedRNG[198] = LFSRcolor2[284];
    UnbiasedRNG[199] = LFSRcolor2[338];
    UnbiasedRNG[200] = LFSRcolor2[229];
    UnbiasedRNG[201] = LFSRcolor2[100];
    UnbiasedRNG[202] = LFSRcolor2[314];
    UnbiasedRNG[203] = LFSRcolor2[174];
    UnbiasedRNG[204] = LFSRcolor2[142];
    UnbiasedRNG[205] = LFSRcolor2[409];
    UnbiasedRNG[206] = LFSRcolor2[3];
    UnbiasedRNG[207] = LFSRcolor2[185];
    UnbiasedRNG[208] = LFSRcolor2[291];
    UnbiasedRNG[209] = LFSRcolor2[364];
    UnbiasedRNG[210] = LFSRcolor2[349];
    UnbiasedRNG[211] = LFSRcolor2[301];
    UnbiasedRNG[212] = LFSRcolor2[343];
    UnbiasedRNG[213] = LFSRcolor2[298];
    UnbiasedRNG[214] = LFSRcolor2[97];
    UnbiasedRNG[215] = LFSRcolor2[37];
    UnbiasedRNG[216] = LFSRcolor2[220];
    UnbiasedRNG[217] = LFSRcolor2[227];
    UnbiasedRNG[218] = LFSRcolor2[277];
    UnbiasedRNG[219] = LFSRcolor2[201];
    UnbiasedRNG[220] = LFSRcolor2[88];
    UnbiasedRNG[221] = LFSRcolor2[33];
    UnbiasedRNG[222] = LFSRcolor2[177];
    UnbiasedRNG[223] = LFSRcolor2[368];
    UnbiasedRNG[224] = LFSRcolor2[471];
    UnbiasedRNG[225] = LFSRcolor2[501];
    UnbiasedRNG[226] = LFSRcolor2[454];
    UnbiasedRNG[227] = LFSRcolor2[156];
    UnbiasedRNG[228] = LFSRcolor2[106];
    UnbiasedRNG[229] = LFSRcolor2[29];
    UnbiasedRNG[230] = LFSRcolor2[456];
    UnbiasedRNG[231] = LFSRcolor2[463];
    UnbiasedRNG[232] = LFSRcolor2[44];
    UnbiasedRNG[233] = LFSRcolor2[217];
    UnbiasedRNG[234] = LFSRcolor2[376];
    UnbiasedRNG[235] = LFSRcolor2[218];
    UnbiasedRNG[236] = LFSRcolor2[286];
    UnbiasedRNG[237] = LFSRcolor2[320];
    UnbiasedRNG[238] = LFSRcolor2[488];
    UnbiasedRNG[239] = LFSRcolor2[403];
    UnbiasedRNG[240] = LFSRcolor2[166];
    UnbiasedRNG[241] = LFSRcolor2[334];
    UnbiasedRNG[242] = LFSRcolor2[261];
    UnbiasedRNG[243] = LFSRcolor2[443];
    UnbiasedRNG[244] = LFSRcolor2[430];
    UnbiasedRNG[245] = LFSRcolor2[110];
    UnbiasedRNG[246] = LFSRcolor2[129];
    UnbiasedRNG[247] = LFSRcolor2[1];
    UnbiasedRNG[248] = LFSRcolor2[406];
    UnbiasedRNG[249] = LFSRcolor2[68];
    UnbiasedRNG[250] = LFSRcolor2[182];
    UnbiasedRNG[251] = LFSRcolor2[397];
    UnbiasedRNG[252] = LFSRcolor2[243];
    UnbiasedRNG[253] = LFSRcolor2[165];
    UnbiasedRNG[254] = LFSRcolor2[448];
    UnbiasedRNG[255] = LFSRcolor2[264];
    UnbiasedRNG[256] = LFSRcolor2[419];
    UnbiasedRNG[257] = LFSRcolor2[489];
    UnbiasedRNG[258] = LFSRcolor2[192];
    UnbiasedRNG[259] = LFSRcolor2[394];
    UnbiasedRNG[260] = LFSRcolor2[31];
    UnbiasedRNG[261] = LFSRcolor2[139];
    UnbiasedRNG[262] = LFSRcolor2[52];
    UnbiasedRNG[263] = LFSRcolor2[370];
    UnbiasedRNG[264] = LFSRcolor2[325];
    UnbiasedRNG[265] = LFSRcolor2[497];
    UnbiasedRNG[266] = LFSRcolor2[137];
    UnbiasedRNG[267] = LFSRcolor2[210];
    UnbiasedRNG[268] = LFSRcolor2[183];
    UnbiasedRNG[269] = LFSRcolor2[83];
    UnbiasedRNG[270] = LFSRcolor2[34];
    UnbiasedRNG[271] = LFSRcolor2[0];
    UnbiasedRNG[272] = LFSRcolor2[276];
    UnbiasedRNG[273] = LFSRcolor2[153];
    UnbiasedRNG[274] = LFSRcolor2[383];
    UnbiasedRNG[275] = LFSRcolor2[11];
    UnbiasedRNG[276] = LFSRcolor2[126];
    UnbiasedRNG[277] = LFSRcolor2[71];
    UnbiasedRNG[278] = LFSRcolor2[283];
    UnbiasedRNG[279] = LFSRcolor2[223];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[280] = LFSRcolor3[43];
    UnbiasedRNG[281] = LFSRcolor3[59];
    UnbiasedRNG[282] = LFSRcolor3[37];
    UnbiasedRNG[283] = LFSRcolor3[50];
    UnbiasedRNG[284] = LFSRcolor3[16];
    UnbiasedRNG[285] = LFSRcolor3[31];
    UnbiasedRNG[286] = LFSRcolor3[63];
    UnbiasedRNG[287] = LFSRcolor3[3];
    UnbiasedRNG[288] = LFSRcolor3[66];
    UnbiasedRNG[289] = LFSRcolor3[13];
    UnbiasedRNG[290] = LFSRcolor3[27];
    UnbiasedRNG[291] = LFSRcolor3[28];
    UnbiasedRNG[292] = LFSRcolor3[10];
    UnbiasedRNG[293] = LFSRcolor3[19];
    UnbiasedRNG[294] = LFSRcolor3[84];
    UnbiasedRNG[295] = LFSRcolor3[88];
    UnbiasedRNG[296] = LFSRcolor3[56];
    UnbiasedRNG[297] = LFSRcolor3[33];
    UnbiasedRNG[298] = LFSRcolor3[82];
    UnbiasedRNG[299] = LFSRcolor3[73];
    UnbiasedRNG[300] = LFSRcolor3[85];
    UnbiasedRNG[301] = LFSRcolor3[2];
    UnbiasedRNG[302] = LFSRcolor3[38];
    UnbiasedRNG[303] = LFSRcolor3[90];
    UnbiasedRNG[304] = LFSRcolor3[34];
    UnbiasedRNG[305] = LFSRcolor3[67];
    UnbiasedRNG[306] = LFSRcolor3[46];
    UnbiasedRNG[307] = LFSRcolor3[0];
    UnbiasedRNG[308] = LFSRcolor3[25];
    UnbiasedRNG[309] = LFSRcolor3[1];
    UnbiasedRNG[310] = LFSRcolor3[18];
    UnbiasedRNG[311] = LFSRcolor3[7];
    UnbiasedRNG[312] = LFSRcolor3[52];
    UnbiasedRNG[313] = LFSRcolor3[41];
    UnbiasedRNG[314] = LFSRcolor3[49];
    UnbiasedRNG[315] = LFSRcolor3[36];
    UnbiasedRNG[316] = LFSRcolor3[57];
    UnbiasedRNG[317] = LFSRcolor3[83];
    UnbiasedRNG[318] = LFSRcolor3[11];
    UnbiasedRNG[319] = LFSRcolor3[86];
    UnbiasedRNG[320] = LFSRcolor3[79];
    UnbiasedRNG[321] = LFSRcolor3[80];
    UnbiasedRNG[322] = LFSRcolor3[58];
    UnbiasedRNG[323] = LFSRcolor3[8];
    UnbiasedRNG[324] = LFSRcolor3[17];
    UnbiasedRNG[325] = LFSRcolor3[14];
    UnbiasedRNG[326] = LFSRcolor3[44];
    UnbiasedRNG[327] = LFSRcolor3[21];
    UnbiasedRNG[328] = LFSRcolor3[39];
    UnbiasedRNG[329] = LFSRcolor3[4];
    UnbiasedRNG[330] = LFSRcolor3[76];
    UnbiasedRNG[331] = LFSRcolor3[89];
    UnbiasedRNG[332] = LFSRcolor3[9];
    UnbiasedRNG[333] = LFSRcolor3[15];
    UnbiasedRNG[334] = LFSRcolor3[64];
    UnbiasedRNG[335] = LFSRcolor3[62];
    UnbiasedRNG[336] = LFSRcolor3[45];
    UnbiasedRNG[337] = LFSRcolor3[78];
    UnbiasedRNG[338] = LFSRcolor3[24];
    UnbiasedRNG[339] = LFSRcolor3[12];
    UnbiasedRNG[340] = LFSRcolor3[40];
    UnbiasedRNG[341] = LFSRcolor3[30];
    UnbiasedRNG[342] = LFSRcolor3[72];
    UnbiasedRNG[343] = LFSRcolor3[51];
    UnbiasedRNG[344] = LFSRcolor3[87];
    UnbiasedRNG[345] = LFSRcolor3[48];
    UnbiasedRNG[346] = LFSRcolor3[22];
    UnbiasedRNG[347] = LFSRcolor3[32];
    UnbiasedRNG[348] = LFSRcolor3[60];
    UnbiasedRNG[349] = LFSRcolor3[5];
    UnbiasedRNG[350] = LFSRcolor3[77];
    UnbiasedRNG[351] = LFSRcolor3[65];
end

always @(posedge color3_clk) begin
    BiasedRNG[339] = (LFSRcolor4[305]&LFSRcolor4[128]&LFSRcolor4[23]&LFSRcolor4[66]);
    BiasedRNG[340] = (LFSRcolor4[205]&LFSRcolor4[22]&LFSRcolor4[283]&LFSRcolor4[90]);
    BiasedRNG[341] = (LFSRcolor4[189]&LFSRcolor4[224]&LFSRcolor4[56]&LFSRcolor4[149]);
    BiasedRNG[342] = (LFSRcolor4[315]&LFSRcolor4[327]&LFSRcolor4[30]&LFSRcolor4[304]);
    BiasedRNG[343] = (LFSRcolor4[320]&LFSRcolor4[300]&LFSRcolor4[72]&LFSRcolor4[177]);
    BiasedRNG[344] = (LFSRcolor4[36]&LFSRcolor4[250]&LFSRcolor4[272]&LFSRcolor4[136]);
    BiasedRNG[345] = (LFSRcolor4[234]&LFSRcolor4[311]&LFSRcolor4[242]&LFSRcolor4[8]);
    BiasedRNG[346] = (LFSRcolor4[193]&LFSRcolor4[277]&LFSRcolor4[285]&LFSRcolor4[27]);
    BiasedRNG[347] = (LFSRcolor4[41]&LFSRcolor4[130]&LFSRcolor4[29]&LFSRcolor4[171]);
    BiasedRNG[348] = (LFSRcolor4[338]&LFSRcolor4[31]&LFSRcolor4[25]&LFSRcolor4[5]);
    BiasedRNG[349] = (LFSRcolor4[297]&LFSRcolor4[20]&LFSRcolor4[109]&LFSRcolor4[70]);
    BiasedRNG[350] = (LFSRcolor4[59]&LFSRcolor4[170]&LFSRcolor4[160]&LFSRcolor4[54]);
    BiasedRNG[351] = (LFSRcolor4[119]&LFSRcolor4[11]&LFSRcolor4[214]&LFSRcolor4[166]);
    BiasedRNG[352] = (LFSRcolor4[58]&LFSRcolor4[239]&LFSRcolor4[192]&LFSRcolor4[264]);
    BiasedRNG[353] = (LFSRcolor4[196]&LFSRcolor4[347]&LFSRcolor4[209]&LFSRcolor4[52]);
    BiasedRNG[354] = (LFSRcolor4[269]&LFSRcolor4[256]&LFSRcolor4[75]&LFSRcolor4[69]);
    BiasedRNG[355] = (LFSRcolor4[176]&LFSRcolor4[340]&LFSRcolor4[115]&LFSRcolor4[76]);
    BiasedRNG[356] = (LFSRcolor4[203]&LFSRcolor4[275]&LFSRcolor4[138]&LFSRcolor4[350]);
    BiasedRNG[357] = (LFSRcolor4[181]&LFSRcolor4[85]&LFSRcolor4[53]&LFSRcolor4[122]);
    BiasedRNG[358] = (LFSRcolor4[162]&LFSRcolor4[245]&LFSRcolor4[169]&LFSRcolor4[310]);
    BiasedRNG[359] = (LFSRcolor4[6]&LFSRcolor4[299]&LFSRcolor4[38]&LFSRcolor4[291]);
    BiasedRNG[360] = (LFSRcolor4[204]&LFSRcolor4[306]&LFSRcolor4[78]&LFSRcolor4[164]);
    BiasedRNG[361] = (LFSRcolor4[336]&LFSRcolor4[173]&LFSRcolor4[137]&LFSRcolor4[108]);
    BiasedRNG[362] = (LFSRcolor4[290]&LFSRcolor4[295]&LFSRcolor4[167]&LFSRcolor4[187]);
    BiasedRNG[363] = (LFSRcolor4[81]&LFSRcolor4[334]&LFSRcolor4[47]&LFSRcolor4[141]);
    BiasedRNG[364] = (LFSRcolor4[324]&LFSRcolor4[319]&LFSRcolor4[280]&LFSRcolor4[229]);
    BiasedRNG[365] = (LFSRcolor4[281]&LFSRcolor4[117]&LFSRcolor4[49]&LFSRcolor4[263]);
    BiasedRNG[366] = (LFSRcolor4[211]&LFSRcolor4[116]&LFSRcolor4[216]&LFSRcolor4[57]);
    BiasedRNG[367] = (LFSRcolor4[344]&LFSRcolor4[37]&LFSRcolor4[325]&LFSRcolor4[126]);
    BiasedRNG[368] = (LFSRcolor4[352]&LFSRcolor4[332]&LFSRcolor4[80]&LFSRcolor4[287]);
    BiasedRNG[369] = (LFSRcolor4[63]&LFSRcolor4[91]&LFSRcolor4[301]&LFSRcolor4[147]);
    BiasedRNG[370] = (LFSRcolor4[261]&LFSRcolor4[221]&LFSRcolor4[270]&LFSRcolor4[55]);
    BiasedRNG[371] = (LFSRcolor4[73]&LFSRcolor4[174]&LFSRcolor4[180]&LFSRcolor4[257]);
    BiasedRNG[372] = (LFSRcolor4[97]&LFSRcolor4[267]&LFSRcolor4[271]&LFSRcolor4[105]);
    BiasedRNG[373] = (LFSRcolor4[19]&LFSRcolor4[168]&LFSRcolor4[129]&LFSRcolor4[346]);
    BiasedRNG[374] = (LFSRcolor4[161]&LFSRcolor4[212]&LFSRcolor4[150]&LFSRcolor4[293]);
    BiasedRNG[375] = (LFSRcolor4[102]&LFSRcolor4[335]&LFSRcolor4[121]&LFSRcolor4[142]);
    BiasedRNG[376] = (LFSRcolor4[84]&LFSRcolor4[237]&LFSRcolor4[246]&LFSRcolor4[228]);
    BiasedRNG[377] = (LFSRcolor4[201]&LFSRcolor4[159]&LFSRcolor4[248]&LFSRcolor4[175]);
    BiasedRNG[378] = (LFSRcolor4[292]&LFSRcolor4[14]&LFSRcolor4[223]&LFSRcolor4[326]);
    BiasedRNG[379] = (LFSRcolor4[104]&LFSRcolor4[207]&LFSRcolor4[13]&LFSRcolor4[26]);
    BiasedRNG[380] = (LFSRcolor4[226]&LFSRcolor4[241]&LFSRcolor4[183]&LFSRcolor4[131]);
    BiasedRNG[381] = (LFSRcolor4[240]&LFSRcolor4[17]&LFSRcolor4[339]&LFSRcolor4[64]);
    BiasedRNG[382] = (LFSRcolor4[233]&LFSRcolor4[154]&LFSRcolor4[92]&LFSRcolor4[43]);
    BiasedRNG[383] = (LFSRcolor4[185]&LFSRcolor4[32]&LFSRcolor4[114]&LFSRcolor4[83]);
    BiasedRNG[384] = (LFSRcolor4[230]&LFSRcolor4[244]&LFSRcolor4[12]&LFSRcolor4[15]);
    BiasedRNG[385] = (LFSRcolor4[77]&LFSRcolor4[313]&LFSRcolor4[62]&LFSRcolor4[98]);
    BiasedRNG[386] = (LFSRcolor4[123]&LFSRcolor4[50]&LFSRcolor4[262]&LFSRcolor4[360]);
    BiasedRNG[387] = (LFSRcolor4[134]&LFSRcolor4[86]&LFSRcolor4[302]&LFSRcolor4[132]);
    BiasedRNG[388] = (LFSRcolor4[39]&LFSRcolor4[111]&LFSRcolor4[95]&LFSRcolor4[156]);
    BiasedRNG[389] = (LFSRcolor4[34]&LFSRcolor4[144]&LFSRcolor4[289]&LFSRcolor4[243]);
    BiasedRNG[390] = (LFSRcolor4[274]&LFSRcolor4[16]&LFSRcolor4[273]&LFSRcolor4[7]);
    BiasedRNG[391] = (LFSRcolor4[345]&LFSRcolor4[365]&LFSRcolor4[284]&LFSRcolor4[140]);
    BiasedRNG[392] = (LFSRcolor4[79]&LFSRcolor4[158]&LFSRcolor4[312]&LFSRcolor4[318]);
    BiasedRNG[393] = (LFSRcolor4[182]&LFSRcolor4[46]&LFSRcolor4[220]&LFSRcolor4[74]);
    BiasedRNG[394] = (LFSRcolor4[44]&LFSRcolor4[282]&LFSRcolor4[266]&LFSRcolor4[355]);
    BiasedRNG[395] = (LFSRcolor4[188]&LFSRcolor4[165]&LFSRcolor4[82]&LFSRcolor4[279]);
    BiasedRNG[396] = (LFSRcolor4[321]&LFSRcolor4[197]&LFSRcolor4[199]&LFSRcolor4[247]);
    BiasedRNG[397] = (LFSRcolor4[100]&LFSRcolor4[342]&LFSRcolor4[296]&LFSRcolor4[343]);
    BiasedRNG[398] = (LFSRcolor4[139]&LFSRcolor4[198]&LFSRcolor4[35]&LFSRcolor4[10]);
    BiasedRNG[399] = (LFSRcolor4[367]&LFSRcolor4[260]&LFSRcolor4[18]&LFSRcolor4[323]);
    BiasedRNG[400] = (LFSRcolor4[101]&LFSRcolor4[191]&LFSRcolor4[236]&LFSRcolor4[178]);
    BiasedRNG[401] = (LFSRcolor4[276]&LFSRcolor4[225]&LFSRcolor4[87]&LFSRcolor4[113]);
    BiasedRNG[402] = (LFSRcolor4[48]&LFSRcolor4[143]&LFSRcolor4[9]&LFSRcolor4[96]);
    BiasedRNG[403] = (LFSRcolor4[120]&LFSRcolor4[93]&LFSRcolor4[51]&LFSRcolor4[2]);
    BiasedRNG[404] = (LFSRcolor4[24]&LFSRcolor4[45]&LFSRcolor4[303]&LFSRcolor4[298]);
    BiasedRNG[405] = (LFSRcolor4[1]&LFSRcolor4[330]&LFSRcolor4[232]&LFSRcolor4[251]);
    BiasedRNG[406] = (LFSRcolor4[333]&LFSRcolor4[238]&LFSRcolor4[67]&LFSRcolor4[153]);
    BiasedRNG[407] = (LFSRcolor4[124]&LFSRcolor4[107]&LFSRcolor4[252]&LFSRcolor4[210]);
    BiasedRNG[408] = (LFSRcolor4[366]&LFSRcolor4[307]&LFSRcolor4[206]&LFSRcolor4[356]);
    BiasedRNG[409] = (LFSRcolor4[329]&LFSRcolor4[348]&LFSRcolor4[222]&LFSRcolor4[145]);
    BiasedRNG[410] = (LFSRcolor4[337]&LFSRcolor4[194]&LFSRcolor4[268]&LFSRcolor4[219]);
    BiasedRNG[411] = (LFSRcolor4[249]&LFSRcolor4[322]&LFSRcolor4[71]&LFSRcolor4[146]);
    BiasedRNG[412] = (LFSRcolor4[65]&LFSRcolor4[361]&LFSRcolor4[351]&LFSRcolor4[202]);
    BiasedRNG[413] = (LFSRcolor4[195]&LFSRcolor4[217]&LFSRcolor4[118]&LFSRcolor4[112]);
    BiasedRNG[414] = (LFSRcolor4[200]&LFSRcolor4[157]&LFSRcolor4[110]&LFSRcolor4[133]);
    BiasedRNG[415] = (LFSRcolor4[215]&LFSRcolor4[308]&LFSRcolor4[235]&LFSRcolor4[314]);
    BiasedRNG[416] = (LFSRcolor4[359]&LFSRcolor4[40]&LFSRcolor4[190]&LFSRcolor4[357]);
    BiasedRNG[417] = (LFSRcolor4[354]&LFSRcolor4[364]&LFSRcolor4[218]&LFSRcolor4[184]);
    BiasedRNG[418] = (LFSRcolor4[213]&LFSRcolor4[99]&LFSRcolor4[28]&LFSRcolor4[33]);
    BiasedRNG[419] = (LFSRcolor4[259]&LFSRcolor4[155]&LFSRcolor4[125]&LFSRcolor4[106]);
    BiasedRNG[420] = (LFSRcolor4[208]&LFSRcolor4[127]&LFSRcolor4[331]&LFSRcolor4[341]);
    BiasedRNG[421] = (LFSRcolor4[363]&LFSRcolor4[227]&LFSRcolor4[148]&LFSRcolor4[286]);
    BiasedRNG[422] = (LFSRcolor4[288]&LFSRcolor4[231]&LFSRcolor4[328]&LFSRcolor4[60]);
    BiasedRNG[423] = (LFSRcolor4[3]&LFSRcolor4[4]&LFSRcolor4[68]&LFSRcolor4[21]);
    BiasedRNG[424] = (LFSRcolor4[152]&LFSRcolor4[278]&LFSRcolor4[88]&LFSRcolor4[362]);
    BiasedRNG[425] = (LFSRcolor4[172]&LFSRcolor4[253]&LFSRcolor4[258]&LFSRcolor4[61]);
    BiasedRNG[426] = (LFSRcolor4[265]&LFSRcolor4[358]&LFSRcolor4[317]&LFSRcolor4[151]);
    BiasedRNG[427] = (LFSRcolor4[186]&LFSRcolor4[94]&LFSRcolor4[316]&LFSRcolor4[179]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule