//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [11:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [229:0] LFSRcolor0;
wire [229:0] LFSRcolor1;
wire [183:0] LFSRcolor2;
wire [45:0] LFSRcolor3;
wire [137:0] LFSRcolor4;
reg [159:0] BiasedRNG;       //For I=+/-1 cases
reg [103:0] UnbiasedRNG;   //For I=0 cases
reg [0:281] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[96] = 1'b1;
initial m[135] = 1'b0;
initial m[145] = 1'b0;
initial m[160] = 1'b0;
initial m[180] = 1'b0;
initial m[205] = 1'b1;
initial m[230] = 1'b0;
initial m[250] = 1'b1;
initial m[265] = 1'b0;
initial m[275] = 1'b0;
initial m[280] = 1'b1;
initial m[281] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[134] = 1'b0;
initial m[144] = 1'b0;
initial m[159] = 1'b0;
initial m[179] = 1'b0;
initial m[204] = 1'b0;
initial m[207] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 1;
initial m[1] = 0;
initial m[2] = 1;
initial m[3] = 0;
initial m[4] = 1;
initial m[5] = 0;
initial m[6] = 0;
initial m[7] = 0;
initial m[8] = 1;
initial m[9] = 0;
initial m[10] = 0;
initial m[11] = 1;
initial m[12] = 0;
initial m[13] = 0;
initial m[14] = 1;
initial m[15] = 1;
initial m[16] = 1;
initial m[17] = 0;
initial m[18] = 1;
initial m[19] = 0;
initial m[20] = 1;
initial m[21] = 0;
initial m[22] = 1;
initial m[23] = 1;
initial m[24] = 0;
initial m[25] = 1;
initial m[26] = 1;
initial m[27] = 0;
initial m[28] = 0;
initial m[29] = 0;
initial m[30] = 1;
initial m[31] = 1;
initial m[32] = 0;
initial m[33] = 0;
initial m[34] = 0;
initial m[35] = 0;
initial m[36] = 0;
initial m[37] = 1;
initial m[38] = 0;
initial m[39] = 1;
initial m[40] = 1;
initial m[41] = 0;
initial m[42] = 0;
initial m[43] = 1;
initial m[44] = 0;
initial m[45] = 1;
initial m[46] = 0;
initial m[47] = 0;
initial m[48] = 0;
initial m[49] = 1;
initial m[50] = 0;
initial m[51] = 0;
initial m[52] = 0;
initial m[53] = 0;
initial m[54] = 1;
initial m[55] = 1;
initial m[56] = 1;
initial m[57] = 0;
initial m[58] = 1;
initial m[59] = 0;
initial m[60] = 0;
initial m[61] = 1;
initial m[62] = 1;
initial m[63] = 1;
initial m[64] = 1;
initial m[65] = 1;
initial m[66] = 1;
initial m[67] = 1;
initial m[68] = 0;
initial m[69] = 0;
initial m[70] = 0;
initial m[71] = 0;
initial m[72] = 0;
initial m[73] = 1;
initial m[74] = 0;
initial m[75] = 0;
initial m[76] = 1;
initial m[77] = 0;
initial m[78] = 1;
initial m[79] = 0;
initial m[80] = 0;
initial m[81] = 1;
initial m[82] = 0;
initial m[83] = 0;
initial m[84] = 0;
initial m[85] = 0;
initial m[86] = 0;
initial m[87] = 0;
initial m[88] = 0;
initial m[89] = 0;
initial m[90] = 1;
initial m[91] = 0;
initial m[92] = 1;
initial m[93] = 0;
initial m[94] = 1;
initial m[95] = 1;
initial m[97] = 0;
initial m[98] = 0;
initial m[99] = 1;
initial m[100] = 0;
initial m[101] = 0;
initial m[102] = 1;
initial m[103] = 1;
initial m[104] = 1;
initial m[105] = 1;
initial m[106] = 0;
initial m[107] = 0;
initial m[108] = 0;
initial m[109] = 1;
initial m[110] = 0;
initial m[111] = 1;
initial m[112] = 1;
initial m[113] = 0;
initial m[114] = 1;
initial m[115] = 1;
initial m[116] = 1;
initial m[117] = 1;
initial m[118] = 1;
initial m[119] = 0;
initial m[120] = 1;
initial m[121] = 1;
initial m[122] = 0;
initial m[123] = 0;
initial m[124] = 0;
initial m[125] = 1;
initial m[126] = 1;
initial m[127] = 1;
initial m[128] = 1;
initial m[129] = 0;
initial m[130] = 1;
initial m[131] = 1;
initial m[132] = 1;
initial m[133] = 1;
initial m[136] = 1;
initial m[137] = 1;
initial m[138] = 0;
initial m[139] = 1;
initial m[140] = 1;
initial m[141] = 1;
initial m[142] = 0;
initial m[143] = 1;
initial m[146] = 0;
initial m[147] = 1;
initial m[148] = 0;
initial m[149] = 0;
initial m[150] = 1;
initial m[151] = 0;
initial m[152] = 1;
initial m[153] = 0;
initial m[154] = 1;
initial m[155] = 0;
initial m[156] = 1;
initial m[157] = 0;
initial m[158] = 1;
initial m[161] = 0;
initial m[162] = 0;
initial m[163] = 1;
initial m[164] = 1;
initial m[165] = 0;
initial m[166] = 0;
initial m[167] = 1;
initial m[168] = 1;
initial m[169] = 0;
initial m[170] = 1;
initial m[171] = 0;
initial m[172] = 1;
initial m[173] = 0;
initial m[174] = 0;
initial m[175] = 1;
initial m[176] = 1;
initial m[177] = 1;
initial m[178] = 0;
initial m[181] = 0;
initial m[182] = 0;
initial m[183] = 0;
initial m[184] = 1;
initial m[185] = 0;
initial m[186] = 1;
initial m[187] = 1;
initial m[188] = 0;
initial m[189] = 0;
initial m[190] = 0;
initial m[191] = 0;
initial m[192] = 0;
initial m[193] = 0;
initial m[194] = 0;
initial m[195] = 1;
initial m[196] = 0;
initial m[197] = 0;
initial m[198] = 0;
initial m[199] = 0;
initial m[200] = 0;
initial m[201] = 1;
initial m[202] = 1;
initial m[203] = 1;
initial m[206] = 1;
initial m[208] = 1;
initial m[209] = 0;
initial m[210] = 1;
initial m[211] = 0;
initial m[212] = 0;
initial m[213] = 0;
initial m[214] = 1;
initial m[215] = 0;
initial m[216] = 1;
initial m[217] = 1;
initial m[218] = 0;
initial m[219] = 0;
initial m[220] = 1;
initial m[221] = 0;
initial m[222] = 1;
initial m[223] = 0;
initial m[224] = 1;
initial m[225] = 1;
initial m[226] = 0;
initial m[227] = 0;
initial m[228] = 1;
initial m[229] = 0;
initial m[231] = 0;
initial m[232] = 1;
initial m[233] = 0;
initial m[234] = 0;
initial m[235] = 0;
initial m[236] = 0;
initial m[237] = 1;
initial m[238] = 1;
initial m[239] = 0;
initial m[240] = 1;
initial m[241] = 0;
initial m[242] = 1;
initial m[243] = 0;
initial m[244] = 1;
initial m[245] = 0;
initial m[246] = 1;
initial m[247] = 0;
initial m[248] = 1;
initial m[249] = 1;
initial m[251] = 0;
initial m[252] = 0;
initial m[253] = 1;
initial m[254] = 1;
initial m[255] = 1;
initial m[256] = 1;
initial m[257] = 1;
initial m[258] = 0;
initial m[259] = 1;
initial m[260] = 1;
initial m[261] = 0;
initial m[262] = 0;
initial m[263] = 1;
initial m[264] = 0;
initial m[266] = 1;
initial m[267] = 1;
initial m[268] = 1;
initial m[269] = 0;
initial m[270] = 1;
initial m[271] = 1;
initial m[272] = 1;
initial m[273] = 0;
initial m[274] = 1;
initial m[276] = 1;
initial m[277] = 0;
initial m[278] = 0;
initial m[279] = 1;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[5],m[4],m[3],m[2],m[1],m[0]}*{m[11],m[10],m[9],m[8],m[7],m[6]};
end

always @(negedge sample_clk) begin
    if (solution == 12'b110010100001)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[12]&~m[24]&~m[25])|(~m[12]&m[24]&~m[25])|(~m[12]&~m[24]&m[25]))&BiasedRNG[0])|(((m[12]&m[24]&~m[25])|(m[12]&~m[24]&m[25])|(~m[12]&m[24]&m[25]))&~BiasedRNG[0])|((m[12]&m[24]&m[25]));
    m[1] = (((m[13]&~m[30]&~m[31])|(~m[13]&m[30]&~m[31])|(~m[13]&~m[30]&m[31]))&BiasedRNG[1])|(((m[13]&m[30]&~m[31])|(m[13]&~m[30]&m[31])|(~m[13]&m[30]&m[31]))&~BiasedRNG[1])|((m[13]&m[30]&m[31]));
    m[2] = (((m[14]&~m[36]&~m[37])|(~m[14]&m[36]&~m[37])|(~m[14]&~m[36]&m[37]))&BiasedRNG[2])|(((m[14]&m[36]&~m[37])|(m[14]&~m[36]&m[37])|(~m[14]&m[36]&m[37]))&~BiasedRNG[2])|((m[14]&m[36]&m[37]));
    m[3] = (((m[15]&~m[42]&~m[43])|(~m[15]&m[42]&~m[43])|(~m[15]&~m[42]&m[43]))&BiasedRNG[3])|(((m[15]&m[42]&~m[43])|(m[15]&~m[42]&m[43])|(~m[15]&m[42]&m[43]))&~BiasedRNG[3])|((m[15]&m[42]&m[43]));
    m[4] = (((m[16]&~m[48]&~m[49])|(~m[16]&m[48]&~m[49])|(~m[16]&~m[48]&m[49]))&BiasedRNG[4])|(((m[16]&m[48]&~m[49])|(m[16]&~m[48]&m[49])|(~m[16]&m[48]&m[49]))&~BiasedRNG[4])|((m[16]&m[48]&m[49]));
    m[5] = (((m[17]&~m[54]&~m[55])|(~m[17]&m[54]&~m[55])|(~m[17]&~m[54]&m[55]))&BiasedRNG[5])|(((m[17]&m[54]&~m[55])|(m[17]&~m[54]&m[55])|(~m[17]&m[54]&m[55]))&~BiasedRNG[5])|((m[17]&m[54]&m[55]));
    m[6] = (((m[18]&~m[60]&~m[61])|(~m[18]&m[60]&~m[61])|(~m[18]&~m[60]&m[61]))&BiasedRNG[6])|(((m[18]&m[60]&~m[61])|(m[18]&~m[60]&m[61])|(~m[18]&m[60]&m[61]))&~BiasedRNG[6])|((m[18]&m[60]&m[61]));
    m[7] = (((m[19]&~m[66]&~m[67])|(~m[19]&m[66]&~m[67])|(~m[19]&~m[66]&m[67]))&BiasedRNG[7])|(((m[19]&m[66]&~m[67])|(m[19]&~m[66]&m[67])|(~m[19]&m[66]&m[67]))&~BiasedRNG[7])|((m[19]&m[66]&m[67]));
    m[8] = (((m[20]&~m[72]&~m[73])|(~m[20]&m[72]&~m[73])|(~m[20]&~m[72]&m[73]))&BiasedRNG[8])|(((m[20]&m[72]&~m[73])|(m[20]&~m[72]&m[73])|(~m[20]&m[72]&m[73]))&~BiasedRNG[8])|((m[20]&m[72]&m[73]));
    m[9] = (((m[21]&~m[78]&~m[79])|(~m[21]&m[78]&~m[79])|(~m[21]&~m[78]&m[79]))&BiasedRNG[9])|(((m[21]&m[78]&~m[79])|(m[21]&~m[78]&m[79])|(~m[21]&m[78]&m[79]))&~BiasedRNG[9])|((m[21]&m[78]&m[79]));
    m[10] = (((m[22]&~m[84]&~m[85])|(~m[22]&m[84]&~m[85])|(~m[22]&~m[84]&m[85]))&BiasedRNG[10])|(((m[22]&m[84]&~m[85])|(m[22]&~m[84]&m[85])|(~m[22]&m[84]&m[85]))&~BiasedRNG[10])|((m[22]&m[84]&m[85]));
    m[11] = (((m[23]&~m[90]&~m[91])|(~m[23]&m[90]&~m[91])|(~m[23]&~m[90]&m[91]))&BiasedRNG[11])|(((m[23]&m[90]&~m[91])|(m[23]&~m[90]&m[91])|(~m[23]&m[90]&m[91]))&~BiasedRNG[11])|((m[23]&m[90]&m[91]));
    m[26] = (((~m[12]&~m[72]&~m[108])|(m[12]&m[72]&~m[108]))&BiasedRNG[12])|(((m[12]&~m[72]&~m[108])|(~m[12]&m[72]&m[108]))&~BiasedRNG[12])|((~m[12]&~m[72]&m[108])|(m[12]&~m[72]&m[108])|(m[12]&m[72]&m[108]));
    m[27] = (((~m[12]&~m[78]&~m[114])|(m[12]&m[78]&~m[114]))&BiasedRNG[13])|(((m[12]&~m[78]&~m[114])|(~m[12]&m[78]&m[114]))&~BiasedRNG[13])|((~m[12]&~m[78]&m[114])|(m[12]&~m[78]&m[114])|(m[12]&m[78]&m[114]));
    m[28] = (((~m[12]&~m[84]&~m[120])|(m[12]&m[84]&~m[120]))&BiasedRNG[14])|(((m[12]&~m[84]&~m[120])|(~m[12]&m[84]&m[120]))&~BiasedRNG[14])|((~m[12]&~m[84]&m[120])|(m[12]&~m[84]&m[120])|(m[12]&m[84]&m[120]));
    m[29] = (((~m[12]&~m[90]&~m[126])|(m[12]&m[90]&~m[126]))&BiasedRNG[15])|(((m[12]&~m[90]&~m[126])|(~m[12]&m[90]&m[126]))&~BiasedRNG[15])|((~m[12]&~m[90]&m[126])|(m[12]&~m[90]&m[126])|(m[12]&m[90]&m[126]));
    m[32] = (((~m[13]&~m[73]&~m[109])|(m[13]&m[73]&~m[109]))&BiasedRNG[16])|(((m[13]&~m[73]&~m[109])|(~m[13]&m[73]&m[109]))&~BiasedRNG[16])|((~m[13]&~m[73]&m[109])|(m[13]&~m[73]&m[109])|(m[13]&m[73]&m[109]));
    m[33] = (((~m[13]&~m[79]&~m[115])|(m[13]&m[79]&~m[115]))&BiasedRNG[17])|(((m[13]&~m[79]&~m[115])|(~m[13]&m[79]&m[115]))&~BiasedRNG[17])|((~m[13]&~m[79]&m[115])|(m[13]&~m[79]&m[115])|(m[13]&m[79]&m[115]));
    m[34] = (((~m[13]&~m[85]&~m[121])|(m[13]&m[85]&~m[121]))&BiasedRNG[18])|(((m[13]&~m[85]&~m[121])|(~m[13]&m[85]&m[121]))&~BiasedRNG[18])|((~m[13]&~m[85]&m[121])|(m[13]&~m[85]&m[121])|(m[13]&m[85]&m[121]));
    m[35] = (((~m[13]&~m[91]&~m[127])|(m[13]&m[91]&~m[127]))&BiasedRNG[19])|(((m[13]&~m[91]&~m[127])|(~m[13]&m[91]&m[127]))&~BiasedRNG[19])|((~m[13]&~m[91]&m[127])|(m[13]&~m[91]&m[127])|(m[13]&m[91]&m[127]));
    m[38] = (((~m[14]&~m[74]&~m[110])|(m[14]&m[74]&~m[110]))&BiasedRNG[20])|(((m[14]&~m[74]&~m[110])|(~m[14]&m[74]&m[110]))&~BiasedRNG[20])|((~m[14]&~m[74]&m[110])|(m[14]&~m[74]&m[110])|(m[14]&m[74]&m[110]));
    m[39] = (((~m[14]&~m[80]&~m[116])|(m[14]&m[80]&~m[116]))&BiasedRNG[21])|(((m[14]&~m[80]&~m[116])|(~m[14]&m[80]&m[116]))&~BiasedRNG[21])|((~m[14]&~m[80]&m[116])|(m[14]&~m[80]&m[116])|(m[14]&m[80]&m[116]));
    m[40] = (((~m[14]&~m[86]&~m[122])|(m[14]&m[86]&~m[122]))&BiasedRNG[22])|(((m[14]&~m[86]&~m[122])|(~m[14]&m[86]&m[122]))&~BiasedRNG[22])|((~m[14]&~m[86]&m[122])|(m[14]&~m[86]&m[122])|(m[14]&m[86]&m[122]));
    m[41] = (((~m[14]&~m[92]&~m[128])|(m[14]&m[92]&~m[128]))&BiasedRNG[23])|(((m[14]&~m[92]&~m[128])|(~m[14]&m[92]&m[128]))&~BiasedRNG[23])|((~m[14]&~m[92]&m[128])|(m[14]&~m[92]&m[128])|(m[14]&m[92]&m[128]));
    m[44] = (((~m[15]&~m[75]&~m[111])|(m[15]&m[75]&~m[111]))&BiasedRNG[24])|(((m[15]&~m[75]&~m[111])|(~m[15]&m[75]&m[111]))&~BiasedRNG[24])|((~m[15]&~m[75]&m[111])|(m[15]&~m[75]&m[111])|(m[15]&m[75]&m[111]));
    m[45] = (((~m[15]&~m[81]&~m[117])|(m[15]&m[81]&~m[117]))&BiasedRNG[25])|(((m[15]&~m[81]&~m[117])|(~m[15]&m[81]&m[117]))&~BiasedRNG[25])|((~m[15]&~m[81]&m[117])|(m[15]&~m[81]&m[117])|(m[15]&m[81]&m[117]));
    m[46] = (((~m[15]&~m[87]&~m[123])|(m[15]&m[87]&~m[123]))&BiasedRNG[26])|(((m[15]&~m[87]&~m[123])|(~m[15]&m[87]&m[123]))&~BiasedRNG[26])|((~m[15]&~m[87]&m[123])|(m[15]&~m[87]&m[123])|(m[15]&m[87]&m[123]));
    m[47] = (((~m[15]&~m[93]&~m[129])|(m[15]&m[93]&~m[129]))&BiasedRNG[27])|(((m[15]&~m[93]&~m[129])|(~m[15]&m[93]&m[129]))&~BiasedRNG[27])|((~m[15]&~m[93]&m[129])|(m[15]&~m[93]&m[129])|(m[15]&m[93]&m[129]));
    m[50] = (((~m[16]&~m[76]&~m[112])|(m[16]&m[76]&~m[112]))&BiasedRNG[28])|(((m[16]&~m[76]&~m[112])|(~m[16]&m[76]&m[112]))&~BiasedRNG[28])|((~m[16]&~m[76]&m[112])|(m[16]&~m[76]&m[112])|(m[16]&m[76]&m[112]));
    m[51] = (((~m[16]&~m[82]&~m[118])|(m[16]&m[82]&~m[118]))&BiasedRNG[29])|(((m[16]&~m[82]&~m[118])|(~m[16]&m[82]&m[118]))&~BiasedRNG[29])|((~m[16]&~m[82]&m[118])|(m[16]&~m[82]&m[118])|(m[16]&m[82]&m[118]));
    m[52] = (((~m[16]&~m[88]&~m[124])|(m[16]&m[88]&~m[124]))&BiasedRNG[30])|(((m[16]&~m[88]&~m[124])|(~m[16]&m[88]&m[124]))&~BiasedRNG[30])|((~m[16]&~m[88]&m[124])|(m[16]&~m[88]&m[124])|(m[16]&m[88]&m[124]));
    m[53] = (((~m[16]&~m[94]&~m[130])|(m[16]&m[94]&~m[130]))&BiasedRNG[31])|(((m[16]&~m[94]&~m[130])|(~m[16]&m[94]&m[130]))&~BiasedRNG[31])|((~m[16]&~m[94]&m[130])|(m[16]&~m[94]&m[130])|(m[16]&m[94]&m[130]));
    m[56] = (((~m[17]&~m[77]&~m[113])|(m[17]&m[77]&~m[113]))&BiasedRNG[32])|(((m[17]&~m[77]&~m[113])|(~m[17]&m[77]&m[113]))&~BiasedRNG[32])|((~m[17]&~m[77]&m[113])|(m[17]&~m[77]&m[113])|(m[17]&m[77]&m[113]));
    m[57] = (((~m[17]&~m[83]&~m[119])|(m[17]&m[83]&~m[119]))&BiasedRNG[33])|(((m[17]&~m[83]&~m[119])|(~m[17]&m[83]&m[119]))&~BiasedRNG[33])|((~m[17]&~m[83]&m[119])|(m[17]&~m[83]&m[119])|(m[17]&m[83]&m[119]));
    m[58] = (((~m[17]&~m[89]&~m[125])|(m[17]&m[89]&~m[125]))&BiasedRNG[34])|(((m[17]&~m[89]&~m[125])|(~m[17]&m[89]&m[125]))&~BiasedRNG[34])|((~m[17]&~m[89]&m[125])|(m[17]&~m[89]&m[125])|(m[17]&m[89]&m[125]));
    m[59] = (((~m[17]&~m[95]&~m[131])|(m[17]&m[95]&~m[131]))&BiasedRNG[35])|(((m[17]&~m[95]&~m[131])|(~m[17]&m[95]&m[131]))&~BiasedRNG[35])|((~m[17]&~m[95]&m[131])|(m[17]&~m[95]&m[131])|(m[17]&m[95]&m[131]));
    m[62] = (((~m[18]&~m[36]&~m[98])|(m[18]&m[36]&~m[98]))&BiasedRNG[36])|(((m[18]&~m[36]&~m[98])|(~m[18]&m[36]&m[98]))&~BiasedRNG[36])|((~m[18]&~m[36]&m[98])|(m[18]&~m[36]&m[98])|(m[18]&m[36]&m[98]));
    m[63] = (((~m[18]&~m[42]&~m[99])|(m[18]&m[42]&~m[99]))&BiasedRNG[37])|(((m[18]&~m[42]&~m[99])|(~m[18]&m[42]&m[99]))&~BiasedRNG[37])|((~m[18]&~m[42]&m[99])|(m[18]&~m[42]&m[99])|(m[18]&m[42]&m[99]));
    m[64] = (((~m[18]&~m[48]&~m[100])|(m[18]&m[48]&~m[100]))&BiasedRNG[38])|(((m[18]&~m[48]&~m[100])|(~m[18]&m[48]&m[100]))&~BiasedRNG[38])|((~m[18]&~m[48]&m[100])|(m[18]&~m[48]&m[100])|(m[18]&m[48]&m[100]));
    m[65] = (((~m[18]&~m[54]&~m[101])|(m[18]&m[54]&~m[101]))&BiasedRNG[39])|(((m[18]&~m[54]&~m[101])|(~m[18]&m[54]&m[101]))&~BiasedRNG[39])|((~m[18]&~m[54]&m[101])|(m[18]&~m[54]&m[101])|(m[18]&m[54]&m[101]));
    m[68] = (((~m[19]&~m[37]&~m[104])|(m[19]&m[37]&~m[104]))&BiasedRNG[40])|(((m[19]&~m[37]&~m[104])|(~m[19]&m[37]&m[104]))&~BiasedRNG[40])|((~m[19]&~m[37]&m[104])|(m[19]&~m[37]&m[104])|(m[19]&m[37]&m[104]));
    m[69] = (((~m[19]&~m[43]&~m[105])|(m[19]&m[43]&~m[105]))&BiasedRNG[41])|(((m[19]&~m[43]&~m[105])|(~m[19]&m[43]&m[105]))&~BiasedRNG[41])|((~m[19]&~m[43]&m[105])|(m[19]&~m[43]&m[105])|(m[19]&m[43]&m[105]));
    m[70] = (((~m[19]&~m[49]&~m[106])|(m[19]&m[49]&~m[106]))&BiasedRNG[42])|(((m[19]&~m[49]&~m[106])|(~m[19]&m[49]&m[106]))&~BiasedRNG[42])|((~m[19]&~m[49]&m[106])|(m[19]&~m[49]&m[106])|(m[19]&m[49]&m[106]));
    m[71] = (((~m[19]&~m[55]&~m[107])|(m[19]&m[55]&~m[107]))&BiasedRNG[43])|(((m[19]&~m[55]&~m[107])|(~m[19]&m[55]&m[107]))&~BiasedRNG[43])|((~m[19]&~m[55]&m[107])|(m[19]&~m[55]&m[107])|(m[19]&m[55]&m[107]));
    m[97] = (((m[30]&~m[61]&m[132])|(~m[30]&m[61]&m[132]))&BiasedRNG[44])|(((m[30]&m[61]&~m[132]))&~BiasedRNG[44])|((m[30]&m[61]&m[132]));
    m[102] = (((m[25]&~m[66]&m[133])|(~m[25]&m[66]&m[133]))&BiasedRNG[45])|(((m[25]&m[66]&~m[133]))&~BiasedRNG[45])|((m[25]&m[66]&m[133]));
    m[103] = (((m[31]&~m[67]&m[138])|(~m[31]&m[67]&m[138]))&BiasedRNG[46])|(((m[31]&m[67]&~m[138]))&~BiasedRNG[46])|((m[31]&m[67]&m[138]));
    m[137] = (((m[98]&~m[138]&~m[139]&~m[140]&~m[141])|(~m[98]&~m[138]&~m[139]&m[140]&~m[141])|(m[98]&m[138]&~m[139]&m[140]&~m[141])|(m[98]&~m[138]&m[139]&m[140]&~m[141])|(~m[98]&m[138]&~m[139]&~m[140]&m[141])|(~m[98]&~m[138]&m[139]&~m[140]&m[141])|(m[98]&m[138]&m[139]&~m[140]&m[141])|(~m[98]&m[138]&m[139]&m[140]&m[141]))&UnbiasedRNG[0])|((m[98]&~m[138]&~m[139]&m[140]&~m[141])|(~m[98]&~m[138]&~m[139]&~m[140]&m[141])|(m[98]&~m[138]&~m[139]&~m[140]&m[141])|(m[98]&m[138]&~m[139]&~m[140]&m[141])|(m[98]&~m[138]&m[139]&~m[140]&m[141])|(~m[98]&~m[138]&~m[139]&m[140]&m[141])|(m[98]&~m[138]&~m[139]&m[140]&m[141])|(~m[98]&m[138]&~m[139]&m[140]&m[141])|(m[98]&m[138]&~m[139]&m[140]&m[141])|(~m[98]&~m[138]&m[139]&m[140]&m[141])|(m[98]&~m[138]&m[139]&m[140]&m[141])|(m[98]&m[138]&m[139]&m[140]&m[141]));
    m[142] = (((m[140]&~m[143]&~m[144]&~m[145]&~m[146])|(~m[140]&~m[143]&~m[144]&m[145]&~m[146])|(m[140]&m[143]&~m[144]&m[145]&~m[146])|(m[140]&~m[143]&m[144]&m[145]&~m[146])|(~m[140]&m[143]&~m[144]&~m[145]&m[146])|(~m[140]&~m[143]&m[144]&~m[145]&m[146])|(m[140]&m[143]&m[144]&~m[145]&m[146])|(~m[140]&m[143]&m[144]&m[145]&m[146]))&UnbiasedRNG[1])|((m[140]&~m[143]&~m[144]&m[145]&~m[146])|(~m[140]&~m[143]&~m[144]&~m[145]&m[146])|(m[140]&~m[143]&~m[144]&~m[145]&m[146])|(m[140]&m[143]&~m[144]&~m[145]&m[146])|(m[140]&~m[143]&m[144]&~m[145]&m[146])|(~m[140]&~m[143]&~m[144]&m[145]&m[146])|(m[140]&~m[143]&~m[144]&m[145]&m[146])|(~m[140]&m[143]&~m[144]&m[145]&m[146])|(m[140]&m[143]&~m[144]&m[145]&m[146])|(~m[140]&~m[143]&m[144]&m[145]&m[146])|(m[140]&~m[143]&m[144]&m[145]&m[146])|(m[140]&m[143]&m[144]&m[145]&m[146]));
    m[147] = (((m[99]&~m[148]&~m[149]&~m[150]&~m[151])|(~m[99]&~m[148]&~m[149]&m[150]&~m[151])|(m[99]&m[148]&~m[149]&m[150]&~m[151])|(m[99]&~m[148]&m[149]&m[150]&~m[151])|(~m[99]&m[148]&~m[149]&~m[150]&m[151])|(~m[99]&~m[148]&m[149]&~m[150]&m[151])|(m[99]&m[148]&m[149]&~m[150]&m[151])|(~m[99]&m[148]&m[149]&m[150]&m[151]))&UnbiasedRNG[2])|((m[99]&~m[148]&~m[149]&m[150]&~m[151])|(~m[99]&~m[148]&~m[149]&~m[150]&m[151])|(m[99]&~m[148]&~m[149]&~m[150]&m[151])|(m[99]&m[148]&~m[149]&~m[150]&m[151])|(m[99]&~m[148]&m[149]&~m[150]&m[151])|(~m[99]&~m[148]&~m[149]&m[150]&m[151])|(m[99]&~m[148]&~m[149]&m[150]&m[151])|(~m[99]&m[148]&~m[149]&m[150]&m[151])|(m[99]&m[148]&~m[149]&m[150]&m[151])|(~m[99]&~m[148]&m[149]&m[150]&m[151])|(m[99]&~m[148]&m[149]&m[150]&m[151])|(m[99]&m[148]&m[149]&m[150]&m[151]));
    m[152] = (((m[150]&~m[153]&~m[154]&~m[155]&~m[156])|(~m[150]&~m[153]&~m[154]&m[155]&~m[156])|(m[150]&m[153]&~m[154]&m[155]&~m[156])|(m[150]&~m[153]&m[154]&m[155]&~m[156])|(~m[150]&m[153]&~m[154]&~m[155]&m[156])|(~m[150]&~m[153]&m[154]&~m[155]&m[156])|(m[150]&m[153]&m[154]&~m[155]&m[156])|(~m[150]&m[153]&m[154]&m[155]&m[156]))&UnbiasedRNG[3])|((m[150]&~m[153]&~m[154]&m[155]&~m[156])|(~m[150]&~m[153]&~m[154]&~m[155]&m[156])|(m[150]&~m[153]&~m[154]&~m[155]&m[156])|(m[150]&m[153]&~m[154]&~m[155]&m[156])|(m[150]&~m[153]&m[154]&~m[155]&m[156])|(~m[150]&~m[153]&~m[154]&m[155]&m[156])|(m[150]&~m[153]&~m[154]&m[155]&m[156])|(~m[150]&m[153]&~m[154]&m[155]&m[156])|(m[150]&m[153]&~m[154]&m[155]&m[156])|(~m[150]&~m[153]&m[154]&m[155]&m[156])|(m[150]&~m[153]&m[154]&m[155]&m[156])|(m[150]&m[153]&m[154]&m[155]&m[156]));
    m[157] = (((m[155]&~m[158]&~m[159]&~m[160]&~m[161])|(~m[155]&~m[158]&~m[159]&m[160]&~m[161])|(m[155]&m[158]&~m[159]&m[160]&~m[161])|(m[155]&~m[158]&m[159]&m[160]&~m[161])|(~m[155]&m[158]&~m[159]&~m[160]&m[161])|(~m[155]&~m[158]&m[159]&~m[160]&m[161])|(m[155]&m[158]&m[159]&~m[160]&m[161])|(~m[155]&m[158]&m[159]&m[160]&m[161]))&UnbiasedRNG[4])|((m[155]&~m[158]&~m[159]&m[160]&~m[161])|(~m[155]&~m[158]&~m[159]&~m[160]&m[161])|(m[155]&~m[158]&~m[159]&~m[160]&m[161])|(m[155]&m[158]&~m[159]&~m[160]&m[161])|(m[155]&~m[158]&m[159]&~m[160]&m[161])|(~m[155]&~m[158]&~m[159]&m[160]&m[161])|(m[155]&~m[158]&~m[159]&m[160]&m[161])|(~m[155]&m[158]&~m[159]&m[160]&m[161])|(m[155]&m[158]&~m[159]&m[160]&m[161])|(~m[155]&~m[158]&m[159]&m[160]&m[161])|(m[155]&~m[158]&m[159]&m[160]&m[161])|(m[155]&m[158]&m[159]&m[160]&m[161]));
    m[162] = (((m[100]&~m[163]&~m[164]&~m[165]&~m[166])|(~m[100]&~m[163]&~m[164]&m[165]&~m[166])|(m[100]&m[163]&~m[164]&m[165]&~m[166])|(m[100]&~m[163]&m[164]&m[165]&~m[166])|(~m[100]&m[163]&~m[164]&~m[165]&m[166])|(~m[100]&~m[163]&m[164]&~m[165]&m[166])|(m[100]&m[163]&m[164]&~m[165]&m[166])|(~m[100]&m[163]&m[164]&m[165]&m[166]))&UnbiasedRNG[5])|((m[100]&~m[163]&~m[164]&m[165]&~m[166])|(~m[100]&~m[163]&~m[164]&~m[165]&m[166])|(m[100]&~m[163]&~m[164]&~m[165]&m[166])|(m[100]&m[163]&~m[164]&~m[165]&m[166])|(m[100]&~m[163]&m[164]&~m[165]&m[166])|(~m[100]&~m[163]&~m[164]&m[165]&m[166])|(m[100]&~m[163]&~m[164]&m[165]&m[166])|(~m[100]&m[163]&~m[164]&m[165]&m[166])|(m[100]&m[163]&~m[164]&m[165]&m[166])|(~m[100]&~m[163]&m[164]&m[165]&m[166])|(m[100]&~m[163]&m[164]&m[165]&m[166])|(m[100]&m[163]&m[164]&m[165]&m[166]));
    m[167] = (((m[165]&~m[168]&~m[169]&~m[170]&~m[171])|(~m[165]&~m[168]&~m[169]&m[170]&~m[171])|(m[165]&m[168]&~m[169]&m[170]&~m[171])|(m[165]&~m[168]&m[169]&m[170]&~m[171])|(~m[165]&m[168]&~m[169]&~m[170]&m[171])|(~m[165]&~m[168]&m[169]&~m[170]&m[171])|(m[165]&m[168]&m[169]&~m[170]&m[171])|(~m[165]&m[168]&m[169]&m[170]&m[171]))&UnbiasedRNG[6])|((m[165]&~m[168]&~m[169]&m[170]&~m[171])|(~m[165]&~m[168]&~m[169]&~m[170]&m[171])|(m[165]&~m[168]&~m[169]&~m[170]&m[171])|(m[165]&m[168]&~m[169]&~m[170]&m[171])|(m[165]&~m[168]&m[169]&~m[170]&m[171])|(~m[165]&~m[168]&~m[169]&m[170]&m[171])|(m[165]&~m[168]&~m[169]&m[170]&m[171])|(~m[165]&m[168]&~m[169]&m[170]&m[171])|(m[165]&m[168]&~m[169]&m[170]&m[171])|(~m[165]&~m[168]&m[169]&m[170]&m[171])|(m[165]&~m[168]&m[169]&m[170]&m[171])|(m[165]&m[168]&m[169]&m[170]&m[171]));
    m[172] = (((m[170]&~m[173]&~m[174]&~m[175]&~m[176])|(~m[170]&~m[173]&~m[174]&m[175]&~m[176])|(m[170]&m[173]&~m[174]&m[175]&~m[176])|(m[170]&~m[173]&m[174]&m[175]&~m[176])|(~m[170]&m[173]&~m[174]&~m[175]&m[176])|(~m[170]&~m[173]&m[174]&~m[175]&m[176])|(m[170]&m[173]&m[174]&~m[175]&m[176])|(~m[170]&m[173]&m[174]&m[175]&m[176]))&UnbiasedRNG[7])|((m[170]&~m[173]&~m[174]&m[175]&~m[176])|(~m[170]&~m[173]&~m[174]&~m[175]&m[176])|(m[170]&~m[173]&~m[174]&~m[175]&m[176])|(m[170]&m[173]&~m[174]&~m[175]&m[176])|(m[170]&~m[173]&m[174]&~m[175]&m[176])|(~m[170]&~m[173]&~m[174]&m[175]&m[176])|(m[170]&~m[173]&~m[174]&m[175]&m[176])|(~m[170]&m[173]&~m[174]&m[175]&m[176])|(m[170]&m[173]&~m[174]&m[175]&m[176])|(~m[170]&~m[173]&m[174]&m[175]&m[176])|(m[170]&~m[173]&m[174]&m[175]&m[176])|(m[170]&m[173]&m[174]&m[175]&m[176]));
    m[177] = (((m[175]&~m[178]&~m[179]&~m[180]&~m[181])|(~m[175]&~m[178]&~m[179]&m[180]&~m[181])|(m[175]&m[178]&~m[179]&m[180]&~m[181])|(m[175]&~m[178]&m[179]&m[180]&~m[181])|(~m[175]&m[178]&~m[179]&~m[180]&m[181])|(~m[175]&~m[178]&m[179]&~m[180]&m[181])|(m[175]&m[178]&m[179]&~m[180]&m[181])|(~m[175]&m[178]&m[179]&m[180]&m[181]))&UnbiasedRNG[8])|((m[175]&~m[178]&~m[179]&m[180]&~m[181])|(~m[175]&~m[178]&~m[179]&~m[180]&m[181])|(m[175]&~m[178]&~m[179]&~m[180]&m[181])|(m[175]&m[178]&~m[179]&~m[180]&m[181])|(m[175]&~m[178]&m[179]&~m[180]&m[181])|(~m[175]&~m[178]&~m[179]&m[180]&m[181])|(m[175]&~m[178]&~m[179]&m[180]&m[181])|(~m[175]&m[178]&~m[179]&m[180]&m[181])|(m[175]&m[178]&~m[179]&m[180]&m[181])|(~m[175]&~m[178]&m[179]&m[180]&m[181])|(m[175]&~m[178]&m[179]&m[180]&m[181])|(m[175]&m[178]&m[179]&m[180]&m[181]));
    m[182] = (((m[101]&~m[183]&~m[184]&~m[185]&~m[186])|(~m[101]&~m[183]&~m[184]&m[185]&~m[186])|(m[101]&m[183]&~m[184]&m[185]&~m[186])|(m[101]&~m[183]&m[184]&m[185]&~m[186])|(~m[101]&m[183]&~m[184]&~m[185]&m[186])|(~m[101]&~m[183]&m[184]&~m[185]&m[186])|(m[101]&m[183]&m[184]&~m[185]&m[186])|(~m[101]&m[183]&m[184]&m[185]&m[186]))&UnbiasedRNG[9])|((m[101]&~m[183]&~m[184]&m[185]&~m[186])|(~m[101]&~m[183]&~m[184]&~m[185]&m[186])|(m[101]&~m[183]&~m[184]&~m[185]&m[186])|(m[101]&m[183]&~m[184]&~m[185]&m[186])|(m[101]&~m[183]&m[184]&~m[185]&m[186])|(~m[101]&~m[183]&~m[184]&m[185]&m[186])|(m[101]&~m[183]&~m[184]&m[185]&m[186])|(~m[101]&m[183]&~m[184]&m[185]&m[186])|(m[101]&m[183]&~m[184]&m[185]&m[186])|(~m[101]&~m[183]&m[184]&m[185]&m[186])|(m[101]&~m[183]&m[184]&m[185]&m[186])|(m[101]&m[183]&m[184]&m[185]&m[186]));
    m[187] = (((m[185]&~m[188]&~m[189]&~m[190]&~m[191])|(~m[185]&~m[188]&~m[189]&m[190]&~m[191])|(m[185]&m[188]&~m[189]&m[190]&~m[191])|(m[185]&~m[188]&m[189]&m[190]&~m[191])|(~m[185]&m[188]&~m[189]&~m[190]&m[191])|(~m[185]&~m[188]&m[189]&~m[190]&m[191])|(m[185]&m[188]&m[189]&~m[190]&m[191])|(~m[185]&m[188]&m[189]&m[190]&m[191]))&UnbiasedRNG[10])|((m[185]&~m[188]&~m[189]&m[190]&~m[191])|(~m[185]&~m[188]&~m[189]&~m[190]&m[191])|(m[185]&~m[188]&~m[189]&~m[190]&m[191])|(m[185]&m[188]&~m[189]&~m[190]&m[191])|(m[185]&~m[188]&m[189]&~m[190]&m[191])|(~m[185]&~m[188]&~m[189]&m[190]&m[191])|(m[185]&~m[188]&~m[189]&m[190]&m[191])|(~m[185]&m[188]&~m[189]&m[190]&m[191])|(m[185]&m[188]&~m[189]&m[190]&m[191])|(~m[185]&~m[188]&m[189]&m[190]&m[191])|(m[185]&~m[188]&m[189]&m[190]&m[191])|(m[185]&m[188]&m[189]&m[190]&m[191]));
    m[192] = (((m[190]&~m[193]&~m[194]&~m[195]&~m[196])|(~m[190]&~m[193]&~m[194]&m[195]&~m[196])|(m[190]&m[193]&~m[194]&m[195]&~m[196])|(m[190]&~m[193]&m[194]&m[195]&~m[196])|(~m[190]&m[193]&~m[194]&~m[195]&m[196])|(~m[190]&~m[193]&m[194]&~m[195]&m[196])|(m[190]&m[193]&m[194]&~m[195]&m[196])|(~m[190]&m[193]&m[194]&m[195]&m[196]))&UnbiasedRNG[11])|((m[190]&~m[193]&~m[194]&m[195]&~m[196])|(~m[190]&~m[193]&~m[194]&~m[195]&m[196])|(m[190]&~m[193]&~m[194]&~m[195]&m[196])|(m[190]&m[193]&~m[194]&~m[195]&m[196])|(m[190]&~m[193]&m[194]&~m[195]&m[196])|(~m[190]&~m[193]&~m[194]&m[195]&m[196])|(m[190]&~m[193]&~m[194]&m[195]&m[196])|(~m[190]&m[193]&~m[194]&m[195]&m[196])|(m[190]&m[193]&~m[194]&m[195]&m[196])|(~m[190]&~m[193]&m[194]&m[195]&m[196])|(m[190]&~m[193]&m[194]&m[195]&m[196])|(m[190]&m[193]&m[194]&m[195]&m[196]));
    m[197] = (((m[195]&~m[198]&~m[199]&~m[200]&~m[201])|(~m[195]&~m[198]&~m[199]&m[200]&~m[201])|(m[195]&m[198]&~m[199]&m[200]&~m[201])|(m[195]&~m[198]&m[199]&m[200]&~m[201])|(~m[195]&m[198]&~m[199]&~m[200]&m[201])|(~m[195]&~m[198]&m[199]&~m[200]&m[201])|(m[195]&m[198]&m[199]&~m[200]&m[201])|(~m[195]&m[198]&m[199]&m[200]&m[201]))&UnbiasedRNG[12])|((m[195]&~m[198]&~m[199]&m[200]&~m[201])|(~m[195]&~m[198]&~m[199]&~m[200]&m[201])|(m[195]&~m[198]&~m[199]&~m[200]&m[201])|(m[195]&m[198]&~m[199]&~m[200]&m[201])|(m[195]&~m[198]&m[199]&~m[200]&m[201])|(~m[195]&~m[198]&~m[199]&m[200]&m[201])|(m[195]&~m[198]&~m[199]&m[200]&m[201])|(~m[195]&m[198]&~m[199]&m[200]&m[201])|(m[195]&m[198]&~m[199]&m[200]&m[201])|(~m[195]&~m[198]&m[199]&m[200]&m[201])|(m[195]&~m[198]&m[199]&m[200]&m[201])|(m[195]&m[198]&m[199]&m[200]&m[201]));
    m[202] = (((m[200]&~m[203]&~m[204]&~m[205]&~m[206])|(~m[200]&~m[203]&~m[204]&m[205]&~m[206])|(m[200]&m[203]&~m[204]&m[205]&~m[206])|(m[200]&~m[203]&m[204]&m[205]&~m[206])|(~m[200]&m[203]&~m[204]&~m[205]&m[206])|(~m[200]&~m[203]&m[204]&~m[205]&m[206])|(m[200]&m[203]&m[204]&~m[205]&m[206])|(~m[200]&m[203]&m[204]&m[205]&m[206]))&UnbiasedRNG[13])|((m[200]&~m[203]&~m[204]&m[205]&~m[206])|(~m[200]&~m[203]&~m[204]&~m[205]&m[206])|(m[200]&~m[203]&~m[204]&~m[205]&m[206])|(m[200]&m[203]&~m[204]&~m[205]&m[206])|(m[200]&~m[203]&m[204]&~m[205]&m[206])|(~m[200]&~m[203]&~m[204]&m[205]&m[206])|(m[200]&~m[203]&~m[204]&m[205]&m[206])|(~m[200]&m[203]&~m[204]&m[205]&m[206])|(m[200]&m[203]&~m[204]&m[205]&m[206])|(~m[200]&~m[203]&m[204]&m[205]&m[206])|(m[200]&~m[203]&m[204]&m[205]&m[206])|(m[200]&m[203]&m[204]&m[205]&m[206]));
    m[212] = (((m[210]&~m[213]&~m[214]&~m[215]&~m[216])|(~m[210]&~m[213]&~m[214]&m[215]&~m[216])|(m[210]&m[213]&~m[214]&m[215]&~m[216])|(m[210]&~m[213]&m[214]&m[215]&~m[216])|(~m[210]&m[213]&~m[214]&~m[215]&m[216])|(~m[210]&~m[213]&m[214]&~m[215]&m[216])|(m[210]&m[213]&m[214]&~m[215]&m[216])|(~m[210]&m[213]&m[214]&m[215]&m[216]))&UnbiasedRNG[14])|((m[210]&~m[213]&~m[214]&m[215]&~m[216])|(~m[210]&~m[213]&~m[214]&~m[215]&m[216])|(m[210]&~m[213]&~m[214]&~m[215]&m[216])|(m[210]&m[213]&~m[214]&~m[215]&m[216])|(m[210]&~m[213]&m[214]&~m[215]&m[216])|(~m[210]&~m[213]&~m[214]&m[215]&m[216])|(m[210]&~m[213]&~m[214]&m[215]&m[216])|(~m[210]&m[213]&~m[214]&m[215]&m[216])|(m[210]&m[213]&~m[214]&m[215]&m[216])|(~m[210]&~m[213]&m[214]&m[215]&m[216])|(m[210]&~m[213]&m[214]&m[215]&m[216])|(m[210]&m[213]&m[214]&m[215]&m[216]));
    m[217] = (((m[215]&~m[218]&~m[219]&~m[220]&~m[221])|(~m[215]&~m[218]&~m[219]&m[220]&~m[221])|(m[215]&m[218]&~m[219]&m[220]&~m[221])|(m[215]&~m[218]&m[219]&m[220]&~m[221])|(~m[215]&m[218]&~m[219]&~m[220]&m[221])|(~m[215]&~m[218]&m[219]&~m[220]&m[221])|(m[215]&m[218]&m[219]&~m[220]&m[221])|(~m[215]&m[218]&m[219]&m[220]&m[221]))&UnbiasedRNG[15])|((m[215]&~m[218]&~m[219]&m[220]&~m[221])|(~m[215]&~m[218]&~m[219]&~m[220]&m[221])|(m[215]&~m[218]&~m[219]&~m[220]&m[221])|(m[215]&m[218]&~m[219]&~m[220]&m[221])|(m[215]&~m[218]&m[219]&~m[220]&m[221])|(~m[215]&~m[218]&~m[219]&m[220]&m[221])|(m[215]&~m[218]&~m[219]&m[220]&m[221])|(~m[215]&m[218]&~m[219]&m[220]&m[221])|(m[215]&m[218]&~m[219]&m[220]&m[221])|(~m[215]&~m[218]&m[219]&m[220]&m[221])|(m[215]&~m[218]&m[219]&m[220]&m[221])|(m[215]&m[218]&m[219]&m[220]&m[221]));
    m[222] = (((m[220]&~m[223]&~m[224]&~m[225]&~m[226])|(~m[220]&~m[223]&~m[224]&m[225]&~m[226])|(m[220]&m[223]&~m[224]&m[225]&~m[226])|(m[220]&~m[223]&m[224]&m[225]&~m[226])|(~m[220]&m[223]&~m[224]&~m[225]&m[226])|(~m[220]&~m[223]&m[224]&~m[225]&m[226])|(m[220]&m[223]&m[224]&~m[225]&m[226])|(~m[220]&m[223]&m[224]&m[225]&m[226]))&UnbiasedRNG[16])|((m[220]&~m[223]&~m[224]&m[225]&~m[226])|(~m[220]&~m[223]&~m[224]&~m[225]&m[226])|(m[220]&~m[223]&~m[224]&~m[225]&m[226])|(m[220]&m[223]&~m[224]&~m[225]&m[226])|(m[220]&~m[223]&m[224]&~m[225]&m[226])|(~m[220]&~m[223]&~m[224]&m[225]&m[226])|(m[220]&~m[223]&~m[224]&m[225]&m[226])|(~m[220]&m[223]&~m[224]&m[225]&m[226])|(m[220]&m[223]&~m[224]&m[225]&m[226])|(~m[220]&~m[223]&m[224]&m[225]&m[226])|(m[220]&~m[223]&m[224]&m[225]&m[226])|(m[220]&m[223]&m[224]&m[225]&m[226]));
    m[227] = (((m[225]&~m[228]&~m[229]&~m[230]&~m[231])|(~m[225]&~m[228]&~m[229]&m[230]&~m[231])|(m[225]&m[228]&~m[229]&m[230]&~m[231])|(m[225]&~m[228]&m[229]&m[230]&~m[231])|(~m[225]&m[228]&~m[229]&~m[230]&m[231])|(~m[225]&~m[228]&m[229]&~m[230]&m[231])|(m[225]&m[228]&m[229]&~m[230]&m[231])|(~m[225]&m[228]&m[229]&m[230]&m[231]))&UnbiasedRNG[17])|((m[225]&~m[228]&~m[229]&m[230]&~m[231])|(~m[225]&~m[228]&~m[229]&~m[230]&m[231])|(m[225]&~m[228]&~m[229]&~m[230]&m[231])|(m[225]&m[228]&~m[229]&~m[230]&m[231])|(m[225]&~m[228]&m[229]&~m[230]&m[231])|(~m[225]&~m[228]&~m[229]&m[230]&m[231])|(m[225]&~m[228]&~m[229]&m[230]&m[231])|(~m[225]&m[228]&~m[229]&m[230]&m[231])|(m[225]&m[228]&~m[229]&m[230]&m[231])|(~m[225]&~m[228]&m[229]&m[230]&m[231])|(m[225]&~m[228]&m[229]&m[230]&m[231])|(m[225]&m[228]&m[229]&m[230]&m[231]));
    m[232] = (((m[211]&~m[233]&~m[234]&~m[235]&~m[236])|(~m[211]&~m[233]&~m[234]&m[235]&~m[236])|(m[211]&m[233]&~m[234]&m[235]&~m[236])|(m[211]&~m[233]&m[234]&m[235]&~m[236])|(~m[211]&m[233]&~m[234]&~m[235]&m[236])|(~m[211]&~m[233]&m[234]&~m[235]&m[236])|(m[211]&m[233]&m[234]&~m[235]&m[236])|(~m[211]&m[233]&m[234]&m[235]&m[236]))&UnbiasedRNG[18])|((m[211]&~m[233]&~m[234]&m[235]&~m[236])|(~m[211]&~m[233]&~m[234]&~m[235]&m[236])|(m[211]&~m[233]&~m[234]&~m[235]&m[236])|(m[211]&m[233]&~m[234]&~m[235]&m[236])|(m[211]&~m[233]&m[234]&~m[235]&m[236])|(~m[211]&~m[233]&~m[234]&m[235]&m[236])|(m[211]&~m[233]&~m[234]&m[235]&m[236])|(~m[211]&m[233]&~m[234]&m[235]&m[236])|(m[211]&m[233]&~m[234]&m[235]&m[236])|(~m[211]&~m[233]&m[234]&m[235]&m[236])|(m[211]&~m[233]&m[234]&m[235]&m[236])|(m[211]&m[233]&m[234]&m[235]&m[236]));
    m[237] = (((m[235]&~m[238]&~m[239]&~m[240]&~m[241])|(~m[235]&~m[238]&~m[239]&m[240]&~m[241])|(m[235]&m[238]&~m[239]&m[240]&~m[241])|(m[235]&~m[238]&m[239]&m[240]&~m[241])|(~m[235]&m[238]&~m[239]&~m[240]&m[241])|(~m[235]&~m[238]&m[239]&~m[240]&m[241])|(m[235]&m[238]&m[239]&~m[240]&m[241])|(~m[235]&m[238]&m[239]&m[240]&m[241]))&UnbiasedRNG[19])|((m[235]&~m[238]&~m[239]&m[240]&~m[241])|(~m[235]&~m[238]&~m[239]&~m[240]&m[241])|(m[235]&~m[238]&~m[239]&~m[240]&m[241])|(m[235]&m[238]&~m[239]&~m[240]&m[241])|(m[235]&~m[238]&m[239]&~m[240]&m[241])|(~m[235]&~m[238]&~m[239]&m[240]&m[241])|(m[235]&~m[238]&~m[239]&m[240]&m[241])|(~m[235]&m[238]&~m[239]&m[240]&m[241])|(m[235]&m[238]&~m[239]&m[240]&m[241])|(~m[235]&~m[238]&m[239]&m[240]&m[241])|(m[235]&~m[238]&m[239]&m[240]&m[241])|(m[235]&m[238]&m[239]&m[240]&m[241]));
    m[242] = (((m[240]&~m[243]&~m[244]&~m[245]&~m[246])|(~m[240]&~m[243]&~m[244]&m[245]&~m[246])|(m[240]&m[243]&~m[244]&m[245]&~m[246])|(m[240]&~m[243]&m[244]&m[245]&~m[246])|(~m[240]&m[243]&~m[244]&~m[245]&m[246])|(~m[240]&~m[243]&m[244]&~m[245]&m[246])|(m[240]&m[243]&m[244]&~m[245]&m[246])|(~m[240]&m[243]&m[244]&m[245]&m[246]))&UnbiasedRNG[20])|((m[240]&~m[243]&~m[244]&m[245]&~m[246])|(~m[240]&~m[243]&~m[244]&~m[245]&m[246])|(m[240]&~m[243]&~m[244]&~m[245]&m[246])|(m[240]&m[243]&~m[244]&~m[245]&m[246])|(m[240]&~m[243]&m[244]&~m[245]&m[246])|(~m[240]&~m[243]&~m[244]&m[245]&m[246])|(m[240]&~m[243]&~m[244]&m[245]&m[246])|(~m[240]&m[243]&~m[244]&m[245]&m[246])|(m[240]&m[243]&~m[244]&m[245]&m[246])|(~m[240]&~m[243]&m[244]&m[245]&m[246])|(m[240]&~m[243]&m[244]&m[245]&m[246])|(m[240]&m[243]&m[244]&m[245]&m[246]));
    m[247] = (((m[245]&~m[248]&~m[249]&~m[250]&~m[251])|(~m[245]&~m[248]&~m[249]&m[250]&~m[251])|(m[245]&m[248]&~m[249]&m[250]&~m[251])|(m[245]&~m[248]&m[249]&m[250]&~m[251])|(~m[245]&m[248]&~m[249]&~m[250]&m[251])|(~m[245]&~m[248]&m[249]&~m[250]&m[251])|(m[245]&m[248]&m[249]&~m[250]&m[251])|(~m[245]&m[248]&m[249]&m[250]&m[251]))&UnbiasedRNG[21])|((m[245]&~m[248]&~m[249]&m[250]&~m[251])|(~m[245]&~m[248]&~m[249]&~m[250]&m[251])|(m[245]&~m[248]&~m[249]&~m[250]&m[251])|(m[245]&m[248]&~m[249]&~m[250]&m[251])|(m[245]&~m[248]&m[249]&~m[250]&m[251])|(~m[245]&~m[248]&~m[249]&m[250]&m[251])|(m[245]&~m[248]&~m[249]&m[250]&m[251])|(~m[245]&m[248]&~m[249]&m[250]&m[251])|(m[245]&m[248]&~m[249]&m[250]&m[251])|(~m[245]&~m[248]&m[249]&m[250]&m[251])|(m[245]&~m[248]&m[249]&m[250]&m[251])|(m[245]&m[248]&m[249]&m[250]&m[251]));
    m[252] = (((m[236]&~m[253]&~m[254]&~m[255]&~m[256])|(~m[236]&~m[253]&~m[254]&m[255]&~m[256])|(m[236]&m[253]&~m[254]&m[255]&~m[256])|(m[236]&~m[253]&m[254]&m[255]&~m[256])|(~m[236]&m[253]&~m[254]&~m[255]&m[256])|(~m[236]&~m[253]&m[254]&~m[255]&m[256])|(m[236]&m[253]&m[254]&~m[255]&m[256])|(~m[236]&m[253]&m[254]&m[255]&m[256]))&UnbiasedRNG[22])|((m[236]&~m[253]&~m[254]&m[255]&~m[256])|(~m[236]&~m[253]&~m[254]&~m[255]&m[256])|(m[236]&~m[253]&~m[254]&~m[255]&m[256])|(m[236]&m[253]&~m[254]&~m[255]&m[256])|(m[236]&~m[253]&m[254]&~m[255]&m[256])|(~m[236]&~m[253]&~m[254]&m[255]&m[256])|(m[236]&~m[253]&~m[254]&m[255]&m[256])|(~m[236]&m[253]&~m[254]&m[255]&m[256])|(m[236]&m[253]&~m[254]&m[255]&m[256])|(~m[236]&~m[253]&m[254]&m[255]&m[256])|(m[236]&~m[253]&m[254]&m[255]&m[256])|(m[236]&m[253]&m[254]&m[255]&m[256]));
    m[257] = (((m[255]&~m[258]&~m[259]&~m[260]&~m[261])|(~m[255]&~m[258]&~m[259]&m[260]&~m[261])|(m[255]&m[258]&~m[259]&m[260]&~m[261])|(m[255]&~m[258]&m[259]&m[260]&~m[261])|(~m[255]&m[258]&~m[259]&~m[260]&m[261])|(~m[255]&~m[258]&m[259]&~m[260]&m[261])|(m[255]&m[258]&m[259]&~m[260]&m[261])|(~m[255]&m[258]&m[259]&m[260]&m[261]))&UnbiasedRNG[23])|((m[255]&~m[258]&~m[259]&m[260]&~m[261])|(~m[255]&~m[258]&~m[259]&~m[260]&m[261])|(m[255]&~m[258]&~m[259]&~m[260]&m[261])|(m[255]&m[258]&~m[259]&~m[260]&m[261])|(m[255]&~m[258]&m[259]&~m[260]&m[261])|(~m[255]&~m[258]&~m[259]&m[260]&m[261])|(m[255]&~m[258]&~m[259]&m[260]&m[261])|(~m[255]&m[258]&~m[259]&m[260]&m[261])|(m[255]&m[258]&~m[259]&m[260]&m[261])|(~m[255]&~m[258]&m[259]&m[260]&m[261])|(m[255]&~m[258]&m[259]&m[260]&m[261])|(m[255]&m[258]&m[259]&m[260]&m[261]));
    m[262] = (((m[260]&~m[263]&~m[264]&~m[265]&~m[266])|(~m[260]&~m[263]&~m[264]&m[265]&~m[266])|(m[260]&m[263]&~m[264]&m[265]&~m[266])|(m[260]&~m[263]&m[264]&m[265]&~m[266])|(~m[260]&m[263]&~m[264]&~m[265]&m[266])|(~m[260]&~m[263]&m[264]&~m[265]&m[266])|(m[260]&m[263]&m[264]&~m[265]&m[266])|(~m[260]&m[263]&m[264]&m[265]&m[266]))&UnbiasedRNG[24])|((m[260]&~m[263]&~m[264]&m[265]&~m[266])|(~m[260]&~m[263]&~m[264]&~m[265]&m[266])|(m[260]&~m[263]&~m[264]&~m[265]&m[266])|(m[260]&m[263]&~m[264]&~m[265]&m[266])|(m[260]&~m[263]&m[264]&~m[265]&m[266])|(~m[260]&~m[263]&~m[264]&m[265]&m[266])|(m[260]&~m[263]&~m[264]&m[265]&m[266])|(~m[260]&m[263]&~m[264]&m[265]&m[266])|(m[260]&m[263]&~m[264]&m[265]&m[266])|(~m[260]&~m[263]&m[264]&m[265]&m[266])|(m[260]&~m[263]&m[264]&m[265]&m[266])|(m[260]&m[263]&m[264]&m[265]&m[266]));
    m[267] = (((m[256]&~m[268]&~m[269]&~m[270]&~m[271])|(~m[256]&~m[268]&~m[269]&m[270]&~m[271])|(m[256]&m[268]&~m[269]&m[270]&~m[271])|(m[256]&~m[268]&m[269]&m[270]&~m[271])|(~m[256]&m[268]&~m[269]&~m[270]&m[271])|(~m[256]&~m[268]&m[269]&~m[270]&m[271])|(m[256]&m[268]&m[269]&~m[270]&m[271])|(~m[256]&m[268]&m[269]&m[270]&m[271]))&UnbiasedRNG[25])|((m[256]&~m[268]&~m[269]&m[270]&~m[271])|(~m[256]&~m[268]&~m[269]&~m[270]&m[271])|(m[256]&~m[268]&~m[269]&~m[270]&m[271])|(m[256]&m[268]&~m[269]&~m[270]&m[271])|(m[256]&~m[268]&m[269]&~m[270]&m[271])|(~m[256]&~m[268]&~m[269]&m[270]&m[271])|(m[256]&~m[268]&~m[269]&m[270]&m[271])|(~m[256]&m[268]&~m[269]&m[270]&m[271])|(m[256]&m[268]&~m[269]&m[270]&m[271])|(~m[256]&~m[268]&m[269]&m[270]&m[271])|(m[256]&~m[268]&m[269]&m[270]&m[271])|(m[256]&m[268]&m[269]&m[270]&m[271]));
    m[272] = (((m[270]&~m[273]&~m[274]&~m[275]&~m[276])|(~m[270]&~m[273]&~m[274]&m[275]&~m[276])|(m[270]&m[273]&~m[274]&m[275]&~m[276])|(m[270]&~m[273]&m[274]&m[275]&~m[276])|(~m[270]&m[273]&~m[274]&~m[275]&m[276])|(~m[270]&~m[273]&m[274]&~m[275]&m[276])|(m[270]&m[273]&m[274]&~m[275]&m[276])|(~m[270]&m[273]&m[274]&m[275]&m[276]))&UnbiasedRNG[26])|((m[270]&~m[273]&~m[274]&m[275]&~m[276])|(~m[270]&~m[273]&~m[274]&~m[275]&m[276])|(m[270]&~m[273]&~m[274]&~m[275]&m[276])|(m[270]&m[273]&~m[274]&~m[275]&m[276])|(m[270]&~m[273]&m[274]&~m[275]&m[276])|(~m[270]&~m[273]&~m[274]&m[275]&m[276])|(m[270]&~m[273]&~m[274]&m[275]&m[276])|(~m[270]&m[273]&~m[274]&m[275]&m[276])|(m[270]&m[273]&~m[274]&m[275]&m[276])|(~m[270]&~m[273]&m[274]&m[275]&m[276])|(m[270]&~m[273]&m[274]&m[275]&m[276])|(m[270]&m[273]&m[274]&m[275]&m[276]));
    m[277] = (((m[271]&~m[278]&~m[279]&~m[280]&~m[281])|(~m[271]&~m[278]&~m[279]&m[280]&~m[281])|(m[271]&m[278]&~m[279]&m[280]&~m[281])|(m[271]&~m[278]&m[279]&m[280]&~m[281])|(~m[271]&m[278]&~m[279]&~m[280]&m[281])|(~m[271]&~m[278]&m[279]&~m[280]&m[281])|(m[271]&m[278]&m[279]&~m[280]&m[281])|(~m[271]&m[278]&m[279]&m[280]&m[281]))&UnbiasedRNG[27])|((m[271]&~m[278]&~m[279]&m[280]&~m[281])|(~m[271]&~m[278]&~m[279]&~m[280]&m[281])|(m[271]&~m[278]&~m[279]&~m[280]&m[281])|(m[271]&m[278]&~m[279]&~m[280]&m[281])|(m[271]&~m[278]&m[279]&~m[280]&m[281])|(~m[271]&~m[278]&~m[279]&m[280]&m[281])|(m[271]&~m[278]&~m[279]&m[280]&m[281])|(~m[271]&m[278]&~m[279]&m[280]&m[281])|(m[271]&m[278]&~m[279]&m[280]&m[281])|(~m[271]&~m[278]&m[279]&m[280]&m[281])|(m[271]&~m[278]&m[279]&m[280]&m[281])|(m[271]&m[278]&m[279]&m[280]&m[281]));
end

always @(posedge color1_clk) begin
    m[12] = (((m[0]&m[26]&~m[27]&~m[28]&~m[29])|(m[0]&~m[26]&m[27]&~m[28]&~m[29])|(~m[0]&m[26]&m[27]&~m[28]&~m[29])|(m[0]&~m[26]&~m[27]&m[28]&~m[29])|(~m[0]&m[26]&~m[27]&m[28]&~m[29])|(~m[0]&~m[26]&m[27]&m[28]&~m[29])|(m[0]&~m[26]&~m[27]&~m[28]&m[29])|(~m[0]&m[26]&~m[27]&~m[28]&m[29])|(~m[0]&~m[26]&m[27]&~m[28]&m[29])|(~m[0]&~m[26]&~m[27]&m[28]&m[29]))&BiasedRNG[47])|(((m[0]&m[26]&m[27]&~m[28]&~m[29])|(m[0]&m[26]&~m[27]&m[28]&~m[29])|(m[0]&~m[26]&m[27]&m[28]&~m[29])|(~m[0]&m[26]&m[27]&m[28]&~m[29])|(m[0]&m[26]&~m[27]&~m[28]&m[29])|(m[0]&~m[26]&m[27]&~m[28]&m[29])|(~m[0]&m[26]&m[27]&~m[28]&m[29])|(m[0]&~m[26]&~m[27]&m[28]&m[29])|(~m[0]&m[26]&~m[27]&m[28]&m[29])|(~m[0]&~m[26]&m[27]&m[28]&m[29]))&~BiasedRNG[47])|((m[0]&m[26]&m[27]&m[28]&~m[29])|(m[0]&m[26]&m[27]&~m[28]&m[29])|(m[0]&m[26]&~m[27]&m[28]&m[29])|(m[0]&~m[26]&m[27]&m[28]&m[29])|(~m[0]&m[26]&m[27]&m[28]&m[29])|(m[0]&m[26]&m[27]&m[28]&m[29]));
    m[13] = (((m[1]&m[32]&~m[33]&~m[34]&~m[35])|(m[1]&~m[32]&m[33]&~m[34]&~m[35])|(~m[1]&m[32]&m[33]&~m[34]&~m[35])|(m[1]&~m[32]&~m[33]&m[34]&~m[35])|(~m[1]&m[32]&~m[33]&m[34]&~m[35])|(~m[1]&~m[32]&m[33]&m[34]&~m[35])|(m[1]&~m[32]&~m[33]&~m[34]&m[35])|(~m[1]&m[32]&~m[33]&~m[34]&m[35])|(~m[1]&~m[32]&m[33]&~m[34]&m[35])|(~m[1]&~m[32]&~m[33]&m[34]&m[35]))&BiasedRNG[48])|(((m[1]&m[32]&m[33]&~m[34]&~m[35])|(m[1]&m[32]&~m[33]&m[34]&~m[35])|(m[1]&~m[32]&m[33]&m[34]&~m[35])|(~m[1]&m[32]&m[33]&m[34]&~m[35])|(m[1]&m[32]&~m[33]&~m[34]&m[35])|(m[1]&~m[32]&m[33]&~m[34]&m[35])|(~m[1]&m[32]&m[33]&~m[34]&m[35])|(m[1]&~m[32]&~m[33]&m[34]&m[35])|(~m[1]&m[32]&~m[33]&m[34]&m[35])|(~m[1]&~m[32]&m[33]&m[34]&m[35]))&~BiasedRNG[48])|((m[1]&m[32]&m[33]&m[34]&~m[35])|(m[1]&m[32]&m[33]&~m[34]&m[35])|(m[1]&m[32]&~m[33]&m[34]&m[35])|(m[1]&~m[32]&m[33]&m[34]&m[35])|(~m[1]&m[32]&m[33]&m[34]&m[35])|(m[1]&m[32]&m[33]&m[34]&m[35]));
    m[14] = (((m[2]&m[38]&~m[39]&~m[40]&~m[41])|(m[2]&~m[38]&m[39]&~m[40]&~m[41])|(~m[2]&m[38]&m[39]&~m[40]&~m[41])|(m[2]&~m[38]&~m[39]&m[40]&~m[41])|(~m[2]&m[38]&~m[39]&m[40]&~m[41])|(~m[2]&~m[38]&m[39]&m[40]&~m[41])|(m[2]&~m[38]&~m[39]&~m[40]&m[41])|(~m[2]&m[38]&~m[39]&~m[40]&m[41])|(~m[2]&~m[38]&m[39]&~m[40]&m[41])|(~m[2]&~m[38]&~m[39]&m[40]&m[41]))&BiasedRNG[49])|(((m[2]&m[38]&m[39]&~m[40]&~m[41])|(m[2]&m[38]&~m[39]&m[40]&~m[41])|(m[2]&~m[38]&m[39]&m[40]&~m[41])|(~m[2]&m[38]&m[39]&m[40]&~m[41])|(m[2]&m[38]&~m[39]&~m[40]&m[41])|(m[2]&~m[38]&m[39]&~m[40]&m[41])|(~m[2]&m[38]&m[39]&~m[40]&m[41])|(m[2]&~m[38]&~m[39]&m[40]&m[41])|(~m[2]&m[38]&~m[39]&m[40]&m[41])|(~m[2]&~m[38]&m[39]&m[40]&m[41]))&~BiasedRNG[49])|((m[2]&m[38]&m[39]&m[40]&~m[41])|(m[2]&m[38]&m[39]&~m[40]&m[41])|(m[2]&m[38]&~m[39]&m[40]&m[41])|(m[2]&~m[38]&m[39]&m[40]&m[41])|(~m[2]&m[38]&m[39]&m[40]&m[41])|(m[2]&m[38]&m[39]&m[40]&m[41]));
    m[15] = (((m[3]&m[44]&~m[45]&~m[46]&~m[47])|(m[3]&~m[44]&m[45]&~m[46]&~m[47])|(~m[3]&m[44]&m[45]&~m[46]&~m[47])|(m[3]&~m[44]&~m[45]&m[46]&~m[47])|(~m[3]&m[44]&~m[45]&m[46]&~m[47])|(~m[3]&~m[44]&m[45]&m[46]&~m[47])|(m[3]&~m[44]&~m[45]&~m[46]&m[47])|(~m[3]&m[44]&~m[45]&~m[46]&m[47])|(~m[3]&~m[44]&m[45]&~m[46]&m[47])|(~m[3]&~m[44]&~m[45]&m[46]&m[47]))&BiasedRNG[50])|(((m[3]&m[44]&m[45]&~m[46]&~m[47])|(m[3]&m[44]&~m[45]&m[46]&~m[47])|(m[3]&~m[44]&m[45]&m[46]&~m[47])|(~m[3]&m[44]&m[45]&m[46]&~m[47])|(m[3]&m[44]&~m[45]&~m[46]&m[47])|(m[3]&~m[44]&m[45]&~m[46]&m[47])|(~m[3]&m[44]&m[45]&~m[46]&m[47])|(m[3]&~m[44]&~m[45]&m[46]&m[47])|(~m[3]&m[44]&~m[45]&m[46]&m[47])|(~m[3]&~m[44]&m[45]&m[46]&m[47]))&~BiasedRNG[50])|((m[3]&m[44]&m[45]&m[46]&~m[47])|(m[3]&m[44]&m[45]&~m[46]&m[47])|(m[3]&m[44]&~m[45]&m[46]&m[47])|(m[3]&~m[44]&m[45]&m[46]&m[47])|(~m[3]&m[44]&m[45]&m[46]&m[47])|(m[3]&m[44]&m[45]&m[46]&m[47]));
    m[16] = (((m[4]&m[50]&~m[51]&~m[52]&~m[53])|(m[4]&~m[50]&m[51]&~m[52]&~m[53])|(~m[4]&m[50]&m[51]&~m[52]&~m[53])|(m[4]&~m[50]&~m[51]&m[52]&~m[53])|(~m[4]&m[50]&~m[51]&m[52]&~m[53])|(~m[4]&~m[50]&m[51]&m[52]&~m[53])|(m[4]&~m[50]&~m[51]&~m[52]&m[53])|(~m[4]&m[50]&~m[51]&~m[52]&m[53])|(~m[4]&~m[50]&m[51]&~m[52]&m[53])|(~m[4]&~m[50]&~m[51]&m[52]&m[53]))&BiasedRNG[51])|(((m[4]&m[50]&m[51]&~m[52]&~m[53])|(m[4]&m[50]&~m[51]&m[52]&~m[53])|(m[4]&~m[50]&m[51]&m[52]&~m[53])|(~m[4]&m[50]&m[51]&m[52]&~m[53])|(m[4]&m[50]&~m[51]&~m[52]&m[53])|(m[4]&~m[50]&m[51]&~m[52]&m[53])|(~m[4]&m[50]&m[51]&~m[52]&m[53])|(m[4]&~m[50]&~m[51]&m[52]&m[53])|(~m[4]&m[50]&~m[51]&m[52]&m[53])|(~m[4]&~m[50]&m[51]&m[52]&m[53]))&~BiasedRNG[51])|((m[4]&m[50]&m[51]&m[52]&~m[53])|(m[4]&m[50]&m[51]&~m[52]&m[53])|(m[4]&m[50]&~m[51]&m[52]&m[53])|(m[4]&~m[50]&m[51]&m[52]&m[53])|(~m[4]&m[50]&m[51]&m[52]&m[53])|(m[4]&m[50]&m[51]&m[52]&m[53]));
    m[17] = (((m[5]&m[56]&~m[57]&~m[58]&~m[59])|(m[5]&~m[56]&m[57]&~m[58]&~m[59])|(~m[5]&m[56]&m[57]&~m[58]&~m[59])|(m[5]&~m[56]&~m[57]&m[58]&~m[59])|(~m[5]&m[56]&~m[57]&m[58]&~m[59])|(~m[5]&~m[56]&m[57]&m[58]&~m[59])|(m[5]&~m[56]&~m[57]&~m[58]&m[59])|(~m[5]&m[56]&~m[57]&~m[58]&m[59])|(~m[5]&~m[56]&m[57]&~m[58]&m[59])|(~m[5]&~m[56]&~m[57]&m[58]&m[59]))&BiasedRNG[52])|(((m[5]&m[56]&m[57]&~m[58]&~m[59])|(m[5]&m[56]&~m[57]&m[58]&~m[59])|(m[5]&~m[56]&m[57]&m[58]&~m[59])|(~m[5]&m[56]&m[57]&m[58]&~m[59])|(m[5]&m[56]&~m[57]&~m[58]&m[59])|(m[5]&~m[56]&m[57]&~m[58]&m[59])|(~m[5]&m[56]&m[57]&~m[58]&m[59])|(m[5]&~m[56]&~m[57]&m[58]&m[59])|(~m[5]&m[56]&~m[57]&m[58]&m[59])|(~m[5]&~m[56]&m[57]&m[58]&m[59]))&~BiasedRNG[52])|((m[5]&m[56]&m[57]&m[58]&~m[59])|(m[5]&m[56]&m[57]&~m[58]&m[59])|(m[5]&m[56]&~m[57]&m[58]&m[59])|(m[5]&~m[56]&m[57]&m[58]&m[59])|(~m[5]&m[56]&m[57]&m[58]&m[59])|(m[5]&m[56]&m[57]&m[58]&m[59]));
    m[18] = (((m[6]&m[62]&~m[63]&~m[64]&~m[65])|(m[6]&~m[62]&m[63]&~m[64]&~m[65])|(~m[6]&m[62]&m[63]&~m[64]&~m[65])|(m[6]&~m[62]&~m[63]&m[64]&~m[65])|(~m[6]&m[62]&~m[63]&m[64]&~m[65])|(~m[6]&~m[62]&m[63]&m[64]&~m[65])|(m[6]&~m[62]&~m[63]&~m[64]&m[65])|(~m[6]&m[62]&~m[63]&~m[64]&m[65])|(~m[6]&~m[62]&m[63]&~m[64]&m[65])|(~m[6]&~m[62]&~m[63]&m[64]&m[65]))&BiasedRNG[53])|(((m[6]&m[62]&m[63]&~m[64]&~m[65])|(m[6]&m[62]&~m[63]&m[64]&~m[65])|(m[6]&~m[62]&m[63]&m[64]&~m[65])|(~m[6]&m[62]&m[63]&m[64]&~m[65])|(m[6]&m[62]&~m[63]&~m[64]&m[65])|(m[6]&~m[62]&m[63]&~m[64]&m[65])|(~m[6]&m[62]&m[63]&~m[64]&m[65])|(m[6]&~m[62]&~m[63]&m[64]&m[65])|(~m[6]&m[62]&~m[63]&m[64]&m[65])|(~m[6]&~m[62]&m[63]&m[64]&m[65]))&~BiasedRNG[53])|((m[6]&m[62]&m[63]&m[64]&~m[65])|(m[6]&m[62]&m[63]&~m[64]&m[65])|(m[6]&m[62]&~m[63]&m[64]&m[65])|(m[6]&~m[62]&m[63]&m[64]&m[65])|(~m[6]&m[62]&m[63]&m[64]&m[65])|(m[6]&m[62]&m[63]&m[64]&m[65]));
    m[19] = (((m[7]&m[68]&~m[69]&~m[70]&~m[71])|(m[7]&~m[68]&m[69]&~m[70]&~m[71])|(~m[7]&m[68]&m[69]&~m[70]&~m[71])|(m[7]&~m[68]&~m[69]&m[70]&~m[71])|(~m[7]&m[68]&~m[69]&m[70]&~m[71])|(~m[7]&~m[68]&m[69]&m[70]&~m[71])|(m[7]&~m[68]&~m[69]&~m[70]&m[71])|(~m[7]&m[68]&~m[69]&~m[70]&m[71])|(~m[7]&~m[68]&m[69]&~m[70]&m[71])|(~m[7]&~m[68]&~m[69]&m[70]&m[71]))&BiasedRNG[54])|(((m[7]&m[68]&m[69]&~m[70]&~m[71])|(m[7]&m[68]&~m[69]&m[70]&~m[71])|(m[7]&~m[68]&m[69]&m[70]&~m[71])|(~m[7]&m[68]&m[69]&m[70]&~m[71])|(m[7]&m[68]&~m[69]&~m[70]&m[71])|(m[7]&~m[68]&m[69]&~m[70]&m[71])|(~m[7]&m[68]&m[69]&~m[70]&m[71])|(m[7]&~m[68]&~m[69]&m[70]&m[71])|(~m[7]&m[68]&~m[69]&m[70]&m[71])|(~m[7]&~m[68]&m[69]&m[70]&m[71]))&~BiasedRNG[54])|((m[7]&m[68]&m[69]&m[70]&~m[71])|(m[7]&m[68]&m[69]&~m[70]&m[71])|(m[7]&m[68]&~m[69]&m[70]&m[71])|(m[7]&~m[68]&m[69]&m[70]&m[71])|(~m[7]&m[68]&m[69]&m[70]&m[71])|(m[7]&m[68]&m[69]&m[70]&m[71]));
    m[20] = (((m[8]&m[74]&~m[75]&~m[76]&~m[77])|(m[8]&~m[74]&m[75]&~m[76]&~m[77])|(~m[8]&m[74]&m[75]&~m[76]&~m[77])|(m[8]&~m[74]&~m[75]&m[76]&~m[77])|(~m[8]&m[74]&~m[75]&m[76]&~m[77])|(~m[8]&~m[74]&m[75]&m[76]&~m[77])|(m[8]&~m[74]&~m[75]&~m[76]&m[77])|(~m[8]&m[74]&~m[75]&~m[76]&m[77])|(~m[8]&~m[74]&m[75]&~m[76]&m[77])|(~m[8]&~m[74]&~m[75]&m[76]&m[77]))&BiasedRNG[55])|(((m[8]&m[74]&m[75]&~m[76]&~m[77])|(m[8]&m[74]&~m[75]&m[76]&~m[77])|(m[8]&~m[74]&m[75]&m[76]&~m[77])|(~m[8]&m[74]&m[75]&m[76]&~m[77])|(m[8]&m[74]&~m[75]&~m[76]&m[77])|(m[8]&~m[74]&m[75]&~m[76]&m[77])|(~m[8]&m[74]&m[75]&~m[76]&m[77])|(m[8]&~m[74]&~m[75]&m[76]&m[77])|(~m[8]&m[74]&~m[75]&m[76]&m[77])|(~m[8]&~m[74]&m[75]&m[76]&m[77]))&~BiasedRNG[55])|((m[8]&m[74]&m[75]&m[76]&~m[77])|(m[8]&m[74]&m[75]&~m[76]&m[77])|(m[8]&m[74]&~m[75]&m[76]&m[77])|(m[8]&~m[74]&m[75]&m[76]&m[77])|(~m[8]&m[74]&m[75]&m[76]&m[77])|(m[8]&m[74]&m[75]&m[76]&m[77]));
    m[21] = (((m[9]&m[80]&~m[81]&~m[82]&~m[83])|(m[9]&~m[80]&m[81]&~m[82]&~m[83])|(~m[9]&m[80]&m[81]&~m[82]&~m[83])|(m[9]&~m[80]&~m[81]&m[82]&~m[83])|(~m[9]&m[80]&~m[81]&m[82]&~m[83])|(~m[9]&~m[80]&m[81]&m[82]&~m[83])|(m[9]&~m[80]&~m[81]&~m[82]&m[83])|(~m[9]&m[80]&~m[81]&~m[82]&m[83])|(~m[9]&~m[80]&m[81]&~m[82]&m[83])|(~m[9]&~m[80]&~m[81]&m[82]&m[83]))&BiasedRNG[56])|(((m[9]&m[80]&m[81]&~m[82]&~m[83])|(m[9]&m[80]&~m[81]&m[82]&~m[83])|(m[9]&~m[80]&m[81]&m[82]&~m[83])|(~m[9]&m[80]&m[81]&m[82]&~m[83])|(m[9]&m[80]&~m[81]&~m[82]&m[83])|(m[9]&~m[80]&m[81]&~m[82]&m[83])|(~m[9]&m[80]&m[81]&~m[82]&m[83])|(m[9]&~m[80]&~m[81]&m[82]&m[83])|(~m[9]&m[80]&~m[81]&m[82]&m[83])|(~m[9]&~m[80]&m[81]&m[82]&m[83]))&~BiasedRNG[56])|((m[9]&m[80]&m[81]&m[82]&~m[83])|(m[9]&m[80]&m[81]&~m[82]&m[83])|(m[9]&m[80]&~m[81]&m[82]&m[83])|(m[9]&~m[80]&m[81]&m[82]&m[83])|(~m[9]&m[80]&m[81]&m[82]&m[83])|(m[9]&m[80]&m[81]&m[82]&m[83]));
    m[22] = (((m[10]&m[86]&~m[87]&~m[88]&~m[89])|(m[10]&~m[86]&m[87]&~m[88]&~m[89])|(~m[10]&m[86]&m[87]&~m[88]&~m[89])|(m[10]&~m[86]&~m[87]&m[88]&~m[89])|(~m[10]&m[86]&~m[87]&m[88]&~m[89])|(~m[10]&~m[86]&m[87]&m[88]&~m[89])|(m[10]&~m[86]&~m[87]&~m[88]&m[89])|(~m[10]&m[86]&~m[87]&~m[88]&m[89])|(~m[10]&~m[86]&m[87]&~m[88]&m[89])|(~m[10]&~m[86]&~m[87]&m[88]&m[89]))&BiasedRNG[57])|(((m[10]&m[86]&m[87]&~m[88]&~m[89])|(m[10]&m[86]&~m[87]&m[88]&~m[89])|(m[10]&~m[86]&m[87]&m[88]&~m[89])|(~m[10]&m[86]&m[87]&m[88]&~m[89])|(m[10]&m[86]&~m[87]&~m[88]&m[89])|(m[10]&~m[86]&m[87]&~m[88]&m[89])|(~m[10]&m[86]&m[87]&~m[88]&m[89])|(m[10]&~m[86]&~m[87]&m[88]&m[89])|(~m[10]&m[86]&~m[87]&m[88]&m[89])|(~m[10]&~m[86]&m[87]&m[88]&m[89]))&~BiasedRNG[57])|((m[10]&m[86]&m[87]&m[88]&~m[89])|(m[10]&m[86]&m[87]&~m[88]&m[89])|(m[10]&m[86]&~m[87]&m[88]&m[89])|(m[10]&~m[86]&m[87]&m[88]&m[89])|(~m[10]&m[86]&m[87]&m[88]&m[89])|(m[10]&m[86]&m[87]&m[88]&m[89]));
    m[23] = (((m[11]&m[92]&~m[93]&~m[94]&~m[95])|(m[11]&~m[92]&m[93]&~m[94]&~m[95])|(~m[11]&m[92]&m[93]&~m[94]&~m[95])|(m[11]&~m[92]&~m[93]&m[94]&~m[95])|(~m[11]&m[92]&~m[93]&m[94]&~m[95])|(~m[11]&~m[92]&m[93]&m[94]&~m[95])|(m[11]&~m[92]&~m[93]&~m[94]&m[95])|(~m[11]&m[92]&~m[93]&~m[94]&m[95])|(~m[11]&~m[92]&m[93]&~m[94]&m[95])|(~m[11]&~m[92]&~m[93]&m[94]&m[95]))&BiasedRNG[58])|(((m[11]&m[92]&m[93]&~m[94]&~m[95])|(m[11]&m[92]&~m[93]&m[94]&~m[95])|(m[11]&~m[92]&m[93]&m[94]&~m[95])|(~m[11]&m[92]&m[93]&m[94]&~m[95])|(m[11]&m[92]&~m[93]&~m[94]&m[95])|(m[11]&~m[92]&m[93]&~m[94]&m[95])|(~m[11]&m[92]&m[93]&~m[94]&m[95])|(m[11]&~m[92]&~m[93]&m[94]&m[95])|(~m[11]&m[92]&~m[93]&m[94]&m[95])|(~m[11]&~m[92]&m[93]&m[94]&m[95]))&~BiasedRNG[58])|((m[11]&m[92]&m[93]&m[94]&~m[95])|(m[11]&m[92]&m[93]&~m[94]&m[95])|(m[11]&m[92]&~m[93]&m[94]&m[95])|(m[11]&~m[92]&m[93]&m[94]&m[95])|(~m[11]&m[92]&m[93]&m[94]&m[95])|(m[11]&m[92]&m[93]&m[94]&m[95]));
    m[24] = (((~m[0]&~m[60]&~m[96])|(m[0]&m[60]&~m[96]))&BiasedRNG[59])|(((m[0]&~m[60]&~m[96])|(~m[0]&m[60]&m[96]))&~BiasedRNG[59])|((~m[0]&~m[60]&m[96])|(m[0]&~m[60]&m[96])|(m[0]&m[60]&m[96]));
    m[25] = (((~m[0]&~m[66]&~m[102])|(m[0]&m[66]&~m[102]))&BiasedRNG[60])|(((m[0]&~m[66]&~m[102])|(~m[0]&m[66]&m[102]))&~BiasedRNG[60])|((~m[0]&~m[66]&m[102])|(m[0]&~m[66]&m[102])|(m[0]&m[66]&m[102]));
    m[30] = (((~m[1]&~m[61]&~m[97])|(m[1]&m[61]&~m[97]))&BiasedRNG[61])|(((m[1]&~m[61]&~m[97])|(~m[1]&m[61]&m[97]))&~BiasedRNG[61])|((~m[1]&~m[61]&m[97])|(m[1]&~m[61]&m[97])|(m[1]&m[61]&m[97]));
    m[31] = (((~m[1]&~m[67]&~m[103])|(m[1]&m[67]&~m[103]))&BiasedRNG[62])|(((m[1]&~m[67]&~m[103])|(~m[1]&m[67]&m[103]))&~BiasedRNG[62])|((~m[1]&~m[67]&m[103])|(m[1]&~m[67]&m[103])|(m[1]&m[67]&m[103]));
    m[36] = (((~m[2]&~m[62]&~m[98])|(m[2]&m[62]&~m[98]))&BiasedRNG[63])|(((m[2]&~m[62]&~m[98])|(~m[2]&m[62]&m[98]))&~BiasedRNG[63])|((~m[2]&~m[62]&m[98])|(m[2]&~m[62]&m[98])|(m[2]&m[62]&m[98]));
    m[37] = (((~m[2]&~m[68]&~m[104])|(m[2]&m[68]&~m[104]))&BiasedRNG[64])|(((m[2]&~m[68]&~m[104])|(~m[2]&m[68]&m[104]))&~BiasedRNG[64])|((~m[2]&~m[68]&m[104])|(m[2]&~m[68]&m[104])|(m[2]&m[68]&m[104]));
    m[42] = (((~m[3]&~m[63]&~m[99])|(m[3]&m[63]&~m[99]))&BiasedRNG[65])|(((m[3]&~m[63]&~m[99])|(~m[3]&m[63]&m[99]))&~BiasedRNG[65])|((~m[3]&~m[63]&m[99])|(m[3]&~m[63]&m[99])|(m[3]&m[63]&m[99]));
    m[43] = (((~m[3]&~m[69]&~m[105])|(m[3]&m[69]&~m[105]))&BiasedRNG[66])|(((m[3]&~m[69]&~m[105])|(~m[3]&m[69]&m[105]))&~BiasedRNG[66])|((~m[3]&~m[69]&m[105])|(m[3]&~m[69]&m[105])|(m[3]&m[69]&m[105]));
    m[48] = (((~m[4]&~m[64]&~m[100])|(m[4]&m[64]&~m[100]))&BiasedRNG[67])|(((m[4]&~m[64]&~m[100])|(~m[4]&m[64]&m[100]))&~BiasedRNG[67])|((~m[4]&~m[64]&m[100])|(m[4]&~m[64]&m[100])|(m[4]&m[64]&m[100]));
    m[49] = (((~m[4]&~m[70]&~m[106])|(m[4]&m[70]&~m[106]))&BiasedRNG[68])|(((m[4]&~m[70]&~m[106])|(~m[4]&m[70]&m[106]))&~BiasedRNG[68])|((~m[4]&~m[70]&m[106])|(m[4]&~m[70]&m[106])|(m[4]&m[70]&m[106]));
    m[54] = (((~m[5]&~m[65]&~m[101])|(m[5]&m[65]&~m[101]))&BiasedRNG[69])|(((m[5]&~m[65]&~m[101])|(~m[5]&m[65]&m[101]))&~BiasedRNG[69])|((~m[5]&~m[65]&m[101])|(m[5]&~m[65]&m[101])|(m[5]&m[65]&m[101]));
    m[55] = (((~m[5]&~m[71]&~m[107])|(m[5]&m[71]&~m[107]))&BiasedRNG[70])|(((m[5]&~m[71]&~m[107])|(~m[5]&m[71]&m[107]))&~BiasedRNG[70])|((~m[5]&~m[71]&m[107])|(m[5]&~m[71]&m[107])|(m[5]&m[71]&m[107]));
    m[72] = (((~m[8]&~m[26]&~m[108])|(m[8]&m[26]&~m[108]))&BiasedRNG[71])|(((m[8]&~m[26]&~m[108])|(~m[8]&m[26]&m[108]))&~BiasedRNG[71])|((~m[8]&~m[26]&m[108])|(m[8]&~m[26]&m[108])|(m[8]&m[26]&m[108]));
    m[73] = (((~m[8]&~m[32]&~m[109])|(m[8]&m[32]&~m[109]))&BiasedRNG[72])|(((m[8]&~m[32]&~m[109])|(~m[8]&m[32]&m[109]))&~BiasedRNG[72])|((~m[8]&~m[32]&m[109])|(m[8]&~m[32]&m[109])|(m[8]&m[32]&m[109]));
    m[78] = (((~m[9]&~m[27]&~m[114])|(m[9]&m[27]&~m[114]))&BiasedRNG[73])|(((m[9]&~m[27]&~m[114])|(~m[9]&m[27]&m[114]))&~BiasedRNG[73])|((~m[9]&~m[27]&m[114])|(m[9]&~m[27]&m[114])|(m[9]&m[27]&m[114]));
    m[79] = (((~m[9]&~m[33]&~m[115])|(m[9]&m[33]&~m[115]))&BiasedRNG[74])|(((m[9]&~m[33]&~m[115])|(~m[9]&m[33]&m[115]))&~BiasedRNG[74])|((~m[9]&~m[33]&m[115])|(m[9]&~m[33]&m[115])|(m[9]&m[33]&m[115]));
    m[84] = (((~m[10]&~m[28]&~m[120])|(m[10]&m[28]&~m[120]))&BiasedRNG[75])|(((m[10]&~m[28]&~m[120])|(~m[10]&m[28]&m[120]))&~BiasedRNG[75])|((~m[10]&~m[28]&m[120])|(m[10]&~m[28]&m[120])|(m[10]&m[28]&m[120]));
    m[85] = (((~m[10]&~m[34]&~m[121])|(m[10]&m[34]&~m[121]))&BiasedRNG[76])|(((m[10]&~m[34]&~m[121])|(~m[10]&m[34]&m[121]))&~BiasedRNG[76])|((~m[10]&~m[34]&m[121])|(m[10]&~m[34]&m[121])|(m[10]&m[34]&m[121]));
    m[90] = (((~m[11]&~m[29]&~m[126])|(m[11]&m[29]&~m[126]))&BiasedRNG[77])|(((m[11]&~m[29]&~m[126])|(~m[11]&m[29]&m[126]))&~BiasedRNG[77])|((~m[11]&~m[29]&m[126])|(m[11]&~m[29]&m[126])|(m[11]&m[29]&m[126]));
    m[91] = (((~m[11]&~m[35]&~m[127])|(m[11]&m[35]&~m[127]))&BiasedRNG[78])|(((m[11]&~m[35]&~m[127])|(~m[11]&m[35]&m[127]))&~BiasedRNG[78])|((~m[11]&~m[35]&m[127])|(m[11]&~m[35]&m[127])|(m[11]&m[35]&m[127]));
    m[110] = (((m[38]&~m[74]&m[168])|(~m[38]&m[74]&m[168]))&BiasedRNG[79])|(((m[38]&m[74]&~m[168]))&~BiasedRNG[79])|((m[38]&m[74]&m[168]));
    m[111] = (((m[44]&~m[75]&m[188])|(~m[44]&m[75]&m[188]))&BiasedRNG[80])|(((m[44]&m[75]&~m[188]))&~BiasedRNG[80])|((m[44]&m[75]&m[188]));
    m[112] = (((m[50]&~m[76]&m[213])|(~m[50]&m[76]&m[213]))&BiasedRNG[81])|(((m[50]&m[76]&~m[213]))&~BiasedRNG[81])|((m[50]&m[76]&m[213]));
    m[113] = (((m[56]&~m[77]&m[233])|(~m[56]&m[77]&m[233]))&BiasedRNG[82])|(((m[56]&m[77]&~m[233]))&~BiasedRNG[82])|((m[56]&m[77]&m[233]));
    m[116] = (((m[39]&~m[80]&m[193])|(~m[39]&m[80]&m[193]))&BiasedRNG[83])|(((m[39]&m[80]&~m[193]))&~BiasedRNG[83])|((m[39]&m[80]&m[193]));
    m[117] = (((m[45]&~m[81]&m[218])|(~m[45]&m[81]&m[218]))&BiasedRNG[84])|(((m[45]&m[81]&~m[218]))&~BiasedRNG[84])|((m[45]&m[81]&m[218]));
    m[118] = (((m[51]&~m[82]&m[238])|(~m[51]&m[82]&m[238]))&BiasedRNG[85])|(((m[51]&m[82]&~m[238]))&~BiasedRNG[85])|((m[51]&m[82]&m[238]));
    m[119] = (((m[57]&~m[83]&m[253])|(~m[57]&m[83]&m[253]))&BiasedRNG[86])|(((m[57]&m[83]&~m[253]))&~BiasedRNG[86])|((m[57]&m[83]&m[253]));
    m[122] = (((m[40]&~m[86]&m[223])|(~m[40]&m[86]&m[223]))&BiasedRNG[87])|(((m[40]&m[86]&~m[223]))&~BiasedRNG[87])|((m[40]&m[86]&m[223]));
    m[123] = (((m[46]&~m[87]&m[243])|(~m[46]&m[87]&m[243]))&BiasedRNG[88])|(((m[46]&m[87]&~m[243]))&~BiasedRNG[88])|((m[46]&m[87]&m[243]));
    m[124] = (((m[52]&~m[88]&m[258])|(~m[52]&m[88]&m[258]))&BiasedRNG[89])|(((m[52]&m[88]&~m[258]))&~BiasedRNG[89])|((m[52]&m[88]&m[258]));
    m[125] = (((m[58]&~m[89]&m[268])|(~m[58]&m[89]&m[268]))&BiasedRNG[90])|(((m[58]&m[89]&~m[268]))&~BiasedRNG[90])|((m[58]&m[89]&m[268]));
    m[128] = (((m[41]&~m[92]&m[248])|(~m[41]&m[92]&m[248]))&BiasedRNG[91])|(((m[41]&m[92]&~m[248]))&~BiasedRNG[91])|((m[41]&m[92]&m[248]));
    m[129] = (((m[47]&~m[93]&m[263])|(~m[47]&m[93]&m[263]))&BiasedRNG[92])|(((m[47]&m[93]&~m[263]))&~BiasedRNG[92])|((m[47]&m[93]&m[263]));
    m[130] = (((m[53]&~m[94]&m[273])|(~m[53]&m[94]&m[273]))&BiasedRNG[93])|(((m[53]&m[94]&~m[273]))&~BiasedRNG[93])|((m[53]&m[94]&m[273]));
    m[131] = (((m[59]&~m[95]&m[278])|(~m[59]&m[95]&m[278]))&BiasedRNG[94])|(((m[59]&m[95]&~m[278]))&~BiasedRNG[94])|((m[59]&m[95]&m[278]));
    m[132] = (((m[97]&~m[133]&~m[134]&~m[135]&~m[136])|(~m[97]&~m[133]&~m[134]&m[135]&~m[136])|(m[97]&m[133]&~m[134]&m[135]&~m[136])|(m[97]&~m[133]&m[134]&m[135]&~m[136])|(~m[97]&m[133]&~m[134]&~m[135]&m[136])|(~m[97]&~m[133]&m[134]&~m[135]&m[136])|(m[97]&m[133]&m[134]&~m[135]&m[136])|(~m[97]&m[133]&m[134]&m[135]&m[136]))&UnbiasedRNG[28])|((m[97]&~m[133]&~m[134]&m[135]&~m[136])|(~m[97]&~m[133]&~m[134]&~m[135]&m[136])|(m[97]&~m[133]&~m[134]&~m[135]&m[136])|(m[97]&m[133]&~m[134]&~m[135]&m[136])|(m[97]&~m[133]&m[134]&~m[135]&m[136])|(~m[97]&~m[133]&~m[134]&m[135]&m[136])|(m[97]&~m[133]&~m[134]&m[135]&m[136])|(~m[97]&m[133]&~m[134]&m[135]&m[136])|(m[97]&m[133]&~m[134]&m[135]&m[136])|(~m[97]&~m[133]&m[134]&m[135]&m[136])|(m[97]&~m[133]&m[134]&m[135]&m[136])|(m[97]&m[133]&m[134]&m[135]&m[136]));
    m[138] = (((m[103]&~m[137]&~m[139]&~m[140]&~m[141])|(~m[103]&~m[137]&~m[139]&m[140]&~m[141])|(m[103]&m[137]&~m[139]&m[140]&~m[141])|(m[103]&~m[137]&m[139]&m[140]&~m[141])|(~m[103]&m[137]&~m[139]&~m[140]&m[141])|(~m[103]&~m[137]&m[139]&~m[140]&m[141])|(m[103]&m[137]&m[139]&~m[140]&m[141])|(~m[103]&m[137]&m[139]&m[140]&m[141]))&UnbiasedRNG[29])|((m[103]&~m[137]&~m[139]&m[140]&~m[141])|(~m[103]&~m[137]&~m[139]&~m[140]&m[141])|(m[103]&~m[137]&~m[139]&~m[140]&m[141])|(m[103]&m[137]&~m[139]&~m[140]&m[141])|(m[103]&~m[137]&m[139]&~m[140]&m[141])|(~m[103]&~m[137]&~m[139]&m[140]&m[141])|(m[103]&~m[137]&~m[139]&m[140]&m[141])|(~m[103]&m[137]&~m[139]&m[140]&m[141])|(m[103]&m[137]&~m[139]&m[140]&m[141])|(~m[103]&~m[137]&m[139]&m[140]&m[141])|(m[103]&~m[137]&m[139]&m[140]&m[141])|(m[103]&m[137]&m[139]&m[140]&m[141]));
    m[143] = (((m[108]&~m[142]&~m[144]&~m[145]&~m[146])|(~m[108]&~m[142]&~m[144]&m[145]&~m[146])|(m[108]&m[142]&~m[144]&m[145]&~m[146])|(m[108]&~m[142]&m[144]&m[145]&~m[146])|(~m[108]&m[142]&~m[144]&~m[145]&m[146])|(~m[108]&~m[142]&m[144]&~m[145]&m[146])|(m[108]&m[142]&m[144]&~m[145]&m[146])|(~m[108]&m[142]&m[144]&m[145]&m[146]))&UnbiasedRNG[30])|((m[108]&~m[142]&~m[144]&m[145]&~m[146])|(~m[108]&~m[142]&~m[144]&~m[145]&m[146])|(m[108]&~m[142]&~m[144]&~m[145]&m[146])|(m[108]&m[142]&~m[144]&~m[145]&m[146])|(m[108]&~m[142]&m[144]&~m[145]&m[146])|(~m[108]&~m[142]&~m[144]&m[145]&m[146])|(m[108]&~m[142]&~m[144]&m[145]&m[146])|(~m[108]&m[142]&~m[144]&m[145]&m[146])|(m[108]&m[142]&~m[144]&m[145]&m[146])|(~m[108]&~m[142]&m[144]&m[145]&m[146])|(m[108]&~m[142]&m[144]&m[145]&m[146])|(m[108]&m[142]&m[144]&m[145]&m[146]));
    m[148] = (((m[104]&~m[147]&~m[149]&~m[150]&~m[151])|(~m[104]&~m[147]&~m[149]&m[150]&~m[151])|(m[104]&m[147]&~m[149]&m[150]&~m[151])|(m[104]&~m[147]&m[149]&m[150]&~m[151])|(~m[104]&m[147]&~m[149]&~m[150]&m[151])|(~m[104]&~m[147]&m[149]&~m[150]&m[151])|(m[104]&m[147]&m[149]&~m[150]&m[151])|(~m[104]&m[147]&m[149]&m[150]&m[151]))&UnbiasedRNG[31])|((m[104]&~m[147]&~m[149]&m[150]&~m[151])|(~m[104]&~m[147]&~m[149]&~m[150]&m[151])|(m[104]&~m[147]&~m[149]&~m[150]&m[151])|(m[104]&m[147]&~m[149]&~m[150]&m[151])|(m[104]&~m[147]&m[149]&~m[150]&m[151])|(~m[104]&~m[147]&~m[149]&m[150]&m[151])|(m[104]&~m[147]&~m[149]&m[150]&m[151])|(~m[104]&m[147]&~m[149]&m[150]&m[151])|(m[104]&m[147]&~m[149]&m[150]&m[151])|(~m[104]&~m[147]&m[149]&m[150]&m[151])|(m[104]&~m[147]&m[149]&m[150]&m[151])|(m[104]&m[147]&m[149]&m[150]&m[151]));
    m[153] = (((m[109]&~m[152]&~m[154]&~m[155]&~m[156])|(~m[109]&~m[152]&~m[154]&m[155]&~m[156])|(m[109]&m[152]&~m[154]&m[155]&~m[156])|(m[109]&~m[152]&m[154]&m[155]&~m[156])|(~m[109]&m[152]&~m[154]&~m[155]&m[156])|(~m[109]&~m[152]&m[154]&~m[155]&m[156])|(m[109]&m[152]&m[154]&~m[155]&m[156])|(~m[109]&m[152]&m[154]&m[155]&m[156]))&UnbiasedRNG[32])|((m[109]&~m[152]&~m[154]&m[155]&~m[156])|(~m[109]&~m[152]&~m[154]&~m[155]&m[156])|(m[109]&~m[152]&~m[154]&~m[155]&m[156])|(m[109]&m[152]&~m[154]&~m[155]&m[156])|(m[109]&~m[152]&m[154]&~m[155]&m[156])|(~m[109]&~m[152]&~m[154]&m[155]&m[156])|(m[109]&~m[152]&~m[154]&m[155]&m[156])|(~m[109]&m[152]&~m[154]&m[155]&m[156])|(m[109]&m[152]&~m[154]&m[155]&m[156])|(~m[109]&~m[152]&m[154]&m[155]&m[156])|(m[109]&~m[152]&m[154]&m[155]&m[156])|(m[109]&m[152]&m[154]&m[155]&m[156]));
    m[158] = (((m[114]&~m[157]&~m[159]&~m[160]&~m[161])|(~m[114]&~m[157]&~m[159]&m[160]&~m[161])|(m[114]&m[157]&~m[159]&m[160]&~m[161])|(m[114]&~m[157]&m[159]&m[160]&~m[161])|(~m[114]&m[157]&~m[159]&~m[160]&m[161])|(~m[114]&~m[157]&m[159]&~m[160]&m[161])|(m[114]&m[157]&m[159]&~m[160]&m[161])|(~m[114]&m[157]&m[159]&m[160]&m[161]))&UnbiasedRNG[33])|((m[114]&~m[157]&~m[159]&m[160]&~m[161])|(~m[114]&~m[157]&~m[159]&~m[160]&m[161])|(m[114]&~m[157]&~m[159]&~m[160]&m[161])|(m[114]&m[157]&~m[159]&~m[160]&m[161])|(m[114]&~m[157]&m[159]&~m[160]&m[161])|(~m[114]&~m[157]&~m[159]&m[160]&m[161])|(m[114]&~m[157]&~m[159]&m[160]&m[161])|(~m[114]&m[157]&~m[159]&m[160]&m[161])|(m[114]&m[157]&~m[159]&m[160]&m[161])|(~m[114]&~m[157]&m[159]&m[160]&m[161])|(m[114]&~m[157]&m[159]&m[160]&m[161])|(m[114]&m[157]&m[159]&m[160]&m[161]));
    m[163] = (((m[105]&~m[162]&~m[164]&~m[165]&~m[166])|(~m[105]&~m[162]&~m[164]&m[165]&~m[166])|(m[105]&m[162]&~m[164]&m[165]&~m[166])|(m[105]&~m[162]&m[164]&m[165]&~m[166])|(~m[105]&m[162]&~m[164]&~m[165]&m[166])|(~m[105]&~m[162]&m[164]&~m[165]&m[166])|(m[105]&m[162]&m[164]&~m[165]&m[166])|(~m[105]&m[162]&m[164]&m[165]&m[166]))&UnbiasedRNG[34])|((m[105]&~m[162]&~m[164]&m[165]&~m[166])|(~m[105]&~m[162]&~m[164]&~m[165]&m[166])|(m[105]&~m[162]&~m[164]&~m[165]&m[166])|(m[105]&m[162]&~m[164]&~m[165]&m[166])|(m[105]&~m[162]&m[164]&~m[165]&m[166])|(~m[105]&~m[162]&~m[164]&m[165]&m[166])|(m[105]&~m[162]&~m[164]&m[165]&m[166])|(~m[105]&m[162]&~m[164]&m[165]&m[166])|(m[105]&m[162]&~m[164]&m[165]&m[166])|(~m[105]&~m[162]&m[164]&m[165]&m[166])|(m[105]&~m[162]&m[164]&m[165]&m[166])|(m[105]&m[162]&m[164]&m[165]&m[166]));
    m[169] = (((m[156]&~m[167]&~m[168]&~m[170]&~m[171])|(~m[156]&~m[167]&~m[168]&m[170]&~m[171])|(m[156]&m[167]&~m[168]&m[170]&~m[171])|(m[156]&~m[167]&m[168]&m[170]&~m[171])|(~m[156]&m[167]&~m[168]&~m[170]&m[171])|(~m[156]&~m[167]&m[168]&~m[170]&m[171])|(m[156]&m[167]&m[168]&~m[170]&m[171])|(~m[156]&m[167]&m[168]&m[170]&m[171]))&UnbiasedRNG[35])|((m[156]&~m[167]&~m[168]&m[170]&~m[171])|(~m[156]&~m[167]&~m[168]&~m[170]&m[171])|(m[156]&~m[167]&~m[168]&~m[170]&m[171])|(m[156]&m[167]&~m[168]&~m[170]&m[171])|(m[156]&~m[167]&m[168]&~m[170]&m[171])|(~m[156]&~m[167]&~m[168]&m[170]&m[171])|(m[156]&~m[167]&~m[168]&m[170]&m[171])|(~m[156]&m[167]&~m[168]&m[170]&m[171])|(m[156]&m[167]&~m[168]&m[170]&m[171])|(~m[156]&~m[167]&m[168]&m[170]&m[171])|(m[156]&~m[167]&m[168]&m[170]&m[171])|(m[156]&m[167]&m[168]&m[170]&m[171]));
    m[173] = (((m[115]&~m[172]&~m[174]&~m[175]&~m[176])|(~m[115]&~m[172]&~m[174]&m[175]&~m[176])|(m[115]&m[172]&~m[174]&m[175]&~m[176])|(m[115]&~m[172]&m[174]&m[175]&~m[176])|(~m[115]&m[172]&~m[174]&~m[175]&m[176])|(~m[115]&~m[172]&m[174]&~m[175]&m[176])|(m[115]&m[172]&m[174]&~m[175]&m[176])|(~m[115]&m[172]&m[174]&m[175]&m[176]))&UnbiasedRNG[36])|((m[115]&~m[172]&~m[174]&m[175]&~m[176])|(~m[115]&~m[172]&~m[174]&~m[175]&m[176])|(m[115]&~m[172]&~m[174]&~m[175]&m[176])|(m[115]&m[172]&~m[174]&~m[175]&m[176])|(m[115]&~m[172]&m[174]&~m[175]&m[176])|(~m[115]&~m[172]&~m[174]&m[175]&m[176])|(m[115]&~m[172]&~m[174]&m[175]&m[176])|(~m[115]&m[172]&~m[174]&m[175]&m[176])|(m[115]&m[172]&~m[174]&m[175]&m[176])|(~m[115]&~m[172]&m[174]&m[175]&m[176])|(m[115]&~m[172]&m[174]&m[175]&m[176])|(m[115]&m[172]&m[174]&m[175]&m[176]));
    m[178] = (((m[120]&~m[177]&~m[179]&~m[180]&~m[181])|(~m[120]&~m[177]&~m[179]&m[180]&~m[181])|(m[120]&m[177]&~m[179]&m[180]&~m[181])|(m[120]&~m[177]&m[179]&m[180]&~m[181])|(~m[120]&m[177]&~m[179]&~m[180]&m[181])|(~m[120]&~m[177]&m[179]&~m[180]&m[181])|(m[120]&m[177]&m[179]&~m[180]&m[181])|(~m[120]&m[177]&m[179]&m[180]&m[181]))&UnbiasedRNG[37])|((m[120]&~m[177]&~m[179]&m[180]&~m[181])|(~m[120]&~m[177]&~m[179]&~m[180]&m[181])|(m[120]&~m[177]&~m[179]&~m[180]&m[181])|(m[120]&m[177]&~m[179]&~m[180]&m[181])|(m[120]&~m[177]&m[179]&~m[180]&m[181])|(~m[120]&~m[177]&~m[179]&m[180]&m[181])|(m[120]&~m[177]&~m[179]&m[180]&m[181])|(~m[120]&m[177]&~m[179]&m[180]&m[181])|(m[120]&m[177]&~m[179]&m[180]&m[181])|(~m[120]&~m[177]&m[179]&m[180]&m[181])|(m[120]&~m[177]&m[179]&m[180]&m[181])|(m[120]&m[177]&m[179]&m[180]&m[181]));
    m[183] = (((m[106]&~m[182]&~m[184]&~m[185]&~m[186])|(~m[106]&~m[182]&~m[184]&m[185]&~m[186])|(m[106]&m[182]&~m[184]&m[185]&~m[186])|(m[106]&~m[182]&m[184]&m[185]&~m[186])|(~m[106]&m[182]&~m[184]&~m[185]&m[186])|(~m[106]&~m[182]&m[184]&~m[185]&m[186])|(m[106]&m[182]&m[184]&~m[185]&m[186])|(~m[106]&m[182]&m[184]&m[185]&m[186]))&UnbiasedRNG[38])|((m[106]&~m[182]&~m[184]&m[185]&~m[186])|(~m[106]&~m[182]&~m[184]&~m[185]&m[186])|(m[106]&~m[182]&~m[184]&~m[185]&m[186])|(m[106]&m[182]&~m[184]&~m[185]&m[186])|(m[106]&~m[182]&m[184]&~m[185]&m[186])|(~m[106]&~m[182]&~m[184]&m[185]&m[186])|(m[106]&~m[182]&~m[184]&m[185]&m[186])|(~m[106]&m[182]&~m[184]&m[185]&m[186])|(m[106]&m[182]&~m[184]&m[185]&m[186])|(~m[106]&~m[182]&m[184]&m[185]&m[186])|(m[106]&~m[182]&m[184]&m[185]&m[186])|(m[106]&m[182]&m[184]&m[185]&m[186]));
    m[189] = (((m[171]&~m[187]&~m[188]&~m[190]&~m[191])|(~m[171]&~m[187]&~m[188]&m[190]&~m[191])|(m[171]&m[187]&~m[188]&m[190]&~m[191])|(m[171]&~m[187]&m[188]&m[190]&~m[191])|(~m[171]&m[187]&~m[188]&~m[190]&m[191])|(~m[171]&~m[187]&m[188]&~m[190]&m[191])|(m[171]&m[187]&m[188]&~m[190]&m[191])|(~m[171]&m[187]&m[188]&m[190]&m[191]))&UnbiasedRNG[39])|((m[171]&~m[187]&~m[188]&m[190]&~m[191])|(~m[171]&~m[187]&~m[188]&~m[190]&m[191])|(m[171]&~m[187]&~m[188]&~m[190]&m[191])|(m[171]&m[187]&~m[188]&~m[190]&m[191])|(m[171]&~m[187]&m[188]&~m[190]&m[191])|(~m[171]&~m[187]&~m[188]&m[190]&m[191])|(m[171]&~m[187]&~m[188]&m[190]&m[191])|(~m[171]&m[187]&~m[188]&m[190]&m[191])|(m[171]&m[187]&~m[188]&m[190]&m[191])|(~m[171]&~m[187]&m[188]&m[190]&m[191])|(m[171]&~m[187]&m[188]&m[190]&m[191])|(m[171]&m[187]&m[188]&m[190]&m[191]));
    m[194] = (((m[176]&~m[192]&~m[193]&~m[195]&~m[196])|(~m[176]&~m[192]&~m[193]&m[195]&~m[196])|(m[176]&m[192]&~m[193]&m[195]&~m[196])|(m[176]&~m[192]&m[193]&m[195]&~m[196])|(~m[176]&m[192]&~m[193]&~m[195]&m[196])|(~m[176]&~m[192]&m[193]&~m[195]&m[196])|(m[176]&m[192]&m[193]&~m[195]&m[196])|(~m[176]&m[192]&m[193]&m[195]&m[196]))&UnbiasedRNG[40])|((m[176]&~m[192]&~m[193]&m[195]&~m[196])|(~m[176]&~m[192]&~m[193]&~m[195]&m[196])|(m[176]&~m[192]&~m[193]&~m[195]&m[196])|(m[176]&m[192]&~m[193]&~m[195]&m[196])|(m[176]&~m[192]&m[193]&~m[195]&m[196])|(~m[176]&~m[192]&~m[193]&m[195]&m[196])|(m[176]&~m[192]&~m[193]&m[195]&m[196])|(~m[176]&m[192]&~m[193]&m[195]&m[196])|(m[176]&m[192]&~m[193]&m[195]&m[196])|(~m[176]&~m[192]&m[193]&m[195]&m[196])|(m[176]&~m[192]&m[193]&m[195]&m[196])|(m[176]&m[192]&m[193]&m[195]&m[196]));
    m[198] = (((m[121]&~m[197]&~m[199]&~m[200]&~m[201])|(~m[121]&~m[197]&~m[199]&m[200]&~m[201])|(m[121]&m[197]&~m[199]&m[200]&~m[201])|(m[121]&~m[197]&m[199]&m[200]&~m[201])|(~m[121]&m[197]&~m[199]&~m[200]&m[201])|(~m[121]&~m[197]&m[199]&~m[200]&m[201])|(m[121]&m[197]&m[199]&~m[200]&m[201])|(~m[121]&m[197]&m[199]&m[200]&m[201]))&UnbiasedRNG[41])|((m[121]&~m[197]&~m[199]&m[200]&~m[201])|(~m[121]&~m[197]&~m[199]&~m[200]&m[201])|(m[121]&~m[197]&~m[199]&~m[200]&m[201])|(m[121]&m[197]&~m[199]&~m[200]&m[201])|(m[121]&~m[197]&m[199]&~m[200]&m[201])|(~m[121]&~m[197]&~m[199]&m[200]&m[201])|(m[121]&~m[197]&~m[199]&m[200]&m[201])|(~m[121]&m[197]&~m[199]&m[200]&m[201])|(m[121]&m[197]&~m[199]&m[200]&m[201])|(~m[121]&~m[197]&m[199]&m[200]&m[201])|(m[121]&~m[197]&m[199]&m[200]&m[201])|(m[121]&m[197]&m[199]&m[200]&m[201]));
    m[203] = (((m[126]&~m[202]&~m[204]&~m[205]&~m[206])|(~m[126]&~m[202]&~m[204]&m[205]&~m[206])|(m[126]&m[202]&~m[204]&m[205]&~m[206])|(m[126]&~m[202]&m[204]&m[205]&~m[206])|(~m[126]&m[202]&~m[204]&~m[205]&m[206])|(~m[126]&~m[202]&m[204]&~m[205]&m[206])|(m[126]&m[202]&m[204]&~m[205]&m[206])|(~m[126]&m[202]&m[204]&m[205]&m[206]))&UnbiasedRNG[42])|((m[126]&~m[202]&~m[204]&m[205]&~m[206])|(~m[126]&~m[202]&~m[204]&~m[205]&m[206])|(m[126]&~m[202]&~m[204]&~m[205]&m[206])|(m[126]&m[202]&~m[204]&~m[205]&m[206])|(m[126]&~m[202]&m[204]&~m[205]&m[206])|(~m[126]&~m[202]&~m[204]&m[205]&m[206])|(m[126]&~m[202]&~m[204]&m[205]&m[206])|(~m[126]&m[202]&~m[204]&m[205]&m[206])|(m[126]&m[202]&~m[204]&m[205]&m[206])|(~m[126]&~m[202]&m[204]&m[205]&m[206])|(m[126]&~m[202]&m[204]&m[205]&m[206])|(m[126]&m[202]&m[204]&m[205]&m[206]));
    m[208] = (((m[107]&~m[207]&~m[209]&~m[210]&~m[211])|(~m[107]&~m[207]&~m[209]&m[210]&~m[211])|(m[107]&m[207]&~m[209]&m[210]&~m[211])|(m[107]&~m[207]&m[209]&m[210]&~m[211])|(~m[107]&m[207]&~m[209]&~m[210]&m[211])|(~m[107]&~m[207]&m[209]&~m[210]&m[211])|(m[107]&m[207]&m[209]&~m[210]&m[211])|(~m[107]&m[207]&m[209]&m[210]&m[211]))&UnbiasedRNG[43])|((m[107]&~m[207]&~m[209]&m[210]&~m[211])|(~m[107]&~m[207]&~m[209]&~m[210]&m[211])|(m[107]&~m[207]&~m[209]&~m[210]&m[211])|(m[107]&m[207]&~m[209]&~m[210]&m[211])|(m[107]&~m[207]&m[209]&~m[210]&m[211])|(~m[107]&~m[207]&~m[209]&m[210]&m[211])|(m[107]&~m[207]&~m[209]&m[210]&m[211])|(~m[107]&m[207]&~m[209]&m[210]&m[211])|(m[107]&m[207]&~m[209]&m[210]&m[211])|(~m[107]&~m[207]&m[209]&m[210]&m[211])|(m[107]&~m[207]&m[209]&m[210]&m[211])|(m[107]&m[207]&m[209]&m[210]&m[211]));
    m[214] = (((m[191]&~m[212]&~m[213]&~m[215]&~m[216])|(~m[191]&~m[212]&~m[213]&m[215]&~m[216])|(m[191]&m[212]&~m[213]&m[215]&~m[216])|(m[191]&~m[212]&m[213]&m[215]&~m[216])|(~m[191]&m[212]&~m[213]&~m[215]&m[216])|(~m[191]&~m[212]&m[213]&~m[215]&m[216])|(m[191]&m[212]&m[213]&~m[215]&m[216])|(~m[191]&m[212]&m[213]&m[215]&m[216]))&UnbiasedRNG[44])|((m[191]&~m[212]&~m[213]&m[215]&~m[216])|(~m[191]&~m[212]&~m[213]&~m[215]&m[216])|(m[191]&~m[212]&~m[213]&~m[215]&m[216])|(m[191]&m[212]&~m[213]&~m[215]&m[216])|(m[191]&~m[212]&m[213]&~m[215]&m[216])|(~m[191]&~m[212]&~m[213]&m[215]&m[216])|(m[191]&~m[212]&~m[213]&m[215]&m[216])|(~m[191]&m[212]&~m[213]&m[215]&m[216])|(m[191]&m[212]&~m[213]&m[215]&m[216])|(~m[191]&~m[212]&m[213]&m[215]&m[216])|(m[191]&~m[212]&m[213]&m[215]&m[216])|(m[191]&m[212]&m[213]&m[215]&m[216]));
    m[219] = (((m[196]&~m[217]&~m[218]&~m[220]&~m[221])|(~m[196]&~m[217]&~m[218]&m[220]&~m[221])|(m[196]&m[217]&~m[218]&m[220]&~m[221])|(m[196]&~m[217]&m[218]&m[220]&~m[221])|(~m[196]&m[217]&~m[218]&~m[220]&m[221])|(~m[196]&~m[217]&m[218]&~m[220]&m[221])|(m[196]&m[217]&m[218]&~m[220]&m[221])|(~m[196]&m[217]&m[218]&m[220]&m[221]))&UnbiasedRNG[45])|((m[196]&~m[217]&~m[218]&m[220]&~m[221])|(~m[196]&~m[217]&~m[218]&~m[220]&m[221])|(m[196]&~m[217]&~m[218]&~m[220]&m[221])|(m[196]&m[217]&~m[218]&~m[220]&m[221])|(m[196]&~m[217]&m[218]&~m[220]&m[221])|(~m[196]&~m[217]&~m[218]&m[220]&m[221])|(m[196]&~m[217]&~m[218]&m[220]&m[221])|(~m[196]&m[217]&~m[218]&m[220]&m[221])|(m[196]&m[217]&~m[218]&m[220]&m[221])|(~m[196]&~m[217]&m[218]&m[220]&m[221])|(m[196]&~m[217]&m[218]&m[220]&m[221])|(m[196]&m[217]&m[218]&m[220]&m[221]));
    m[224] = (((m[201]&~m[222]&~m[223]&~m[225]&~m[226])|(~m[201]&~m[222]&~m[223]&m[225]&~m[226])|(m[201]&m[222]&~m[223]&m[225]&~m[226])|(m[201]&~m[222]&m[223]&m[225]&~m[226])|(~m[201]&m[222]&~m[223]&~m[225]&m[226])|(~m[201]&~m[222]&m[223]&~m[225]&m[226])|(m[201]&m[222]&m[223]&~m[225]&m[226])|(~m[201]&m[222]&m[223]&m[225]&m[226]))&UnbiasedRNG[46])|((m[201]&~m[222]&~m[223]&m[225]&~m[226])|(~m[201]&~m[222]&~m[223]&~m[225]&m[226])|(m[201]&~m[222]&~m[223]&~m[225]&m[226])|(m[201]&m[222]&~m[223]&~m[225]&m[226])|(m[201]&~m[222]&m[223]&~m[225]&m[226])|(~m[201]&~m[222]&~m[223]&m[225]&m[226])|(m[201]&~m[222]&~m[223]&m[225]&m[226])|(~m[201]&m[222]&~m[223]&m[225]&m[226])|(m[201]&m[222]&~m[223]&m[225]&m[226])|(~m[201]&~m[222]&m[223]&m[225]&m[226])|(m[201]&~m[222]&m[223]&m[225]&m[226])|(m[201]&m[222]&m[223]&m[225]&m[226]));
    m[228] = (((m[127]&~m[227]&~m[229]&~m[230]&~m[231])|(~m[127]&~m[227]&~m[229]&m[230]&~m[231])|(m[127]&m[227]&~m[229]&m[230]&~m[231])|(m[127]&~m[227]&m[229]&m[230]&~m[231])|(~m[127]&m[227]&~m[229]&~m[230]&m[231])|(~m[127]&~m[227]&m[229]&~m[230]&m[231])|(m[127]&m[227]&m[229]&~m[230]&m[231])|(~m[127]&m[227]&m[229]&m[230]&m[231]))&UnbiasedRNG[47])|((m[127]&~m[227]&~m[229]&m[230]&~m[231])|(~m[127]&~m[227]&~m[229]&~m[230]&m[231])|(m[127]&~m[227]&~m[229]&~m[230]&m[231])|(m[127]&m[227]&~m[229]&~m[230]&m[231])|(m[127]&~m[227]&m[229]&~m[230]&m[231])|(~m[127]&~m[227]&~m[229]&m[230]&m[231])|(m[127]&~m[227]&~m[229]&m[230]&m[231])|(~m[127]&m[227]&~m[229]&m[230]&m[231])|(m[127]&m[227]&~m[229]&m[230]&m[231])|(~m[127]&~m[227]&m[229]&m[230]&m[231])|(m[127]&~m[227]&m[229]&m[230]&m[231])|(m[127]&m[227]&m[229]&m[230]&m[231]));
    m[234] = (((m[216]&~m[232]&~m[233]&~m[235]&~m[236])|(~m[216]&~m[232]&~m[233]&m[235]&~m[236])|(m[216]&m[232]&~m[233]&m[235]&~m[236])|(m[216]&~m[232]&m[233]&m[235]&~m[236])|(~m[216]&m[232]&~m[233]&~m[235]&m[236])|(~m[216]&~m[232]&m[233]&~m[235]&m[236])|(m[216]&m[232]&m[233]&~m[235]&m[236])|(~m[216]&m[232]&m[233]&m[235]&m[236]))&UnbiasedRNG[48])|((m[216]&~m[232]&~m[233]&m[235]&~m[236])|(~m[216]&~m[232]&~m[233]&~m[235]&m[236])|(m[216]&~m[232]&~m[233]&~m[235]&m[236])|(m[216]&m[232]&~m[233]&~m[235]&m[236])|(m[216]&~m[232]&m[233]&~m[235]&m[236])|(~m[216]&~m[232]&~m[233]&m[235]&m[236])|(m[216]&~m[232]&~m[233]&m[235]&m[236])|(~m[216]&m[232]&~m[233]&m[235]&m[236])|(m[216]&m[232]&~m[233]&m[235]&m[236])|(~m[216]&~m[232]&m[233]&m[235]&m[236])|(m[216]&~m[232]&m[233]&m[235]&m[236])|(m[216]&m[232]&m[233]&m[235]&m[236]));
    m[239] = (((m[221]&~m[237]&~m[238]&~m[240]&~m[241])|(~m[221]&~m[237]&~m[238]&m[240]&~m[241])|(m[221]&m[237]&~m[238]&m[240]&~m[241])|(m[221]&~m[237]&m[238]&m[240]&~m[241])|(~m[221]&m[237]&~m[238]&~m[240]&m[241])|(~m[221]&~m[237]&m[238]&~m[240]&m[241])|(m[221]&m[237]&m[238]&~m[240]&m[241])|(~m[221]&m[237]&m[238]&m[240]&m[241]))&UnbiasedRNG[49])|((m[221]&~m[237]&~m[238]&m[240]&~m[241])|(~m[221]&~m[237]&~m[238]&~m[240]&m[241])|(m[221]&~m[237]&~m[238]&~m[240]&m[241])|(m[221]&m[237]&~m[238]&~m[240]&m[241])|(m[221]&~m[237]&m[238]&~m[240]&m[241])|(~m[221]&~m[237]&~m[238]&m[240]&m[241])|(m[221]&~m[237]&~m[238]&m[240]&m[241])|(~m[221]&m[237]&~m[238]&m[240]&m[241])|(m[221]&m[237]&~m[238]&m[240]&m[241])|(~m[221]&~m[237]&m[238]&m[240]&m[241])|(m[221]&~m[237]&m[238]&m[240]&m[241])|(m[221]&m[237]&m[238]&m[240]&m[241]));
    m[244] = (((m[226]&~m[242]&~m[243]&~m[245]&~m[246])|(~m[226]&~m[242]&~m[243]&m[245]&~m[246])|(m[226]&m[242]&~m[243]&m[245]&~m[246])|(m[226]&~m[242]&m[243]&m[245]&~m[246])|(~m[226]&m[242]&~m[243]&~m[245]&m[246])|(~m[226]&~m[242]&m[243]&~m[245]&m[246])|(m[226]&m[242]&m[243]&~m[245]&m[246])|(~m[226]&m[242]&m[243]&m[245]&m[246]))&UnbiasedRNG[50])|((m[226]&~m[242]&~m[243]&m[245]&~m[246])|(~m[226]&~m[242]&~m[243]&~m[245]&m[246])|(m[226]&~m[242]&~m[243]&~m[245]&m[246])|(m[226]&m[242]&~m[243]&~m[245]&m[246])|(m[226]&~m[242]&m[243]&~m[245]&m[246])|(~m[226]&~m[242]&~m[243]&m[245]&m[246])|(m[226]&~m[242]&~m[243]&m[245]&m[246])|(~m[226]&m[242]&~m[243]&m[245]&m[246])|(m[226]&m[242]&~m[243]&m[245]&m[246])|(~m[226]&~m[242]&m[243]&m[245]&m[246])|(m[226]&~m[242]&m[243]&m[245]&m[246])|(m[226]&m[242]&m[243]&m[245]&m[246]));
    m[249] = (((m[231]&~m[247]&~m[248]&~m[250]&~m[251])|(~m[231]&~m[247]&~m[248]&m[250]&~m[251])|(m[231]&m[247]&~m[248]&m[250]&~m[251])|(m[231]&~m[247]&m[248]&m[250]&~m[251])|(~m[231]&m[247]&~m[248]&~m[250]&m[251])|(~m[231]&~m[247]&m[248]&~m[250]&m[251])|(m[231]&m[247]&m[248]&~m[250]&m[251])|(~m[231]&m[247]&m[248]&m[250]&m[251]))&UnbiasedRNG[51])|((m[231]&~m[247]&~m[248]&m[250]&~m[251])|(~m[231]&~m[247]&~m[248]&~m[250]&m[251])|(m[231]&~m[247]&~m[248]&~m[250]&m[251])|(m[231]&m[247]&~m[248]&~m[250]&m[251])|(m[231]&~m[247]&m[248]&~m[250]&m[251])|(~m[231]&~m[247]&~m[248]&m[250]&m[251])|(m[231]&~m[247]&~m[248]&m[250]&m[251])|(~m[231]&m[247]&~m[248]&m[250]&m[251])|(m[231]&m[247]&~m[248]&m[250]&m[251])|(~m[231]&~m[247]&m[248]&m[250]&m[251])|(m[231]&~m[247]&m[248]&m[250]&m[251])|(m[231]&m[247]&m[248]&m[250]&m[251]));
    m[254] = (((m[241]&~m[252]&~m[253]&~m[255]&~m[256])|(~m[241]&~m[252]&~m[253]&m[255]&~m[256])|(m[241]&m[252]&~m[253]&m[255]&~m[256])|(m[241]&~m[252]&m[253]&m[255]&~m[256])|(~m[241]&m[252]&~m[253]&~m[255]&m[256])|(~m[241]&~m[252]&m[253]&~m[255]&m[256])|(m[241]&m[252]&m[253]&~m[255]&m[256])|(~m[241]&m[252]&m[253]&m[255]&m[256]))&UnbiasedRNG[52])|((m[241]&~m[252]&~m[253]&m[255]&~m[256])|(~m[241]&~m[252]&~m[253]&~m[255]&m[256])|(m[241]&~m[252]&~m[253]&~m[255]&m[256])|(m[241]&m[252]&~m[253]&~m[255]&m[256])|(m[241]&~m[252]&m[253]&~m[255]&m[256])|(~m[241]&~m[252]&~m[253]&m[255]&m[256])|(m[241]&~m[252]&~m[253]&m[255]&m[256])|(~m[241]&m[252]&~m[253]&m[255]&m[256])|(m[241]&m[252]&~m[253]&m[255]&m[256])|(~m[241]&~m[252]&m[253]&m[255]&m[256])|(m[241]&~m[252]&m[253]&m[255]&m[256])|(m[241]&m[252]&m[253]&m[255]&m[256]));
    m[259] = (((m[246]&~m[257]&~m[258]&~m[260]&~m[261])|(~m[246]&~m[257]&~m[258]&m[260]&~m[261])|(m[246]&m[257]&~m[258]&m[260]&~m[261])|(m[246]&~m[257]&m[258]&m[260]&~m[261])|(~m[246]&m[257]&~m[258]&~m[260]&m[261])|(~m[246]&~m[257]&m[258]&~m[260]&m[261])|(m[246]&m[257]&m[258]&~m[260]&m[261])|(~m[246]&m[257]&m[258]&m[260]&m[261]))&UnbiasedRNG[53])|((m[246]&~m[257]&~m[258]&m[260]&~m[261])|(~m[246]&~m[257]&~m[258]&~m[260]&m[261])|(m[246]&~m[257]&~m[258]&~m[260]&m[261])|(m[246]&m[257]&~m[258]&~m[260]&m[261])|(m[246]&~m[257]&m[258]&~m[260]&m[261])|(~m[246]&~m[257]&~m[258]&m[260]&m[261])|(m[246]&~m[257]&~m[258]&m[260]&m[261])|(~m[246]&m[257]&~m[258]&m[260]&m[261])|(m[246]&m[257]&~m[258]&m[260]&m[261])|(~m[246]&~m[257]&m[258]&m[260]&m[261])|(m[246]&~m[257]&m[258]&m[260]&m[261])|(m[246]&m[257]&m[258]&m[260]&m[261]));
    m[264] = (((m[251]&~m[262]&~m[263]&~m[265]&~m[266])|(~m[251]&~m[262]&~m[263]&m[265]&~m[266])|(m[251]&m[262]&~m[263]&m[265]&~m[266])|(m[251]&~m[262]&m[263]&m[265]&~m[266])|(~m[251]&m[262]&~m[263]&~m[265]&m[266])|(~m[251]&~m[262]&m[263]&~m[265]&m[266])|(m[251]&m[262]&m[263]&~m[265]&m[266])|(~m[251]&m[262]&m[263]&m[265]&m[266]))&UnbiasedRNG[54])|((m[251]&~m[262]&~m[263]&m[265]&~m[266])|(~m[251]&~m[262]&~m[263]&~m[265]&m[266])|(m[251]&~m[262]&~m[263]&~m[265]&m[266])|(m[251]&m[262]&~m[263]&~m[265]&m[266])|(m[251]&~m[262]&m[263]&~m[265]&m[266])|(~m[251]&~m[262]&~m[263]&m[265]&m[266])|(m[251]&~m[262]&~m[263]&m[265]&m[266])|(~m[251]&m[262]&~m[263]&m[265]&m[266])|(m[251]&m[262]&~m[263]&m[265]&m[266])|(~m[251]&~m[262]&m[263]&m[265]&m[266])|(m[251]&~m[262]&m[263]&m[265]&m[266])|(m[251]&m[262]&m[263]&m[265]&m[266]));
    m[269] = (((m[261]&~m[267]&~m[268]&~m[270]&~m[271])|(~m[261]&~m[267]&~m[268]&m[270]&~m[271])|(m[261]&m[267]&~m[268]&m[270]&~m[271])|(m[261]&~m[267]&m[268]&m[270]&~m[271])|(~m[261]&m[267]&~m[268]&~m[270]&m[271])|(~m[261]&~m[267]&m[268]&~m[270]&m[271])|(m[261]&m[267]&m[268]&~m[270]&m[271])|(~m[261]&m[267]&m[268]&m[270]&m[271]))&UnbiasedRNG[55])|((m[261]&~m[267]&~m[268]&m[270]&~m[271])|(~m[261]&~m[267]&~m[268]&~m[270]&m[271])|(m[261]&~m[267]&~m[268]&~m[270]&m[271])|(m[261]&m[267]&~m[268]&~m[270]&m[271])|(m[261]&~m[267]&m[268]&~m[270]&m[271])|(~m[261]&~m[267]&~m[268]&m[270]&m[271])|(m[261]&~m[267]&~m[268]&m[270]&m[271])|(~m[261]&m[267]&~m[268]&m[270]&m[271])|(m[261]&m[267]&~m[268]&m[270]&m[271])|(~m[261]&~m[267]&m[268]&m[270]&m[271])|(m[261]&~m[267]&m[268]&m[270]&m[271])|(m[261]&m[267]&m[268]&m[270]&m[271]));
    m[274] = (((m[266]&~m[272]&~m[273]&~m[275]&~m[276])|(~m[266]&~m[272]&~m[273]&m[275]&~m[276])|(m[266]&m[272]&~m[273]&m[275]&~m[276])|(m[266]&~m[272]&m[273]&m[275]&~m[276])|(~m[266]&m[272]&~m[273]&~m[275]&m[276])|(~m[266]&~m[272]&m[273]&~m[275]&m[276])|(m[266]&m[272]&m[273]&~m[275]&m[276])|(~m[266]&m[272]&m[273]&m[275]&m[276]))&UnbiasedRNG[56])|((m[266]&~m[272]&~m[273]&m[275]&~m[276])|(~m[266]&~m[272]&~m[273]&~m[275]&m[276])|(m[266]&~m[272]&~m[273]&~m[275]&m[276])|(m[266]&m[272]&~m[273]&~m[275]&m[276])|(m[266]&~m[272]&m[273]&~m[275]&m[276])|(~m[266]&~m[272]&~m[273]&m[275]&m[276])|(m[266]&~m[272]&~m[273]&m[275]&m[276])|(~m[266]&m[272]&~m[273]&m[275]&m[276])|(m[266]&m[272]&~m[273]&m[275]&m[276])|(~m[266]&~m[272]&m[273]&m[275]&m[276])|(m[266]&~m[272]&m[273]&m[275]&m[276])|(m[266]&m[272]&m[273]&m[275]&m[276]));
    m[279] = (((m[276]&~m[277]&~m[278]&~m[280]&~m[281])|(~m[276]&~m[277]&~m[278]&m[280]&~m[281])|(m[276]&m[277]&~m[278]&m[280]&~m[281])|(m[276]&~m[277]&m[278]&m[280]&~m[281])|(~m[276]&m[277]&~m[278]&~m[280]&m[281])|(~m[276]&~m[277]&m[278]&~m[280]&m[281])|(m[276]&m[277]&m[278]&~m[280]&m[281])|(~m[276]&m[277]&m[278]&m[280]&m[281]))&UnbiasedRNG[57])|((m[276]&~m[277]&~m[278]&m[280]&~m[281])|(~m[276]&~m[277]&~m[278]&~m[280]&m[281])|(m[276]&~m[277]&~m[278]&~m[280]&m[281])|(m[276]&m[277]&~m[278]&~m[280]&m[281])|(m[276]&~m[277]&m[278]&~m[280]&m[281])|(~m[276]&~m[277]&~m[278]&m[280]&m[281])|(m[276]&~m[277]&~m[278]&m[280]&m[281])|(~m[276]&m[277]&~m[278]&m[280]&m[281])|(m[276]&m[277]&~m[278]&m[280]&m[281])|(~m[276]&~m[277]&m[278]&m[280]&m[281])|(m[276]&~m[277]&m[278]&m[280]&m[281])|(m[276]&m[277]&m[278]&m[280]&m[281]));
end

always @(posedge color2_clk) begin
    m[60] = (((~m[6]&~m[24]&~m[96])|(m[6]&m[24]&~m[96]))&BiasedRNG[95])|(((m[6]&~m[24]&~m[96])|(~m[6]&m[24]&m[96]))&~BiasedRNG[95])|((~m[6]&~m[24]&m[96])|(m[6]&~m[24]&m[96])|(m[6]&m[24]&m[96]));
    m[61] = (((~m[6]&~m[30]&~m[97])|(m[6]&m[30]&~m[97]))&BiasedRNG[96])|(((m[6]&~m[30]&~m[97])|(~m[6]&m[30]&m[97]))&~BiasedRNG[96])|((~m[6]&~m[30]&m[97])|(m[6]&~m[30]&m[97])|(m[6]&m[30]&m[97]));
    m[66] = (((~m[7]&~m[25]&~m[102])|(m[7]&m[25]&~m[102]))&BiasedRNG[97])|(((m[7]&~m[25]&~m[102])|(~m[7]&m[25]&m[102]))&~BiasedRNG[97])|((~m[7]&~m[25]&m[102])|(m[7]&~m[25]&m[102])|(m[7]&m[25]&m[102]));
    m[67] = (((~m[7]&~m[31]&~m[103])|(m[7]&m[31]&~m[103]))&BiasedRNG[98])|(((m[7]&~m[31]&~m[103])|(~m[7]&m[31]&m[103]))&~BiasedRNG[98])|((~m[7]&~m[31]&m[103])|(m[7]&~m[31]&m[103])|(m[7]&m[31]&m[103]));
    m[74] = (((~m[20]&~m[38]&~m[110])|(m[20]&m[38]&~m[110]))&BiasedRNG[99])|(((m[20]&~m[38]&~m[110])|(~m[20]&m[38]&m[110]))&~BiasedRNG[99])|((~m[20]&~m[38]&m[110])|(m[20]&~m[38]&m[110])|(m[20]&m[38]&m[110]));
    m[75] = (((~m[20]&~m[44]&~m[111])|(m[20]&m[44]&~m[111]))&BiasedRNG[100])|(((m[20]&~m[44]&~m[111])|(~m[20]&m[44]&m[111]))&~BiasedRNG[100])|((~m[20]&~m[44]&m[111])|(m[20]&~m[44]&m[111])|(m[20]&m[44]&m[111]));
    m[76] = (((~m[20]&~m[50]&~m[112])|(m[20]&m[50]&~m[112]))&BiasedRNG[101])|(((m[20]&~m[50]&~m[112])|(~m[20]&m[50]&m[112]))&~BiasedRNG[101])|((~m[20]&~m[50]&m[112])|(m[20]&~m[50]&m[112])|(m[20]&m[50]&m[112]));
    m[77] = (((~m[20]&~m[56]&~m[113])|(m[20]&m[56]&~m[113]))&BiasedRNG[102])|(((m[20]&~m[56]&~m[113])|(~m[20]&m[56]&m[113]))&~BiasedRNG[102])|((~m[20]&~m[56]&m[113])|(m[20]&~m[56]&m[113])|(m[20]&m[56]&m[113]));
    m[80] = (((~m[21]&~m[39]&~m[116])|(m[21]&m[39]&~m[116]))&BiasedRNG[103])|(((m[21]&~m[39]&~m[116])|(~m[21]&m[39]&m[116]))&~BiasedRNG[103])|((~m[21]&~m[39]&m[116])|(m[21]&~m[39]&m[116])|(m[21]&m[39]&m[116]));
    m[81] = (((~m[21]&~m[45]&~m[117])|(m[21]&m[45]&~m[117]))&BiasedRNG[104])|(((m[21]&~m[45]&~m[117])|(~m[21]&m[45]&m[117]))&~BiasedRNG[104])|((~m[21]&~m[45]&m[117])|(m[21]&~m[45]&m[117])|(m[21]&m[45]&m[117]));
    m[82] = (((~m[21]&~m[51]&~m[118])|(m[21]&m[51]&~m[118]))&BiasedRNG[105])|(((m[21]&~m[51]&~m[118])|(~m[21]&m[51]&m[118]))&~BiasedRNG[105])|((~m[21]&~m[51]&m[118])|(m[21]&~m[51]&m[118])|(m[21]&m[51]&m[118]));
    m[83] = (((~m[21]&~m[57]&~m[119])|(m[21]&m[57]&~m[119]))&BiasedRNG[106])|(((m[21]&~m[57]&~m[119])|(~m[21]&m[57]&m[119]))&~BiasedRNG[106])|((~m[21]&~m[57]&m[119])|(m[21]&~m[57]&m[119])|(m[21]&m[57]&m[119]));
    m[86] = (((~m[22]&~m[40]&~m[122])|(m[22]&m[40]&~m[122]))&BiasedRNG[107])|(((m[22]&~m[40]&~m[122])|(~m[22]&m[40]&m[122]))&~BiasedRNG[107])|((~m[22]&~m[40]&m[122])|(m[22]&~m[40]&m[122])|(m[22]&m[40]&m[122]));
    m[87] = (((~m[22]&~m[46]&~m[123])|(m[22]&m[46]&~m[123]))&BiasedRNG[108])|(((m[22]&~m[46]&~m[123])|(~m[22]&m[46]&m[123]))&~BiasedRNG[108])|((~m[22]&~m[46]&m[123])|(m[22]&~m[46]&m[123])|(m[22]&m[46]&m[123]));
    m[88] = (((~m[22]&~m[52]&~m[124])|(m[22]&m[52]&~m[124]))&BiasedRNG[109])|(((m[22]&~m[52]&~m[124])|(~m[22]&m[52]&m[124]))&~BiasedRNG[109])|((~m[22]&~m[52]&m[124])|(m[22]&~m[52]&m[124])|(m[22]&m[52]&m[124]));
    m[89] = (((~m[22]&~m[58]&~m[125])|(m[22]&m[58]&~m[125]))&BiasedRNG[110])|(((m[22]&~m[58]&~m[125])|(~m[22]&m[58]&m[125]))&~BiasedRNG[110])|((~m[22]&~m[58]&m[125])|(m[22]&~m[58]&m[125])|(m[22]&m[58]&m[125]));
    m[92] = (((~m[23]&~m[41]&~m[128])|(m[23]&m[41]&~m[128]))&BiasedRNG[111])|(((m[23]&~m[41]&~m[128])|(~m[23]&m[41]&m[128]))&~BiasedRNG[111])|((~m[23]&~m[41]&m[128])|(m[23]&~m[41]&m[128])|(m[23]&m[41]&m[128]));
    m[93] = (((~m[23]&~m[47]&~m[129])|(m[23]&m[47]&~m[129]))&BiasedRNG[112])|(((m[23]&~m[47]&~m[129])|(~m[23]&m[47]&m[129]))&~BiasedRNG[112])|((~m[23]&~m[47]&m[129])|(m[23]&~m[47]&m[129])|(m[23]&m[47]&m[129]));
    m[94] = (((~m[23]&~m[53]&~m[130])|(m[23]&m[53]&~m[130]))&BiasedRNG[113])|(((m[23]&~m[53]&~m[130])|(~m[23]&m[53]&m[130]))&~BiasedRNG[113])|((~m[23]&~m[53]&m[130])|(m[23]&~m[53]&m[130])|(m[23]&m[53]&m[130]));
    m[95] = (((~m[23]&~m[59]&~m[131])|(m[23]&m[59]&~m[131]))&BiasedRNG[114])|(((m[23]&~m[59]&~m[131])|(~m[23]&m[59]&m[131]))&~BiasedRNG[114])|((~m[23]&~m[59]&m[131])|(m[23]&~m[59]&m[131])|(m[23]&m[59]&m[131]));
    m[98] = (((m[36]&~m[62]&m[137])|(~m[36]&m[62]&m[137]))&BiasedRNG[115])|(((m[36]&m[62]&~m[137]))&~BiasedRNG[115])|((m[36]&m[62]&m[137]));
    m[99] = (((m[42]&~m[63]&m[147])|(~m[42]&m[63]&m[147]))&BiasedRNG[116])|(((m[42]&m[63]&~m[147]))&~BiasedRNG[116])|((m[42]&m[63]&m[147]));
    m[100] = (((m[48]&~m[64]&m[162])|(~m[48]&m[64]&m[162]))&BiasedRNG[117])|(((m[48]&m[64]&~m[162]))&~BiasedRNG[117])|((m[48]&m[64]&m[162]));
    m[101] = (((m[54]&~m[65]&m[182])|(~m[54]&m[65]&m[182]))&BiasedRNG[118])|(((m[54]&m[65]&~m[182]))&~BiasedRNG[118])|((m[54]&m[65]&m[182]));
    m[104] = (((m[37]&~m[68]&m[148])|(~m[37]&m[68]&m[148]))&BiasedRNG[119])|(((m[37]&m[68]&~m[148]))&~BiasedRNG[119])|((m[37]&m[68]&m[148]));
    m[105] = (((m[43]&~m[69]&m[163])|(~m[43]&m[69]&m[163]))&BiasedRNG[120])|(((m[43]&m[69]&~m[163]))&~BiasedRNG[120])|((m[43]&m[69]&m[163]));
    m[106] = (((m[49]&~m[70]&m[183])|(~m[49]&m[70]&m[183]))&BiasedRNG[121])|(((m[49]&m[70]&~m[183]))&~BiasedRNG[121])|((m[49]&m[70]&m[183]));
    m[107] = (((m[55]&~m[71]&m[208])|(~m[55]&m[71]&m[208]))&BiasedRNG[122])|(((m[55]&m[71]&~m[208]))&~BiasedRNG[122])|((m[55]&m[71]&m[208]));
    m[108] = (((m[26]&~m[72]&m[143])|(~m[26]&m[72]&m[143]))&BiasedRNG[123])|(((m[26]&m[72]&~m[143]))&~BiasedRNG[123])|((m[26]&m[72]&m[143]));
    m[109] = (((m[32]&~m[73]&m[153])|(~m[32]&m[73]&m[153]))&BiasedRNG[124])|(((m[32]&m[73]&~m[153]))&~BiasedRNG[124])|((m[32]&m[73]&m[153]));
    m[114] = (((m[27]&~m[78]&m[158])|(~m[27]&m[78]&m[158]))&BiasedRNG[125])|(((m[27]&m[78]&~m[158]))&~BiasedRNG[125])|((m[27]&m[78]&m[158]));
    m[115] = (((m[33]&~m[79]&m[173])|(~m[33]&m[79]&m[173]))&BiasedRNG[126])|(((m[33]&m[79]&~m[173]))&~BiasedRNG[126])|((m[33]&m[79]&m[173]));
    m[120] = (((m[28]&~m[84]&m[178])|(~m[28]&m[84]&m[178]))&BiasedRNG[127])|(((m[28]&m[84]&~m[178]))&~BiasedRNG[127])|((m[28]&m[84]&m[178]));
    m[121] = (((m[34]&~m[85]&m[198])|(~m[34]&m[85]&m[198]))&BiasedRNG[128])|(((m[34]&m[85]&~m[198]))&~BiasedRNG[128])|((m[34]&m[85]&m[198]));
    m[126] = (((m[29]&~m[90]&m[203])|(~m[29]&m[90]&m[203]))&BiasedRNG[129])|(((m[29]&m[90]&~m[203]))&~BiasedRNG[129])|((m[29]&m[90]&m[203]));
    m[127] = (((m[35]&~m[91]&m[228])|(~m[35]&m[91]&m[228]))&BiasedRNG[130])|(((m[35]&m[91]&~m[228]))&~BiasedRNG[130])|((m[35]&m[91]&m[228]));
    m[133] = (((m[102]&~m[132]&~m[134]&~m[135]&~m[136])|(~m[102]&~m[132]&~m[134]&m[135]&~m[136])|(m[102]&m[132]&~m[134]&m[135]&~m[136])|(m[102]&~m[132]&m[134]&m[135]&~m[136])|(~m[102]&m[132]&~m[134]&~m[135]&m[136])|(~m[102]&~m[132]&m[134]&~m[135]&m[136])|(m[102]&m[132]&m[134]&~m[135]&m[136])|(~m[102]&m[132]&m[134]&m[135]&m[136]))&UnbiasedRNG[58])|((m[102]&~m[132]&~m[134]&m[135]&~m[136])|(~m[102]&~m[132]&~m[134]&~m[135]&m[136])|(m[102]&~m[132]&~m[134]&~m[135]&m[136])|(m[102]&m[132]&~m[134]&~m[135]&m[136])|(m[102]&~m[132]&m[134]&~m[135]&m[136])|(~m[102]&~m[132]&~m[134]&m[135]&m[136])|(m[102]&~m[132]&~m[134]&m[135]&m[136])|(~m[102]&m[132]&~m[134]&m[135]&m[136])|(m[102]&m[132]&~m[134]&m[135]&m[136])|(~m[102]&~m[132]&m[134]&m[135]&m[136])|(m[102]&~m[132]&m[134]&m[135]&m[136])|(m[102]&m[132]&m[134]&m[135]&m[136]));
    m[139] = (((m[136]&~m[137]&~m[138]&~m[140]&~m[141])|(~m[136]&~m[137]&~m[138]&m[140]&~m[141])|(m[136]&m[137]&~m[138]&m[140]&~m[141])|(m[136]&~m[137]&m[138]&m[140]&~m[141])|(~m[136]&m[137]&~m[138]&~m[140]&m[141])|(~m[136]&~m[137]&m[138]&~m[140]&m[141])|(m[136]&m[137]&m[138]&~m[140]&m[141])|(~m[136]&m[137]&m[138]&m[140]&m[141]))&UnbiasedRNG[59])|((m[136]&~m[137]&~m[138]&m[140]&~m[141])|(~m[136]&~m[137]&~m[138]&~m[140]&m[141])|(m[136]&~m[137]&~m[138]&~m[140]&m[141])|(m[136]&m[137]&~m[138]&~m[140]&m[141])|(m[136]&~m[137]&m[138]&~m[140]&m[141])|(~m[136]&~m[137]&~m[138]&m[140]&m[141])|(m[136]&~m[137]&~m[138]&m[140]&m[141])|(~m[136]&m[137]&~m[138]&m[140]&m[141])|(m[136]&m[137]&~m[138]&m[140]&m[141])|(~m[136]&~m[137]&m[138]&m[140]&m[141])|(m[136]&~m[137]&m[138]&m[140]&m[141])|(m[136]&m[137]&m[138]&m[140]&m[141]));
    m[149] = (((m[141]&~m[147]&~m[148]&~m[150]&~m[151])|(~m[141]&~m[147]&~m[148]&m[150]&~m[151])|(m[141]&m[147]&~m[148]&m[150]&~m[151])|(m[141]&~m[147]&m[148]&m[150]&~m[151])|(~m[141]&m[147]&~m[148]&~m[150]&m[151])|(~m[141]&~m[147]&m[148]&~m[150]&m[151])|(m[141]&m[147]&m[148]&~m[150]&m[151])|(~m[141]&m[147]&m[148]&m[150]&m[151]))&UnbiasedRNG[60])|((m[141]&~m[147]&~m[148]&m[150]&~m[151])|(~m[141]&~m[147]&~m[148]&~m[150]&m[151])|(m[141]&~m[147]&~m[148]&~m[150]&m[151])|(m[141]&m[147]&~m[148]&~m[150]&m[151])|(m[141]&~m[147]&m[148]&~m[150]&m[151])|(~m[141]&~m[147]&~m[148]&m[150]&m[151])|(m[141]&~m[147]&~m[148]&m[150]&m[151])|(~m[141]&m[147]&~m[148]&m[150]&m[151])|(m[141]&m[147]&~m[148]&m[150]&m[151])|(~m[141]&~m[147]&m[148]&m[150]&m[151])|(m[141]&~m[147]&m[148]&m[150]&m[151])|(m[141]&m[147]&m[148]&m[150]&m[151]));
    m[154] = (((m[146]&~m[152]&~m[153]&~m[155]&~m[156])|(~m[146]&~m[152]&~m[153]&m[155]&~m[156])|(m[146]&m[152]&~m[153]&m[155]&~m[156])|(m[146]&~m[152]&m[153]&m[155]&~m[156])|(~m[146]&m[152]&~m[153]&~m[155]&m[156])|(~m[146]&~m[152]&m[153]&~m[155]&m[156])|(m[146]&m[152]&m[153]&~m[155]&m[156])|(~m[146]&m[152]&m[153]&m[155]&m[156]))&UnbiasedRNG[61])|((m[146]&~m[152]&~m[153]&m[155]&~m[156])|(~m[146]&~m[152]&~m[153]&~m[155]&m[156])|(m[146]&~m[152]&~m[153]&~m[155]&m[156])|(m[146]&m[152]&~m[153]&~m[155]&m[156])|(m[146]&~m[152]&m[153]&~m[155]&m[156])|(~m[146]&~m[152]&~m[153]&m[155]&m[156])|(m[146]&~m[152]&~m[153]&m[155]&m[156])|(~m[146]&m[152]&~m[153]&m[155]&m[156])|(m[146]&m[152]&~m[153]&m[155]&m[156])|(~m[146]&~m[152]&m[153]&m[155]&m[156])|(m[146]&~m[152]&m[153]&m[155]&m[156])|(m[146]&m[152]&m[153]&m[155]&m[156]));
    m[164] = (((m[151]&~m[162]&~m[163]&~m[165]&~m[166])|(~m[151]&~m[162]&~m[163]&m[165]&~m[166])|(m[151]&m[162]&~m[163]&m[165]&~m[166])|(m[151]&~m[162]&m[163]&m[165]&~m[166])|(~m[151]&m[162]&~m[163]&~m[165]&m[166])|(~m[151]&~m[162]&m[163]&~m[165]&m[166])|(m[151]&m[162]&m[163]&~m[165]&m[166])|(~m[151]&m[162]&m[163]&m[165]&m[166]))&UnbiasedRNG[62])|((m[151]&~m[162]&~m[163]&m[165]&~m[166])|(~m[151]&~m[162]&~m[163]&~m[165]&m[166])|(m[151]&~m[162]&~m[163]&~m[165]&m[166])|(m[151]&m[162]&~m[163]&~m[165]&m[166])|(m[151]&~m[162]&m[163]&~m[165]&m[166])|(~m[151]&~m[162]&~m[163]&m[165]&m[166])|(m[151]&~m[162]&~m[163]&m[165]&m[166])|(~m[151]&m[162]&~m[163]&m[165]&m[166])|(m[151]&m[162]&~m[163]&m[165]&m[166])|(~m[151]&~m[162]&m[163]&m[165]&m[166])|(m[151]&~m[162]&m[163]&m[165]&m[166])|(m[151]&m[162]&m[163]&m[165]&m[166]));
    m[168] = (((m[110]&~m[167]&~m[169]&~m[170]&~m[171])|(~m[110]&~m[167]&~m[169]&m[170]&~m[171])|(m[110]&m[167]&~m[169]&m[170]&~m[171])|(m[110]&~m[167]&m[169]&m[170]&~m[171])|(~m[110]&m[167]&~m[169]&~m[170]&m[171])|(~m[110]&~m[167]&m[169]&~m[170]&m[171])|(m[110]&m[167]&m[169]&~m[170]&m[171])|(~m[110]&m[167]&m[169]&m[170]&m[171]))&UnbiasedRNG[63])|((m[110]&~m[167]&~m[169]&m[170]&~m[171])|(~m[110]&~m[167]&~m[169]&~m[170]&m[171])|(m[110]&~m[167]&~m[169]&~m[170]&m[171])|(m[110]&m[167]&~m[169]&~m[170]&m[171])|(m[110]&~m[167]&m[169]&~m[170]&m[171])|(~m[110]&~m[167]&~m[169]&m[170]&m[171])|(m[110]&~m[167]&~m[169]&m[170]&m[171])|(~m[110]&m[167]&~m[169]&m[170]&m[171])|(m[110]&m[167]&~m[169]&m[170]&m[171])|(~m[110]&~m[167]&m[169]&m[170]&m[171])|(m[110]&~m[167]&m[169]&m[170]&m[171])|(m[110]&m[167]&m[169]&m[170]&m[171]));
    m[174] = (((m[161]&~m[172]&~m[173]&~m[175]&~m[176])|(~m[161]&~m[172]&~m[173]&m[175]&~m[176])|(m[161]&m[172]&~m[173]&m[175]&~m[176])|(m[161]&~m[172]&m[173]&m[175]&~m[176])|(~m[161]&m[172]&~m[173]&~m[175]&m[176])|(~m[161]&~m[172]&m[173]&~m[175]&m[176])|(m[161]&m[172]&m[173]&~m[175]&m[176])|(~m[161]&m[172]&m[173]&m[175]&m[176]))&UnbiasedRNG[64])|((m[161]&~m[172]&~m[173]&m[175]&~m[176])|(~m[161]&~m[172]&~m[173]&~m[175]&m[176])|(m[161]&~m[172]&~m[173]&~m[175]&m[176])|(m[161]&m[172]&~m[173]&~m[175]&m[176])|(m[161]&~m[172]&m[173]&~m[175]&m[176])|(~m[161]&~m[172]&~m[173]&m[175]&m[176])|(m[161]&~m[172]&~m[173]&m[175]&m[176])|(~m[161]&m[172]&~m[173]&m[175]&m[176])|(m[161]&m[172]&~m[173]&m[175]&m[176])|(~m[161]&~m[172]&m[173]&m[175]&m[176])|(m[161]&~m[172]&m[173]&m[175]&m[176])|(m[161]&m[172]&m[173]&m[175]&m[176]));
    m[184] = (((m[166]&~m[182]&~m[183]&~m[185]&~m[186])|(~m[166]&~m[182]&~m[183]&m[185]&~m[186])|(m[166]&m[182]&~m[183]&m[185]&~m[186])|(m[166]&~m[182]&m[183]&m[185]&~m[186])|(~m[166]&m[182]&~m[183]&~m[185]&m[186])|(~m[166]&~m[182]&m[183]&~m[185]&m[186])|(m[166]&m[182]&m[183]&~m[185]&m[186])|(~m[166]&m[182]&m[183]&m[185]&m[186]))&UnbiasedRNG[65])|((m[166]&~m[182]&~m[183]&m[185]&~m[186])|(~m[166]&~m[182]&~m[183]&~m[185]&m[186])|(m[166]&~m[182]&~m[183]&~m[185]&m[186])|(m[166]&m[182]&~m[183]&~m[185]&m[186])|(m[166]&~m[182]&m[183]&~m[185]&m[186])|(~m[166]&~m[182]&~m[183]&m[185]&m[186])|(m[166]&~m[182]&~m[183]&m[185]&m[186])|(~m[166]&m[182]&~m[183]&m[185]&m[186])|(m[166]&m[182]&~m[183]&m[185]&m[186])|(~m[166]&~m[182]&m[183]&m[185]&m[186])|(m[166]&~m[182]&m[183]&m[185]&m[186])|(m[166]&m[182]&m[183]&m[185]&m[186]));
    m[188] = (((m[111]&~m[187]&~m[189]&~m[190]&~m[191])|(~m[111]&~m[187]&~m[189]&m[190]&~m[191])|(m[111]&m[187]&~m[189]&m[190]&~m[191])|(m[111]&~m[187]&m[189]&m[190]&~m[191])|(~m[111]&m[187]&~m[189]&~m[190]&m[191])|(~m[111]&~m[187]&m[189]&~m[190]&m[191])|(m[111]&m[187]&m[189]&~m[190]&m[191])|(~m[111]&m[187]&m[189]&m[190]&m[191]))&UnbiasedRNG[66])|((m[111]&~m[187]&~m[189]&m[190]&~m[191])|(~m[111]&~m[187]&~m[189]&~m[190]&m[191])|(m[111]&~m[187]&~m[189]&~m[190]&m[191])|(m[111]&m[187]&~m[189]&~m[190]&m[191])|(m[111]&~m[187]&m[189]&~m[190]&m[191])|(~m[111]&~m[187]&~m[189]&m[190]&m[191])|(m[111]&~m[187]&~m[189]&m[190]&m[191])|(~m[111]&m[187]&~m[189]&m[190]&m[191])|(m[111]&m[187]&~m[189]&m[190]&m[191])|(~m[111]&~m[187]&m[189]&m[190]&m[191])|(m[111]&~m[187]&m[189]&m[190]&m[191])|(m[111]&m[187]&m[189]&m[190]&m[191]));
    m[193] = (((m[116]&~m[192]&~m[194]&~m[195]&~m[196])|(~m[116]&~m[192]&~m[194]&m[195]&~m[196])|(m[116]&m[192]&~m[194]&m[195]&~m[196])|(m[116]&~m[192]&m[194]&m[195]&~m[196])|(~m[116]&m[192]&~m[194]&~m[195]&m[196])|(~m[116]&~m[192]&m[194]&~m[195]&m[196])|(m[116]&m[192]&m[194]&~m[195]&m[196])|(~m[116]&m[192]&m[194]&m[195]&m[196]))&UnbiasedRNG[67])|((m[116]&~m[192]&~m[194]&m[195]&~m[196])|(~m[116]&~m[192]&~m[194]&~m[195]&m[196])|(m[116]&~m[192]&~m[194]&~m[195]&m[196])|(m[116]&m[192]&~m[194]&~m[195]&m[196])|(m[116]&~m[192]&m[194]&~m[195]&m[196])|(~m[116]&~m[192]&~m[194]&m[195]&m[196])|(m[116]&~m[192]&~m[194]&m[195]&m[196])|(~m[116]&m[192]&~m[194]&m[195]&m[196])|(m[116]&m[192]&~m[194]&m[195]&m[196])|(~m[116]&~m[192]&m[194]&m[195]&m[196])|(m[116]&~m[192]&m[194]&m[195]&m[196])|(m[116]&m[192]&m[194]&m[195]&m[196]));
    m[199] = (((m[181]&~m[197]&~m[198]&~m[200]&~m[201])|(~m[181]&~m[197]&~m[198]&m[200]&~m[201])|(m[181]&m[197]&~m[198]&m[200]&~m[201])|(m[181]&~m[197]&m[198]&m[200]&~m[201])|(~m[181]&m[197]&~m[198]&~m[200]&m[201])|(~m[181]&~m[197]&m[198]&~m[200]&m[201])|(m[181]&m[197]&m[198]&~m[200]&m[201])|(~m[181]&m[197]&m[198]&m[200]&m[201]))&UnbiasedRNG[68])|((m[181]&~m[197]&~m[198]&m[200]&~m[201])|(~m[181]&~m[197]&~m[198]&~m[200]&m[201])|(m[181]&~m[197]&~m[198]&~m[200]&m[201])|(m[181]&m[197]&~m[198]&~m[200]&m[201])|(m[181]&~m[197]&m[198]&~m[200]&m[201])|(~m[181]&~m[197]&~m[198]&m[200]&m[201])|(m[181]&~m[197]&~m[198]&m[200]&m[201])|(~m[181]&m[197]&~m[198]&m[200]&m[201])|(m[181]&m[197]&~m[198]&m[200]&m[201])|(~m[181]&~m[197]&m[198]&m[200]&m[201])|(m[181]&~m[197]&m[198]&m[200]&m[201])|(m[181]&m[197]&m[198]&m[200]&m[201]));
    m[209] = (((m[186]&~m[207]&~m[208]&~m[210]&~m[211])|(~m[186]&~m[207]&~m[208]&m[210]&~m[211])|(m[186]&m[207]&~m[208]&m[210]&~m[211])|(m[186]&~m[207]&m[208]&m[210]&~m[211])|(~m[186]&m[207]&~m[208]&~m[210]&m[211])|(~m[186]&~m[207]&m[208]&~m[210]&m[211])|(m[186]&m[207]&m[208]&~m[210]&m[211])|(~m[186]&m[207]&m[208]&m[210]&m[211]))&UnbiasedRNG[69])|((m[186]&~m[207]&~m[208]&m[210]&~m[211])|(~m[186]&~m[207]&~m[208]&~m[210]&m[211])|(m[186]&~m[207]&~m[208]&~m[210]&m[211])|(m[186]&m[207]&~m[208]&~m[210]&m[211])|(m[186]&~m[207]&m[208]&~m[210]&m[211])|(~m[186]&~m[207]&~m[208]&m[210]&m[211])|(m[186]&~m[207]&~m[208]&m[210]&m[211])|(~m[186]&m[207]&~m[208]&m[210]&m[211])|(m[186]&m[207]&~m[208]&m[210]&m[211])|(~m[186]&~m[207]&m[208]&m[210]&m[211])|(m[186]&~m[207]&m[208]&m[210]&m[211])|(m[186]&m[207]&m[208]&m[210]&m[211]));
    m[213] = (((m[112]&~m[212]&~m[214]&~m[215]&~m[216])|(~m[112]&~m[212]&~m[214]&m[215]&~m[216])|(m[112]&m[212]&~m[214]&m[215]&~m[216])|(m[112]&~m[212]&m[214]&m[215]&~m[216])|(~m[112]&m[212]&~m[214]&~m[215]&m[216])|(~m[112]&~m[212]&m[214]&~m[215]&m[216])|(m[112]&m[212]&m[214]&~m[215]&m[216])|(~m[112]&m[212]&m[214]&m[215]&m[216]))&UnbiasedRNG[70])|((m[112]&~m[212]&~m[214]&m[215]&~m[216])|(~m[112]&~m[212]&~m[214]&~m[215]&m[216])|(m[112]&~m[212]&~m[214]&~m[215]&m[216])|(m[112]&m[212]&~m[214]&~m[215]&m[216])|(m[112]&~m[212]&m[214]&~m[215]&m[216])|(~m[112]&~m[212]&~m[214]&m[215]&m[216])|(m[112]&~m[212]&~m[214]&m[215]&m[216])|(~m[112]&m[212]&~m[214]&m[215]&m[216])|(m[112]&m[212]&~m[214]&m[215]&m[216])|(~m[112]&~m[212]&m[214]&m[215]&m[216])|(m[112]&~m[212]&m[214]&m[215]&m[216])|(m[112]&m[212]&m[214]&m[215]&m[216]));
    m[218] = (((m[117]&~m[217]&~m[219]&~m[220]&~m[221])|(~m[117]&~m[217]&~m[219]&m[220]&~m[221])|(m[117]&m[217]&~m[219]&m[220]&~m[221])|(m[117]&~m[217]&m[219]&m[220]&~m[221])|(~m[117]&m[217]&~m[219]&~m[220]&m[221])|(~m[117]&~m[217]&m[219]&~m[220]&m[221])|(m[117]&m[217]&m[219]&~m[220]&m[221])|(~m[117]&m[217]&m[219]&m[220]&m[221]))&UnbiasedRNG[71])|((m[117]&~m[217]&~m[219]&m[220]&~m[221])|(~m[117]&~m[217]&~m[219]&~m[220]&m[221])|(m[117]&~m[217]&~m[219]&~m[220]&m[221])|(m[117]&m[217]&~m[219]&~m[220]&m[221])|(m[117]&~m[217]&m[219]&~m[220]&m[221])|(~m[117]&~m[217]&~m[219]&m[220]&m[221])|(m[117]&~m[217]&~m[219]&m[220]&m[221])|(~m[117]&m[217]&~m[219]&m[220]&m[221])|(m[117]&m[217]&~m[219]&m[220]&m[221])|(~m[117]&~m[217]&m[219]&m[220]&m[221])|(m[117]&~m[217]&m[219]&m[220]&m[221])|(m[117]&m[217]&m[219]&m[220]&m[221]));
    m[223] = (((m[122]&~m[222]&~m[224]&~m[225]&~m[226])|(~m[122]&~m[222]&~m[224]&m[225]&~m[226])|(m[122]&m[222]&~m[224]&m[225]&~m[226])|(m[122]&~m[222]&m[224]&m[225]&~m[226])|(~m[122]&m[222]&~m[224]&~m[225]&m[226])|(~m[122]&~m[222]&m[224]&~m[225]&m[226])|(m[122]&m[222]&m[224]&~m[225]&m[226])|(~m[122]&m[222]&m[224]&m[225]&m[226]))&UnbiasedRNG[72])|((m[122]&~m[222]&~m[224]&m[225]&~m[226])|(~m[122]&~m[222]&~m[224]&~m[225]&m[226])|(m[122]&~m[222]&~m[224]&~m[225]&m[226])|(m[122]&m[222]&~m[224]&~m[225]&m[226])|(m[122]&~m[222]&m[224]&~m[225]&m[226])|(~m[122]&~m[222]&~m[224]&m[225]&m[226])|(m[122]&~m[222]&~m[224]&m[225]&m[226])|(~m[122]&m[222]&~m[224]&m[225]&m[226])|(m[122]&m[222]&~m[224]&m[225]&m[226])|(~m[122]&~m[222]&m[224]&m[225]&m[226])|(m[122]&~m[222]&m[224]&m[225]&m[226])|(m[122]&m[222]&m[224]&m[225]&m[226]));
    m[229] = (((m[206]&~m[227]&~m[228]&~m[230]&~m[231])|(~m[206]&~m[227]&~m[228]&m[230]&~m[231])|(m[206]&m[227]&~m[228]&m[230]&~m[231])|(m[206]&~m[227]&m[228]&m[230]&~m[231])|(~m[206]&m[227]&~m[228]&~m[230]&m[231])|(~m[206]&~m[227]&m[228]&~m[230]&m[231])|(m[206]&m[227]&m[228]&~m[230]&m[231])|(~m[206]&m[227]&m[228]&m[230]&m[231]))&UnbiasedRNG[73])|((m[206]&~m[227]&~m[228]&m[230]&~m[231])|(~m[206]&~m[227]&~m[228]&~m[230]&m[231])|(m[206]&~m[227]&~m[228]&~m[230]&m[231])|(m[206]&m[227]&~m[228]&~m[230]&m[231])|(m[206]&~m[227]&m[228]&~m[230]&m[231])|(~m[206]&~m[227]&~m[228]&m[230]&m[231])|(m[206]&~m[227]&~m[228]&m[230]&m[231])|(~m[206]&m[227]&~m[228]&m[230]&m[231])|(m[206]&m[227]&~m[228]&m[230]&m[231])|(~m[206]&~m[227]&m[228]&m[230]&m[231])|(m[206]&~m[227]&m[228]&m[230]&m[231])|(m[206]&m[227]&m[228]&m[230]&m[231]));
    m[233] = (((m[113]&~m[232]&~m[234]&~m[235]&~m[236])|(~m[113]&~m[232]&~m[234]&m[235]&~m[236])|(m[113]&m[232]&~m[234]&m[235]&~m[236])|(m[113]&~m[232]&m[234]&m[235]&~m[236])|(~m[113]&m[232]&~m[234]&~m[235]&m[236])|(~m[113]&~m[232]&m[234]&~m[235]&m[236])|(m[113]&m[232]&m[234]&~m[235]&m[236])|(~m[113]&m[232]&m[234]&m[235]&m[236]))&UnbiasedRNG[74])|((m[113]&~m[232]&~m[234]&m[235]&~m[236])|(~m[113]&~m[232]&~m[234]&~m[235]&m[236])|(m[113]&~m[232]&~m[234]&~m[235]&m[236])|(m[113]&m[232]&~m[234]&~m[235]&m[236])|(m[113]&~m[232]&m[234]&~m[235]&m[236])|(~m[113]&~m[232]&~m[234]&m[235]&m[236])|(m[113]&~m[232]&~m[234]&m[235]&m[236])|(~m[113]&m[232]&~m[234]&m[235]&m[236])|(m[113]&m[232]&~m[234]&m[235]&m[236])|(~m[113]&~m[232]&m[234]&m[235]&m[236])|(m[113]&~m[232]&m[234]&m[235]&m[236])|(m[113]&m[232]&m[234]&m[235]&m[236]));
    m[238] = (((m[118]&~m[237]&~m[239]&~m[240]&~m[241])|(~m[118]&~m[237]&~m[239]&m[240]&~m[241])|(m[118]&m[237]&~m[239]&m[240]&~m[241])|(m[118]&~m[237]&m[239]&m[240]&~m[241])|(~m[118]&m[237]&~m[239]&~m[240]&m[241])|(~m[118]&~m[237]&m[239]&~m[240]&m[241])|(m[118]&m[237]&m[239]&~m[240]&m[241])|(~m[118]&m[237]&m[239]&m[240]&m[241]))&UnbiasedRNG[75])|((m[118]&~m[237]&~m[239]&m[240]&~m[241])|(~m[118]&~m[237]&~m[239]&~m[240]&m[241])|(m[118]&~m[237]&~m[239]&~m[240]&m[241])|(m[118]&m[237]&~m[239]&~m[240]&m[241])|(m[118]&~m[237]&m[239]&~m[240]&m[241])|(~m[118]&~m[237]&~m[239]&m[240]&m[241])|(m[118]&~m[237]&~m[239]&m[240]&m[241])|(~m[118]&m[237]&~m[239]&m[240]&m[241])|(m[118]&m[237]&~m[239]&m[240]&m[241])|(~m[118]&~m[237]&m[239]&m[240]&m[241])|(m[118]&~m[237]&m[239]&m[240]&m[241])|(m[118]&m[237]&m[239]&m[240]&m[241]));
    m[243] = (((m[123]&~m[242]&~m[244]&~m[245]&~m[246])|(~m[123]&~m[242]&~m[244]&m[245]&~m[246])|(m[123]&m[242]&~m[244]&m[245]&~m[246])|(m[123]&~m[242]&m[244]&m[245]&~m[246])|(~m[123]&m[242]&~m[244]&~m[245]&m[246])|(~m[123]&~m[242]&m[244]&~m[245]&m[246])|(m[123]&m[242]&m[244]&~m[245]&m[246])|(~m[123]&m[242]&m[244]&m[245]&m[246]))&UnbiasedRNG[76])|((m[123]&~m[242]&~m[244]&m[245]&~m[246])|(~m[123]&~m[242]&~m[244]&~m[245]&m[246])|(m[123]&~m[242]&~m[244]&~m[245]&m[246])|(m[123]&m[242]&~m[244]&~m[245]&m[246])|(m[123]&~m[242]&m[244]&~m[245]&m[246])|(~m[123]&~m[242]&~m[244]&m[245]&m[246])|(m[123]&~m[242]&~m[244]&m[245]&m[246])|(~m[123]&m[242]&~m[244]&m[245]&m[246])|(m[123]&m[242]&~m[244]&m[245]&m[246])|(~m[123]&~m[242]&m[244]&m[245]&m[246])|(m[123]&~m[242]&m[244]&m[245]&m[246])|(m[123]&m[242]&m[244]&m[245]&m[246]));
    m[248] = (((m[128]&~m[247]&~m[249]&~m[250]&~m[251])|(~m[128]&~m[247]&~m[249]&m[250]&~m[251])|(m[128]&m[247]&~m[249]&m[250]&~m[251])|(m[128]&~m[247]&m[249]&m[250]&~m[251])|(~m[128]&m[247]&~m[249]&~m[250]&m[251])|(~m[128]&~m[247]&m[249]&~m[250]&m[251])|(m[128]&m[247]&m[249]&~m[250]&m[251])|(~m[128]&m[247]&m[249]&m[250]&m[251]))&UnbiasedRNG[77])|((m[128]&~m[247]&~m[249]&m[250]&~m[251])|(~m[128]&~m[247]&~m[249]&~m[250]&m[251])|(m[128]&~m[247]&~m[249]&~m[250]&m[251])|(m[128]&m[247]&~m[249]&~m[250]&m[251])|(m[128]&~m[247]&m[249]&~m[250]&m[251])|(~m[128]&~m[247]&~m[249]&m[250]&m[251])|(m[128]&~m[247]&~m[249]&m[250]&m[251])|(~m[128]&m[247]&~m[249]&m[250]&m[251])|(m[128]&m[247]&~m[249]&m[250]&m[251])|(~m[128]&~m[247]&m[249]&m[250]&m[251])|(m[128]&~m[247]&m[249]&m[250]&m[251])|(m[128]&m[247]&m[249]&m[250]&m[251]));
    m[253] = (((m[119]&~m[252]&~m[254]&~m[255]&~m[256])|(~m[119]&~m[252]&~m[254]&m[255]&~m[256])|(m[119]&m[252]&~m[254]&m[255]&~m[256])|(m[119]&~m[252]&m[254]&m[255]&~m[256])|(~m[119]&m[252]&~m[254]&~m[255]&m[256])|(~m[119]&~m[252]&m[254]&~m[255]&m[256])|(m[119]&m[252]&m[254]&~m[255]&m[256])|(~m[119]&m[252]&m[254]&m[255]&m[256]))&UnbiasedRNG[78])|((m[119]&~m[252]&~m[254]&m[255]&~m[256])|(~m[119]&~m[252]&~m[254]&~m[255]&m[256])|(m[119]&~m[252]&~m[254]&~m[255]&m[256])|(m[119]&m[252]&~m[254]&~m[255]&m[256])|(m[119]&~m[252]&m[254]&~m[255]&m[256])|(~m[119]&~m[252]&~m[254]&m[255]&m[256])|(m[119]&~m[252]&~m[254]&m[255]&m[256])|(~m[119]&m[252]&~m[254]&m[255]&m[256])|(m[119]&m[252]&~m[254]&m[255]&m[256])|(~m[119]&~m[252]&m[254]&m[255]&m[256])|(m[119]&~m[252]&m[254]&m[255]&m[256])|(m[119]&m[252]&m[254]&m[255]&m[256]));
    m[258] = (((m[124]&~m[257]&~m[259]&~m[260]&~m[261])|(~m[124]&~m[257]&~m[259]&m[260]&~m[261])|(m[124]&m[257]&~m[259]&m[260]&~m[261])|(m[124]&~m[257]&m[259]&m[260]&~m[261])|(~m[124]&m[257]&~m[259]&~m[260]&m[261])|(~m[124]&~m[257]&m[259]&~m[260]&m[261])|(m[124]&m[257]&m[259]&~m[260]&m[261])|(~m[124]&m[257]&m[259]&m[260]&m[261]))&UnbiasedRNG[79])|((m[124]&~m[257]&~m[259]&m[260]&~m[261])|(~m[124]&~m[257]&~m[259]&~m[260]&m[261])|(m[124]&~m[257]&~m[259]&~m[260]&m[261])|(m[124]&m[257]&~m[259]&~m[260]&m[261])|(m[124]&~m[257]&m[259]&~m[260]&m[261])|(~m[124]&~m[257]&~m[259]&m[260]&m[261])|(m[124]&~m[257]&~m[259]&m[260]&m[261])|(~m[124]&m[257]&~m[259]&m[260]&m[261])|(m[124]&m[257]&~m[259]&m[260]&m[261])|(~m[124]&~m[257]&m[259]&m[260]&m[261])|(m[124]&~m[257]&m[259]&m[260]&m[261])|(m[124]&m[257]&m[259]&m[260]&m[261]));
    m[263] = (((m[129]&~m[262]&~m[264]&~m[265]&~m[266])|(~m[129]&~m[262]&~m[264]&m[265]&~m[266])|(m[129]&m[262]&~m[264]&m[265]&~m[266])|(m[129]&~m[262]&m[264]&m[265]&~m[266])|(~m[129]&m[262]&~m[264]&~m[265]&m[266])|(~m[129]&~m[262]&m[264]&~m[265]&m[266])|(m[129]&m[262]&m[264]&~m[265]&m[266])|(~m[129]&m[262]&m[264]&m[265]&m[266]))&UnbiasedRNG[80])|((m[129]&~m[262]&~m[264]&m[265]&~m[266])|(~m[129]&~m[262]&~m[264]&~m[265]&m[266])|(m[129]&~m[262]&~m[264]&~m[265]&m[266])|(m[129]&m[262]&~m[264]&~m[265]&m[266])|(m[129]&~m[262]&m[264]&~m[265]&m[266])|(~m[129]&~m[262]&~m[264]&m[265]&m[266])|(m[129]&~m[262]&~m[264]&m[265]&m[266])|(~m[129]&m[262]&~m[264]&m[265]&m[266])|(m[129]&m[262]&~m[264]&m[265]&m[266])|(~m[129]&~m[262]&m[264]&m[265]&m[266])|(m[129]&~m[262]&m[264]&m[265]&m[266])|(m[129]&m[262]&m[264]&m[265]&m[266]));
    m[268] = (((m[125]&~m[267]&~m[269]&~m[270]&~m[271])|(~m[125]&~m[267]&~m[269]&m[270]&~m[271])|(m[125]&m[267]&~m[269]&m[270]&~m[271])|(m[125]&~m[267]&m[269]&m[270]&~m[271])|(~m[125]&m[267]&~m[269]&~m[270]&m[271])|(~m[125]&~m[267]&m[269]&~m[270]&m[271])|(m[125]&m[267]&m[269]&~m[270]&m[271])|(~m[125]&m[267]&m[269]&m[270]&m[271]))&UnbiasedRNG[81])|((m[125]&~m[267]&~m[269]&m[270]&~m[271])|(~m[125]&~m[267]&~m[269]&~m[270]&m[271])|(m[125]&~m[267]&~m[269]&~m[270]&m[271])|(m[125]&m[267]&~m[269]&~m[270]&m[271])|(m[125]&~m[267]&m[269]&~m[270]&m[271])|(~m[125]&~m[267]&~m[269]&m[270]&m[271])|(m[125]&~m[267]&~m[269]&m[270]&m[271])|(~m[125]&m[267]&~m[269]&m[270]&m[271])|(m[125]&m[267]&~m[269]&m[270]&m[271])|(~m[125]&~m[267]&m[269]&m[270]&m[271])|(m[125]&~m[267]&m[269]&m[270]&m[271])|(m[125]&m[267]&m[269]&m[270]&m[271]));
    m[273] = (((m[130]&~m[272]&~m[274]&~m[275]&~m[276])|(~m[130]&~m[272]&~m[274]&m[275]&~m[276])|(m[130]&m[272]&~m[274]&m[275]&~m[276])|(m[130]&~m[272]&m[274]&m[275]&~m[276])|(~m[130]&m[272]&~m[274]&~m[275]&m[276])|(~m[130]&~m[272]&m[274]&~m[275]&m[276])|(m[130]&m[272]&m[274]&~m[275]&m[276])|(~m[130]&m[272]&m[274]&m[275]&m[276]))&UnbiasedRNG[82])|((m[130]&~m[272]&~m[274]&m[275]&~m[276])|(~m[130]&~m[272]&~m[274]&~m[275]&m[276])|(m[130]&~m[272]&~m[274]&~m[275]&m[276])|(m[130]&m[272]&~m[274]&~m[275]&m[276])|(m[130]&~m[272]&m[274]&~m[275]&m[276])|(~m[130]&~m[272]&~m[274]&m[275]&m[276])|(m[130]&~m[272]&~m[274]&m[275]&m[276])|(~m[130]&m[272]&~m[274]&m[275]&m[276])|(m[130]&m[272]&~m[274]&m[275]&m[276])|(~m[130]&~m[272]&m[274]&m[275]&m[276])|(m[130]&~m[272]&m[274]&m[275]&m[276])|(m[130]&m[272]&m[274]&m[275]&m[276]));
    m[278] = (((m[131]&~m[277]&~m[279]&~m[280]&~m[281])|(~m[131]&~m[277]&~m[279]&m[280]&~m[281])|(m[131]&m[277]&~m[279]&m[280]&~m[281])|(m[131]&~m[277]&m[279]&m[280]&~m[281])|(~m[131]&m[277]&~m[279]&~m[280]&m[281])|(~m[131]&~m[277]&m[279]&~m[280]&m[281])|(m[131]&m[277]&m[279]&~m[280]&m[281])|(~m[131]&m[277]&m[279]&m[280]&m[281]))&UnbiasedRNG[83])|((m[131]&~m[277]&~m[279]&m[280]&~m[281])|(~m[131]&~m[277]&~m[279]&~m[280]&m[281])|(m[131]&~m[277]&~m[279]&~m[280]&m[281])|(m[131]&m[277]&~m[279]&~m[280]&m[281])|(m[131]&~m[277]&m[279]&~m[280]&m[281])|(~m[131]&~m[277]&~m[279]&m[280]&m[281])|(m[131]&~m[277]&~m[279]&m[280]&m[281])|(~m[131]&m[277]&~m[279]&m[280]&m[281])|(m[131]&m[277]&~m[279]&m[280]&m[281])|(~m[131]&~m[277]&m[279]&m[280]&m[281])|(m[131]&~m[277]&m[279]&m[280]&m[281])|(m[131]&m[277]&m[279]&m[280]&m[281]));
end

always @(posedge color3_clk) begin
    m[140] = (((m[137]&~m[138]&~m[139]&~m[141]&~m[142])|(~m[137]&m[138]&~m[139]&~m[141]&~m[142])|(~m[137]&~m[138]&m[139]&~m[141]&~m[142])|(m[137]&m[138]&m[139]&m[141]&~m[142])|(~m[137]&~m[138]&~m[139]&~m[141]&m[142])|(m[137]&m[138]&~m[139]&m[141]&m[142])|(m[137]&~m[138]&m[139]&m[141]&m[142])|(~m[137]&m[138]&m[139]&m[141]&m[142]))&UnbiasedRNG[84])|((m[137]&m[138]&~m[139]&~m[141]&~m[142])|(m[137]&~m[138]&m[139]&~m[141]&~m[142])|(~m[137]&m[138]&m[139]&~m[141]&~m[142])|(m[137]&m[138]&m[139]&~m[141]&~m[142])|(m[137]&~m[138]&~m[139]&~m[141]&m[142])|(~m[137]&m[138]&~m[139]&~m[141]&m[142])|(m[137]&m[138]&~m[139]&~m[141]&m[142])|(~m[137]&~m[138]&m[139]&~m[141]&m[142])|(m[137]&~m[138]&m[139]&~m[141]&m[142])|(~m[137]&m[138]&m[139]&~m[141]&m[142])|(m[137]&m[138]&m[139]&~m[141]&m[142])|(m[137]&m[138]&m[139]&m[141]&m[142]));
    m[150] = (((m[147]&~m[148]&~m[149]&~m[151]&~m[152])|(~m[147]&m[148]&~m[149]&~m[151]&~m[152])|(~m[147]&~m[148]&m[149]&~m[151]&~m[152])|(m[147]&m[148]&m[149]&m[151]&~m[152])|(~m[147]&~m[148]&~m[149]&~m[151]&m[152])|(m[147]&m[148]&~m[149]&m[151]&m[152])|(m[147]&~m[148]&m[149]&m[151]&m[152])|(~m[147]&m[148]&m[149]&m[151]&m[152]))&UnbiasedRNG[85])|((m[147]&m[148]&~m[149]&~m[151]&~m[152])|(m[147]&~m[148]&m[149]&~m[151]&~m[152])|(~m[147]&m[148]&m[149]&~m[151]&~m[152])|(m[147]&m[148]&m[149]&~m[151]&~m[152])|(m[147]&~m[148]&~m[149]&~m[151]&m[152])|(~m[147]&m[148]&~m[149]&~m[151]&m[152])|(m[147]&m[148]&~m[149]&~m[151]&m[152])|(~m[147]&~m[148]&m[149]&~m[151]&m[152])|(m[147]&~m[148]&m[149]&~m[151]&m[152])|(~m[147]&m[148]&m[149]&~m[151]&m[152])|(m[147]&m[148]&m[149]&~m[151]&m[152])|(m[147]&m[148]&m[149]&m[151]&m[152]));
    m[155] = (((m[152]&~m[153]&~m[154]&~m[156]&~m[157])|(~m[152]&m[153]&~m[154]&~m[156]&~m[157])|(~m[152]&~m[153]&m[154]&~m[156]&~m[157])|(m[152]&m[153]&m[154]&m[156]&~m[157])|(~m[152]&~m[153]&~m[154]&~m[156]&m[157])|(m[152]&m[153]&~m[154]&m[156]&m[157])|(m[152]&~m[153]&m[154]&m[156]&m[157])|(~m[152]&m[153]&m[154]&m[156]&m[157]))&UnbiasedRNG[86])|((m[152]&m[153]&~m[154]&~m[156]&~m[157])|(m[152]&~m[153]&m[154]&~m[156]&~m[157])|(~m[152]&m[153]&m[154]&~m[156]&~m[157])|(m[152]&m[153]&m[154]&~m[156]&~m[157])|(m[152]&~m[153]&~m[154]&~m[156]&m[157])|(~m[152]&m[153]&~m[154]&~m[156]&m[157])|(m[152]&m[153]&~m[154]&~m[156]&m[157])|(~m[152]&~m[153]&m[154]&~m[156]&m[157])|(m[152]&~m[153]&m[154]&~m[156]&m[157])|(~m[152]&m[153]&m[154]&~m[156]&m[157])|(m[152]&m[153]&m[154]&~m[156]&m[157])|(m[152]&m[153]&m[154]&m[156]&m[157]));
    m[165] = (((m[162]&~m[163]&~m[164]&~m[166]&~m[167])|(~m[162]&m[163]&~m[164]&~m[166]&~m[167])|(~m[162]&~m[163]&m[164]&~m[166]&~m[167])|(m[162]&m[163]&m[164]&m[166]&~m[167])|(~m[162]&~m[163]&~m[164]&~m[166]&m[167])|(m[162]&m[163]&~m[164]&m[166]&m[167])|(m[162]&~m[163]&m[164]&m[166]&m[167])|(~m[162]&m[163]&m[164]&m[166]&m[167]))&UnbiasedRNG[87])|((m[162]&m[163]&~m[164]&~m[166]&~m[167])|(m[162]&~m[163]&m[164]&~m[166]&~m[167])|(~m[162]&m[163]&m[164]&~m[166]&~m[167])|(m[162]&m[163]&m[164]&~m[166]&~m[167])|(m[162]&~m[163]&~m[164]&~m[166]&m[167])|(~m[162]&m[163]&~m[164]&~m[166]&m[167])|(m[162]&m[163]&~m[164]&~m[166]&m[167])|(~m[162]&~m[163]&m[164]&~m[166]&m[167])|(m[162]&~m[163]&m[164]&~m[166]&m[167])|(~m[162]&m[163]&m[164]&~m[166]&m[167])|(m[162]&m[163]&m[164]&~m[166]&m[167])|(m[162]&m[163]&m[164]&m[166]&m[167]));
    m[170] = (((m[167]&~m[168]&~m[169]&~m[171]&~m[172])|(~m[167]&m[168]&~m[169]&~m[171]&~m[172])|(~m[167]&~m[168]&m[169]&~m[171]&~m[172])|(m[167]&m[168]&m[169]&m[171]&~m[172])|(~m[167]&~m[168]&~m[169]&~m[171]&m[172])|(m[167]&m[168]&~m[169]&m[171]&m[172])|(m[167]&~m[168]&m[169]&m[171]&m[172])|(~m[167]&m[168]&m[169]&m[171]&m[172]))&UnbiasedRNG[88])|((m[167]&m[168]&~m[169]&~m[171]&~m[172])|(m[167]&~m[168]&m[169]&~m[171]&~m[172])|(~m[167]&m[168]&m[169]&~m[171]&~m[172])|(m[167]&m[168]&m[169]&~m[171]&~m[172])|(m[167]&~m[168]&~m[169]&~m[171]&m[172])|(~m[167]&m[168]&~m[169]&~m[171]&m[172])|(m[167]&m[168]&~m[169]&~m[171]&m[172])|(~m[167]&~m[168]&m[169]&~m[171]&m[172])|(m[167]&~m[168]&m[169]&~m[171]&m[172])|(~m[167]&m[168]&m[169]&~m[171]&m[172])|(m[167]&m[168]&m[169]&~m[171]&m[172])|(m[167]&m[168]&m[169]&m[171]&m[172]));
    m[175] = (((m[172]&~m[173]&~m[174]&~m[176]&~m[177])|(~m[172]&m[173]&~m[174]&~m[176]&~m[177])|(~m[172]&~m[173]&m[174]&~m[176]&~m[177])|(m[172]&m[173]&m[174]&m[176]&~m[177])|(~m[172]&~m[173]&~m[174]&~m[176]&m[177])|(m[172]&m[173]&~m[174]&m[176]&m[177])|(m[172]&~m[173]&m[174]&m[176]&m[177])|(~m[172]&m[173]&m[174]&m[176]&m[177]))&UnbiasedRNG[89])|((m[172]&m[173]&~m[174]&~m[176]&~m[177])|(m[172]&~m[173]&m[174]&~m[176]&~m[177])|(~m[172]&m[173]&m[174]&~m[176]&~m[177])|(m[172]&m[173]&m[174]&~m[176]&~m[177])|(m[172]&~m[173]&~m[174]&~m[176]&m[177])|(~m[172]&m[173]&~m[174]&~m[176]&m[177])|(m[172]&m[173]&~m[174]&~m[176]&m[177])|(~m[172]&~m[173]&m[174]&~m[176]&m[177])|(m[172]&~m[173]&m[174]&~m[176]&m[177])|(~m[172]&m[173]&m[174]&~m[176]&m[177])|(m[172]&m[173]&m[174]&~m[176]&m[177])|(m[172]&m[173]&m[174]&m[176]&m[177]));
    m[185] = (((m[182]&~m[183]&~m[184]&~m[186]&~m[187])|(~m[182]&m[183]&~m[184]&~m[186]&~m[187])|(~m[182]&~m[183]&m[184]&~m[186]&~m[187])|(m[182]&m[183]&m[184]&m[186]&~m[187])|(~m[182]&~m[183]&~m[184]&~m[186]&m[187])|(m[182]&m[183]&~m[184]&m[186]&m[187])|(m[182]&~m[183]&m[184]&m[186]&m[187])|(~m[182]&m[183]&m[184]&m[186]&m[187]))&UnbiasedRNG[90])|((m[182]&m[183]&~m[184]&~m[186]&~m[187])|(m[182]&~m[183]&m[184]&~m[186]&~m[187])|(~m[182]&m[183]&m[184]&~m[186]&~m[187])|(m[182]&m[183]&m[184]&~m[186]&~m[187])|(m[182]&~m[183]&~m[184]&~m[186]&m[187])|(~m[182]&m[183]&~m[184]&~m[186]&m[187])|(m[182]&m[183]&~m[184]&~m[186]&m[187])|(~m[182]&~m[183]&m[184]&~m[186]&m[187])|(m[182]&~m[183]&m[184]&~m[186]&m[187])|(~m[182]&m[183]&m[184]&~m[186]&m[187])|(m[182]&m[183]&m[184]&~m[186]&m[187])|(m[182]&m[183]&m[184]&m[186]&m[187]));
    m[190] = (((m[187]&~m[188]&~m[189]&~m[191]&~m[192])|(~m[187]&m[188]&~m[189]&~m[191]&~m[192])|(~m[187]&~m[188]&m[189]&~m[191]&~m[192])|(m[187]&m[188]&m[189]&m[191]&~m[192])|(~m[187]&~m[188]&~m[189]&~m[191]&m[192])|(m[187]&m[188]&~m[189]&m[191]&m[192])|(m[187]&~m[188]&m[189]&m[191]&m[192])|(~m[187]&m[188]&m[189]&m[191]&m[192]))&UnbiasedRNG[91])|((m[187]&m[188]&~m[189]&~m[191]&~m[192])|(m[187]&~m[188]&m[189]&~m[191]&~m[192])|(~m[187]&m[188]&m[189]&~m[191]&~m[192])|(m[187]&m[188]&m[189]&~m[191]&~m[192])|(m[187]&~m[188]&~m[189]&~m[191]&m[192])|(~m[187]&m[188]&~m[189]&~m[191]&m[192])|(m[187]&m[188]&~m[189]&~m[191]&m[192])|(~m[187]&~m[188]&m[189]&~m[191]&m[192])|(m[187]&~m[188]&m[189]&~m[191]&m[192])|(~m[187]&m[188]&m[189]&~m[191]&m[192])|(m[187]&m[188]&m[189]&~m[191]&m[192])|(m[187]&m[188]&m[189]&m[191]&m[192]));
    m[195] = (((m[192]&~m[193]&~m[194]&~m[196]&~m[197])|(~m[192]&m[193]&~m[194]&~m[196]&~m[197])|(~m[192]&~m[193]&m[194]&~m[196]&~m[197])|(m[192]&m[193]&m[194]&m[196]&~m[197])|(~m[192]&~m[193]&~m[194]&~m[196]&m[197])|(m[192]&m[193]&~m[194]&m[196]&m[197])|(m[192]&~m[193]&m[194]&m[196]&m[197])|(~m[192]&m[193]&m[194]&m[196]&m[197]))&UnbiasedRNG[92])|((m[192]&m[193]&~m[194]&~m[196]&~m[197])|(m[192]&~m[193]&m[194]&~m[196]&~m[197])|(~m[192]&m[193]&m[194]&~m[196]&~m[197])|(m[192]&m[193]&m[194]&~m[196]&~m[197])|(m[192]&~m[193]&~m[194]&~m[196]&m[197])|(~m[192]&m[193]&~m[194]&~m[196]&m[197])|(m[192]&m[193]&~m[194]&~m[196]&m[197])|(~m[192]&~m[193]&m[194]&~m[196]&m[197])|(m[192]&~m[193]&m[194]&~m[196]&m[197])|(~m[192]&m[193]&m[194]&~m[196]&m[197])|(m[192]&m[193]&m[194]&~m[196]&m[197])|(m[192]&m[193]&m[194]&m[196]&m[197]));
    m[200] = (((m[197]&~m[198]&~m[199]&~m[201]&~m[202])|(~m[197]&m[198]&~m[199]&~m[201]&~m[202])|(~m[197]&~m[198]&m[199]&~m[201]&~m[202])|(m[197]&m[198]&m[199]&m[201]&~m[202])|(~m[197]&~m[198]&~m[199]&~m[201]&m[202])|(m[197]&m[198]&~m[199]&m[201]&m[202])|(m[197]&~m[198]&m[199]&m[201]&m[202])|(~m[197]&m[198]&m[199]&m[201]&m[202]))&UnbiasedRNG[93])|((m[197]&m[198]&~m[199]&~m[201]&~m[202])|(m[197]&~m[198]&m[199]&~m[201]&~m[202])|(~m[197]&m[198]&m[199]&~m[201]&~m[202])|(m[197]&m[198]&m[199]&~m[201]&~m[202])|(m[197]&~m[198]&~m[199]&~m[201]&m[202])|(~m[197]&m[198]&~m[199]&~m[201]&m[202])|(m[197]&m[198]&~m[199]&~m[201]&m[202])|(~m[197]&~m[198]&m[199]&~m[201]&m[202])|(m[197]&~m[198]&m[199]&~m[201]&m[202])|(~m[197]&m[198]&m[199]&~m[201]&m[202])|(m[197]&m[198]&m[199]&~m[201]&m[202])|(m[197]&m[198]&m[199]&m[201]&m[202]));
    m[210] = (((m[207]&~m[208]&~m[209]&~m[211]&~m[212])|(~m[207]&m[208]&~m[209]&~m[211]&~m[212])|(~m[207]&~m[208]&m[209]&~m[211]&~m[212])|(m[207]&m[208]&m[209]&m[211]&~m[212])|(~m[207]&~m[208]&~m[209]&~m[211]&m[212])|(m[207]&m[208]&~m[209]&m[211]&m[212])|(m[207]&~m[208]&m[209]&m[211]&m[212])|(~m[207]&m[208]&m[209]&m[211]&m[212]))&UnbiasedRNG[94])|((m[207]&m[208]&~m[209]&~m[211]&~m[212])|(m[207]&~m[208]&m[209]&~m[211]&~m[212])|(~m[207]&m[208]&m[209]&~m[211]&~m[212])|(m[207]&m[208]&m[209]&~m[211]&~m[212])|(m[207]&~m[208]&~m[209]&~m[211]&m[212])|(~m[207]&m[208]&~m[209]&~m[211]&m[212])|(m[207]&m[208]&~m[209]&~m[211]&m[212])|(~m[207]&~m[208]&m[209]&~m[211]&m[212])|(m[207]&~m[208]&m[209]&~m[211]&m[212])|(~m[207]&m[208]&m[209]&~m[211]&m[212])|(m[207]&m[208]&m[209]&~m[211]&m[212])|(m[207]&m[208]&m[209]&m[211]&m[212]));
    m[215] = (((m[212]&~m[213]&~m[214]&~m[216]&~m[217])|(~m[212]&m[213]&~m[214]&~m[216]&~m[217])|(~m[212]&~m[213]&m[214]&~m[216]&~m[217])|(m[212]&m[213]&m[214]&m[216]&~m[217])|(~m[212]&~m[213]&~m[214]&~m[216]&m[217])|(m[212]&m[213]&~m[214]&m[216]&m[217])|(m[212]&~m[213]&m[214]&m[216]&m[217])|(~m[212]&m[213]&m[214]&m[216]&m[217]))&UnbiasedRNG[95])|((m[212]&m[213]&~m[214]&~m[216]&~m[217])|(m[212]&~m[213]&m[214]&~m[216]&~m[217])|(~m[212]&m[213]&m[214]&~m[216]&~m[217])|(m[212]&m[213]&m[214]&~m[216]&~m[217])|(m[212]&~m[213]&~m[214]&~m[216]&m[217])|(~m[212]&m[213]&~m[214]&~m[216]&m[217])|(m[212]&m[213]&~m[214]&~m[216]&m[217])|(~m[212]&~m[213]&m[214]&~m[216]&m[217])|(m[212]&~m[213]&m[214]&~m[216]&m[217])|(~m[212]&m[213]&m[214]&~m[216]&m[217])|(m[212]&m[213]&m[214]&~m[216]&m[217])|(m[212]&m[213]&m[214]&m[216]&m[217]));
    m[220] = (((m[217]&~m[218]&~m[219]&~m[221]&~m[222])|(~m[217]&m[218]&~m[219]&~m[221]&~m[222])|(~m[217]&~m[218]&m[219]&~m[221]&~m[222])|(m[217]&m[218]&m[219]&m[221]&~m[222])|(~m[217]&~m[218]&~m[219]&~m[221]&m[222])|(m[217]&m[218]&~m[219]&m[221]&m[222])|(m[217]&~m[218]&m[219]&m[221]&m[222])|(~m[217]&m[218]&m[219]&m[221]&m[222]))&UnbiasedRNG[96])|((m[217]&m[218]&~m[219]&~m[221]&~m[222])|(m[217]&~m[218]&m[219]&~m[221]&~m[222])|(~m[217]&m[218]&m[219]&~m[221]&~m[222])|(m[217]&m[218]&m[219]&~m[221]&~m[222])|(m[217]&~m[218]&~m[219]&~m[221]&m[222])|(~m[217]&m[218]&~m[219]&~m[221]&m[222])|(m[217]&m[218]&~m[219]&~m[221]&m[222])|(~m[217]&~m[218]&m[219]&~m[221]&m[222])|(m[217]&~m[218]&m[219]&~m[221]&m[222])|(~m[217]&m[218]&m[219]&~m[221]&m[222])|(m[217]&m[218]&m[219]&~m[221]&m[222])|(m[217]&m[218]&m[219]&m[221]&m[222]));
    m[225] = (((m[222]&~m[223]&~m[224]&~m[226]&~m[227])|(~m[222]&m[223]&~m[224]&~m[226]&~m[227])|(~m[222]&~m[223]&m[224]&~m[226]&~m[227])|(m[222]&m[223]&m[224]&m[226]&~m[227])|(~m[222]&~m[223]&~m[224]&~m[226]&m[227])|(m[222]&m[223]&~m[224]&m[226]&m[227])|(m[222]&~m[223]&m[224]&m[226]&m[227])|(~m[222]&m[223]&m[224]&m[226]&m[227]))&UnbiasedRNG[97])|((m[222]&m[223]&~m[224]&~m[226]&~m[227])|(m[222]&~m[223]&m[224]&~m[226]&~m[227])|(~m[222]&m[223]&m[224]&~m[226]&~m[227])|(m[222]&m[223]&m[224]&~m[226]&~m[227])|(m[222]&~m[223]&~m[224]&~m[226]&m[227])|(~m[222]&m[223]&~m[224]&~m[226]&m[227])|(m[222]&m[223]&~m[224]&~m[226]&m[227])|(~m[222]&~m[223]&m[224]&~m[226]&m[227])|(m[222]&~m[223]&m[224]&~m[226]&m[227])|(~m[222]&m[223]&m[224]&~m[226]&m[227])|(m[222]&m[223]&m[224]&~m[226]&m[227])|(m[222]&m[223]&m[224]&m[226]&m[227]));
    m[235] = (((m[232]&~m[233]&~m[234]&~m[236]&~m[237])|(~m[232]&m[233]&~m[234]&~m[236]&~m[237])|(~m[232]&~m[233]&m[234]&~m[236]&~m[237])|(m[232]&m[233]&m[234]&m[236]&~m[237])|(~m[232]&~m[233]&~m[234]&~m[236]&m[237])|(m[232]&m[233]&~m[234]&m[236]&m[237])|(m[232]&~m[233]&m[234]&m[236]&m[237])|(~m[232]&m[233]&m[234]&m[236]&m[237]))&UnbiasedRNG[98])|((m[232]&m[233]&~m[234]&~m[236]&~m[237])|(m[232]&~m[233]&m[234]&~m[236]&~m[237])|(~m[232]&m[233]&m[234]&~m[236]&~m[237])|(m[232]&m[233]&m[234]&~m[236]&~m[237])|(m[232]&~m[233]&~m[234]&~m[236]&m[237])|(~m[232]&m[233]&~m[234]&~m[236]&m[237])|(m[232]&m[233]&~m[234]&~m[236]&m[237])|(~m[232]&~m[233]&m[234]&~m[236]&m[237])|(m[232]&~m[233]&m[234]&~m[236]&m[237])|(~m[232]&m[233]&m[234]&~m[236]&m[237])|(m[232]&m[233]&m[234]&~m[236]&m[237])|(m[232]&m[233]&m[234]&m[236]&m[237]));
    m[240] = (((m[237]&~m[238]&~m[239]&~m[241]&~m[242])|(~m[237]&m[238]&~m[239]&~m[241]&~m[242])|(~m[237]&~m[238]&m[239]&~m[241]&~m[242])|(m[237]&m[238]&m[239]&m[241]&~m[242])|(~m[237]&~m[238]&~m[239]&~m[241]&m[242])|(m[237]&m[238]&~m[239]&m[241]&m[242])|(m[237]&~m[238]&m[239]&m[241]&m[242])|(~m[237]&m[238]&m[239]&m[241]&m[242]))&UnbiasedRNG[99])|((m[237]&m[238]&~m[239]&~m[241]&~m[242])|(m[237]&~m[238]&m[239]&~m[241]&~m[242])|(~m[237]&m[238]&m[239]&~m[241]&~m[242])|(m[237]&m[238]&m[239]&~m[241]&~m[242])|(m[237]&~m[238]&~m[239]&~m[241]&m[242])|(~m[237]&m[238]&~m[239]&~m[241]&m[242])|(m[237]&m[238]&~m[239]&~m[241]&m[242])|(~m[237]&~m[238]&m[239]&~m[241]&m[242])|(m[237]&~m[238]&m[239]&~m[241]&m[242])|(~m[237]&m[238]&m[239]&~m[241]&m[242])|(m[237]&m[238]&m[239]&~m[241]&m[242])|(m[237]&m[238]&m[239]&m[241]&m[242]));
    m[245] = (((m[242]&~m[243]&~m[244]&~m[246]&~m[247])|(~m[242]&m[243]&~m[244]&~m[246]&~m[247])|(~m[242]&~m[243]&m[244]&~m[246]&~m[247])|(m[242]&m[243]&m[244]&m[246]&~m[247])|(~m[242]&~m[243]&~m[244]&~m[246]&m[247])|(m[242]&m[243]&~m[244]&m[246]&m[247])|(m[242]&~m[243]&m[244]&m[246]&m[247])|(~m[242]&m[243]&m[244]&m[246]&m[247]))&UnbiasedRNG[100])|((m[242]&m[243]&~m[244]&~m[246]&~m[247])|(m[242]&~m[243]&m[244]&~m[246]&~m[247])|(~m[242]&m[243]&m[244]&~m[246]&~m[247])|(m[242]&m[243]&m[244]&~m[246]&~m[247])|(m[242]&~m[243]&~m[244]&~m[246]&m[247])|(~m[242]&m[243]&~m[244]&~m[246]&m[247])|(m[242]&m[243]&~m[244]&~m[246]&m[247])|(~m[242]&~m[243]&m[244]&~m[246]&m[247])|(m[242]&~m[243]&m[244]&~m[246]&m[247])|(~m[242]&m[243]&m[244]&~m[246]&m[247])|(m[242]&m[243]&m[244]&~m[246]&m[247])|(m[242]&m[243]&m[244]&m[246]&m[247]));
    m[255] = (((m[252]&~m[253]&~m[254]&~m[256]&~m[257])|(~m[252]&m[253]&~m[254]&~m[256]&~m[257])|(~m[252]&~m[253]&m[254]&~m[256]&~m[257])|(m[252]&m[253]&m[254]&m[256]&~m[257])|(~m[252]&~m[253]&~m[254]&~m[256]&m[257])|(m[252]&m[253]&~m[254]&m[256]&m[257])|(m[252]&~m[253]&m[254]&m[256]&m[257])|(~m[252]&m[253]&m[254]&m[256]&m[257]))&UnbiasedRNG[101])|((m[252]&m[253]&~m[254]&~m[256]&~m[257])|(m[252]&~m[253]&m[254]&~m[256]&~m[257])|(~m[252]&m[253]&m[254]&~m[256]&~m[257])|(m[252]&m[253]&m[254]&~m[256]&~m[257])|(m[252]&~m[253]&~m[254]&~m[256]&m[257])|(~m[252]&m[253]&~m[254]&~m[256]&m[257])|(m[252]&m[253]&~m[254]&~m[256]&m[257])|(~m[252]&~m[253]&m[254]&~m[256]&m[257])|(m[252]&~m[253]&m[254]&~m[256]&m[257])|(~m[252]&m[253]&m[254]&~m[256]&m[257])|(m[252]&m[253]&m[254]&~m[256]&m[257])|(m[252]&m[253]&m[254]&m[256]&m[257]));
    m[260] = (((m[257]&~m[258]&~m[259]&~m[261]&~m[262])|(~m[257]&m[258]&~m[259]&~m[261]&~m[262])|(~m[257]&~m[258]&m[259]&~m[261]&~m[262])|(m[257]&m[258]&m[259]&m[261]&~m[262])|(~m[257]&~m[258]&~m[259]&~m[261]&m[262])|(m[257]&m[258]&~m[259]&m[261]&m[262])|(m[257]&~m[258]&m[259]&m[261]&m[262])|(~m[257]&m[258]&m[259]&m[261]&m[262]))&UnbiasedRNG[102])|((m[257]&m[258]&~m[259]&~m[261]&~m[262])|(m[257]&~m[258]&m[259]&~m[261]&~m[262])|(~m[257]&m[258]&m[259]&~m[261]&~m[262])|(m[257]&m[258]&m[259]&~m[261]&~m[262])|(m[257]&~m[258]&~m[259]&~m[261]&m[262])|(~m[257]&m[258]&~m[259]&~m[261]&m[262])|(m[257]&m[258]&~m[259]&~m[261]&m[262])|(~m[257]&~m[258]&m[259]&~m[261]&m[262])|(m[257]&~m[258]&m[259]&~m[261]&m[262])|(~m[257]&m[258]&m[259]&~m[261]&m[262])|(m[257]&m[258]&m[259]&~m[261]&m[262])|(m[257]&m[258]&m[259]&m[261]&m[262]));
    m[270] = (((m[267]&~m[268]&~m[269]&~m[271]&~m[272])|(~m[267]&m[268]&~m[269]&~m[271]&~m[272])|(~m[267]&~m[268]&m[269]&~m[271]&~m[272])|(m[267]&m[268]&m[269]&m[271]&~m[272])|(~m[267]&~m[268]&~m[269]&~m[271]&m[272])|(m[267]&m[268]&~m[269]&m[271]&m[272])|(m[267]&~m[268]&m[269]&m[271]&m[272])|(~m[267]&m[268]&m[269]&m[271]&m[272]))&UnbiasedRNG[103])|((m[267]&m[268]&~m[269]&~m[271]&~m[272])|(m[267]&~m[268]&m[269]&~m[271]&~m[272])|(~m[267]&m[268]&m[269]&~m[271]&~m[272])|(m[267]&m[268]&m[269]&~m[271]&~m[272])|(m[267]&~m[268]&~m[269]&~m[271]&m[272])|(~m[267]&m[268]&~m[269]&~m[271]&m[272])|(m[267]&m[268]&~m[269]&~m[271]&m[272])|(~m[267]&~m[268]&m[269]&~m[271]&m[272])|(m[267]&~m[268]&m[269]&~m[271]&m[272])|(~m[267]&m[268]&m[269]&~m[271]&m[272])|(m[267]&m[268]&m[269]&~m[271]&m[272])|(m[267]&m[268]&m[269]&m[271]&m[272]));
end

always @(posedge color4_clk) begin
    m[136] = (((m[132]&~m[133]&~m[134]&~m[135]&~m[139])|(~m[132]&m[133]&~m[134]&~m[135]&~m[139])|(~m[132]&~m[133]&m[134]&~m[135]&~m[139])|(m[132]&m[133]&~m[134]&m[135]&~m[139])|(m[132]&~m[133]&m[134]&m[135]&~m[139])|(~m[132]&m[133]&m[134]&m[135]&~m[139]))&BiasedRNG[131])|(((m[132]&~m[133]&~m[134]&~m[135]&m[139])|(~m[132]&m[133]&~m[134]&~m[135]&m[139])|(~m[132]&~m[133]&m[134]&~m[135]&m[139])|(m[132]&m[133]&~m[134]&m[135]&m[139])|(m[132]&~m[133]&m[134]&m[135]&m[139])|(~m[132]&m[133]&m[134]&m[135]&m[139]))&~BiasedRNG[131])|((m[132]&m[133]&~m[134]&~m[135]&~m[139])|(m[132]&~m[133]&m[134]&~m[135]&~m[139])|(~m[132]&m[133]&m[134]&~m[135]&~m[139])|(m[132]&m[133]&m[134]&~m[135]&~m[139])|(m[132]&m[133]&m[134]&m[135]&~m[139])|(m[132]&m[133]&~m[134]&~m[135]&m[139])|(m[132]&~m[133]&m[134]&~m[135]&m[139])|(~m[132]&m[133]&m[134]&~m[135]&m[139])|(m[132]&m[133]&m[134]&~m[135]&m[139])|(m[132]&m[133]&m[134]&m[135]&m[139]));
    m[141] = (((m[137]&~m[138]&~m[139]&~m[140]&~m[149])|(~m[137]&m[138]&~m[139]&~m[140]&~m[149])|(~m[137]&~m[138]&m[139]&~m[140]&~m[149])|(m[137]&m[138]&~m[139]&m[140]&~m[149])|(m[137]&~m[138]&m[139]&m[140]&~m[149])|(~m[137]&m[138]&m[139]&m[140]&~m[149]))&BiasedRNG[132])|(((m[137]&~m[138]&~m[139]&~m[140]&m[149])|(~m[137]&m[138]&~m[139]&~m[140]&m[149])|(~m[137]&~m[138]&m[139]&~m[140]&m[149])|(m[137]&m[138]&~m[139]&m[140]&m[149])|(m[137]&~m[138]&m[139]&m[140]&m[149])|(~m[137]&m[138]&m[139]&m[140]&m[149]))&~BiasedRNG[132])|((m[137]&m[138]&~m[139]&~m[140]&~m[149])|(m[137]&~m[138]&m[139]&~m[140]&~m[149])|(~m[137]&m[138]&m[139]&~m[140]&~m[149])|(m[137]&m[138]&m[139]&~m[140]&~m[149])|(m[137]&m[138]&m[139]&m[140]&~m[149])|(m[137]&m[138]&~m[139]&~m[140]&m[149])|(m[137]&~m[138]&m[139]&~m[140]&m[149])|(~m[137]&m[138]&m[139]&~m[140]&m[149])|(m[137]&m[138]&m[139]&~m[140]&m[149])|(m[137]&m[138]&m[139]&m[140]&m[149]));
    m[146] = (((m[142]&~m[143]&~m[144]&~m[145]&~m[154])|(~m[142]&m[143]&~m[144]&~m[145]&~m[154])|(~m[142]&~m[143]&m[144]&~m[145]&~m[154])|(m[142]&m[143]&~m[144]&m[145]&~m[154])|(m[142]&~m[143]&m[144]&m[145]&~m[154])|(~m[142]&m[143]&m[144]&m[145]&~m[154]))&BiasedRNG[133])|(((m[142]&~m[143]&~m[144]&~m[145]&m[154])|(~m[142]&m[143]&~m[144]&~m[145]&m[154])|(~m[142]&~m[143]&m[144]&~m[145]&m[154])|(m[142]&m[143]&~m[144]&m[145]&m[154])|(m[142]&~m[143]&m[144]&m[145]&m[154])|(~m[142]&m[143]&m[144]&m[145]&m[154]))&~BiasedRNG[133])|((m[142]&m[143]&~m[144]&~m[145]&~m[154])|(m[142]&~m[143]&m[144]&~m[145]&~m[154])|(~m[142]&m[143]&m[144]&~m[145]&~m[154])|(m[142]&m[143]&m[144]&~m[145]&~m[154])|(m[142]&m[143]&m[144]&m[145]&~m[154])|(m[142]&m[143]&~m[144]&~m[145]&m[154])|(m[142]&~m[143]&m[144]&~m[145]&m[154])|(~m[142]&m[143]&m[144]&~m[145]&m[154])|(m[142]&m[143]&m[144]&~m[145]&m[154])|(m[142]&m[143]&m[144]&m[145]&m[154]));
    m[151] = (((m[147]&~m[148]&~m[149]&~m[150]&~m[164])|(~m[147]&m[148]&~m[149]&~m[150]&~m[164])|(~m[147]&~m[148]&m[149]&~m[150]&~m[164])|(m[147]&m[148]&~m[149]&m[150]&~m[164])|(m[147]&~m[148]&m[149]&m[150]&~m[164])|(~m[147]&m[148]&m[149]&m[150]&~m[164]))&BiasedRNG[134])|(((m[147]&~m[148]&~m[149]&~m[150]&m[164])|(~m[147]&m[148]&~m[149]&~m[150]&m[164])|(~m[147]&~m[148]&m[149]&~m[150]&m[164])|(m[147]&m[148]&~m[149]&m[150]&m[164])|(m[147]&~m[148]&m[149]&m[150]&m[164])|(~m[147]&m[148]&m[149]&m[150]&m[164]))&~BiasedRNG[134])|((m[147]&m[148]&~m[149]&~m[150]&~m[164])|(m[147]&~m[148]&m[149]&~m[150]&~m[164])|(~m[147]&m[148]&m[149]&~m[150]&~m[164])|(m[147]&m[148]&m[149]&~m[150]&~m[164])|(m[147]&m[148]&m[149]&m[150]&~m[164])|(m[147]&m[148]&~m[149]&~m[150]&m[164])|(m[147]&~m[148]&m[149]&~m[150]&m[164])|(~m[147]&m[148]&m[149]&~m[150]&m[164])|(m[147]&m[148]&m[149]&~m[150]&m[164])|(m[147]&m[148]&m[149]&m[150]&m[164]));
    m[156] = (((m[152]&~m[153]&~m[154]&~m[155]&~m[169])|(~m[152]&m[153]&~m[154]&~m[155]&~m[169])|(~m[152]&~m[153]&m[154]&~m[155]&~m[169])|(m[152]&m[153]&~m[154]&m[155]&~m[169])|(m[152]&~m[153]&m[154]&m[155]&~m[169])|(~m[152]&m[153]&m[154]&m[155]&~m[169]))&BiasedRNG[135])|(((m[152]&~m[153]&~m[154]&~m[155]&m[169])|(~m[152]&m[153]&~m[154]&~m[155]&m[169])|(~m[152]&~m[153]&m[154]&~m[155]&m[169])|(m[152]&m[153]&~m[154]&m[155]&m[169])|(m[152]&~m[153]&m[154]&m[155]&m[169])|(~m[152]&m[153]&m[154]&m[155]&m[169]))&~BiasedRNG[135])|((m[152]&m[153]&~m[154]&~m[155]&~m[169])|(m[152]&~m[153]&m[154]&~m[155]&~m[169])|(~m[152]&m[153]&m[154]&~m[155]&~m[169])|(m[152]&m[153]&m[154]&~m[155]&~m[169])|(m[152]&m[153]&m[154]&m[155]&~m[169])|(m[152]&m[153]&~m[154]&~m[155]&m[169])|(m[152]&~m[153]&m[154]&~m[155]&m[169])|(~m[152]&m[153]&m[154]&~m[155]&m[169])|(m[152]&m[153]&m[154]&~m[155]&m[169])|(m[152]&m[153]&m[154]&m[155]&m[169]));
    m[161] = (((m[157]&~m[158]&~m[159]&~m[160]&~m[174])|(~m[157]&m[158]&~m[159]&~m[160]&~m[174])|(~m[157]&~m[158]&m[159]&~m[160]&~m[174])|(m[157]&m[158]&~m[159]&m[160]&~m[174])|(m[157]&~m[158]&m[159]&m[160]&~m[174])|(~m[157]&m[158]&m[159]&m[160]&~m[174]))&BiasedRNG[136])|(((m[157]&~m[158]&~m[159]&~m[160]&m[174])|(~m[157]&m[158]&~m[159]&~m[160]&m[174])|(~m[157]&~m[158]&m[159]&~m[160]&m[174])|(m[157]&m[158]&~m[159]&m[160]&m[174])|(m[157]&~m[158]&m[159]&m[160]&m[174])|(~m[157]&m[158]&m[159]&m[160]&m[174]))&~BiasedRNG[136])|((m[157]&m[158]&~m[159]&~m[160]&~m[174])|(m[157]&~m[158]&m[159]&~m[160]&~m[174])|(~m[157]&m[158]&m[159]&~m[160]&~m[174])|(m[157]&m[158]&m[159]&~m[160]&~m[174])|(m[157]&m[158]&m[159]&m[160]&~m[174])|(m[157]&m[158]&~m[159]&~m[160]&m[174])|(m[157]&~m[158]&m[159]&~m[160]&m[174])|(~m[157]&m[158]&m[159]&~m[160]&m[174])|(m[157]&m[158]&m[159]&~m[160]&m[174])|(m[157]&m[158]&m[159]&m[160]&m[174]));
    m[166] = (((m[162]&~m[163]&~m[164]&~m[165]&~m[184])|(~m[162]&m[163]&~m[164]&~m[165]&~m[184])|(~m[162]&~m[163]&m[164]&~m[165]&~m[184])|(m[162]&m[163]&~m[164]&m[165]&~m[184])|(m[162]&~m[163]&m[164]&m[165]&~m[184])|(~m[162]&m[163]&m[164]&m[165]&~m[184]))&BiasedRNG[137])|(((m[162]&~m[163]&~m[164]&~m[165]&m[184])|(~m[162]&m[163]&~m[164]&~m[165]&m[184])|(~m[162]&~m[163]&m[164]&~m[165]&m[184])|(m[162]&m[163]&~m[164]&m[165]&m[184])|(m[162]&~m[163]&m[164]&m[165]&m[184])|(~m[162]&m[163]&m[164]&m[165]&m[184]))&~BiasedRNG[137])|((m[162]&m[163]&~m[164]&~m[165]&~m[184])|(m[162]&~m[163]&m[164]&~m[165]&~m[184])|(~m[162]&m[163]&m[164]&~m[165]&~m[184])|(m[162]&m[163]&m[164]&~m[165]&~m[184])|(m[162]&m[163]&m[164]&m[165]&~m[184])|(m[162]&m[163]&~m[164]&~m[165]&m[184])|(m[162]&~m[163]&m[164]&~m[165]&m[184])|(~m[162]&m[163]&m[164]&~m[165]&m[184])|(m[162]&m[163]&m[164]&~m[165]&m[184])|(m[162]&m[163]&m[164]&m[165]&m[184]));
    m[171] = (((m[167]&~m[168]&~m[169]&~m[170]&~m[189])|(~m[167]&m[168]&~m[169]&~m[170]&~m[189])|(~m[167]&~m[168]&m[169]&~m[170]&~m[189])|(m[167]&m[168]&~m[169]&m[170]&~m[189])|(m[167]&~m[168]&m[169]&m[170]&~m[189])|(~m[167]&m[168]&m[169]&m[170]&~m[189]))&BiasedRNG[138])|(((m[167]&~m[168]&~m[169]&~m[170]&m[189])|(~m[167]&m[168]&~m[169]&~m[170]&m[189])|(~m[167]&~m[168]&m[169]&~m[170]&m[189])|(m[167]&m[168]&~m[169]&m[170]&m[189])|(m[167]&~m[168]&m[169]&m[170]&m[189])|(~m[167]&m[168]&m[169]&m[170]&m[189]))&~BiasedRNG[138])|((m[167]&m[168]&~m[169]&~m[170]&~m[189])|(m[167]&~m[168]&m[169]&~m[170]&~m[189])|(~m[167]&m[168]&m[169]&~m[170]&~m[189])|(m[167]&m[168]&m[169]&~m[170]&~m[189])|(m[167]&m[168]&m[169]&m[170]&~m[189])|(m[167]&m[168]&~m[169]&~m[170]&m[189])|(m[167]&~m[168]&m[169]&~m[170]&m[189])|(~m[167]&m[168]&m[169]&~m[170]&m[189])|(m[167]&m[168]&m[169]&~m[170]&m[189])|(m[167]&m[168]&m[169]&m[170]&m[189]));
    m[176] = (((m[172]&~m[173]&~m[174]&~m[175]&~m[194])|(~m[172]&m[173]&~m[174]&~m[175]&~m[194])|(~m[172]&~m[173]&m[174]&~m[175]&~m[194])|(m[172]&m[173]&~m[174]&m[175]&~m[194])|(m[172]&~m[173]&m[174]&m[175]&~m[194])|(~m[172]&m[173]&m[174]&m[175]&~m[194]))&BiasedRNG[139])|(((m[172]&~m[173]&~m[174]&~m[175]&m[194])|(~m[172]&m[173]&~m[174]&~m[175]&m[194])|(~m[172]&~m[173]&m[174]&~m[175]&m[194])|(m[172]&m[173]&~m[174]&m[175]&m[194])|(m[172]&~m[173]&m[174]&m[175]&m[194])|(~m[172]&m[173]&m[174]&m[175]&m[194]))&~BiasedRNG[139])|((m[172]&m[173]&~m[174]&~m[175]&~m[194])|(m[172]&~m[173]&m[174]&~m[175]&~m[194])|(~m[172]&m[173]&m[174]&~m[175]&~m[194])|(m[172]&m[173]&m[174]&~m[175]&~m[194])|(m[172]&m[173]&m[174]&m[175]&~m[194])|(m[172]&m[173]&~m[174]&~m[175]&m[194])|(m[172]&~m[173]&m[174]&~m[175]&m[194])|(~m[172]&m[173]&m[174]&~m[175]&m[194])|(m[172]&m[173]&m[174]&~m[175]&m[194])|(m[172]&m[173]&m[174]&m[175]&m[194]));
    m[181] = (((m[177]&~m[178]&~m[179]&~m[180]&~m[199])|(~m[177]&m[178]&~m[179]&~m[180]&~m[199])|(~m[177]&~m[178]&m[179]&~m[180]&~m[199])|(m[177]&m[178]&~m[179]&m[180]&~m[199])|(m[177]&~m[178]&m[179]&m[180]&~m[199])|(~m[177]&m[178]&m[179]&m[180]&~m[199]))&BiasedRNG[140])|(((m[177]&~m[178]&~m[179]&~m[180]&m[199])|(~m[177]&m[178]&~m[179]&~m[180]&m[199])|(~m[177]&~m[178]&m[179]&~m[180]&m[199])|(m[177]&m[178]&~m[179]&m[180]&m[199])|(m[177]&~m[178]&m[179]&m[180]&m[199])|(~m[177]&m[178]&m[179]&m[180]&m[199]))&~BiasedRNG[140])|((m[177]&m[178]&~m[179]&~m[180]&~m[199])|(m[177]&~m[178]&m[179]&~m[180]&~m[199])|(~m[177]&m[178]&m[179]&~m[180]&~m[199])|(m[177]&m[178]&m[179]&~m[180]&~m[199])|(m[177]&m[178]&m[179]&m[180]&~m[199])|(m[177]&m[178]&~m[179]&~m[180]&m[199])|(m[177]&~m[178]&m[179]&~m[180]&m[199])|(~m[177]&m[178]&m[179]&~m[180]&m[199])|(m[177]&m[178]&m[179]&~m[180]&m[199])|(m[177]&m[178]&m[179]&m[180]&m[199]));
    m[186] = (((m[182]&~m[183]&~m[184]&~m[185]&~m[209])|(~m[182]&m[183]&~m[184]&~m[185]&~m[209])|(~m[182]&~m[183]&m[184]&~m[185]&~m[209])|(m[182]&m[183]&~m[184]&m[185]&~m[209])|(m[182]&~m[183]&m[184]&m[185]&~m[209])|(~m[182]&m[183]&m[184]&m[185]&~m[209]))&BiasedRNG[141])|(((m[182]&~m[183]&~m[184]&~m[185]&m[209])|(~m[182]&m[183]&~m[184]&~m[185]&m[209])|(~m[182]&~m[183]&m[184]&~m[185]&m[209])|(m[182]&m[183]&~m[184]&m[185]&m[209])|(m[182]&~m[183]&m[184]&m[185]&m[209])|(~m[182]&m[183]&m[184]&m[185]&m[209]))&~BiasedRNG[141])|((m[182]&m[183]&~m[184]&~m[185]&~m[209])|(m[182]&~m[183]&m[184]&~m[185]&~m[209])|(~m[182]&m[183]&m[184]&~m[185]&~m[209])|(m[182]&m[183]&m[184]&~m[185]&~m[209])|(m[182]&m[183]&m[184]&m[185]&~m[209])|(m[182]&m[183]&~m[184]&~m[185]&m[209])|(m[182]&~m[183]&m[184]&~m[185]&m[209])|(~m[182]&m[183]&m[184]&~m[185]&m[209])|(m[182]&m[183]&m[184]&~m[185]&m[209])|(m[182]&m[183]&m[184]&m[185]&m[209]));
    m[191] = (((m[187]&~m[188]&~m[189]&~m[190]&~m[214])|(~m[187]&m[188]&~m[189]&~m[190]&~m[214])|(~m[187]&~m[188]&m[189]&~m[190]&~m[214])|(m[187]&m[188]&~m[189]&m[190]&~m[214])|(m[187]&~m[188]&m[189]&m[190]&~m[214])|(~m[187]&m[188]&m[189]&m[190]&~m[214]))&BiasedRNG[142])|(((m[187]&~m[188]&~m[189]&~m[190]&m[214])|(~m[187]&m[188]&~m[189]&~m[190]&m[214])|(~m[187]&~m[188]&m[189]&~m[190]&m[214])|(m[187]&m[188]&~m[189]&m[190]&m[214])|(m[187]&~m[188]&m[189]&m[190]&m[214])|(~m[187]&m[188]&m[189]&m[190]&m[214]))&~BiasedRNG[142])|((m[187]&m[188]&~m[189]&~m[190]&~m[214])|(m[187]&~m[188]&m[189]&~m[190]&~m[214])|(~m[187]&m[188]&m[189]&~m[190]&~m[214])|(m[187]&m[188]&m[189]&~m[190]&~m[214])|(m[187]&m[188]&m[189]&m[190]&~m[214])|(m[187]&m[188]&~m[189]&~m[190]&m[214])|(m[187]&~m[188]&m[189]&~m[190]&m[214])|(~m[187]&m[188]&m[189]&~m[190]&m[214])|(m[187]&m[188]&m[189]&~m[190]&m[214])|(m[187]&m[188]&m[189]&m[190]&m[214]));
    m[196] = (((m[192]&~m[193]&~m[194]&~m[195]&~m[219])|(~m[192]&m[193]&~m[194]&~m[195]&~m[219])|(~m[192]&~m[193]&m[194]&~m[195]&~m[219])|(m[192]&m[193]&~m[194]&m[195]&~m[219])|(m[192]&~m[193]&m[194]&m[195]&~m[219])|(~m[192]&m[193]&m[194]&m[195]&~m[219]))&BiasedRNG[143])|(((m[192]&~m[193]&~m[194]&~m[195]&m[219])|(~m[192]&m[193]&~m[194]&~m[195]&m[219])|(~m[192]&~m[193]&m[194]&~m[195]&m[219])|(m[192]&m[193]&~m[194]&m[195]&m[219])|(m[192]&~m[193]&m[194]&m[195]&m[219])|(~m[192]&m[193]&m[194]&m[195]&m[219]))&~BiasedRNG[143])|((m[192]&m[193]&~m[194]&~m[195]&~m[219])|(m[192]&~m[193]&m[194]&~m[195]&~m[219])|(~m[192]&m[193]&m[194]&~m[195]&~m[219])|(m[192]&m[193]&m[194]&~m[195]&~m[219])|(m[192]&m[193]&m[194]&m[195]&~m[219])|(m[192]&m[193]&~m[194]&~m[195]&m[219])|(m[192]&~m[193]&m[194]&~m[195]&m[219])|(~m[192]&m[193]&m[194]&~m[195]&m[219])|(m[192]&m[193]&m[194]&~m[195]&m[219])|(m[192]&m[193]&m[194]&m[195]&m[219]));
    m[201] = (((m[197]&~m[198]&~m[199]&~m[200]&~m[224])|(~m[197]&m[198]&~m[199]&~m[200]&~m[224])|(~m[197]&~m[198]&m[199]&~m[200]&~m[224])|(m[197]&m[198]&~m[199]&m[200]&~m[224])|(m[197]&~m[198]&m[199]&m[200]&~m[224])|(~m[197]&m[198]&m[199]&m[200]&~m[224]))&BiasedRNG[144])|(((m[197]&~m[198]&~m[199]&~m[200]&m[224])|(~m[197]&m[198]&~m[199]&~m[200]&m[224])|(~m[197]&~m[198]&m[199]&~m[200]&m[224])|(m[197]&m[198]&~m[199]&m[200]&m[224])|(m[197]&~m[198]&m[199]&m[200]&m[224])|(~m[197]&m[198]&m[199]&m[200]&m[224]))&~BiasedRNG[144])|((m[197]&m[198]&~m[199]&~m[200]&~m[224])|(m[197]&~m[198]&m[199]&~m[200]&~m[224])|(~m[197]&m[198]&m[199]&~m[200]&~m[224])|(m[197]&m[198]&m[199]&~m[200]&~m[224])|(m[197]&m[198]&m[199]&m[200]&~m[224])|(m[197]&m[198]&~m[199]&~m[200]&m[224])|(m[197]&~m[198]&m[199]&~m[200]&m[224])|(~m[197]&m[198]&m[199]&~m[200]&m[224])|(m[197]&m[198]&m[199]&~m[200]&m[224])|(m[197]&m[198]&m[199]&m[200]&m[224]));
    m[206] = (((m[202]&~m[203]&~m[204]&~m[205]&~m[229])|(~m[202]&m[203]&~m[204]&~m[205]&~m[229])|(~m[202]&~m[203]&m[204]&~m[205]&~m[229])|(m[202]&m[203]&~m[204]&m[205]&~m[229])|(m[202]&~m[203]&m[204]&m[205]&~m[229])|(~m[202]&m[203]&m[204]&m[205]&~m[229]))&BiasedRNG[145])|(((m[202]&~m[203]&~m[204]&~m[205]&m[229])|(~m[202]&m[203]&~m[204]&~m[205]&m[229])|(~m[202]&~m[203]&m[204]&~m[205]&m[229])|(m[202]&m[203]&~m[204]&m[205]&m[229])|(m[202]&~m[203]&m[204]&m[205]&m[229])|(~m[202]&m[203]&m[204]&m[205]&m[229]))&~BiasedRNG[145])|((m[202]&m[203]&~m[204]&~m[205]&~m[229])|(m[202]&~m[203]&m[204]&~m[205]&~m[229])|(~m[202]&m[203]&m[204]&~m[205]&~m[229])|(m[202]&m[203]&m[204]&~m[205]&~m[229])|(m[202]&m[203]&m[204]&m[205]&~m[229])|(m[202]&m[203]&~m[204]&~m[205]&m[229])|(m[202]&~m[203]&m[204]&~m[205]&m[229])|(~m[202]&m[203]&m[204]&~m[205]&m[229])|(m[202]&m[203]&m[204]&~m[205]&m[229])|(m[202]&m[203]&m[204]&m[205]&m[229]));
    m[211] = (((m[207]&~m[208]&~m[209]&~m[210]&~m[232])|(~m[207]&m[208]&~m[209]&~m[210]&~m[232])|(~m[207]&~m[208]&m[209]&~m[210]&~m[232])|(m[207]&m[208]&~m[209]&m[210]&~m[232])|(m[207]&~m[208]&m[209]&m[210]&~m[232])|(~m[207]&m[208]&m[209]&m[210]&~m[232]))&BiasedRNG[146])|(((m[207]&~m[208]&~m[209]&~m[210]&m[232])|(~m[207]&m[208]&~m[209]&~m[210]&m[232])|(~m[207]&~m[208]&m[209]&~m[210]&m[232])|(m[207]&m[208]&~m[209]&m[210]&m[232])|(m[207]&~m[208]&m[209]&m[210]&m[232])|(~m[207]&m[208]&m[209]&m[210]&m[232]))&~BiasedRNG[146])|((m[207]&m[208]&~m[209]&~m[210]&~m[232])|(m[207]&~m[208]&m[209]&~m[210]&~m[232])|(~m[207]&m[208]&m[209]&~m[210]&~m[232])|(m[207]&m[208]&m[209]&~m[210]&~m[232])|(m[207]&m[208]&m[209]&m[210]&~m[232])|(m[207]&m[208]&~m[209]&~m[210]&m[232])|(m[207]&~m[208]&m[209]&~m[210]&m[232])|(~m[207]&m[208]&m[209]&~m[210]&m[232])|(m[207]&m[208]&m[209]&~m[210]&m[232])|(m[207]&m[208]&m[209]&m[210]&m[232]));
    m[216] = (((m[212]&~m[213]&~m[214]&~m[215]&~m[234])|(~m[212]&m[213]&~m[214]&~m[215]&~m[234])|(~m[212]&~m[213]&m[214]&~m[215]&~m[234])|(m[212]&m[213]&~m[214]&m[215]&~m[234])|(m[212]&~m[213]&m[214]&m[215]&~m[234])|(~m[212]&m[213]&m[214]&m[215]&~m[234]))&BiasedRNG[147])|(((m[212]&~m[213]&~m[214]&~m[215]&m[234])|(~m[212]&m[213]&~m[214]&~m[215]&m[234])|(~m[212]&~m[213]&m[214]&~m[215]&m[234])|(m[212]&m[213]&~m[214]&m[215]&m[234])|(m[212]&~m[213]&m[214]&m[215]&m[234])|(~m[212]&m[213]&m[214]&m[215]&m[234]))&~BiasedRNG[147])|((m[212]&m[213]&~m[214]&~m[215]&~m[234])|(m[212]&~m[213]&m[214]&~m[215]&~m[234])|(~m[212]&m[213]&m[214]&~m[215]&~m[234])|(m[212]&m[213]&m[214]&~m[215]&~m[234])|(m[212]&m[213]&m[214]&m[215]&~m[234])|(m[212]&m[213]&~m[214]&~m[215]&m[234])|(m[212]&~m[213]&m[214]&~m[215]&m[234])|(~m[212]&m[213]&m[214]&~m[215]&m[234])|(m[212]&m[213]&m[214]&~m[215]&m[234])|(m[212]&m[213]&m[214]&m[215]&m[234]));
    m[221] = (((m[217]&~m[218]&~m[219]&~m[220]&~m[239])|(~m[217]&m[218]&~m[219]&~m[220]&~m[239])|(~m[217]&~m[218]&m[219]&~m[220]&~m[239])|(m[217]&m[218]&~m[219]&m[220]&~m[239])|(m[217]&~m[218]&m[219]&m[220]&~m[239])|(~m[217]&m[218]&m[219]&m[220]&~m[239]))&BiasedRNG[148])|(((m[217]&~m[218]&~m[219]&~m[220]&m[239])|(~m[217]&m[218]&~m[219]&~m[220]&m[239])|(~m[217]&~m[218]&m[219]&~m[220]&m[239])|(m[217]&m[218]&~m[219]&m[220]&m[239])|(m[217]&~m[218]&m[219]&m[220]&m[239])|(~m[217]&m[218]&m[219]&m[220]&m[239]))&~BiasedRNG[148])|((m[217]&m[218]&~m[219]&~m[220]&~m[239])|(m[217]&~m[218]&m[219]&~m[220]&~m[239])|(~m[217]&m[218]&m[219]&~m[220]&~m[239])|(m[217]&m[218]&m[219]&~m[220]&~m[239])|(m[217]&m[218]&m[219]&m[220]&~m[239])|(m[217]&m[218]&~m[219]&~m[220]&m[239])|(m[217]&~m[218]&m[219]&~m[220]&m[239])|(~m[217]&m[218]&m[219]&~m[220]&m[239])|(m[217]&m[218]&m[219]&~m[220]&m[239])|(m[217]&m[218]&m[219]&m[220]&m[239]));
    m[226] = (((m[222]&~m[223]&~m[224]&~m[225]&~m[244])|(~m[222]&m[223]&~m[224]&~m[225]&~m[244])|(~m[222]&~m[223]&m[224]&~m[225]&~m[244])|(m[222]&m[223]&~m[224]&m[225]&~m[244])|(m[222]&~m[223]&m[224]&m[225]&~m[244])|(~m[222]&m[223]&m[224]&m[225]&~m[244]))&BiasedRNG[149])|(((m[222]&~m[223]&~m[224]&~m[225]&m[244])|(~m[222]&m[223]&~m[224]&~m[225]&m[244])|(~m[222]&~m[223]&m[224]&~m[225]&m[244])|(m[222]&m[223]&~m[224]&m[225]&m[244])|(m[222]&~m[223]&m[224]&m[225]&m[244])|(~m[222]&m[223]&m[224]&m[225]&m[244]))&~BiasedRNG[149])|((m[222]&m[223]&~m[224]&~m[225]&~m[244])|(m[222]&~m[223]&m[224]&~m[225]&~m[244])|(~m[222]&m[223]&m[224]&~m[225]&~m[244])|(m[222]&m[223]&m[224]&~m[225]&~m[244])|(m[222]&m[223]&m[224]&m[225]&~m[244])|(m[222]&m[223]&~m[224]&~m[225]&m[244])|(m[222]&~m[223]&m[224]&~m[225]&m[244])|(~m[222]&m[223]&m[224]&~m[225]&m[244])|(m[222]&m[223]&m[224]&~m[225]&m[244])|(m[222]&m[223]&m[224]&m[225]&m[244]));
    m[231] = (((m[227]&~m[228]&~m[229]&~m[230]&~m[249])|(~m[227]&m[228]&~m[229]&~m[230]&~m[249])|(~m[227]&~m[228]&m[229]&~m[230]&~m[249])|(m[227]&m[228]&~m[229]&m[230]&~m[249])|(m[227]&~m[228]&m[229]&m[230]&~m[249])|(~m[227]&m[228]&m[229]&m[230]&~m[249]))&BiasedRNG[150])|(((m[227]&~m[228]&~m[229]&~m[230]&m[249])|(~m[227]&m[228]&~m[229]&~m[230]&m[249])|(~m[227]&~m[228]&m[229]&~m[230]&m[249])|(m[227]&m[228]&~m[229]&m[230]&m[249])|(m[227]&~m[228]&m[229]&m[230]&m[249])|(~m[227]&m[228]&m[229]&m[230]&m[249]))&~BiasedRNG[150])|((m[227]&m[228]&~m[229]&~m[230]&~m[249])|(m[227]&~m[228]&m[229]&~m[230]&~m[249])|(~m[227]&m[228]&m[229]&~m[230]&~m[249])|(m[227]&m[228]&m[229]&~m[230]&~m[249])|(m[227]&m[228]&m[229]&m[230]&~m[249])|(m[227]&m[228]&~m[229]&~m[230]&m[249])|(m[227]&~m[228]&m[229]&~m[230]&m[249])|(~m[227]&m[228]&m[229]&~m[230]&m[249])|(m[227]&m[228]&m[229]&~m[230]&m[249])|(m[227]&m[228]&m[229]&m[230]&m[249]));
    m[236] = (((m[232]&~m[233]&~m[234]&~m[235]&~m[252])|(~m[232]&m[233]&~m[234]&~m[235]&~m[252])|(~m[232]&~m[233]&m[234]&~m[235]&~m[252])|(m[232]&m[233]&~m[234]&m[235]&~m[252])|(m[232]&~m[233]&m[234]&m[235]&~m[252])|(~m[232]&m[233]&m[234]&m[235]&~m[252]))&BiasedRNG[151])|(((m[232]&~m[233]&~m[234]&~m[235]&m[252])|(~m[232]&m[233]&~m[234]&~m[235]&m[252])|(~m[232]&~m[233]&m[234]&~m[235]&m[252])|(m[232]&m[233]&~m[234]&m[235]&m[252])|(m[232]&~m[233]&m[234]&m[235]&m[252])|(~m[232]&m[233]&m[234]&m[235]&m[252]))&~BiasedRNG[151])|((m[232]&m[233]&~m[234]&~m[235]&~m[252])|(m[232]&~m[233]&m[234]&~m[235]&~m[252])|(~m[232]&m[233]&m[234]&~m[235]&~m[252])|(m[232]&m[233]&m[234]&~m[235]&~m[252])|(m[232]&m[233]&m[234]&m[235]&~m[252])|(m[232]&m[233]&~m[234]&~m[235]&m[252])|(m[232]&~m[233]&m[234]&~m[235]&m[252])|(~m[232]&m[233]&m[234]&~m[235]&m[252])|(m[232]&m[233]&m[234]&~m[235]&m[252])|(m[232]&m[233]&m[234]&m[235]&m[252]));
    m[241] = (((m[237]&~m[238]&~m[239]&~m[240]&~m[254])|(~m[237]&m[238]&~m[239]&~m[240]&~m[254])|(~m[237]&~m[238]&m[239]&~m[240]&~m[254])|(m[237]&m[238]&~m[239]&m[240]&~m[254])|(m[237]&~m[238]&m[239]&m[240]&~m[254])|(~m[237]&m[238]&m[239]&m[240]&~m[254]))&BiasedRNG[152])|(((m[237]&~m[238]&~m[239]&~m[240]&m[254])|(~m[237]&m[238]&~m[239]&~m[240]&m[254])|(~m[237]&~m[238]&m[239]&~m[240]&m[254])|(m[237]&m[238]&~m[239]&m[240]&m[254])|(m[237]&~m[238]&m[239]&m[240]&m[254])|(~m[237]&m[238]&m[239]&m[240]&m[254]))&~BiasedRNG[152])|((m[237]&m[238]&~m[239]&~m[240]&~m[254])|(m[237]&~m[238]&m[239]&~m[240]&~m[254])|(~m[237]&m[238]&m[239]&~m[240]&~m[254])|(m[237]&m[238]&m[239]&~m[240]&~m[254])|(m[237]&m[238]&m[239]&m[240]&~m[254])|(m[237]&m[238]&~m[239]&~m[240]&m[254])|(m[237]&~m[238]&m[239]&~m[240]&m[254])|(~m[237]&m[238]&m[239]&~m[240]&m[254])|(m[237]&m[238]&m[239]&~m[240]&m[254])|(m[237]&m[238]&m[239]&m[240]&m[254]));
    m[246] = (((m[242]&~m[243]&~m[244]&~m[245]&~m[259])|(~m[242]&m[243]&~m[244]&~m[245]&~m[259])|(~m[242]&~m[243]&m[244]&~m[245]&~m[259])|(m[242]&m[243]&~m[244]&m[245]&~m[259])|(m[242]&~m[243]&m[244]&m[245]&~m[259])|(~m[242]&m[243]&m[244]&m[245]&~m[259]))&BiasedRNG[153])|(((m[242]&~m[243]&~m[244]&~m[245]&m[259])|(~m[242]&m[243]&~m[244]&~m[245]&m[259])|(~m[242]&~m[243]&m[244]&~m[245]&m[259])|(m[242]&m[243]&~m[244]&m[245]&m[259])|(m[242]&~m[243]&m[244]&m[245]&m[259])|(~m[242]&m[243]&m[244]&m[245]&m[259]))&~BiasedRNG[153])|((m[242]&m[243]&~m[244]&~m[245]&~m[259])|(m[242]&~m[243]&m[244]&~m[245]&~m[259])|(~m[242]&m[243]&m[244]&~m[245]&~m[259])|(m[242]&m[243]&m[244]&~m[245]&~m[259])|(m[242]&m[243]&m[244]&m[245]&~m[259])|(m[242]&m[243]&~m[244]&~m[245]&m[259])|(m[242]&~m[243]&m[244]&~m[245]&m[259])|(~m[242]&m[243]&m[244]&~m[245]&m[259])|(m[242]&m[243]&m[244]&~m[245]&m[259])|(m[242]&m[243]&m[244]&m[245]&m[259]));
    m[251] = (((m[247]&~m[248]&~m[249]&~m[250]&~m[264])|(~m[247]&m[248]&~m[249]&~m[250]&~m[264])|(~m[247]&~m[248]&m[249]&~m[250]&~m[264])|(m[247]&m[248]&~m[249]&m[250]&~m[264])|(m[247]&~m[248]&m[249]&m[250]&~m[264])|(~m[247]&m[248]&m[249]&m[250]&~m[264]))&BiasedRNG[154])|(((m[247]&~m[248]&~m[249]&~m[250]&m[264])|(~m[247]&m[248]&~m[249]&~m[250]&m[264])|(~m[247]&~m[248]&m[249]&~m[250]&m[264])|(m[247]&m[248]&~m[249]&m[250]&m[264])|(m[247]&~m[248]&m[249]&m[250]&m[264])|(~m[247]&m[248]&m[249]&m[250]&m[264]))&~BiasedRNG[154])|((m[247]&m[248]&~m[249]&~m[250]&~m[264])|(m[247]&~m[248]&m[249]&~m[250]&~m[264])|(~m[247]&m[248]&m[249]&~m[250]&~m[264])|(m[247]&m[248]&m[249]&~m[250]&~m[264])|(m[247]&m[248]&m[249]&m[250]&~m[264])|(m[247]&m[248]&~m[249]&~m[250]&m[264])|(m[247]&~m[248]&m[249]&~m[250]&m[264])|(~m[247]&m[248]&m[249]&~m[250]&m[264])|(m[247]&m[248]&m[249]&~m[250]&m[264])|(m[247]&m[248]&m[249]&m[250]&m[264]));
    m[256] = (((m[252]&~m[253]&~m[254]&~m[255]&~m[267])|(~m[252]&m[253]&~m[254]&~m[255]&~m[267])|(~m[252]&~m[253]&m[254]&~m[255]&~m[267])|(m[252]&m[253]&~m[254]&m[255]&~m[267])|(m[252]&~m[253]&m[254]&m[255]&~m[267])|(~m[252]&m[253]&m[254]&m[255]&~m[267]))&BiasedRNG[155])|(((m[252]&~m[253]&~m[254]&~m[255]&m[267])|(~m[252]&m[253]&~m[254]&~m[255]&m[267])|(~m[252]&~m[253]&m[254]&~m[255]&m[267])|(m[252]&m[253]&~m[254]&m[255]&m[267])|(m[252]&~m[253]&m[254]&m[255]&m[267])|(~m[252]&m[253]&m[254]&m[255]&m[267]))&~BiasedRNG[155])|((m[252]&m[253]&~m[254]&~m[255]&~m[267])|(m[252]&~m[253]&m[254]&~m[255]&~m[267])|(~m[252]&m[253]&m[254]&~m[255]&~m[267])|(m[252]&m[253]&m[254]&~m[255]&~m[267])|(m[252]&m[253]&m[254]&m[255]&~m[267])|(m[252]&m[253]&~m[254]&~m[255]&m[267])|(m[252]&~m[253]&m[254]&~m[255]&m[267])|(~m[252]&m[253]&m[254]&~m[255]&m[267])|(m[252]&m[253]&m[254]&~m[255]&m[267])|(m[252]&m[253]&m[254]&m[255]&m[267]));
    m[261] = (((m[257]&~m[258]&~m[259]&~m[260]&~m[269])|(~m[257]&m[258]&~m[259]&~m[260]&~m[269])|(~m[257]&~m[258]&m[259]&~m[260]&~m[269])|(m[257]&m[258]&~m[259]&m[260]&~m[269])|(m[257]&~m[258]&m[259]&m[260]&~m[269])|(~m[257]&m[258]&m[259]&m[260]&~m[269]))&BiasedRNG[156])|(((m[257]&~m[258]&~m[259]&~m[260]&m[269])|(~m[257]&m[258]&~m[259]&~m[260]&m[269])|(~m[257]&~m[258]&m[259]&~m[260]&m[269])|(m[257]&m[258]&~m[259]&m[260]&m[269])|(m[257]&~m[258]&m[259]&m[260]&m[269])|(~m[257]&m[258]&m[259]&m[260]&m[269]))&~BiasedRNG[156])|((m[257]&m[258]&~m[259]&~m[260]&~m[269])|(m[257]&~m[258]&m[259]&~m[260]&~m[269])|(~m[257]&m[258]&m[259]&~m[260]&~m[269])|(m[257]&m[258]&m[259]&~m[260]&~m[269])|(m[257]&m[258]&m[259]&m[260]&~m[269])|(m[257]&m[258]&~m[259]&~m[260]&m[269])|(m[257]&~m[258]&m[259]&~m[260]&m[269])|(~m[257]&m[258]&m[259]&~m[260]&m[269])|(m[257]&m[258]&m[259]&~m[260]&m[269])|(m[257]&m[258]&m[259]&m[260]&m[269]));
    m[266] = (((m[262]&~m[263]&~m[264]&~m[265]&~m[274])|(~m[262]&m[263]&~m[264]&~m[265]&~m[274])|(~m[262]&~m[263]&m[264]&~m[265]&~m[274])|(m[262]&m[263]&~m[264]&m[265]&~m[274])|(m[262]&~m[263]&m[264]&m[265]&~m[274])|(~m[262]&m[263]&m[264]&m[265]&~m[274]))&BiasedRNG[157])|(((m[262]&~m[263]&~m[264]&~m[265]&m[274])|(~m[262]&m[263]&~m[264]&~m[265]&m[274])|(~m[262]&~m[263]&m[264]&~m[265]&m[274])|(m[262]&m[263]&~m[264]&m[265]&m[274])|(m[262]&~m[263]&m[264]&m[265]&m[274])|(~m[262]&m[263]&m[264]&m[265]&m[274]))&~BiasedRNG[157])|((m[262]&m[263]&~m[264]&~m[265]&~m[274])|(m[262]&~m[263]&m[264]&~m[265]&~m[274])|(~m[262]&m[263]&m[264]&~m[265]&~m[274])|(m[262]&m[263]&m[264]&~m[265]&~m[274])|(m[262]&m[263]&m[264]&m[265]&~m[274])|(m[262]&m[263]&~m[264]&~m[265]&m[274])|(m[262]&~m[263]&m[264]&~m[265]&m[274])|(~m[262]&m[263]&m[264]&~m[265]&m[274])|(m[262]&m[263]&m[264]&~m[265]&m[274])|(m[262]&m[263]&m[264]&m[265]&m[274]));
    m[271] = (((m[267]&~m[268]&~m[269]&~m[270]&~m[277])|(~m[267]&m[268]&~m[269]&~m[270]&~m[277])|(~m[267]&~m[268]&m[269]&~m[270]&~m[277])|(m[267]&m[268]&~m[269]&m[270]&~m[277])|(m[267]&~m[268]&m[269]&m[270]&~m[277])|(~m[267]&m[268]&m[269]&m[270]&~m[277]))&BiasedRNG[158])|(((m[267]&~m[268]&~m[269]&~m[270]&m[277])|(~m[267]&m[268]&~m[269]&~m[270]&m[277])|(~m[267]&~m[268]&m[269]&~m[270]&m[277])|(m[267]&m[268]&~m[269]&m[270]&m[277])|(m[267]&~m[268]&m[269]&m[270]&m[277])|(~m[267]&m[268]&m[269]&m[270]&m[277]))&~BiasedRNG[158])|((m[267]&m[268]&~m[269]&~m[270]&~m[277])|(m[267]&~m[268]&m[269]&~m[270]&~m[277])|(~m[267]&m[268]&m[269]&~m[270]&~m[277])|(m[267]&m[268]&m[269]&~m[270]&~m[277])|(m[267]&m[268]&m[269]&m[270]&~m[277])|(m[267]&m[268]&~m[269]&~m[270]&m[277])|(m[267]&~m[268]&m[269]&~m[270]&m[277])|(~m[267]&m[268]&m[269]&~m[270]&m[277])|(m[267]&m[268]&m[269]&~m[270]&m[277])|(m[267]&m[268]&m[269]&m[270]&m[277]));
    m[276] = (((m[272]&~m[273]&~m[274]&~m[275]&~m[279])|(~m[272]&m[273]&~m[274]&~m[275]&~m[279])|(~m[272]&~m[273]&m[274]&~m[275]&~m[279])|(m[272]&m[273]&~m[274]&m[275]&~m[279])|(m[272]&~m[273]&m[274]&m[275]&~m[279])|(~m[272]&m[273]&m[274]&m[275]&~m[279]))&BiasedRNG[159])|(((m[272]&~m[273]&~m[274]&~m[275]&m[279])|(~m[272]&m[273]&~m[274]&~m[275]&m[279])|(~m[272]&~m[273]&m[274]&~m[275]&m[279])|(m[272]&m[273]&~m[274]&m[275]&m[279])|(m[272]&~m[273]&m[274]&m[275]&m[279])|(~m[272]&m[273]&m[274]&m[275]&m[279]))&~BiasedRNG[159])|((m[272]&m[273]&~m[274]&~m[275]&~m[279])|(m[272]&~m[273]&m[274]&~m[275]&~m[279])|(~m[272]&m[273]&m[274]&~m[275]&~m[279])|(m[272]&m[273]&m[274]&~m[275]&~m[279])|(m[272]&m[273]&m[274]&m[275]&~m[279])|(m[272]&m[273]&~m[274]&~m[275]&m[279])|(m[272]&~m[273]&m[274]&~m[275]&m[279])|(~m[272]&m[273]&m[274]&~m[275]&m[279])|(m[272]&m[273]&m[274]&~m[275]&m[279])|(m[272]&m[273]&m[274]&m[275]&m[279]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[100]&LFSRcolor0[77]&LFSRcolor0[195]&LFSRcolor0[123]);
    BiasedRNG[1] = (LFSRcolor0[54]&LFSRcolor0[150]&LFSRcolor0[16]&LFSRcolor0[119]);
    BiasedRNG[2] = (LFSRcolor0[220]&LFSRcolor0[223]&LFSRcolor0[226]&LFSRcolor0[126]);
    BiasedRNG[3] = (LFSRcolor0[189]&LFSRcolor0[227]&LFSRcolor0[83]&LFSRcolor0[107]);
    BiasedRNG[4] = (LFSRcolor0[94]&LFSRcolor0[0]&LFSRcolor0[229]&LFSRcolor0[72]);
    BiasedRNG[5] = (LFSRcolor0[22]&LFSRcolor0[86]&LFSRcolor0[180]&LFSRcolor0[112]);
    BiasedRNG[6] = (LFSRcolor0[157]&LFSRcolor0[103]&LFSRcolor0[127]&LFSRcolor0[146]);
    BiasedRNG[7] = (LFSRcolor0[89]&LFSRcolor0[202]&LFSRcolor0[166]&LFSRcolor0[183]);
    BiasedRNG[8] = (LFSRcolor0[164]&LFSRcolor0[49]&LFSRcolor0[40]&LFSRcolor0[169]);
    BiasedRNG[9] = (LFSRcolor0[163]&LFSRcolor0[25]&LFSRcolor0[196]&LFSRcolor0[9]);
    BiasedRNG[10] = (LFSRcolor0[44]&LFSRcolor0[214]&LFSRcolor0[186]&LFSRcolor0[70]);
    BiasedRNG[11] = (LFSRcolor0[219]&LFSRcolor0[47]&LFSRcolor0[133]&LFSRcolor0[97]);
    BiasedRNG[12] = (LFSRcolor0[52]&LFSRcolor0[24]&LFSRcolor0[41]&LFSRcolor0[34]);
    BiasedRNG[13] = (LFSRcolor0[177]&LFSRcolor0[68]&LFSRcolor0[7]&LFSRcolor0[198]);
    BiasedRNG[14] = (LFSRcolor0[206]&LFSRcolor0[228]&LFSRcolor0[147]&LFSRcolor0[57]);
    BiasedRNG[15] = (LFSRcolor0[185]&LFSRcolor0[170]&LFSRcolor0[73]&LFSRcolor0[79]);
    BiasedRNG[16] = (LFSRcolor0[4]&LFSRcolor0[74]&LFSRcolor0[55]&LFSRcolor0[28]);
    BiasedRNG[17] = (LFSRcolor0[218]&LFSRcolor0[209]&LFSRcolor0[207]&LFSRcolor0[144]);
    BiasedRNG[18] = (LFSRcolor0[225]&LFSRcolor0[155]&LFSRcolor0[101]&LFSRcolor0[36]);
    BiasedRNG[19] = (LFSRcolor0[125]&LFSRcolor0[29]&LFSRcolor0[20]&LFSRcolor0[203]);
    BiasedRNG[20] = (LFSRcolor0[33]&LFSRcolor0[201]&LFSRcolor0[182]&LFSRcolor0[176]);
    BiasedRNG[21] = (LFSRcolor0[131]&LFSRcolor0[106]&LFSRcolor0[187]&LFSRcolor0[161]);
    BiasedRNG[22] = (LFSRcolor0[224]&LFSRcolor0[14]&LFSRcolor0[15]&LFSRcolor0[95]);
    BiasedRNG[23] = (LFSRcolor0[140]&LFSRcolor0[158]&LFSRcolor0[204]&LFSRcolor0[118]);
    BiasedRNG[24] = (LFSRcolor0[60]&LFSRcolor0[173]&LFSRcolor0[152]&LFSRcolor0[137]);
    BiasedRNG[25] = (LFSRcolor0[62]&LFSRcolor0[138]&LFSRcolor0[134]&LFSRcolor0[154]);
    BiasedRNG[26] = (LFSRcolor0[165]&LFSRcolor0[102]&LFSRcolor0[21]&LFSRcolor0[67]);
    BiasedRNG[27] = (LFSRcolor0[171]&LFSRcolor0[8]&LFSRcolor0[213]&LFSRcolor0[193]);
    BiasedRNG[28] = (LFSRcolor0[181]&LFSRcolor0[75]&LFSRcolor0[87]&LFSRcolor0[114]);
    BiasedRNG[29] = (LFSRcolor0[160]&LFSRcolor0[58]&LFSRcolor0[184]&LFSRcolor0[12]);
    BiasedRNG[30] = (LFSRcolor0[1]&LFSRcolor0[132]&LFSRcolor0[135]&LFSRcolor0[190]);
    BiasedRNG[31] = (LFSRcolor0[145]&LFSRcolor0[85]&LFSRcolor0[26]&LFSRcolor0[63]);
    BiasedRNG[32] = (LFSRcolor0[13]&LFSRcolor0[64]&LFSRcolor0[156]&LFSRcolor0[98]);
    BiasedRNG[33] = (LFSRcolor0[172]&LFSRcolor0[116]&LFSRcolor0[136]&LFSRcolor0[148]);
    BiasedRNG[34] = (LFSRcolor0[215]&LFSRcolor0[222]&LFSRcolor0[168]&LFSRcolor0[82]);
    BiasedRNG[35] = (LFSRcolor0[38]&LFSRcolor0[211]&LFSRcolor0[197]&LFSRcolor0[121]);
    BiasedRNG[36] = (LFSRcolor0[110]&LFSRcolor0[93]&LFSRcolor0[2]&LFSRcolor0[5]);
    BiasedRNG[37] = (LFSRcolor0[42]&LFSRcolor0[53]&LFSRcolor0[96]&LFSRcolor0[65]);
    BiasedRNG[38] = (LFSRcolor0[80]&LFSRcolor0[105]&LFSRcolor0[124]&LFSRcolor0[84]);
    BiasedRNG[39] = (LFSRcolor0[167]&LFSRcolor0[30]&LFSRcolor0[23]&LFSRcolor0[192]);
    BiasedRNG[40] = (LFSRcolor0[162]&LFSRcolor0[17]&LFSRcolor0[130]&LFSRcolor0[71]);
    BiasedRNG[41] = (LFSRcolor0[179]&LFSRcolor0[191]&LFSRcolor0[81]&LFSRcolor0[27]);
    BiasedRNG[42] = (LFSRcolor0[217]&LFSRcolor0[32]&LFSRcolor0[128]&LFSRcolor0[142]);
    BiasedRNG[43] = (LFSRcolor0[141]&LFSRcolor0[149]&LFSRcolor0[117]&LFSRcolor0[88]);
    BiasedRNG[44] = (LFSRcolor0[111]&LFSRcolor0[120]&LFSRcolor0[76]&LFSRcolor0[129]);
    BiasedRNG[45] = (LFSRcolor0[59]&LFSRcolor0[31]&LFSRcolor0[91]&LFSRcolor0[159]);
    BiasedRNG[46] = (LFSRcolor0[37]&LFSRcolor0[113]&LFSRcolor0[153]&LFSRcolor0[51]);
    UnbiasedRNG[0] = LFSRcolor0[210];
    UnbiasedRNG[1] = LFSRcolor0[10];
    UnbiasedRNG[2] = LFSRcolor0[19];
    UnbiasedRNG[3] = LFSRcolor0[115];
    UnbiasedRNG[4] = LFSRcolor0[39];
    UnbiasedRNG[5] = LFSRcolor0[175];
    UnbiasedRNG[6] = LFSRcolor0[56];
    UnbiasedRNG[7] = LFSRcolor0[208];
    UnbiasedRNG[8] = LFSRcolor0[48];
    UnbiasedRNG[9] = LFSRcolor0[61];
    UnbiasedRNG[10] = LFSRcolor0[104];
    UnbiasedRNG[11] = LFSRcolor0[109];
    UnbiasedRNG[12] = LFSRcolor0[92];
    UnbiasedRNG[13] = LFSRcolor0[35];
    UnbiasedRNG[14] = LFSRcolor0[66];
    UnbiasedRNG[15] = LFSRcolor0[11];
    UnbiasedRNG[16] = LFSRcolor0[188];
    UnbiasedRNG[17] = LFSRcolor0[221];
    UnbiasedRNG[18] = LFSRcolor0[205];
    UnbiasedRNG[19] = LFSRcolor0[194];
    UnbiasedRNG[20] = LFSRcolor0[151];
    UnbiasedRNG[21] = LFSRcolor0[212];
    UnbiasedRNG[22] = LFSRcolor0[143];
    UnbiasedRNG[23] = LFSRcolor0[45];
    UnbiasedRNG[24] = LFSRcolor0[178];
    UnbiasedRNG[25] = LFSRcolor0[216];
    UnbiasedRNG[26] = LFSRcolor0[43];
    UnbiasedRNG[27] = LFSRcolor0[199];
end

always @(posedge color0_clk) begin
    BiasedRNG[47] = (LFSRcolor1[197]&LFSRcolor1[201]&LFSRcolor1[76]&LFSRcolor1[103]);
    BiasedRNG[48] = (LFSRcolor1[19]&LFSRcolor1[3]&LFSRcolor1[162]&LFSRcolor1[193]);
    BiasedRNG[49] = (LFSRcolor1[149]&LFSRcolor1[57]&LFSRcolor1[111]&LFSRcolor1[188]);
    BiasedRNG[50] = (LFSRcolor1[35]&LFSRcolor1[228]&LFSRcolor1[10]&LFSRcolor1[26]);
    BiasedRNG[51] = (LFSRcolor1[71]&LFSRcolor1[28]&LFSRcolor1[166]&LFSRcolor1[150]);
    BiasedRNG[52] = (LFSRcolor1[80]&LFSRcolor1[94]&LFSRcolor1[47]&LFSRcolor1[181]);
    BiasedRNG[53] = (LFSRcolor1[114]&LFSRcolor1[93]&LFSRcolor1[189]&LFSRcolor1[78]);
    BiasedRNG[54] = (LFSRcolor1[209]&LFSRcolor1[116]&LFSRcolor1[216]&LFSRcolor1[92]);
    BiasedRNG[55] = (LFSRcolor1[0]&LFSRcolor1[32]&LFSRcolor1[63]&LFSRcolor1[7]);
    BiasedRNG[56] = (LFSRcolor1[64]&LFSRcolor1[65]&LFSRcolor1[185]&LFSRcolor1[203]);
    BiasedRNG[57] = (LFSRcolor1[138]&LFSRcolor1[139]&LFSRcolor1[213]&LFSRcolor1[70]);
    BiasedRNG[58] = (LFSRcolor1[74]&LFSRcolor1[42]&LFSRcolor1[210]&LFSRcolor1[115]);
    BiasedRNG[59] = (LFSRcolor1[202]&LFSRcolor1[58]&LFSRcolor1[50]&LFSRcolor1[153]);
    BiasedRNG[60] = (LFSRcolor1[164]&LFSRcolor1[100]&LFSRcolor1[88]&LFSRcolor1[204]);
    BiasedRNG[61] = (LFSRcolor1[37]&LFSRcolor1[211]&LFSRcolor1[99]&LFSRcolor1[128]);
    BiasedRNG[62] = (LFSRcolor1[220]&LFSRcolor1[91]&LFSRcolor1[134]&LFSRcolor1[196]);
    BiasedRNG[63] = (LFSRcolor1[159]&LFSRcolor1[120]&LFSRcolor1[27]&LFSRcolor1[172]);
    BiasedRNG[64] = (LFSRcolor1[77]&LFSRcolor1[182]&LFSRcolor1[148]&LFSRcolor1[158]);
    BiasedRNG[65] = (LFSRcolor1[133]&LFSRcolor1[137]&LFSRcolor1[72]&LFSRcolor1[156]);
    BiasedRNG[66] = (LFSRcolor1[68]&LFSRcolor1[96]&LFSRcolor1[67]&LFSRcolor1[180]);
    BiasedRNG[67] = (LFSRcolor1[85]&LFSRcolor1[25]&LFSRcolor1[143]&LFSRcolor1[60]);
    BiasedRNG[68] = (LFSRcolor1[1]&LFSRcolor1[105]&LFSRcolor1[176]&LFSRcolor1[110]);
    BiasedRNG[69] = (LFSRcolor1[229]&LFSRcolor1[223]&LFSRcolor1[39]&LFSRcolor1[227]);
    BiasedRNG[70] = (LFSRcolor1[132]&LFSRcolor1[84]&LFSRcolor1[140]&LFSRcolor1[146]);
    BiasedRNG[71] = (LFSRcolor1[121]&LFSRcolor1[89]&LFSRcolor1[36]&LFSRcolor1[2]);
    BiasedRNG[72] = (LFSRcolor1[151]&LFSRcolor1[160]&LFSRcolor1[199]&LFSRcolor1[127]);
    BiasedRNG[73] = (LFSRcolor1[31]&LFSRcolor1[11]&LFSRcolor1[14]&LFSRcolor1[200]);
    BiasedRNG[74] = (LFSRcolor1[48]&LFSRcolor1[55]&LFSRcolor1[101]&LFSRcolor1[45]);
    BiasedRNG[75] = (LFSRcolor1[23]&LFSRcolor1[119]&LFSRcolor1[215]&LFSRcolor1[41]);
    BiasedRNG[76] = (LFSRcolor1[191]&LFSRcolor1[218]&LFSRcolor1[117]&LFSRcolor1[161]);
    BiasedRNG[77] = (LFSRcolor1[107]&LFSRcolor1[174]&LFSRcolor1[56]&LFSRcolor1[187]);
    BiasedRNG[78] = (LFSRcolor1[147]&LFSRcolor1[167]&LFSRcolor1[18]&LFSRcolor1[212]);
    BiasedRNG[79] = (LFSRcolor1[219]&LFSRcolor1[214]&LFSRcolor1[198]&LFSRcolor1[20]);
    BiasedRNG[80] = (LFSRcolor1[113]&LFSRcolor1[168]&LFSRcolor1[123]&LFSRcolor1[24]);
    BiasedRNG[81] = (LFSRcolor1[224]&LFSRcolor1[186]&LFSRcolor1[142]&LFSRcolor1[124]);
    BiasedRNG[82] = (LFSRcolor1[97]&LFSRcolor1[9]&LFSRcolor1[15]&LFSRcolor1[87]);
    BiasedRNG[83] = (LFSRcolor1[62]&LFSRcolor1[192]&LFSRcolor1[169]&LFSRcolor1[125]);
    BiasedRNG[84] = (LFSRcolor1[118]&LFSRcolor1[90]&LFSRcolor1[83]&LFSRcolor1[129]);
    BiasedRNG[85] = (LFSRcolor1[205]&LFSRcolor1[184]&LFSRcolor1[183]&LFSRcolor1[190]);
    BiasedRNG[86] = (LFSRcolor1[217]&LFSRcolor1[178]&LFSRcolor1[75]&LFSRcolor1[173]);
    BiasedRNG[87] = (LFSRcolor1[112]&LFSRcolor1[21]&LFSRcolor1[6]&LFSRcolor1[221]);
    BiasedRNG[88] = (LFSRcolor1[122]&LFSRcolor1[12]&LFSRcolor1[222]&LFSRcolor1[38]);
    BiasedRNG[89] = (LFSRcolor1[86]&LFSRcolor1[126]&LFSRcolor1[82]&LFSRcolor1[108]);
    BiasedRNG[90] = (LFSRcolor1[177]&LFSRcolor1[157]&LFSRcolor1[17]&LFSRcolor1[33]);
    BiasedRNG[91] = (LFSRcolor1[59]&LFSRcolor1[66]&LFSRcolor1[44]&LFSRcolor1[30]);
    BiasedRNG[92] = (LFSRcolor1[152]&LFSRcolor1[95]&LFSRcolor1[51]&LFSRcolor1[175]);
    BiasedRNG[93] = (LFSRcolor1[16]&LFSRcolor1[61]&LFSRcolor1[145]&LFSRcolor1[102]);
    BiasedRNG[94] = (LFSRcolor1[13]&LFSRcolor1[226]&LFSRcolor1[4]&LFSRcolor1[170]);
    UnbiasedRNG[28] = LFSRcolor1[43];
    UnbiasedRNG[29] = LFSRcolor1[104];
    UnbiasedRNG[30] = LFSRcolor1[144];
    UnbiasedRNG[31] = LFSRcolor1[154];
    UnbiasedRNG[32] = LFSRcolor1[22];
    UnbiasedRNG[33] = LFSRcolor1[208];
    UnbiasedRNG[34] = LFSRcolor1[40];
    UnbiasedRNG[35] = LFSRcolor1[136];
    UnbiasedRNG[36] = LFSRcolor1[49];
    UnbiasedRNG[37] = LFSRcolor1[5];
    UnbiasedRNG[38] = LFSRcolor1[165];
    UnbiasedRNG[39] = LFSRcolor1[163];
    UnbiasedRNG[40] = LFSRcolor1[131];
    UnbiasedRNG[41] = LFSRcolor1[8];
    UnbiasedRNG[42] = LFSRcolor1[179];
    UnbiasedRNG[43] = LFSRcolor1[141];
    UnbiasedRNG[44] = LFSRcolor1[135];
    UnbiasedRNG[45] = LFSRcolor1[54];
    UnbiasedRNG[46] = LFSRcolor1[46];
    UnbiasedRNG[47] = LFSRcolor1[171];
    UnbiasedRNG[48] = LFSRcolor1[79];
    UnbiasedRNG[49] = LFSRcolor1[207];
    UnbiasedRNG[50] = LFSRcolor1[109];
    UnbiasedRNG[51] = LFSRcolor1[69];
    UnbiasedRNG[52] = LFSRcolor1[130];
    UnbiasedRNG[53] = LFSRcolor1[155];
    UnbiasedRNG[54] = LFSRcolor1[106];
    UnbiasedRNG[55] = LFSRcolor1[73];
    UnbiasedRNG[56] = LFSRcolor1[195];
    UnbiasedRNG[57] = LFSRcolor1[206];
end

always @(posedge color1_clk) begin
    BiasedRNG[95] = (LFSRcolor2[18]&LFSRcolor2[177]&LFSRcolor2[170]&LFSRcolor2[12]);
    BiasedRNG[96] = (LFSRcolor2[72]&LFSRcolor2[8]&LFSRcolor2[57]&LFSRcolor2[59]);
    BiasedRNG[97] = (LFSRcolor2[73]&LFSRcolor2[142]&LFSRcolor2[100]&LFSRcolor2[19]);
    BiasedRNG[98] = (LFSRcolor2[125]&LFSRcolor2[7]&LFSRcolor2[115]&LFSRcolor2[69]);
    BiasedRNG[99] = (LFSRcolor2[124]&LFSRcolor2[37]&LFSRcolor2[151]&LFSRcolor2[26]);
    BiasedRNG[100] = (LFSRcolor2[3]&LFSRcolor2[76]&LFSRcolor2[153]&LFSRcolor2[121]);
    BiasedRNG[101] = (LFSRcolor2[60]&LFSRcolor2[134]&LFSRcolor2[65]&LFSRcolor2[145]);
    BiasedRNG[102] = (LFSRcolor2[93]&LFSRcolor2[77]&LFSRcolor2[67]&LFSRcolor2[181]);
    BiasedRNG[103] = (LFSRcolor2[123]&LFSRcolor2[103]&LFSRcolor2[2]&LFSRcolor2[111]);
    BiasedRNG[104] = (LFSRcolor2[54]&LFSRcolor2[140]&LFSRcolor2[45]&LFSRcolor2[135]);
    BiasedRNG[105] = (LFSRcolor2[71]&LFSRcolor2[35]&LFSRcolor2[162]&LFSRcolor2[127]);
    BiasedRNG[106] = (LFSRcolor2[97]&LFSRcolor2[156]&LFSRcolor2[139]&LFSRcolor2[126]);
    BiasedRNG[107] = (LFSRcolor2[152]&LFSRcolor2[83]&LFSRcolor2[17]&LFSRcolor2[74]);
    BiasedRNG[108] = (LFSRcolor2[183]&LFSRcolor2[44]&LFSRcolor2[41]&LFSRcolor2[53]);
    BiasedRNG[109] = (LFSRcolor2[165]&LFSRcolor2[95]&LFSRcolor2[82]&LFSRcolor2[149]);
    BiasedRNG[110] = (LFSRcolor2[89]&LFSRcolor2[128]&LFSRcolor2[174]&LFSRcolor2[30]);
    BiasedRNG[111] = (LFSRcolor2[113]&LFSRcolor2[179]&LFSRcolor2[175]&LFSRcolor2[90]);
    BiasedRNG[112] = (LFSRcolor2[64]&LFSRcolor2[40]&LFSRcolor2[51]&LFSRcolor2[178]);
    BiasedRNG[113] = (LFSRcolor2[105]&LFSRcolor2[86]&LFSRcolor2[46]&LFSRcolor2[104]);
    BiasedRNG[114] = (LFSRcolor2[0]&LFSRcolor2[48]&LFSRcolor2[91]&LFSRcolor2[87]);
    BiasedRNG[115] = (LFSRcolor2[137]&LFSRcolor2[148]&LFSRcolor2[122]&LFSRcolor2[21]);
    BiasedRNG[116] = (LFSRcolor2[49]&LFSRcolor2[85]&LFSRcolor2[11]&LFSRcolor2[42]);
    BiasedRNG[117] = (LFSRcolor2[101]&LFSRcolor2[78]&LFSRcolor2[180]&LFSRcolor2[22]);
    BiasedRNG[118] = (LFSRcolor2[68]&LFSRcolor2[38]&LFSRcolor2[171]&LFSRcolor2[52]);
    BiasedRNG[119] = (LFSRcolor2[79]&LFSRcolor2[15]&LFSRcolor2[4]&LFSRcolor2[130]);
    BiasedRNG[120] = (LFSRcolor2[169]&LFSRcolor2[157]&LFSRcolor2[144]&LFSRcolor2[147]);
    BiasedRNG[121] = (LFSRcolor2[55]&LFSRcolor2[47]&LFSRcolor2[80]&LFSRcolor2[5]);
    BiasedRNG[122] = (LFSRcolor2[150]&LFSRcolor2[176]&LFSRcolor2[159]&LFSRcolor2[61]);
    BiasedRNG[123] = (LFSRcolor2[96]&LFSRcolor2[120]&LFSRcolor2[102]&LFSRcolor2[164]);
    BiasedRNG[124] = (LFSRcolor2[161]&LFSRcolor2[6]&LFSRcolor2[143]&LFSRcolor2[24]);
    BiasedRNG[125] = (LFSRcolor2[88]&LFSRcolor2[62]&LFSRcolor2[13]&LFSRcolor2[70]);
    BiasedRNG[126] = (LFSRcolor2[114]&LFSRcolor2[39]&LFSRcolor2[154]&LFSRcolor2[167]);
    BiasedRNG[127] = (LFSRcolor2[158]&LFSRcolor2[10]&LFSRcolor2[138]&LFSRcolor2[14]);
    BiasedRNG[128] = (LFSRcolor2[50]&LFSRcolor2[56]&LFSRcolor2[146]&LFSRcolor2[29]);
    BiasedRNG[129] = (LFSRcolor2[108]&LFSRcolor2[116]&LFSRcolor2[25]&LFSRcolor2[43]);
    BiasedRNG[130] = (LFSRcolor2[163]&LFSRcolor2[9]&LFSRcolor2[166]&LFSRcolor2[28]);
    UnbiasedRNG[58] = LFSRcolor2[99];
    UnbiasedRNG[59] = LFSRcolor2[27];
    UnbiasedRNG[60] = LFSRcolor2[20];
    UnbiasedRNG[61] = LFSRcolor2[112];
    UnbiasedRNG[62] = LFSRcolor2[106];
    UnbiasedRNG[63] = LFSRcolor2[107];
    UnbiasedRNG[64] = LFSRcolor2[132];
    UnbiasedRNG[65] = LFSRcolor2[133];
    UnbiasedRNG[66] = LFSRcolor2[84];
    UnbiasedRNG[67] = LFSRcolor2[173];
    UnbiasedRNG[68] = LFSRcolor2[98];
    UnbiasedRNG[69] = LFSRcolor2[131];
    UnbiasedRNG[70] = LFSRcolor2[136];
    UnbiasedRNG[71] = LFSRcolor2[75];
    UnbiasedRNG[72] = LFSRcolor2[92];
    UnbiasedRNG[73] = LFSRcolor2[110];
    UnbiasedRNG[74] = LFSRcolor2[118];
    UnbiasedRNG[75] = LFSRcolor2[172];
    UnbiasedRNG[76] = LFSRcolor2[58];
    UnbiasedRNG[77] = LFSRcolor2[31];
    UnbiasedRNG[78] = LFSRcolor2[141];
    UnbiasedRNG[79] = LFSRcolor2[16];
    UnbiasedRNG[80] = LFSRcolor2[32];
    UnbiasedRNG[81] = LFSRcolor2[1];
    UnbiasedRNG[82] = LFSRcolor2[94];
    UnbiasedRNG[83] = LFSRcolor2[33];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[84] = LFSRcolor3[29];
    UnbiasedRNG[85] = LFSRcolor3[39];
    UnbiasedRNG[86] = LFSRcolor3[21];
    UnbiasedRNG[87] = LFSRcolor3[9];
    UnbiasedRNG[88] = LFSRcolor3[32];
    UnbiasedRNG[89] = LFSRcolor3[25];
    UnbiasedRNG[90] = LFSRcolor3[33];
    UnbiasedRNG[91] = LFSRcolor3[40];
    UnbiasedRNG[92] = LFSRcolor3[20];
    UnbiasedRNG[93] = LFSRcolor3[44];
    UnbiasedRNG[94] = LFSRcolor3[4];
    UnbiasedRNG[95] = LFSRcolor3[35];
    UnbiasedRNG[96] = LFSRcolor3[11];
    UnbiasedRNG[97] = LFSRcolor3[27];
    UnbiasedRNG[98] = LFSRcolor3[16];
    UnbiasedRNG[99] = LFSRcolor3[30];
    UnbiasedRNG[100] = LFSRcolor3[6];
    UnbiasedRNG[101] = LFSRcolor3[7];
    UnbiasedRNG[102] = LFSRcolor3[28];
    UnbiasedRNG[103] = LFSRcolor3[14];
end

always @(posedge color3_clk) begin
    BiasedRNG[131] = (LFSRcolor4[97]&LFSRcolor4[49]&LFSRcolor4[112]&LFSRcolor4[58]);
    BiasedRNG[132] = (LFSRcolor4[99]&LFSRcolor4[68]&LFSRcolor4[13]&LFSRcolor4[27]);
    BiasedRNG[133] = (LFSRcolor4[89]&LFSRcolor4[69]&LFSRcolor4[116]&LFSRcolor4[55]);
    BiasedRNG[134] = (LFSRcolor4[90]&LFSRcolor4[24]&LFSRcolor4[83]&LFSRcolor4[71]);
    BiasedRNG[135] = (LFSRcolor4[41]&LFSRcolor4[2]&LFSRcolor4[3]&LFSRcolor4[134]);
    BiasedRNG[136] = (LFSRcolor4[73]&LFSRcolor4[35]&LFSRcolor4[130]&LFSRcolor4[38]);
    BiasedRNG[137] = (LFSRcolor4[46]&LFSRcolor4[115]&LFSRcolor4[59]&LFSRcolor4[113]);
    BiasedRNG[138] = (LFSRcolor4[126]&LFSRcolor4[136]&LFSRcolor4[50]&LFSRcolor4[10]);
    BiasedRNG[139] = (LFSRcolor4[12]&LFSRcolor4[94]&LFSRcolor4[114]&LFSRcolor4[70]);
    BiasedRNG[140] = (LFSRcolor4[76]&LFSRcolor4[78]&LFSRcolor4[119]&LFSRcolor4[45]);
    BiasedRNG[141] = (LFSRcolor4[100]&LFSRcolor4[108]&LFSRcolor4[4]&LFSRcolor4[104]);
    BiasedRNG[142] = (LFSRcolor4[37]&LFSRcolor4[77]&LFSRcolor4[51]&LFSRcolor4[42]);
    BiasedRNG[143] = (LFSRcolor4[127]&LFSRcolor4[96]&LFSRcolor4[102]&LFSRcolor4[137]);
    BiasedRNG[144] = (LFSRcolor4[84]&LFSRcolor4[54]&LFSRcolor4[91]&LFSRcolor4[1]);
    BiasedRNG[145] = (LFSRcolor4[43]&LFSRcolor4[105]&LFSRcolor4[56]&LFSRcolor4[87]);
    BiasedRNG[146] = (LFSRcolor4[61]&LFSRcolor4[6]&LFSRcolor4[19]&LFSRcolor4[85]);
    BiasedRNG[147] = (LFSRcolor4[120]&LFSRcolor4[103]&LFSRcolor4[32]&LFSRcolor4[53]);
    BiasedRNG[148] = (LFSRcolor4[133]&LFSRcolor4[135]&LFSRcolor4[93]&LFSRcolor4[66]);
    BiasedRNG[149] = (LFSRcolor4[98]&LFSRcolor4[65]&LFSRcolor4[122]&LFSRcolor4[86]);
    BiasedRNG[150] = (LFSRcolor4[79]&LFSRcolor4[101]&LFSRcolor4[22]&LFSRcolor4[26]);
    BiasedRNG[151] = (LFSRcolor4[106]&LFSRcolor4[11]&LFSRcolor4[132]&LFSRcolor4[131]);
    BiasedRNG[152] = (LFSRcolor4[20]&LFSRcolor4[111]&LFSRcolor4[40]&LFSRcolor4[30]);
    BiasedRNG[153] = (LFSRcolor4[9]&LFSRcolor4[123]&LFSRcolor4[57]&LFSRcolor4[15]);
    BiasedRNG[154] = (LFSRcolor4[47]&LFSRcolor4[72]&LFSRcolor4[7]&LFSRcolor4[14]);
    BiasedRNG[155] = (LFSRcolor4[18]&LFSRcolor4[28]&LFSRcolor4[75]&LFSRcolor4[31]);
    BiasedRNG[156] = (LFSRcolor4[17]&LFSRcolor4[125]&LFSRcolor4[80]&LFSRcolor4[34]);
    BiasedRNG[157] = (LFSRcolor4[121]&LFSRcolor4[82]&LFSRcolor4[60]&LFSRcolor4[23]);
    BiasedRNG[158] = (LFSRcolor4[128]&LFSRcolor4[88]&LFSRcolor4[107]&LFSRcolor4[67]);
    BiasedRNG[159] = (LFSRcolor4[16]&LFSRcolor4[5]&LFSRcolor4[29]&LFSRcolor4[8]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule