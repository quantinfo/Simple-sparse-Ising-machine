//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [31:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [1333:0] LFSRcolor0;
wire [1793:0] LFSRcolor1;
wire [1287:0] LFSRcolor2;
wire [229:0] LFSRcolor3;
wire [965:0] LFSRcolor4;
reg [1133:0] BiasedRNG;       //For I=+/-1 cases
reg [945:0] UnbiasedRNG;   //For I=0 cases
reg [0:2127] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[672] = 1'b1;
initial m[931] = 1'b0;
initial m[941] = 1'b0;
initial m[956] = 1'b0;
initial m[976] = 1'b1;
initial m[1001] = 1'b0;
initial m[1031] = 1'b1;
initial m[1066] = 1'b0;
initial m[1106] = 1'b1;
initial m[1151] = 1'b1;
initial m[1201] = 1'b0;
initial m[1256] = 1'b0;
initial m[1316] = 1'b0;
initial m[1381] = 1'b0;
initial m[1451] = 1'b1;
initial m[1526] = 1'b0;
initial m[1601] = 1'b1;
initial m[1671] = 1'b0;
initial m[1736] = 1'b0;
initial m[1796] = 1'b1;
initial m[1851] = 1'b1;
initial m[1901] = 1'b1;
initial m[1946] = 1'b0;
initial m[1986] = 1'b1;
initial m[2021] = 1'b1;
initial m[2051] = 1'b1;
initial m[2076] = 1'b0;
initial m[2096] = 1'b1;
initial m[2111] = 1'b0;
initial m[2121] = 1'b1;
initial m[2126] = 1'b1;
initial m[2127] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[930] = 1'b0;
initial m[940] = 1'b0;
initial m[955] = 1'b0;
initial m[975] = 1'b0;
initial m[1000] = 1'b0;
initial m[1030] = 1'b0;
initial m[1065] = 1'b0;
initial m[1105] = 1'b0;
initial m[1150] = 1'b0;
initial m[1200] = 1'b0;
initial m[1255] = 1'b0;
initial m[1315] = 1'b0;
initial m[1380] = 1'b0;
initial m[1450] = 1'b0;
initial m[1525] = 1'b0;
initial m[1528] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR0_11(.LFSRregister(LFSRcolor0[551:506]),.clk(sample_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR0_12(.LFSRregister(LFSRcolor0[597:552]),.clk(sample_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR0_13(.LFSRregister(LFSRcolor0[643:598]),.clk(sample_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR0_14(.LFSRregister(LFSRcolor0[689:644]),.clk(sample_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR0_15(.LFSRregister(LFSRcolor0[735:690]),.clk(sample_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR0_16(.LFSRregister(LFSRcolor0[781:736]),.clk(sample_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR0_17(.LFSRregister(LFSRcolor0[827:782]),.clk(sample_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR0_18(.LFSRregister(LFSRcolor0[873:828]),.clk(sample_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR0_19(.LFSRregister(LFSRcolor0[919:874]),.clk(sample_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR0_20(.LFSRregister(LFSRcolor0[965:920]),.clk(sample_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR0_21(.LFSRregister(LFSRcolor0[1011:966]),.clk(sample_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR0_22(.LFSRregister(LFSRcolor0[1057:1012]),.clk(sample_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR0_23(.LFSRregister(LFSRcolor0[1103:1058]),.clk(sample_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR0_24(.LFSRregister(LFSRcolor0[1149:1104]),.clk(sample_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR0_25(.LFSRregister(LFSRcolor0[1195:1150]),.clk(sample_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR0_26(.LFSRregister(LFSRcolor0[1241:1196]),.clk(sample_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR0_27(.LFSRregister(LFSRcolor0[1287:1242]),.clk(sample_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR0_28(.LFSRregister(LFSRcolor0[1333:1288]),.clk(sample_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR1_15(.LFSRregister(LFSRcolor1[735:690]),.clk(color0_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR1_16(.LFSRregister(LFSRcolor1[781:736]),.clk(color0_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR1_17(.LFSRregister(LFSRcolor1[827:782]),.clk(color0_clk));
lfsr #(.seed(46'b0011001000010001001111001110101111011111000110)) LFSR1_18(.LFSRregister(LFSRcolor1[873:828]),.clk(color0_clk));
lfsr #(.seed(46'b0101000110100000010101001000010000101101100110)) LFSR1_19(.LFSRregister(LFSRcolor1[919:874]),.clk(color0_clk));
lfsr #(.seed(46'b1110011010010011001010111010100101111111100000)) LFSR1_20(.LFSRregister(LFSRcolor1[965:920]),.clk(color0_clk));
lfsr #(.seed(46'b1001111000010100100001100010110000001111101011)) LFSR1_21(.LFSRregister(LFSRcolor1[1011:966]),.clk(color0_clk));
lfsr #(.seed(46'b0011101001111100110111000000010000101100111110)) LFSR1_22(.LFSRregister(LFSRcolor1[1057:1012]),.clk(color0_clk));
lfsr #(.seed(46'b1010111010001100001100010110010011100100101100)) LFSR1_23(.LFSRregister(LFSRcolor1[1103:1058]),.clk(color0_clk));
lfsr #(.seed(46'b1101010000110001000001011010110100010000110101)) LFSR1_24(.LFSRregister(LFSRcolor1[1149:1104]),.clk(color0_clk));
lfsr #(.seed(46'b0111111000001001010001100011001110110101101001)) LFSR1_25(.LFSRregister(LFSRcolor1[1195:1150]),.clk(color0_clk));
lfsr #(.seed(46'b0111011110101100100001111000001001111001010010)) LFSR1_26(.LFSRregister(LFSRcolor1[1241:1196]),.clk(color0_clk));
lfsr #(.seed(46'b0110010001011011111100000000110011011110000100)) LFSR1_27(.LFSRregister(LFSRcolor1[1287:1242]),.clk(color0_clk));
lfsr #(.seed(46'b1100101101001001110010011101110000001110111111)) LFSR1_28(.LFSRregister(LFSRcolor1[1333:1288]),.clk(color0_clk));
lfsr #(.seed(46'b1110010100000011100111110011000001001000000101)) LFSR1_29(.LFSRregister(LFSRcolor1[1379:1334]),.clk(color0_clk));
lfsr #(.seed(46'b1100111110111110000101110101010111111010101000)) LFSR1_30(.LFSRregister(LFSRcolor1[1425:1380]),.clk(color0_clk));
lfsr #(.seed(46'b1101101000110111001110111111011011100011111101)) LFSR1_31(.LFSRregister(LFSRcolor1[1471:1426]),.clk(color0_clk));
lfsr #(.seed(46'b1011100111101011110000001101111100001111100011)) LFSR1_32(.LFSRregister(LFSRcolor1[1517:1472]),.clk(color0_clk));
lfsr #(.seed(46'b1000011101010100110111010000000111000111010111)) LFSR1_33(.LFSRregister(LFSRcolor1[1563:1518]),.clk(color0_clk));
lfsr #(.seed(46'b0011001001101100101110110001011100100100110000)) LFSR1_34(.LFSRregister(LFSRcolor1[1609:1564]),.clk(color0_clk));
lfsr #(.seed(46'b0011110010011101000111111110100110110100101000)) LFSR1_35(.LFSRregister(LFSRcolor1[1655:1610]),.clk(color0_clk));
lfsr #(.seed(46'b1100000100011100010111001011000000101100110100)) LFSR1_36(.LFSRregister(LFSRcolor1[1701:1656]),.clk(color0_clk));
lfsr #(.seed(46'b1001101001101101001001111001110100110001100010)) LFSR1_37(.LFSRregister(LFSRcolor1[1747:1702]),.clk(color0_clk));
lfsr #(.seed(46'b1000000000001101011011010100000001101001001111)) LFSR1_38(.LFSRregister(LFSRcolor1[1793:1748]),.clk(color0_clk));
lfsr #(.seed(46'b1000011000100000010011100100110100001010000001)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0101000011110010010110011011111101010101011010)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0011111001110010110000110100101000000000100010)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0011101001110100101101111100101010101100110000)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1100111100001111010111011100011110001010110011)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0101101111111000101111101010111101100011110011)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1100101101101111100100111011110111010010100100)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b0110001110010011010100101010010010100100011000)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b0010101111101011001110100001110011000100001001)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b0100110100101000110001000110101010001110100101)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b1111010011010001011111110011011111011111011010)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b0011000010001101011100101011111101010001010111)) LFSR2_11(.LFSRregister(LFSRcolor2[551:506]),.clk(color1_clk));
lfsr #(.seed(46'b0011010011011000100111011100010000001110001110)) LFSR2_12(.LFSRregister(LFSRcolor2[597:552]),.clk(color1_clk));
lfsr #(.seed(46'b0010110000011111111111101000111101111100101000)) LFSR2_13(.LFSRregister(LFSRcolor2[643:598]),.clk(color1_clk));
lfsr #(.seed(46'b1110000110010010100110000110010000011111100110)) LFSR2_14(.LFSRregister(LFSRcolor2[689:644]),.clk(color1_clk));
lfsr #(.seed(46'b0011101100010010111110000100001011000110001101)) LFSR2_15(.LFSRregister(LFSRcolor2[735:690]),.clk(color1_clk));
lfsr #(.seed(46'b0010001010111001000011110110110110100001001011)) LFSR2_16(.LFSRregister(LFSRcolor2[781:736]),.clk(color1_clk));
lfsr #(.seed(46'b1010111110010100100000100111111111101010101011)) LFSR2_17(.LFSRregister(LFSRcolor2[827:782]),.clk(color1_clk));
lfsr #(.seed(46'b0000001101010010101110010000001110111100000000)) LFSR2_18(.LFSRregister(LFSRcolor2[873:828]),.clk(color1_clk));
lfsr #(.seed(46'b0001101011110001101001101001111111011101001010)) LFSR2_19(.LFSRregister(LFSRcolor2[919:874]),.clk(color1_clk));
lfsr #(.seed(46'b1010111010011010101000111010001000010011110111)) LFSR2_20(.LFSRregister(LFSRcolor2[965:920]),.clk(color1_clk));
lfsr #(.seed(46'b0001100101111110101010111111100101111000000011)) LFSR2_21(.LFSRregister(LFSRcolor2[1011:966]),.clk(color1_clk));
lfsr #(.seed(46'b1110110011101111100000001011100011010010100101)) LFSR2_22(.LFSRregister(LFSRcolor2[1057:1012]),.clk(color1_clk));
lfsr #(.seed(46'b1110101011011010101011001110110110100100110110)) LFSR2_23(.LFSRregister(LFSRcolor2[1103:1058]),.clk(color1_clk));
lfsr #(.seed(46'b0011111111100000000000011101001000101110111011)) LFSR2_24(.LFSRregister(LFSRcolor2[1149:1104]),.clk(color1_clk));
lfsr #(.seed(46'b0111111111000000001010100101100111000000010111)) LFSR2_25(.LFSRregister(LFSRcolor2[1195:1150]),.clk(color1_clk));
lfsr #(.seed(46'b0010111000110010000000110100011011001101000000)) LFSR2_26(.LFSRregister(LFSRcolor2[1241:1196]),.clk(color1_clk));
lfsr #(.seed(46'b1101101011000110111100101001100011010100111001)) LFSR2_27(.LFSRregister(LFSRcolor2[1287:1242]),.clk(color1_clk));
lfsr #(.seed(46'b1111011111010000011011010110110000011100001001)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1111101011000001010101111101111100010010110011)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b0101100101110001001001001101011110111001010010)) LFSR3_2(.LFSRregister(LFSRcolor3[137:92]),.clk(color2_clk));
lfsr #(.seed(46'b1101101001111010000010010010000100111110010001)) LFSR3_3(.LFSRregister(LFSRcolor3[183:138]),.clk(color2_clk));
lfsr #(.seed(46'b1111000000101100101101011010011110000100110011)) LFSR3_4(.LFSRregister(LFSRcolor3[229:184]),.clk(color2_clk));
lfsr #(.seed(46'b1101010101111111011100011001110101100110111001)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1000011111100100101011011011111000001100000011)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1011001100010110101100000111011111101000010100)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0100111111000101011011111100100110100001010010)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b1000111010001010000011110001100111110100110110)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b1100000100111011010101010100011010010011010000)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b0101010110001011110100001010110111000011000110)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b0110100110100010111000101000100010110011001010)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));
lfsr #(.seed(46'b1101101011000111110111100100101001001000001000)) LFSR4_8(.LFSRregister(LFSRcolor4[413:368]),.clk(color3_clk));
lfsr #(.seed(46'b0100101010101111111110001111100100100100000010)) LFSR4_9(.LFSRregister(LFSRcolor4[459:414]),.clk(color3_clk));
lfsr #(.seed(46'b0000001011001111100011100101111110011111110011)) LFSR4_10(.LFSRregister(LFSRcolor4[505:460]),.clk(color3_clk));
lfsr #(.seed(46'b0000011001011000001100001011001111011010110000)) LFSR4_11(.LFSRregister(LFSRcolor4[551:506]),.clk(color3_clk));
lfsr #(.seed(46'b0011010001101000011011101101001100000111110001)) LFSR4_12(.LFSRregister(LFSRcolor4[597:552]),.clk(color3_clk));
lfsr #(.seed(46'b1110101010010001010111100100100011110001110111)) LFSR4_13(.LFSRregister(LFSRcolor4[643:598]),.clk(color3_clk));
lfsr #(.seed(46'b0000101001010111110000010011110000110111101011)) LFSR4_14(.LFSRregister(LFSRcolor4[689:644]),.clk(color3_clk));
lfsr #(.seed(46'b0000011110001011011000010010101101101001100100)) LFSR4_15(.LFSRregister(LFSRcolor4[735:690]),.clk(color3_clk));
lfsr #(.seed(46'b0011110010101101111001000000011110000111110110)) LFSR4_16(.LFSRregister(LFSRcolor4[781:736]),.clk(color3_clk));
lfsr #(.seed(46'b0001011110001010011011010001010011100001100111)) LFSR4_17(.LFSRregister(LFSRcolor4[827:782]),.clk(color3_clk));
lfsr #(.seed(46'b0010011001101010001000101001001010101010110000)) LFSR4_18(.LFSRregister(LFSRcolor4[873:828]),.clk(color3_clk));
lfsr #(.seed(46'b1010001011001110001110110010000010100011011000)) LFSR4_19(.LFSRregister(LFSRcolor4[919:874]),.clk(color3_clk));
lfsr #(.seed(46'b1001101010011110100011110100010110011001110001)) LFSR4_20(.LFSRregister(LFSRcolor4[965:920]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 1;
initial m[1] = 1;
initial m[2] = 1;
initial m[3] = 0;
initial m[4] = 0;
initial m[5] = 0;
initial m[6] = 0;
initial m[7] = 0;
initial m[8] = 0;
initial m[9] = 1;
initial m[10] = 0;
initial m[11] = 1;
initial m[12] = 1;
initial m[13] = 0;
initial m[14] = 0;
initial m[15] = 0;
initial m[16] = 1;
initial m[17] = 0;
initial m[18] = 1;
initial m[19] = 1;
initial m[20] = 1;
initial m[21] = 1;
initial m[22] = 1;
initial m[23] = 1;
initial m[24] = 1;
initial m[25] = 1;
initial m[26] = 0;
initial m[27] = 0;
initial m[28] = 1;
initial m[29] = 0;
initial m[30] = 1;
initial m[31] = 1;
initial m[32] = 1;
initial m[33] = 1;
initial m[34] = 1;
initial m[35] = 1;
initial m[36] = 1;
initial m[37] = 1;
initial m[38] = 0;
initial m[39] = 1;
initial m[40] = 0;
initial m[41] = 1;
initial m[42] = 1;
initial m[43] = 1;
initial m[44] = 1;
initial m[45] = 0;
initial m[46] = 1;
initial m[47] = 1;
initial m[48] = 0;
initial m[49] = 1;
initial m[50] = 0;
initial m[51] = 0;
initial m[52] = 0;
initial m[53] = 0;
initial m[54] = 1;
initial m[55] = 1;
initial m[56] = 1;
initial m[57] = 1;
initial m[58] = 1;
initial m[59] = 0;
initial m[60] = 1;
initial m[61] = 1;
initial m[62] = 1;
initial m[63] = 1;
initial m[64] = 1;
initial m[65] = 1;
initial m[66] = 1;
initial m[67] = 1;
initial m[68] = 1;
initial m[69] = 0;
initial m[70] = 1;
initial m[71] = 0;
initial m[72] = 1;
initial m[73] = 1;
initial m[74] = 1;
initial m[75] = 0;
initial m[76] = 0;
initial m[77] = 0;
initial m[78] = 0;
initial m[79] = 1;
initial m[80] = 1;
initial m[81] = 1;
initial m[82] = 1;
initial m[83] = 0;
initial m[84] = 0;
initial m[85] = 0;
initial m[86] = 1;
initial m[87] = 1;
initial m[88] = 0;
initial m[89] = 0;
initial m[90] = 1;
initial m[91] = 0;
initial m[92] = 1;
initial m[93] = 1;
initial m[94] = 1;
initial m[95] = 0;
initial m[96] = 0;
initial m[97] = 1;
initial m[98] = 0;
initial m[99] = 1;
initial m[100] = 0;
initial m[101] = 1;
initial m[102] = 0;
initial m[103] = 1;
initial m[104] = 1;
initial m[105] = 1;
initial m[106] = 0;
initial m[107] = 0;
initial m[108] = 1;
initial m[109] = 0;
initial m[110] = 0;
initial m[111] = 0;
initial m[112] = 1;
initial m[113] = 1;
initial m[114] = 0;
initial m[115] = 1;
initial m[116] = 1;
initial m[117] = 1;
initial m[118] = 0;
initial m[119] = 1;
initial m[120] = 0;
initial m[121] = 1;
initial m[122] = 1;
initial m[123] = 1;
initial m[124] = 0;
initial m[125] = 0;
initial m[126] = 0;
initial m[127] = 0;
initial m[128] = 0;
initial m[129] = 1;
initial m[130] = 1;
initial m[131] = 1;
initial m[132] = 0;
initial m[133] = 0;
initial m[134] = 1;
initial m[135] = 0;
initial m[136] = 1;
initial m[137] = 0;
initial m[138] = 1;
initial m[139] = 1;
initial m[140] = 0;
initial m[141] = 1;
initial m[142] = 1;
initial m[143] = 1;
initial m[144] = 0;
initial m[145] = 1;
initial m[146] = 1;
initial m[147] = 1;
initial m[148] = 1;
initial m[149] = 1;
initial m[150] = 0;
initial m[151] = 0;
initial m[152] = 0;
initial m[153] = 0;
initial m[154] = 0;
initial m[155] = 1;
initial m[156] = 0;
initial m[157] = 0;
initial m[158] = 1;
initial m[159] = 1;
initial m[160] = 0;
initial m[161] = 1;
initial m[162] = 0;
initial m[163] = 1;
initial m[164] = 0;
initial m[165] = 1;
initial m[166] = 1;
initial m[167] = 1;
initial m[168] = 0;
initial m[169] = 0;
initial m[170] = 0;
initial m[171] = 1;
initial m[172] = 0;
initial m[173] = 0;
initial m[174] = 1;
initial m[175] = 1;
initial m[176] = 1;
initial m[177] = 1;
initial m[178] = 0;
initial m[179] = 1;
initial m[180] = 0;
initial m[181] = 1;
initial m[182] = 0;
initial m[183] = 1;
initial m[184] = 1;
initial m[185] = 0;
initial m[186] = 1;
initial m[187] = 1;
initial m[188] = 0;
initial m[189] = 0;
initial m[190] = 1;
initial m[191] = 1;
initial m[192] = 1;
initial m[193] = 1;
initial m[194] = 1;
initial m[195] = 0;
initial m[196] = 0;
initial m[197] = 0;
initial m[198] = 1;
initial m[199] = 1;
initial m[200] = 1;
initial m[201] = 1;
initial m[202] = 0;
initial m[203] = 0;
initial m[204] = 0;
initial m[205] = 1;
initial m[206] = 1;
initial m[207] = 1;
initial m[208] = 1;
initial m[209] = 0;
initial m[210] = 1;
initial m[211] = 0;
initial m[212] = 1;
initial m[213] = 0;
initial m[214] = 0;
initial m[215] = 0;
initial m[216] = 1;
initial m[217] = 1;
initial m[218] = 1;
initial m[219] = 1;
initial m[220] = 1;
initial m[221] = 1;
initial m[222] = 0;
initial m[223] = 0;
initial m[224] = 1;
initial m[225] = 1;
initial m[226] = 0;
initial m[227] = 0;
initial m[228] = 1;
initial m[229] = 1;
initial m[230] = 1;
initial m[231] = 0;
initial m[232] = 0;
initial m[233] = 0;
initial m[234] = 1;
initial m[235] = 1;
initial m[236] = 1;
initial m[237] = 1;
initial m[238] = 0;
initial m[239] = 1;
initial m[240] = 1;
initial m[241] = 0;
initial m[242] = 1;
initial m[243] = 0;
initial m[244] = 1;
initial m[245] = 1;
initial m[246] = 1;
initial m[247] = 0;
initial m[248] = 1;
initial m[249] = 1;
initial m[250] = 0;
initial m[251] = 1;
initial m[252] = 1;
initial m[253] = 0;
initial m[254] = 0;
initial m[255] = 1;
initial m[256] = 1;
initial m[257] = 0;
initial m[258] = 1;
initial m[259] = 0;
initial m[260] = 1;
initial m[261] = 1;
initial m[262] = 0;
initial m[263] = 0;
initial m[264] = 1;
initial m[265] = 1;
initial m[266] = 0;
initial m[267] = 1;
initial m[268] = 1;
initial m[269] = 1;
initial m[270] = 0;
initial m[271] = 1;
initial m[272] = 0;
initial m[273] = 0;
initial m[274] = 0;
initial m[275] = 0;
initial m[276] = 1;
initial m[277] = 0;
initial m[278] = 0;
initial m[279] = 0;
initial m[280] = 0;
initial m[281] = 0;
initial m[282] = 1;
initial m[283] = 0;
initial m[284] = 0;
initial m[285] = 0;
initial m[286] = 0;
initial m[287] = 0;
initial m[288] = 1;
initial m[289] = 0;
initial m[290] = 0;
initial m[291] = 1;
initial m[292] = 0;
initial m[293] = 1;
initial m[294] = 0;
initial m[295] = 1;
initial m[296] = 0;
initial m[297] = 0;
initial m[298] = 1;
initial m[299] = 1;
initial m[300] = 1;
initial m[301] = 0;
initial m[302] = 1;
initial m[303] = 0;
initial m[304] = 1;
initial m[305] = 1;
initial m[306] = 1;
initial m[307] = 0;
initial m[308] = 1;
initial m[309] = 0;
initial m[310] = 1;
initial m[311] = 1;
initial m[312] = 0;
initial m[313] = 0;
initial m[314] = 1;
initial m[315] = 0;
initial m[316] = 0;
initial m[317] = 0;
initial m[318] = 1;
initial m[319] = 0;
initial m[320] = 0;
initial m[321] = 0;
initial m[322] = 0;
initial m[323] = 0;
initial m[324] = 0;
initial m[325] = 1;
initial m[326] = 1;
initial m[327] = 1;
initial m[328] = 0;
initial m[329] = 1;
initial m[330] = 0;
initial m[331] = 1;
initial m[332] = 1;
initial m[333] = 0;
initial m[334] = 0;
initial m[335] = 0;
initial m[336] = 0;
initial m[337] = 0;
initial m[338] = 0;
initial m[339] = 0;
initial m[340] = 0;
initial m[341] = 1;
initial m[342] = 1;
initial m[343] = 1;
initial m[344] = 1;
initial m[345] = 1;
initial m[346] = 1;
initial m[347] = 0;
initial m[348] = 0;
initial m[349] = 0;
initial m[350] = 1;
initial m[351] = 1;
initial m[352] = 1;
initial m[353] = 0;
initial m[354] = 0;
initial m[355] = 0;
initial m[356] = 0;
initial m[357] = 0;
initial m[358] = 1;
initial m[359] = 1;
initial m[360] = 1;
initial m[361] = 1;
initial m[362] = 0;
initial m[363] = 0;
initial m[364] = 0;
initial m[365] = 1;
initial m[366] = 0;
initial m[367] = 0;
initial m[368] = 0;
initial m[369] = 0;
initial m[370] = 1;
initial m[371] = 1;
initial m[372] = 0;
initial m[373] = 0;
initial m[374] = 0;
initial m[375] = 0;
initial m[376] = 0;
initial m[377] = 1;
initial m[378] = 0;
initial m[379] = 1;
initial m[380] = 0;
initial m[381] = 0;
initial m[382] = 0;
initial m[383] = 1;
initial m[384] = 0;
initial m[385] = 1;
initial m[386] = 0;
initial m[387] = 1;
initial m[388] = 1;
initial m[389] = 1;
initial m[390] = 1;
initial m[391] = 0;
initial m[392] = 1;
initial m[393] = 1;
initial m[394] = 0;
initial m[395] = 0;
initial m[396] = 1;
initial m[397] = 1;
initial m[398] = 0;
initial m[399] = 0;
initial m[400] = 1;
initial m[401] = 0;
initial m[402] = 0;
initial m[403] = 1;
initial m[404] = 1;
initial m[405] = 1;
initial m[406] = 1;
initial m[407] = 1;
initial m[408] = 1;
initial m[409] = 1;
initial m[410] = 0;
initial m[411] = 0;
initial m[412] = 1;
initial m[413] = 0;
initial m[414] = 1;
initial m[415] = 0;
initial m[416] = 0;
initial m[417] = 0;
initial m[418] = 0;
initial m[419] = 0;
initial m[420] = 1;
initial m[421] = 1;
initial m[422] = 1;
initial m[423] = 1;
initial m[424] = 0;
initial m[425] = 0;
initial m[426] = 1;
initial m[427] = 1;
initial m[428] = 1;
initial m[429] = 0;
initial m[430] = 1;
initial m[431] = 0;
initial m[432] = 1;
initial m[433] = 0;
initial m[434] = 1;
initial m[435] = 0;
initial m[436] = 1;
initial m[437] = 1;
initial m[438] = 0;
initial m[439] = 1;
initial m[440] = 0;
initial m[441] = 0;
initial m[442] = 1;
initial m[443] = 0;
initial m[444] = 0;
initial m[445] = 1;
initial m[446] = 1;
initial m[447] = 1;
initial m[448] = 1;
initial m[449] = 0;
initial m[450] = 0;
initial m[451] = 1;
initial m[452] = 0;
initial m[453] = 0;
initial m[454] = 1;
initial m[455] = 0;
initial m[456] = 0;
initial m[457] = 1;
initial m[458] = 1;
initial m[459] = 1;
initial m[460] = 1;
initial m[461] = 1;
initial m[462] = 0;
initial m[463] = 1;
initial m[464] = 0;
initial m[465] = 1;
initial m[466] = 0;
initial m[467] = 0;
initial m[468] = 1;
initial m[469] = 0;
initial m[470] = 1;
initial m[471] = 0;
initial m[472] = 0;
initial m[473] = 1;
initial m[474] = 1;
initial m[475] = 1;
initial m[476] = 0;
initial m[477] = 1;
initial m[478] = 0;
initial m[479] = 1;
initial m[480] = 1;
initial m[481] = 0;
initial m[482] = 1;
initial m[483] = 1;
initial m[484] = 0;
initial m[485] = 1;
initial m[486] = 1;
initial m[487] = 1;
initial m[488] = 1;
initial m[489] = 1;
initial m[490] = 0;
initial m[491] = 0;
initial m[492] = 0;
initial m[493] = 0;
initial m[494] = 1;
initial m[495] = 0;
initial m[496] = 1;
initial m[497] = 0;
initial m[498] = 1;
initial m[499] = 0;
initial m[500] = 1;
initial m[501] = 1;
initial m[502] = 1;
initial m[503] = 1;
initial m[504] = 1;
initial m[505] = 1;
initial m[506] = 0;
initial m[507] = 1;
initial m[508] = 0;
initial m[509] = 1;
initial m[510] = 0;
initial m[511] = 0;
initial m[512] = 0;
initial m[513] = 1;
initial m[514] = 0;
initial m[515] = 0;
initial m[516] = 0;
initial m[517] = 1;
initial m[518] = 0;
initial m[519] = 0;
initial m[520] = 1;
initial m[521] = 0;
initial m[522] = 0;
initial m[523] = 0;
initial m[524] = 1;
initial m[525] = 1;
initial m[526] = 0;
initial m[527] = 0;
initial m[528] = 1;
initial m[529] = 1;
initial m[530] = 0;
initial m[531] = 0;
initial m[532] = 0;
initial m[533] = 0;
initial m[534] = 0;
initial m[535] = 1;
initial m[536] = 1;
initial m[537] = 0;
initial m[538] = 0;
initial m[539] = 1;
initial m[540] = 0;
initial m[541] = 1;
initial m[542] = 0;
initial m[543] = 0;
initial m[544] = 0;
initial m[545] = 0;
initial m[546] = 0;
initial m[547] = 0;
initial m[548] = 0;
initial m[549] = 1;
initial m[550] = 0;
initial m[551] = 1;
initial m[552] = 1;
initial m[553] = 0;
initial m[554] = 0;
initial m[555] = 1;
initial m[556] = 0;
initial m[557] = 1;
initial m[558] = 0;
initial m[559] = 0;
initial m[560] = 0;
initial m[561] = 1;
initial m[562] = 1;
initial m[563] = 0;
initial m[564] = 0;
initial m[565] = 1;
initial m[566] = 0;
initial m[567] = 0;
initial m[568] = 0;
initial m[569] = 0;
initial m[570] = 1;
initial m[571] = 0;
initial m[572] = 0;
initial m[573] = 0;
initial m[574] = 1;
initial m[575] = 1;
initial m[576] = 0;
initial m[577] = 0;
initial m[578] = 1;
initial m[579] = 1;
initial m[580] = 1;
initial m[581] = 1;
initial m[582] = 1;
initial m[583] = 1;
initial m[584] = 0;
initial m[585] = 0;
initial m[586] = 0;
initial m[587] = 1;
initial m[588] = 1;
initial m[589] = 0;
initial m[590] = 0;
initial m[591] = 0;
initial m[592] = 0;
initial m[593] = 0;
initial m[594] = 0;
initial m[595] = 0;
initial m[596] = 1;
initial m[597] = 0;
initial m[598] = 0;
initial m[599] = 1;
initial m[600] = 1;
initial m[601] = 1;
initial m[602] = 0;
initial m[603] = 1;
initial m[604] = 1;
initial m[605] = 0;
initial m[606] = 0;
initial m[607] = 0;
initial m[608] = 0;
initial m[609] = 1;
initial m[610] = 0;
initial m[611] = 0;
initial m[612] = 0;
initial m[613] = 1;
initial m[614] = 0;
initial m[615] = 0;
initial m[616] = 0;
initial m[617] = 1;
initial m[618] = 0;
initial m[619] = 1;
initial m[620] = 0;
initial m[621] = 0;
initial m[622] = 0;
initial m[623] = 0;
initial m[624] = 0;
initial m[625] = 0;
initial m[626] = 1;
initial m[627] = 1;
initial m[628] = 0;
initial m[629] = 1;
initial m[630] = 1;
initial m[631] = 1;
initial m[632] = 0;
initial m[633] = 1;
initial m[634] = 1;
initial m[635] = 0;
initial m[636] = 1;
initial m[637] = 0;
initial m[638] = 0;
initial m[639] = 1;
initial m[640] = 0;
initial m[641] = 0;
initial m[642] = 0;
initial m[643] = 1;
initial m[644] = 0;
initial m[645] = 1;
initial m[646] = 1;
initial m[647] = 1;
initial m[648] = 1;
initial m[649] = 0;
initial m[650] = 0;
initial m[651] = 0;
initial m[652] = 1;
initial m[653] = 1;
initial m[654] = 0;
initial m[655] = 0;
initial m[656] = 0;
initial m[657] = 1;
initial m[658] = 0;
initial m[659] = 0;
initial m[660] = 0;
initial m[661] = 0;
initial m[662] = 0;
initial m[663] = 0;
initial m[664] = 1;
initial m[665] = 1;
initial m[666] = 0;
initial m[667] = 0;
initial m[668] = 0;
initial m[669] = 1;
initial m[670] = 0;
initial m[671] = 1;
initial m[673] = 1;
initial m[674] = 0;
initial m[675] = 0;
initial m[676] = 1;
initial m[677] = 0;
initial m[678] = 1;
initial m[679] = 1;
initial m[680] = 1;
initial m[681] = 1;
initial m[682] = 1;
initial m[683] = 0;
initial m[684] = 1;
initial m[685] = 0;
initial m[686] = 1;
initial m[687] = 0;
initial m[688] = 1;
initial m[689] = 1;
initial m[690] = 0;
initial m[691] = 1;
initial m[692] = 0;
initial m[693] = 1;
initial m[694] = 1;
initial m[695] = 0;
initial m[696] = 0;
initial m[697] = 0;
initial m[698] = 1;
initial m[699] = 0;
initial m[700] = 0;
initial m[701] = 1;
initial m[702] = 0;
initial m[703] = 1;
initial m[704] = 0;
initial m[705] = 0;
initial m[706] = 1;
initial m[707] = 1;
initial m[708] = 0;
initial m[709] = 1;
initial m[710] = 1;
initial m[711] = 1;
initial m[712] = 1;
initial m[713] = 0;
initial m[714] = 0;
initial m[715] = 1;
initial m[716] = 1;
initial m[717] = 0;
initial m[718] = 1;
initial m[719] = 0;
initial m[720] = 1;
initial m[721] = 1;
initial m[722] = 1;
initial m[723] = 1;
initial m[724] = 0;
initial m[725] = 0;
initial m[726] = 1;
initial m[727] = 0;
initial m[728] = 1;
initial m[729] = 0;
initial m[730] = 1;
initial m[731] = 0;
initial m[732] = 1;
initial m[733] = 0;
initial m[734] = 1;
initial m[735] = 0;
initial m[736] = 0;
initial m[737] = 1;
initial m[738] = 0;
initial m[739] = 1;
initial m[740] = 1;
initial m[741] = 0;
initial m[742] = 0;
initial m[743] = 0;
initial m[744] = 1;
initial m[745] = 1;
initial m[746] = 1;
initial m[747] = 1;
initial m[748] = 1;
initial m[749] = 1;
initial m[750] = 0;
initial m[751] = 0;
initial m[752] = 0;
initial m[753] = 1;
initial m[754] = 0;
initial m[755] = 0;
initial m[756] = 0;
initial m[757] = 1;
initial m[758] = 1;
initial m[759] = 1;
initial m[760] = 1;
initial m[761] = 1;
initial m[762] = 1;
initial m[763] = 0;
initial m[764] = 0;
initial m[765] = 1;
initial m[766] = 1;
initial m[767] = 1;
initial m[768] = 0;
initial m[769] = 1;
initial m[770] = 1;
initial m[771] = 0;
initial m[772] = 0;
initial m[773] = 1;
initial m[774] = 1;
initial m[775] = 1;
initial m[776] = 1;
initial m[777] = 1;
initial m[778] = 1;
initial m[779] = 1;
initial m[780] = 1;
initial m[781] = 1;
initial m[782] = 1;
initial m[783] = 0;
initial m[784] = 0;
initial m[785] = 1;
initial m[786] = 1;
initial m[787] = 0;
initial m[788] = 1;
initial m[789] = 1;
initial m[790] = 1;
initial m[791] = 1;
initial m[792] = 1;
initial m[793] = 1;
initial m[794] = 0;
initial m[795] = 0;
initial m[796] = 0;
initial m[797] = 1;
initial m[798] = 1;
initial m[799] = 1;
initial m[800] = 1;
initial m[801] = 0;
initial m[802] = 0;
initial m[803] = 1;
initial m[804] = 1;
initial m[805] = 0;
initial m[806] = 1;
initial m[807] = 0;
initial m[808] = 0;
initial m[809] = 1;
initial m[810] = 1;
initial m[811] = 1;
initial m[812] = 0;
initial m[813] = 0;
initial m[814] = 1;
initial m[815] = 0;
initial m[816] = 1;
initial m[817] = 1;
initial m[818] = 0;
initial m[819] = 0;
initial m[820] = 0;
initial m[821] = 1;
initial m[822] = 1;
initial m[823] = 1;
initial m[824] = 1;
initial m[825] = 0;
initial m[826] = 0;
initial m[827] = 1;
initial m[828] = 0;
initial m[829] = 1;
initial m[830] = 0;
initial m[831] = 0;
initial m[832] = 0;
initial m[833] = 1;
initial m[834] = 1;
initial m[835] = 0;
initial m[836] = 1;
initial m[837] = 0;
initial m[838] = 1;
initial m[839] = 1;
initial m[840] = 0;
initial m[841] = 1;
initial m[842] = 1;
initial m[843] = 0;
initial m[844] = 1;
initial m[845] = 1;
initial m[846] = 1;
initial m[847] = 1;
initial m[848] = 1;
initial m[849] = 0;
initial m[850] = 1;
initial m[851] = 0;
initial m[852] = 0;
initial m[853] = 1;
initial m[854] = 0;
initial m[855] = 0;
initial m[856] = 0;
initial m[857] = 0;
initial m[858] = 0;
initial m[859] = 1;
initial m[860] = 1;
initial m[861] = 1;
initial m[862] = 0;
initial m[863] = 1;
initial m[864] = 0;
initial m[865] = 0;
initial m[866] = 0;
initial m[867] = 1;
initial m[868] = 0;
initial m[869] = 0;
initial m[870] = 1;
initial m[871] = 1;
initial m[872] = 0;
initial m[873] = 0;
initial m[874] = 1;
initial m[875] = 0;
initial m[876] = 0;
initial m[877] = 0;
initial m[878] = 0;
initial m[879] = 0;
initial m[880] = 0;
initial m[881] = 1;
initial m[882] = 1;
initial m[883] = 0;
initial m[884] = 0;
initial m[885] = 1;
initial m[886] = 1;
initial m[887] = 1;
initial m[888] = 0;
initial m[889] = 1;
initial m[890] = 1;
initial m[891] = 1;
initial m[892] = 1;
initial m[893] = 0;
initial m[894] = 1;
initial m[895] = 1;
initial m[896] = 0;
initial m[897] = 1;
initial m[898] = 0;
initial m[899] = 1;
initial m[900] = 0;
initial m[901] = 1;
initial m[902] = 0;
initial m[903] = 1;
initial m[904] = 1;
initial m[905] = 0;
initial m[906] = 1;
initial m[907] = 0;
initial m[908] = 1;
initial m[909] = 1;
initial m[910] = 0;
initial m[911] = 1;
initial m[912] = 0;
initial m[913] = 1;
initial m[914] = 1;
initial m[915] = 1;
initial m[916] = 1;
initial m[917] = 0;
initial m[918] = 1;
initial m[919] = 1;
initial m[920] = 0;
initial m[921] = 1;
initial m[922] = 1;
initial m[923] = 0;
initial m[924] = 0;
initial m[925] = 0;
initial m[926] = 0;
initial m[927] = 0;
initial m[928] = 0;
initial m[929] = 1;
initial m[932] = 0;
initial m[933] = 1;
initial m[934] = 0;
initial m[935] = 1;
initial m[936] = 1;
initial m[937] = 1;
initial m[938] = 1;
initial m[939] = 0;
initial m[942] = 1;
initial m[943] = 0;
initial m[944] = 0;
initial m[945] = 0;
initial m[946] = 0;
initial m[947] = 0;
initial m[948] = 0;
initial m[949] = 0;
initial m[950] = 0;
initial m[951] = 1;
initial m[952] = 0;
initial m[953] = 0;
initial m[954] = 1;
initial m[957] = 1;
initial m[958] = 1;
initial m[959] = 1;
initial m[960] = 0;
initial m[961] = 1;
initial m[962] = 0;
initial m[963] = 0;
initial m[964] = 1;
initial m[965] = 1;
initial m[966] = 1;
initial m[967] = 0;
initial m[968] = 0;
initial m[969] = 0;
initial m[970] = 0;
initial m[971] = 1;
initial m[972] = 1;
initial m[973] = 1;
initial m[974] = 0;
initial m[977] = 1;
initial m[978] = 1;
initial m[979] = 0;
initial m[980] = 1;
initial m[981] = 1;
initial m[982] = 0;
initial m[983] = 0;
initial m[984] = 1;
initial m[985] = 1;
initial m[986] = 1;
initial m[987] = 0;
initial m[988] = 0;
initial m[989] = 1;
initial m[990] = 0;
initial m[991] = 1;
initial m[992] = 0;
initial m[993] = 0;
initial m[994] = 0;
initial m[995] = 1;
initial m[996] = 1;
initial m[997] = 1;
initial m[998] = 0;
initial m[999] = 1;
initial m[1002] = 0;
initial m[1003] = 0;
initial m[1004] = 0;
initial m[1005] = 1;
initial m[1006] = 0;
initial m[1007] = 0;
initial m[1008] = 1;
initial m[1009] = 1;
initial m[1010] = 0;
initial m[1011] = 1;
initial m[1012] = 1;
initial m[1013] = 1;
initial m[1014] = 0;
initial m[1015] = 0;
initial m[1016] = 1;
initial m[1017] = 1;
initial m[1018] = 1;
initial m[1019] = 0;
initial m[1020] = 1;
initial m[1021] = 1;
initial m[1022] = 1;
initial m[1023] = 1;
initial m[1024] = 0;
initial m[1025] = 0;
initial m[1026] = 1;
initial m[1027] = 1;
initial m[1028] = 1;
initial m[1029] = 1;
initial m[1032] = 1;
initial m[1033] = 1;
initial m[1034] = 0;
initial m[1035] = 1;
initial m[1036] = 1;
initial m[1037] = 0;
initial m[1038] = 1;
initial m[1039] = 1;
initial m[1040] = 1;
initial m[1041] = 1;
initial m[1042] = 1;
initial m[1043] = 1;
initial m[1044] = 0;
initial m[1045] = 0;
initial m[1046] = 0;
initial m[1047] = 0;
initial m[1048] = 0;
initial m[1049] = 1;
initial m[1050] = 0;
initial m[1051] = 1;
initial m[1052] = 0;
initial m[1053] = 0;
initial m[1054] = 1;
initial m[1055] = 1;
initial m[1056] = 1;
initial m[1057] = 0;
initial m[1058] = 1;
initial m[1059] = 0;
initial m[1060] = 0;
initial m[1061] = 1;
initial m[1062] = 1;
initial m[1063] = 0;
initial m[1064] = 0;
initial m[1067] = 1;
initial m[1068] = 0;
initial m[1069] = 1;
initial m[1070] = 1;
initial m[1071] = 1;
initial m[1072] = 1;
initial m[1073] = 0;
initial m[1074] = 0;
initial m[1075] = 1;
initial m[1076] = 0;
initial m[1077] = 1;
initial m[1078] = 0;
initial m[1079] = 1;
initial m[1080] = 1;
initial m[1081] = 1;
initial m[1082] = 0;
initial m[1083] = 0;
initial m[1084] = 0;
initial m[1085] = 1;
initial m[1086] = 1;
initial m[1087] = 0;
initial m[1088] = 0;
initial m[1089] = 1;
initial m[1090] = 1;
initial m[1091] = 0;
initial m[1092] = 0;
initial m[1093] = 1;
initial m[1094] = 1;
initial m[1095] = 1;
initial m[1096] = 1;
initial m[1097] = 0;
initial m[1098] = 1;
initial m[1099] = 1;
initial m[1100] = 0;
initial m[1101] = 1;
initial m[1102] = 0;
initial m[1103] = 1;
initial m[1104] = 1;
initial m[1107] = 0;
initial m[1108] = 1;
initial m[1109] = 0;
initial m[1110] = 1;
initial m[1111] = 0;
initial m[1112] = 1;
initial m[1113] = 1;
initial m[1114] = 1;
initial m[1115] = 0;
initial m[1116] = 1;
initial m[1117] = 0;
initial m[1118] = 0;
initial m[1119] = 1;
initial m[1120] = 1;
initial m[1121] = 0;
initial m[1122] = 1;
initial m[1123] = 0;
initial m[1124] = 1;
initial m[1125] = 0;
initial m[1126] = 0;
initial m[1127] = 0;
initial m[1128] = 0;
initial m[1129] = 1;
initial m[1130] = 1;
initial m[1131] = 1;
initial m[1132] = 1;
initial m[1133] = 1;
initial m[1134] = 0;
initial m[1135] = 1;
initial m[1136] = 0;
initial m[1137] = 0;
initial m[1138] = 0;
initial m[1139] = 0;
initial m[1140] = 1;
initial m[1141] = 0;
initial m[1142] = 0;
initial m[1143] = 1;
initial m[1144] = 1;
initial m[1145] = 0;
initial m[1146] = 1;
initial m[1147] = 0;
initial m[1148] = 0;
initial m[1149] = 1;
initial m[1152] = 0;
initial m[1153] = 1;
initial m[1154] = 0;
initial m[1155] = 1;
initial m[1156] = 0;
initial m[1157] = 1;
initial m[1158] = 1;
initial m[1159] = 1;
initial m[1160] = 1;
initial m[1161] = 1;
initial m[1162] = 1;
initial m[1163] = 1;
initial m[1164] = 0;
initial m[1165] = 0;
initial m[1166] = 1;
initial m[1167] = 0;
initial m[1168] = 0;
initial m[1169] = 1;
initial m[1170] = 1;
initial m[1171] = 0;
initial m[1172] = 1;
initial m[1173] = 1;
initial m[1174] = 0;
initial m[1175] = 1;
initial m[1176] = 0;
initial m[1177] = 0;
initial m[1178] = 1;
initial m[1179] = 1;
initial m[1180] = 0;
initial m[1181] = 0;
initial m[1182] = 1;
initial m[1183] = 1;
initial m[1184] = 0;
initial m[1185] = 1;
initial m[1186] = 1;
initial m[1187] = 0;
initial m[1188] = 0;
initial m[1189] = 0;
initial m[1190] = 1;
initial m[1191] = 0;
initial m[1192] = 1;
initial m[1193] = 0;
initial m[1194] = 1;
initial m[1195] = 0;
initial m[1196] = 0;
initial m[1197] = 0;
initial m[1198] = 0;
initial m[1199] = 0;
initial m[1202] = 1;
initial m[1203] = 1;
initial m[1204] = 1;
initial m[1205] = 1;
initial m[1206] = 1;
initial m[1207] = 0;
initial m[1208] = 1;
initial m[1209] = 0;
initial m[1210] = 0;
initial m[1211] = 1;
initial m[1212] = 0;
initial m[1213] = 1;
initial m[1214] = 1;
initial m[1215] = 1;
initial m[1216] = 1;
initial m[1217] = 0;
initial m[1218] = 0;
initial m[1219] = 0;
initial m[1220] = 1;
initial m[1221] = 0;
initial m[1222] = 0;
initial m[1223] = 1;
initial m[1224] = 1;
initial m[1225] = 0;
initial m[1226] = 0;
initial m[1227] = 0;
initial m[1228] = 0;
initial m[1229] = 0;
initial m[1230] = 1;
initial m[1231] = 1;
initial m[1232] = 1;
initial m[1233] = 1;
initial m[1234] = 0;
initial m[1235] = 1;
initial m[1236] = 0;
initial m[1237] = 1;
initial m[1238] = 1;
initial m[1239] = 1;
initial m[1240] = 1;
initial m[1241] = 1;
initial m[1242] = 0;
initial m[1243] = 1;
initial m[1244] = 1;
initial m[1245] = 0;
initial m[1246] = 0;
initial m[1247] = 1;
initial m[1248] = 1;
initial m[1249] = 1;
initial m[1250] = 0;
initial m[1251] = 0;
initial m[1252] = 0;
initial m[1253] = 0;
initial m[1254] = 0;
initial m[1257] = 1;
initial m[1258] = 1;
initial m[1259] = 0;
initial m[1260] = 0;
initial m[1261] = 0;
initial m[1262] = 0;
initial m[1263] = 1;
initial m[1264] = 0;
initial m[1265] = 1;
initial m[1266] = 1;
initial m[1267] = 1;
initial m[1268] = 1;
initial m[1269] = 0;
initial m[1270] = 0;
initial m[1271] = 0;
initial m[1272] = 0;
initial m[1273] = 1;
initial m[1274] = 1;
initial m[1275] = 0;
initial m[1276] = 1;
initial m[1277] = 1;
initial m[1278] = 0;
initial m[1279] = 1;
initial m[1280] = 1;
initial m[1281] = 1;
initial m[1282] = 1;
initial m[1283] = 1;
initial m[1284] = 0;
initial m[1285] = 0;
initial m[1286] = 1;
initial m[1287] = 1;
initial m[1288] = 1;
initial m[1289] = 1;
initial m[1290] = 0;
initial m[1291] = 1;
initial m[1292] = 0;
initial m[1293] = 0;
initial m[1294] = 0;
initial m[1295] = 1;
initial m[1296] = 1;
initial m[1297] = 0;
initial m[1298] = 1;
initial m[1299] = 1;
initial m[1300] = 0;
initial m[1301] = 1;
initial m[1302] = 0;
initial m[1303] = 1;
initial m[1304] = 1;
initial m[1305] = 0;
initial m[1306] = 1;
initial m[1307] = 1;
initial m[1308] = 0;
initial m[1309] = 0;
initial m[1310] = 0;
initial m[1311] = 0;
initial m[1312] = 1;
initial m[1313] = 0;
initial m[1314] = 1;
initial m[1317] = 1;
initial m[1318] = 0;
initial m[1319] = 0;
initial m[1320] = 1;
initial m[1321] = 0;
initial m[1322] = 1;
initial m[1323] = 1;
initial m[1324] = 1;
initial m[1325] = 0;
initial m[1326] = 0;
initial m[1327] = 1;
initial m[1328] = 1;
initial m[1329] = 0;
initial m[1330] = 1;
initial m[1331] = 0;
initial m[1332] = 0;
initial m[1333] = 1;
initial m[1334] = 0;
initial m[1335] = 1;
initial m[1336] = 1;
initial m[1337] = 1;
initial m[1338] = 1;
initial m[1339] = 1;
initial m[1340] = 1;
initial m[1341] = 0;
initial m[1342] = 0;
initial m[1343] = 1;
initial m[1344] = 0;
initial m[1345] = 0;
initial m[1346] = 0;
initial m[1347] = 0;
initial m[1348] = 0;
initial m[1349] = 0;
initial m[1350] = 1;
initial m[1351] = 0;
initial m[1352] = 0;
initial m[1353] = 0;
initial m[1354] = 0;
initial m[1355] = 0;
initial m[1356] = 1;
initial m[1357] = 0;
initial m[1358] = 1;
initial m[1359] = 0;
initial m[1360] = 1;
initial m[1361] = 1;
initial m[1362] = 1;
initial m[1363] = 0;
initial m[1364] = 0;
initial m[1365] = 0;
initial m[1366] = 0;
initial m[1367] = 1;
initial m[1368] = 0;
initial m[1369] = 1;
initial m[1370] = 1;
initial m[1371] = 1;
initial m[1372] = 0;
initial m[1373] = 0;
initial m[1374] = 1;
initial m[1375] = 1;
initial m[1376] = 0;
initial m[1377] = 0;
initial m[1378] = 1;
initial m[1379] = 1;
initial m[1382] = 0;
initial m[1383] = 1;
initial m[1384] = 0;
initial m[1385] = 1;
initial m[1386] = 0;
initial m[1387] = 0;
initial m[1388] = 1;
initial m[1389] = 0;
initial m[1390] = 1;
initial m[1391] = 0;
initial m[1392] = 0;
initial m[1393] = 1;
initial m[1394] = 1;
initial m[1395] = 0;
initial m[1396] = 1;
initial m[1397] = 1;
initial m[1398] = 1;
initial m[1399] = 0;
initial m[1400] = 0;
initial m[1401] = 0;
initial m[1402] = 1;
initial m[1403] = 1;
initial m[1404] = 1;
initial m[1405] = 0;
initial m[1406] = 0;
initial m[1407] = 1;
initial m[1408] = 1;
initial m[1409] = 1;
initial m[1410] = 0;
initial m[1411] = 1;
initial m[1412] = 1;
initial m[1413] = 0;
initial m[1414] = 1;
initial m[1415] = 0;
initial m[1416] = 1;
initial m[1417] = 1;
initial m[1418] = 0;
initial m[1419] = 1;
initial m[1420] = 1;
initial m[1421] = 0;
initial m[1422] = 1;
initial m[1423] = 0;
initial m[1424] = 1;
initial m[1425] = 1;
initial m[1426] = 0;
initial m[1427] = 0;
initial m[1428] = 0;
initial m[1429] = 0;
initial m[1430] = 1;
initial m[1431] = 1;
initial m[1432] = 0;
initial m[1433] = 1;
initial m[1434] = 0;
initial m[1435] = 0;
initial m[1436] = 0;
initial m[1437] = 1;
initial m[1438] = 0;
initial m[1439] = 1;
initial m[1440] = 1;
initial m[1441] = 1;
initial m[1442] = 0;
initial m[1443] = 1;
initial m[1444] = 1;
initial m[1445] = 0;
initial m[1446] = 1;
initial m[1447] = 0;
initial m[1448] = 0;
initial m[1449] = 0;
initial m[1452] = 0;
initial m[1453] = 0;
initial m[1454] = 0;
initial m[1455] = 1;
initial m[1456] = 1;
initial m[1457] = 1;
initial m[1458] = 1;
initial m[1459] = 1;
initial m[1460] = 1;
initial m[1461] = 1;
initial m[1462] = 1;
initial m[1463] = 1;
initial m[1464] = 1;
initial m[1465] = 0;
initial m[1466] = 0;
initial m[1467] = 0;
initial m[1468] = 0;
initial m[1469] = 0;
initial m[1470] = 0;
initial m[1471] = 0;
initial m[1472] = 0;
initial m[1473] = 0;
initial m[1474] = 1;
initial m[1475] = 1;
initial m[1476] = 1;
initial m[1477] = 1;
initial m[1478] = 0;
initial m[1479] = 0;
initial m[1480] = 0;
initial m[1481] = 1;
initial m[1482] = 0;
initial m[1483] = 0;
initial m[1484] = 0;
initial m[1485] = 1;
initial m[1486] = 0;
initial m[1487] = 0;
initial m[1488] = 1;
initial m[1489] = 0;
initial m[1490] = 0;
initial m[1491] = 0;
initial m[1492] = 0;
initial m[1493] = 0;
initial m[1494] = 0;
initial m[1495] = 1;
initial m[1496] = 1;
initial m[1497] = 1;
initial m[1498] = 0;
initial m[1499] = 1;
initial m[1500] = 1;
initial m[1501] = 1;
initial m[1502] = 0;
initial m[1503] = 1;
initial m[1504] = 1;
initial m[1505] = 1;
initial m[1506] = 0;
initial m[1507] = 0;
initial m[1508] = 1;
initial m[1509] = 1;
initial m[1510] = 1;
initial m[1511] = 1;
initial m[1512] = 1;
initial m[1513] = 0;
initial m[1514] = 1;
initial m[1515] = 1;
initial m[1516] = 1;
initial m[1517] = 1;
initial m[1518] = 1;
initial m[1519] = 1;
initial m[1520] = 0;
initial m[1521] = 1;
initial m[1522] = 0;
initial m[1523] = 0;
initial m[1524] = 0;
initial m[1527] = 1;
initial m[1529] = 0;
initial m[1530] = 0;
initial m[1531] = 0;
initial m[1532] = 1;
initial m[1533] = 0;
initial m[1534] = 0;
initial m[1535] = 1;
initial m[1536] = 1;
initial m[1537] = 0;
initial m[1538] = 1;
initial m[1539] = 1;
initial m[1540] = 1;
initial m[1541] = 1;
initial m[1542] = 0;
initial m[1543] = 1;
initial m[1544] = 0;
initial m[1545] = 0;
initial m[1546] = 1;
initial m[1547] = 0;
initial m[1548] = 0;
initial m[1549] = 0;
initial m[1550] = 0;
initial m[1551] = 0;
initial m[1552] = 1;
initial m[1553] = 1;
initial m[1554] = 1;
initial m[1555] = 1;
initial m[1556] = 1;
initial m[1557] = 1;
initial m[1558] = 0;
initial m[1559] = 1;
initial m[1560] = 1;
initial m[1561] = 0;
initial m[1562] = 1;
initial m[1563] = 1;
initial m[1564] = 0;
initial m[1565] = 0;
initial m[1566] = 1;
initial m[1567] = 1;
initial m[1568] = 0;
initial m[1569] = 1;
initial m[1570] = 1;
initial m[1571] = 0;
initial m[1572] = 1;
initial m[1573] = 0;
initial m[1574] = 0;
initial m[1575] = 1;
initial m[1576] = 1;
initial m[1577] = 1;
initial m[1578] = 1;
initial m[1579] = 1;
initial m[1580] = 0;
initial m[1581] = 1;
initial m[1582] = 0;
initial m[1583] = 0;
initial m[1584] = 0;
initial m[1585] = 0;
initial m[1586] = 0;
initial m[1587] = 0;
initial m[1588] = 1;
initial m[1589] = 0;
initial m[1590] = 1;
initial m[1591] = 0;
initial m[1592] = 0;
initial m[1593] = 1;
initial m[1594] = 1;
initial m[1595] = 0;
initial m[1596] = 1;
initial m[1597] = 1;
initial m[1598] = 1;
initial m[1599] = 0;
initial m[1600] = 1;
initial m[1602] = 0;
initial m[1603] = 1;
initial m[1604] = 0;
initial m[1605] = 0;
initial m[1606] = 0;
initial m[1607] = 1;
initial m[1608] = 0;
initial m[1609] = 1;
initial m[1610] = 0;
initial m[1611] = 1;
initial m[1612] = 0;
initial m[1613] = 1;
initial m[1614] = 1;
initial m[1615] = 1;
initial m[1616] = 1;
initial m[1617] = 1;
initial m[1618] = 0;
initial m[1619] = 0;
initial m[1620] = 0;
initial m[1621] = 0;
initial m[1622] = 0;
initial m[1623] = 1;
initial m[1624] = 1;
initial m[1625] = 0;
initial m[1626] = 1;
initial m[1627] = 0;
initial m[1628] = 0;
initial m[1629] = 0;
initial m[1630] = 1;
initial m[1631] = 0;
initial m[1632] = 1;
initial m[1633] = 1;
initial m[1634] = 1;
initial m[1635] = 0;
initial m[1636] = 0;
initial m[1637] = 0;
initial m[1638] = 1;
initial m[1639] = 1;
initial m[1640] = 0;
initial m[1641] = 1;
initial m[1642] = 1;
initial m[1643] = 1;
initial m[1644] = 0;
initial m[1645] = 1;
initial m[1646] = 1;
initial m[1647] = 0;
initial m[1648] = 0;
initial m[1649] = 0;
initial m[1650] = 0;
initial m[1651] = 1;
initial m[1652] = 1;
initial m[1653] = 0;
initial m[1654] = 0;
initial m[1655] = 1;
initial m[1656] = 1;
initial m[1657] = 1;
initial m[1658] = 0;
initial m[1659] = 0;
initial m[1660] = 1;
initial m[1661] = 0;
initial m[1662] = 0;
initial m[1663] = 1;
initial m[1664] = 0;
initial m[1665] = 0;
initial m[1666] = 1;
initial m[1667] = 0;
initial m[1668] = 1;
initial m[1669] = 0;
initial m[1670] = 1;
initial m[1672] = 1;
initial m[1673] = 0;
initial m[1674] = 1;
initial m[1675] = 0;
initial m[1676] = 0;
initial m[1677] = 1;
initial m[1678] = 0;
initial m[1679] = 1;
initial m[1680] = 0;
initial m[1681] = 0;
initial m[1682] = 0;
initial m[1683] = 0;
initial m[1684] = 0;
initial m[1685] = 0;
initial m[1686] = 0;
initial m[1687] = 1;
initial m[1688] = 0;
initial m[1689] = 0;
initial m[1690] = 1;
initial m[1691] = 0;
initial m[1692] = 1;
initial m[1693] = 0;
initial m[1694] = 0;
initial m[1695] = 1;
initial m[1696] = 1;
initial m[1697] = 0;
initial m[1698] = 0;
initial m[1699] = 1;
initial m[1700] = 1;
initial m[1701] = 1;
initial m[1702] = 0;
initial m[1703] = 1;
initial m[1704] = 1;
initial m[1705] = 1;
initial m[1706] = 0;
initial m[1707] = 1;
initial m[1708] = 1;
initial m[1709] = 1;
initial m[1710] = 1;
initial m[1711] = 0;
initial m[1712] = 0;
initial m[1713] = 0;
initial m[1714] = 1;
initial m[1715] = 1;
initial m[1716] = 0;
initial m[1717] = 1;
initial m[1718] = 1;
initial m[1719] = 0;
initial m[1720] = 0;
initial m[1721] = 0;
initial m[1722] = 1;
initial m[1723] = 0;
initial m[1724] = 1;
initial m[1725] = 1;
initial m[1726] = 1;
initial m[1727] = 0;
initial m[1728] = 0;
initial m[1729] = 1;
initial m[1730] = 1;
initial m[1731] = 0;
initial m[1732] = 1;
initial m[1733] = 0;
initial m[1734] = 1;
initial m[1735] = 0;
initial m[1737] = 1;
initial m[1738] = 1;
initial m[1739] = 0;
initial m[1740] = 0;
initial m[1741] = 1;
initial m[1742] = 1;
initial m[1743] = 0;
initial m[1744] = 1;
initial m[1745] = 1;
initial m[1746] = 1;
initial m[1747] = 1;
initial m[1748] = 0;
initial m[1749] = 1;
initial m[1750] = 1;
initial m[1751] = 1;
initial m[1752] = 0;
initial m[1753] = 1;
initial m[1754] = 1;
initial m[1755] = 1;
initial m[1756] = 0;
initial m[1757] = 1;
initial m[1758] = 1;
initial m[1759] = 0;
initial m[1760] = 1;
initial m[1761] = 1;
initial m[1762] = 1;
initial m[1763] = 0;
initial m[1764] = 0;
initial m[1765] = 1;
initial m[1766] = 0;
initial m[1767] = 0;
initial m[1768] = 0;
initial m[1769] = 0;
initial m[1770] = 0;
initial m[1771] = 1;
initial m[1772] = 0;
initial m[1773] = 0;
initial m[1774] = 0;
initial m[1775] = 0;
initial m[1776] = 0;
initial m[1777] = 0;
initial m[1778] = 0;
initial m[1779] = 0;
initial m[1780] = 0;
initial m[1781] = 0;
initial m[1782] = 1;
initial m[1783] = 0;
initial m[1784] = 0;
initial m[1785] = 0;
initial m[1786] = 1;
initial m[1787] = 0;
initial m[1788] = 1;
initial m[1789] = 1;
initial m[1790] = 1;
initial m[1791] = 1;
initial m[1792] = 1;
initial m[1793] = 0;
initial m[1794] = 1;
initial m[1795] = 1;
initial m[1797] = 1;
initial m[1798] = 0;
initial m[1799] = 1;
initial m[1800] = 1;
initial m[1801] = 0;
initial m[1802] = 1;
initial m[1803] = 0;
initial m[1804] = 0;
initial m[1805] = 1;
initial m[1806] = 1;
initial m[1807] = 1;
initial m[1808] = 0;
initial m[1809] = 1;
initial m[1810] = 0;
initial m[1811] = 0;
initial m[1812] = 1;
initial m[1813] = 1;
initial m[1814] = 1;
initial m[1815] = 0;
initial m[1816] = 0;
initial m[1817] = 1;
initial m[1818] = 1;
initial m[1819] = 1;
initial m[1820] = 1;
initial m[1821] = 1;
initial m[1822] = 1;
initial m[1823] = 0;
initial m[1824] = 0;
initial m[1825] = 1;
initial m[1826] = 0;
initial m[1827] = 0;
initial m[1828] = 0;
initial m[1829] = 1;
initial m[1830] = 0;
initial m[1831] = 0;
initial m[1832] = 1;
initial m[1833] = 1;
initial m[1834] = 0;
initial m[1835] = 0;
initial m[1836] = 1;
initial m[1837] = 1;
initial m[1838] = 0;
initial m[1839] = 0;
initial m[1840] = 1;
initial m[1841] = 1;
initial m[1842] = 0;
initial m[1843] = 0;
initial m[1844] = 1;
initial m[1845] = 0;
initial m[1846] = 1;
initial m[1847] = 1;
initial m[1848] = 0;
initial m[1849] = 0;
initial m[1850] = 1;
initial m[1852] = 1;
initial m[1853] = 1;
initial m[1854] = 0;
initial m[1855] = 1;
initial m[1856] = 0;
initial m[1857] = 0;
initial m[1858] = 1;
initial m[1859] = 0;
initial m[1860] = 0;
initial m[1861] = 0;
initial m[1862] = 1;
initial m[1863] = 0;
initial m[1864] = 0;
initial m[1865] = 1;
initial m[1866] = 1;
initial m[1867] = 1;
initial m[1868] = 1;
initial m[1869] = 0;
initial m[1870] = 0;
initial m[1871] = 1;
initial m[1872] = 1;
initial m[1873] = 0;
initial m[1874] = 0;
initial m[1875] = 0;
initial m[1876] = 0;
initial m[1877] = 0;
initial m[1878] = 1;
initial m[1879] = 1;
initial m[1880] = 0;
initial m[1881] = 0;
initial m[1882] = 1;
initial m[1883] = 0;
initial m[1884] = 0;
initial m[1885] = 0;
initial m[1886] = 0;
initial m[1887] = 0;
initial m[1888] = 0;
initial m[1889] = 1;
initial m[1890] = 1;
initial m[1891] = 1;
initial m[1892] = 1;
initial m[1893] = 0;
initial m[1894] = 0;
initial m[1895] = 0;
initial m[1896] = 1;
initial m[1897] = 1;
initial m[1898] = 1;
initial m[1899] = 1;
initial m[1900] = 0;
initial m[1902] = 0;
initial m[1903] = 1;
initial m[1904] = 0;
initial m[1905] = 1;
initial m[1906] = 1;
initial m[1907] = 0;
initial m[1908] = 0;
initial m[1909] = 1;
initial m[1910] = 0;
initial m[1911] = 0;
initial m[1912] = 1;
initial m[1913] = 0;
initial m[1914] = 1;
initial m[1915] = 0;
initial m[1916] = 0;
initial m[1917] = 0;
initial m[1918] = 1;
initial m[1919] = 0;
initial m[1920] = 1;
initial m[1921] = 0;
initial m[1922] = 0;
initial m[1923] = 1;
initial m[1924] = 0;
initial m[1925] = 1;
initial m[1926] = 1;
initial m[1927] = 1;
initial m[1928] = 0;
initial m[1929] = 1;
initial m[1930] = 0;
initial m[1931] = 0;
initial m[1932] = 1;
initial m[1933] = 1;
initial m[1934] = 1;
initial m[1935] = 0;
initial m[1936] = 0;
initial m[1937] = 0;
initial m[1938] = 0;
initial m[1939] = 0;
initial m[1940] = 1;
initial m[1941] = 1;
initial m[1942] = 1;
initial m[1943] = 1;
initial m[1944] = 0;
initial m[1945] = 1;
initial m[1947] = 1;
initial m[1948] = 1;
initial m[1949] = 1;
initial m[1950] = 1;
initial m[1951] = 0;
initial m[1952] = 0;
initial m[1953] = 0;
initial m[1954] = 1;
initial m[1955] = 1;
initial m[1956] = 1;
initial m[1957] = 0;
initial m[1958] = 1;
initial m[1959] = 0;
initial m[1960] = 0;
initial m[1961] = 0;
initial m[1962] = 0;
initial m[1963] = 1;
initial m[1964] = 0;
initial m[1965] = 0;
initial m[1966] = 0;
initial m[1967] = 0;
initial m[1968] = 1;
initial m[1969] = 1;
initial m[1970] = 0;
initial m[1971] = 0;
initial m[1972] = 0;
initial m[1973] = 0;
initial m[1974] = 0;
initial m[1975] = 0;
initial m[1976] = 1;
initial m[1977] = 1;
initial m[1978] = 0;
initial m[1979] = 0;
initial m[1980] = 1;
initial m[1981] = 0;
initial m[1982] = 0;
initial m[1983] = 0;
initial m[1984] = 0;
initial m[1985] = 0;
initial m[1987] = 1;
initial m[1988] = 0;
initial m[1989] = 1;
initial m[1990] = 0;
initial m[1991] = 0;
initial m[1992] = 0;
initial m[1993] = 0;
initial m[1994] = 0;
initial m[1995] = 1;
initial m[1996] = 0;
initial m[1997] = 0;
initial m[1998] = 1;
initial m[1999] = 1;
initial m[2000] = 0;
initial m[2001] = 1;
initial m[2002] = 0;
initial m[2003] = 0;
initial m[2004] = 1;
initial m[2005] = 1;
initial m[2006] = 1;
initial m[2007] = 1;
initial m[2008] = 0;
initial m[2009] = 1;
initial m[2010] = 1;
initial m[2011] = 1;
initial m[2012] = 1;
initial m[2013] = 0;
initial m[2014] = 1;
initial m[2015] = 0;
initial m[2016] = 1;
initial m[2017] = 1;
initial m[2018] = 0;
initial m[2019] = 1;
initial m[2020] = 1;
initial m[2022] = 0;
initial m[2023] = 1;
initial m[2024] = 0;
initial m[2025] = 0;
initial m[2026] = 1;
initial m[2027] = 0;
initial m[2028] = 0;
initial m[2029] = 0;
initial m[2030] = 0;
initial m[2031] = 0;
initial m[2032] = 1;
initial m[2033] = 0;
initial m[2034] = 0;
initial m[2035] = 1;
initial m[2036] = 0;
initial m[2037] = 0;
initial m[2038] = 0;
initial m[2039] = 0;
initial m[2040] = 1;
initial m[2041] = 0;
initial m[2042] = 0;
initial m[2043] = 0;
initial m[2044] = 1;
initial m[2045] = 1;
initial m[2046] = 1;
initial m[2047] = 1;
initial m[2048] = 1;
initial m[2049] = 1;
initial m[2050] = 1;
initial m[2052] = 1;
initial m[2053] = 0;
initial m[2054] = 0;
initial m[2055] = 1;
initial m[2056] = 1;
initial m[2057] = 1;
initial m[2058] = 1;
initial m[2059] = 0;
initial m[2060] = 1;
initial m[2061] = 0;
initial m[2062] = 1;
initial m[2063] = 0;
initial m[2064] = 0;
initial m[2065] = 1;
initial m[2066] = 0;
initial m[2067] = 1;
initial m[2068] = 1;
initial m[2069] = 0;
initial m[2070] = 0;
initial m[2071] = 0;
initial m[2072] = 0;
initial m[2073] = 0;
initial m[2074] = 1;
initial m[2075] = 0;
initial m[2077] = 0;
initial m[2078] = 0;
initial m[2079] = 1;
initial m[2080] = 0;
initial m[2081] = 0;
initial m[2082] = 0;
initial m[2083] = 1;
initial m[2084] = 0;
initial m[2085] = 1;
initial m[2086] = 1;
initial m[2087] = 0;
initial m[2088] = 0;
initial m[2089] = 0;
initial m[2090] = 0;
initial m[2091] = 0;
initial m[2092] = 0;
initial m[2093] = 0;
initial m[2094] = 1;
initial m[2095] = 0;
initial m[2097] = 1;
initial m[2098] = 1;
initial m[2099] = 1;
initial m[2100] = 0;
initial m[2101] = 1;
initial m[2102] = 1;
initial m[2103] = 0;
initial m[2104] = 1;
initial m[2105] = 0;
initial m[2106] = 1;
initial m[2107] = 1;
initial m[2108] = 1;
initial m[2109] = 1;
initial m[2110] = 1;
initial m[2112] = 1;
initial m[2113] = 0;
initial m[2114] = 0;
initial m[2115] = 1;
initial m[2116] = 0;
initial m[2117] = 0;
initial m[2118] = 0;
initial m[2119] = 0;
initial m[2120] = 1;
initial m[2122] = 0;
initial m[2123] = 0;
initial m[2124] = 0;
initial m[2125] = 0;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[15],m[14],m[13],m[12],m[11],m[10],m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[31],m[30],m[29],m[28],m[27],m[26],m[25],m[24],m[23],m[22],m[21],m[20],m[19],m[18],m[17],m[16]};
end

always @(negedge sample_clk) begin
    if (solution == 32'b11101011101110010100001101010001)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[32]&m[33]&~m[34]&~m[35])|(m[32]&~m[33]&m[34]&~m[35])|(~m[32]&m[33]&m[34]&~m[35])|(m[32]&~m[33]&~m[34]&m[35])|(~m[32]&m[33]&~m[34]&m[35])|(~m[32]&~m[33]&m[34]&m[35]))&UnbiasedRNG[0])|((m[32]&m[33]&m[34]&~m[35])|(m[32]&m[33]&~m[34]&m[35])|(m[32]&~m[33]&m[34]&m[35])|(~m[32]&m[33]&m[34]&m[35])|(m[32]&m[33]&m[34]&m[35]));
    m[1] = (((m[36]&m[37]&~m[38]&~m[39])|(m[36]&~m[37]&m[38]&~m[39])|(~m[36]&m[37]&m[38]&~m[39])|(m[36]&~m[37]&~m[38]&m[39])|(~m[36]&m[37]&~m[38]&m[39])|(~m[36]&~m[37]&m[38]&m[39]))&UnbiasedRNG[1])|((m[36]&m[37]&m[38]&~m[39])|(m[36]&m[37]&~m[38]&m[39])|(m[36]&~m[37]&m[38]&m[39])|(~m[36]&m[37]&m[38]&m[39])|(m[36]&m[37]&m[38]&m[39]));
    m[2] = (((m[40]&m[41]&~m[42]&~m[43])|(m[40]&~m[41]&m[42]&~m[43])|(~m[40]&m[41]&m[42]&~m[43])|(m[40]&~m[41]&~m[42]&m[43])|(~m[40]&m[41]&~m[42]&m[43])|(~m[40]&~m[41]&m[42]&m[43]))&UnbiasedRNG[2])|((m[40]&m[41]&m[42]&~m[43])|(m[40]&m[41]&~m[42]&m[43])|(m[40]&~m[41]&m[42]&m[43])|(~m[40]&m[41]&m[42]&m[43])|(m[40]&m[41]&m[42]&m[43]));
    m[3] = (((m[44]&m[45]&~m[46]&~m[47])|(m[44]&~m[45]&m[46]&~m[47])|(~m[44]&m[45]&m[46]&~m[47])|(m[44]&~m[45]&~m[46]&m[47])|(~m[44]&m[45]&~m[46]&m[47])|(~m[44]&~m[45]&m[46]&m[47]))&UnbiasedRNG[3])|((m[44]&m[45]&m[46]&~m[47])|(m[44]&m[45]&~m[46]&m[47])|(m[44]&~m[45]&m[46]&m[47])|(~m[44]&m[45]&m[46]&m[47])|(m[44]&m[45]&m[46]&m[47]));
    m[4] = (((m[48]&m[49]&~m[50]&~m[51])|(m[48]&~m[49]&m[50]&~m[51])|(~m[48]&m[49]&m[50]&~m[51])|(m[48]&~m[49]&~m[50]&m[51])|(~m[48]&m[49]&~m[50]&m[51])|(~m[48]&~m[49]&m[50]&m[51]))&UnbiasedRNG[4])|((m[48]&m[49]&m[50]&~m[51])|(m[48]&m[49]&~m[50]&m[51])|(m[48]&~m[49]&m[50]&m[51])|(~m[48]&m[49]&m[50]&m[51])|(m[48]&m[49]&m[50]&m[51]));
    m[5] = (((m[52]&m[53]&~m[54]&~m[55])|(m[52]&~m[53]&m[54]&~m[55])|(~m[52]&m[53]&m[54]&~m[55])|(m[52]&~m[53]&~m[54]&m[55])|(~m[52]&m[53]&~m[54]&m[55])|(~m[52]&~m[53]&m[54]&m[55]))&UnbiasedRNG[5])|((m[52]&m[53]&m[54]&~m[55])|(m[52]&m[53]&~m[54]&m[55])|(m[52]&~m[53]&m[54]&m[55])|(~m[52]&m[53]&m[54]&m[55])|(m[52]&m[53]&m[54]&m[55]));
    m[6] = (((m[56]&m[57]&~m[58]&~m[59])|(m[56]&~m[57]&m[58]&~m[59])|(~m[56]&m[57]&m[58]&~m[59])|(m[56]&~m[57]&~m[58]&m[59])|(~m[56]&m[57]&~m[58]&m[59])|(~m[56]&~m[57]&m[58]&m[59]))&UnbiasedRNG[6])|((m[56]&m[57]&m[58]&~m[59])|(m[56]&m[57]&~m[58]&m[59])|(m[56]&~m[57]&m[58]&m[59])|(~m[56]&m[57]&m[58]&m[59])|(m[56]&m[57]&m[58]&m[59]));
    m[7] = (((m[60]&m[61]&~m[62]&~m[63])|(m[60]&~m[61]&m[62]&~m[63])|(~m[60]&m[61]&m[62]&~m[63])|(m[60]&~m[61]&~m[62]&m[63])|(~m[60]&m[61]&~m[62]&m[63])|(~m[60]&~m[61]&m[62]&m[63]))&UnbiasedRNG[7])|((m[60]&m[61]&m[62]&~m[63])|(m[60]&m[61]&~m[62]&m[63])|(m[60]&~m[61]&m[62]&m[63])|(~m[60]&m[61]&m[62]&m[63])|(m[60]&m[61]&m[62]&m[63]));
    m[8] = (((m[64]&m[65]&~m[66]&~m[67])|(m[64]&~m[65]&m[66]&~m[67])|(~m[64]&m[65]&m[66]&~m[67])|(m[64]&~m[65]&~m[66]&m[67])|(~m[64]&m[65]&~m[66]&m[67])|(~m[64]&~m[65]&m[66]&m[67]))&UnbiasedRNG[8])|((m[64]&m[65]&m[66]&~m[67])|(m[64]&m[65]&~m[66]&m[67])|(m[64]&~m[65]&m[66]&m[67])|(~m[64]&m[65]&m[66]&m[67])|(m[64]&m[65]&m[66]&m[67]));
    m[9] = (((m[68]&m[69]&~m[70]&~m[71])|(m[68]&~m[69]&m[70]&~m[71])|(~m[68]&m[69]&m[70]&~m[71])|(m[68]&~m[69]&~m[70]&m[71])|(~m[68]&m[69]&~m[70]&m[71])|(~m[68]&~m[69]&m[70]&m[71]))&UnbiasedRNG[9])|((m[68]&m[69]&m[70]&~m[71])|(m[68]&m[69]&~m[70]&m[71])|(m[68]&~m[69]&m[70]&m[71])|(~m[68]&m[69]&m[70]&m[71])|(m[68]&m[69]&m[70]&m[71]));
    m[10] = (((m[72]&m[73]&~m[74]&~m[75])|(m[72]&~m[73]&m[74]&~m[75])|(~m[72]&m[73]&m[74]&~m[75])|(m[72]&~m[73]&~m[74]&m[75])|(~m[72]&m[73]&~m[74]&m[75])|(~m[72]&~m[73]&m[74]&m[75]))&UnbiasedRNG[10])|((m[72]&m[73]&m[74]&~m[75])|(m[72]&m[73]&~m[74]&m[75])|(m[72]&~m[73]&m[74]&m[75])|(~m[72]&m[73]&m[74]&m[75])|(m[72]&m[73]&m[74]&m[75]));
    m[11] = (((m[76]&m[77]&~m[78]&~m[79])|(m[76]&~m[77]&m[78]&~m[79])|(~m[76]&m[77]&m[78]&~m[79])|(m[76]&~m[77]&~m[78]&m[79])|(~m[76]&m[77]&~m[78]&m[79])|(~m[76]&~m[77]&m[78]&m[79]))&UnbiasedRNG[11])|((m[76]&m[77]&m[78]&~m[79])|(m[76]&m[77]&~m[78]&m[79])|(m[76]&~m[77]&m[78]&m[79])|(~m[76]&m[77]&m[78]&m[79])|(m[76]&m[77]&m[78]&m[79]));
    m[12] = (((m[80]&m[81]&~m[82]&~m[83])|(m[80]&~m[81]&m[82]&~m[83])|(~m[80]&m[81]&m[82]&~m[83])|(m[80]&~m[81]&~m[82]&m[83])|(~m[80]&m[81]&~m[82]&m[83])|(~m[80]&~m[81]&m[82]&m[83]))&UnbiasedRNG[12])|((m[80]&m[81]&m[82]&~m[83])|(m[80]&m[81]&~m[82]&m[83])|(m[80]&~m[81]&m[82]&m[83])|(~m[80]&m[81]&m[82]&m[83])|(m[80]&m[81]&m[82]&m[83]));
    m[13] = (((m[84]&m[85]&~m[86]&~m[87])|(m[84]&~m[85]&m[86]&~m[87])|(~m[84]&m[85]&m[86]&~m[87])|(m[84]&~m[85]&~m[86]&m[87])|(~m[84]&m[85]&~m[86]&m[87])|(~m[84]&~m[85]&m[86]&m[87]))&UnbiasedRNG[13])|((m[84]&m[85]&m[86]&~m[87])|(m[84]&m[85]&~m[86]&m[87])|(m[84]&~m[85]&m[86]&m[87])|(~m[84]&m[85]&m[86]&m[87])|(m[84]&m[85]&m[86]&m[87]));
    m[14] = (((m[88]&m[89]&~m[90]&~m[91])|(m[88]&~m[89]&m[90]&~m[91])|(~m[88]&m[89]&m[90]&~m[91])|(m[88]&~m[89]&~m[90]&m[91])|(~m[88]&m[89]&~m[90]&m[91])|(~m[88]&~m[89]&m[90]&m[91]))&UnbiasedRNG[14])|((m[88]&m[89]&m[90]&~m[91])|(m[88]&m[89]&~m[90]&m[91])|(m[88]&~m[89]&m[90]&m[91])|(~m[88]&m[89]&m[90]&m[91])|(m[88]&m[89]&m[90]&m[91]));
    m[15] = (((m[92]&m[93]&~m[94]&~m[95])|(m[92]&~m[93]&m[94]&~m[95])|(~m[92]&m[93]&m[94]&~m[95])|(m[92]&~m[93]&~m[94]&m[95])|(~m[92]&m[93]&~m[94]&m[95])|(~m[92]&~m[93]&m[94]&m[95]))&UnbiasedRNG[15])|((m[92]&m[93]&m[94]&~m[95])|(m[92]&m[93]&~m[94]&m[95])|(m[92]&~m[93]&m[94]&m[95])|(~m[92]&m[93]&m[94]&m[95])|(m[92]&m[93]&m[94]&m[95]));
    m[16] = (((m[96]&m[97]&~m[98]&~m[99])|(m[96]&~m[97]&m[98]&~m[99])|(~m[96]&m[97]&m[98]&~m[99])|(m[96]&~m[97]&~m[98]&m[99])|(~m[96]&m[97]&~m[98]&m[99])|(~m[96]&~m[97]&m[98]&m[99]))&UnbiasedRNG[16])|((m[96]&m[97]&m[98]&~m[99])|(m[96]&m[97]&~m[98]&m[99])|(m[96]&~m[97]&m[98]&m[99])|(~m[96]&m[97]&m[98]&m[99])|(m[96]&m[97]&m[98]&m[99]));
    m[17] = (((m[100]&m[101]&~m[102]&~m[103])|(m[100]&~m[101]&m[102]&~m[103])|(~m[100]&m[101]&m[102]&~m[103])|(m[100]&~m[101]&~m[102]&m[103])|(~m[100]&m[101]&~m[102]&m[103])|(~m[100]&~m[101]&m[102]&m[103]))&UnbiasedRNG[17])|((m[100]&m[101]&m[102]&~m[103])|(m[100]&m[101]&~m[102]&m[103])|(m[100]&~m[101]&m[102]&m[103])|(~m[100]&m[101]&m[102]&m[103])|(m[100]&m[101]&m[102]&m[103]));
    m[18] = (((m[104]&m[105]&~m[106]&~m[107])|(m[104]&~m[105]&m[106]&~m[107])|(~m[104]&m[105]&m[106]&~m[107])|(m[104]&~m[105]&~m[106]&m[107])|(~m[104]&m[105]&~m[106]&m[107])|(~m[104]&~m[105]&m[106]&m[107]))&UnbiasedRNG[18])|((m[104]&m[105]&m[106]&~m[107])|(m[104]&m[105]&~m[106]&m[107])|(m[104]&~m[105]&m[106]&m[107])|(~m[104]&m[105]&m[106]&m[107])|(m[104]&m[105]&m[106]&m[107]));
    m[19] = (((m[108]&m[109]&~m[110]&~m[111])|(m[108]&~m[109]&m[110]&~m[111])|(~m[108]&m[109]&m[110]&~m[111])|(m[108]&~m[109]&~m[110]&m[111])|(~m[108]&m[109]&~m[110]&m[111])|(~m[108]&~m[109]&m[110]&m[111]))&UnbiasedRNG[19])|((m[108]&m[109]&m[110]&~m[111])|(m[108]&m[109]&~m[110]&m[111])|(m[108]&~m[109]&m[110]&m[111])|(~m[108]&m[109]&m[110]&m[111])|(m[108]&m[109]&m[110]&m[111]));
    m[20] = (((m[112]&m[113]&~m[114]&~m[115])|(m[112]&~m[113]&m[114]&~m[115])|(~m[112]&m[113]&m[114]&~m[115])|(m[112]&~m[113]&~m[114]&m[115])|(~m[112]&m[113]&~m[114]&m[115])|(~m[112]&~m[113]&m[114]&m[115]))&UnbiasedRNG[20])|((m[112]&m[113]&m[114]&~m[115])|(m[112]&m[113]&~m[114]&m[115])|(m[112]&~m[113]&m[114]&m[115])|(~m[112]&m[113]&m[114]&m[115])|(m[112]&m[113]&m[114]&m[115]));
    m[21] = (((m[116]&m[117]&~m[118]&~m[119])|(m[116]&~m[117]&m[118]&~m[119])|(~m[116]&m[117]&m[118]&~m[119])|(m[116]&~m[117]&~m[118]&m[119])|(~m[116]&m[117]&~m[118]&m[119])|(~m[116]&~m[117]&m[118]&m[119]))&UnbiasedRNG[21])|((m[116]&m[117]&m[118]&~m[119])|(m[116]&m[117]&~m[118]&m[119])|(m[116]&~m[117]&m[118]&m[119])|(~m[116]&m[117]&m[118]&m[119])|(m[116]&m[117]&m[118]&m[119]));
    m[22] = (((m[120]&m[121]&~m[122]&~m[123])|(m[120]&~m[121]&m[122]&~m[123])|(~m[120]&m[121]&m[122]&~m[123])|(m[120]&~m[121]&~m[122]&m[123])|(~m[120]&m[121]&~m[122]&m[123])|(~m[120]&~m[121]&m[122]&m[123]))&UnbiasedRNG[22])|((m[120]&m[121]&m[122]&~m[123])|(m[120]&m[121]&~m[122]&m[123])|(m[120]&~m[121]&m[122]&m[123])|(~m[120]&m[121]&m[122]&m[123])|(m[120]&m[121]&m[122]&m[123]));
    m[23] = (((m[124]&m[125]&~m[126]&~m[127])|(m[124]&~m[125]&m[126]&~m[127])|(~m[124]&m[125]&m[126]&~m[127])|(m[124]&~m[125]&~m[126]&m[127])|(~m[124]&m[125]&~m[126]&m[127])|(~m[124]&~m[125]&m[126]&m[127]))&UnbiasedRNG[23])|((m[124]&m[125]&m[126]&~m[127])|(m[124]&m[125]&~m[126]&m[127])|(m[124]&~m[125]&m[126]&m[127])|(~m[124]&m[125]&m[126]&m[127])|(m[124]&m[125]&m[126]&m[127]));
    m[24] = (((m[128]&m[129]&~m[130]&~m[131])|(m[128]&~m[129]&m[130]&~m[131])|(~m[128]&m[129]&m[130]&~m[131])|(m[128]&~m[129]&~m[130]&m[131])|(~m[128]&m[129]&~m[130]&m[131])|(~m[128]&~m[129]&m[130]&m[131]))&UnbiasedRNG[24])|((m[128]&m[129]&m[130]&~m[131])|(m[128]&m[129]&~m[130]&m[131])|(m[128]&~m[129]&m[130]&m[131])|(~m[128]&m[129]&m[130]&m[131])|(m[128]&m[129]&m[130]&m[131]));
    m[25] = (((m[132]&m[133]&~m[134]&~m[135])|(m[132]&~m[133]&m[134]&~m[135])|(~m[132]&m[133]&m[134]&~m[135])|(m[132]&~m[133]&~m[134]&m[135])|(~m[132]&m[133]&~m[134]&m[135])|(~m[132]&~m[133]&m[134]&m[135]))&UnbiasedRNG[25])|((m[132]&m[133]&m[134]&~m[135])|(m[132]&m[133]&~m[134]&m[135])|(m[132]&~m[133]&m[134]&m[135])|(~m[132]&m[133]&m[134]&m[135])|(m[132]&m[133]&m[134]&m[135]));
    m[26] = (((m[136]&m[137]&~m[138]&~m[139])|(m[136]&~m[137]&m[138]&~m[139])|(~m[136]&m[137]&m[138]&~m[139])|(m[136]&~m[137]&~m[138]&m[139])|(~m[136]&m[137]&~m[138]&m[139])|(~m[136]&~m[137]&m[138]&m[139]))&UnbiasedRNG[26])|((m[136]&m[137]&m[138]&~m[139])|(m[136]&m[137]&~m[138]&m[139])|(m[136]&~m[137]&m[138]&m[139])|(~m[136]&m[137]&m[138]&m[139])|(m[136]&m[137]&m[138]&m[139]));
    m[27] = (((m[140]&m[141]&~m[142]&~m[143])|(m[140]&~m[141]&m[142]&~m[143])|(~m[140]&m[141]&m[142]&~m[143])|(m[140]&~m[141]&~m[142]&m[143])|(~m[140]&m[141]&~m[142]&m[143])|(~m[140]&~m[141]&m[142]&m[143]))&UnbiasedRNG[27])|((m[140]&m[141]&m[142]&~m[143])|(m[140]&m[141]&~m[142]&m[143])|(m[140]&~m[141]&m[142]&m[143])|(~m[140]&m[141]&m[142]&m[143])|(m[140]&m[141]&m[142]&m[143]));
    m[28] = (((m[144]&m[145]&~m[146]&~m[147])|(m[144]&~m[145]&m[146]&~m[147])|(~m[144]&m[145]&m[146]&~m[147])|(m[144]&~m[145]&~m[146]&m[147])|(~m[144]&m[145]&~m[146]&m[147])|(~m[144]&~m[145]&m[146]&m[147]))&UnbiasedRNG[28])|((m[144]&m[145]&m[146]&~m[147])|(m[144]&m[145]&~m[146]&m[147])|(m[144]&~m[145]&m[146]&m[147])|(~m[144]&m[145]&m[146]&m[147])|(m[144]&m[145]&m[146]&m[147]));
    m[29] = (((m[148]&m[149]&~m[150]&~m[151])|(m[148]&~m[149]&m[150]&~m[151])|(~m[148]&m[149]&m[150]&~m[151])|(m[148]&~m[149]&~m[150]&m[151])|(~m[148]&m[149]&~m[150]&m[151])|(~m[148]&~m[149]&m[150]&m[151]))&UnbiasedRNG[29])|((m[148]&m[149]&m[150]&~m[151])|(m[148]&m[149]&~m[150]&m[151])|(m[148]&~m[149]&m[150]&m[151])|(~m[148]&m[149]&m[150]&m[151])|(m[148]&m[149]&m[150]&m[151]));
    m[30] = (((m[152]&m[153]&~m[154]&~m[155])|(m[152]&~m[153]&m[154]&~m[155])|(~m[152]&m[153]&m[154]&~m[155])|(m[152]&~m[153]&~m[154]&m[155])|(~m[152]&m[153]&~m[154]&m[155])|(~m[152]&~m[153]&m[154]&m[155]))&UnbiasedRNG[30])|((m[152]&m[153]&m[154]&~m[155])|(m[152]&m[153]&~m[154]&m[155])|(m[152]&~m[153]&m[154]&m[155])|(~m[152]&m[153]&m[154]&m[155])|(m[152]&m[153]&m[154]&m[155]));
    m[31] = (((m[156]&m[157]&~m[158]&~m[159])|(m[156]&~m[157]&m[158]&~m[159])|(~m[156]&m[157]&m[158]&~m[159])|(m[156]&~m[157]&~m[158]&m[159])|(~m[156]&m[157]&~m[158]&m[159])|(~m[156]&~m[157]&m[158]&m[159]))&UnbiasedRNG[31])|((m[156]&m[157]&m[158]&~m[159])|(m[156]&m[157]&~m[158]&m[159])|(m[156]&~m[157]&m[158]&m[159])|(~m[156]&m[157]&m[158]&m[159])|(m[156]&m[157]&m[158]&m[159]));
    m[160] = (((~m[32]&~m[416]&~m[672])|(m[32]&m[416]&~m[672]))&BiasedRNG[0])|(((m[32]&~m[416]&~m[672])|(~m[32]&m[416]&m[672]))&~BiasedRNG[0])|((~m[32]&~m[416]&m[672])|(m[32]&~m[416]&m[672])|(m[32]&m[416]&m[672]));
    m[161] = (((~m[32]&~m[432]&~m[688])|(m[32]&m[432]&~m[688]))&BiasedRNG[1])|(((m[32]&~m[432]&~m[688])|(~m[32]&m[432]&m[688]))&~BiasedRNG[1])|((~m[32]&~m[432]&m[688])|(m[32]&~m[432]&m[688])|(m[32]&m[432]&m[688]));
    m[162] = (((~m[32]&~m[448]&~m[704])|(m[32]&m[448]&~m[704]))&BiasedRNG[2])|(((m[32]&~m[448]&~m[704])|(~m[32]&m[448]&m[704]))&~BiasedRNG[2])|((~m[32]&~m[448]&m[704])|(m[32]&~m[448]&m[704])|(m[32]&m[448]&m[704]));
    m[163] = (((~m[32]&~m[464]&~m[720])|(m[32]&m[464]&~m[720]))&BiasedRNG[3])|(((m[32]&~m[464]&~m[720])|(~m[32]&m[464]&m[720]))&~BiasedRNG[3])|((~m[32]&~m[464]&m[720])|(m[32]&~m[464]&m[720])|(m[32]&m[464]&m[720]));
    m[164] = (((~m[33]&~m[480]&~m[736])|(m[33]&m[480]&~m[736]))&BiasedRNG[4])|(((m[33]&~m[480]&~m[736])|(~m[33]&m[480]&m[736]))&~BiasedRNG[4])|((~m[33]&~m[480]&m[736])|(m[33]&~m[480]&m[736])|(m[33]&m[480]&m[736]));
    m[165] = (((~m[33]&~m[496]&~m[752])|(m[33]&m[496]&~m[752]))&BiasedRNG[5])|(((m[33]&~m[496]&~m[752])|(~m[33]&m[496]&m[752]))&~BiasedRNG[5])|((~m[33]&~m[496]&m[752])|(m[33]&~m[496]&m[752])|(m[33]&m[496]&m[752]));
    m[166] = (((~m[33]&~m[512]&~m[768])|(m[33]&m[512]&~m[768]))&BiasedRNG[6])|(((m[33]&~m[512]&~m[768])|(~m[33]&m[512]&m[768]))&~BiasedRNG[6])|((~m[33]&~m[512]&m[768])|(m[33]&~m[512]&m[768])|(m[33]&m[512]&m[768]));
    m[167] = (((~m[33]&~m[528]&~m[784])|(m[33]&m[528]&~m[784]))&BiasedRNG[7])|(((m[33]&~m[528]&~m[784])|(~m[33]&m[528]&m[784]))&~BiasedRNG[7])|((~m[33]&~m[528]&m[784])|(m[33]&~m[528]&m[784])|(m[33]&m[528]&m[784]));
    m[168] = (((~m[34]&~m[544]&~m[800])|(m[34]&m[544]&~m[800]))&BiasedRNG[8])|(((m[34]&~m[544]&~m[800])|(~m[34]&m[544]&m[800]))&~BiasedRNG[8])|((~m[34]&~m[544]&m[800])|(m[34]&~m[544]&m[800])|(m[34]&m[544]&m[800]));
    m[169] = (((~m[34]&~m[560]&~m[816])|(m[34]&m[560]&~m[816]))&BiasedRNG[9])|(((m[34]&~m[560]&~m[816])|(~m[34]&m[560]&m[816]))&~BiasedRNG[9])|((~m[34]&~m[560]&m[816])|(m[34]&~m[560]&m[816])|(m[34]&m[560]&m[816]));
    m[170] = (((~m[34]&~m[576]&~m[832])|(m[34]&m[576]&~m[832]))&BiasedRNG[10])|(((m[34]&~m[576]&~m[832])|(~m[34]&m[576]&m[832]))&~BiasedRNG[10])|((~m[34]&~m[576]&m[832])|(m[34]&~m[576]&m[832])|(m[34]&m[576]&m[832]));
    m[171] = (((~m[34]&~m[592]&~m[848])|(m[34]&m[592]&~m[848]))&BiasedRNG[11])|(((m[34]&~m[592]&~m[848])|(~m[34]&m[592]&m[848]))&~BiasedRNG[11])|((~m[34]&~m[592]&m[848])|(m[34]&~m[592]&m[848])|(m[34]&m[592]&m[848]));
    m[172] = (((~m[35]&~m[608]&~m[864])|(m[35]&m[608]&~m[864]))&BiasedRNG[12])|(((m[35]&~m[608]&~m[864])|(~m[35]&m[608]&m[864]))&~BiasedRNG[12])|((~m[35]&~m[608]&m[864])|(m[35]&~m[608]&m[864])|(m[35]&m[608]&m[864]));
    m[173] = (((~m[35]&~m[624]&~m[880])|(m[35]&m[624]&~m[880]))&BiasedRNG[13])|(((m[35]&~m[624]&~m[880])|(~m[35]&m[624]&m[880]))&~BiasedRNG[13])|((~m[35]&~m[624]&m[880])|(m[35]&~m[624]&m[880])|(m[35]&m[624]&m[880]));
    m[174] = (((~m[35]&~m[640]&~m[896])|(m[35]&m[640]&~m[896]))&BiasedRNG[14])|(((m[35]&~m[640]&~m[896])|(~m[35]&m[640]&m[896]))&~BiasedRNG[14])|((~m[35]&~m[640]&m[896])|(m[35]&~m[640]&m[896])|(m[35]&m[640]&m[896]));
    m[175] = (((~m[35]&~m[656]&~m[912])|(m[35]&m[656]&~m[912]))&BiasedRNG[15])|(((m[35]&~m[656]&~m[912])|(~m[35]&m[656]&m[912]))&~BiasedRNG[15])|((~m[35]&~m[656]&m[912])|(m[35]&~m[656]&m[912])|(m[35]&m[656]&m[912]));
    m[176] = (((~m[36]&~m[417]&~m[673])|(m[36]&m[417]&~m[673]))&BiasedRNG[16])|(((m[36]&~m[417]&~m[673])|(~m[36]&m[417]&m[673]))&~BiasedRNG[16])|((~m[36]&~m[417]&m[673])|(m[36]&~m[417]&m[673])|(m[36]&m[417]&m[673]));
    m[177] = (((~m[36]&~m[433]&~m[689])|(m[36]&m[433]&~m[689]))&BiasedRNG[17])|(((m[36]&~m[433]&~m[689])|(~m[36]&m[433]&m[689]))&~BiasedRNG[17])|((~m[36]&~m[433]&m[689])|(m[36]&~m[433]&m[689])|(m[36]&m[433]&m[689]));
    m[178] = (((~m[36]&~m[449]&~m[705])|(m[36]&m[449]&~m[705]))&BiasedRNG[18])|(((m[36]&~m[449]&~m[705])|(~m[36]&m[449]&m[705]))&~BiasedRNG[18])|((~m[36]&~m[449]&m[705])|(m[36]&~m[449]&m[705])|(m[36]&m[449]&m[705]));
    m[179] = (((~m[36]&~m[465]&~m[721])|(m[36]&m[465]&~m[721]))&BiasedRNG[19])|(((m[36]&~m[465]&~m[721])|(~m[36]&m[465]&m[721]))&~BiasedRNG[19])|((~m[36]&~m[465]&m[721])|(m[36]&~m[465]&m[721])|(m[36]&m[465]&m[721]));
    m[180] = (((~m[37]&~m[481]&~m[737])|(m[37]&m[481]&~m[737]))&BiasedRNG[20])|(((m[37]&~m[481]&~m[737])|(~m[37]&m[481]&m[737]))&~BiasedRNG[20])|((~m[37]&~m[481]&m[737])|(m[37]&~m[481]&m[737])|(m[37]&m[481]&m[737]));
    m[181] = (((~m[37]&~m[497]&~m[753])|(m[37]&m[497]&~m[753]))&BiasedRNG[21])|(((m[37]&~m[497]&~m[753])|(~m[37]&m[497]&m[753]))&~BiasedRNG[21])|((~m[37]&~m[497]&m[753])|(m[37]&~m[497]&m[753])|(m[37]&m[497]&m[753]));
    m[182] = (((~m[37]&~m[513]&~m[769])|(m[37]&m[513]&~m[769]))&BiasedRNG[22])|(((m[37]&~m[513]&~m[769])|(~m[37]&m[513]&m[769]))&~BiasedRNG[22])|((~m[37]&~m[513]&m[769])|(m[37]&~m[513]&m[769])|(m[37]&m[513]&m[769]));
    m[183] = (((~m[37]&~m[529]&~m[785])|(m[37]&m[529]&~m[785]))&BiasedRNG[23])|(((m[37]&~m[529]&~m[785])|(~m[37]&m[529]&m[785]))&~BiasedRNG[23])|((~m[37]&~m[529]&m[785])|(m[37]&~m[529]&m[785])|(m[37]&m[529]&m[785]));
    m[184] = (((~m[38]&~m[545]&~m[801])|(m[38]&m[545]&~m[801]))&BiasedRNG[24])|(((m[38]&~m[545]&~m[801])|(~m[38]&m[545]&m[801]))&~BiasedRNG[24])|((~m[38]&~m[545]&m[801])|(m[38]&~m[545]&m[801])|(m[38]&m[545]&m[801]));
    m[185] = (((~m[38]&~m[561]&~m[817])|(m[38]&m[561]&~m[817]))&BiasedRNG[25])|(((m[38]&~m[561]&~m[817])|(~m[38]&m[561]&m[817]))&~BiasedRNG[25])|((~m[38]&~m[561]&m[817])|(m[38]&~m[561]&m[817])|(m[38]&m[561]&m[817]));
    m[186] = (((~m[38]&~m[577]&~m[833])|(m[38]&m[577]&~m[833]))&BiasedRNG[26])|(((m[38]&~m[577]&~m[833])|(~m[38]&m[577]&m[833]))&~BiasedRNG[26])|((~m[38]&~m[577]&m[833])|(m[38]&~m[577]&m[833])|(m[38]&m[577]&m[833]));
    m[187] = (((~m[38]&~m[593]&~m[849])|(m[38]&m[593]&~m[849]))&BiasedRNG[27])|(((m[38]&~m[593]&~m[849])|(~m[38]&m[593]&m[849]))&~BiasedRNG[27])|((~m[38]&~m[593]&m[849])|(m[38]&~m[593]&m[849])|(m[38]&m[593]&m[849]));
    m[188] = (((~m[39]&~m[609]&~m[865])|(m[39]&m[609]&~m[865]))&BiasedRNG[28])|(((m[39]&~m[609]&~m[865])|(~m[39]&m[609]&m[865]))&~BiasedRNG[28])|((~m[39]&~m[609]&m[865])|(m[39]&~m[609]&m[865])|(m[39]&m[609]&m[865]));
    m[189] = (((~m[39]&~m[625]&~m[881])|(m[39]&m[625]&~m[881]))&BiasedRNG[29])|(((m[39]&~m[625]&~m[881])|(~m[39]&m[625]&m[881]))&~BiasedRNG[29])|((~m[39]&~m[625]&m[881])|(m[39]&~m[625]&m[881])|(m[39]&m[625]&m[881]));
    m[190] = (((~m[39]&~m[641]&~m[897])|(m[39]&m[641]&~m[897]))&BiasedRNG[30])|(((m[39]&~m[641]&~m[897])|(~m[39]&m[641]&m[897]))&~BiasedRNG[30])|((~m[39]&~m[641]&m[897])|(m[39]&~m[641]&m[897])|(m[39]&m[641]&m[897]));
    m[191] = (((~m[39]&~m[657]&~m[913])|(m[39]&m[657]&~m[913]))&BiasedRNG[31])|(((m[39]&~m[657]&~m[913])|(~m[39]&m[657]&m[913]))&~BiasedRNG[31])|((~m[39]&~m[657]&m[913])|(m[39]&~m[657]&m[913])|(m[39]&m[657]&m[913]));
    m[192] = (((~m[40]&~m[418]&~m[674])|(m[40]&m[418]&~m[674]))&BiasedRNG[32])|(((m[40]&~m[418]&~m[674])|(~m[40]&m[418]&m[674]))&~BiasedRNG[32])|((~m[40]&~m[418]&m[674])|(m[40]&~m[418]&m[674])|(m[40]&m[418]&m[674]));
    m[193] = (((~m[40]&~m[434]&~m[690])|(m[40]&m[434]&~m[690]))&BiasedRNG[33])|(((m[40]&~m[434]&~m[690])|(~m[40]&m[434]&m[690]))&~BiasedRNG[33])|((~m[40]&~m[434]&m[690])|(m[40]&~m[434]&m[690])|(m[40]&m[434]&m[690]));
    m[194] = (((~m[40]&~m[450]&~m[706])|(m[40]&m[450]&~m[706]))&BiasedRNG[34])|(((m[40]&~m[450]&~m[706])|(~m[40]&m[450]&m[706]))&~BiasedRNG[34])|((~m[40]&~m[450]&m[706])|(m[40]&~m[450]&m[706])|(m[40]&m[450]&m[706]));
    m[195] = (((~m[40]&~m[466]&~m[722])|(m[40]&m[466]&~m[722]))&BiasedRNG[35])|(((m[40]&~m[466]&~m[722])|(~m[40]&m[466]&m[722]))&~BiasedRNG[35])|((~m[40]&~m[466]&m[722])|(m[40]&~m[466]&m[722])|(m[40]&m[466]&m[722]));
    m[196] = (((~m[41]&~m[482]&~m[738])|(m[41]&m[482]&~m[738]))&BiasedRNG[36])|(((m[41]&~m[482]&~m[738])|(~m[41]&m[482]&m[738]))&~BiasedRNG[36])|((~m[41]&~m[482]&m[738])|(m[41]&~m[482]&m[738])|(m[41]&m[482]&m[738]));
    m[197] = (((~m[41]&~m[498]&~m[754])|(m[41]&m[498]&~m[754]))&BiasedRNG[37])|(((m[41]&~m[498]&~m[754])|(~m[41]&m[498]&m[754]))&~BiasedRNG[37])|((~m[41]&~m[498]&m[754])|(m[41]&~m[498]&m[754])|(m[41]&m[498]&m[754]));
    m[198] = (((~m[41]&~m[514]&~m[770])|(m[41]&m[514]&~m[770]))&BiasedRNG[38])|(((m[41]&~m[514]&~m[770])|(~m[41]&m[514]&m[770]))&~BiasedRNG[38])|((~m[41]&~m[514]&m[770])|(m[41]&~m[514]&m[770])|(m[41]&m[514]&m[770]));
    m[199] = (((~m[41]&~m[530]&~m[786])|(m[41]&m[530]&~m[786]))&BiasedRNG[39])|(((m[41]&~m[530]&~m[786])|(~m[41]&m[530]&m[786]))&~BiasedRNG[39])|((~m[41]&~m[530]&m[786])|(m[41]&~m[530]&m[786])|(m[41]&m[530]&m[786]));
    m[200] = (((~m[42]&~m[546]&~m[802])|(m[42]&m[546]&~m[802]))&BiasedRNG[40])|(((m[42]&~m[546]&~m[802])|(~m[42]&m[546]&m[802]))&~BiasedRNG[40])|((~m[42]&~m[546]&m[802])|(m[42]&~m[546]&m[802])|(m[42]&m[546]&m[802]));
    m[201] = (((~m[42]&~m[562]&~m[818])|(m[42]&m[562]&~m[818]))&BiasedRNG[41])|(((m[42]&~m[562]&~m[818])|(~m[42]&m[562]&m[818]))&~BiasedRNG[41])|((~m[42]&~m[562]&m[818])|(m[42]&~m[562]&m[818])|(m[42]&m[562]&m[818]));
    m[202] = (((~m[42]&~m[578]&~m[834])|(m[42]&m[578]&~m[834]))&BiasedRNG[42])|(((m[42]&~m[578]&~m[834])|(~m[42]&m[578]&m[834]))&~BiasedRNG[42])|((~m[42]&~m[578]&m[834])|(m[42]&~m[578]&m[834])|(m[42]&m[578]&m[834]));
    m[203] = (((~m[42]&~m[594]&~m[850])|(m[42]&m[594]&~m[850]))&BiasedRNG[43])|(((m[42]&~m[594]&~m[850])|(~m[42]&m[594]&m[850]))&~BiasedRNG[43])|((~m[42]&~m[594]&m[850])|(m[42]&~m[594]&m[850])|(m[42]&m[594]&m[850]));
    m[204] = (((~m[43]&~m[610]&~m[866])|(m[43]&m[610]&~m[866]))&BiasedRNG[44])|(((m[43]&~m[610]&~m[866])|(~m[43]&m[610]&m[866]))&~BiasedRNG[44])|((~m[43]&~m[610]&m[866])|(m[43]&~m[610]&m[866])|(m[43]&m[610]&m[866]));
    m[205] = (((~m[43]&~m[626]&~m[882])|(m[43]&m[626]&~m[882]))&BiasedRNG[45])|(((m[43]&~m[626]&~m[882])|(~m[43]&m[626]&m[882]))&~BiasedRNG[45])|((~m[43]&~m[626]&m[882])|(m[43]&~m[626]&m[882])|(m[43]&m[626]&m[882]));
    m[206] = (((~m[43]&~m[642]&~m[898])|(m[43]&m[642]&~m[898]))&BiasedRNG[46])|(((m[43]&~m[642]&~m[898])|(~m[43]&m[642]&m[898]))&~BiasedRNG[46])|((~m[43]&~m[642]&m[898])|(m[43]&~m[642]&m[898])|(m[43]&m[642]&m[898]));
    m[207] = (((~m[43]&~m[658]&~m[914])|(m[43]&m[658]&~m[914]))&BiasedRNG[47])|(((m[43]&~m[658]&~m[914])|(~m[43]&m[658]&m[914]))&~BiasedRNG[47])|((~m[43]&~m[658]&m[914])|(m[43]&~m[658]&m[914])|(m[43]&m[658]&m[914]));
    m[208] = (((~m[44]&~m[419]&~m[675])|(m[44]&m[419]&~m[675]))&BiasedRNG[48])|(((m[44]&~m[419]&~m[675])|(~m[44]&m[419]&m[675]))&~BiasedRNG[48])|((~m[44]&~m[419]&m[675])|(m[44]&~m[419]&m[675])|(m[44]&m[419]&m[675]));
    m[209] = (((~m[44]&~m[435]&~m[691])|(m[44]&m[435]&~m[691]))&BiasedRNG[49])|(((m[44]&~m[435]&~m[691])|(~m[44]&m[435]&m[691]))&~BiasedRNG[49])|((~m[44]&~m[435]&m[691])|(m[44]&~m[435]&m[691])|(m[44]&m[435]&m[691]));
    m[210] = (((~m[44]&~m[451]&~m[707])|(m[44]&m[451]&~m[707]))&BiasedRNG[50])|(((m[44]&~m[451]&~m[707])|(~m[44]&m[451]&m[707]))&~BiasedRNG[50])|((~m[44]&~m[451]&m[707])|(m[44]&~m[451]&m[707])|(m[44]&m[451]&m[707]));
    m[211] = (((~m[44]&~m[467]&~m[723])|(m[44]&m[467]&~m[723]))&BiasedRNG[51])|(((m[44]&~m[467]&~m[723])|(~m[44]&m[467]&m[723]))&~BiasedRNG[51])|((~m[44]&~m[467]&m[723])|(m[44]&~m[467]&m[723])|(m[44]&m[467]&m[723]));
    m[212] = (((~m[45]&~m[483]&~m[739])|(m[45]&m[483]&~m[739]))&BiasedRNG[52])|(((m[45]&~m[483]&~m[739])|(~m[45]&m[483]&m[739]))&~BiasedRNG[52])|((~m[45]&~m[483]&m[739])|(m[45]&~m[483]&m[739])|(m[45]&m[483]&m[739]));
    m[213] = (((~m[45]&~m[499]&~m[755])|(m[45]&m[499]&~m[755]))&BiasedRNG[53])|(((m[45]&~m[499]&~m[755])|(~m[45]&m[499]&m[755]))&~BiasedRNG[53])|((~m[45]&~m[499]&m[755])|(m[45]&~m[499]&m[755])|(m[45]&m[499]&m[755]));
    m[214] = (((~m[45]&~m[515]&~m[771])|(m[45]&m[515]&~m[771]))&BiasedRNG[54])|(((m[45]&~m[515]&~m[771])|(~m[45]&m[515]&m[771]))&~BiasedRNG[54])|((~m[45]&~m[515]&m[771])|(m[45]&~m[515]&m[771])|(m[45]&m[515]&m[771]));
    m[215] = (((~m[45]&~m[531]&~m[787])|(m[45]&m[531]&~m[787]))&BiasedRNG[55])|(((m[45]&~m[531]&~m[787])|(~m[45]&m[531]&m[787]))&~BiasedRNG[55])|((~m[45]&~m[531]&m[787])|(m[45]&~m[531]&m[787])|(m[45]&m[531]&m[787]));
    m[216] = (((~m[46]&~m[547]&~m[803])|(m[46]&m[547]&~m[803]))&BiasedRNG[56])|(((m[46]&~m[547]&~m[803])|(~m[46]&m[547]&m[803]))&~BiasedRNG[56])|((~m[46]&~m[547]&m[803])|(m[46]&~m[547]&m[803])|(m[46]&m[547]&m[803]));
    m[217] = (((~m[46]&~m[563]&~m[819])|(m[46]&m[563]&~m[819]))&BiasedRNG[57])|(((m[46]&~m[563]&~m[819])|(~m[46]&m[563]&m[819]))&~BiasedRNG[57])|((~m[46]&~m[563]&m[819])|(m[46]&~m[563]&m[819])|(m[46]&m[563]&m[819]));
    m[218] = (((~m[46]&~m[579]&~m[835])|(m[46]&m[579]&~m[835]))&BiasedRNG[58])|(((m[46]&~m[579]&~m[835])|(~m[46]&m[579]&m[835]))&~BiasedRNG[58])|((~m[46]&~m[579]&m[835])|(m[46]&~m[579]&m[835])|(m[46]&m[579]&m[835]));
    m[219] = (((~m[46]&~m[595]&~m[851])|(m[46]&m[595]&~m[851]))&BiasedRNG[59])|(((m[46]&~m[595]&~m[851])|(~m[46]&m[595]&m[851]))&~BiasedRNG[59])|((~m[46]&~m[595]&m[851])|(m[46]&~m[595]&m[851])|(m[46]&m[595]&m[851]));
    m[220] = (((~m[47]&~m[611]&~m[867])|(m[47]&m[611]&~m[867]))&BiasedRNG[60])|(((m[47]&~m[611]&~m[867])|(~m[47]&m[611]&m[867]))&~BiasedRNG[60])|((~m[47]&~m[611]&m[867])|(m[47]&~m[611]&m[867])|(m[47]&m[611]&m[867]));
    m[221] = (((~m[47]&~m[627]&~m[883])|(m[47]&m[627]&~m[883]))&BiasedRNG[61])|(((m[47]&~m[627]&~m[883])|(~m[47]&m[627]&m[883]))&~BiasedRNG[61])|((~m[47]&~m[627]&m[883])|(m[47]&~m[627]&m[883])|(m[47]&m[627]&m[883]));
    m[222] = (((~m[47]&~m[643]&~m[899])|(m[47]&m[643]&~m[899]))&BiasedRNG[62])|(((m[47]&~m[643]&~m[899])|(~m[47]&m[643]&m[899]))&~BiasedRNG[62])|((~m[47]&~m[643]&m[899])|(m[47]&~m[643]&m[899])|(m[47]&m[643]&m[899]));
    m[223] = (((~m[47]&~m[659]&~m[915])|(m[47]&m[659]&~m[915]))&BiasedRNG[63])|(((m[47]&~m[659]&~m[915])|(~m[47]&m[659]&m[915]))&~BiasedRNG[63])|((~m[47]&~m[659]&m[915])|(m[47]&~m[659]&m[915])|(m[47]&m[659]&m[915]));
    m[224] = (((~m[48]&~m[420]&~m[676])|(m[48]&m[420]&~m[676]))&BiasedRNG[64])|(((m[48]&~m[420]&~m[676])|(~m[48]&m[420]&m[676]))&~BiasedRNG[64])|((~m[48]&~m[420]&m[676])|(m[48]&~m[420]&m[676])|(m[48]&m[420]&m[676]));
    m[225] = (((~m[48]&~m[436]&~m[692])|(m[48]&m[436]&~m[692]))&BiasedRNG[65])|(((m[48]&~m[436]&~m[692])|(~m[48]&m[436]&m[692]))&~BiasedRNG[65])|((~m[48]&~m[436]&m[692])|(m[48]&~m[436]&m[692])|(m[48]&m[436]&m[692]));
    m[226] = (((~m[48]&~m[452]&~m[708])|(m[48]&m[452]&~m[708]))&BiasedRNG[66])|(((m[48]&~m[452]&~m[708])|(~m[48]&m[452]&m[708]))&~BiasedRNG[66])|((~m[48]&~m[452]&m[708])|(m[48]&~m[452]&m[708])|(m[48]&m[452]&m[708]));
    m[227] = (((~m[48]&~m[468]&~m[724])|(m[48]&m[468]&~m[724]))&BiasedRNG[67])|(((m[48]&~m[468]&~m[724])|(~m[48]&m[468]&m[724]))&~BiasedRNG[67])|((~m[48]&~m[468]&m[724])|(m[48]&~m[468]&m[724])|(m[48]&m[468]&m[724]));
    m[228] = (((~m[49]&~m[484]&~m[740])|(m[49]&m[484]&~m[740]))&BiasedRNG[68])|(((m[49]&~m[484]&~m[740])|(~m[49]&m[484]&m[740]))&~BiasedRNG[68])|((~m[49]&~m[484]&m[740])|(m[49]&~m[484]&m[740])|(m[49]&m[484]&m[740]));
    m[229] = (((~m[49]&~m[500]&~m[756])|(m[49]&m[500]&~m[756]))&BiasedRNG[69])|(((m[49]&~m[500]&~m[756])|(~m[49]&m[500]&m[756]))&~BiasedRNG[69])|((~m[49]&~m[500]&m[756])|(m[49]&~m[500]&m[756])|(m[49]&m[500]&m[756]));
    m[230] = (((~m[49]&~m[516]&~m[772])|(m[49]&m[516]&~m[772]))&BiasedRNG[70])|(((m[49]&~m[516]&~m[772])|(~m[49]&m[516]&m[772]))&~BiasedRNG[70])|((~m[49]&~m[516]&m[772])|(m[49]&~m[516]&m[772])|(m[49]&m[516]&m[772]));
    m[231] = (((~m[49]&~m[532]&~m[788])|(m[49]&m[532]&~m[788]))&BiasedRNG[71])|(((m[49]&~m[532]&~m[788])|(~m[49]&m[532]&m[788]))&~BiasedRNG[71])|((~m[49]&~m[532]&m[788])|(m[49]&~m[532]&m[788])|(m[49]&m[532]&m[788]));
    m[232] = (((~m[50]&~m[548]&~m[804])|(m[50]&m[548]&~m[804]))&BiasedRNG[72])|(((m[50]&~m[548]&~m[804])|(~m[50]&m[548]&m[804]))&~BiasedRNG[72])|((~m[50]&~m[548]&m[804])|(m[50]&~m[548]&m[804])|(m[50]&m[548]&m[804]));
    m[233] = (((~m[50]&~m[564]&~m[820])|(m[50]&m[564]&~m[820]))&BiasedRNG[73])|(((m[50]&~m[564]&~m[820])|(~m[50]&m[564]&m[820]))&~BiasedRNG[73])|((~m[50]&~m[564]&m[820])|(m[50]&~m[564]&m[820])|(m[50]&m[564]&m[820]));
    m[234] = (((~m[50]&~m[580]&~m[836])|(m[50]&m[580]&~m[836]))&BiasedRNG[74])|(((m[50]&~m[580]&~m[836])|(~m[50]&m[580]&m[836]))&~BiasedRNG[74])|((~m[50]&~m[580]&m[836])|(m[50]&~m[580]&m[836])|(m[50]&m[580]&m[836]));
    m[235] = (((~m[50]&~m[596]&~m[852])|(m[50]&m[596]&~m[852]))&BiasedRNG[75])|(((m[50]&~m[596]&~m[852])|(~m[50]&m[596]&m[852]))&~BiasedRNG[75])|((~m[50]&~m[596]&m[852])|(m[50]&~m[596]&m[852])|(m[50]&m[596]&m[852]));
    m[236] = (((~m[51]&~m[612]&~m[868])|(m[51]&m[612]&~m[868]))&BiasedRNG[76])|(((m[51]&~m[612]&~m[868])|(~m[51]&m[612]&m[868]))&~BiasedRNG[76])|((~m[51]&~m[612]&m[868])|(m[51]&~m[612]&m[868])|(m[51]&m[612]&m[868]));
    m[237] = (((~m[51]&~m[628]&~m[884])|(m[51]&m[628]&~m[884]))&BiasedRNG[77])|(((m[51]&~m[628]&~m[884])|(~m[51]&m[628]&m[884]))&~BiasedRNG[77])|((~m[51]&~m[628]&m[884])|(m[51]&~m[628]&m[884])|(m[51]&m[628]&m[884]));
    m[238] = (((~m[51]&~m[644]&~m[900])|(m[51]&m[644]&~m[900]))&BiasedRNG[78])|(((m[51]&~m[644]&~m[900])|(~m[51]&m[644]&m[900]))&~BiasedRNG[78])|((~m[51]&~m[644]&m[900])|(m[51]&~m[644]&m[900])|(m[51]&m[644]&m[900]));
    m[239] = (((~m[51]&~m[660]&~m[916])|(m[51]&m[660]&~m[916]))&BiasedRNG[79])|(((m[51]&~m[660]&~m[916])|(~m[51]&m[660]&m[916]))&~BiasedRNG[79])|((~m[51]&~m[660]&m[916])|(m[51]&~m[660]&m[916])|(m[51]&m[660]&m[916]));
    m[240] = (((~m[52]&~m[421]&~m[677])|(m[52]&m[421]&~m[677]))&BiasedRNG[80])|(((m[52]&~m[421]&~m[677])|(~m[52]&m[421]&m[677]))&~BiasedRNG[80])|((~m[52]&~m[421]&m[677])|(m[52]&~m[421]&m[677])|(m[52]&m[421]&m[677]));
    m[241] = (((~m[52]&~m[437]&~m[693])|(m[52]&m[437]&~m[693]))&BiasedRNG[81])|(((m[52]&~m[437]&~m[693])|(~m[52]&m[437]&m[693]))&~BiasedRNG[81])|((~m[52]&~m[437]&m[693])|(m[52]&~m[437]&m[693])|(m[52]&m[437]&m[693]));
    m[242] = (((~m[52]&~m[453]&~m[709])|(m[52]&m[453]&~m[709]))&BiasedRNG[82])|(((m[52]&~m[453]&~m[709])|(~m[52]&m[453]&m[709]))&~BiasedRNG[82])|((~m[52]&~m[453]&m[709])|(m[52]&~m[453]&m[709])|(m[52]&m[453]&m[709]));
    m[243] = (((~m[52]&~m[469]&~m[725])|(m[52]&m[469]&~m[725]))&BiasedRNG[83])|(((m[52]&~m[469]&~m[725])|(~m[52]&m[469]&m[725]))&~BiasedRNG[83])|((~m[52]&~m[469]&m[725])|(m[52]&~m[469]&m[725])|(m[52]&m[469]&m[725]));
    m[244] = (((~m[53]&~m[485]&~m[741])|(m[53]&m[485]&~m[741]))&BiasedRNG[84])|(((m[53]&~m[485]&~m[741])|(~m[53]&m[485]&m[741]))&~BiasedRNG[84])|((~m[53]&~m[485]&m[741])|(m[53]&~m[485]&m[741])|(m[53]&m[485]&m[741]));
    m[245] = (((~m[53]&~m[501]&~m[757])|(m[53]&m[501]&~m[757]))&BiasedRNG[85])|(((m[53]&~m[501]&~m[757])|(~m[53]&m[501]&m[757]))&~BiasedRNG[85])|((~m[53]&~m[501]&m[757])|(m[53]&~m[501]&m[757])|(m[53]&m[501]&m[757]));
    m[246] = (((~m[53]&~m[517]&~m[773])|(m[53]&m[517]&~m[773]))&BiasedRNG[86])|(((m[53]&~m[517]&~m[773])|(~m[53]&m[517]&m[773]))&~BiasedRNG[86])|((~m[53]&~m[517]&m[773])|(m[53]&~m[517]&m[773])|(m[53]&m[517]&m[773]));
    m[247] = (((~m[53]&~m[533]&~m[789])|(m[53]&m[533]&~m[789]))&BiasedRNG[87])|(((m[53]&~m[533]&~m[789])|(~m[53]&m[533]&m[789]))&~BiasedRNG[87])|((~m[53]&~m[533]&m[789])|(m[53]&~m[533]&m[789])|(m[53]&m[533]&m[789]));
    m[248] = (((~m[54]&~m[549]&~m[805])|(m[54]&m[549]&~m[805]))&BiasedRNG[88])|(((m[54]&~m[549]&~m[805])|(~m[54]&m[549]&m[805]))&~BiasedRNG[88])|((~m[54]&~m[549]&m[805])|(m[54]&~m[549]&m[805])|(m[54]&m[549]&m[805]));
    m[249] = (((~m[54]&~m[565]&~m[821])|(m[54]&m[565]&~m[821]))&BiasedRNG[89])|(((m[54]&~m[565]&~m[821])|(~m[54]&m[565]&m[821]))&~BiasedRNG[89])|((~m[54]&~m[565]&m[821])|(m[54]&~m[565]&m[821])|(m[54]&m[565]&m[821]));
    m[250] = (((~m[54]&~m[581]&~m[837])|(m[54]&m[581]&~m[837]))&BiasedRNG[90])|(((m[54]&~m[581]&~m[837])|(~m[54]&m[581]&m[837]))&~BiasedRNG[90])|((~m[54]&~m[581]&m[837])|(m[54]&~m[581]&m[837])|(m[54]&m[581]&m[837]));
    m[251] = (((~m[54]&~m[597]&~m[853])|(m[54]&m[597]&~m[853]))&BiasedRNG[91])|(((m[54]&~m[597]&~m[853])|(~m[54]&m[597]&m[853]))&~BiasedRNG[91])|((~m[54]&~m[597]&m[853])|(m[54]&~m[597]&m[853])|(m[54]&m[597]&m[853]));
    m[252] = (((~m[55]&~m[613]&~m[869])|(m[55]&m[613]&~m[869]))&BiasedRNG[92])|(((m[55]&~m[613]&~m[869])|(~m[55]&m[613]&m[869]))&~BiasedRNG[92])|((~m[55]&~m[613]&m[869])|(m[55]&~m[613]&m[869])|(m[55]&m[613]&m[869]));
    m[253] = (((~m[55]&~m[629]&~m[885])|(m[55]&m[629]&~m[885]))&BiasedRNG[93])|(((m[55]&~m[629]&~m[885])|(~m[55]&m[629]&m[885]))&~BiasedRNG[93])|((~m[55]&~m[629]&m[885])|(m[55]&~m[629]&m[885])|(m[55]&m[629]&m[885]));
    m[254] = (((~m[55]&~m[645]&~m[901])|(m[55]&m[645]&~m[901]))&BiasedRNG[94])|(((m[55]&~m[645]&~m[901])|(~m[55]&m[645]&m[901]))&~BiasedRNG[94])|((~m[55]&~m[645]&m[901])|(m[55]&~m[645]&m[901])|(m[55]&m[645]&m[901]));
    m[255] = (((~m[55]&~m[661]&~m[917])|(m[55]&m[661]&~m[917]))&BiasedRNG[95])|(((m[55]&~m[661]&~m[917])|(~m[55]&m[661]&m[917]))&~BiasedRNG[95])|((~m[55]&~m[661]&m[917])|(m[55]&~m[661]&m[917])|(m[55]&m[661]&m[917]));
    m[256] = (((~m[56]&~m[422]&~m[678])|(m[56]&m[422]&~m[678]))&BiasedRNG[96])|(((m[56]&~m[422]&~m[678])|(~m[56]&m[422]&m[678]))&~BiasedRNG[96])|((~m[56]&~m[422]&m[678])|(m[56]&~m[422]&m[678])|(m[56]&m[422]&m[678]));
    m[257] = (((~m[56]&~m[438]&~m[694])|(m[56]&m[438]&~m[694]))&BiasedRNG[97])|(((m[56]&~m[438]&~m[694])|(~m[56]&m[438]&m[694]))&~BiasedRNG[97])|((~m[56]&~m[438]&m[694])|(m[56]&~m[438]&m[694])|(m[56]&m[438]&m[694]));
    m[258] = (((~m[56]&~m[454]&~m[710])|(m[56]&m[454]&~m[710]))&BiasedRNG[98])|(((m[56]&~m[454]&~m[710])|(~m[56]&m[454]&m[710]))&~BiasedRNG[98])|((~m[56]&~m[454]&m[710])|(m[56]&~m[454]&m[710])|(m[56]&m[454]&m[710]));
    m[259] = (((~m[56]&~m[470]&~m[726])|(m[56]&m[470]&~m[726]))&BiasedRNG[99])|(((m[56]&~m[470]&~m[726])|(~m[56]&m[470]&m[726]))&~BiasedRNG[99])|((~m[56]&~m[470]&m[726])|(m[56]&~m[470]&m[726])|(m[56]&m[470]&m[726]));
    m[260] = (((~m[57]&~m[486]&~m[742])|(m[57]&m[486]&~m[742]))&BiasedRNG[100])|(((m[57]&~m[486]&~m[742])|(~m[57]&m[486]&m[742]))&~BiasedRNG[100])|((~m[57]&~m[486]&m[742])|(m[57]&~m[486]&m[742])|(m[57]&m[486]&m[742]));
    m[261] = (((~m[57]&~m[502]&~m[758])|(m[57]&m[502]&~m[758]))&BiasedRNG[101])|(((m[57]&~m[502]&~m[758])|(~m[57]&m[502]&m[758]))&~BiasedRNG[101])|((~m[57]&~m[502]&m[758])|(m[57]&~m[502]&m[758])|(m[57]&m[502]&m[758]));
    m[262] = (((~m[57]&~m[518]&~m[774])|(m[57]&m[518]&~m[774]))&BiasedRNG[102])|(((m[57]&~m[518]&~m[774])|(~m[57]&m[518]&m[774]))&~BiasedRNG[102])|((~m[57]&~m[518]&m[774])|(m[57]&~m[518]&m[774])|(m[57]&m[518]&m[774]));
    m[263] = (((~m[57]&~m[534]&~m[790])|(m[57]&m[534]&~m[790]))&BiasedRNG[103])|(((m[57]&~m[534]&~m[790])|(~m[57]&m[534]&m[790]))&~BiasedRNG[103])|((~m[57]&~m[534]&m[790])|(m[57]&~m[534]&m[790])|(m[57]&m[534]&m[790]));
    m[264] = (((~m[58]&~m[550]&~m[806])|(m[58]&m[550]&~m[806]))&BiasedRNG[104])|(((m[58]&~m[550]&~m[806])|(~m[58]&m[550]&m[806]))&~BiasedRNG[104])|((~m[58]&~m[550]&m[806])|(m[58]&~m[550]&m[806])|(m[58]&m[550]&m[806]));
    m[265] = (((~m[58]&~m[566]&~m[822])|(m[58]&m[566]&~m[822]))&BiasedRNG[105])|(((m[58]&~m[566]&~m[822])|(~m[58]&m[566]&m[822]))&~BiasedRNG[105])|((~m[58]&~m[566]&m[822])|(m[58]&~m[566]&m[822])|(m[58]&m[566]&m[822]));
    m[266] = (((~m[58]&~m[582]&~m[838])|(m[58]&m[582]&~m[838]))&BiasedRNG[106])|(((m[58]&~m[582]&~m[838])|(~m[58]&m[582]&m[838]))&~BiasedRNG[106])|((~m[58]&~m[582]&m[838])|(m[58]&~m[582]&m[838])|(m[58]&m[582]&m[838]));
    m[267] = (((~m[58]&~m[598]&~m[854])|(m[58]&m[598]&~m[854]))&BiasedRNG[107])|(((m[58]&~m[598]&~m[854])|(~m[58]&m[598]&m[854]))&~BiasedRNG[107])|((~m[58]&~m[598]&m[854])|(m[58]&~m[598]&m[854])|(m[58]&m[598]&m[854]));
    m[268] = (((~m[59]&~m[614]&~m[870])|(m[59]&m[614]&~m[870]))&BiasedRNG[108])|(((m[59]&~m[614]&~m[870])|(~m[59]&m[614]&m[870]))&~BiasedRNG[108])|((~m[59]&~m[614]&m[870])|(m[59]&~m[614]&m[870])|(m[59]&m[614]&m[870]));
    m[269] = (((~m[59]&~m[630]&~m[886])|(m[59]&m[630]&~m[886]))&BiasedRNG[109])|(((m[59]&~m[630]&~m[886])|(~m[59]&m[630]&m[886]))&~BiasedRNG[109])|((~m[59]&~m[630]&m[886])|(m[59]&~m[630]&m[886])|(m[59]&m[630]&m[886]));
    m[270] = (((~m[59]&~m[646]&~m[902])|(m[59]&m[646]&~m[902]))&BiasedRNG[110])|(((m[59]&~m[646]&~m[902])|(~m[59]&m[646]&m[902]))&~BiasedRNG[110])|((~m[59]&~m[646]&m[902])|(m[59]&~m[646]&m[902])|(m[59]&m[646]&m[902]));
    m[271] = (((~m[59]&~m[662]&~m[918])|(m[59]&m[662]&~m[918]))&BiasedRNG[111])|(((m[59]&~m[662]&~m[918])|(~m[59]&m[662]&m[918]))&~BiasedRNG[111])|((~m[59]&~m[662]&m[918])|(m[59]&~m[662]&m[918])|(m[59]&m[662]&m[918]));
    m[272] = (((~m[60]&~m[423]&~m[679])|(m[60]&m[423]&~m[679]))&BiasedRNG[112])|(((m[60]&~m[423]&~m[679])|(~m[60]&m[423]&m[679]))&~BiasedRNG[112])|((~m[60]&~m[423]&m[679])|(m[60]&~m[423]&m[679])|(m[60]&m[423]&m[679]));
    m[273] = (((~m[60]&~m[439]&~m[695])|(m[60]&m[439]&~m[695]))&BiasedRNG[113])|(((m[60]&~m[439]&~m[695])|(~m[60]&m[439]&m[695]))&~BiasedRNG[113])|((~m[60]&~m[439]&m[695])|(m[60]&~m[439]&m[695])|(m[60]&m[439]&m[695]));
    m[274] = (((~m[60]&~m[455]&~m[711])|(m[60]&m[455]&~m[711]))&BiasedRNG[114])|(((m[60]&~m[455]&~m[711])|(~m[60]&m[455]&m[711]))&~BiasedRNG[114])|((~m[60]&~m[455]&m[711])|(m[60]&~m[455]&m[711])|(m[60]&m[455]&m[711]));
    m[275] = (((~m[60]&~m[471]&~m[727])|(m[60]&m[471]&~m[727]))&BiasedRNG[115])|(((m[60]&~m[471]&~m[727])|(~m[60]&m[471]&m[727]))&~BiasedRNG[115])|((~m[60]&~m[471]&m[727])|(m[60]&~m[471]&m[727])|(m[60]&m[471]&m[727]));
    m[276] = (((~m[61]&~m[487]&~m[743])|(m[61]&m[487]&~m[743]))&BiasedRNG[116])|(((m[61]&~m[487]&~m[743])|(~m[61]&m[487]&m[743]))&~BiasedRNG[116])|((~m[61]&~m[487]&m[743])|(m[61]&~m[487]&m[743])|(m[61]&m[487]&m[743]));
    m[277] = (((~m[61]&~m[503]&~m[759])|(m[61]&m[503]&~m[759]))&BiasedRNG[117])|(((m[61]&~m[503]&~m[759])|(~m[61]&m[503]&m[759]))&~BiasedRNG[117])|((~m[61]&~m[503]&m[759])|(m[61]&~m[503]&m[759])|(m[61]&m[503]&m[759]));
    m[278] = (((~m[61]&~m[519]&~m[775])|(m[61]&m[519]&~m[775]))&BiasedRNG[118])|(((m[61]&~m[519]&~m[775])|(~m[61]&m[519]&m[775]))&~BiasedRNG[118])|((~m[61]&~m[519]&m[775])|(m[61]&~m[519]&m[775])|(m[61]&m[519]&m[775]));
    m[279] = (((~m[61]&~m[535]&~m[791])|(m[61]&m[535]&~m[791]))&BiasedRNG[119])|(((m[61]&~m[535]&~m[791])|(~m[61]&m[535]&m[791]))&~BiasedRNG[119])|((~m[61]&~m[535]&m[791])|(m[61]&~m[535]&m[791])|(m[61]&m[535]&m[791]));
    m[280] = (((~m[62]&~m[551]&~m[807])|(m[62]&m[551]&~m[807]))&BiasedRNG[120])|(((m[62]&~m[551]&~m[807])|(~m[62]&m[551]&m[807]))&~BiasedRNG[120])|((~m[62]&~m[551]&m[807])|(m[62]&~m[551]&m[807])|(m[62]&m[551]&m[807]));
    m[281] = (((~m[62]&~m[567]&~m[823])|(m[62]&m[567]&~m[823]))&BiasedRNG[121])|(((m[62]&~m[567]&~m[823])|(~m[62]&m[567]&m[823]))&~BiasedRNG[121])|((~m[62]&~m[567]&m[823])|(m[62]&~m[567]&m[823])|(m[62]&m[567]&m[823]));
    m[282] = (((~m[62]&~m[583]&~m[839])|(m[62]&m[583]&~m[839]))&BiasedRNG[122])|(((m[62]&~m[583]&~m[839])|(~m[62]&m[583]&m[839]))&~BiasedRNG[122])|((~m[62]&~m[583]&m[839])|(m[62]&~m[583]&m[839])|(m[62]&m[583]&m[839]));
    m[283] = (((~m[62]&~m[599]&~m[855])|(m[62]&m[599]&~m[855]))&BiasedRNG[123])|(((m[62]&~m[599]&~m[855])|(~m[62]&m[599]&m[855]))&~BiasedRNG[123])|((~m[62]&~m[599]&m[855])|(m[62]&~m[599]&m[855])|(m[62]&m[599]&m[855]));
    m[284] = (((~m[63]&~m[615]&~m[871])|(m[63]&m[615]&~m[871]))&BiasedRNG[124])|(((m[63]&~m[615]&~m[871])|(~m[63]&m[615]&m[871]))&~BiasedRNG[124])|((~m[63]&~m[615]&m[871])|(m[63]&~m[615]&m[871])|(m[63]&m[615]&m[871]));
    m[285] = (((~m[63]&~m[631]&~m[887])|(m[63]&m[631]&~m[887]))&BiasedRNG[125])|(((m[63]&~m[631]&~m[887])|(~m[63]&m[631]&m[887]))&~BiasedRNG[125])|((~m[63]&~m[631]&m[887])|(m[63]&~m[631]&m[887])|(m[63]&m[631]&m[887]));
    m[286] = (((~m[63]&~m[647]&~m[903])|(m[63]&m[647]&~m[903]))&BiasedRNG[126])|(((m[63]&~m[647]&~m[903])|(~m[63]&m[647]&m[903]))&~BiasedRNG[126])|((~m[63]&~m[647]&m[903])|(m[63]&~m[647]&m[903])|(m[63]&m[647]&m[903]));
    m[287] = (((~m[63]&~m[663]&~m[919])|(m[63]&m[663]&~m[919]))&BiasedRNG[127])|(((m[63]&~m[663]&~m[919])|(~m[63]&m[663]&m[919]))&~BiasedRNG[127])|((~m[63]&~m[663]&m[919])|(m[63]&~m[663]&m[919])|(m[63]&m[663]&m[919]));
    m[288] = (((~m[64]&~m[424]&~m[680])|(m[64]&m[424]&~m[680]))&BiasedRNG[128])|(((m[64]&~m[424]&~m[680])|(~m[64]&m[424]&m[680]))&~BiasedRNG[128])|((~m[64]&~m[424]&m[680])|(m[64]&~m[424]&m[680])|(m[64]&m[424]&m[680]));
    m[289] = (((~m[64]&~m[440]&~m[696])|(m[64]&m[440]&~m[696]))&BiasedRNG[129])|(((m[64]&~m[440]&~m[696])|(~m[64]&m[440]&m[696]))&~BiasedRNG[129])|((~m[64]&~m[440]&m[696])|(m[64]&~m[440]&m[696])|(m[64]&m[440]&m[696]));
    m[290] = (((~m[64]&~m[456]&~m[712])|(m[64]&m[456]&~m[712]))&BiasedRNG[130])|(((m[64]&~m[456]&~m[712])|(~m[64]&m[456]&m[712]))&~BiasedRNG[130])|((~m[64]&~m[456]&m[712])|(m[64]&~m[456]&m[712])|(m[64]&m[456]&m[712]));
    m[291] = (((~m[64]&~m[472]&~m[728])|(m[64]&m[472]&~m[728]))&BiasedRNG[131])|(((m[64]&~m[472]&~m[728])|(~m[64]&m[472]&m[728]))&~BiasedRNG[131])|((~m[64]&~m[472]&m[728])|(m[64]&~m[472]&m[728])|(m[64]&m[472]&m[728]));
    m[292] = (((~m[65]&~m[488]&~m[744])|(m[65]&m[488]&~m[744]))&BiasedRNG[132])|(((m[65]&~m[488]&~m[744])|(~m[65]&m[488]&m[744]))&~BiasedRNG[132])|((~m[65]&~m[488]&m[744])|(m[65]&~m[488]&m[744])|(m[65]&m[488]&m[744]));
    m[293] = (((~m[65]&~m[504]&~m[760])|(m[65]&m[504]&~m[760]))&BiasedRNG[133])|(((m[65]&~m[504]&~m[760])|(~m[65]&m[504]&m[760]))&~BiasedRNG[133])|((~m[65]&~m[504]&m[760])|(m[65]&~m[504]&m[760])|(m[65]&m[504]&m[760]));
    m[294] = (((~m[65]&~m[520]&~m[776])|(m[65]&m[520]&~m[776]))&BiasedRNG[134])|(((m[65]&~m[520]&~m[776])|(~m[65]&m[520]&m[776]))&~BiasedRNG[134])|((~m[65]&~m[520]&m[776])|(m[65]&~m[520]&m[776])|(m[65]&m[520]&m[776]));
    m[295] = (((~m[65]&~m[536]&~m[792])|(m[65]&m[536]&~m[792]))&BiasedRNG[135])|(((m[65]&~m[536]&~m[792])|(~m[65]&m[536]&m[792]))&~BiasedRNG[135])|((~m[65]&~m[536]&m[792])|(m[65]&~m[536]&m[792])|(m[65]&m[536]&m[792]));
    m[296] = (((~m[66]&~m[552]&~m[808])|(m[66]&m[552]&~m[808]))&BiasedRNG[136])|(((m[66]&~m[552]&~m[808])|(~m[66]&m[552]&m[808]))&~BiasedRNG[136])|((~m[66]&~m[552]&m[808])|(m[66]&~m[552]&m[808])|(m[66]&m[552]&m[808]));
    m[297] = (((~m[66]&~m[568]&~m[824])|(m[66]&m[568]&~m[824]))&BiasedRNG[137])|(((m[66]&~m[568]&~m[824])|(~m[66]&m[568]&m[824]))&~BiasedRNG[137])|((~m[66]&~m[568]&m[824])|(m[66]&~m[568]&m[824])|(m[66]&m[568]&m[824]));
    m[298] = (((~m[66]&~m[584]&~m[840])|(m[66]&m[584]&~m[840]))&BiasedRNG[138])|(((m[66]&~m[584]&~m[840])|(~m[66]&m[584]&m[840]))&~BiasedRNG[138])|((~m[66]&~m[584]&m[840])|(m[66]&~m[584]&m[840])|(m[66]&m[584]&m[840]));
    m[299] = (((~m[66]&~m[600]&~m[856])|(m[66]&m[600]&~m[856]))&BiasedRNG[139])|(((m[66]&~m[600]&~m[856])|(~m[66]&m[600]&m[856]))&~BiasedRNG[139])|((~m[66]&~m[600]&m[856])|(m[66]&~m[600]&m[856])|(m[66]&m[600]&m[856]));
    m[300] = (((~m[67]&~m[616]&~m[872])|(m[67]&m[616]&~m[872]))&BiasedRNG[140])|(((m[67]&~m[616]&~m[872])|(~m[67]&m[616]&m[872]))&~BiasedRNG[140])|((~m[67]&~m[616]&m[872])|(m[67]&~m[616]&m[872])|(m[67]&m[616]&m[872]));
    m[301] = (((~m[67]&~m[632]&~m[888])|(m[67]&m[632]&~m[888]))&BiasedRNG[141])|(((m[67]&~m[632]&~m[888])|(~m[67]&m[632]&m[888]))&~BiasedRNG[141])|((~m[67]&~m[632]&m[888])|(m[67]&~m[632]&m[888])|(m[67]&m[632]&m[888]));
    m[302] = (((~m[67]&~m[648]&~m[904])|(m[67]&m[648]&~m[904]))&BiasedRNG[142])|(((m[67]&~m[648]&~m[904])|(~m[67]&m[648]&m[904]))&~BiasedRNG[142])|((~m[67]&~m[648]&m[904])|(m[67]&~m[648]&m[904])|(m[67]&m[648]&m[904]));
    m[303] = (((~m[67]&~m[664]&~m[920])|(m[67]&m[664]&~m[920]))&BiasedRNG[143])|(((m[67]&~m[664]&~m[920])|(~m[67]&m[664]&m[920]))&~BiasedRNG[143])|((~m[67]&~m[664]&m[920])|(m[67]&~m[664]&m[920])|(m[67]&m[664]&m[920]));
    m[304] = (((~m[68]&~m[425]&~m[681])|(m[68]&m[425]&~m[681]))&BiasedRNG[144])|(((m[68]&~m[425]&~m[681])|(~m[68]&m[425]&m[681]))&~BiasedRNG[144])|((~m[68]&~m[425]&m[681])|(m[68]&~m[425]&m[681])|(m[68]&m[425]&m[681]));
    m[305] = (((~m[68]&~m[441]&~m[697])|(m[68]&m[441]&~m[697]))&BiasedRNG[145])|(((m[68]&~m[441]&~m[697])|(~m[68]&m[441]&m[697]))&~BiasedRNG[145])|((~m[68]&~m[441]&m[697])|(m[68]&~m[441]&m[697])|(m[68]&m[441]&m[697]));
    m[306] = (((~m[68]&~m[457]&~m[713])|(m[68]&m[457]&~m[713]))&BiasedRNG[146])|(((m[68]&~m[457]&~m[713])|(~m[68]&m[457]&m[713]))&~BiasedRNG[146])|((~m[68]&~m[457]&m[713])|(m[68]&~m[457]&m[713])|(m[68]&m[457]&m[713]));
    m[307] = (((~m[68]&~m[473]&~m[729])|(m[68]&m[473]&~m[729]))&BiasedRNG[147])|(((m[68]&~m[473]&~m[729])|(~m[68]&m[473]&m[729]))&~BiasedRNG[147])|((~m[68]&~m[473]&m[729])|(m[68]&~m[473]&m[729])|(m[68]&m[473]&m[729]));
    m[308] = (((~m[69]&~m[489]&~m[745])|(m[69]&m[489]&~m[745]))&BiasedRNG[148])|(((m[69]&~m[489]&~m[745])|(~m[69]&m[489]&m[745]))&~BiasedRNG[148])|((~m[69]&~m[489]&m[745])|(m[69]&~m[489]&m[745])|(m[69]&m[489]&m[745]));
    m[309] = (((~m[69]&~m[505]&~m[761])|(m[69]&m[505]&~m[761]))&BiasedRNG[149])|(((m[69]&~m[505]&~m[761])|(~m[69]&m[505]&m[761]))&~BiasedRNG[149])|((~m[69]&~m[505]&m[761])|(m[69]&~m[505]&m[761])|(m[69]&m[505]&m[761]));
    m[310] = (((~m[69]&~m[521]&~m[777])|(m[69]&m[521]&~m[777]))&BiasedRNG[150])|(((m[69]&~m[521]&~m[777])|(~m[69]&m[521]&m[777]))&~BiasedRNG[150])|((~m[69]&~m[521]&m[777])|(m[69]&~m[521]&m[777])|(m[69]&m[521]&m[777]));
    m[311] = (((~m[69]&~m[537]&~m[793])|(m[69]&m[537]&~m[793]))&BiasedRNG[151])|(((m[69]&~m[537]&~m[793])|(~m[69]&m[537]&m[793]))&~BiasedRNG[151])|((~m[69]&~m[537]&m[793])|(m[69]&~m[537]&m[793])|(m[69]&m[537]&m[793]));
    m[312] = (((~m[70]&~m[553]&~m[809])|(m[70]&m[553]&~m[809]))&BiasedRNG[152])|(((m[70]&~m[553]&~m[809])|(~m[70]&m[553]&m[809]))&~BiasedRNG[152])|((~m[70]&~m[553]&m[809])|(m[70]&~m[553]&m[809])|(m[70]&m[553]&m[809]));
    m[313] = (((~m[70]&~m[569]&~m[825])|(m[70]&m[569]&~m[825]))&BiasedRNG[153])|(((m[70]&~m[569]&~m[825])|(~m[70]&m[569]&m[825]))&~BiasedRNG[153])|((~m[70]&~m[569]&m[825])|(m[70]&~m[569]&m[825])|(m[70]&m[569]&m[825]));
    m[314] = (((~m[70]&~m[585]&~m[841])|(m[70]&m[585]&~m[841]))&BiasedRNG[154])|(((m[70]&~m[585]&~m[841])|(~m[70]&m[585]&m[841]))&~BiasedRNG[154])|((~m[70]&~m[585]&m[841])|(m[70]&~m[585]&m[841])|(m[70]&m[585]&m[841]));
    m[315] = (((~m[70]&~m[601]&~m[857])|(m[70]&m[601]&~m[857]))&BiasedRNG[155])|(((m[70]&~m[601]&~m[857])|(~m[70]&m[601]&m[857]))&~BiasedRNG[155])|((~m[70]&~m[601]&m[857])|(m[70]&~m[601]&m[857])|(m[70]&m[601]&m[857]));
    m[316] = (((~m[71]&~m[617]&~m[873])|(m[71]&m[617]&~m[873]))&BiasedRNG[156])|(((m[71]&~m[617]&~m[873])|(~m[71]&m[617]&m[873]))&~BiasedRNG[156])|((~m[71]&~m[617]&m[873])|(m[71]&~m[617]&m[873])|(m[71]&m[617]&m[873]));
    m[317] = (((~m[71]&~m[633]&~m[889])|(m[71]&m[633]&~m[889]))&BiasedRNG[157])|(((m[71]&~m[633]&~m[889])|(~m[71]&m[633]&m[889]))&~BiasedRNG[157])|((~m[71]&~m[633]&m[889])|(m[71]&~m[633]&m[889])|(m[71]&m[633]&m[889]));
    m[318] = (((~m[71]&~m[649]&~m[905])|(m[71]&m[649]&~m[905]))&BiasedRNG[158])|(((m[71]&~m[649]&~m[905])|(~m[71]&m[649]&m[905]))&~BiasedRNG[158])|((~m[71]&~m[649]&m[905])|(m[71]&~m[649]&m[905])|(m[71]&m[649]&m[905]));
    m[319] = (((~m[71]&~m[665]&~m[921])|(m[71]&m[665]&~m[921]))&BiasedRNG[159])|(((m[71]&~m[665]&~m[921])|(~m[71]&m[665]&m[921]))&~BiasedRNG[159])|((~m[71]&~m[665]&m[921])|(m[71]&~m[665]&m[921])|(m[71]&m[665]&m[921]));
    m[320] = (((~m[72]&~m[426]&~m[682])|(m[72]&m[426]&~m[682]))&BiasedRNG[160])|(((m[72]&~m[426]&~m[682])|(~m[72]&m[426]&m[682]))&~BiasedRNG[160])|((~m[72]&~m[426]&m[682])|(m[72]&~m[426]&m[682])|(m[72]&m[426]&m[682]));
    m[321] = (((~m[72]&~m[442]&~m[698])|(m[72]&m[442]&~m[698]))&BiasedRNG[161])|(((m[72]&~m[442]&~m[698])|(~m[72]&m[442]&m[698]))&~BiasedRNG[161])|((~m[72]&~m[442]&m[698])|(m[72]&~m[442]&m[698])|(m[72]&m[442]&m[698]));
    m[322] = (((~m[72]&~m[458]&~m[714])|(m[72]&m[458]&~m[714]))&BiasedRNG[162])|(((m[72]&~m[458]&~m[714])|(~m[72]&m[458]&m[714]))&~BiasedRNG[162])|((~m[72]&~m[458]&m[714])|(m[72]&~m[458]&m[714])|(m[72]&m[458]&m[714]));
    m[323] = (((~m[72]&~m[474]&~m[730])|(m[72]&m[474]&~m[730]))&BiasedRNG[163])|(((m[72]&~m[474]&~m[730])|(~m[72]&m[474]&m[730]))&~BiasedRNG[163])|((~m[72]&~m[474]&m[730])|(m[72]&~m[474]&m[730])|(m[72]&m[474]&m[730]));
    m[324] = (((~m[73]&~m[490]&~m[746])|(m[73]&m[490]&~m[746]))&BiasedRNG[164])|(((m[73]&~m[490]&~m[746])|(~m[73]&m[490]&m[746]))&~BiasedRNG[164])|((~m[73]&~m[490]&m[746])|(m[73]&~m[490]&m[746])|(m[73]&m[490]&m[746]));
    m[325] = (((~m[73]&~m[506]&~m[762])|(m[73]&m[506]&~m[762]))&BiasedRNG[165])|(((m[73]&~m[506]&~m[762])|(~m[73]&m[506]&m[762]))&~BiasedRNG[165])|((~m[73]&~m[506]&m[762])|(m[73]&~m[506]&m[762])|(m[73]&m[506]&m[762]));
    m[326] = (((~m[73]&~m[522]&~m[778])|(m[73]&m[522]&~m[778]))&BiasedRNG[166])|(((m[73]&~m[522]&~m[778])|(~m[73]&m[522]&m[778]))&~BiasedRNG[166])|((~m[73]&~m[522]&m[778])|(m[73]&~m[522]&m[778])|(m[73]&m[522]&m[778]));
    m[327] = (((~m[73]&~m[538]&~m[794])|(m[73]&m[538]&~m[794]))&BiasedRNG[167])|(((m[73]&~m[538]&~m[794])|(~m[73]&m[538]&m[794]))&~BiasedRNG[167])|((~m[73]&~m[538]&m[794])|(m[73]&~m[538]&m[794])|(m[73]&m[538]&m[794]));
    m[328] = (((~m[74]&~m[554]&~m[810])|(m[74]&m[554]&~m[810]))&BiasedRNG[168])|(((m[74]&~m[554]&~m[810])|(~m[74]&m[554]&m[810]))&~BiasedRNG[168])|((~m[74]&~m[554]&m[810])|(m[74]&~m[554]&m[810])|(m[74]&m[554]&m[810]));
    m[329] = (((~m[74]&~m[570]&~m[826])|(m[74]&m[570]&~m[826]))&BiasedRNG[169])|(((m[74]&~m[570]&~m[826])|(~m[74]&m[570]&m[826]))&~BiasedRNG[169])|((~m[74]&~m[570]&m[826])|(m[74]&~m[570]&m[826])|(m[74]&m[570]&m[826]));
    m[330] = (((~m[74]&~m[586]&~m[842])|(m[74]&m[586]&~m[842]))&BiasedRNG[170])|(((m[74]&~m[586]&~m[842])|(~m[74]&m[586]&m[842]))&~BiasedRNG[170])|((~m[74]&~m[586]&m[842])|(m[74]&~m[586]&m[842])|(m[74]&m[586]&m[842]));
    m[331] = (((~m[74]&~m[602]&~m[858])|(m[74]&m[602]&~m[858]))&BiasedRNG[171])|(((m[74]&~m[602]&~m[858])|(~m[74]&m[602]&m[858]))&~BiasedRNG[171])|((~m[74]&~m[602]&m[858])|(m[74]&~m[602]&m[858])|(m[74]&m[602]&m[858]));
    m[332] = (((~m[75]&~m[618]&~m[874])|(m[75]&m[618]&~m[874]))&BiasedRNG[172])|(((m[75]&~m[618]&~m[874])|(~m[75]&m[618]&m[874]))&~BiasedRNG[172])|((~m[75]&~m[618]&m[874])|(m[75]&~m[618]&m[874])|(m[75]&m[618]&m[874]));
    m[333] = (((~m[75]&~m[634]&~m[890])|(m[75]&m[634]&~m[890]))&BiasedRNG[173])|(((m[75]&~m[634]&~m[890])|(~m[75]&m[634]&m[890]))&~BiasedRNG[173])|((~m[75]&~m[634]&m[890])|(m[75]&~m[634]&m[890])|(m[75]&m[634]&m[890]));
    m[334] = (((~m[75]&~m[650]&~m[906])|(m[75]&m[650]&~m[906]))&BiasedRNG[174])|(((m[75]&~m[650]&~m[906])|(~m[75]&m[650]&m[906]))&~BiasedRNG[174])|((~m[75]&~m[650]&m[906])|(m[75]&~m[650]&m[906])|(m[75]&m[650]&m[906]));
    m[335] = (((~m[75]&~m[666]&~m[922])|(m[75]&m[666]&~m[922]))&BiasedRNG[175])|(((m[75]&~m[666]&~m[922])|(~m[75]&m[666]&m[922]))&~BiasedRNG[175])|((~m[75]&~m[666]&m[922])|(m[75]&~m[666]&m[922])|(m[75]&m[666]&m[922]));
    m[336] = (((~m[76]&~m[427]&~m[683])|(m[76]&m[427]&~m[683]))&BiasedRNG[176])|(((m[76]&~m[427]&~m[683])|(~m[76]&m[427]&m[683]))&~BiasedRNG[176])|((~m[76]&~m[427]&m[683])|(m[76]&~m[427]&m[683])|(m[76]&m[427]&m[683]));
    m[337] = (((~m[76]&~m[443]&~m[699])|(m[76]&m[443]&~m[699]))&BiasedRNG[177])|(((m[76]&~m[443]&~m[699])|(~m[76]&m[443]&m[699]))&~BiasedRNG[177])|((~m[76]&~m[443]&m[699])|(m[76]&~m[443]&m[699])|(m[76]&m[443]&m[699]));
    m[338] = (((~m[76]&~m[459]&~m[715])|(m[76]&m[459]&~m[715]))&BiasedRNG[178])|(((m[76]&~m[459]&~m[715])|(~m[76]&m[459]&m[715]))&~BiasedRNG[178])|((~m[76]&~m[459]&m[715])|(m[76]&~m[459]&m[715])|(m[76]&m[459]&m[715]));
    m[339] = (((~m[76]&~m[475]&~m[731])|(m[76]&m[475]&~m[731]))&BiasedRNG[179])|(((m[76]&~m[475]&~m[731])|(~m[76]&m[475]&m[731]))&~BiasedRNG[179])|((~m[76]&~m[475]&m[731])|(m[76]&~m[475]&m[731])|(m[76]&m[475]&m[731]));
    m[340] = (((~m[77]&~m[491]&~m[747])|(m[77]&m[491]&~m[747]))&BiasedRNG[180])|(((m[77]&~m[491]&~m[747])|(~m[77]&m[491]&m[747]))&~BiasedRNG[180])|((~m[77]&~m[491]&m[747])|(m[77]&~m[491]&m[747])|(m[77]&m[491]&m[747]));
    m[341] = (((~m[77]&~m[507]&~m[763])|(m[77]&m[507]&~m[763]))&BiasedRNG[181])|(((m[77]&~m[507]&~m[763])|(~m[77]&m[507]&m[763]))&~BiasedRNG[181])|((~m[77]&~m[507]&m[763])|(m[77]&~m[507]&m[763])|(m[77]&m[507]&m[763]));
    m[342] = (((~m[77]&~m[523]&~m[779])|(m[77]&m[523]&~m[779]))&BiasedRNG[182])|(((m[77]&~m[523]&~m[779])|(~m[77]&m[523]&m[779]))&~BiasedRNG[182])|((~m[77]&~m[523]&m[779])|(m[77]&~m[523]&m[779])|(m[77]&m[523]&m[779]));
    m[343] = (((~m[77]&~m[539]&~m[795])|(m[77]&m[539]&~m[795]))&BiasedRNG[183])|(((m[77]&~m[539]&~m[795])|(~m[77]&m[539]&m[795]))&~BiasedRNG[183])|((~m[77]&~m[539]&m[795])|(m[77]&~m[539]&m[795])|(m[77]&m[539]&m[795]));
    m[344] = (((~m[78]&~m[555]&~m[811])|(m[78]&m[555]&~m[811]))&BiasedRNG[184])|(((m[78]&~m[555]&~m[811])|(~m[78]&m[555]&m[811]))&~BiasedRNG[184])|((~m[78]&~m[555]&m[811])|(m[78]&~m[555]&m[811])|(m[78]&m[555]&m[811]));
    m[345] = (((~m[78]&~m[571]&~m[827])|(m[78]&m[571]&~m[827]))&BiasedRNG[185])|(((m[78]&~m[571]&~m[827])|(~m[78]&m[571]&m[827]))&~BiasedRNG[185])|((~m[78]&~m[571]&m[827])|(m[78]&~m[571]&m[827])|(m[78]&m[571]&m[827]));
    m[346] = (((~m[78]&~m[587]&~m[843])|(m[78]&m[587]&~m[843]))&BiasedRNG[186])|(((m[78]&~m[587]&~m[843])|(~m[78]&m[587]&m[843]))&~BiasedRNG[186])|((~m[78]&~m[587]&m[843])|(m[78]&~m[587]&m[843])|(m[78]&m[587]&m[843]));
    m[347] = (((~m[78]&~m[603]&~m[859])|(m[78]&m[603]&~m[859]))&BiasedRNG[187])|(((m[78]&~m[603]&~m[859])|(~m[78]&m[603]&m[859]))&~BiasedRNG[187])|((~m[78]&~m[603]&m[859])|(m[78]&~m[603]&m[859])|(m[78]&m[603]&m[859]));
    m[348] = (((~m[79]&~m[619]&~m[875])|(m[79]&m[619]&~m[875]))&BiasedRNG[188])|(((m[79]&~m[619]&~m[875])|(~m[79]&m[619]&m[875]))&~BiasedRNG[188])|((~m[79]&~m[619]&m[875])|(m[79]&~m[619]&m[875])|(m[79]&m[619]&m[875]));
    m[349] = (((~m[79]&~m[635]&~m[891])|(m[79]&m[635]&~m[891]))&BiasedRNG[189])|(((m[79]&~m[635]&~m[891])|(~m[79]&m[635]&m[891]))&~BiasedRNG[189])|((~m[79]&~m[635]&m[891])|(m[79]&~m[635]&m[891])|(m[79]&m[635]&m[891]));
    m[350] = (((~m[79]&~m[651]&~m[907])|(m[79]&m[651]&~m[907]))&BiasedRNG[190])|(((m[79]&~m[651]&~m[907])|(~m[79]&m[651]&m[907]))&~BiasedRNG[190])|((~m[79]&~m[651]&m[907])|(m[79]&~m[651]&m[907])|(m[79]&m[651]&m[907]));
    m[351] = (((~m[79]&~m[667]&~m[923])|(m[79]&m[667]&~m[923]))&BiasedRNG[191])|(((m[79]&~m[667]&~m[923])|(~m[79]&m[667]&m[923]))&~BiasedRNG[191])|((~m[79]&~m[667]&m[923])|(m[79]&~m[667]&m[923])|(m[79]&m[667]&m[923]));
    m[352] = (((~m[80]&~m[428]&~m[684])|(m[80]&m[428]&~m[684]))&BiasedRNG[192])|(((m[80]&~m[428]&~m[684])|(~m[80]&m[428]&m[684]))&~BiasedRNG[192])|((~m[80]&~m[428]&m[684])|(m[80]&~m[428]&m[684])|(m[80]&m[428]&m[684]));
    m[353] = (((~m[80]&~m[444]&~m[700])|(m[80]&m[444]&~m[700]))&BiasedRNG[193])|(((m[80]&~m[444]&~m[700])|(~m[80]&m[444]&m[700]))&~BiasedRNG[193])|((~m[80]&~m[444]&m[700])|(m[80]&~m[444]&m[700])|(m[80]&m[444]&m[700]));
    m[354] = (((~m[80]&~m[460]&~m[716])|(m[80]&m[460]&~m[716]))&BiasedRNG[194])|(((m[80]&~m[460]&~m[716])|(~m[80]&m[460]&m[716]))&~BiasedRNG[194])|((~m[80]&~m[460]&m[716])|(m[80]&~m[460]&m[716])|(m[80]&m[460]&m[716]));
    m[355] = (((~m[80]&~m[476]&~m[732])|(m[80]&m[476]&~m[732]))&BiasedRNG[195])|(((m[80]&~m[476]&~m[732])|(~m[80]&m[476]&m[732]))&~BiasedRNG[195])|((~m[80]&~m[476]&m[732])|(m[80]&~m[476]&m[732])|(m[80]&m[476]&m[732]));
    m[356] = (((~m[81]&~m[492]&~m[748])|(m[81]&m[492]&~m[748]))&BiasedRNG[196])|(((m[81]&~m[492]&~m[748])|(~m[81]&m[492]&m[748]))&~BiasedRNG[196])|((~m[81]&~m[492]&m[748])|(m[81]&~m[492]&m[748])|(m[81]&m[492]&m[748]));
    m[357] = (((~m[81]&~m[508]&~m[764])|(m[81]&m[508]&~m[764]))&BiasedRNG[197])|(((m[81]&~m[508]&~m[764])|(~m[81]&m[508]&m[764]))&~BiasedRNG[197])|((~m[81]&~m[508]&m[764])|(m[81]&~m[508]&m[764])|(m[81]&m[508]&m[764]));
    m[358] = (((~m[81]&~m[524]&~m[780])|(m[81]&m[524]&~m[780]))&BiasedRNG[198])|(((m[81]&~m[524]&~m[780])|(~m[81]&m[524]&m[780]))&~BiasedRNG[198])|((~m[81]&~m[524]&m[780])|(m[81]&~m[524]&m[780])|(m[81]&m[524]&m[780]));
    m[359] = (((~m[81]&~m[540]&~m[796])|(m[81]&m[540]&~m[796]))&BiasedRNG[199])|(((m[81]&~m[540]&~m[796])|(~m[81]&m[540]&m[796]))&~BiasedRNG[199])|((~m[81]&~m[540]&m[796])|(m[81]&~m[540]&m[796])|(m[81]&m[540]&m[796]));
    m[360] = (((~m[82]&~m[556]&~m[812])|(m[82]&m[556]&~m[812]))&BiasedRNG[200])|(((m[82]&~m[556]&~m[812])|(~m[82]&m[556]&m[812]))&~BiasedRNG[200])|((~m[82]&~m[556]&m[812])|(m[82]&~m[556]&m[812])|(m[82]&m[556]&m[812]));
    m[361] = (((~m[82]&~m[572]&~m[828])|(m[82]&m[572]&~m[828]))&BiasedRNG[201])|(((m[82]&~m[572]&~m[828])|(~m[82]&m[572]&m[828]))&~BiasedRNG[201])|((~m[82]&~m[572]&m[828])|(m[82]&~m[572]&m[828])|(m[82]&m[572]&m[828]));
    m[362] = (((~m[82]&~m[588]&~m[844])|(m[82]&m[588]&~m[844]))&BiasedRNG[202])|(((m[82]&~m[588]&~m[844])|(~m[82]&m[588]&m[844]))&~BiasedRNG[202])|((~m[82]&~m[588]&m[844])|(m[82]&~m[588]&m[844])|(m[82]&m[588]&m[844]));
    m[363] = (((~m[82]&~m[604]&~m[860])|(m[82]&m[604]&~m[860]))&BiasedRNG[203])|(((m[82]&~m[604]&~m[860])|(~m[82]&m[604]&m[860]))&~BiasedRNG[203])|((~m[82]&~m[604]&m[860])|(m[82]&~m[604]&m[860])|(m[82]&m[604]&m[860]));
    m[364] = (((~m[83]&~m[620]&~m[876])|(m[83]&m[620]&~m[876]))&BiasedRNG[204])|(((m[83]&~m[620]&~m[876])|(~m[83]&m[620]&m[876]))&~BiasedRNG[204])|((~m[83]&~m[620]&m[876])|(m[83]&~m[620]&m[876])|(m[83]&m[620]&m[876]));
    m[365] = (((~m[83]&~m[636]&~m[892])|(m[83]&m[636]&~m[892]))&BiasedRNG[205])|(((m[83]&~m[636]&~m[892])|(~m[83]&m[636]&m[892]))&~BiasedRNG[205])|((~m[83]&~m[636]&m[892])|(m[83]&~m[636]&m[892])|(m[83]&m[636]&m[892]));
    m[366] = (((~m[83]&~m[652]&~m[908])|(m[83]&m[652]&~m[908]))&BiasedRNG[206])|(((m[83]&~m[652]&~m[908])|(~m[83]&m[652]&m[908]))&~BiasedRNG[206])|((~m[83]&~m[652]&m[908])|(m[83]&~m[652]&m[908])|(m[83]&m[652]&m[908]));
    m[367] = (((~m[83]&~m[668]&~m[924])|(m[83]&m[668]&~m[924]))&BiasedRNG[207])|(((m[83]&~m[668]&~m[924])|(~m[83]&m[668]&m[924]))&~BiasedRNG[207])|((~m[83]&~m[668]&m[924])|(m[83]&~m[668]&m[924])|(m[83]&m[668]&m[924]));
    m[368] = (((~m[84]&~m[429]&~m[685])|(m[84]&m[429]&~m[685]))&BiasedRNG[208])|(((m[84]&~m[429]&~m[685])|(~m[84]&m[429]&m[685]))&~BiasedRNG[208])|((~m[84]&~m[429]&m[685])|(m[84]&~m[429]&m[685])|(m[84]&m[429]&m[685]));
    m[369] = (((~m[84]&~m[445]&~m[701])|(m[84]&m[445]&~m[701]))&BiasedRNG[209])|(((m[84]&~m[445]&~m[701])|(~m[84]&m[445]&m[701]))&~BiasedRNG[209])|((~m[84]&~m[445]&m[701])|(m[84]&~m[445]&m[701])|(m[84]&m[445]&m[701]));
    m[370] = (((~m[84]&~m[461]&~m[717])|(m[84]&m[461]&~m[717]))&BiasedRNG[210])|(((m[84]&~m[461]&~m[717])|(~m[84]&m[461]&m[717]))&~BiasedRNG[210])|((~m[84]&~m[461]&m[717])|(m[84]&~m[461]&m[717])|(m[84]&m[461]&m[717]));
    m[371] = (((~m[84]&~m[477]&~m[733])|(m[84]&m[477]&~m[733]))&BiasedRNG[211])|(((m[84]&~m[477]&~m[733])|(~m[84]&m[477]&m[733]))&~BiasedRNG[211])|((~m[84]&~m[477]&m[733])|(m[84]&~m[477]&m[733])|(m[84]&m[477]&m[733]));
    m[372] = (((~m[85]&~m[493]&~m[749])|(m[85]&m[493]&~m[749]))&BiasedRNG[212])|(((m[85]&~m[493]&~m[749])|(~m[85]&m[493]&m[749]))&~BiasedRNG[212])|((~m[85]&~m[493]&m[749])|(m[85]&~m[493]&m[749])|(m[85]&m[493]&m[749]));
    m[373] = (((~m[85]&~m[509]&~m[765])|(m[85]&m[509]&~m[765]))&BiasedRNG[213])|(((m[85]&~m[509]&~m[765])|(~m[85]&m[509]&m[765]))&~BiasedRNG[213])|((~m[85]&~m[509]&m[765])|(m[85]&~m[509]&m[765])|(m[85]&m[509]&m[765]));
    m[374] = (((~m[85]&~m[525]&~m[781])|(m[85]&m[525]&~m[781]))&BiasedRNG[214])|(((m[85]&~m[525]&~m[781])|(~m[85]&m[525]&m[781]))&~BiasedRNG[214])|((~m[85]&~m[525]&m[781])|(m[85]&~m[525]&m[781])|(m[85]&m[525]&m[781]));
    m[375] = (((~m[85]&~m[541]&~m[797])|(m[85]&m[541]&~m[797]))&BiasedRNG[215])|(((m[85]&~m[541]&~m[797])|(~m[85]&m[541]&m[797]))&~BiasedRNG[215])|((~m[85]&~m[541]&m[797])|(m[85]&~m[541]&m[797])|(m[85]&m[541]&m[797]));
    m[376] = (((~m[86]&~m[557]&~m[813])|(m[86]&m[557]&~m[813]))&BiasedRNG[216])|(((m[86]&~m[557]&~m[813])|(~m[86]&m[557]&m[813]))&~BiasedRNG[216])|((~m[86]&~m[557]&m[813])|(m[86]&~m[557]&m[813])|(m[86]&m[557]&m[813]));
    m[377] = (((~m[86]&~m[573]&~m[829])|(m[86]&m[573]&~m[829]))&BiasedRNG[217])|(((m[86]&~m[573]&~m[829])|(~m[86]&m[573]&m[829]))&~BiasedRNG[217])|((~m[86]&~m[573]&m[829])|(m[86]&~m[573]&m[829])|(m[86]&m[573]&m[829]));
    m[378] = (((~m[86]&~m[589]&~m[845])|(m[86]&m[589]&~m[845]))&BiasedRNG[218])|(((m[86]&~m[589]&~m[845])|(~m[86]&m[589]&m[845]))&~BiasedRNG[218])|((~m[86]&~m[589]&m[845])|(m[86]&~m[589]&m[845])|(m[86]&m[589]&m[845]));
    m[379] = (((~m[86]&~m[605]&~m[861])|(m[86]&m[605]&~m[861]))&BiasedRNG[219])|(((m[86]&~m[605]&~m[861])|(~m[86]&m[605]&m[861]))&~BiasedRNG[219])|((~m[86]&~m[605]&m[861])|(m[86]&~m[605]&m[861])|(m[86]&m[605]&m[861]));
    m[380] = (((~m[87]&~m[621]&~m[877])|(m[87]&m[621]&~m[877]))&BiasedRNG[220])|(((m[87]&~m[621]&~m[877])|(~m[87]&m[621]&m[877]))&~BiasedRNG[220])|((~m[87]&~m[621]&m[877])|(m[87]&~m[621]&m[877])|(m[87]&m[621]&m[877]));
    m[381] = (((~m[87]&~m[637]&~m[893])|(m[87]&m[637]&~m[893]))&BiasedRNG[221])|(((m[87]&~m[637]&~m[893])|(~m[87]&m[637]&m[893]))&~BiasedRNG[221])|((~m[87]&~m[637]&m[893])|(m[87]&~m[637]&m[893])|(m[87]&m[637]&m[893]));
    m[382] = (((~m[87]&~m[653]&~m[909])|(m[87]&m[653]&~m[909]))&BiasedRNG[222])|(((m[87]&~m[653]&~m[909])|(~m[87]&m[653]&m[909]))&~BiasedRNG[222])|((~m[87]&~m[653]&m[909])|(m[87]&~m[653]&m[909])|(m[87]&m[653]&m[909]));
    m[383] = (((~m[87]&~m[669]&~m[925])|(m[87]&m[669]&~m[925]))&BiasedRNG[223])|(((m[87]&~m[669]&~m[925])|(~m[87]&m[669]&m[925]))&~BiasedRNG[223])|((~m[87]&~m[669]&m[925])|(m[87]&~m[669]&m[925])|(m[87]&m[669]&m[925]));
    m[384] = (((~m[88]&~m[430]&~m[686])|(m[88]&m[430]&~m[686]))&BiasedRNG[224])|(((m[88]&~m[430]&~m[686])|(~m[88]&m[430]&m[686]))&~BiasedRNG[224])|((~m[88]&~m[430]&m[686])|(m[88]&~m[430]&m[686])|(m[88]&m[430]&m[686]));
    m[385] = (((~m[88]&~m[446]&~m[702])|(m[88]&m[446]&~m[702]))&BiasedRNG[225])|(((m[88]&~m[446]&~m[702])|(~m[88]&m[446]&m[702]))&~BiasedRNG[225])|((~m[88]&~m[446]&m[702])|(m[88]&~m[446]&m[702])|(m[88]&m[446]&m[702]));
    m[386] = (((~m[88]&~m[462]&~m[718])|(m[88]&m[462]&~m[718]))&BiasedRNG[226])|(((m[88]&~m[462]&~m[718])|(~m[88]&m[462]&m[718]))&~BiasedRNG[226])|((~m[88]&~m[462]&m[718])|(m[88]&~m[462]&m[718])|(m[88]&m[462]&m[718]));
    m[387] = (((~m[88]&~m[478]&~m[734])|(m[88]&m[478]&~m[734]))&BiasedRNG[227])|(((m[88]&~m[478]&~m[734])|(~m[88]&m[478]&m[734]))&~BiasedRNG[227])|((~m[88]&~m[478]&m[734])|(m[88]&~m[478]&m[734])|(m[88]&m[478]&m[734]));
    m[388] = (((~m[89]&~m[494]&~m[750])|(m[89]&m[494]&~m[750]))&BiasedRNG[228])|(((m[89]&~m[494]&~m[750])|(~m[89]&m[494]&m[750]))&~BiasedRNG[228])|((~m[89]&~m[494]&m[750])|(m[89]&~m[494]&m[750])|(m[89]&m[494]&m[750]));
    m[389] = (((~m[89]&~m[510]&~m[766])|(m[89]&m[510]&~m[766]))&BiasedRNG[229])|(((m[89]&~m[510]&~m[766])|(~m[89]&m[510]&m[766]))&~BiasedRNG[229])|((~m[89]&~m[510]&m[766])|(m[89]&~m[510]&m[766])|(m[89]&m[510]&m[766]));
    m[390] = (((~m[89]&~m[526]&~m[782])|(m[89]&m[526]&~m[782]))&BiasedRNG[230])|(((m[89]&~m[526]&~m[782])|(~m[89]&m[526]&m[782]))&~BiasedRNG[230])|((~m[89]&~m[526]&m[782])|(m[89]&~m[526]&m[782])|(m[89]&m[526]&m[782]));
    m[391] = (((~m[89]&~m[542]&~m[798])|(m[89]&m[542]&~m[798]))&BiasedRNG[231])|(((m[89]&~m[542]&~m[798])|(~m[89]&m[542]&m[798]))&~BiasedRNG[231])|((~m[89]&~m[542]&m[798])|(m[89]&~m[542]&m[798])|(m[89]&m[542]&m[798]));
    m[392] = (((~m[90]&~m[558]&~m[814])|(m[90]&m[558]&~m[814]))&BiasedRNG[232])|(((m[90]&~m[558]&~m[814])|(~m[90]&m[558]&m[814]))&~BiasedRNG[232])|((~m[90]&~m[558]&m[814])|(m[90]&~m[558]&m[814])|(m[90]&m[558]&m[814]));
    m[393] = (((~m[90]&~m[574]&~m[830])|(m[90]&m[574]&~m[830]))&BiasedRNG[233])|(((m[90]&~m[574]&~m[830])|(~m[90]&m[574]&m[830]))&~BiasedRNG[233])|((~m[90]&~m[574]&m[830])|(m[90]&~m[574]&m[830])|(m[90]&m[574]&m[830]));
    m[394] = (((~m[90]&~m[590]&~m[846])|(m[90]&m[590]&~m[846]))&BiasedRNG[234])|(((m[90]&~m[590]&~m[846])|(~m[90]&m[590]&m[846]))&~BiasedRNG[234])|((~m[90]&~m[590]&m[846])|(m[90]&~m[590]&m[846])|(m[90]&m[590]&m[846]));
    m[395] = (((~m[90]&~m[606]&~m[862])|(m[90]&m[606]&~m[862]))&BiasedRNG[235])|(((m[90]&~m[606]&~m[862])|(~m[90]&m[606]&m[862]))&~BiasedRNG[235])|((~m[90]&~m[606]&m[862])|(m[90]&~m[606]&m[862])|(m[90]&m[606]&m[862]));
    m[396] = (((~m[91]&~m[622]&~m[878])|(m[91]&m[622]&~m[878]))&BiasedRNG[236])|(((m[91]&~m[622]&~m[878])|(~m[91]&m[622]&m[878]))&~BiasedRNG[236])|((~m[91]&~m[622]&m[878])|(m[91]&~m[622]&m[878])|(m[91]&m[622]&m[878]));
    m[397] = (((~m[91]&~m[638]&~m[894])|(m[91]&m[638]&~m[894]))&BiasedRNG[237])|(((m[91]&~m[638]&~m[894])|(~m[91]&m[638]&m[894]))&~BiasedRNG[237])|((~m[91]&~m[638]&m[894])|(m[91]&~m[638]&m[894])|(m[91]&m[638]&m[894]));
    m[398] = (((~m[91]&~m[654]&~m[910])|(m[91]&m[654]&~m[910]))&BiasedRNG[238])|(((m[91]&~m[654]&~m[910])|(~m[91]&m[654]&m[910]))&~BiasedRNG[238])|((~m[91]&~m[654]&m[910])|(m[91]&~m[654]&m[910])|(m[91]&m[654]&m[910]));
    m[399] = (((~m[91]&~m[670]&~m[926])|(m[91]&m[670]&~m[926]))&BiasedRNG[239])|(((m[91]&~m[670]&~m[926])|(~m[91]&m[670]&m[926]))&~BiasedRNG[239])|((~m[91]&~m[670]&m[926])|(m[91]&~m[670]&m[926])|(m[91]&m[670]&m[926]));
    m[400] = (((~m[92]&~m[431]&~m[687])|(m[92]&m[431]&~m[687]))&BiasedRNG[240])|(((m[92]&~m[431]&~m[687])|(~m[92]&m[431]&m[687]))&~BiasedRNG[240])|((~m[92]&~m[431]&m[687])|(m[92]&~m[431]&m[687])|(m[92]&m[431]&m[687]));
    m[401] = (((~m[92]&~m[447]&~m[703])|(m[92]&m[447]&~m[703]))&BiasedRNG[241])|(((m[92]&~m[447]&~m[703])|(~m[92]&m[447]&m[703]))&~BiasedRNG[241])|((~m[92]&~m[447]&m[703])|(m[92]&~m[447]&m[703])|(m[92]&m[447]&m[703]));
    m[402] = (((~m[92]&~m[463]&~m[719])|(m[92]&m[463]&~m[719]))&BiasedRNG[242])|(((m[92]&~m[463]&~m[719])|(~m[92]&m[463]&m[719]))&~BiasedRNG[242])|((~m[92]&~m[463]&m[719])|(m[92]&~m[463]&m[719])|(m[92]&m[463]&m[719]));
    m[403] = (((~m[92]&~m[479]&~m[735])|(m[92]&m[479]&~m[735]))&BiasedRNG[243])|(((m[92]&~m[479]&~m[735])|(~m[92]&m[479]&m[735]))&~BiasedRNG[243])|((~m[92]&~m[479]&m[735])|(m[92]&~m[479]&m[735])|(m[92]&m[479]&m[735]));
    m[404] = (((~m[93]&~m[495]&~m[751])|(m[93]&m[495]&~m[751]))&BiasedRNG[244])|(((m[93]&~m[495]&~m[751])|(~m[93]&m[495]&m[751]))&~BiasedRNG[244])|((~m[93]&~m[495]&m[751])|(m[93]&~m[495]&m[751])|(m[93]&m[495]&m[751]));
    m[405] = (((~m[93]&~m[511]&~m[767])|(m[93]&m[511]&~m[767]))&BiasedRNG[245])|(((m[93]&~m[511]&~m[767])|(~m[93]&m[511]&m[767]))&~BiasedRNG[245])|((~m[93]&~m[511]&m[767])|(m[93]&~m[511]&m[767])|(m[93]&m[511]&m[767]));
    m[406] = (((~m[93]&~m[527]&~m[783])|(m[93]&m[527]&~m[783]))&BiasedRNG[246])|(((m[93]&~m[527]&~m[783])|(~m[93]&m[527]&m[783]))&~BiasedRNG[246])|((~m[93]&~m[527]&m[783])|(m[93]&~m[527]&m[783])|(m[93]&m[527]&m[783]));
    m[407] = (((~m[93]&~m[543]&~m[799])|(m[93]&m[543]&~m[799]))&BiasedRNG[247])|(((m[93]&~m[543]&~m[799])|(~m[93]&m[543]&m[799]))&~BiasedRNG[247])|((~m[93]&~m[543]&m[799])|(m[93]&~m[543]&m[799])|(m[93]&m[543]&m[799]));
    m[408] = (((~m[94]&~m[559]&~m[815])|(m[94]&m[559]&~m[815]))&BiasedRNG[248])|(((m[94]&~m[559]&~m[815])|(~m[94]&m[559]&m[815]))&~BiasedRNG[248])|((~m[94]&~m[559]&m[815])|(m[94]&~m[559]&m[815])|(m[94]&m[559]&m[815]));
    m[409] = (((~m[94]&~m[575]&~m[831])|(m[94]&m[575]&~m[831]))&BiasedRNG[249])|(((m[94]&~m[575]&~m[831])|(~m[94]&m[575]&m[831]))&~BiasedRNG[249])|((~m[94]&~m[575]&m[831])|(m[94]&~m[575]&m[831])|(m[94]&m[575]&m[831]));
    m[410] = (((~m[94]&~m[591]&~m[847])|(m[94]&m[591]&~m[847]))&BiasedRNG[250])|(((m[94]&~m[591]&~m[847])|(~m[94]&m[591]&m[847]))&~BiasedRNG[250])|((~m[94]&~m[591]&m[847])|(m[94]&~m[591]&m[847])|(m[94]&m[591]&m[847]));
    m[411] = (((~m[94]&~m[607]&~m[863])|(m[94]&m[607]&~m[863]))&BiasedRNG[251])|(((m[94]&~m[607]&~m[863])|(~m[94]&m[607]&m[863]))&~BiasedRNG[251])|((~m[94]&~m[607]&m[863])|(m[94]&~m[607]&m[863])|(m[94]&m[607]&m[863]));
    m[412] = (((~m[95]&~m[623]&~m[879])|(m[95]&m[623]&~m[879]))&BiasedRNG[252])|(((m[95]&~m[623]&~m[879])|(~m[95]&m[623]&m[879]))&~BiasedRNG[252])|((~m[95]&~m[623]&m[879])|(m[95]&~m[623]&m[879])|(m[95]&m[623]&m[879]));
    m[413] = (((~m[95]&~m[639]&~m[895])|(m[95]&m[639]&~m[895]))&BiasedRNG[253])|(((m[95]&~m[639]&~m[895])|(~m[95]&m[639]&m[895]))&~BiasedRNG[253])|((~m[95]&~m[639]&m[895])|(m[95]&~m[639]&m[895])|(m[95]&m[639]&m[895]));
    m[414] = (((~m[95]&~m[655]&~m[911])|(m[95]&m[655]&~m[911]))&BiasedRNG[254])|(((m[95]&~m[655]&~m[911])|(~m[95]&m[655]&m[911]))&~BiasedRNG[254])|((~m[95]&~m[655]&m[911])|(m[95]&~m[655]&m[911])|(m[95]&m[655]&m[911]));
    m[415] = (((~m[95]&~m[671]&~m[927])|(m[95]&m[671]&~m[927]))&BiasedRNG[255])|(((m[95]&~m[671]&~m[927])|(~m[95]&m[671]&m[927]))&~BiasedRNG[255])|((~m[95]&~m[671]&m[927])|(m[95]&~m[671]&m[927])|(m[95]&m[671]&m[927]));
    m[928] = (((m[673]&~m[929]&~m[930]&~m[931]&~m[932])|(~m[673]&~m[929]&~m[930]&m[931]&~m[932])|(m[673]&m[929]&~m[930]&m[931]&~m[932])|(m[673]&~m[929]&m[930]&m[931]&~m[932])|(~m[673]&m[929]&~m[930]&~m[931]&m[932])|(~m[673]&~m[929]&m[930]&~m[931]&m[932])|(m[673]&m[929]&m[930]&~m[931]&m[932])|(~m[673]&m[929]&m[930]&m[931]&m[932]))&UnbiasedRNG[32])|((m[673]&~m[929]&~m[930]&m[931]&~m[932])|(~m[673]&~m[929]&~m[930]&~m[931]&m[932])|(m[673]&~m[929]&~m[930]&~m[931]&m[932])|(m[673]&m[929]&~m[930]&~m[931]&m[932])|(m[673]&~m[929]&m[930]&~m[931]&m[932])|(~m[673]&~m[929]&~m[930]&m[931]&m[932])|(m[673]&~m[929]&~m[930]&m[931]&m[932])|(~m[673]&m[929]&~m[930]&m[931]&m[932])|(m[673]&m[929]&~m[930]&m[931]&m[932])|(~m[673]&~m[929]&m[930]&m[931]&m[932])|(m[673]&~m[929]&m[930]&m[931]&m[932])|(m[673]&m[929]&m[930]&m[931]&m[932]));
    m[933] = (((m[674]&~m[934]&~m[935]&~m[936]&~m[937])|(~m[674]&~m[934]&~m[935]&m[936]&~m[937])|(m[674]&m[934]&~m[935]&m[936]&~m[937])|(m[674]&~m[934]&m[935]&m[936]&~m[937])|(~m[674]&m[934]&~m[935]&~m[936]&m[937])|(~m[674]&~m[934]&m[935]&~m[936]&m[937])|(m[674]&m[934]&m[935]&~m[936]&m[937])|(~m[674]&m[934]&m[935]&m[936]&m[937]))&UnbiasedRNG[33])|((m[674]&~m[934]&~m[935]&m[936]&~m[937])|(~m[674]&~m[934]&~m[935]&~m[936]&m[937])|(m[674]&~m[934]&~m[935]&~m[936]&m[937])|(m[674]&m[934]&~m[935]&~m[936]&m[937])|(m[674]&~m[934]&m[935]&~m[936]&m[937])|(~m[674]&~m[934]&~m[935]&m[936]&m[937])|(m[674]&~m[934]&~m[935]&m[936]&m[937])|(~m[674]&m[934]&~m[935]&m[936]&m[937])|(m[674]&m[934]&~m[935]&m[936]&m[937])|(~m[674]&~m[934]&m[935]&m[936]&m[937])|(m[674]&~m[934]&m[935]&m[936]&m[937])|(m[674]&m[934]&m[935]&m[936]&m[937]));
    m[938] = (((m[936]&~m[939]&~m[940]&~m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&m[941]&~m[942])|(m[936]&m[939]&~m[940]&m[941]&~m[942])|(m[936]&~m[939]&m[940]&m[941]&~m[942])|(~m[936]&m[939]&~m[940]&~m[941]&m[942])|(~m[936]&~m[939]&m[940]&~m[941]&m[942])|(m[936]&m[939]&m[940]&~m[941]&m[942])|(~m[936]&m[939]&m[940]&m[941]&m[942]))&UnbiasedRNG[34])|((m[936]&~m[939]&~m[940]&m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&m[940]&~m[941]&m[942])|(~m[936]&~m[939]&~m[940]&m[941]&m[942])|(m[936]&~m[939]&~m[940]&m[941]&m[942])|(~m[936]&m[939]&~m[940]&m[941]&m[942])|(m[936]&m[939]&~m[940]&m[941]&m[942])|(~m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&m[939]&m[940]&m[941]&m[942]));
    m[943] = (((m[675]&~m[944]&~m[945]&~m[946]&~m[947])|(~m[675]&~m[944]&~m[945]&m[946]&~m[947])|(m[675]&m[944]&~m[945]&m[946]&~m[947])|(m[675]&~m[944]&m[945]&m[946]&~m[947])|(~m[675]&m[944]&~m[945]&~m[946]&m[947])|(~m[675]&~m[944]&m[945]&~m[946]&m[947])|(m[675]&m[944]&m[945]&~m[946]&m[947])|(~m[675]&m[944]&m[945]&m[946]&m[947]))&UnbiasedRNG[35])|((m[675]&~m[944]&~m[945]&m[946]&~m[947])|(~m[675]&~m[944]&~m[945]&~m[946]&m[947])|(m[675]&~m[944]&~m[945]&~m[946]&m[947])|(m[675]&m[944]&~m[945]&~m[946]&m[947])|(m[675]&~m[944]&m[945]&~m[946]&m[947])|(~m[675]&~m[944]&~m[945]&m[946]&m[947])|(m[675]&~m[944]&~m[945]&m[946]&m[947])|(~m[675]&m[944]&~m[945]&m[946]&m[947])|(m[675]&m[944]&~m[945]&m[946]&m[947])|(~m[675]&~m[944]&m[945]&m[946]&m[947])|(m[675]&~m[944]&m[945]&m[946]&m[947])|(m[675]&m[944]&m[945]&m[946]&m[947]));
    m[948] = (((m[946]&~m[949]&~m[950]&~m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&m[951]&~m[952])|(m[946]&m[949]&~m[950]&m[951]&~m[952])|(m[946]&~m[949]&m[950]&m[951]&~m[952])|(~m[946]&m[949]&~m[950]&~m[951]&m[952])|(~m[946]&~m[949]&m[950]&~m[951]&m[952])|(m[946]&m[949]&m[950]&~m[951]&m[952])|(~m[946]&m[949]&m[950]&m[951]&m[952]))&UnbiasedRNG[36])|((m[946]&~m[949]&~m[950]&m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&m[950]&~m[951]&m[952])|(~m[946]&~m[949]&~m[950]&m[951]&m[952])|(m[946]&~m[949]&~m[950]&m[951]&m[952])|(~m[946]&m[949]&~m[950]&m[951]&m[952])|(m[946]&m[949]&~m[950]&m[951]&m[952])|(~m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&m[949]&m[950]&m[951]&m[952]));
    m[953] = (((m[951]&~m[954]&~m[955]&~m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&m[956]&~m[957])|(m[951]&m[954]&~m[955]&m[956]&~m[957])|(m[951]&~m[954]&m[955]&m[956]&~m[957])|(~m[951]&m[954]&~m[955]&~m[956]&m[957])|(~m[951]&~m[954]&m[955]&~m[956]&m[957])|(m[951]&m[954]&m[955]&~m[956]&m[957])|(~m[951]&m[954]&m[955]&m[956]&m[957]))&UnbiasedRNG[37])|((m[951]&~m[954]&~m[955]&m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&m[955]&~m[956]&m[957])|(~m[951]&~m[954]&~m[955]&m[956]&m[957])|(m[951]&~m[954]&~m[955]&m[956]&m[957])|(~m[951]&m[954]&~m[955]&m[956]&m[957])|(m[951]&m[954]&~m[955]&m[956]&m[957])|(~m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&m[954]&m[955]&m[956]&m[957]));
    m[958] = (((m[676]&~m[959]&~m[960]&~m[961]&~m[962])|(~m[676]&~m[959]&~m[960]&m[961]&~m[962])|(m[676]&m[959]&~m[960]&m[961]&~m[962])|(m[676]&~m[959]&m[960]&m[961]&~m[962])|(~m[676]&m[959]&~m[960]&~m[961]&m[962])|(~m[676]&~m[959]&m[960]&~m[961]&m[962])|(m[676]&m[959]&m[960]&~m[961]&m[962])|(~m[676]&m[959]&m[960]&m[961]&m[962]))&UnbiasedRNG[38])|((m[676]&~m[959]&~m[960]&m[961]&~m[962])|(~m[676]&~m[959]&~m[960]&~m[961]&m[962])|(m[676]&~m[959]&~m[960]&~m[961]&m[962])|(m[676]&m[959]&~m[960]&~m[961]&m[962])|(m[676]&~m[959]&m[960]&~m[961]&m[962])|(~m[676]&~m[959]&~m[960]&m[961]&m[962])|(m[676]&~m[959]&~m[960]&m[961]&m[962])|(~m[676]&m[959]&~m[960]&m[961]&m[962])|(m[676]&m[959]&~m[960]&m[961]&m[962])|(~m[676]&~m[959]&m[960]&m[961]&m[962])|(m[676]&~m[959]&m[960]&m[961]&m[962])|(m[676]&m[959]&m[960]&m[961]&m[962]));
    m[963] = (((m[961]&~m[964]&~m[965]&~m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&m[966]&~m[967])|(m[961]&m[964]&~m[965]&m[966]&~m[967])|(m[961]&~m[964]&m[965]&m[966]&~m[967])|(~m[961]&m[964]&~m[965]&~m[966]&m[967])|(~m[961]&~m[964]&m[965]&~m[966]&m[967])|(m[961]&m[964]&m[965]&~m[966]&m[967])|(~m[961]&m[964]&m[965]&m[966]&m[967]))&UnbiasedRNG[39])|((m[961]&~m[964]&~m[965]&m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&m[965]&~m[966]&m[967])|(~m[961]&~m[964]&~m[965]&m[966]&m[967])|(m[961]&~m[964]&~m[965]&m[966]&m[967])|(~m[961]&m[964]&~m[965]&m[966]&m[967])|(m[961]&m[964]&~m[965]&m[966]&m[967])|(~m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&m[964]&m[965]&m[966]&m[967]));
    m[968] = (((m[966]&~m[969]&~m[970]&~m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&m[971]&~m[972])|(m[966]&m[969]&~m[970]&m[971]&~m[972])|(m[966]&~m[969]&m[970]&m[971]&~m[972])|(~m[966]&m[969]&~m[970]&~m[971]&m[972])|(~m[966]&~m[969]&m[970]&~m[971]&m[972])|(m[966]&m[969]&m[970]&~m[971]&m[972])|(~m[966]&m[969]&m[970]&m[971]&m[972]))&UnbiasedRNG[40])|((m[966]&~m[969]&~m[970]&m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&m[970]&~m[971]&m[972])|(~m[966]&~m[969]&~m[970]&m[971]&m[972])|(m[966]&~m[969]&~m[970]&m[971]&m[972])|(~m[966]&m[969]&~m[970]&m[971]&m[972])|(m[966]&m[969]&~m[970]&m[971]&m[972])|(~m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&m[969]&m[970]&m[971]&m[972]));
    m[973] = (((m[971]&~m[974]&~m[975]&~m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&m[976]&~m[977])|(m[971]&m[974]&~m[975]&m[976]&~m[977])|(m[971]&~m[974]&m[975]&m[976]&~m[977])|(~m[971]&m[974]&~m[975]&~m[976]&m[977])|(~m[971]&~m[974]&m[975]&~m[976]&m[977])|(m[971]&m[974]&m[975]&~m[976]&m[977])|(~m[971]&m[974]&m[975]&m[976]&m[977]))&UnbiasedRNG[41])|((m[971]&~m[974]&~m[975]&m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&m[975]&~m[976]&m[977])|(~m[971]&~m[974]&~m[975]&m[976]&m[977])|(m[971]&~m[974]&~m[975]&m[976]&m[977])|(~m[971]&m[974]&~m[975]&m[976]&m[977])|(m[971]&m[974]&~m[975]&m[976]&m[977])|(~m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&m[974]&m[975]&m[976]&m[977]));
    m[978] = (((m[677]&~m[979]&~m[980]&~m[981]&~m[982])|(~m[677]&~m[979]&~m[980]&m[981]&~m[982])|(m[677]&m[979]&~m[980]&m[981]&~m[982])|(m[677]&~m[979]&m[980]&m[981]&~m[982])|(~m[677]&m[979]&~m[980]&~m[981]&m[982])|(~m[677]&~m[979]&m[980]&~m[981]&m[982])|(m[677]&m[979]&m[980]&~m[981]&m[982])|(~m[677]&m[979]&m[980]&m[981]&m[982]))&UnbiasedRNG[42])|((m[677]&~m[979]&~m[980]&m[981]&~m[982])|(~m[677]&~m[979]&~m[980]&~m[981]&m[982])|(m[677]&~m[979]&~m[980]&~m[981]&m[982])|(m[677]&m[979]&~m[980]&~m[981]&m[982])|(m[677]&~m[979]&m[980]&~m[981]&m[982])|(~m[677]&~m[979]&~m[980]&m[981]&m[982])|(m[677]&~m[979]&~m[980]&m[981]&m[982])|(~m[677]&m[979]&~m[980]&m[981]&m[982])|(m[677]&m[979]&~m[980]&m[981]&m[982])|(~m[677]&~m[979]&m[980]&m[981]&m[982])|(m[677]&~m[979]&m[980]&m[981]&m[982])|(m[677]&m[979]&m[980]&m[981]&m[982]));
    m[983] = (((m[981]&~m[984]&~m[985]&~m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&m[986]&~m[987])|(m[981]&m[984]&~m[985]&m[986]&~m[987])|(m[981]&~m[984]&m[985]&m[986]&~m[987])|(~m[981]&m[984]&~m[985]&~m[986]&m[987])|(~m[981]&~m[984]&m[985]&~m[986]&m[987])|(m[981]&m[984]&m[985]&~m[986]&m[987])|(~m[981]&m[984]&m[985]&m[986]&m[987]))&UnbiasedRNG[43])|((m[981]&~m[984]&~m[985]&m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&m[985]&~m[986]&m[987])|(~m[981]&~m[984]&~m[985]&m[986]&m[987])|(m[981]&~m[984]&~m[985]&m[986]&m[987])|(~m[981]&m[984]&~m[985]&m[986]&m[987])|(m[981]&m[984]&~m[985]&m[986]&m[987])|(~m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&m[984]&m[985]&m[986]&m[987]));
    m[988] = (((m[986]&~m[989]&~m[990]&~m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&m[991]&~m[992])|(m[986]&m[989]&~m[990]&m[991]&~m[992])|(m[986]&~m[989]&m[990]&m[991]&~m[992])|(~m[986]&m[989]&~m[990]&~m[991]&m[992])|(~m[986]&~m[989]&m[990]&~m[991]&m[992])|(m[986]&m[989]&m[990]&~m[991]&m[992])|(~m[986]&m[989]&m[990]&m[991]&m[992]))&UnbiasedRNG[44])|((m[986]&~m[989]&~m[990]&m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&m[990]&~m[991]&m[992])|(~m[986]&~m[989]&~m[990]&m[991]&m[992])|(m[986]&~m[989]&~m[990]&m[991]&m[992])|(~m[986]&m[989]&~m[990]&m[991]&m[992])|(m[986]&m[989]&~m[990]&m[991]&m[992])|(~m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&m[989]&m[990]&m[991]&m[992]));
    m[993] = (((m[991]&~m[994]&~m[995]&~m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&m[996]&~m[997])|(m[991]&m[994]&~m[995]&m[996]&~m[997])|(m[991]&~m[994]&m[995]&m[996]&~m[997])|(~m[991]&m[994]&~m[995]&~m[996]&m[997])|(~m[991]&~m[994]&m[995]&~m[996]&m[997])|(m[991]&m[994]&m[995]&~m[996]&m[997])|(~m[991]&m[994]&m[995]&m[996]&m[997]))&UnbiasedRNG[45])|((m[991]&~m[994]&~m[995]&m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&m[995]&~m[996]&m[997])|(~m[991]&~m[994]&~m[995]&m[996]&m[997])|(m[991]&~m[994]&~m[995]&m[996]&m[997])|(~m[991]&m[994]&~m[995]&m[996]&m[997])|(m[991]&m[994]&~m[995]&m[996]&m[997])|(~m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&m[994]&m[995]&m[996]&m[997]));
    m[998] = (((m[996]&~m[999]&~m[1000]&~m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&~m[1002])|(~m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&m[999]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[46])|((m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&m[999]&m[1000]&m[1001]&m[1002]));
    m[1003] = (((m[678]&~m[1004]&~m[1005]&~m[1006]&~m[1007])|(~m[678]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(m[678]&m[1004]&~m[1005]&m[1006]&~m[1007])|(m[678]&~m[1004]&m[1005]&m[1006]&~m[1007])|(~m[678]&m[1004]&~m[1005]&~m[1006]&m[1007])|(~m[678]&~m[1004]&m[1005]&~m[1006]&m[1007])|(m[678]&m[1004]&m[1005]&~m[1006]&m[1007])|(~m[678]&m[1004]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[47])|((m[678]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(~m[678]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[678]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[678]&m[1004]&~m[1005]&~m[1006]&m[1007])|(m[678]&~m[1004]&m[1005]&~m[1006]&m[1007])|(~m[678]&~m[1004]&~m[1005]&m[1006]&m[1007])|(m[678]&~m[1004]&~m[1005]&m[1006]&m[1007])|(~m[678]&m[1004]&~m[1005]&m[1006]&m[1007])|(m[678]&m[1004]&~m[1005]&m[1006]&m[1007])|(~m[678]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[678]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[678]&m[1004]&m[1005]&m[1006]&m[1007]));
    m[1008] = (((m[1006]&~m[1009]&~m[1010]&~m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&~m[1012])|(~m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&m[1009]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[48])|((m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&m[1011]&m[1012]));
    m[1013] = (((m[1011]&~m[1014]&~m[1015]&~m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&~m[1017])|(~m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[49])|((m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&m[1016]&m[1017]));
    m[1018] = (((m[1016]&~m[1019]&~m[1020]&~m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&~m[1022])|(~m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[50])|((m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&m[1021]&m[1022]));
    m[1023] = (((m[1021]&~m[1024]&~m[1025]&~m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&~m[1027])|(~m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[51])|((m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&m[1026]&m[1027]));
    m[1028] = (((m[1026]&~m[1029]&~m[1030]&~m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&~m[1032])|(~m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[52])|((m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&m[1031]&m[1032]));
    m[1033] = (((m[679]&~m[1034]&~m[1035]&~m[1036]&~m[1037])|(~m[679]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(m[679]&m[1034]&~m[1035]&m[1036]&~m[1037])|(m[679]&~m[1034]&m[1035]&m[1036]&~m[1037])|(~m[679]&m[1034]&~m[1035]&~m[1036]&m[1037])|(~m[679]&~m[1034]&m[1035]&~m[1036]&m[1037])|(m[679]&m[1034]&m[1035]&~m[1036]&m[1037])|(~m[679]&m[1034]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[53])|((m[679]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(~m[679]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[679]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[679]&m[1034]&~m[1035]&~m[1036]&m[1037])|(m[679]&~m[1034]&m[1035]&~m[1036]&m[1037])|(~m[679]&~m[1034]&~m[1035]&m[1036]&m[1037])|(m[679]&~m[1034]&~m[1035]&m[1036]&m[1037])|(~m[679]&m[1034]&~m[1035]&m[1036]&m[1037])|(m[679]&m[1034]&~m[1035]&m[1036]&m[1037])|(~m[679]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[679]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[679]&m[1034]&m[1035]&m[1036]&m[1037]));
    m[1038] = (((m[1036]&~m[1039]&~m[1040]&~m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&~m[1042])|(~m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[54])|((m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&m[1041]&m[1042]));
    m[1043] = (((m[1041]&~m[1044]&~m[1045]&~m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&~m[1047])|(~m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[55])|((m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&m[1046]&m[1047]));
    m[1048] = (((m[1046]&~m[1049]&~m[1050]&~m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&~m[1052])|(~m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&m[1049]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[56])|((m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&m[1051]&m[1052]));
    m[1053] = (((m[1051]&~m[1054]&~m[1055]&~m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&~m[1057])|(~m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[57])|((m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&m[1056]&m[1057]));
    m[1058] = (((m[1056]&~m[1059]&~m[1060]&~m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&~m[1062])|(~m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&m[1059]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[58])|((m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&m[1061]&m[1062]));
    m[1063] = (((m[1061]&~m[1064]&~m[1065]&~m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&~m[1067])|(~m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[59])|((m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&m[1066]&m[1067]));
    m[1068] = (((m[680]&~m[1069]&~m[1070]&~m[1071]&~m[1072])|(~m[680]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(m[680]&m[1069]&~m[1070]&m[1071]&~m[1072])|(m[680]&~m[1069]&m[1070]&m[1071]&~m[1072])|(~m[680]&m[1069]&~m[1070]&~m[1071]&m[1072])|(~m[680]&~m[1069]&m[1070]&~m[1071]&m[1072])|(m[680]&m[1069]&m[1070]&~m[1071]&m[1072])|(~m[680]&m[1069]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[60])|((m[680]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(~m[680]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[680]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[680]&m[1069]&~m[1070]&~m[1071]&m[1072])|(m[680]&~m[1069]&m[1070]&~m[1071]&m[1072])|(~m[680]&~m[1069]&~m[1070]&m[1071]&m[1072])|(m[680]&~m[1069]&~m[1070]&m[1071]&m[1072])|(~m[680]&m[1069]&~m[1070]&m[1071]&m[1072])|(m[680]&m[1069]&~m[1070]&m[1071]&m[1072])|(~m[680]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[680]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[680]&m[1069]&m[1070]&m[1071]&m[1072]));
    m[1073] = (((m[1071]&~m[1074]&~m[1075]&~m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&~m[1077])|(~m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[61])|((m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&m[1076]&m[1077]));
    m[1078] = (((m[1076]&~m[1079]&~m[1080]&~m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&~m[1082])|(~m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[62])|((m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&m[1081]&m[1082]));
    m[1083] = (((m[1081]&~m[1084]&~m[1085]&~m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&~m[1087])|(~m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&m[1084]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[63])|((m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&m[1086]&m[1087]));
    m[1088] = (((m[1086]&~m[1089]&~m[1090]&~m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&~m[1092])|(~m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[64])|((m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&m[1091]&m[1092]));
    m[1093] = (((m[1091]&~m[1094]&~m[1095]&~m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&~m[1097])|(~m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[65])|((m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&m[1096]&m[1097]));
    m[1098] = (((m[1096]&~m[1099]&~m[1100]&~m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&~m[1102])|(~m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[66])|((m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&m[1101]&m[1102]));
    m[1103] = (((m[1101]&~m[1104]&~m[1105]&~m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&~m[1107])|(~m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[67])|((m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&m[1106]&m[1107]));
    m[1108] = (((m[681]&~m[1109]&~m[1110]&~m[1111]&~m[1112])|(~m[681]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(m[681]&m[1109]&~m[1110]&m[1111]&~m[1112])|(m[681]&~m[1109]&m[1110]&m[1111]&~m[1112])|(~m[681]&m[1109]&~m[1110]&~m[1111]&m[1112])|(~m[681]&~m[1109]&m[1110]&~m[1111]&m[1112])|(m[681]&m[1109]&m[1110]&~m[1111]&m[1112])|(~m[681]&m[1109]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[68])|((m[681]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(~m[681]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[681]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[681]&m[1109]&~m[1110]&~m[1111]&m[1112])|(m[681]&~m[1109]&m[1110]&~m[1111]&m[1112])|(~m[681]&~m[1109]&~m[1110]&m[1111]&m[1112])|(m[681]&~m[1109]&~m[1110]&m[1111]&m[1112])|(~m[681]&m[1109]&~m[1110]&m[1111]&m[1112])|(m[681]&m[1109]&~m[1110]&m[1111]&m[1112])|(~m[681]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[681]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[681]&m[1109]&m[1110]&m[1111]&m[1112]));
    m[1113] = (((m[1111]&~m[1114]&~m[1115]&~m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&~m[1117])|(~m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&m[1114]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[69])|((m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&m[1116]&m[1117]));
    m[1118] = (((m[1116]&~m[1119]&~m[1120]&~m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&~m[1122])|(~m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&m[1119]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[70])|((m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&m[1121]&m[1122]));
    m[1123] = (((m[1121]&~m[1124]&~m[1125]&~m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&~m[1127])|(~m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[71])|((m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&m[1126]&m[1127]));
    m[1128] = (((m[1126]&~m[1129]&~m[1130]&~m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&~m[1132])|(~m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[72])|((m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&m[1131]&m[1132]));
    m[1133] = (((m[1131]&~m[1134]&~m[1135]&~m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&~m[1137])|(~m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[73])|((m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&m[1136]&m[1137]));
    m[1138] = (((m[1136]&~m[1139]&~m[1140]&~m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&~m[1142])|(~m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&m[1139]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[74])|((m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&m[1141]&m[1142]));
    m[1143] = (((m[1141]&~m[1144]&~m[1145]&~m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&~m[1147])|(~m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[75])|((m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&m[1146]&m[1147]));
    m[1148] = (((m[1146]&~m[1149]&~m[1150]&~m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&~m[1152])|(~m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[76])|((m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&m[1151]&m[1152]));
    m[1153] = (((m[682]&~m[1154]&~m[1155]&~m[1156]&~m[1157])|(~m[682]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(m[682]&m[1154]&~m[1155]&m[1156]&~m[1157])|(m[682]&~m[1154]&m[1155]&m[1156]&~m[1157])|(~m[682]&m[1154]&~m[1155]&~m[1156]&m[1157])|(~m[682]&~m[1154]&m[1155]&~m[1156]&m[1157])|(m[682]&m[1154]&m[1155]&~m[1156]&m[1157])|(~m[682]&m[1154]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[77])|((m[682]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(~m[682]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[682]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[682]&m[1154]&~m[1155]&~m[1156]&m[1157])|(m[682]&~m[1154]&m[1155]&~m[1156]&m[1157])|(~m[682]&~m[1154]&~m[1155]&m[1156]&m[1157])|(m[682]&~m[1154]&~m[1155]&m[1156]&m[1157])|(~m[682]&m[1154]&~m[1155]&m[1156]&m[1157])|(m[682]&m[1154]&~m[1155]&m[1156]&m[1157])|(~m[682]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[682]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[682]&m[1154]&m[1155]&m[1156]&m[1157]));
    m[1158] = (((m[1156]&~m[1159]&~m[1160]&~m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&~m[1162])|(~m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&m[1159]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[78])|((m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&m[1161]&m[1162]));
    m[1163] = (((m[1161]&~m[1164]&~m[1165]&~m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&~m[1167])|(~m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[79])|((m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&m[1166]&m[1167]));
    m[1168] = (((m[1166]&~m[1169]&~m[1170]&~m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&~m[1172])|(~m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[80])|((m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&m[1171]&m[1172]));
    m[1173] = (((m[1171]&~m[1174]&~m[1175]&~m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&~m[1177])|(~m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&m[1174]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[81])|((m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&m[1176]&m[1177]));
    m[1178] = (((m[1176]&~m[1179]&~m[1180]&~m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&~m[1182])|(~m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[82])|((m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&m[1181]&m[1182]));
    m[1183] = (((m[1181]&~m[1184]&~m[1185]&~m[1186]&~m[1187])|(~m[1181]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1181]&m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1181]&~m[1184]&m[1185]&m[1186]&~m[1187])|(~m[1181]&m[1184]&~m[1185]&~m[1186]&m[1187])|(~m[1181]&~m[1184]&m[1185]&~m[1186]&m[1187])|(m[1181]&m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1181]&m[1184]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[83])|((m[1181]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(~m[1181]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1181]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1181]&m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1181]&~m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1181]&~m[1184]&~m[1185]&m[1186]&m[1187])|(m[1181]&~m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1181]&m[1184]&~m[1185]&m[1186]&m[1187])|(m[1181]&m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1181]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1181]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1181]&m[1184]&m[1185]&m[1186]&m[1187]));
    m[1188] = (((m[1186]&~m[1189]&~m[1190]&~m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&~m[1192])|(~m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&m[1189]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[84])|((m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&m[1191]&m[1192]));
    m[1193] = (((m[1191]&~m[1194]&~m[1195]&~m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&~m[1197])|(~m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&m[1194]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[85])|((m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&m[1196]&m[1197]));
    m[1198] = (((m[1196]&~m[1199]&~m[1200]&~m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&~m[1202])|(~m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&m[1199]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[86])|((m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&m[1201]&m[1202]));
    m[1203] = (((m[683]&~m[1204]&~m[1205]&~m[1206]&~m[1207])|(~m[683]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(m[683]&m[1204]&~m[1205]&m[1206]&~m[1207])|(m[683]&~m[1204]&m[1205]&m[1206]&~m[1207])|(~m[683]&m[1204]&~m[1205]&~m[1206]&m[1207])|(~m[683]&~m[1204]&m[1205]&~m[1206]&m[1207])|(m[683]&m[1204]&m[1205]&~m[1206]&m[1207])|(~m[683]&m[1204]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[87])|((m[683]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(~m[683]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[683]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[683]&m[1204]&~m[1205]&~m[1206]&m[1207])|(m[683]&~m[1204]&m[1205]&~m[1206]&m[1207])|(~m[683]&~m[1204]&~m[1205]&m[1206]&m[1207])|(m[683]&~m[1204]&~m[1205]&m[1206]&m[1207])|(~m[683]&m[1204]&~m[1205]&m[1206]&m[1207])|(m[683]&m[1204]&~m[1205]&m[1206]&m[1207])|(~m[683]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[683]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[683]&m[1204]&m[1205]&m[1206]&m[1207]));
    m[1208] = (((m[1206]&~m[1209]&~m[1210]&~m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&~m[1212])|(~m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&m[1209]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[88])|((m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&m[1211]&m[1212]));
    m[1213] = (((m[1211]&~m[1214]&~m[1215]&~m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&~m[1217])|(~m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&m[1214]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[89])|((m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&m[1216]&m[1217]));
    m[1218] = (((m[1216]&~m[1219]&~m[1220]&~m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&~m[1222])|(~m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&m[1219]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[90])|((m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&m[1221]&m[1222]));
    m[1223] = (((m[1221]&~m[1224]&~m[1225]&~m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&~m[1227])|(~m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&m[1224]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[91])|((m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&m[1226]&m[1227]));
    m[1228] = (((m[1226]&~m[1229]&~m[1230]&~m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&~m[1232])|(~m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&m[1229]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[92])|((m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&m[1231]&m[1232]));
    m[1233] = (((m[1231]&~m[1234]&~m[1235]&~m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&~m[1237])|(~m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&m[1234]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[93])|((m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&m[1236]&m[1237]));
    m[1238] = (((m[1236]&~m[1239]&~m[1240]&~m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&~m[1242])|(~m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&m[1239]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[94])|((m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&m[1241]&m[1242]));
    m[1243] = (((m[1241]&~m[1244]&~m[1245]&~m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&~m[1247])|(~m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&m[1244]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[95])|((m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&m[1246]&m[1247]));
    m[1248] = (((m[1246]&~m[1249]&~m[1250]&~m[1251]&~m[1252])|(~m[1246]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1246]&m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1246]&~m[1249]&m[1250]&m[1251]&~m[1252])|(~m[1246]&m[1249]&~m[1250]&~m[1251]&m[1252])|(~m[1246]&~m[1249]&m[1250]&~m[1251]&m[1252])|(m[1246]&m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1246]&m[1249]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[96])|((m[1246]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(~m[1246]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1246]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1246]&m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1246]&~m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1246]&~m[1249]&~m[1250]&m[1251]&m[1252])|(m[1246]&~m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1246]&m[1249]&~m[1250]&m[1251]&m[1252])|(m[1246]&m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1246]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1246]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1246]&m[1249]&m[1250]&m[1251]&m[1252]));
    m[1253] = (((m[1251]&~m[1254]&~m[1255]&~m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&~m[1257])|(~m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&m[1254]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[97])|((m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&m[1256]&m[1257]));
    m[1258] = (((m[684]&~m[1259]&~m[1260]&~m[1261]&~m[1262])|(~m[684]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(m[684]&m[1259]&~m[1260]&m[1261]&~m[1262])|(m[684]&~m[1259]&m[1260]&m[1261]&~m[1262])|(~m[684]&m[1259]&~m[1260]&~m[1261]&m[1262])|(~m[684]&~m[1259]&m[1260]&~m[1261]&m[1262])|(m[684]&m[1259]&m[1260]&~m[1261]&m[1262])|(~m[684]&m[1259]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[98])|((m[684]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(~m[684]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[684]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[684]&m[1259]&~m[1260]&~m[1261]&m[1262])|(m[684]&~m[1259]&m[1260]&~m[1261]&m[1262])|(~m[684]&~m[1259]&~m[1260]&m[1261]&m[1262])|(m[684]&~m[1259]&~m[1260]&m[1261]&m[1262])|(~m[684]&m[1259]&~m[1260]&m[1261]&m[1262])|(m[684]&m[1259]&~m[1260]&m[1261]&m[1262])|(~m[684]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[684]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[684]&m[1259]&m[1260]&m[1261]&m[1262]));
    m[1263] = (((m[1261]&~m[1264]&~m[1265]&~m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&~m[1267])|(~m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&m[1264]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[99])|((m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&m[1266]&m[1267]));
    m[1268] = (((m[1266]&~m[1269]&~m[1270]&~m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&~m[1272])|(~m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&m[1269]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[100])|((m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&m[1271]&m[1272]));
    m[1273] = (((m[1271]&~m[1274]&~m[1275]&~m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&~m[1277])|(~m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&m[1274]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[101])|((m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&m[1276]&m[1277]));
    m[1278] = (((m[1276]&~m[1279]&~m[1280]&~m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&~m[1282])|(~m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&m[1279]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[102])|((m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&m[1281]&m[1282]));
    m[1283] = (((m[1281]&~m[1284]&~m[1285]&~m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&~m[1287])|(~m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&m[1284]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[103])|((m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&m[1286]&m[1287]));
    m[1288] = (((m[1286]&~m[1289]&~m[1290]&~m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&~m[1292])|(~m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&m[1289]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[104])|((m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&m[1291]&m[1292]));
    m[1293] = (((m[1291]&~m[1294]&~m[1295]&~m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&~m[1297])|(~m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&m[1294]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[105])|((m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&m[1296]&m[1297]));
    m[1298] = (((m[1296]&~m[1299]&~m[1300]&~m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&~m[1302])|(~m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&m[1299]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[106])|((m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&m[1301]&m[1302]));
    m[1303] = (((m[1301]&~m[1304]&~m[1305]&~m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&~m[1307])|(~m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&m[1304]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[107])|((m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&m[1306]&m[1307]));
    m[1308] = (((m[1306]&~m[1309]&~m[1310]&~m[1311]&~m[1312])|(~m[1306]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1306]&m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1306]&~m[1309]&m[1310]&m[1311]&~m[1312])|(~m[1306]&m[1309]&~m[1310]&~m[1311]&m[1312])|(~m[1306]&~m[1309]&m[1310]&~m[1311]&m[1312])|(m[1306]&m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1306]&m[1309]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[108])|((m[1306]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(~m[1306]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1306]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1306]&m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1306]&~m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1306]&~m[1309]&~m[1310]&m[1311]&m[1312])|(m[1306]&~m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1306]&m[1309]&~m[1310]&m[1311]&m[1312])|(m[1306]&m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1306]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1306]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1306]&m[1309]&m[1310]&m[1311]&m[1312]));
    m[1313] = (((m[1311]&~m[1314]&~m[1315]&~m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&~m[1317])|(~m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&m[1314]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[109])|((m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&m[1316]&m[1317]));
    m[1318] = (((m[685]&~m[1319]&~m[1320]&~m[1321]&~m[1322])|(~m[685]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(m[685]&m[1319]&~m[1320]&m[1321]&~m[1322])|(m[685]&~m[1319]&m[1320]&m[1321]&~m[1322])|(~m[685]&m[1319]&~m[1320]&~m[1321]&m[1322])|(~m[685]&~m[1319]&m[1320]&~m[1321]&m[1322])|(m[685]&m[1319]&m[1320]&~m[1321]&m[1322])|(~m[685]&m[1319]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[110])|((m[685]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(~m[685]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[685]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[685]&m[1319]&~m[1320]&~m[1321]&m[1322])|(m[685]&~m[1319]&m[1320]&~m[1321]&m[1322])|(~m[685]&~m[1319]&~m[1320]&m[1321]&m[1322])|(m[685]&~m[1319]&~m[1320]&m[1321]&m[1322])|(~m[685]&m[1319]&~m[1320]&m[1321]&m[1322])|(m[685]&m[1319]&~m[1320]&m[1321]&m[1322])|(~m[685]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[685]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[685]&m[1319]&m[1320]&m[1321]&m[1322]));
    m[1323] = (((m[1321]&~m[1324]&~m[1325]&~m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&~m[1327])|(~m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&m[1324]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[111])|((m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&m[1326]&m[1327]));
    m[1328] = (((m[1326]&~m[1329]&~m[1330]&~m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&~m[1332])|(~m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&m[1329]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[112])|((m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&m[1331]&m[1332]));
    m[1333] = (((m[1331]&~m[1334]&~m[1335]&~m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&~m[1337])|(~m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&m[1334]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[113])|((m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&m[1336]&m[1337]));
    m[1338] = (((m[1336]&~m[1339]&~m[1340]&~m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&~m[1342])|(~m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&m[1339]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[114])|((m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&m[1341]&m[1342]));
    m[1343] = (((m[1341]&~m[1344]&~m[1345]&~m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&~m[1347])|(~m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&m[1344]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[115])|((m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&m[1346]&m[1347]));
    m[1348] = (((m[1346]&~m[1349]&~m[1350]&~m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&~m[1352])|(~m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&m[1349]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[116])|((m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&m[1351]&m[1352]));
    m[1353] = (((m[1351]&~m[1354]&~m[1355]&~m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&~m[1357])|(~m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&m[1354]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[117])|((m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&m[1356]&m[1357]));
    m[1358] = (((m[1356]&~m[1359]&~m[1360]&~m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&~m[1362])|(~m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&m[1359]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[118])|((m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&m[1361]&m[1362]));
    m[1363] = (((m[1361]&~m[1364]&~m[1365]&~m[1366]&~m[1367])|(~m[1361]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1361]&m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1361]&~m[1364]&m[1365]&m[1366]&~m[1367])|(~m[1361]&m[1364]&~m[1365]&~m[1366]&m[1367])|(~m[1361]&~m[1364]&m[1365]&~m[1366]&m[1367])|(m[1361]&m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1361]&m[1364]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[119])|((m[1361]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(~m[1361]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1361]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1361]&m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1361]&~m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1361]&~m[1364]&~m[1365]&m[1366]&m[1367])|(m[1361]&~m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1361]&m[1364]&~m[1365]&m[1366]&m[1367])|(m[1361]&m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1361]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1361]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1361]&m[1364]&m[1365]&m[1366]&m[1367]));
    m[1368] = (((m[1366]&~m[1369]&~m[1370]&~m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&~m[1372])|(~m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&m[1369]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[120])|((m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&m[1371]&m[1372]));
    m[1373] = (((m[1371]&~m[1374]&~m[1375]&~m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&~m[1377])|(~m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&m[1374]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[121])|((m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&m[1376]&m[1377]));
    m[1378] = (((m[1376]&~m[1379]&~m[1380]&~m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&~m[1382])|(~m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&m[1379]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[122])|((m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&m[1381]&m[1382]));
    m[1383] = (((m[686]&~m[1384]&~m[1385]&~m[1386]&~m[1387])|(~m[686]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(m[686]&m[1384]&~m[1385]&m[1386]&~m[1387])|(m[686]&~m[1384]&m[1385]&m[1386]&~m[1387])|(~m[686]&m[1384]&~m[1385]&~m[1386]&m[1387])|(~m[686]&~m[1384]&m[1385]&~m[1386]&m[1387])|(m[686]&m[1384]&m[1385]&~m[1386]&m[1387])|(~m[686]&m[1384]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[123])|((m[686]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(~m[686]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[686]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[686]&m[1384]&~m[1385]&~m[1386]&m[1387])|(m[686]&~m[1384]&m[1385]&~m[1386]&m[1387])|(~m[686]&~m[1384]&~m[1385]&m[1386]&m[1387])|(m[686]&~m[1384]&~m[1385]&m[1386]&m[1387])|(~m[686]&m[1384]&~m[1385]&m[1386]&m[1387])|(m[686]&m[1384]&~m[1385]&m[1386]&m[1387])|(~m[686]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[686]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[686]&m[1384]&m[1385]&m[1386]&m[1387]));
    m[1388] = (((m[1386]&~m[1389]&~m[1390]&~m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&~m[1392])|(~m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&m[1389]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[124])|((m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&m[1391]&m[1392]));
    m[1393] = (((m[1391]&~m[1394]&~m[1395]&~m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&~m[1397])|(~m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&m[1394]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[125])|((m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&m[1396]&m[1397]));
    m[1398] = (((m[1396]&~m[1399]&~m[1400]&~m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&~m[1402])|(~m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&m[1399]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[126])|((m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&m[1401]&m[1402]));
    m[1403] = (((m[1401]&~m[1404]&~m[1405]&~m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&~m[1407])|(~m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&m[1404]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[127])|((m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&m[1406]&m[1407]));
    m[1408] = (((m[1406]&~m[1409]&~m[1410]&~m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&~m[1412])|(~m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&m[1409]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[128])|((m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&m[1411]&m[1412]));
    m[1413] = (((m[1411]&~m[1414]&~m[1415]&~m[1416]&~m[1417])|(~m[1411]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1411]&m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1411]&~m[1414]&m[1415]&m[1416]&~m[1417])|(~m[1411]&m[1414]&~m[1415]&~m[1416]&m[1417])|(~m[1411]&~m[1414]&m[1415]&~m[1416]&m[1417])|(m[1411]&m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1411]&m[1414]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[129])|((m[1411]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(~m[1411]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1411]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1411]&m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1411]&~m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1411]&~m[1414]&~m[1415]&m[1416]&m[1417])|(m[1411]&~m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1411]&m[1414]&~m[1415]&m[1416]&m[1417])|(m[1411]&m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1411]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1411]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1411]&m[1414]&m[1415]&m[1416]&m[1417]));
    m[1418] = (((m[1416]&~m[1419]&~m[1420]&~m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&~m[1422])|(~m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&m[1419]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[130])|((m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&m[1421]&m[1422]));
    m[1423] = (((m[1421]&~m[1424]&~m[1425]&~m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&~m[1427])|(~m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&m[1424]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[131])|((m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&m[1426]&m[1427]));
    m[1428] = (((m[1426]&~m[1429]&~m[1430]&~m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&~m[1432])|(~m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&m[1429]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[132])|((m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&m[1431]&m[1432]));
    m[1433] = (((m[1431]&~m[1434]&~m[1435]&~m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&~m[1437])|(~m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&m[1434]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[133])|((m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&m[1436]&m[1437]));
    m[1438] = (((m[1436]&~m[1439]&~m[1440]&~m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&~m[1442])|(~m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&m[1439]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[134])|((m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&m[1441]&m[1442]));
    m[1443] = (((m[1441]&~m[1444]&~m[1445]&~m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&~m[1447])|(~m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&m[1444]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[135])|((m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&m[1446]&m[1447]));
    m[1448] = (((m[1446]&~m[1449]&~m[1450]&~m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&~m[1452])|(~m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&m[1449]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[136])|((m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&m[1451]&m[1452]));
    m[1453] = (((m[687]&~m[1454]&~m[1455]&~m[1456]&~m[1457])|(~m[687]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(m[687]&m[1454]&~m[1455]&m[1456]&~m[1457])|(m[687]&~m[1454]&m[1455]&m[1456]&~m[1457])|(~m[687]&m[1454]&~m[1455]&~m[1456]&m[1457])|(~m[687]&~m[1454]&m[1455]&~m[1456]&m[1457])|(m[687]&m[1454]&m[1455]&~m[1456]&m[1457])|(~m[687]&m[1454]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[137])|((m[687]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(~m[687]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[687]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[687]&m[1454]&~m[1455]&~m[1456]&m[1457])|(m[687]&~m[1454]&m[1455]&~m[1456]&m[1457])|(~m[687]&~m[1454]&~m[1455]&m[1456]&m[1457])|(m[687]&~m[1454]&~m[1455]&m[1456]&m[1457])|(~m[687]&m[1454]&~m[1455]&m[1456]&m[1457])|(m[687]&m[1454]&~m[1455]&m[1456]&m[1457])|(~m[687]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[687]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[687]&m[1454]&m[1455]&m[1456]&m[1457]));
    m[1458] = (((m[1456]&~m[1459]&~m[1460]&~m[1461]&~m[1462])|(~m[1456]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1456]&m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1456]&~m[1459]&m[1460]&m[1461]&~m[1462])|(~m[1456]&m[1459]&~m[1460]&~m[1461]&m[1462])|(~m[1456]&~m[1459]&m[1460]&~m[1461]&m[1462])|(m[1456]&m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1456]&m[1459]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[138])|((m[1456]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(~m[1456]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1456]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1456]&m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1456]&~m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1456]&~m[1459]&~m[1460]&m[1461]&m[1462])|(m[1456]&~m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1456]&m[1459]&~m[1460]&m[1461]&m[1462])|(m[1456]&m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1456]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1456]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1456]&m[1459]&m[1460]&m[1461]&m[1462]));
    m[1463] = (((m[1461]&~m[1464]&~m[1465]&~m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&~m[1467])|(~m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&m[1464]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[139])|((m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&m[1466]&m[1467]));
    m[1468] = (((m[1466]&~m[1469]&~m[1470]&~m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&~m[1472])|(~m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&m[1469]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[140])|((m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&m[1471]&m[1472]));
    m[1473] = (((m[1471]&~m[1474]&~m[1475]&~m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&~m[1477])|(~m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&m[1474]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[141])|((m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&m[1476]&m[1477]));
    m[1478] = (((m[1476]&~m[1479]&~m[1480]&~m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&~m[1482])|(~m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&m[1479]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[142])|((m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&m[1481]&m[1482]));
    m[1483] = (((m[1481]&~m[1484]&~m[1485]&~m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&~m[1487])|(~m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&m[1484]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[143])|((m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&m[1486]&m[1487]));
    m[1488] = (((m[1486]&~m[1489]&~m[1490]&~m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&~m[1492])|(~m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&m[1489]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[144])|((m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&m[1491]&m[1492]));
    m[1493] = (((m[1491]&~m[1494]&~m[1495]&~m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&~m[1497])|(~m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&m[1494]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[145])|((m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&m[1496]&m[1497]));
    m[1498] = (((m[1496]&~m[1499]&~m[1500]&~m[1501]&~m[1502])|(~m[1496]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1496]&m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1496]&~m[1499]&m[1500]&m[1501]&~m[1502])|(~m[1496]&m[1499]&~m[1500]&~m[1501]&m[1502])|(~m[1496]&~m[1499]&m[1500]&~m[1501]&m[1502])|(m[1496]&m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1496]&m[1499]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[146])|((m[1496]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(~m[1496]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1496]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1496]&m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1496]&~m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1496]&~m[1499]&~m[1500]&m[1501]&m[1502])|(m[1496]&~m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1496]&m[1499]&~m[1500]&m[1501]&m[1502])|(m[1496]&m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1496]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1496]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1496]&m[1499]&m[1500]&m[1501]&m[1502]));
    m[1503] = (((m[1501]&~m[1504]&~m[1505]&~m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&~m[1507])|(~m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&m[1504]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[147])|((m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&m[1506]&m[1507]));
    m[1508] = (((m[1506]&~m[1509]&~m[1510]&~m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&~m[1512])|(~m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&m[1509]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[148])|((m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&m[1511]&m[1512]));
    m[1513] = (((m[1511]&~m[1514]&~m[1515]&~m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&~m[1517])|(~m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&m[1514]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[149])|((m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&m[1516]&m[1517]));
    m[1518] = (((m[1516]&~m[1519]&~m[1520]&~m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&~m[1522])|(~m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&m[1519]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[150])|((m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&m[1521]&m[1522]));
    m[1523] = (((m[1521]&~m[1524]&~m[1525]&~m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&~m[1527])|(~m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&m[1524]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[151])|((m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&m[1526]&m[1527]));
    m[1533] = (((m[1531]&~m[1534]&~m[1535]&~m[1536]&~m[1537])|(~m[1531]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1531]&m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1531]&~m[1534]&m[1535]&m[1536]&~m[1537])|(~m[1531]&m[1534]&~m[1535]&~m[1536]&m[1537])|(~m[1531]&~m[1534]&m[1535]&~m[1536]&m[1537])|(m[1531]&m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1531]&m[1534]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[152])|((m[1531]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(~m[1531]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1531]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1531]&m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1531]&~m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1531]&~m[1534]&~m[1535]&m[1536]&m[1537])|(m[1531]&~m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1531]&m[1534]&~m[1535]&m[1536]&m[1537])|(m[1531]&m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1531]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1531]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1531]&m[1534]&m[1535]&m[1536]&m[1537]));
    m[1538] = (((m[1536]&~m[1539]&~m[1540]&~m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&~m[1542])|(~m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&m[1539]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[153])|((m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&m[1541]&m[1542]));
    m[1543] = (((m[1541]&~m[1544]&~m[1545]&~m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&~m[1547])|(~m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&m[1544]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[154])|((m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&m[1546]&m[1547]));
    m[1548] = (((m[1546]&~m[1549]&~m[1550]&~m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&~m[1552])|(~m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&m[1549]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[155])|((m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&m[1551]&m[1552]));
    m[1553] = (((m[1551]&~m[1554]&~m[1555]&~m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&~m[1557])|(~m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&m[1554]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[156])|((m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&m[1556]&m[1557]));
    m[1558] = (((m[1556]&~m[1559]&~m[1560]&~m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&~m[1562])|(~m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&m[1559]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[157])|((m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&m[1561]&m[1562]));
    m[1563] = (((m[1561]&~m[1564]&~m[1565]&~m[1566]&~m[1567])|(~m[1561]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1561]&m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1561]&~m[1564]&m[1565]&m[1566]&~m[1567])|(~m[1561]&m[1564]&~m[1565]&~m[1566]&m[1567])|(~m[1561]&~m[1564]&m[1565]&~m[1566]&m[1567])|(m[1561]&m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1561]&m[1564]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[158])|((m[1561]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(~m[1561]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1561]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1561]&m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1561]&~m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1561]&~m[1564]&~m[1565]&m[1566]&m[1567])|(m[1561]&~m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1561]&m[1564]&~m[1565]&m[1566]&m[1567])|(m[1561]&m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1561]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1561]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1561]&m[1564]&m[1565]&m[1566]&m[1567]));
    m[1568] = (((m[1566]&~m[1569]&~m[1570]&~m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&~m[1572])|(~m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&m[1569]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[159])|((m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&m[1571]&m[1572]));
    m[1573] = (((m[1571]&~m[1574]&~m[1575]&~m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&~m[1577])|(~m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&m[1574]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[160])|((m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&m[1576]&m[1577]));
    m[1578] = (((m[1576]&~m[1579]&~m[1580]&~m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&~m[1582])|(~m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&m[1579]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[161])|((m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&m[1581]&m[1582]));
    m[1583] = (((m[1581]&~m[1584]&~m[1585]&~m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&~m[1587])|(~m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&m[1584]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[162])|((m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&m[1586]&m[1587]));
    m[1588] = (((m[1586]&~m[1589]&~m[1590]&~m[1591]&~m[1592])|(~m[1586]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1586]&m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1586]&~m[1589]&m[1590]&m[1591]&~m[1592])|(~m[1586]&m[1589]&~m[1590]&~m[1591]&m[1592])|(~m[1586]&~m[1589]&m[1590]&~m[1591]&m[1592])|(m[1586]&m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1586]&m[1589]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[163])|((m[1586]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(~m[1586]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1586]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1586]&m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1586]&~m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1586]&~m[1589]&~m[1590]&m[1591]&m[1592])|(m[1586]&~m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1586]&m[1589]&~m[1590]&m[1591]&m[1592])|(m[1586]&m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1586]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1586]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1586]&m[1589]&m[1590]&m[1591]&m[1592]));
    m[1593] = (((m[1591]&~m[1594]&~m[1595]&~m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&~m[1597])|(~m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&m[1594]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[164])|((m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&m[1596]&m[1597]));
    m[1598] = (((m[1596]&~m[1599]&~m[1600]&~m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&~m[1602])|(~m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&m[1599]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[165])|((m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&m[1601]&m[1602]));
    m[1603] = (((m[1532]&~m[1604]&~m[1605]&~m[1606]&~m[1607])|(~m[1532]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1532]&m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1532]&~m[1604]&m[1605]&m[1606]&~m[1607])|(~m[1532]&m[1604]&~m[1605]&~m[1606]&m[1607])|(~m[1532]&~m[1604]&m[1605]&~m[1606]&m[1607])|(m[1532]&m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1532]&m[1604]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[166])|((m[1532]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(~m[1532]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1532]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1532]&m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1532]&~m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1532]&~m[1604]&~m[1605]&m[1606]&m[1607])|(m[1532]&~m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1532]&m[1604]&~m[1605]&m[1606]&m[1607])|(m[1532]&m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1532]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1532]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1532]&m[1604]&m[1605]&m[1606]&m[1607]));
    m[1608] = (((m[1606]&~m[1609]&~m[1610]&~m[1611]&~m[1612])|(~m[1606]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1606]&m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1606]&~m[1609]&m[1610]&m[1611]&~m[1612])|(~m[1606]&m[1609]&~m[1610]&~m[1611]&m[1612])|(~m[1606]&~m[1609]&m[1610]&~m[1611]&m[1612])|(m[1606]&m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1606]&m[1609]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[167])|((m[1606]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(~m[1606]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1606]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1606]&m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1606]&~m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1606]&~m[1609]&~m[1610]&m[1611]&m[1612])|(m[1606]&~m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1606]&m[1609]&~m[1610]&m[1611]&m[1612])|(m[1606]&m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1606]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1606]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1606]&m[1609]&m[1610]&m[1611]&m[1612]));
    m[1613] = (((m[1611]&~m[1614]&~m[1615]&~m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&~m[1617])|(~m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&m[1614]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[168])|((m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&m[1616]&m[1617]));
    m[1618] = (((m[1616]&~m[1619]&~m[1620]&~m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&~m[1622])|(~m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&m[1619]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[169])|((m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&m[1621]&m[1622]));
    m[1623] = (((m[1621]&~m[1624]&~m[1625]&~m[1626]&~m[1627])|(~m[1621]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1621]&m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1621]&~m[1624]&m[1625]&m[1626]&~m[1627])|(~m[1621]&m[1624]&~m[1625]&~m[1626]&m[1627])|(~m[1621]&~m[1624]&m[1625]&~m[1626]&m[1627])|(m[1621]&m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1621]&m[1624]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[170])|((m[1621]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(~m[1621]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1621]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1621]&m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1621]&~m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1621]&~m[1624]&~m[1625]&m[1626]&m[1627])|(m[1621]&~m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1621]&m[1624]&~m[1625]&m[1626]&m[1627])|(m[1621]&m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1621]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1621]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1621]&m[1624]&m[1625]&m[1626]&m[1627]));
    m[1628] = (((m[1626]&~m[1629]&~m[1630]&~m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&~m[1632])|(~m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&m[1629]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[171])|((m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&m[1631]&m[1632]));
    m[1633] = (((m[1631]&~m[1634]&~m[1635]&~m[1636]&~m[1637])|(~m[1631]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1631]&m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1631]&~m[1634]&m[1635]&m[1636]&~m[1637])|(~m[1631]&m[1634]&~m[1635]&~m[1636]&m[1637])|(~m[1631]&~m[1634]&m[1635]&~m[1636]&m[1637])|(m[1631]&m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1631]&m[1634]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[172])|((m[1631]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(~m[1631]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1631]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1631]&m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1631]&~m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1631]&~m[1634]&~m[1635]&m[1636]&m[1637])|(m[1631]&~m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1631]&m[1634]&~m[1635]&m[1636]&m[1637])|(m[1631]&m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1631]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1631]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1631]&m[1634]&m[1635]&m[1636]&m[1637]));
    m[1638] = (((m[1636]&~m[1639]&~m[1640]&~m[1641]&~m[1642])|(~m[1636]&~m[1639]&~m[1640]&m[1641]&~m[1642])|(m[1636]&m[1639]&~m[1640]&m[1641]&~m[1642])|(m[1636]&~m[1639]&m[1640]&m[1641]&~m[1642])|(~m[1636]&m[1639]&~m[1640]&~m[1641]&m[1642])|(~m[1636]&~m[1639]&m[1640]&~m[1641]&m[1642])|(m[1636]&m[1639]&m[1640]&~m[1641]&m[1642])|(~m[1636]&m[1639]&m[1640]&m[1641]&m[1642]))&UnbiasedRNG[173])|((m[1636]&~m[1639]&~m[1640]&m[1641]&~m[1642])|(~m[1636]&~m[1639]&~m[1640]&~m[1641]&m[1642])|(m[1636]&~m[1639]&~m[1640]&~m[1641]&m[1642])|(m[1636]&m[1639]&~m[1640]&~m[1641]&m[1642])|(m[1636]&~m[1639]&m[1640]&~m[1641]&m[1642])|(~m[1636]&~m[1639]&~m[1640]&m[1641]&m[1642])|(m[1636]&~m[1639]&~m[1640]&m[1641]&m[1642])|(~m[1636]&m[1639]&~m[1640]&m[1641]&m[1642])|(m[1636]&m[1639]&~m[1640]&m[1641]&m[1642])|(~m[1636]&~m[1639]&m[1640]&m[1641]&m[1642])|(m[1636]&~m[1639]&m[1640]&m[1641]&m[1642])|(m[1636]&m[1639]&m[1640]&m[1641]&m[1642]));
    m[1643] = (((m[1641]&~m[1644]&~m[1645]&~m[1646]&~m[1647])|(~m[1641]&~m[1644]&~m[1645]&m[1646]&~m[1647])|(m[1641]&m[1644]&~m[1645]&m[1646]&~m[1647])|(m[1641]&~m[1644]&m[1645]&m[1646]&~m[1647])|(~m[1641]&m[1644]&~m[1645]&~m[1646]&m[1647])|(~m[1641]&~m[1644]&m[1645]&~m[1646]&m[1647])|(m[1641]&m[1644]&m[1645]&~m[1646]&m[1647])|(~m[1641]&m[1644]&m[1645]&m[1646]&m[1647]))&UnbiasedRNG[174])|((m[1641]&~m[1644]&~m[1645]&m[1646]&~m[1647])|(~m[1641]&~m[1644]&~m[1645]&~m[1646]&m[1647])|(m[1641]&~m[1644]&~m[1645]&~m[1646]&m[1647])|(m[1641]&m[1644]&~m[1645]&~m[1646]&m[1647])|(m[1641]&~m[1644]&m[1645]&~m[1646]&m[1647])|(~m[1641]&~m[1644]&~m[1645]&m[1646]&m[1647])|(m[1641]&~m[1644]&~m[1645]&m[1646]&m[1647])|(~m[1641]&m[1644]&~m[1645]&m[1646]&m[1647])|(m[1641]&m[1644]&~m[1645]&m[1646]&m[1647])|(~m[1641]&~m[1644]&m[1645]&m[1646]&m[1647])|(m[1641]&~m[1644]&m[1645]&m[1646]&m[1647])|(m[1641]&m[1644]&m[1645]&m[1646]&m[1647]));
    m[1648] = (((m[1646]&~m[1649]&~m[1650]&~m[1651]&~m[1652])|(~m[1646]&~m[1649]&~m[1650]&m[1651]&~m[1652])|(m[1646]&m[1649]&~m[1650]&m[1651]&~m[1652])|(m[1646]&~m[1649]&m[1650]&m[1651]&~m[1652])|(~m[1646]&m[1649]&~m[1650]&~m[1651]&m[1652])|(~m[1646]&~m[1649]&m[1650]&~m[1651]&m[1652])|(m[1646]&m[1649]&m[1650]&~m[1651]&m[1652])|(~m[1646]&m[1649]&m[1650]&m[1651]&m[1652]))&UnbiasedRNG[175])|((m[1646]&~m[1649]&~m[1650]&m[1651]&~m[1652])|(~m[1646]&~m[1649]&~m[1650]&~m[1651]&m[1652])|(m[1646]&~m[1649]&~m[1650]&~m[1651]&m[1652])|(m[1646]&m[1649]&~m[1650]&~m[1651]&m[1652])|(m[1646]&~m[1649]&m[1650]&~m[1651]&m[1652])|(~m[1646]&~m[1649]&~m[1650]&m[1651]&m[1652])|(m[1646]&~m[1649]&~m[1650]&m[1651]&m[1652])|(~m[1646]&m[1649]&~m[1650]&m[1651]&m[1652])|(m[1646]&m[1649]&~m[1650]&m[1651]&m[1652])|(~m[1646]&~m[1649]&m[1650]&m[1651]&m[1652])|(m[1646]&~m[1649]&m[1650]&m[1651]&m[1652])|(m[1646]&m[1649]&m[1650]&m[1651]&m[1652]));
    m[1653] = (((m[1651]&~m[1654]&~m[1655]&~m[1656]&~m[1657])|(~m[1651]&~m[1654]&~m[1655]&m[1656]&~m[1657])|(m[1651]&m[1654]&~m[1655]&m[1656]&~m[1657])|(m[1651]&~m[1654]&m[1655]&m[1656]&~m[1657])|(~m[1651]&m[1654]&~m[1655]&~m[1656]&m[1657])|(~m[1651]&~m[1654]&m[1655]&~m[1656]&m[1657])|(m[1651]&m[1654]&m[1655]&~m[1656]&m[1657])|(~m[1651]&m[1654]&m[1655]&m[1656]&m[1657]))&UnbiasedRNG[176])|((m[1651]&~m[1654]&~m[1655]&m[1656]&~m[1657])|(~m[1651]&~m[1654]&~m[1655]&~m[1656]&m[1657])|(m[1651]&~m[1654]&~m[1655]&~m[1656]&m[1657])|(m[1651]&m[1654]&~m[1655]&~m[1656]&m[1657])|(m[1651]&~m[1654]&m[1655]&~m[1656]&m[1657])|(~m[1651]&~m[1654]&~m[1655]&m[1656]&m[1657])|(m[1651]&~m[1654]&~m[1655]&m[1656]&m[1657])|(~m[1651]&m[1654]&~m[1655]&m[1656]&m[1657])|(m[1651]&m[1654]&~m[1655]&m[1656]&m[1657])|(~m[1651]&~m[1654]&m[1655]&m[1656]&m[1657])|(m[1651]&~m[1654]&m[1655]&m[1656]&m[1657])|(m[1651]&m[1654]&m[1655]&m[1656]&m[1657]));
    m[1658] = (((m[1656]&~m[1659]&~m[1660]&~m[1661]&~m[1662])|(~m[1656]&~m[1659]&~m[1660]&m[1661]&~m[1662])|(m[1656]&m[1659]&~m[1660]&m[1661]&~m[1662])|(m[1656]&~m[1659]&m[1660]&m[1661]&~m[1662])|(~m[1656]&m[1659]&~m[1660]&~m[1661]&m[1662])|(~m[1656]&~m[1659]&m[1660]&~m[1661]&m[1662])|(m[1656]&m[1659]&m[1660]&~m[1661]&m[1662])|(~m[1656]&m[1659]&m[1660]&m[1661]&m[1662]))&UnbiasedRNG[177])|((m[1656]&~m[1659]&~m[1660]&m[1661]&~m[1662])|(~m[1656]&~m[1659]&~m[1660]&~m[1661]&m[1662])|(m[1656]&~m[1659]&~m[1660]&~m[1661]&m[1662])|(m[1656]&m[1659]&~m[1660]&~m[1661]&m[1662])|(m[1656]&~m[1659]&m[1660]&~m[1661]&m[1662])|(~m[1656]&~m[1659]&~m[1660]&m[1661]&m[1662])|(m[1656]&~m[1659]&~m[1660]&m[1661]&m[1662])|(~m[1656]&m[1659]&~m[1660]&m[1661]&m[1662])|(m[1656]&m[1659]&~m[1660]&m[1661]&m[1662])|(~m[1656]&~m[1659]&m[1660]&m[1661]&m[1662])|(m[1656]&~m[1659]&m[1660]&m[1661]&m[1662])|(m[1656]&m[1659]&m[1660]&m[1661]&m[1662]));
    m[1663] = (((m[1661]&~m[1664]&~m[1665]&~m[1666]&~m[1667])|(~m[1661]&~m[1664]&~m[1665]&m[1666]&~m[1667])|(m[1661]&m[1664]&~m[1665]&m[1666]&~m[1667])|(m[1661]&~m[1664]&m[1665]&m[1666]&~m[1667])|(~m[1661]&m[1664]&~m[1665]&~m[1666]&m[1667])|(~m[1661]&~m[1664]&m[1665]&~m[1666]&m[1667])|(m[1661]&m[1664]&m[1665]&~m[1666]&m[1667])|(~m[1661]&m[1664]&m[1665]&m[1666]&m[1667]))&UnbiasedRNG[178])|((m[1661]&~m[1664]&~m[1665]&m[1666]&~m[1667])|(~m[1661]&~m[1664]&~m[1665]&~m[1666]&m[1667])|(m[1661]&~m[1664]&~m[1665]&~m[1666]&m[1667])|(m[1661]&m[1664]&~m[1665]&~m[1666]&m[1667])|(m[1661]&~m[1664]&m[1665]&~m[1666]&m[1667])|(~m[1661]&~m[1664]&~m[1665]&m[1666]&m[1667])|(m[1661]&~m[1664]&~m[1665]&m[1666]&m[1667])|(~m[1661]&m[1664]&~m[1665]&m[1666]&m[1667])|(m[1661]&m[1664]&~m[1665]&m[1666]&m[1667])|(~m[1661]&~m[1664]&m[1665]&m[1666]&m[1667])|(m[1661]&~m[1664]&m[1665]&m[1666]&m[1667])|(m[1661]&m[1664]&m[1665]&m[1666]&m[1667]));
    m[1668] = (((m[1666]&~m[1669]&~m[1670]&~m[1671]&~m[1672])|(~m[1666]&~m[1669]&~m[1670]&m[1671]&~m[1672])|(m[1666]&m[1669]&~m[1670]&m[1671]&~m[1672])|(m[1666]&~m[1669]&m[1670]&m[1671]&~m[1672])|(~m[1666]&m[1669]&~m[1670]&~m[1671]&m[1672])|(~m[1666]&~m[1669]&m[1670]&~m[1671]&m[1672])|(m[1666]&m[1669]&m[1670]&~m[1671]&m[1672])|(~m[1666]&m[1669]&m[1670]&m[1671]&m[1672]))&UnbiasedRNG[179])|((m[1666]&~m[1669]&~m[1670]&m[1671]&~m[1672])|(~m[1666]&~m[1669]&~m[1670]&~m[1671]&m[1672])|(m[1666]&~m[1669]&~m[1670]&~m[1671]&m[1672])|(m[1666]&m[1669]&~m[1670]&~m[1671]&m[1672])|(m[1666]&~m[1669]&m[1670]&~m[1671]&m[1672])|(~m[1666]&~m[1669]&~m[1670]&m[1671]&m[1672])|(m[1666]&~m[1669]&~m[1670]&m[1671]&m[1672])|(~m[1666]&m[1669]&~m[1670]&m[1671]&m[1672])|(m[1666]&m[1669]&~m[1670]&m[1671]&m[1672])|(~m[1666]&~m[1669]&m[1670]&m[1671]&m[1672])|(m[1666]&~m[1669]&m[1670]&m[1671]&m[1672])|(m[1666]&m[1669]&m[1670]&m[1671]&m[1672]));
    m[1673] = (((m[1607]&~m[1674]&~m[1675]&~m[1676]&~m[1677])|(~m[1607]&~m[1674]&~m[1675]&m[1676]&~m[1677])|(m[1607]&m[1674]&~m[1675]&m[1676]&~m[1677])|(m[1607]&~m[1674]&m[1675]&m[1676]&~m[1677])|(~m[1607]&m[1674]&~m[1675]&~m[1676]&m[1677])|(~m[1607]&~m[1674]&m[1675]&~m[1676]&m[1677])|(m[1607]&m[1674]&m[1675]&~m[1676]&m[1677])|(~m[1607]&m[1674]&m[1675]&m[1676]&m[1677]))&UnbiasedRNG[180])|((m[1607]&~m[1674]&~m[1675]&m[1676]&~m[1677])|(~m[1607]&~m[1674]&~m[1675]&~m[1676]&m[1677])|(m[1607]&~m[1674]&~m[1675]&~m[1676]&m[1677])|(m[1607]&m[1674]&~m[1675]&~m[1676]&m[1677])|(m[1607]&~m[1674]&m[1675]&~m[1676]&m[1677])|(~m[1607]&~m[1674]&~m[1675]&m[1676]&m[1677])|(m[1607]&~m[1674]&~m[1675]&m[1676]&m[1677])|(~m[1607]&m[1674]&~m[1675]&m[1676]&m[1677])|(m[1607]&m[1674]&~m[1675]&m[1676]&m[1677])|(~m[1607]&~m[1674]&m[1675]&m[1676]&m[1677])|(m[1607]&~m[1674]&m[1675]&m[1676]&m[1677])|(m[1607]&m[1674]&m[1675]&m[1676]&m[1677]));
    m[1678] = (((m[1676]&~m[1679]&~m[1680]&~m[1681]&~m[1682])|(~m[1676]&~m[1679]&~m[1680]&m[1681]&~m[1682])|(m[1676]&m[1679]&~m[1680]&m[1681]&~m[1682])|(m[1676]&~m[1679]&m[1680]&m[1681]&~m[1682])|(~m[1676]&m[1679]&~m[1680]&~m[1681]&m[1682])|(~m[1676]&~m[1679]&m[1680]&~m[1681]&m[1682])|(m[1676]&m[1679]&m[1680]&~m[1681]&m[1682])|(~m[1676]&m[1679]&m[1680]&m[1681]&m[1682]))&UnbiasedRNG[181])|((m[1676]&~m[1679]&~m[1680]&m[1681]&~m[1682])|(~m[1676]&~m[1679]&~m[1680]&~m[1681]&m[1682])|(m[1676]&~m[1679]&~m[1680]&~m[1681]&m[1682])|(m[1676]&m[1679]&~m[1680]&~m[1681]&m[1682])|(m[1676]&~m[1679]&m[1680]&~m[1681]&m[1682])|(~m[1676]&~m[1679]&~m[1680]&m[1681]&m[1682])|(m[1676]&~m[1679]&~m[1680]&m[1681]&m[1682])|(~m[1676]&m[1679]&~m[1680]&m[1681]&m[1682])|(m[1676]&m[1679]&~m[1680]&m[1681]&m[1682])|(~m[1676]&~m[1679]&m[1680]&m[1681]&m[1682])|(m[1676]&~m[1679]&m[1680]&m[1681]&m[1682])|(m[1676]&m[1679]&m[1680]&m[1681]&m[1682]));
    m[1683] = (((m[1681]&~m[1684]&~m[1685]&~m[1686]&~m[1687])|(~m[1681]&~m[1684]&~m[1685]&m[1686]&~m[1687])|(m[1681]&m[1684]&~m[1685]&m[1686]&~m[1687])|(m[1681]&~m[1684]&m[1685]&m[1686]&~m[1687])|(~m[1681]&m[1684]&~m[1685]&~m[1686]&m[1687])|(~m[1681]&~m[1684]&m[1685]&~m[1686]&m[1687])|(m[1681]&m[1684]&m[1685]&~m[1686]&m[1687])|(~m[1681]&m[1684]&m[1685]&m[1686]&m[1687]))&UnbiasedRNG[182])|((m[1681]&~m[1684]&~m[1685]&m[1686]&~m[1687])|(~m[1681]&~m[1684]&~m[1685]&~m[1686]&m[1687])|(m[1681]&~m[1684]&~m[1685]&~m[1686]&m[1687])|(m[1681]&m[1684]&~m[1685]&~m[1686]&m[1687])|(m[1681]&~m[1684]&m[1685]&~m[1686]&m[1687])|(~m[1681]&~m[1684]&~m[1685]&m[1686]&m[1687])|(m[1681]&~m[1684]&~m[1685]&m[1686]&m[1687])|(~m[1681]&m[1684]&~m[1685]&m[1686]&m[1687])|(m[1681]&m[1684]&~m[1685]&m[1686]&m[1687])|(~m[1681]&~m[1684]&m[1685]&m[1686]&m[1687])|(m[1681]&~m[1684]&m[1685]&m[1686]&m[1687])|(m[1681]&m[1684]&m[1685]&m[1686]&m[1687]));
    m[1688] = (((m[1686]&~m[1689]&~m[1690]&~m[1691]&~m[1692])|(~m[1686]&~m[1689]&~m[1690]&m[1691]&~m[1692])|(m[1686]&m[1689]&~m[1690]&m[1691]&~m[1692])|(m[1686]&~m[1689]&m[1690]&m[1691]&~m[1692])|(~m[1686]&m[1689]&~m[1690]&~m[1691]&m[1692])|(~m[1686]&~m[1689]&m[1690]&~m[1691]&m[1692])|(m[1686]&m[1689]&m[1690]&~m[1691]&m[1692])|(~m[1686]&m[1689]&m[1690]&m[1691]&m[1692]))&UnbiasedRNG[183])|((m[1686]&~m[1689]&~m[1690]&m[1691]&~m[1692])|(~m[1686]&~m[1689]&~m[1690]&~m[1691]&m[1692])|(m[1686]&~m[1689]&~m[1690]&~m[1691]&m[1692])|(m[1686]&m[1689]&~m[1690]&~m[1691]&m[1692])|(m[1686]&~m[1689]&m[1690]&~m[1691]&m[1692])|(~m[1686]&~m[1689]&~m[1690]&m[1691]&m[1692])|(m[1686]&~m[1689]&~m[1690]&m[1691]&m[1692])|(~m[1686]&m[1689]&~m[1690]&m[1691]&m[1692])|(m[1686]&m[1689]&~m[1690]&m[1691]&m[1692])|(~m[1686]&~m[1689]&m[1690]&m[1691]&m[1692])|(m[1686]&~m[1689]&m[1690]&m[1691]&m[1692])|(m[1686]&m[1689]&m[1690]&m[1691]&m[1692]));
    m[1693] = (((m[1691]&~m[1694]&~m[1695]&~m[1696]&~m[1697])|(~m[1691]&~m[1694]&~m[1695]&m[1696]&~m[1697])|(m[1691]&m[1694]&~m[1695]&m[1696]&~m[1697])|(m[1691]&~m[1694]&m[1695]&m[1696]&~m[1697])|(~m[1691]&m[1694]&~m[1695]&~m[1696]&m[1697])|(~m[1691]&~m[1694]&m[1695]&~m[1696]&m[1697])|(m[1691]&m[1694]&m[1695]&~m[1696]&m[1697])|(~m[1691]&m[1694]&m[1695]&m[1696]&m[1697]))&UnbiasedRNG[184])|((m[1691]&~m[1694]&~m[1695]&m[1696]&~m[1697])|(~m[1691]&~m[1694]&~m[1695]&~m[1696]&m[1697])|(m[1691]&~m[1694]&~m[1695]&~m[1696]&m[1697])|(m[1691]&m[1694]&~m[1695]&~m[1696]&m[1697])|(m[1691]&~m[1694]&m[1695]&~m[1696]&m[1697])|(~m[1691]&~m[1694]&~m[1695]&m[1696]&m[1697])|(m[1691]&~m[1694]&~m[1695]&m[1696]&m[1697])|(~m[1691]&m[1694]&~m[1695]&m[1696]&m[1697])|(m[1691]&m[1694]&~m[1695]&m[1696]&m[1697])|(~m[1691]&~m[1694]&m[1695]&m[1696]&m[1697])|(m[1691]&~m[1694]&m[1695]&m[1696]&m[1697])|(m[1691]&m[1694]&m[1695]&m[1696]&m[1697]));
    m[1698] = (((m[1696]&~m[1699]&~m[1700]&~m[1701]&~m[1702])|(~m[1696]&~m[1699]&~m[1700]&m[1701]&~m[1702])|(m[1696]&m[1699]&~m[1700]&m[1701]&~m[1702])|(m[1696]&~m[1699]&m[1700]&m[1701]&~m[1702])|(~m[1696]&m[1699]&~m[1700]&~m[1701]&m[1702])|(~m[1696]&~m[1699]&m[1700]&~m[1701]&m[1702])|(m[1696]&m[1699]&m[1700]&~m[1701]&m[1702])|(~m[1696]&m[1699]&m[1700]&m[1701]&m[1702]))&UnbiasedRNG[185])|((m[1696]&~m[1699]&~m[1700]&m[1701]&~m[1702])|(~m[1696]&~m[1699]&~m[1700]&~m[1701]&m[1702])|(m[1696]&~m[1699]&~m[1700]&~m[1701]&m[1702])|(m[1696]&m[1699]&~m[1700]&~m[1701]&m[1702])|(m[1696]&~m[1699]&m[1700]&~m[1701]&m[1702])|(~m[1696]&~m[1699]&~m[1700]&m[1701]&m[1702])|(m[1696]&~m[1699]&~m[1700]&m[1701]&m[1702])|(~m[1696]&m[1699]&~m[1700]&m[1701]&m[1702])|(m[1696]&m[1699]&~m[1700]&m[1701]&m[1702])|(~m[1696]&~m[1699]&m[1700]&m[1701]&m[1702])|(m[1696]&~m[1699]&m[1700]&m[1701]&m[1702])|(m[1696]&m[1699]&m[1700]&m[1701]&m[1702]));
    m[1703] = (((m[1701]&~m[1704]&~m[1705]&~m[1706]&~m[1707])|(~m[1701]&~m[1704]&~m[1705]&m[1706]&~m[1707])|(m[1701]&m[1704]&~m[1705]&m[1706]&~m[1707])|(m[1701]&~m[1704]&m[1705]&m[1706]&~m[1707])|(~m[1701]&m[1704]&~m[1705]&~m[1706]&m[1707])|(~m[1701]&~m[1704]&m[1705]&~m[1706]&m[1707])|(m[1701]&m[1704]&m[1705]&~m[1706]&m[1707])|(~m[1701]&m[1704]&m[1705]&m[1706]&m[1707]))&UnbiasedRNG[186])|((m[1701]&~m[1704]&~m[1705]&m[1706]&~m[1707])|(~m[1701]&~m[1704]&~m[1705]&~m[1706]&m[1707])|(m[1701]&~m[1704]&~m[1705]&~m[1706]&m[1707])|(m[1701]&m[1704]&~m[1705]&~m[1706]&m[1707])|(m[1701]&~m[1704]&m[1705]&~m[1706]&m[1707])|(~m[1701]&~m[1704]&~m[1705]&m[1706]&m[1707])|(m[1701]&~m[1704]&~m[1705]&m[1706]&m[1707])|(~m[1701]&m[1704]&~m[1705]&m[1706]&m[1707])|(m[1701]&m[1704]&~m[1705]&m[1706]&m[1707])|(~m[1701]&~m[1704]&m[1705]&m[1706]&m[1707])|(m[1701]&~m[1704]&m[1705]&m[1706]&m[1707])|(m[1701]&m[1704]&m[1705]&m[1706]&m[1707]));
    m[1708] = (((m[1706]&~m[1709]&~m[1710]&~m[1711]&~m[1712])|(~m[1706]&~m[1709]&~m[1710]&m[1711]&~m[1712])|(m[1706]&m[1709]&~m[1710]&m[1711]&~m[1712])|(m[1706]&~m[1709]&m[1710]&m[1711]&~m[1712])|(~m[1706]&m[1709]&~m[1710]&~m[1711]&m[1712])|(~m[1706]&~m[1709]&m[1710]&~m[1711]&m[1712])|(m[1706]&m[1709]&m[1710]&~m[1711]&m[1712])|(~m[1706]&m[1709]&m[1710]&m[1711]&m[1712]))&UnbiasedRNG[187])|((m[1706]&~m[1709]&~m[1710]&m[1711]&~m[1712])|(~m[1706]&~m[1709]&~m[1710]&~m[1711]&m[1712])|(m[1706]&~m[1709]&~m[1710]&~m[1711]&m[1712])|(m[1706]&m[1709]&~m[1710]&~m[1711]&m[1712])|(m[1706]&~m[1709]&m[1710]&~m[1711]&m[1712])|(~m[1706]&~m[1709]&~m[1710]&m[1711]&m[1712])|(m[1706]&~m[1709]&~m[1710]&m[1711]&m[1712])|(~m[1706]&m[1709]&~m[1710]&m[1711]&m[1712])|(m[1706]&m[1709]&~m[1710]&m[1711]&m[1712])|(~m[1706]&~m[1709]&m[1710]&m[1711]&m[1712])|(m[1706]&~m[1709]&m[1710]&m[1711]&m[1712])|(m[1706]&m[1709]&m[1710]&m[1711]&m[1712]));
    m[1713] = (((m[1711]&~m[1714]&~m[1715]&~m[1716]&~m[1717])|(~m[1711]&~m[1714]&~m[1715]&m[1716]&~m[1717])|(m[1711]&m[1714]&~m[1715]&m[1716]&~m[1717])|(m[1711]&~m[1714]&m[1715]&m[1716]&~m[1717])|(~m[1711]&m[1714]&~m[1715]&~m[1716]&m[1717])|(~m[1711]&~m[1714]&m[1715]&~m[1716]&m[1717])|(m[1711]&m[1714]&m[1715]&~m[1716]&m[1717])|(~m[1711]&m[1714]&m[1715]&m[1716]&m[1717]))&UnbiasedRNG[188])|((m[1711]&~m[1714]&~m[1715]&m[1716]&~m[1717])|(~m[1711]&~m[1714]&~m[1715]&~m[1716]&m[1717])|(m[1711]&~m[1714]&~m[1715]&~m[1716]&m[1717])|(m[1711]&m[1714]&~m[1715]&~m[1716]&m[1717])|(m[1711]&~m[1714]&m[1715]&~m[1716]&m[1717])|(~m[1711]&~m[1714]&~m[1715]&m[1716]&m[1717])|(m[1711]&~m[1714]&~m[1715]&m[1716]&m[1717])|(~m[1711]&m[1714]&~m[1715]&m[1716]&m[1717])|(m[1711]&m[1714]&~m[1715]&m[1716]&m[1717])|(~m[1711]&~m[1714]&m[1715]&m[1716]&m[1717])|(m[1711]&~m[1714]&m[1715]&m[1716]&m[1717])|(m[1711]&m[1714]&m[1715]&m[1716]&m[1717]));
    m[1718] = (((m[1716]&~m[1719]&~m[1720]&~m[1721]&~m[1722])|(~m[1716]&~m[1719]&~m[1720]&m[1721]&~m[1722])|(m[1716]&m[1719]&~m[1720]&m[1721]&~m[1722])|(m[1716]&~m[1719]&m[1720]&m[1721]&~m[1722])|(~m[1716]&m[1719]&~m[1720]&~m[1721]&m[1722])|(~m[1716]&~m[1719]&m[1720]&~m[1721]&m[1722])|(m[1716]&m[1719]&m[1720]&~m[1721]&m[1722])|(~m[1716]&m[1719]&m[1720]&m[1721]&m[1722]))&UnbiasedRNG[189])|((m[1716]&~m[1719]&~m[1720]&m[1721]&~m[1722])|(~m[1716]&~m[1719]&~m[1720]&~m[1721]&m[1722])|(m[1716]&~m[1719]&~m[1720]&~m[1721]&m[1722])|(m[1716]&m[1719]&~m[1720]&~m[1721]&m[1722])|(m[1716]&~m[1719]&m[1720]&~m[1721]&m[1722])|(~m[1716]&~m[1719]&~m[1720]&m[1721]&m[1722])|(m[1716]&~m[1719]&~m[1720]&m[1721]&m[1722])|(~m[1716]&m[1719]&~m[1720]&m[1721]&m[1722])|(m[1716]&m[1719]&~m[1720]&m[1721]&m[1722])|(~m[1716]&~m[1719]&m[1720]&m[1721]&m[1722])|(m[1716]&~m[1719]&m[1720]&m[1721]&m[1722])|(m[1716]&m[1719]&m[1720]&m[1721]&m[1722]));
    m[1723] = (((m[1721]&~m[1724]&~m[1725]&~m[1726]&~m[1727])|(~m[1721]&~m[1724]&~m[1725]&m[1726]&~m[1727])|(m[1721]&m[1724]&~m[1725]&m[1726]&~m[1727])|(m[1721]&~m[1724]&m[1725]&m[1726]&~m[1727])|(~m[1721]&m[1724]&~m[1725]&~m[1726]&m[1727])|(~m[1721]&~m[1724]&m[1725]&~m[1726]&m[1727])|(m[1721]&m[1724]&m[1725]&~m[1726]&m[1727])|(~m[1721]&m[1724]&m[1725]&m[1726]&m[1727]))&UnbiasedRNG[190])|((m[1721]&~m[1724]&~m[1725]&m[1726]&~m[1727])|(~m[1721]&~m[1724]&~m[1725]&~m[1726]&m[1727])|(m[1721]&~m[1724]&~m[1725]&~m[1726]&m[1727])|(m[1721]&m[1724]&~m[1725]&~m[1726]&m[1727])|(m[1721]&~m[1724]&m[1725]&~m[1726]&m[1727])|(~m[1721]&~m[1724]&~m[1725]&m[1726]&m[1727])|(m[1721]&~m[1724]&~m[1725]&m[1726]&m[1727])|(~m[1721]&m[1724]&~m[1725]&m[1726]&m[1727])|(m[1721]&m[1724]&~m[1725]&m[1726]&m[1727])|(~m[1721]&~m[1724]&m[1725]&m[1726]&m[1727])|(m[1721]&~m[1724]&m[1725]&m[1726]&m[1727])|(m[1721]&m[1724]&m[1725]&m[1726]&m[1727]));
    m[1728] = (((m[1726]&~m[1729]&~m[1730]&~m[1731]&~m[1732])|(~m[1726]&~m[1729]&~m[1730]&m[1731]&~m[1732])|(m[1726]&m[1729]&~m[1730]&m[1731]&~m[1732])|(m[1726]&~m[1729]&m[1730]&m[1731]&~m[1732])|(~m[1726]&m[1729]&~m[1730]&~m[1731]&m[1732])|(~m[1726]&~m[1729]&m[1730]&~m[1731]&m[1732])|(m[1726]&m[1729]&m[1730]&~m[1731]&m[1732])|(~m[1726]&m[1729]&m[1730]&m[1731]&m[1732]))&UnbiasedRNG[191])|((m[1726]&~m[1729]&~m[1730]&m[1731]&~m[1732])|(~m[1726]&~m[1729]&~m[1730]&~m[1731]&m[1732])|(m[1726]&~m[1729]&~m[1730]&~m[1731]&m[1732])|(m[1726]&m[1729]&~m[1730]&~m[1731]&m[1732])|(m[1726]&~m[1729]&m[1730]&~m[1731]&m[1732])|(~m[1726]&~m[1729]&~m[1730]&m[1731]&m[1732])|(m[1726]&~m[1729]&~m[1730]&m[1731]&m[1732])|(~m[1726]&m[1729]&~m[1730]&m[1731]&m[1732])|(m[1726]&m[1729]&~m[1730]&m[1731]&m[1732])|(~m[1726]&~m[1729]&m[1730]&m[1731]&m[1732])|(m[1726]&~m[1729]&m[1730]&m[1731]&m[1732])|(m[1726]&m[1729]&m[1730]&m[1731]&m[1732]));
    m[1733] = (((m[1731]&~m[1734]&~m[1735]&~m[1736]&~m[1737])|(~m[1731]&~m[1734]&~m[1735]&m[1736]&~m[1737])|(m[1731]&m[1734]&~m[1735]&m[1736]&~m[1737])|(m[1731]&~m[1734]&m[1735]&m[1736]&~m[1737])|(~m[1731]&m[1734]&~m[1735]&~m[1736]&m[1737])|(~m[1731]&~m[1734]&m[1735]&~m[1736]&m[1737])|(m[1731]&m[1734]&m[1735]&~m[1736]&m[1737])|(~m[1731]&m[1734]&m[1735]&m[1736]&m[1737]))&UnbiasedRNG[192])|((m[1731]&~m[1734]&~m[1735]&m[1736]&~m[1737])|(~m[1731]&~m[1734]&~m[1735]&~m[1736]&m[1737])|(m[1731]&~m[1734]&~m[1735]&~m[1736]&m[1737])|(m[1731]&m[1734]&~m[1735]&~m[1736]&m[1737])|(m[1731]&~m[1734]&m[1735]&~m[1736]&m[1737])|(~m[1731]&~m[1734]&~m[1735]&m[1736]&m[1737])|(m[1731]&~m[1734]&~m[1735]&m[1736]&m[1737])|(~m[1731]&m[1734]&~m[1735]&m[1736]&m[1737])|(m[1731]&m[1734]&~m[1735]&m[1736]&m[1737])|(~m[1731]&~m[1734]&m[1735]&m[1736]&m[1737])|(m[1731]&~m[1734]&m[1735]&m[1736]&m[1737])|(m[1731]&m[1734]&m[1735]&m[1736]&m[1737]));
    m[1738] = (((m[1677]&~m[1739]&~m[1740]&~m[1741]&~m[1742])|(~m[1677]&~m[1739]&~m[1740]&m[1741]&~m[1742])|(m[1677]&m[1739]&~m[1740]&m[1741]&~m[1742])|(m[1677]&~m[1739]&m[1740]&m[1741]&~m[1742])|(~m[1677]&m[1739]&~m[1740]&~m[1741]&m[1742])|(~m[1677]&~m[1739]&m[1740]&~m[1741]&m[1742])|(m[1677]&m[1739]&m[1740]&~m[1741]&m[1742])|(~m[1677]&m[1739]&m[1740]&m[1741]&m[1742]))&UnbiasedRNG[193])|((m[1677]&~m[1739]&~m[1740]&m[1741]&~m[1742])|(~m[1677]&~m[1739]&~m[1740]&~m[1741]&m[1742])|(m[1677]&~m[1739]&~m[1740]&~m[1741]&m[1742])|(m[1677]&m[1739]&~m[1740]&~m[1741]&m[1742])|(m[1677]&~m[1739]&m[1740]&~m[1741]&m[1742])|(~m[1677]&~m[1739]&~m[1740]&m[1741]&m[1742])|(m[1677]&~m[1739]&~m[1740]&m[1741]&m[1742])|(~m[1677]&m[1739]&~m[1740]&m[1741]&m[1742])|(m[1677]&m[1739]&~m[1740]&m[1741]&m[1742])|(~m[1677]&~m[1739]&m[1740]&m[1741]&m[1742])|(m[1677]&~m[1739]&m[1740]&m[1741]&m[1742])|(m[1677]&m[1739]&m[1740]&m[1741]&m[1742]));
    m[1743] = (((m[1741]&~m[1744]&~m[1745]&~m[1746]&~m[1747])|(~m[1741]&~m[1744]&~m[1745]&m[1746]&~m[1747])|(m[1741]&m[1744]&~m[1745]&m[1746]&~m[1747])|(m[1741]&~m[1744]&m[1745]&m[1746]&~m[1747])|(~m[1741]&m[1744]&~m[1745]&~m[1746]&m[1747])|(~m[1741]&~m[1744]&m[1745]&~m[1746]&m[1747])|(m[1741]&m[1744]&m[1745]&~m[1746]&m[1747])|(~m[1741]&m[1744]&m[1745]&m[1746]&m[1747]))&UnbiasedRNG[194])|((m[1741]&~m[1744]&~m[1745]&m[1746]&~m[1747])|(~m[1741]&~m[1744]&~m[1745]&~m[1746]&m[1747])|(m[1741]&~m[1744]&~m[1745]&~m[1746]&m[1747])|(m[1741]&m[1744]&~m[1745]&~m[1746]&m[1747])|(m[1741]&~m[1744]&m[1745]&~m[1746]&m[1747])|(~m[1741]&~m[1744]&~m[1745]&m[1746]&m[1747])|(m[1741]&~m[1744]&~m[1745]&m[1746]&m[1747])|(~m[1741]&m[1744]&~m[1745]&m[1746]&m[1747])|(m[1741]&m[1744]&~m[1745]&m[1746]&m[1747])|(~m[1741]&~m[1744]&m[1745]&m[1746]&m[1747])|(m[1741]&~m[1744]&m[1745]&m[1746]&m[1747])|(m[1741]&m[1744]&m[1745]&m[1746]&m[1747]));
    m[1748] = (((m[1746]&~m[1749]&~m[1750]&~m[1751]&~m[1752])|(~m[1746]&~m[1749]&~m[1750]&m[1751]&~m[1752])|(m[1746]&m[1749]&~m[1750]&m[1751]&~m[1752])|(m[1746]&~m[1749]&m[1750]&m[1751]&~m[1752])|(~m[1746]&m[1749]&~m[1750]&~m[1751]&m[1752])|(~m[1746]&~m[1749]&m[1750]&~m[1751]&m[1752])|(m[1746]&m[1749]&m[1750]&~m[1751]&m[1752])|(~m[1746]&m[1749]&m[1750]&m[1751]&m[1752]))&UnbiasedRNG[195])|((m[1746]&~m[1749]&~m[1750]&m[1751]&~m[1752])|(~m[1746]&~m[1749]&~m[1750]&~m[1751]&m[1752])|(m[1746]&~m[1749]&~m[1750]&~m[1751]&m[1752])|(m[1746]&m[1749]&~m[1750]&~m[1751]&m[1752])|(m[1746]&~m[1749]&m[1750]&~m[1751]&m[1752])|(~m[1746]&~m[1749]&~m[1750]&m[1751]&m[1752])|(m[1746]&~m[1749]&~m[1750]&m[1751]&m[1752])|(~m[1746]&m[1749]&~m[1750]&m[1751]&m[1752])|(m[1746]&m[1749]&~m[1750]&m[1751]&m[1752])|(~m[1746]&~m[1749]&m[1750]&m[1751]&m[1752])|(m[1746]&~m[1749]&m[1750]&m[1751]&m[1752])|(m[1746]&m[1749]&m[1750]&m[1751]&m[1752]));
    m[1753] = (((m[1751]&~m[1754]&~m[1755]&~m[1756]&~m[1757])|(~m[1751]&~m[1754]&~m[1755]&m[1756]&~m[1757])|(m[1751]&m[1754]&~m[1755]&m[1756]&~m[1757])|(m[1751]&~m[1754]&m[1755]&m[1756]&~m[1757])|(~m[1751]&m[1754]&~m[1755]&~m[1756]&m[1757])|(~m[1751]&~m[1754]&m[1755]&~m[1756]&m[1757])|(m[1751]&m[1754]&m[1755]&~m[1756]&m[1757])|(~m[1751]&m[1754]&m[1755]&m[1756]&m[1757]))&UnbiasedRNG[196])|((m[1751]&~m[1754]&~m[1755]&m[1756]&~m[1757])|(~m[1751]&~m[1754]&~m[1755]&~m[1756]&m[1757])|(m[1751]&~m[1754]&~m[1755]&~m[1756]&m[1757])|(m[1751]&m[1754]&~m[1755]&~m[1756]&m[1757])|(m[1751]&~m[1754]&m[1755]&~m[1756]&m[1757])|(~m[1751]&~m[1754]&~m[1755]&m[1756]&m[1757])|(m[1751]&~m[1754]&~m[1755]&m[1756]&m[1757])|(~m[1751]&m[1754]&~m[1755]&m[1756]&m[1757])|(m[1751]&m[1754]&~m[1755]&m[1756]&m[1757])|(~m[1751]&~m[1754]&m[1755]&m[1756]&m[1757])|(m[1751]&~m[1754]&m[1755]&m[1756]&m[1757])|(m[1751]&m[1754]&m[1755]&m[1756]&m[1757]));
    m[1758] = (((m[1756]&~m[1759]&~m[1760]&~m[1761]&~m[1762])|(~m[1756]&~m[1759]&~m[1760]&m[1761]&~m[1762])|(m[1756]&m[1759]&~m[1760]&m[1761]&~m[1762])|(m[1756]&~m[1759]&m[1760]&m[1761]&~m[1762])|(~m[1756]&m[1759]&~m[1760]&~m[1761]&m[1762])|(~m[1756]&~m[1759]&m[1760]&~m[1761]&m[1762])|(m[1756]&m[1759]&m[1760]&~m[1761]&m[1762])|(~m[1756]&m[1759]&m[1760]&m[1761]&m[1762]))&UnbiasedRNG[197])|((m[1756]&~m[1759]&~m[1760]&m[1761]&~m[1762])|(~m[1756]&~m[1759]&~m[1760]&~m[1761]&m[1762])|(m[1756]&~m[1759]&~m[1760]&~m[1761]&m[1762])|(m[1756]&m[1759]&~m[1760]&~m[1761]&m[1762])|(m[1756]&~m[1759]&m[1760]&~m[1761]&m[1762])|(~m[1756]&~m[1759]&~m[1760]&m[1761]&m[1762])|(m[1756]&~m[1759]&~m[1760]&m[1761]&m[1762])|(~m[1756]&m[1759]&~m[1760]&m[1761]&m[1762])|(m[1756]&m[1759]&~m[1760]&m[1761]&m[1762])|(~m[1756]&~m[1759]&m[1760]&m[1761]&m[1762])|(m[1756]&~m[1759]&m[1760]&m[1761]&m[1762])|(m[1756]&m[1759]&m[1760]&m[1761]&m[1762]));
    m[1763] = (((m[1761]&~m[1764]&~m[1765]&~m[1766]&~m[1767])|(~m[1761]&~m[1764]&~m[1765]&m[1766]&~m[1767])|(m[1761]&m[1764]&~m[1765]&m[1766]&~m[1767])|(m[1761]&~m[1764]&m[1765]&m[1766]&~m[1767])|(~m[1761]&m[1764]&~m[1765]&~m[1766]&m[1767])|(~m[1761]&~m[1764]&m[1765]&~m[1766]&m[1767])|(m[1761]&m[1764]&m[1765]&~m[1766]&m[1767])|(~m[1761]&m[1764]&m[1765]&m[1766]&m[1767]))&UnbiasedRNG[198])|((m[1761]&~m[1764]&~m[1765]&m[1766]&~m[1767])|(~m[1761]&~m[1764]&~m[1765]&~m[1766]&m[1767])|(m[1761]&~m[1764]&~m[1765]&~m[1766]&m[1767])|(m[1761]&m[1764]&~m[1765]&~m[1766]&m[1767])|(m[1761]&~m[1764]&m[1765]&~m[1766]&m[1767])|(~m[1761]&~m[1764]&~m[1765]&m[1766]&m[1767])|(m[1761]&~m[1764]&~m[1765]&m[1766]&m[1767])|(~m[1761]&m[1764]&~m[1765]&m[1766]&m[1767])|(m[1761]&m[1764]&~m[1765]&m[1766]&m[1767])|(~m[1761]&~m[1764]&m[1765]&m[1766]&m[1767])|(m[1761]&~m[1764]&m[1765]&m[1766]&m[1767])|(m[1761]&m[1764]&m[1765]&m[1766]&m[1767]));
    m[1768] = (((m[1766]&~m[1769]&~m[1770]&~m[1771]&~m[1772])|(~m[1766]&~m[1769]&~m[1770]&m[1771]&~m[1772])|(m[1766]&m[1769]&~m[1770]&m[1771]&~m[1772])|(m[1766]&~m[1769]&m[1770]&m[1771]&~m[1772])|(~m[1766]&m[1769]&~m[1770]&~m[1771]&m[1772])|(~m[1766]&~m[1769]&m[1770]&~m[1771]&m[1772])|(m[1766]&m[1769]&m[1770]&~m[1771]&m[1772])|(~m[1766]&m[1769]&m[1770]&m[1771]&m[1772]))&UnbiasedRNG[199])|((m[1766]&~m[1769]&~m[1770]&m[1771]&~m[1772])|(~m[1766]&~m[1769]&~m[1770]&~m[1771]&m[1772])|(m[1766]&~m[1769]&~m[1770]&~m[1771]&m[1772])|(m[1766]&m[1769]&~m[1770]&~m[1771]&m[1772])|(m[1766]&~m[1769]&m[1770]&~m[1771]&m[1772])|(~m[1766]&~m[1769]&~m[1770]&m[1771]&m[1772])|(m[1766]&~m[1769]&~m[1770]&m[1771]&m[1772])|(~m[1766]&m[1769]&~m[1770]&m[1771]&m[1772])|(m[1766]&m[1769]&~m[1770]&m[1771]&m[1772])|(~m[1766]&~m[1769]&m[1770]&m[1771]&m[1772])|(m[1766]&~m[1769]&m[1770]&m[1771]&m[1772])|(m[1766]&m[1769]&m[1770]&m[1771]&m[1772]));
    m[1773] = (((m[1771]&~m[1774]&~m[1775]&~m[1776]&~m[1777])|(~m[1771]&~m[1774]&~m[1775]&m[1776]&~m[1777])|(m[1771]&m[1774]&~m[1775]&m[1776]&~m[1777])|(m[1771]&~m[1774]&m[1775]&m[1776]&~m[1777])|(~m[1771]&m[1774]&~m[1775]&~m[1776]&m[1777])|(~m[1771]&~m[1774]&m[1775]&~m[1776]&m[1777])|(m[1771]&m[1774]&m[1775]&~m[1776]&m[1777])|(~m[1771]&m[1774]&m[1775]&m[1776]&m[1777]))&UnbiasedRNG[200])|((m[1771]&~m[1774]&~m[1775]&m[1776]&~m[1777])|(~m[1771]&~m[1774]&~m[1775]&~m[1776]&m[1777])|(m[1771]&~m[1774]&~m[1775]&~m[1776]&m[1777])|(m[1771]&m[1774]&~m[1775]&~m[1776]&m[1777])|(m[1771]&~m[1774]&m[1775]&~m[1776]&m[1777])|(~m[1771]&~m[1774]&~m[1775]&m[1776]&m[1777])|(m[1771]&~m[1774]&~m[1775]&m[1776]&m[1777])|(~m[1771]&m[1774]&~m[1775]&m[1776]&m[1777])|(m[1771]&m[1774]&~m[1775]&m[1776]&m[1777])|(~m[1771]&~m[1774]&m[1775]&m[1776]&m[1777])|(m[1771]&~m[1774]&m[1775]&m[1776]&m[1777])|(m[1771]&m[1774]&m[1775]&m[1776]&m[1777]));
    m[1778] = (((m[1776]&~m[1779]&~m[1780]&~m[1781]&~m[1782])|(~m[1776]&~m[1779]&~m[1780]&m[1781]&~m[1782])|(m[1776]&m[1779]&~m[1780]&m[1781]&~m[1782])|(m[1776]&~m[1779]&m[1780]&m[1781]&~m[1782])|(~m[1776]&m[1779]&~m[1780]&~m[1781]&m[1782])|(~m[1776]&~m[1779]&m[1780]&~m[1781]&m[1782])|(m[1776]&m[1779]&m[1780]&~m[1781]&m[1782])|(~m[1776]&m[1779]&m[1780]&m[1781]&m[1782]))&UnbiasedRNG[201])|((m[1776]&~m[1779]&~m[1780]&m[1781]&~m[1782])|(~m[1776]&~m[1779]&~m[1780]&~m[1781]&m[1782])|(m[1776]&~m[1779]&~m[1780]&~m[1781]&m[1782])|(m[1776]&m[1779]&~m[1780]&~m[1781]&m[1782])|(m[1776]&~m[1779]&m[1780]&~m[1781]&m[1782])|(~m[1776]&~m[1779]&~m[1780]&m[1781]&m[1782])|(m[1776]&~m[1779]&~m[1780]&m[1781]&m[1782])|(~m[1776]&m[1779]&~m[1780]&m[1781]&m[1782])|(m[1776]&m[1779]&~m[1780]&m[1781]&m[1782])|(~m[1776]&~m[1779]&m[1780]&m[1781]&m[1782])|(m[1776]&~m[1779]&m[1780]&m[1781]&m[1782])|(m[1776]&m[1779]&m[1780]&m[1781]&m[1782]));
    m[1783] = (((m[1781]&~m[1784]&~m[1785]&~m[1786]&~m[1787])|(~m[1781]&~m[1784]&~m[1785]&m[1786]&~m[1787])|(m[1781]&m[1784]&~m[1785]&m[1786]&~m[1787])|(m[1781]&~m[1784]&m[1785]&m[1786]&~m[1787])|(~m[1781]&m[1784]&~m[1785]&~m[1786]&m[1787])|(~m[1781]&~m[1784]&m[1785]&~m[1786]&m[1787])|(m[1781]&m[1784]&m[1785]&~m[1786]&m[1787])|(~m[1781]&m[1784]&m[1785]&m[1786]&m[1787]))&UnbiasedRNG[202])|((m[1781]&~m[1784]&~m[1785]&m[1786]&~m[1787])|(~m[1781]&~m[1784]&~m[1785]&~m[1786]&m[1787])|(m[1781]&~m[1784]&~m[1785]&~m[1786]&m[1787])|(m[1781]&m[1784]&~m[1785]&~m[1786]&m[1787])|(m[1781]&~m[1784]&m[1785]&~m[1786]&m[1787])|(~m[1781]&~m[1784]&~m[1785]&m[1786]&m[1787])|(m[1781]&~m[1784]&~m[1785]&m[1786]&m[1787])|(~m[1781]&m[1784]&~m[1785]&m[1786]&m[1787])|(m[1781]&m[1784]&~m[1785]&m[1786]&m[1787])|(~m[1781]&~m[1784]&m[1785]&m[1786]&m[1787])|(m[1781]&~m[1784]&m[1785]&m[1786]&m[1787])|(m[1781]&m[1784]&m[1785]&m[1786]&m[1787]));
    m[1788] = (((m[1786]&~m[1789]&~m[1790]&~m[1791]&~m[1792])|(~m[1786]&~m[1789]&~m[1790]&m[1791]&~m[1792])|(m[1786]&m[1789]&~m[1790]&m[1791]&~m[1792])|(m[1786]&~m[1789]&m[1790]&m[1791]&~m[1792])|(~m[1786]&m[1789]&~m[1790]&~m[1791]&m[1792])|(~m[1786]&~m[1789]&m[1790]&~m[1791]&m[1792])|(m[1786]&m[1789]&m[1790]&~m[1791]&m[1792])|(~m[1786]&m[1789]&m[1790]&m[1791]&m[1792]))&UnbiasedRNG[203])|((m[1786]&~m[1789]&~m[1790]&m[1791]&~m[1792])|(~m[1786]&~m[1789]&~m[1790]&~m[1791]&m[1792])|(m[1786]&~m[1789]&~m[1790]&~m[1791]&m[1792])|(m[1786]&m[1789]&~m[1790]&~m[1791]&m[1792])|(m[1786]&~m[1789]&m[1790]&~m[1791]&m[1792])|(~m[1786]&~m[1789]&~m[1790]&m[1791]&m[1792])|(m[1786]&~m[1789]&~m[1790]&m[1791]&m[1792])|(~m[1786]&m[1789]&~m[1790]&m[1791]&m[1792])|(m[1786]&m[1789]&~m[1790]&m[1791]&m[1792])|(~m[1786]&~m[1789]&m[1790]&m[1791]&m[1792])|(m[1786]&~m[1789]&m[1790]&m[1791]&m[1792])|(m[1786]&m[1789]&m[1790]&m[1791]&m[1792]));
    m[1793] = (((m[1791]&~m[1794]&~m[1795]&~m[1796]&~m[1797])|(~m[1791]&~m[1794]&~m[1795]&m[1796]&~m[1797])|(m[1791]&m[1794]&~m[1795]&m[1796]&~m[1797])|(m[1791]&~m[1794]&m[1795]&m[1796]&~m[1797])|(~m[1791]&m[1794]&~m[1795]&~m[1796]&m[1797])|(~m[1791]&~m[1794]&m[1795]&~m[1796]&m[1797])|(m[1791]&m[1794]&m[1795]&~m[1796]&m[1797])|(~m[1791]&m[1794]&m[1795]&m[1796]&m[1797]))&UnbiasedRNG[204])|((m[1791]&~m[1794]&~m[1795]&m[1796]&~m[1797])|(~m[1791]&~m[1794]&~m[1795]&~m[1796]&m[1797])|(m[1791]&~m[1794]&~m[1795]&~m[1796]&m[1797])|(m[1791]&m[1794]&~m[1795]&~m[1796]&m[1797])|(m[1791]&~m[1794]&m[1795]&~m[1796]&m[1797])|(~m[1791]&~m[1794]&~m[1795]&m[1796]&m[1797])|(m[1791]&~m[1794]&~m[1795]&m[1796]&m[1797])|(~m[1791]&m[1794]&~m[1795]&m[1796]&m[1797])|(m[1791]&m[1794]&~m[1795]&m[1796]&m[1797])|(~m[1791]&~m[1794]&m[1795]&m[1796]&m[1797])|(m[1791]&~m[1794]&m[1795]&m[1796]&m[1797])|(m[1791]&m[1794]&m[1795]&m[1796]&m[1797]));
    m[1798] = (((m[1742]&~m[1799]&~m[1800]&~m[1801]&~m[1802])|(~m[1742]&~m[1799]&~m[1800]&m[1801]&~m[1802])|(m[1742]&m[1799]&~m[1800]&m[1801]&~m[1802])|(m[1742]&~m[1799]&m[1800]&m[1801]&~m[1802])|(~m[1742]&m[1799]&~m[1800]&~m[1801]&m[1802])|(~m[1742]&~m[1799]&m[1800]&~m[1801]&m[1802])|(m[1742]&m[1799]&m[1800]&~m[1801]&m[1802])|(~m[1742]&m[1799]&m[1800]&m[1801]&m[1802]))&UnbiasedRNG[205])|((m[1742]&~m[1799]&~m[1800]&m[1801]&~m[1802])|(~m[1742]&~m[1799]&~m[1800]&~m[1801]&m[1802])|(m[1742]&~m[1799]&~m[1800]&~m[1801]&m[1802])|(m[1742]&m[1799]&~m[1800]&~m[1801]&m[1802])|(m[1742]&~m[1799]&m[1800]&~m[1801]&m[1802])|(~m[1742]&~m[1799]&~m[1800]&m[1801]&m[1802])|(m[1742]&~m[1799]&~m[1800]&m[1801]&m[1802])|(~m[1742]&m[1799]&~m[1800]&m[1801]&m[1802])|(m[1742]&m[1799]&~m[1800]&m[1801]&m[1802])|(~m[1742]&~m[1799]&m[1800]&m[1801]&m[1802])|(m[1742]&~m[1799]&m[1800]&m[1801]&m[1802])|(m[1742]&m[1799]&m[1800]&m[1801]&m[1802]));
    m[1803] = (((m[1801]&~m[1804]&~m[1805]&~m[1806]&~m[1807])|(~m[1801]&~m[1804]&~m[1805]&m[1806]&~m[1807])|(m[1801]&m[1804]&~m[1805]&m[1806]&~m[1807])|(m[1801]&~m[1804]&m[1805]&m[1806]&~m[1807])|(~m[1801]&m[1804]&~m[1805]&~m[1806]&m[1807])|(~m[1801]&~m[1804]&m[1805]&~m[1806]&m[1807])|(m[1801]&m[1804]&m[1805]&~m[1806]&m[1807])|(~m[1801]&m[1804]&m[1805]&m[1806]&m[1807]))&UnbiasedRNG[206])|((m[1801]&~m[1804]&~m[1805]&m[1806]&~m[1807])|(~m[1801]&~m[1804]&~m[1805]&~m[1806]&m[1807])|(m[1801]&~m[1804]&~m[1805]&~m[1806]&m[1807])|(m[1801]&m[1804]&~m[1805]&~m[1806]&m[1807])|(m[1801]&~m[1804]&m[1805]&~m[1806]&m[1807])|(~m[1801]&~m[1804]&~m[1805]&m[1806]&m[1807])|(m[1801]&~m[1804]&~m[1805]&m[1806]&m[1807])|(~m[1801]&m[1804]&~m[1805]&m[1806]&m[1807])|(m[1801]&m[1804]&~m[1805]&m[1806]&m[1807])|(~m[1801]&~m[1804]&m[1805]&m[1806]&m[1807])|(m[1801]&~m[1804]&m[1805]&m[1806]&m[1807])|(m[1801]&m[1804]&m[1805]&m[1806]&m[1807]));
    m[1808] = (((m[1806]&~m[1809]&~m[1810]&~m[1811]&~m[1812])|(~m[1806]&~m[1809]&~m[1810]&m[1811]&~m[1812])|(m[1806]&m[1809]&~m[1810]&m[1811]&~m[1812])|(m[1806]&~m[1809]&m[1810]&m[1811]&~m[1812])|(~m[1806]&m[1809]&~m[1810]&~m[1811]&m[1812])|(~m[1806]&~m[1809]&m[1810]&~m[1811]&m[1812])|(m[1806]&m[1809]&m[1810]&~m[1811]&m[1812])|(~m[1806]&m[1809]&m[1810]&m[1811]&m[1812]))&UnbiasedRNG[207])|((m[1806]&~m[1809]&~m[1810]&m[1811]&~m[1812])|(~m[1806]&~m[1809]&~m[1810]&~m[1811]&m[1812])|(m[1806]&~m[1809]&~m[1810]&~m[1811]&m[1812])|(m[1806]&m[1809]&~m[1810]&~m[1811]&m[1812])|(m[1806]&~m[1809]&m[1810]&~m[1811]&m[1812])|(~m[1806]&~m[1809]&~m[1810]&m[1811]&m[1812])|(m[1806]&~m[1809]&~m[1810]&m[1811]&m[1812])|(~m[1806]&m[1809]&~m[1810]&m[1811]&m[1812])|(m[1806]&m[1809]&~m[1810]&m[1811]&m[1812])|(~m[1806]&~m[1809]&m[1810]&m[1811]&m[1812])|(m[1806]&~m[1809]&m[1810]&m[1811]&m[1812])|(m[1806]&m[1809]&m[1810]&m[1811]&m[1812]));
    m[1813] = (((m[1811]&~m[1814]&~m[1815]&~m[1816]&~m[1817])|(~m[1811]&~m[1814]&~m[1815]&m[1816]&~m[1817])|(m[1811]&m[1814]&~m[1815]&m[1816]&~m[1817])|(m[1811]&~m[1814]&m[1815]&m[1816]&~m[1817])|(~m[1811]&m[1814]&~m[1815]&~m[1816]&m[1817])|(~m[1811]&~m[1814]&m[1815]&~m[1816]&m[1817])|(m[1811]&m[1814]&m[1815]&~m[1816]&m[1817])|(~m[1811]&m[1814]&m[1815]&m[1816]&m[1817]))&UnbiasedRNG[208])|((m[1811]&~m[1814]&~m[1815]&m[1816]&~m[1817])|(~m[1811]&~m[1814]&~m[1815]&~m[1816]&m[1817])|(m[1811]&~m[1814]&~m[1815]&~m[1816]&m[1817])|(m[1811]&m[1814]&~m[1815]&~m[1816]&m[1817])|(m[1811]&~m[1814]&m[1815]&~m[1816]&m[1817])|(~m[1811]&~m[1814]&~m[1815]&m[1816]&m[1817])|(m[1811]&~m[1814]&~m[1815]&m[1816]&m[1817])|(~m[1811]&m[1814]&~m[1815]&m[1816]&m[1817])|(m[1811]&m[1814]&~m[1815]&m[1816]&m[1817])|(~m[1811]&~m[1814]&m[1815]&m[1816]&m[1817])|(m[1811]&~m[1814]&m[1815]&m[1816]&m[1817])|(m[1811]&m[1814]&m[1815]&m[1816]&m[1817]));
    m[1818] = (((m[1816]&~m[1819]&~m[1820]&~m[1821]&~m[1822])|(~m[1816]&~m[1819]&~m[1820]&m[1821]&~m[1822])|(m[1816]&m[1819]&~m[1820]&m[1821]&~m[1822])|(m[1816]&~m[1819]&m[1820]&m[1821]&~m[1822])|(~m[1816]&m[1819]&~m[1820]&~m[1821]&m[1822])|(~m[1816]&~m[1819]&m[1820]&~m[1821]&m[1822])|(m[1816]&m[1819]&m[1820]&~m[1821]&m[1822])|(~m[1816]&m[1819]&m[1820]&m[1821]&m[1822]))&UnbiasedRNG[209])|((m[1816]&~m[1819]&~m[1820]&m[1821]&~m[1822])|(~m[1816]&~m[1819]&~m[1820]&~m[1821]&m[1822])|(m[1816]&~m[1819]&~m[1820]&~m[1821]&m[1822])|(m[1816]&m[1819]&~m[1820]&~m[1821]&m[1822])|(m[1816]&~m[1819]&m[1820]&~m[1821]&m[1822])|(~m[1816]&~m[1819]&~m[1820]&m[1821]&m[1822])|(m[1816]&~m[1819]&~m[1820]&m[1821]&m[1822])|(~m[1816]&m[1819]&~m[1820]&m[1821]&m[1822])|(m[1816]&m[1819]&~m[1820]&m[1821]&m[1822])|(~m[1816]&~m[1819]&m[1820]&m[1821]&m[1822])|(m[1816]&~m[1819]&m[1820]&m[1821]&m[1822])|(m[1816]&m[1819]&m[1820]&m[1821]&m[1822]));
    m[1823] = (((m[1821]&~m[1824]&~m[1825]&~m[1826]&~m[1827])|(~m[1821]&~m[1824]&~m[1825]&m[1826]&~m[1827])|(m[1821]&m[1824]&~m[1825]&m[1826]&~m[1827])|(m[1821]&~m[1824]&m[1825]&m[1826]&~m[1827])|(~m[1821]&m[1824]&~m[1825]&~m[1826]&m[1827])|(~m[1821]&~m[1824]&m[1825]&~m[1826]&m[1827])|(m[1821]&m[1824]&m[1825]&~m[1826]&m[1827])|(~m[1821]&m[1824]&m[1825]&m[1826]&m[1827]))&UnbiasedRNG[210])|((m[1821]&~m[1824]&~m[1825]&m[1826]&~m[1827])|(~m[1821]&~m[1824]&~m[1825]&~m[1826]&m[1827])|(m[1821]&~m[1824]&~m[1825]&~m[1826]&m[1827])|(m[1821]&m[1824]&~m[1825]&~m[1826]&m[1827])|(m[1821]&~m[1824]&m[1825]&~m[1826]&m[1827])|(~m[1821]&~m[1824]&~m[1825]&m[1826]&m[1827])|(m[1821]&~m[1824]&~m[1825]&m[1826]&m[1827])|(~m[1821]&m[1824]&~m[1825]&m[1826]&m[1827])|(m[1821]&m[1824]&~m[1825]&m[1826]&m[1827])|(~m[1821]&~m[1824]&m[1825]&m[1826]&m[1827])|(m[1821]&~m[1824]&m[1825]&m[1826]&m[1827])|(m[1821]&m[1824]&m[1825]&m[1826]&m[1827]));
    m[1828] = (((m[1826]&~m[1829]&~m[1830]&~m[1831]&~m[1832])|(~m[1826]&~m[1829]&~m[1830]&m[1831]&~m[1832])|(m[1826]&m[1829]&~m[1830]&m[1831]&~m[1832])|(m[1826]&~m[1829]&m[1830]&m[1831]&~m[1832])|(~m[1826]&m[1829]&~m[1830]&~m[1831]&m[1832])|(~m[1826]&~m[1829]&m[1830]&~m[1831]&m[1832])|(m[1826]&m[1829]&m[1830]&~m[1831]&m[1832])|(~m[1826]&m[1829]&m[1830]&m[1831]&m[1832]))&UnbiasedRNG[211])|((m[1826]&~m[1829]&~m[1830]&m[1831]&~m[1832])|(~m[1826]&~m[1829]&~m[1830]&~m[1831]&m[1832])|(m[1826]&~m[1829]&~m[1830]&~m[1831]&m[1832])|(m[1826]&m[1829]&~m[1830]&~m[1831]&m[1832])|(m[1826]&~m[1829]&m[1830]&~m[1831]&m[1832])|(~m[1826]&~m[1829]&~m[1830]&m[1831]&m[1832])|(m[1826]&~m[1829]&~m[1830]&m[1831]&m[1832])|(~m[1826]&m[1829]&~m[1830]&m[1831]&m[1832])|(m[1826]&m[1829]&~m[1830]&m[1831]&m[1832])|(~m[1826]&~m[1829]&m[1830]&m[1831]&m[1832])|(m[1826]&~m[1829]&m[1830]&m[1831]&m[1832])|(m[1826]&m[1829]&m[1830]&m[1831]&m[1832]));
    m[1833] = (((m[1831]&~m[1834]&~m[1835]&~m[1836]&~m[1837])|(~m[1831]&~m[1834]&~m[1835]&m[1836]&~m[1837])|(m[1831]&m[1834]&~m[1835]&m[1836]&~m[1837])|(m[1831]&~m[1834]&m[1835]&m[1836]&~m[1837])|(~m[1831]&m[1834]&~m[1835]&~m[1836]&m[1837])|(~m[1831]&~m[1834]&m[1835]&~m[1836]&m[1837])|(m[1831]&m[1834]&m[1835]&~m[1836]&m[1837])|(~m[1831]&m[1834]&m[1835]&m[1836]&m[1837]))&UnbiasedRNG[212])|((m[1831]&~m[1834]&~m[1835]&m[1836]&~m[1837])|(~m[1831]&~m[1834]&~m[1835]&~m[1836]&m[1837])|(m[1831]&~m[1834]&~m[1835]&~m[1836]&m[1837])|(m[1831]&m[1834]&~m[1835]&~m[1836]&m[1837])|(m[1831]&~m[1834]&m[1835]&~m[1836]&m[1837])|(~m[1831]&~m[1834]&~m[1835]&m[1836]&m[1837])|(m[1831]&~m[1834]&~m[1835]&m[1836]&m[1837])|(~m[1831]&m[1834]&~m[1835]&m[1836]&m[1837])|(m[1831]&m[1834]&~m[1835]&m[1836]&m[1837])|(~m[1831]&~m[1834]&m[1835]&m[1836]&m[1837])|(m[1831]&~m[1834]&m[1835]&m[1836]&m[1837])|(m[1831]&m[1834]&m[1835]&m[1836]&m[1837]));
    m[1838] = (((m[1836]&~m[1839]&~m[1840]&~m[1841]&~m[1842])|(~m[1836]&~m[1839]&~m[1840]&m[1841]&~m[1842])|(m[1836]&m[1839]&~m[1840]&m[1841]&~m[1842])|(m[1836]&~m[1839]&m[1840]&m[1841]&~m[1842])|(~m[1836]&m[1839]&~m[1840]&~m[1841]&m[1842])|(~m[1836]&~m[1839]&m[1840]&~m[1841]&m[1842])|(m[1836]&m[1839]&m[1840]&~m[1841]&m[1842])|(~m[1836]&m[1839]&m[1840]&m[1841]&m[1842]))&UnbiasedRNG[213])|((m[1836]&~m[1839]&~m[1840]&m[1841]&~m[1842])|(~m[1836]&~m[1839]&~m[1840]&~m[1841]&m[1842])|(m[1836]&~m[1839]&~m[1840]&~m[1841]&m[1842])|(m[1836]&m[1839]&~m[1840]&~m[1841]&m[1842])|(m[1836]&~m[1839]&m[1840]&~m[1841]&m[1842])|(~m[1836]&~m[1839]&~m[1840]&m[1841]&m[1842])|(m[1836]&~m[1839]&~m[1840]&m[1841]&m[1842])|(~m[1836]&m[1839]&~m[1840]&m[1841]&m[1842])|(m[1836]&m[1839]&~m[1840]&m[1841]&m[1842])|(~m[1836]&~m[1839]&m[1840]&m[1841]&m[1842])|(m[1836]&~m[1839]&m[1840]&m[1841]&m[1842])|(m[1836]&m[1839]&m[1840]&m[1841]&m[1842]));
    m[1843] = (((m[1841]&~m[1844]&~m[1845]&~m[1846]&~m[1847])|(~m[1841]&~m[1844]&~m[1845]&m[1846]&~m[1847])|(m[1841]&m[1844]&~m[1845]&m[1846]&~m[1847])|(m[1841]&~m[1844]&m[1845]&m[1846]&~m[1847])|(~m[1841]&m[1844]&~m[1845]&~m[1846]&m[1847])|(~m[1841]&~m[1844]&m[1845]&~m[1846]&m[1847])|(m[1841]&m[1844]&m[1845]&~m[1846]&m[1847])|(~m[1841]&m[1844]&m[1845]&m[1846]&m[1847]))&UnbiasedRNG[214])|((m[1841]&~m[1844]&~m[1845]&m[1846]&~m[1847])|(~m[1841]&~m[1844]&~m[1845]&~m[1846]&m[1847])|(m[1841]&~m[1844]&~m[1845]&~m[1846]&m[1847])|(m[1841]&m[1844]&~m[1845]&~m[1846]&m[1847])|(m[1841]&~m[1844]&m[1845]&~m[1846]&m[1847])|(~m[1841]&~m[1844]&~m[1845]&m[1846]&m[1847])|(m[1841]&~m[1844]&~m[1845]&m[1846]&m[1847])|(~m[1841]&m[1844]&~m[1845]&m[1846]&m[1847])|(m[1841]&m[1844]&~m[1845]&m[1846]&m[1847])|(~m[1841]&~m[1844]&m[1845]&m[1846]&m[1847])|(m[1841]&~m[1844]&m[1845]&m[1846]&m[1847])|(m[1841]&m[1844]&m[1845]&m[1846]&m[1847]));
    m[1848] = (((m[1846]&~m[1849]&~m[1850]&~m[1851]&~m[1852])|(~m[1846]&~m[1849]&~m[1850]&m[1851]&~m[1852])|(m[1846]&m[1849]&~m[1850]&m[1851]&~m[1852])|(m[1846]&~m[1849]&m[1850]&m[1851]&~m[1852])|(~m[1846]&m[1849]&~m[1850]&~m[1851]&m[1852])|(~m[1846]&~m[1849]&m[1850]&~m[1851]&m[1852])|(m[1846]&m[1849]&m[1850]&~m[1851]&m[1852])|(~m[1846]&m[1849]&m[1850]&m[1851]&m[1852]))&UnbiasedRNG[215])|((m[1846]&~m[1849]&~m[1850]&m[1851]&~m[1852])|(~m[1846]&~m[1849]&~m[1850]&~m[1851]&m[1852])|(m[1846]&~m[1849]&~m[1850]&~m[1851]&m[1852])|(m[1846]&m[1849]&~m[1850]&~m[1851]&m[1852])|(m[1846]&~m[1849]&m[1850]&~m[1851]&m[1852])|(~m[1846]&~m[1849]&~m[1850]&m[1851]&m[1852])|(m[1846]&~m[1849]&~m[1850]&m[1851]&m[1852])|(~m[1846]&m[1849]&~m[1850]&m[1851]&m[1852])|(m[1846]&m[1849]&~m[1850]&m[1851]&m[1852])|(~m[1846]&~m[1849]&m[1850]&m[1851]&m[1852])|(m[1846]&~m[1849]&m[1850]&m[1851]&m[1852])|(m[1846]&m[1849]&m[1850]&m[1851]&m[1852]));
    m[1853] = (((m[1802]&~m[1854]&~m[1855]&~m[1856]&~m[1857])|(~m[1802]&~m[1854]&~m[1855]&m[1856]&~m[1857])|(m[1802]&m[1854]&~m[1855]&m[1856]&~m[1857])|(m[1802]&~m[1854]&m[1855]&m[1856]&~m[1857])|(~m[1802]&m[1854]&~m[1855]&~m[1856]&m[1857])|(~m[1802]&~m[1854]&m[1855]&~m[1856]&m[1857])|(m[1802]&m[1854]&m[1855]&~m[1856]&m[1857])|(~m[1802]&m[1854]&m[1855]&m[1856]&m[1857]))&UnbiasedRNG[216])|((m[1802]&~m[1854]&~m[1855]&m[1856]&~m[1857])|(~m[1802]&~m[1854]&~m[1855]&~m[1856]&m[1857])|(m[1802]&~m[1854]&~m[1855]&~m[1856]&m[1857])|(m[1802]&m[1854]&~m[1855]&~m[1856]&m[1857])|(m[1802]&~m[1854]&m[1855]&~m[1856]&m[1857])|(~m[1802]&~m[1854]&~m[1855]&m[1856]&m[1857])|(m[1802]&~m[1854]&~m[1855]&m[1856]&m[1857])|(~m[1802]&m[1854]&~m[1855]&m[1856]&m[1857])|(m[1802]&m[1854]&~m[1855]&m[1856]&m[1857])|(~m[1802]&~m[1854]&m[1855]&m[1856]&m[1857])|(m[1802]&~m[1854]&m[1855]&m[1856]&m[1857])|(m[1802]&m[1854]&m[1855]&m[1856]&m[1857]));
    m[1858] = (((m[1856]&~m[1859]&~m[1860]&~m[1861]&~m[1862])|(~m[1856]&~m[1859]&~m[1860]&m[1861]&~m[1862])|(m[1856]&m[1859]&~m[1860]&m[1861]&~m[1862])|(m[1856]&~m[1859]&m[1860]&m[1861]&~m[1862])|(~m[1856]&m[1859]&~m[1860]&~m[1861]&m[1862])|(~m[1856]&~m[1859]&m[1860]&~m[1861]&m[1862])|(m[1856]&m[1859]&m[1860]&~m[1861]&m[1862])|(~m[1856]&m[1859]&m[1860]&m[1861]&m[1862]))&UnbiasedRNG[217])|((m[1856]&~m[1859]&~m[1860]&m[1861]&~m[1862])|(~m[1856]&~m[1859]&~m[1860]&~m[1861]&m[1862])|(m[1856]&~m[1859]&~m[1860]&~m[1861]&m[1862])|(m[1856]&m[1859]&~m[1860]&~m[1861]&m[1862])|(m[1856]&~m[1859]&m[1860]&~m[1861]&m[1862])|(~m[1856]&~m[1859]&~m[1860]&m[1861]&m[1862])|(m[1856]&~m[1859]&~m[1860]&m[1861]&m[1862])|(~m[1856]&m[1859]&~m[1860]&m[1861]&m[1862])|(m[1856]&m[1859]&~m[1860]&m[1861]&m[1862])|(~m[1856]&~m[1859]&m[1860]&m[1861]&m[1862])|(m[1856]&~m[1859]&m[1860]&m[1861]&m[1862])|(m[1856]&m[1859]&m[1860]&m[1861]&m[1862]));
    m[1863] = (((m[1861]&~m[1864]&~m[1865]&~m[1866]&~m[1867])|(~m[1861]&~m[1864]&~m[1865]&m[1866]&~m[1867])|(m[1861]&m[1864]&~m[1865]&m[1866]&~m[1867])|(m[1861]&~m[1864]&m[1865]&m[1866]&~m[1867])|(~m[1861]&m[1864]&~m[1865]&~m[1866]&m[1867])|(~m[1861]&~m[1864]&m[1865]&~m[1866]&m[1867])|(m[1861]&m[1864]&m[1865]&~m[1866]&m[1867])|(~m[1861]&m[1864]&m[1865]&m[1866]&m[1867]))&UnbiasedRNG[218])|((m[1861]&~m[1864]&~m[1865]&m[1866]&~m[1867])|(~m[1861]&~m[1864]&~m[1865]&~m[1866]&m[1867])|(m[1861]&~m[1864]&~m[1865]&~m[1866]&m[1867])|(m[1861]&m[1864]&~m[1865]&~m[1866]&m[1867])|(m[1861]&~m[1864]&m[1865]&~m[1866]&m[1867])|(~m[1861]&~m[1864]&~m[1865]&m[1866]&m[1867])|(m[1861]&~m[1864]&~m[1865]&m[1866]&m[1867])|(~m[1861]&m[1864]&~m[1865]&m[1866]&m[1867])|(m[1861]&m[1864]&~m[1865]&m[1866]&m[1867])|(~m[1861]&~m[1864]&m[1865]&m[1866]&m[1867])|(m[1861]&~m[1864]&m[1865]&m[1866]&m[1867])|(m[1861]&m[1864]&m[1865]&m[1866]&m[1867]));
    m[1868] = (((m[1866]&~m[1869]&~m[1870]&~m[1871]&~m[1872])|(~m[1866]&~m[1869]&~m[1870]&m[1871]&~m[1872])|(m[1866]&m[1869]&~m[1870]&m[1871]&~m[1872])|(m[1866]&~m[1869]&m[1870]&m[1871]&~m[1872])|(~m[1866]&m[1869]&~m[1870]&~m[1871]&m[1872])|(~m[1866]&~m[1869]&m[1870]&~m[1871]&m[1872])|(m[1866]&m[1869]&m[1870]&~m[1871]&m[1872])|(~m[1866]&m[1869]&m[1870]&m[1871]&m[1872]))&UnbiasedRNG[219])|((m[1866]&~m[1869]&~m[1870]&m[1871]&~m[1872])|(~m[1866]&~m[1869]&~m[1870]&~m[1871]&m[1872])|(m[1866]&~m[1869]&~m[1870]&~m[1871]&m[1872])|(m[1866]&m[1869]&~m[1870]&~m[1871]&m[1872])|(m[1866]&~m[1869]&m[1870]&~m[1871]&m[1872])|(~m[1866]&~m[1869]&~m[1870]&m[1871]&m[1872])|(m[1866]&~m[1869]&~m[1870]&m[1871]&m[1872])|(~m[1866]&m[1869]&~m[1870]&m[1871]&m[1872])|(m[1866]&m[1869]&~m[1870]&m[1871]&m[1872])|(~m[1866]&~m[1869]&m[1870]&m[1871]&m[1872])|(m[1866]&~m[1869]&m[1870]&m[1871]&m[1872])|(m[1866]&m[1869]&m[1870]&m[1871]&m[1872]));
    m[1873] = (((m[1871]&~m[1874]&~m[1875]&~m[1876]&~m[1877])|(~m[1871]&~m[1874]&~m[1875]&m[1876]&~m[1877])|(m[1871]&m[1874]&~m[1875]&m[1876]&~m[1877])|(m[1871]&~m[1874]&m[1875]&m[1876]&~m[1877])|(~m[1871]&m[1874]&~m[1875]&~m[1876]&m[1877])|(~m[1871]&~m[1874]&m[1875]&~m[1876]&m[1877])|(m[1871]&m[1874]&m[1875]&~m[1876]&m[1877])|(~m[1871]&m[1874]&m[1875]&m[1876]&m[1877]))&UnbiasedRNG[220])|((m[1871]&~m[1874]&~m[1875]&m[1876]&~m[1877])|(~m[1871]&~m[1874]&~m[1875]&~m[1876]&m[1877])|(m[1871]&~m[1874]&~m[1875]&~m[1876]&m[1877])|(m[1871]&m[1874]&~m[1875]&~m[1876]&m[1877])|(m[1871]&~m[1874]&m[1875]&~m[1876]&m[1877])|(~m[1871]&~m[1874]&~m[1875]&m[1876]&m[1877])|(m[1871]&~m[1874]&~m[1875]&m[1876]&m[1877])|(~m[1871]&m[1874]&~m[1875]&m[1876]&m[1877])|(m[1871]&m[1874]&~m[1875]&m[1876]&m[1877])|(~m[1871]&~m[1874]&m[1875]&m[1876]&m[1877])|(m[1871]&~m[1874]&m[1875]&m[1876]&m[1877])|(m[1871]&m[1874]&m[1875]&m[1876]&m[1877]));
    m[1878] = (((m[1876]&~m[1879]&~m[1880]&~m[1881]&~m[1882])|(~m[1876]&~m[1879]&~m[1880]&m[1881]&~m[1882])|(m[1876]&m[1879]&~m[1880]&m[1881]&~m[1882])|(m[1876]&~m[1879]&m[1880]&m[1881]&~m[1882])|(~m[1876]&m[1879]&~m[1880]&~m[1881]&m[1882])|(~m[1876]&~m[1879]&m[1880]&~m[1881]&m[1882])|(m[1876]&m[1879]&m[1880]&~m[1881]&m[1882])|(~m[1876]&m[1879]&m[1880]&m[1881]&m[1882]))&UnbiasedRNG[221])|((m[1876]&~m[1879]&~m[1880]&m[1881]&~m[1882])|(~m[1876]&~m[1879]&~m[1880]&~m[1881]&m[1882])|(m[1876]&~m[1879]&~m[1880]&~m[1881]&m[1882])|(m[1876]&m[1879]&~m[1880]&~m[1881]&m[1882])|(m[1876]&~m[1879]&m[1880]&~m[1881]&m[1882])|(~m[1876]&~m[1879]&~m[1880]&m[1881]&m[1882])|(m[1876]&~m[1879]&~m[1880]&m[1881]&m[1882])|(~m[1876]&m[1879]&~m[1880]&m[1881]&m[1882])|(m[1876]&m[1879]&~m[1880]&m[1881]&m[1882])|(~m[1876]&~m[1879]&m[1880]&m[1881]&m[1882])|(m[1876]&~m[1879]&m[1880]&m[1881]&m[1882])|(m[1876]&m[1879]&m[1880]&m[1881]&m[1882]));
    m[1883] = (((m[1881]&~m[1884]&~m[1885]&~m[1886]&~m[1887])|(~m[1881]&~m[1884]&~m[1885]&m[1886]&~m[1887])|(m[1881]&m[1884]&~m[1885]&m[1886]&~m[1887])|(m[1881]&~m[1884]&m[1885]&m[1886]&~m[1887])|(~m[1881]&m[1884]&~m[1885]&~m[1886]&m[1887])|(~m[1881]&~m[1884]&m[1885]&~m[1886]&m[1887])|(m[1881]&m[1884]&m[1885]&~m[1886]&m[1887])|(~m[1881]&m[1884]&m[1885]&m[1886]&m[1887]))&UnbiasedRNG[222])|((m[1881]&~m[1884]&~m[1885]&m[1886]&~m[1887])|(~m[1881]&~m[1884]&~m[1885]&~m[1886]&m[1887])|(m[1881]&~m[1884]&~m[1885]&~m[1886]&m[1887])|(m[1881]&m[1884]&~m[1885]&~m[1886]&m[1887])|(m[1881]&~m[1884]&m[1885]&~m[1886]&m[1887])|(~m[1881]&~m[1884]&~m[1885]&m[1886]&m[1887])|(m[1881]&~m[1884]&~m[1885]&m[1886]&m[1887])|(~m[1881]&m[1884]&~m[1885]&m[1886]&m[1887])|(m[1881]&m[1884]&~m[1885]&m[1886]&m[1887])|(~m[1881]&~m[1884]&m[1885]&m[1886]&m[1887])|(m[1881]&~m[1884]&m[1885]&m[1886]&m[1887])|(m[1881]&m[1884]&m[1885]&m[1886]&m[1887]));
    m[1888] = (((m[1886]&~m[1889]&~m[1890]&~m[1891]&~m[1892])|(~m[1886]&~m[1889]&~m[1890]&m[1891]&~m[1892])|(m[1886]&m[1889]&~m[1890]&m[1891]&~m[1892])|(m[1886]&~m[1889]&m[1890]&m[1891]&~m[1892])|(~m[1886]&m[1889]&~m[1890]&~m[1891]&m[1892])|(~m[1886]&~m[1889]&m[1890]&~m[1891]&m[1892])|(m[1886]&m[1889]&m[1890]&~m[1891]&m[1892])|(~m[1886]&m[1889]&m[1890]&m[1891]&m[1892]))&UnbiasedRNG[223])|((m[1886]&~m[1889]&~m[1890]&m[1891]&~m[1892])|(~m[1886]&~m[1889]&~m[1890]&~m[1891]&m[1892])|(m[1886]&~m[1889]&~m[1890]&~m[1891]&m[1892])|(m[1886]&m[1889]&~m[1890]&~m[1891]&m[1892])|(m[1886]&~m[1889]&m[1890]&~m[1891]&m[1892])|(~m[1886]&~m[1889]&~m[1890]&m[1891]&m[1892])|(m[1886]&~m[1889]&~m[1890]&m[1891]&m[1892])|(~m[1886]&m[1889]&~m[1890]&m[1891]&m[1892])|(m[1886]&m[1889]&~m[1890]&m[1891]&m[1892])|(~m[1886]&~m[1889]&m[1890]&m[1891]&m[1892])|(m[1886]&~m[1889]&m[1890]&m[1891]&m[1892])|(m[1886]&m[1889]&m[1890]&m[1891]&m[1892]));
    m[1893] = (((m[1891]&~m[1894]&~m[1895]&~m[1896]&~m[1897])|(~m[1891]&~m[1894]&~m[1895]&m[1896]&~m[1897])|(m[1891]&m[1894]&~m[1895]&m[1896]&~m[1897])|(m[1891]&~m[1894]&m[1895]&m[1896]&~m[1897])|(~m[1891]&m[1894]&~m[1895]&~m[1896]&m[1897])|(~m[1891]&~m[1894]&m[1895]&~m[1896]&m[1897])|(m[1891]&m[1894]&m[1895]&~m[1896]&m[1897])|(~m[1891]&m[1894]&m[1895]&m[1896]&m[1897]))&UnbiasedRNG[224])|((m[1891]&~m[1894]&~m[1895]&m[1896]&~m[1897])|(~m[1891]&~m[1894]&~m[1895]&~m[1896]&m[1897])|(m[1891]&~m[1894]&~m[1895]&~m[1896]&m[1897])|(m[1891]&m[1894]&~m[1895]&~m[1896]&m[1897])|(m[1891]&~m[1894]&m[1895]&~m[1896]&m[1897])|(~m[1891]&~m[1894]&~m[1895]&m[1896]&m[1897])|(m[1891]&~m[1894]&~m[1895]&m[1896]&m[1897])|(~m[1891]&m[1894]&~m[1895]&m[1896]&m[1897])|(m[1891]&m[1894]&~m[1895]&m[1896]&m[1897])|(~m[1891]&~m[1894]&m[1895]&m[1896]&m[1897])|(m[1891]&~m[1894]&m[1895]&m[1896]&m[1897])|(m[1891]&m[1894]&m[1895]&m[1896]&m[1897]));
    m[1898] = (((m[1896]&~m[1899]&~m[1900]&~m[1901]&~m[1902])|(~m[1896]&~m[1899]&~m[1900]&m[1901]&~m[1902])|(m[1896]&m[1899]&~m[1900]&m[1901]&~m[1902])|(m[1896]&~m[1899]&m[1900]&m[1901]&~m[1902])|(~m[1896]&m[1899]&~m[1900]&~m[1901]&m[1902])|(~m[1896]&~m[1899]&m[1900]&~m[1901]&m[1902])|(m[1896]&m[1899]&m[1900]&~m[1901]&m[1902])|(~m[1896]&m[1899]&m[1900]&m[1901]&m[1902]))&UnbiasedRNG[225])|((m[1896]&~m[1899]&~m[1900]&m[1901]&~m[1902])|(~m[1896]&~m[1899]&~m[1900]&~m[1901]&m[1902])|(m[1896]&~m[1899]&~m[1900]&~m[1901]&m[1902])|(m[1896]&m[1899]&~m[1900]&~m[1901]&m[1902])|(m[1896]&~m[1899]&m[1900]&~m[1901]&m[1902])|(~m[1896]&~m[1899]&~m[1900]&m[1901]&m[1902])|(m[1896]&~m[1899]&~m[1900]&m[1901]&m[1902])|(~m[1896]&m[1899]&~m[1900]&m[1901]&m[1902])|(m[1896]&m[1899]&~m[1900]&m[1901]&m[1902])|(~m[1896]&~m[1899]&m[1900]&m[1901]&m[1902])|(m[1896]&~m[1899]&m[1900]&m[1901]&m[1902])|(m[1896]&m[1899]&m[1900]&m[1901]&m[1902]));
    m[1903] = (((m[1857]&~m[1904]&~m[1905]&~m[1906]&~m[1907])|(~m[1857]&~m[1904]&~m[1905]&m[1906]&~m[1907])|(m[1857]&m[1904]&~m[1905]&m[1906]&~m[1907])|(m[1857]&~m[1904]&m[1905]&m[1906]&~m[1907])|(~m[1857]&m[1904]&~m[1905]&~m[1906]&m[1907])|(~m[1857]&~m[1904]&m[1905]&~m[1906]&m[1907])|(m[1857]&m[1904]&m[1905]&~m[1906]&m[1907])|(~m[1857]&m[1904]&m[1905]&m[1906]&m[1907]))&UnbiasedRNG[226])|((m[1857]&~m[1904]&~m[1905]&m[1906]&~m[1907])|(~m[1857]&~m[1904]&~m[1905]&~m[1906]&m[1907])|(m[1857]&~m[1904]&~m[1905]&~m[1906]&m[1907])|(m[1857]&m[1904]&~m[1905]&~m[1906]&m[1907])|(m[1857]&~m[1904]&m[1905]&~m[1906]&m[1907])|(~m[1857]&~m[1904]&~m[1905]&m[1906]&m[1907])|(m[1857]&~m[1904]&~m[1905]&m[1906]&m[1907])|(~m[1857]&m[1904]&~m[1905]&m[1906]&m[1907])|(m[1857]&m[1904]&~m[1905]&m[1906]&m[1907])|(~m[1857]&~m[1904]&m[1905]&m[1906]&m[1907])|(m[1857]&~m[1904]&m[1905]&m[1906]&m[1907])|(m[1857]&m[1904]&m[1905]&m[1906]&m[1907]));
    m[1908] = (((m[1906]&~m[1909]&~m[1910]&~m[1911]&~m[1912])|(~m[1906]&~m[1909]&~m[1910]&m[1911]&~m[1912])|(m[1906]&m[1909]&~m[1910]&m[1911]&~m[1912])|(m[1906]&~m[1909]&m[1910]&m[1911]&~m[1912])|(~m[1906]&m[1909]&~m[1910]&~m[1911]&m[1912])|(~m[1906]&~m[1909]&m[1910]&~m[1911]&m[1912])|(m[1906]&m[1909]&m[1910]&~m[1911]&m[1912])|(~m[1906]&m[1909]&m[1910]&m[1911]&m[1912]))&UnbiasedRNG[227])|((m[1906]&~m[1909]&~m[1910]&m[1911]&~m[1912])|(~m[1906]&~m[1909]&~m[1910]&~m[1911]&m[1912])|(m[1906]&~m[1909]&~m[1910]&~m[1911]&m[1912])|(m[1906]&m[1909]&~m[1910]&~m[1911]&m[1912])|(m[1906]&~m[1909]&m[1910]&~m[1911]&m[1912])|(~m[1906]&~m[1909]&~m[1910]&m[1911]&m[1912])|(m[1906]&~m[1909]&~m[1910]&m[1911]&m[1912])|(~m[1906]&m[1909]&~m[1910]&m[1911]&m[1912])|(m[1906]&m[1909]&~m[1910]&m[1911]&m[1912])|(~m[1906]&~m[1909]&m[1910]&m[1911]&m[1912])|(m[1906]&~m[1909]&m[1910]&m[1911]&m[1912])|(m[1906]&m[1909]&m[1910]&m[1911]&m[1912]));
    m[1913] = (((m[1911]&~m[1914]&~m[1915]&~m[1916]&~m[1917])|(~m[1911]&~m[1914]&~m[1915]&m[1916]&~m[1917])|(m[1911]&m[1914]&~m[1915]&m[1916]&~m[1917])|(m[1911]&~m[1914]&m[1915]&m[1916]&~m[1917])|(~m[1911]&m[1914]&~m[1915]&~m[1916]&m[1917])|(~m[1911]&~m[1914]&m[1915]&~m[1916]&m[1917])|(m[1911]&m[1914]&m[1915]&~m[1916]&m[1917])|(~m[1911]&m[1914]&m[1915]&m[1916]&m[1917]))&UnbiasedRNG[228])|((m[1911]&~m[1914]&~m[1915]&m[1916]&~m[1917])|(~m[1911]&~m[1914]&~m[1915]&~m[1916]&m[1917])|(m[1911]&~m[1914]&~m[1915]&~m[1916]&m[1917])|(m[1911]&m[1914]&~m[1915]&~m[1916]&m[1917])|(m[1911]&~m[1914]&m[1915]&~m[1916]&m[1917])|(~m[1911]&~m[1914]&~m[1915]&m[1916]&m[1917])|(m[1911]&~m[1914]&~m[1915]&m[1916]&m[1917])|(~m[1911]&m[1914]&~m[1915]&m[1916]&m[1917])|(m[1911]&m[1914]&~m[1915]&m[1916]&m[1917])|(~m[1911]&~m[1914]&m[1915]&m[1916]&m[1917])|(m[1911]&~m[1914]&m[1915]&m[1916]&m[1917])|(m[1911]&m[1914]&m[1915]&m[1916]&m[1917]));
    m[1918] = (((m[1916]&~m[1919]&~m[1920]&~m[1921]&~m[1922])|(~m[1916]&~m[1919]&~m[1920]&m[1921]&~m[1922])|(m[1916]&m[1919]&~m[1920]&m[1921]&~m[1922])|(m[1916]&~m[1919]&m[1920]&m[1921]&~m[1922])|(~m[1916]&m[1919]&~m[1920]&~m[1921]&m[1922])|(~m[1916]&~m[1919]&m[1920]&~m[1921]&m[1922])|(m[1916]&m[1919]&m[1920]&~m[1921]&m[1922])|(~m[1916]&m[1919]&m[1920]&m[1921]&m[1922]))&UnbiasedRNG[229])|((m[1916]&~m[1919]&~m[1920]&m[1921]&~m[1922])|(~m[1916]&~m[1919]&~m[1920]&~m[1921]&m[1922])|(m[1916]&~m[1919]&~m[1920]&~m[1921]&m[1922])|(m[1916]&m[1919]&~m[1920]&~m[1921]&m[1922])|(m[1916]&~m[1919]&m[1920]&~m[1921]&m[1922])|(~m[1916]&~m[1919]&~m[1920]&m[1921]&m[1922])|(m[1916]&~m[1919]&~m[1920]&m[1921]&m[1922])|(~m[1916]&m[1919]&~m[1920]&m[1921]&m[1922])|(m[1916]&m[1919]&~m[1920]&m[1921]&m[1922])|(~m[1916]&~m[1919]&m[1920]&m[1921]&m[1922])|(m[1916]&~m[1919]&m[1920]&m[1921]&m[1922])|(m[1916]&m[1919]&m[1920]&m[1921]&m[1922]));
    m[1923] = (((m[1921]&~m[1924]&~m[1925]&~m[1926]&~m[1927])|(~m[1921]&~m[1924]&~m[1925]&m[1926]&~m[1927])|(m[1921]&m[1924]&~m[1925]&m[1926]&~m[1927])|(m[1921]&~m[1924]&m[1925]&m[1926]&~m[1927])|(~m[1921]&m[1924]&~m[1925]&~m[1926]&m[1927])|(~m[1921]&~m[1924]&m[1925]&~m[1926]&m[1927])|(m[1921]&m[1924]&m[1925]&~m[1926]&m[1927])|(~m[1921]&m[1924]&m[1925]&m[1926]&m[1927]))&UnbiasedRNG[230])|((m[1921]&~m[1924]&~m[1925]&m[1926]&~m[1927])|(~m[1921]&~m[1924]&~m[1925]&~m[1926]&m[1927])|(m[1921]&~m[1924]&~m[1925]&~m[1926]&m[1927])|(m[1921]&m[1924]&~m[1925]&~m[1926]&m[1927])|(m[1921]&~m[1924]&m[1925]&~m[1926]&m[1927])|(~m[1921]&~m[1924]&~m[1925]&m[1926]&m[1927])|(m[1921]&~m[1924]&~m[1925]&m[1926]&m[1927])|(~m[1921]&m[1924]&~m[1925]&m[1926]&m[1927])|(m[1921]&m[1924]&~m[1925]&m[1926]&m[1927])|(~m[1921]&~m[1924]&m[1925]&m[1926]&m[1927])|(m[1921]&~m[1924]&m[1925]&m[1926]&m[1927])|(m[1921]&m[1924]&m[1925]&m[1926]&m[1927]));
    m[1928] = (((m[1926]&~m[1929]&~m[1930]&~m[1931]&~m[1932])|(~m[1926]&~m[1929]&~m[1930]&m[1931]&~m[1932])|(m[1926]&m[1929]&~m[1930]&m[1931]&~m[1932])|(m[1926]&~m[1929]&m[1930]&m[1931]&~m[1932])|(~m[1926]&m[1929]&~m[1930]&~m[1931]&m[1932])|(~m[1926]&~m[1929]&m[1930]&~m[1931]&m[1932])|(m[1926]&m[1929]&m[1930]&~m[1931]&m[1932])|(~m[1926]&m[1929]&m[1930]&m[1931]&m[1932]))&UnbiasedRNG[231])|((m[1926]&~m[1929]&~m[1930]&m[1931]&~m[1932])|(~m[1926]&~m[1929]&~m[1930]&~m[1931]&m[1932])|(m[1926]&~m[1929]&~m[1930]&~m[1931]&m[1932])|(m[1926]&m[1929]&~m[1930]&~m[1931]&m[1932])|(m[1926]&~m[1929]&m[1930]&~m[1931]&m[1932])|(~m[1926]&~m[1929]&~m[1930]&m[1931]&m[1932])|(m[1926]&~m[1929]&~m[1930]&m[1931]&m[1932])|(~m[1926]&m[1929]&~m[1930]&m[1931]&m[1932])|(m[1926]&m[1929]&~m[1930]&m[1931]&m[1932])|(~m[1926]&~m[1929]&m[1930]&m[1931]&m[1932])|(m[1926]&~m[1929]&m[1930]&m[1931]&m[1932])|(m[1926]&m[1929]&m[1930]&m[1931]&m[1932]));
    m[1933] = (((m[1931]&~m[1934]&~m[1935]&~m[1936]&~m[1937])|(~m[1931]&~m[1934]&~m[1935]&m[1936]&~m[1937])|(m[1931]&m[1934]&~m[1935]&m[1936]&~m[1937])|(m[1931]&~m[1934]&m[1935]&m[1936]&~m[1937])|(~m[1931]&m[1934]&~m[1935]&~m[1936]&m[1937])|(~m[1931]&~m[1934]&m[1935]&~m[1936]&m[1937])|(m[1931]&m[1934]&m[1935]&~m[1936]&m[1937])|(~m[1931]&m[1934]&m[1935]&m[1936]&m[1937]))&UnbiasedRNG[232])|((m[1931]&~m[1934]&~m[1935]&m[1936]&~m[1937])|(~m[1931]&~m[1934]&~m[1935]&~m[1936]&m[1937])|(m[1931]&~m[1934]&~m[1935]&~m[1936]&m[1937])|(m[1931]&m[1934]&~m[1935]&~m[1936]&m[1937])|(m[1931]&~m[1934]&m[1935]&~m[1936]&m[1937])|(~m[1931]&~m[1934]&~m[1935]&m[1936]&m[1937])|(m[1931]&~m[1934]&~m[1935]&m[1936]&m[1937])|(~m[1931]&m[1934]&~m[1935]&m[1936]&m[1937])|(m[1931]&m[1934]&~m[1935]&m[1936]&m[1937])|(~m[1931]&~m[1934]&m[1935]&m[1936]&m[1937])|(m[1931]&~m[1934]&m[1935]&m[1936]&m[1937])|(m[1931]&m[1934]&m[1935]&m[1936]&m[1937]));
    m[1938] = (((m[1936]&~m[1939]&~m[1940]&~m[1941]&~m[1942])|(~m[1936]&~m[1939]&~m[1940]&m[1941]&~m[1942])|(m[1936]&m[1939]&~m[1940]&m[1941]&~m[1942])|(m[1936]&~m[1939]&m[1940]&m[1941]&~m[1942])|(~m[1936]&m[1939]&~m[1940]&~m[1941]&m[1942])|(~m[1936]&~m[1939]&m[1940]&~m[1941]&m[1942])|(m[1936]&m[1939]&m[1940]&~m[1941]&m[1942])|(~m[1936]&m[1939]&m[1940]&m[1941]&m[1942]))&UnbiasedRNG[233])|((m[1936]&~m[1939]&~m[1940]&m[1941]&~m[1942])|(~m[1936]&~m[1939]&~m[1940]&~m[1941]&m[1942])|(m[1936]&~m[1939]&~m[1940]&~m[1941]&m[1942])|(m[1936]&m[1939]&~m[1940]&~m[1941]&m[1942])|(m[1936]&~m[1939]&m[1940]&~m[1941]&m[1942])|(~m[1936]&~m[1939]&~m[1940]&m[1941]&m[1942])|(m[1936]&~m[1939]&~m[1940]&m[1941]&m[1942])|(~m[1936]&m[1939]&~m[1940]&m[1941]&m[1942])|(m[1936]&m[1939]&~m[1940]&m[1941]&m[1942])|(~m[1936]&~m[1939]&m[1940]&m[1941]&m[1942])|(m[1936]&~m[1939]&m[1940]&m[1941]&m[1942])|(m[1936]&m[1939]&m[1940]&m[1941]&m[1942]));
    m[1943] = (((m[1941]&~m[1944]&~m[1945]&~m[1946]&~m[1947])|(~m[1941]&~m[1944]&~m[1945]&m[1946]&~m[1947])|(m[1941]&m[1944]&~m[1945]&m[1946]&~m[1947])|(m[1941]&~m[1944]&m[1945]&m[1946]&~m[1947])|(~m[1941]&m[1944]&~m[1945]&~m[1946]&m[1947])|(~m[1941]&~m[1944]&m[1945]&~m[1946]&m[1947])|(m[1941]&m[1944]&m[1945]&~m[1946]&m[1947])|(~m[1941]&m[1944]&m[1945]&m[1946]&m[1947]))&UnbiasedRNG[234])|((m[1941]&~m[1944]&~m[1945]&m[1946]&~m[1947])|(~m[1941]&~m[1944]&~m[1945]&~m[1946]&m[1947])|(m[1941]&~m[1944]&~m[1945]&~m[1946]&m[1947])|(m[1941]&m[1944]&~m[1945]&~m[1946]&m[1947])|(m[1941]&~m[1944]&m[1945]&~m[1946]&m[1947])|(~m[1941]&~m[1944]&~m[1945]&m[1946]&m[1947])|(m[1941]&~m[1944]&~m[1945]&m[1946]&m[1947])|(~m[1941]&m[1944]&~m[1945]&m[1946]&m[1947])|(m[1941]&m[1944]&~m[1945]&m[1946]&m[1947])|(~m[1941]&~m[1944]&m[1945]&m[1946]&m[1947])|(m[1941]&~m[1944]&m[1945]&m[1946]&m[1947])|(m[1941]&m[1944]&m[1945]&m[1946]&m[1947]));
    m[1948] = (((m[1907]&~m[1949]&~m[1950]&~m[1951]&~m[1952])|(~m[1907]&~m[1949]&~m[1950]&m[1951]&~m[1952])|(m[1907]&m[1949]&~m[1950]&m[1951]&~m[1952])|(m[1907]&~m[1949]&m[1950]&m[1951]&~m[1952])|(~m[1907]&m[1949]&~m[1950]&~m[1951]&m[1952])|(~m[1907]&~m[1949]&m[1950]&~m[1951]&m[1952])|(m[1907]&m[1949]&m[1950]&~m[1951]&m[1952])|(~m[1907]&m[1949]&m[1950]&m[1951]&m[1952]))&UnbiasedRNG[235])|((m[1907]&~m[1949]&~m[1950]&m[1951]&~m[1952])|(~m[1907]&~m[1949]&~m[1950]&~m[1951]&m[1952])|(m[1907]&~m[1949]&~m[1950]&~m[1951]&m[1952])|(m[1907]&m[1949]&~m[1950]&~m[1951]&m[1952])|(m[1907]&~m[1949]&m[1950]&~m[1951]&m[1952])|(~m[1907]&~m[1949]&~m[1950]&m[1951]&m[1952])|(m[1907]&~m[1949]&~m[1950]&m[1951]&m[1952])|(~m[1907]&m[1949]&~m[1950]&m[1951]&m[1952])|(m[1907]&m[1949]&~m[1950]&m[1951]&m[1952])|(~m[1907]&~m[1949]&m[1950]&m[1951]&m[1952])|(m[1907]&~m[1949]&m[1950]&m[1951]&m[1952])|(m[1907]&m[1949]&m[1950]&m[1951]&m[1952]));
    m[1953] = (((m[1951]&~m[1954]&~m[1955]&~m[1956]&~m[1957])|(~m[1951]&~m[1954]&~m[1955]&m[1956]&~m[1957])|(m[1951]&m[1954]&~m[1955]&m[1956]&~m[1957])|(m[1951]&~m[1954]&m[1955]&m[1956]&~m[1957])|(~m[1951]&m[1954]&~m[1955]&~m[1956]&m[1957])|(~m[1951]&~m[1954]&m[1955]&~m[1956]&m[1957])|(m[1951]&m[1954]&m[1955]&~m[1956]&m[1957])|(~m[1951]&m[1954]&m[1955]&m[1956]&m[1957]))&UnbiasedRNG[236])|((m[1951]&~m[1954]&~m[1955]&m[1956]&~m[1957])|(~m[1951]&~m[1954]&~m[1955]&~m[1956]&m[1957])|(m[1951]&~m[1954]&~m[1955]&~m[1956]&m[1957])|(m[1951]&m[1954]&~m[1955]&~m[1956]&m[1957])|(m[1951]&~m[1954]&m[1955]&~m[1956]&m[1957])|(~m[1951]&~m[1954]&~m[1955]&m[1956]&m[1957])|(m[1951]&~m[1954]&~m[1955]&m[1956]&m[1957])|(~m[1951]&m[1954]&~m[1955]&m[1956]&m[1957])|(m[1951]&m[1954]&~m[1955]&m[1956]&m[1957])|(~m[1951]&~m[1954]&m[1955]&m[1956]&m[1957])|(m[1951]&~m[1954]&m[1955]&m[1956]&m[1957])|(m[1951]&m[1954]&m[1955]&m[1956]&m[1957]));
    m[1958] = (((m[1956]&~m[1959]&~m[1960]&~m[1961]&~m[1962])|(~m[1956]&~m[1959]&~m[1960]&m[1961]&~m[1962])|(m[1956]&m[1959]&~m[1960]&m[1961]&~m[1962])|(m[1956]&~m[1959]&m[1960]&m[1961]&~m[1962])|(~m[1956]&m[1959]&~m[1960]&~m[1961]&m[1962])|(~m[1956]&~m[1959]&m[1960]&~m[1961]&m[1962])|(m[1956]&m[1959]&m[1960]&~m[1961]&m[1962])|(~m[1956]&m[1959]&m[1960]&m[1961]&m[1962]))&UnbiasedRNG[237])|((m[1956]&~m[1959]&~m[1960]&m[1961]&~m[1962])|(~m[1956]&~m[1959]&~m[1960]&~m[1961]&m[1962])|(m[1956]&~m[1959]&~m[1960]&~m[1961]&m[1962])|(m[1956]&m[1959]&~m[1960]&~m[1961]&m[1962])|(m[1956]&~m[1959]&m[1960]&~m[1961]&m[1962])|(~m[1956]&~m[1959]&~m[1960]&m[1961]&m[1962])|(m[1956]&~m[1959]&~m[1960]&m[1961]&m[1962])|(~m[1956]&m[1959]&~m[1960]&m[1961]&m[1962])|(m[1956]&m[1959]&~m[1960]&m[1961]&m[1962])|(~m[1956]&~m[1959]&m[1960]&m[1961]&m[1962])|(m[1956]&~m[1959]&m[1960]&m[1961]&m[1962])|(m[1956]&m[1959]&m[1960]&m[1961]&m[1962]));
    m[1963] = (((m[1961]&~m[1964]&~m[1965]&~m[1966]&~m[1967])|(~m[1961]&~m[1964]&~m[1965]&m[1966]&~m[1967])|(m[1961]&m[1964]&~m[1965]&m[1966]&~m[1967])|(m[1961]&~m[1964]&m[1965]&m[1966]&~m[1967])|(~m[1961]&m[1964]&~m[1965]&~m[1966]&m[1967])|(~m[1961]&~m[1964]&m[1965]&~m[1966]&m[1967])|(m[1961]&m[1964]&m[1965]&~m[1966]&m[1967])|(~m[1961]&m[1964]&m[1965]&m[1966]&m[1967]))&UnbiasedRNG[238])|((m[1961]&~m[1964]&~m[1965]&m[1966]&~m[1967])|(~m[1961]&~m[1964]&~m[1965]&~m[1966]&m[1967])|(m[1961]&~m[1964]&~m[1965]&~m[1966]&m[1967])|(m[1961]&m[1964]&~m[1965]&~m[1966]&m[1967])|(m[1961]&~m[1964]&m[1965]&~m[1966]&m[1967])|(~m[1961]&~m[1964]&~m[1965]&m[1966]&m[1967])|(m[1961]&~m[1964]&~m[1965]&m[1966]&m[1967])|(~m[1961]&m[1964]&~m[1965]&m[1966]&m[1967])|(m[1961]&m[1964]&~m[1965]&m[1966]&m[1967])|(~m[1961]&~m[1964]&m[1965]&m[1966]&m[1967])|(m[1961]&~m[1964]&m[1965]&m[1966]&m[1967])|(m[1961]&m[1964]&m[1965]&m[1966]&m[1967]));
    m[1968] = (((m[1966]&~m[1969]&~m[1970]&~m[1971]&~m[1972])|(~m[1966]&~m[1969]&~m[1970]&m[1971]&~m[1972])|(m[1966]&m[1969]&~m[1970]&m[1971]&~m[1972])|(m[1966]&~m[1969]&m[1970]&m[1971]&~m[1972])|(~m[1966]&m[1969]&~m[1970]&~m[1971]&m[1972])|(~m[1966]&~m[1969]&m[1970]&~m[1971]&m[1972])|(m[1966]&m[1969]&m[1970]&~m[1971]&m[1972])|(~m[1966]&m[1969]&m[1970]&m[1971]&m[1972]))&UnbiasedRNG[239])|((m[1966]&~m[1969]&~m[1970]&m[1971]&~m[1972])|(~m[1966]&~m[1969]&~m[1970]&~m[1971]&m[1972])|(m[1966]&~m[1969]&~m[1970]&~m[1971]&m[1972])|(m[1966]&m[1969]&~m[1970]&~m[1971]&m[1972])|(m[1966]&~m[1969]&m[1970]&~m[1971]&m[1972])|(~m[1966]&~m[1969]&~m[1970]&m[1971]&m[1972])|(m[1966]&~m[1969]&~m[1970]&m[1971]&m[1972])|(~m[1966]&m[1969]&~m[1970]&m[1971]&m[1972])|(m[1966]&m[1969]&~m[1970]&m[1971]&m[1972])|(~m[1966]&~m[1969]&m[1970]&m[1971]&m[1972])|(m[1966]&~m[1969]&m[1970]&m[1971]&m[1972])|(m[1966]&m[1969]&m[1970]&m[1971]&m[1972]));
    m[1973] = (((m[1971]&~m[1974]&~m[1975]&~m[1976]&~m[1977])|(~m[1971]&~m[1974]&~m[1975]&m[1976]&~m[1977])|(m[1971]&m[1974]&~m[1975]&m[1976]&~m[1977])|(m[1971]&~m[1974]&m[1975]&m[1976]&~m[1977])|(~m[1971]&m[1974]&~m[1975]&~m[1976]&m[1977])|(~m[1971]&~m[1974]&m[1975]&~m[1976]&m[1977])|(m[1971]&m[1974]&m[1975]&~m[1976]&m[1977])|(~m[1971]&m[1974]&m[1975]&m[1976]&m[1977]))&UnbiasedRNG[240])|((m[1971]&~m[1974]&~m[1975]&m[1976]&~m[1977])|(~m[1971]&~m[1974]&~m[1975]&~m[1976]&m[1977])|(m[1971]&~m[1974]&~m[1975]&~m[1976]&m[1977])|(m[1971]&m[1974]&~m[1975]&~m[1976]&m[1977])|(m[1971]&~m[1974]&m[1975]&~m[1976]&m[1977])|(~m[1971]&~m[1974]&~m[1975]&m[1976]&m[1977])|(m[1971]&~m[1974]&~m[1975]&m[1976]&m[1977])|(~m[1971]&m[1974]&~m[1975]&m[1976]&m[1977])|(m[1971]&m[1974]&~m[1975]&m[1976]&m[1977])|(~m[1971]&~m[1974]&m[1975]&m[1976]&m[1977])|(m[1971]&~m[1974]&m[1975]&m[1976]&m[1977])|(m[1971]&m[1974]&m[1975]&m[1976]&m[1977]));
    m[1978] = (((m[1976]&~m[1979]&~m[1980]&~m[1981]&~m[1982])|(~m[1976]&~m[1979]&~m[1980]&m[1981]&~m[1982])|(m[1976]&m[1979]&~m[1980]&m[1981]&~m[1982])|(m[1976]&~m[1979]&m[1980]&m[1981]&~m[1982])|(~m[1976]&m[1979]&~m[1980]&~m[1981]&m[1982])|(~m[1976]&~m[1979]&m[1980]&~m[1981]&m[1982])|(m[1976]&m[1979]&m[1980]&~m[1981]&m[1982])|(~m[1976]&m[1979]&m[1980]&m[1981]&m[1982]))&UnbiasedRNG[241])|((m[1976]&~m[1979]&~m[1980]&m[1981]&~m[1982])|(~m[1976]&~m[1979]&~m[1980]&~m[1981]&m[1982])|(m[1976]&~m[1979]&~m[1980]&~m[1981]&m[1982])|(m[1976]&m[1979]&~m[1980]&~m[1981]&m[1982])|(m[1976]&~m[1979]&m[1980]&~m[1981]&m[1982])|(~m[1976]&~m[1979]&~m[1980]&m[1981]&m[1982])|(m[1976]&~m[1979]&~m[1980]&m[1981]&m[1982])|(~m[1976]&m[1979]&~m[1980]&m[1981]&m[1982])|(m[1976]&m[1979]&~m[1980]&m[1981]&m[1982])|(~m[1976]&~m[1979]&m[1980]&m[1981]&m[1982])|(m[1976]&~m[1979]&m[1980]&m[1981]&m[1982])|(m[1976]&m[1979]&m[1980]&m[1981]&m[1982]));
    m[1983] = (((m[1981]&~m[1984]&~m[1985]&~m[1986]&~m[1987])|(~m[1981]&~m[1984]&~m[1985]&m[1986]&~m[1987])|(m[1981]&m[1984]&~m[1985]&m[1986]&~m[1987])|(m[1981]&~m[1984]&m[1985]&m[1986]&~m[1987])|(~m[1981]&m[1984]&~m[1985]&~m[1986]&m[1987])|(~m[1981]&~m[1984]&m[1985]&~m[1986]&m[1987])|(m[1981]&m[1984]&m[1985]&~m[1986]&m[1987])|(~m[1981]&m[1984]&m[1985]&m[1986]&m[1987]))&UnbiasedRNG[242])|((m[1981]&~m[1984]&~m[1985]&m[1986]&~m[1987])|(~m[1981]&~m[1984]&~m[1985]&~m[1986]&m[1987])|(m[1981]&~m[1984]&~m[1985]&~m[1986]&m[1987])|(m[1981]&m[1984]&~m[1985]&~m[1986]&m[1987])|(m[1981]&~m[1984]&m[1985]&~m[1986]&m[1987])|(~m[1981]&~m[1984]&~m[1985]&m[1986]&m[1987])|(m[1981]&~m[1984]&~m[1985]&m[1986]&m[1987])|(~m[1981]&m[1984]&~m[1985]&m[1986]&m[1987])|(m[1981]&m[1984]&~m[1985]&m[1986]&m[1987])|(~m[1981]&~m[1984]&m[1985]&m[1986]&m[1987])|(m[1981]&~m[1984]&m[1985]&m[1986]&m[1987])|(m[1981]&m[1984]&m[1985]&m[1986]&m[1987]));
    m[1988] = (((m[1952]&~m[1989]&~m[1990]&~m[1991]&~m[1992])|(~m[1952]&~m[1989]&~m[1990]&m[1991]&~m[1992])|(m[1952]&m[1989]&~m[1990]&m[1991]&~m[1992])|(m[1952]&~m[1989]&m[1990]&m[1991]&~m[1992])|(~m[1952]&m[1989]&~m[1990]&~m[1991]&m[1992])|(~m[1952]&~m[1989]&m[1990]&~m[1991]&m[1992])|(m[1952]&m[1989]&m[1990]&~m[1991]&m[1992])|(~m[1952]&m[1989]&m[1990]&m[1991]&m[1992]))&UnbiasedRNG[243])|((m[1952]&~m[1989]&~m[1990]&m[1991]&~m[1992])|(~m[1952]&~m[1989]&~m[1990]&~m[1991]&m[1992])|(m[1952]&~m[1989]&~m[1990]&~m[1991]&m[1992])|(m[1952]&m[1989]&~m[1990]&~m[1991]&m[1992])|(m[1952]&~m[1989]&m[1990]&~m[1991]&m[1992])|(~m[1952]&~m[1989]&~m[1990]&m[1991]&m[1992])|(m[1952]&~m[1989]&~m[1990]&m[1991]&m[1992])|(~m[1952]&m[1989]&~m[1990]&m[1991]&m[1992])|(m[1952]&m[1989]&~m[1990]&m[1991]&m[1992])|(~m[1952]&~m[1989]&m[1990]&m[1991]&m[1992])|(m[1952]&~m[1989]&m[1990]&m[1991]&m[1992])|(m[1952]&m[1989]&m[1990]&m[1991]&m[1992]));
    m[1993] = (((m[1991]&~m[1994]&~m[1995]&~m[1996]&~m[1997])|(~m[1991]&~m[1994]&~m[1995]&m[1996]&~m[1997])|(m[1991]&m[1994]&~m[1995]&m[1996]&~m[1997])|(m[1991]&~m[1994]&m[1995]&m[1996]&~m[1997])|(~m[1991]&m[1994]&~m[1995]&~m[1996]&m[1997])|(~m[1991]&~m[1994]&m[1995]&~m[1996]&m[1997])|(m[1991]&m[1994]&m[1995]&~m[1996]&m[1997])|(~m[1991]&m[1994]&m[1995]&m[1996]&m[1997]))&UnbiasedRNG[244])|((m[1991]&~m[1994]&~m[1995]&m[1996]&~m[1997])|(~m[1991]&~m[1994]&~m[1995]&~m[1996]&m[1997])|(m[1991]&~m[1994]&~m[1995]&~m[1996]&m[1997])|(m[1991]&m[1994]&~m[1995]&~m[1996]&m[1997])|(m[1991]&~m[1994]&m[1995]&~m[1996]&m[1997])|(~m[1991]&~m[1994]&~m[1995]&m[1996]&m[1997])|(m[1991]&~m[1994]&~m[1995]&m[1996]&m[1997])|(~m[1991]&m[1994]&~m[1995]&m[1996]&m[1997])|(m[1991]&m[1994]&~m[1995]&m[1996]&m[1997])|(~m[1991]&~m[1994]&m[1995]&m[1996]&m[1997])|(m[1991]&~m[1994]&m[1995]&m[1996]&m[1997])|(m[1991]&m[1994]&m[1995]&m[1996]&m[1997]));
    m[1998] = (((m[1996]&~m[1999]&~m[2000]&~m[2001]&~m[2002])|(~m[1996]&~m[1999]&~m[2000]&m[2001]&~m[2002])|(m[1996]&m[1999]&~m[2000]&m[2001]&~m[2002])|(m[1996]&~m[1999]&m[2000]&m[2001]&~m[2002])|(~m[1996]&m[1999]&~m[2000]&~m[2001]&m[2002])|(~m[1996]&~m[1999]&m[2000]&~m[2001]&m[2002])|(m[1996]&m[1999]&m[2000]&~m[2001]&m[2002])|(~m[1996]&m[1999]&m[2000]&m[2001]&m[2002]))&UnbiasedRNG[245])|((m[1996]&~m[1999]&~m[2000]&m[2001]&~m[2002])|(~m[1996]&~m[1999]&~m[2000]&~m[2001]&m[2002])|(m[1996]&~m[1999]&~m[2000]&~m[2001]&m[2002])|(m[1996]&m[1999]&~m[2000]&~m[2001]&m[2002])|(m[1996]&~m[1999]&m[2000]&~m[2001]&m[2002])|(~m[1996]&~m[1999]&~m[2000]&m[2001]&m[2002])|(m[1996]&~m[1999]&~m[2000]&m[2001]&m[2002])|(~m[1996]&m[1999]&~m[2000]&m[2001]&m[2002])|(m[1996]&m[1999]&~m[2000]&m[2001]&m[2002])|(~m[1996]&~m[1999]&m[2000]&m[2001]&m[2002])|(m[1996]&~m[1999]&m[2000]&m[2001]&m[2002])|(m[1996]&m[1999]&m[2000]&m[2001]&m[2002]));
    m[2003] = (((m[2001]&~m[2004]&~m[2005]&~m[2006]&~m[2007])|(~m[2001]&~m[2004]&~m[2005]&m[2006]&~m[2007])|(m[2001]&m[2004]&~m[2005]&m[2006]&~m[2007])|(m[2001]&~m[2004]&m[2005]&m[2006]&~m[2007])|(~m[2001]&m[2004]&~m[2005]&~m[2006]&m[2007])|(~m[2001]&~m[2004]&m[2005]&~m[2006]&m[2007])|(m[2001]&m[2004]&m[2005]&~m[2006]&m[2007])|(~m[2001]&m[2004]&m[2005]&m[2006]&m[2007]))&UnbiasedRNG[246])|((m[2001]&~m[2004]&~m[2005]&m[2006]&~m[2007])|(~m[2001]&~m[2004]&~m[2005]&~m[2006]&m[2007])|(m[2001]&~m[2004]&~m[2005]&~m[2006]&m[2007])|(m[2001]&m[2004]&~m[2005]&~m[2006]&m[2007])|(m[2001]&~m[2004]&m[2005]&~m[2006]&m[2007])|(~m[2001]&~m[2004]&~m[2005]&m[2006]&m[2007])|(m[2001]&~m[2004]&~m[2005]&m[2006]&m[2007])|(~m[2001]&m[2004]&~m[2005]&m[2006]&m[2007])|(m[2001]&m[2004]&~m[2005]&m[2006]&m[2007])|(~m[2001]&~m[2004]&m[2005]&m[2006]&m[2007])|(m[2001]&~m[2004]&m[2005]&m[2006]&m[2007])|(m[2001]&m[2004]&m[2005]&m[2006]&m[2007]));
    m[2008] = (((m[2006]&~m[2009]&~m[2010]&~m[2011]&~m[2012])|(~m[2006]&~m[2009]&~m[2010]&m[2011]&~m[2012])|(m[2006]&m[2009]&~m[2010]&m[2011]&~m[2012])|(m[2006]&~m[2009]&m[2010]&m[2011]&~m[2012])|(~m[2006]&m[2009]&~m[2010]&~m[2011]&m[2012])|(~m[2006]&~m[2009]&m[2010]&~m[2011]&m[2012])|(m[2006]&m[2009]&m[2010]&~m[2011]&m[2012])|(~m[2006]&m[2009]&m[2010]&m[2011]&m[2012]))&UnbiasedRNG[247])|((m[2006]&~m[2009]&~m[2010]&m[2011]&~m[2012])|(~m[2006]&~m[2009]&~m[2010]&~m[2011]&m[2012])|(m[2006]&~m[2009]&~m[2010]&~m[2011]&m[2012])|(m[2006]&m[2009]&~m[2010]&~m[2011]&m[2012])|(m[2006]&~m[2009]&m[2010]&~m[2011]&m[2012])|(~m[2006]&~m[2009]&~m[2010]&m[2011]&m[2012])|(m[2006]&~m[2009]&~m[2010]&m[2011]&m[2012])|(~m[2006]&m[2009]&~m[2010]&m[2011]&m[2012])|(m[2006]&m[2009]&~m[2010]&m[2011]&m[2012])|(~m[2006]&~m[2009]&m[2010]&m[2011]&m[2012])|(m[2006]&~m[2009]&m[2010]&m[2011]&m[2012])|(m[2006]&m[2009]&m[2010]&m[2011]&m[2012]));
    m[2013] = (((m[2011]&~m[2014]&~m[2015]&~m[2016]&~m[2017])|(~m[2011]&~m[2014]&~m[2015]&m[2016]&~m[2017])|(m[2011]&m[2014]&~m[2015]&m[2016]&~m[2017])|(m[2011]&~m[2014]&m[2015]&m[2016]&~m[2017])|(~m[2011]&m[2014]&~m[2015]&~m[2016]&m[2017])|(~m[2011]&~m[2014]&m[2015]&~m[2016]&m[2017])|(m[2011]&m[2014]&m[2015]&~m[2016]&m[2017])|(~m[2011]&m[2014]&m[2015]&m[2016]&m[2017]))&UnbiasedRNG[248])|((m[2011]&~m[2014]&~m[2015]&m[2016]&~m[2017])|(~m[2011]&~m[2014]&~m[2015]&~m[2016]&m[2017])|(m[2011]&~m[2014]&~m[2015]&~m[2016]&m[2017])|(m[2011]&m[2014]&~m[2015]&~m[2016]&m[2017])|(m[2011]&~m[2014]&m[2015]&~m[2016]&m[2017])|(~m[2011]&~m[2014]&~m[2015]&m[2016]&m[2017])|(m[2011]&~m[2014]&~m[2015]&m[2016]&m[2017])|(~m[2011]&m[2014]&~m[2015]&m[2016]&m[2017])|(m[2011]&m[2014]&~m[2015]&m[2016]&m[2017])|(~m[2011]&~m[2014]&m[2015]&m[2016]&m[2017])|(m[2011]&~m[2014]&m[2015]&m[2016]&m[2017])|(m[2011]&m[2014]&m[2015]&m[2016]&m[2017]));
    m[2018] = (((m[2016]&~m[2019]&~m[2020]&~m[2021]&~m[2022])|(~m[2016]&~m[2019]&~m[2020]&m[2021]&~m[2022])|(m[2016]&m[2019]&~m[2020]&m[2021]&~m[2022])|(m[2016]&~m[2019]&m[2020]&m[2021]&~m[2022])|(~m[2016]&m[2019]&~m[2020]&~m[2021]&m[2022])|(~m[2016]&~m[2019]&m[2020]&~m[2021]&m[2022])|(m[2016]&m[2019]&m[2020]&~m[2021]&m[2022])|(~m[2016]&m[2019]&m[2020]&m[2021]&m[2022]))&UnbiasedRNG[249])|((m[2016]&~m[2019]&~m[2020]&m[2021]&~m[2022])|(~m[2016]&~m[2019]&~m[2020]&~m[2021]&m[2022])|(m[2016]&~m[2019]&~m[2020]&~m[2021]&m[2022])|(m[2016]&m[2019]&~m[2020]&~m[2021]&m[2022])|(m[2016]&~m[2019]&m[2020]&~m[2021]&m[2022])|(~m[2016]&~m[2019]&~m[2020]&m[2021]&m[2022])|(m[2016]&~m[2019]&~m[2020]&m[2021]&m[2022])|(~m[2016]&m[2019]&~m[2020]&m[2021]&m[2022])|(m[2016]&m[2019]&~m[2020]&m[2021]&m[2022])|(~m[2016]&~m[2019]&m[2020]&m[2021]&m[2022])|(m[2016]&~m[2019]&m[2020]&m[2021]&m[2022])|(m[2016]&m[2019]&m[2020]&m[2021]&m[2022]));
    m[2023] = (((m[1992]&~m[2024]&~m[2025]&~m[2026]&~m[2027])|(~m[1992]&~m[2024]&~m[2025]&m[2026]&~m[2027])|(m[1992]&m[2024]&~m[2025]&m[2026]&~m[2027])|(m[1992]&~m[2024]&m[2025]&m[2026]&~m[2027])|(~m[1992]&m[2024]&~m[2025]&~m[2026]&m[2027])|(~m[1992]&~m[2024]&m[2025]&~m[2026]&m[2027])|(m[1992]&m[2024]&m[2025]&~m[2026]&m[2027])|(~m[1992]&m[2024]&m[2025]&m[2026]&m[2027]))&UnbiasedRNG[250])|((m[1992]&~m[2024]&~m[2025]&m[2026]&~m[2027])|(~m[1992]&~m[2024]&~m[2025]&~m[2026]&m[2027])|(m[1992]&~m[2024]&~m[2025]&~m[2026]&m[2027])|(m[1992]&m[2024]&~m[2025]&~m[2026]&m[2027])|(m[1992]&~m[2024]&m[2025]&~m[2026]&m[2027])|(~m[1992]&~m[2024]&~m[2025]&m[2026]&m[2027])|(m[1992]&~m[2024]&~m[2025]&m[2026]&m[2027])|(~m[1992]&m[2024]&~m[2025]&m[2026]&m[2027])|(m[1992]&m[2024]&~m[2025]&m[2026]&m[2027])|(~m[1992]&~m[2024]&m[2025]&m[2026]&m[2027])|(m[1992]&~m[2024]&m[2025]&m[2026]&m[2027])|(m[1992]&m[2024]&m[2025]&m[2026]&m[2027]));
    m[2028] = (((m[2026]&~m[2029]&~m[2030]&~m[2031]&~m[2032])|(~m[2026]&~m[2029]&~m[2030]&m[2031]&~m[2032])|(m[2026]&m[2029]&~m[2030]&m[2031]&~m[2032])|(m[2026]&~m[2029]&m[2030]&m[2031]&~m[2032])|(~m[2026]&m[2029]&~m[2030]&~m[2031]&m[2032])|(~m[2026]&~m[2029]&m[2030]&~m[2031]&m[2032])|(m[2026]&m[2029]&m[2030]&~m[2031]&m[2032])|(~m[2026]&m[2029]&m[2030]&m[2031]&m[2032]))&UnbiasedRNG[251])|((m[2026]&~m[2029]&~m[2030]&m[2031]&~m[2032])|(~m[2026]&~m[2029]&~m[2030]&~m[2031]&m[2032])|(m[2026]&~m[2029]&~m[2030]&~m[2031]&m[2032])|(m[2026]&m[2029]&~m[2030]&~m[2031]&m[2032])|(m[2026]&~m[2029]&m[2030]&~m[2031]&m[2032])|(~m[2026]&~m[2029]&~m[2030]&m[2031]&m[2032])|(m[2026]&~m[2029]&~m[2030]&m[2031]&m[2032])|(~m[2026]&m[2029]&~m[2030]&m[2031]&m[2032])|(m[2026]&m[2029]&~m[2030]&m[2031]&m[2032])|(~m[2026]&~m[2029]&m[2030]&m[2031]&m[2032])|(m[2026]&~m[2029]&m[2030]&m[2031]&m[2032])|(m[2026]&m[2029]&m[2030]&m[2031]&m[2032]));
    m[2033] = (((m[2031]&~m[2034]&~m[2035]&~m[2036]&~m[2037])|(~m[2031]&~m[2034]&~m[2035]&m[2036]&~m[2037])|(m[2031]&m[2034]&~m[2035]&m[2036]&~m[2037])|(m[2031]&~m[2034]&m[2035]&m[2036]&~m[2037])|(~m[2031]&m[2034]&~m[2035]&~m[2036]&m[2037])|(~m[2031]&~m[2034]&m[2035]&~m[2036]&m[2037])|(m[2031]&m[2034]&m[2035]&~m[2036]&m[2037])|(~m[2031]&m[2034]&m[2035]&m[2036]&m[2037]))&UnbiasedRNG[252])|((m[2031]&~m[2034]&~m[2035]&m[2036]&~m[2037])|(~m[2031]&~m[2034]&~m[2035]&~m[2036]&m[2037])|(m[2031]&~m[2034]&~m[2035]&~m[2036]&m[2037])|(m[2031]&m[2034]&~m[2035]&~m[2036]&m[2037])|(m[2031]&~m[2034]&m[2035]&~m[2036]&m[2037])|(~m[2031]&~m[2034]&~m[2035]&m[2036]&m[2037])|(m[2031]&~m[2034]&~m[2035]&m[2036]&m[2037])|(~m[2031]&m[2034]&~m[2035]&m[2036]&m[2037])|(m[2031]&m[2034]&~m[2035]&m[2036]&m[2037])|(~m[2031]&~m[2034]&m[2035]&m[2036]&m[2037])|(m[2031]&~m[2034]&m[2035]&m[2036]&m[2037])|(m[2031]&m[2034]&m[2035]&m[2036]&m[2037]));
    m[2038] = (((m[2036]&~m[2039]&~m[2040]&~m[2041]&~m[2042])|(~m[2036]&~m[2039]&~m[2040]&m[2041]&~m[2042])|(m[2036]&m[2039]&~m[2040]&m[2041]&~m[2042])|(m[2036]&~m[2039]&m[2040]&m[2041]&~m[2042])|(~m[2036]&m[2039]&~m[2040]&~m[2041]&m[2042])|(~m[2036]&~m[2039]&m[2040]&~m[2041]&m[2042])|(m[2036]&m[2039]&m[2040]&~m[2041]&m[2042])|(~m[2036]&m[2039]&m[2040]&m[2041]&m[2042]))&UnbiasedRNG[253])|((m[2036]&~m[2039]&~m[2040]&m[2041]&~m[2042])|(~m[2036]&~m[2039]&~m[2040]&~m[2041]&m[2042])|(m[2036]&~m[2039]&~m[2040]&~m[2041]&m[2042])|(m[2036]&m[2039]&~m[2040]&~m[2041]&m[2042])|(m[2036]&~m[2039]&m[2040]&~m[2041]&m[2042])|(~m[2036]&~m[2039]&~m[2040]&m[2041]&m[2042])|(m[2036]&~m[2039]&~m[2040]&m[2041]&m[2042])|(~m[2036]&m[2039]&~m[2040]&m[2041]&m[2042])|(m[2036]&m[2039]&~m[2040]&m[2041]&m[2042])|(~m[2036]&~m[2039]&m[2040]&m[2041]&m[2042])|(m[2036]&~m[2039]&m[2040]&m[2041]&m[2042])|(m[2036]&m[2039]&m[2040]&m[2041]&m[2042]));
    m[2043] = (((m[2041]&~m[2044]&~m[2045]&~m[2046]&~m[2047])|(~m[2041]&~m[2044]&~m[2045]&m[2046]&~m[2047])|(m[2041]&m[2044]&~m[2045]&m[2046]&~m[2047])|(m[2041]&~m[2044]&m[2045]&m[2046]&~m[2047])|(~m[2041]&m[2044]&~m[2045]&~m[2046]&m[2047])|(~m[2041]&~m[2044]&m[2045]&~m[2046]&m[2047])|(m[2041]&m[2044]&m[2045]&~m[2046]&m[2047])|(~m[2041]&m[2044]&m[2045]&m[2046]&m[2047]))&UnbiasedRNG[254])|((m[2041]&~m[2044]&~m[2045]&m[2046]&~m[2047])|(~m[2041]&~m[2044]&~m[2045]&~m[2046]&m[2047])|(m[2041]&~m[2044]&~m[2045]&~m[2046]&m[2047])|(m[2041]&m[2044]&~m[2045]&~m[2046]&m[2047])|(m[2041]&~m[2044]&m[2045]&~m[2046]&m[2047])|(~m[2041]&~m[2044]&~m[2045]&m[2046]&m[2047])|(m[2041]&~m[2044]&~m[2045]&m[2046]&m[2047])|(~m[2041]&m[2044]&~m[2045]&m[2046]&m[2047])|(m[2041]&m[2044]&~m[2045]&m[2046]&m[2047])|(~m[2041]&~m[2044]&m[2045]&m[2046]&m[2047])|(m[2041]&~m[2044]&m[2045]&m[2046]&m[2047])|(m[2041]&m[2044]&m[2045]&m[2046]&m[2047]));
    m[2048] = (((m[2046]&~m[2049]&~m[2050]&~m[2051]&~m[2052])|(~m[2046]&~m[2049]&~m[2050]&m[2051]&~m[2052])|(m[2046]&m[2049]&~m[2050]&m[2051]&~m[2052])|(m[2046]&~m[2049]&m[2050]&m[2051]&~m[2052])|(~m[2046]&m[2049]&~m[2050]&~m[2051]&m[2052])|(~m[2046]&~m[2049]&m[2050]&~m[2051]&m[2052])|(m[2046]&m[2049]&m[2050]&~m[2051]&m[2052])|(~m[2046]&m[2049]&m[2050]&m[2051]&m[2052]))&UnbiasedRNG[255])|((m[2046]&~m[2049]&~m[2050]&m[2051]&~m[2052])|(~m[2046]&~m[2049]&~m[2050]&~m[2051]&m[2052])|(m[2046]&~m[2049]&~m[2050]&~m[2051]&m[2052])|(m[2046]&m[2049]&~m[2050]&~m[2051]&m[2052])|(m[2046]&~m[2049]&m[2050]&~m[2051]&m[2052])|(~m[2046]&~m[2049]&~m[2050]&m[2051]&m[2052])|(m[2046]&~m[2049]&~m[2050]&m[2051]&m[2052])|(~m[2046]&m[2049]&~m[2050]&m[2051]&m[2052])|(m[2046]&m[2049]&~m[2050]&m[2051]&m[2052])|(~m[2046]&~m[2049]&m[2050]&m[2051]&m[2052])|(m[2046]&~m[2049]&m[2050]&m[2051]&m[2052])|(m[2046]&m[2049]&m[2050]&m[2051]&m[2052]));
    m[2053] = (((m[2027]&~m[2054]&~m[2055]&~m[2056]&~m[2057])|(~m[2027]&~m[2054]&~m[2055]&m[2056]&~m[2057])|(m[2027]&m[2054]&~m[2055]&m[2056]&~m[2057])|(m[2027]&~m[2054]&m[2055]&m[2056]&~m[2057])|(~m[2027]&m[2054]&~m[2055]&~m[2056]&m[2057])|(~m[2027]&~m[2054]&m[2055]&~m[2056]&m[2057])|(m[2027]&m[2054]&m[2055]&~m[2056]&m[2057])|(~m[2027]&m[2054]&m[2055]&m[2056]&m[2057]))&UnbiasedRNG[256])|((m[2027]&~m[2054]&~m[2055]&m[2056]&~m[2057])|(~m[2027]&~m[2054]&~m[2055]&~m[2056]&m[2057])|(m[2027]&~m[2054]&~m[2055]&~m[2056]&m[2057])|(m[2027]&m[2054]&~m[2055]&~m[2056]&m[2057])|(m[2027]&~m[2054]&m[2055]&~m[2056]&m[2057])|(~m[2027]&~m[2054]&~m[2055]&m[2056]&m[2057])|(m[2027]&~m[2054]&~m[2055]&m[2056]&m[2057])|(~m[2027]&m[2054]&~m[2055]&m[2056]&m[2057])|(m[2027]&m[2054]&~m[2055]&m[2056]&m[2057])|(~m[2027]&~m[2054]&m[2055]&m[2056]&m[2057])|(m[2027]&~m[2054]&m[2055]&m[2056]&m[2057])|(m[2027]&m[2054]&m[2055]&m[2056]&m[2057]));
    m[2058] = (((m[2056]&~m[2059]&~m[2060]&~m[2061]&~m[2062])|(~m[2056]&~m[2059]&~m[2060]&m[2061]&~m[2062])|(m[2056]&m[2059]&~m[2060]&m[2061]&~m[2062])|(m[2056]&~m[2059]&m[2060]&m[2061]&~m[2062])|(~m[2056]&m[2059]&~m[2060]&~m[2061]&m[2062])|(~m[2056]&~m[2059]&m[2060]&~m[2061]&m[2062])|(m[2056]&m[2059]&m[2060]&~m[2061]&m[2062])|(~m[2056]&m[2059]&m[2060]&m[2061]&m[2062]))&UnbiasedRNG[257])|((m[2056]&~m[2059]&~m[2060]&m[2061]&~m[2062])|(~m[2056]&~m[2059]&~m[2060]&~m[2061]&m[2062])|(m[2056]&~m[2059]&~m[2060]&~m[2061]&m[2062])|(m[2056]&m[2059]&~m[2060]&~m[2061]&m[2062])|(m[2056]&~m[2059]&m[2060]&~m[2061]&m[2062])|(~m[2056]&~m[2059]&~m[2060]&m[2061]&m[2062])|(m[2056]&~m[2059]&~m[2060]&m[2061]&m[2062])|(~m[2056]&m[2059]&~m[2060]&m[2061]&m[2062])|(m[2056]&m[2059]&~m[2060]&m[2061]&m[2062])|(~m[2056]&~m[2059]&m[2060]&m[2061]&m[2062])|(m[2056]&~m[2059]&m[2060]&m[2061]&m[2062])|(m[2056]&m[2059]&m[2060]&m[2061]&m[2062]));
    m[2063] = (((m[2061]&~m[2064]&~m[2065]&~m[2066]&~m[2067])|(~m[2061]&~m[2064]&~m[2065]&m[2066]&~m[2067])|(m[2061]&m[2064]&~m[2065]&m[2066]&~m[2067])|(m[2061]&~m[2064]&m[2065]&m[2066]&~m[2067])|(~m[2061]&m[2064]&~m[2065]&~m[2066]&m[2067])|(~m[2061]&~m[2064]&m[2065]&~m[2066]&m[2067])|(m[2061]&m[2064]&m[2065]&~m[2066]&m[2067])|(~m[2061]&m[2064]&m[2065]&m[2066]&m[2067]))&UnbiasedRNG[258])|((m[2061]&~m[2064]&~m[2065]&m[2066]&~m[2067])|(~m[2061]&~m[2064]&~m[2065]&~m[2066]&m[2067])|(m[2061]&~m[2064]&~m[2065]&~m[2066]&m[2067])|(m[2061]&m[2064]&~m[2065]&~m[2066]&m[2067])|(m[2061]&~m[2064]&m[2065]&~m[2066]&m[2067])|(~m[2061]&~m[2064]&~m[2065]&m[2066]&m[2067])|(m[2061]&~m[2064]&~m[2065]&m[2066]&m[2067])|(~m[2061]&m[2064]&~m[2065]&m[2066]&m[2067])|(m[2061]&m[2064]&~m[2065]&m[2066]&m[2067])|(~m[2061]&~m[2064]&m[2065]&m[2066]&m[2067])|(m[2061]&~m[2064]&m[2065]&m[2066]&m[2067])|(m[2061]&m[2064]&m[2065]&m[2066]&m[2067]));
    m[2068] = (((m[2066]&~m[2069]&~m[2070]&~m[2071]&~m[2072])|(~m[2066]&~m[2069]&~m[2070]&m[2071]&~m[2072])|(m[2066]&m[2069]&~m[2070]&m[2071]&~m[2072])|(m[2066]&~m[2069]&m[2070]&m[2071]&~m[2072])|(~m[2066]&m[2069]&~m[2070]&~m[2071]&m[2072])|(~m[2066]&~m[2069]&m[2070]&~m[2071]&m[2072])|(m[2066]&m[2069]&m[2070]&~m[2071]&m[2072])|(~m[2066]&m[2069]&m[2070]&m[2071]&m[2072]))&UnbiasedRNG[259])|((m[2066]&~m[2069]&~m[2070]&m[2071]&~m[2072])|(~m[2066]&~m[2069]&~m[2070]&~m[2071]&m[2072])|(m[2066]&~m[2069]&~m[2070]&~m[2071]&m[2072])|(m[2066]&m[2069]&~m[2070]&~m[2071]&m[2072])|(m[2066]&~m[2069]&m[2070]&~m[2071]&m[2072])|(~m[2066]&~m[2069]&~m[2070]&m[2071]&m[2072])|(m[2066]&~m[2069]&~m[2070]&m[2071]&m[2072])|(~m[2066]&m[2069]&~m[2070]&m[2071]&m[2072])|(m[2066]&m[2069]&~m[2070]&m[2071]&m[2072])|(~m[2066]&~m[2069]&m[2070]&m[2071]&m[2072])|(m[2066]&~m[2069]&m[2070]&m[2071]&m[2072])|(m[2066]&m[2069]&m[2070]&m[2071]&m[2072]));
    m[2073] = (((m[2071]&~m[2074]&~m[2075]&~m[2076]&~m[2077])|(~m[2071]&~m[2074]&~m[2075]&m[2076]&~m[2077])|(m[2071]&m[2074]&~m[2075]&m[2076]&~m[2077])|(m[2071]&~m[2074]&m[2075]&m[2076]&~m[2077])|(~m[2071]&m[2074]&~m[2075]&~m[2076]&m[2077])|(~m[2071]&~m[2074]&m[2075]&~m[2076]&m[2077])|(m[2071]&m[2074]&m[2075]&~m[2076]&m[2077])|(~m[2071]&m[2074]&m[2075]&m[2076]&m[2077]))&UnbiasedRNG[260])|((m[2071]&~m[2074]&~m[2075]&m[2076]&~m[2077])|(~m[2071]&~m[2074]&~m[2075]&~m[2076]&m[2077])|(m[2071]&~m[2074]&~m[2075]&~m[2076]&m[2077])|(m[2071]&m[2074]&~m[2075]&~m[2076]&m[2077])|(m[2071]&~m[2074]&m[2075]&~m[2076]&m[2077])|(~m[2071]&~m[2074]&~m[2075]&m[2076]&m[2077])|(m[2071]&~m[2074]&~m[2075]&m[2076]&m[2077])|(~m[2071]&m[2074]&~m[2075]&m[2076]&m[2077])|(m[2071]&m[2074]&~m[2075]&m[2076]&m[2077])|(~m[2071]&~m[2074]&m[2075]&m[2076]&m[2077])|(m[2071]&~m[2074]&m[2075]&m[2076]&m[2077])|(m[2071]&m[2074]&m[2075]&m[2076]&m[2077]));
    m[2078] = (((m[2057]&~m[2079]&~m[2080]&~m[2081]&~m[2082])|(~m[2057]&~m[2079]&~m[2080]&m[2081]&~m[2082])|(m[2057]&m[2079]&~m[2080]&m[2081]&~m[2082])|(m[2057]&~m[2079]&m[2080]&m[2081]&~m[2082])|(~m[2057]&m[2079]&~m[2080]&~m[2081]&m[2082])|(~m[2057]&~m[2079]&m[2080]&~m[2081]&m[2082])|(m[2057]&m[2079]&m[2080]&~m[2081]&m[2082])|(~m[2057]&m[2079]&m[2080]&m[2081]&m[2082]))&UnbiasedRNG[261])|((m[2057]&~m[2079]&~m[2080]&m[2081]&~m[2082])|(~m[2057]&~m[2079]&~m[2080]&~m[2081]&m[2082])|(m[2057]&~m[2079]&~m[2080]&~m[2081]&m[2082])|(m[2057]&m[2079]&~m[2080]&~m[2081]&m[2082])|(m[2057]&~m[2079]&m[2080]&~m[2081]&m[2082])|(~m[2057]&~m[2079]&~m[2080]&m[2081]&m[2082])|(m[2057]&~m[2079]&~m[2080]&m[2081]&m[2082])|(~m[2057]&m[2079]&~m[2080]&m[2081]&m[2082])|(m[2057]&m[2079]&~m[2080]&m[2081]&m[2082])|(~m[2057]&~m[2079]&m[2080]&m[2081]&m[2082])|(m[2057]&~m[2079]&m[2080]&m[2081]&m[2082])|(m[2057]&m[2079]&m[2080]&m[2081]&m[2082]));
    m[2083] = (((m[2081]&~m[2084]&~m[2085]&~m[2086]&~m[2087])|(~m[2081]&~m[2084]&~m[2085]&m[2086]&~m[2087])|(m[2081]&m[2084]&~m[2085]&m[2086]&~m[2087])|(m[2081]&~m[2084]&m[2085]&m[2086]&~m[2087])|(~m[2081]&m[2084]&~m[2085]&~m[2086]&m[2087])|(~m[2081]&~m[2084]&m[2085]&~m[2086]&m[2087])|(m[2081]&m[2084]&m[2085]&~m[2086]&m[2087])|(~m[2081]&m[2084]&m[2085]&m[2086]&m[2087]))&UnbiasedRNG[262])|((m[2081]&~m[2084]&~m[2085]&m[2086]&~m[2087])|(~m[2081]&~m[2084]&~m[2085]&~m[2086]&m[2087])|(m[2081]&~m[2084]&~m[2085]&~m[2086]&m[2087])|(m[2081]&m[2084]&~m[2085]&~m[2086]&m[2087])|(m[2081]&~m[2084]&m[2085]&~m[2086]&m[2087])|(~m[2081]&~m[2084]&~m[2085]&m[2086]&m[2087])|(m[2081]&~m[2084]&~m[2085]&m[2086]&m[2087])|(~m[2081]&m[2084]&~m[2085]&m[2086]&m[2087])|(m[2081]&m[2084]&~m[2085]&m[2086]&m[2087])|(~m[2081]&~m[2084]&m[2085]&m[2086]&m[2087])|(m[2081]&~m[2084]&m[2085]&m[2086]&m[2087])|(m[2081]&m[2084]&m[2085]&m[2086]&m[2087]));
    m[2088] = (((m[2086]&~m[2089]&~m[2090]&~m[2091]&~m[2092])|(~m[2086]&~m[2089]&~m[2090]&m[2091]&~m[2092])|(m[2086]&m[2089]&~m[2090]&m[2091]&~m[2092])|(m[2086]&~m[2089]&m[2090]&m[2091]&~m[2092])|(~m[2086]&m[2089]&~m[2090]&~m[2091]&m[2092])|(~m[2086]&~m[2089]&m[2090]&~m[2091]&m[2092])|(m[2086]&m[2089]&m[2090]&~m[2091]&m[2092])|(~m[2086]&m[2089]&m[2090]&m[2091]&m[2092]))&UnbiasedRNG[263])|((m[2086]&~m[2089]&~m[2090]&m[2091]&~m[2092])|(~m[2086]&~m[2089]&~m[2090]&~m[2091]&m[2092])|(m[2086]&~m[2089]&~m[2090]&~m[2091]&m[2092])|(m[2086]&m[2089]&~m[2090]&~m[2091]&m[2092])|(m[2086]&~m[2089]&m[2090]&~m[2091]&m[2092])|(~m[2086]&~m[2089]&~m[2090]&m[2091]&m[2092])|(m[2086]&~m[2089]&~m[2090]&m[2091]&m[2092])|(~m[2086]&m[2089]&~m[2090]&m[2091]&m[2092])|(m[2086]&m[2089]&~m[2090]&m[2091]&m[2092])|(~m[2086]&~m[2089]&m[2090]&m[2091]&m[2092])|(m[2086]&~m[2089]&m[2090]&m[2091]&m[2092])|(m[2086]&m[2089]&m[2090]&m[2091]&m[2092]));
    m[2093] = (((m[2091]&~m[2094]&~m[2095]&~m[2096]&~m[2097])|(~m[2091]&~m[2094]&~m[2095]&m[2096]&~m[2097])|(m[2091]&m[2094]&~m[2095]&m[2096]&~m[2097])|(m[2091]&~m[2094]&m[2095]&m[2096]&~m[2097])|(~m[2091]&m[2094]&~m[2095]&~m[2096]&m[2097])|(~m[2091]&~m[2094]&m[2095]&~m[2096]&m[2097])|(m[2091]&m[2094]&m[2095]&~m[2096]&m[2097])|(~m[2091]&m[2094]&m[2095]&m[2096]&m[2097]))&UnbiasedRNG[264])|((m[2091]&~m[2094]&~m[2095]&m[2096]&~m[2097])|(~m[2091]&~m[2094]&~m[2095]&~m[2096]&m[2097])|(m[2091]&~m[2094]&~m[2095]&~m[2096]&m[2097])|(m[2091]&m[2094]&~m[2095]&~m[2096]&m[2097])|(m[2091]&~m[2094]&m[2095]&~m[2096]&m[2097])|(~m[2091]&~m[2094]&~m[2095]&m[2096]&m[2097])|(m[2091]&~m[2094]&~m[2095]&m[2096]&m[2097])|(~m[2091]&m[2094]&~m[2095]&m[2096]&m[2097])|(m[2091]&m[2094]&~m[2095]&m[2096]&m[2097])|(~m[2091]&~m[2094]&m[2095]&m[2096]&m[2097])|(m[2091]&~m[2094]&m[2095]&m[2096]&m[2097])|(m[2091]&m[2094]&m[2095]&m[2096]&m[2097]));
    m[2098] = (((m[2082]&~m[2099]&~m[2100]&~m[2101]&~m[2102])|(~m[2082]&~m[2099]&~m[2100]&m[2101]&~m[2102])|(m[2082]&m[2099]&~m[2100]&m[2101]&~m[2102])|(m[2082]&~m[2099]&m[2100]&m[2101]&~m[2102])|(~m[2082]&m[2099]&~m[2100]&~m[2101]&m[2102])|(~m[2082]&~m[2099]&m[2100]&~m[2101]&m[2102])|(m[2082]&m[2099]&m[2100]&~m[2101]&m[2102])|(~m[2082]&m[2099]&m[2100]&m[2101]&m[2102]))&UnbiasedRNG[265])|((m[2082]&~m[2099]&~m[2100]&m[2101]&~m[2102])|(~m[2082]&~m[2099]&~m[2100]&~m[2101]&m[2102])|(m[2082]&~m[2099]&~m[2100]&~m[2101]&m[2102])|(m[2082]&m[2099]&~m[2100]&~m[2101]&m[2102])|(m[2082]&~m[2099]&m[2100]&~m[2101]&m[2102])|(~m[2082]&~m[2099]&~m[2100]&m[2101]&m[2102])|(m[2082]&~m[2099]&~m[2100]&m[2101]&m[2102])|(~m[2082]&m[2099]&~m[2100]&m[2101]&m[2102])|(m[2082]&m[2099]&~m[2100]&m[2101]&m[2102])|(~m[2082]&~m[2099]&m[2100]&m[2101]&m[2102])|(m[2082]&~m[2099]&m[2100]&m[2101]&m[2102])|(m[2082]&m[2099]&m[2100]&m[2101]&m[2102]));
    m[2103] = (((m[2101]&~m[2104]&~m[2105]&~m[2106]&~m[2107])|(~m[2101]&~m[2104]&~m[2105]&m[2106]&~m[2107])|(m[2101]&m[2104]&~m[2105]&m[2106]&~m[2107])|(m[2101]&~m[2104]&m[2105]&m[2106]&~m[2107])|(~m[2101]&m[2104]&~m[2105]&~m[2106]&m[2107])|(~m[2101]&~m[2104]&m[2105]&~m[2106]&m[2107])|(m[2101]&m[2104]&m[2105]&~m[2106]&m[2107])|(~m[2101]&m[2104]&m[2105]&m[2106]&m[2107]))&UnbiasedRNG[266])|((m[2101]&~m[2104]&~m[2105]&m[2106]&~m[2107])|(~m[2101]&~m[2104]&~m[2105]&~m[2106]&m[2107])|(m[2101]&~m[2104]&~m[2105]&~m[2106]&m[2107])|(m[2101]&m[2104]&~m[2105]&~m[2106]&m[2107])|(m[2101]&~m[2104]&m[2105]&~m[2106]&m[2107])|(~m[2101]&~m[2104]&~m[2105]&m[2106]&m[2107])|(m[2101]&~m[2104]&~m[2105]&m[2106]&m[2107])|(~m[2101]&m[2104]&~m[2105]&m[2106]&m[2107])|(m[2101]&m[2104]&~m[2105]&m[2106]&m[2107])|(~m[2101]&~m[2104]&m[2105]&m[2106]&m[2107])|(m[2101]&~m[2104]&m[2105]&m[2106]&m[2107])|(m[2101]&m[2104]&m[2105]&m[2106]&m[2107]));
    m[2108] = (((m[2106]&~m[2109]&~m[2110]&~m[2111]&~m[2112])|(~m[2106]&~m[2109]&~m[2110]&m[2111]&~m[2112])|(m[2106]&m[2109]&~m[2110]&m[2111]&~m[2112])|(m[2106]&~m[2109]&m[2110]&m[2111]&~m[2112])|(~m[2106]&m[2109]&~m[2110]&~m[2111]&m[2112])|(~m[2106]&~m[2109]&m[2110]&~m[2111]&m[2112])|(m[2106]&m[2109]&m[2110]&~m[2111]&m[2112])|(~m[2106]&m[2109]&m[2110]&m[2111]&m[2112]))&UnbiasedRNG[267])|((m[2106]&~m[2109]&~m[2110]&m[2111]&~m[2112])|(~m[2106]&~m[2109]&~m[2110]&~m[2111]&m[2112])|(m[2106]&~m[2109]&~m[2110]&~m[2111]&m[2112])|(m[2106]&m[2109]&~m[2110]&~m[2111]&m[2112])|(m[2106]&~m[2109]&m[2110]&~m[2111]&m[2112])|(~m[2106]&~m[2109]&~m[2110]&m[2111]&m[2112])|(m[2106]&~m[2109]&~m[2110]&m[2111]&m[2112])|(~m[2106]&m[2109]&~m[2110]&m[2111]&m[2112])|(m[2106]&m[2109]&~m[2110]&m[2111]&m[2112])|(~m[2106]&~m[2109]&m[2110]&m[2111]&m[2112])|(m[2106]&~m[2109]&m[2110]&m[2111]&m[2112])|(m[2106]&m[2109]&m[2110]&m[2111]&m[2112]));
    m[2113] = (((m[2102]&~m[2114]&~m[2115]&~m[2116]&~m[2117])|(~m[2102]&~m[2114]&~m[2115]&m[2116]&~m[2117])|(m[2102]&m[2114]&~m[2115]&m[2116]&~m[2117])|(m[2102]&~m[2114]&m[2115]&m[2116]&~m[2117])|(~m[2102]&m[2114]&~m[2115]&~m[2116]&m[2117])|(~m[2102]&~m[2114]&m[2115]&~m[2116]&m[2117])|(m[2102]&m[2114]&m[2115]&~m[2116]&m[2117])|(~m[2102]&m[2114]&m[2115]&m[2116]&m[2117]))&UnbiasedRNG[268])|((m[2102]&~m[2114]&~m[2115]&m[2116]&~m[2117])|(~m[2102]&~m[2114]&~m[2115]&~m[2116]&m[2117])|(m[2102]&~m[2114]&~m[2115]&~m[2116]&m[2117])|(m[2102]&m[2114]&~m[2115]&~m[2116]&m[2117])|(m[2102]&~m[2114]&m[2115]&~m[2116]&m[2117])|(~m[2102]&~m[2114]&~m[2115]&m[2116]&m[2117])|(m[2102]&~m[2114]&~m[2115]&m[2116]&m[2117])|(~m[2102]&m[2114]&~m[2115]&m[2116]&m[2117])|(m[2102]&m[2114]&~m[2115]&m[2116]&m[2117])|(~m[2102]&~m[2114]&m[2115]&m[2116]&m[2117])|(m[2102]&~m[2114]&m[2115]&m[2116]&m[2117])|(m[2102]&m[2114]&m[2115]&m[2116]&m[2117]));
    m[2118] = (((m[2116]&~m[2119]&~m[2120]&~m[2121]&~m[2122])|(~m[2116]&~m[2119]&~m[2120]&m[2121]&~m[2122])|(m[2116]&m[2119]&~m[2120]&m[2121]&~m[2122])|(m[2116]&~m[2119]&m[2120]&m[2121]&~m[2122])|(~m[2116]&m[2119]&~m[2120]&~m[2121]&m[2122])|(~m[2116]&~m[2119]&m[2120]&~m[2121]&m[2122])|(m[2116]&m[2119]&m[2120]&~m[2121]&m[2122])|(~m[2116]&m[2119]&m[2120]&m[2121]&m[2122]))&UnbiasedRNG[269])|((m[2116]&~m[2119]&~m[2120]&m[2121]&~m[2122])|(~m[2116]&~m[2119]&~m[2120]&~m[2121]&m[2122])|(m[2116]&~m[2119]&~m[2120]&~m[2121]&m[2122])|(m[2116]&m[2119]&~m[2120]&~m[2121]&m[2122])|(m[2116]&~m[2119]&m[2120]&~m[2121]&m[2122])|(~m[2116]&~m[2119]&~m[2120]&m[2121]&m[2122])|(m[2116]&~m[2119]&~m[2120]&m[2121]&m[2122])|(~m[2116]&m[2119]&~m[2120]&m[2121]&m[2122])|(m[2116]&m[2119]&~m[2120]&m[2121]&m[2122])|(~m[2116]&~m[2119]&m[2120]&m[2121]&m[2122])|(m[2116]&~m[2119]&m[2120]&m[2121]&m[2122])|(m[2116]&m[2119]&m[2120]&m[2121]&m[2122]));
    m[2123] = (((m[2117]&~m[2124]&~m[2125]&~m[2126]&~m[2127])|(~m[2117]&~m[2124]&~m[2125]&m[2126]&~m[2127])|(m[2117]&m[2124]&~m[2125]&m[2126]&~m[2127])|(m[2117]&~m[2124]&m[2125]&m[2126]&~m[2127])|(~m[2117]&m[2124]&~m[2125]&~m[2126]&m[2127])|(~m[2117]&~m[2124]&m[2125]&~m[2126]&m[2127])|(m[2117]&m[2124]&m[2125]&~m[2126]&m[2127])|(~m[2117]&m[2124]&m[2125]&m[2126]&m[2127]))&UnbiasedRNG[270])|((m[2117]&~m[2124]&~m[2125]&m[2126]&~m[2127])|(~m[2117]&~m[2124]&~m[2125]&~m[2126]&m[2127])|(m[2117]&~m[2124]&~m[2125]&~m[2126]&m[2127])|(m[2117]&m[2124]&~m[2125]&~m[2126]&m[2127])|(m[2117]&~m[2124]&m[2125]&~m[2126]&m[2127])|(~m[2117]&~m[2124]&~m[2125]&m[2126]&m[2127])|(m[2117]&~m[2124]&~m[2125]&m[2126]&m[2127])|(~m[2117]&m[2124]&~m[2125]&m[2126]&m[2127])|(m[2117]&m[2124]&~m[2125]&m[2126]&m[2127])|(~m[2117]&~m[2124]&m[2125]&m[2126]&m[2127])|(m[2117]&~m[2124]&m[2125]&m[2126]&m[2127])|(m[2117]&m[2124]&m[2125]&m[2126]&m[2127]));
end

always @(posedge color1_clk) begin
    m[32] = (((m[0]&m[160]&~m[161]&~m[162]&~m[163])|(m[0]&~m[160]&m[161]&~m[162]&~m[163])|(~m[0]&m[160]&m[161]&~m[162]&~m[163])|(m[0]&~m[160]&~m[161]&m[162]&~m[163])|(~m[0]&m[160]&~m[161]&m[162]&~m[163])|(~m[0]&~m[160]&m[161]&m[162]&~m[163])|(m[0]&~m[160]&~m[161]&~m[162]&m[163])|(~m[0]&m[160]&~m[161]&~m[162]&m[163])|(~m[0]&~m[160]&m[161]&~m[162]&m[163])|(~m[0]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[256])|(((m[0]&m[160]&m[161]&~m[162]&~m[163])|(m[0]&m[160]&~m[161]&m[162]&~m[163])|(m[0]&~m[160]&m[161]&m[162]&~m[163])|(~m[0]&m[160]&m[161]&m[162]&~m[163])|(m[0]&m[160]&~m[161]&~m[162]&m[163])|(m[0]&~m[160]&m[161]&~m[162]&m[163])|(~m[0]&m[160]&m[161]&~m[162]&m[163])|(m[0]&~m[160]&~m[161]&m[162]&m[163])|(~m[0]&m[160]&~m[161]&m[162]&m[163])|(~m[0]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[256])|((m[0]&m[160]&m[161]&m[162]&~m[163])|(m[0]&m[160]&m[161]&~m[162]&m[163])|(m[0]&m[160]&~m[161]&m[162]&m[163])|(m[0]&~m[160]&m[161]&m[162]&m[163])|(~m[0]&m[160]&m[161]&m[162]&m[163])|(m[0]&m[160]&m[161]&m[162]&m[163]));
    m[33] = (((m[0]&m[164]&~m[165]&~m[166]&~m[167])|(m[0]&~m[164]&m[165]&~m[166]&~m[167])|(~m[0]&m[164]&m[165]&~m[166]&~m[167])|(m[0]&~m[164]&~m[165]&m[166]&~m[167])|(~m[0]&m[164]&~m[165]&m[166]&~m[167])|(~m[0]&~m[164]&m[165]&m[166]&~m[167])|(m[0]&~m[164]&~m[165]&~m[166]&m[167])|(~m[0]&m[164]&~m[165]&~m[166]&m[167])|(~m[0]&~m[164]&m[165]&~m[166]&m[167])|(~m[0]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[257])|(((m[0]&m[164]&m[165]&~m[166]&~m[167])|(m[0]&m[164]&~m[165]&m[166]&~m[167])|(m[0]&~m[164]&m[165]&m[166]&~m[167])|(~m[0]&m[164]&m[165]&m[166]&~m[167])|(m[0]&m[164]&~m[165]&~m[166]&m[167])|(m[0]&~m[164]&m[165]&~m[166]&m[167])|(~m[0]&m[164]&m[165]&~m[166]&m[167])|(m[0]&~m[164]&~m[165]&m[166]&m[167])|(~m[0]&m[164]&~m[165]&m[166]&m[167])|(~m[0]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[257])|((m[0]&m[164]&m[165]&m[166]&~m[167])|(m[0]&m[164]&m[165]&~m[166]&m[167])|(m[0]&m[164]&~m[165]&m[166]&m[167])|(m[0]&~m[164]&m[165]&m[166]&m[167])|(~m[0]&m[164]&m[165]&m[166]&m[167])|(m[0]&m[164]&m[165]&m[166]&m[167]));
    m[34] = (((m[0]&m[168]&~m[169]&~m[170]&~m[171])|(m[0]&~m[168]&m[169]&~m[170]&~m[171])|(~m[0]&m[168]&m[169]&~m[170]&~m[171])|(m[0]&~m[168]&~m[169]&m[170]&~m[171])|(~m[0]&m[168]&~m[169]&m[170]&~m[171])|(~m[0]&~m[168]&m[169]&m[170]&~m[171])|(m[0]&~m[168]&~m[169]&~m[170]&m[171])|(~m[0]&m[168]&~m[169]&~m[170]&m[171])|(~m[0]&~m[168]&m[169]&~m[170]&m[171])|(~m[0]&~m[168]&~m[169]&m[170]&m[171]))&BiasedRNG[258])|(((m[0]&m[168]&m[169]&~m[170]&~m[171])|(m[0]&m[168]&~m[169]&m[170]&~m[171])|(m[0]&~m[168]&m[169]&m[170]&~m[171])|(~m[0]&m[168]&m[169]&m[170]&~m[171])|(m[0]&m[168]&~m[169]&~m[170]&m[171])|(m[0]&~m[168]&m[169]&~m[170]&m[171])|(~m[0]&m[168]&m[169]&~m[170]&m[171])|(m[0]&~m[168]&~m[169]&m[170]&m[171])|(~m[0]&m[168]&~m[169]&m[170]&m[171])|(~m[0]&~m[168]&m[169]&m[170]&m[171]))&~BiasedRNG[258])|((m[0]&m[168]&m[169]&m[170]&~m[171])|(m[0]&m[168]&m[169]&~m[170]&m[171])|(m[0]&m[168]&~m[169]&m[170]&m[171])|(m[0]&~m[168]&m[169]&m[170]&m[171])|(~m[0]&m[168]&m[169]&m[170]&m[171])|(m[0]&m[168]&m[169]&m[170]&m[171]));
    m[35] = (((m[0]&m[172]&~m[173]&~m[174]&~m[175])|(m[0]&~m[172]&m[173]&~m[174]&~m[175])|(~m[0]&m[172]&m[173]&~m[174]&~m[175])|(m[0]&~m[172]&~m[173]&m[174]&~m[175])|(~m[0]&m[172]&~m[173]&m[174]&~m[175])|(~m[0]&~m[172]&m[173]&m[174]&~m[175])|(m[0]&~m[172]&~m[173]&~m[174]&m[175])|(~m[0]&m[172]&~m[173]&~m[174]&m[175])|(~m[0]&~m[172]&m[173]&~m[174]&m[175])|(~m[0]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[259])|(((m[0]&m[172]&m[173]&~m[174]&~m[175])|(m[0]&m[172]&~m[173]&m[174]&~m[175])|(m[0]&~m[172]&m[173]&m[174]&~m[175])|(~m[0]&m[172]&m[173]&m[174]&~m[175])|(m[0]&m[172]&~m[173]&~m[174]&m[175])|(m[0]&~m[172]&m[173]&~m[174]&m[175])|(~m[0]&m[172]&m[173]&~m[174]&m[175])|(m[0]&~m[172]&~m[173]&m[174]&m[175])|(~m[0]&m[172]&~m[173]&m[174]&m[175])|(~m[0]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[259])|((m[0]&m[172]&m[173]&m[174]&~m[175])|(m[0]&m[172]&m[173]&~m[174]&m[175])|(m[0]&m[172]&~m[173]&m[174]&m[175])|(m[0]&~m[172]&m[173]&m[174]&m[175])|(~m[0]&m[172]&m[173]&m[174]&m[175])|(m[0]&m[172]&m[173]&m[174]&m[175]));
    m[36] = (((m[1]&m[176]&~m[177]&~m[178]&~m[179])|(m[1]&~m[176]&m[177]&~m[178]&~m[179])|(~m[1]&m[176]&m[177]&~m[178]&~m[179])|(m[1]&~m[176]&~m[177]&m[178]&~m[179])|(~m[1]&m[176]&~m[177]&m[178]&~m[179])|(~m[1]&~m[176]&m[177]&m[178]&~m[179])|(m[1]&~m[176]&~m[177]&~m[178]&m[179])|(~m[1]&m[176]&~m[177]&~m[178]&m[179])|(~m[1]&~m[176]&m[177]&~m[178]&m[179])|(~m[1]&~m[176]&~m[177]&m[178]&m[179]))&BiasedRNG[260])|(((m[1]&m[176]&m[177]&~m[178]&~m[179])|(m[1]&m[176]&~m[177]&m[178]&~m[179])|(m[1]&~m[176]&m[177]&m[178]&~m[179])|(~m[1]&m[176]&m[177]&m[178]&~m[179])|(m[1]&m[176]&~m[177]&~m[178]&m[179])|(m[1]&~m[176]&m[177]&~m[178]&m[179])|(~m[1]&m[176]&m[177]&~m[178]&m[179])|(m[1]&~m[176]&~m[177]&m[178]&m[179])|(~m[1]&m[176]&~m[177]&m[178]&m[179])|(~m[1]&~m[176]&m[177]&m[178]&m[179]))&~BiasedRNG[260])|((m[1]&m[176]&m[177]&m[178]&~m[179])|(m[1]&m[176]&m[177]&~m[178]&m[179])|(m[1]&m[176]&~m[177]&m[178]&m[179])|(m[1]&~m[176]&m[177]&m[178]&m[179])|(~m[1]&m[176]&m[177]&m[178]&m[179])|(m[1]&m[176]&m[177]&m[178]&m[179]));
    m[37] = (((m[1]&m[180]&~m[181]&~m[182]&~m[183])|(m[1]&~m[180]&m[181]&~m[182]&~m[183])|(~m[1]&m[180]&m[181]&~m[182]&~m[183])|(m[1]&~m[180]&~m[181]&m[182]&~m[183])|(~m[1]&m[180]&~m[181]&m[182]&~m[183])|(~m[1]&~m[180]&m[181]&m[182]&~m[183])|(m[1]&~m[180]&~m[181]&~m[182]&m[183])|(~m[1]&m[180]&~m[181]&~m[182]&m[183])|(~m[1]&~m[180]&m[181]&~m[182]&m[183])|(~m[1]&~m[180]&~m[181]&m[182]&m[183]))&BiasedRNG[261])|(((m[1]&m[180]&m[181]&~m[182]&~m[183])|(m[1]&m[180]&~m[181]&m[182]&~m[183])|(m[1]&~m[180]&m[181]&m[182]&~m[183])|(~m[1]&m[180]&m[181]&m[182]&~m[183])|(m[1]&m[180]&~m[181]&~m[182]&m[183])|(m[1]&~m[180]&m[181]&~m[182]&m[183])|(~m[1]&m[180]&m[181]&~m[182]&m[183])|(m[1]&~m[180]&~m[181]&m[182]&m[183])|(~m[1]&m[180]&~m[181]&m[182]&m[183])|(~m[1]&~m[180]&m[181]&m[182]&m[183]))&~BiasedRNG[261])|((m[1]&m[180]&m[181]&m[182]&~m[183])|(m[1]&m[180]&m[181]&~m[182]&m[183])|(m[1]&m[180]&~m[181]&m[182]&m[183])|(m[1]&~m[180]&m[181]&m[182]&m[183])|(~m[1]&m[180]&m[181]&m[182]&m[183])|(m[1]&m[180]&m[181]&m[182]&m[183]));
    m[38] = (((m[1]&m[184]&~m[185]&~m[186]&~m[187])|(m[1]&~m[184]&m[185]&~m[186]&~m[187])|(~m[1]&m[184]&m[185]&~m[186]&~m[187])|(m[1]&~m[184]&~m[185]&m[186]&~m[187])|(~m[1]&m[184]&~m[185]&m[186]&~m[187])|(~m[1]&~m[184]&m[185]&m[186]&~m[187])|(m[1]&~m[184]&~m[185]&~m[186]&m[187])|(~m[1]&m[184]&~m[185]&~m[186]&m[187])|(~m[1]&~m[184]&m[185]&~m[186]&m[187])|(~m[1]&~m[184]&~m[185]&m[186]&m[187]))&BiasedRNG[262])|(((m[1]&m[184]&m[185]&~m[186]&~m[187])|(m[1]&m[184]&~m[185]&m[186]&~m[187])|(m[1]&~m[184]&m[185]&m[186]&~m[187])|(~m[1]&m[184]&m[185]&m[186]&~m[187])|(m[1]&m[184]&~m[185]&~m[186]&m[187])|(m[1]&~m[184]&m[185]&~m[186]&m[187])|(~m[1]&m[184]&m[185]&~m[186]&m[187])|(m[1]&~m[184]&~m[185]&m[186]&m[187])|(~m[1]&m[184]&~m[185]&m[186]&m[187])|(~m[1]&~m[184]&m[185]&m[186]&m[187]))&~BiasedRNG[262])|((m[1]&m[184]&m[185]&m[186]&~m[187])|(m[1]&m[184]&m[185]&~m[186]&m[187])|(m[1]&m[184]&~m[185]&m[186]&m[187])|(m[1]&~m[184]&m[185]&m[186]&m[187])|(~m[1]&m[184]&m[185]&m[186]&m[187])|(m[1]&m[184]&m[185]&m[186]&m[187]));
    m[39] = (((m[1]&m[188]&~m[189]&~m[190]&~m[191])|(m[1]&~m[188]&m[189]&~m[190]&~m[191])|(~m[1]&m[188]&m[189]&~m[190]&~m[191])|(m[1]&~m[188]&~m[189]&m[190]&~m[191])|(~m[1]&m[188]&~m[189]&m[190]&~m[191])|(~m[1]&~m[188]&m[189]&m[190]&~m[191])|(m[1]&~m[188]&~m[189]&~m[190]&m[191])|(~m[1]&m[188]&~m[189]&~m[190]&m[191])|(~m[1]&~m[188]&m[189]&~m[190]&m[191])|(~m[1]&~m[188]&~m[189]&m[190]&m[191]))&BiasedRNG[263])|(((m[1]&m[188]&m[189]&~m[190]&~m[191])|(m[1]&m[188]&~m[189]&m[190]&~m[191])|(m[1]&~m[188]&m[189]&m[190]&~m[191])|(~m[1]&m[188]&m[189]&m[190]&~m[191])|(m[1]&m[188]&~m[189]&~m[190]&m[191])|(m[1]&~m[188]&m[189]&~m[190]&m[191])|(~m[1]&m[188]&m[189]&~m[190]&m[191])|(m[1]&~m[188]&~m[189]&m[190]&m[191])|(~m[1]&m[188]&~m[189]&m[190]&m[191])|(~m[1]&~m[188]&m[189]&m[190]&m[191]))&~BiasedRNG[263])|((m[1]&m[188]&m[189]&m[190]&~m[191])|(m[1]&m[188]&m[189]&~m[190]&m[191])|(m[1]&m[188]&~m[189]&m[190]&m[191])|(m[1]&~m[188]&m[189]&m[190]&m[191])|(~m[1]&m[188]&m[189]&m[190]&m[191])|(m[1]&m[188]&m[189]&m[190]&m[191]));
    m[40] = (((m[2]&m[192]&~m[193]&~m[194]&~m[195])|(m[2]&~m[192]&m[193]&~m[194]&~m[195])|(~m[2]&m[192]&m[193]&~m[194]&~m[195])|(m[2]&~m[192]&~m[193]&m[194]&~m[195])|(~m[2]&m[192]&~m[193]&m[194]&~m[195])|(~m[2]&~m[192]&m[193]&m[194]&~m[195])|(m[2]&~m[192]&~m[193]&~m[194]&m[195])|(~m[2]&m[192]&~m[193]&~m[194]&m[195])|(~m[2]&~m[192]&m[193]&~m[194]&m[195])|(~m[2]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[264])|(((m[2]&m[192]&m[193]&~m[194]&~m[195])|(m[2]&m[192]&~m[193]&m[194]&~m[195])|(m[2]&~m[192]&m[193]&m[194]&~m[195])|(~m[2]&m[192]&m[193]&m[194]&~m[195])|(m[2]&m[192]&~m[193]&~m[194]&m[195])|(m[2]&~m[192]&m[193]&~m[194]&m[195])|(~m[2]&m[192]&m[193]&~m[194]&m[195])|(m[2]&~m[192]&~m[193]&m[194]&m[195])|(~m[2]&m[192]&~m[193]&m[194]&m[195])|(~m[2]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[264])|((m[2]&m[192]&m[193]&m[194]&~m[195])|(m[2]&m[192]&m[193]&~m[194]&m[195])|(m[2]&m[192]&~m[193]&m[194]&m[195])|(m[2]&~m[192]&m[193]&m[194]&m[195])|(~m[2]&m[192]&m[193]&m[194]&m[195])|(m[2]&m[192]&m[193]&m[194]&m[195]));
    m[41] = (((m[2]&m[196]&~m[197]&~m[198]&~m[199])|(m[2]&~m[196]&m[197]&~m[198]&~m[199])|(~m[2]&m[196]&m[197]&~m[198]&~m[199])|(m[2]&~m[196]&~m[197]&m[198]&~m[199])|(~m[2]&m[196]&~m[197]&m[198]&~m[199])|(~m[2]&~m[196]&m[197]&m[198]&~m[199])|(m[2]&~m[196]&~m[197]&~m[198]&m[199])|(~m[2]&m[196]&~m[197]&~m[198]&m[199])|(~m[2]&~m[196]&m[197]&~m[198]&m[199])|(~m[2]&~m[196]&~m[197]&m[198]&m[199]))&BiasedRNG[265])|(((m[2]&m[196]&m[197]&~m[198]&~m[199])|(m[2]&m[196]&~m[197]&m[198]&~m[199])|(m[2]&~m[196]&m[197]&m[198]&~m[199])|(~m[2]&m[196]&m[197]&m[198]&~m[199])|(m[2]&m[196]&~m[197]&~m[198]&m[199])|(m[2]&~m[196]&m[197]&~m[198]&m[199])|(~m[2]&m[196]&m[197]&~m[198]&m[199])|(m[2]&~m[196]&~m[197]&m[198]&m[199])|(~m[2]&m[196]&~m[197]&m[198]&m[199])|(~m[2]&~m[196]&m[197]&m[198]&m[199]))&~BiasedRNG[265])|((m[2]&m[196]&m[197]&m[198]&~m[199])|(m[2]&m[196]&m[197]&~m[198]&m[199])|(m[2]&m[196]&~m[197]&m[198]&m[199])|(m[2]&~m[196]&m[197]&m[198]&m[199])|(~m[2]&m[196]&m[197]&m[198]&m[199])|(m[2]&m[196]&m[197]&m[198]&m[199]));
    m[42] = (((m[2]&m[200]&~m[201]&~m[202]&~m[203])|(m[2]&~m[200]&m[201]&~m[202]&~m[203])|(~m[2]&m[200]&m[201]&~m[202]&~m[203])|(m[2]&~m[200]&~m[201]&m[202]&~m[203])|(~m[2]&m[200]&~m[201]&m[202]&~m[203])|(~m[2]&~m[200]&m[201]&m[202]&~m[203])|(m[2]&~m[200]&~m[201]&~m[202]&m[203])|(~m[2]&m[200]&~m[201]&~m[202]&m[203])|(~m[2]&~m[200]&m[201]&~m[202]&m[203])|(~m[2]&~m[200]&~m[201]&m[202]&m[203]))&BiasedRNG[266])|(((m[2]&m[200]&m[201]&~m[202]&~m[203])|(m[2]&m[200]&~m[201]&m[202]&~m[203])|(m[2]&~m[200]&m[201]&m[202]&~m[203])|(~m[2]&m[200]&m[201]&m[202]&~m[203])|(m[2]&m[200]&~m[201]&~m[202]&m[203])|(m[2]&~m[200]&m[201]&~m[202]&m[203])|(~m[2]&m[200]&m[201]&~m[202]&m[203])|(m[2]&~m[200]&~m[201]&m[202]&m[203])|(~m[2]&m[200]&~m[201]&m[202]&m[203])|(~m[2]&~m[200]&m[201]&m[202]&m[203]))&~BiasedRNG[266])|((m[2]&m[200]&m[201]&m[202]&~m[203])|(m[2]&m[200]&m[201]&~m[202]&m[203])|(m[2]&m[200]&~m[201]&m[202]&m[203])|(m[2]&~m[200]&m[201]&m[202]&m[203])|(~m[2]&m[200]&m[201]&m[202]&m[203])|(m[2]&m[200]&m[201]&m[202]&m[203]));
    m[43] = (((m[2]&m[204]&~m[205]&~m[206]&~m[207])|(m[2]&~m[204]&m[205]&~m[206]&~m[207])|(~m[2]&m[204]&m[205]&~m[206]&~m[207])|(m[2]&~m[204]&~m[205]&m[206]&~m[207])|(~m[2]&m[204]&~m[205]&m[206]&~m[207])|(~m[2]&~m[204]&m[205]&m[206]&~m[207])|(m[2]&~m[204]&~m[205]&~m[206]&m[207])|(~m[2]&m[204]&~m[205]&~m[206]&m[207])|(~m[2]&~m[204]&m[205]&~m[206]&m[207])|(~m[2]&~m[204]&~m[205]&m[206]&m[207]))&BiasedRNG[267])|(((m[2]&m[204]&m[205]&~m[206]&~m[207])|(m[2]&m[204]&~m[205]&m[206]&~m[207])|(m[2]&~m[204]&m[205]&m[206]&~m[207])|(~m[2]&m[204]&m[205]&m[206]&~m[207])|(m[2]&m[204]&~m[205]&~m[206]&m[207])|(m[2]&~m[204]&m[205]&~m[206]&m[207])|(~m[2]&m[204]&m[205]&~m[206]&m[207])|(m[2]&~m[204]&~m[205]&m[206]&m[207])|(~m[2]&m[204]&~m[205]&m[206]&m[207])|(~m[2]&~m[204]&m[205]&m[206]&m[207]))&~BiasedRNG[267])|((m[2]&m[204]&m[205]&m[206]&~m[207])|(m[2]&m[204]&m[205]&~m[206]&m[207])|(m[2]&m[204]&~m[205]&m[206]&m[207])|(m[2]&~m[204]&m[205]&m[206]&m[207])|(~m[2]&m[204]&m[205]&m[206]&m[207])|(m[2]&m[204]&m[205]&m[206]&m[207]));
    m[44] = (((m[3]&m[208]&~m[209]&~m[210]&~m[211])|(m[3]&~m[208]&m[209]&~m[210]&~m[211])|(~m[3]&m[208]&m[209]&~m[210]&~m[211])|(m[3]&~m[208]&~m[209]&m[210]&~m[211])|(~m[3]&m[208]&~m[209]&m[210]&~m[211])|(~m[3]&~m[208]&m[209]&m[210]&~m[211])|(m[3]&~m[208]&~m[209]&~m[210]&m[211])|(~m[3]&m[208]&~m[209]&~m[210]&m[211])|(~m[3]&~m[208]&m[209]&~m[210]&m[211])|(~m[3]&~m[208]&~m[209]&m[210]&m[211]))&BiasedRNG[268])|(((m[3]&m[208]&m[209]&~m[210]&~m[211])|(m[3]&m[208]&~m[209]&m[210]&~m[211])|(m[3]&~m[208]&m[209]&m[210]&~m[211])|(~m[3]&m[208]&m[209]&m[210]&~m[211])|(m[3]&m[208]&~m[209]&~m[210]&m[211])|(m[3]&~m[208]&m[209]&~m[210]&m[211])|(~m[3]&m[208]&m[209]&~m[210]&m[211])|(m[3]&~m[208]&~m[209]&m[210]&m[211])|(~m[3]&m[208]&~m[209]&m[210]&m[211])|(~m[3]&~m[208]&m[209]&m[210]&m[211]))&~BiasedRNG[268])|((m[3]&m[208]&m[209]&m[210]&~m[211])|(m[3]&m[208]&m[209]&~m[210]&m[211])|(m[3]&m[208]&~m[209]&m[210]&m[211])|(m[3]&~m[208]&m[209]&m[210]&m[211])|(~m[3]&m[208]&m[209]&m[210]&m[211])|(m[3]&m[208]&m[209]&m[210]&m[211]));
    m[45] = (((m[3]&m[212]&~m[213]&~m[214]&~m[215])|(m[3]&~m[212]&m[213]&~m[214]&~m[215])|(~m[3]&m[212]&m[213]&~m[214]&~m[215])|(m[3]&~m[212]&~m[213]&m[214]&~m[215])|(~m[3]&m[212]&~m[213]&m[214]&~m[215])|(~m[3]&~m[212]&m[213]&m[214]&~m[215])|(m[3]&~m[212]&~m[213]&~m[214]&m[215])|(~m[3]&m[212]&~m[213]&~m[214]&m[215])|(~m[3]&~m[212]&m[213]&~m[214]&m[215])|(~m[3]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[269])|(((m[3]&m[212]&m[213]&~m[214]&~m[215])|(m[3]&m[212]&~m[213]&m[214]&~m[215])|(m[3]&~m[212]&m[213]&m[214]&~m[215])|(~m[3]&m[212]&m[213]&m[214]&~m[215])|(m[3]&m[212]&~m[213]&~m[214]&m[215])|(m[3]&~m[212]&m[213]&~m[214]&m[215])|(~m[3]&m[212]&m[213]&~m[214]&m[215])|(m[3]&~m[212]&~m[213]&m[214]&m[215])|(~m[3]&m[212]&~m[213]&m[214]&m[215])|(~m[3]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[269])|((m[3]&m[212]&m[213]&m[214]&~m[215])|(m[3]&m[212]&m[213]&~m[214]&m[215])|(m[3]&m[212]&~m[213]&m[214]&m[215])|(m[3]&~m[212]&m[213]&m[214]&m[215])|(~m[3]&m[212]&m[213]&m[214]&m[215])|(m[3]&m[212]&m[213]&m[214]&m[215]));
    m[46] = (((m[3]&m[216]&~m[217]&~m[218]&~m[219])|(m[3]&~m[216]&m[217]&~m[218]&~m[219])|(~m[3]&m[216]&m[217]&~m[218]&~m[219])|(m[3]&~m[216]&~m[217]&m[218]&~m[219])|(~m[3]&m[216]&~m[217]&m[218]&~m[219])|(~m[3]&~m[216]&m[217]&m[218]&~m[219])|(m[3]&~m[216]&~m[217]&~m[218]&m[219])|(~m[3]&m[216]&~m[217]&~m[218]&m[219])|(~m[3]&~m[216]&m[217]&~m[218]&m[219])|(~m[3]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[270])|(((m[3]&m[216]&m[217]&~m[218]&~m[219])|(m[3]&m[216]&~m[217]&m[218]&~m[219])|(m[3]&~m[216]&m[217]&m[218]&~m[219])|(~m[3]&m[216]&m[217]&m[218]&~m[219])|(m[3]&m[216]&~m[217]&~m[218]&m[219])|(m[3]&~m[216]&m[217]&~m[218]&m[219])|(~m[3]&m[216]&m[217]&~m[218]&m[219])|(m[3]&~m[216]&~m[217]&m[218]&m[219])|(~m[3]&m[216]&~m[217]&m[218]&m[219])|(~m[3]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[270])|((m[3]&m[216]&m[217]&m[218]&~m[219])|(m[3]&m[216]&m[217]&~m[218]&m[219])|(m[3]&m[216]&~m[217]&m[218]&m[219])|(m[3]&~m[216]&m[217]&m[218]&m[219])|(~m[3]&m[216]&m[217]&m[218]&m[219])|(m[3]&m[216]&m[217]&m[218]&m[219]));
    m[47] = (((m[3]&m[220]&~m[221]&~m[222]&~m[223])|(m[3]&~m[220]&m[221]&~m[222]&~m[223])|(~m[3]&m[220]&m[221]&~m[222]&~m[223])|(m[3]&~m[220]&~m[221]&m[222]&~m[223])|(~m[3]&m[220]&~m[221]&m[222]&~m[223])|(~m[3]&~m[220]&m[221]&m[222]&~m[223])|(m[3]&~m[220]&~m[221]&~m[222]&m[223])|(~m[3]&m[220]&~m[221]&~m[222]&m[223])|(~m[3]&~m[220]&m[221]&~m[222]&m[223])|(~m[3]&~m[220]&~m[221]&m[222]&m[223]))&BiasedRNG[271])|(((m[3]&m[220]&m[221]&~m[222]&~m[223])|(m[3]&m[220]&~m[221]&m[222]&~m[223])|(m[3]&~m[220]&m[221]&m[222]&~m[223])|(~m[3]&m[220]&m[221]&m[222]&~m[223])|(m[3]&m[220]&~m[221]&~m[222]&m[223])|(m[3]&~m[220]&m[221]&~m[222]&m[223])|(~m[3]&m[220]&m[221]&~m[222]&m[223])|(m[3]&~m[220]&~m[221]&m[222]&m[223])|(~m[3]&m[220]&~m[221]&m[222]&m[223])|(~m[3]&~m[220]&m[221]&m[222]&m[223]))&~BiasedRNG[271])|((m[3]&m[220]&m[221]&m[222]&~m[223])|(m[3]&m[220]&m[221]&~m[222]&m[223])|(m[3]&m[220]&~m[221]&m[222]&m[223])|(m[3]&~m[220]&m[221]&m[222]&m[223])|(~m[3]&m[220]&m[221]&m[222]&m[223])|(m[3]&m[220]&m[221]&m[222]&m[223]));
    m[48] = (((m[4]&m[224]&~m[225]&~m[226]&~m[227])|(m[4]&~m[224]&m[225]&~m[226]&~m[227])|(~m[4]&m[224]&m[225]&~m[226]&~m[227])|(m[4]&~m[224]&~m[225]&m[226]&~m[227])|(~m[4]&m[224]&~m[225]&m[226]&~m[227])|(~m[4]&~m[224]&m[225]&m[226]&~m[227])|(m[4]&~m[224]&~m[225]&~m[226]&m[227])|(~m[4]&m[224]&~m[225]&~m[226]&m[227])|(~m[4]&~m[224]&m[225]&~m[226]&m[227])|(~m[4]&~m[224]&~m[225]&m[226]&m[227]))&BiasedRNG[272])|(((m[4]&m[224]&m[225]&~m[226]&~m[227])|(m[4]&m[224]&~m[225]&m[226]&~m[227])|(m[4]&~m[224]&m[225]&m[226]&~m[227])|(~m[4]&m[224]&m[225]&m[226]&~m[227])|(m[4]&m[224]&~m[225]&~m[226]&m[227])|(m[4]&~m[224]&m[225]&~m[226]&m[227])|(~m[4]&m[224]&m[225]&~m[226]&m[227])|(m[4]&~m[224]&~m[225]&m[226]&m[227])|(~m[4]&m[224]&~m[225]&m[226]&m[227])|(~m[4]&~m[224]&m[225]&m[226]&m[227]))&~BiasedRNG[272])|((m[4]&m[224]&m[225]&m[226]&~m[227])|(m[4]&m[224]&m[225]&~m[226]&m[227])|(m[4]&m[224]&~m[225]&m[226]&m[227])|(m[4]&~m[224]&m[225]&m[226]&m[227])|(~m[4]&m[224]&m[225]&m[226]&m[227])|(m[4]&m[224]&m[225]&m[226]&m[227]));
    m[49] = (((m[4]&m[228]&~m[229]&~m[230]&~m[231])|(m[4]&~m[228]&m[229]&~m[230]&~m[231])|(~m[4]&m[228]&m[229]&~m[230]&~m[231])|(m[4]&~m[228]&~m[229]&m[230]&~m[231])|(~m[4]&m[228]&~m[229]&m[230]&~m[231])|(~m[4]&~m[228]&m[229]&m[230]&~m[231])|(m[4]&~m[228]&~m[229]&~m[230]&m[231])|(~m[4]&m[228]&~m[229]&~m[230]&m[231])|(~m[4]&~m[228]&m[229]&~m[230]&m[231])|(~m[4]&~m[228]&~m[229]&m[230]&m[231]))&BiasedRNG[273])|(((m[4]&m[228]&m[229]&~m[230]&~m[231])|(m[4]&m[228]&~m[229]&m[230]&~m[231])|(m[4]&~m[228]&m[229]&m[230]&~m[231])|(~m[4]&m[228]&m[229]&m[230]&~m[231])|(m[4]&m[228]&~m[229]&~m[230]&m[231])|(m[4]&~m[228]&m[229]&~m[230]&m[231])|(~m[4]&m[228]&m[229]&~m[230]&m[231])|(m[4]&~m[228]&~m[229]&m[230]&m[231])|(~m[4]&m[228]&~m[229]&m[230]&m[231])|(~m[4]&~m[228]&m[229]&m[230]&m[231]))&~BiasedRNG[273])|((m[4]&m[228]&m[229]&m[230]&~m[231])|(m[4]&m[228]&m[229]&~m[230]&m[231])|(m[4]&m[228]&~m[229]&m[230]&m[231])|(m[4]&~m[228]&m[229]&m[230]&m[231])|(~m[4]&m[228]&m[229]&m[230]&m[231])|(m[4]&m[228]&m[229]&m[230]&m[231]));
    m[50] = (((m[4]&m[232]&~m[233]&~m[234]&~m[235])|(m[4]&~m[232]&m[233]&~m[234]&~m[235])|(~m[4]&m[232]&m[233]&~m[234]&~m[235])|(m[4]&~m[232]&~m[233]&m[234]&~m[235])|(~m[4]&m[232]&~m[233]&m[234]&~m[235])|(~m[4]&~m[232]&m[233]&m[234]&~m[235])|(m[4]&~m[232]&~m[233]&~m[234]&m[235])|(~m[4]&m[232]&~m[233]&~m[234]&m[235])|(~m[4]&~m[232]&m[233]&~m[234]&m[235])|(~m[4]&~m[232]&~m[233]&m[234]&m[235]))&BiasedRNG[274])|(((m[4]&m[232]&m[233]&~m[234]&~m[235])|(m[4]&m[232]&~m[233]&m[234]&~m[235])|(m[4]&~m[232]&m[233]&m[234]&~m[235])|(~m[4]&m[232]&m[233]&m[234]&~m[235])|(m[4]&m[232]&~m[233]&~m[234]&m[235])|(m[4]&~m[232]&m[233]&~m[234]&m[235])|(~m[4]&m[232]&m[233]&~m[234]&m[235])|(m[4]&~m[232]&~m[233]&m[234]&m[235])|(~m[4]&m[232]&~m[233]&m[234]&m[235])|(~m[4]&~m[232]&m[233]&m[234]&m[235]))&~BiasedRNG[274])|((m[4]&m[232]&m[233]&m[234]&~m[235])|(m[4]&m[232]&m[233]&~m[234]&m[235])|(m[4]&m[232]&~m[233]&m[234]&m[235])|(m[4]&~m[232]&m[233]&m[234]&m[235])|(~m[4]&m[232]&m[233]&m[234]&m[235])|(m[4]&m[232]&m[233]&m[234]&m[235]));
    m[51] = (((m[4]&m[236]&~m[237]&~m[238]&~m[239])|(m[4]&~m[236]&m[237]&~m[238]&~m[239])|(~m[4]&m[236]&m[237]&~m[238]&~m[239])|(m[4]&~m[236]&~m[237]&m[238]&~m[239])|(~m[4]&m[236]&~m[237]&m[238]&~m[239])|(~m[4]&~m[236]&m[237]&m[238]&~m[239])|(m[4]&~m[236]&~m[237]&~m[238]&m[239])|(~m[4]&m[236]&~m[237]&~m[238]&m[239])|(~m[4]&~m[236]&m[237]&~m[238]&m[239])|(~m[4]&~m[236]&~m[237]&m[238]&m[239]))&BiasedRNG[275])|(((m[4]&m[236]&m[237]&~m[238]&~m[239])|(m[4]&m[236]&~m[237]&m[238]&~m[239])|(m[4]&~m[236]&m[237]&m[238]&~m[239])|(~m[4]&m[236]&m[237]&m[238]&~m[239])|(m[4]&m[236]&~m[237]&~m[238]&m[239])|(m[4]&~m[236]&m[237]&~m[238]&m[239])|(~m[4]&m[236]&m[237]&~m[238]&m[239])|(m[4]&~m[236]&~m[237]&m[238]&m[239])|(~m[4]&m[236]&~m[237]&m[238]&m[239])|(~m[4]&~m[236]&m[237]&m[238]&m[239]))&~BiasedRNG[275])|((m[4]&m[236]&m[237]&m[238]&~m[239])|(m[4]&m[236]&m[237]&~m[238]&m[239])|(m[4]&m[236]&~m[237]&m[238]&m[239])|(m[4]&~m[236]&m[237]&m[238]&m[239])|(~m[4]&m[236]&m[237]&m[238]&m[239])|(m[4]&m[236]&m[237]&m[238]&m[239]));
    m[52] = (((m[5]&m[240]&~m[241]&~m[242]&~m[243])|(m[5]&~m[240]&m[241]&~m[242]&~m[243])|(~m[5]&m[240]&m[241]&~m[242]&~m[243])|(m[5]&~m[240]&~m[241]&m[242]&~m[243])|(~m[5]&m[240]&~m[241]&m[242]&~m[243])|(~m[5]&~m[240]&m[241]&m[242]&~m[243])|(m[5]&~m[240]&~m[241]&~m[242]&m[243])|(~m[5]&m[240]&~m[241]&~m[242]&m[243])|(~m[5]&~m[240]&m[241]&~m[242]&m[243])|(~m[5]&~m[240]&~m[241]&m[242]&m[243]))&BiasedRNG[276])|(((m[5]&m[240]&m[241]&~m[242]&~m[243])|(m[5]&m[240]&~m[241]&m[242]&~m[243])|(m[5]&~m[240]&m[241]&m[242]&~m[243])|(~m[5]&m[240]&m[241]&m[242]&~m[243])|(m[5]&m[240]&~m[241]&~m[242]&m[243])|(m[5]&~m[240]&m[241]&~m[242]&m[243])|(~m[5]&m[240]&m[241]&~m[242]&m[243])|(m[5]&~m[240]&~m[241]&m[242]&m[243])|(~m[5]&m[240]&~m[241]&m[242]&m[243])|(~m[5]&~m[240]&m[241]&m[242]&m[243]))&~BiasedRNG[276])|((m[5]&m[240]&m[241]&m[242]&~m[243])|(m[5]&m[240]&m[241]&~m[242]&m[243])|(m[5]&m[240]&~m[241]&m[242]&m[243])|(m[5]&~m[240]&m[241]&m[242]&m[243])|(~m[5]&m[240]&m[241]&m[242]&m[243])|(m[5]&m[240]&m[241]&m[242]&m[243]));
    m[53] = (((m[5]&m[244]&~m[245]&~m[246]&~m[247])|(m[5]&~m[244]&m[245]&~m[246]&~m[247])|(~m[5]&m[244]&m[245]&~m[246]&~m[247])|(m[5]&~m[244]&~m[245]&m[246]&~m[247])|(~m[5]&m[244]&~m[245]&m[246]&~m[247])|(~m[5]&~m[244]&m[245]&m[246]&~m[247])|(m[5]&~m[244]&~m[245]&~m[246]&m[247])|(~m[5]&m[244]&~m[245]&~m[246]&m[247])|(~m[5]&~m[244]&m[245]&~m[246]&m[247])|(~m[5]&~m[244]&~m[245]&m[246]&m[247]))&BiasedRNG[277])|(((m[5]&m[244]&m[245]&~m[246]&~m[247])|(m[5]&m[244]&~m[245]&m[246]&~m[247])|(m[5]&~m[244]&m[245]&m[246]&~m[247])|(~m[5]&m[244]&m[245]&m[246]&~m[247])|(m[5]&m[244]&~m[245]&~m[246]&m[247])|(m[5]&~m[244]&m[245]&~m[246]&m[247])|(~m[5]&m[244]&m[245]&~m[246]&m[247])|(m[5]&~m[244]&~m[245]&m[246]&m[247])|(~m[5]&m[244]&~m[245]&m[246]&m[247])|(~m[5]&~m[244]&m[245]&m[246]&m[247]))&~BiasedRNG[277])|((m[5]&m[244]&m[245]&m[246]&~m[247])|(m[5]&m[244]&m[245]&~m[246]&m[247])|(m[5]&m[244]&~m[245]&m[246]&m[247])|(m[5]&~m[244]&m[245]&m[246]&m[247])|(~m[5]&m[244]&m[245]&m[246]&m[247])|(m[5]&m[244]&m[245]&m[246]&m[247]));
    m[54] = (((m[5]&m[248]&~m[249]&~m[250]&~m[251])|(m[5]&~m[248]&m[249]&~m[250]&~m[251])|(~m[5]&m[248]&m[249]&~m[250]&~m[251])|(m[5]&~m[248]&~m[249]&m[250]&~m[251])|(~m[5]&m[248]&~m[249]&m[250]&~m[251])|(~m[5]&~m[248]&m[249]&m[250]&~m[251])|(m[5]&~m[248]&~m[249]&~m[250]&m[251])|(~m[5]&m[248]&~m[249]&~m[250]&m[251])|(~m[5]&~m[248]&m[249]&~m[250]&m[251])|(~m[5]&~m[248]&~m[249]&m[250]&m[251]))&BiasedRNG[278])|(((m[5]&m[248]&m[249]&~m[250]&~m[251])|(m[5]&m[248]&~m[249]&m[250]&~m[251])|(m[5]&~m[248]&m[249]&m[250]&~m[251])|(~m[5]&m[248]&m[249]&m[250]&~m[251])|(m[5]&m[248]&~m[249]&~m[250]&m[251])|(m[5]&~m[248]&m[249]&~m[250]&m[251])|(~m[5]&m[248]&m[249]&~m[250]&m[251])|(m[5]&~m[248]&~m[249]&m[250]&m[251])|(~m[5]&m[248]&~m[249]&m[250]&m[251])|(~m[5]&~m[248]&m[249]&m[250]&m[251]))&~BiasedRNG[278])|((m[5]&m[248]&m[249]&m[250]&~m[251])|(m[5]&m[248]&m[249]&~m[250]&m[251])|(m[5]&m[248]&~m[249]&m[250]&m[251])|(m[5]&~m[248]&m[249]&m[250]&m[251])|(~m[5]&m[248]&m[249]&m[250]&m[251])|(m[5]&m[248]&m[249]&m[250]&m[251]));
    m[55] = (((m[5]&m[252]&~m[253]&~m[254]&~m[255])|(m[5]&~m[252]&m[253]&~m[254]&~m[255])|(~m[5]&m[252]&m[253]&~m[254]&~m[255])|(m[5]&~m[252]&~m[253]&m[254]&~m[255])|(~m[5]&m[252]&~m[253]&m[254]&~m[255])|(~m[5]&~m[252]&m[253]&m[254]&~m[255])|(m[5]&~m[252]&~m[253]&~m[254]&m[255])|(~m[5]&m[252]&~m[253]&~m[254]&m[255])|(~m[5]&~m[252]&m[253]&~m[254]&m[255])|(~m[5]&~m[252]&~m[253]&m[254]&m[255]))&BiasedRNG[279])|(((m[5]&m[252]&m[253]&~m[254]&~m[255])|(m[5]&m[252]&~m[253]&m[254]&~m[255])|(m[5]&~m[252]&m[253]&m[254]&~m[255])|(~m[5]&m[252]&m[253]&m[254]&~m[255])|(m[5]&m[252]&~m[253]&~m[254]&m[255])|(m[5]&~m[252]&m[253]&~m[254]&m[255])|(~m[5]&m[252]&m[253]&~m[254]&m[255])|(m[5]&~m[252]&~m[253]&m[254]&m[255])|(~m[5]&m[252]&~m[253]&m[254]&m[255])|(~m[5]&~m[252]&m[253]&m[254]&m[255]))&~BiasedRNG[279])|((m[5]&m[252]&m[253]&m[254]&~m[255])|(m[5]&m[252]&m[253]&~m[254]&m[255])|(m[5]&m[252]&~m[253]&m[254]&m[255])|(m[5]&~m[252]&m[253]&m[254]&m[255])|(~m[5]&m[252]&m[253]&m[254]&m[255])|(m[5]&m[252]&m[253]&m[254]&m[255]));
    m[56] = (((m[6]&m[256]&~m[257]&~m[258]&~m[259])|(m[6]&~m[256]&m[257]&~m[258]&~m[259])|(~m[6]&m[256]&m[257]&~m[258]&~m[259])|(m[6]&~m[256]&~m[257]&m[258]&~m[259])|(~m[6]&m[256]&~m[257]&m[258]&~m[259])|(~m[6]&~m[256]&m[257]&m[258]&~m[259])|(m[6]&~m[256]&~m[257]&~m[258]&m[259])|(~m[6]&m[256]&~m[257]&~m[258]&m[259])|(~m[6]&~m[256]&m[257]&~m[258]&m[259])|(~m[6]&~m[256]&~m[257]&m[258]&m[259]))&BiasedRNG[280])|(((m[6]&m[256]&m[257]&~m[258]&~m[259])|(m[6]&m[256]&~m[257]&m[258]&~m[259])|(m[6]&~m[256]&m[257]&m[258]&~m[259])|(~m[6]&m[256]&m[257]&m[258]&~m[259])|(m[6]&m[256]&~m[257]&~m[258]&m[259])|(m[6]&~m[256]&m[257]&~m[258]&m[259])|(~m[6]&m[256]&m[257]&~m[258]&m[259])|(m[6]&~m[256]&~m[257]&m[258]&m[259])|(~m[6]&m[256]&~m[257]&m[258]&m[259])|(~m[6]&~m[256]&m[257]&m[258]&m[259]))&~BiasedRNG[280])|((m[6]&m[256]&m[257]&m[258]&~m[259])|(m[6]&m[256]&m[257]&~m[258]&m[259])|(m[6]&m[256]&~m[257]&m[258]&m[259])|(m[6]&~m[256]&m[257]&m[258]&m[259])|(~m[6]&m[256]&m[257]&m[258]&m[259])|(m[6]&m[256]&m[257]&m[258]&m[259]));
    m[57] = (((m[6]&m[260]&~m[261]&~m[262]&~m[263])|(m[6]&~m[260]&m[261]&~m[262]&~m[263])|(~m[6]&m[260]&m[261]&~m[262]&~m[263])|(m[6]&~m[260]&~m[261]&m[262]&~m[263])|(~m[6]&m[260]&~m[261]&m[262]&~m[263])|(~m[6]&~m[260]&m[261]&m[262]&~m[263])|(m[6]&~m[260]&~m[261]&~m[262]&m[263])|(~m[6]&m[260]&~m[261]&~m[262]&m[263])|(~m[6]&~m[260]&m[261]&~m[262]&m[263])|(~m[6]&~m[260]&~m[261]&m[262]&m[263]))&BiasedRNG[281])|(((m[6]&m[260]&m[261]&~m[262]&~m[263])|(m[6]&m[260]&~m[261]&m[262]&~m[263])|(m[6]&~m[260]&m[261]&m[262]&~m[263])|(~m[6]&m[260]&m[261]&m[262]&~m[263])|(m[6]&m[260]&~m[261]&~m[262]&m[263])|(m[6]&~m[260]&m[261]&~m[262]&m[263])|(~m[6]&m[260]&m[261]&~m[262]&m[263])|(m[6]&~m[260]&~m[261]&m[262]&m[263])|(~m[6]&m[260]&~m[261]&m[262]&m[263])|(~m[6]&~m[260]&m[261]&m[262]&m[263]))&~BiasedRNG[281])|((m[6]&m[260]&m[261]&m[262]&~m[263])|(m[6]&m[260]&m[261]&~m[262]&m[263])|(m[6]&m[260]&~m[261]&m[262]&m[263])|(m[6]&~m[260]&m[261]&m[262]&m[263])|(~m[6]&m[260]&m[261]&m[262]&m[263])|(m[6]&m[260]&m[261]&m[262]&m[263]));
    m[58] = (((m[6]&m[264]&~m[265]&~m[266]&~m[267])|(m[6]&~m[264]&m[265]&~m[266]&~m[267])|(~m[6]&m[264]&m[265]&~m[266]&~m[267])|(m[6]&~m[264]&~m[265]&m[266]&~m[267])|(~m[6]&m[264]&~m[265]&m[266]&~m[267])|(~m[6]&~m[264]&m[265]&m[266]&~m[267])|(m[6]&~m[264]&~m[265]&~m[266]&m[267])|(~m[6]&m[264]&~m[265]&~m[266]&m[267])|(~m[6]&~m[264]&m[265]&~m[266]&m[267])|(~m[6]&~m[264]&~m[265]&m[266]&m[267]))&BiasedRNG[282])|(((m[6]&m[264]&m[265]&~m[266]&~m[267])|(m[6]&m[264]&~m[265]&m[266]&~m[267])|(m[6]&~m[264]&m[265]&m[266]&~m[267])|(~m[6]&m[264]&m[265]&m[266]&~m[267])|(m[6]&m[264]&~m[265]&~m[266]&m[267])|(m[6]&~m[264]&m[265]&~m[266]&m[267])|(~m[6]&m[264]&m[265]&~m[266]&m[267])|(m[6]&~m[264]&~m[265]&m[266]&m[267])|(~m[6]&m[264]&~m[265]&m[266]&m[267])|(~m[6]&~m[264]&m[265]&m[266]&m[267]))&~BiasedRNG[282])|((m[6]&m[264]&m[265]&m[266]&~m[267])|(m[6]&m[264]&m[265]&~m[266]&m[267])|(m[6]&m[264]&~m[265]&m[266]&m[267])|(m[6]&~m[264]&m[265]&m[266]&m[267])|(~m[6]&m[264]&m[265]&m[266]&m[267])|(m[6]&m[264]&m[265]&m[266]&m[267]));
    m[59] = (((m[6]&m[268]&~m[269]&~m[270]&~m[271])|(m[6]&~m[268]&m[269]&~m[270]&~m[271])|(~m[6]&m[268]&m[269]&~m[270]&~m[271])|(m[6]&~m[268]&~m[269]&m[270]&~m[271])|(~m[6]&m[268]&~m[269]&m[270]&~m[271])|(~m[6]&~m[268]&m[269]&m[270]&~m[271])|(m[6]&~m[268]&~m[269]&~m[270]&m[271])|(~m[6]&m[268]&~m[269]&~m[270]&m[271])|(~m[6]&~m[268]&m[269]&~m[270]&m[271])|(~m[6]&~m[268]&~m[269]&m[270]&m[271]))&BiasedRNG[283])|(((m[6]&m[268]&m[269]&~m[270]&~m[271])|(m[6]&m[268]&~m[269]&m[270]&~m[271])|(m[6]&~m[268]&m[269]&m[270]&~m[271])|(~m[6]&m[268]&m[269]&m[270]&~m[271])|(m[6]&m[268]&~m[269]&~m[270]&m[271])|(m[6]&~m[268]&m[269]&~m[270]&m[271])|(~m[6]&m[268]&m[269]&~m[270]&m[271])|(m[6]&~m[268]&~m[269]&m[270]&m[271])|(~m[6]&m[268]&~m[269]&m[270]&m[271])|(~m[6]&~m[268]&m[269]&m[270]&m[271]))&~BiasedRNG[283])|((m[6]&m[268]&m[269]&m[270]&~m[271])|(m[6]&m[268]&m[269]&~m[270]&m[271])|(m[6]&m[268]&~m[269]&m[270]&m[271])|(m[6]&~m[268]&m[269]&m[270]&m[271])|(~m[6]&m[268]&m[269]&m[270]&m[271])|(m[6]&m[268]&m[269]&m[270]&m[271]));
    m[60] = (((m[7]&m[272]&~m[273]&~m[274]&~m[275])|(m[7]&~m[272]&m[273]&~m[274]&~m[275])|(~m[7]&m[272]&m[273]&~m[274]&~m[275])|(m[7]&~m[272]&~m[273]&m[274]&~m[275])|(~m[7]&m[272]&~m[273]&m[274]&~m[275])|(~m[7]&~m[272]&m[273]&m[274]&~m[275])|(m[7]&~m[272]&~m[273]&~m[274]&m[275])|(~m[7]&m[272]&~m[273]&~m[274]&m[275])|(~m[7]&~m[272]&m[273]&~m[274]&m[275])|(~m[7]&~m[272]&~m[273]&m[274]&m[275]))&BiasedRNG[284])|(((m[7]&m[272]&m[273]&~m[274]&~m[275])|(m[7]&m[272]&~m[273]&m[274]&~m[275])|(m[7]&~m[272]&m[273]&m[274]&~m[275])|(~m[7]&m[272]&m[273]&m[274]&~m[275])|(m[7]&m[272]&~m[273]&~m[274]&m[275])|(m[7]&~m[272]&m[273]&~m[274]&m[275])|(~m[7]&m[272]&m[273]&~m[274]&m[275])|(m[7]&~m[272]&~m[273]&m[274]&m[275])|(~m[7]&m[272]&~m[273]&m[274]&m[275])|(~m[7]&~m[272]&m[273]&m[274]&m[275]))&~BiasedRNG[284])|((m[7]&m[272]&m[273]&m[274]&~m[275])|(m[7]&m[272]&m[273]&~m[274]&m[275])|(m[7]&m[272]&~m[273]&m[274]&m[275])|(m[7]&~m[272]&m[273]&m[274]&m[275])|(~m[7]&m[272]&m[273]&m[274]&m[275])|(m[7]&m[272]&m[273]&m[274]&m[275]));
    m[61] = (((m[7]&m[276]&~m[277]&~m[278]&~m[279])|(m[7]&~m[276]&m[277]&~m[278]&~m[279])|(~m[7]&m[276]&m[277]&~m[278]&~m[279])|(m[7]&~m[276]&~m[277]&m[278]&~m[279])|(~m[7]&m[276]&~m[277]&m[278]&~m[279])|(~m[7]&~m[276]&m[277]&m[278]&~m[279])|(m[7]&~m[276]&~m[277]&~m[278]&m[279])|(~m[7]&m[276]&~m[277]&~m[278]&m[279])|(~m[7]&~m[276]&m[277]&~m[278]&m[279])|(~m[7]&~m[276]&~m[277]&m[278]&m[279]))&BiasedRNG[285])|(((m[7]&m[276]&m[277]&~m[278]&~m[279])|(m[7]&m[276]&~m[277]&m[278]&~m[279])|(m[7]&~m[276]&m[277]&m[278]&~m[279])|(~m[7]&m[276]&m[277]&m[278]&~m[279])|(m[7]&m[276]&~m[277]&~m[278]&m[279])|(m[7]&~m[276]&m[277]&~m[278]&m[279])|(~m[7]&m[276]&m[277]&~m[278]&m[279])|(m[7]&~m[276]&~m[277]&m[278]&m[279])|(~m[7]&m[276]&~m[277]&m[278]&m[279])|(~m[7]&~m[276]&m[277]&m[278]&m[279]))&~BiasedRNG[285])|((m[7]&m[276]&m[277]&m[278]&~m[279])|(m[7]&m[276]&m[277]&~m[278]&m[279])|(m[7]&m[276]&~m[277]&m[278]&m[279])|(m[7]&~m[276]&m[277]&m[278]&m[279])|(~m[7]&m[276]&m[277]&m[278]&m[279])|(m[7]&m[276]&m[277]&m[278]&m[279]));
    m[62] = (((m[7]&m[280]&~m[281]&~m[282]&~m[283])|(m[7]&~m[280]&m[281]&~m[282]&~m[283])|(~m[7]&m[280]&m[281]&~m[282]&~m[283])|(m[7]&~m[280]&~m[281]&m[282]&~m[283])|(~m[7]&m[280]&~m[281]&m[282]&~m[283])|(~m[7]&~m[280]&m[281]&m[282]&~m[283])|(m[7]&~m[280]&~m[281]&~m[282]&m[283])|(~m[7]&m[280]&~m[281]&~m[282]&m[283])|(~m[7]&~m[280]&m[281]&~m[282]&m[283])|(~m[7]&~m[280]&~m[281]&m[282]&m[283]))&BiasedRNG[286])|(((m[7]&m[280]&m[281]&~m[282]&~m[283])|(m[7]&m[280]&~m[281]&m[282]&~m[283])|(m[7]&~m[280]&m[281]&m[282]&~m[283])|(~m[7]&m[280]&m[281]&m[282]&~m[283])|(m[7]&m[280]&~m[281]&~m[282]&m[283])|(m[7]&~m[280]&m[281]&~m[282]&m[283])|(~m[7]&m[280]&m[281]&~m[282]&m[283])|(m[7]&~m[280]&~m[281]&m[282]&m[283])|(~m[7]&m[280]&~m[281]&m[282]&m[283])|(~m[7]&~m[280]&m[281]&m[282]&m[283]))&~BiasedRNG[286])|((m[7]&m[280]&m[281]&m[282]&~m[283])|(m[7]&m[280]&m[281]&~m[282]&m[283])|(m[7]&m[280]&~m[281]&m[282]&m[283])|(m[7]&~m[280]&m[281]&m[282]&m[283])|(~m[7]&m[280]&m[281]&m[282]&m[283])|(m[7]&m[280]&m[281]&m[282]&m[283]));
    m[63] = (((m[7]&m[284]&~m[285]&~m[286]&~m[287])|(m[7]&~m[284]&m[285]&~m[286]&~m[287])|(~m[7]&m[284]&m[285]&~m[286]&~m[287])|(m[7]&~m[284]&~m[285]&m[286]&~m[287])|(~m[7]&m[284]&~m[285]&m[286]&~m[287])|(~m[7]&~m[284]&m[285]&m[286]&~m[287])|(m[7]&~m[284]&~m[285]&~m[286]&m[287])|(~m[7]&m[284]&~m[285]&~m[286]&m[287])|(~m[7]&~m[284]&m[285]&~m[286]&m[287])|(~m[7]&~m[284]&~m[285]&m[286]&m[287]))&BiasedRNG[287])|(((m[7]&m[284]&m[285]&~m[286]&~m[287])|(m[7]&m[284]&~m[285]&m[286]&~m[287])|(m[7]&~m[284]&m[285]&m[286]&~m[287])|(~m[7]&m[284]&m[285]&m[286]&~m[287])|(m[7]&m[284]&~m[285]&~m[286]&m[287])|(m[7]&~m[284]&m[285]&~m[286]&m[287])|(~m[7]&m[284]&m[285]&~m[286]&m[287])|(m[7]&~m[284]&~m[285]&m[286]&m[287])|(~m[7]&m[284]&~m[285]&m[286]&m[287])|(~m[7]&~m[284]&m[285]&m[286]&m[287]))&~BiasedRNG[287])|((m[7]&m[284]&m[285]&m[286]&~m[287])|(m[7]&m[284]&m[285]&~m[286]&m[287])|(m[7]&m[284]&~m[285]&m[286]&m[287])|(m[7]&~m[284]&m[285]&m[286]&m[287])|(~m[7]&m[284]&m[285]&m[286]&m[287])|(m[7]&m[284]&m[285]&m[286]&m[287]));
    m[64] = (((m[8]&m[288]&~m[289]&~m[290]&~m[291])|(m[8]&~m[288]&m[289]&~m[290]&~m[291])|(~m[8]&m[288]&m[289]&~m[290]&~m[291])|(m[8]&~m[288]&~m[289]&m[290]&~m[291])|(~m[8]&m[288]&~m[289]&m[290]&~m[291])|(~m[8]&~m[288]&m[289]&m[290]&~m[291])|(m[8]&~m[288]&~m[289]&~m[290]&m[291])|(~m[8]&m[288]&~m[289]&~m[290]&m[291])|(~m[8]&~m[288]&m[289]&~m[290]&m[291])|(~m[8]&~m[288]&~m[289]&m[290]&m[291]))&BiasedRNG[288])|(((m[8]&m[288]&m[289]&~m[290]&~m[291])|(m[8]&m[288]&~m[289]&m[290]&~m[291])|(m[8]&~m[288]&m[289]&m[290]&~m[291])|(~m[8]&m[288]&m[289]&m[290]&~m[291])|(m[8]&m[288]&~m[289]&~m[290]&m[291])|(m[8]&~m[288]&m[289]&~m[290]&m[291])|(~m[8]&m[288]&m[289]&~m[290]&m[291])|(m[8]&~m[288]&~m[289]&m[290]&m[291])|(~m[8]&m[288]&~m[289]&m[290]&m[291])|(~m[8]&~m[288]&m[289]&m[290]&m[291]))&~BiasedRNG[288])|((m[8]&m[288]&m[289]&m[290]&~m[291])|(m[8]&m[288]&m[289]&~m[290]&m[291])|(m[8]&m[288]&~m[289]&m[290]&m[291])|(m[8]&~m[288]&m[289]&m[290]&m[291])|(~m[8]&m[288]&m[289]&m[290]&m[291])|(m[8]&m[288]&m[289]&m[290]&m[291]));
    m[65] = (((m[8]&m[292]&~m[293]&~m[294]&~m[295])|(m[8]&~m[292]&m[293]&~m[294]&~m[295])|(~m[8]&m[292]&m[293]&~m[294]&~m[295])|(m[8]&~m[292]&~m[293]&m[294]&~m[295])|(~m[8]&m[292]&~m[293]&m[294]&~m[295])|(~m[8]&~m[292]&m[293]&m[294]&~m[295])|(m[8]&~m[292]&~m[293]&~m[294]&m[295])|(~m[8]&m[292]&~m[293]&~m[294]&m[295])|(~m[8]&~m[292]&m[293]&~m[294]&m[295])|(~m[8]&~m[292]&~m[293]&m[294]&m[295]))&BiasedRNG[289])|(((m[8]&m[292]&m[293]&~m[294]&~m[295])|(m[8]&m[292]&~m[293]&m[294]&~m[295])|(m[8]&~m[292]&m[293]&m[294]&~m[295])|(~m[8]&m[292]&m[293]&m[294]&~m[295])|(m[8]&m[292]&~m[293]&~m[294]&m[295])|(m[8]&~m[292]&m[293]&~m[294]&m[295])|(~m[8]&m[292]&m[293]&~m[294]&m[295])|(m[8]&~m[292]&~m[293]&m[294]&m[295])|(~m[8]&m[292]&~m[293]&m[294]&m[295])|(~m[8]&~m[292]&m[293]&m[294]&m[295]))&~BiasedRNG[289])|((m[8]&m[292]&m[293]&m[294]&~m[295])|(m[8]&m[292]&m[293]&~m[294]&m[295])|(m[8]&m[292]&~m[293]&m[294]&m[295])|(m[8]&~m[292]&m[293]&m[294]&m[295])|(~m[8]&m[292]&m[293]&m[294]&m[295])|(m[8]&m[292]&m[293]&m[294]&m[295]));
    m[66] = (((m[8]&m[296]&~m[297]&~m[298]&~m[299])|(m[8]&~m[296]&m[297]&~m[298]&~m[299])|(~m[8]&m[296]&m[297]&~m[298]&~m[299])|(m[8]&~m[296]&~m[297]&m[298]&~m[299])|(~m[8]&m[296]&~m[297]&m[298]&~m[299])|(~m[8]&~m[296]&m[297]&m[298]&~m[299])|(m[8]&~m[296]&~m[297]&~m[298]&m[299])|(~m[8]&m[296]&~m[297]&~m[298]&m[299])|(~m[8]&~m[296]&m[297]&~m[298]&m[299])|(~m[8]&~m[296]&~m[297]&m[298]&m[299]))&BiasedRNG[290])|(((m[8]&m[296]&m[297]&~m[298]&~m[299])|(m[8]&m[296]&~m[297]&m[298]&~m[299])|(m[8]&~m[296]&m[297]&m[298]&~m[299])|(~m[8]&m[296]&m[297]&m[298]&~m[299])|(m[8]&m[296]&~m[297]&~m[298]&m[299])|(m[8]&~m[296]&m[297]&~m[298]&m[299])|(~m[8]&m[296]&m[297]&~m[298]&m[299])|(m[8]&~m[296]&~m[297]&m[298]&m[299])|(~m[8]&m[296]&~m[297]&m[298]&m[299])|(~m[8]&~m[296]&m[297]&m[298]&m[299]))&~BiasedRNG[290])|((m[8]&m[296]&m[297]&m[298]&~m[299])|(m[8]&m[296]&m[297]&~m[298]&m[299])|(m[8]&m[296]&~m[297]&m[298]&m[299])|(m[8]&~m[296]&m[297]&m[298]&m[299])|(~m[8]&m[296]&m[297]&m[298]&m[299])|(m[8]&m[296]&m[297]&m[298]&m[299]));
    m[67] = (((m[8]&m[300]&~m[301]&~m[302]&~m[303])|(m[8]&~m[300]&m[301]&~m[302]&~m[303])|(~m[8]&m[300]&m[301]&~m[302]&~m[303])|(m[8]&~m[300]&~m[301]&m[302]&~m[303])|(~m[8]&m[300]&~m[301]&m[302]&~m[303])|(~m[8]&~m[300]&m[301]&m[302]&~m[303])|(m[8]&~m[300]&~m[301]&~m[302]&m[303])|(~m[8]&m[300]&~m[301]&~m[302]&m[303])|(~m[8]&~m[300]&m[301]&~m[302]&m[303])|(~m[8]&~m[300]&~m[301]&m[302]&m[303]))&BiasedRNG[291])|(((m[8]&m[300]&m[301]&~m[302]&~m[303])|(m[8]&m[300]&~m[301]&m[302]&~m[303])|(m[8]&~m[300]&m[301]&m[302]&~m[303])|(~m[8]&m[300]&m[301]&m[302]&~m[303])|(m[8]&m[300]&~m[301]&~m[302]&m[303])|(m[8]&~m[300]&m[301]&~m[302]&m[303])|(~m[8]&m[300]&m[301]&~m[302]&m[303])|(m[8]&~m[300]&~m[301]&m[302]&m[303])|(~m[8]&m[300]&~m[301]&m[302]&m[303])|(~m[8]&~m[300]&m[301]&m[302]&m[303]))&~BiasedRNG[291])|((m[8]&m[300]&m[301]&m[302]&~m[303])|(m[8]&m[300]&m[301]&~m[302]&m[303])|(m[8]&m[300]&~m[301]&m[302]&m[303])|(m[8]&~m[300]&m[301]&m[302]&m[303])|(~m[8]&m[300]&m[301]&m[302]&m[303])|(m[8]&m[300]&m[301]&m[302]&m[303]));
    m[68] = (((m[9]&m[304]&~m[305]&~m[306]&~m[307])|(m[9]&~m[304]&m[305]&~m[306]&~m[307])|(~m[9]&m[304]&m[305]&~m[306]&~m[307])|(m[9]&~m[304]&~m[305]&m[306]&~m[307])|(~m[9]&m[304]&~m[305]&m[306]&~m[307])|(~m[9]&~m[304]&m[305]&m[306]&~m[307])|(m[9]&~m[304]&~m[305]&~m[306]&m[307])|(~m[9]&m[304]&~m[305]&~m[306]&m[307])|(~m[9]&~m[304]&m[305]&~m[306]&m[307])|(~m[9]&~m[304]&~m[305]&m[306]&m[307]))&BiasedRNG[292])|(((m[9]&m[304]&m[305]&~m[306]&~m[307])|(m[9]&m[304]&~m[305]&m[306]&~m[307])|(m[9]&~m[304]&m[305]&m[306]&~m[307])|(~m[9]&m[304]&m[305]&m[306]&~m[307])|(m[9]&m[304]&~m[305]&~m[306]&m[307])|(m[9]&~m[304]&m[305]&~m[306]&m[307])|(~m[9]&m[304]&m[305]&~m[306]&m[307])|(m[9]&~m[304]&~m[305]&m[306]&m[307])|(~m[9]&m[304]&~m[305]&m[306]&m[307])|(~m[9]&~m[304]&m[305]&m[306]&m[307]))&~BiasedRNG[292])|((m[9]&m[304]&m[305]&m[306]&~m[307])|(m[9]&m[304]&m[305]&~m[306]&m[307])|(m[9]&m[304]&~m[305]&m[306]&m[307])|(m[9]&~m[304]&m[305]&m[306]&m[307])|(~m[9]&m[304]&m[305]&m[306]&m[307])|(m[9]&m[304]&m[305]&m[306]&m[307]));
    m[69] = (((m[9]&m[308]&~m[309]&~m[310]&~m[311])|(m[9]&~m[308]&m[309]&~m[310]&~m[311])|(~m[9]&m[308]&m[309]&~m[310]&~m[311])|(m[9]&~m[308]&~m[309]&m[310]&~m[311])|(~m[9]&m[308]&~m[309]&m[310]&~m[311])|(~m[9]&~m[308]&m[309]&m[310]&~m[311])|(m[9]&~m[308]&~m[309]&~m[310]&m[311])|(~m[9]&m[308]&~m[309]&~m[310]&m[311])|(~m[9]&~m[308]&m[309]&~m[310]&m[311])|(~m[9]&~m[308]&~m[309]&m[310]&m[311]))&BiasedRNG[293])|(((m[9]&m[308]&m[309]&~m[310]&~m[311])|(m[9]&m[308]&~m[309]&m[310]&~m[311])|(m[9]&~m[308]&m[309]&m[310]&~m[311])|(~m[9]&m[308]&m[309]&m[310]&~m[311])|(m[9]&m[308]&~m[309]&~m[310]&m[311])|(m[9]&~m[308]&m[309]&~m[310]&m[311])|(~m[9]&m[308]&m[309]&~m[310]&m[311])|(m[9]&~m[308]&~m[309]&m[310]&m[311])|(~m[9]&m[308]&~m[309]&m[310]&m[311])|(~m[9]&~m[308]&m[309]&m[310]&m[311]))&~BiasedRNG[293])|((m[9]&m[308]&m[309]&m[310]&~m[311])|(m[9]&m[308]&m[309]&~m[310]&m[311])|(m[9]&m[308]&~m[309]&m[310]&m[311])|(m[9]&~m[308]&m[309]&m[310]&m[311])|(~m[9]&m[308]&m[309]&m[310]&m[311])|(m[9]&m[308]&m[309]&m[310]&m[311]));
    m[70] = (((m[9]&m[312]&~m[313]&~m[314]&~m[315])|(m[9]&~m[312]&m[313]&~m[314]&~m[315])|(~m[9]&m[312]&m[313]&~m[314]&~m[315])|(m[9]&~m[312]&~m[313]&m[314]&~m[315])|(~m[9]&m[312]&~m[313]&m[314]&~m[315])|(~m[9]&~m[312]&m[313]&m[314]&~m[315])|(m[9]&~m[312]&~m[313]&~m[314]&m[315])|(~m[9]&m[312]&~m[313]&~m[314]&m[315])|(~m[9]&~m[312]&m[313]&~m[314]&m[315])|(~m[9]&~m[312]&~m[313]&m[314]&m[315]))&BiasedRNG[294])|(((m[9]&m[312]&m[313]&~m[314]&~m[315])|(m[9]&m[312]&~m[313]&m[314]&~m[315])|(m[9]&~m[312]&m[313]&m[314]&~m[315])|(~m[9]&m[312]&m[313]&m[314]&~m[315])|(m[9]&m[312]&~m[313]&~m[314]&m[315])|(m[9]&~m[312]&m[313]&~m[314]&m[315])|(~m[9]&m[312]&m[313]&~m[314]&m[315])|(m[9]&~m[312]&~m[313]&m[314]&m[315])|(~m[9]&m[312]&~m[313]&m[314]&m[315])|(~m[9]&~m[312]&m[313]&m[314]&m[315]))&~BiasedRNG[294])|((m[9]&m[312]&m[313]&m[314]&~m[315])|(m[9]&m[312]&m[313]&~m[314]&m[315])|(m[9]&m[312]&~m[313]&m[314]&m[315])|(m[9]&~m[312]&m[313]&m[314]&m[315])|(~m[9]&m[312]&m[313]&m[314]&m[315])|(m[9]&m[312]&m[313]&m[314]&m[315]));
    m[71] = (((m[9]&m[316]&~m[317]&~m[318]&~m[319])|(m[9]&~m[316]&m[317]&~m[318]&~m[319])|(~m[9]&m[316]&m[317]&~m[318]&~m[319])|(m[9]&~m[316]&~m[317]&m[318]&~m[319])|(~m[9]&m[316]&~m[317]&m[318]&~m[319])|(~m[9]&~m[316]&m[317]&m[318]&~m[319])|(m[9]&~m[316]&~m[317]&~m[318]&m[319])|(~m[9]&m[316]&~m[317]&~m[318]&m[319])|(~m[9]&~m[316]&m[317]&~m[318]&m[319])|(~m[9]&~m[316]&~m[317]&m[318]&m[319]))&BiasedRNG[295])|(((m[9]&m[316]&m[317]&~m[318]&~m[319])|(m[9]&m[316]&~m[317]&m[318]&~m[319])|(m[9]&~m[316]&m[317]&m[318]&~m[319])|(~m[9]&m[316]&m[317]&m[318]&~m[319])|(m[9]&m[316]&~m[317]&~m[318]&m[319])|(m[9]&~m[316]&m[317]&~m[318]&m[319])|(~m[9]&m[316]&m[317]&~m[318]&m[319])|(m[9]&~m[316]&~m[317]&m[318]&m[319])|(~m[9]&m[316]&~m[317]&m[318]&m[319])|(~m[9]&~m[316]&m[317]&m[318]&m[319]))&~BiasedRNG[295])|((m[9]&m[316]&m[317]&m[318]&~m[319])|(m[9]&m[316]&m[317]&~m[318]&m[319])|(m[9]&m[316]&~m[317]&m[318]&m[319])|(m[9]&~m[316]&m[317]&m[318]&m[319])|(~m[9]&m[316]&m[317]&m[318]&m[319])|(m[9]&m[316]&m[317]&m[318]&m[319]));
    m[72] = (((m[10]&m[320]&~m[321]&~m[322]&~m[323])|(m[10]&~m[320]&m[321]&~m[322]&~m[323])|(~m[10]&m[320]&m[321]&~m[322]&~m[323])|(m[10]&~m[320]&~m[321]&m[322]&~m[323])|(~m[10]&m[320]&~m[321]&m[322]&~m[323])|(~m[10]&~m[320]&m[321]&m[322]&~m[323])|(m[10]&~m[320]&~m[321]&~m[322]&m[323])|(~m[10]&m[320]&~m[321]&~m[322]&m[323])|(~m[10]&~m[320]&m[321]&~m[322]&m[323])|(~m[10]&~m[320]&~m[321]&m[322]&m[323]))&BiasedRNG[296])|(((m[10]&m[320]&m[321]&~m[322]&~m[323])|(m[10]&m[320]&~m[321]&m[322]&~m[323])|(m[10]&~m[320]&m[321]&m[322]&~m[323])|(~m[10]&m[320]&m[321]&m[322]&~m[323])|(m[10]&m[320]&~m[321]&~m[322]&m[323])|(m[10]&~m[320]&m[321]&~m[322]&m[323])|(~m[10]&m[320]&m[321]&~m[322]&m[323])|(m[10]&~m[320]&~m[321]&m[322]&m[323])|(~m[10]&m[320]&~m[321]&m[322]&m[323])|(~m[10]&~m[320]&m[321]&m[322]&m[323]))&~BiasedRNG[296])|((m[10]&m[320]&m[321]&m[322]&~m[323])|(m[10]&m[320]&m[321]&~m[322]&m[323])|(m[10]&m[320]&~m[321]&m[322]&m[323])|(m[10]&~m[320]&m[321]&m[322]&m[323])|(~m[10]&m[320]&m[321]&m[322]&m[323])|(m[10]&m[320]&m[321]&m[322]&m[323]));
    m[73] = (((m[10]&m[324]&~m[325]&~m[326]&~m[327])|(m[10]&~m[324]&m[325]&~m[326]&~m[327])|(~m[10]&m[324]&m[325]&~m[326]&~m[327])|(m[10]&~m[324]&~m[325]&m[326]&~m[327])|(~m[10]&m[324]&~m[325]&m[326]&~m[327])|(~m[10]&~m[324]&m[325]&m[326]&~m[327])|(m[10]&~m[324]&~m[325]&~m[326]&m[327])|(~m[10]&m[324]&~m[325]&~m[326]&m[327])|(~m[10]&~m[324]&m[325]&~m[326]&m[327])|(~m[10]&~m[324]&~m[325]&m[326]&m[327]))&BiasedRNG[297])|(((m[10]&m[324]&m[325]&~m[326]&~m[327])|(m[10]&m[324]&~m[325]&m[326]&~m[327])|(m[10]&~m[324]&m[325]&m[326]&~m[327])|(~m[10]&m[324]&m[325]&m[326]&~m[327])|(m[10]&m[324]&~m[325]&~m[326]&m[327])|(m[10]&~m[324]&m[325]&~m[326]&m[327])|(~m[10]&m[324]&m[325]&~m[326]&m[327])|(m[10]&~m[324]&~m[325]&m[326]&m[327])|(~m[10]&m[324]&~m[325]&m[326]&m[327])|(~m[10]&~m[324]&m[325]&m[326]&m[327]))&~BiasedRNG[297])|((m[10]&m[324]&m[325]&m[326]&~m[327])|(m[10]&m[324]&m[325]&~m[326]&m[327])|(m[10]&m[324]&~m[325]&m[326]&m[327])|(m[10]&~m[324]&m[325]&m[326]&m[327])|(~m[10]&m[324]&m[325]&m[326]&m[327])|(m[10]&m[324]&m[325]&m[326]&m[327]));
    m[74] = (((m[10]&m[328]&~m[329]&~m[330]&~m[331])|(m[10]&~m[328]&m[329]&~m[330]&~m[331])|(~m[10]&m[328]&m[329]&~m[330]&~m[331])|(m[10]&~m[328]&~m[329]&m[330]&~m[331])|(~m[10]&m[328]&~m[329]&m[330]&~m[331])|(~m[10]&~m[328]&m[329]&m[330]&~m[331])|(m[10]&~m[328]&~m[329]&~m[330]&m[331])|(~m[10]&m[328]&~m[329]&~m[330]&m[331])|(~m[10]&~m[328]&m[329]&~m[330]&m[331])|(~m[10]&~m[328]&~m[329]&m[330]&m[331]))&BiasedRNG[298])|(((m[10]&m[328]&m[329]&~m[330]&~m[331])|(m[10]&m[328]&~m[329]&m[330]&~m[331])|(m[10]&~m[328]&m[329]&m[330]&~m[331])|(~m[10]&m[328]&m[329]&m[330]&~m[331])|(m[10]&m[328]&~m[329]&~m[330]&m[331])|(m[10]&~m[328]&m[329]&~m[330]&m[331])|(~m[10]&m[328]&m[329]&~m[330]&m[331])|(m[10]&~m[328]&~m[329]&m[330]&m[331])|(~m[10]&m[328]&~m[329]&m[330]&m[331])|(~m[10]&~m[328]&m[329]&m[330]&m[331]))&~BiasedRNG[298])|((m[10]&m[328]&m[329]&m[330]&~m[331])|(m[10]&m[328]&m[329]&~m[330]&m[331])|(m[10]&m[328]&~m[329]&m[330]&m[331])|(m[10]&~m[328]&m[329]&m[330]&m[331])|(~m[10]&m[328]&m[329]&m[330]&m[331])|(m[10]&m[328]&m[329]&m[330]&m[331]));
    m[75] = (((m[10]&m[332]&~m[333]&~m[334]&~m[335])|(m[10]&~m[332]&m[333]&~m[334]&~m[335])|(~m[10]&m[332]&m[333]&~m[334]&~m[335])|(m[10]&~m[332]&~m[333]&m[334]&~m[335])|(~m[10]&m[332]&~m[333]&m[334]&~m[335])|(~m[10]&~m[332]&m[333]&m[334]&~m[335])|(m[10]&~m[332]&~m[333]&~m[334]&m[335])|(~m[10]&m[332]&~m[333]&~m[334]&m[335])|(~m[10]&~m[332]&m[333]&~m[334]&m[335])|(~m[10]&~m[332]&~m[333]&m[334]&m[335]))&BiasedRNG[299])|(((m[10]&m[332]&m[333]&~m[334]&~m[335])|(m[10]&m[332]&~m[333]&m[334]&~m[335])|(m[10]&~m[332]&m[333]&m[334]&~m[335])|(~m[10]&m[332]&m[333]&m[334]&~m[335])|(m[10]&m[332]&~m[333]&~m[334]&m[335])|(m[10]&~m[332]&m[333]&~m[334]&m[335])|(~m[10]&m[332]&m[333]&~m[334]&m[335])|(m[10]&~m[332]&~m[333]&m[334]&m[335])|(~m[10]&m[332]&~m[333]&m[334]&m[335])|(~m[10]&~m[332]&m[333]&m[334]&m[335]))&~BiasedRNG[299])|((m[10]&m[332]&m[333]&m[334]&~m[335])|(m[10]&m[332]&m[333]&~m[334]&m[335])|(m[10]&m[332]&~m[333]&m[334]&m[335])|(m[10]&~m[332]&m[333]&m[334]&m[335])|(~m[10]&m[332]&m[333]&m[334]&m[335])|(m[10]&m[332]&m[333]&m[334]&m[335]));
    m[76] = (((m[11]&m[336]&~m[337]&~m[338]&~m[339])|(m[11]&~m[336]&m[337]&~m[338]&~m[339])|(~m[11]&m[336]&m[337]&~m[338]&~m[339])|(m[11]&~m[336]&~m[337]&m[338]&~m[339])|(~m[11]&m[336]&~m[337]&m[338]&~m[339])|(~m[11]&~m[336]&m[337]&m[338]&~m[339])|(m[11]&~m[336]&~m[337]&~m[338]&m[339])|(~m[11]&m[336]&~m[337]&~m[338]&m[339])|(~m[11]&~m[336]&m[337]&~m[338]&m[339])|(~m[11]&~m[336]&~m[337]&m[338]&m[339]))&BiasedRNG[300])|(((m[11]&m[336]&m[337]&~m[338]&~m[339])|(m[11]&m[336]&~m[337]&m[338]&~m[339])|(m[11]&~m[336]&m[337]&m[338]&~m[339])|(~m[11]&m[336]&m[337]&m[338]&~m[339])|(m[11]&m[336]&~m[337]&~m[338]&m[339])|(m[11]&~m[336]&m[337]&~m[338]&m[339])|(~m[11]&m[336]&m[337]&~m[338]&m[339])|(m[11]&~m[336]&~m[337]&m[338]&m[339])|(~m[11]&m[336]&~m[337]&m[338]&m[339])|(~m[11]&~m[336]&m[337]&m[338]&m[339]))&~BiasedRNG[300])|((m[11]&m[336]&m[337]&m[338]&~m[339])|(m[11]&m[336]&m[337]&~m[338]&m[339])|(m[11]&m[336]&~m[337]&m[338]&m[339])|(m[11]&~m[336]&m[337]&m[338]&m[339])|(~m[11]&m[336]&m[337]&m[338]&m[339])|(m[11]&m[336]&m[337]&m[338]&m[339]));
    m[77] = (((m[11]&m[340]&~m[341]&~m[342]&~m[343])|(m[11]&~m[340]&m[341]&~m[342]&~m[343])|(~m[11]&m[340]&m[341]&~m[342]&~m[343])|(m[11]&~m[340]&~m[341]&m[342]&~m[343])|(~m[11]&m[340]&~m[341]&m[342]&~m[343])|(~m[11]&~m[340]&m[341]&m[342]&~m[343])|(m[11]&~m[340]&~m[341]&~m[342]&m[343])|(~m[11]&m[340]&~m[341]&~m[342]&m[343])|(~m[11]&~m[340]&m[341]&~m[342]&m[343])|(~m[11]&~m[340]&~m[341]&m[342]&m[343]))&BiasedRNG[301])|(((m[11]&m[340]&m[341]&~m[342]&~m[343])|(m[11]&m[340]&~m[341]&m[342]&~m[343])|(m[11]&~m[340]&m[341]&m[342]&~m[343])|(~m[11]&m[340]&m[341]&m[342]&~m[343])|(m[11]&m[340]&~m[341]&~m[342]&m[343])|(m[11]&~m[340]&m[341]&~m[342]&m[343])|(~m[11]&m[340]&m[341]&~m[342]&m[343])|(m[11]&~m[340]&~m[341]&m[342]&m[343])|(~m[11]&m[340]&~m[341]&m[342]&m[343])|(~m[11]&~m[340]&m[341]&m[342]&m[343]))&~BiasedRNG[301])|((m[11]&m[340]&m[341]&m[342]&~m[343])|(m[11]&m[340]&m[341]&~m[342]&m[343])|(m[11]&m[340]&~m[341]&m[342]&m[343])|(m[11]&~m[340]&m[341]&m[342]&m[343])|(~m[11]&m[340]&m[341]&m[342]&m[343])|(m[11]&m[340]&m[341]&m[342]&m[343]));
    m[78] = (((m[11]&m[344]&~m[345]&~m[346]&~m[347])|(m[11]&~m[344]&m[345]&~m[346]&~m[347])|(~m[11]&m[344]&m[345]&~m[346]&~m[347])|(m[11]&~m[344]&~m[345]&m[346]&~m[347])|(~m[11]&m[344]&~m[345]&m[346]&~m[347])|(~m[11]&~m[344]&m[345]&m[346]&~m[347])|(m[11]&~m[344]&~m[345]&~m[346]&m[347])|(~m[11]&m[344]&~m[345]&~m[346]&m[347])|(~m[11]&~m[344]&m[345]&~m[346]&m[347])|(~m[11]&~m[344]&~m[345]&m[346]&m[347]))&BiasedRNG[302])|(((m[11]&m[344]&m[345]&~m[346]&~m[347])|(m[11]&m[344]&~m[345]&m[346]&~m[347])|(m[11]&~m[344]&m[345]&m[346]&~m[347])|(~m[11]&m[344]&m[345]&m[346]&~m[347])|(m[11]&m[344]&~m[345]&~m[346]&m[347])|(m[11]&~m[344]&m[345]&~m[346]&m[347])|(~m[11]&m[344]&m[345]&~m[346]&m[347])|(m[11]&~m[344]&~m[345]&m[346]&m[347])|(~m[11]&m[344]&~m[345]&m[346]&m[347])|(~m[11]&~m[344]&m[345]&m[346]&m[347]))&~BiasedRNG[302])|((m[11]&m[344]&m[345]&m[346]&~m[347])|(m[11]&m[344]&m[345]&~m[346]&m[347])|(m[11]&m[344]&~m[345]&m[346]&m[347])|(m[11]&~m[344]&m[345]&m[346]&m[347])|(~m[11]&m[344]&m[345]&m[346]&m[347])|(m[11]&m[344]&m[345]&m[346]&m[347]));
    m[79] = (((m[11]&m[348]&~m[349]&~m[350]&~m[351])|(m[11]&~m[348]&m[349]&~m[350]&~m[351])|(~m[11]&m[348]&m[349]&~m[350]&~m[351])|(m[11]&~m[348]&~m[349]&m[350]&~m[351])|(~m[11]&m[348]&~m[349]&m[350]&~m[351])|(~m[11]&~m[348]&m[349]&m[350]&~m[351])|(m[11]&~m[348]&~m[349]&~m[350]&m[351])|(~m[11]&m[348]&~m[349]&~m[350]&m[351])|(~m[11]&~m[348]&m[349]&~m[350]&m[351])|(~m[11]&~m[348]&~m[349]&m[350]&m[351]))&BiasedRNG[303])|(((m[11]&m[348]&m[349]&~m[350]&~m[351])|(m[11]&m[348]&~m[349]&m[350]&~m[351])|(m[11]&~m[348]&m[349]&m[350]&~m[351])|(~m[11]&m[348]&m[349]&m[350]&~m[351])|(m[11]&m[348]&~m[349]&~m[350]&m[351])|(m[11]&~m[348]&m[349]&~m[350]&m[351])|(~m[11]&m[348]&m[349]&~m[350]&m[351])|(m[11]&~m[348]&~m[349]&m[350]&m[351])|(~m[11]&m[348]&~m[349]&m[350]&m[351])|(~m[11]&~m[348]&m[349]&m[350]&m[351]))&~BiasedRNG[303])|((m[11]&m[348]&m[349]&m[350]&~m[351])|(m[11]&m[348]&m[349]&~m[350]&m[351])|(m[11]&m[348]&~m[349]&m[350]&m[351])|(m[11]&~m[348]&m[349]&m[350]&m[351])|(~m[11]&m[348]&m[349]&m[350]&m[351])|(m[11]&m[348]&m[349]&m[350]&m[351]));
    m[80] = (((m[12]&m[352]&~m[353]&~m[354]&~m[355])|(m[12]&~m[352]&m[353]&~m[354]&~m[355])|(~m[12]&m[352]&m[353]&~m[354]&~m[355])|(m[12]&~m[352]&~m[353]&m[354]&~m[355])|(~m[12]&m[352]&~m[353]&m[354]&~m[355])|(~m[12]&~m[352]&m[353]&m[354]&~m[355])|(m[12]&~m[352]&~m[353]&~m[354]&m[355])|(~m[12]&m[352]&~m[353]&~m[354]&m[355])|(~m[12]&~m[352]&m[353]&~m[354]&m[355])|(~m[12]&~m[352]&~m[353]&m[354]&m[355]))&BiasedRNG[304])|(((m[12]&m[352]&m[353]&~m[354]&~m[355])|(m[12]&m[352]&~m[353]&m[354]&~m[355])|(m[12]&~m[352]&m[353]&m[354]&~m[355])|(~m[12]&m[352]&m[353]&m[354]&~m[355])|(m[12]&m[352]&~m[353]&~m[354]&m[355])|(m[12]&~m[352]&m[353]&~m[354]&m[355])|(~m[12]&m[352]&m[353]&~m[354]&m[355])|(m[12]&~m[352]&~m[353]&m[354]&m[355])|(~m[12]&m[352]&~m[353]&m[354]&m[355])|(~m[12]&~m[352]&m[353]&m[354]&m[355]))&~BiasedRNG[304])|((m[12]&m[352]&m[353]&m[354]&~m[355])|(m[12]&m[352]&m[353]&~m[354]&m[355])|(m[12]&m[352]&~m[353]&m[354]&m[355])|(m[12]&~m[352]&m[353]&m[354]&m[355])|(~m[12]&m[352]&m[353]&m[354]&m[355])|(m[12]&m[352]&m[353]&m[354]&m[355]));
    m[81] = (((m[12]&m[356]&~m[357]&~m[358]&~m[359])|(m[12]&~m[356]&m[357]&~m[358]&~m[359])|(~m[12]&m[356]&m[357]&~m[358]&~m[359])|(m[12]&~m[356]&~m[357]&m[358]&~m[359])|(~m[12]&m[356]&~m[357]&m[358]&~m[359])|(~m[12]&~m[356]&m[357]&m[358]&~m[359])|(m[12]&~m[356]&~m[357]&~m[358]&m[359])|(~m[12]&m[356]&~m[357]&~m[358]&m[359])|(~m[12]&~m[356]&m[357]&~m[358]&m[359])|(~m[12]&~m[356]&~m[357]&m[358]&m[359]))&BiasedRNG[305])|(((m[12]&m[356]&m[357]&~m[358]&~m[359])|(m[12]&m[356]&~m[357]&m[358]&~m[359])|(m[12]&~m[356]&m[357]&m[358]&~m[359])|(~m[12]&m[356]&m[357]&m[358]&~m[359])|(m[12]&m[356]&~m[357]&~m[358]&m[359])|(m[12]&~m[356]&m[357]&~m[358]&m[359])|(~m[12]&m[356]&m[357]&~m[358]&m[359])|(m[12]&~m[356]&~m[357]&m[358]&m[359])|(~m[12]&m[356]&~m[357]&m[358]&m[359])|(~m[12]&~m[356]&m[357]&m[358]&m[359]))&~BiasedRNG[305])|((m[12]&m[356]&m[357]&m[358]&~m[359])|(m[12]&m[356]&m[357]&~m[358]&m[359])|(m[12]&m[356]&~m[357]&m[358]&m[359])|(m[12]&~m[356]&m[357]&m[358]&m[359])|(~m[12]&m[356]&m[357]&m[358]&m[359])|(m[12]&m[356]&m[357]&m[358]&m[359]));
    m[82] = (((m[12]&m[360]&~m[361]&~m[362]&~m[363])|(m[12]&~m[360]&m[361]&~m[362]&~m[363])|(~m[12]&m[360]&m[361]&~m[362]&~m[363])|(m[12]&~m[360]&~m[361]&m[362]&~m[363])|(~m[12]&m[360]&~m[361]&m[362]&~m[363])|(~m[12]&~m[360]&m[361]&m[362]&~m[363])|(m[12]&~m[360]&~m[361]&~m[362]&m[363])|(~m[12]&m[360]&~m[361]&~m[362]&m[363])|(~m[12]&~m[360]&m[361]&~m[362]&m[363])|(~m[12]&~m[360]&~m[361]&m[362]&m[363]))&BiasedRNG[306])|(((m[12]&m[360]&m[361]&~m[362]&~m[363])|(m[12]&m[360]&~m[361]&m[362]&~m[363])|(m[12]&~m[360]&m[361]&m[362]&~m[363])|(~m[12]&m[360]&m[361]&m[362]&~m[363])|(m[12]&m[360]&~m[361]&~m[362]&m[363])|(m[12]&~m[360]&m[361]&~m[362]&m[363])|(~m[12]&m[360]&m[361]&~m[362]&m[363])|(m[12]&~m[360]&~m[361]&m[362]&m[363])|(~m[12]&m[360]&~m[361]&m[362]&m[363])|(~m[12]&~m[360]&m[361]&m[362]&m[363]))&~BiasedRNG[306])|((m[12]&m[360]&m[361]&m[362]&~m[363])|(m[12]&m[360]&m[361]&~m[362]&m[363])|(m[12]&m[360]&~m[361]&m[362]&m[363])|(m[12]&~m[360]&m[361]&m[362]&m[363])|(~m[12]&m[360]&m[361]&m[362]&m[363])|(m[12]&m[360]&m[361]&m[362]&m[363]));
    m[83] = (((m[12]&m[364]&~m[365]&~m[366]&~m[367])|(m[12]&~m[364]&m[365]&~m[366]&~m[367])|(~m[12]&m[364]&m[365]&~m[366]&~m[367])|(m[12]&~m[364]&~m[365]&m[366]&~m[367])|(~m[12]&m[364]&~m[365]&m[366]&~m[367])|(~m[12]&~m[364]&m[365]&m[366]&~m[367])|(m[12]&~m[364]&~m[365]&~m[366]&m[367])|(~m[12]&m[364]&~m[365]&~m[366]&m[367])|(~m[12]&~m[364]&m[365]&~m[366]&m[367])|(~m[12]&~m[364]&~m[365]&m[366]&m[367]))&BiasedRNG[307])|(((m[12]&m[364]&m[365]&~m[366]&~m[367])|(m[12]&m[364]&~m[365]&m[366]&~m[367])|(m[12]&~m[364]&m[365]&m[366]&~m[367])|(~m[12]&m[364]&m[365]&m[366]&~m[367])|(m[12]&m[364]&~m[365]&~m[366]&m[367])|(m[12]&~m[364]&m[365]&~m[366]&m[367])|(~m[12]&m[364]&m[365]&~m[366]&m[367])|(m[12]&~m[364]&~m[365]&m[366]&m[367])|(~m[12]&m[364]&~m[365]&m[366]&m[367])|(~m[12]&~m[364]&m[365]&m[366]&m[367]))&~BiasedRNG[307])|((m[12]&m[364]&m[365]&m[366]&~m[367])|(m[12]&m[364]&m[365]&~m[366]&m[367])|(m[12]&m[364]&~m[365]&m[366]&m[367])|(m[12]&~m[364]&m[365]&m[366]&m[367])|(~m[12]&m[364]&m[365]&m[366]&m[367])|(m[12]&m[364]&m[365]&m[366]&m[367]));
    m[84] = (((m[13]&m[368]&~m[369]&~m[370]&~m[371])|(m[13]&~m[368]&m[369]&~m[370]&~m[371])|(~m[13]&m[368]&m[369]&~m[370]&~m[371])|(m[13]&~m[368]&~m[369]&m[370]&~m[371])|(~m[13]&m[368]&~m[369]&m[370]&~m[371])|(~m[13]&~m[368]&m[369]&m[370]&~m[371])|(m[13]&~m[368]&~m[369]&~m[370]&m[371])|(~m[13]&m[368]&~m[369]&~m[370]&m[371])|(~m[13]&~m[368]&m[369]&~m[370]&m[371])|(~m[13]&~m[368]&~m[369]&m[370]&m[371]))&BiasedRNG[308])|(((m[13]&m[368]&m[369]&~m[370]&~m[371])|(m[13]&m[368]&~m[369]&m[370]&~m[371])|(m[13]&~m[368]&m[369]&m[370]&~m[371])|(~m[13]&m[368]&m[369]&m[370]&~m[371])|(m[13]&m[368]&~m[369]&~m[370]&m[371])|(m[13]&~m[368]&m[369]&~m[370]&m[371])|(~m[13]&m[368]&m[369]&~m[370]&m[371])|(m[13]&~m[368]&~m[369]&m[370]&m[371])|(~m[13]&m[368]&~m[369]&m[370]&m[371])|(~m[13]&~m[368]&m[369]&m[370]&m[371]))&~BiasedRNG[308])|((m[13]&m[368]&m[369]&m[370]&~m[371])|(m[13]&m[368]&m[369]&~m[370]&m[371])|(m[13]&m[368]&~m[369]&m[370]&m[371])|(m[13]&~m[368]&m[369]&m[370]&m[371])|(~m[13]&m[368]&m[369]&m[370]&m[371])|(m[13]&m[368]&m[369]&m[370]&m[371]));
    m[85] = (((m[13]&m[372]&~m[373]&~m[374]&~m[375])|(m[13]&~m[372]&m[373]&~m[374]&~m[375])|(~m[13]&m[372]&m[373]&~m[374]&~m[375])|(m[13]&~m[372]&~m[373]&m[374]&~m[375])|(~m[13]&m[372]&~m[373]&m[374]&~m[375])|(~m[13]&~m[372]&m[373]&m[374]&~m[375])|(m[13]&~m[372]&~m[373]&~m[374]&m[375])|(~m[13]&m[372]&~m[373]&~m[374]&m[375])|(~m[13]&~m[372]&m[373]&~m[374]&m[375])|(~m[13]&~m[372]&~m[373]&m[374]&m[375]))&BiasedRNG[309])|(((m[13]&m[372]&m[373]&~m[374]&~m[375])|(m[13]&m[372]&~m[373]&m[374]&~m[375])|(m[13]&~m[372]&m[373]&m[374]&~m[375])|(~m[13]&m[372]&m[373]&m[374]&~m[375])|(m[13]&m[372]&~m[373]&~m[374]&m[375])|(m[13]&~m[372]&m[373]&~m[374]&m[375])|(~m[13]&m[372]&m[373]&~m[374]&m[375])|(m[13]&~m[372]&~m[373]&m[374]&m[375])|(~m[13]&m[372]&~m[373]&m[374]&m[375])|(~m[13]&~m[372]&m[373]&m[374]&m[375]))&~BiasedRNG[309])|((m[13]&m[372]&m[373]&m[374]&~m[375])|(m[13]&m[372]&m[373]&~m[374]&m[375])|(m[13]&m[372]&~m[373]&m[374]&m[375])|(m[13]&~m[372]&m[373]&m[374]&m[375])|(~m[13]&m[372]&m[373]&m[374]&m[375])|(m[13]&m[372]&m[373]&m[374]&m[375]));
    m[86] = (((m[13]&m[376]&~m[377]&~m[378]&~m[379])|(m[13]&~m[376]&m[377]&~m[378]&~m[379])|(~m[13]&m[376]&m[377]&~m[378]&~m[379])|(m[13]&~m[376]&~m[377]&m[378]&~m[379])|(~m[13]&m[376]&~m[377]&m[378]&~m[379])|(~m[13]&~m[376]&m[377]&m[378]&~m[379])|(m[13]&~m[376]&~m[377]&~m[378]&m[379])|(~m[13]&m[376]&~m[377]&~m[378]&m[379])|(~m[13]&~m[376]&m[377]&~m[378]&m[379])|(~m[13]&~m[376]&~m[377]&m[378]&m[379]))&BiasedRNG[310])|(((m[13]&m[376]&m[377]&~m[378]&~m[379])|(m[13]&m[376]&~m[377]&m[378]&~m[379])|(m[13]&~m[376]&m[377]&m[378]&~m[379])|(~m[13]&m[376]&m[377]&m[378]&~m[379])|(m[13]&m[376]&~m[377]&~m[378]&m[379])|(m[13]&~m[376]&m[377]&~m[378]&m[379])|(~m[13]&m[376]&m[377]&~m[378]&m[379])|(m[13]&~m[376]&~m[377]&m[378]&m[379])|(~m[13]&m[376]&~m[377]&m[378]&m[379])|(~m[13]&~m[376]&m[377]&m[378]&m[379]))&~BiasedRNG[310])|((m[13]&m[376]&m[377]&m[378]&~m[379])|(m[13]&m[376]&m[377]&~m[378]&m[379])|(m[13]&m[376]&~m[377]&m[378]&m[379])|(m[13]&~m[376]&m[377]&m[378]&m[379])|(~m[13]&m[376]&m[377]&m[378]&m[379])|(m[13]&m[376]&m[377]&m[378]&m[379]));
    m[87] = (((m[13]&m[380]&~m[381]&~m[382]&~m[383])|(m[13]&~m[380]&m[381]&~m[382]&~m[383])|(~m[13]&m[380]&m[381]&~m[382]&~m[383])|(m[13]&~m[380]&~m[381]&m[382]&~m[383])|(~m[13]&m[380]&~m[381]&m[382]&~m[383])|(~m[13]&~m[380]&m[381]&m[382]&~m[383])|(m[13]&~m[380]&~m[381]&~m[382]&m[383])|(~m[13]&m[380]&~m[381]&~m[382]&m[383])|(~m[13]&~m[380]&m[381]&~m[382]&m[383])|(~m[13]&~m[380]&~m[381]&m[382]&m[383]))&BiasedRNG[311])|(((m[13]&m[380]&m[381]&~m[382]&~m[383])|(m[13]&m[380]&~m[381]&m[382]&~m[383])|(m[13]&~m[380]&m[381]&m[382]&~m[383])|(~m[13]&m[380]&m[381]&m[382]&~m[383])|(m[13]&m[380]&~m[381]&~m[382]&m[383])|(m[13]&~m[380]&m[381]&~m[382]&m[383])|(~m[13]&m[380]&m[381]&~m[382]&m[383])|(m[13]&~m[380]&~m[381]&m[382]&m[383])|(~m[13]&m[380]&~m[381]&m[382]&m[383])|(~m[13]&~m[380]&m[381]&m[382]&m[383]))&~BiasedRNG[311])|((m[13]&m[380]&m[381]&m[382]&~m[383])|(m[13]&m[380]&m[381]&~m[382]&m[383])|(m[13]&m[380]&~m[381]&m[382]&m[383])|(m[13]&~m[380]&m[381]&m[382]&m[383])|(~m[13]&m[380]&m[381]&m[382]&m[383])|(m[13]&m[380]&m[381]&m[382]&m[383]));
    m[88] = (((m[14]&m[384]&~m[385]&~m[386]&~m[387])|(m[14]&~m[384]&m[385]&~m[386]&~m[387])|(~m[14]&m[384]&m[385]&~m[386]&~m[387])|(m[14]&~m[384]&~m[385]&m[386]&~m[387])|(~m[14]&m[384]&~m[385]&m[386]&~m[387])|(~m[14]&~m[384]&m[385]&m[386]&~m[387])|(m[14]&~m[384]&~m[385]&~m[386]&m[387])|(~m[14]&m[384]&~m[385]&~m[386]&m[387])|(~m[14]&~m[384]&m[385]&~m[386]&m[387])|(~m[14]&~m[384]&~m[385]&m[386]&m[387]))&BiasedRNG[312])|(((m[14]&m[384]&m[385]&~m[386]&~m[387])|(m[14]&m[384]&~m[385]&m[386]&~m[387])|(m[14]&~m[384]&m[385]&m[386]&~m[387])|(~m[14]&m[384]&m[385]&m[386]&~m[387])|(m[14]&m[384]&~m[385]&~m[386]&m[387])|(m[14]&~m[384]&m[385]&~m[386]&m[387])|(~m[14]&m[384]&m[385]&~m[386]&m[387])|(m[14]&~m[384]&~m[385]&m[386]&m[387])|(~m[14]&m[384]&~m[385]&m[386]&m[387])|(~m[14]&~m[384]&m[385]&m[386]&m[387]))&~BiasedRNG[312])|((m[14]&m[384]&m[385]&m[386]&~m[387])|(m[14]&m[384]&m[385]&~m[386]&m[387])|(m[14]&m[384]&~m[385]&m[386]&m[387])|(m[14]&~m[384]&m[385]&m[386]&m[387])|(~m[14]&m[384]&m[385]&m[386]&m[387])|(m[14]&m[384]&m[385]&m[386]&m[387]));
    m[89] = (((m[14]&m[388]&~m[389]&~m[390]&~m[391])|(m[14]&~m[388]&m[389]&~m[390]&~m[391])|(~m[14]&m[388]&m[389]&~m[390]&~m[391])|(m[14]&~m[388]&~m[389]&m[390]&~m[391])|(~m[14]&m[388]&~m[389]&m[390]&~m[391])|(~m[14]&~m[388]&m[389]&m[390]&~m[391])|(m[14]&~m[388]&~m[389]&~m[390]&m[391])|(~m[14]&m[388]&~m[389]&~m[390]&m[391])|(~m[14]&~m[388]&m[389]&~m[390]&m[391])|(~m[14]&~m[388]&~m[389]&m[390]&m[391]))&BiasedRNG[313])|(((m[14]&m[388]&m[389]&~m[390]&~m[391])|(m[14]&m[388]&~m[389]&m[390]&~m[391])|(m[14]&~m[388]&m[389]&m[390]&~m[391])|(~m[14]&m[388]&m[389]&m[390]&~m[391])|(m[14]&m[388]&~m[389]&~m[390]&m[391])|(m[14]&~m[388]&m[389]&~m[390]&m[391])|(~m[14]&m[388]&m[389]&~m[390]&m[391])|(m[14]&~m[388]&~m[389]&m[390]&m[391])|(~m[14]&m[388]&~m[389]&m[390]&m[391])|(~m[14]&~m[388]&m[389]&m[390]&m[391]))&~BiasedRNG[313])|((m[14]&m[388]&m[389]&m[390]&~m[391])|(m[14]&m[388]&m[389]&~m[390]&m[391])|(m[14]&m[388]&~m[389]&m[390]&m[391])|(m[14]&~m[388]&m[389]&m[390]&m[391])|(~m[14]&m[388]&m[389]&m[390]&m[391])|(m[14]&m[388]&m[389]&m[390]&m[391]));
    m[90] = (((m[14]&m[392]&~m[393]&~m[394]&~m[395])|(m[14]&~m[392]&m[393]&~m[394]&~m[395])|(~m[14]&m[392]&m[393]&~m[394]&~m[395])|(m[14]&~m[392]&~m[393]&m[394]&~m[395])|(~m[14]&m[392]&~m[393]&m[394]&~m[395])|(~m[14]&~m[392]&m[393]&m[394]&~m[395])|(m[14]&~m[392]&~m[393]&~m[394]&m[395])|(~m[14]&m[392]&~m[393]&~m[394]&m[395])|(~m[14]&~m[392]&m[393]&~m[394]&m[395])|(~m[14]&~m[392]&~m[393]&m[394]&m[395]))&BiasedRNG[314])|(((m[14]&m[392]&m[393]&~m[394]&~m[395])|(m[14]&m[392]&~m[393]&m[394]&~m[395])|(m[14]&~m[392]&m[393]&m[394]&~m[395])|(~m[14]&m[392]&m[393]&m[394]&~m[395])|(m[14]&m[392]&~m[393]&~m[394]&m[395])|(m[14]&~m[392]&m[393]&~m[394]&m[395])|(~m[14]&m[392]&m[393]&~m[394]&m[395])|(m[14]&~m[392]&~m[393]&m[394]&m[395])|(~m[14]&m[392]&~m[393]&m[394]&m[395])|(~m[14]&~m[392]&m[393]&m[394]&m[395]))&~BiasedRNG[314])|((m[14]&m[392]&m[393]&m[394]&~m[395])|(m[14]&m[392]&m[393]&~m[394]&m[395])|(m[14]&m[392]&~m[393]&m[394]&m[395])|(m[14]&~m[392]&m[393]&m[394]&m[395])|(~m[14]&m[392]&m[393]&m[394]&m[395])|(m[14]&m[392]&m[393]&m[394]&m[395]));
    m[91] = (((m[14]&m[396]&~m[397]&~m[398]&~m[399])|(m[14]&~m[396]&m[397]&~m[398]&~m[399])|(~m[14]&m[396]&m[397]&~m[398]&~m[399])|(m[14]&~m[396]&~m[397]&m[398]&~m[399])|(~m[14]&m[396]&~m[397]&m[398]&~m[399])|(~m[14]&~m[396]&m[397]&m[398]&~m[399])|(m[14]&~m[396]&~m[397]&~m[398]&m[399])|(~m[14]&m[396]&~m[397]&~m[398]&m[399])|(~m[14]&~m[396]&m[397]&~m[398]&m[399])|(~m[14]&~m[396]&~m[397]&m[398]&m[399]))&BiasedRNG[315])|(((m[14]&m[396]&m[397]&~m[398]&~m[399])|(m[14]&m[396]&~m[397]&m[398]&~m[399])|(m[14]&~m[396]&m[397]&m[398]&~m[399])|(~m[14]&m[396]&m[397]&m[398]&~m[399])|(m[14]&m[396]&~m[397]&~m[398]&m[399])|(m[14]&~m[396]&m[397]&~m[398]&m[399])|(~m[14]&m[396]&m[397]&~m[398]&m[399])|(m[14]&~m[396]&~m[397]&m[398]&m[399])|(~m[14]&m[396]&~m[397]&m[398]&m[399])|(~m[14]&~m[396]&m[397]&m[398]&m[399]))&~BiasedRNG[315])|((m[14]&m[396]&m[397]&m[398]&~m[399])|(m[14]&m[396]&m[397]&~m[398]&m[399])|(m[14]&m[396]&~m[397]&m[398]&m[399])|(m[14]&~m[396]&m[397]&m[398]&m[399])|(~m[14]&m[396]&m[397]&m[398]&m[399])|(m[14]&m[396]&m[397]&m[398]&m[399]));
    m[92] = (((m[15]&m[400]&~m[401]&~m[402]&~m[403])|(m[15]&~m[400]&m[401]&~m[402]&~m[403])|(~m[15]&m[400]&m[401]&~m[402]&~m[403])|(m[15]&~m[400]&~m[401]&m[402]&~m[403])|(~m[15]&m[400]&~m[401]&m[402]&~m[403])|(~m[15]&~m[400]&m[401]&m[402]&~m[403])|(m[15]&~m[400]&~m[401]&~m[402]&m[403])|(~m[15]&m[400]&~m[401]&~m[402]&m[403])|(~m[15]&~m[400]&m[401]&~m[402]&m[403])|(~m[15]&~m[400]&~m[401]&m[402]&m[403]))&BiasedRNG[316])|(((m[15]&m[400]&m[401]&~m[402]&~m[403])|(m[15]&m[400]&~m[401]&m[402]&~m[403])|(m[15]&~m[400]&m[401]&m[402]&~m[403])|(~m[15]&m[400]&m[401]&m[402]&~m[403])|(m[15]&m[400]&~m[401]&~m[402]&m[403])|(m[15]&~m[400]&m[401]&~m[402]&m[403])|(~m[15]&m[400]&m[401]&~m[402]&m[403])|(m[15]&~m[400]&~m[401]&m[402]&m[403])|(~m[15]&m[400]&~m[401]&m[402]&m[403])|(~m[15]&~m[400]&m[401]&m[402]&m[403]))&~BiasedRNG[316])|((m[15]&m[400]&m[401]&m[402]&~m[403])|(m[15]&m[400]&m[401]&~m[402]&m[403])|(m[15]&m[400]&~m[401]&m[402]&m[403])|(m[15]&~m[400]&m[401]&m[402]&m[403])|(~m[15]&m[400]&m[401]&m[402]&m[403])|(m[15]&m[400]&m[401]&m[402]&m[403]));
    m[93] = (((m[15]&m[404]&~m[405]&~m[406]&~m[407])|(m[15]&~m[404]&m[405]&~m[406]&~m[407])|(~m[15]&m[404]&m[405]&~m[406]&~m[407])|(m[15]&~m[404]&~m[405]&m[406]&~m[407])|(~m[15]&m[404]&~m[405]&m[406]&~m[407])|(~m[15]&~m[404]&m[405]&m[406]&~m[407])|(m[15]&~m[404]&~m[405]&~m[406]&m[407])|(~m[15]&m[404]&~m[405]&~m[406]&m[407])|(~m[15]&~m[404]&m[405]&~m[406]&m[407])|(~m[15]&~m[404]&~m[405]&m[406]&m[407]))&BiasedRNG[317])|(((m[15]&m[404]&m[405]&~m[406]&~m[407])|(m[15]&m[404]&~m[405]&m[406]&~m[407])|(m[15]&~m[404]&m[405]&m[406]&~m[407])|(~m[15]&m[404]&m[405]&m[406]&~m[407])|(m[15]&m[404]&~m[405]&~m[406]&m[407])|(m[15]&~m[404]&m[405]&~m[406]&m[407])|(~m[15]&m[404]&m[405]&~m[406]&m[407])|(m[15]&~m[404]&~m[405]&m[406]&m[407])|(~m[15]&m[404]&~m[405]&m[406]&m[407])|(~m[15]&~m[404]&m[405]&m[406]&m[407]))&~BiasedRNG[317])|((m[15]&m[404]&m[405]&m[406]&~m[407])|(m[15]&m[404]&m[405]&~m[406]&m[407])|(m[15]&m[404]&~m[405]&m[406]&m[407])|(m[15]&~m[404]&m[405]&m[406]&m[407])|(~m[15]&m[404]&m[405]&m[406]&m[407])|(m[15]&m[404]&m[405]&m[406]&m[407]));
    m[94] = (((m[15]&m[408]&~m[409]&~m[410]&~m[411])|(m[15]&~m[408]&m[409]&~m[410]&~m[411])|(~m[15]&m[408]&m[409]&~m[410]&~m[411])|(m[15]&~m[408]&~m[409]&m[410]&~m[411])|(~m[15]&m[408]&~m[409]&m[410]&~m[411])|(~m[15]&~m[408]&m[409]&m[410]&~m[411])|(m[15]&~m[408]&~m[409]&~m[410]&m[411])|(~m[15]&m[408]&~m[409]&~m[410]&m[411])|(~m[15]&~m[408]&m[409]&~m[410]&m[411])|(~m[15]&~m[408]&~m[409]&m[410]&m[411]))&BiasedRNG[318])|(((m[15]&m[408]&m[409]&~m[410]&~m[411])|(m[15]&m[408]&~m[409]&m[410]&~m[411])|(m[15]&~m[408]&m[409]&m[410]&~m[411])|(~m[15]&m[408]&m[409]&m[410]&~m[411])|(m[15]&m[408]&~m[409]&~m[410]&m[411])|(m[15]&~m[408]&m[409]&~m[410]&m[411])|(~m[15]&m[408]&m[409]&~m[410]&m[411])|(m[15]&~m[408]&~m[409]&m[410]&m[411])|(~m[15]&m[408]&~m[409]&m[410]&m[411])|(~m[15]&~m[408]&m[409]&m[410]&m[411]))&~BiasedRNG[318])|((m[15]&m[408]&m[409]&m[410]&~m[411])|(m[15]&m[408]&m[409]&~m[410]&m[411])|(m[15]&m[408]&~m[409]&m[410]&m[411])|(m[15]&~m[408]&m[409]&m[410]&m[411])|(~m[15]&m[408]&m[409]&m[410]&m[411])|(m[15]&m[408]&m[409]&m[410]&m[411]));
    m[95] = (((m[15]&m[412]&~m[413]&~m[414]&~m[415])|(m[15]&~m[412]&m[413]&~m[414]&~m[415])|(~m[15]&m[412]&m[413]&~m[414]&~m[415])|(m[15]&~m[412]&~m[413]&m[414]&~m[415])|(~m[15]&m[412]&~m[413]&m[414]&~m[415])|(~m[15]&~m[412]&m[413]&m[414]&~m[415])|(m[15]&~m[412]&~m[413]&~m[414]&m[415])|(~m[15]&m[412]&~m[413]&~m[414]&m[415])|(~m[15]&~m[412]&m[413]&~m[414]&m[415])|(~m[15]&~m[412]&~m[413]&m[414]&m[415]))&BiasedRNG[319])|(((m[15]&m[412]&m[413]&~m[414]&~m[415])|(m[15]&m[412]&~m[413]&m[414]&~m[415])|(m[15]&~m[412]&m[413]&m[414]&~m[415])|(~m[15]&m[412]&m[413]&m[414]&~m[415])|(m[15]&m[412]&~m[413]&~m[414]&m[415])|(m[15]&~m[412]&m[413]&~m[414]&m[415])|(~m[15]&m[412]&m[413]&~m[414]&m[415])|(m[15]&~m[412]&~m[413]&m[414]&m[415])|(~m[15]&m[412]&~m[413]&m[414]&m[415])|(~m[15]&~m[412]&m[413]&m[414]&m[415]))&~BiasedRNG[319])|((m[15]&m[412]&m[413]&m[414]&~m[415])|(m[15]&m[412]&m[413]&~m[414]&m[415])|(m[15]&m[412]&~m[413]&m[414]&m[415])|(m[15]&~m[412]&m[413]&m[414]&m[415])|(~m[15]&m[412]&m[413]&m[414]&m[415])|(m[15]&m[412]&m[413]&m[414]&m[415]));
    m[96] = (((m[16]&m[416]&~m[417]&~m[418]&~m[419])|(m[16]&~m[416]&m[417]&~m[418]&~m[419])|(~m[16]&m[416]&m[417]&~m[418]&~m[419])|(m[16]&~m[416]&~m[417]&m[418]&~m[419])|(~m[16]&m[416]&~m[417]&m[418]&~m[419])|(~m[16]&~m[416]&m[417]&m[418]&~m[419])|(m[16]&~m[416]&~m[417]&~m[418]&m[419])|(~m[16]&m[416]&~m[417]&~m[418]&m[419])|(~m[16]&~m[416]&m[417]&~m[418]&m[419])|(~m[16]&~m[416]&~m[417]&m[418]&m[419]))&BiasedRNG[320])|(((m[16]&m[416]&m[417]&~m[418]&~m[419])|(m[16]&m[416]&~m[417]&m[418]&~m[419])|(m[16]&~m[416]&m[417]&m[418]&~m[419])|(~m[16]&m[416]&m[417]&m[418]&~m[419])|(m[16]&m[416]&~m[417]&~m[418]&m[419])|(m[16]&~m[416]&m[417]&~m[418]&m[419])|(~m[16]&m[416]&m[417]&~m[418]&m[419])|(m[16]&~m[416]&~m[417]&m[418]&m[419])|(~m[16]&m[416]&~m[417]&m[418]&m[419])|(~m[16]&~m[416]&m[417]&m[418]&m[419]))&~BiasedRNG[320])|((m[16]&m[416]&m[417]&m[418]&~m[419])|(m[16]&m[416]&m[417]&~m[418]&m[419])|(m[16]&m[416]&~m[417]&m[418]&m[419])|(m[16]&~m[416]&m[417]&m[418]&m[419])|(~m[16]&m[416]&m[417]&m[418]&m[419])|(m[16]&m[416]&m[417]&m[418]&m[419]));
    m[97] = (((m[16]&m[420]&~m[421]&~m[422]&~m[423])|(m[16]&~m[420]&m[421]&~m[422]&~m[423])|(~m[16]&m[420]&m[421]&~m[422]&~m[423])|(m[16]&~m[420]&~m[421]&m[422]&~m[423])|(~m[16]&m[420]&~m[421]&m[422]&~m[423])|(~m[16]&~m[420]&m[421]&m[422]&~m[423])|(m[16]&~m[420]&~m[421]&~m[422]&m[423])|(~m[16]&m[420]&~m[421]&~m[422]&m[423])|(~m[16]&~m[420]&m[421]&~m[422]&m[423])|(~m[16]&~m[420]&~m[421]&m[422]&m[423]))&BiasedRNG[321])|(((m[16]&m[420]&m[421]&~m[422]&~m[423])|(m[16]&m[420]&~m[421]&m[422]&~m[423])|(m[16]&~m[420]&m[421]&m[422]&~m[423])|(~m[16]&m[420]&m[421]&m[422]&~m[423])|(m[16]&m[420]&~m[421]&~m[422]&m[423])|(m[16]&~m[420]&m[421]&~m[422]&m[423])|(~m[16]&m[420]&m[421]&~m[422]&m[423])|(m[16]&~m[420]&~m[421]&m[422]&m[423])|(~m[16]&m[420]&~m[421]&m[422]&m[423])|(~m[16]&~m[420]&m[421]&m[422]&m[423]))&~BiasedRNG[321])|((m[16]&m[420]&m[421]&m[422]&~m[423])|(m[16]&m[420]&m[421]&~m[422]&m[423])|(m[16]&m[420]&~m[421]&m[422]&m[423])|(m[16]&~m[420]&m[421]&m[422]&m[423])|(~m[16]&m[420]&m[421]&m[422]&m[423])|(m[16]&m[420]&m[421]&m[422]&m[423]));
    m[98] = (((m[16]&m[424]&~m[425]&~m[426]&~m[427])|(m[16]&~m[424]&m[425]&~m[426]&~m[427])|(~m[16]&m[424]&m[425]&~m[426]&~m[427])|(m[16]&~m[424]&~m[425]&m[426]&~m[427])|(~m[16]&m[424]&~m[425]&m[426]&~m[427])|(~m[16]&~m[424]&m[425]&m[426]&~m[427])|(m[16]&~m[424]&~m[425]&~m[426]&m[427])|(~m[16]&m[424]&~m[425]&~m[426]&m[427])|(~m[16]&~m[424]&m[425]&~m[426]&m[427])|(~m[16]&~m[424]&~m[425]&m[426]&m[427]))&BiasedRNG[322])|(((m[16]&m[424]&m[425]&~m[426]&~m[427])|(m[16]&m[424]&~m[425]&m[426]&~m[427])|(m[16]&~m[424]&m[425]&m[426]&~m[427])|(~m[16]&m[424]&m[425]&m[426]&~m[427])|(m[16]&m[424]&~m[425]&~m[426]&m[427])|(m[16]&~m[424]&m[425]&~m[426]&m[427])|(~m[16]&m[424]&m[425]&~m[426]&m[427])|(m[16]&~m[424]&~m[425]&m[426]&m[427])|(~m[16]&m[424]&~m[425]&m[426]&m[427])|(~m[16]&~m[424]&m[425]&m[426]&m[427]))&~BiasedRNG[322])|((m[16]&m[424]&m[425]&m[426]&~m[427])|(m[16]&m[424]&m[425]&~m[426]&m[427])|(m[16]&m[424]&~m[425]&m[426]&m[427])|(m[16]&~m[424]&m[425]&m[426]&m[427])|(~m[16]&m[424]&m[425]&m[426]&m[427])|(m[16]&m[424]&m[425]&m[426]&m[427]));
    m[99] = (((m[16]&m[428]&~m[429]&~m[430]&~m[431])|(m[16]&~m[428]&m[429]&~m[430]&~m[431])|(~m[16]&m[428]&m[429]&~m[430]&~m[431])|(m[16]&~m[428]&~m[429]&m[430]&~m[431])|(~m[16]&m[428]&~m[429]&m[430]&~m[431])|(~m[16]&~m[428]&m[429]&m[430]&~m[431])|(m[16]&~m[428]&~m[429]&~m[430]&m[431])|(~m[16]&m[428]&~m[429]&~m[430]&m[431])|(~m[16]&~m[428]&m[429]&~m[430]&m[431])|(~m[16]&~m[428]&~m[429]&m[430]&m[431]))&BiasedRNG[323])|(((m[16]&m[428]&m[429]&~m[430]&~m[431])|(m[16]&m[428]&~m[429]&m[430]&~m[431])|(m[16]&~m[428]&m[429]&m[430]&~m[431])|(~m[16]&m[428]&m[429]&m[430]&~m[431])|(m[16]&m[428]&~m[429]&~m[430]&m[431])|(m[16]&~m[428]&m[429]&~m[430]&m[431])|(~m[16]&m[428]&m[429]&~m[430]&m[431])|(m[16]&~m[428]&~m[429]&m[430]&m[431])|(~m[16]&m[428]&~m[429]&m[430]&m[431])|(~m[16]&~m[428]&m[429]&m[430]&m[431]))&~BiasedRNG[323])|((m[16]&m[428]&m[429]&m[430]&~m[431])|(m[16]&m[428]&m[429]&~m[430]&m[431])|(m[16]&m[428]&~m[429]&m[430]&m[431])|(m[16]&~m[428]&m[429]&m[430]&m[431])|(~m[16]&m[428]&m[429]&m[430]&m[431])|(m[16]&m[428]&m[429]&m[430]&m[431]));
    m[100] = (((m[17]&m[432]&~m[433]&~m[434]&~m[435])|(m[17]&~m[432]&m[433]&~m[434]&~m[435])|(~m[17]&m[432]&m[433]&~m[434]&~m[435])|(m[17]&~m[432]&~m[433]&m[434]&~m[435])|(~m[17]&m[432]&~m[433]&m[434]&~m[435])|(~m[17]&~m[432]&m[433]&m[434]&~m[435])|(m[17]&~m[432]&~m[433]&~m[434]&m[435])|(~m[17]&m[432]&~m[433]&~m[434]&m[435])|(~m[17]&~m[432]&m[433]&~m[434]&m[435])|(~m[17]&~m[432]&~m[433]&m[434]&m[435]))&BiasedRNG[324])|(((m[17]&m[432]&m[433]&~m[434]&~m[435])|(m[17]&m[432]&~m[433]&m[434]&~m[435])|(m[17]&~m[432]&m[433]&m[434]&~m[435])|(~m[17]&m[432]&m[433]&m[434]&~m[435])|(m[17]&m[432]&~m[433]&~m[434]&m[435])|(m[17]&~m[432]&m[433]&~m[434]&m[435])|(~m[17]&m[432]&m[433]&~m[434]&m[435])|(m[17]&~m[432]&~m[433]&m[434]&m[435])|(~m[17]&m[432]&~m[433]&m[434]&m[435])|(~m[17]&~m[432]&m[433]&m[434]&m[435]))&~BiasedRNG[324])|((m[17]&m[432]&m[433]&m[434]&~m[435])|(m[17]&m[432]&m[433]&~m[434]&m[435])|(m[17]&m[432]&~m[433]&m[434]&m[435])|(m[17]&~m[432]&m[433]&m[434]&m[435])|(~m[17]&m[432]&m[433]&m[434]&m[435])|(m[17]&m[432]&m[433]&m[434]&m[435]));
    m[101] = (((m[17]&m[436]&~m[437]&~m[438]&~m[439])|(m[17]&~m[436]&m[437]&~m[438]&~m[439])|(~m[17]&m[436]&m[437]&~m[438]&~m[439])|(m[17]&~m[436]&~m[437]&m[438]&~m[439])|(~m[17]&m[436]&~m[437]&m[438]&~m[439])|(~m[17]&~m[436]&m[437]&m[438]&~m[439])|(m[17]&~m[436]&~m[437]&~m[438]&m[439])|(~m[17]&m[436]&~m[437]&~m[438]&m[439])|(~m[17]&~m[436]&m[437]&~m[438]&m[439])|(~m[17]&~m[436]&~m[437]&m[438]&m[439]))&BiasedRNG[325])|(((m[17]&m[436]&m[437]&~m[438]&~m[439])|(m[17]&m[436]&~m[437]&m[438]&~m[439])|(m[17]&~m[436]&m[437]&m[438]&~m[439])|(~m[17]&m[436]&m[437]&m[438]&~m[439])|(m[17]&m[436]&~m[437]&~m[438]&m[439])|(m[17]&~m[436]&m[437]&~m[438]&m[439])|(~m[17]&m[436]&m[437]&~m[438]&m[439])|(m[17]&~m[436]&~m[437]&m[438]&m[439])|(~m[17]&m[436]&~m[437]&m[438]&m[439])|(~m[17]&~m[436]&m[437]&m[438]&m[439]))&~BiasedRNG[325])|((m[17]&m[436]&m[437]&m[438]&~m[439])|(m[17]&m[436]&m[437]&~m[438]&m[439])|(m[17]&m[436]&~m[437]&m[438]&m[439])|(m[17]&~m[436]&m[437]&m[438]&m[439])|(~m[17]&m[436]&m[437]&m[438]&m[439])|(m[17]&m[436]&m[437]&m[438]&m[439]));
    m[102] = (((m[17]&m[440]&~m[441]&~m[442]&~m[443])|(m[17]&~m[440]&m[441]&~m[442]&~m[443])|(~m[17]&m[440]&m[441]&~m[442]&~m[443])|(m[17]&~m[440]&~m[441]&m[442]&~m[443])|(~m[17]&m[440]&~m[441]&m[442]&~m[443])|(~m[17]&~m[440]&m[441]&m[442]&~m[443])|(m[17]&~m[440]&~m[441]&~m[442]&m[443])|(~m[17]&m[440]&~m[441]&~m[442]&m[443])|(~m[17]&~m[440]&m[441]&~m[442]&m[443])|(~m[17]&~m[440]&~m[441]&m[442]&m[443]))&BiasedRNG[326])|(((m[17]&m[440]&m[441]&~m[442]&~m[443])|(m[17]&m[440]&~m[441]&m[442]&~m[443])|(m[17]&~m[440]&m[441]&m[442]&~m[443])|(~m[17]&m[440]&m[441]&m[442]&~m[443])|(m[17]&m[440]&~m[441]&~m[442]&m[443])|(m[17]&~m[440]&m[441]&~m[442]&m[443])|(~m[17]&m[440]&m[441]&~m[442]&m[443])|(m[17]&~m[440]&~m[441]&m[442]&m[443])|(~m[17]&m[440]&~m[441]&m[442]&m[443])|(~m[17]&~m[440]&m[441]&m[442]&m[443]))&~BiasedRNG[326])|((m[17]&m[440]&m[441]&m[442]&~m[443])|(m[17]&m[440]&m[441]&~m[442]&m[443])|(m[17]&m[440]&~m[441]&m[442]&m[443])|(m[17]&~m[440]&m[441]&m[442]&m[443])|(~m[17]&m[440]&m[441]&m[442]&m[443])|(m[17]&m[440]&m[441]&m[442]&m[443]));
    m[103] = (((m[17]&m[444]&~m[445]&~m[446]&~m[447])|(m[17]&~m[444]&m[445]&~m[446]&~m[447])|(~m[17]&m[444]&m[445]&~m[446]&~m[447])|(m[17]&~m[444]&~m[445]&m[446]&~m[447])|(~m[17]&m[444]&~m[445]&m[446]&~m[447])|(~m[17]&~m[444]&m[445]&m[446]&~m[447])|(m[17]&~m[444]&~m[445]&~m[446]&m[447])|(~m[17]&m[444]&~m[445]&~m[446]&m[447])|(~m[17]&~m[444]&m[445]&~m[446]&m[447])|(~m[17]&~m[444]&~m[445]&m[446]&m[447]))&BiasedRNG[327])|(((m[17]&m[444]&m[445]&~m[446]&~m[447])|(m[17]&m[444]&~m[445]&m[446]&~m[447])|(m[17]&~m[444]&m[445]&m[446]&~m[447])|(~m[17]&m[444]&m[445]&m[446]&~m[447])|(m[17]&m[444]&~m[445]&~m[446]&m[447])|(m[17]&~m[444]&m[445]&~m[446]&m[447])|(~m[17]&m[444]&m[445]&~m[446]&m[447])|(m[17]&~m[444]&~m[445]&m[446]&m[447])|(~m[17]&m[444]&~m[445]&m[446]&m[447])|(~m[17]&~m[444]&m[445]&m[446]&m[447]))&~BiasedRNG[327])|((m[17]&m[444]&m[445]&m[446]&~m[447])|(m[17]&m[444]&m[445]&~m[446]&m[447])|(m[17]&m[444]&~m[445]&m[446]&m[447])|(m[17]&~m[444]&m[445]&m[446]&m[447])|(~m[17]&m[444]&m[445]&m[446]&m[447])|(m[17]&m[444]&m[445]&m[446]&m[447]));
    m[104] = (((m[18]&m[448]&~m[449]&~m[450]&~m[451])|(m[18]&~m[448]&m[449]&~m[450]&~m[451])|(~m[18]&m[448]&m[449]&~m[450]&~m[451])|(m[18]&~m[448]&~m[449]&m[450]&~m[451])|(~m[18]&m[448]&~m[449]&m[450]&~m[451])|(~m[18]&~m[448]&m[449]&m[450]&~m[451])|(m[18]&~m[448]&~m[449]&~m[450]&m[451])|(~m[18]&m[448]&~m[449]&~m[450]&m[451])|(~m[18]&~m[448]&m[449]&~m[450]&m[451])|(~m[18]&~m[448]&~m[449]&m[450]&m[451]))&BiasedRNG[328])|(((m[18]&m[448]&m[449]&~m[450]&~m[451])|(m[18]&m[448]&~m[449]&m[450]&~m[451])|(m[18]&~m[448]&m[449]&m[450]&~m[451])|(~m[18]&m[448]&m[449]&m[450]&~m[451])|(m[18]&m[448]&~m[449]&~m[450]&m[451])|(m[18]&~m[448]&m[449]&~m[450]&m[451])|(~m[18]&m[448]&m[449]&~m[450]&m[451])|(m[18]&~m[448]&~m[449]&m[450]&m[451])|(~m[18]&m[448]&~m[449]&m[450]&m[451])|(~m[18]&~m[448]&m[449]&m[450]&m[451]))&~BiasedRNG[328])|((m[18]&m[448]&m[449]&m[450]&~m[451])|(m[18]&m[448]&m[449]&~m[450]&m[451])|(m[18]&m[448]&~m[449]&m[450]&m[451])|(m[18]&~m[448]&m[449]&m[450]&m[451])|(~m[18]&m[448]&m[449]&m[450]&m[451])|(m[18]&m[448]&m[449]&m[450]&m[451]));
    m[105] = (((m[18]&m[452]&~m[453]&~m[454]&~m[455])|(m[18]&~m[452]&m[453]&~m[454]&~m[455])|(~m[18]&m[452]&m[453]&~m[454]&~m[455])|(m[18]&~m[452]&~m[453]&m[454]&~m[455])|(~m[18]&m[452]&~m[453]&m[454]&~m[455])|(~m[18]&~m[452]&m[453]&m[454]&~m[455])|(m[18]&~m[452]&~m[453]&~m[454]&m[455])|(~m[18]&m[452]&~m[453]&~m[454]&m[455])|(~m[18]&~m[452]&m[453]&~m[454]&m[455])|(~m[18]&~m[452]&~m[453]&m[454]&m[455]))&BiasedRNG[329])|(((m[18]&m[452]&m[453]&~m[454]&~m[455])|(m[18]&m[452]&~m[453]&m[454]&~m[455])|(m[18]&~m[452]&m[453]&m[454]&~m[455])|(~m[18]&m[452]&m[453]&m[454]&~m[455])|(m[18]&m[452]&~m[453]&~m[454]&m[455])|(m[18]&~m[452]&m[453]&~m[454]&m[455])|(~m[18]&m[452]&m[453]&~m[454]&m[455])|(m[18]&~m[452]&~m[453]&m[454]&m[455])|(~m[18]&m[452]&~m[453]&m[454]&m[455])|(~m[18]&~m[452]&m[453]&m[454]&m[455]))&~BiasedRNG[329])|((m[18]&m[452]&m[453]&m[454]&~m[455])|(m[18]&m[452]&m[453]&~m[454]&m[455])|(m[18]&m[452]&~m[453]&m[454]&m[455])|(m[18]&~m[452]&m[453]&m[454]&m[455])|(~m[18]&m[452]&m[453]&m[454]&m[455])|(m[18]&m[452]&m[453]&m[454]&m[455]));
    m[106] = (((m[18]&m[456]&~m[457]&~m[458]&~m[459])|(m[18]&~m[456]&m[457]&~m[458]&~m[459])|(~m[18]&m[456]&m[457]&~m[458]&~m[459])|(m[18]&~m[456]&~m[457]&m[458]&~m[459])|(~m[18]&m[456]&~m[457]&m[458]&~m[459])|(~m[18]&~m[456]&m[457]&m[458]&~m[459])|(m[18]&~m[456]&~m[457]&~m[458]&m[459])|(~m[18]&m[456]&~m[457]&~m[458]&m[459])|(~m[18]&~m[456]&m[457]&~m[458]&m[459])|(~m[18]&~m[456]&~m[457]&m[458]&m[459]))&BiasedRNG[330])|(((m[18]&m[456]&m[457]&~m[458]&~m[459])|(m[18]&m[456]&~m[457]&m[458]&~m[459])|(m[18]&~m[456]&m[457]&m[458]&~m[459])|(~m[18]&m[456]&m[457]&m[458]&~m[459])|(m[18]&m[456]&~m[457]&~m[458]&m[459])|(m[18]&~m[456]&m[457]&~m[458]&m[459])|(~m[18]&m[456]&m[457]&~m[458]&m[459])|(m[18]&~m[456]&~m[457]&m[458]&m[459])|(~m[18]&m[456]&~m[457]&m[458]&m[459])|(~m[18]&~m[456]&m[457]&m[458]&m[459]))&~BiasedRNG[330])|((m[18]&m[456]&m[457]&m[458]&~m[459])|(m[18]&m[456]&m[457]&~m[458]&m[459])|(m[18]&m[456]&~m[457]&m[458]&m[459])|(m[18]&~m[456]&m[457]&m[458]&m[459])|(~m[18]&m[456]&m[457]&m[458]&m[459])|(m[18]&m[456]&m[457]&m[458]&m[459]));
    m[107] = (((m[18]&m[460]&~m[461]&~m[462]&~m[463])|(m[18]&~m[460]&m[461]&~m[462]&~m[463])|(~m[18]&m[460]&m[461]&~m[462]&~m[463])|(m[18]&~m[460]&~m[461]&m[462]&~m[463])|(~m[18]&m[460]&~m[461]&m[462]&~m[463])|(~m[18]&~m[460]&m[461]&m[462]&~m[463])|(m[18]&~m[460]&~m[461]&~m[462]&m[463])|(~m[18]&m[460]&~m[461]&~m[462]&m[463])|(~m[18]&~m[460]&m[461]&~m[462]&m[463])|(~m[18]&~m[460]&~m[461]&m[462]&m[463]))&BiasedRNG[331])|(((m[18]&m[460]&m[461]&~m[462]&~m[463])|(m[18]&m[460]&~m[461]&m[462]&~m[463])|(m[18]&~m[460]&m[461]&m[462]&~m[463])|(~m[18]&m[460]&m[461]&m[462]&~m[463])|(m[18]&m[460]&~m[461]&~m[462]&m[463])|(m[18]&~m[460]&m[461]&~m[462]&m[463])|(~m[18]&m[460]&m[461]&~m[462]&m[463])|(m[18]&~m[460]&~m[461]&m[462]&m[463])|(~m[18]&m[460]&~m[461]&m[462]&m[463])|(~m[18]&~m[460]&m[461]&m[462]&m[463]))&~BiasedRNG[331])|((m[18]&m[460]&m[461]&m[462]&~m[463])|(m[18]&m[460]&m[461]&~m[462]&m[463])|(m[18]&m[460]&~m[461]&m[462]&m[463])|(m[18]&~m[460]&m[461]&m[462]&m[463])|(~m[18]&m[460]&m[461]&m[462]&m[463])|(m[18]&m[460]&m[461]&m[462]&m[463]));
    m[108] = (((m[19]&m[464]&~m[465]&~m[466]&~m[467])|(m[19]&~m[464]&m[465]&~m[466]&~m[467])|(~m[19]&m[464]&m[465]&~m[466]&~m[467])|(m[19]&~m[464]&~m[465]&m[466]&~m[467])|(~m[19]&m[464]&~m[465]&m[466]&~m[467])|(~m[19]&~m[464]&m[465]&m[466]&~m[467])|(m[19]&~m[464]&~m[465]&~m[466]&m[467])|(~m[19]&m[464]&~m[465]&~m[466]&m[467])|(~m[19]&~m[464]&m[465]&~m[466]&m[467])|(~m[19]&~m[464]&~m[465]&m[466]&m[467]))&BiasedRNG[332])|(((m[19]&m[464]&m[465]&~m[466]&~m[467])|(m[19]&m[464]&~m[465]&m[466]&~m[467])|(m[19]&~m[464]&m[465]&m[466]&~m[467])|(~m[19]&m[464]&m[465]&m[466]&~m[467])|(m[19]&m[464]&~m[465]&~m[466]&m[467])|(m[19]&~m[464]&m[465]&~m[466]&m[467])|(~m[19]&m[464]&m[465]&~m[466]&m[467])|(m[19]&~m[464]&~m[465]&m[466]&m[467])|(~m[19]&m[464]&~m[465]&m[466]&m[467])|(~m[19]&~m[464]&m[465]&m[466]&m[467]))&~BiasedRNG[332])|((m[19]&m[464]&m[465]&m[466]&~m[467])|(m[19]&m[464]&m[465]&~m[466]&m[467])|(m[19]&m[464]&~m[465]&m[466]&m[467])|(m[19]&~m[464]&m[465]&m[466]&m[467])|(~m[19]&m[464]&m[465]&m[466]&m[467])|(m[19]&m[464]&m[465]&m[466]&m[467]));
    m[109] = (((m[19]&m[468]&~m[469]&~m[470]&~m[471])|(m[19]&~m[468]&m[469]&~m[470]&~m[471])|(~m[19]&m[468]&m[469]&~m[470]&~m[471])|(m[19]&~m[468]&~m[469]&m[470]&~m[471])|(~m[19]&m[468]&~m[469]&m[470]&~m[471])|(~m[19]&~m[468]&m[469]&m[470]&~m[471])|(m[19]&~m[468]&~m[469]&~m[470]&m[471])|(~m[19]&m[468]&~m[469]&~m[470]&m[471])|(~m[19]&~m[468]&m[469]&~m[470]&m[471])|(~m[19]&~m[468]&~m[469]&m[470]&m[471]))&BiasedRNG[333])|(((m[19]&m[468]&m[469]&~m[470]&~m[471])|(m[19]&m[468]&~m[469]&m[470]&~m[471])|(m[19]&~m[468]&m[469]&m[470]&~m[471])|(~m[19]&m[468]&m[469]&m[470]&~m[471])|(m[19]&m[468]&~m[469]&~m[470]&m[471])|(m[19]&~m[468]&m[469]&~m[470]&m[471])|(~m[19]&m[468]&m[469]&~m[470]&m[471])|(m[19]&~m[468]&~m[469]&m[470]&m[471])|(~m[19]&m[468]&~m[469]&m[470]&m[471])|(~m[19]&~m[468]&m[469]&m[470]&m[471]))&~BiasedRNG[333])|((m[19]&m[468]&m[469]&m[470]&~m[471])|(m[19]&m[468]&m[469]&~m[470]&m[471])|(m[19]&m[468]&~m[469]&m[470]&m[471])|(m[19]&~m[468]&m[469]&m[470]&m[471])|(~m[19]&m[468]&m[469]&m[470]&m[471])|(m[19]&m[468]&m[469]&m[470]&m[471]));
    m[110] = (((m[19]&m[472]&~m[473]&~m[474]&~m[475])|(m[19]&~m[472]&m[473]&~m[474]&~m[475])|(~m[19]&m[472]&m[473]&~m[474]&~m[475])|(m[19]&~m[472]&~m[473]&m[474]&~m[475])|(~m[19]&m[472]&~m[473]&m[474]&~m[475])|(~m[19]&~m[472]&m[473]&m[474]&~m[475])|(m[19]&~m[472]&~m[473]&~m[474]&m[475])|(~m[19]&m[472]&~m[473]&~m[474]&m[475])|(~m[19]&~m[472]&m[473]&~m[474]&m[475])|(~m[19]&~m[472]&~m[473]&m[474]&m[475]))&BiasedRNG[334])|(((m[19]&m[472]&m[473]&~m[474]&~m[475])|(m[19]&m[472]&~m[473]&m[474]&~m[475])|(m[19]&~m[472]&m[473]&m[474]&~m[475])|(~m[19]&m[472]&m[473]&m[474]&~m[475])|(m[19]&m[472]&~m[473]&~m[474]&m[475])|(m[19]&~m[472]&m[473]&~m[474]&m[475])|(~m[19]&m[472]&m[473]&~m[474]&m[475])|(m[19]&~m[472]&~m[473]&m[474]&m[475])|(~m[19]&m[472]&~m[473]&m[474]&m[475])|(~m[19]&~m[472]&m[473]&m[474]&m[475]))&~BiasedRNG[334])|((m[19]&m[472]&m[473]&m[474]&~m[475])|(m[19]&m[472]&m[473]&~m[474]&m[475])|(m[19]&m[472]&~m[473]&m[474]&m[475])|(m[19]&~m[472]&m[473]&m[474]&m[475])|(~m[19]&m[472]&m[473]&m[474]&m[475])|(m[19]&m[472]&m[473]&m[474]&m[475]));
    m[111] = (((m[19]&m[476]&~m[477]&~m[478]&~m[479])|(m[19]&~m[476]&m[477]&~m[478]&~m[479])|(~m[19]&m[476]&m[477]&~m[478]&~m[479])|(m[19]&~m[476]&~m[477]&m[478]&~m[479])|(~m[19]&m[476]&~m[477]&m[478]&~m[479])|(~m[19]&~m[476]&m[477]&m[478]&~m[479])|(m[19]&~m[476]&~m[477]&~m[478]&m[479])|(~m[19]&m[476]&~m[477]&~m[478]&m[479])|(~m[19]&~m[476]&m[477]&~m[478]&m[479])|(~m[19]&~m[476]&~m[477]&m[478]&m[479]))&BiasedRNG[335])|(((m[19]&m[476]&m[477]&~m[478]&~m[479])|(m[19]&m[476]&~m[477]&m[478]&~m[479])|(m[19]&~m[476]&m[477]&m[478]&~m[479])|(~m[19]&m[476]&m[477]&m[478]&~m[479])|(m[19]&m[476]&~m[477]&~m[478]&m[479])|(m[19]&~m[476]&m[477]&~m[478]&m[479])|(~m[19]&m[476]&m[477]&~m[478]&m[479])|(m[19]&~m[476]&~m[477]&m[478]&m[479])|(~m[19]&m[476]&~m[477]&m[478]&m[479])|(~m[19]&~m[476]&m[477]&m[478]&m[479]))&~BiasedRNG[335])|((m[19]&m[476]&m[477]&m[478]&~m[479])|(m[19]&m[476]&m[477]&~m[478]&m[479])|(m[19]&m[476]&~m[477]&m[478]&m[479])|(m[19]&~m[476]&m[477]&m[478]&m[479])|(~m[19]&m[476]&m[477]&m[478]&m[479])|(m[19]&m[476]&m[477]&m[478]&m[479]));
    m[112] = (((m[20]&m[480]&~m[481]&~m[482]&~m[483])|(m[20]&~m[480]&m[481]&~m[482]&~m[483])|(~m[20]&m[480]&m[481]&~m[482]&~m[483])|(m[20]&~m[480]&~m[481]&m[482]&~m[483])|(~m[20]&m[480]&~m[481]&m[482]&~m[483])|(~m[20]&~m[480]&m[481]&m[482]&~m[483])|(m[20]&~m[480]&~m[481]&~m[482]&m[483])|(~m[20]&m[480]&~m[481]&~m[482]&m[483])|(~m[20]&~m[480]&m[481]&~m[482]&m[483])|(~m[20]&~m[480]&~m[481]&m[482]&m[483]))&BiasedRNG[336])|(((m[20]&m[480]&m[481]&~m[482]&~m[483])|(m[20]&m[480]&~m[481]&m[482]&~m[483])|(m[20]&~m[480]&m[481]&m[482]&~m[483])|(~m[20]&m[480]&m[481]&m[482]&~m[483])|(m[20]&m[480]&~m[481]&~m[482]&m[483])|(m[20]&~m[480]&m[481]&~m[482]&m[483])|(~m[20]&m[480]&m[481]&~m[482]&m[483])|(m[20]&~m[480]&~m[481]&m[482]&m[483])|(~m[20]&m[480]&~m[481]&m[482]&m[483])|(~m[20]&~m[480]&m[481]&m[482]&m[483]))&~BiasedRNG[336])|((m[20]&m[480]&m[481]&m[482]&~m[483])|(m[20]&m[480]&m[481]&~m[482]&m[483])|(m[20]&m[480]&~m[481]&m[482]&m[483])|(m[20]&~m[480]&m[481]&m[482]&m[483])|(~m[20]&m[480]&m[481]&m[482]&m[483])|(m[20]&m[480]&m[481]&m[482]&m[483]));
    m[113] = (((m[20]&m[484]&~m[485]&~m[486]&~m[487])|(m[20]&~m[484]&m[485]&~m[486]&~m[487])|(~m[20]&m[484]&m[485]&~m[486]&~m[487])|(m[20]&~m[484]&~m[485]&m[486]&~m[487])|(~m[20]&m[484]&~m[485]&m[486]&~m[487])|(~m[20]&~m[484]&m[485]&m[486]&~m[487])|(m[20]&~m[484]&~m[485]&~m[486]&m[487])|(~m[20]&m[484]&~m[485]&~m[486]&m[487])|(~m[20]&~m[484]&m[485]&~m[486]&m[487])|(~m[20]&~m[484]&~m[485]&m[486]&m[487]))&BiasedRNG[337])|(((m[20]&m[484]&m[485]&~m[486]&~m[487])|(m[20]&m[484]&~m[485]&m[486]&~m[487])|(m[20]&~m[484]&m[485]&m[486]&~m[487])|(~m[20]&m[484]&m[485]&m[486]&~m[487])|(m[20]&m[484]&~m[485]&~m[486]&m[487])|(m[20]&~m[484]&m[485]&~m[486]&m[487])|(~m[20]&m[484]&m[485]&~m[486]&m[487])|(m[20]&~m[484]&~m[485]&m[486]&m[487])|(~m[20]&m[484]&~m[485]&m[486]&m[487])|(~m[20]&~m[484]&m[485]&m[486]&m[487]))&~BiasedRNG[337])|((m[20]&m[484]&m[485]&m[486]&~m[487])|(m[20]&m[484]&m[485]&~m[486]&m[487])|(m[20]&m[484]&~m[485]&m[486]&m[487])|(m[20]&~m[484]&m[485]&m[486]&m[487])|(~m[20]&m[484]&m[485]&m[486]&m[487])|(m[20]&m[484]&m[485]&m[486]&m[487]));
    m[114] = (((m[20]&m[488]&~m[489]&~m[490]&~m[491])|(m[20]&~m[488]&m[489]&~m[490]&~m[491])|(~m[20]&m[488]&m[489]&~m[490]&~m[491])|(m[20]&~m[488]&~m[489]&m[490]&~m[491])|(~m[20]&m[488]&~m[489]&m[490]&~m[491])|(~m[20]&~m[488]&m[489]&m[490]&~m[491])|(m[20]&~m[488]&~m[489]&~m[490]&m[491])|(~m[20]&m[488]&~m[489]&~m[490]&m[491])|(~m[20]&~m[488]&m[489]&~m[490]&m[491])|(~m[20]&~m[488]&~m[489]&m[490]&m[491]))&BiasedRNG[338])|(((m[20]&m[488]&m[489]&~m[490]&~m[491])|(m[20]&m[488]&~m[489]&m[490]&~m[491])|(m[20]&~m[488]&m[489]&m[490]&~m[491])|(~m[20]&m[488]&m[489]&m[490]&~m[491])|(m[20]&m[488]&~m[489]&~m[490]&m[491])|(m[20]&~m[488]&m[489]&~m[490]&m[491])|(~m[20]&m[488]&m[489]&~m[490]&m[491])|(m[20]&~m[488]&~m[489]&m[490]&m[491])|(~m[20]&m[488]&~m[489]&m[490]&m[491])|(~m[20]&~m[488]&m[489]&m[490]&m[491]))&~BiasedRNG[338])|((m[20]&m[488]&m[489]&m[490]&~m[491])|(m[20]&m[488]&m[489]&~m[490]&m[491])|(m[20]&m[488]&~m[489]&m[490]&m[491])|(m[20]&~m[488]&m[489]&m[490]&m[491])|(~m[20]&m[488]&m[489]&m[490]&m[491])|(m[20]&m[488]&m[489]&m[490]&m[491]));
    m[115] = (((m[20]&m[492]&~m[493]&~m[494]&~m[495])|(m[20]&~m[492]&m[493]&~m[494]&~m[495])|(~m[20]&m[492]&m[493]&~m[494]&~m[495])|(m[20]&~m[492]&~m[493]&m[494]&~m[495])|(~m[20]&m[492]&~m[493]&m[494]&~m[495])|(~m[20]&~m[492]&m[493]&m[494]&~m[495])|(m[20]&~m[492]&~m[493]&~m[494]&m[495])|(~m[20]&m[492]&~m[493]&~m[494]&m[495])|(~m[20]&~m[492]&m[493]&~m[494]&m[495])|(~m[20]&~m[492]&~m[493]&m[494]&m[495]))&BiasedRNG[339])|(((m[20]&m[492]&m[493]&~m[494]&~m[495])|(m[20]&m[492]&~m[493]&m[494]&~m[495])|(m[20]&~m[492]&m[493]&m[494]&~m[495])|(~m[20]&m[492]&m[493]&m[494]&~m[495])|(m[20]&m[492]&~m[493]&~m[494]&m[495])|(m[20]&~m[492]&m[493]&~m[494]&m[495])|(~m[20]&m[492]&m[493]&~m[494]&m[495])|(m[20]&~m[492]&~m[493]&m[494]&m[495])|(~m[20]&m[492]&~m[493]&m[494]&m[495])|(~m[20]&~m[492]&m[493]&m[494]&m[495]))&~BiasedRNG[339])|((m[20]&m[492]&m[493]&m[494]&~m[495])|(m[20]&m[492]&m[493]&~m[494]&m[495])|(m[20]&m[492]&~m[493]&m[494]&m[495])|(m[20]&~m[492]&m[493]&m[494]&m[495])|(~m[20]&m[492]&m[493]&m[494]&m[495])|(m[20]&m[492]&m[493]&m[494]&m[495]));
    m[116] = (((m[21]&m[496]&~m[497]&~m[498]&~m[499])|(m[21]&~m[496]&m[497]&~m[498]&~m[499])|(~m[21]&m[496]&m[497]&~m[498]&~m[499])|(m[21]&~m[496]&~m[497]&m[498]&~m[499])|(~m[21]&m[496]&~m[497]&m[498]&~m[499])|(~m[21]&~m[496]&m[497]&m[498]&~m[499])|(m[21]&~m[496]&~m[497]&~m[498]&m[499])|(~m[21]&m[496]&~m[497]&~m[498]&m[499])|(~m[21]&~m[496]&m[497]&~m[498]&m[499])|(~m[21]&~m[496]&~m[497]&m[498]&m[499]))&BiasedRNG[340])|(((m[21]&m[496]&m[497]&~m[498]&~m[499])|(m[21]&m[496]&~m[497]&m[498]&~m[499])|(m[21]&~m[496]&m[497]&m[498]&~m[499])|(~m[21]&m[496]&m[497]&m[498]&~m[499])|(m[21]&m[496]&~m[497]&~m[498]&m[499])|(m[21]&~m[496]&m[497]&~m[498]&m[499])|(~m[21]&m[496]&m[497]&~m[498]&m[499])|(m[21]&~m[496]&~m[497]&m[498]&m[499])|(~m[21]&m[496]&~m[497]&m[498]&m[499])|(~m[21]&~m[496]&m[497]&m[498]&m[499]))&~BiasedRNG[340])|((m[21]&m[496]&m[497]&m[498]&~m[499])|(m[21]&m[496]&m[497]&~m[498]&m[499])|(m[21]&m[496]&~m[497]&m[498]&m[499])|(m[21]&~m[496]&m[497]&m[498]&m[499])|(~m[21]&m[496]&m[497]&m[498]&m[499])|(m[21]&m[496]&m[497]&m[498]&m[499]));
    m[117] = (((m[21]&m[500]&~m[501]&~m[502]&~m[503])|(m[21]&~m[500]&m[501]&~m[502]&~m[503])|(~m[21]&m[500]&m[501]&~m[502]&~m[503])|(m[21]&~m[500]&~m[501]&m[502]&~m[503])|(~m[21]&m[500]&~m[501]&m[502]&~m[503])|(~m[21]&~m[500]&m[501]&m[502]&~m[503])|(m[21]&~m[500]&~m[501]&~m[502]&m[503])|(~m[21]&m[500]&~m[501]&~m[502]&m[503])|(~m[21]&~m[500]&m[501]&~m[502]&m[503])|(~m[21]&~m[500]&~m[501]&m[502]&m[503]))&BiasedRNG[341])|(((m[21]&m[500]&m[501]&~m[502]&~m[503])|(m[21]&m[500]&~m[501]&m[502]&~m[503])|(m[21]&~m[500]&m[501]&m[502]&~m[503])|(~m[21]&m[500]&m[501]&m[502]&~m[503])|(m[21]&m[500]&~m[501]&~m[502]&m[503])|(m[21]&~m[500]&m[501]&~m[502]&m[503])|(~m[21]&m[500]&m[501]&~m[502]&m[503])|(m[21]&~m[500]&~m[501]&m[502]&m[503])|(~m[21]&m[500]&~m[501]&m[502]&m[503])|(~m[21]&~m[500]&m[501]&m[502]&m[503]))&~BiasedRNG[341])|((m[21]&m[500]&m[501]&m[502]&~m[503])|(m[21]&m[500]&m[501]&~m[502]&m[503])|(m[21]&m[500]&~m[501]&m[502]&m[503])|(m[21]&~m[500]&m[501]&m[502]&m[503])|(~m[21]&m[500]&m[501]&m[502]&m[503])|(m[21]&m[500]&m[501]&m[502]&m[503]));
    m[118] = (((m[21]&m[504]&~m[505]&~m[506]&~m[507])|(m[21]&~m[504]&m[505]&~m[506]&~m[507])|(~m[21]&m[504]&m[505]&~m[506]&~m[507])|(m[21]&~m[504]&~m[505]&m[506]&~m[507])|(~m[21]&m[504]&~m[505]&m[506]&~m[507])|(~m[21]&~m[504]&m[505]&m[506]&~m[507])|(m[21]&~m[504]&~m[505]&~m[506]&m[507])|(~m[21]&m[504]&~m[505]&~m[506]&m[507])|(~m[21]&~m[504]&m[505]&~m[506]&m[507])|(~m[21]&~m[504]&~m[505]&m[506]&m[507]))&BiasedRNG[342])|(((m[21]&m[504]&m[505]&~m[506]&~m[507])|(m[21]&m[504]&~m[505]&m[506]&~m[507])|(m[21]&~m[504]&m[505]&m[506]&~m[507])|(~m[21]&m[504]&m[505]&m[506]&~m[507])|(m[21]&m[504]&~m[505]&~m[506]&m[507])|(m[21]&~m[504]&m[505]&~m[506]&m[507])|(~m[21]&m[504]&m[505]&~m[506]&m[507])|(m[21]&~m[504]&~m[505]&m[506]&m[507])|(~m[21]&m[504]&~m[505]&m[506]&m[507])|(~m[21]&~m[504]&m[505]&m[506]&m[507]))&~BiasedRNG[342])|((m[21]&m[504]&m[505]&m[506]&~m[507])|(m[21]&m[504]&m[505]&~m[506]&m[507])|(m[21]&m[504]&~m[505]&m[506]&m[507])|(m[21]&~m[504]&m[505]&m[506]&m[507])|(~m[21]&m[504]&m[505]&m[506]&m[507])|(m[21]&m[504]&m[505]&m[506]&m[507]));
    m[119] = (((m[21]&m[508]&~m[509]&~m[510]&~m[511])|(m[21]&~m[508]&m[509]&~m[510]&~m[511])|(~m[21]&m[508]&m[509]&~m[510]&~m[511])|(m[21]&~m[508]&~m[509]&m[510]&~m[511])|(~m[21]&m[508]&~m[509]&m[510]&~m[511])|(~m[21]&~m[508]&m[509]&m[510]&~m[511])|(m[21]&~m[508]&~m[509]&~m[510]&m[511])|(~m[21]&m[508]&~m[509]&~m[510]&m[511])|(~m[21]&~m[508]&m[509]&~m[510]&m[511])|(~m[21]&~m[508]&~m[509]&m[510]&m[511]))&BiasedRNG[343])|(((m[21]&m[508]&m[509]&~m[510]&~m[511])|(m[21]&m[508]&~m[509]&m[510]&~m[511])|(m[21]&~m[508]&m[509]&m[510]&~m[511])|(~m[21]&m[508]&m[509]&m[510]&~m[511])|(m[21]&m[508]&~m[509]&~m[510]&m[511])|(m[21]&~m[508]&m[509]&~m[510]&m[511])|(~m[21]&m[508]&m[509]&~m[510]&m[511])|(m[21]&~m[508]&~m[509]&m[510]&m[511])|(~m[21]&m[508]&~m[509]&m[510]&m[511])|(~m[21]&~m[508]&m[509]&m[510]&m[511]))&~BiasedRNG[343])|((m[21]&m[508]&m[509]&m[510]&~m[511])|(m[21]&m[508]&m[509]&~m[510]&m[511])|(m[21]&m[508]&~m[509]&m[510]&m[511])|(m[21]&~m[508]&m[509]&m[510]&m[511])|(~m[21]&m[508]&m[509]&m[510]&m[511])|(m[21]&m[508]&m[509]&m[510]&m[511]));
    m[120] = (((m[22]&m[512]&~m[513]&~m[514]&~m[515])|(m[22]&~m[512]&m[513]&~m[514]&~m[515])|(~m[22]&m[512]&m[513]&~m[514]&~m[515])|(m[22]&~m[512]&~m[513]&m[514]&~m[515])|(~m[22]&m[512]&~m[513]&m[514]&~m[515])|(~m[22]&~m[512]&m[513]&m[514]&~m[515])|(m[22]&~m[512]&~m[513]&~m[514]&m[515])|(~m[22]&m[512]&~m[513]&~m[514]&m[515])|(~m[22]&~m[512]&m[513]&~m[514]&m[515])|(~m[22]&~m[512]&~m[513]&m[514]&m[515]))&BiasedRNG[344])|(((m[22]&m[512]&m[513]&~m[514]&~m[515])|(m[22]&m[512]&~m[513]&m[514]&~m[515])|(m[22]&~m[512]&m[513]&m[514]&~m[515])|(~m[22]&m[512]&m[513]&m[514]&~m[515])|(m[22]&m[512]&~m[513]&~m[514]&m[515])|(m[22]&~m[512]&m[513]&~m[514]&m[515])|(~m[22]&m[512]&m[513]&~m[514]&m[515])|(m[22]&~m[512]&~m[513]&m[514]&m[515])|(~m[22]&m[512]&~m[513]&m[514]&m[515])|(~m[22]&~m[512]&m[513]&m[514]&m[515]))&~BiasedRNG[344])|((m[22]&m[512]&m[513]&m[514]&~m[515])|(m[22]&m[512]&m[513]&~m[514]&m[515])|(m[22]&m[512]&~m[513]&m[514]&m[515])|(m[22]&~m[512]&m[513]&m[514]&m[515])|(~m[22]&m[512]&m[513]&m[514]&m[515])|(m[22]&m[512]&m[513]&m[514]&m[515]));
    m[121] = (((m[22]&m[516]&~m[517]&~m[518]&~m[519])|(m[22]&~m[516]&m[517]&~m[518]&~m[519])|(~m[22]&m[516]&m[517]&~m[518]&~m[519])|(m[22]&~m[516]&~m[517]&m[518]&~m[519])|(~m[22]&m[516]&~m[517]&m[518]&~m[519])|(~m[22]&~m[516]&m[517]&m[518]&~m[519])|(m[22]&~m[516]&~m[517]&~m[518]&m[519])|(~m[22]&m[516]&~m[517]&~m[518]&m[519])|(~m[22]&~m[516]&m[517]&~m[518]&m[519])|(~m[22]&~m[516]&~m[517]&m[518]&m[519]))&BiasedRNG[345])|(((m[22]&m[516]&m[517]&~m[518]&~m[519])|(m[22]&m[516]&~m[517]&m[518]&~m[519])|(m[22]&~m[516]&m[517]&m[518]&~m[519])|(~m[22]&m[516]&m[517]&m[518]&~m[519])|(m[22]&m[516]&~m[517]&~m[518]&m[519])|(m[22]&~m[516]&m[517]&~m[518]&m[519])|(~m[22]&m[516]&m[517]&~m[518]&m[519])|(m[22]&~m[516]&~m[517]&m[518]&m[519])|(~m[22]&m[516]&~m[517]&m[518]&m[519])|(~m[22]&~m[516]&m[517]&m[518]&m[519]))&~BiasedRNG[345])|((m[22]&m[516]&m[517]&m[518]&~m[519])|(m[22]&m[516]&m[517]&~m[518]&m[519])|(m[22]&m[516]&~m[517]&m[518]&m[519])|(m[22]&~m[516]&m[517]&m[518]&m[519])|(~m[22]&m[516]&m[517]&m[518]&m[519])|(m[22]&m[516]&m[517]&m[518]&m[519]));
    m[122] = (((m[22]&m[520]&~m[521]&~m[522]&~m[523])|(m[22]&~m[520]&m[521]&~m[522]&~m[523])|(~m[22]&m[520]&m[521]&~m[522]&~m[523])|(m[22]&~m[520]&~m[521]&m[522]&~m[523])|(~m[22]&m[520]&~m[521]&m[522]&~m[523])|(~m[22]&~m[520]&m[521]&m[522]&~m[523])|(m[22]&~m[520]&~m[521]&~m[522]&m[523])|(~m[22]&m[520]&~m[521]&~m[522]&m[523])|(~m[22]&~m[520]&m[521]&~m[522]&m[523])|(~m[22]&~m[520]&~m[521]&m[522]&m[523]))&BiasedRNG[346])|(((m[22]&m[520]&m[521]&~m[522]&~m[523])|(m[22]&m[520]&~m[521]&m[522]&~m[523])|(m[22]&~m[520]&m[521]&m[522]&~m[523])|(~m[22]&m[520]&m[521]&m[522]&~m[523])|(m[22]&m[520]&~m[521]&~m[522]&m[523])|(m[22]&~m[520]&m[521]&~m[522]&m[523])|(~m[22]&m[520]&m[521]&~m[522]&m[523])|(m[22]&~m[520]&~m[521]&m[522]&m[523])|(~m[22]&m[520]&~m[521]&m[522]&m[523])|(~m[22]&~m[520]&m[521]&m[522]&m[523]))&~BiasedRNG[346])|((m[22]&m[520]&m[521]&m[522]&~m[523])|(m[22]&m[520]&m[521]&~m[522]&m[523])|(m[22]&m[520]&~m[521]&m[522]&m[523])|(m[22]&~m[520]&m[521]&m[522]&m[523])|(~m[22]&m[520]&m[521]&m[522]&m[523])|(m[22]&m[520]&m[521]&m[522]&m[523]));
    m[123] = (((m[22]&m[524]&~m[525]&~m[526]&~m[527])|(m[22]&~m[524]&m[525]&~m[526]&~m[527])|(~m[22]&m[524]&m[525]&~m[526]&~m[527])|(m[22]&~m[524]&~m[525]&m[526]&~m[527])|(~m[22]&m[524]&~m[525]&m[526]&~m[527])|(~m[22]&~m[524]&m[525]&m[526]&~m[527])|(m[22]&~m[524]&~m[525]&~m[526]&m[527])|(~m[22]&m[524]&~m[525]&~m[526]&m[527])|(~m[22]&~m[524]&m[525]&~m[526]&m[527])|(~m[22]&~m[524]&~m[525]&m[526]&m[527]))&BiasedRNG[347])|(((m[22]&m[524]&m[525]&~m[526]&~m[527])|(m[22]&m[524]&~m[525]&m[526]&~m[527])|(m[22]&~m[524]&m[525]&m[526]&~m[527])|(~m[22]&m[524]&m[525]&m[526]&~m[527])|(m[22]&m[524]&~m[525]&~m[526]&m[527])|(m[22]&~m[524]&m[525]&~m[526]&m[527])|(~m[22]&m[524]&m[525]&~m[526]&m[527])|(m[22]&~m[524]&~m[525]&m[526]&m[527])|(~m[22]&m[524]&~m[525]&m[526]&m[527])|(~m[22]&~m[524]&m[525]&m[526]&m[527]))&~BiasedRNG[347])|((m[22]&m[524]&m[525]&m[526]&~m[527])|(m[22]&m[524]&m[525]&~m[526]&m[527])|(m[22]&m[524]&~m[525]&m[526]&m[527])|(m[22]&~m[524]&m[525]&m[526]&m[527])|(~m[22]&m[524]&m[525]&m[526]&m[527])|(m[22]&m[524]&m[525]&m[526]&m[527]));
    m[124] = (((m[23]&m[528]&~m[529]&~m[530]&~m[531])|(m[23]&~m[528]&m[529]&~m[530]&~m[531])|(~m[23]&m[528]&m[529]&~m[530]&~m[531])|(m[23]&~m[528]&~m[529]&m[530]&~m[531])|(~m[23]&m[528]&~m[529]&m[530]&~m[531])|(~m[23]&~m[528]&m[529]&m[530]&~m[531])|(m[23]&~m[528]&~m[529]&~m[530]&m[531])|(~m[23]&m[528]&~m[529]&~m[530]&m[531])|(~m[23]&~m[528]&m[529]&~m[530]&m[531])|(~m[23]&~m[528]&~m[529]&m[530]&m[531]))&BiasedRNG[348])|(((m[23]&m[528]&m[529]&~m[530]&~m[531])|(m[23]&m[528]&~m[529]&m[530]&~m[531])|(m[23]&~m[528]&m[529]&m[530]&~m[531])|(~m[23]&m[528]&m[529]&m[530]&~m[531])|(m[23]&m[528]&~m[529]&~m[530]&m[531])|(m[23]&~m[528]&m[529]&~m[530]&m[531])|(~m[23]&m[528]&m[529]&~m[530]&m[531])|(m[23]&~m[528]&~m[529]&m[530]&m[531])|(~m[23]&m[528]&~m[529]&m[530]&m[531])|(~m[23]&~m[528]&m[529]&m[530]&m[531]))&~BiasedRNG[348])|((m[23]&m[528]&m[529]&m[530]&~m[531])|(m[23]&m[528]&m[529]&~m[530]&m[531])|(m[23]&m[528]&~m[529]&m[530]&m[531])|(m[23]&~m[528]&m[529]&m[530]&m[531])|(~m[23]&m[528]&m[529]&m[530]&m[531])|(m[23]&m[528]&m[529]&m[530]&m[531]));
    m[125] = (((m[23]&m[532]&~m[533]&~m[534]&~m[535])|(m[23]&~m[532]&m[533]&~m[534]&~m[535])|(~m[23]&m[532]&m[533]&~m[534]&~m[535])|(m[23]&~m[532]&~m[533]&m[534]&~m[535])|(~m[23]&m[532]&~m[533]&m[534]&~m[535])|(~m[23]&~m[532]&m[533]&m[534]&~m[535])|(m[23]&~m[532]&~m[533]&~m[534]&m[535])|(~m[23]&m[532]&~m[533]&~m[534]&m[535])|(~m[23]&~m[532]&m[533]&~m[534]&m[535])|(~m[23]&~m[532]&~m[533]&m[534]&m[535]))&BiasedRNG[349])|(((m[23]&m[532]&m[533]&~m[534]&~m[535])|(m[23]&m[532]&~m[533]&m[534]&~m[535])|(m[23]&~m[532]&m[533]&m[534]&~m[535])|(~m[23]&m[532]&m[533]&m[534]&~m[535])|(m[23]&m[532]&~m[533]&~m[534]&m[535])|(m[23]&~m[532]&m[533]&~m[534]&m[535])|(~m[23]&m[532]&m[533]&~m[534]&m[535])|(m[23]&~m[532]&~m[533]&m[534]&m[535])|(~m[23]&m[532]&~m[533]&m[534]&m[535])|(~m[23]&~m[532]&m[533]&m[534]&m[535]))&~BiasedRNG[349])|((m[23]&m[532]&m[533]&m[534]&~m[535])|(m[23]&m[532]&m[533]&~m[534]&m[535])|(m[23]&m[532]&~m[533]&m[534]&m[535])|(m[23]&~m[532]&m[533]&m[534]&m[535])|(~m[23]&m[532]&m[533]&m[534]&m[535])|(m[23]&m[532]&m[533]&m[534]&m[535]));
    m[126] = (((m[23]&m[536]&~m[537]&~m[538]&~m[539])|(m[23]&~m[536]&m[537]&~m[538]&~m[539])|(~m[23]&m[536]&m[537]&~m[538]&~m[539])|(m[23]&~m[536]&~m[537]&m[538]&~m[539])|(~m[23]&m[536]&~m[537]&m[538]&~m[539])|(~m[23]&~m[536]&m[537]&m[538]&~m[539])|(m[23]&~m[536]&~m[537]&~m[538]&m[539])|(~m[23]&m[536]&~m[537]&~m[538]&m[539])|(~m[23]&~m[536]&m[537]&~m[538]&m[539])|(~m[23]&~m[536]&~m[537]&m[538]&m[539]))&BiasedRNG[350])|(((m[23]&m[536]&m[537]&~m[538]&~m[539])|(m[23]&m[536]&~m[537]&m[538]&~m[539])|(m[23]&~m[536]&m[537]&m[538]&~m[539])|(~m[23]&m[536]&m[537]&m[538]&~m[539])|(m[23]&m[536]&~m[537]&~m[538]&m[539])|(m[23]&~m[536]&m[537]&~m[538]&m[539])|(~m[23]&m[536]&m[537]&~m[538]&m[539])|(m[23]&~m[536]&~m[537]&m[538]&m[539])|(~m[23]&m[536]&~m[537]&m[538]&m[539])|(~m[23]&~m[536]&m[537]&m[538]&m[539]))&~BiasedRNG[350])|((m[23]&m[536]&m[537]&m[538]&~m[539])|(m[23]&m[536]&m[537]&~m[538]&m[539])|(m[23]&m[536]&~m[537]&m[538]&m[539])|(m[23]&~m[536]&m[537]&m[538]&m[539])|(~m[23]&m[536]&m[537]&m[538]&m[539])|(m[23]&m[536]&m[537]&m[538]&m[539]));
    m[127] = (((m[23]&m[540]&~m[541]&~m[542]&~m[543])|(m[23]&~m[540]&m[541]&~m[542]&~m[543])|(~m[23]&m[540]&m[541]&~m[542]&~m[543])|(m[23]&~m[540]&~m[541]&m[542]&~m[543])|(~m[23]&m[540]&~m[541]&m[542]&~m[543])|(~m[23]&~m[540]&m[541]&m[542]&~m[543])|(m[23]&~m[540]&~m[541]&~m[542]&m[543])|(~m[23]&m[540]&~m[541]&~m[542]&m[543])|(~m[23]&~m[540]&m[541]&~m[542]&m[543])|(~m[23]&~m[540]&~m[541]&m[542]&m[543]))&BiasedRNG[351])|(((m[23]&m[540]&m[541]&~m[542]&~m[543])|(m[23]&m[540]&~m[541]&m[542]&~m[543])|(m[23]&~m[540]&m[541]&m[542]&~m[543])|(~m[23]&m[540]&m[541]&m[542]&~m[543])|(m[23]&m[540]&~m[541]&~m[542]&m[543])|(m[23]&~m[540]&m[541]&~m[542]&m[543])|(~m[23]&m[540]&m[541]&~m[542]&m[543])|(m[23]&~m[540]&~m[541]&m[542]&m[543])|(~m[23]&m[540]&~m[541]&m[542]&m[543])|(~m[23]&~m[540]&m[541]&m[542]&m[543]))&~BiasedRNG[351])|((m[23]&m[540]&m[541]&m[542]&~m[543])|(m[23]&m[540]&m[541]&~m[542]&m[543])|(m[23]&m[540]&~m[541]&m[542]&m[543])|(m[23]&~m[540]&m[541]&m[542]&m[543])|(~m[23]&m[540]&m[541]&m[542]&m[543])|(m[23]&m[540]&m[541]&m[542]&m[543]));
    m[128] = (((m[24]&m[544]&~m[545]&~m[546]&~m[547])|(m[24]&~m[544]&m[545]&~m[546]&~m[547])|(~m[24]&m[544]&m[545]&~m[546]&~m[547])|(m[24]&~m[544]&~m[545]&m[546]&~m[547])|(~m[24]&m[544]&~m[545]&m[546]&~m[547])|(~m[24]&~m[544]&m[545]&m[546]&~m[547])|(m[24]&~m[544]&~m[545]&~m[546]&m[547])|(~m[24]&m[544]&~m[545]&~m[546]&m[547])|(~m[24]&~m[544]&m[545]&~m[546]&m[547])|(~m[24]&~m[544]&~m[545]&m[546]&m[547]))&BiasedRNG[352])|(((m[24]&m[544]&m[545]&~m[546]&~m[547])|(m[24]&m[544]&~m[545]&m[546]&~m[547])|(m[24]&~m[544]&m[545]&m[546]&~m[547])|(~m[24]&m[544]&m[545]&m[546]&~m[547])|(m[24]&m[544]&~m[545]&~m[546]&m[547])|(m[24]&~m[544]&m[545]&~m[546]&m[547])|(~m[24]&m[544]&m[545]&~m[546]&m[547])|(m[24]&~m[544]&~m[545]&m[546]&m[547])|(~m[24]&m[544]&~m[545]&m[546]&m[547])|(~m[24]&~m[544]&m[545]&m[546]&m[547]))&~BiasedRNG[352])|((m[24]&m[544]&m[545]&m[546]&~m[547])|(m[24]&m[544]&m[545]&~m[546]&m[547])|(m[24]&m[544]&~m[545]&m[546]&m[547])|(m[24]&~m[544]&m[545]&m[546]&m[547])|(~m[24]&m[544]&m[545]&m[546]&m[547])|(m[24]&m[544]&m[545]&m[546]&m[547]));
    m[129] = (((m[24]&m[548]&~m[549]&~m[550]&~m[551])|(m[24]&~m[548]&m[549]&~m[550]&~m[551])|(~m[24]&m[548]&m[549]&~m[550]&~m[551])|(m[24]&~m[548]&~m[549]&m[550]&~m[551])|(~m[24]&m[548]&~m[549]&m[550]&~m[551])|(~m[24]&~m[548]&m[549]&m[550]&~m[551])|(m[24]&~m[548]&~m[549]&~m[550]&m[551])|(~m[24]&m[548]&~m[549]&~m[550]&m[551])|(~m[24]&~m[548]&m[549]&~m[550]&m[551])|(~m[24]&~m[548]&~m[549]&m[550]&m[551]))&BiasedRNG[353])|(((m[24]&m[548]&m[549]&~m[550]&~m[551])|(m[24]&m[548]&~m[549]&m[550]&~m[551])|(m[24]&~m[548]&m[549]&m[550]&~m[551])|(~m[24]&m[548]&m[549]&m[550]&~m[551])|(m[24]&m[548]&~m[549]&~m[550]&m[551])|(m[24]&~m[548]&m[549]&~m[550]&m[551])|(~m[24]&m[548]&m[549]&~m[550]&m[551])|(m[24]&~m[548]&~m[549]&m[550]&m[551])|(~m[24]&m[548]&~m[549]&m[550]&m[551])|(~m[24]&~m[548]&m[549]&m[550]&m[551]))&~BiasedRNG[353])|((m[24]&m[548]&m[549]&m[550]&~m[551])|(m[24]&m[548]&m[549]&~m[550]&m[551])|(m[24]&m[548]&~m[549]&m[550]&m[551])|(m[24]&~m[548]&m[549]&m[550]&m[551])|(~m[24]&m[548]&m[549]&m[550]&m[551])|(m[24]&m[548]&m[549]&m[550]&m[551]));
    m[130] = (((m[24]&m[552]&~m[553]&~m[554]&~m[555])|(m[24]&~m[552]&m[553]&~m[554]&~m[555])|(~m[24]&m[552]&m[553]&~m[554]&~m[555])|(m[24]&~m[552]&~m[553]&m[554]&~m[555])|(~m[24]&m[552]&~m[553]&m[554]&~m[555])|(~m[24]&~m[552]&m[553]&m[554]&~m[555])|(m[24]&~m[552]&~m[553]&~m[554]&m[555])|(~m[24]&m[552]&~m[553]&~m[554]&m[555])|(~m[24]&~m[552]&m[553]&~m[554]&m[555])|(~m[24]&~m[552]&~m[553]&m[554]&m[555]))&BiasedRNG[354])|(((m[24]&m[552]&m[553]&~m[554]&~m[555])|(m[24]&m[552]&~m[553]&m[554]&~m[555])|(m[24]&~m[552]&m[553]&m[554]&~m[555])|(~m[24]&m[552]&m[553]&m[554]&~m[555])|(m[24]&m[552]&~m[553]&~m[554]&m[555])|(m[24]&~m[552]&m[553]&~m[554]&m[555])|(~m[24]&m[552]&m[553]&~m[554]&m[555])|(m[24]&~m[552]&~m[553]&m[554]&m[555])|(~m[24]&m[552]&~m[553]&m[554]&m[555])|(~m[24]&~m[552]&m[553]&m[554]&m[555]))&~BiasedRNG[354])|((m[24]&m[552]&m[553]&m[554]&~m[555])|(m[24]&m[552]&m[553]&~m[554]&m[555])|(m[24]&m[552]&~m[553]&m[554]&m[555])|(m[24]&~m[552]&m[553]&m[554]&m[555])|(~m[24]&m[552]&m[553]&m[554]&m[555])|(m[24]&m[552]&m[553]&m[554]&m[555]));
    m[131] = (((m[24]&m[556]&~m[557]&~m[558]&~m[559])|(m[24]&~m[556]&m[557]&~m[558]&~m[559])|(~m[24]&m[556]&m[557]&~m[558]&~m[559])|(m[24]&~m[556]&~m[557]&m[558]&~m[559])|(~m[24]&m[556]&~m[557]&m[558]&~m[559])|(~m[24]&~m[556]&m[557]&m[558]&~m[559])|(m[24]&~m[556]&~m[557]&~m[558]&m[559])|(~m[24]&m[556]&~m[557]&~m[558]&m[559])|(~m[24]&~m[556]&m[557]&~m[558]&m[559])|(~m[24]&~m[556]&~m[557]&m[558]&m[559]))&BiasedRNG[355])|(((m[24]&m[556]&m[557]&~m[558]&~m[559])|(m[24]&m[556]&~m[557]&m[558]&~m[559])|(m[24]&~m[556]&m[557]&m[558]&~m[559])|(~m[24]&m[556]&m[557]&m[558]&~m[559])|(m[24]&m[556]&~m[557]&~m[558]&m[559])|(m[24]&~m[556]&m[557]&~m[558]&m[559])|(~m[24]&m[556]&m[557]&~m[558]&m[559])|(m[24]&~m[556]&~m[557]&m[558]&m[559])|(~m[24]&m[556]&~m[557]&m[558]&m[559])|(~m[24]&~m[556]&m[557]&m[558]&m[559]))&~BiasedRNG[355])|((m[24]&m[556]&m[557]&m[558]&~m[559])|(m[24]&m[556]&m[557]&~m[558]&m[559])|(m[24]&m[556]&~m[557]&m[558]&m[559])|(m[24]&~m[556]&m[557]&m[558]&m[559])|(~m[24]&m[556]&m[557]&m[558]&m[559])|(m[24]&m[556]&m[557]&m[558]&m[559]));
    m[132] = (((m[25]&m[560]&~m[561]&~m[562]&~m[563])|(m[25]&~m[560]&m[561]&~m[562]&~m[563])|(~m[25]&m[560]&m[561]&~m[562]&~m[563])|(m[25]&~m[560]&~m[561]&m[562]&~m[563])|(~m[25]&m[560]&~m[561]&m[562]&~m[563])|(~m[25]&~m[560]&m[561]&m[562]&~m[563])|(m[25]&~m[560]&~m[561]&~m[562]&m[563])|(~m[25]&m[560]&~m[561]&~m[562]&m[563])|(~m[25]&~m[560]&m[561]&~m[562]&m[563])|(~m[25]&~m[560]&~m[561]&m[562]&m[563]))&BiasedRNG[356])|(((m[25]&m[560]&m[561]&~m[562]&~m[563])|(m[25]&m[560]&~m[561]&m[562]&~m[563])|(m[25]&~m[560]&m[561]&m[562]&~m[563])|(~m[25]&m[560]&m[561]&m[562]&~m[563])|(m[25]&m[560]&~m[561]&~m[562]&m[563])|(m[25]&~m[560]&m[561]&~m[562]&m[563])|(~m[25]&m[560]&m[561]&~m[562]&m[563])|(m[25]&~m[560]&~m[561]&m[562]&m[563])|(~m[25]&m[560]&~m[561]&m[562]&m[563])|(~m[25]&~m[560]&m[561]&m[562]&m[563]))&~BiasedRNG[356])|((m[25]&m[560]&m[561]&m[562]&~m[563])|(m[25]&m[560]&m[561]&~m[562]&m[563])|(m[25]&m[560]&~m[561]&m[562]&m[563])|(m[25]&~m[560]&m[561]&m[562]&m[563])|(~m[25]&m[560]&m[561]&m[562]&m[563])|(m[25]&m[560]&m[561]&m[562]&m[563]));
    m[133] = (((m[25]&m[564]&~m[565]&~m[566]&~m[567])|(m[25]&~m[564]&m[565]&~m[566]&~m[567])|(~m[25]&m[564]&m[565]&~m[566]&~m[567])|(m[25]&~m[564]&~m[565]&m[566]&~m[567])|(~m[25]&m[564]&~m[565]&m[566]&~m[567])|(~m[25]&~m[564]&m[565]&m[566]&~m[567])|(m[25]&~m[564]&~m[565]&~m[566]&m[567])|(~m[25]&m[564]&~m[565]&~m[566]&m[567])|(~m[25]&~m[564]&m[565]&~m[566]&m[567])|(~m[25]&~m[564]&~m[565]&m[566]&m[567]))&BiasedRNG[357])|(((m[25]&m[564]&m[565]&~m[566]&~m[567])|(m[25]&m[564]&~m[565]&m[566]&~m[567])|(m[25]&~m[564]&m[565]&m[566]&~m[567])|(~m[25]&m[564]&m[565]&m[566]&~m[567])|(m[25]&m[564]&~m[565]&~m[566]&m[567])|(m[25]&~m[564]&m[565]&~m[566]&m[567])|(~m[25]&m[564]&m[565]&~m[566]&m[567])|(m[25]&~m[564]&~m[565]&m[566]&m[567])|(~m[25]&m[564]&~m[565]&m[566]&m[567])|(~m[25]&~m[564]&m[565]&m[566]&m[567]))&~BiasedRNG[357])|((m[25]&m[564]&m[565]&m[566]&~m[567])|(m[25]&m[564]&m[565]&~m[566]&m[567])|(m[25]&m[564]&~m[565]&m[566]&m[567])|(m[25]&~m[564]&m[565]&m[566]&m[567])|(~m[25]&m[564]&m[565]&m[566]&m[567])|(m[25]&m[564]&m[565]&m[566]&m[567]));
    m[134] = (((m[25]&m[568]&~m[569]&~m[570]&~m[571])|(m[25]&~m[568]&m[569]&~m[570]&~m[571])|(~m[25]&m[568]&m[569]&~m[570]&~m[571])|(m[25]&~m[568]&~m[569]&m[570]&~m[571])|(~m[25]&m[568]&~m[569]&m[570]&~m[571])|(~m[25]&~m[568]&m[569]&m[570]&~m[571])|(m[25]&~m[568]&~m[569]&~m[570]&m[571])|(~m[25]&m[568]&~m[569]&~m[570]&m[571])|(~m[25]&~m[568]&m[569]&~m[570]&m[571])|(~m[25]&~m[568]&~m[569]&m[570]&m[571]))&BiasedRNG[358])|(((m[25]&m[568]&m[569]&~m[570]&~m[571])|(m[25]&m[568]&~m[569]&m[570]&~m[571])|(m[25]&~m[568]&m[569]&m[570]&~m[571])|(~m[25]&m[568]&m[569]&m[570]&~m[571])|(m[25]&m[568]&~m[569]&~m[570]&m[571])|(m[25]&~m[568]&m[569]&~m[570]&m[571])|(~m[25]&m[568]&m[569]&~m[570]&m[571])|(m[25]&~m[568]&~m[569]&m[570]&m[571])|(~m[25]&m[568]&~m[569]&m[570]&m[571])|(~m[25]&~m[568]&m[569]&m[570]&m[571]))&~BiasedRNG[358])|((m[25]&m[568]&m[569]&m[570]&~m[571])|(m[25]&m[568]&m[569]&~m[570]&m[571])|(m[25]&m[568]&~m[569]&m[570]&m[571])|(m[25]&~m[568]&m[569]&m[570]&m[571])|(~m[25]&m[568]&m[569]&m[570]&m[571])|(m[25]&m[568]&m[569]&m[570]&m[571]));
    m[135] = (((m[25]&m[572]&~m[573]&~m[574]&~m[575])|(m[25]&~m[572]&m[573]&~m[574]&~m[575])|(~m[25]&m[572]&m[573]&~m[574]&~m[575])|(m[25]&~m[572]&~m[573]&m[574]&~m[575])|(~m[25]&m[572]&~m[573]&m[574]&~m[575])|(~m[25]&~m[572]&m[573]&m[574]&~m[575])|(m[25]&~m[572]&~m[573]&~m[574]&m[575])|(~m[25]&m[572]&~m[573]&~m[574]&m[575])|(~m[25]&~m[572]&m[573]&~m[574]&m[575])|(~m[25]&~m[572]&~m[573]&m[574]&m[575]))&BiasedRNG[359])|(((m[25]&m[572]&m[573]&~m[574]&~m[575])|(m[25]&m[572]&~m[573]&m[574]&~m[575])|(m[25]&~m[572]&m[573]&m[574]&~m[575])|(~m[25]&m[572]&m[573]&m[574]&~m[575])|(m[25]&m[572]&~m[573]&~m[574]&m[575])|(m[25]&~m[572]&m[573]&~m[574]&m[575])|(~m[25]&m[572]&m[573]&~m[574]&m[575])|(m[25]&~m[572]&~m[573]&m[574]&m[575])|(~m[25]&m[572]&~m[573]&m[574]&m[575])|(~m[25]&~m[572]&m[573]&m[574]&m[575]))&~BiasedRNG[359])|((m[25]&m[572]&m[573]&m[574]&~m[575])|(m[25]&m[572]&m[573]&~m[574]&m[575])|(m[25]&m[572]&~m[573]&m[574]&m[575])|(m[25]&~m[572]&m[573]&m[574]&m[575])|(~m[25]&m[572]&m[573]&m[574]&m[575])|(m[25]&m[572]&m[573]&m[574]&m[575]));
    m[136] = (((m[26]&m[576]&~m[577]&~m[578]&~m[579])|(m[26]&~m[576]&m[577]&~m[578]&~m[579])|(~m[26]&m[576]&m[577]&~m[578]&~m[579])|(m[26]&~m[576]&~m[577]&m[578]&~m[579])|(~m[26]&m[576]&~m[577]&m[578]&~m[579])|(~m[26]&~m[576]&m[577]&m[578]&~m[579])|(m[26]&~m[576]&~m[577]&~m[578]&m[579])|(~m[26]&m[576]&~m[577]&~m[578]&m[579])|(~m[26]&~m[576]&m[577]&~m[578]&m[579])|(~m[26]&~m[576]&~m[577]&m[578]&m[579]))&BiasedRNG[360])|(((m[26]&m[576]&m[577]&~m[578]&~m[579])|(m[26]&m[576]&~m[577]&m[578]&~m[579])|(m[26]&~m[576]&m[577]&m[578]&~m[579])|(~m[26]&m[576]&m[577]&m[578]&~m[579])|(m[26]&m[576]&~m[577]&~m[578]&m[579])|(m[26]&~m[576]&m[577]&~m[578]&m[579])|(~m[26]&m[576]&m[577]&~m[578]&m[579])|(m[26]&~m[576]&~m[577]&m[578]&m[579])|(~m[26]&m[576]&~m[577]&m[578]&m[579])|(~m[26]&~m[576]&m[577]&m[578]&m[579]))&~BiasedRNG[360])|((m[26]&m[576]&m[577]&m[578]&~m[579])|(m[26]&m[576]&m[577]&~m[578]&m[579])|(m[26]&m[576]&~m[577]&m[578]&m[579])|(m[26]&~m[576]&m[577]&m[578]&m[579])|(~m[26]&m[576]&m[577]&m[578]&m[579])|(m[26]&m[576]&m[577]&m[578]&m[579]));
    m[137] = (((m[26]&m[580]&~m[581]&~m[582]&~m[583])|(m[26]&~m[580]&m[581]&~m[582]&~m[583])|(~m[26]&m[580]&m[581]&~m[582]&~m[583])|(m[26]&~m[580]&~m[581]&m[582]&~m[583])|(~m[26]&m[580]&~m[581]&m[582]&~m[583])|(~m[26]&~m[580]&m[581]&m[582]&~m[583])|(m[26]&~m[580]&~m[581]&~m[582]&m[583])|(~m[26]&m[580]&~m[581]&~m[582]&m[583])|(~m[26]&~m[580]&m[581]&~m[582]&m[583])|(~m[26]&~m[580]&~m[581]&m[582]&m[583]))&BiasedRNG[361])|(((m[26]&m[580]&m[581]&~m[582]&~m[583])|(m[26]&m[580]&~m[581]&m[582]&~m[583])|(m[26]&~m[580]&m[581]&m[582]&~m[583])|(~m[26]&m[580]&m[581]&m[582]&~m[583])|(m[26]&m[580]&~m[581]&~m[582]&m[583])|(m[26]&~m[580]&m[581]&~m[582]&m[583])|(~m[26]&m[580]&m[581]&~m[582]&m[583])|(m[26]&~m[580]&~m[581]&m[582]&m[583])|(~m[26]&m[580]&~m[581]&m[582]&m[583])|(~m[26]&~m[580]&m[581]&m[582]&m[583]))&~BiasedRNG[361])|((m[26]&m[580]&m[581]&m[582]&~m[583])|(m[26]&m[580]&m[581]&~m[582]&m[583])|(m[26]&m[580]&~m[581]&m[582]&m[583])|(m[26]&~m[580]&m[581]&m[582]&m[583])|(~m[26]&m[580]&m[581]&m[582]&m[583])|(m[26]&m[580]&m[581]&m[582]&m[583]));
    m[138] = (((m[26]&m[584]&~m[585]&~m[586]&~m[587])|(m[26]&~m[584]&m[585]&~m[586]&~m[587])|(~m[26]&m[584]&m[585]&~m[586]&~m[587])|(m[26]&~m[584]&~m[585]&m[586]&~m[587])|(~m[26]&m[584]&~m[585]&m[586]&~m[587])|(~m[26]&~m[584]&m[585]&m[586]&~m[587])|(m[26]&~m[584]&~m[585]&~m[586]&m[587])|(~m[26]&m[584]&~m[585]&~m[586]&m[587])|(~m[26]&~m[584]&m[585]&~m[586]&m[587])|(~m[26]&~m[584]&~m[585]&m[586]&m[587]))&BiasedRNG[362])|(((m[26]&m[584]&m[585]&~m[586]&~m[587])|(m[26]&m[584]&~m[585]&m[586]&~m[587])|(m[26]&~m[584]&m[585]&m[586]&~m[587])|(~m[26]&m[584]&m[585]&m[586]&~m[587])|(m[26]&m[584]&~m[585]&~m[586]&m[587])|(m[26]&~m[584]&m[585]&~m[586]&m[587])|(~m[26]&m[584]&m[585]&~m[586]&m[587])|(m[26]&~m[584]&~m[585]&m[586]&m[587])|(~m[26]&m[584]&~m[585]&m[586]&m[587])|(~m[26]&~m[584]&m[585]&m[586]&m[587]))&~BiasedRNG[362])|((m[26]&m[584]&m[585]&m[586]&~m[587])|(m[26]&m[584]&m[585]&~m[586]&m[587])|(m[26]&m[584]&~m[585]&m[586]&m[587])|(m[26]&~m[584]&m[585]&m[586]&m[587])|(~m[26]&m[584]&m[585]&m[586]&m[587])|(m[26]&m[584]&m[585]&m[586]&m[587]));
    m[139] = (((m[26]&m[588]&~m[589]&~m[590]&~m[591])|(m[26]&~m[588]&m[589]&~m[590]&~m[591])|(~m[26]&m[588]&m[589]&~m[590]&~m[591])|(m[26]&~m[588]&~m[589]&m[590]&~m[591])|(~m[26]&m[588]&~m[589]&m[590]&~m[591])|(~m[26]&~m[588]&m[589]&m[590]&~m[591])|(m[26]&~m[588]&~m[589]&~m[590]&m[591])|(~m[26]&m[588]&~m[589]&~m[590]&m[591])|(~m[26]&~m[588]&m[589]&~m[590]&m[591])|(~m[26]&~m[588]&~m[589]&m[590]&m[591]))&BiasedRNG[363])|(((m[26]&m[588]&m[589]&~m[590]&~m[591])|(m[26]&m[588]&~m[589]&m[590]&~m[591])|(m[26]&~m[588]&m[589]&m[590]&~m[591])|(~m[26]&m[588]&m[589]&m[590]&~m[591])|(m[26]&m[588]&~m[589]&~m[590]&m[591])|(m[26]&~m[588]&m[589]&~m[590]&m[591])|(~m[26]&m[588]&m[589]&~m[590]&m[591])|(m[26]&~m[588]&~m[589]&m[590]&m[591])|(~m[26]&m[588]&~m[589]&m[590]&m[591])|(~m[26]&~m[588]&m[589]&m[590]&m[591]))&~BiasedRNG[363])|((m[26]&m[588]&m[589]&m[590]&~m[591])|(m[26]&m[588]&m[589]&~m[590]&m[591])|(m[26]&m[588]&~m[589]&m[590]&m[591])|(m[26]&~m[588]&m[589]&m[590]&m[591])|(~m[26]&m[588]&m[589]&m[590]&m[591])|(m[26]&m[588]&m[589]&m[590]&m[591]));
    m[140] = (((m[27]&m[592]&~m[593]&~m[594]&~m[595])|(m[27]&~m[592]&m[593]&~m[594]&~m[595])|(~m[27]&m[592]&m[593]&~m[594]&~m[595])|(m[27]&~m[592]&~m[593]&m[594]&~m[595])|(~m[27]&m[592]&~m[593]&m[594]&~m[595])|(~m[27]&~m[592]&m[593]&m[594]&~m[595])|(m[27]&~m[592]&~m[593]&~m[594]&m[595])|(~m[27]&m[592]&~m[593]&~m[594]&m[595])|(~m[27]&~m[592]&m[593]&~m[594]&m[595])|(~m[27]&~m[592]&~m[593]&m[594]&m[595]))&BiasedRNG[364])|(((m[27]&m[592]&m[593]&~m[594]&~m[595])|(m[27]&m[592]&~m[593]&m[594]&~m[595])|(m[27]&~m[592]&m[593]&m[594]&~m[595])|(~m[27]&m[592]&m[593]&m[594]&~m[595])|(m[27]&m[592]&~m[593]&~m[594]&m[595])|(m[27]&~m[592]&m[593]&~m[594]&m[595])|(~m[27]&m[592]&m[593]&~m[594]&m[595])|(m[27]&~m[592]&~m[593]&m[594]&m[595])|(~m[27]&m[592]&~m[593]&m[594]&m[595])|(~m[27]&~m[592]&m[593]&m[594]&m[595]))&~BiasedRNG[364])|((m[27]&m[592]&m[593]&m[594]&~m[595])|(m[27]&m[592]&m[593]&~m[594]&m[595])|(m[27]&m[592]&~m[593]&m[594]&m[595])|(m[27]&~m[592]&m[593]&m[594]&m[595])|(~m[27]&m[592]&m[593]&m[594]&m[595])|(m[27]&m[592]&m[593]&m[594]&m[595]));
    m[141] = (((m[27]&m[596]&~m[597]&~m[598]&~m[599])|(m[27]&~m[596]&m[597]&~m[598]&~m[599])|(~m[27]&m[596]&m[597]&~m[598]&~m[599])|(m[27]&~m[596]&~m[597]&m[598]&~m[599])|(~m[27]&m[596]&~m[597]&m[598]&~m[599])|(~m[27]&~m[596]&m[597]&m[598]&~m[599])|(m[27]&~m[596]&~m[597]&~m[598]&m[599])|(~m[27]&m[596]&~m[597]&~m[598]&m[599])|(~m[27]&~m[596]&m[597]&~m[598]&m[599])|(~m[27]&~m[596]&~m[597]&m[598]&m[599]))&BiasedRNG[365])|(((m[27]&m[596]&m[597]&~m[598]&~m[599])|(m[27]&m[596]&~m[597]&m[598]&~m[599])|(m[27]&~m[596]&m[597]&m[598]&~m[599])|(~m[27]&m[596]&m[597]&m[598]&~m[599])|(m[27]&m[596]&~m[597]&~m[598]&m[599])|(m[27]&~m[596]&m[597]&~m[598]&m[599])|(~m[27]&m[596]&m[597]&~m[598]&m[599])|(m[27]&~m[596]&~m[597]&m[598]&m[599])|(~m[27]&m[596]&~m[597]&m[598]&m[599])|(~m[27]&~m[596]&m[597]&m[598]&m[599]))&~BiasedRNG[365])|((m[27]&m[596]&m[597]&m[598]&~m[599])|(m[27]&m[596]&m[597]&~m[598]&m[599])|(m[27]&m[596]&~m[597]&m[598]&m[599])|(m[27]&~m[596]&m[597]&m[598]&m[599])|(~m[27]&m[596]&m[597]&m[598]&m[599])|(m[27]&m[596]&m[597]&m[598]&m[599]));
    m[142] = (((m[27]&m[600]&~m[601]&~m[602]&~m[603])|(m[27]&~m[600]&m[601]&~m[602]&~m[603])|(~m[27]&m[600]&m[601]&~m[602]&~m[603])|(m[27]&~m[600]&~m[601]&m[602]&~m[603])|(~m[27]&m[600]&~m[601]&m[602]&~m[603])|(~m[27]&~m[600]&m[601]&m[602]&~m[603])|(m[27]&~m[600]&~m[601]&~m[602]&m[603])|(~m[27]&m[600]&~m[601]&~m[602]&m[603])|(~m[27]&~m[600]&m[601]&~m[602]&m[603])|(~m[27]&~m[600]&~m[601]&m[602]&m[603]))&BiasedRNG[366])|(((m[27]&m[600]&m[601]&~m[602]&~m[603])|(m[27]&m[600]&~m[601]&m[602]&~m[603])|(m[27]&~m[600]&m[601]&m[602]&~m[603])|(~m[27]&m[600]&m[601]&m[602]&~m[603])|(m[27]&m[600]&~m[601]&~m[602]&m[603])|(m[27]&~m[600]&m[601]&~m[602]&m[603])|(~m[27]&m[600]&m[601]&~m[602]&m[603])|(m[27]&~m[600]&~m[601]&m[602]&m[603])|(~m[27]&m[600]&~m[601]&m[602]&m[603])|(~m[27]&~m[600]&m[601]&m[602]&m[603]))&~BiasedRNG[366])|((m[27]&m[600]&m[601]&m[602]&~m[603])|(m[27]&m[600]&m[601]&~m[602]&m[603])|(m[27]&m[600]&~m[601]&m[602]&m[603])|(m[27]&~m[600]&m[601]&m[602]&m[603])|(~m[27]&m[600]&m[601]&m[602]&m[603])|(m[27]&m[600]&m[601]&m[602]&m[603]));
    m[143] = (((m[27]&m[604]&~m[605]&~m[606]&~m[607])|(m[27]&~m[604]&m[605]&~m[606]&~m[607])|(~m[27]&m[604]&m[605]&~m[606]&~m[607])|(m[27]&~m[604]&~m[605]&m[606]&~m[607])|(~m[27]&m[604]&~m[605]&m[606]&~m[607])|(~m[27]&~m[604]&m[605]&m[606]&~m[607])|(m[27]&~m[604]&~m[605]&~m[606]&m[607])|(~m[27]&m[604]&~m[605]&~m[606]&m[607])|(~m[27]&~m[604]&m[605]&~m[606]&m[607])|(~m[27]&~m[604]&~m[605]&m[606]&m[607]))&BiasedRNG[367])|(((m[27]&m[604]&m[605]&~m[606]&~m[607])|(m[27]&m[604]&~m[605]&m[606]&~m[607])|(m[27]&~m[604]&m[605]&m[606]&~m[607])|(~m[27]&m[604]&m[605]&m[606]&~m[607])|(m[27]&m[604]&~m[605]&~m[606]&m[607])|(m[27]&~m[604]&m[605]&~m[606]&m[607])|(~m[27]&m[604]&m[605]&~m[606]&m[607])|(m[27]&~m[604]&~m[605]&m[606]&m[607])|(~m[27]&m[604]&~m[605]&m[606]&m[607])|(~m[27]&~m[604]&m[605]&m[606]&m[607]))&~BiasedRNG[367])|((m[27]&m[604]&m[605]&m[606]&~m[607])|(m[27]&m[604]&m[605]&~m[606]&m[607])|(m[27]&m[604]&~m[605]&m[606]&m[607])|(m[27]&~m[604]&m[605]&m[606]&m[607])|(~m[27]&m[604]&m[605]&m[606]&m[607])|(m[27]&m[604]&m[605]&m[606]&m[607]));
    m[144] = (((m[28]&m[608]&~m[609]&~m[610]&~m[611])|(m[28]&~m[608]&m[609]&~m[610]&~m[611])|(~m[28]&m[608]&m[609]&~m[610]&~m[611])|(m[28]&~m[608]&~m[609]&m[610]&~m[611])|(~m[28]&m[608]&~m[609]&m[610]&~m[611])|(~m[28]&~m[608]&m[609]&m[610]&~m[611])|(m[28]&~m[608]&~m[609]&~m[610]&m[611])|(~m[28]&m[608]&~m[609]&~m[610]&m[611])|(~m[28]&~m[608]&m[609]&~m[610]&m[611])|(~m[28]&~m[608]&~m[609]&m[610]&m[611]))&BiasedRNG[368])|(((m[28]&m[608]&m[609]&~m[610]&~m[611])|(m[28]&m[608]&~m[609]&m[610]&~m[611])|(m[28]&~m[608]&m[609]&m[610]&~m[611])|(~m[28]&m[608]&m[609]&m[610]&~m[611])|(m[28]&m[608]&~m[609]&~m[610]&m[611])|(m[28]&~m[608]&m[609]&~m[610]&m[611])|(~m[28]&m[608]&m[609]&~m[610]&m[611])|(m[28]&~m[608]&~m[609]&m[610]&m[611])|(~m[28]&m[608]&~m[609]&m[610]&m[611])|(~m[28]&~m[608]&m[609]&m[610]&m[611]))&~BiasedRNG[368])|((m[28]&m[608]&m[609]&m[610]&~m[611])|(m[28]&m[608]&m[609]&~m[610]&m[611])|(m[28]&m[608]&~m[609]&m[610]&m[611])|(m[28]&~m[608]&m[609]&m[610]&m[611])|(~m[28]&m[608]&m[609]&m[610]&m[611])|(m[28]&m[608]&m[609]&m[610]&m[611]));
    m[145] = (((m[28]&m[612]&~m[613]&~m[614]&~m[615])|(m[28]&~m[612]&m[613]&~m[614]&~m[615])|(~m[28]&m[612]&m[613]&~m[614]&~m[615])|(m[28]&~m[612]&~m[613]&m[614]&~m[615])|(~m[28]&m[612]&~m[613]&m[614]&~m[615])|(~m[28]&~m[612]&m[613]&m[614]&~m[615])|(m[28]&~m[612]&~m[613]&~m[614]&m[615])|(~m[28]&m[612]&~m[613]&~m[614]&m[615])|(~m[28]&~m[612]&m[613]&~m[614]&m[615])|(~m[28]&~m[612]&~m[613]&m[614]&m[615]))&BiasedRNG[369])|(((m[28]&m[612]&m[613]&~m[614]&~m[615])|(m[28]&m[612]&~m[613]&m[614]&~m[615])|(m[28]&~m[612]&m[613]&m[614]&~m[615])|(~m[28]&m[612]&m[613]&m[614]&~m[615])|(m[28]&m[612]&~m[613]&~m[614]&m[615])|(m[28]&~m[612]&m[613]&~m[614]&m[615])|(~m[28]&m[612]&m[613]&~m[614]&m[615])|(m[28]&~m[612]&~m[613]&m[614]&m[615])|(~m[28]&m[612]&~m[613]&m[614]&m[615])|(~m[28]&~m[612]&m[613]&m[614]&m[615]))&~BiasedRNG[369])|((m[28]&m[612]&m[613]&m[614]&~m[615])|(m[28]&m[612]&m[613]&~m[614]&m[615])|(m[28]&m[612]&~m[613]&m[614]&m[615])|(m[28]&~m[612]&m[613]&m[614]&m[615])|(~m[28]&m[612]&m[613]&m[614]&m[615])|(m[28]&m[612]&m[613]&m[614]&m[615]));
    m[146] = (((m[28]&m[616]&~m[617]&~m[618]&~m[619])|(m[28]&~m[616]&m[617]&~m[618]&~m[619])|(~m[28]&m[616]&m[617]&~m[618]&~m[619])|(m[28]&~m[616]&~m[617]&m[618]&~m[619])|(~m[28]&m[616]&~m[617]&m[618]&~m[619])|(~m[28]&~m[616]&m[617]&m[618]&~m[619])|(m[28]&~m[616]&~m[617]&~m[618]&m[619])|(~m[28]&m[616]&~m[617]&~m[618]&m[619])|(~m[28]&~m[616]&m[617]&~m[618]&m[619])|(~m[28]&~m[616]&~m[617]&m[618]&m[619]))&BiasedRNG[370])|(((m[28]&m[616]&m[617]&~m[618]&~m[619])|(m[28]&m[616]&~m[617]&m[618]&~m[619])|(m[28]&~m[616]&m[617]&m[618]&~m[619])|(~m[28]&m[616]&m[617]&m[618]&~m[619])|(m[28]&m[616]&~m[617]&~m[618]&m[619])|(m[28]&~m[616]&m[617]&~m[618]&m[619])|(~m[28]&m[616]&m[617]&~m[618]&m[619])|(m[28]&~m[616]&~m[617]&m[618]&m[619])|(~m[28]&m[616]&~m[617]&m[618]&m[619])|(~m[28]&~m[616]&m[617]&m[618]&m[619]))&~BiasedRNG[370])|((m[28]&m[616]&m[617]&m[618]&~m[619])|(m[28]&m[616]&m[617]&~m[618]&m[619])|(m[28]&m[616]&~m[617]&m[618]&m[619])|(m[28]&~m[616]&m[617]&m[618]&m[619])|(~m[28]&m[616]&m[617]&m[618]&m[619])|(m[28]&m[616]&m[617]&m[618]&m[619]));
    m[147] = (((m[28]&m[620]&~m[621]&~m[622]&~m[623])|(m[28]&~m[620]&m[621]&~m[622]&~m[623])|(~m[28]&m[620]&m[621]&~m[622]&~m[623])|(m[28]&~m[620]&~m[621]&m[622]&~m[623])|(~m[28]&m[620]&~m[621]&m[622]&~m[623])|(~m[28]&~m[620]&m[621]&m[622]&~m[623])|(m[28]&~m[620]&~m[621]&~m[622]&m[623])|(~m[28]&m[620]&~m[621]&~m[622]&m[623])|(~m[28]&~m[620]&m[621]&~m[622]&m[623])|(~m[28]&~m[620]&~m[621]&m[622]&m[623]))&BiasedRNG[371])|(((m[28]&m[620]&m[621]&~m[622]&~m[623])|(m[28]&m[620]&~m[621]&m[622]&~m[623])|(m[28]&~m[620]&m[621]&m[622]&~m[623])|(~m[28]&m[620]&m[621]&m[622]&~m[623])|(m[28]&m[620]&~m[621]&~m[622]&m[623])|(m[28]&~m[620]&m[621]&~m[622]&m[623])|(~m[28]&m[620]&m[621]&~m[622]&m[623])|(m[28]&~m[620]&~m[621]&m[622]&m[623])|(~m[28]&m[620]&~m[621]&m[622]&m[623])|(~m[28]&~m[620]&m[621]&m[622]&m[623]))&~BiasedRNG[371])|((m[28]&m[620]&m[621]&m[622]&~m[623])|(m[28]&m[620]&m[621]&~m[622]&m[623])|(m[28]&m[620]&~m[621]&m[622]&m[623])|(m[28]&~m[620]&m[621]&m[622]&m[623])|(~m[28]&m[620]&m[621]&m[622]&m[623])|(m[28]&m[620]&m[621]&m[622]&m[623]));
    m[148] = (((m[29]&m[624]&~m[625]&~m[626]&~m[627])|(m[29]&~m[624]&m[625]&~m[626]&~m[627])|(~m[29]&m[624]&m[625]&~m[626]&~m[627])|(m[29]&~m[624]&~m[625]&m[626]&~m[627])|(~m[29]&m[624]&~m[625]&m[626]&~m[627])|(~m[29]&~m[624]&m[625]&m[626]&~m[627])|(m[29]&~m[624]&~m[625]&~m[626]&m[627])|(~m[29]&m[624]&~m[625]&~m[626]&m[627])|(~m[29]&~m[624]&m[625]&~m[626]&m[627])|(~m[29]&~m[624]&~m[625]&m[626]&m[627]))&BiasedRNG[372])|(((m[29]&m[624]&m[625]&~m[626]&~m[627])|(m[29]&m[624]&~m[625]&m[626]&~m[627])|(m[29]&~m[624]&m[625]&m[626]&~m[627])|(~m[29]&m[624]&m[625]&m[626]&~m[627])|(m[29]&m[624]&~m[625]&~m[626]&m[627])|(m[29]&~m[624]&m[625]&~m[626]&m[627])|(~m[29]&m[624]&m[625]&~m[626]&m[627])|(m[29]&~m[624]&~m[625]&m[626]&m[627])|(~m[29]&m[624]&~m[625]&m[626]&m[627])|(~m[29]&~m[624]&m[625]&m[626]&m[627]))&~BiasedRNG[372])|((m[29]&m[624]&m[625]&m[626]&~m[627])|(m[29]&m[624]&m[625]&~m[626]&m[627])|(m[29]&m[624]&~m[625]&m[626]&m[627])|(m[29]&~m[624]&m[625]&m[626]&m[627])|(~m[29]&m[624]&m[625]&m[626]&m[627])|(m[29]&m[624]&m[625]&m[626]&m[627]));
    m[149] = (((m[29]&m[628]&~m[629]&~m[630]&~m[631])|(m[29]&~m[628]&m[629]&~m[630]&~m[631])|(~m[29]&m[628]&m[629]&~m[630]&~m[631])|(m[29]&~m[628]&~m[629]&m[630]&~m[631])|(~m[29]&m[628]&~m[629]&m[630]&~m[631])|(~m[29]&~m[628]&m[629]&m[630]&~m[631])|(m[29]&~m[628]&~m[629]&~m[630]&m[631])|(~m[29]&m[628]&~m[629]&~m[630]&m[631])|(~m[29]&~m[628]&m[629]&~m[630]&m[631])|(~m[29]&~m[628]&~m[629]&m[630]&m[631]))&BiasedRNG[373])|(((m[29]&m[628]&m[629]&~m[630]&~m[631])|(m[29]&m[628]&~m[629]&m[630]&~m[631])|(m[29]&~m[628]&m[629]&m[630]&~m[631])|(~m[29]&m[628]&m[629]&m[630]&~m[631])|(m[29]&m[628]&~m[629]&~m[630]&m[631])|(m[29]&~m[628]&m[629]&~m[630]&m[631])|(~m[29]&m[628]&m[629]&~m[630]&m[631])|(m[29]&~m[628]&~m[629]&m[630]&m[631])|(~m[29]&m[628]&~m[629]&m[630]&m[631])|(~m[29]&~m[628]&m[629]&m[630]&m[631]))&~BiasedRNG[373])|((m[29]&m[628]&m[629]&m[630]&~m[631])|(m[29]&m[628]&m[629]&~m[630]&m[631])|(m[29]&m[628]&~m[629]&m[630]&m[631])|(m[29]&~m[628]&m[629]&m[630]&m[631])|(~m[29]&m[628]&m[629]&m[630]&m[631])|(m[29]&m[628]&m[629]&m[630]&m[631]));
    m[150] = (((m[29]&m[632]&~m[633]&~m[634]&~m[635])|(m[29]&~m[632]&m[633]&~m[634]&~m[635])|(~m[29]&m[632]&m[633]&~m[634]&~m[635])|(m[29]&~m[632]&~m[633]&m[634]&~m[635])|(~m[29]&m[632]&~m[633]&m[634]&~m[635])|(~m[29]&~m[632]&m[633]&m[634]&~m[635])|(m[29]&~m[632]&~m[633]&~m[634]&m[635])|(~m[29]&m[632]&~m[633]&~m[634]&m[635])|(~m[29]&~m[632]&m[633]&~m[634]&m[635])|(~m[29]&~m[632]&~m[633]&m[634]&m[635]))&BiasedRNG[374])|(((m[29]&m[632]&m[633]&~m[634]&~m[635])|(m[29]&m[632]&~m[633]&m[634]&~m[635])|(m[29]&~m[632]&m[633]&m[634]&~m[635])|(~m[29]&m[632]&m[633]&m[634]&~m[635])|(m[29]&m[632]&~m[633]&~m[634]&m[635])|(m[29]&~m[632]&m[633]&~m[634]&m[635])|(~m[29]&m[632]&m[633]&~m[634]&m[635])|(m[29]&~m[632]&~m[633]&m[634]&m[635])|(~m[29]&m[632]&~m[633]&m[634]&m[635])|(~m[29]&~m[632]&m[633]&m[634]&m[635]))&~BiasedRNG[374])|((m[29]&m[632]&m[633]&m[634]&~m[635])|(m[29]&m[632]&m[633]&~m[634]&m[635])|(m[29]&m[632]&~m[633]&m[634]&m[635])|(m[29]&~m[632]&m[633]&m[634]&m[635])|(~m[29]&m[632]&m[633]&m[634]&m[635])|(m[29]&m[632]&m[633]&m[634]&m[635]));
    m[151] = (((m[29]&m[636]&~m[637]&~m[638]&~m[639])|(m[29]&~m[636]&m[637]&~m[638]&~m[639])|(~m[29]&m[636]&m[637]&~m[638]&~m[639])|(m[29]&~m[636]&~m[637]&m[638]&~m[639])|(~m[29]&m[636]&~m[637]&m[638]&~m[639])|(~m[29]&~m[636]&m[637]&m[638]&~m[639])|(m[29]&~m[636]&~m[637]&~m[638]&m[639])|(~m[29]&m[636]&~m[637]&~m[638]&m[639])|(~m[29]&~m[636]&m[637]&~m[638]&m[639])|(~m[29]&~m[636]&~m[637]&m[638]&m[639]))&BiasedRNG[375])|(((m[29]&m[636]&m[637]&~m[638]&~m[639])|(m[29]&m[636]&~m[637]&m[638]&~m[639])|(m[29]&~m[636]&m[637]&m[638]&~m[639])|(~m[29]&m[636]&m[637]&m[638]&~m[639])|(m[29]&m[636]&~m[637]&~m[638]&m[639])|(m[29]&~m[636]&m[637]&~m[638]&m[639])|(~m[29]&m[636]&m[637]&~m[638]&m[639])|(m[29]&~m[636]&~m[637]&m[638]&m[639])|(~m[29]&m[636]&~m[637]&m[638]&m[639])|(~m[29]&~m[636]&m[637]&m[638]&m[639]))&~BiasedRNG[375])|((m[29]&m[636]&m[637]&m[638]&~m[639])|(m[29]&m[636]&m[637]&~m[638]&m[639])|(m[29]&m[636]&~m[637]&m[638]&m[639])|(m[29]&~m[636]&m[637]&m[638]&m[639])|(~m[29]&m[636]&m[637]&m[638]&m[639])|(m[29]&m[636]&m[637]&m[638]&m[639]));
    m[152] = (((m[30]&m[640]&~m[641]&~m[642]&~m[643])|(m[30]&~m[640]&m[641]&~m[642]&~m[643])|(~m[30]&m[640]&m[641]&~m[642]&~m[643])|(m[30]&~m[640]&~m[641]&m[642]&~m[643])|(~m[30]&m[640]&~m[641]&m[642]&~m[643])|(~m[30]&~m[640]&m[641]&m[642]&~m[643])|(m[30]&~m[640]&~m[641]&~m[642]&m[643])|(~m[30]&m[640]&~m[641]&~m[642]&m[643])|(~m[30]&~m[640]&m[641]&~m[642]&m[643])|(~m[30]&~m[640]&~m[641]&m[642]&m[643]))&BiasedRNG[376])|(((m[30]&m[640]&m[641]&~m[642]&~m[643])|(m[30]&m[640]&~m[641]&m[642]&~m[643])|(m[30]&~m[640]&m[641]&m[642]&~m[643])|(~m[30]&m[640]&m[641]&m[642]&~m[643])|(m[30]&m[640]&~m[641]&~m[642]&m[643])|(m[30]&~m[640]&m[641]&~m[642]&m[643])|(~m[30]&m[640]&m[641]&~m[642]&m[643])|(m[30]&~m[640]&~m[641]&m[642]&m[643])|(~m[30]&m[640]&~m[641]&m[642]&m[643])|(~m[30]&~m[640]&m[641]&m[642]&m[643]))&~BiasedRNG[376])|((m[30]&m[640]&m[641]&m[642]&~m[643])|(m[30]&m[640]&m[641]&~m[642]&m[643])|(m[30]&m[640]&~m[641]&m[642]&m[643])|(m[30]&~m[640]&m[641]&m[642]&m[643])|(~m[30]&m[640]&m[641]&m[642]&m[643])|(m[30]&m[640]&m[641]&m[642]&m[643]));
    m[153] = (((m[30]&m[644]&~m[645]&~m[646]&~m[647])|(m[30]&~m[644]&m[645]&~m[646]&~m[647])|(~m[30]&m[644]&m[645]&~m[646]&~m[647])|(m[30]&~m[644]&~m[645]&m[646]&~m[647])|(~m[30]&m[644]&~m[645]&m[646]&~m[647])|(~m[30]&~m[644]&m[645]&m[646]&~m[647])|(m[30]&~m[644]&~m[645]&~m[646]&m[647])|(~m[30]&m[644]&~m[645]&~m[646]&m[647])|(~m[30]&~m[644]&m[645]&~m[646]&m[647])|(~m[30]&~m[644]&~m[645]&m[646]&m[647]))&BiasedRNG[377])|(((m[30]&m[644]&m[645]&~m[646]&~m[647])|(m[30]&m[644]&~m[645]&m[646]&~m[647])|(m[30]&~m[644]&m[645]&m[646]&~m[647])|(~m[30]&m[644]&m[645]&m[646]&~m[647])|(m[30]&m[644]&~m[645]&~m[646]&m[647])|(m[30]&~m[644]&m[645]&~m[646]&m[647])|(~m[30]&m[644]&m[645]&~m[646]&m[647])|(m[30]&~m[644]&~m[645]&m[646]&m[647])|(~m[30]&m[644]&~m[645]&m[646]&m[647])|(~m[30]&~m[644]&m[645]&m[646]&m[647]))&~BiasedRNG[377])|((m[30]&m[644]&m[645]&m[646]&~m[647])|(m[30]&m[644]&m[645]&~m[646]&m[647])|(m[30]&m[644]&~m[645]&m[646]&m[647])|(m[30]&~m[644]&m[645]&m[646]&m[647])|(~m[30]&m[644]&m[645]&m[646]&m[647])|(m[30]&m[644]&m[645]&m[646]&m[647]));
    m[154] = (((m[30]&m[648]&~m[649]&~m[650]&~m[651])|(m[30]&~m[648]&m[649]&~m[650]&~m[651])|(~m[30]&m[648]&m[649]&~m[650]&~m[651])|(m[30]&~m[648]&~m[649]&m[650]&~m[651])|(~m[30]&m[648]&~m[649]&m[650]&~m[651])|(~m[30]&~m[648]&m[649]&m[650]&~m[651])|(m[30]&~m[648]&~m[649]&~m[650]&m[651])|(~m[30]&m[648]&~m[649]&~m[650]&m[651])|(~m[30]&~m[648]&m[649]&~m[650]&m[651])|(~m[30]&~m[648]&~m[649]&m[650]&m[651]))&BiasedRNG[378])|(((m[30]&m[648]&m[649]&~m[650]&~m[651])|(m[30]&m[648]&~m[649]&m[650]&~m[651])|(m[30]&~m[648]&m[649]&m[650]&~m[651])|(~m[30]&m[648]&m[649]&m[650]&~m[651])|(m[30]&m[648]&~m[649]&~m[650]&m[651])|(m[30]&~m[648]&m[649]&~m[650]&m[651])|(~m[30]&m[648]&m[649]&~m[650]&m[651])|(m[30]&~m[648]&~m[649]&m[650]&m[651])|(~m[30]&m[648]&~m[649]&m[650]&m[651])|(~m[30]&~m[648]&m[649]&m[650]&m[651]))&~BiasedRNG[378])|((m[30]&m[648]&m[649]&m[650]&~m[651])|(m[30]&m[648]&m[649]&~m[650]&m[651])|(m[30]&m[648]&~m[649]&m[650]&m[651])|(m[30]&~m[648]&m[649]&m[650]&m[651])|(~m[30]&m[648]&m[649]&m[650]&m[651])|(m[30]&m[648]&m[649]&m[650]&m[651]));
    m[155] = (((m[30]&m[652]&~m[653]&~m[654]&~m[655])|(m[30]&~m[652]&m[653]&~m[654]&~m[655])|(~m[30]&m[652]&m[653]&~m[654]&~m[655])|(m[30]&~m[652]&~m[653]&m[654]&~m[655])|(~m[30]&m[652]&~m[653]&m[654]&~m[655])|(~m[30]&~m[652]&m[653]&m[654]&~m[655])|(m[30]&~m[652]&~m[653]&~m[654]&m[655])|(~m[30]&m[652]&~m[653]&~m[654]&m[655])|(~m[30]&~m[652]&m[653]&~m[654]&m[655])|(~m[30]&~m[652]&~m[653]&m[654]&m[655]))&BiasedRNG[379])|(((m[30]&m[652]&m[653]&~m[654]&~m[655])|(m[30]&m[652]&~m[653]&m[654]&~m[655])|(m[30]&~m[652]&m[653]&m[654]&~m[655])|(~m[30]&m[652]&m[653]&m[654]&~m[655])|(m[30]&m[652]&~m[653]&~m[654]&m[655])|(m[30]&~m[652]&m[653]&~m[654]&m[655])|(~m[30]&m[652]&m[653]&~m[654]&m[655])|(m[30]&~m[652]&~m[653]&m[654]&m[655])|(~m[30]&m[652]&~m[653]&m[654]&m[655])|(~m[30]&~m[652]&m[653]&m[654]&m[655]))&~BiasedRNG[379])|((m[30]&m[652]&m[653]&m[654]&~m[655])|(m[30]&m[652]&m[653]&~m[654]&m[655])|(m[30]&m[652]&~m[653]&m[654]&m[655])|(m[30]&~m[652]&m[653]&m[654]&m[655])|(~m[30]&m[652]&m[653]&m[654]&m[655])|(m[30]&m[652]&m[653]&m[654]&m[655]));
    m[156] = (((m[31]&m[656]&~m[657]&~m[658]&~m[659])|(m[31]&~m[656]&m[657]&~m[658]&~m[659])|(~m[31]&m[656]&m[657]&~m[658]&~m[659])|(m[31]&~m[656]&~m[657]&m[658]&~m[659])|(~m[31]&m[656]&~m[657]&m[658]&~m[659])|(~m[31]&~m[656]&m[657]&m[658]&~m[659])|(m[31]&~m[656]&~m[657]&~m[658]&m[659])|(~m[31]&m[656]&~m[657]&~m[658]&m[659])|(~m[31]&~m[656]&m[657]&~m[658]&m[659])|(~m[31]&~m[656]&~m[657]&m[658]&m[659]))&BiasedRNG[380])|(((m[31]&m[656]&m[657]&~m[658]&~m[659])|(m[31]&m[656]&~m[657]&m[658]&~m[659])|(m[31]&~m[656]&m[657]&m[658]&~m[659])|(~m[31]&m[656]&m[657]&m[658]&~m[659])|(m[31]&m[656]&~m[657]&~m[658]&m[659])|(m[31]&~m[656]&m[657]&~m[658]&m[659])|(~m[31]&m[656]&m[657]&~m[658]&m[659])|(m[31]&~m[656]&~m[657]&m[658]&m[659])|(~m[31]&m[656]&~m[657]&m[658]&m[659])|(~m[31]&~m[656]&m[657]&m[658]&m[659]))&~BiasedRNG[380])|((m[31]&m[656]&m[657]&m[658]&~m[659])|(m[31]&m[656]&m[657]&~m[658]&m[659])|(m[31]&m[656]&~m[657]&m[658]&m[659])|(m[31]&~m[656]&m[657]&m[658]&m[659])|(~m[31]&m[656]&m[657]&m[658]&m[659])|(m[31]&m[656]&m[657]&m[658]&m[659]));
    m[157] = (((m[31]&m[660]&~m[661]&~m[662]&~m[663])|(m[31]&~m[660]&m[661]&~m[662]&~m[663])|(~m[31]&m[660]&m[661]&~m[662]&~m[663])|(m[31]&~m[660]&~m[661]&m[662]&~m[663])|(~m[31]&m[660]&~m[661]&m[662]&~m[663])|(~m[31]&~m[660]&m[661]&m[662]&~m[663])|(m[31]&~m[660]&~m[661]&~m[662]&m[663])|(~m[31]&m[660]&~m[661]&~m[662]&m[663])|(~m[31]&~m[660]&m[661]&~m[662]&m[663])|(~m[31]&~m[660]&~m[661]&m[662]&m[663]))&BiasedRNG[381])|(((m[31]&m[660]&m[661]&~m[662]&~m[663])|(m[31]&m[660]&~m[661]&m[662]&~m[663])|(m[31]&~m[660]&m[661]&m[662]&~m[663])|(~m[31]&m[660]&m[661]&m[662]&~m[663])|(m[31]&m[660]&~m[661]&~m[662]&m[663])|(m[31]&~m[660]&m[661]&~m[662]&m[663])|(~m[31]&m[660]&m[661]&~m[662]&m[663])|(m[31]&~m[660]&~m[661]&m[662]&m[663])|(~m[31]&m[660]&~m[661]&m[662]&m[663])|(~m[31]&~m[660]&m[661]&m[662]&m[663]))&~BiasedRNG[381])|((m[31]&m[660]&m[661]&m[662]&~m[663])|(m[31]&m[660]&m[661]&~m[662]&m[663])|(m[31]&m[660]&~m[661]&m[662]&m[663])|(m[31]&~m[660]&m[661]&m[662]&m[663])|(~m[31]&m[660]&m[661]&m[662]&m[663])|(m[31]&m[660]&m[661]&m[662]&m[663]));
    m[158] = (((m[31]&m[664]&~m[665]&~m[666]&~m[667])|(m[31]&~m[664]&m[665]&~m[666]&~m[667])|(~m[31]&m[664]&m[665]&~m[666]&~m[667])|(m[31]&~m[664]&~m[665]&m[666]&~m[667])|(~m[31]&m[664]&~m[665]&m[666]&~m[667])|(~m[31]&~m[664]&m[665]&m[666]&~m[667])|(m[31]&~m[664]&~m[665]&~m[666]&m[667])|(~m[31]&m[664]&~m[665]&~m[666]&m[667])|(~m[31]&~m[664]&m[665]&~m[666]&m[667])|(~m[31]&~m[664]&~m[665]&m[666]&m[667]))&BiasedRNG[382])|(((m[31]&m[664]&m[665]&~m[666]&~m[667])|(m[31]&m[664]&~m[665]&m[666]&~m[667])|(m[31]&~m[664]&m[665]&m[666]&~m[667])|(~m[31]&m[664]&m[665]&m[666]&~m[667])|(m[31]&m[664]&~m[665]&~m[666]&m[667])|(m[31]&~m[664]&m[665]&~m[666]&m[667])|(~m[31]&m[664]&m[665]&~m[666]&m[667])|(m[31]&~m[664]&~m[665]&m[666]&m[667])|(~m[31]&m[664]&~m[665]&m[666]&m[667])|(~m[31]&~m[664]&m[665]&m[666]&m[667]))&~BiasedRNG[382])|((m[31]&m[664]&m[665]&m[666]&~m[667])|(m[31]&m[664]&m[665]&~m[666]&m[667])|(m[31]&m[664]&~m[665]&m[666]&m[667])|(m[31]&~m[664]&m[665]&m[666]&m[667])|(~m[31]&m[664]&m[665]&m[666]&m[667])|(m[31]&m[664]&m[665]&m[666]&m[667]));
    m[159] = (((m[31]&m[668]&~m[669]&~m[670]&~m[671])|(m[31]&~m[668]&m[669]&~m[670]&~m[671])|(~m[31]&m[668]&m[669]&~m[670]&~m[671])|(m[31]&~m[668]&~m[669]&m[670]&~m[671])|(~m[31]&m[668]&~m[669]&m[670]&~m[671])|(~m[31]&~m[668]&m[669]&m[670]&~m[671])|(m[31]&~m[668]&~m[669]&~m[670]&m[671])|(~m[31]&m[668]&~m[669]&~m[670]&m[671])|(~m[31]&~m[668]&m[669]&~m[670]&m[671])|(~m[31]&~m[668]&~m[669]&m[670]&m[671]))&BiasedRNG[383])|(((m[31]&m[668]&m[669]&~m[670]&~m[671])|(m[31]&m[668]&~m[669]&m[670]&~m[671])|(m[31]&~m[668]&m[669]&m[670]&~m[671])|(~m[31]&m[668]&m[669]&m[670]&~m[671])|(m[31]&m[668]&~m[669]&~m[670]&m[671])|(m[31]&~m[668]&m[669]&~m[670]&m[671])|(~m[31]&m[668]&m[669]&~m[670]&m[671])|(m[31]&~m[668]&~m[669]&m[670]&m[671])|(~m[31]&m[668]&~m[669]&m[670]&m[671])|(~m[31]&~m[668]&m[669]&m[670]&m[671]))&~BiasedRNG[383])|((m[31]&m[668]&m[669]&m[670]&~m[671])|(m[31]&m[668]&m[669]&~m[670]&m[671])|(m[31]&m[668]&~m[669]&m[670]&m[671])|(m[31]&~m[668]&m[669]&m[670]&m[671])|(~m[31]&m[668]&m[669]&m[670]&m[671])|(m[31]&m[668]&m[669]&m[670]&m[671]));
    m[673] = (((m[176]&~m[417]&m[928])|(~m[176]&m[417]&m[928]))&BiasedRNG[384])|(((m[176]&m[417]&~m[928]))&~BiasedRNG[384])|((m[176]&m[417]&m[928]));
    m[674] = (((m[192]&~m[418]&m[933])|(~m[192]&m[418]&m[933]))&BiasedRNG[385])|(((m[192]&m[418]&~m[933]))&~BiasedRNG[385])|((m[192]&m[418]&m[933]));
    m[675] = (((m[208]&~m[419]&m[943])|(~m[208]&m[419]&m[943]))&BiasedRNG[386])|(((m[208]&m[419]&~m[943]))&~BiasedRNG[386])|((m[208]&m[419]&m[943]));
    m[676] = (((m[224]&~m[420]&m[958])|(~m[224]&m[420]&m[958]))&BiasedRNG[387])|(((m[224]&m[420]&~m[958]))&~BiasedRNG[387])|((m[224]&m[420]&m[958]));
    m[677] = (((m[240]&~m[421]&m[978])|(~m[240]&m[421]&m[978]))&BiasedRNG[388])|(((m[240]&m[421]&~m[978]))&~BiasedRNG[388])|((m[240]&m[421]&m[978]));
    m[678] = (((m[256]&~m[422]&m[1003])|(~m[256]&m[422]&m[1003]))&BiasedRNG[389])|(((m[256]&m[422]&~m[1003]))&~BiasedRNG[389])|((m[256]&m[422]&m[1003]));
    m[679] = (((m[272]&~m[423]&m[1033])|(~m[272]&m[423]&m[1033]))&BiasedRNG[390])|(((m[272]&m[423]&~m[1033]))&~BiasedRNG[390])|((m[272]&m[423]&m[1033]));
    m[680] = (((m[288]&~m[424]&m[1068])|(~m[288]&m[424]&m[1068]))&BiasedRNG[391])|(((m[288]&m[424]&~m[1068]))&~BiasedRNG[391])|((m[288]&m[424]&m[1068]));
    m[681] = (((m[304]&~m[425]&m[1108])|(~m[304]&m[425]&m[1108]))&BiasedRNG[392])|(((m[304]&m[425]&~m[1108]))&~BiasedRNG[392])|((m[304]&m[425]&m[1108]));
    m[682] = (((m[320]&~m[426]&m[1153])|(~m[320]&m[426]&m[1153]))&BiasedRNG[393])|(((m[320]&m[426]&~m[1153]))&~BiasedRNG[393])|((m[320]&m[426]&m[1153]));
    m[683] = (((m[336]&~m[427]&m[1203])|(~m[336]&m[427]&m[1203]))&BiasedRNG[394])|(((m[336]&m[427]&~m[1203]))&~BiasedRNG[394])|((m[336]&m[427]&m[1203]));
    m[684] = (((m[352]&~m[428]&m[1258])|(~m[352]&m[428]&m[1258]))&BiasedRNG[395])|(((m[352]&m[428]&~m[1258]))&~BiasedRNG[395])|((m[352]&m[428]&m[1258]));
    m[685] = (((m[368]&~m[429]&m[1318])|(~m[368]&m[429]&m[1318]))&BiasedRNG[396])|(((m[368]&m[429]&~m[1318]))&~BiasedRNG[396])|((m[368]&m[429]&m[1318]));
    m[686] = (((m[384]&~m[430]&m[1383])|(~m[384]&m[430]&m[1383]))&BiasedRNG[397])|(((m[384]&m[430]&~m[1383]))&~BiasedRNG[397])|((m[384]&m[430]&m[1383]));
    m[687] = (((m[400]&~m[431]&m[1453])|(~m[400]&m[431]&m[1453]))&BiasedRNG[398])|(((m[400]&m[431]&~m[1453]))&~BiasedRNG[398])|((m[400]&m[431]&m[1453]));
    m[688] = (((m[161]&~m[432]&m[929])|(~m[161]&m[432]&m[929]))&BiasedRNG[399])|(((m[161]&m[432]&~m[929]))&~BiasedRNG[399])|((m[161]&m[432]&m[929]));
    m[689] = (((m[177]&~m[433]&m[934])|(~m[177]&m[433]&m[934]))&BiasedRNG[400])|(((m[177]&m[433]&~m[934]))&~BiasedRNG[400])|((m[177]&m[433]&m[934]));
    m[690] = (((m[193]&~m[434]&m[944])|(~m[193]&m[434]&m[944]))&BiasedRNG[401])|(((m[193]&m[434]&~m[944]))&~BiasedRNG[401])|((m[193]&m[434]&m[944]));
    m[691] = (((m[209]&~m[435]&m[959])|(~m[209]&m[435]&m[959]))&BiasedRNG[402])|(((m[209]&m[435]&~m[959]))&~BiasedRNG[402])|((m[209]&m[435]&m[959]));
    m[692] = (((m[225]&~m[436]&m[979])|(~m[225]&m[436]&m[979]))&BiasedRNG[403])|(((m[225]&m[436]&~m[979]))&~BiasedRNG[403])|((m[225]&m[436]&m[979]));
    m[693] = (((m[241]&~m[437]&m[1004])|(~m[241]&m[437]&m[1004]))&BiasedRNG[404])|(((m[241]&m[437]&~m[1004]))&~BiasedRNG[404])|((m[241]&m[437]&m[1004]));
    m[694] = (((m[257]&~m[438]&m[1034])|(~m[257]&m[438]&m[1034]))&BiasedRNG[405])|(((m[257]&m[438]&~m[1034]))&~BiasedRNG[405])|((m[257]&m[438]&m[1034]));
    m[695] = (((m[273]&~m[439]&m[1069])|(~m[273]&m[439]&m[1069]))&BiasedRNG[406])|(((m[273]&m[439]&~m[1069]))&~BiasedRNG[406])|((m[273]&m[439]&m[1069]));
    m[696] = (((m[289]&~m[440]&m[1109])|(~m[289]&m[440]&m[1109]))&BiasedRNG[407])|(((m[289]&m[440]&~m[1109]))&~BiasedRNG[407])|((m[289]&m[440]&m[1109]));
    m[697] = (((m[305]&~m[441]&m[1154])|(~m[305]&m[441]&m[1154]))&BiasedRNG[408])|(((m[305]&m[441]&~m[1154]))&~BiasedRNG[408])|((m[305]&m[441]&m[1154]));
    m[698] = (((m[321]&~m[442]&m[1204])|(~m[321]&m[442]&m[1204]))&BiasedRNG[409])|(((m[321]&m[442]&~m[1204]))&~BiasedRNG[409])|((m[321]&m[442]&m[1204]));
    m[699] = (((m[337]&~m[443]&m[1259])|(~m[337]&m[443]&m[1259]))&BiasedRNG[410])|(((m[337]&m[443]&~m[1259]))&~BiasedRNG[410])|((m[337]&m[443]&m[1259]));
    m[700] = (((m[353]&~m[444]&m[1319])|(~m[353]&m[444]&m[1319]))&BiasedRNG[411])|(((m[353]&m[444]&~m[1319]))&~BiasedRNG[411])|((m[353]&m[444]&m[1319]));
    m[701] = (((m[369]&~m[445]&m[1384])|(~m[369]&m[445]&m[1384]))&BiasedRNG[412])|(((m[369]&m[445]&~m[1384]))&~BiasedRNG[412])|((m[369]&m[445]&m[1384]));
    m[702] = (((m[385]&~m[446]&m[1454])|(~m[385]&m[446]&m[1454]))&BiasedRNG[413])|(((m[385]&m[446]&~m[1454]))&~BiasedRNG[413])|((m[385]&m[446]&m[1454]));
    m[703] = (((m[401]&~m[447]&m[1529])|(~m[401]&m[447]&m[1529]))&BiasedRNG[414])|(((m[401]&m[447]&~m[1529]))&~BiasedRNG[414])|((m[401]&m[447]&m[1529]));
    m[704] = (((m[162]&~m[448]&m[939])|(~m[162]&m[448]&m[939]))&BiasedRNG[415])|(((m[162]&m[448]&~m[939]))&~BiasedRNG[415])|((m[162]&m[448]&m[939]));
    m[705] = (((m[178]&~m[449]&m[949])|(~m[178]&m[449]&m[949]))&BiasedRNG[416])|(((m[178]&m[449]&~m[949]))&~BiasedRNG[416])|((m[178]&m[449]&m[949]));
    m[706] = (((m[194]&~m[450]&m[964])|(~m[194]&m[450]&m[964]))&BiasedRNG[417])|(((m[194]&m[450]&~m[964]))&~BiasedRNG[417])|((m[194]&m[450]&m[964]));
    m[707] = (((m[210]&~m[451]&m[984])|(~m[210]&m[451]&m[984]))&BiasedRNG[418])|(((m[210]&m[451]&~m[984]))&~BiasedRNG[418])|((m[210]&m[451]&m[984]));
    m[708] = (((m[226]&~m[452]&m[1009])|(~m[226]&m[452]&m[1009]))&BiasedRNG[419])|(((m[226]&m[452]&~m[1009]))&~BiasedRNG[419])|((m[226]&m[452]&m[1009]));
    m[709] = (((m[242]&~m[453]&m[1039])|(~m[242]&m[453]&m[1039]))&BiasedRNG[420])|(((m[242]&m[453]&~m[1039]))&~BiasedRNG[420])|((m[242]&m[453]&m[1039]));
    m[710] = (((m[258]&~m[454]&m[1074])|(~m[258]&m[454]&m[1074]))&BiasedRNG[421])|(((m[258]&m[454]&~m[1074]))&~BiasedRNG[421])|((m[258]&m[454]&m[1074]));
    m[711] = (((m[274]&~m[455]&m[1114])|(~m[274]&m[455]&m[1114]))&BiasedRNG[422])|(((m[274]&m[455]&~m[1114]))&~BiasedRNG[422])|((m[274]&m[455]&m[1114]));
    m[712] = (((m[290]&~m[456]&m[1159])|(~m[290]&m[456]&m[1159]))&BiasedRNG[423])|(((m[290]&m[456]&~m[1159]))&~BiasedRNG[423])|((m[290]&m[456]&m[1159]));
    m[713] = (((m[306]&~m[457]&m[1209])|(~m[306]&m[457]&m[1209]))&BiasedRNG[424])|(((m[306]&m[457]&~m[1209]))&~BiasedRNG[424])|((m[306]&m[457]&m[1209]));
    m[714] = (((m[322]&~m[458]&m[1264])|(~m[322]&m[458]&m[1264]))&BiasedRNG[425])|(((m[322]&m[458]&~m[1264]))&~BiasedRNG[425])|((m[322]&m[458]&m[1264]));
    m[715] = (((m[338]&~m[459]&m[1324])|(~m[338]&m[459]&m[1324]))&BiasedRNG[426])|(((m[338]&m[459]&~m[1324]))&~BiasedRNG[426])|((m[338]&m[459]&m[1324]));
    m[716] = (((m[354]&~m[460]&m[1389])|(~m[354]&m[460]&m[1389]))&BiasedRNG[427])|(((m[354]&m[460]&~m[1389]))&~BiasedRNG[427])|((m[354]&m[460]&m[1389]));
    m[717] = (((m[370]&~m[461]&m[1459])|(~m[370]&m[461]&m[1459]))&BiasedRNG[428])|(((m[370]&m[461]&~m[1459]))&~BiasedRNG[428])|((m[370]&m[461]&m[1459]));
    m[718] = (((m[386]&~m[462]&m[1534])|(~m[386]&m[462]&m[1534]))&BiasedRNG[429])|(((m[386]&m[462]&~m[1534]))&~BiasedRNG[429])|((m[386]&m[462]&m[1534]));
    m[719] = (((m[402]&~m[463]&m[1604])|(~m[402]&m[463]&m[1604]))&BiasedRNG[430])|(((m[402]&m[463]&~m[1604]))&~BiasedRNG[430])|((m[402]&m[463]&m[1604]));
    m[720] = (((m[163]&~m[464]&m[954])|(~m[163]&m[464]&m[954]))&BiasedRNG[431])|(((m[163]&m[464]&~m[954]))&~BiasedRNG[431])|((m[163]&m[464]&m[954]));
    m[721] = (((m[179]&~m[465]&m[969])|(~m[179]&m[465]&m[969]))&BiasedRNG[432])|(((m[179]&m[465]&~m[969]))&~BiasedRNG[432])|((m[179]&m[465]&m[969]));
    m[722] = (((m[195]&~m[466]&m[989])|(~m[195]&m[466]&m[989]))&BiasedRNG[433])|(((m[195]&m[466]&~m[989]))&~BiasedRNG[433])|((m[195]&m[466]&m[989]));
    m[723] = (((m[211]&~m[467]&m[1014])|(~m[211]&m[467]&m[1014]))&BiasedRNG[434])|(((m[211]&m[467]&~m[1014]))&~BiasedRNG[434])|((m[211]&m[467]&m[1014]));
    m[724] = (((m[227]&~m[468]&m[1044])|(~m[227]&m[468]&m[1044]))&BiasedRNG[435])|(((m[227]&m[468]&~m[1044]))&~BiasedRNG[435])|((m[227]&m[468]&m[1044]));
    m[725] = (((m[243]&~m[469]&m[1079])|(~m[243]&m[469]&m[1079]))&BiasedRNG[436])|(((m[243]&m[469]&~m[1079]))&~BiasedRNG[436])|((m[243]&m[469]&m[1079]));
    m[726] = (((m[259]&~m[470]&m[1119])|(~m[259]&m[470]&m[1119]))&BiasedRNG[437])|(((m[259]&m[470]&~m[1119]))&~BiasedRNG[437])|((m[259]&m[470]&m[1119]));
    m[727] = (((m[275]&~m[471]&m[1164])|(~m[275]&m[471]&m[1164]))&BiasedRNG[438])|(((m[275]&m[471]&~m[1164]))&~BiasedRNG[438])|((m[275]&m[471]&m[1164]));
    m[728] = (((m[291]&~m[472]&m[1214])|(~m[291]&m[472]&m[1214]))&BiasedRNG[439])|(((m[291]&m[472]&~m[1214]))&~BiasedRNG[439])|((m[291]&m[472]&m[1214]));
    m[729] = (((m[307]&~m[473]&m[1269])|(~m[307]&m[473]&m[1269]))&BiasedRNG[440])|(((m[307]&m[473]&~m[1269]))&~BiasedRNG[440])|((m[307]&m[473]&m[1269]));
    m[730] = (((m[323]&~m[474]&m[1329])|(~m[323]&m[474]&m[1329]))&BiasedRNG[441])|(((m[323]&m[474]&~m[1329]))&~BiasedRNG[441])|((m[323]&m[474]&m[1329]));
    m[731] = (((m[339]&~m[475]&m[1394])|(~m[339]&m[475]&m[1394]))&BiasedRNG[442])|(((m[339]&m[475]&~m[1394]))&~BiasedRNG[442])|((m[339]&m[475]&m[1394]));
    m[732] = (((m[355]&~m[476]&m[1464])|(~m[355]&m[476]&m[1464]))&BiasedRNG[443])|(((m[355]&m[476]&~m[1464]))&~BiasedRNG[443])|((m[355]&m[476]&m[1464]));
    m[733] = (((m[371]&~m[477]&m[1539])|(~m[371]&m[477]&m[1539]))&BiasedRNG[444])|(((m[371]&m[477]&~m[1539]))&~BiasedRNG[444])|((m[371]&m[477]&m[1539]));
    m[734] = (((m[387]&~m[478]&m[1609])|(~m[387]&m[478]&m[1609]))&BiasedRNG[445])|(((m[387]&m[478]&~m[1609]))&~BiasedRNG[445])|((m[387]&m[478]&m[1609]));
    m[735] = (((m[403]&~m[479]&m[1674])|(~m[403]&m[479]&m[1674]))&BiasedRNG[446])|(((m[403]&m[479]&~m[1674]))&~BiasedRNG[446])|((m[403]&m[479]&m[1674]));
    m[736] = (((m[164]&~m[480]&m[974])|(~m[164]&m[480]&m[974]))&BiasedRNG[447])|(((m[164]&m[480]&~m[974]))&~BiasedRNG[447])|((m[164]&m[480]&m[974]));
    m[737] = (((m[180]&~m[481]&m[994])|(~m[180]&m[481]&m[994]))&BiasedRNG[448])|(((m[180]&m[481]&~m[994]))&~BiasedRNG[448])|((m[180]&m[481]&m[994]));
    m[738] = (((m[196]&~m[482]&m[1019])|(~m[196]&m[482]&m[1019]))&BiasedRNG[449])|(((m[196]&m[482]&~m[1019]))&~BiasedRNG[449])|((m[196]&m[482]&m[1019]));
    m[739] = (((m[212]&~m[483]&m[1049])|(~m[212]&m[483]&m[1049]))&BiasedRNG[450])|(((m[212]&m[483]&~m[1049]))&~BiasedRNG[450])|((m[212]&m[483]&m[1049]));
    m[740] = (((m[228]&~m[484]&m[1084])|(~m[228]&m[484]&m[1084]))&BiasedRNG[451])|(((m[228]&m[484]&~m[1084]))&~BiasedRNG[451])|((m[228]&m[484]&m[1084]));
    m[741] = (((m[244]&~m[485]&m[1124])|(~m[244]&m[485]&m[1124]))&BiasedRNG[452])|(((m[244]&m[485]&~m[1124]))&~BiasedRNG[452])|((m[244]&m[485]&m[1124]));
    m[742] = (((m[260]&~m[486]&m[1169])|(~m[260]&m[486]&m[1169]))&BiasedRNG[453])|(((m[260]&m[486]&~m[1169]))&~BiasedRNG[453])|((m[260]&m[486]&m[1169]));
    m[743] = (((m[276]&~m[487]&m[1219])|(~m[276]&m[487]&m[1219]))&BiasedRNG[454])|(((m[276]&m[487]&~m[1219]))&~BiasedRNG[454])|((m[276]&m[487]&m[1219]));
    m[744] = (((m[292]&~m[488]&m[1274])|(~m[292]&m[488]&m[1274]))&BiasedRNG[455])|(((m[292]&m[488]&~m[1274]))&~BiasedRNG[455])|((m[292]&m[488]&m[1274]));
    m[745] = (((m[308]&~m[489]&m[1334])|(~m[308]&m[489]&m[1334]))&BiasedRNG[456])|(((m[308]&m[489]&~m[1334]))&~BiasedRNG[456])|((m[308]&m[489]&m[1334]));
    m[746] = (((m[324]&~m[490]&m[1399])|(~m[324]&m[490]&m[1399]))&BiasedRNG[457])|(((m[324]&m[490]&~m[1399]))&~BiasedRNG[457])|((m[324]&m[490]&m[1399]));
    m[747] = (((m[340]&~m[491]&m[1469])|(~m[340]&m[491]&m[1469]))&BiasedRNG[458])|(((m[340]&m[491]&~m[1469]))&~BiasedRNG[458])|((m[340]&m[491]&m[1469]));
    m[748] = (((m[356]&~m[492]&m[1544])|(~m[356]&m[492]&m[1544]))&BiasedRNG[459])|(((m[356]&m[492]&~m[1544]))&~BiasedRNG[459])|((m[356]&m[492]&m[1544]));
    m[749] = (((m[372]&~m[493]&m[1614])|(~m[372]&m[493]&m[1614]))&BiasedRNG[460])|(((m[372]&m[493]&~m[1614]))&~BiasedRNG[460])|((m[372]&m[493]&m[1614]));
    m[750] = (((m[388]&~m[494]&m[1679])|(~m[388]&m[494]&m[1679]))&BiasedRNG[461])|(((m[388]&m[494]&~m[1679]))&~BiasedRNG[461])|((m[388]&m[494]&m[1679]));
    m[751] = (((m[404]&~m[495]&m[1739])|(~m[404]&m[495]&m[1739]))&BiasedRNG[462])|(((m[404]&m[495]&~m[1739]))&~BiasedRNG[462])|((m[404]&m[495]&m[1739]));
    m[752] = (((m[165]&~m[496]&m[999])|(~m[165]&m[496]&m[999]))&BiasedRNG[463])|(((m[165]&m[496]&~m[999]))&~BiasedRNG[463])|((m[165]&m[496]&m[999]));
    m[753] = (((m[181]&~m[497]&m[1024])|(~m[181]&m[497]&m[1024]))&BiasedRNG[464])|(((m[181]&m[497]&~m[1024]))&~BiasedRNG[464])|((m[181]&m[497]&m[1024]));
    m[754] = (((m[197]&~m[498]&m[1054])|(~m[197]&m[498]&m[1054]))&BiasedRNG[465])|(((m[197]&m[498]&~m[1054]))&~BiasedRNG[465])|((m[197]&m[498]&m[1054]));
    m[755] = (((m[213]&~m[499]&m[1089])|(~m[213]&m[499]&m[1089]))&BiasedRNG[466])|(((m[213]&m[499]&~m[1089]))&~BiasedRNG[466])|((m[213]&m[499]&m[1089]));
    m[756] = (((m[229]&~m[500]&m[1129])|(~m[229]&m[500]&m[1129]))&BiasedRNG[467])|(((m[229]&m[500]&~m[1129]))&~BiasedRNG[467])|((m[229]&m[500]&m[1129]));
    m[757] = (((m[245]&~m[501]&m[1174])|(~m[245]&m[501]&m[1174]))&BiasedRNG[468])|(((m[245]&m[501]&~m[1174]))&~BiasedRNG[468])|((m[245]&m[501]&m[1174]));
    m[758] = (((m[261]&~m[502]&m[1224])|(~m[261]&m[502]&m[1224]))&BiasedRNG[469])|(((m[261]&m[502]&~m[1224]))&~BiasedRNG[469])|((m[261]&m[502]&m[1224]));
    m[759] = (((m[277]&~m[503]&m[1279])|(~m[277]&m[503]&m[1279]))&BiasedRNG[470])|(((m[277]&m[503]&~m[1279]))&~BiasedRNG[470])|((m[277]&m[503]&m[1279]));
    m[760] = (((m[293]&~m[504]&m[1339])|(~m[293]&m[504]&m[1339]))&BiasedRNG[471])|(((m[293]&m[504]&~m[1339]))&~BiasedRNG[471])|((m[293]&m[504]&m[1339]));
    m[761] = (((m[309]&~m[505]&m[1404])|(~m[309]&m[505]&m[1404]))&BiasedRNG[472])|(((m[309]&m[505]&~m[1404]))&~BiasedRNG[472])|((m[309]&m[505]&m[1404]));
    m[762] = (((m[325]&~m[506]&m[1474])|(~m[325]&m[506]&m[1474]))&BiasedRNG[473])|(((m[325]&m[506]&~m[1474]))&~BiasedRNG[473])|((m[325]&m[506]&m[1474]));
    m[763] = (((m[341]&~m[507]&m[1549])|(~m[341]&m[507]&m[1549]))&BiasedRNG[474])|(((m[341]&m[507]&~m[1549]))&~BiasedRNG[474])|((m[341]&m[507]&m[1549]));
    m[764] = (((m[357]&~m[508]&m[1619])|(~m[357]&m[508]&m[1619]))&BiasedRNG[475])|(((m[357]&m[508]&~m[1619]))&~BiasedRNG[475])|((m[357]&m[508]&m[1619]));
    m[765] = (((m[373]&~m[509]&m[1684])|(~m[373]&m[509]&m[1684]))&BiasedRNG[476])|(((m[373]&m[509]&~m[1684]))&~BiasedRNG[476])|((m[373]&m[509]&m[1684]));
    m[766] = (((m[389]&~m[510]&m[1744])|(~m[389]&m[510]&m[1744]))&BiasedRNG[477])|(((m[389]&m[510]&~m[1744]))&~BiasedRNG[477])|((m[389]&m[510]&m[1744]));
    m[767] = (((m[405]&~m[511]&m[1799])|(~m[405]&m[511]&m[1799]))&BiasedRNG[478])|(((m[405]&m[511]&~m[1799]))&~BiasedRNG[478])|((m[405]&m[511]&m[1799]));
    m[768] = (((m[166]&~m[512]&m[1029])|(~m[166]&m[512]&m[1029]))&BiasedRNG[479])|(((m[166]&m[512]&~m[1029]))&~BiasedRNG[479])|((m[166]&m[512]&m[1029]));
    m[769] = (((m[182]&~m[513]&m[1059])|(~m[182]&m[513]&m[1059]))&BiasedRNG[480])|(((m[182]&m[513]&~m[1059]))&~BiasedRNG[480])|((m[182]&m[513]&m[1059]));
    m[770] = (((m[198]&~m[514]&m[1094])|(~m[198]&m[514]&m[1094]))&BiasedRNG[481])|(((m[198]&m[514]&~m[1094]))&~BiasedRNG[481])|((m[198]&m[514]&m[1094]));
    m[771] = (((m[214]&~m[515]&m[1134])|(~m[214]&m[515]&m[1134]))&BiasedRNG[482])|(((m[214]&m[515]&~m[1134]))&~BiasedRNG[482])|((m[214]&m[515]&m[1134]));
    m[772] = (((m[230]&~m[516]&m[1179])|(~m[230]&m[516]&m[1179]))&BiasedRNG[483])|(((m[230]&m[516]&~m[1179]))&~BiasedRNG[483])|((m[230]&m[516]&m[1179]));
    m[773] = (((m[246]&~m[517]&m[1229])|(~m[246]&m[517]&m[1229]))&BiasedRNG[484])|(((m[246]&m[517]&~m[1229]))&~BiasedRNG[484])|((m[246]&m[517]&m[1229]));
    m[774] = (((m[262]&~m[518]&m[1284])|(~m[262]&m[518]&m[1284]))&BiasedRNG[485])|(((m[262]&m[518]&~m[1284]))&~BiasedRNG[485])|((m[262]&m[518]&m[1284]));
    m[775] = (((m[278]&~m[519]&m[1344])|(~m[278]&m[519]&m[1344]))&BiasedRNG[486])|(((m[278]&m[519]&~m[1344]))&~BiasedRNG[486])|((m[278]&m[519]&m[1344]));
    m[776] = (((m[294]&~m[520]&m[1409])|(~m[294]&m[520]&m[1409]))&BiasedRNG[487])|(((m[294]&m[520]&~m[1409]))&~BiasedRNG[487])|((m[294]&m[520]&m[1409]));
    m[777] = (((m[310]&~m[521]&m[1479])|(~m[310]&m[521]&m[1479]))&BiasedRNG[488])|(((m[310]&m[521]&~m[1479]))&~BiasedRNG[488])|((m[310]&m[521]&m[1479]));
    m[778] = (((m[326]&~m[522]&m[1554])|(~m[326]&m[522]&m[1554]))&BiasedRNG[489])|(((m[326]&m[522]&~m[1554]))&~BiasedRNG[489])|((m[326]&m[522]&m[1554]));
    m[779] = (((m[342]&~m[523]&m[1624])|(~m[342]&m[523]&m[1624]))&BiasedRNG[490])|(((m[342]&m[523]&~m[1624]))&~BiasedRNG[490])|((m[342]&m[523]&m[1624]));
    m[780] = (((m[358]&~m[524]&m[1689])|(~m[358]&m[524]&m[1689]))&BiasedRNG[491])|(((m[358]&m[524]&~m[1689]))&~BiasedRNG[491])|((m[358]&m[524]&m[1689]));
    m[781] = (((m[374]&~m[525]&m[1749])|(~m[374]&m[525]&m[1749]))&BiasedRNG[492])|(((m[374]&m[525]&~m[1749]))&~BiasedRNG[492])|((m[374]&m[525]&m[1749]));
    m[782] = (((m[390]&~m[526]&m[1804])|(~m[390]&m[526]&m[1804]))&BiasedRNG[493])|(((m[390]&m[526]&~m[1804]))&~BiasedRNG[493])|((m[390]&m[526]&m[1804]));
    m[783] = (((m[406]&~m[527]&m[1854])|(~m[406]&m[527]&m[1854]))&BiasedRNG[494])|(((m[406]&m[527]&~m[1854]))&~BiasedRNG[494])|((m[406]&m[527]&m[1854]));
    m[784] = (((m[167]&~m[528]&m[1064])|(~m[167]&m[528]&m[1064]))&BiasedRNG[495])|(((m[167]&m[528]&~m[1064]))&~BiasedRNG[495])|((m[167]&m[528]&m[1064]));
    m[785] = (((m[183]&~m[529]&m[1099])|(~m[183]&m[529]&m[1099]))&BiasedRNG[496])|(((m[183]&m[529]&~m[1099]))&~BiasedRNG[496])|((m[183]&m[529]&m[1099]));
    m[786] = (((m[199]&~m[530]&m[1139])|(~m[199]&m[530]&m[1139]))&BiasedRNG[497])|(((m[199]&m[530]&~m[1139]))&~BiasedRNG[497])|((m[199]&m[530]&m[1139]));
    m[787] = (((m[215]&~m[531]&m[1184])|(~m[215]&m[531]&m[1184]))&BiasedRNG[498])|(((m[215]&m[531]&~m[1184]))&~BiasedRNG[498])|((m[215]&m[531]&m[1184]));
    m[788] = (((m[231]&~m[532]&m[1234])|(~m[231]&m[532]&m[1234]))&BiasedRNG[499])|(((m[231]&m[532]&~m[1234]))&~BiasedRNG[499])|((m[231]&m[532]&m[1234]));
    m[789] = (((m[247]&~m[533]&m[1289])|(~m[247]&m[533]&m[1289]))&BiasedRNG[500])|(((m[247]&m[533]&~m[1289]))&~BiasedRNG[500])|((m[247]&m[533]&m[1289]));
    m[790] = (((m[263]&~m[534]&m[1349])|(~m[263]&m[534]&m[1349]))&BiasedRNG[501])|(((m[263]&m[534]&~m[1349]))&~BiasedRNG[501])|((m[263]&m[534]&m[1349]));
    m[791] = (((m[279]&~m[535]&m[1414])|(~m[279]&m[535]&m[1414]))&BiasedRNG[502])|(((m[279]&m[535]&~m[1414]))&~BiasedRNG[502])|((m[279]&m[535]&m[1414]));
    m[792] = (((m[295]&~m[536]&m[1484])|(~m[295]&m[536]&m[1484]))&BiasedRNG[503])|(((m[295]&m[536]&~m[1484]))&~BiasedRNG[503])|((m[295]&m[536]&m[1484]));
    m[793] = (((m[311]&~m[537]&m[1559])|(~m[311]&m[537]&m[1559]))&BiasedRNG[504])|(((m[311]&m[537]&~m[1559]))&~BiasedRNG[504])|((m[311]&m[537]&m[1559]));
    m[794] = (((m[327]&~m[538]&m[1629])|(~m[327]&m[538]&m[1629]))&BiasedRNG[505])|(((m[327]&m[538]&~m[1629]))&~BiasedRNG[505])|((m[327]&m[538]&m[1629]));
    m[795] = (((m[343]&~m[539]&m[1694])|(~m[343]&m[539]&m[1694]))&BiasedRNG[506])|(((m[343]&m[539]&~m[1694]))&~BiasedRNG[506])|((m[343]&m[539]&m[1694]));
    m[796] = (((m[359]&~m[540]&m[1754])|(~m[359]&m[540]&m[1754]))&BiasedRNG[507])|(((m[359]&m[540]&~m[1754]))&~BiasedRNG[507])|((m[359]&m[540]&m[1754]));
    m[797] = (((m[375]&~m[541]&m[1809])|(~m[375]&m[541]&m[1809]))&BiasedRNG[508])|(((m[375]&m[541]&~m[1809]))&~BiasedRNG[508])|((m[375]&m[541]&m[1809]));
    m[798] = (((m[391]&~m[542]&m[1859])|(~m[391]&m[542]&m[1859]))&BiasedRNG[509])|(((m[391]&m[542]&~m[1859]))&~BiasedRNG[509])|((m[391]&m[542]&m[1859]));
    m[799] = (((m[407]&~m[543]&m[1904])|(~m[407]&m[543]&m[1904]))&BiasedRNG[510])|(((m[407]&m[543]&~m[1904]))&~BiasedRNG[510])|((m[407]&m[543]&m[1904]));
    m[800] = (((m[168]&~m[544]&m[1104])|(~m[168]&m[544]&m[1104]))&BiasedRNG[511])|(((m[168]&m[544]&~m[1104]))&~BiasedRNG[511])|((m[168]&m[544]&m[1104]));
    m[801] = (((m[184]&~m[545]&m[1144])|(~m[184]&m[545]&m[1144]))&BiasedRNG[512])|(((m[184]&m[545]&~m[1144]))&~BiasedRNG[512])|((m[184]&m[545]&m[1144]));
    m[802] = (((m[200]&~m[546]&m[1189])|(~m[200]&m[546]&m[1189]))&BiasedRNG[513])|(((m[200]&m[546]&~m[1189]))&~BiasedRNG[513])|((m[200]&m[546]&m[1189]));
    m[803] = (((m[216]&~m[547]&m[1239])|(~m[216]&m[547]&m[1239]))&BiasedRNG[514])|(((m[216]&m[547]&~m[1239]))&~BiasedRNG[514])|((m[216]&m[547]&m[1239]));
    m[804] = (((m[232]&~m[548]&m[1294])|(~m[232]&m[548]&m[1294]))&BiasedRNG[515])|(((m[232]&m[548]&~m[1294]))&~BiasedRNG[515])|((m[232]&m[548]&m[1294]));
    m[805] = (((m[248]&~m[549]&m[1354])|(~m[248]&m[549]&m[1354]))&BiasedRNG[516])|(((m[248]&m[549]&~m[1354]))&~BiasedRNG[516])|((m[248]&m[549]&m[1354]));
    m[806] = (((m[264]&~m[550]&m[1419])|(~m[264]&m[550]&m[1419]))&BiasedRNG[517])|(((m[264]&m[550]&~m[1419]))&~BiasedRNG[517])|((m[264]&m[550]&m[1419]));
    m[807] = (((m[280]&~m[551]&m[1489])|(~m[280]&m[551]&m[1489]))&BiasedRNG[518])|(((m[280]&m[551]&~m[1489]))&~BiasedRNG[518])|((m[280]&m[551]&m[1489]));
    m[808] = (((m[296]&~m[552]&m[1564])|(~m[296]&m[552]&m[1564]))&BiasedRNG[519])|(((m[296]&m[552]&~m[1564]))&~BiasedRNG[519])|((m[296]&m[552]&m[1564]));
    m[809] = (((m[312]&~m[553]&m[1634])|(~m[312]&m[553]&m[1634]))&BiasedRNG[520])|(((m[312]&m[553]&~m[1634]))&~BiasedRNG[520])|((m[312]&m[553]&m[1634]));
    m[810] = (((m[328]&~m[554]&m[1699])|(~m[328]&m[554]&m[1699]))&BiasedRNG[521])|(((m[328]&m[554]&~m[1699]))&~BiasedRNG[521])|((m[328]&m[554]&m[1699]));
    m[811] = (((m[344]&~m[555]&m[1759])|(~m[344]&m[555]&m[1759]))&BiasedRNG[522])|(((m[344]&m[555]&~m[1759]))&~BiasedRNG[522])|((m[344]&m[555]&m[1759]));
    m[812] = (((m[360]&~m[556]&m[1814])|(~m[360]&m[556]&m[1814]))&BiasedRNG[523])|(((m[360]&m[556]&~m[1814]))&~BiasedRNG[523])|((m[360]&m[556]&m[1814]));
    m[813] = (((m[376]&~m[557]&m[1864])|(~m[376]&m[557]&m[1864]))&BiasedRNG[524])|(((m[376]&m[557]&~m[1864]))&~BiasedRNG[524])|((m[376]&m[557]&m[1864]));
    m[814] = (((m[392]&~m[558]&m[1909])|(~m[392]&m[558]&m[1909]))&BiasedRNG[525])|(((m[392]&m[558]&~m[1909]))&~BiasedRNG[525])|((m[392]&m[558]&m[1909]));
    m[815] = (((m[408]&~m[559]&m[1949])|(~m[408]&m[559]&m[1949]))&BiasedRNG[526])|(((m[408]&m[559]&~m[1949]))&~BiasedRNG[526])|((m[408]&m[559]&m[1949]));
    m[816] = (((m[169]&~m[560]&m[1149])|(~m[169]&m[560]&m[1149]))&BiasedRNG[527])|(((m[169]&m[560]&~m[1149]))&~BiasedRNG[527])|((m[169]&m[560]&m[1149]));
    m[817] = (((m[185]&~m[561]&m[1194])|(~m[185]&m[561]&m[1194]))&BiasedRNG[528])|(((m[185]&m[561]&~m[1194]))&~BiasedRNG[528])|((m[185]&m[561]&m[1194]));
    m[818] = (((m[201]&~m[562]&m[1244])|(~m[201]&m[562]&m[1244]))&BiasedRNG[529])|(((m[201]&m[562]&~m[1244]))&~BiasedRNG[529])|((m[201]&m[562]&m[1244]));
    m[819] = (((m[217]&~m[563]&m[1299])|(~m[217]&m[563]&m[1299]))&BiasedRNG[530])|(((m[217]&m[563]&~m[1299]))&~BiasedRNG[530])|((m[217]&m[563]&m[1299]));
    m[820] = (((m[233]&~m[564]&m[1359])|(~m[233]&m[564]&m[1359]))&BiasedRNG[531])|(((m[233]&m[564]&~m[1359]))&~BiasedRNG[531])|((m[233]&m[564]&m[1359]));
    m[821] = (((m[249]&~m[565]&m[1424])|(~m[249]&m[565]&m[1424]))&BiasedRNG[532])|(((m[249]&m[565]&~m[1424]))&~BiasedRNG[532])|((m[249]&m[565]&m[1424]));
    m[822] = (((m[265]&~m[566]&m[1494])|(~m[265]&m[566]&m[1494]))&BiasedRNG[533])|(((m[265]&m[566]&~m[1494]))&~BiasedRNG[533])|((m[265]&m[566]&m[1494]));
    m[823] = (((m[281]&~m[567]&m[1569])|(~m[281]&m[567]&m[1569]))&BiasedRNG[534])|(((m[281]&m[567]&~m[1569]))&~BiasedRNG[534])|((m[281]&m[567]&m[1569]));
    m[824] = (((m[297]&~m[568]&m[1639])|(~m[297]&m[568]&m[1639]))&BiasedRNG[535])|(((m[297]&m[568]&~m[1639]))&~BiasedRNG[535])|((m[297]&m[568]&m[1639]));
    m[825] = (((m[313]&~m[569]&m[1704])|(~m[313]&m[569]&m[1704]))&BiasedRNG[536])|(((m[313]&m[569]&~m[1704]))&~BiasedRNG[536])|((m[313]&m[569]&m[1704]));
    m[826] = (((m[329]&~m[570]&m[1764])|(~m[329]&m[570]&m[1764]))&BiasedRNG[537])|(((m[329]&m[570]&~m[1764]))&~BiasedRNG[537])|((m[329]&m[570]&m[1764]));
    m[827] = (((m[345]&~m[571]&m[1819])|(~m[345]&m[571]&m[1819]))&BiasedRNG[538])|(((m[345]&m[571]&~m[1819]))&~BiasedRNG[538])|((m[345]&m[571]&m[1819]));
    m[828] = (((m[361]&~m[572]&m[1869])|(~m[361]&m[572]&m[1869]))&BiasedRNG[539])|(((m[361]&m[572]&~m[1869]))&~BiasedRNG[539])|((m[361]&m[572]&m[1869]));
    m[829] = (((m[377]&~m[573]&m[1914])|(~m[377]&m[573]&m[1914]))&BiasedRNG[540])|(((m[377]&m[573]&~m[1914]))&~BiasedRNG[540])|((m[377]&m[573]&m[1914]));
    m[830] = (((m[393]&~m[574]&m[1954])|(~m[393]&m[574]&m[1954]))&BiasedRNG[541])|(((m[393]&m[574]&~m[1954]))&~BiasedRNG[541])|((m[393]&m[574]&m[1954]));
    m[831] = (((m[409]&~m[575]&m[1989])|(~m[409]&m[575]&m[1989]))&BiasedRNG[542])|(((m[409]&m[575]&~m[1989]))&~BiasedRNG[542])|((m[409]&m[575]&m[1989]));
    m[832] = (((m[170]&~m[576]&m[1199])|(~m[170]&m[576]&m[1199]))&BiasedRNG[543])|(((m[170]&m[576]&~m[1199]))&~BiasedRNG[543])|((m[170]&m[576]&m[1199]));
    m[833] = (((m[186]&~m[577]&m[1249])|(~m[186]&m[577]&m[1249]))&BiasedRNG[544])|(((m[186]&m[577]&~m[1249]))&~BiasedRNG[544])|((m[186]&m[577]&m[1249]));
    m[834] = (((m[202]&~m[578]&m[1304])|(~m[202]&m[578]&m[1304]))&BiasedRNG[545])|(((m[202]&m[578]&~m[1304]))&~BiasedRNG[545])|((m[202]&m[578]&m[1304]));
    m[835] = (((m[218]&~m[579]&m[1364])|(~m[218]&m[579]&m[1364]))&BiasedRNG[546])|(((m[218]&m[579]&~m[1364]))&~BiasedRNG[546])|((m[218]&m[579]&m[1364]));
    m[836] = (((m[234]&~m[580]&m[1429])|(~m[234]&m[580]&m[1429]))&BiasedRNG[547])|(((m[234]&m[580]&~m[1429]))&~BiasedRNG[547])|((m[234]&m[580]&m[1429]));
    m[837] = (((m[250]&~m[581]&m[1499])|(~m[250]&m[581]&m[1499]))&BiasedRNG[548])|(((m[250]&m[581]&~m[1499]))&~BiasedRNG[548])|((m[250]&m[581]&m[1499]));
    m[838] = (((m[266]&~m[582]&m[1574])|(~m[266]&m[582]&m[1574]))&BiasedRNG[549])|(((m[266]&m[582]&~m[1574]))&~BiasedRNG[549])|((m[266]&m[582]&m[1574]));
    m[839] = (((m[282]&~m[583]&m[1644])|(~m[282]&m[583]&m[1644]))&BiasedRNG[550])|(((m[282]&m[583]&~m[1644]))&~BiasedRNG[550])|((m[282]&m[583]&m[1644]));
    m[840] = (((m[298]&~m[584]&m[1709])|(~m[298]&m[584]&m[1709]))&BiasedRNG[551])|(((m[298]&m[584]&~m[1709]))&~BiasedRNG[551])|((m[298]&m[584]&m[1709]));
    m[841] = (((m[314]&~m[585]&m[1769])|(~m[314]&m[585]&m[1769]))&BiasedRNG[552])|(((m[314]&m[585]&~m[1769]))&~BiasedRNG[552])|((m[314]&m[585]&m[1769]));
    m[842] = (((m[330]&~m[586]&m[1824])|(~m[330]&m[586]&m[1824]))&BiasedRNG[553])|(((m[330]&m[586]&~m[1824]))&~BiasedRNG[553])|((m[330]&m[586]&m[1824]));
    m[843] = (((m[346]&~m[587]&m[1874])|(~m[346]&m[587]&m[1874]))&BiasedRNG[554])|(((m[346]&m[587]&~m[1874]))&~BiasedRNG[554])|((m[346]&m[587]&m[1874]));
    m[844] = (((m[362]&~m[588]&m[1919])|(~m[362]&m[588]&m[1919]))&BiasedRNG[555])|(((m[362]&m[588]&~m[1919]))&~BiasedRNG[555])|((m[362]&m[588]&m[1919]));
    m[845] = (((m[378]&~m[589]&m[1959])|(~m[378]&m[589]&m[1959]))&BiasedRNG[556])|(((m[378]&m[589]&~m[1959]))&~BiasedRNG[556])|((m[378]&m[589]&m[1959]));
    m[846] = (((m[394]&~m[590]&m[1994])|(~m[394]&m[590]&m[1994]))&BiasedRNG[557])|(((m[394]&m[590]&~m[1994]))&~BiasedRNG[557])|((m[394]&m[590]&m[1994]));
    m[847] = (((m[410]&~m[591]&m[2024])|(~m[410]&m[591]&m[2024]))&BiasedRNG[558])|(((m[410]&m[591]&~m[2024]))&~BiasedRNG[558])|((m[410]&m[591]&m[2024]));
    m[848] = (((m[171]&~m[592]&m[1254])|(~m[171]&m[592]&m[1254]))&BiasedRNG[559])|(((m[171]&m[592]&~m[1254]))&~BiasedRNG[559])|((m[171]&m[592]&m[1254]));
    m[849] = (((m[187]&~m[593]&m[1309])|(~m[187]&m[593]&m[1309]))&BiasedRNG[560])|(((m[187]&m[593]&~m[1309]))&~BiasedRNG[560])|((m[187]&m[593]&m[1309]));
    m[850] = (((m[203]&~m[594]&m[1369])|(~m[203]&m[594]&m[1369]))&BiasedRNG[561])|(((m[203]&m[594]&~m[1369]))&~BiasedRNG[561])|((m[203]&m[594]&m[1369]));
    m[851] = (((m[219]&~m[595]&m[1434])|(~m[219]&m[595]&m[1434]))&BiasedRNG[562])|(((m[219]&m[595]&~m[1434]))&~BiasedRNG[562])|((m[219]&m[595]&m[1434]));
    m[852] = (((m[235]&~m[596]&m[1504])|(~m[235]&m[596]&m[1504]))&BiasedRNG[563])|(((m[235]&m[596]&~m[1504]))&~BiasedRNG[563])|((m[235]&m[596]&m[1504]));
    m[853] = (((m[251]&~m[597]&m[1579])|(~m[251]&m[597]&m[1579]))&BiasedRNG[564])|(((m[251]&m[597]&~m[1579]))&~BiasedRNG[564])|((m[251]&m[597]&m[1579]));
    m[854] = (((m[267]&~m[598]&m[1649])|(~m[267]&m[598]&m[1649]))&BiasedRNG[565])|(((m[267]&m[598]&~m[1649]))&~BiasedRNG[565])|((m[267]&m[598]&m[1649]));
    m[855] = (((m[283]&~m[599]&m[1714])|(~m[283]&m[599]&m[1714]))&BiasedRNG[566])|(((m[283]&m[599]&~m[1714]))&~BiasedRNG[566])|((m[283]&m[599]&m[1714]));
    m[856] = (((m[299]&~m[600]&m[1774])|(~m[299]&m[600]&m[1774]))&BiasedRNG[567])|(((m[299]&m[600]&~m[1774]))&~BiasedRNG[567])|((m[299]&m[600]&m[1774]));
    m[857] = (((m[315]&~m[601]&m[1829])|(~m[315]&m[601]&m[1829]))&BiasedRNG[568])|(((m[315]&m[601]&~m[1829]))&~BiasedRNG[568])|((m[315]&m[601]&m[1829]));
    m[858] = (((m[331]&~m[602]&m[1879])|(~m[331]&m[602]&m[1879]))&BiasedRNG[569])|(((m[331]&m[602]&~m[1879]))&~BiasedRNG[569])|((m[331]&m[602]&m[1879]));
    m[859] = (((m[347]&~m[603]&m[1924])|(~m[347]&m[603]&m[1924]))&BiasedRNG[570])|(((m[347]&m[603]&~m[1924]))&~BiasedRNG[570])|((m[347]&m[603]&m[1924]));
    m[860] = (((m[363]&~m[604]&m[1964])|(~m[363]&m[604]&m[1964]))&BiasedRNG[571])|(((m[363]&m[604]&~m[1964]))&~BiasedRNG[571])|((m[363]&m[604]&m[1964]));
    m[861] = (((m[379]&~m[605]&m[1999])|(~m[379]&m[605]&m[1999]))&BiasedRNG[572])|(((m[379]&m[605]&~m[1999]))&~BiasedRNG[572])|((m[379]&m[605]&m[1999]));
    m[862] = (((m[395]&~m[606]&m[2029])|(~m[395]&m[606]&m[2029]))&BiasedRNG[573])|(((m[395]&m[606]&~m[2029]))&~BiasedRNG[573])|((m[395]&m[606]&m[2029]));
    m[863] = (((m[411]&~m[607]&m[2054])|(~m[411]&m[607]&m[2054]))&BiasedRNG[574])|(((m[411]&m[607]&~m[2054]))&~BiasedRNG[574])|((m[411]&m[607]&m[2054]));
    m[864] = (((m[172]&~m[608]&m[1314])|(~m[172]&m[608]&m[1314]))&BiasedRNG[575])|(((m[172]&m[608]&~m[1314]))&~BiasedRNG[575])|((m[172]&m[608]&m[1314]));
    m[865] = (((m[188]&~m[609]&m[1374])|(~m[188]&m[609]&m[1374]))&BiasedRNG[576])|(((m[188]&m[609]&~m[1374]))&~BiasedRNG[576])|((m[188]&m[609]&m[1374]));
    m[866] = (((m[204]&~m[610]&m[1439])|(~m[204]&m[610]&m[1439]))&BiasedRNG[577])|(((m[204]&m[610]&~m[1439]))&~BiasedRNG[577])|((m[204]&m[610]&m[1439]));
    m[867] = (((m[220]&~m[611]&m[1509])|(~m[220]&m[611]&m[1509]))&BiasedRNG[578])|(((m[220]&m[611]&~m[1509]))&~BiasedRNG[578])|((m[220]&m[611]&m[1509]));
    m[868] = (((m[236]&~m[612]&m[1584])|(~m[236]&m[612]&m[1584]))&BiasedRNG[579])|(((m[236]&m[612]&~m[1584]))&~BiasedRNG[579])|((m[236]&m[612]&m[1584]));
    m[869] = (((m[252]&~m[613]&m[1654])|(~m[252]&m[613]&m[1654]))&BiasedRNG[580])|(((m[252]&m[613]&~m[1654]))&~BiasedRNG[580])|((m[252]&m[613]&m[1654]));
    m[870] = (((m[268]&~m[614]&m[1719])|(~m[268]&m[614]&m[1719]))&BiasedRNG[581])|(((m[268]&m[614]&~m[1719]))&~BiasedRNG[581])|((m[268]&m[614]&m[1719]));
    m[871] = (((m[284]&~m[615]&m[1779])|(~m[284]&m[615]&m[1779]))&BiasedRNG[582])|(((m[284]&m[615]&~m[1779]))&~BiasedRNG[582])|((m[284]&m[615]&m[1779]));
    m[872] = (((m[300]&~m[616]&m[1834])|(~m[300]&m[616]&m[1834]))&BiasedRNG[583])|(((m[300]&m[616]&~m[1834]))&~BiasedRNG[583])|((m[300]&m[616]&m[1834]));
    m[873] = (((m[316]&~m[617]&m[1884])|(~m[316]&m[617]&m[1884]))&BiasedRNG[584])|(((m[316]&m[617]&~m[1884]))&~BiasedRNG[584])|((m[316]&m[617]&m[1884]));
    m[874] = (((m[332]&~m[618]&m[1929])|(~m[332]&m[618]&m[1929]))&BiasedRNG[585])|(((m[332]&m[618]&~m[1929]))&~BiasedRNG[585])|((m[332]&m[618]&m[1929]));
    m[875] = (((m[348]&~m[619]&m[1969])|(~m[348]&m[619]&m[1969]))&BiasedRNG[586])|(((m[348]&m[619]&~m[1969]))&~BiasedRNG[586])|((m[348]&m[619]&m[1969]));
    m[876] = (((m[364]&~m[620]&m[2004])|(~m[364]&m[620]&m[2004]))&BiasedRNG[587])|(((m[364]&m[620]&~m[2004]))&~BiasedRNG[587])|((m[364]&m[620]&m[2004]));
    m[877] = (((m[380]&~m[621]&m[2034])|(~m[380]&m[621]&m[2034]))&BiasedRNG[588])|(((m[380]&m[621]&~m[2034]))&~BiasedRNG[588])|((m[380]&m[621]&m[2034]));
    m[878] = (((m[396]&~m[622]&m[2059])|(~m[396]&m[622]&m[2059]))&BiasedRNG[589])|(((m[396]&m[622]&~m[2059]))&~BiasedRNG[589])|((m[396]&m[622]&m[2059]));
    m[879] = (((m[412]&~m[623]&m[2079])|(~m[412]&m[623]&m[2079]))&BiasedRNG[590])|(((m[412]&m[623]&~m[2079]))&~BiasedRNG[590])|((m[412]&m[623]&m[2079]));
    m[880] = (((m[173]&~m[624]&m[1379])|(~m[173]&m[624]&m[1379]))&BiasedRNG[591])|(((m[173]&m[624]&~m[1379]))&~BiasedRNG[591])|((m[173]&m[624]&m[1379]));
    m[881] = (((m[189]&~m[625]&m[1444])|(~m[189]&m[625]&m[1444]))&BiasedRNG[592])|(((m[189]&m[625]&~m[1444]))&~BiasedRNG[592])|((m[189]&m[625]&m[1444]));
    m[882] = (((m[205]&~m[626]&m[1514])|(~m[205]&m[626]&m[1514]))&BiasedRNG[593])|(((m[205]&m[626]&~m[1514]))&~BiasedRNG[593])|((m[205]&m[626]&m[1514]));
    m[883] = (((m[221]&~m[627]&m[1589])|(~m[221]&m[627]&m[1589]))&BiasedRNG[594])|(((m[221]&m[627]&~m[1589]))&~BiasedRNG[594])|((m[221]&m[627]&m[1589]));
    m[884] = (((m[237]&~m[628]&m[1659])|(~m[237]&m[628]&m[1659]))&BiasedRNG[595])|(((m[237]&m[628]&~m[1659]))&~BiasedRNG[595])|((m[237]&m[628]&m[1659]));
    m[885] = (((m[253]&~m[629]&m[1724])|(~m[253]&m[629]&m[1724]))&BiasedRNG[596])|(((m[253]&m[629]&~m[1724]))&~BiasedRNG[596])|((m[253]&m[629]&m[1724]));
    m[886] = (((m[269]&~m[630]&m[1784])|(~m[269]&m[630]&m[1784]))&BiasedRNG[597])|(((m[269]&m[630]&~m[1784]))&~BiasedRNG[597])|((m[269]&m[630]&m[1784]));
    m[887] = (((m[285]&~m[631]&m[1839])|(~m[285]&m[631]&m[1839]))&BiasedRNG[598])|(((m[285]&m[631]&~m[1839]))&~BiasedRNG[598])|((m[285]&m[631]&m[1839]));
    m[888] = (((m[301]&~m[632]&m[1889])|(~m[301]&m[632]&m[1889]))&BiasedRNG[599])|(((m[301]&m[632]&~m[1889]))&~BiasedRNG[599])|((m[301]&m[632]&m[1889]));
    m[889] = (((m[317]&~m[633]&m[1934])|(~m[317]&m[633]&m[1934]))&BiasedRNG[600])|(((m[317]&m[633]&~m[1934]))&~BiasedRNG[600])|((m[317]&m[633]&m[1934]));
    m[890] = (((m[333]&~m[634]&m[1974])|(~m[333]&m[634]&m[1974]))&BiasedRNG[601])|(((m[333]&m[634]&~m[1974]))&~BiasedRNG[601])|((m[333]&m[634]&m[1974]));
    m[891] = (((m[349]&~m[635]&m[2009])|(~m[349]&m[635]&m[2009]))&BiasedRNG[602])|(((m[349]&m[635]&~m[2009]))&~BiasedRNG[602])|((m[349]&m[635]&m[2009]));
    m[892] = (((m[365]&~m[636]&m[2039])|(~m[365]&m[636]&m[2039]))&BiasedRNG[603])|(((m[365]&m[636]&~m[2039]))&~BiasedRNG[603])|((m[365]&m[636]&m[2039]));
    m[893] = (((m[381]&~m[637]&m[2064])|(~m[381]&m[637]&m[2064]))&BiasedRNG[604])|(((m[381]&m[637]&~m[2064]))&~BiasedRNG[604])|((m[381]&m[637]&m[2064]));
    m[894] = (((m[397]&~m[638]&m[2084])|(~m[397]&m[638]&m[2084]))&BiasedRNG[605])|(((m[397]&m[638]&~m[2084]))&~BiasedRNG[605])|((m[397]&m[638]&m[2084]));
    m[895] = (((m[413]&~m[639]&m[2099])|(~m[413]&m[639]&m[2099]))&BiasedRNG[606])|(((m[413]&m[639]&~m[2099]))&~BiasedRNG[606])|((m[413]&m[639]&m[2099]));
    m[896] = (((m[174]&~m[640]&m[1449])|(~m[174]&m[640]&m[1449]))&BiasedRNG[607])|(((m[174]&m[640]&~m[1449]))&~BiasedRNG[607])|((m[174]&m[640]&m[1449]));
    m[897] = (((m[190]&~m[641]&m[1519])|(~m[190]&m[641]&m[1519]))&BiasedRNG[608])|(((m[190]&m[641]&~m[1519]))&~BiasedRNG[608])|((m[190]&m[641]&m[1519]));
    m[898] = (((m[206]&~m[642]&m[1594])|(~m[206]&m[642]&m[1594]))&BiasedRNG[609])|(((m[206]&m[642]&~m[1594]))&~BiasedRNG[609])|((m[206]&m[642]&m[1594]));
    m[899] = (((m[222]&~m[643]&m[1664])|(~m[222]&m[643]&m[1664]))&BiasedRNG[610])|(((m[222]&m[643]&~m[1664]))&~BiasedRNG[610])|((m[222]&m[643]&m[1664]));
    m[900] = (((m[238]&~m[644]&m[1729])|(~m[238]&m[644]&m[1729]))&BiasedRNG[611])|(((m[238]&m[644]&~m[1729]))&~BiasedRNG[611])|((m[238]&m[644]&m[1729]));
    m[901] = (((m[254]&~m[645]&m[1789])|(~m[254]&m[645]&m[1789]))&BiasedRNG[612])|(((m[254]&m[645]&~m[1789]))&~BiasedRNG[612])|((m[254]&m[645]&m[1789]));
    m[902] = (((m[270]&~m[646]&m[1844])|(~m[270]&m[646]&m[1844]))&BiasedRNG[613])|(((m[270]&m[646]&~m[1844]))&~BiasedRNG[613])|((m[270]&m[646]&m[1844]));
    m[903] = (((m[286]&~m[647]&m[1894])|(~m[286]&m[647]&m[1894]))&BiasedRNG[614])|(((m[286]&m[647]&~m[1894]))&~BiasedRNG[614])|((m[286]&m[647]&m[1894]));
    m[904] = (((m[302]&~m[648]&m[1939])|(~m[302]&m[648]&m[1939]))&BiasedRNG[615])|(((m[302]&m[648]&~m[1939]))&~BiasedRNG[615])|((m[302]&m[648]&m[1939]));
    m[905] = (((m[318]&~m[649]&m[1979])|(~m[318]&m[649]&m[1979]))&BiasedRNG[616])|(((m[318]&m[649]&~m[1979]))&~BiasedRNG[616])|((m[318]&m[649]&m[1979]));
    m[906] = (((m[334]&~m[650]&m[2014])|(~m[334]&m[650]&m[2014]))&BiasedRNG[617])|(((m[334]&m[650]&~m[2014]))&~BiasedRNG[617])|((m[334]&m[650]&m[2014]));
    m[907] = (((m[350]&~m[651]&m[2044])|(~m[350]&m[651]&m[2044]))&BiasedRNG[618])|(((m[350]&m[651]&~m[2044]))&~BiasedRNG[618])|((m[350]&m[651]&m[2044]));
    m[908] = (((m[366]&~m[652]&m[2069])|(~m[366]&m[652]&m[2069]))&BiasedRNG[619])|(((m[366]&m[652]&~m[2069]))&~BiasedRNG[619])|((m[366]&m[652]&m[2069]));
    m[909] = (((m[382]&~m[653]&m[2089])|(~m[382]&m[653]&m[2089]))&BiasedRNG[620])|(((m[382]&m[653]&~m[2089]))&~BiasedRNG[620])|((m[382]&m[653]&m[2089]));
    m[910] = (((m[398]&~m[654]&m[2104])|(~m[398]&m[654]&m[2104]))&BiasedRNG[621])|(((m[398]&m[654]&~m[2104]))&~BiasedRNG[621])|((m[398]&m[654]&m[2104]));
    m[911] = (((m[414]&~m[655]&m[2114])|(~m[414]&m[655]&m[2114]))&BiasedRNG[622])|(((m[414]&m[655]&~m[2114]))&~BiasedRNG[622])|((m[414]&m[655]&m[2114]));
    m[912] = (((m[175]&~m[656]&m[1524])|(~m[175]&m[656]&m[1524]))&BiasedRNG[623])|(((m[175]&m[656]&~m[1524]))&~BiasedRNG[623])|((m[175]&m[656]&m[1524]));
    m[913] = (((m[191]&~m[657]&m[1599])|(~m[191]&m[657]&m[1599]))&BiasedRNG[624])|(((m[191]&m[657]&~m[1599]))&~BiasedRNG[624])|((m[191]&m[657]&m[1599]));
    m[914] = (((m[207]&~m[658]&m[1669])|(~m[207]&m[658]&m[1669]))&BiasedRNG[625])|(((m[207]&m[658]&~m[1669]))&~BiasedRNG[625])|((m[207]&m[658]&m[1669]));
    m[915] = (((m[223]&~m[659]&m[1734])|(~m[223]&m[659]&m[1734]))&BiasedRNG[626])|(((m[223]&m[659]&~m[1734]))&~BiasedRNG[626])|((m[223]&m[659]&m[1734]));
    m[916] = (((m[239]&~m[660]&m[1794])|(~m[239]&m[660]&m[1794]))&BiasedRNG[627])|(((m[239]&m[660]&~m[1794]))&~BiasedRNG[627])|((m[239]&m[660]&m[1794]));
    m[917] = (((m[255]&~m[661]&m[1849])|(~m[255]&m[661]&m[1849]))&BiasedRNG[628])|(((m[255]&m[661]&~m[1849]))&~BiasedRNG[628])|((m[255]&m[661]&m[1849]));
    m[918] = (((m[271]&~m[662]&m[1899])|(~m[271]&m[662]&m[1899]))&BiasedRNG[629])|(((m[271]&m[662]&~m[1899]))&~BiasedRNG[629])|((m[271]&m[662]&m[1899]));
    m[919] = (((m[287]&~m[663]&m[1944])|(~m[287]&m[663]&m[1944]))&BiasedRNG[630])|(((m[287]&m[663]&~m[1944]))&~BiasedRNG[630])|((m[287]&m[663]&m[1944]));
    m[920] = (((m[303]&~m[664]&m[1984])|(~m[303]&m[664]&m[1984]))&BiasedRNG[631])|(((m[303]&m[664]&~m[1984]))&~BiasedRNG[631])|((m[303]&m[664]&m[1984]));
    m[921] = (((m[319]&~m[665]&m[2019])|(~m[319]&m[665]&m[2019]))&BiasedRNG[632])|(((m[319]&m[665]&~m[2019]))&~BiasedRNG[632])|((m[319]&m[665]&m[2019]));
    m[922] = (((m[335]&~m[666]&m[2049])|(~m[335]&m[666]&m[2049]))&BiasedRNG[633])|(((m[335]&m[666]&~m[2049]))&~BiasedRNG[633])|((m[335]&m[666]&m[2049]));
    m[923] = (((m[351]&~m[667]&m[2074])|(~m[351]&m[667]&m[2074]))&BiasedRNG[634])|(((m[351]&m[667]&~m[2074]))&~BiasedRNG[634])|((m[351]&m[667]&m[2074]));
    m[924] = (((m[367]&~m[668]&m[2094])|(~m[367]&m[668]&m[2094]))&BiasedRNG[635])|(((m[367]&m[668]&~m[2094]))&~BiasedRNG[635])|((m[367]&m[668]&m[2094]));
    m[925] = (((m[383]&~m[669]&m[2109])|(~m[383]&m[669]&m[2109]))&BiasedRNG[636])|(((m[383]&m[669]&~m[2109]))&~BiasedRNG[636])|((m[383]&m[669]&m[2109]));
    m[926] = (((m[399]&~m[670]&m[2119])|(~m[399]&m[670]&m[2119]))&BiasedRNG[637])|(((m[399]&m[670]&~m[2119]))&~BiasedRNG[637])|((m[399]&m[670]&m[2119]));
    m[927] = (((m[415]&~m[671]&m[2124])|(~m[415]&m[671]&m[2124]))&BiasedRNG[638])|(((m[415]&m[671]&~m[2124]))&~BiasedRNG[638])|((m[415]&m[671]&m[2124]));
    m[935] = (((m[932]&~m[933]&~m[934]&~m[936]&~m[937])|(~m[932]&~m[933]&~m[934]&m[936]&~m[937])|(m[932]&m[933]&~m[934]&m[936]&~m[937])|(m[932]&~m[933]&m[934]&m[936]&~m[937])|(~m[932]&m[933]&~m[934]&~m[936]&m[937])|(~m[932]&~m[933]&m[934]&~m[936]&m[937])|(m[932]&m[933]&m[934]&~m[936]&m[937])|(~m[932]&m[933]&m[934]&m[936]&m[937]))&UnbiasedRNG[271])|((m[932]&~m[933]&~m[934]&m[936]&~m[937])|(~m[932]&~m[933]&~m[934]&~m[936]&m[937])|(m[932]&~m[933]&~m[934]&~m[936]&m[937])|(m[932]&m[933]&~m[934]&~m[936]&m[937])|(m[932]&~m[933]&m[934]&~m[936]&m[937])|(~m[932]&~m[933]&~m[934]&m[936]&m[937])|(m[932]&~m[933]&~m[934]&m[936]&m[937])|(~m[932]&m[933]&~m[934]&m[936]&m[937])|(m[932]&m[933]&~m[934]&m[936]&m[937])|(~m[932]&~m[933]&m[934]&m[936]&m[937])|(m[932]&~m[933]&m[934]&m[936]&m[937])|(m[932]&m[933]&m[934]&m[936]&m[937]));
    m[945] = (((m[937]&~m[943]&~m[944]&~m[946]&~m[947])|(~m[937]&~m[943]&~m[944]&m[946]&~m[947])|(m[937]&m[943]&~m[944]&m[946]&~m[947])|(m[937]&~m[943]&m[944]&m[946]&~m[947])|(~m[937]&m[943]&~m[944]&~m[946]&m[947])|(~m[937]&~m[943]&m[944]&~m[946]&m[947])|(m[937]&m[943]&m[944]&~m[946]&m[947])|(~m[937]&m[943]&m[944]&m[946]&m[947]))&UnbiasedRNG[272])|((m[937]&~m[943]&~m[944]&m[946]&~m[947])|(~m[937]&~m[943]&~m[944]&~m[946]&m[947])|(m[937]&~m[943]&~m[944]&~m[946]&m[947])|(m[937]&m[943]&~m[944]&~m[946]&m[947])|(m[937]&~m[943]&m[944]&~m[946]&m[947])|(~m[937]&~m[943]&~m[944]&m[946]&m[947])|(m[937]&~m[943]&~m[944]&m[946]&m[947])|(~m[937]&m[943]&~m[944]&m[946]&m[947])|(m[937]&m[943]&~m[944]&m[946]&m[947])|(~m[937]&~m[943]&m[944]&m[946]&m[947])|(m[937]&~m[943]&m[944]&m[946]&m[947])|(m[937]&m[943]&m[944]&m[946]&m[947]));
    m[950] = (((m[942]&~m[948]&~m[949]&~m[951]&~m[952])|(~m[942]&~m[948]&~m[949]&m[951]&~m[952])|(m[942]&m[948]&~m[949]&m[951]&~m[952])|(m[942]&~m[948]&m[949]&m[951]&~m[952])|(~m[942]&m[948]&~m[949]&~m[951]&m[952])|(~m[942]&~m[948]&m[949]&~m[951]&m[952])|(m[942]&m[948]&m[949]&~m[951]&m[952])|(~m[942]&m[948]&m[949]&m[951]&m[952]))&UnbiasedRNG[273])|((m[942]&~m[948]&~m[949]&m[951]&~m[952])|(~m[942]&~m[948]&~m[949]&~m[951]&m[952])|(m[942]&~m[948]&~m[949]&~m[951]&m[952])|(m[942]&m[948]&~m[949]&~m[951]&m[952])|(m[942]&~m[948]&m[949]&~m[951]&m[952])|(~m[942]&~m[948]&~m[949]&m[951]&m[952])|(m[942]&~m[948]&~m[949]&m[951]&m[952])|(~m[942]&m[948]&~m[949]&m[951]&m[952])|(m[942]&m[948]&~m[949]&m[951]&m[952])|(~m[942]&~m[948]&m[949]&m[951]&m[952])|(m[942]&~m[948]&m[949]&m[951]&m[952])|(m[942]&m[948]&m[949]&m[951]&m[952]));
    m[960] = (((m[947]&~m[958]&~m[959]&~m[961]&~m[962])|(~m[947]&~m[958]&~m[959]&m[961]&~m[962])|(m[947]&m[958]&~m[959]&m[961]&~m[962])|(m[947]&~m[958]&m[959]&m[961]&~m[962])|(~m[947]&m[958]&~m[959]&~m[961]&m[962])|(~m[947]&~m[958]&m[959]&~m[961]&m[962])|(m[947]&m[958]&m[959]&~m[961]&m[962])|(~m[947]&m[958]&m[959]&m[961]&m[962]))&UnbiasedRNG[274])|((m[947]&~m[958]&~m[959]&m[961]&~m[962])|(~m[947]&~m[958]&~m[959]&~m[961]&m[962])|(m[947]&~m[958]&~m[959]&~m[961]&m[962])|(m[947]&m[958]&~m[959]&~m[961]&m[962])|(m[947]&~m[958]&m[959]&~m[961]&m[962])|(~m[947]&~m[958]&~m[959]&m[961]&m[962])|(m[947]&~m[958]&~m[959]&m[961]&m[962])|(~m[947]&m[958]&~m[959]&m[961]&m[962])|(m[947]&m[958]&~m[959]&m[961]&m[962])|(~m[947]&~m[958]&m[959]&m[961]&m[962])|(m[947]&~m[958]&m[959]&m[961]&m[962])|(m[947]&m[958]&m[959]&m[961]&m[962]));
    m[965] = (((m[952]&~m[963]&~m[964]&~m[966]&~m[967])|(~m[952]&~m[963]&~m[964]&m[966]&~m[967])|(m[952]&m[963]&~m[964]&m[966]&~m[967])|(m[952]&~m[963]&m[964]&m[966]&~m[967])|(~m[952]&m[963]&~m[964]&~m[966]&m[967])|(~m[952]&~m[963]&m[964]&~m[966]&m[967])|(m[952]&m[963]&m[964]&~m[966]&m[967])|(~m[952]&m[963]&m[964]&m[966]&m[967]))&UnbiasedRNG[275])|((m[952]&~m[963]&~m[964]&m[966]&~m[967])|(~m[952]&~m[963]&~m[964]&~m[966]&m[967])|(m[952]&~m[963]&~m[964]&~m[966]&m[967])|(m[952]&m[963]&~m[964]&~m[966]&m[967])|(m[952]&~m[963]&m[964]&~m[966]&m[967])|(~m[952]&~m[963]&~m[964]&m[966]&m[967])|(m[952]&~m[963]&~m[964]&m[966]&m[967])|(~m[952]&m[963]&~m[964]&m[966]&m[967])|(m[952]&m[963]&~m[964]&m[966]&m[967])|(~m[952]&~m[963]&m[964]&m[966]&m[967])|(m[952]&~m[963]&m[964]&m[966]&m[967])|(m[952]&m[963]&m[964]&m[966]&m[967]));
    m[970] = (((m[957]&~m[968]&~m[969]&~m[971]&~m[972])|(~m[957]&~m[968]&~m[969]&m[971]&~m[972])|(m[957]&m[968]&~m[969]&m[971]&~m[972])|(m[957]&~m[968]&m[969]&m[971]&~m[972])|(~m[957]&m[968]&~m[969]&~m[971]&m[972])|(~m[957]&~m[968]&m[969]&~m[971]&m[972])|(m[957]&m[968]&m[969]&~m[971]&m[972])|(~m[957]&m[968]&m[969]&m[971]&m[972]))&UnbiasedRNG[276])|((m[957]&~m[968]&~m[969]&m[971]&~m[972])|(~m[957]&~m[968]&~m[969]&~m[971]&m[972])|(m[957]&~m[968]&~m[969]&~m[971]&m[972])|(m[957]&m[968]&~m[969]&~m[971]&m[972])|(m[957]&~m[968]&m[969]&~m[971]&m[972])|(~m[957]&~m[968]&~m[969]&m[971]&m[972])|(m[957]&~m[968]&~m[969]&m[971]&m[972])|(~m[957]&m[968]&~m[969]&m[971]&m[972])|(m[957]&m[968]&~m[969]&m[971]&m[972])|(~m[957]&~m[968]&m[969]&m[971]&m[972])|(m[957]&~m[968]&m[969]&m[971]&m[972])|(m[957]&m[968]&m[969]&m[971]&m[972]));
    m[980] = (((m[962]&~m[978]&~m[979]&~m[981]&~m[982])|(~m[962]&~m[978]&~m[979]&m[981]&~m[982])|(m[962]&m[978]&~m[979]&m[981]&~m[982])|(m[962]&~m[978]&m[979]&m[981]&~m[982])|(~m[962]&m[978]&~m[979]&~m[981]&m[982])|(~m[962]&~m[978]&m[979]&~m[981]&m[982])|(m[962]&m[978]&m[979]&~m[981]&m[982])|(~m[962]&m[978]&m[979]&m[981]&m[982]))&UnbiasedRNG[277])|((m[962]&~m[978]&~m[979]&m[981]&~m[982])|(~m[962]&~m[978]&~m[979]&~m[981]&m[982])|(m[962]&~m[978]&~m[979]&~m[981]&m[982])|(m[962]&m[978]&~m[979]&~m[981]&m[982])|(m[962]&~m[978]&m[979]&~m[981]&m[982])|(~m[962]&~m[978]&~m[979]&m[981]&m[982])|(m[962]&~m[978]&~m[979]&m[981]&m[982])|(~m[962]&m[978]&~m[979]&m[981]&m[982])|(m[962]&m[978]&~m[979]&m[981]&m[982])|(~m[962]&~m[978]&m[979]&m[981]&m[982])|(m[962]&~m[978]&m[979]&m[981]&m[982])|(m[962]&m[978]&m[979]&m[981]&m[982]));
    m[985] = (((m[967]&~m[983]&~m[984]&~m[986]&~m[987])|(~m[967]&~m[983]&~m[984]&m[986]&~m[987])|(m[967]&m[983]&~m[984]&m[986]&~m[987])|(m[967]&~m[983]&m[984]&m[986]&~m[987])|(~m[967]&m[983]&~m[984]&~m[986]&m[987])|(~m[967]&~m[983]&m[984]&~m[986]&m[987])|(m[967]&m[983]&m[984]&~m[986]&m[987])|(~m[967]&m[983]&m[984]&m[986]&m[987]))&UnbiasedRNG[278])|((m[967]&~m[983]&~m[984]&m[986]&~m[987])|(~m[967]&~m[983]&~m[984]&~m[986]&m[987])|(m[967]&~m[983]&~m[984]&~m[986]&m[987])|(m[967]&m[983]&~m[984]&~m[986]&m[987])|(m[967]&~m[983]&m[984]&~m[986]&m[987])|(~m[967]&~m[983]&~m[984]&m[986]&m[987])|(m[967]&~m[983]&~m[984]&m[986]&m[987])|(~m[967]&m[983]&~m[984]&m[986]&m[987])|(m[967]&m[983]&~m[984]&m[986]&m[987])|(~m[967]&~m[983]&m[984]&m[986]&m[987])|(m[967]&~m[983]&m[984]&m[986]&m[987])|(m[967]&m[983]&m[984]&m[986]&m[987]));
    m[990] = (((m[972]&~m[988]&~m[989]&~m[991]&~m[992])|(~m[972]&~m[988]&~m[989]&m[991]&~m[992])|(m[972]&m[988]&~m[989]&m[991]&~m[992])|(m[972]&~m[988]&m[989]&m[991]&~m[992])|(~m[972]&m[988]&~m[989]&~m[991]&m[992])|(~m[972]&~m[988]&m[989]&~m[991]&m[992])|(m[972]&m[988]&m[989]&~m[991]&m[992])|(~m[972]&m[988]&m[989]&m[991]&m[992]))&UnbiasedRNG[279])|((m[972]&~m[988]&~m[989]&m[991]&~m[992])|(~m[972]&~m[988]&~m[989]&~m[991]&m[992])|(m[972]&~m[988]&~m[989]&~m[991]&m[992])|(m[972]&m[988]&~m[989]&~m[991]&m[992])|(m[972]&~m[988]&m[989]&~m[991]&m[992])|(~m[972]&~m[988]&~m[989]&m[991]&m[992])|(m[972]&~m[988]&~m[989]&m[991]&m[992])|(~m[972]&m[988]&~m[989]&m[991]&m[992])|(m[972]&m[988]&~m[989]&m[991]&m[992])|(~m[972]&~m[988]&m[989]&m[991]&m[992])|(m[972]&~m[988]&m[989]&m[991]&m[992])|(m[972]&m[988]&m[989]&m[991]&m[992]));
    m[995] = (((m[977]&~m[993]&~m[994]&~m[996]&~m[997])|(~m[977]&~m[993]&~m[994]&m[996]&~m[997])|(m[977]&m[993]&~m[994]&m[996]&~m[997])|(m[977]&~m[993]&m[994]&m[996]&~m[997])|(~m[977]&m[993]&~m[994]&~m[996]&m[997])|(~m[977]&~m[993]&m[994]&~m[996]&m[997])|(m[977]&m[993]&m[994]&~m[996]&m[997])|(~m[977]&m[993]&m[994]&m[996]&m[997]))&UnbiasedRNG[280])|((m[977]&~m[993]&~m[994]&m[996]&~m[997])|(~m[977]&~m[993]&~m[994]&~m[996]&m[997])|(m[977]&~m[993]&~m[994]&~m[996]&m[997])|(m[977]&m[993]&~m[994]&~m[996]&m[997])|(m[977]&~m[993]&m[994]&~m[996]&m[997])|(~m[977]&~m[993]&~m[994]&m[996]&m[997])|(m[977]&~m[993]&~m[994]&m[996]&m[997])|(~m[977]&m[993]&~m[994]&m[996]&m[997])|(m[977]&m[993]&~m[994]&m[996]&m[997])|(~m[977]&~m[993]&m[994]&m[996]&m[997])|(m[977]&~m[993]&m[994]&m[996]&m[997])|(m[977]&m[993]&m[994]&m[996]&m[997]));
    m[1005] = (((m[982]&~m[1003]&~m[1004]&~m[1006]&~m[1007])|(~m[982]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(m[982]&m[1003]&~m[1004]&m[1006]&~m[1007])|(m[982]&~m[1003]&m[1004]&m[1006]&~m[1007])|(~m[982]&m[1003]&~m[1004]&~m[1006]&m[1007])|(~m[982]&~m[1003]&m[1004]&~m[1006]&m[1007])|(m[982]&m[1003]&m[1004]&~m[1006]&m[1007])|(~m[982]&m[1003]&m[1004]&m[1006]&m[1007]))&UnbiasedRNG[281])|((m[982]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(~m[982]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[982]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[982]&m[1003]&~m[1004]&~m[1006]&m[1007])|(m[982]&~m[1003]&m[1004]&~m[1006]&m[1007])|(~m[982]&~m[1003]&~m[1004]&m[1006]&m[1007])|(m[982]&~m[1003]&~m[1004]&m[1006]&m[1007])|(~m[982]&m[1003]&~m[1004]&m[1006]&m[1007])|(m[982]&m[1003]&~m[1004]&m[1006]&m[1007])|(~m[982]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[982]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[982]&m[1003]&m[1004]&m[1006]&m[1007]));
    m[1010] = (((m[987]&~m[1008]&~m[1009]&~m[1011]&~m[1012])|(~m[987]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(m[987]&m[1008]&~m[1009]&m[1011]&~m[1012])|(m[987]&~m[1008]&m[1009]&m[1011]&~m[1012])|(~m[987]&m[1008]&~m[1009]&~m[1011]&m[1012])|(~m[987]&~m[1008]&m[1009]&~m[1011]&m[1012])|(m[987]&m[1008]&m[1009]&~m[1011]&m[1012])|(~m[987]&m[1008]&m[1009]&m[1011]&m[1012]))&UnbiasedRNG[282])|((m[987]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(~m[987]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[987]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[987]&m[1008]&~m[1009]&~m[1011]&m[1012])|(m[987]&~m[1008]&m[1009]&~m[1011]&m[1012])|(~m[987]&~m[1008]&~m[1009]&m[1011]&m[1012])|(m[987]&~m[1008]&~m[1009]&m[1011]&m[1012])|(~m[987]&m[1008]&~m[1009]&m[1011]&m[1012])|(m[987]&m[1008]&~m[1009]&m[1011]&m[1012])|(~m[987]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[987]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[987]&m[1008]&m[1009]&m[1011]&m[1012]));
    m[1015] = (((m[992]&~m[1013]&~m[1014]&~m[1016]&~m[1017])|(~m[992]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(m[992]&m[1013]&~m[1014]&m[1016]&~m[1017])|(m[992]&~m[1013]&m[1014]&m[1016]&~m[1017])|(~m[992]&m[1013]&~m[1014]&~m[1016]&m[1017])|(~m[992]&~m[1013]&m[1014]&~m[1016]&m[1017])|(m[992]&m[1013]&m[1014]&~m[1016]&m[1017])|(~m[992]&m[1013]&m[1014]&m[1016]&m[1017]))&UnbiasedRNG[283])|((m[992]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(~m[992]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[992]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[992]&m[1013]&~m[1014]&~m[1016]&m[1017])|(m[992]&~m[1013]&m[1014]&~m[1016]&m[1017])|(~m[992]&~m[1013]&~m[1014]&m[1016]&m[1017])|(m[992]&~m[1013]&~m[1014]&m[1016]&m[1017])|(~m[992]&m[1013]&~m[1014]&m[1016]&m[1017])|(m[992]&m[1013]&~m[1014]&m[1016]&m[1017])|(~m[992]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[992]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[992]&m[1013]&m[1014]&m[1016]&m[1017]));
    m[1020] = (((m[997]&~m[1018]&~m[1019]&~m[1021]&~m[1022])|(~m[997]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(m[997]&m[1018]&~m[1019]&m[1021]&~m[1022])|(m[997]&~m[1018]&m[1019]&m[1021]&~m[1022])|(~m[997]&m[1018]&~m[1019]&~m[1021]&m[1022])|(~m[997]&~m[1018]&m[1019]&~m[1021]&m[1022])|(m[997]&m[1018]&m[1019]&~m[1021]&m[1022])|(~m[997]&m[1018]&m[1019]&m[1021]&m[1022]))&UnbiasedRNG[284])|((m[997]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(~m[997]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[997]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[997]&m[1018]&~m[1019]&~m[1021]&m[1022])|(m[997]&~m[1018]&m[1019]&~m[1021]&m[1022])|(~m[997]&~m[1018]&~m[1019]&m[1021]&m[1022])|(m[997]&~m[1018]&~m[1019]&m[1021]&m[1022])|(~m[997]&m[1018]&~m[1019]&m[1021]&m[1022])|(m[997]&m[1018]&~m[1019]&m[1021]&m[1022])|(~m[997]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[997]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[997]&m[1018]&m[1019]&m[1021]&m[1022]));
    m[1025] = (((m[1002]&~m[1023]&~m[1024]&~m[1026]&~m[1027])|(~m[1002]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(m[1002]&m[1023]&~m[1024]&m[1026]&~m[1027])|(m[1002]&~m[1023]&m[1024]&m[1026]&~m[1027])|(~m[1002]&m[1023]&~m[1024]&~m[1026]&m[1027])|(~m[1002]&~m[1023]&m[1024]&~m[1026]&m[1027])|(m[1002]&m[1023]&m[1024]&~m[1026]&m[1027])|(~m[1002]&m[1023]&m[1024]&m[1026]&m[1027]))&UnbiasedRNG[285])|((m[1002]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(~m[1002]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[1002]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[1002]&m[1023]&~m[1024]&~m[1026]&m[1027])|(m[1002]&~m[1023]&m[1024]&~m[1026]&m[1027])|(~m[1002]&~m[1023]&~m[1024]&m[1026]&m[1027])|(m[1002]&~m[1023]&~m[1024]&m[1026]&m[1027])|(~m[1002]&m[1023]&~m[1024]&m[1026]&m[1027])|(m[1002]&m[1023]&~m[1024]&m[1026]&m[1027])|(~m[1002]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[1002]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[1002]&m[1023]&m[1024]&m[1026]&m[1027]));
    m[1035] = (((m[1007]&~m[1033]&~m[1034]&~m[1036]&~m[1037])|(~m[1007]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(m[1007]&m[1033]&~m[1034]&m[1036]&~m[1037])|(m[1007]&~m[1033]&m[1034]&m[1036]&~m[1037])|(~m[1007]&m[1033]&~m[1034]&~m[1036]&m[1037])|(~m[1007]&~m[1033]&m[1034]&~m[1036]&m[1037])|(m[1007]&m[1033]&m[1034]&~m[1036]&m[1037])|(~m[1007]&m[1033]&m[1034]&m[1036]&m[1037]))&UnbiasedRNG[286])|((m[1007]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(~m[1007]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[1007]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[1007]&m[1033]&~m[1034]&~m[1036]&m[1037])|(m[1007]&~m[1033]&m[1034]&~m[1036]&m[1037])|(~m[1007]&~m[1033]&~m[1034]&m[1036]&m[1037])|(m[1007]&~m[1033]&~m[1034]&m[1036]&m[1037])|(~m[1007]&m[1033]&~m[1034]&m[1036]&m[1037])|(m[1007]&m[1033]&~m[1034]&m[1036]&m[1037])|(~m[1007]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[1007]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[1007]&m[1033]&m[1034]&m[1036]&m[1037]));
    m[1040] = (((m[1012]&~m[1038]&~m[1039]&~m[1041]&~m[1042])|(~m[1012]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1012]&m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1012]&~m[1038]&m[1039]&m[1041]&~m[1042])|(~m[1012]&m[1038]&~m[1039]&~m[1041]&m[1042])|(~m[1012]&~m[1038]&m[1039]&~m[1041]&m[1042])|(m[1012]&m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1012]&m[1038]&m[1039]&m[1041]&m[1042]))&UnbiasedRNG[287])|((m[1012]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(~m[1012]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1012]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1012]&m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1012]&~m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1012]&~m[1038]&~m[1039]&m[1041]&m[1042])|(m[1012]&~m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1012]&m[1038]&~m[1039]&m[1041]&m[1042])|(m[1012]&m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1012]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1012]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1012]&m[1038]&m[1039]&m[1041]&m[1042]));
    m[1045] = (((m[1017]&~m[1043]&~m[1044]&~m[1046]&~m[1047])|(~m[1017]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1017]&m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1017]&~m[1043]&m[1044]&m[1046]&~m[1047])|(~m[1017]&m[1043]&~m[1044]&~m[1046]&m[1047])|(~m[1017]&~m[1043]&m[1044]&~m[1046]&m[1047])|(m[1017]&m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1017]&m[1043]&m[1044]&m[1046]&m[1047]))&UnbiasedRNG[288])|((m[1017]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(~m[1017]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1017]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1017]&m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1017]&~m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1017]&~m[1043]&~m[1044]&m[1046]&m[1047])|(m[1017]&~m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1017]&m[1043]&~m[1044]&m[1046]&m[1047])|(m[1017]&m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1017]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1017]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1017]&m[1043]&m[1044]&m[1046]&m[1047]));
    m[1050] = (((m[1022]&~m[1048]&~m[1049]&~m[1051]&~m[1052])|(~m[1022]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1022]&m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1022]&~m[1048]&m[1049]&m[1051]&~m[1052])|(~m[1022]&m[1048]&~m[1049]&~m[1051]&m[1052])|(~m[1022]&~m[1048]&m[1049]&~m[1051]&m[1052])|(m[1022]&m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1022]&m[1048]&m[1049]&m[1051]&m[1052]))&UnbiasedRNG[289])|((m[1022]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(~m[1022]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1022]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1022]&m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1022]&~m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1022]&~m[1048]&~m[1049]&m[1051]&m[1052])|(m[1022]&~m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1022]&m[1048]&~m[1049]&m[1051]&m[1052])|(m[1022]&m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1022]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1022]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1022]&m[1048]&m[1049]&m[1051]&m[1052]));
    m[1055] = (((m[1027]&~m[1053]&~m[1054]&~m[1056]&~m[1057])|(~m[1027]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1027]&m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1027]&~m[1053]&m[1054]&m[1056]&~m[1057])|(~m[1027]&m[1053]&~m[1054]&~m[1056]&m[1057])|(~m[1027]&~m[1053]&m[1054]&~m[1056]&m[1057])|(m[1027]&m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1027]&m[1053]&m[1054]&m[1056]&m[1057]))&UnbiasedRNG[290])|((m[1027]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(~m[1027]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1027]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1027]&m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1027]&~m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1027]&~m[1053]&~m[1054]&m[1056]&m[1057])|(m[1027]&~m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1027]&m[1053]&~m[1054]&m[1056]&m[1057])|(m[1027]&m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1027]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1027]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1027]&m[1053]&m[1054]&m[1056]&m[1057]));
    m[1060] = (((m[1032]&~m[1058]&~m[1059]&~m[1061]&~m[1062])|(~m[1032]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1032]&m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1032]&~m[1058]&m[1059]&m[1061]&~m[1062])|(~m[1032]&m[1058]&~m[1059]&~m[1061]&m[1062])|(~m[1032]&~m[1058]&m[1059]&~m[1061]&m[1062])|(m[1032]&m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1032]&m[1058]&m[1059]&m[1061]&m[1062]))&UnbiasedRNG[291])|((m[1032]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(~m[1032]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1032]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1032]&m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1032]&~m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1032]&~m[1058]&~m[1059]&m[1061]&m[1062])|(m[1032]&~m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1032]&m[1058]&~m[1059]&m[1061]&m[1062])|(m[1032]&m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1032]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1032]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1032]&m[1058]&m[1059]&m[1061]&m[1062]));
    m[1070] = (((m[1037]&~m[1068]&~m[1069]&~m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&~m[1072])|(~m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&m[1068]&m[1069]&m[1071]&m[1072]))&UnbiasedRNG[292])|((m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&m[1071]&m[1072]));
    m[1075] = (((m[1042]&~m[1073]&~m[1074]&~m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&~m[1077])|(~m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&m[1073]&m[1074]&m[1076]&m[1077]))&UnbiasedRNG[293])|((m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&m[1076]&m[1077]));
    m[1080] = (((m[1047]&~m[1078]&~m[1079]&~m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&~m[1082])|(~m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&m[1078]&m[1079]&m[1081]&m[1082]))&UnbiasedRNG[294])|((m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&m[1081]&m[1082]));
    m[1085] = (((m[1052]&~m[1083]&~m[1084]&~m[1086]&~m[1087])|(~m[1052]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1052]&m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1052]&~m[1083]&m[1084]&m[1086]&~m[1087])|(~m[1052]&m[1083]&~m[1084]&~m[1086]&m[1087])|(~m[1052]&~m[1083]&m[1084]&~m[1086]&m[1087])|(m[1052]&m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1052]&m[1083]&m[1084]&m[1086]&m[1087]))&UnbiasedRNG[295])|((m[1052]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(~m[1052]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1052]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1052]&m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1052]&~m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1052]&~m[1083]&~m[1084]&m[1086]&m[1087])|(m[1052]&~m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1052]&m[1083]&~m[1084]&m[1086]&m[1087])|(m[1052]&m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1052]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1052]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1052]&m[1083]&m[1084]&m[1086]&m[1087]));
    m[1090] = (((m[1057]&~m[1088]&~m[1089]&~m[1091]&~m[1092])|(~m[1057]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1057]&m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1057]&~m[1088]&m[1089]&m[1091]&~m[1092])|(~m[1057]&m[1088]&~m[1089]&~m[1091]&m[1092])|(~m[1057]&~m[1088]&m[1089]&~m[1091]&m[1092])|(m[1057]&m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1057]&m[1088]&m[1089]&m[1091]&m[1092]))&UnbiasedRNG[296])|((m[1057]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(~m[1057]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1057]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1057]&m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1057]&~m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1057]&~m[1088]&~m[1089]&m[1091]&m[1092])|(m[1057]&~m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1057]&m[1088]&~m[1089]&m[1091]&m[1092])|(m[1057]&m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1057]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1057]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1057]&m[1088]&m[1089]&m[1091]&m[1092]));
    m[1095] = (((m[1062]&~m[1093]&~m[1094]&~m[1096]&~m[1097])|(~m[1062]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1062]&m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1062]&~m[1093]&m[1094]&m[1096]&~m[1097])|(~m[1062]&m[1093]&~m[1094]&~m[1096]&m[1097])|(~m[1062]&~m[1093]&m[1094]&~m[1096]&m[1097])|(m[1062]&m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1062]&m[1093]&m[1094]&m[1096]&m[1097]))&UnbiasedRNG[297])|((m[1062]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(~m[1062]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1062]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1062]&m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1062]&~m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1062]&~m[1093]&~m[1094]&m[1096]&m[1097])|(m[1062]&~m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1062]&m[1093]&~m[1094]&m[1096]&m[1097])|(m[1062]&m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1062]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1062]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1062]&m[1093]&m[1094]&m[1096]&m[1097]));
    m[1100] = (((m[1067]&~m[1098]&~m[1099]&~m[1101]&~m[1102])|(~m[1067]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1067]&m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1067]&~m[1098]&m[1099]&m[1101]&~m[1102])|(~m[1067]&m[1098]&~m[1099]&~m[1101]&m[1102])|(~m[1067]&~m[1098]&m[1099]&~m[1101]&m[1102])|(m[1067]&m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1067]&m[1098]&m[1099]&m[1101]&m[1102]))&UnbiasedRNG[298])|((m[1067]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(~m[1067]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1067]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1067]&m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1067]&~m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1067]&~m[1098]&~m[1099]&m[1101]&m[1102])|(m[1067]&~m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1067]&m[1098]&~m[1099]&m[1101]&m[1102])|(m[1067]&m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1067]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1067]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1067]&m[1098]&m[1099]&m[1101]&m[1102]));
    m[1110] = (((m[1072]&~m[1108]&~m[1109]&~m[1111]&~m[1112])|(~m[1072]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1072]&m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1072]&~m[1108]&m[1109]&m[1111]&~m[1112])|(~m[1072]&m[1108]&~m[1109]&~m[1111]&m[1112])|(~m[1072]&~m[1108]&m[1109]&~m[1111]&m[1112])|(m[1072]&m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1072]&m[1108]&m[1109]&m[1111]&m[1112]))&UnbiasedRNG[299])|((m[1072]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(~m[1072]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1072]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1072]&m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1072]&~m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1072]&~m[1108]&~m[1109]&m[1111]&m[1112])|(m[1072]&~m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1072]&m[1108]&~m[1109]&m[1111]&m[1112])|(m[1072]&m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1072]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1072]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1072]&m[1108]&m[1109]&m[1111]&m[1112]));
    m[1115] = (((m[1077]&~m[1113]&~m[1114]&~m[1116]&~m[1117])|(~m[1077]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1077]&m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1077]&~m[1113]&m[1114]&m[1116]&~m[1117])|(~m[1077]&m[1113]&~m[1114]&~m[1116]&m[1117])|(~m[1077]&~m[1113]&m[1114]&~m[1116]&m[1117])|(m[1077]&m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1077]&m[1113]&m[1114]&m[1116]&m[1117]))&UnbiasedRNG[300])|((m[1077]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(~m[1077]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1077]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1077]&m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1077]&~m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1077]&~m[1113]&~m[1114]&m[1116]&m[1117])|(m[1077]&~m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1077]&m[1113]&~m[1114]&m[1116]&m[1117])|(m[1077]&m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1077]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1077]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1077]&m[1113]&m[1114]&m[1116]&m[1117]));
    m[1120] = (((m[1082]&~m[1118]&~m[1119]&~m[1121]&~m[1122])|(~m[1082]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1082]&m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1082]&~m[1118]&m[1119]&m[1121]&~m[1122])|(~m[1082]&m[1118]&~m[1119]&~m[1121]&m[1122])|(~m[1082]&~m[1118]&m[1119]&~m[1121]&m[1122])|(m[1082]&m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1082]&m[1118]&m[1119]&m[1121]&m[1122]))&UnbiasedRNG[301])|((m[1082]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(~m[1082]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1082]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1082]&m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1082]&~m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1082]&~m[1118]&~m[1119]&m[1121]&m[1122])|(m[1082]&~m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1082]&m[1118]&~m[1119]&m[1121]&m[1122])|(m[1082]&m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1082]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1082]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1082]&m[1118]&m[1119]&m[1121]&m[1122]));
    m[1125] = (((m[1087]&~m[1123]&~m[1124]&~m[1126]&~m[1127])|(~m[1087]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1087]&m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1087]&~m[1123]&m[1124]&m[1126]&~m[1127])|(~m[1087]&m[1123]&~m[1124]&~m[1126]&m[1127])|(~m[1087]&~m[1123]&m[1124]&~m[1126]&m[1127])|(m[1087]&m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1087]&m[1123]&m[1124]&m[1126]&m[1127]))&UnbiasedRNG[302])|((m[1087]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(~m[1087]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1087]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1087]&m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1087]&~m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1087]&~m[1123]&~m[1124]&m[1126]&m[1127])|(m[1087]&~m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1087]&m[1123]&~m[1124]&m[1126]&m[1127])|(m[1087]&m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1087]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1087]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1087]&m[1123]&m[1124]&m[1126]&m[1127]));
    m[1130] = (((m[1092]&~m[1128]&~m[1129]&~m[1131]&~m[1132])|(~m[1092]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1092]&m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1092]&~m[1128]&m[1129]&m[1131]&~m[1132])|(~m[1092]&m[1128]&~m[1129]&~m[1131]&m[1132])|(~m[1092]&~m[1128]&m[1129]&~m[1131]&m[1132])|(m[1092]&m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1092]&m[1128]&m[1129]&m[1131]&m[1132]))&UnbiasedRNG[303])|((m[1092]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(~m[1092]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1092]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1092]&m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1092]&~m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1092]&~m[1128]&~m[1129]&m[1131]&m[1132])|(m[1092]&~m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1092]&m[1128]&~m[1129]&m[1131]&m[1132])|(m[1092]&m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1092]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1092]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1092]&m[1128]&m[1129]&m[1131]&m[1132]));
    m[1135] = (((m[1097]&~m[1133]&~m[1134]&~m[1136]&~m[1137])|(~m[1097]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1097]&m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1097]&~m[1133]&m[1134]&m[1136]&~m[1137])|(~m[1097]&m[1133]&~m[1134]&~m[1136]&m[1137])|(~m[1097]&~m[1133]&m[1134]&~m[1136]&m[1137])|(m[1097]&m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1097]&m[1133]&m[1134]&m[1136]&m[1137]))&UnbiasedRNG[304])|((m[1097]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(~m[1097]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1097]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1097]&m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1097]&~m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1097]&~m[1133]&~m[1134]&m[1136]&m[1137])|(m[1097]&~m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1097]&m[1133]&~m[1134]&m[1136]&m[1137])|(m[1097]&m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1097]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1097]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1097]&m[1133]&m[1134]&m[1136]&m[1137]));
    m[1140] = (((m[1102]&~m[1138]&~m[1139]&~m[1141]&~m[1142])|(~m[1102]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1102]&m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1102]&~m[1138]&m[1139]&m[1141]&~m[1142])|(~m[1102]&m[1138]&~m[1139]&~m[1141]&m[1142])|(~m[1102]&~m[1138]&m[1139]&~m[1141]&m[1142])|(m[1102]&m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1102]&m[1138]&m[1139]&m[1141]&m[1142]))&UnbiasedRNG[305])|((m[1102]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(~m[1102]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1102]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1102]&m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1102]&~m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1102]&~m[1138]&~m[1139]&m[1141]&m[1142])|(m[1102]&~m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1102]&m[1138]&~m[1139]&m[1141]&m[1142])|(m[1102]&m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1102]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1102]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1102]&m[1138]&m[1139]&m[1141]&m[1142]));
    m[1145] = (((m[1107]&~m[1143]&~m[1144]&~m[1146]&~m[1147])|(~m[1107]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1107]&m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1107]&~m[1143]&m[1144]&m[1146]&~m[1147])|(~m[1107]&m[1143]&~m[1144]&~m[1146]&m[1147])|(~m[1107]&~m[1143]&m[1144]&~m[1146]&m[1147])|(m[1107]&m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1107]&m[1143]&m[1144]&m[1146]&m[1147]))&UnbiasedRNG[306])|((m[1107]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(~m[1107]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1107]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1107]&m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1107]&~m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1107]&~m[1143]&~m[1144]&m[1146]&m[1147])|(m[1107]&~m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1107]&m[1143]&~m[1144]&m[1146]&m[1147])|(m[1107]&m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1107]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1107]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1107]&m[1143]&m[1144]&m[1146]&m[1147]));
    m[1155] = (((m[1112]&~m[1153]&~m[1154]&~m[1156]&~m[1157])|(~m[1112]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1112]&m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1112]&~m[1153]&m[1154]&m[1156]&~m[1157])|(~m[1112]&m[1153]&~m[1154]&~m[1156]&m[1157])|(~m[1112]&~m[1153]&m[1154]&~m[1156]&m[1157])|(m[1112]&m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1112]&m[1153]&m[1154]&m[1156]&m[1157]))&UnbiasedRNG[307])|((m[1112]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(~m[1112]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1112]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1112]&m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1112]&~m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1112]&~m[1153]&~m[1154]&m[1156]&m[1157])|(m[1112]&~m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1112]&m[1153]&~m[1154]&m[1156]&m[1157])|(m[1112]&m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1112]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1112]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1112]&m[1153]&m[1154]&m[1156]&m[1157]));
    m[1160] = (((m[1117]&~m[1158]&~m[1159]&~m[1161]&~m[1162])|(~m[1117]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1117]&m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1117]&~m[1158]&m[1159]&m[1161]&~m[1162])|(~m[1117]&m[1158]&~m[1159]&~m[1161]&m[1162])|(~m[1117]&~m[1158]&m[1159]&~m[1161]&m[1162])|(m[1117]&m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1117]&m[1158]&m[1159]&m[1161]&m[1162]))&UnbiasedRNG[308])|((m[1117]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(~m[1117]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1117]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1117]&m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1117]&~m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1117]&~m[1158]&~m[1159]&m[1161]&m[1162])|(m[1117]&~m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1117]&m[1158]&~m[1159]&m[1161]&m[1162])|(m[1117]&m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1117]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1117]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1117]&m[1158]&m[1159]&m[1161]&m[1162]));
    m[1165] = (((m[1122]&~m[1163]&~m[1164]&~m[1166]&~m[1167])|(~m[1122]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1122]&m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1122]&~m[1163]&m[1164]&m[1166]&~m[1167])|(~m[1122]&m[1163]&~m[1164]&~m[1166]&m[1167])|(~m[1122]&~m[1163]&m[1164]&~m[1166]&m[1167])|(m[1122]&m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1122]&m[1163]&m[1164]&m[1166]&m[1167]))&UnbiasedRNG[309])|((m[1122]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(~m[1122]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1122]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1122]&m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1122]&~m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1122]&~m[1163]&~m[1164]&m[1166]&m[1167])|(m[1122]&~m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1122]&m[1163]&~m[1164]&m[1166]&m[1167])|(m[1122]&m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1122]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1122]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1122]&m[1163]&m[1164]&m[1166]&m[1167]));
    m[1170] = (((m[1127]&~m[1168]&~m[1169]&~m[1171]&~m[1172])|(~m[1127]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1127]&m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1127]&~m[1168]&m[1169]&m[1171]&~m[1172])|(~m[1127]&m[1168]&~m[1169]&~m[1171]&m[1172])|(~m[1127]&~m[1168]&m[1169]&~m[1171]&m[1172])|(m[1127]&m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1127]&m[1168]&m[1169]&m[1171]&m[1172]))&UnbiasedRNG[310])|((m[1127]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(~m[1127]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1127]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1127]&m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1127]&~m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1127]&~m[1168]&~m[1169]&m[1171]&m[1172])|(m[1127]&~m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1127]&m[1168]&~m[1169]&m[1171]&m[1172])|(m[1127]&m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1127]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1127]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1127]&m[1168]&m[1169]&m[1171]&m[1172]));
    m[1175] = (((m[1132]&~m[1173]&~m[1174]&~m[1176]&~m[1177])|(~m[1132]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1132]&m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1132]&~m[1173]&m[1174]&m[1176]&~m[1177])|(~m[1132]&m[1173]&~m[1174]&~m[1176]&m[1177])|(~m[1132]&~m[1173]&m[1174]&~m[1176]&m[1177])|(m[1132]&m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1132]&m[1173]&m[1174]&m[1176]&m[1177]))&UnbiasedRNG[311])|((m[1132]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(~m[1132]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1132]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1132]&m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1132]&~m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1132]&~m[1173]&~m[1174]&m[1176]&m[1177])|(m[1132]&~m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1132]&m[1173]&~m[1174]&m[1176]&m[1177])|(m[1132]&m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1132]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1132]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1132]&m[1173]&m[1174]&m[1176]&m[1177]));
    m[1180] = (((m[1137]&~m[1178]&~m[1179]&~m[1181]&~m[1182])|(~m[1137]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1137]&m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1137]&~m[1178]&m[1179]&m[1181]&~m[1182])|(~m[1137]&m[1178]&~m[1179]&~m[1181]&m[1182])|(~m[1137]&~m[1178]&m[1179]&~m[1181]&m[1182])|(m[1137]&m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1137]&m[1178]&m[1179]&m[1181]&m[1182]))&UnbiasedRNG[312])|((m[1137]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(~m[1137]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1137]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1137]&m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1137]&~m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1137]&~m[1178]&~m[1179]&m[1181]&m[1182])|(m[1137]&~m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1137]&m[1178]&~m[1179]&m[1181]&m[1182])|(m[1137]&m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1137]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1137]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1137]&m[1178]&m[1179]&m[1181]&m[1182]));
    m[1185] = (((m[1142]&~m[1183]&~m[1184]&~m[1186]&~m[1187])|(~m[1142]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1142]&m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1142]&~m[1183]&m[1184]&m[1186]&~m[1187])|(~m[1142]&m[1183]&~m[1184]&~m[1186]&m[1187])|(~m[1142]&~m[1183]&m[1184]&~m[1186]&m[1187])|(m[1142]&m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1142]&m[1183]&m[1184]&m[1186]&m[1187]))&UnbiasedRNG[313])|((m[1142]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(~m[1142]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1142]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1142]&m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1142]&~m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1142]&~m[1183]&~m[1184]&m[1186]&m[1187])|(m[1142]&~m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1142]&m[1183]&~m[1184]&m[1186]&m[1187])|(m[1142]&m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1142]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1142]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1142]&m[1183]&m[1184]&m[1186]&m[1187]));
    m[1190] = (((m[1147]&~m[1188]&~m[1189]&~m[1191]&~m[1192])|(~m[1147]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1147]&m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1147]&~m[1188]&m[1189]&m[1191]&~m[1192])|(~m[1147]&m[1188]&~m[1189]&~m[1191]&m[1192])|(~m[1147]&~m[1188]&m[1189]&~m[1191]&m[1192])|(m[1147]&m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1147]&m[1188]&m[1189]&m[1191]&m[1192]))&UnbiasedRNG[314])|((m[1147]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(~m[1147]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1147]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1147]&m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1147]&~m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1147]&~m[1188]&~m[1189]&m[1191]&m[1192])|(m[1147]&~m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1147]&m[1188]&~m[1189]&m[1191]&m[1192])|(m[1147]&m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1147]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1147]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1147]&m[1188]&m[1189]&m[1191]&m[1192]));
    m[1195] = (((m[1152]&~m[1193]&~m[1194]&~m[1196]&~m[1197])|(~m[1152]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1152]&m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1152]&~m[1193]&m[1194]&m[1196]&~m[1197])|(~m[1152]&m[1193]&~m[1194]&~m[1196]&m[1197])|(~m[1152]&~m[1193]&m[1194]&~m[1196]&m[1197])|(m[1152]&m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1152]&m[1193]&m[1194]&m[1196]&m[1197]))&UnbiasedRNG[315])|((m[1152]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(~m[1152]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1152]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1152]&m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1152]&~m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1152]&~m[1193]&~m[1194]&m[1196]&m[1197])|(m[1152]&~m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1152]&m[1193]&~m[1194]&m[1196]&m[1197])|(m[1152]&m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1152]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1152]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1152]&m[1193]&m[1194]&m[1196]&m[1197]));
    m[1205] = (((m[1157]&~m[1203]&~m[1204]&~m[1206]&~m[1207])|(~m[1157]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1157]&m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1157]&~m[1203]&m[1204]&m[1206]&~m[1207])|(~m[1157]&m[1203]&~m[1204]&~m[1206]&m[1207])|(~m[1157]&~m[1203]&m[1204]&~m[1206]&m[1207])|(m[1157]&m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1157]&m[1203]&m[1204]&m[1206]&m[1207]))&UnbiasedRNG[316])|((m[1157]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(~m[1157]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1157]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1157]&m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1157]&~m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1157]&~m[1203]&~m[1204]&m[1206]&m[1207])|(m[1157]&~m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1157]&m[1203]&~m[1204]&m[1206]&m[1207])|(m[1157]&m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1157]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1157]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1157]&m[1203]&m[1204]&m[1206]&m[1207]));
    m[1210] = (((m[1162]&~m[1208]&~m[1209]&~m[1211]&~m[1212])|(~m[1162]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1162]&m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1162]&~m[1208]&m[1209]&m[1211]&~m[1212])|(~m[1162]&m[1208]&~m[1209]&~m[1211]&m[1212])|(~m[1162]&~m[1208]&m[1209]&~m[1211]&m[1212])|(m[1162]&m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1162]&m[1208]&m[1209]&m[1211]&m[1212]))&UnbiasedRNG[317])|((m[1162]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(~m[1162]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1162]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1162]&m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1162]&~m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1162]&~m[1208]&~m[1209]&m[1211]&m[1212])|(m[1162]&~m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1162]&m[1208]&~m[1209]&m[1211]&m[1212])|(m[1162]&m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1162]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1162]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1162]&m[1208]&m[1209]&m[1211]&m[1212]));
    m[1215] = (((m[1167]&~m[1213]&~m[1214]&~m[1216]&~m[1217])|(~m[1167]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1167]&m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1167]&~m[1213]&m[1214]&m[1216]&~m[1217])|(~m[1167]&m[1213]&~m[1214]&~m[1216]&m[1217])|(~m[1167]&~m[1213]&m[1214]&~m[1216]&m[1217])|(m[1167]&m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1167]&m[1213]&m[1214]&m[1216]&m[1217]))&UnbiasedRNG[318])|((m[1167]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(~m[1167]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1167]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1167]&m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1167]&~m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1167]&~m[1213]&~m[1214]&m[1216]&m[1217])|(m[1167]&~m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1167]&m[1213]&~m[1214]&m[1216]&m[1217])|(m[1167]&m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1167]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1167]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1167]&m[1213]&m[1214]&m[1216]&m[1217]));
    m[1220] = (((m[1172]&~m[1218]&~m[1219]&~m[1221]&~m[1222])|(~m[1172]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1172]&m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1172]&~m[1218]&m[1219]&m[1221]&~m[1222])|(~m[1172]&m[1218]&~m[1219]&~m[1221]&m[1222])|(~m[1172]&~m[1218]&m[1219]&~m[1221]&m[1222])|(m[1172]&m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1172]&m[1218]&m[1219]&m[1221]&m[1222]))&UnbiasedRNG[319])|((m[1172]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(~m[1172]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1172]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1172]&m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1172]&~m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1172]&~m[1218]&~m[1219]&m[1221]&m[1222])|(m[1172]&~m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1172]&m[1218]&~m[1219]&m[1221]&m[1222])|(m[1172]&m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1172]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1172]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1172]&m[1218]&m[1219]&m[1221]&m[1222]));
    m[1225] = (((m[1177]&~m[1223]&~m[1224]&~m[1226]&~m[1227])|(~m[1177]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1177]&m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1177]&~m[1223]&m[1224]&m[1226]&~m[1227])|(~m[1177]&m[1223]&~m[1224]&~m[1226]&m[1227])|(~m[1177]&~m[1223]&m[1224]&~m[1226]&m[1227])|(m[1177]&m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1177]&m[1223]&m[1224]&m[1226]&m[1227]))&UnbiasedRNG[320])|((m[1177]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(~m[1177]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1177]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1177]&m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1177]&~m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1177]&~m[1223]&~m[1224]&m[1226]&m[1227])|(m[1177]&~m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1177]&m[1223]&~m[1224]&m[1226]&m[1227])|(m[1177]&m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1177]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1177]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1177]&m[1223]&m[1224]&m[1226]&m[1227]));
    m[1230] = (((m[1182]&~m[1228]&~m[1229]&~m[1231]&~m[1232])|(~m[1182]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1182]&m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1182]&~m[1228]&m[1229]&m[1231]&~m[1232])|(~m[1182]&m[1228]&~m[1229]&~m[1231]&m[1232])|(~m[1182]&~m[1228]&m[1229]&~m[1231]&m[1232])|(m[1182]&m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1182]&m[1228]&m[1229]&m[1231]&m[1232]))&UnbiasedRNG[321])|((m[1182]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(~m[1182]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1182]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1182]&m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1182]&~m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1182]&~m[1228]&~m[1229]&m[1231]&m[1232])|(m[1182]&~m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1182]&m[1228]&~m[1229]&m[1231]&m[1232])|(m[1182]&m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1182]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1182]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1182]&m[1228]&m[1229]&m[1231]&m[1232]));
    m[1235] = (((m[1187]&~m[1233]&~m[1234]&~m[1236]&~m[1237])|(~m[1187]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1187]&m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1187]&~m[1233]&m[1234]&m[1236]&~m[1237])|(~m[1187]&m[1233]&~m[1234]&~m[1236]&m[1237])|(~m[1187]&~m[1233]&m[1234]&~m[1236]&m[1237])|(m[1187]&m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1187]&m[1233]&m[1234]&m[1236]&m[1237]))&UnbiasedRNG[322])|((m[1187]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(~m[1187]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1187]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1187]&m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1187]&~m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1187]&~m[1233]&~m[1234]&m[1236]&m[1237])|(m[1187]&~m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1187]&m[1233]&~m[1234]&m[1236]&m[1237])|(m[1187]&m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1187]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1187]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1187]&m[1233]&m[1234]&m[1236]&m[1237]));
    m[1240] = (((m[1192]&~m[1238]&~m[1239]&~m[1241]&~m[1242])|(~m[1192]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1192]&m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1192]&~m[1238]&m[1239]&m[1241]&~m[1242])|(~m[1192]&m[1238]&~m[1239]&~m[1241]&m[1242])|(~m[1192]&~m[1238]&m[1239]&~m[1241]&m[1242])|(m[1192]&m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1192]&m[1238]&m[1239]&m[1241]&m[1242]))&UnbiasedRNG[323])|((m[1192]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(~m[1192]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1192]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1192]&m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1192]&~m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1192]&~m[1238]&~m[1239]&m[1241]&m[1242])|(m[1192]&~m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1192]&m[1238]&~m[1239]&m[1241]&m[1242])|(m[1192]&m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1192]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1192]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1192]&m[1238]&m[1239]&m[1241]&m[1242]));
    m[1245] = (((m[1197]&~m[1243]&~m[1244]&~m[1246]&~m[1247])|(~m[1197]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1197]&m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1197]&~m[1243]&m[1244]&m[1246]&~m[1247])|(~m[1197]&m[1243]&~m[1244]&~m[1246]&m[1247])|(~m[1197]&~m[1243]&m[1244]&~m[1246]&m[1247])|(m[1197]&m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1197]&m[1243]&m[1244]&m[1246]&m[1247]))&UnbiasedRNG[324])|((m[1197]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(~m[1197]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1197]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1197]&m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1197]&~m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1197]&~m[1243]&~m[1244]&m[1246]&m[1247])|(m[1197]&~m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1197]&m[1243]&~m[1244]&m[1246]&m[1247])|(m[1197]&m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1197]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1197]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1197]&m[1243]&m[1244]&m[1246]&m[1247]));
    m[1250] = (((m[1202]&~m[1248]&~m[1249]&~m[1251]&~m[1252])|(~m[1202]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1202]&m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1202]&~m[1248]&m[1249]&m[1251]&~m[1252])|(~m[1202]&m[1248]&~m[1249]&~m[1251]&m[1252])|(~m[1202]&~m[1248]&m[1249]&~m[1251]&m[1252])|(m[1202]&m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1202]&m[1248]&m[1249]&m[1251]&m[1252]))&UnbiasedRNG[325])|((m[1202]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(~m[1202]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1202]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1202]&m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1202]&~m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1202]&~m[1248]&~m[1249]&m[1251]&m[1252])|(m[1202]&~m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1202]&m[1248]&~m[1249]&m[1251]&m[1252])|(m[1202]&m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1202]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1202]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1202]&m[1248]&m[1249]&m[1251]&m[1252]));
    m[1260] = (((m[1207]&~m[1258]&~m[1259]&~m[1261]&~m[1262])|(~m[1207]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1207]&m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1207]&~m[1258]&m[1259]&m[1261]&~m[1262])|(~m[1207]&m[1258]&~m[1259]&~m[1261]&m[1262])|(~m[1207]&~m[1258]&m[1259]&~m[1261]&m[1262])|(m[1207]&m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1207]&m[1258]&m[1259]&m[1261]&m[1262]))&UnbiasedRNG[326])|((m[1207]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(~m[1207]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1207]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1207]&m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1207]&~m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1207]&~m[1258]&~m[1259]&m[1261]&m[1262])|(m[1207]&~m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1207]&m[1258]&~m[1259]&m[1261]&m[1262])|(m[1207]&m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1207]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1207]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1207]&m[1258]&m[1259]&m[1261]&m[1262]));
    m[1265] = (((m[1212]&~m[1263]&~m[1264]&~m[1266]&~m[1267])|(~m[1212]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1212]&m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1212]&~m[1263]&m[1264]&m[1266]&~m[1267])|(~m[1212]&m[1263]&~m[1264]&~m[1266]&m[1267])|(~m[1212]&~m[1263]&m[1264]&~m[1266]&m[1267])|(m[1212]&m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1212]&m[1263]&m[1264]&m[1266]&m[1267]))&UnbiasedRNG[327])|((m[1212]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(~m[1212]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1212]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1212]&m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1212]&~m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1212]&~m[1263]&~m[1264]&m[1266]&m[1267])|(m[1212]&~m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1212]&m[1263]&~m[1264]&m[1266]&m[1267])|(m[1212]&m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1212]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1212]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1212]&m[1263]&m[1264]&m[1266]&m[1267]));
    m[1270] = (((m[1217]&~m[1268]&~m[1269]&~m[1271]&~m[1272])|(~m[1217]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1217]&m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1217]&~m[1268]&m[1269]&m[1271]&~m[1272])|(~m[1217]&m[1268]&~m[1269]&~m[1271]&m[1272])|(~m[1217]&~m[1268]&m[1269]&~m[1271]&m[1272])|(m[1217]&m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1217]&m[1268]&m[1269]&m[1271]&m[1272]))&UnbiasedRNG[328])|((m[1217]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(~m[1217]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1217]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1217]&m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1217]&~m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1217]&~m[1268]&~m[1269]&m[1271]&m[1272])|(m[1217]&~m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1217]&m[1268]&~m[1269]&m[1271]&m[1272])|(m[1217]&m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1217]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1217]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1217]&m[1268]&m[1269]&m[1271]&m[1272]));
    m[1275] = (((m[1222]&~m[1273]&~m[1274]&~m[1276]&~m[1277])|(~m[1222]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1222]&m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1222]&~m[1273]&m[1274]&m[1276]&~m[1277])|(~m[1222]&m[1273]&~m[1274]&~m[1276]&m[1277])|(~m[1222]&~m[1273]&m[1274]&~m[1276]&m[1277])|(m[1222]&m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1222]&m[1273]&m[1274]&m[1276]&m[1277]))&UnbiasedRNG[329])|((m[1222]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(~m[1222]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1222]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1222]&m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1222]&~m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1222]&~m[1273]&~m[1274]&m[1276]&m[1277])|(m[1222]&~m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1222]&m[1273]&~m[1274]&m[1276]&m[1277])|(m[1222]&m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1222]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1222]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1222]&m[1273]&m[1274]&m[1276]&m[1277]));
    m[1280] = (((m[1227]&~m[1278]&~m[1279]&~m[1281]&~m[1282])|(~m[1227]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1227]&m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1227]&~m[1278]&m[1279]&m[1281]&~m[1282])|(~m[1227]&m[1278]&~m[1279]&~m[1281]&m[1282])|(~m[1227]&~m[1278]&m[1279]&~m[1281]&m[1282])|(m[1227]&m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1227]&m[1278]&m[1279]&m[1281]&m[1282]))&UnbiasedRNG[330])|((m[1227]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(~m[1227]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1227]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1227]&m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1227]&~m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1227]&~m[1278]&~m[1279]&m[1281]&m[1282])|(m[1227]&~m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1227]&m[1278]&~m[1279]&m[1281]&m[1282])|(m[1227]&m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1227]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1227]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1227]&m[1278]&m[1279]&m[1281]&m[1282]));
    m[1285] = (((m[1232]&~m[1283]&~m[1284]&~m[1286]&~m[1287])|(~m[1232]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1232]&m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1232]&~m[1283]&m[1284]&m[1286]&~m[1287])|(~m[1232]&m[1283]&~m[1284]&~m[1286]&m[1287])|(~m[1232]&~m[1283]&m[1284]&~m[1286]&m[1287])|(m[1232]&m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1232]&m[1283]&m[1284]&m[1286]&m[1287]))&UnbiasedRNG[331])|((m[1232]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(~m[1232]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1232]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1232]&m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1232]&~m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1232]&~m[1283]&~m[1284]&m[1286]&m[1287])|(m[1232]&~m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1232]&m[1283]&~m[1284]&m[1286]&m[1287])|(m[1232]&m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1232]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1232]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1232]&m[1283]&m[1284]&m[1286]&m[1287]));
    m[1290] = (((m[1237]&~m[1288]&~m[1289]&~m[1291]&~m[1292])|(~m[1237]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1237]&m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1237]&~m[1288]&m[1289]&m[1291]&~m[1292])|(~m[1237]&m[1288]&~m[1289]&~m[1291]&m[1292])|(~m[1237]&~m[1288]&m[1289]&~m[1291]&m[1292])|(m[1237]&m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1237]&m[1288]&m[1289]&m[1291]&m[1292]))&UnbiasedRNG[332])|((m[1237]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(~m[1237]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1237]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1237]&m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1237]&~m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1237]&~m[1288]&~m[1289]&m[1291]&m[1292])|(m[1237]&~m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1237]&m[1288]&~m[1289]&m[1291]&m[1292])|(m[1237]&m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1237]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1237]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1237]&m[1288]&m[1289]&m[1291]&m[1292]));
    m[1295] = (((m[1242]&~m[1293]&~m[1294]&~m[1296]&~m[1297])|(~m[1242]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1242]&m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1242]&~m[1293]&m[1294]&m[1296]&~m[1297])|(~m[1242]&m[1293]&~m[1294]&~m[1296]&m[1297])|(~m[1242]&~m[1293]&m[1294]&~m[1296]&m[1297])|(m[1242]&m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1242]&m[1293]&m[1294]&m[1296]&m[1297]))&UnbiasedRNG[333])|((m[1242]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(~m[1242]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1242]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1242]&m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1242]&~m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1242]&~m[1293]&~m[1294]&m[1296]&m[1297])|(m[1242]&~m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1242]&m[1293]&~m[1294]&m[1296]&m[1297])|(m[1242]&m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1242]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1242]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1242]&m[1293]&m[1294]&m[1296]&m[1297]));
    m[1300] = (((m[1247]&~m[1298]&~m[1299]&~m[1301]&~m[1302])|(~m[1247]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1247]&m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1247]&~m[1298]&m[1299]&m[1301]&~m[1302])|(~m[1247]&m[1298]&~m[1299]&~m[1301]&m[1302])|(~m[1247]&~m[1298]&m[1299]&~m[1301]&m[1302])|(m[1247]&m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1247]&m[1298]&m[1299]&m[1301]&m[1302]))&UnbiasedRNG[334])|((m[1247]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(~m[1247]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1247]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1247]&m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1247]&~m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1247]&~m[1298]&~m[1299]&m[1301]&m[1302])|(m[1247]&~m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1247]&m[1298]&~m[1299]&m[1301]&m[1302])|(m[1247]&m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1247]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1247]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1247]&m[1298]&m[1299]&m[1301]&m[1302]));
    m[1305] = (((m[1252]&~m[1303]&~m[1304]&~m[1306]&~m[1307])|(~m[1252]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1252]&m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1252]&~m[1303]&m[1304]&m[1306]&~m[1307])|(~m[1252]&m[1303]&~m[1304]&~m[1306]&m[1307])|(~m[1252]&~m[1303]&m[1304]&~m[1306]&m[1307])|(m[1252]&m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1252]&m[1303]&m[1304]&m[1306]&m[1307]))&UnbiasedRNG[335])|((m[1252]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(~m[1252]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1252]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1252]&m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1252]&~m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1252]&~m[1303]&~m[1304]&m[1306]&m[1307])|(m[1252]&~m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1252]&m[1303]&~m[1304]&m[1306]&m[1307])|(m[1252]&m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1252]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1252]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1252]&m[1303]&m[1304]&m[1306]&m[1307]));
    m[1310] = (((m[1257]&~m[1308]&~m[1309]&~m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&~m[1312])|(~m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&m[1308]&m[1309]&m[1311]&m[1312]))&UnbiasedRNG[336])|((m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&m[1311]&m[1312]));
    m[1320] = (((m[1262]&~m[1318]&~m[1319]&~m[1321]&~m[1322])|(~m[1262]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1262]&m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1262]&~m[1318]&m[1319]&m[1321]&~m[1322])|(~m[1262]&m[1318]&~m[1319]&~m[1321]&m[1322])|(~m[1262]&~m[1318]&m[1319]&~m[1321]&m[1322])|(m[1262]&m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1262]&m[1318]&m[1319]&m[1321]&m[1322]))&UnbiasedRNG[337])|((m[1262]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(~m[1262]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1262]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1262]&m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1262]&~m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1262]&~m[1318]&~m[1319]&m[1321]&m[1322])|(m[1262]&~m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1262]&m[1318]&~m[1319]&m[1321]&m[1322])|(m[1262]&m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1262]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1262]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1262]&m[1318]&m[1319]&m[1321]&m[1322]));
    m[1325] = (((m[1267]&~m[1323]&~m[1324]&~m[1326]&~m[1327])|(~m[1267]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1267]&m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1267]&~m[1323]&m[1324]&m[1326]&~m[1327])|(~m[1267]&m[1323]&~m[1324]&~m[1326]&m[1327])|(~m[1267]&~m[1323]&m[1324]&~m[1326]&m[1327])|(m[1267]&m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1267]&m[1323]&m[1324]&m[1326]&m[1327]))&UnbiasedRNG[338])|((m[1267]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(~m[1267]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1267]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1267]&m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1267]&~m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1267]&~m[1323]&~m[1324]&m[1326]&m[1327])|(m[1267]&~m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1267]&m[1323]&~m[1324]&m[1326]&m[1327])|(m[1267]&m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1267]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1267]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1267]&m[1323]&m[1324]&m[1326]&m[1327]));
    m[1330] = (((m[1272]&~m[1328]&~m[1329]&~m[1331]&~m[1332])|(~m[1272]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1272]&m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1272]&~m[1328]&m[1329]&m[1331]&~m[1332])|(~m[1272]&m[1328]&~m[1329]&~m[1331]&m[1332])|(~m[1272]&~m[1328]&m[1329]&~m[1331]&m[1332])|(m[1272]&m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1272]&m[1328]&m[1329]&m[1331]&m[1332]))&UnbiasedRNG[339])|((m[1272]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(~m[1272]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1272]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1272]&m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1272]&~m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1272]&~m[1328]&~m[1329]&m[1331]&m[1332])|(m[1272]&~m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1272]&m[1328]&~m[1329]&m[1331]&m[1332])|(m[1272]&m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1272]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1272]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1272]&m[1328]&m[1329]&m[1331]&m[1332]));
    m[1335] = (((m[1277]&~m[1333]&~m[1334]&~m[1336]&~m[1337])|(~m[1277]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1277]&m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1277]&~m[1333]&m[1334]&m[1336]&~m[1337])|(~m[1277]&m[1333]&~m[1334]&~m[1336]&m[1337])|(~m[1277]&~m[1333]&m[1334]&~m[1336]&m[1337])|(m[1277]&m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1277]&m[1333]&m[1334]&m[1336]&m[1337]))&UnbiasedRNG[340])|((m[1277]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(~m[1277]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1277]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1277]&m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1277]&~m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1277]&~m[1333]&~m[1334]&m[1336]&m[1337])|(m[1277]&~m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1277]&m[1333]&~m[1334]&m[1336]&m[1337])|(m[1277]&m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1277]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1277]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1277]&m[1333]&m[1334]&m[1336]&m[1337]));
    m[1340] = (((m[1282]&~m[1338]&~m[1339]&~m[1341]&~m[1342])|(~m[1282]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1282]&m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1282]&~m[1338]&m[1339]&m[1341]&~m[1342])|(~m[1282]&m[1338]&~m[1339]&~m[1341]&m[1342])|(~m[1282]&~m[1338]&m[1339]&~m[1341]&m[1342])|(m[1282]&m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1282]&m[1338]&m[1339]&m[1341]&m[1342]))&UnbiasedRNG[341])|((m[1282]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(~m[1282]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1282]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1282]&m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1282]&~m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1282]&~m[1338]&~m[1339]&m[1341]&m[1342])|(m[1282]&~m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1282]&m[1338]&~m[1339]&m[1341]&m[1342])|(m[1282]&m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1282]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1282]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1282]&m[1338]&m[1339]&m[1341]&m[1342]));
    m[1345] = (((m[1287]&~m[1343]&~m[1344]&~m[1346]&~m[1347])|(~m[1287]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1287]&m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1287]&~m[1343]&m[1344]&m[1346]&~m[1347])|(~m[1287]&m[1343]&~m[1344]&~m[1346]&m[1347])|(~m[1287]&~m[1343]&m[1344]&~m[1346]&m[1347])|(m[1287]&m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1287]&m[1343]&m[1344]&m[1346]&m[1347]))&UnbiasedRNG[342])|((m[1287]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(~m[1287]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1287]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1287]&m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1287]&~m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1287]&~m[1343]&~m[1344]&m[1346]&m[1347])|(m[1287]&~m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1287]&m[1343]&~m[1344]&m[1346]&m[1347])|(m[1287]&m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1287]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1287]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1287]&m[1343]&m[1344]&m[1346]&m[1347]));
    m[1350] = (((m[1292]&~m[1348]&~m[1349]&~m[1351]&~m[1352])|(~m[1292]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1292]&m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1292]&~m[1348]&m[1349]&m[1351]&~m[1352])|(~m[1292]&m[1348]&~m[1349]&~m[1351]&m[1352])|(~m[1292]&~m[1348]&m[1349]&~m[1351]&m[1352])|(m[1292]&m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1292]&m[1348]&m[1349]&m[1351]&m[1352]))&UnbiasedRNG[343])|((m[1292]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(~m[1292]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1292]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1292]&m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1292]&~m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1292]&~m[1348]&~m[1349]&m[1351]&m[1352])|(m[1292]&~m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1292]&m[1348]&~m[1349]&m[1351]&m[1352])|(m[1292]&m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1292]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1292]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1292]&m[1348]&m[1349]&m[1351]&m[1352]));
    m[1355] = (((m[1297]&~m[1353]&~m[1354]&~m[1356]&~m[1357])|(~m[1297]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1297]&m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1297]&~m[1353]&m[1354]&m[1356]&~m[1357])|(~m[1297]&m[1353]&~m[1354]&~m[1356]&m[1357])|(~m[1297]&~m[1353]&m[1354]&~m[1356]&m[1357])|(m[1297]&m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1297]&m[1353]&m[1354]&m[1356]&m[1357]))&UnbiasedRNG[344])|((m[1297]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(~m[1297]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1297]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1297]&m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1297]&~m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1297]&~m[1353]&~m[1354]&m[1356]&m[1357])|(m[1297]&~m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1297]&m[1353]&~m[1354]&m[1356]&m[1357])|(m[1297]&m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1297]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1297]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1297]&m[1353]&m[1354]&m[1356]&m[1357]));
    m[1360] = (((m[1302]&~m[1358]&~m[1359]&~m[1361]&~m[1362])|(~m[1302]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1302]&m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1302]&~m[1358]&m[1359]&m[1361]&~m[1362])|(~m[1302]&m[1358]&~m[1359]&~m[1361]&m[1362])|(~m[1302]&~m[1358]&m[1359]&~m[1361]&m[1362])|(m[1302]&m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1302]&m[1358]&m[1359]&m[1361]&m[1362]))&UnbiasedRNG[345])|((m[1302]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(~m[1302]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1302]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1302]&m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1302]&~m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1302]&~m[1358]&~m[1359]&m[1361]&m[1362])|(m[1302]&~m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1302]&m[1358]&~m[1359]&m[1361]&m[1362])|(m[1302]&m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1302]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1302]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1302]&m[1358]&m[1359]&m[1361]&m[1362]));
    m[1365] = (((m[1307]&~m[1363]&~m[1364]&~m[1366]&~m[1367])|(~m[1307]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1307]&m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1307]&~m[1363]&m[1364]&m[1366]&~m[1367])|(~m[1307]&m[1363]&~m[1364]&~m[1366]&m[1367])|(~m[1307]&~m[1363]&m[1364]&~m[1366]&m[1367])|(m[1307]&m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1307]&m[1363]&m[1364]&m[1366]&m[1367]))&UnbiasedRNG[346])|((m[1307]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(~m[1307]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1307]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1307]&m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1307]&~m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1307]&~m[1363]&~m[1364]&m[1366]&m[1367])|(m[1307]&~m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1307]&m[1363]&~m[1364]&m[1366]&m[1367])|(m[1307]&m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1307]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1307]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1307]&m[1363]&m[1364]&m[1366]&m[1367]));
    m[1370] = (((m[1312]&~m[1368]&~m[1369]&~m[1371]&~m[1372])|(~m[1312]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1312]&m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1312]&~m[1368]&m[1369]&m[1371]&~m[1372])|(~m[1312]&m[1368]&~m[1369]&~m[1371]&m[1372])|(~m[1312]&~m[1368]&m[1369]&~m[1371]&m[1372])|(m[1312]&m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1312]&m[1368]&m[1369]&m[1371]&m[1372]))&UnbiasedRNG[347])|((m[1312]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(~m[1312]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1312]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1312]&m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1312]&~m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1312]&~m[1368]&~m[1369]&m[1371]&m[1372])|(m[1312]&~m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1312]&m[1368]&~m[1369]&m[1371]&m[1372])|(m[1312]&m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1312]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1312]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1312]&m[1368]&m[1369]&m[1371]&m[1372]));
    m[1375] = (((m[1317]&~m[1373]&~m[1374]&~m[1376]&~m[1377])|(~m[1317]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1317]&m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1317]&~m[1373]&m[1374]&m[1376]&~m[1377])|(~m[1317]&m[1373]&~m[1374]&~m[1376]&m[1377])|(~m[1317]&~m[1373]&m[1374]&~m[1376]&m[1377])|(m[1317]&m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1317]&m[1373]&m[1374]&m[1376]&m[1377]))&UnbiasedRNG[348])|((m[1317]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(~m[1317]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1317]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1317]&m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1317]&~m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1317]&~m[1373]&~m[1374]&m[1376]&m[1377])|(m[1317]&~m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1317]&m[1373]&~m[1374]&m[1376]&m[1377])|(m[1317]&m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1317]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1317]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1317]&m[1373]&m[1374]&m[1376]&m[1377]));
    m[1385] = (((m[1322]&~m[1383]&~m[1384]&~m[1386]&~m[1387])|(~m[1322]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1322]&m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1322]&~m[1383]&m[1384]&m[1386]&~m[1387])|(~m[1322]&m[1383]&~m[1384]&~m[1386]&m[1387])|(~m[1322]&~m[1383]&m[1384]&~m[1386]&m[1387])|(m[1322]&m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1322]&m[1383]&m[1384]&m[1386]&m[1387]))&UnbiasedRNG[349])|((m[1322]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(~m[1322]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1322]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1322]&m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1322]&~m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1322]&~m[1383]&~m[1384]&m[1386]&m[1387])|(m[1322]&~m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1322]&m[1383]&~m[1384]&m[1386]&m[1387])|(m[1322]&m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1322]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1322]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1322]&m[1383]&m[1384]&m[1386]&m[1387]));
    m[1390] = (((m[1327]&~m[1388]&~m[1389]&~m[1391]&~m[1392])|(~m[1327]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1327]&m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1327]&~m[1388]&m[1389]&m[1391]&~m[1392])|(~m[1327]&m[1388]&~m[1389]&~m[1391]&m[1392])|(~m[1327]&~m[1388]&m[1389]&~m[1391]&m[1392])|(m[1327]&m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1327]&m[1388]&m[1389]&m[1391]&m[1392]))&UnbiasedRNG[350])|((m[1327]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(~m[1327]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1327]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1327]&m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1327]&~m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1327]&~m[1388]&~m[1389]&m[1391]&m[1392])|(m[1327]&~m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1327]&m[1388]&~m[1389]&m[1391]&m[1392])|(m[1327]&m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1327]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1327]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1327]&m[1388]&m[1389]&m[1391]&m[1392]));
    m[1395] = (((m[1332]&~m[1393]&~m[1394]&~m[1396]&~m[1397])|(~m[1332]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1332]&m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1332]&~m[1393]&m[1394]&m[1396]&~m[1397])|(~m[1332]&m[1393]&~m[1394]&~m[1396]&m[1397])|(~m[1332]&~m[1393]&m[1394]&~m[1396]&m[1397])|(m[1332]&m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1332]&m[1393]&m[1394]&m[1396]&m[1397]))&UnbiasedRNG[351])|((m[1332]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(~m[1332]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1332]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1332]&m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1332]&~m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1332]&~m[1393]&~m[1394]&m[1396]&m[1397])|(m[1332]&~m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1332]&m[1393]&~m[1394]&m[1396]&m[1397])|(m[1332]&m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1332]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1332]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1332]&m[1393]&m[1394]&m[1396]&m[1397]));
    m[1400] = (((m[1337]&~m[1398]&~m[1399]&~m[1401]&~m[1402])|(~m[1337]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1337]&m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1337]&~m[1398]&m[1399]&m[1401]&~m[1402])|(~m[1337]&m[1398]&~m[1399]&~m[1401]&m[1402])|(~m[1337]&~m[1398]&m[1399]&~m[1401]&m[1402])|(m[1337]&m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1337]&m[1398]&m[1399]&m[1401]&m[1402]))&UnbiasedRNG[352])|((m[1337]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(~m[1337]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1337]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1337]&m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1337]&~m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1337]&~m[1398]&~m[1399]&m[1401]&m[1402])|(m[1337]&~m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1337]&m[1398]&~m[1399]&m[1401]&m[1402])|(m[1337]&m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1337]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1337]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1337]&m[1398]&m[1399]&m[1401]&m[1402]));
    m[1405] = (((m[1342]&~m[1403]&~m[1404]&~m[1406]&~m[1407])|(~m[1342]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1342]&m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1342]&~m[1403]&m[1404]&m[1406]&~m[1407])|(~m[1342]&m[1403]&~m[1404]&~m[1406]&m[1407])|(~m[1342]&~m[1403]&m[1404]&~m[1406]&m[1407])|(m[1342]&m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1342]&m[1403]&m[1404]&m[1406]&m[1407]))&UnbiasedRNG[353])|((m[1342]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(~m[1342]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1342]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1342]&m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1342]&~m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1342]&~m[1403]&~m[1404]&m[1406]&m[1407])|(m[1342]&~m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1342]&m[1403]&~m[1404]&m[1406]&m[1407])|(m[1342]&m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1342]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1342]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1342]&m[1403]&m[1404]&m[1406]&m[1407]));
    m[1410] = (((m[1347]&~m[1408]&~m[1409]&~m[1411]&~m[1412])|(~m[1347]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1347]&m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1347]&~m[1408]&m[1409]&m[1411]&~m[1412])|(~m[1347]&m[1408]&~m[1409]&~m[1411]&m[1412])|(~m[1347]&~m[1408]&m[1409]&~m[1411]&m[1412])|(m[1347]&m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1347]&m[1408]&m[1409]&m[1411]&m[1412]))&UnbiasedRNG[354])|((m[1347]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(~m[1347]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1347]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1347]&m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1347]&~m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1347]&~m[1408]&~m[1409]&m[1411]&m[1412])|(m[1347]&~m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1347]&m[1408]&~m[1409]&m[1411]&m[1412])|(m[1347]&m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1347]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1347]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1347]&m[1408]&m[1409]&m[1411]&m[1412]));
    m[1415] = (((m[1352]&~m[1413]&~m[1414]&~m[1416]&~m[1417])|(~m[1352]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1352]&m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1352]&~m[1413]&m[1414]&m[1416]&~m[1417])|(~m[1352]&m[1413]&~m[1414]&~m[1416]&m[1417])|(~m[1352]&~m[1413]&m[1414]&~m[1416]&m[1417])|(m[1352]&m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1352]&m[1413]&m[1414]&m[1416]&m[1417]))&UnbiasedRNG[355])|((m[1352]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(~m[1352]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1352]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1352]&m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1352]&~m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1352]&~m[1413]&~m[1414]&m[1416]&m[1417])|(m[1352]&~m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1352]&m[1413]&~m[1414]&m[1416]&m[1417])|(m[1352]&m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1352]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1352]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1352]&m[1413]&m[1414]&m[1416]&m[1417]));
    m[1420] = (((m[1357]&~m[1418]&~m[1419]&~m[1421]&~m[1422])|(~m[1357]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1357]&m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1357]&~m[1418]&m[1419]&m[1421]&~m[1422])|(~m[1357]&m[1418]&~m[1419]&~m[1421]&m[1422])|(~m[1357]&~m[1418]&m[1419]&~m[1421]&m[1422])|(m[1357]&m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1357]&m[1418]&m[1419]&m[1421]&m[1422]))&UnbiasedRNG[356])|((m[1357]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(~m[1357]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1357]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1357]&m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1357]&~m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1357]&~m[1418]&~m[1419]&m[1421]&m[1422])|(m[1357]&~m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1357]&m[1418]&~m[1419]&m[1421]&m[1422])|(m[1357]&m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1357]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1357]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1357]&m[1418]&m[1419]&m[1421]&m[1422]));
    m[1425] = (((m[1362]&~m[1423]&~m[1424]&~m[1426]&~m[1427])|(~m[1362]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1362]&m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1362]&~m[1423]&m[1424]&m[1426]&~m[1427])|(~m[1362]&m[1423]&~m[1424]&~m[1426]&m[1427])|(~m[1362]&~m[1423]&m[1424]&~m[1426]&m[1427])|(m[1362]&m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1362]&m[1423]&m[1424]&m[1426]&m[1427]))&UnbiasedRNG[357])|((m[1362]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(~m[1362]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1362]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1362]&m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1362]&~m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1362]&~m[1423]&~m[1424]&m[1426]&m[1427])|(m[1362]&~m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1362]&m[1423]&~m[1424]&m[1426]&m[1427])|(m[1362]&m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1362]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1362]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1362]&m[1423]&m[1424]&m[1426]&m[1427]));
    m[1430] = (((m[1367]&~m[1428]&~m[1429]&~m[1431]&~m[1432])|(~m[1367]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1367]&m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1367]&~m[1428]&m[1429]&m[1431]&~m[1432])|(~m[1367]&m[1428]&~m[1429]&~m[1431]&m[1432])|(~m[1367]&~m[1428]&m[1429]&~m[1431]&m[1432])|(m[1367]&m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1367]&m[1428]&m[1429]&m[1431]&m[1432]))&UnbiasedRNG[358])|((m[1367]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(~m[1367]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1367]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1367]&m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1367]&~m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1367]&~m[1428]&~m[1429]&m[1431]&m[1432])|(m[1367]&~m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1367]&m[1428]&~m[1429]&m[1431]&m[1432])|(m[1367]&m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1367]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1367]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1367]&m[1428]&m[1429]&m[1431]&m[1432]));
    m[1435] = (((m[1372]&~m[1433]&~m[1434]&~m[1436]&~m[1437])|(~m[1372]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1372]&m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1372]&~m[1433]&m[1434]&m[1436]&~m[1437])|(~m[1372]&m[1433]&~m[1434]&~m[1436]&m[1437])|(~m[1372]&~m[1433]&m[1434]&~m[1436]&m[1437])|(m[1372]&m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1372]&m[1433]&m[1434]&m[1436]&m[1437]))&UnbiasedRNG[359])|((m[1372]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(~m[1372]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1372]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1372]&m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1372]&~m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1372]&~m[1433]&~m[1434]&m[1436]&m[1437])|(m[1372]&~m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1372]&m[1433]&~m[1434]&m[1436]&m[1437])|(m[1372]&m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1372]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1372]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1372]&m[1433]&m[1434]&m[1436]&m[1437]));
    m[1440] = (((m[1377]&~m[1438]&~m[1439]&~m[1441]&~m[1442])|(~m[1377]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1377]&m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1377]&~m[1438]&m[1439]&m[1441]&~m[1442])|(~m[1377]&m[1438]&~m[1439]&~m[1441]&m[1442])|(~m[1377]&~m[1438]&m[1439]&~m[1441]&m[1442])|(m[1377]&m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1377]&m[1438]&m[1439]&m[1441]&m[1442]))&UnbiasedRNG[360])|((m[1377]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(~m[1377]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1377]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1377]&m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1377]&~m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1377]&~m[1438]&~m[1439]&m[1441]&m[1442])|(m[1377]&~m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1377]&m[1438]&~m[1439]&m[1441]&m[1442])|(m[1377]&m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1377]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1377]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1377]&m[1438]&m[1439]&m[1441]&m[1442]));
    m[1445] = (((m[1382]&~m[1443]&~m[1444]&~m[1446]&~m[1447])|(~m[1382]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1382]&m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1382]&~m[1443]&m[1444]&m[1446]&~m[1447])|(~m[1382]&m[1443]&~m[1444]&~m[1446]&m[1447])|(~m[1382]&~m[1443]&m[1444]&~m[1446]&m[1447])|(m[1382]&m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1382]&m[1443]&m[1444]&m[1446]&m[1447]))&UnbiasedRNG[361])|((m[1382]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(~m[1382]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1382]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1382]&m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1382]&~m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1382]&~m[1443]&~m[1444]&m[1446]&m[1447])|(m[1382]&~m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1382]&m[1443]&~m[1444]&m[1446]&m[1447])|(m[1382]&m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1382]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1382]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1382]&m[1443]&m[1444]&m[1446]&m[1447]));
    m[1455] = (((m[1387]&~m[1453]&~m[1454]&~m[1456]&~m[1457])|(~m[1387]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1387]&m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1387]&~m[1453]&m[1454]&m[1456]&~m[1457])|(~m[1387]&m[1453]&~m[1454]&~m[1456]&m[1457])|(~m[1387]&~m[1453]&m[1454]&~m[1456]&m[1457])|(m[1387]&m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1387]&m[1453]&m[1454]&m[1456]&m[1457]))&UnbiasedRNG[362])|((m[1387]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(~m[1387]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1387]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1387]&m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1387]&~m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1387]&~m[1453]&~m[1454]&m[1456]&m[1457])|(m[1387]&~m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1387]&m[1453]&~m[1454]&m[1456]&m[1457])|(m[1387]&m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1387]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1387]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1387]&m[1453]&m[1454]&m[1456]&m[1457]));
    m[1460] = (((m[1392]&~m[1458]&~m[1459]&~m[1461]&~m[1462])|(~m[1392]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1392]&m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1392]&~m[1458]&m[1459]&m[1461]&~m[1462])|(~m[1392]&m[1458]&~m[1459]&~m[1461]&m[1462])|(~m[1392]&~m[1458]&m[1459]&~m[1461]&m[1462])|(m[1392]&m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1392]&m[1458]&m[1459]&m[1461]&m[1462]))&UnbiasedRNG[363])|((m[1392]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(~m[1392]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1392]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1392]&m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1392]&~m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1392]&~m[1458]&~m[1459]&m[1461]&m[1462])|(m[1392]&~m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1392]&m[1458]&~m[1459]&m[1461]&m[1462])|(m[1392]&m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1392]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1392]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1392]&m[1458]&m[1459]&m[1461]&m[1462]));
    m[1465] = (((m[1397]&~m[1463]&~m[1464]&~m[1466]&~m[1467])|(~m[1397]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1397]&m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1397]&~m[1463]&m[1464]&m[1466]&~m[1467])|(~m[1397]&m[1463]&~m[1464]&~m[1466]&m[1467])|(~m[1397]&~m[1463]&m[1464]&~m[1466]&m[1467])|(m[1397]&m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1397]&m[1463]&m[1464]&m[1466]&m[1467]))&UnbiasedRNG[364])|((m[1397]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(~m[1397]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1397]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1397]&m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1397]&~m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1397]&~m[1463]&~m[1464]&m[1466]&m[1467])|(m[1397]&~m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1397]&m[1463]&~m[1464]&m[1466]&m[1467])|(m[1397]&m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1397]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1397]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1397]&m[1463]&m[1464]&m[1466]&m[1467]));
    m[1470] = (((m[1402]&~m[1468]&~m[1469]&~m[1471]&~m[1472])|(~m[1402]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1402]&m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1402]&~m[1468]&m[1469]&m[1471]&~m[1472])|(~m[1402]&m[1468]&~m[1469]&~m[1471]&m[1472])|(~m[1402]&~m[1468]&m[1469]&~m[1471]&m[1472])|(m[1402]&m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1402]&m[1468]&m[1469]&m[1471]&m[1472]))&UnbiasedRNG[365])|((m[1402]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(~m[1402]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1402]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1402]&m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1402]&~m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1402]&~m[1468]&~m[1469]&m[1471]&m[1472])|(m[1402]&~m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1402]&m[1468]&~m[1469]&m[1471]&m[1472])|(m[1402]&m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1402]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1402]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1402]&m[1468]&m[1469]&m[1471]&m[1472]));
    m[1475] = (((m[1407]&~m[1473]&~m[1474]&~m[1476]&~m[1477])|(~m[1407]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1407]&m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1407]&~m[1473]&m[1474]&m[1476]&~m[1477])|(~m[1407]&m[1473]&~m[1474]&~m[1476]&m[1477])|(~m[1407]&~m[1473]&m[1474]&~m[1476]&m[1477])|(m[1407]&m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1407]&m[1473]&m[1474]&m[1476]&m[1477]))&UnbiasedRNG[366])|((m[1407]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(~m[1407]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1407]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1407]&m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1407]&~m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1407]&~m[1473]&~m[1474]&m[1476]&m[1477])|(m[1407]&~m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1407]&m[1473]&~m[1474]&m[1476]&m[1477])|(m[1407]&m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1407]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1407]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1407]&m[1473]&m[1474]&m[1476]&m[1477]));
    m[1480] = (((m[1412]&~m[1478]&~m[1479]&~m[1481]&~m[1482])|(~m[1412]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1412]&m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1412]&~m[1478]&m[1479]&m[1481]&~m[1482])|(~m[1412]&m[1478]&~m[1479]&~m[1481]&m[1482])|(~m[1412]&~m[1478]&m[1479]&~m[1481]&m[1482])|(m[1412]&m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1412]&m[1478]&m[1479]&m[1481]&m[1482]))&UnbiasedRNG[367])|((m[1412]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(~m[1412]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1412]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1412]&m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1412]&~m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1412]&~m[1478]&~m[1479]&m[1481]&m[1482])|(m[1412]&~m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1412]&m[1478]&~m[1479]&m[1481]&m[1482])|(m[1412]&m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1412]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1412]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1412]&m[1478]&m[1479]&m[1481]&m[1482]));
    m[1485] = (((m[1417]&~m[1483]&~m[1484]&~m[1486]&~m[1487])|(~m[1417]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1417]&m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1417]&~m[1483]&m[1484]&m[1486]&~m[1487])|(~m[1417]&m[1483]&~m[1484]&~m[1486]&m[1487])|(~m[1417]&~m[1483]&m[1484]&~m[1486]&m[1487])|(m[1417]&m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1417]&m[1483]&m[1484]&m[1486]&m[1487]))&UnbiasedRNG[368])|((m[1417]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(~m[1417]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1417]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1417]&m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1417]&~m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1417]&~m[1483]&~m[1484]&m[1486]&m[1487])|(m[1417]&~m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1417]&m[1483]&~m[1484]&m[1486]&m[1487])|(m[1417]&m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1417]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1417]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1417]&m[1483]&m[1484]&m[1486]&m[1487]));
    m[1490] = (((m[1422]&~m[1488]&~m[1489]&~m[1491]&~m[1492])|(~m[1422]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1422]&m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1422]&~m[1488]&m[1489]&m[1491]&~m[1492])|(~m[1422]&m[1488]&~m[1489]&~m[1491]&m[1492])|(~m[1422]&~m[1488]&m[1489]&~m[1491]&m[1492])|(m[1422]&m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1422]&m[1488]&m[1489]&m[1491]&m[1492]))&UnbiasedRNG[369])|((m[1422]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(~m[1422]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1422]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1422]&m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1422]&~m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1422]&~m[1488]&~m[1489]&m[1491]&m[1492])|(m[1422]&~m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1422]&m[1488]&~m[1489]&m[1491]&m[1492])|(m[1422]&m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1422]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1422]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1422]&m[1488]&m[1489]&m[1491]&m[1492]));
    m[1495] = (((m[1427]&~m[1493]&~m[1494]&~m[1496]&~m[1497])|(~m[1427]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1427]&m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1427]&~m[1493]&m[1494]&m[1496]&~m[1497])|(~m[1427]&m[1493]&~m[1494]&~m[1496]&m[1497])|(~m[1427]&~m[1493]&m[1494]&~m[1496]&m[1497])|(m[1427]&m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1427]&m[1493]&m[1494]&m[1496]&m[1497]))&UnbiasedRNG[370])|((m[1427]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(~m[1427]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1427]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1427]&m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1427]&~m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1427]&~m[1493]&~m[1494]&m[1496]&m[1497])|(m[1427]&~m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1427]&m[1493]&~m[1494]&m[1496]&m[1497])|(m[1427]&m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1427]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1427]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1427]&m[1493]&m[1494]&m[1496]&m[1497]));
    m[1500] = (((m[1432]&~m[1498]&~m[1499]&~m[1501]&~m[1502])|(~m[1432]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1432]&m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1432]&~m[1498]&m[1499]&m[1501]&~m[1502])|(~m[1432]&m[1498]&~m[1499]&~m[1501]&m[1502])|(~m[1432]&~m[1498]&m[1499]&~m[1501]&m[1502])|(m[1432]&m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1432]&m[1498]&m[1499]&m[1501]&m[1502]))&UnbiasedRNG[371])|((m[1432]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(~m[1432]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1432]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1432]&m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1432]&~m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1432]&~m[1498]&~m[1499]&m[1501]&m[1502])|(m[1432]&~m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1432]&m[1498]&~m[1499]&m[1501]&m[1502])|(m[1432]&m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1432]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1432]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1432]&m[1498]&m[1499]&m[1501]&m[1502]));
    m[1505] = (((m[1437]&~m[1503]&~m[1504]&~m[1506]&~m[1507])|(~m[1437]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1437]&m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1437]&~m[1503]&m[1504]&m[1506]&~m[1507])|(~m[1437]&m[1503]&~m[1504]&~m[1506]&m[1507])|(~m[1437]&~m[1503]&m[1504]&~m[1506]&m[1507])|(m[1437]&m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1437]&m[1503]&m[1504]&m[1506]&m[1507]))&UnbiasedRNG[372])|((m[1437]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(~m[1437]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1437]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1437]&m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1437]&~m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1437]&~m[1503]&~m[1504]&m[1506]&m[1507])|(m[1437]&~m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1437]&m[1503]&~m[1504]&m[1506]&m[1507])|(m[1437]&m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1437]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1437]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1437]&m[1503]&m[1504]&m[1506]&m[1507]));
    m[1510] = (((m[1442]&~m[1508]&~m[1509]&~m[1511]&~m[1512])|(~m[1442]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1442]&m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1442]&~m[1508]&m[1509]&m[1511]&~m[1512])|(~m[1442]&m[1508]&~m[1509]&~m[1511]&m[1512])|(~m[1442]&~m[1508]&m[1509]&~m[1511]&m[1512])|(m[1442]&m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1442]&m[1508]&m[1509]&m[1511]&m[1512]))&UnbiasedRNG[373])|((m[1442]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(~m[1442]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1442]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1442]&m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1442]&~m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1442]&~m[1508]&~m[1509]&m[1511]&m[1512])|(m[1442]&~m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1442]&m[1508]&~m[1509]&m[1511]&m[1512])|(m[1442]&m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1442]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1442]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1442]&m[1508]&m[1509]&m[1511]&m[1512]));
    m[1515] = (((m[1447]&~m[1513]&~m[1514]&~m[1516]&~m[1517])|(~m[1447]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1447]&m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1447]&~m[1513]&m[1514]&m[1516]&~m[1517])|(~m[1447]&m[1513]&~m[1514]&~m[1516]&m[1517])|(~m[1447]&~m[1513]&m[1514]&~m[1516]&m[1517])|(m[1447]&m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1447]&m[1513]&m[1514]&m[1516]&m[1517]))&UnbiasedRNG[374])|((m[1447]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(~m[1447]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1447]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1447]&m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1447]&~m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1447]&~m[1513]&~m[1514]&m[1516]&m[1517])|(m[1447]&~m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1447]&m[1513]&~m[1514]&m[1516]&m[1517])|(m[1447]&m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1447]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1447]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1447]&m[1513]&m[1514]&m[1516]&m[1517]));
    m[1520] = (((m[1452]&~m[1518]&~m[1519]&~m[1521]&~m[1522])|(~m[1452]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1452]&m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1452]&~m[1518]&m[1519]&m[1521]&~m[1522])|(~m[1452]&m[1518]&~m[1519]&~m[1521]&m[1522])|(~m[1452]&~m[1518]&m[1519]&~m[1521]&m[1522])|(m[1452]&m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1452]&m[1518]&m[1519]&m[1521]&m[1522]))&UnbiasedRNG[375])|((m[1452]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(~m[1452]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1452]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1452]&m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1452]&~m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1452]&~m[1518]&~m[1519]&m[1521]&m[1522])|(m[1452]&~m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1452]&m[1518]&~m[1519]&m[1521]&m[1522])|(m[1452]&m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1452]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1452]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1452]&m[1518]&m[1519]&m[1521]&m[1522]));
    m[1530] = (((m[1457]&~m[1528]&~m[1529]&~m[1531]&~m[1532])|(~m[1457]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1457]&m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1457]&~m[1528]&m[1529]&m[1531]&~m[1532])|(~m[1457]&m[1528]&~m[1529]&~m[1531]&m[1532])|(~m[1457]&~m[1528]&m[1529]&~m[1531]&m[1532])|(m[1457]&m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1457]&m[1528]&m[1529]&m[1531]&m[1532]))&UnbiasedRNG[376])|((m[1457]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(~m[1457]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1457]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1457]&m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1457]&~m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1457]&~m[1528]&~m[1529]&m[1531]&m[1532])|(m[1457]&~m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1457]&m[1528]&~m[1529]&m[1531]&m[1532])|(m[1457]&m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1457]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1457]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1457]&m[1528]&m[1529]&m[1531]&m[1532]));
    m[1535] = (((m[1462]&~m[1533]&~m[1534]&~m[1536]&~m[1537])|(~m[1462]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1462]&m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1462]&~m[1533]&m[1534]&m[1536]&~m[1537])|(~m[1462]&m[1533]&~m[1534]&~m[1536]&m[1537])|(~m[1462]&~m[1533]&m[1534]&~m[1536]&m[1537])|(m[1462]&m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1462]&m[1533]&m[1534]&m[1536]&m[1537]))&UnbiasedRNG[377])|((m[1462]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(~m[1462]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1462]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1462]&m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1462]&~m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1462]&~m[1533]&~m[1534]&m[1536]&m[1537])|(m[1462]&~m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1462]&m[1533]&~m[1534]&m[1536]&m[1537])|(m[1462]&m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1462]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1462]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1462]&m[1533]&m[1534]&m[1536]&m[1537]));
    m[1540] = (((m[1467]&~m[1538]&~m[1539]&~m[1541]&~m[1542])|(~m[1467]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1467]&m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1467]&~m[1538]&m[1539]&m[1541]&~m[1542])|(~m[1467]&m[1538]&~m[1539]&~m[1541]&m[1542])|(~m[1467]&~m[1538]&m[1539]&~m[1541]&m[1542])|(m[1467]&m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1467]&m[1538]&m[1539]&m[1541]&m[1542]))&UnbiasedRNG[378])|((m[1467]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(~m[1467]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1467]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1467]&m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1467]&~m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1467]&~m[1538]&~m[1539]&m[1541]&m[1542])|(m[1467]&~m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1467]&m[1538]&~m[1539]&m[1541]&m[1542])|(m[1467]&m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1467]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1467]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1467]&m[1538]&m[1539]&m[1541]&m[1542]));
    m[1545] = (((m[1472]&~m[1543]&~m[1544]&~m[1546]&~m[1547])|(~m[1472]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1472]&m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1472]&~m[1543]&m[1544]&m[1546]&~m[1547])|(~m[1472]&m[1543]&~m[1544]&~m[1546]&m[1547])|(~m[1472]&~m[1543]&m[1544]&~m[1546]&m[1547])|(m[1472]&m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1472]&m[1543]&m[1544]&m[1546]&m[1547]))&UnbiasedRNG[379])|((m[1472]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(~m[1472]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1472]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1472]&m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1472]&~m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1472]&~m[1543]&~m[1544]&m[1546]&m[1547])|(m[1472]&~m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1472]&m[1543]&~m[1544]&m[1546]&m[1547])|(m[1472]&m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1472]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1472]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1472]&m[1543]&m[1544]&m[1546]&m[1547]));
    m[1550] = (((m[1477]&~m[1548]&~m[1549]&~m[1551]&~m[1552])|(~m[1477]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1477]&m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1477]&~m[1548]&m[1549]&m[1551]&~m[1552])|(~m[1477]&m[1548]&~m[1549]&~m[1551]&m[1552])|(~m[1477]&~m[1548]&m[1549]&~m[1551]&m[1552])|(m[1477]&m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1477]&m[1548]&m[1549]&m[1551]&m[1552]))&UnbiasedRNG[380])|((m[1477]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(~m[1477]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1477]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1477]&m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1477]&~m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1477]&~m[1548]&~m[1549]&m[1551]&m[1552])|(m[1477]&~m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1477]&m[1548]&~m[1549]&m[1551]&m[1552])|(m[1477]&m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1477]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1477]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1477]&m[1548]&m[1549]&m[1551]&m[1552]));
    m[1555] = (((m[1482]&~m[1553]&~m[1554]&~m[1556]&~m[1557])|(~m[1482]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1482]&m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1482]&~m[1553]&m[1554]&m[1556]&~m[1557])|(~m[1482]&m[1553]&~m[1554]&~m[1556]&m[1557])|(~m[1482]&~m[1553]&m[1554]&~m[1556]&m[1557])|(m[1482]&m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1482]&m[1553]&m[1554]&m[1556]&m[1557]))&UnbiasedRNG[381])|((m[1482]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(~m[1482]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1482]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1482]&m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1482]&~m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1482]&~m[1553]&~m[1554]&m[1556]&m[1557])|(m[1482]&~m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1482]&m[1553]&~m[1554]&m[1556]&m[1557])|(m[1482]&m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1482]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1482]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1482]&m[1553]&m[1554]&m[1556]&m[1557]));
    m[1560] = (((m[1487]&~m[1558]&~m[1559]&~m[1561]&~m[1562])|(~m[1487]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1487]&m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1487]&~m[1558]&m[1559]&m[1561]&~m[1562])|(~m[1487]&m[1558]&~m[1559]&~m[1561]&m[1562])|(~m[1487]&~m[1558]&m[1559]&~m[1561]&m[1562])|(m[1487]&m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1487]&m[1558]&m[1559]&m[1561]&m[1562]))&UnbiasedRNG[382])|((m[1487]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(~m[1487]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1487]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1487]&m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1487]&~m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1487]&~m[1558]&~m[1559]&m[1561]&m[1562])|(m[1487]&~m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1487]&m[1558]&~m[1559]&m[1561]&m[1562])|(m[1487]&m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1487]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1487]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1487]&m[1558]&m[1559]&m[1561]&m[1562]));
    m[1565] = (((m[1492]&~m[1563]&~m[1564]&~m[1566]&~m[1567])|(~m[1492]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1492]&m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1492]&~m[1563]&m[1564]&m[1566]&~m[1567])|(~m[1492]&m[1563]&~m[1564]&~m[1566]&m[1567])|(~m[1492]&~m[1563]&m[1564]&~m[1566]&m[1567])|(m[1492]&m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1492]&m[1563]&m[1564]&m[1566]&m[1567]))&UnbiasedRNG[383])|((m[1492]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(~m[1492]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1492]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1492]&m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1492]&~m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1492]&~m[1563]&~m[1564]&m[1566]&m[1567])|(m[1492]&~m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1492]&m[1563]&~m[1564]&m[1566]&m[1567])|(m[1492]&m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1492]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1492]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1492]&m[1563]&m[1564]&m[1566]&m[1567]));
    m[1570] = (((m[1497]&~m[1568]&~m[1569]&~m[1571]&~m[1572])|(~m[1497]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1497]&m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1497]&~m[1568]&m[1569]&m[1571]&~m[1572])|(~m[1497]&m[1568]&~m[1569]&~m[1571]&m[1572])|(~m[1497]&~m[1568]&m[1569]&~m[1571]&m[1572])|(m[1497]&m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1497]&m[1568]&m[1569]&m[1571]&m[1572]))&UnbiasedRNG[384])|((m[1497]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(~m[1497]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1497]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1497]&m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1497]&~m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1497]&~m[1568]&~m[1569]&m[1571]&m[1572])|(m[1497]&~m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1497]&m[1568]&~m[1569]&m[1571]&m[1572])|(m[1497]&m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1497]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1497]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1497]&m[1568]&m[1569]&m[1571]&m[1572]));
    m[1575] = (((m[1502]&~m[1573]&~m[1574]&~m[1576]&~m[1577])|(~m[1502]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1502]&m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1502]&~m[1573]&m[1574]&m[1576]&~m[1577])|(~m[1502]&m[1573]&~m[1574]&~m[1576]&m[1577])|(~m[1502]&~m[1573]&m[1574]&~m[1576]&m[1577])|(m[1502]&m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1502]&m[1573]&m[1574]&m[1576]&m[1577]))&UnbiasedRNG[385])|((m[1502]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(~m[1502]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1502]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1502]&m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1502]&~m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1502]&~m[1573]&~m[1574]&m[1576]&m[1577])|(m[1502]&~m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1502]&m[1573]&~m[1574]&m[1576]&m[1577])|(m[1502]&m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1502]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1502]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1502]&m[1573]&m[1574]&m[1576]&m[1577]));
    m[1580] = (((m[1507]&~m[1578]&~m[1579]&~m[1581]&~m[1582])|(~m[1507]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1507]&m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1507]&~m[1578]&m[1579]&m[1581]&~m[1582])|(~m[1507]&m[1578]&~m[1579]&~m[1581]&m[1582])|(~m[1507]&~m[1578]&m[1579]&~m[1581]&m[1582])|(m[1507]&m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1507]&m[1578]&m[1579]&m[1581]&m[1582]))&UnbiasedRNG[386])|((m[1507]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(~m[1507]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1507]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1507]&m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1507]&~m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1507]&~m[1578]&~m[1579]&m[1581]&m[1582])|(m[1507]&~m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1507]&m[1578]&~m[1579]&m[1581]&m[1582])|(m[1507]&m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1507]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1507]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1507]&m[1578]&m[1579]&m[1581]&m[1582]));
    m[1585] = (((m[1512]&~m[1583]&~m[1584]&~m[1586]&~m[1587])|(~m[1512]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1512]&m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1512]&~m[1583]&m[1584]&m[1586]&~m[1587])|(~m[1512]&m[1583]&~m[1584]&~m[1586]&m[1587])|(~m[1512]&~m[1583]&m[1584]&~m[1586]&m[1587])|(m[1512]&m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1512]&m[1583]&m[1584]&m[1586]&m[1587]))&UnbiasedRNG[387])|((m[1512]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(~m[1512]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1512]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1512]&m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1512]&~m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1512]&~m[1583]&~m[1584]&m[1586]&m[1587])|(m[1512]&~m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1512]&m[1583]&~m[1584]&m[1586]&m[1587])|(m[1512]&m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1512]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1512]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1512]&m[1583]&m[1584]&m[1586]&m[1587]));
    m[1590] = (((m[1517]&~m[1588]&~m[1589]&~m[1591]&~m[1592])|(~m[1517]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1517]&m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1517]&~m[1588]&m[1589]&m[1591]&~m[1592])|(~m[1517]&m[1588]&~m[1589]&~m[1591]&m[1592])|(~m[1517]&~m[1588]&m[1589]&~m[1591]&m[1592])|(m[1517]&m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1517]&m[1588]&m[1589]&m[1591]&m[1592]))&UnbiasedRNG[388])|((m[1517]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(~m[1517]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1517]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1517]&m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1517]&~m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1517]&~m[1588]&~m[1589]&m[1591]&m[1592])|(m[1517]&~m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1517]&m[1588]&~m[1589]&m[1591]&m[1592])|(m[1517]&m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1517]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1517]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1517]&m[1588]&m[1589]&m[1591]&m[1592]));
    m[1595] = (((m[1522]&~m[1593]&~m[1594]&~m[1596]&~m[1597])|(~m[1522]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1522]&m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1522]&~m[1593]&m[1594]&m[1596]&~m[1597])|(~m[1522]&m[1593]&~m[1594]&~m[1596]&m[1597])|(~m[1522]&~m[1593]&m[1594]&~m[1596]&m[1597])|(m[1522]&m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1522]&m[1593]&m[1594]&m[1596]&m[1597]))&UnbiasedRNG[389])|((m[1522]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(~m[1522]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1522]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1522]&m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1522]&~m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1522]&~m[1593]&~m[1594]&m[1596]&m[1597])|(m[1522]&~m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1522]&m[1593]&~m[1594]&m[1596]&m[1597])|(m[1522]&m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1522]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1522]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1522]&m[1593]&m[1594]&m[1596]&m[1597]));
    m[1600] = (((m[1527]&~m[1598]&~m[1599]&~m[1601]&~m[1602])|(~m[1527]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1527]&m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1527]&~m[1598]&m[1599]&m[1601]&~m[1602])|(~m[1527]&m[1598]&~m[1599]&~m[1601]&m[1602])|(~m[1527]&~m[1598]&m[1599]&~m[1601]&m[1602])|(m[1527]&m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1527]&m[1598]&m[1599]&m[1601]&m[1602]))&UnbiasedRNG[390])|((m[1527]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(~m[1527]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1527]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1527]&m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1527]&~m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1527]&~m[1598]&~m[1599]&m[1601]&m[1602])|(m[1527]&~m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1527]&m[1598]&~m[1599]&m[1601]&m[1602])|(m[1527]&m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1527]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1527]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1527]&m[1598]&m[1599]&m[1601]&m[1602]));
    m[1605] = (((m[1537]&~m[1603]&~m[1604]&~m[1606]&~m[1607])|(~m[1537]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1537]&m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1537]&~m[1603]&m[1604]&m[1606]&~m[1607])|(~m[1537]&m[1603]&~m[1604]&~m[1606]&m[1607])|(~m[1537]&~m[1603]&m[1604]&~m[1606]&m[1607])|(m[1537]&m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1537]&m[1603]&m[1604]&m[1606]&m[1607]))&UnbiasedRNG[391])|((m[1537]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(~m[1537]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1537]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1537]&m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1537]&~m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1537]&~m[1603]&~m[1604]&m[1606]&m[1607])|(m[1537]&~m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1537]&m[1603]&~m[1604]&m[1606]&m[1607])|(m[1537]&m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1537]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1537]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1537]&m[1603]&m[1604]&m[1606]&m[1607]));
    m[1610] = (((m[1542]&~m[1608]&~m[1609]&~m[1611]&~m[1612])|(~m[1542]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1542]&m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1542]&~m[1608]&m[1609]&m[1611]&~m[1612])|(~m[1542]&m[1608]&~m[1609]&~m[1611]&m[1612])|(~m[1542]&~m[1608]&m[1609]&~m[1611]&m[1612])|(m[1542]&m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1542]&m[1608]&m[1609]&m[1611]&m[1612]))&UnbiasedRNG[392])|((m[1542]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(~m[1542]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1542]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1542]&m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1542]&~m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1542]&~m[1608]&~m[1609]&m[1611]&m[1612])|(m[1542]&~m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1542]&m[1608]&~m[1609]&m[1611]&m[1612])|(m[1542]&m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1542]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1542]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1542]&m[1608]&m[1609]&m[1611]&m[1612]));
    m[1615] = (((m[1547]&~m[1613]&~m[1614]&~m[1616]&~m[1617])|(~m[1547]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1547]&m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1547]&~m[1613]&m[1614]&m[1616]&~m[1617])|(~m[1547]&m[1613]&~m[1614]&~m[1616]&m[1617])|(~m[1547]&~m[1613]&m[1614]&~m[1616]&m[1617])|(m[1547]&m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1547]&m[1613]&m[1614]&m[1616]&m[1617]))&UnbiasedRNG[393])|((m[1547]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(~m[1547]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1547]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1547]&m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1547]&~m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1547]&~m[1613]&~m[1614]&m[1616]&m[1617])|(m[1547]&~m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1547]&m[1613]&~m[1614]&m[1616]&m[1617])|(m[1547]&m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1547]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1547]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1547]&m[1613]&m[1614]&m[1616]&m[1617]));
    m[1620] = (((m[1552]&~m[1618]&~m[1619]&~m[1621]&~m[1622])|(~m[1552]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1552]&m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1552]&~m[1618]&m[1619]&m[1621]&~m[1622])|(~m[1552]&m[1618]&~m[1619]&~m[1621]&m[1622])|(~m[1552]&~m[1618]&m[1619]&~m[1621]&m[1622])|(m[1552]&m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1552]&m[1618]&m[1619]&m[1621]&m[1622]))&UnbiasedRNG[394])|((m[1552]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(~m[1552]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1552]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1552]&m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1552]&~m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1552]&~m[1618]&~m[1619]&m[1621]&m[1622])|(m[1552]&~m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1552]&m[1618]&~m[1619]&m[1621]&m[1622])|(m[1552]&m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1552]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1552]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1552]&m[1618]&m[1619]&m[1621]&m[1622]));
    m[1625] = (((m[1557]&~m[1623]&~m[1624]&~m[1626]&~m[1627])|(~m[1557]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1557]&m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1557]&~m[1623]&m[1624]&m[1626]&~m[1627])|(~m[1557]&m[1623]&~m[1624]&~m[1626]&m[1627])|(~m[1557]&~m[1623]&m[1624]&~m[1626]&m[1627])|(m[1557]&m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1557]&m[1623]&m[1624]&m[1626]&m[1627]))&UnbiasedRNG[395])|((m[1557]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(~m[1557]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1557]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1557]&m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1557]&~m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1557]&~m[1623]&~m[1624]&m[1626]&m[1627])|(m[1557]&~m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1557]&m[1623]&~m[1624]&m[1626]&m[1627])|(m[1557]&m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1557]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1557]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1557]&m[1623]&m[1624]&m[1626]&m[1627]));
    m[1630] = (((m[1562]&~m[1628]&~m[1629]&~m[1631]&~m[1632])|(~m[1562]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1562]&m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1562]&~m[1628]&m[1629]&m[1631]&~m[1632])|(~m[1562]&m[1628]&~m[1629]&~m[1631]&m[1632])|(~m[1562]&~m[1628]&m[1629]&~m[1631]&m[1632])|(m[1562]&m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1562]&m[1628]&m[1629]&m[1631]&m[1632]))&UnbiasedRNG[396])|((m[1562]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(~m[1562]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1562]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1562]&m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1562]&~m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1562]&~m[1628]&~m[1629]&m[1631]&m[1632])|(m[1562]&~m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1562]&m[1628]&~m[1629]&m[1631]&m[1632])|(m[1562]&m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1562]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1562]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1562]&m[1628]&m[1629]&m[1631]&m[1632]));
    m[1635] = (((m[1567]&~m[1633]&~m[1634]&~m[1636]&~m[1637])|(~m[1567]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1567]&m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1567]&~m[1633]&m[1634]&m[1636]&~m[1637])|(~m[1567]&m[1633]&~m[1634]&~m[1636]&m[1637])|(~m[1567]&~m[1633]&m[1634]&~m[1636]&m[1637])|(m[1567]&m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1567]&m[1633]&m[1634]&m[1636]&m[1637]))&UnbiasedRNG[397])|((m[1567]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(~m[1567]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1567]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1567]&m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1567]&~m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1567]&~m[1633]&~m[1634]&m[1636]&m[1637])|(m[1567]&~m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1567]&m[1633]&~m[1634]&m[1636]&m[1637])|(m[1567]&m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1567]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1567]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1567]&m[1633]&m[1634]&m[1636]&m[1637]));
    m[1640] = (((m[1572]&~m[1638]&~m[1639]&~m[1641]&~m[1642])|(~m[1572]&~m[1638]&~m[1639]&m[1641]&~m[1642])|(m[1572]&m[1638]&~m[1639]&m[1641]&~m[1642])|(m[1572]&~m[1638]&m[1639]&m[1641]&~m[1642])|(~m[1572]&m[1638]&~m[1639]&~m[1641]&m[1642])|(~m[1572]&~m[1638]&m[1639]&~m[1641]&m[1642])|(m[1572]&m[1638]&m[1639]&~m[1641]&m[1642])|(~m[1572]&m[1638]&m[1639]&m[1641]&m[1642]))&UnbiasedRNG[398])|((m[1572]&~m[1638]&~m[1639]&m[1641]&~m[1642])|(~m[1572]&~m[1638]&~m[1639]&~m[1641]&m[1642])|(m[1572]&~m[1638]&~m[1639]&~m[1641]&m[1642])|(m[1572]&m[1638]&~m[1639]&~m[1641]&m[1642])|(m[1572]&~m[1638]&m[1639]&~m[1641]&m[1642])|(~m[1572]&~m[1638]&~m[1639]&m[1641]&m[1642])|(m[1572]&~m[1638]&~m[1639]&m[1641]&m[1642])|(~m[1572]&m[1638]&~m[1639]&m[1641]&m[1642])|(m[1572]&m[1638]&~m[1639]&m[1641]&m[1642])|(~m[1572]&~m[1638]&m[1639]&m[1641]&m[1642])|(m[1572]&~m[1638]&m[1639]&m[1641]&m[1642])|(m[1572]&m[1638]&m[1639]&m[1641]&m[1642]));
    m[1645] = (((m[1577]&~m[1643]&~m[1644]&~m[1646]&~m[1647])|(~m[1577]&~m[1643]&~m[1644]&m[1646]&~m[1647])|(m[1577]&m[1643]&~m[1644]&m[1646]&~m[1647])|(m[1577]&~m[1643]&m[1644]&m[1646]&~m[1647])|(~m[1577]&m[1643]&~m[1644]&~m[1646]&m[1647])|(~m[1577]&~m[1643]&m[1644]&~m[1646]&m[1647])|(m[1577]&m[1643]&m[1644]&~m[1646]&m[1647])|(~m[1577]&m[1643]&m[1644]&m[1646]&m[1647]))&UnbiasedRNG[399])|((m[1577]&~m[1643]&~m[1644]&m[1646]&~m[1647])|(~m[1577]&~m[1643]&~m[1644]&~m[1646]&m[1647])|(m[1577]&~m[1643]&~m[1644]&~m[1646]&m[1647])|(m[1577]&m[1643]&~m[1644]&~m[1646]&m[1647])|(m[1577]&~m[1643]&m[1644]&~m[1646]&m[1647])|(~m[1577]&~m[1643]&~m[1644]&m[1646]&m[1647])|(m[1577]&~m[1643]&~m[1644]&m[1646]&m[1647])|(~m[1577]&m[1643]&~m[1644]&m[1646]&m[1647])|(m[1577]&m[1643]&~m[1644]&m[1646]&m[1647])|(~m[1577]&~m[1643]&m[1644]&m[1646]&m[1647])|(m[1577]&~m[1643]&m[1644]&m[1646]&m[1647])|(m[1577]&m[1643]&m[1644]&m[1646]&m[1647]));
    m[1650] = (((m[1582]&~m[1648]&~m[1649]&~m[1651]&~m[1652])|(~m[1582]&~m[1648]&~m[1649]&m[1651]&~m[1652])|(m[1582]&m[1648]&~m[1649]&m[1651]&~m[1652])|(m[1582]&~m[1648]&m[1649]&m[1651]&~m[1652])|(~m[1582]&m[1648]&~m[1649]&~m[1651]&m[1652])|(~m[1582]&~m[1648]&m[1649]&~m[1651]&m[1652])|(m[1582]&m[1648]&m[1649]&~m[1651]&m[1652])|(~m[1582]&m[1648]&m[1649]&m[1651]&m[1652]))&UnbiasedRNG[400])|((m[1582]&~m[1648]&~m[1649]&m[1651]&~m[1652])|(~m[1582]&~m[1648]&~m[1649]&~m[1651]&m[1652])|(m[1582]&~m[1648]&~m[1649]&~m[1651]&m[1652])|(m[1582]&m[1648]&~m[1649]&~m[1651]&m[1652])|(m[1582]&~m[1648]&m[1649]&~m[1651]&m[1652])|(~m[1582]&~m[1648]&~m[1649]&m[1651]&m[1652])|(m[1582]&~m[1648]&~m[1649]&m[1651]&m[1652])|(~m[1582]&m[1648]&~m[1649]&m[1651]&m[1652])|(m[1582]&m[1648]&~m[1649]&m[1651]&m[1652])|(~m[1582]&~m[1648]&m[1649]&m[1651]&m[1652])|(m[1582]&~m[1648]&m[1649]&m[1651]&m[1652])|(m[1582]&m[1648]&m[1649]&m[1651]&m[1652]));
    m[1655] = (((m[1587]&~m[1653]&~m[1654]&~m[1656]&~m[1657])|(~m[1587]&~m[1653]&~m[1654]&m[1656]&~m[1657])|(m[1587]&m[1653]&~m[1654]&m[1656]&~m[1657])|(m[1587]&~m[1653]&m[1654]&m[1656]&~m[1657])|(~m[1587]&m[1653]&~m[1654]&~m[1656]&m[1657])|(~m[1587]&~m[1653]&m[1654]&~m[1656]&m[1657])|(m[1587]&m[1653]&m[1654]&~m[1656]&m[1657])|(~m[1587]&m[1653]&m[1654]&m[1656]&m[1657]))&UnbiasedRNG[401])|((m[1587]&~m[1653]&~m[1654]&m[1656]&~m[1657])|(~m[1587]&~m[1653]&~m[1654]&~m[1656]&m[1657])|(m[1587]&~m[1653]&~m[1654]&~m[1656]&m[1657])|(m[1587]&m[1653]&~m[1654]&~m[1656]&m[1657])|(m[1587]&~m[1653]&m[1654]&~m[1656]&m[1657])|(~m[1587]&~m[1653]&~m[1654]&m[1656]&m[1657])|(m[1587]&~m[1653]&~m[1654]&m[1656]&m[1657])|(~m[1587]&m[1653]&~m[1654]&m[1656]&m[1657])|(m[1587]&m[1653]&~m[1654]&m[1656]&m[1657])|(~m[1587]&~m[1653]&m[1654]&m[1656]&m[1657])|(m[1587]&~m[1653]&m[1654]&m[1656]&m[1657])|(m[1587]&m[1653]&m[1654]&m[1656]&m[1657]));
    m[1660] = (((m[1592]&~m[1658]&~m[1659]&~m[1661]&~m[1662])|(~m[1592]&~m[1658]&~m[1659]&m[1661]&~m[1662])|(m[1592]&m[1658]&~m[1659]&m[1661]&~m[1662])|(m[1592]&~m[1658]&m[1659]&m[1661]&~m[1662])|(~m[1592]&m[1658]&~m[1659]&~m[1661]&m[1662])|(~m[1592]&~m[1658]&m[1659]&~m[1661]&m[1662])|(m[1592]&m[1658]&m[1659]&~m[1661]&m[1662])|(~m[1592]&m[1658]&m[1659]&m[1661]&m[1662]))&UnbiasedRNG[402])|((m[1592]&~m[1658]&~m[1659]&m[1661]&~m[1662])|(~m[1592]&~m[1658]&~m[1659]&~m[1661]&m[1662])|(m[1592]&~m[1658]&~m[1659]&~m[1661]&m[1662])|(m[1592]&m[1658]&~m[1659]&~m[1661]&m[1662])|(m[1592]&~m[1658]&m[1659]&~m[1661]&m[1662])|(~m[1592]&~m[1658]&~m[1659]&m[1661]&m[1662])|(m[1592]&~m[1658]&~m[1659]&m[1661]&m[1662])|(~m[1592]&m[1658]&~m[1659]&m[1661]&m[1662])|(m[1592]&m[1658]&~m[1659]&m[1661]&m[1662])|(~m[1592]&~m[1658]&m[1659]&m[1661]&m[1662])|(m[1592]&~m[1658]&m[1659]&m[1661]&m[1662])|(m[1592]&m[1658]&m[1659]&m[1661]&m[1662]));
    m[1665] = (((m[1597]&~m[1663]&~m[1664]&~m[1666]&~m[1667])|(~m[1597]&~m[1663]&~m[1664]&m[1666]&~m[1667])|(m[1597]&m[1663]&~m[1664]&m[1666]&~m[1667])|(m[1597]&~m[1663]&m[1664]&m[1666]&~m[1667])|(~m[1597]&m[1663]&~m[1664]&~m[1666]&m[1667])|(~m[1597]&~m[1663]&m[1664]&~m[1666]&m[1667])|(m[1597]&m[1663]&m[1664]&~m[1666]&m[1667])|(~m[1597]&m[1663]&m[1664]&m[1666]&m[1667]))&UnbiasedRNG[403])|((m[1597]&~m[1663]&~m[1664]&m[1666]&~m[1667])|(~m[1597]&~m[1663]&~m[1664]&~m[1666]&m[1667])|(m[1597]&~m[1663]&~m[1664]&~m[1666]&m[1667])|(m[1597]&m[1663]&~m[1664]&~m[1666]&m[1667])|(m[1597]&~m[1663]&m[1664]&~m[1666]&m[1667])|(~m[1597]&~m[1663]&~m[1664]&m[1666]&m[1667])|(m[1597]&~m[1663]&~m[1664]&m[1666]&m[1667])|(~m[1597]&m[1663]&~m[1664]&m[1666]&m[1667])|(m[1597]&m[1663]&~m[1664]&m[1666]&m[1667])|(~m[1597]&~m[1663]&m[1664]&m[1666]&m[1667])|(m[1597]&~m[1663]&m[1664]&m[1666]&m[1667])|(m[1597]&m[1663]&m[1664]&m[1666]&m[1667]));
    m[1670] = (((m[1602]&~m[1668]&~m[1669]&~m[1671]&~m[1672])|(~m[1602]&~m[1668]&~m[1669]&m[1671]&~m[1672])|(m[1602]&m[1668]&~m[1669]&m[1671]&~m[1672])|(m[1602]&~m[1668]&m[1669]&m[1671]&~m[1672])|(~m[1602]&m[1668]&~m[1669]&~m[1671]&m[1672])|(~m[1602]&~m[1668]&m[1669]&~m[1671]&m[1672])|(m[1602]&m[1668]&m[1669]&~m[1671]&m[1672])|(~m[1602]&m[1668]&m[1669]&m[1671]&m[1672]))&UnbiasedRNG[404])|((m[1602]&~m[1668]&~m[1669]&m[1671]&~m[1672])|(~m[1602]&~m[1668]&~m[1669]&~m[1671]&m[1672])|(m[1602]&~m[1668]&~m[1669]&~m[1671]&m[1672])|(m[1602]&m[1668]&~m[1669]&~m[1671]&m[1672])|(m[1602]&~m[1668]&m[1669]&~m[1671]&m[1672])|(~m[1602]&~m[1668]&~m[1669]&m[1671]&m[1672])|(m[1602]&~m[1668]&~m[1669]&m[1671]&m[1672])|(~m[1602]&m[1668]&~m[1669]&m[1671]&m[1672])|(m[1602]&m[1668]&~m[1669]&m[1671]&m[1672])|(~m[1602]&~m[1668]&m[1669]&m[1671]&m[1672])|(m[1602]&~m[1668]&m[1669]&m[1671]&m[1672])|(m[1602]&m[1668]&m[1669]&m[1671]&m[1672]));
    m[1675] = (((m[1612]&~m[1673]&~m[1674]&~m[1676]&~m[1677])|(~m[1612]&~m[1673]&~m[1674]&m[1676]&~m[1677])|(m[1612]&m[1673]&~m[1674]&m[1676]&~m[1677])|(m[1612]&~m[1673]&m[1674]&m[1676]&~m[1677])|(~m[1612]&m[1673]&~m[1674]&~m[1676]&m[1677])|(~m[1612]&~m[1673]&m[1674]&~m[1676]&m[1677])|(m[1612]&m[1673]&m[1674]&~m[1676]&m[1677])|(~m[1612]&m[1673]&m[1674]&m[1676]&m[1677]))&UnbiasedRNG[405])|((m[1612]&~m[1673]&~m[1674]&m[1676]&~m[1677])|(~m[1612]&~m[1673]&~m[1674]&~m[1676]&m[1677])|(m[1612]&~m[1673]&~m[1674]&~m[1676]&m[1677])|(m[1612]&m[1673]&~m[1674]&~m[1676]&m[1677])|(m[1612]&~m[1673]&m[1674]&~m[1676]&m[1677])|(~m[1612]&~m[1673]&~m[1674]&m[1676]&m[1677])|(m[1612]&~m[1673]&~m[1674]&m[1676]&m[1677])|(~m[1612]&m[1673]&~m[1674]&m[1676]&m[1677])|(m[1612]&m[1673]&~m[1674]&m[1676]&m[1677])|(~m[1612]&~m[1673]&m[1674]&m[1676]&m[1677])|(m[1612]&~m[1673]&m[1674]&m[1676]&m[1677])|(m[1612]&m[1673]&m[1674]&m[1676]&m[1677]));
    m[1680] = (((m[1617]&~m[1678]&~m[1679]&~m[1681]&~m[1682])|(~m[1617]&~m[1678]&~m[1679]&m[1681]&~m[1682])|(m[1617]&m[1678]&~m[1679]&m[1681]&~m[1682])|(m[1617]&~m[1678]&m[1679]&m[1681]&~m[1682])|(~m[1617]&m[1678]&~m[1679]&~m[1681]&m[1682])|(~m[1617]&~m[1678]&m[1679]&~m[1681]&m[1682])|(m[1617]&m[1678]&m[1679]&~m[1681]&m[1682])|(~m[1617]&m[1678]&m[1679]&m[1681]&m[1682]))&UnbiasedRNG[406])|((m[1617]&~m[1678]&~m[1679]&m[1681]&~m[1682])|(~m[1617]&~m[1678]&~m[1679]&~m[1681]&m[1682])|(m[1617]&~m[1678]&~m[1679]&~m[1681]&m[1682])|(m[1617]&m[1678]&~m[1679]&~m[1681]&m[1682])|(m[1617]&~m[1678]&m[1679]&~m[1681]&m[1682])|(~m[1617]&~m[1678]&~m[1679]&m[1681]&m[1682])|(m[1617]&~m[1678]&~m[1679]&m[1681]&m[1682])|(~m[1617]&m[1678]&~m[1679]&m[1681]&m[1682])|(m[1617]&m[1678]&~m[1679]&m[1681]&m[1682])|(~m[1617]&~m[1678]&m[1679]&m[1681]&m[1682])|(m[1617]&~m[1678]&m[1679]&m[1681]&m[1682])|(m[1617]&m[1678]&m[1679]&m[1681]&m[1682]));
    m[1685] = (((m[1622]&~m[1683]&~m[1684]&~m[1686]&~m[1687])|(~m[1622]&~m[1683]&~m[1684]&m[1686]&~m[1687])|(m[1622]&m[1683]&~m[1684]&m[1686]&~m[1687])|(m[1622]&~m[1683]&m[1684]&m[1686]&~m[1687])|(~m[1622]&m[1683]&~m[1684]&~m[1686]&m[1687])|(~m[1622]&~m[1683]&m[1684]&~m[1686]&m[1687])|(m[1622]&m[1683]&m[1684]&~m[1686]&m[1687])|(~m[1622]&m[1683]&m[1684]&m[1686]&m[1687]))&UnbiasedRNG[407])|((m[1622]&~m[1683]&~m[1684]&m[1686]&~m[1687])|(~m[1622]&~m[1683]&~m[1684]&~m[1686]&m[1687])|(m[1622]&~m[1683]&~m[1684]&~m[1686]&m[1687])|(m[1622]&m[1683]&~m[1684]&~m[1686]&m[1687])|(m[1622]&~m[1683]&m[1684]&~m[1686]&m[1687])|(~m[1622]&~m[1683]&~m[1684]&m[1686]&m[1687])|(m[1622]&~m[1683]&~m[1684]&m[1686]&m[1687])|(~m[1622]&m[1683]&~m[1684]&m[1686]&m[1687])|(m[1622]&m[1683]&~m[1684]&m[1686]&m[1687])|(~m[1622]&~m[1683]&m[1684]&m[1686]&m[1687])|(m[1622]&~m[1683]&m[1684]&m[1686]&m[1687])|(m[1622]&m[1683]&m[1684]&m[1686]&m[1687]));
    m[1690] = (((m[1627]&~m[1688]&~m[1689]&~m[1691]&~m[1692])|(~m[1627]&~m[1688]&~m[1689]&m[1691]&~m[1692])|(m[1627]&m[1688]&~m[1689]&m[1691]&~m[1692])|(m[1627]&~m[1688]&m[1689]&m[1691]&~m[1692])|(~m[1627]&m[1688]&~m[1689]&~m[1691]&m[1692])|(~m[1627]&~m[1688]&m[1689]&~m[1691]&m[1692])|(m[1627]&m[1688]&m[1689]&~m[1691]&m[1692])|(~m[1627]&m[1688]&m[1689]&m[1691]&m[1692]))&UnbiasedRNG[408])|((m[1627]&~m[1688]&~m[1689]&m[1691]&~m[1692])|(~m[1627]&~m[1688]&~m[1689]&~m[1691]&m[1692])|(m[1627]&~m[1688]&~m[1689]&~m[1691]&m[1692])|(m[1627]&m[1688]&~m[1689]&~m[1691]&m[1692])|(m[1627]&~m[1688]&m[1689]&~m[1691]&m[1692])|(~m[1627]&~m[1688]&~m[1689]&m[1691]&m[1692])|(m[1627]&~m[1688]&~m[1689]&m[1691]&m[1692])|(~m[1627]&m[1688]&~m[1689]&m[1691]&m[1692])|(m[1627]&m[1688]&~m[1689]&m[1691]&m[1692])|(~m[1627]&~m[1688]&m[1689]&m[1691]&m[1692])|(m[1627]&~m[1688]&m[1689]&m[1691]&m[1692])|(m[1627]&m[1688]&m[1689]&m[1691]&m[1692]));
    m[1695] = (((m[1632]&~m[1693]&~m[1694]&~m[1696]&~m[1697])|(~m[1632]&~m[1693]&~m[1694]&m[1696]&~m[1697])|(m[1632]&m[1693]&~m[1694]&m[1696]&~m[1697])|(m[1632]&~m[1693]&m[1694]&m[1696]&~m[1697])|(~m[1632]&m[1693]&~m[1694]&~m[1696]&m[1697])|(~m[1632]&~m[1693]&m[1694]&~m[1696]&m[1697])|(m[1632]&m[1693]&m[1694]&~m[1696]&m[1697])|(~m[1632]&m[1693]&m[1694]&m[1696]&m[1697]))&UnbiasedRNG[409])|((m[1632]&~m[1693]&~m[1694]&m[1696]&~m[1697])|(~m[1632]&~m[1693]&~m[1694]&~m[1696]&m[1697])|(m[1632]&~m[1693]&~m[1694]&~m[1696]&m[1697])|(m[1632]&m[1693]&~m[1694]&~m[1696]&m[1697])|(m[1632]&~m[1693]&m[1694]&~m[1696]&m[1697])|(~m[1632]&~m[1693]&~m[1694]&m[1696]&m[1697])|(m[1632]&~m[1693]&~m[1694]&m[1696]&m[1697])|(~m[1632]&m[1693]&~m[1694]&m[1696]&m[1697])|(m[1632]&m[1693]&~m[1694]&m[1696]&m[1697])|(~m[1632]&~m[1693]&m[1694]&m[1696]&m[1697])|(m[1632]&~m[1693]&m[1694]&m[1696]&m[1697])|(m[1632]&m[1693]&m[1694]&m[1696]&m[1697]));
    m[1700] = (((m[1637]&~m[1698]&~m[1699]&~m[1701]&~m[1702])|(~m[1637]&~m[1698]&~m[1699]&m[1701]&~m[1702])|(m[1637]&m[1698]&~m[1699]&m[1701]&~m[1702])|(m[1637]&~m[1698]&m[1699]&m[1701]&~m[1702])|(~m[1637]&m[1698]&~m[1699]&~m[1701]&m[1702])|(~m[1637]&~m[1698]&m[1699]&~m[1701]&m[1702])|(m[1637]&m[1698]&m[1699]&~m[1701]&m[1702])|(~m[1637]&m[1698]&m[1699]&m[1701]&m[1702]))&UnbiasedRNG[410])|((m[1637]&~m[1698]&~m[1699]&m[1701]&~m[1702])|(~m[1637]&~m[1698]&~m[1699]&~m[1701]&m[1702])|(m[1637]&~m[1698]&~m[1699]&~m[1701]&m[1702])|(m[1637]&m[1698]&~m[1699]&~m[1701]&m[1702])|(m[1637]&~m[1698]&m[1699]&~m[1701]&m[1702])|(~m[1637]&~m[1698]&~m[1699]&m[1701]&m[1702])|(m[1637]&~m[1698]&~m[1699]&m[1701]&m[1702])|(~m[1637]&m[1698]&~m[1699]&m[1701]&m[1702])|(m[1637]&m[1698]&~m[1699]&m[1701]&m[1702])|(~m[1637]&~m[1698]&m[1699]&m[1701]&m[1702])|(m[1637]&~m[1698]&m[1699]&m[1701]&m[1702])|(m[1637]&m[1698]&m[1699]&m[1701]&m[1702]));
    m[1705] = (((m[1642]&~m[1703]&~m[1704]&~m[1706]&~m[1707])|(~m[1642]&~m[1703]&~m[1704]&m[1706]&~m[1707])|(m[1642]&m[1703]&~m[1704]&m[1706]&~m[1707])|(m[1642]&~m[1703]&m[1704]&m[1706]&~m[1707])|(~m[1642]&m[1703]&~m[1704]&~m[1706]&m[1707])|(~m[1642]&~m[1703]&m[1704]&~m[1706]&m[1707])|(m[1642]&m[1703]&m[1704]&~m[1706]&m[1707])|(~m[1642]&m[1703]&m[1704]&m[1706]&m[1707]))&UnbiasedRNG[411])|((m[1642]&~m[1703]&~m[1704]&m[1706]&~m[1707])|(~m[1642]&~m[1703]&~m[1704]&~m[1706]&m[1707])|(m[1642]&~m[1703]&~m[1704]&~m[1706]&m[1707])|(m[1642]&m[1703]&~m[1704]&~m[1706]&m[1707])|(m[1642]&~m[1703]&m[1704]&~m[1706]&m[1707])|(~m[1642]&~m[1703]&~m[1704]&m[1706]&m[1707])|(m[1642]&~m[1703]&~m[1704]&m[1706]&m[1707])|(~m[1642]&m[1703]&~m[1704]&m[1706]&m[1707])|(m[1642]&m[1703]&~m[1704]&m[1706]&m[1707])|(~m[1642]&~m[1703]&m[1704]&m[1706]&m[1707])|(m[1642]&~m[1703]&m[1704]&m[1706]&m[1707])|(m[1642]&m[1703]&m[1704]&m[1706]&m[1707]));
    m[1710] = (((m[1647]&~m[1708]&~m[1709]&~m[1711]&~m[1712])|(~m[1647]&~m[1708]&~m[1709]&m[1711]&~m[1712])|(m[1647]&m[1708]&~m[1709]&m[1711]&~m[1712])|(m[1647]&~m[1708]&m[1709]&m[1711]&~m[1712])|(~m[1647]&m[1708]&~m[1709]&~m[1711]&m[1712])|(~m[1647]&~m[1708]&m[1709]&~m[1711]&m[1712])|(m[1647]&m[1708]&m[1709]&~m[1711]&m[1712])|(~m[1647]&m[1708]&m[1709]&m[1711]&m[1712]))&UnbiasedRNG[412])|((m[1647]&~m[1708]&~m[1709]&m[1711]&~m[1712])|(~m[1647]&~m[1708]&~m[1709]&~m[1711]&m[1712])|(m[1647]&~m[1708]&~m[1709]&~m[1711]&m[1712])|(m[1647]&m[1708]&~m[1709]&~m[1711]&m[1712])|(m[1647]&~m[1708]&m[1709]&~m[1711]&m[1712])|(~m[1647]&~m[1708]&~m[1709]&m[1711]&m[1712])|(m[1647]&~m[1708]&~m[1709]&m[1711]&m[1712])|(~m[1647]&m[1708]&~m[1709]&m[1711]&m[1712])|(m[1647]&m[1708]&~m[1709]&m[1711]&m[1712])|(~m[1647]&~m[1708]&m[1709]&m[1711]&m[1712])|(m[1647]&~m[1708]&m[1709]&m[1711]&m[1712])|(m[1647]&m[1708]&m[1709]&m[1711]&m[1712]));
    m[1715] = (((m[1652]&~m[1713]&~m[1714]&~m[1716]&~m[1717])|(~m[1652]&~m[1713]&~m[1714]&m[1716]&~m[1717])|(m[1652]&m[1713]&~m[1714]&m[1716]&~m[1717])|(m[1652]&~m[1713]&m[1714]&m[1716]&~m[1717])|(~m[1652]&m[1713]&~m[1714]&~m[1716]&m[1717])|(~m[1652]&~m[1713]&m[1714]&~m[1716]&m[1717])|(m[1652]&m[1713]&m[1714]&~m[1716]&m[1717])|(~m[1652]&m[1713]&m[1714]&m[1716]&m[1717]))&UnbiasedRNG[413])|((m[1652]&~m[1713]&~m[1714]&m[1716]&~m[1717])|(~m[1652]&~m[1713]&~m[1714]&~m[1716]&m[1717])|(m[1652]&~m[1713]&~m[1714]&~m[1716]&m[1717])|(m[1652]&m[1713]&~m[1714]&~m[1716]&m[1717])|(m[1652]&~m[1713]&m[1714]&~m[1716]&m[1717])|(~m[1652]&~m[1713]&~m[1714]&m[1716]&m[1717])|(m[1652]&~m[1713]&~m[1714]&m[1716]&m[1717])|(~m[1652]&m[1713]&~m[1714]&m[1716]&m[1717])|(m[1652]&m[1713]&~m[1714]&m[1716]&m[1717])|(~m[1652]&~m[1713]&m[1714]&m[1716]&m[1717])|(m[1652]&~m[1713]&m[1714]&m[1716]&m[1717])|(m[1652]&m[1713]&m[1714]&m[1716]&m[1717]));
    m[1720] = (((m[1657]&~m[1718]&~m[1719]&~m[1721]&~m[1722])|(~m[1657]&~m[1718]&~m[1719]&m[1721]&~m[1722])|(m[1657]&m[1718]&~m[1719]&m[1721]&~m[1722])|(m[1657]&~m[1718]&m[1719]&m[1721]&~m[1722])|(~m[1657]&m[1718]&~m[1719]&~m[1721]&m[1722])|(~m[1657]&~m[1718]&m[1719]&~m[1721]&m[1722])|(m[1657]&m[1718]&m[1719]&~m[1721]&m[1722])|(~m[1657]&m[1718]&m[1719]&m[1721]&m[1722]))&UnbiasedRNG[414])|((m[1657]&~m[1718]&~m[1719]&m[1721]&~m[1722])|(~m[1657]&~m[1718]&~m[1719]&~m[1721]&m[1722])|(m[1657]&~m[1718]&~m[1719]&~m[1721]&m[1722])|(m[1657]&m[1718]&~m[1719]&~m[1721]&m[1722])|(m[1657]&~m[1718]&m[1719]&~m[1721]&m[1722])|(~m[1657]&~m[1718]&~m[1719]&m[1721]&m[1722])|(m[1657]&~m[1718]&~m[1719]&m[1721]&m[1722])|(~m[1657]&m[1718]&~m[1719]&m[1721]&m[1722])|(m[1657]&m[1718]&~m[1719]&m[1721]&m[1722])|(~m[1657]&~m[1718]&m[1719]&m[1721]&m[1722])|(m[1657]&~m[1718]&m[1719]&m[1721]&m[1722])|(m[1657]&m[1718]&m[1719]&m[1721]&m[1722]));
    m[1725] = (((m[1662]&~m[1723]&~m[1724]&~m[1726]&~m[1727])|(~m[1662]&~m[1723]&~m[1724]&m[1726]&~m[1727])|(m[1662]&m[1723]&~m[1724]&m[1726]&~m[1727])|(m[1662]&~m[1723]&m[1724]&m[1726]&~m[1727])|(~m[1662]&m[1723]&~m[1724]&~m[1726]&m[1727])|(~m[1662]&~m[1723]&m[1724]&~m[1726]&m[1727])|(m[1662]&m[1723]&m[1724]&~m[1726]&m[1727])|(~m[1662]&m[1723]&m[1724]&m[1726]&m[1727]))&UnbiasedRNG[415])|((m[1662]&~m[1723]&~m[1724]&m[1726]&~m[1727])|(~m[1662]&~m[1723]&~m[1724]&~m[1726]&m[1727])|(m[1662]&~m[1723]&~m[1724]&~m[1726]&m[1727])|(m[1662]&m[1723]&~m[1724]&~m[1726]&m[1727])|(m[1662]&~m[1723]&m[1724]&~m[1726]&m[1727])|(~m[1662]&~m[1723]&~m[1724]&m[1726]&m[1727])|(m[1662]&~m[1723]&~m[1724]&m[1726]&m[1727])|(~m[1662]&m[1723]&~m[1724]&m[1726]&m[1727])|(m[1662]&m[1723]&~m[1724]&m[1726]&m[1727])|(~m[1662]&~m[1723]&m[1724]&m[1726]&m[1727])|(m[1662]&~m[1723]&m[1724]&m[1726]&m[1727])|(m[1662]&m[1723]&m[1724]&m[1726]&m[1727]));
    m[1730] = (((m[1667]&~m[1728]&~m[1729]&~m[1731]&~m[1732])|(~m[1667]&~m[1728]&~m[1729]&m[1731]&~m[1732])|(m[1667]&m[1728]&~m[1729]&m[1731]&~m[1732])|(m[1667]&~m[1728]&m[1729]&m[1731]&~m[1732])|(~m[1667]&m[1728]&~m[1729]&~m[1731]&m[1732])|(~m[1667]&~m[1728]&m[1729]&~m[1731]&m[1732])|(m[1667]&m[1728]&m[1729]&~m[1731]&m[1732])|(~m[1667]&m[1728]&m[1729]&m[1731]&m[1732]))&UnbiasedRNG[416])|((m[1667]&~m[1728]&~m[1729]&m[1731]&~m[1732])|(~m[1667]&~m[1728]&~m[1729]&~m[1731]&m[1732])|(m[1667]&~m[1728]&~m[1729]&~m[1731]&m[1732])|(m[1667]&m[1728]&~m[1729]&~m[1731]&m[1732])|(m[1667]&~m[1728]&m[1729]&~m[1731]&m[1732])|(~m[1667]&~m[1728]&~m[1729]&m[1731]&m[1732])|(m[1667]&~m[1728]&~m[1729]&m[1731]&m[1732])|(~m[1667]&m[1728]&~m[1729]&m[1731]&m[1732])|(m[1667]&m[1728]&~m[1729]&m[1731]&m[1732])|(~m[1667]&~m[1728]&m[1729]&m[1731]&m[1732])|(m[1667]&~m[1728]&m[1729]&m[1731]&m[1732])|(m[1667]&m[1728]&m[1729]&m[1731]&m[1732]));
    m[1735] = (((m[1672]&~m[1733]&~m[1734]&~m[1736]&~m[1737])|(~m[1672]&~m[1733]&~m[1734]&m[1736]&~m[1737])|(m[1672]&m[1733]&~m[1734]&m[1736]&~m[1737])|(m[1672]&~m[1733]&m[1734]&m[1736]&~m[1737])|(~m[1672]&m[1733]&~m[1734]&~m[1736]&m[1737])|(~m[1672]&~m[1733]&m[1734]&~m[1736]&m[1737])|(m[1672]&m[1733]&m[1734]&~m[1736]&m[1737])|(~m[1672]&m[1733]&m[1734]&m[1736]&m[1737]))&UnbiasedRNG[417])|((m[1672]&~m[1733]&~m[1734]&m[1736]&~m[1737])|(~m[1672]&~m[1733]&~m[1734]&~m[1736]&m[1737])|(m[1672]&~m[1733]&~m[1734]&~m[1736]&m[1737])|(m[1672]&m[1733]&~m[1734]&~m[1736]&m[1737])|(m[1672]&~m[1733]&m[1734]&~m[1736]&m[1737])|(~m[1672]&~m[1733]&~m[1734]&m[1736]&m[1737])|(m[1672]&~m[1733]&~m[1734]&m[1736]&m[1737])|(~m[1672]&m[1733]&~m[1734]&m[1736]&m[1737])|(m[1672]&m[1733]&~m[1734]&m[1736]&m[1737])|(~m[1672]&~m[1733]&m[1734]&m[1736]&m[1737])|(m[1672]&~m[1733]&m[1734]&m[1736]&m[1737])|(m[1672]&m[1733]&m[1734]&m[1736]&m[1737]));
    m[1740] = (((m[1682]&~m[1738]&~m[1739]&~m[1741]&~m[1742])|(~m[1682]&~m[1738]&~m[1739]&m[1741]&~m[1742])|(m[1682]&m[1738]&~m[1739]&m[1741]&~m[1742])|(m[1682]&~m[1738]&m[1739]&m[1741]&~m[1742])|(~m[1682]&m[1738]&~m[1739]&~m[1741]&m[1742])|(~m[1682]&~m[1738]&m[1739]&~m[1741]&m[1742])|(m[1682]&m[1738]&m[1739]&~m[1741]&m[1742])|(~m[1682]&m[1738]&m[1739]&m[1741]&m[1742]))&UnbiasedRNG[418])|((m[1682]&~m[1738]&~m[1739]&m[1741]&~m[1742])|(~m[1682]&~m[1738]&~m[1739]&~m[1741]&m[1742])|(m[1682]&~m[1738]&~m[1739]&~m[1741]&m[1742])|(m[1682]&m[1738]&~m[1739]&~m[1741]&m[1742])|(m[1682]&~m[1738]&m[1739]&~m[1741]&m[1742])|(~m[1682]&~m[1738]&~m[1739]&m[1741]&m[1742])|(m[1682]&~m[1738]&~m[1739]&m[1741]&m[1742])|(~m[1682]&m[1738]&~m[1739]&m[1741]&m[1742])|(m[1682]&m[1738]&~m[1739]&m[1741]&m[1742])|(~m[1682]&~m[1738]&m[1739]&m[1741]&m[1742])|(m[1682]&~m[1738]&m[1739]&m[1741]&m[1742])|(m[1682]&m[1738]&m[1739]&m[1741]&m[1742]));
    m[1745] = (((m[1687]&~m[1743]&~m[1744]&~m[1746]&~m[1747])|(~m[1687]&~m[1743]&~m[1744]&m[1746]&~m[1747])|(m[1687]&m[1743]&~m[1744]&m[1746]&~m[1747])|(m[1687]&~m[1743]&m[1744]&m[1746]&~m[1747])|(~m[1687]&m[1743]&~m[1744]&~m[1746]&m[1747])|(~m[1687]&~m[1743]&m[1744]&~m[1746]&m[1747])|(m[1687]&m[1743]&m[1744]&~m[1746]&m[1747])|(~m[1687]&m[1743]&m[1744]&m[1746]&m[1747]))&UnbiasedRNG[419])|((m[1687]&~m[1743]&~m[1744]&m[1746]&~m[1747])|(~m[1687]&~m[1743]&~m[1744]&~m[1746]&m[1747])|(m[1687]&~m[1743]&~m[1744]&~m[1746]&m[1747])|(m[1687]&m[1743]&~m[1744]&~m[1746]&m[1747])|(m[1687]&~m[1743]&m[1744]&~m[1746]&m[1747])|(~m[1687]&~m[1743]&~m[1744]&m[1746]&m[1747])|(m[1687]&~m[1743]&~m[1744]&m[1746]&m[1747])|(~m[1687]&m[1743]&~m[1744]&m[1746]&m[1747])|(m[1687]&m[1743]&~m[1744]&m[1746]&m[1747])|(~m[1687]&~m[1743]&m[1744]&m[1746]&m[1747])|(m[1687]&~m[1743]&m[1744]&m[1746]&m[1747])|(m[1687]&m[1743]&m[1744]&m[1746]&m[1747]));
    m[1750] = (((m[1692]&~m[1748]&~m[1749]&~m[1751]&~m[1752])|(~m[1692]&~m[1748]&~m[1749]&m[1751]&~m[1752])|(m[1692]&m[1748]&~m[1749]&m[1751]&~m[1752])|(m[1692]&~m[1748]&m[1749]&m[1751]&~m[1752])|(~m[1692]&m[1748]&~m[1749]&~m[1751]&m[1752])|(~m[1692]&~m[1748]&m[1749]&~m[1751]&m[1752])|(m[1692]&m[1748]&m[1749]&~m[1751]&m[1752])|(~m[1692]&m[1748]&m[1749]&m[1751]&m[1752]))&UnbiasedRNG[420])|((m[1692]&~m[1748]&~m[1749]&m[1751]&~m[1752])|(~m[1692]&~m[1748]&~m[1749]&~m[1751]&m[1752])|(m[1692]&~m[1748]&~m[1749]&~m[1751]&m[1752])|(m[1692]&m[1748]&~m[1749]&~m[1751]&m[1752])|(m[1692]&~m[1748]&m[1749]&~m[1751]&m[1752])|(~m[1692]&~m[1748]&~m[1749]&m[1751]&m[1752])|(m[1692]&~m[1748]&~m[1749]&m[1751]&m[1752])|(~m[1692]&m[1748]&~m[1749]&m[1751]&m[1752])|(m[1692]&m[1748]&~m[1749]&m[1751]&m[1752])|(~m[1692]&~m[1748]&m[1749]&m[1751]&m[1752])|(m[1692]&~m[1748]&m[1749]&m[1751]&m[1752])|(m[1692]&m[1748]&m[1749]&m[1751]&m[1752]));
    m[1755] = (((m[1697]&~m[1753]&~m[1754]&~m[1756]&~m[1757])|(~m[1697]&~m[1753]&~m[1754]&m[1756]&~m[1757])|(m[1697]&m[1753]&~m[1754]&m[1756]&~m[1757])|(m[1697]&~m[1753]&m[1754]&m[1756]&~m[1757])|(~m[1697]&m[1753]&~m[1754]&~m[1756]&m[1757])|(~m[1697]&~m[1753]&m[1754]&~m[1756]&m[1757])|(m[1697]&m[1753]&m[1754]&~m[1756]&m[1757])|(~m[1697]&m[1753]&m[1754]&m[1756]&m[1757]))&UnbiasedRNG[421])|((m[1697]&~m[1753]&~m[1754]&m[1756]&~m[1757])|(~m[1697]&~m[1753]&~m[1754]&~m[1756]&m[1757])|(m[1697]&~m[1753]&~m[1754]&~m[1756]&m[1757])|(m[1697]&m[1753]&~m[1754]&~m[1756]&m[1757])|(m[1697]&~m[1753]&m[1754]&~m[1756]&m[1757])|(~m[1697]&~m[1753]&~m[1754]&m[1756]&m[1757])|(m[1697]&~m[1753]&~m[1754]&m[1756]&m[1757])|(~m[1697]&m[1753]&~m[1754]&m[1756]&m[1757])|(m[1697]&m[1753]&~m[1754]&m[1756]&m[1757])|(~m[1697]&~m[1753]&m[1754]&m[1756]&m[1757])|(m[1697]&~m[1753]&m[1754]&m[1756]&m[1757])|(m[1697]&m[1753]&m[1754]&m[1756]&m[1757]));
    m[1760] = (((m[1702]&~m[1758]&~m[1759]&~m[1761]&~m[1762])|(~m[1702]&~m[1758]&~m[1759]&m[1761]&~m[1762])|(m[1702]&m[1758]&~m[1759]&m[1761]&~m[1762])|(m[1702]&~m[1758]&m[1759]&m[1761]&~m[1762])|(~m[1702]&m[1758]&~m[1759]&~m[1761]&m[1762])|(~m[1702]&~m[1758]&m[1759]&~m[1761]&m[1762])|(m[1702]&m[1758]&m[1759]&~m[1761]&m[1762])|(~m[1702]&m[1758]&m[1759]&m[1761]&m[1762]))&UnbiasedRNG[422])|((m[1702]&~m[1758]&~m[1759]&m[1761]&~m[1762])|(~m[1702]&~m[1758]&~m[1759]&~m[1761]&m[1762])|(m[1702]&~m[1758]&~m[1759]&~m[1761]&m[1762])|(m[1702]&m[1758]&~m[1759]&~m[1761]&m[1762])|(m[1702]&~m[1758]&m[1759]&~m[1761]&m[1762])|(~m[1702]&~m[1758]&~m[1759]&m[1761]&m[1762])|(m[1702]&~m[1758]&~m[1759]&m[1761]&m[1762])|(~m[1702]&m[1758]&~m[1759]&m[1761]&m[1762])|(m[1702]&m[1758]&~m[1759]&m[1761]&m[1762])|(~m[1702]&~m[1758]&m[1759]&m[1761]&m[1762])|(m[1702]&~m[1758]&m[1759]&m[1761]&m[1762])|(m[1702]&m[1758]&m[1759]&m[1761]&m[1762]));
    m[1765] = (((m[1707]&~m[1763]&~m[1764]&~m[1766]&~m[1767])|(~m[1707]&~m[1763]&~m[1764]&m[1766]&~m[1767])|(m[1707]&m[1763]&~m[1764]&m[1766]&~m[1767])|(m[1707]&~m[1763]&m[1764]&m[1766]&~m[1767])|(~m[1707]&m[1763]&~m[1764]&~m[1766]&m[1767])|(~m[1707]&~m[1763]&m[1764]&~m[1766]&m[1767])|(m[1707]&m[1763]&m[1764]&~m[1766]&m[1767])|(~m[1707]&m[1763]&m[1764]&m[1766]&m[1767]))&UnbiasedRNG[423])|((m[1707]&~m[1763]&~m[1764]&m[1766]&~m[1767])|(~m[1707]&~m[1763]&~m[1764]&~m[1766]&m[1767])|(m[1707]&~m[1763]&~m[1764]&~m[1766]&m[1767])|(m[1707]&m[1763]&~m[1764]&~m[1766]&m[1767])|(m[1707]&~m[1763]&m[1764]&~m[1766]&m[1767])|(~m[1707]&~m[1763]&~m[1764]&m[1766]&m[1767])|(m[1707]&~m[1763]&~m[1764]&m[1766]&m[1767])|(~m[1707]&m[1763]&~m[1764]&m[1766]&m[1767])|(m[1707]&m[1763]&~m[1764]&m[1766]&m[1767])|(~m[1707]&~m[1763]&m[1764]&m[1766]&m[1767])|(m[1707]&~m[1763]&m[1764]&m[1766]&m[1767])|(m[1707]&m[1763]&m[1764]&m[1766]&m[1767]));
    m[1770] = (((m[1712]&~m[1768]&~m[1769]&~m[1771]&~m[1772])|(~m[1712]&~m[1768]&~m[1769]&m[1771]&~m[1772])|(m[1712]&m[1768]&~m[1769]&m[1771]&~m[1772])|(m[1712]&~m[1768]&m[1769]&m[1771]&~m[1772])|(~m[1712]&m[1768]&~m[1769]&~m[1771]&m[1772])|(~m[1712]&~m[1768]&m[1769]&~m[1771]&m[1772])|(m[1712]&m[1768]&m[1769]&~m[1771]&m[1772])|(~m[1712]&m[1768]&m[1769]&m[1771]&m[1772]))&UnbiasedRNG[424])|((m[1712]&~m[1768]&~m[1769]&m[1771]&~m[1772])|(~m[1712]&~m[1768]&~m[1769]&~m[1771]&m[1772])|(m[1712]&~m[1768]&~m[1769]&~m[1771]&m[1772])|(m[1712]&m[1768]&~m[1769]&~m[1771]&m[1772])|(m[1712]&~m[1768]&m[1769]&~m[1771]&m[1772])|(~m[1712]&~m[1768]&~m[1769]&m[1771]&m[1772])|(m[1712]&~m[1768]&~m[1769]&m[1771]&m[1772])|(~m[1712]&m[1768]&~m[1769]&m[1771]&m[1772])|(m[1712]&m[1768]&~m[1769]&m[1771]&m[1772])|(~m[1712]&~m[1768]&m[1769]&m[1771]&m[1772])|(m[1712]&~m[1768]&m[1769]&m[1771]&m[1772])|(m[1712]&m[1768]&m[1769]&m[1771]&m[1772]));
    m[1775] = (((m[1717]&~m[1773]&~m[1774]&~m[1776]&~m[1777])|(~m[1717]&~m[1773]&~m[1774]&m[1776]&~m[1777])|(m[1717]&m[1773]&~m[1774]&m[1776]&~m[1777])|(m[1717]&~m[1773]&m[1774]&m[1776]&~m[1777])|(~m[1717]&m[1773]&~m[1774]&~m[1776]&m[1777])|(~m[1717]&~m[1773]&m[1774]&~m[1776]&m[1777])|(m[1717]&m[1773]&m[1774]&~m[1776]&m[1777])|(~m[1717]&m[1773]&m[1774]&m[1776]&m[1777]))&UnbiasedRNG[425])|((m[1717]&~m[1773]&~m[1774]&m[1776]&~m[1777])|(~m[1717]&~m[1773]&~m[1774]&~m[1776]&m[1777])|(m[1717]&~m[1773]&~m[1774]&~m[1776]&m[1777])|(m[1717]&m[1773]&~m[1774]&~m[1776]&m[1777])|(m[1717]&~m[1773]&m[1774]&~m[1776]&m[1777])|(~m[1717]&~m[1773]&~m[1774]&m[1776]&m[1777])|(m[1717]&~m[1773]&~m[1774]&m[1776]&m[1777])|(~m[1717]&m[1773]&~m[1774]&m[1776]&m[1777])|(m[1717]&m[1773]&~m[1774]&m[1776]&m[1777])|(~m[1717]&~m[1773]&m[1774]&m[1776]&m[1777])|(m[1717]&~m[1773]&m[1774]&m[1776]&m[1777])|(m[1717]&m[1773]&m[1774]&m[1776]&m[1777]));
    m[1780] = (((m[1722]&~m[1778]&~m[1779]&~m[1781]&~m[1782])|(~m[1722]&~m[1778]&~m[1779]&m[1781]&~m[1782])|(m[1722]&m[1778]&~m[1779]&m[1781]&~m[1782])|(m[1722]&~m[1778]&m[1779]&m[1781]&~m[1782])|(~m[1722]&m[1778]&~m[1779]&~m[1781]&m[1782])|(~m[1722]&~m[1778]&m[1779]&~m[1781]&m[1782])|(m[1722]&m[1778]&m[1779]&~m[1781]&m[1782])|(~m[1722]&m[1778]&m[1779]&m[1781]&m[1782]))&UnbiasedRNG[426])|((m[1722]&~m[1778]&~m[1779]&m[1781]&~m[1782])|(~m[1722]&~m[1778]&~m[1779]&~m[1781]&m[1782])|(m[1722]&~m[1778]&~m[1779]&~m[1781]&m[1782])|(m[1722]&m[1778]&~m[1779]&~m[1781]&m[1782])|(m[1722]&~m[1778]&m[1779]&~m[1781]&m[1782])|(~m[1722]&~m[1778]&~m[1779]&m[1781]&m[1782])|(m[1722]&~m[1778]&~m[1779]&m[1781]&m[1782])|(~m[1722]&m[1778]&~m[1779]&m[1781]&m[1782])|(m[1722]&m[1778]&~m[1779]&m[1781]&m[1782])|(~m[1722]&~m[1778]&m[1779]&m[1781]&m[1782])|(m[1722]&~m[1778]&m[1779]&m[1781]&m[1782])|(m[1722]&m[1778]&m[1779]&m[1781]&m[1782]));
    m[1785] = (((m[1727]&~m[1783]&~m[1784]&~m[1786]&~m[1787])|(~m[1727]&~m[1783]&~m[1784]&m[1786]&~m[1787])|(m[1727]&m[1783]&~m[1784]&m[1786]&~m[1787])|(m[1727]&~m[1783]&m[1784]&m[1786]&~m[1787])|(~m[1727]&m[1783]&~m[1784]&~m[1786]&m[1787])|(~m[1727]&~m[1783]&m[1784]&~m[1786]&m[1787])|(m[1727]&m[1783]&m[1784]&~m[1786]&m[1787])|(~m[1727]&m[1783]&m[1784]&m[1786]&m[1787]))&UnbiasedRNG[427])|((m[1727]&~m[1783]&~m[1784]&m[1786]&~m[1787])|(~m[1727]&~m[1783]&~m[1784]&~m[1786]&m[1787])|(m[1727]&~m[1783]&~m[1784]&~m[1786]&m[1787])|(m[1727]&m[1783]&~m[1784]&~m[1786]&m[1787])|(m[1727]&~m[1783]&m[1784]&~m[1786]&m[1787])|(~m[1727]&~m[1783]&~m[1784]&m[1786]&m[1787])|(m[1727]&~m[1783]&~m[1784]&m[1786]&m[1787])|(~m[1727]&m[1783]&~m[1784]&m[1786]&m[1787])|(m[1727]&m[1783]&~m[1784]&m[1786]&m[1787])|(~m[1727]&~m[1783]&m[1784]&m[1786]&m[1787])|(m[1727]&~m[1783]&m[1784]&m[1786]&m[1787])|(m[1727]&m[1783]&m[1784]&m[1786]&m[1787]));
    m[1790] = (((m[1732]&~m[1788]&~m[1789]&~m[1791]&~m[1792])|(~m[1732]&~m[1788]&~m[1789]&m[1791]&~m[1792])|(m[1732]&m[1788]&~m[1789]&m[1791]&~m[1792])|(m[1732]&~m[1788]&m[1789]&m[1791]&~m[1792])|(~m[1732]&m[1788]&~m[1789]&~m[1791]&m[1792])|(~m[1732]&~m[1788]&m[1789]&~m[1791]&m[1792])|(m[1732]&m[1788]&m[1789]&~m[1791]&m[1792])|(~m[1732]&m[1788]&m[1789]&m[1791]&m[1792]))&UnbiasedRNG[428])|((m[1732]&~m[1788]&~m[1789]&m[1791]&~m[1792])|(~m[1732]&~m[1788]&~m[1789]&~m[1791]&m[1792])|(m[1732]&~m[1788]&~m[1789]&~m[1791]&m[1792])|(m[1732]&m[1788]&~m[1789]&~m[1791]&m[1792])|(m[1732]&~m[1788]&m[1789]&~m[1791]&m[1792])|(~m[1732]&~m[1788]&~m[1789]&m[1791]&m[1792])|(m[1732]&~m[1788]&~m[1789]&m[1791]&m[1792])|(~m[1732]&m[1788]&~m[1789]&m[1791]&m[1792])|(m[1732]&m[1788]&~m[1789]&m[1791]&m[1792])|(~m[1732]&~m[1788]&m[1789]&m[1791]&m[1792])|(m[1732]&~m[1788]&m[1789]&m[1791]&m[1792])|(m[1732]&m[1788]&m[1789]&m[1791]&m[1792]));
    m[1795] = (((m[1737]&~m[1793]&~m[1794]&~m[1796]&~m[1797])|(~m[1737]&~m[1793]&~m[1794]&m[1796]&~m[1797])|(m[1737]&m[1793]&~m[1794]&m[1796]&~m[1797])|(m[1737]&~m[1793]&m[1794]&m[1796]&~m[1797])|(~m[1737]&m[1793]&~m[1794]&~m[1796]&m[1797])|(~m[1737]&~m[1793]&m[1794]&~m[1796]&m[1797])|(m[1737]&m[1793]&m[1794]&~m[1796]&m[1797])|(~m[1737]&m[1793]&m[1794]&m[1796]&m[1797]))&UnbiasedRNG[429])|((m[1737]&~m[1793]&~m[1794]&m[1796]&~m[1797])|(~m[1737]&~m[1793]&~m[1794]&~m[1796]&m[1797])|(m[1737]&~m[1793]&~m[1794]&~m[1796]&m[1797])|(m[1737]&m[1793]&~m[1794]&~m[1796]&m[1797])|(m[1737]&~m[1793]&m[1794]&~m[1796]&m[1797])|(~m[1737]&~m[1793]&~m[1794]&m[1796]&m[1797])|(m[1737]&~m[1793]&~m[1794]&m[1796]&m[1797])|(~m[1737]&m[1793]&~m[1794]&m[1796]&m[1797])|(m[1737]&m[1793]&~m[1794]&m[1796]&m[1797])|(~m[1737]&~m[1793]&m[1794]&m[1796]&m[1797])|(m[1737]&~m[1793]&m[1794]&m[1796]&m[1797])|(m[1737]&m[1793]&m[1794]&m[1796]&m[1797]));
    m[1800] = (((m[1747]&~m[1798]&~m[1799]&~m[1801]&~m[1802])|(~m[1747]&~m[1798]&~m[1799]&m[1801]&~m[1802])|(m[1747]&m[1798]&~m[1799]&m[1801]&~m[1802])|(m[1747]&~m[1798]&m[1799]&m[1801]&~m[1802])|(~m[1747]&m[1798]&~m[1799]&~m[1801]&m[1802])|(~m[1747]&~m[1798]&m[1799]&~m[1801]&m[1802])|(m[1747]&m[1798]&m[1799]&~m[1801]&m[1802])|(~m[1747]&m[1798]&m[1799]&m[1801]&m[1802]))&UnbiasedRNG[430])|((m[1747]&~m[1798]&~m[1799]&m[1801]&~m[1802])|(~m[1747]&~m[1798]&~m[1799]&~m[1801]&m[1802])|(m[1747]&~m[1798]&~m[1799]&~m[1801]&m[1802])|(m[1747]&m[1798]&~m[1799]&~m[1801]&m[1802])|(m[1747]&~m[1798]&m[1799]&~m[1801]&m[1802])|(~m[1747]&~m[1798]&~m[1799]&m[1801]&m[1802])|(m[1747]&~m[1798]&~m[1799]&m[1801]&m[1802])|(~m[1747]&m[1798]&~m[1799]&m[1801]&m[1802])|(m[1747]&m[1798]&~m[1799]&m[1801]&m[1802])|(~m[1747]&~m[1798]&m[1799]&m[1801]&m[1802])|(m[1747]&~m[1798]&m[1799]&m[1801]&m[1802])|(m[1747]&m[1798]&m[1799]&m[1801]&m[1802]));
    m[1805] = (((m[1752]&~m[1803]&~m[1804]&~m[1806]&~m[1807])|(~m[1752]&~m[1803]&~m[1804]&m[1806]&~m[1807])|(m[1752]&m[1803]&~m[1804]&m[1806]&~m[1807])|(m[1752]&~m[1803]&m[1804]&m[1806]&~m[1807])|(~m[1752]&m[1803]&~m[1804]&~m[1806]&m[1807])|(~m[1752]&~m[1803]&m[1804]&~m[1806]&m[1807])|(m[1752]&m[1803]&m[1804]&~m[1806]&m[1807])|(~m[1752]&m[1803]&m[1804]&m[1806]&m[1807]))&UnbiasedRNG[431])|((m[1752]&~m[1803]&~m[1804]&m[1806]&~m[1807])|(~m[1752]&~m[1803]&~m[1804]&~m[1806]&m[1807])|(m[1752]&~m[1803]&~m[1804]&~m[1806]&m[1807])|(m[1752]&m[1803]&~m[1804]&~m[1806]&m[1807])|(m[1752]&~m[1803]&m[1804]&~m[1806]&m[1807])|(~m[1752]&~m[1803]&~m[1804]&m[1806]&m[1807])|(m[1752]&~m[1803]&~m[1804]&m[1806]&m[1807])|(~m[1752]&m[1803]&~m[1804]&m[1806]&m[1807])|(m[1752]&m[1803]&~m[1804]&m[1806]&m[1807])|(~m[1752]&~m[1803]&m[1804]&m[1806]&m[1807])|(m[1752]&~m[1803]&m[1804]&m[1806]&m[1807])|(m[1752]&m[1803]&m[1804]&m[1806]&m[1807]));
    m[1810] = (((m[1757]&~m[1808]&~m[1809]&~m[1811]&~m[1812])|(~m[1757]&~m[1808]&~m[1809]&m[1811]&~m[1812])|(m[1757]&m[1808]&~m[1809]&m[1811]&~m[1812])|(m[1757]&~m[1808]&m[1809]&m[1811]&~m[1812])|(~m[1757]&m[1808]&~m[1809]&~m[1811]&m[1812])|(~m[1757]&~m[1808]&m[1809]&~m[1811]&m[1812])|(m[1757]&m[1808]&m[1809]&~m[1811]&m[1812])|(~m[1757]&m[1808]&m[1809]&m[1811]&m[1812]))&UnbiasedRNG[432])|((m[1757]&~m[1808]&~m[1809]&m[1811]&~m[1812])|(~m[1757]&~m[1808]&~m[1809]&~m[1811]&m[1812])|(m[1757]&~m[1808]&~m[1809]&~m[1811]&m[1812])|(m[1757]&m[1808]&~m[1809]&~m[1811]&m[1812])|(m[1757]&~m[1808]&m[1809]&~m[1811]&m[1812])|(~m[1757]&~m[1808]&~m[1809]&m[1811]&m[1812])|(m[1757]&~m[1808]&~m[1809]&m[1811]&m[1812])|(~m[1757]&m[1808]&~m[1809]&m[1811]&m[1812])|(m[1757]&m[1808]&~m[1809]&m[1811]&m[1812])|(~m[1757]&~m[1808]&m[1809]&m[1811]&m[1812])|(m[1757]&~m[1808]&m[1809]&m[1811]&m[1812])|(m[1757]&m[1808]&m[1809]&m[1811]&m[1812]));
    m[1815] = (((m[1762]&~m[1813]&~m[1814]&~m[1816]&~m[1817])|(~m[1762]&~m[1813]&~m[1814]&m[1816]&~m[1817])|(m[1762]&m[1813]&~m[1814]&m[1816]&~m[1817])|(m[1762]&~m[1813]&m[1814]&m[1816]&~m[1817])|(~m[1762]&m[1813]&~m[1814]&~m[1816]&m[1817])|(~m[1762]&~m[1813]&m[1814]&~m[1816]&m[1817])|(m[1762]&m[1813]&m[1814]&~m[1816]&m[1817])|(~m[1762]&m[1813]&m[1814]&m[1816]&m[1817]))&UnbiasedRNG[433])|((m[1762]&~m[1813]&~m[1814]&m[1816]&~m[1817])|(~m[1762]&~m[1813]&~m[1814]&~m[1816]&m[1817])|(m[1762]&~m[1813]&~m[1814]&~m[1816]&m[1817])|(m[1762]&m[1813]&~m[1814]&~m[1816]&m[1817])|(m[1762]&~m[1813]&m[1814]&~m[1816]&m[1817])|(~m[1762]&~m[1813]&~m[1814]&m[1816]&m[1817])|(m[1762]&~m[1813]&~m[1814]&m[1816]&m[1817])|(~m[1762]&m[1813]&~m[1814]&m[1816]&m[1817])|(m[1762]&m[1813]&~m[1814]&m[1816]&m[1817])|(~m[1762]&~m[1813]&m[1814]&m[1816]&m[1817])|(m[1762]&~m[1813]&m[1814]&m[1816]&m[1817])|(m[1762]&m[1813]&m[1814]&m[1816]&m[1817]));
    m[1820] = (((m[1767]&~m[1818]&~m[1819]&~m[1821]&~m[1822])|(~m[1767]&~m[1818]&~m[1819]&m[1821]&~m[1822])|(m[1767]&m[1818]&~m[1819]&m[1821]&~m[1822])|(m[1767]&~m[1818]&m[1819]&m[1821]&~m[1822])|(~m[1767]&m[1818]&~m[1819]&~m[1821]&m[1822])|(~m[1767]&~m[1818]&m[1819]&~m[1821]&m[1822])|(m[1767]&m[1818]&m[1819]&~m[1821]&m[1822])|(~m[1767]&m[1818]&m[1819]&m[1821]&m[1822]))&UnbiasedRNG[434])|((m[1767]&~m[1818]&~m[1819]&m[1821]&~m[1822])|(~m[1767]&~m[1818]&~m[1819]&~m[1821]&m[1822])|(m[1767]&~m[1818]&~m[1819]&~m[1821]&m[1822])|(m[1767]&m[1818]&~m[1819]&~m[1821]&m[1822])|(m[1767]&~m[1818]&m[1819]&~m[1821]&m[1822])|(~m[1767]&~m[1818]&~m[1819]&m[1821]&m[1822])|(m[1767]&~m[1818]&~m[1819]&m[1821]&m[1822])|(~m[1767]&m[1818]&~m[1819]&m[1821]&m[1822])|(m[1767]&m[1818]&~m[1819]&m[1821]&m[1822])|(~m[1767]&~m[1818]&m[1819]&m[1821]&m[1822])|(m[1767]&~m[1818]&m[1819]&m[1821]&m[1822])|(m[1767]&m[1818]&m[1819]&m[1821]&m[1822]));
    m[1825] = (((m[1772]&~m[1823]&~m[1824]&~m[1826]&~m[1827])|(~m[1772]&~m[1823]&~m[1824]&m[1826]&~m[1827])|(m[1772]&m[1823]&~m[1824]&m[1826]&~m[1827])|(m[1772]&~m[1823]&m[1824]&m[1826]&~m[1827])|(~m[1772]&m[1823]&~m[1824]&~m[1826]&m[1827])|(~m[1772]&~m[1823]&m[1824]&~m[1826]&m[1827])|(m[1772]&m[1823]&m[1824]&~m[1826]&m[1827])|(~m[1772]&m[1823]&m[1824]&m[1826]&m[1827]))&UnbiasedRNG[435])|((m[1772]&~m[1823]&~m[1824]&m[1826]&~m[1827])|(~m[1772]&~m[1823]&~m[1824]&~m[1826]&m[1827])|(m[1772]&~m[1823]&~m[1824]&~m[1826]&m[1827])|(m[1772]&m[1823]&~m[1824]&~m[1826]&m[1827])|(m[1772]&~m[1823]&m[1824]&~m[1826]&m[1827])|(~m[1772]&~m[1823]&~m[1824]&m[1826]&m[1827])|(m[1772]&~m[1823]&~m[1824]&m[1826]&m[1827])|(~m[1772]&m[1823]&~m[1824]&m[1826]&m[1827])|(m[1772]&m[1823]&~m[1824]&m[1826]&m[1827])|(~m[1772]&~m[1823]&m[1824]&m[1826]&m[1827])|(m[1772]&~m[1823]&m[1824]&m[1826]&m[1827])|(m[1772]&m[1823]&m[1824]&m[1826]&m[1827]));
    m[1830] = (((m[1777]&~m[1828]&~m[1829]&~m[1831]&~m[1832])|(~m[1777]&~m[1828]&~m[1829]&m[1831]&~m[1832])|(m[1777]&m[1828]&~m[1829]&m[1831]&~m[1832])|(m[1777]&~m[1828]&m[1829]&m[1831]&~m[1832])|(~m[1777]&m[1828]&~m[1829]&~m[1831]&m[1832])|(~m[1777]&~m[1828]&m[1829]&~m[1831]&m[1832])|(m[1777]&m[1828]&m[1829]&~m[1831]&m[1832])|(~m[1777]&m[1828]&m[1829]&m[1831]&m[1832]))&UnbiasedRNG[436])|((m[1777]&~m[1828]&~m[1829]&m[1831]&~m[1832])|(~m[1777]&~m[1828]&~m[1829]&~m[1831]&m[1832])|(m[1777]&~m[1828]&~m[1829]&~m[1831]&m[1832])|(m[1777]&m[1828]&~m[1829]&~m[1831]&m[1832])|(m[1777]&~m[1828]&m[1829]&~m[1831]&m[1832])|(~m[1777]&~m[1828]&~m[1829]&m[1831]&m[1832])|(m[1777]&~m[1828]&~m[1829]&m[1831]&m[1832])|(~m[1777]&m[1828]&~m[1829]&m[1831]&m[1832])|(m[1777]&m[1828]&~m[1829]&m[1831]&m[1832])|(~m[1777]&~m[1828]&m[1829]&m[1831]&m[1832])|(m[1777]&~m[1828]&m[1829]&m[1831]&m[1832])|(m[1777]&m[1828]&m[1829]&m[1831]&m[1832]));
    m[1835] = (((m[1782]&~m[1833]&~m[1834]&~m[1836]&~m[1837])|(~m[1782]&~m[1833]&~m[1834]&m[1836]&~m[1837])|(m[1782]&m[1833]&~m[1834]&m[1836]&~m[1837])|(m[1782]&~m[1833]&m[1834]&m[1836]&~m[1837])|(~m[1782]&m[1833]&~m[1834]&~m[1836]&m[1837])|(~m[1782]&~m[1833]&m[1834]&~m[1836]&m[1837])|(m[1782]&m[1833]&m[1834]&~m[1836]&m[1837])|(~m[1782]&m[1833]&m[1834]&m[1836]&m[1837]))&UnbiasedRNG[437])|((m[1782]&~m[1833]&~m[1834]&m[1836]&~m[1837])|(~m[1782]&~m[1833]&~m[1834]&~m[1836]&m[1837])|(m[1782]&~m[1833]&~m[1834]&~m[1836]&m[1837])|(m[1782]&m[1833]&~m[1834]&~m[1836]&m[1837])|(m[1782]&~m[1833]&m[1834]&~m[1836]&m[1837])|(~m[1782]&~m[1833]&~m[1834]&m[1836]&m[1837])|(m[1782]&~m[1833]&~m[1834]&m[1836]&m[1837])|(~m[1782]&m[1833]&~m[1834]&m[1836]&m[1837])|(m[1782]&m[1833]&~m[1834]&m[1836]&m[1837])|(~m[1782]&~m[1833]&m[1834]&m[1836]&m[1837])|(m[1782]&~m[1833]&m[1834]&m[1836]&m[1837])|(m[1782]&m[1833]&m[1834]&m[1836]&m[1837]));
    m[1840] = (((m[1787]&~m[1838]&~m[1839]&~m[1841]&~m[1842])|(~m[1787]&~m[1838]&~m[1839]&m[1841]&~m[1842])|(m[1787]&m[1838]&~m[1839]&m[1841]&~m[1842])|(m[1787]&~m[1838]&m[1839]&m[1841]&~m[1842])|(~m[1787]&m[1838]&~m[1839]&~m[1841]&m[1842])|(~m[1787]&~m[1838]&m[1839]&~m[1841]&m[1842])|(m[1787]&m[1838]&m[1839]&~m[1841]&m[1842])|(~m[1787]&m[1838]&m[1839]&m[1841]&m[1842]))&UnbiasedRNG[438])|((m[1787]&~m[1838]&~m[1839]&m[1841]&~m[1842])|(~m[1787]&~m[1838]&~m[1839]&~m[1841]&m[1842])|(m[1787]&~m[1838]&~m[1839]&~m[1841]&m[1842])|(m[1787]&m[1838]&~m[1839]&~m[1841]&m[1842])|(m[1787]&~m[1838]&m[1839]&~m[1841]&m[1842])|(~m[1787]&~m[1838]&~m[1839]&m[1841]&m[1842])|(m[1787]&~m[1838]&~m[1839]&m[1841]&m[1842])|(~m[1787]&m[1838]&~m[1839]&m[1841]&m[1842])|(m[1787]&m[1838]&~m[1839]&m[1841]&m[1842])|(~m[1787]&~m[1838]&m[1839]&m[1841]&m[1842])|(m[1787]&~m[1838]&m[1839]&m[1841]&m[1842])|(m[1787]&m[1838]&m[1839]&m[1841]&m[1842]));
    m[1845] = (((m[1792]&~m[1843]&~m[1844]&~m[1846]&~m[1847])|(~m[1792]&~m[1843]&~m[1844]&m[1846]&~m[1847])|(m[1792]&m[1843]&~m[1844]&m[1846]&~m[1847])|(m[1792]&~m[1843]&m[1844]&m[1846]&~m[1847])|(~m[1792]&m[1843]&~m[1844]&~m[1846]&m[1847])|(~m[1792]&~m[1843]&m[1844]&~m[1846]&m[1847])|(m[1792]&m[1843]&m[1844]&~m[1846]&m[1847])|(~m[1792]&m[1843]&m[1844]&m[1846]&m[1847]))&UnbiasedRNG[439])|((m[1792]&~m[1843]&~m[1844]&m[1846]&~m[1847])|(~m[1792]&~m[1843]&~m[1844]&~m[1846]&m[1847])|(m[1792]&~m[1843]&~m[1844]&~m[1846]&m[1847])|(m[1792]&m[1843]&~m[1844]&~m[1846]&m[1847])|(m[1792]&~m[1843]&m[1844]&~m[1846]&m[1847])|(~m[1792]&~m[1843]&~m[1844]&m[1846]&m[1847])|(m[1792]&~m[1843]&~m[1844]&m[1846]&m[1847])|(~m[1792]&m[1843]&~m[1844]&m[1846]&m[1847])|(m[1792]&m[1843]&~m[1844]&m[1846]&m[1847])|(~m[1792]&~m[1843]&m[1844]&m[1846]&m[1847])|(m[1792]&~m[1843]&m[1844]&m[1846]&m[1847])|(m[1792]&m[1843]&m[1844]&m[1846]&m[1847]));
    m[1850] = (((m[1797]&~m[1848]&~m[1849]&~m[1851]&~m[1852])|(~m[1797]&~m[1848]&~m[1849]&m[1851]&~m[1852])|(m[1797]&m[1848]&~m[1849]&m[1851]&~m[1852])|(m[1797]&~m[1848]&m[1849]&m[1851]&~m[1852])|(~m[1797]&m[1848]&~m[1849]&~m[1851]&m[1852])|(~m[1797]&~m[1848]&m[1849]&~m[1851]&m[1852])|(m[1797]&m[1848]&m[1849]&~m[1851]&m[1852])|(~m[1797]&m[1848]&m[1849]&m[1851]&m[1852]))&UnbiasedRNG[440])|((m[1797]&~m[1848]&~m[1849]&m[1851]&~m[1852])|(~m[1797]&~m[1848]&~m[1849]&~m[1851]&m[1852])|(m[1797]&~m[1848]&~m[1849]&~m[1851]&m[1852])|(m[1797]&m[1848]&~m[1849]&~m[1851]&m[1852])|(m[1797]&~m[1848]&m[1849]&~m[1851]&m[1852])|(~m[1797]&~m[1848]&~m[1849]&m[1851]&m[1852])|(m[1797]&~m[1848]&~m[1849]&m[1851]&m[1852])|(~m[1797]&m[1848]&~m[1849]&m[1851]&m[1852])|(m[1797]&m[1848]&~m[1849]&m[1851]&m[1852])|(~m[1797]&~m[1848]&m[1849]&m[1851]&m[1852])|(m[1797]&~m[1848]&m[1849]&m[1851]&m[1852])|(m[1797]&m[1848]&m[1849]&m[1851]&m[1852]));
    m[1855] = (((m[1807]&~m[1853]&~m[1854]&~m[1856]&~m[1857])|(~m[1807]&~m[1853]&~m[1854]&m[1856]&~m[1857])|(m[1807]&m[1853]&~m[1854]&m[1856]&~m[1857])|(m[1807]&~m[1853]&m[1854]&m[1856]&~m[1857])|(~m[1807]&m[1853]&~m[1854]&~m[1856]&m[1857])|(~m[1807]&~m[1853]&m[1854]&~m[1856]&m[1857])|(m[1807]&m[1853]&m[1854]&~m[1856]&m[1857])|(~m[1807]&m[1853]&m[1854]&m[1856]&m[1857]))&UnbiasedRNG[441])|((m[1807]&~m[1853]&~m[1854]&m[1856]&~m[1857])|(~m[1807]&~m[1853]&~m[1854]&~m[1856]&m[1857])|(m[1807]&~m[1853]&~m[1854]&~m[1856]&m[1857])|(m[1807]&m[1853]&~m[1854]&~m[1856]&m[1857])|(m[1807]&~m[1853]&m[1854]&~m[1856]&m[1857])|(~m[1807]&~m[1853]&~m[1854]&m[1856]&m[1857])|(m[1807]&~m[1853]&~m[1854]&m[1856]&m[1857])|(~m[1807]&m[1853]&~m[1854]&m[1856]&m[1857])|(m[1807]&m[1853]&~m[1854]&m[1856]&m[1857])|(~m[1807]&~m[1853]&m[1854]&m[1856]&m[1857])|(m[1807]&~m[1853]&m[1854]&m[1856]&m[1857])|(m[1807]&m[1853]&m[1854]&m[1856]&m[1857]));
    m[1860] = (((m[1812]&~m[1858]&~m[1859]&~m[1861]&~m[1862])|(~m[1812]&~m[1858]&~m[1859]&m[1861]&~m[1862])|(m[1812]&m[1858]&~m[1859]&m[1861]&~m[1862])|(m[1812]&~m[1858]&m[1859]&m[1861]&~m[1862])|(~m[1812]&m[1858]&~m[1859]&~m[1861]&m[1862])|(~m[1812]&~m[1858]&m[1859]&~m[1861]&m[1862])|(m[1812]&m[1858]&m[1859]&~m[1861]&m[1862])|(~m[1812]&m[1858]&m[1859]&m[1861]&m[1862]))&UnbiasedRNG[442])|((m[1812]&~m[1858]&~m[1859]&m[1861]&~m[1862])|(~m[1812]&~m[1858]&~m[1859]&~m[1861]&m[1862])|(m[1812]&~m[1858]&~m[1859]&~m[1861]&m[1862])|(m[1812]&m[1858]&~m[1859]&~m[1861]&m[1862])|(m[1812]&~m[1858]&m[1859]&~m[1861]&m[1862])|(~m[1812]&~m[1858]&~m[1859]&m[1861]&m[1862])|(m[1812]&~m[1858]&~m[1859]&m[1861]&m[1862])|(~m[1812]&m[1858]&~m[1859]&m[1861]&m[1862])|(m[1812]&m[1858]&~m[1859]&m[1861]&m[1862])|(~m[1812]&~m[1858]&m[1859]&m[1861]&m[1862])|(m[1812]&~m[1858]&m[1859]&m[1861]&m[1862])|(m[1812]&m[1858]&m[1859]&m[1861]&m[1862]));
    m[1865] = (((m[1817]&~m[1863]&~m[1864]&~m[1866]&~m[1867])|(~m[1817]&~m[1863]&~m[1864]&m[1866]&~m[1867])|(m[1817]&m[1863]&~m[1864]&m[1866]&~m[1867])|(m[1817]&~m[1863]&m[1864]&m[1866]&~m[1867])|(~m[1817]&m[1863]&~m[1864]&~m[1866]&m[1867])|(~m[1817]&~m[1863]&m[1864]&~m[1866]&m[1867])|(m[1817]&m[1863]&m[1864]&~m[1866]&m[1867])|(~m[1817]&m[1863]&m[1864]&m[1866]&m[1867]))&UnbiasedRNG[443])|((m[1817]&~m[1863]&~m[1864]&m[1866]&~m[1867])|(~m[1817]&~m[1863]&~m[1864]&~m[1866]&m[1867])|(m[1817]&~m[1863]&~m[1864]&~m[1866]&m[1867])|(m[1817]&m[1863]&~m[1864]&~m[1866]&m[1867])|(m[1817]&~m[1863]&m[1864]&~m[1866]&m[1867])|(~m[1817]&~m[1863]&~m[1864]&m[1866]&m[1867])|(m[1817]&~m[1863]&~m[1864]&m[1866]&m[1867])|(~m[1817]&m[1863]&~m[1864]&m[1866]&m[1867])|(m[1817]&m[1863]&~m[1864]&m[1866]&m[1867])|(~m[1817]&~m[1863]&m[1864]&m[1866]&m[1867])|(m[1817]&~m[1863]&m[1864]&m[1866]&m[1867])|(m[1817]&m[1863]&m[1864]&m[1866]&m[1867]));
    m[1870] = (((m[1822]&~m[1868]&~m[1869]&~m[1871]&~m[1872])|(~m[1822]&~m[1868]&~m[1869]&m[1871]&~m[1872])|(m[1822]&m[1868]&~m[1869]&m[1871]&~m[1872])|(m[1822]&~m[1868]&m[1869]&m[1871]&~m[1872])|(~m[1822]&m[1868]&~m[1869]&~m[1871]&m[1872])|(~m[1822]&~m[1868]&m[1869]&~m[1871]&m[1872])|(m[1822]&m[1868]&m[1869]&~m[1871]&m[1872])|(~m[1822]&m[1868]&m[1869]&m[1871]&m[1872]))&UnbiasedRNG[444])|((m[1822]&~m[1868]&~m[1869]&m[1871]&~m[1872])|(~m[1822]&~m[1868]&~m[1869]&~m[1871]&m[1872])|(m[1822]&~m[1868]&~m[1869]&~m[1871]&m[1872])|(m[1822]&m[1868]&~m[1869]&~m[1871]&m[1872])|(m[1822]&~m[1868]&m[1869]&~m[1871]&m[1872])|(~m[1822]&~m[1868]&~m[1869]&m[1871]&m[1872])|(m[1822]&~m[1868]&~m[1869]&m[1871]&m[1872])|(~m[1822]&m[1868]&~m[1869]&m[1871]&m[1872])|(m[1822]&m[1868]&~m[1869]&m[1871]&m[1872])|(~m[1822]&~m[1868]&m[1869]&m[1871]&m[1872])|(m[1822]&~m[1868]&m[1869]&m[1871]&m[1872])|(m[1822]&m[1868]&m[1869]&m[1871]&m[1872]));
    m[1875] = (((m[1827]&~m[1873]&~m[1874]&~m[1876]&~m[1877])|(~m[1827]&~m[1873]&~m[1874]&m[1876]&~m[1877])|(m[1827]&m[1873]&~m[1874]&m[1876]&~m[1877])|(m[1827]&~m[1873]&m[1874]&m[1876]&~m[1877])|(~m[1827]&m[1873]&~m[1874]&~m[1876]&m[1877])|(~m[1827]&~m[1873]&m[1874]&~m[1876]&m[1877])|(m[1827]&m[1873]&m[1874]&~m[1876]&m[1877])|(~m[1827]&m[1873]&m[1874]&m[1876]&m[1877]))&UnbiasedRNG[445])|((m[1827]&~m[1873]&~m[1874]&m[1876]&~m[1877])|(~m[1827]&~m[1873]&~m[1874]&~m[1876]&m[1877])|(m[1827]&~m[1873]&~m[1874]&~m[1876]&m[1877])|(m[1827]&m[1873]&~m[1874]&~m[1876]&m[1877])|(m[1827]&~m[1873]&m[1874]&~m[1876]&m[1877])|(~m[1827]&~m[1873]&~m[1874]&m[1876]&m[1877])|(m[1827]&~m[1873]&~m[1874]&m[1876]&m[1877])|(~m[1827]&m[1873]&~m[1874]&m[1876]&m[1877])|(m[1827]&m[1873]&~m[1874]&m[1876]&m[1877])|(~m[1827]&~m[1873]&m[1874]&m[1876]&m[1877])|(m[1827]&~m[1873]&m[1874]&m[1876]&m[1877])|(m[1827]&m[1873]&m[1874]&m[1876]&m[1877]));
    m[1880] = (((m[1832]&~m[1878]&~m[1879]&~m[1881]&~m[1882])|(~m[1832]&~m[1878]&~m[1879]&m[1881]&~m[1882])|(m[1832]&m[1878]&~m[1879]&m[1881]&~m[1882])|(m[1832]&~m[1878]&m[1879]&m[1881]&~m[1882])|(~m[1832]&m[1878]&~m[1879]&~m[1881]&m[1882])|(~m[1832]&~m[1878]&m[1879]&~m[1881]&m[1882])|(m[1832]&m[1878]&m[1879]&~m[1881]&m[1882])|(~m[1832]&m[1878]&m[1879]&m[1881]&m[1882]))&UnbiasedRNG[446])|((m[1832]&~m[1878]&~m[1879]&m[1881]&~m[1882])|(~m[1832]&~m[1878]&~m[1879]&~m[1881]&m[1882])|(m[1832]&~m[1878]&~m[1879]&~m[1881]&m[1882])|(m[1832]&m[1878]&~m[1879]&~m[1881]&m[1882])|(m[1832]&~m[1878]&m[1879]&~m[1881]&m[1882])|(~m[1832]&~m[1878]&~m[1879]&m[1881]&m[1882])|(m[1832]&~m[1878]&~m[1879]&m[1881]&m[1882])|(~m[1832]&m[1878]&~m[1879]&m[1881]&m[1882])|(m[1832]&m[1878]&~m[1879]&m[1881]&m[1882])|(~m[1832]&~m[1878]&m[1879]&m[1881]&m[1882])|(m[1832]&~m[1878]&m[1879]&m[1881]&m[1882])|(m[1832]&m[1878]&m[1879]&m[1881]&m[1882]));
    m[1885] = (((m[1837]&~m[1883]&~m[1884]&~m[1886]&~m[1887])|(~m[1837]&~m[1883]&~m[1884]&m[1886]&~m[1887])|(m[1837]&m[1883]&~m[1884]&m[1886]&~m[1887])|(m[1837]&~m[1883]&m[1884]&m[1886]&~m[1887])|(~m[1837]&m[1883]&~m[1884]&~m[1886]&m[1887])|(~m[1837]&~m[1883]&m[1884]&~m[1886]&m[1887])|(m[1837]&m[1883]&m[1884]&~m[1886]&m[1887])|(~m[1837]&m[1883]&m[1884]&m[1886]&m[1887]))&UnbiasedRNG[447])|((m[1837]&~m[1883]&~m[1884]&m[1886]&~m[1887])|(~m[1837]&~m[1883]&~m[1884]&~m[1886]&m[1887])|(m[1837]&~m[1883]&~m[1884]&~m[1886]&m[1887])|(m[1837]&m[1883]&~m[1884]&~m[1886]&m[1887])|(m[1837]&~m[1883]&m[1884]&~m[1886]&m[1887])|(~m[1837]&~m[1883]&~m[1884]&m[1886]&m[1887])|(m[1837]&~m[1883]&~m[1884]&m[1886]&m[1887])|(~m[1837]&m[1883]&~m[1884]&m[1886]&m[1887])|(m[1837]&m[1883]&~m[1884]&m[1886]&m[1887])|(~m[1837]&~m[1883]&m[1884]&m[1886]&m[1887])|(m[1837]&~m[1883]&m[1884]&m[1886]&m[1887])|(m[1837]&m[1883]&m[1884]&m[1886]&m[1887]));
    m[1890] = (((m[1842]&~m[1888]&~m[1889]&~m[1891]&~m[1892])|(~m[1842]&~m[1888]&~m[1889]&m[1891]&~m[1892])|(m[1842]&m[1888]&~m[1889]&m[1891]&~m[1892])|(m[1842]&~m[1888]&m[1889]&m[1891]&~m[1892])|(~m[1842]&m[1888]&~m[1889]&~m[1891]&m[1892])|(~m[1842]&~m[1888]&m[1889]&~m[1891]&m[1892])|(m[1842]&m[1888]&m[1889]&~m[1891]&m[1892])|(~m[1842]&m[1888]&m[1889]&m[1891]&m[1892]))&UnbiasedRNG[448])|((m[1842]&~m[1888]&~m[1889]&m[1891]&~m[1892])|(~m[1842]&~m[1888]&~m[1889]&~m[1891]&m[1892])|(m[1842]&~m[1888]&~m[1889]&~m[1891]&m[1892])|(m[1842]&m[1888]&~m[1889]&~m[1891]&m[1892])|(m[1842]&~m[1888]&m[1889]&~m[1891]&m[1892])|(~m[1842]&~m[1888]&~m[1889]&m[1891]&m[1892])|(m[1842]&~m[1888]&~m[1889]&m[1891]&m[1892])|(~m[1842]&m[1888]&~m[1889]&m[1891]&m[1892])|(m[1842]&m[1888]&~m[1889]&m[1891]&m[1892])|(~m[1842]&~m[1888]&m[1889]&m[1891]&m[1892])|(m[1842]&~m[1888]&m[1889]&m[1891]&m[1892])|(m[1842]&m[1888]&m[1889]&m[1891]&m[1892]));
    m[1895] = (((m[1847]&~m[1893]&~m[1894]&~m[1896]&~m[1897])|(~m[1847]&~m[1893]&~m[1894]&m[1896]&~m[1897])|(m[1847]&m[1893]&~m[1894]&m[1896]&~m[1897])|(m[1847]&~m[1893]&m[1894]&m[1896]&~m[1897])|(~m[1847]&m[1893]&~m[1894]&~m[1896]&m[1897])|(~m[1847]&~m[1893]&m[1894]&~m[1896]&m[1897])|(m[1847]&m[1893]&m[1894]&~m[1896]&m[1897])|(~m[1847]&m[1893]&m[1894]&m[1896]&m[1897]))&UnbiasedRNG[449])|((m[1847]&~m[1893]&~m[1894]&m[1896]&~m[1897])|(~m[1847]&~m[1893]&~m[1894]&~m[1896]&m[1897])|(m[1847]&~m[1893]&~m[1894]&~m[1896]&m[1897])|(m[1847]&m[1893]&~m[1894]&~m[1896]&m[1897])|(m[1847]&~m[1893]&m[1894]&~m[1896]&m[1897])|(~m[1847]&~m[1893]&~m[1894]&m[1896]&m[1897])|(m[1847]&~m[1893]&~m[1894]&m[1896]&m[1897])|(~m[1847]&m[1893]&~m[1894]&m[1896]&m[1897])|(m[1847]&m[1893]&~m[1894]&m[1896]&m[1897])|(~m[1847]&~m[1893]&m[1894]&m[1896]&m[1897])|(m[1847]&~m[1893]&m[1894]&m[1896]&m[1897])|(m[1847]&m[1893]&m[1894]&m[1896]&m[1897]));
    m[1900] = (((m[1852]&~m[1898]&~m[1899]&~m[1901]&~m[1902])|(~m[1852]&~m[1898]&~m[1899]&m[1901]&~m[1902])|(m[1852]&m[1898]&~m[1899]&m[1901]&~m[1902])|(m[1852]&~m[1898]&m[1899]&m[1901]&~m[1902])|(~m[1852]&m[1898]&~m[1899]&~m[1901]&m[1902])|(~m[1852]&~m[1898]&m[1899]&~m[1901]&m[1902])|(m[1852]&m[1898]&m[1899]&~m[1901]&m[1902])|(~m[1852]&m[1898]&m[1899]&m[1901]&m[1902]))&UnbiasedRNG[450])|((m[1852]&~m[1898]&~m[1899]&m[1901]&~m[1902])|(~m[1852]&~m[1898]&~m[1899]&~m[1901]&m[1902])|(m[1852]&~m[1898]&~m[1899]&~m[1901]&m[1902])|(m[1852]&m[1898]&~m[1899]&~m[1901]&m[1902])|(m[1852]&~m[1898]&m[1899]&~m[1901]&m[1902])|(~m[1852]&~m[1898]&~m[1899]&m[1901]&m[1902])|(m[1852]&~m[1898]&~m[1899]&m[1901]&m[1902])|(~m[1852]&m[1898]&~m[1899]&m[1901]&m[1902])|(m[1852]&m[1898]&~m[1899]&m[1901]&m[1902])|(~m[1852]&~m[1898]&m[1899]&m[1901]&m[1902])|(m[1852]&~m[1898]&m[1899]&m[1901]&m[1902])|(m[1852]&m[1898]&m[1899]&m[1901]&m[1902]));
    m[1905] = (((m[1862]&~m[1903]&~m[1904]&~m[1906]&~m[1907])|(~m[1862]&~m[1903]&~m[1904]&m[1906]&~m[1907])|(m[1862]&m[1903]&~m[1904]&m[1906]&~m[1907])|(m[1862]&~m[1903]&m[1904]&m[1906]&~m[1907])|(~m[1862]&m[1903]&~m[1904]&~m[1906]&m[1907])|(~m[1862]&~m[1903]&m[1904]&~m[1906]&m[1907])|(m[1862]&m[1903]&m[1904]&~m[1906]&m[1907])|(~m[1862]&m[1903]&m[1904]&m[1906]&m[1907]))&UnbiasedRNG[451])|((m[1862]&~m[1903]&~m[1904]&m[1906]&~m[1907])|(~m[1862]&~m[1903]&~m[1904]&~m[1906]&m[1907])|(m[1862]&~m[1903]&~m[1904]&~m[1906]&m[1907])|(m[1862]&m[1903]&~m[1904]&~m[1906]&m[1907])|(m[1862]&~m[1903]&m[1904]&~m[1906]&m[1907])|(~m[1862]&~m[1903]&~m[1904]&m[1906]&m[1907])|(m[1862]&~m[1903]&~m[1904]&m[1906]&m[1907])|(~m[1862]&m[1903]&~m[1904]&m[1906]&m[1907])|(m[1862]&m[1903]&~m[1904]&m[1906]&m[1907])|(~m[1862]&~m[1903]&m[1904]&m[1906]&m[1907])|(m[1862]&~m[1903]&m[1904]&m[1906]&m[1907])|(m[1862]&m[1903]&m[1904]&m[1906]&m[1907]));
    m[1910] = (((m[1867]&~m[1908]&~m[1909]&~m[1911]&~m[1912])|(~m[1867]&~m[1908]&~m[1909]&m[1911]&~m[1912])|(m[1867]&m[1908]&~m[1909]&m[1911]&~m[1912])|(m[1867]&~m[1908]&m[1909]&m[1911]&~m[1912])|(~m[1867]&m[1908]&~m[1909]&~m[1911]&m[1912])|(~m[1867]&~m[1908]&m[1909]&~m[1911]&m[1912])|(m[1867]&m[1908]&m[1909]&~m[1911]&m[1912])|(~m[1867]&m[1908]&m[1909]&m[1911]&m[1912]))&UnbiasedRNG[452])|((m[1867]&~m[1908]&~m[1909]&m[1911]&~m[1912])|(~m[1867]&~m[1908]&~m[1909]&~m[1911]&m[1912])|(m[1867]&~m[1908]&~m[1909]&~m[1911]&m[1912])|(m[1867]&m[1908]&~m[1909]&~m[1911]&m[1912])|(m[1867]&~m[1908]&m[1909]&~m[1911]&m[1912])|(~m[1867]&~m[1908]&~m[1909]&m[1911]&m[1912])|(m[1867]&~m[1908]&~m[1909]&m[1911]&m[1912])|(~m[1867]&m[1908]&~m[1909]&m[1911]&m[1912])|(m[1867]&m[1908]&~m[1909]&m[1911]&m[1912])|(~m[1867]&~m[1908]&m[1909]&m[1911]&m[1912])|(m[1867]&~m[1908]&m[1909]&m[1911]&m[1912])|(m[1867]&m[1908]&m[1909]&m[1911]&m[1912]));
    m[1915] = (((m[1872]&~m[1913]&~m[1914]&~m[1916]&~m[1917])|(~m[1872]&~m[1913]&~m[1914]&m[1916]&~m[1917])|(m[1872]&m[1913]&~m[1914]&m[1916]&~m[1917])|(m[1872]&~m[1913]&m[1914]&m[1916]&~m[1917])|(~m[1872]&m[1913]&~m[1914]&~m[1916]&m[1917])|(~m[1872]&~m[1913]&m[1914]&~m[1916]&m[1917])|(m[1872]&m[1913]&m[1914]&~m[1916]&m[1917])|(~m[1872]&m[1913]&m[1914]&m[1916]&m[1917]))&UnbiasedRNG[453])|((m[1872]&~m[1913]&~m[1914]&m[1916]&~m[1917])|(~m[1872]&~m[1913]&~m[1914]&~m[1916]&m[1917])|(m[1872]&~m[1913]&~m[1914]&~m[1916]&m[1917])|(m[1872]&m[1913]&~m[1914]&~m[1916]&m[1917])|(m[1872]&~m[1913]&m[1914]&~m[1916]&m[1917])|(~m[1872]&~m[1913]&~m[1914]&m[1916]&m[1917])|(m[1872]&~m[1913]&~m[1914]&m[1916]&m[1917])|(~m[1872]&m[1913]&~m[1914]&m[1916]&m[1917])|(m[1872]&m[1913]&~m[1914]&m[1916]&m[1917])|(~m[1872]&~m[1913]&m[1914]&m[1916]&m[1917])|(m[1872]&~m[1913]&m[1914]&m[1916]&m[1917])|(m[1872]&m[1913]&m[1914]&m[1916]&m[1917]));
    m[1920] = (((m[1877]&~m[1918]&~m[1919]&~m[1921]&~m[1922])|(~m[1877]&~m[1918]&~m[1919]&m[1921]&~m[1922])|(m[1877]&m[1918]&~m[1919]&m[1921]&~m[1922])|(m[1877]&~m[1918]&m[1919]&m[1921]&~m[1922])|(~m[1877]&m[1918]&~m[1919]&~m[1921]&m[1922])|(~m[1877]&~m[1918]&m[1919]&~m[1921]&m[1922])|(m[1877]&m[1918]&m[1919]&~m[1921]&m[1922])|(~m[1877]&m[1918]&m[1919]&m[1921]&m[1922]))&UnbiasedRNG[454])|((m[1877]&~m[1918]&~m[1919]&m[1921]&~m[1922])|(~m[1877]&~m[1918]&~m[1919]&~m[1921]&m[1922])|(m[1877]&~m[1918]&~m[1919]&~m[1921]&m[1922])|(m[1877]&m[1918]&~m[1919]&~m[1921]&m[1922])|(m[1877]&~m[1918]&m[1919]&~m[1921]&m[1922])|(~m[1877]&~m[1918]&~m[1919]&m[1921]&m[1922])|(m[1877]&~m[1918]&~m[1919]&m[1921]&m[1922])|(~m[1877]&m[1918]&~m[1919]&m[1921]&m[1922])|(m[1877]&m[1918]&~m[1919]&m[1921]&m[1922])|(~m[1877]&~m[1918]&m[1919]&m[1921]&m[1922])|(m[1877]&~m[1918]&m[1919]&m[1921]&m[1922])|(m[1877]&m[1918]&m[1919]&m[1921]&m[1922]));
    m[1925] = (((m[1882]&~m[1923]&~m[1924]&~m[1926]&~m[1927])|(~m[1882]&~m[1923]&~m[1924]&m[1926]&~m[1927])|(m[1882]&m[1923]&~m[1924]&m[1926]&~m[1927])|(m[1882]&~m[1923]&m[1924]&m[1926]&~m[1927])|(~m[1882]&m[1923]&~m[1924]&~m[1926]&m[1927])|(~m[1882]&~m[1923]&m[1924]&~m[1926]&m[1927])|(m[1882]&m[1923]&m[1924]&~m[1926]&m[1927])|(~m[1882]&m[1923]&m[1924]&m[1926]&m[1927]))&UnbiasedRNG[455])|((m[1882]&~m[1923]&~m[1924]&m[1926]&~m[1927])|(~m[1882]&~m[1923]&~m[1924]&~m[1926]&m[1927])|(m[1882]&~m[1923]&~m[1924]&~m[1926]&m[1927])|(m[1882]&m[1923]&~m[1924]&~m[1926]&m[1927])|(m[1882]&~m[1923]&m[1924]&~m[1926]&m[1927])|(~m[1882]&~m[1923]&~m[1924]&m[1926]&m[1927])|(m[1882]&~m[1923]&~m[1924]&m[1926]&m[1927])|(~m[1882]&m[1923]&~m[1924]&m[1926]&m[1927])|(m[1882]&m[1923]&~m[1924]&m[1926]&m[1927])|(~m[1882]&~m[1923]&m[1924]&m[1926]&m[1927])|(m[1882]&~m[1923]&m[1924]&m[1926]&m[1927])|(m[1882]&m[1923]&m[1924]&m[1926]&m[1927]));
    m[1930] = (((m[1887]&~m[1928]&~m[1929]&~m[1931]&~m[1932])|(~m[1887]&~m[1928]&~m[1929]&m[1931]&~m[1932])|(m[1887]&m[1928]&~m[1929]&m[1931]&~m[1932])|(m[1887]&~m[1928]&m[1929]&m[1931]&~m[1932])|(~m[1887]&m[1928]&~m[1929]&~m[1931]&m[1932])|(~m[1887]&~m[1928]&m[1929]&~m[1931]&m[1932])|(m[1887]&m[1928]&m[1929]&~m[1931]&m[1932])|(~m[1887]&m[1928]&m[1929]&m[1931]&m[1932]))&UnbiasedRNG[456])|((m[1887]&~m[1928]&~m[1929]&m[1931]&~m[1932])|(~m[1887]&~m[1928]&~m[1929]&~m[1931]&m[1932])|(m[1887]&~m[1928]&~m[1929]&~m[1931]&m[1932])|(m[1887]&m[1928]&~m[1929]&~m[1931]&m[1932])|(m[1887]&~m[1928]&m[1929]&~m[1931]&m[1932])|(~m[1887]&~m[1928]&~m[1929]&m[1931]&m[1932])|(m[1887]&~m[1928]&~m[1929]&m[1931]&m[1932])|(~m[1887]&m[1928]&~m[1929]&m[1931]&m[1932])|(m[1887]&m[1928]&~m[1929]&m[1931]&m[1932])|(~m[1887]&~m[1928]&m[1929]&m[1931]&m[1932])|(m[1887]&~m[1928]&m[1929]&m[1931]&m[1932])|(m[1887]&m[1928]&m[1929]&m[1931]&m[1932]));
    m[1935] = (((m[1892]&~m[1933]&~m[1934]&~m[1936]&~m[1937])|(~m[1892]&~m[1933]&~m[1934]&m[1936]&~m[1937])|(m[1892]&m[1933]&~m[1934]&m[1936]&~m[1937])|(m[1892]&~m[1933]&m[1934]&m[1936]&~m[1937])|(~m[1892]&m[1933]&~m[1934]&~m[1936]&m[1937])|(~m[1892]&~m[1933]&m[1934]&~m[1936]&m[1937])|(m[1892]&m[1933]&m[1934]&~m[1936]&m[1937])|(~m[1892]&m[1933]&m[1934]&m[1936]&m[1937]))&UnbiasedRNG[457])|((m[1892]&~m[1933]&~m[1934]&m[1936]&~m[1937])|(~m[1892]&~m[1933]&~m[1934]&~m[1936]&m[1937])|(m[1892]&~m[1933]&~m[1934]&~m[1936]&m[1937])|(m[1892]&m[1933]&~m[1934]&~m[1936]&m[1937])|(m[1892]&~m[1933]&m[1934]&~m[1936]&m[1937])|(~m[1892]&~m[1933]&~m[1934]&m[1936]&m[1937])|(m[1892]&~m[1933]&~m[1934]&m[1936]&m[1937])|(~m[1892]&m[1933]&~m[1934]&m[1936]&m[1937])|(m[1892]&m[1933]&~m[1934]&m[1936]&m[1937])|(~m[1892]&~m[1933]&m[1934]&m[1936]&m[1937])|(m[1892]&~m[1933]&m[1934]&m[1936]&m[1937])|(m[1892]&m[1933]&m[1934]&m[1936]&m[1937]));
    m[1940] = (((m[1897]&~m[1938]&~m[1939]&~m[1941]&~m[1942])|(~m[1897]&~m[1938]&~m[1939]&m[1941]&~m[1942])|(m[1897]&m[1938]&~m[1939]&m[1941]&~m[1942])|(m[1897]&~m[1938]&m[1939]&m[1941]&~m[1942])|(~m[1897]&m[1938]&~m[1939]&~m[1941]&m[1942])|(~m[1897]&~m[1938]&m[1939]&~m[1941]&m[1942])|(m[1897]&m[1938]&m[1939]&~m[1941]&m[1942])|(~m[1897]&m[1938]&m[1939]&m[1941]&m[1942]))&UnbiasedRNG[458])|((m[1897]&~m[1938]&~m[1939]&m[1941]&~m[1942])|(~m[1897]&~m[1938]&~m[1939]&~m[1941]&m[1942])|(m[1897]&~m[1938]&~m[1939]&~m[1941]&m[1942])|(m[1897]&m[1938]&~m[1939]&~m[1941]&m[1942])|(m[1897]&~m[1938]&m[1939]&~m[1941]&m[1942])|(~m[1897]&~m[1938]&~m[1939]&m[1941]&m[1942])|(m[1897]&~m[1938]&~m[1939]&m[1941]&m[1942])|(~m[1897]&m[1938]&~m[1939]&m[1941]&m[1942])|(m[1897]&m[1938]&~m[1939]&m[1941]&m[1942])|(~m[1897]&~m[1938]&m[1939]&m[1941]&m[1942])|(m[1897]&~m[1938]&m[1939]&m[1941]&m[1942])|(m[1897]&m[1938]&m[1939]&m[1941]&m[1942]));
    m[1945] = (((m[1902]&~m[1943]&~m[1944]&~m[1946]&~m[1947])|(~m[1902]&~m[1943]&~m[1944]&m[1946]&~m[1947])|(m[1902]&m[1943]&~m[1944]&m[1946]&~m[1947])|(m[1902]&~m[1943]&m[1944]&m[1946]&~m[1947])|(~m[1902]&m[1943]&~m[1944]&~m[1946]&m[1947])|(~m[1902]&~m[1943]&m[1944]&~m[1946]&m[1947])|(m[1902]&m[1943]&m[1944]&~m[1946]&m[1947])|(~m[1902]&m[1943]&m[1944]&m[1946]&m[1947]))&UnbiasedRNG[459])|((m[1902]&~m[1943]&~m[1944]&m[1946]&~m[1947])|(~m[1902]&~m[1943]&~m[1944]&~m[1946]&m[1947])|(m[1902]&~m[1943]&~m[1944]&~m[1946]&m[1947])|(m[1902]&m[1943]&~m[1944]&~m[1946]&m[1947])|(m[1902]&~m[1943]&m[1944]&~m[1946]&m[1947])|(~m[1902]&~m[1943]&~m[1944]&m[1946]&m[1947])|(m[1902]&~m[1943]&~m[1944]&m[1946]&m[1947])|(~m[1902]&m[1943]&~m[1944]&m[1946]&m[1947])|(m[1902]&m[1943]&~m[1944]&m[1946]&m[1947])|(~m[1902]&~m[1943]&m[1944]&m[1946]&m[1947])|(m[1902]&~m[1943]&m[1944]&m[1946]&m[1947])|(m[1902]&m[1943]&m[1944]&m[1946]&m[1947]));
    m[1950] = (((m[1912]&~m[1948]&~m[1949]&~m[1951]&~m[1952])|(~m[1912]&~m[1948]&~m[1949]&m[1951]&~m[1952])|(m[1912]&m[1948]&~m[1949]&m[1951]&~m[1952])|(m[1912]&~m[1948]&m[1949]&m[1951]&~m[1952])|(~m[1912]&m[1948]&~m[1949]&~m[1951]&m[1952])|(~m[1912]&~m[1948]&m[1949]&~m[1951]&m[1952])|(m[1912]&m[1948]&m[1949]&~m[1951]&m[1952])|(~m[1912]&m[1948]&m[1949]&m[1951]&m[1952]))&UnbiasedRNG[460])|((m[1912]&~m[1948]&~m[1949]&m[1951]&~m[1952])|(~m[1912]&~m[1948]&~m[1949]&~m[1951]&m[1952])|(m[1912]&~m[1948]&~m[1949]&~m[1951]&m[1952])|(m[1912]&m[1948]&~m[1949]&~m[1951]&m[1952])|(m[1912]&~m[1948]&m[1949]&~m[1951]&m[1952])|(~m[1912]&~m[1948]&~m[1949]&m[1951]&m[1952])|(m[1912]&~m[1948]&~m[1949]&m[1951]&m[1952])|(~m[1912]&m[1948]&~m[1949]&m[1951]&m[1952])|(m[1912]&m[1948]&~m[1949]&m[1951]&m[1952])|(~m[1912]&~m[1948]&m[1949]&m[1951]&m[1952])|(m[1912]&~m[1948]&m[1949]&m[1951]&m[1952])|(m[1912]&m[1948]&m[1949]&m[1951]&m[1952]));
    m[1955] = (((m[1917]&~m[1953]&~m[1954]&~m[1956]&~m[1957])|(~m[1917]&~m[1953]&~m[1954]&m[1956]&~m[1957])|(m[1917]&m[1953]&~m[1954]&m[1956]&~m[1957])|(m[1917]&~m[1953]&m[1954]&m[1956]&~m[1957])|(~m[1917]&m[1953]&~m[1954]&~m[1956]&m[1957])|(~m[1917]&~m[1953]&m[1954]&~m[1956]&m[1957])|(m[1917]&m[1953]&m[1954]&~m[1956]&m[1957])|(~m[1917]&m[1953]&m[1954]&m[1956]&m[1957]))&UnbiasedRNG[461])|((m[1917]&~m[1953]&~m[1954]&m[1956]&~m[1957])|(~m[1917]&~m[1953]&~m[1954]&~m[1956]&m[1957])|(m[1917]&~m[1953]&~m[1954]&~m[1956]&m[1957])|(m[1917]&m[1953]&~m[1954]&~m[1956]&m[1957])|(m[1917]&~m[1953]&m[1954]&~m[1956]&m[1957])|(~m[1917]&~m[1953]&~m[1954]&m[1956]&m[1957])|(m[1917]&~m[1953]&~m[1954]&m[1956]&m[1957])|(~m[1917]&m[1953]&~m[1954]&m[1956]&m[1957])|(m[1917]&m[1953]&~m[1954]&m[1956]&m[1957])|(~m[1917]&~m[1953]&m[1954]&m[1956]&m[1957])|(m[1917]&~m[1953]&m[1954]&m[1956]&m[1957])|(m[1917]&m[1953]&m[1954]&m[1956]&m[1957]));
    m[1960] = (((m[1922]&~m[1958]&~m[1959]&~m[1961]&~m[1962])|(~m[1922]&~m[1958]&~m[1959]&m[1961]&~m[1962])|(m[1922]&m[1958]&~m[1959]&m[1961]&~m[1962])|(m[1922]&~m[1958]&m[1959]&m[1961]&~m[1962])|(~m[1922]&m[1958]&~m[1959]&~m[1961]&m[1962])|(~m[1922]&~m[1958]&m[1959]&~m[1961]&m[1962])|(m[1922]&m[1958]&m[1959]&~m[1961]&m[1962])|(~m[1922]&m[1958]&m[1959]&m[1961]&m[1962]))&UnbiasedRNG[462])|((m[1922]&~m[1958]&~m[1959]&m[1961]&~m[1962])|(~m[1922]&~m[1958]&~m[1959]&~m[1961]&m[1962])|(m[1922]&~m[1958]&~m[1959]&~m[1961]&m[1962])|(m[1922]&m[1958]&~m[1959]&~m[1961]&m[1962])|(m[1922]&~m[1958]&m[1959]&~m[1961]&m[1962])|(~m[1922]&~m[1958]&~m[1959]&m[1961]&m[1962])|(m[1922]&~m[1958]&~m[1959]&m[1961]&m[1962])|(~m[1922]&m[1958]&~m[1959]&m[1961]&m[1962])|(m[1922]&m[1958]&~m[1959]&m[1961]&m[1962])|(~m[1922]&~m[1958]&m[1959]&m[1961]&m[1962])|(m[1922]&~m[1958]&m[1959]&m[1961]&m[1962])|(m[1922]&m[1958]&m[1959]&m[1961]&m[1962]));
    m[1965] = (((m[1927]&~m[1963]&~m[1964]&~m[1966]&~m[1967])|(~m[1927]&~m[1963]&~m[1964]&m[1966]&~m[1967])|(m[1927]&m[1963]&~m[1964]&m[1966]&~m[1967])|(m[1927]&~m[1963]&m[1964]&m[1966]&~m[1967])|(~m[1927]&m[1963]&~m[1964]&~m[1966]&m[1967])|(~m[1927]&~m[1963]&m[1964]&~m[1966]&m[1967])|(m[1927]&m[1963]&m[1964]&~m[1966]&m[1967])|(~m[1927]&m[1963]&m[1964]&m[1966]&m[1967]))&UnbiasedRNG[463])|((m[1927]&~m[1963]&~m[1964]&m[1966]&~m[1967])|(~m[1927]&~m[1963]&~m[1964]&~m[1966]&m[1967])|(m[1927]&~m[1963]&~m[1964]&~m[1966]&m[1967])|(m[1927]&m[1963]&~m[1964]&~m[1966]&m[1967])|(m[1927]&~m[1963]&m[1964]&~m[1966]&m[1967])|(~m[1927]&~m[1963]&~m[1964]&m[1966]&m[1967])|(m[1927]&~m[1963]&~m[1964]&m[1966]&m[1967])|(~m[1927]&m[1963]&~m[1964]&m[1966]&m[1967])|(m[1927]&m[1963]&~m[1964]&m[1966]&m[1967])|(~m[1927]&~m[1963]&m[1964]&m[1966]&m[1967])|(m[1927]&~m[1963]&m[1964]&m[1966]&m[1967])|(m[1927]&m[1963]&m[1964]&m[1966]&m[1967]));
    m[1970] = (((m[1932]&~m[1968]&~m[1969]&~m[1971]&~m[1972])|(~m[1932]&~m[1968]&~m[1969]&m[1971]&~m[1972])|(m[1932]&m[1968]&~m[1969]&m[1971]&~m[1972])|(m[1932]&~m[1968]&m[1969]&m[1971]&~m[1972])|(~m[1932]&m[1968]&~m[1969]&~m[1971]&m[1972])|(~m[1932]&~m[1968]&m[1969]&~m[1971]&m[1972])|(m[1932]&m[1968]&m[1969]&~m[1971]&m[1972])|(~m[1932]&m[1968]&m[1969]&m[1971]&m[1972]))&UnbiasedRNG[464])|((m[1932]&~m[1968]&~m[1969]&m[1971]&~m[1972])|(~m[1932]&~m[1968]&~m[1969]&~m[1971]&m[1972])|(m[1932]&~m[1968]&~m[1969]&~m[1971]&m[1972])|(m[1932]&m[1968]&~m[1969]&~m[1971]&m[1972])|(m[1932]&~m[1968]&m[1969]&~m[1971]&m[1972])|(~m[1932]&~m[1968]&~m[1969]&m[1971]&m[1972])|(m[1932]&~m[1968]&~m[1969]&m[1971]&m[1972])|(~m[1932]&m[1968]&~m[1969]&m[1971]&m[1972])|(m[1932]&m[1968]&~m[1969]&m[1971]&m[1972])|(~m[1932]&~m[1968]&m[1969]&m[1971]&m[1972])|(m[1932]&~m[1968]&m[1969]&m[1971]&m[1972])|(m[1932]&m[1968]&m[1969]&m[1971]&m[1972]));
    m[1975] = (((m[1937]&~m[1973]&~m[1974]&~m[1976]&~m[1977])|(~m[1937]&~m[1973]&~m[1974]&m[1976]&~m[1977])|(m[1937]&m[1973]&~m[1974]&m[1976]&~m[1977])|(m[1937]&~m[1973]&m[1974]&m[1976]&~m[1977])|(~m[1937]&m[1973]&~m[1974]&~m[1976]&m[1977])|(~m[1937]&~m[1973]&m[1974]&~m[1976]&m[1977])|(m[1937]&m[1973]&m[1974]&~m[1976]&m[1977])|(~m[1937]&m[1973]&m[1974]&m[1976]&m[1977]))&UnbiasedRNG[465])|((m[1937]&~m[1973]&~m[1974]&m[1976]&~m[1977])|(~m[1937]&~m[1973]&~m[1974]&~m[1976]&m[1977])|(m[1937]&~m[1973]&~m[1974]&~m[1976]&m[1977])|(m[1937]&m[1973]&~m[1974]&~m[1976]&m[1977])|(m[1937]&~m[1973]&m[1974]&~m[1976]&m[1977])|(~m[1937]&~m[1973]&~m[1974]&m[1976]&m[1977])|(m[1937]&~m[1973]&~m[1974]&m[1976]&m[1977])|(~m[1937]&m[1973]&~m[1974]&m[1976]&m[1977])|(m[1937]&m[1973]&~m[1974]&m[1976]&m[1977])|(~m[1937]&~m[1973]&m[1974]&m[1976]&m[1977])|(m[1937]&~m[1973]&m[1974]&m[1976]&m[1977])|(m[1937]&m[1973]&m[1974]&m[1976]&m[1977]));
    m[1980] = (((m[1942]&~m[1978]&~m[1979]&~m[1981]&~m[1982])|(~m[1942]&~m[1978]&~m[1979]&m[1981]&~m[1982])|(m[1942]&m[1978]&~m[1979]&m[1981]&~m[1982])|(m[1942]&~m[1978]&m[1979]&m[1981]&~m[1982])|(~m[1942]&m[1978]&~m[1979]&~m[1981]&m[1982])|(~m[1942]&~m[1978]&m[1979]&~m[1981]&m[1982])|(m[1942]&m[1978]&m[1979]&~m[1981]&m[1982])|(~m[1942]&m[1978]&m[1979]&m[1981]&m[1982]))&UnbiasedRNG[466])|((m[1942]&~m[1978]&~m[1979]&m[1981]&~m[1982])|(~m[1942]&~m[1978]&~m[1979]&~m[1981]&m[1982])|(m[1942]&~m[1978]&~m[1979]&~m[1981]&m[1982])|(m[1942]&m[1978]&~m[1979]&~m[1981]&m[1982])|(m[1942]&~m[1978]&m[1979]&~m[1981]&m[1982])|(~m[1942]&~m[1978]&~m[1979]&m[1981]&m[1982])|(m[1942]&~m[1978]&~m[1979]&m[1981]&m[1982])|(~m[1942]&m[1978]&~m[1979]&m[1981]&m[1982])|(m[1942]&m[1978]&~m[1979]&m[1981]&m[1982])|(~m[1942]&~m[1978]&m[1979]&m[1981]&m[1982])|(m[1942]&~m[1978]&m[1979]&m[1981]&m[1982])|(m[1942]&m[1978]&m[1979]&m[1981]&m[1982]));
    m[1985] = (((m[1947]&~m[1983]&~m[1984]&~m[1986]&~m[1987])|(~m[1947]&~m[1983]&~m[1984]&m[1986]&~m[1987])|(m[1947]&m[1983]&~m[1984]&m[1986]&~m[1987])|(m[1947]&~m[1983]&m[1984]&m[1986]&~m[1987])|(~m[1947]&m[1983]&~m[1984]&~m[1986]&m[1987])|(~m[1947]&~m[1983]&m[1984]&~m[1986]&m[1987])|(m[1947]&m[1983]&m[1984]&~m[1986]&m[1987])|(~m[1947]&m[1983]&m[1984]&m[1986]&m[1987]))&UnbiasedRNG[467])|((m[1947]&~m[1983]&~m[1984]&m[1986]&~m[1987])|(~m[1947]&~m[1983]&~m[1984]&~m[1986]&m[1987])|(m[1947]&~m[1983]&~m[1984]&~m[1986]&m[1987])|(m[1947]&m[1983]&~m[1984]&~m[1986]&m[1987])|(m[1947]&~m[1983]&m[1984]&~m[1986]&m[1987])|(~m[1947]&~m[1983]&~m[1984]&m[1986]&m[1987])|(m[1947]&~m[1983]&~m[1984]&m[1986]&m[1987])|(~m[1947]&m[1983]&~m[1984]&m[1986]&m[1987])|(m[1947]&m[1983]&~m[1984]&m[1986]&m[1987])|(~m[1947]&~m[1983]&m[1984]&m[1986]&m[1987])|(m[1947]&~m[1983]&m[1984]&m[1986]&m[1987])|(m[1947]&m[1983]&m[1984]&m[1986]&m[1987]));
    m[1990] = (((m[1957]&~m[1988]&~m[1989]&~m[1991]&~m[1992])|(~m[1957]&~m[1988]&~m[1989]&m[1991]&~m[1992])|(m[1957]&m[1988]&~m[1989]&m[1991]&~m[1992])|(m[1957]&~m[1988]&m[1989]&m[1991]&~m[1992])|(~m[1957]&m[1988]&~m[1989]&~m[1991]&m[1992])|(~m[1957]&~m[1988]&m[1989]&~m[1991]&m[1992])|(m[1957]&m[1988]&m[1989]&~m[1991]&m[1992])|(~m[1957]&m[1988]&m[1989]&m[1991]&m[1992]))&UnbiasedRNG[468])|((m[1957]&~m[1988]&~m[1989]&m[1991]&~m[1992])|(~m[1957]&~m[1988]&~m[1989]&~m[1991]&m[1992])|(m[1957]&~m[1988]&~m[1989]&~m[1991]&m[1992])|(m[1957]&m[1988]&~m[1989]&~m[1991]&m[1992])|(m[1957]&~m[1988]&m[1989]&~m[1991]&m[1992])|(~m[1957]&~m[1988]&~m[1989]&m[1991]&m[1992])|(m[1957]&~m[1988]&~m[1989]&m[1991]&m[1992])|(~m[1957]&m[1988]&~m[1989]&m[1991]&m[1992])|(m[1957]&m[1988]&~m[1989]&m[1991]&m[1992])|(~m[1957]&~m[1988]&m[1989]&m[1991]&m[1992])|(m[1957]&~m[1988]&m[1989]&m[1991]&m[1992])|(m[1957]&m[1988]&m[1989]&m[1991]&m[1992]));
    m[1995] = (((m[1962]&~m[1993]&~m[1994]&~m[1996]&~m[1997])|(~m[1962]&~m[1993]&~m[1994]&m[1996]&~m[1997])|(m[1962]&m[1993]&~m[1994]&m[1996]&~m[1997])|(m[1962]&~m[1993]&m[1994]&m[1996]&~m[1997])|(~m[1962]&m[1993]&~m[1994]&~m[1996]&m[1997])|(~m[1962]&~m[1993]&m[1994]&~m[1996]&m[1997])|(m[1962]&m[1993]&m[1994]&~m[1996]&m[1997])|(~m[1962]&m[1993]&m[1994]&m[1996]&m[1997]))&UnbiasedRNG[469])|((m[1962]&~m[1993]&~m[1994]&m[1996]&~m[1997])|(~m[1962]&~m[1993]&~m[1994]&~m[1996]&m[1997])|(m[1962]&~m[1993]&~m[1994]&~m[1996]&m[1997])|(m[1962]&m[1993]&~m[1994]&~m[1996]&m[1997])|(m[1962]&~m[1993]&m[1994]&~m[1996]&m[1997])|(~m[1962]&~m[1993]&~m[1994]&m[1996]&m[1997])|(m[1962]&~m[1993]&~m[1994]&m[1996]&m[1997])|(~m[1962]&m[1993]&~m[1994]&m[1996]&m[1997])|(m[1962]&m[1993]&~m[1994]&m[1996]&m[1997])|(~m[1962]&~m[1993]&m[1994]&m[1996]&m[1997])|(m[1962]&~m[1993]&m[1994]&m[1996]&m[1997])|(m[1962]&m[1993]&m[1994]&m[1996]&m[1997]));
    m[2000] = (((m[1967]&~m[1998]&~m[1999]&~m[2001]&~m[2002])|(~m[1967]&~m[1998]&~m[1999]&m[2001]&~m[2002])|(m[1967]&m[1998]&~m[1999]&m[2001]&~m[2002])|(m[1967]&~m[1998]&m[1999]&m[2001]&~m[2002])|(~m[1967]&m[1998]&~m[1999]&~m[2001]&m[2002])|(~m[1967]&~m[1998]&m[1999]&~m[2001]&m[2002])|(m[1967]&m[1998]&m[1999]&~m[2001]&m[2002])|(~m[1967]&m[1998]&m[1999]&m[2001]&m[2002]))&UnbiasedRNG[470])|((m[1967]&~m[1998]&~m[1999]&m[2001]&~m[2002])|(~m[1967]&~m[1998]&~m[1999]&~m[2001]&m[2002])|(m[1967]&~m[1998]&~m[1999]&~m[2001]&m[2002])|(m[1967]&m[1998]&~m[1999]&~m[2001]&m[2002])|(m[1967]&~m[1998]&m[1999]&~m[2001]&m[2002])|(~m[1967]&~m[1998]&~m[1999]&m[2001]&m[2002])|(m[1967]&~m[1998]&~m[1999]&m[2001]&m[2002])|(~m[1967]&m[1998]&~m[1999]&m[2001]&m[2002])|(m[1967]&m[1998]&~m[1999]&m[2001]&m[2002])|(~m[1967]&~m[1998]&m[1999]&m[2001]&m[2002])|(m[1967]&~m[1998]&m[1999]&m[2001]&m[2002])|(m[1967]&m[1998]&m[1999]&m[2001]&m[2002]));
    m[2005] = (((m[1972]&~m[2003]&~m[2004]&~m[2006]&~m[2007])|(~m[1972]&~m[2003]&~m[2004]&m[2006]&~m[2007])|(m[1972]&m[2003]&~m[2004]&m[2006]&~m[2007])|(m[1972]&~m[2003]&m[2004]&m[2006]&~m[2007])|(~m[1972]&m[2003]&~m[2004]&~m[2006]&m[2007])|(~m[1972]&~m[2003]&m[2004]&~m[2006]&m[2007])|(m[1972]&m[2003]&m[2004]&~m[2006]&m[2007])|(~m[1972]&m[2003]&m[2004]&m[2006]&m[2007]))&UnbiasedRNG[471])|((m[1972]&~m[2003]&~m[2004]&m[2006]&~m[2007])|(~m[1972]&~m[2003]&~m[2004]&~m[2006]&m[2007])|(m[1972]&~m[2003]&~m[2004]&~m[2006]&m[2007])|(m[1972]&m[2003]&~m[2004]&~m[2006]&m[2007])|(m[1972]&~m[2003]&m[2004]&~m[2006]&m[2007])|(~m[1972]&~m[2003]&~m[2004]&m[2006]&m[2007])|(m[1972]&~m[2003]&~m[2004]&m[2006]&m[2007])|(~m[1972]&m[2003]&~m[2004]&m[2006]&m[2007])|(m[1972]&m[2003]&~m[2004]&m[2006]&m[2007])|(~m[1972]&~m[2003]&m[2004]&m[2006]&m[2007])|(m[1972]&~m[2003]&m[2004]&m[2006]&m[2007])|(m[1972]&m[2003]&m[2004]&m[2006]&m[2007]));
    m[2010] = (((m[1977]&~m[2008]&~m[2009]&~m[2011]&~m[2012])|(~m[1977]&~m[2008]&~m[2009]&m[2011]&~m[2012])|(m[1977]&m[2008]&~m[2009]&m[2011]&~m[2012])|(m[1977]&~m[2008]&m[2009]&m[2011]&~m[2012])|(~m[1977]&m[2008]&~m[2009]&~m[2011]&m[2012])|(~m[1977]&~m[2008]&m[2009]&~m[2011]&m[2012])|(m[1977]&m[2008]&m[2009]&~m[2011]&m[2012])|(~m[1977]&m[2008]&m[2009]&m[2011]&m[2012]))&UnbiasedRNG[472])|((m[1977]&~m[2008]&~m[2009]&m[2011]&~m[2012])|(~m[1977]&~m[2008]&~m[2009]&~m[2011]&m[2012])|(m[1977]&~m[2008]&~m[2009]&~m[2011]&m[2012])|(m[1977]&m[2008]&~m[2009]&~m[2011]&m[2012])|(m[1977]&~m[2008]&m[2009]&~m[2011]&m[2012])|(~m[1977]&~m[2008]&~m[2009]&m[2011]&m[2012])|(m[1977]&~m[2008]&~m[2009]&m[2011]&m[2012])|(~m[1977]&m[2008]&~m[2009]&m[2011]&m[2012])|(m[1977]&m[2008]&~m[2009]&m[2011]&m[2012])|(~m[1977]&~m[2008]&m[2009]&m[2011]&m[2012])|(m[1977]&~m[2008]&m[2009]&m[2011]&m[2012])|(m[1977]&m[2008]&m[2009]&m[2011]&m[2012]));
    m[2015] = (((m[1982]&~m[2013]&~m[2014]&~m[2016]&~m[2017])|(~m[1982]&~m[2013]&~m[2014]&m[2016]&~m[2017])|(m[1982]&m[2013]&~m[2014]&m[2016]&~m[2017])|(m[1982]&~m[2013]&m[2014]&m[2016]&~m[2017])|(~m[1982]&m[2013]&~m[2014]&~m[2016]&m[2017])|(~m[1982]&~m[2013]&m[2014]&~m[2016]&m[2017])|(m[1982]&m[2013]&m[2014]&~m[2016]&m[2017])|(~m[1982]&m[2013]&m[2014]&m[2016]&m[2017]))&UnbiasedRNG[473])|((m[1982]&~m[2013]&~m[2014]&m[2016]&~m[2017])|(~m[1982]&~m[2013]&~m[2014]&~m[2016]&m[2017])|(m[1982]&~m[2013]&~m[2014]&~m[2016]&m[2017])|(m[1982]&m[2013]&~m[2014]&~m[2016]&m[2017])|(m[1982]&~m[2013]&m[2014]&~m[2016]&m[2017])|(~m[1982]&~m[2013]&~m[2014]&m[2016]&m[2017])|(m[1982]&~m[2013]&~m[2014]&m[2016]&m[2017])|(~m[1982]&m[2013]&~m[2014]&m[2016]&m[2017])|(m[1982]&m[2013]&~m[2014]&m[2016]&m[2017])|(~m[1982]&~m[2013]&m[2014]&m[2016]&m[2017])|(m[1982]&~m[2013]&m[2014]&m[2016]&m[2017])|(m[1982]&m[2013]&m[2014]&m[2016]&m[2017]));
    m[2020] = (((m[1987]&~m[2018]&~m[2019]&~m[2021]&~m[2022])|(~m[1987]&~m[2018]&~m[2019]&m[2021]&~m[2022])|(m[1987]&m[2018]&~m[2019]&m[2021]&~m[2022])|(m[1987]&~m[2018]&m[2019]&m[2021]&~m[2022])|(~m[1987]&m[2018]&~m[2019]&~m[2021]&m[2022])|(~m[1987]&~m[2018]&m[2019]&~m[2021]&m[2022])|(m[1987]&m[2018]&m[2019]&~m[2021]&m[2022])|(~m[1987]&m[2018]&m[2019]&m[2021]&m[2022]))&UnbiasedRNG[474])|((m[1987]&~m[2018]&~m[2019]&m[2021]&~m[2022])|(~m[1987]&~m[2018]&~m[2019]&~m[2021]&m[2022])|(m[1987]&~m[2018]&~m[2019]&~m[2021]&m[2022])|(m[1987]&m[2018]&~m[2019]&~m[2021]&m[2022])|(m[1987]&~m[2018]&m[2019]&~m[2021]&m[2022])|(~m[1987]&~m[2018]&~m[2019]&m[2021]&m[2022])|(m[1987]&~m[2018]&~m[2019]&m[2021]&m[2022])|(~m[1987]&m[2018]&~m[2019]&m[2021]&m[2022])|(m[1987]&m[2018]&~m[2019]&m[2021]&m[2022])|(~m[1987]&~m[2018]&m[2019]&m[2021]&m[2022])|(m[1987]&~m[2018]&m[2019]&m[2021]&m[2022])|(m[1987]&m[2018]&m[2019]&m[2021]&m[2022]));
    m[2025] = (((m[1997]&~m[2023]&~m[2024]&~m[2026]&~m[2027])|(~m[1997]&~m[2023]&~m[2024]&m[2026]&~m[2027])|(m[1997]&m[2023]&~m[2024]&m[2026]&~m[2027])|(m[1997]&~m[2023]&m[2024]&m[2026]&~m[2027])|(~m[1997]&m[2023]&~m[2024]&~m[2026]&m[2027])|(~m[1997]&~m[2023]&m[2024]&~m[2026]&m[2027])|(m[1997]&m[2023]&m[2024]&~m[2026]&m[2027])|(~m[1997]&m[2023]&m[2024]&m[2026]&m[2027]))&UnbiasedRNG[475])|((m[1997]&~m[2023]&~m[2024]&m[2026]&~m[2027])|(~m[1997]&~m[2023]&~m[2024]&~m[2026]&m[2027])|(m[1997]&~m[2023]&~m[2024]&~m[2026]&m[2027])|(m[1997]&m[2023]&~m[2024]&~m[2026]&m[2027])|(m[1997]&~m[2023]&m[2024]&~m[2026]&m[2027])|(~m[1997]&~m[2023]&~m[2024]&m[2026]&m[2027])|(m[1997]&~m[2023]&~m[2024]&m[2026]&m[2027])|(~m[1997]&m[2023]&~m[2024]&m[2026]&m[2027])|(m[1997]&m[2023]&~m[2024]&m[2026]&m[2027])|(~m[1997]&~m[2023]&m[2024]&m[2026]&m[2027])|(m[1997]&~m[2023]&m[2024]&m[2026]&m[2027])|(m[1997]&m[2023]&m[2024]&m[2026]&m[2027]));
    m[2030] = (((m[2002]&~m[2028]&~m[2029]&~m[2031]&~m[2032])|(~m[2002]&~m[2028]&~m[2029]&m[2031]&~m[2032])|(m[2002]&m[2028]&~m[2029]&m[2031]&~m[2032])|(m[2002]&~m[2028]&m[2029]&m[2031]&~m[2032])|(~m[2002]&m[2028]&~m[2029]&~m[2031]&m[2032])|(~m[2002]&~m[2028]&m[2029]&~m[2031]&m[2032])|(m[2002]&m[2028]&m[2029]&~m[2031]&m[2032])|(~m[2002]&m[2028]&m[2029]&m[2031]&m[2032]))&UnbiasedRNG[476])|((m[2002]&~m[2028]&~m[2029]&m[2031]&~m[2032])|(~m[2002]&~m[2028]&~m[2029]&~m[2031]&m[2032])|(m[2002]&~m[2028]&~m[2029]&~m[2031]&m[2032])|(m[2002]&m[2028]&~m[2029]&~m[2031]&m[2032])|(m[2002]&~m[2028]&m[2029]&~m[2031]&m[2032])|(~m[2002]&~m[2028]&~m[2029]&m[2031]&m[2032])|(m[2002]&~m[2028]&~m[2029]&m[2031]&m[2032])|(~m[2002]&m[2028]&~m[2029]&m[2031]&m[2032])|(m[2002]&m[2028]&~m[2029]&m[2031]&m[2032])|(~m[2002]&~m[2028]&m[2029]&m[2031]&m[2032])|(m[2002]&~m[2028]&m[2029]&m[2031]&m[2032])|(m[2002]&m[2028]&m[2029]&m[2031]&m[2032]));
    m[2035] = (((m[2007]&~m[2033]&~m[2034]&~m[2036]&~m[2037])|(~m[2007]&~m[2033]&~m[2034]&m[2036]&~m[2037])|(m[2007]&m[2033]&~m[2034]&m[2036]&~m[2037])|(m[2007]&~m[2033]&m[2034]&m[2036]&~m[2037])|(~m[2007]&m[2033]&~m[2034]&~m[2036]&m[2037])|(~m[2007]&~m[2033]&m[2034]&~m[2036]&m[2037])|(m[2007]&m[2033]&m[2034]&~m[2036]&m[2037])|(~m[2007]&m[2033]&m[2034]&m[2036]&m[2037]))&UnbiasedRNG[477])|((m[2007]&~m[2033]&~m[2034]&m[2036]&~m[2037])|(~m[2007]&~m[2033]&~m[2034]&~m[2036]&m[2037])|(m[2007]&~m[2033]&~m[2034]&~m[2036]&m[2037])|(m[2007]&m[2033]&~m[2034]&~m[2036]&m[2037])|(m[2007]&~m[2033]&m[2034]&~m[2036]&m[2037])|(~m[2007]&~m[2033]&~m[2034]&m[2036]&m[2037])|(m[2007]&~m[2033]&~m[2034]&m[2036]&m[2037])|(~m[2007]&m[2033]&~m[2034]&m[2036]&m[2037])|(m[2007]&m[2033]&~m[2034]&m[2036]&m[2037])|(~m[2007]&~m[2033]&m[2034]&m[2036]&m[2037])|(m[2007]&~m[2033]&m[2034]&m[2036]&m[2037])|(m[2007]&m[2033]&m[2034]&m[2036]&m[2037]));
    m[2040] = (((m[2012]&~m[2038]&~m[2039]&~m[2041]&~m[2042])|(~m[2012]&~m[2038]&~m[2039]&m[2041]&~m[2042])|(m[2012]&m[2038]&~m[2039]&m[2041]&~m[2042])|(m[2012]&~m[2038]&m[2039]&m[2041]&~m[2042])|(~m[2012]&m[2038]&~m[2039]&~m[2041]&m[2042])|(~m[2012]&~m[2038]&m[2039]&~m[2041]&m[2042])|(m[2012]&m[2038]&m[2039]&~m[2041]&m[2042])|(~m[2012]&m[2038]&m[2039]&m[2041]&m[2042]))&UnbiasedRNG[478])|((m[2012]&~m[2038]&~m[2039]&m[2041]&~m[2042])|(~m[2012]&~m[2038]&~m[2039]&~m[2041]&m[2042])|(m[2012]&~m[2038]&~m[2039]&~m[2041]&m[2042])|(m[2012]&m[2038]&~m[2039]&~m[2041]&m[2042])|(m[2012]&~m[2038]&m[2039]&~m[2041]&m[2042])|(~m[2012]&~m[2038]&~m[2039]&m[2041]&m[2042])|(m[2012]&~m[2038]&~m[2039]&m[2041]&m[2042])|(~m[2012]&m[2038]&~m[2039]&m[2041]&m[2042])|(m[2012]&m[2038]&~m[2039]&m[2041]&m[2042])|(~m[2012]&~m[2038]&m[2039]&m[2041]&m[2042])|(m[2012]&~m[2038]&m[2039]&m[2041]&m[2042])|(m[2012]&m[2038]&m[2039]&m[2041]&m[2042]));
    m[2045] = (((m[2017]&~m[2043]&~m[2044]&~m[2046]&~m[2047])|(~m[2017]&~m[2043]&~m[2044]&m[2046]&~m[2047])|(m[2017]&m[2043]&~m[2044]&m[2046]&~m[2047])|(m[2017]&~m[2043]&m[2044]&m[2046]&~m[2047])|(~m[2017]&m[2043]&~m[2044]&~m[2046]&m[2047])|(~m[2017]&~m[2043]&m[2044]&~m[2046]&m[2047])|(m[2017]&m[2043]&m[2044]&~m[2046]&m[2047])|(~m[2017]&m[2043]&m[2044]&m[2046]&m[2047]))&UnbiasedRNG[479])|((m[2017]&~m[2043]&~m[2044]&m[2046]&~m[2047])|(~m[2017]&~m[2043]&~m[2044]&~m[2046]&m[2047])|(m[2017]&~m[2043]&~m[2044]&~m[2046]&m[2047])|(m[2017]&m[2043]&~m[2044]&~m[2046]&m[2047])|(m[2017]&~m[2043]&m[2044]&~m[2046]&m[2047])|(~m[2017]&~m[2043]&~m[2044]&m[2046]&m[2047])|(m[2017]&~m[2043]&~m[2044]&m[2046]&m[2047])|(~m[2017]&m[2043]&~m[2044]&m[2046]&m[2047])|(m[2017]&m[2043]&~m[2044]&m[2046]&m[2047])|(~m[2017]&~m[2043]&m[2044]&m[2046]&m[2047])|(m[2017]&~m[2043]&m[2044]&m[2046]&m[2047])|(m[2017]&m[2043]&m[2044]&m[2046]&m[2047]));
    m[2050] = (((m[2022]&~m[2048]&~m[2049]&~m[2051]&~m[2052])|(~m[2022]&~m[2048]&~m[2049]&m[2051]&~m[2052])|(m[2022]&m[2048]&~m[2049]&m[2051]&~m[2052])|(m[2022]&~m[2048]&m[2049]&m[2051]&~m[2052])|(~m[2022]&m[2048]&~m[2049]&~m[2051]&m[2052])|(~m[2022]&~m[2048]&m[2049]&~m[2051]&m[2052])|(m[2022]&m[2048]&m[2049]&~m[2051]&m[2052])|(~m[2022]&m[2048]&m[2049]&m[2051]&m[2052]))&UnbiasedRNG[480])|((m[2022]&~m[2048]&~m[2049]&m[2051]&~m[2052])|(~m[2022]&~m[2048]&~m[2049]&~m[2051]&m[2052])|(m[2022]&~m[2048]&~m[2049]&~m[2051]&m[2052])|(m[2022]&m[2048]&~m[2049]&~m[2051]&m[2052])|(m[2022]&~m[2048]&m[2049]&~m[2051]&m[2052])|(~m[2022]&~m[2048]&~m[2049]&m[2051]&m[2052])|(m[2022]&~m[2048]&~m[2049]&m[2051]&m[2052])|(~m[2022]&m[2048]&~m[2049]&m[2051]&m[2052])|(m[2022]&m[2048]&~m[2049]&m[2051]&m[2052])|(~m[2022]&~m[2048]&m[2049]&m[2051]&m[2052])|(m[2022]&~m[2048]&m[2049]&m[2051]&m[2052])|(m[2022]&m[2048]&m[2049]&m[2051]&m[2052]));
    m[2055] = (((m[2032]&~m[2053]&~m[2054]&~m[2056]&~m[2057])|(~m[2032]&~m[2053]&~m[2054]&m[2056]&~m[2057])|(m[2032]&m[2053]&~m[2054]&m[2056]&~m[2057])|(m[2032]&~m[2053]&m[2054]&m[2056]&~m[2057])|(~m[2032]&m[2053]&~m[2054]&~m[2056]&m[2057])|(~m[2032]&~m[2053]&m[2054]&~m[2056]&m[2057])|(m[2032]&m[2053]&m[2054]&~m[2056]&m[2057])|(~m[2032]&m[2053]&m[2054]&m[2056]&m[2057]))&UnbiasedRNG[481])|((m[2032]&~m[2053]&~m[2054]&m[2056]&~m[2057])|(~m[2032]&~m[2053]&~m[2054]&~m[2056]&m[2057])|(m[2032]&~m[2053]&~m[2054]&~m[2056]&m[2057])|(m[2032]&m[2053]&~m[2054]&~m[2056]&m[2057])|(m[2032]&~m[2053]&m[2054]&~m[2056]&m[2057])|(~m[2032]&~m[2053]&~m[2054]&m[2056]&m[2057])|(m[2032]&~m[2053]&~m[2054]&m[2056]&m[2057])|(~m[2032]&m[2053]&~m[2054]&m[2056]&m[2057])|(m[2032]&m[2053]&~m[2054]&m[2056]&m[2057])|(~m[2032]&~m[2053]&m[2054]&m[2056]&m[2057])|(m[2032]&~m[2053]&m[2054]&m[2056]&m[2057])|(m[2032]&m[2053]&m[2054]&m[2056]&m[2057]));
    m[2060] = (((m[2037]&~m[2058]&~m[2059]&~m[2061]&~m[2062])|(~m[2037]&~m[2058]&~m[2059]&m[2061]&~m[2062])|(m[2037]&m[2058]&~m[2059]&m[2061]&~m[2062])|(m[2037]&~m[2058]&m[2059]&m[2061]&~m[2062])|(~m[2037]&m[2058]&~m[2059]&~m[2061]&m[2062])|(~m[2037]&~m[2058]&m[2059]&~m[2061]&m[2062])|(m[2037]&m[2058]&m[2059]&~m[2061]&m[2062])|(~m[2037]&m[2058]&m[2059]&m[2061]&m[2062]))&UnbiasedRNG[482])|((m[2037]&~m[2058]&~m[2059]&m[2061]&~m[2062])|(~m[2037]&~m[2058]&~m[2059]&~m[2061]&m[2062])|(m[2037]&~m[2058]&~m[2059]&~m[2061]&m[2062])|(m[2037]&m[2058]&~m[2059]&~m[2061]&m[2062])|(m[2037]&~m[2058]&m[2059]&~m[2061]&m[2062])|(~m[2037]&~m[2058]&~m[2059]&m[2061]&m[2062])|(m[2037]&~m[2058]&~m[2059]&m[2061]&m[2062])|(~m[2037]&m[2058]&~m[2059]&m[2061]&m[2062])|(m[2037]&m[2058]&~m[2059]&m[2061]&m[2062])|(~m[2037]&~m[2058]&m[2059]&m[2061]&m[2062])|(m[2037]&~m[2058]&m[2059]&m[2061]&m[2062])|(m[2037]&m[2058]&m[2059]&m[2061]&m[2062]));
    m[2065] = (((m[2042]&~m[2063]&~m[2064]&~m[2066]&~m[2067])|(~m[2042]&~m[2063]&~m[2064]&m[2066]&~m[2067])|(m[2042]&m[2063]&~m[2064]&m[2066]&~m[2067])|(m[2042]&~m[2063]&m[2064]&m[2066]&~m[2067])|(~m[2042]&m[2063]&~m[2064]&~m[2066]&m[2067])|(~m[2042]&~m[2063]&m[2064]&~m[2066]&m[2067])|(m[2042]&m[2063]&m[2064]&~m[2066]&m[2067])|(~m[2042]&m[2063]&m[2064]&m[2066]&m[2067]))&UnbiasedRNG[483])|((m[2042]&~m[2063]&~m[2064]&m[2066]&~m[2067])|(~m[2042]&~m[2063]&~m[2064]&~m[2066]&m[2067])|(m[2042]&~m[2063]&~m[2064]&~m[2066]&m[2067])|(m[2042]&m[2063]&~m[2064]&~m[2066]&m[2067])|(m[2042]&~m[2063]&m[2064]&~m[2066]&m[2067])|(~m[2042]&~m[2063]&~m[2064]&m[2066]&m[2067])|(m[2042]&~m[2063]&~m[2064]&m[2066]&m[2067])|(~m[2042]&m[2063]&~m[2064]&m[2066]&m[2067])|(m[2042]&m[2063]&~m[2064]&m[2066]&m[2067])|(~m[2042]&~m[2063]&m[2064]&m[2066]&m[2067])|(m[2042]&~m[2063]&m[2064]&m[2066]&m[2067])|(m[2042]&m[2063]&m[2064]&m[2066]&m[2067]));
    m[2070] = (((m[2047]&~m[2068]&~m[2069]&~m[2071]&~m[2072])|(~m[2047]&~m[2068]&~m[2069]&m[2071]&~m[2072])|(m[2047]&m[2068]&~m[2069]&m[2071]&~m[2072])|(m[2047]&~m[2068]&m[2069]&m[2071]&~m[2072])|(~m[2047]&m[2068]&~m[2069]&~m[2071]&m[2072])|(~m[2047]&~m[2068]&m[2069]&~m[2071]&m[2072])|(m[2047]&m[2068]&m[2069]&~m[2071]&m[2072])|(~m[2047]&m[2068]&m[2069]&m[2071]&m[2072]))&UnbiasedRNG[484])|((m[2047]&~m[2068]&~m[2069]&m[2071]&~m[2072])|(~m[2047]&~m[2068]&~m[2069]&~m[2071]&m[2072])|(m[2047]&~m[2068]&~m[2069]&~m[2071]&m[2072])|(m[2047]&m[2068]&~m[2069]&~m[2071]&m[2072])|(m[2047]&~m[2068]&m[2069]&~m[2071]&m[2072])|(~m[2047]&~m[2068]&~m[2069]&m[2071]&m[2072])|(m[2047]&~m[2068]&~m[2069]&m[2071]&m[2072])|(~m[2047]&m[2068]&~m[2069]&m[2071]&m[2072])|(m[2047]&m[2068]&~m[2069]&m[2071]&m[2072])|(~m[2047]&~m[2068]&m[2069]&m[2071]&m[2072])|(m[2047]&~m[2068]&m[2069]&m[2071]&m[2072])|(m[2047]&m[2068]&m[2069]&m[2071]&m[2072]));
    m[2075] = (((m[2052]&~m[2073]&~m[2074]&~m[2076]&~m[2077])|(~m[2052]&~m[2073]&~m[2074]&m[2076]&~m[2077])|(m[2052]&m[2073]&~m[2074]&m[2076]&~m[2077])|(m[2052]&~m[2073]&m[2074]&m[2076]&~m[2077])|(~m[2052]&m[2073]&~m[2074]&~m[2076]&m[2077])|(~m[2052]&~m[2073]&m[2074]&~m[2076]&m[2077])|(m[2052]&m[2073]&m[2074]&~m[2076]&m[2077])|(~m[2052]&m[2073]&m[2074]&m[2076]&m[2077]))&UnbiasedRNG[485])|((m[2052]&~m[2073]&~m[2074]&m[2076]&~m[2077])|(~m[2052]&~m[2073]&~m[2074]&~m[2076]&m[2077])|(m[2052]&~m[2073]&~m[2074]&~m[2076]&m[2077])|(m[2052]&m[2073]&~m[2074]&~m[2076]&m[2077])|(m[2052]&~m[2073]&m[2074]&~m[2076]&m[2077])|(~m[2052]&~m[2073]&~m[2074]&m[2076]&m[2077])|(m[2052]&~m[2073]&~m[2074]&m[2076]&m[2077])|(~m[2052]&m[2073]&~m[2074]&m[2076]&m[2077])|(m[2052]&m[2073]&~m[2074]&m[2076]&m[2077])|(~m[2052]&~m[2073]&m[2074]&m[2076]&m[2077])|(m[2052]&~m[2073]&m[2074]&m[2076]&m[2077])|(m[2052]&m[2073]&m[2074]&m[2076]&m[2077]));
    m[2080] = (((m[2062]&~m[2078]&~m[2079]&~m[2081]&~m[2082])|(~m[2062]&~m[2078]&~m[2079]&m[2081]&~m[2082])|(m[2062]&m[2078]&~m[2079]&m[2081]&~m[2082])|(m[2062]&~m[2078]&m[2079]&m[2081]&~m[2082])|(~m[2062]&m[2078]&~m[2079]&~m[2081]&m[2082])|(~m[2062]&~m[2078]&m[2079]&~m[2081]&m[2082])|(m[2062]&m[2078]&m[2079]&~m[2081]&m[2082])|(~m[2062]&m[2078]&m[2079]&m[2081]&m[2082]))&UnbiasedRNG[486])|((m[2062]&~m[2078]&~m[2079]&m[2081]&~m[2082])|(~m[2062]&~m[2078]&~m[2079]&~m[2081]&m[2082])|(m[2062]&~m[2078]&~m[2079]&~m[2081]&m[2082])|(m[2062]&m[2078]&~m[2079]&~m[2081]&m[2082])|(m[2062]&~m[2078]&m[2079]&~m[2081]&m[2082])|(~m[2062]&~m[2078]&~m[2079]&m[2081]&m[2082])|(m[2062]&~m[2078]&~m[2079]&m[2081]&m[2082])|(~m[2062]&m[2078]&~m[2079]&m[2081]&m[2082])|(m[2062]&m[2078]&~m[2079]&m[2081]&m[2082])|(~m[2062]&~m[2078]&m[2079]&m[2081]&m[2082])|(m[2062]&~m[2078]&m[2079]&m[2081]&m[2082])|(m[2062]&m[2078]&m[2079]&m[2081]&m[2082]));
    m[2085] = (((m[2067]&~m[2083]&~m[2084]&~m[2086]&~m[2087])|(~m[2067]&~m[2083]&~m[2084]&m[2086]&~m[2087])|(m[2067]&m[2083]&~m[2084]&m[2086]&~m[2087])|(m[2067]&~m[2083]&m[2084]&m[2086]&~m[2087])|(~m[2067]&m[2083]&~m[2084]&~m[2086]&m[2087])|(~m[2067]&~m[2083]&m[2084]&~m[2086]&m[2087])|(m[2067]&m[2083]&m[2084]&~m[2086]&m[2087])|(~m[2067]&m[2083]&m[2084]&m[2086]&m[2087]))&UnbiasedRNG[487])|((m[2067]&~m[2083]&~m[2084]&m[2086]&~m[2087])|(~m[2067]&~m[2083]&~m[2084]&~m[2086]&m[2087])|(m[2067]&~m[2083]&~m[2084]&~m[2086]&m[2087])|(m[2067]&m[2083]&~m[2084]&~m[2086]&m[2087])|(m[2067]&~m[2083]&m[2084]&~m[2086]&m[2087])|(~m[2067]&~m[2083]&~m[2084]&m[2086]&m[2087])|(m[2067]&~m[2083]&~m[2084]&m[2086]&m[2087])|(~m[2067]&m[2083]&~m[2084]&m[2086]&m[2087])|(m[2067]&m[2083]&~m[2084]&m[2086]&m[2087])|(~m[2067]&~m[2083]&m[2084]&m[2086]&m[2087])|(m[2067]&~m[2083]&m[2084]&m[2086]&m[2087])|(m[2067]&m[2083]&m[2084]&m[2086]&m[2087]));
    m[2090] = (((m[2072]&~m[2088]&~m[2089]&~m[2091]&~m[2092])|(~m[2072]&~m[2088]&~m[2089]&m[2091]&~m[2092])|(m[2072]&m[2088]&~m[2089]&m[2091]&~m[2092])|(m[2072]&~m[2088]&m[2089]&m[2091]&~m[2092])|(~m[2072]&m[2088]&~m[2089]&~m[2091]&m[2092])|(~m[2072]&~m[2088]&m[2089]&~m[2091]&m[2092])|(m[2072]&m[2088]&m[2089]&~m[2091]&m[2092])|(~m[2072]&m[2088]&m[2089]&m[2091]&m[2092]))&UnbiasedRNG[488])|((m[2072]&~m[2088]&~m[2089]&m[2091]&~m[2092])|(~m[2072]&~m[2088]&~m[2089]&~m[2091]&m[2092])|(m[2072]&~m[2088]&~m[2089]&~m[2091]&m[2092])|(m[2072]&m[2088]&~m[2089]&~m[2091]&m[2092])|(m[2072]&~m[2088]&m[2089]&~m[2091]&m[2092])|(~m[2072]&~m[2088]&~m[2089]&m[2091]&m[2092])|(m[2072]&~m[2088]&~m[2089]&m[2091]&m[2092])|(~m[2072]&m[2088]&~m[2089]&m[2091]&m[2092])|(m[2072]&m[2088]&~m[2089]&m[2091]&m[2092])|(~m[2072]&~m[2088]&m[2089]&m[2091]&m[2092])|(m[2072]&~m[2088]&m[2089]&m[2091]&m[2092])|(m[2072]&m[2088]&m[2089]&m[2091]&m[2092]));
    m[2095] = (((m[2077]&~m[2093]&~m[2094]&~m[2096]&~m[2097])|(~m[2077]&~m[2093]&~m[2094]&m[2096]&~m[2097])|(m[2077]&m[2093]&~m[2094]&m[2096]&~m[2097])|(m[2077]&~m[2093]&m[2094]&m[2096]&~m[2097])|(~m[2077]&m[2093]&~m[2094]&~m[2096]&m[2097])|(~m[2077]&~m[2093]&m[2094]&~m[2096]&m[2097])|(m[2077]&m[2093]&m[2094]&~m[2096]&m[2097])|(~m[2077]&m[2093]&m[2094]&m[2096]&m[2097]))&UnbiasedRNG[489])|((m[2077]&~m[2093]&~m[2094]&m[2096]&~m[2097])|(~m[2077]&~m[2093]&~m[2094]&~m[2096]&m[2097])|(m[2077]&~m[2093]&~m[2094]&~m[2096]&m[2097])|(m[2077]&m[2093]&~m[2094]&~m[2096]&m[2097])|(m[2077]&~m[2093]&m[2094]&~m[2096]&m[2097])|(~m[2077]&~m[2093]&~m[2094]&m[2096]&m[2097])|(m[2077]&~m[2093]&~m[2094]&m[2096]&m[2097])|(~m[2077]&m[2093]&~m[2094]&m[2096]&m[2097])|(m[2077]&m[2093]&~m[2094]&m[2096]&m[2097])|(~m[2077]&~m[2093]&m[2094]&m[2096]&m[2097])|(m[2077]&~m[2093]&m[2094]&m[2096]&m[2097])|(m[2077]&m[2093]&m[2094]&m[2096]&m[2097]));
    m[2100] = (((m[2087]&~m[2098]&~m[2099]&~m[2101]&~m[2102])|(~m[2087]&~m[2098]&~m[2099]&m[2101]&~m[2102])|(m[2087]&m[2098]&~m[2099]&m[2101]&~m[2102])|(m[2087]&~m[2098]&m[2099]&m[2101]&~m[2102])|(~m[2087]&m[2098]&~m[2099]&~m[2101]&m[2102])|(~m[2087]&~m[2098]&m[2099]&~m[2101]&m[2102])|(m[2087]&m[2098]&m[2099]&~m[2101]&m[2102])|(~m[2087]&m[2098]&m[2099]&m[2101]&m[2102]))&UnbiasedRNG[490])|((m[2087]&~m[2098]&~m[2099]&m[2101]&~m[2102])|(~m[2087]&~m[2098]&~m[2099]&~m[2101]&m[2102])|(m[2087]&~m[2098]&~m[2099]&~m[2101]&m[2102])|(m[2087]&m[2098]&~m[2099]&~m[2101]&m[2102])|(m[2087]&~m[2098]&m[2099]&~m[2101]&m[2102])|(~m[2087]&~m[2098]&~m[2099]&m[2101]&m[2102])|(m[2087]&~m[2098]&~m[2099]&m[2101]&m[2102])|(~m[2087]&m[2098]&~m[2099]&m[2101]&m[2102])|(m[2087]&m[2098]&~m[2099]&m[2101]&m[2102])|(~m[2087]&~m[2098]&m[2099]&m[2101]&m[2102])|(m[2087]&~m[2098]&m[2099]&m[2101]&m[2102])|(m[2087]&m[2098]&m[2099]&m[2101]&m[2102]));
    m[2105] = (((m[2092]&~m[2103]&~m[2104]&~m[2106]&~m[2107])|(~m[2092]&~m[2103]&~m[2104]&m[2106]&~m[2107])|(m[2092]&m[2103]&~m[2104]&m[2106]&~m[2107])|(m[2092]&~m[2103]&m[2104]&m[2106]&~m[2107])|(~m[2092]&m[2103]&~m[2104]&~m[2106]&m[2107])|(~m[2092]&~m[2103]&m[2104]&~m[2106]&m[2107])|(m[2092]&m[2103]&m[2104]&~m[2106]&m[2107])|(~m[2092]&m[2103]&m[2104]&m[2106]&m[2107]))&UnbiasedRNG[491])|((m[2092]&~m[2103]&~m[2104]&m[2106]&~m[2107])|(~m[2092]&~m[2103]&~m[2104]&~m[2106]&m[2107])|(m[2092]&~m[2103]&~m[2104]&~m[2106]&m[2107])|(m[2092]&m[2103]&~m[2104]&~m[2106]&m[2107])|(m[2092]&~m[2103]&m[2104]&~m[2106]&m[2107])|(~m[2092]&~m[2103]&~m[2104]&m[2106]&m[2107])|(m[2092]&~m[2103]&~m[2104]&m[2106]&m[2107])|(~m[2092]&m[2103]&~m[2104]&m[2106]&m[2107])|(m[2092]&m[2103]&~m[2104]&m[2106]&m[2107])|(~m[2092]&~m[2103]&m[2104]&m[2106]&m[2107])|(m[2092]&~m[2103]&m[2104]&m[2106]&m[2107])|(m[2092]&m[2103]&m[2104]&m[2106]&m[2107]));
    m[2110] = (((m[2097]&~m[2108]&~m[2109]&~m[2111]&~m[2112])|(~m[2097]&~m[2108]&~m[2109]&m[2111]&~m[2112])|(m[2097]&m[2108]&~m[2109]&m[2111]&~m[2112])|(m[2097]&~m[2108]&m[2109]&m[2111]&~m[2112])|(~m[2097]&m[2108]&~m[2109]&~m[2111]&m[2112])|(~m[2097]&~m[2108]&m[2109]&~m[2111]&m[2112])|(m[2097]&m[2108]&m[2109]&~m[2111]&m[2112])|(~m[2097]&m[2108]&m[2109]&m[2111]&m[2112]))&UnbiasedRNG[492])|((m[2097]&~m[2108]&~m[2109]&m[2111]&~m[2112])|(~m[2097]&~m[2108]&~m[2109]&~m[2111]&m[2112])|(m[2097]&~m[2108]&~m[2109]&~m[2111]&m[2112])|(m[2097]&m[2108]&~m[2109]&~m[2111]&m[2112])|(m[2097]&~m[2108]&m[2109]&~m[2111]&m[2112])|(~m[2097]&~m[2108]&~m[2109]&m[2111]&m[2112])|(m[2097]&~m[2108]&~m[2109]&m[2111]&m[2112])|(~m[2097]&m[2108]&~m[2109]&m[2111]&m[2112])|(m[2097]&m[2108]&~m[2109]&m[2111]&m[2112])|(~m[2097]&~m[2108]&m[2109]&m[2111]&m[2112])|(m[2097]&~m[2108]&m[2109]&m[2111]&m[2112])|(m[2097]&m[2108]&m[2109]&m[2111]&m[2112]));
    m[2115] = (((m[2107]&~m[2113]&~m[2114]&~m[2116]&~m[2117])|(~m[2107]&~m[2113]&~m[2114]&m[2116]&~m[2117])|(m[2107]&m[2113]&~m[2114]&m[2116]&~m[2117])|(m[2107]&~m[2113]&m[2114]&m[2116]&~m[2117])|(~m[2107]&m[2113]&~m[2114]&~m[2116]&m[2117])|(~m[2107]&~m[2113]&m[2114]&~m[2116]&m[2117])|(m[2107]&m[2113]&m[2114]&~m[2116]&m[2117])|(~m[2107]&m[2113]&m[2114]&m[2116]&m[2117]))&UnbiasedRNG[493])|((m[2107]&~m[2113]&~m[2114]&m[2116]&~m[2117])|(~m[2107]&~m[2113]&~m[2114]&~m[2116]&m[2117])|(m[2107]&~m[2113]&~m[2114]&~m[2116]&m[2117])|(m[2107]&m[2113]&~m[2114]&~m[2116]&m[2117])|(m[2107]&~m[2113]&m[2114]&~m[2116]&m[2117])|(~m[2107]&~m[2113]&~m[2114]&m[2116]&m[2117])|(m[2107]&~m[2113]&~m[2114]&m[2116]&m[2117])|(~m[2107]&m[2113]&~m[2114]&m[2116]&m[2117])|(m[2107]&m[2113]&~m[2114]&m[2116]&m[2117])|(~m[2107]&~m[2113]&m[2114]&m[2116]&m[2117])|(m[2107]&~m[2113]&m[2114]&m[2116]&m[2117])|(m[2107]&m[2113]&m[2114]&m[2116]&m[2117]));
    m[2120] = (((m[2112]&~m[2118]&~m[2119]&~m[2121]&~m[2122])|(~m[2112]&~m[2118]&~m[2119]&m[2121]&~m[2122])|(m[2112]&m[2118]&~m[2119]&m[2121]&~m[2122])|(m[2112]&~m[2118]&m[2119]&m[2121]&~m[2122])|(~m[2112]&m[2118]&~m[2119]&~m[2121]&m[2122])|(~m[2112]&~m[2118]&m[2119]&~m[2121]&m[2122])|(m[2112]&m[2118]&m[2119]&~m[2121]&m[2122])|(~m[2112]&m[2118]&m[2119]&m[2121]&m[2122]))&UnbiasedRNG[494])|((m[2112]&~m[2118]&~m[2119]&m[2121]&~m[2122])|(~m[2112]&~m[2118]&~m[2119]&~m[2121]&m[2122])|(m[2112]&~m[2118]&~m[2119]&~m[2121]&m[2122])|(m[2112]&m[2118]&~m[2119]&~m[2121]&m[2122])|(m[2112]&~m[2118]&m[2119]&~m[2121]&m[2122])|(~m[2112]&~m[2118]&~m[2119]&m[2121]&m[2122])|(m[2112]&~m[2118]&~m[2119]&m[2121]&m[2122])|(~m[2112]&m[2118]&~m[2119]&m[2121]&m[2122])|(m[2112]&m[2118]&~m[2119]&m[2121]&m[2122])|(~m[2112]&~m[2118]&m[2119]&m[2121]&m[2122])|(m[2112]&~m[2118]&m[2119]&m[2121]&m[2122])|(m[2112]&m[2118]&m[2119]&m[2121]&m[2122]));
    m[2125] = (((m[2122]&~m[2123]&~m[2124]&~m[2126]&~m[2127])|(~m[2122]&~m[2123]&~m[2124]&m[2126]&~m[2127])|(m[2122]&m[2123]&~m[2124]&m[2126]&~m[2127])|(m[2122]&~m[2123]&m[2124]&m[2126]&~m[2127])|(~m[2122]&m[2123]&~m[2124]&~m[2126]&m[2127])|(~m[2122]&~m[2123]&m[2124]&~m[2126]&m[2127])|(m[2122]&m[2123]&m[2124]&~m[2126]&m[2127])|(~m[2122]&m[2123]&m[2124]&m[2126]&m[2127]))&UnbiasedRNG[495])|((m[2122]&~m[2123]&~m[2124]&m[2126]&~m[2127])|(~m[2122]&~m[2123]&~m[2124]&~m[2126]&m[2127])|(m[2122]&~m[2123]&~m[2124]&~m[2126]&m[2127])|(m[2122]&m[2123]&~m[2124]&~m[2126]&m[2127])|(m[2122]&~m[2123]&m[2124]&~m[2126]&m[2127])|(~m[2122]&~m[2123]&~m[2124]&m[2126]&m[2127])|(m[2122]&~m[2123]&~m[2124]&m[2126]&m[2127])|(~m[2122]&m[2123]&~m[2124]&m[2126]&m[2127])|(m[2122]&m[2123]&~m[2124]&m[2126]&m[2127])|(~m[2122]&~m[2123]&m[2124]&m[2126]&m[2127])|(m[2122]&~m[2123]&m[2124]&m[2126]&m[2127])|(m[2122]&m[2123]&m[2124]&m[2126]&m[2127]));
end

always @(posedge color2_clk) begin
    m[416] = (((~m[96]&~m[160]&~m[672])|(m[96]&m[160]&~m[672]))&BiasedRNG[639])|(((m[96]&~m[160]&~m[672])|(~m[96]&m[160]&m[672]))&~BiasedRNG[639])|((~m[96]&~m[160]&m[672])|(m[96]&~m[160]&m[672])|(m[96]&m[160]&m[672]));
    m[417] = (((~m[96]&~m[176]&~m[673])|(m[96]&m[176]&~m[673]))&BiasedRNG[640])|(((m[96]&~m[176]&~m[673])|(~m[96]&m[176]&m[673]))&~BiasedRNG[640])|((~m[96]&~m[176]&m[673])|(m[96]&~m[176]&m[673])|(m[96]&m[176]&m[673]));
    m[418] = (((~m[96]&~m[192]&~m[674])|(m[96]&m[192]&~m[674]))&BiasedRNG[641])|(((m[96]&~m[192]&~m[674])|(~m[96]&m[192]&m[674]))&~BiasedRNG[641])|((~m[96]&~m[192]&m[674])|(m[96]&~m[192]&m[674])|(m[96]&m[192]&m[674]));
    m[419] = (((~m[96]&~m[208]&~m[675])|(m[96]&m[208]&~m[675]))&BiasedRNG[642])|(((m[96]&~m[208]&~m[675])|(~m[96]&m[208]&m[675]))&~BiasedRNG[642])|((~m[96]&~m[208]&m[675])|(m[96]&~m[208]&m[675])|(m[96]&m[208]&m[675]));
    m[420] = (((~m[97]&~m[224]&~m[676])|(m[97]&m[224]&~m[676]))&BiasedRNG[643])|(((m[97]&~m[224]&~m[676])|(~m[97]&m[224]&m[676]))&~BiasedRNG[643])|((~m[97]&~m[224]&m[676])|(m[97]&~m[224]&m[676])|(m[97]&m[224]&m[676]));
    m[421] = (((~m[97]&~m[240]&~m[677])|(m[97]&m[240]&~m[677]))&BiasedRNG[644])|(((m[97]&~m[240]&~m[677])|(~m[97]&m[240]&m[677]))&~BiasedRNG[644])|((~m[97]&~m[240]&m[677])|(m[97]&~m[240]&m[677])|(m[97]&m[240]&m[677]));
    m[422] = (((~m[97]&~m[256]&~m[678])|(m[97]&m[256]&~m[678]))&BiasedRNG[645])|(((m[97]&~m[256]&~m[678])|(~m[97]&m[256]&m[678]))&~BiasedRNG[645])|((~m[97]&~m[256]&m[678])|(m[97]&~m[256]&m[678])|(m[97]&m[256]&m[678]));
    m[423] = (((~m[97]&~m[272]&~m[679])|(m[97]&m[272]&~m[679]))&BiasedRNG[646])|(((m[97]&~m[272]&~m[679])|(~m[97]&m[272]&m[679]))&~BiasedRNG[646])|((~m[97]&~m[272]&m[679])|(m[97]&~m[272]&m[679])|(m[97]&m[272]&m[679]));
    m[424] = (((~m[98]&~m[288]&~m[680])|(m[98]&m[288]&~m[680]))&BiasedRNG[647])|(((m[98]&~m[288]&~m[680])|(~m[98]&m[288]&m[680]))&~BiasedRNG[647])|((~m[98]&~m[288]&m[680])|(m[98]&~m[288]&m[680])|(m[98]&m[288]&m[680]));
    m[425] = (((~m[98]&~m[304]&~m[681])|(m[98]&m[304]&~m[681]))&BiasedRNG[648])|(((m[98]&~m[304]&~m[681])|(~m[98]&m[304]&m[681]))&~BiasedRNG[648])|((~m[98]&~m[304]&m[681])|(m[98]&~m[304]&m[681])|(m[98]&m[304]&m[681]));
    m[426] = (((~m[98]&~m[320]&~m[682])|(m[98]&m[320]&~m[682]))&BiasedRNG[649])|(((m[98]&~m[320]&~m[682])|(~m[98]&m[320]&m[682]))&~BiasedRNG[649])|((~m[98]&~m[320]&m[682])|(m[98]&~m[320]&m[682])|(m[98]&m[320]&m[682]));
    m[427] = (((~m[98]&~m[336]&~m[683])|(m[98]&m[336]&~m[683]))&BiasedRNG[650])|(((m[98]&~m[336]&~m[683])|(~m[98]&m[336]&m[683]))&~BiasedRNG[650])|((~m[98]&~m[336]&m[683])|(m[98]&~m[336]&m[683])|(m[98]&m[336]&m[683]));
    m[428] = (((~m[99]&~m[352]&~m[684])|(m[99]&m[352]&~m[684]))&BiasedRNG[651])|(((m[99]&~m[352]&~m[684])|(~m[99]&m[352]&m[684]))&~BiasedRNG[651])|((~m[99]&~m[352]&m[684])|(m[99]&~m[352]&m[684])|(m[99]&m[352]&m[684]));
    m[429] = (((~m[99]&~m[368]&~m[685])|(m[99]&m[368]&~m[685]))&BiasedRNG[652])|(((m[99]&~m[368]&~m[685])|(~m[99]&m[368]&m[685]))&~BiasedRNG[652])|((~m[99]&~m[368]&m[685])|(m[99]&~m[368]&m[685])|(m[99]&m[368]&m[685]));
    m[430] = (((~m[99]&~m[384]&~m[686])|(m[99]&m[384]&~m[686]))&BiasedRNG[653])|(((m[99]&~m[384]&~m[686])|(~m[99]&m[384]&m[686]))&~BiasedRNG[653])|((~m[99]&~m[384]&m[686])|(m[99]&~m[384]&m[686])|(m[99]&m[384]&m[686]));
    m[431] = (((~m[99]&~m[400]&~m[687])|(m[99]&m[400]&~m[687]))&BiasedRNG[654])|(((m[99]&~m[400]&~m[687])|(~m[99]&m[400]&m[687]))&~BiasedRNG[654])|((~m[99]&~m[400]&m[687])|(m[99]&~m[400]&m[687])|(m[99]&m[400]&m[687]));
    m[432] = (((~m[100]&~m[161]&~m[688])|(m[100]&m[161]&~m[688]))&BiasedRNG[655])|(((m[100]&~m[161]&~m[688])|(~m[100]&m[161]&m[688]))&~BiasedRNG[655])|((~m[100]&~m[161]&m[688])|(m[100]&~m[161]&m[688])|(m[100]&m[161]&m[688]));
    m[433] = (((~m[100]&~m[177]&~m[689])|(m[100]&m[177]&~m[689]))&BiasedRNG[656])|(((m[100]&~m[177]&~m[689])|(~m[100]&m[177]&m[689]))&~BiasedRNG[656])|((~m[100]&~m[177]&m[689])|(m[100]&~m[177]&m[689])|(m[100]&m[177]&m[689]));
    m[434] = (((~m[100]&~m[193]&~m[690])|(m[100]&m[193]&~m[690]))&BiasedRNG[657])|(((m[100]&~m[193]&~m[690])|(~m[100]&m[193]&m[690]))&~BiasedRNG[657])|((~m[100]&~m[193]&m[690])|(m[100]&~m[193]&m[690])|(m[100]&m[193]&m[690]));
    m[435] = (((~m[100]&~m[209]&~m[691])|(m[100]&m[209]&~m[691]))&BiasedRNG[658])|(((m[100]&~m[209]&~m[691])|(~m[100]&m[209]&m[691]))&~BiasedRNG[658])|((~m[100]&~m[209]&m[691])|(m[100]&~m[209]&m[691])|(m[100]&m[209]&m[691]));
    m[436] = (((~m[101]&~m[225]&~m[692])|(m[101]&m[225]&~m[692]))&BiasedRNG[659])|(((m[101]&~m[225]&~m[692])|(~m[101]&m[225]&m[692]))&~BiasedRNG[659])|((~m[101]&~m[225]&m[692])|(m[101]&~m[225]&m[692])|(m[101]&m[225]&m[692]));
    m[437] = (((~m[101]&~m[241]&~m[693])|(m[101]&m[241]&~m[693]))&BiasedRNG[660])|(((m[101]&~m[241]&~m[693])|(~m[101]&m[241]&m[693]))&~BiasedRNG[660])|((~m[101]&~m[241]&m[693])|(m[101]&~m[241]&m[693])|(m[101]&m[241]&m[693]));
    m[438] = (((~m[101]&~m[257]&~m[694])|(m[101]&m[257]&~m[694]))&BiasedRNG[661])|(((m[101]&~m[257]&~m[694])|(~m[101]&m[257]&m[694]))&~BiasedRNG[661])|((~m[101]&~m[257]&m[694])|(m[101]&~m[257]&m[694])|(m[101]&m[257]&m[694]));
    m[439] = (((~m[101]&~m[273]&~m[695])|(m[101]&m[273]&~m[695]))&BiasedRNG[662])|(((m[101]&~m[273]&~m[695])|(~m[101]&m[273]&m[695]))&~BiasedRNG[662])|((~m[101]&~m[273]&m[695])|(m[101]&~m[273]&m[695])|(m[101]&m[273]&m[695]));
    m[440] = (((~m[102]&~m[289]&~m[696])|(m[102]&m[289]&~m[696]))&BiasedRNG[663])|(((m[102]&~m[289]&~m[696])|(~m[102]&m[289]&m[696]))&~BiasedRNG[663])|((~m[102]&~m[289]&m[696])|(m[102]&~m[289]&m[696])|(m[102]&m[289]&m[696]));
    m[441] = (((~m[102]&~m[305]&~m[697])|(m[102]&m[305]&~m[697]))&BiasedRNG[664])|(((m[102]&~m[305]&~m[697])|(~m[102]&m[305]&m[697]))&~BiasedRNG[664])|((~m[102]&~m[305]&m[697])|(m[102]&~m[305]&m[697])|(m[102]&m[305]&m[697]));
    m[442] = (((~m[102]&~m[321]&~m[698])|(m[102]&m[321]&~m[698]))&BiasedRNG[665])|(((m[102]&~m[321]&~m[698])|(~m[102]&m[321]&m[698]))&~BiasedRNG[665])|((~m[102]&~m[321]&m[698])|(m[102]&~m[321]&m[698])|(m[102]&m[321]&m[698]));
    m[443] = (((~m[102]&~m[337]&~m[699])|(m[102]&m[337]&~m[699]))&BiasedRNG[666])|(((m[102]&~m[337]&~m[699])|(~m[102]&m[337]&m[699]))&~BiasedRNG[666])|((~m[102]&~m[337]&m[699])|(m[102]&~m[337]&m[699])|(m[102]&m[337]&m[699]));
    m[444] = (((~m[103]&~m[353]&~m[700])|(m[103]&m[353]&~m[700]))&BiasedRNG[667])|(((m[103]&~m[353]&~m[700])|(~m[103]&m[353]&m[700]))&~BiasedRNG[667])|((~m[103]&~m[353]&m[700])|(m[103]&~m[353]&m[700])|(m[103]&m[353]&m[700]));
    m[445] = (((~m[103]&~m[369]&~m[701])|(m[103]&m[369]&~m[701]))&BiasedRNG[668])|(((m[103]&~m[369]&~m[701])|(~m[103]&m[369]&m[701]))&~BiasedRNG[668])|((~m[103]&~m[369]&m[701])|(m[103]&~m[369]&m[701])|(m[103]&m[369]&m[701]));
    m[446] = (((~m[103]&~m[385]&~m[702])|(m[103]&m[385]&~m[702]))&BiasedRNG[669])|(((m[103]&~m[385]&~m[702])|(~m[103]&m[385]&m[702]))&~BiasedRNG[669])|((~m[103]&~m[385]&m[702])|(m[103]&~m[385]&m[702])|(m[103]&m[385]&m[702]));
    m[447] = (((~m[103]&~m[401]&~m[703])|(m[103]&m[401]&~m[703]))&BiasedRNG[670])|(((m[103]&~m[401]&~m[703])|(~m[103]&m[401]&m[703]))&~BiasedRNG[670])|((~m[103]&~m[401]&m[703])|(m[103]&~m[401]&m[703])|(m[103]&m[401]&m[703]));
    m[448] = (((~m[104]&~m[162]&~m[704])|(m[104]&m[162]&~m[704]))&BiasedRNG[671])|(((m[104]&~m[162]&~m[704])|(~m[104]&m[162]&m[704]))&~BiasedRNG[671])|((~m[104]&~m[162]&m[704])|(m[104]&~m[162]&m[704])|(m[104]&m[162]&m[704]));
    m[449] = (((~m[104]&~m[178]&~m[705])|(m[104]&m[178]&~m[705]))&BiasedRNG[672])|(((m[104]&~m[178]&~m[705])|(~m[104]&m[178]&m[705]))&~BiasedRNG[672])|((~m[104]&~m[178]&m[705])|(m[104]&~m[178]&m[705])|(m[104]&m[178]&m[705]));
    m[450] = (((~m[104]&~m[194]&~m[706])|(m[104]&m[194]&~m[706]))&BiasedRNG[673])|(((m[104]&~m[194]&~m[706])|(~m[104]&m[194]&m[706]))&~BiasedRNG[673])|((~m[104]&~m[194]&m[706])|(m[104]&~m[194]&m[706])|(m[104]&m[194]&m[706]));
    m[451] = (((~m[104]&~m[210]&~m[707])|(m[104]&m[210]&~m[707]))&BiasedRNG[674])|(((m[104]&~m[210]&~m[707])|(~m[104]&m[210]&m[707]))&~BiasedRNG[674])|((~m[104]&~m[210]&m[707])|(m[104]&~m[210]&m[707])|(m[104]&m[210]&m[707]));
    m[452] = (((~m[105]&~m[226]&~m[708])|(m[105]&m[226]&~m[708]))&BiasedRNG[675])|(((m[105]&~m[226]&~m[708])|(~m[105]&m[226]&m[708]))&~BiasedRNG[675])|((~m[105]&~m[226]&m[708])|(m[105]&~m[226]&m[708])|(m[105]&m[226]&m[708]));
    m[453] = (((~m[105]&~m[242]&~m[709])|(m[105]&m[242]&~m[709]))&BiasedRNG[676])|(((m[105]&~m[242]&~m[709])|(~m[105]&m[242]&m[709]))&~BiasedRNG[676])|((~m[105]&~m[242]&m[709])|(m[105]&~m[242]&m[709])|(m[105]&m[242]&m[709]));
    m[454] = (((~m[105]&~m[258]&~m[710])|(m[105]&m[258]&~m[710]))&BiasedRNG[677])|(((m[105]&~m[258]&~m[710])|(~m[105]&m[258]&m[710]))&~BiasedRNG[677])|((~m[105]&~m[258]&m[710])|(m[105]&~m[258]&m[710])|(m[105]&m[258]&m[710]));
    m[455] = (((~m[105]&~m[274]&~m[711])|(m[105]&m[274]&~m[711]))&BiasedRNG[678])|(((m[105]&~m[274]&~m[711])|(~m[105]&m[274]&m[711]))&~BiasedRNG[678])|((~m[105]&~m[274]&m[711])|(m[105]&~m[274]&m[711])|(m[105]&m[274]&m[711]));
    m[456] = (((~m[106]&~m[290]&~m[712])|(m[106]&m[290]&~m[712]))&BiasedRNG[679])|(((m[106]&~m[290]&~m[712])|(~m[106]&m[290]&m[712]))&~BiasedRNG[679])|((~m[106]&~m[290]&m[712])|(m[106]&~m[290]&m[712])|(m[106]&m[290]&m[712]));
    m[457] = (((~m[106]&~m[306]&~m[713])|(m[106]&m[306]&~m[713]))&BiasedRNG[680])|(((m[106]&~m[306]&~m[713])|(~m[106]&m[306]&m[713]))&~BiasedRNG[680])|((~m[106]&~m[306]&m[713])|(m[106]&~m[306]&m[713])|(m[106]&m[306]&m[713]));
    m[458] = (((~m[106]&~m[322]&~m[714])|(m[106]&m[322]&~m[714]))&BiasedRNG[681])|(((m[106]&~m[322]&~m[714])|(~m[106]&m[322]&m[714]))&~BiasedRNG[681])|((~m[106]&~m[322]&m[714])|(m[106]&~m[322]&m[714])|(m[106]&m[322]&m[714]));
    m[459] = (((~m[106]&~m[338]&~m[715])|(m[106]&m[338]&~m[715]))&BiasedRNG[682])|(((m[106]&~m[338]&~m[715])|(~m[106]&m[338]&m[715]))&~BiasedRNG[682])|((~m[106]&~m[338]&m[715])|(m[106]&~m[338]&m[715])|(m[106]&m[338]&m[715]));
    m[460] = (((~m[107]&~m[354]&~m[716])|(m[107]&m[354]&~m[716]))&BiasedRNG[683])|(((m[107]&~m[354]&~m[716])|(~m[107]&m[354]&m[716]))&~BiasedRNG[683])|((~m[107]&~m[354]&m[716])|(m[107]&~m[354]&m[716])|(m[107]&m[354]&m[716]));
    m[461] = (((~m[107]&~m[370]&~m[717])|(m[107]&m[370]&~m[717]))&BiasedRNG[684])|(((m[107]&~m[370]&~m[717])|(~m[107]&m[370]&m[717]))&~BiasedRNG[684])|((~m[107]&~m[370]&m[717])|(m[107]&~m[370]&m[717])|(m[107]&m[370]&m[717]));
    m[462] = (((~m[107]&~m[386]&~m[718])|(m[107]&m[386]&~m[718]))&BiasedRNG[685])|(((m[107]&~m[386]&~m[718])|(~m[107]&m[386]&m[718]))&~BiasedRNG[685])|((~m[107]&~m[386]&m[718])|(m[107]&~m[386]&m[718])|(m[107]&m[386]&m[718]));
    m[463] = (((~m[107]&~m[402]&~m[719])|(m[107]&m[402]&~m[719]))&BiasedRNG[686])|(((m[107]&~m[402]&~m[719])|(~m[107]&m[402]&m[719]))&~BiasedRNG[686])|((~m[107]&~m[402]&m[719])|(m[107]&~m[402]&m[719])|(m[107]&m[402]&m[719]));
    m[464] = (((~m[108]&~m[163]&~m[720])|(m[108]&m[163]&~m[720]))&BiasedRNG[687])|(((m[108]&~m[163]&~m[720])|(~m[108]&m[163]&m[720]))&~BiasedRNG[687])|((~m[108]&~m[163]&m[720])|(m[108]&~m[163]&m[720])|(m[108]&m[163]&m[720]));
    m[465] = (((~m[108]&~m[179]&~m[721])|(m[108]&m[179]&~m[721]))&BiasedRNG[688])|(((m[108]&~m[179]&~m[721])|(~m[108]&m[179]&m[721]))&~BiasedRNG[688])|((~m[108]&~m[179]&m[721])|(m[108]&~m[179]&m[721])|(m[108]&m[179]&m[721]));
    m[466] = (((~m[108]&~m[195]&~m[722])|(m[108]&m[195]&~m[722]))&BiasedRNG[689])|(((m[108]&~m[195]&~m[722])|(~m[108]&m[195]&m[722]))&~BiasedRNG[689])|((~m[108]&~m[195]&m[722])|(m[108]&~m[195]&m[722])|(m[108]&m[195]&m[722]));
    m[467] = (((~m[108]&~m[211]&~m[723])|(m[108]&m[211]&~m[723]))&BiasedRNG[690])|(((m[108]&~m[211]&~m[723])|(~m[108]&m[211]&m[723]))&~BiasedRNG[690])|((~m[108]&~m[211]&m[723])|(m[108]&~m[211]&m[723])|(m[108]&m[211]&m[723]));
    m[468] = (((~m[109]&~m[227]&~m[724])|(m[109]&m[227]&~m[724]))&BiasedRNG[691])|(((m[109]&~m[227]&~m[724])|(~m[109]&m[227]&m[724]))&~BiasedRNG[691])|((~m[109]&~m[227]&m[724])|(m[109]&~m[227]&m[724])|(m[109]&m[227]&m[724]));
    m[469] = (((~m[109]&~m[243]&~m[725])|(m[109]&m[243]&~m[725]))&BiasedRNG[692])|(((m[109]&~m[243]&~m[725])|(~m[109]&m[243]&m[725]))&~BiasedRNG[692])|((~m[109]&~m[243]&m[725])|(m[109]&~m[243]&m[725])|(m[109]&m[243]&m[725]));
    m[470] = (((~m[109]&~m[259]&~m[726])|(m[109]&m[259]&~m[726]))&BiasedRNG[693])|(((m[109]&~m[259]&~m[726])|(~m[109]&m[259]&m[726]))&~BiasedRNG[693])|((~m[109]&~m[259]&m[726])|(m[109]&~m[259]&m[726])|(m[109]&m[259]&m[726]));
    m[471] = (((~m[109]&~m[275]&~m[727])|(m[109]&m[275]&~m[727]))&BiasedRNG[694])|(((m[109]&~m[275]&~m[727])|(~m[109]&m[275]&m[727]))&~BiasedRNG[694])|((~m[109]&~m[275]&m[727])|(m[109]&~m[275]&m[727])|(m[109]&m[275]&m[727]));
    m[472] = (((~m[110]&~m[291]&~m[728])|(m[110]&m[291]&~m[728]))&BiasedRNG[695])|(((m[110]&~m[291]&~m[728])|(~m[110]&m[291]&m[728]))&~BiasedRNG[695])|((~m[110]&~m[291]&m[728])|(m[110]&~m[291]&m[728])|(m[110]&m[291]&m[728]));
    m[473] = (((~m[110]&~m[307]&~m[729])|(m[110]&m[307]&~m[729]))&BiasedRNG[696])|(((m[110]&~m[307]&~m[729])|(~m[110]&m[307]&m[729]))&~BiasedRNG[696])|((~m[110]&~m[307]&m[729])|(m[110]&~m[307]&m[729])|(m[110]&m[307]&m[729]));
    m[474] = (((~m[110]&~m[323]&~m[730])|(m[110]&m[323]&~m[730]))&BiasedRNG[697])|(((m[110]&~m[323]&~m[730])|(~m[110]&m[323]&m[730]))&~BiasedRNG[697])|((~m[110]&~m[323]&m[730])|(m[110]&~m[323]&m[730])|(m[110]&m[323]&m[730]));
    m[475] = (((~m[110]&~m[339]&~m[731])|(m[110]&m[339]&~m[731]))&BiasedRNG[698])|(((m[110]&~m[339]&~m[731])|(~m[110]&m[339]&m[731]))&~BiasedRNG[698])|((~m[110]&~m[339]&m[731])|(m[110]&~m[339]&m[731])|(m[110]&m[339]&m[731]));
    m[476] = (((~m[111]&~m[355]&~m[732])|(m[111]&m[355]&~m[732]))&BiasedRNG[699])|(((m[111]&~m[355]&~m[732])|(~m[111]&m[355]&m[732]))&~BiasedRNG[699])|((~m[111]&~m[355]&m[732])|(m[111]&~m[355]&m[732])|(m[111]&m[355]&m[732]));
    m[477] = (((~m[111]&~m[371]&~m[733])|(m[111]&m[371]&~m[733]))&BiasedRNG[700])|(((m[111]&~m[371]&~m[733])|(~m[111]&m[371]&m[733]))&~BiasedRNG[700])|((~m[111]&~m[371]&m[733])|(m[111]&~m[371]&m[733])|(m[111]&m[371]&m[733]));
    m[478] = (((~m[111]&~m[387]&~m[734])|(m[111]&m[387]&~m[734]))&BiasedRNG[701])|(((m[111]&~m[387]&~m[734])|(~m[111]&m[387]&m[734]))&~BiasedRNG[701])|((~m[111]&~m[387]&m[734])|(m[111]&~m[387]&m[734])|(m[111]&m[387]&m[734]));
    m[479] = (((~m[111]&~m[403]&~m[735])|(m[111]&m[403]&~m[735]))&BiasedRNG[702])|(((m[111]&~m[403]&~m[735])|(~m[111]&m[403]&m[735]))&~BiasedRNG[702])|((~m[111]&~m[403]&m[735])|(m[111]&~m[403]&m[735])|(m[111]&m[403]&m[735]));
    m[480] = (((~m[112]&~m[164]&~m[736])|(m[112]&m[164]&~m[736]))&BiasedRNG[703])|(((m[112]&~m[164]&~m[736])|(~m[112]&m[164]&m[736]))&~BiasedRNG[703])|((~m[112]&~m[164]&m[736])|(m[112]&~m[164]&m[736])|(m[112]&m[164]&m[736]));
    m[481] = (((~m[112]&~m[180]&~m[737])|(m[112]&m[180]&~m[737]))&BiasedRNG[704])|(((m[112]&~m[180]&~m[737])|(~m[112]&m[180]&m[737]))&~BiasedRNG[704])|((~m[112]&~m[180]&m[737])|(m[112]&~m[180]&m[737])|(m[112]&m[180]&m[737]));
    m[482] = (((~m[112]&~m[196]&~m[738])|(m[112]&m[196]&~m[738]))&BiasedRNG[705])|(((m[112]&~m[196]&~m[738])|(~m[112]&m[196]&m[738]))&~BiasedRNG[705])|((~m[112]&~m[196]&m[738])|(m[112]&~m[196]&m[738])|(m[112]&m[196]&m[738]));
    m[483] = (((~m[112]&~m[212]&~m[739])|(m[112]&m[212]&~m[739]))&BiasedRNG[706])|(((m[112]&~m[212]&~m[739])|(~m[112]&m[212]&m[739]))&~BiasedRNG[706])|((~m[112]&~m[212]&m[739])|(m[112]&~m[212]&m[739])|(m[112]&m[212]&m[739]));
    m[484] = (((~m[113]&~m[228]&~m[740])|(m[113]&m[228]&~m[740]))&BiasedRNG[707])|(((m[113]&~m[228]&~m[740])|(~m[113]&m[228]&m[740]))&~BiasedRNG[707])|((~m[113]&~m[228]&m[740])|(m[113]&~m[228]&m[740])|(m[113]&m[228]&m[740]));
    m[485] = (((~m[113]&~m[244]&~m[741])|(m[113]&m[244]&~m[741]))&BiasedRNG[708])|(((m[113]&~m[244]&~m[741])|(~m[113]&m[244]&m[741]))&~BiasedRNG[708])|((~m[113]&~m[244]&m[741])|(m[113]&~m[244]&m[741])|(m[113]&m[244]&m[741]));
    m[486] = (((~m[113]&~m[260]&~m[742])|(m[113]&m[260]&~m[742]))&BiasedRNG[709])|(((m[113]&~m[260]&~m[742])|(~m[113]&m[260]&m[742]))&~BiasedRNG[709])|((~m[113]&~m[260]&m[742])|(m[113]&~m[260]&m[742])|(m[113]&m[260]&m[742]));
    m[487] = (((~m[113]&~m[276]&~m[743])|(m[113]&m[276]&~m[743]))&BiasedRNG[710])|(((m[113]&~m[276]&~m[743])|(~m[113]&m[276]&m[743]))&~BiasedRNG[710])|((~m[113]&~m[276]&m[743])|(m[113]&~m[276]&m[743])|(m[113]&m[276]&m[743]));
    m[488] = (((~m[114]&~m[292]&~m[744])|(m[114]&m[292]&~m[744]))&BiasedRNG[711])|(((m[114]&~m[292]&~m[744])|(~m[114]&m[292]&m[744]))&~BiasedRNG[711])|((~m[114]&~m[292]&m[744])|(m[114]&~m[292]&m[744])|(m[114]&m[292]&m[744]));
    m[489] = (((~m[114]&~m[308]&~m[745])|(m[114]&m[308]&~m[745]))&BiasedRNG[712])|(((m[114]&~m[308]&~m[745])|(~m[114]&m[308]&m[745]))&~BiasedRNG[712])|((~m[114]&~m[308]&m[745])|(m[114]&~m[308]&m[745])|(m[114]&m[308]&m[745]));
    m[490] = (((~m[114]&~m[324]&~m[746])|(m[114]&m[324]&~m[746]))&BiasedRNG[713])|(((m[114]&~m[324]&~m[746])|(~m[114]&m[324]&m[746]))&~BiasedRNG[713])|((~m[114]&~m[324]&m[746])|(m[114]&~m[324]&m[746])|(m[114]&m[324]&m[746]));
    m[491] = (((~m[114]&~m[340]&~m[747])|(m[114]&m[340]&~m[747]))&BiasedRNG[714])|(((m[114]&~m[340]&~m[747])|(~m[114]&m[340]&m[747]))&~BiasedRNG[714])|((~m[114]&~m[340]&m[747])|(m[114]&~m[340]&m[747])|(m[114]&m[340]&m[747]));
    m[492] = (((~m[115]&~m[356]&~m[748])|(m[115]&m[356]&~m[748]))&BiasedRNG[715])|(((m[115]&~m[356]&~m[748])|(~m[115]&m[356]&m[748]))&~BiasedRNG[715])|((~m[115]&~m[356]&m[748])|(m[115]&~m[356]&m[748])|(m[115]&m[356]&m[748]));
    m[493] = (((~m[115]&~m[372]&~m[749])|(m[115]&m[372]&~m[749]))&BiasedRNG[716])|(((m[115]&~m[372]&~m[749])|(~m[115]&m[372]&m[749]))&~BiasedRNG[716])|((~m[115]&~m[372]&m[749])|(m[115]&~m[372]&m[749])|(m[115]&m[372]&m[749]));
    m[494] = (((~m[115]&~m[388]&~m[750])|(m[115]&m[388]&~m[750]))&BiasedRNG[717])|(((m[115]&~m[388]&~m[750])|(~m[115]&m[388]&m[750]))&~BiasedRNG[717])|((~m[115]&~m[388]&m[750])|(m[115]&~m[388]&m[750])|(m[115]&m[388]&m[750]));
    m[495] = (((~m[115]&~m[404]&~m[751])|(m[115]&m[404]&~m[751]))&BiasedRNG[718])|(((m[115]&~m[404]&~m[751])|(~m[115]&m[404]&m[751]))&~BiasedRNG[718])|((~m[115]&~m[404]&m[751])|(m[115]&~m[404]&m[751])|(m[115]&m[404]&m[751]));
    m[496] = (((~m[116]&~m[165]&~m[752])|(m[116]&m[165]&~m[752]))&BiasedRNG[719])|(((m[116]&~m[165]&~m[752])|(~m[116]&m[165]&m[752]))&~BiasedRNG[719])|((~m[116]&~m[165]&m[752])|(m[116]&~m[165]&m[752])|(m[116]&m[165]&m[752]));
    m[497] = (((~m[116]&~m[181]&~m[753])|(m[116]&m[181]&~m[753]))&BiasedRNG[720])|(((m[116]&~m[181]&~m[753])|(~m[116]&m[181]&m[753]))&~BiasedRNG[720])|((~m[116]&~m[181]&m[753])|(m[116]&~m[181]&m[753])|(m[116]&m[181]&m[753]));
    m[498] = (((~m[116]&~m[197]&~m[754])|(m[116]&m[197]&~m[754]))&BiasedRNG[721])|(((m[116]&~m[197]&~m[754])|(~m[116]&m[197]&m[754]))&~BiasedRNG[721])|((~m[116]&~m[197]&m[754])|(m[116]&~m[197]&m[754])|(m[116]&m[197]&m[754]));
    m[499] = (((~m[116]&~m[213]&~m[755])|(m[116]&m[213]&~m[755]))&BiasedRNG[722])|(((m[116]&~m[213]&~m[755])|(~m[116]&m[213]&m[755]))&~BiasedRNG[722])|((~m[116]&~m[213]&m[755])|(m[116]&~m[213]&m[755])|(m[116]&m[213]&m[755]));
    m[500] = (((~m[117]&~m[229]&~m[756])|(m[117]&m[229]&~m[756]))&BiasedRNG[723])|(((m[117]&~m[229]&~m[756])|(~m[117]&m[229]&m[756]))&~BiasedRNG[723])|((~m[117]&~m[229]&m[756])|(m[117]&~m[229]&m[756])|(m[117]&m[229]&m[756]));
    m[501] = (((~m[117]&~m[245]&~m[757])|(m[117]&m[245]&~m[757]))&BiasedRNG[724])|(((m[117]&~m[245]&~m[757])|(~m[117]&m[245]&m[757]))&~BiasedRNG[724])|((~m[117]&~m[245]&m[757])|(m[117]&~m[245]&m[757])|(m[117]&m[245]&m[757]));
    m[502] = (((~m[117]&~m[261]&~m[758])|(m[117]&m[261]&~m[758]))&BiasedRNG[725])|(((m[117]&~m[261]&~m[758])|(~m[117]&m[261]&m[758]))&~BiasedRNG[725])|((~m[117]&~m[261]&m[758])|(m[117]&~m[261]&m[758])|(m[117]&m[261]&m[758]));
    m[503] = (((~m[117]&~m[277]&~m[759])|(m[117]&m[277]&~m[759]))&BiasedRNG[726])|(((m[117]&~m[277]&~m[759])|(~m[117]&m[277]&m[759]))&~BiasedRNG[726])|((~m[117]&~m[277]&m[759])|(m[117]&~m[277]&m[759])|(m[117]&m[277]&m[759]));
    m[504] = (((~m[118]&~m[293]&~m[760])|(m[118]&m[293]&~m[760]))&BiasedRNG[727])|(((m[118]&~m[293]&~m[760])|(~m[118]&m[293]&m[760]))&~BiasedRNG[727])|((~m[118]&~m[293]&m[760])|(m[118]&~m[293]&m[760])|(m[118]&m[293]&m[760]));
    m[505] = (((~m[118]&~m[309]&~m[761])|(m[118]&m[309]&~m[761]))&BiasedRNG[728])|(((m[118]&~m[309]&~m[761])|(~m[118]&m[309]&m[761]))&~BiasedRNG[728])|((~m[118]&~m[309]&m[761])|(m[118]&~m[309]&m[761])|(m[118]&m[309]&m[761]));
    m[506] = (((~m[118]&~m[325]&~m[762])|(m[118]&m[325]&~m[762]))&BiasedRNG[729])|(((m[118]&~m[325]&~m[762])|(~m[118]&m[325]&m[762]))&~BiasedRNG[729])|((~m[118]&~m[325]&m[762])|(m[118]&~m[325]&m[762])|(m[118]&m[325]&m[762]));
    m[507] = (((~m[118]&~m[341]&~m[763])|(m[118]&m[341]&~m[763]))&BiasedRNG[730])|(((m[118]&~m[341]&~m[763])|(~m[118]&m[341]&m[763]))&~BiasedRNG[730])|((~m[118]&~m[341]&m[763])|(m[118]&~m[341]&m[763])|(m[118]&m[341]&m[763]));
    m[508] = (((~m[119]&~m[357]&~m[764])|(m[119]&m[357]&~m[764]))&BiasedRNG[731])|(((m[119]&~m[357]&~m[764])|(~m[119]&m[357]&m[764]))&~BiasedRNG[731])|((~m[119]&~m[357]&m[764])|(m[119]&~m[357]&m[764])|(m[119]&m[357]&m[764]));
    m[509] = (((~m[119]&~m[373]&~m[765])|(m[119]&m[373]&~m[765]))&BiasedRNG[732])|(((m[119]&~m[373]&~m[765])|(~m[119]&m[373]&m[765]))&~BiasedRNG[732])|((~m[119]&~m[373]&m[765])|(m[119]&~m[373]&m[765])|(m[119]&m[373]&m[765]));
    m[510] = (((~m[119]&~m[389]&~m[766])|(m[119]&m[389]&~m[766]))&BiasedRNG[733])|(((m[119]&~m[389]&~m[766])|(~m[119]&m[389]&m[766]))&~BiasedRNG[733])|((~m[119]&~m[389]&m[766])|(m[119]&~m[389]&m[766])|(m[119]&m[389]&m[766]));
    m[511] = (((~m[119]&~m[405]&~m[767])|(m[119]&m[405]&~m[767]))&BiasedRNG[734])|(((m[119]&~m[405]&~m[767])|(~m[119]&m[405]&m[767]))&~BiasedRNG[734])|((~m[119]&~m[405]&m[767])|(m[119]&~m[405]&m[767])|(m[119]&m[405]&m[767]));
    m[512] = (((~m[120]&~m[166]&~m[768])|(m[120]&m[166]&~m[768]))&BiasedRNG[735])|(((m[120]&~m[166]&~m[768])|(~m[120]&m[166]&m[768]))&~BiasedRNG[735])|((~m[120]&~m[166]&m[768])|(m[120]&~m[166]&m[768])|(m[120]&m[166]&m[768]));
    m[513] = (((~m[120]&~m[182]&~m[769])|(m[120]&m[182]&~m[769]))&BiasedRNG[736])|(((m[120]&~m[182]&~m[769])|(~m[120]&m[182]&m[769]))&~BiasedRNG[736])|((~m[120]&~m[182]&m[769])|(m[120]&~m[182]&m[769])|(m[120]&m[182]&m[769]));
    m[514] = (((~m[120]&~m[198]&~m[770])|(m[120]&m[198]&~m[770]))&BiasedRNG[737])|(((m[120]&~m[198]&~m[770])|(~m[120]&m[198]&m[770]))&~BiasedRNG[737])|((~m[120]&~m[198]&m[770])|(m[120]&~m[198]&m[770])|(m[120]&m[198]&m[770]));
    m[515] = (((~m[120]&~m[214]&~m[771])|(m[120]&m[214]&~m[771]))&BiasedRNG[738])|(((m[120]&~m[214]&~m[771])|(~m[120]&m[214]&m[771]))&~BiasedRNG[738])|((~m[120]&~m[214]&m[771])|(m[120]&~m[214]&m[771])|(m[120]&m[214]&m[771]));
    m[516] = (((~m[121]&~m[230]&~m[772])|(m[121]&m[230]&~m[772]))&BiasedRNG[739])|(((m[121]&~m[230]&~m[772])|(~m[121]&m[230]&m[772]))&~BiasedRNG[739])|((~m[121]&~m[230]&m[772])|(m[121]&~m[230]&m[772])|(m[121]&m[230]&m[772]));
    m[517] = (((~m[121]&~m[246]&~m[773])|(m[121]&m[246]&~m[773]))&BiasedRNG[740])|(((m[121]&~m[246]&~m[773])|(~m[121]&m[246]&m[773]))&~BiasedRNG[740])|((~m[121]&~m[246]&m[773])|(m[121]&~m[246]&m[773])|(m[121]&m[246]&m[773]));
    m[518] = (((~m[121]&~m[262]&~m[774])|(m[121]&m[262]&~m[774]))&BiasedRNG[741])|(((m[121]&~m[262]&~m[774])|(~m[121]&m[262]&m[774]))&~BiasedRNG[741])|((~m[121]&~m[262]&m[774])|(m[121]&~m[262]&m[774])|(m[121]&m[262]&m[774]));
    m[519] = (((~m[121]&~m[278]&~m[775])|(m[121]&m[278]&~m[775]))&BiasedRNG[742])|(((m[121]&~m[278]&~m[775])|(~m[121]&m[278]&m[775]))&~BiasedRNG[742])|((~m[121]&~m[278]&m[775])|(m[121]&~m[278]&m[775])|(m[121]&m[278]&m[775]));
    m[520] = (((~m[122]&~m[294]&~m[776])|(m[122]&m[294]&~m[776]))&BiasedRNG[743])|(((m[122]&~m[294]&~m[776])|(~m[122]&m[294]&m[776]))&~BiasedRNG[743])|((~m[122]&~m[294]&m[776])|(m[122]&~m[294]&m[776])|(m[122]&m[294]&m[776]));
    m[521] = (((~m[122]&~m[310]&~m[777])|(m[122]&m[310]&~m[777]))&BiasedRNG[744])|(((m[122]&~m[310]&~m[777])|(~m[122]&m[310]&m[777]))&~BiasedRNG[744])|((~m[122]&~m[310]&m[777])|(m[122]&~m[310]&m[777])|(m[122]&m[310]&m[777]));
    m[522] = (((~m[122]&~m[326]&~m[778])|(m[122]&m[326]&~m[778]))&BiasedRNG[745])|(((m[122]&~m[326]&~m[778])|(~m[122]&m[326]&m[778]))&~BiasedRNG[745])|((~m[122]&~m[326]&m[778])|(m[122]&~m[326]&m[778])|(m[122]&m[326]&m[778]));
    m[523] = (((~m[122]&~m[342]&~m[779])|(m[122]&m[342]&~m[779]))&BiasedRNG[746])|(((m[122]&~m[342]&~m[779])|(~m[122]&m[342]&m[779]))&~BiasedRNG[746])|((~m[122]&~m[342]&m[779])|(m[122]&~m[342]&m[779])|(m[122]&m[342]&m[779]));
    m[524] = (((~m[123]&~m[358]&~m[780])|(m[123]&m[358]&~m[780]))&BiasedRNG[747])|(((m[123]&~m[358]&~m[780])|(~m[123]&m[358]&m[780]))&~BiasedRNG[747])|((~m[123]&~m[358]&m[780])|(m[123]&~m[358]&m[780])|(m[123]&m[358]&m[780]));
    m[525] = (((~m[123]&~m[374]&~m[781])|(m[123]&m[374]&~m[781]))&BiasedRNG[748])|(((m[123]&~m[374]&~m[781])|(~m[123]&m[374]&m[781]))&~BiasedRNG[748])|((~m[123]&~m[374]&m[781])|(m[123]&~m[374]&m[781])|(m[123]&m[374]&m[781]));
    m[526] = (((~m[123]&~m[390]&~m[782])|(m[123]&m[390]&~m[782]))&BiasedRNG[749])|(((m[123]&~m[390]&~m[782])|(~m[123]&m[390]&m[782]))&~BiasedRNG[749])|((~m[123]&~m[390]&m[782])|(m[123]&~m[390]&m[782])|(m[123]&m[390]&m[782]));
    m[527] = (((~m[123]&~m[406]&~m[783])|(m[123]&m[406]&~m[783]))&BiasedRNG[750])|(((m[123]&~m[406]&~m[783])|(~m[123]&m[406]&m[783]))&~BiasedRNG[750])|((~m[123]&~m[406]&m[783])|(m[123]&~m[406]&m[783])|(m[123]&m[406]&m[783]));
    m[528] = (((~m[124]&~m[167]&~m[784])|(m[124]&m[167]&~m[784]))&BiasedRNG[751])|(((m[124]&~m[167]&~m[784])|(~m[124]&m[167]&m[784]))&~BiasedRNG[751])|((~m[124]&~m[167]&m[784])|(m[124]&~m[167]&m[784])|(m[124]&m[167]&m[784]));
    m[529] = (((~m[124]&~m[183]&~m[785])|(m[124]&m[183]&~m[785]))&BiasedRNG[752])|(((m[124]&~m[183]&~m[785])|(~m[124]&m[183]&m[785]))&~BiasedRNG[752])|((~m[124]&~m[183]&m[785])|(m[124]&~m[183]&m[785])|(m[124]&m[183]&m[785]));
    m[530] = (((~m[124]&~m[199]&~m[786])|(m[124]&m[199]&~m[786]))&BiasedRNG[753])|(((m[124]&~m[199]&~m[786])|(~m[124]&m[199]&m[786]))&~BiasedRNG[753])|((~m[124]&~m[199]&m[786])|(m[124]&~m[199]&m[786])|(m[124]&m[199]&m[786]));
    m[531] = (((~m[124]&~m[215]&~m[787])|(m[124]&m[215]&~m[787]))&BiasedRNG[754])|(((m[124]&~m[215]&~m[787])|(~m[124]&m[215]&m[787]))&~BiasedRNG[754])|((~m[124]&~m[215]&m[787])|(m[124]&~m[215]&m[787])|(m[124]&m[215]&m[787]));
    m[532] = (((~m[125]&~m[231]&~m[788])|(m[125]&m[231]&~m[788]))&BiasedRNG[755])|(((m[125]&~m[231]&~m[788])|(~m[125]&m[231]&m[788]))&~BiasedRNG[755])|((~m[125]&~m[231]&m[788])|(m[125]&~m[231]&m[788])|(m[125]&m[231]&m[788]));
    m[533] = (((~m[125]&~m[247]&~m[789])|(m[125]&m[247]&~m[789]))&BiasedRNG[756])|(((m[125]&~m[247]&~m[789])|(~m[125]&m[247]&m[789]))&~BiasedRNG[756])|((~m[125]&~m[247]&m[789])|(m[125]&~m[247]&m[789])|(m[125]&m[247]&m[789]));
    m[534] = (((~m[125]&~m[263]&~m[790])|(m[125]&m[263]&~m[790]))&BiasedRNG[757])|(((m[125]&~m[263]&~m[790])|(~m[125]&m[263]&m[790]))&~BiasedRNG[757])|((~m[125]&~m[263]&m[790])|(m[125]&~m[263]&m[790])|(m[125]&m[263]&m[790]));
    m[535] = (((~m[125]&~m[279]&~m[791])|(m[125]&m[279]&~m[791]))&BiasedRNG[758])|(((m[125]&~m[279]&~m[791])|(~m[125]&m[279]&m[791]))&~BiasedRNG[758])|((~m[125]&~m[279]&m[791])|(m[125]&~m[279]&m[791])|(m[125]&m[279]&m[791]));
    m[536] = (((~m[126]&~m[295]&~m[792])|(m[126]&m[295]&~m[792]))&BiasedRNG[759])|(((m[126]&~m[295]&~m[792])|(~m[126]&m[295]&m[792]))&~BiasedRNG[759])|((~m[126]&~m[295]&m[792])|(m[126]&~m[295]&m[792])|(m[126]&m[295]&m[792]));
    m[537] = (((~m[126]&~m[311]&~m[793])|(m[126]&m[311]&~m[793]))&BiasedRNG[760])|(((m[126]&~m[311]&~m[793])|(~m[126]&m[311]&m[793]))&~BiasedRNG[760])|((~m[126]&~m[311]&m[793])|(m[126]&~m[311]&m[793])|(m[126]&m[311]&m[793]));
    m[538] = (((~m[126]&~m[327]&~m[794])|(m[126]&m[327]&~m[794]))&BiasedRNG[761])|(((m[126]&~m[327]&~m[794])|(~m[126]&m[327]&m[794]))&~BiasedRNG[761])|((~m[126]&~m[327]&m[794])|(m[126]&~m[327]&m[794])|(m[126]&m[327]&m[794]));
    m[539] = (((~m[126]&~m[343]&~m[795])|(m[126]&m[343]&~m[795]))&BiasedRNG[762])|(((m[126]&~m[343]&~m[795])|(~m[126]&m[343]&m[795]))&~BiasedRNG[762])|((~m[126]&~m[343]&m[795])|(m[126]&~m[343]&m[795])|(m[126]&m[343]&m[795]));
    m[540] = (((~m[127]&~m[359]&~m[796])|(m[127]&m[359]&~m[796]))&BiasedRNG[763])|(((m[127]&~m[359]&~m[796])|(~m[127]&m[359]&m[796]))&~BiasedRNG[763])|((~m[127]&~m[359]&m[796])|(m[127]&~m[359]&m[796])|(m[127]&m[359]&m[796]));
    m[541] = (((~m[127]&~m[375]&~m[797])|(m[127]&m[375]&~m[797]))&BiasedRNG[764])|(((m[127]&~m[375]&~m[797])|(~m[127]&m[375]&m[797]))&~BiasedRNG[764])|((~m[127]&~m[375]&m[797])|(m[127]&~m[375]&m[797])|(m[127]&m[375]&m[797]));
    m[542] = (((~m[127]&~m[391]&~m[798])|(m[127]&m[391]&~m[798]))&BiasedRNG[765])|(((m[127]&~m[391]&~m[798])|(~m[127]&m[391]&m[798]))&~BiasedRNG[765])|((~m[127]&~m[391]&m[798])|(m[127]&~m[391]&m[798])|(m[127]&m[391]&m[798]));
    m[543] = (((~m[127]&~m[407]&~m[799])|(m[127]&m[407]&~m[799]))&BiasedRNG[766])|(((m[127]&~m[407]&~m[799])|(~m[127]&m[407]&m[799]))&~BiasedRNG[766])|((~m[127]&~m[407]&m[799])|(m[127]&~m[407]&m[799])|(m[127]&m[407]&m[799]));
    m[544] = (((~m[128]&~m[168]&~m[800])|(m[128]&m[168]&~m[800]))&BiasedRNG[767])|(((m[128]&~m[168]&~m[800])|(~m[128]&m[168]&m[800]))&~BiasedRNG[767])|((~m[128]&~m[168]&m[800])|(m[128]&~m[168]&m[800])|(m[128]&m[168]&m[800]));
    m[545] = (((~m[128]&~m[184]&~m[801])|(m[128]&m[184]&~m[801]))&BiasedRNG[768])|(((m[128]&~m[184]&~m[801])|(~m[128]&m[184]&m[801]))&~BiasedRNG[768])|((~m[128]&~m[184]&m[801])|(m[128]&~m[184]&m[801])|(m[128]&m[184]&m[801]));
    m[546] = (((~m[128]&~m[200]&~m[802])|(m[128]&m[200]&~m[802]))&BiasedRNG[769])|(((m[128]&~m[200]&~m[802])|(~m[128]&m[200]&m[802]))&~BiasedRNG[769])|((~m[128]&~m[200]&m[802])|(m[128]&~m[200]&m[802])|(m[128]&m[200]&m[802]));
    m[547] = (((~m[128]&~m[216]&~m[803])|(m[128]&m[216]&~m[803]))&BiasedRNG[770])|(((m[128]&~m[216]&~m[803])|(~m[128]&m[216]&m[803]))&~BiasedRNG[770])|((~m[128]&~m[216]&m[803])|(m[128]&~m[216]&m[803])|(m[128]&m[216]&m[803]));
    m[548] = (((~m[129]&~m[232]&~m[804])|(m[129]&m[232]&~m[804]))&BiasedRNG[771])|(((m[129]&~m[232]&~m[804])|(~m[129]&m[232]&m[804]))&~BiasedRNG[771])|((~m[129]&~m[232]&m[804])|(m[129]&~m[232]&m[804])|(m[129]&m[232]&m[804]));
    m[549] = (((~m[129]&~m[248]&~m[805])|(m[129]&m[248]&~m[805]))&BiasedRNG[772])|(((m[129]&~m[248]&~m[805])|(~m[129]&m[248]&m[805]))&~BiasedRNG[772])|((~m[129]&~m[248]&m[805])|(m[129]&~m[248]&m[805])|(m[129]&m[248]&m[805]));
    m[550] = (((~m[129]&~m[264]&~m[806])|(m[129]&m[264]&~m[806]))&BiasedRNG[773])|(((m[129]&~m[264]&~m[806])|(~m[129]&m[264]&m[806]))&~BiasedRNG[773])|((~m[129]&~m[264]&m[806])|(m[129]&~m[264]&m[806])|(m[129]&m[264]&m[806]));
    m[551] = (((~m[129]&~m[280]&~m[807])|(m[129]&m[280]&~m[807]))&BiasedRNG[774])|(((m[129]&~m[280]&~m[807])|(~m[129]&m[280]&m[807]))&~BiasedRNG[774])|((~m[129]&~m[280]&m[807])|(m[129]&~m[280]&m[807])|(m[129]&m[280]&m[807]));
    m[552] = (((~m[130]&~m[296]&~m[808])|(m[130]&m[296]&~m[808]))&BiasedRNG[775])|(((m[130]&~m[296]&~m[808])|(~m[130]&m[296]&m[808]))&~BiasedRNG[775])|((~m[130]&~m[296]&m[808])|(m[130]&~m[296]&m[808])|(m[130]&m[296]&m[808]));
    m[553] = (((~m[130]&~m[312]&~m[809])|(m[130]&m[312]&~m[809]))&BiasedRNG[776])|(((m[130]&~m[312]&~m[809])|(~m[130]&m[312]&m[809]))&~BiasedRNG[776])|((~m[130]&~m[312]&m[809])|(m[130]&~m[312]&m[809])|(m[130]&m[312]&m[809]));
    m[554] = (((~m[130]&~m[328]&~m[810])|(m[130]&m[328]&~m[810]))&BiasedRNG[777])|(((m[130]&~m[328]&~m[810])|(~m[130]&m[328]&m[810]))&~BiasedRNG[777])|((~m[130]&~m[328]&m[810])|(m[130]&~m[328]&m[810])|(m[130]&m[328]&m[810]));
    m[555] = (((~m[130]&~m[344]&~m[811])|(m[130]&m[344]&~m[811]))&BiasedRNG[778])|(((m[130]&~m[344]&~m[811])|(~m[130]&m[344]&m[811]))&~BiasedRNG[778])|((~m[130]&~m[344]&m[811])|(m[130]&~m[344]&m[811])|(m[130]&m[344]&m[811]));
    m[556] = (((~m[131]&~m[360]&~m[812])|(m[131]&m[360]&~m[812]))&BiasedRNG[779])|(((m[131]&~m[360]&~m[812])|(~m[131]&m[360]&m[812]))&~BiasedRNG[779])|((~m[131]&~m[360]&m[812])|(m[131]&~m[360]&m[812])|(m[131]&m[360]&m[812]));
    m[557] = (((~m[131]&~m[376]&~m[813])|(m[131]&m[376]&~m[813]))&BiasedRNG[780])|(((m[131]&~m[376]&~m[813])|(~m[131]&m[376]&m[813]))&~BiasedRNG[780])|((~m[131]&~m[376]&m[813])|(m[131]&~m[376]&m[813])|(m[131]&m[376]&m[813]));
    m[558] = (((~m[131]&~m[392]&~m[814])|(m[131]&m[392]&~m[814]))&BiasedRNG[781])|(((m[131]&~m[392]&~m[814])|(~m[131]&m[392]&m[814]))&~BiasedRNG[781])|((~m[131]&~m[392]&m[814])|(m[131]&~m[392]&m[814])|(m[131]&m[392]&m[814]));
    m[559] = (((~m[131]&~m[408]&~m[815])|(m[131]&m[408]&~m[815]))&BiasedRNG[782])|(((m[131]&~m[408]&~m[815])|(~m[131]&m[408]&m[815]))&~BiasedRNG[782])|((~m[131]&~m[408]&m[815])|(m[131]&~m[408]&m[815])|(m[131]&m[408]&m[815]));
    m[560] = (((~m[132]&~m[169]&~m[816])|(m[132]&m[169]&~m[816]))&BiasedRNG[783])|(((m[132]&~m[169]&~m[816])|(~m[132]&m[169]&m[816]))&~BiasedRNG[783])|((~m[132]&~m[169]&m[816])|(m[132]&~m[169]&m[816])|(m[132]&m[169]&m[816]));
    m[561] = (((~m[132]&~m[185]&~m[817])|(m[132]&m[185]&~m[817]))&BiasedRNG[784])|(((m[132]&~m[185]&~m[817])|(~m[132]&m[185]&m[817]))&~BiasedRNG[784])|((~m[132]&~m[185]&m[817])|(m[132]&~m[185]&m[817])|(m[132]&m[185]&m[817]));
    m[562] = (((~m[132]&~m[201]&~m[818])|(m[132]&m[201]&~m[818]))&BiasedRNG[785])|(((m[132]&~m[201]&~m[818])|(~m[132]&m[201]&m[818]))&~BiasedRNG[785])|((~m[132]&~m[201]&m[818])|(m[132]&~m[201]&m[818])|(m[132]&m[201]&m[818]));
    m[563] = (((~m[132]&~m[217]&~m[819])|(m[132]&m[217]&~m[819]))&BiasedRNG[786])|(((m[132]&~m[217]&~m[819])|(~m[132]&m[217]&m[819]))&~BiasedRNG[786])|((~m[132]&~m[217]&m[819])|(m[132]&~m[217]&m[819])|(m[132]&m[217]&m[819]));
    m[564] = (((~m[133]&~m[233]&~m[820])|(m[133]&m[233]&~m[820]))&BiasedRNG[787])|(((m[133]&~m[233]&~m[820])|(~m[133]&m[233]&m[820]))&~BiasedRNG[787])|((~m[133]&~m[233]&m[820])|(m[133]&~m[233]&m[820])|(m[133]&m[233]&m[820]));
    m[565] = (((~m[133]&~m[249]&~m[821])|(m[133]&m[249]&~m[821]))&BiasedRNG[788])|(((m[133]&~m[249]&~m[821])|(~m[133]&m[249]&m[821]))&~BiasedRNG[788])|((~m[133]&~m[249]&m[821])|(m[133]&~m[249]&m[821])|(m[133]&m[249]&m[821]));
    m[566] = (((~m[133]&~m[265]&~m[822])|(m[133]&m[265]&~m[822]))&BiasedRNG[789])|(((m[133]&~m[265]&~m[822])|(~m[133]&m[265]&m[822]))&~BiasedRNG[789])|((~m[133]&~m[265]&m[822])|(m[133]&~m[265]&m[822])|(m[133]&m[265]&m[822]));
    m[567] = (((~m[133]&~m[281]&~m[823])|(m[133]&m[281]&~m[823]))&BiasedRNG[790])|(((m[133]&~m[281]&~m[823])|(~m[133]&m[281]&m[823]))&~BiasedRNG[790])|((~m[133]&~m[281]&m[823])|(m[133]&~m[281]&m[823])|(m[133]&m[281]&m[823]));
    m[568] = (((~m[134]&~m[297]&~m[824])|(m[134]&m[297]&~m[824]))&BiasedRNG[791])|(((m[134]&~m[297]&~m[824])|(~m[134]&m[297]&m[824]))&~BiasedRNG[791])|((~m[134]&~m[297]&m[824])|(m[134]&~m[297]&m[824])|(m[134]&m[297]&m[824]));
    m[569] = (((~m[134]&~m[313]&~m[825])|(m[134]&m[313]&~m[825]))&BiasedRNG[792])|(((m[134]&~m[313]&~m[825])|(~m[134]&m[313]&m[825]))&~BiasedRNG[792])|((~m[134]&~m[313]&m[825])|(m[134]&~m[313]&m[825])|(m[134]&m[313]&m[825]));
    m[570] = (((~m[134]&~m[329]&~m[826])|(m[134]&m[329]&~m[826]))&BiasedRNG[793])|(((m[134]&~m[329]&~m[826])|(~m[134]&m[329]&m[826]))&~BiasedRNG[793])|((~m[134]&~m[329]&m[826])|(m[134]&~m[329]&m[826])|(m[134]&m[329]&m[826]));
    m[571] = (((~m[134]&~m[345]&~m[827])|(m[134]&m[345]&~m[827]))&BiasedRNG[794])|(((m[134]&~m[345]&~m[827])|(~m[134]&m[345]&m[827]))&~BiasedRNG[794])|((~m[134]&~m[345]&m[827])|(m[134]&~m[345]&m[827])|(m[134]&m[345]&m[827]));
    m[572] = (((~m[135]&~m[361]&~m[828])|(m[135]&m[361]&~m[828]))&BiasedRNG[795])|(((m[135]&~m[361]&~m[828])|(~m[135]&m[361]&m[828]))&~BiasedRNG[795])|((~m[135]&~m[361]&m[828])|(m[135]&~m[361]&m[828])|(m[135]&m[361]&m[828]));
    m[573] = (((~m[135]&~m[377]&~m[829])|(m[135]&m[377]&~m[829]))&BiasedRNG[796])|(((m[135]&~m[377]&~m[829])|(~m[135]&m[377]&m[829]))&~BiasedRNG[796])|((~m[135]&~m[377]&m[829])|(m[135]&~m[377]&m[829])|(m[135]&m[377]&m[829]));
    m[574] = (((~m[135]&~m[393]&~m[830])|(m[135]&m[393]&~m[830]))&BiasedRNG[797])|(((m[135]&~m[393]&~m[830])|(~m[135]&m[393]&m[830]))&~BiasedRNG[797])|((~m[135]&~m[393]&m[830])|(m[135]&~m[393]&m[830])|(m[135]&m[393]&m[830]));
    m[575] = (((~m[135]&~m[409]&~m[831])|(m[135]&m[409]&~m[831]))&BiasedRNG[798])|(((m[135]&~m[409]&~m[831])|(~m[135]&m[409]&m[831]))&~BiasedRNG[798])|((~m[135]&~m[409]&m[831])|(m[135]&~m[409]&m[831])|(m[135]&m[409]&m[831]));
    m[576] = (((~m[136]&~m[170]&~m[832])|(m[136]&m[170]&~m[832]))&BiasedRNG[799])|(((m[136]&~m[170]&~m[832])|(~m[136]&m[170]&m[832]))&~BiasedRNG[799])|((~m[136]&~m[170]&m[832])|(m[136]&~m[170]&m[832])|(m[136]&m[170]&m[832]));
    m[577] = (((~m[136]&~m[186]&~m[833])|(m[136]&m[186]&~m[833]))&BiasedRNG[800])|(((m[136]&~m[186]&~m[833])|(~m[136]&m[186]&m[833]))&~BiasedRNG[800])|((~m[136]&~m[186]&m[833])|(m[136]&~m[186]&m[833])|(m[136]&m[186]&m[833]));
    m[578] = (((~m[136]&~m[202]&~m[834])|(m[136]&m[202]&~m[834]))&BiasedRNG[801])|(((m[136]&~m[202]&~m[834])|(~m[136]&m[202]&m[834]))&~BiasedRNG[801])|((~m[136]&~m[202]&m[834])|(m[136]&~m[202]&m[834])|(m[136]&m[202]&m[834]));
    m[579] = (((~m[136]&~m[218]&~m[835])|(m[136]&m[218]&~m[835]))&BiasedRNG[802])|(((m[136]&~m[218]&~m[835])|(~m[136]&m[218]&m[835]))&~BiasedRNG[802])|((~m[136]&~m[218]&m[835])|(m[136]&~m[218]&m[835])|(m[136]&m[218]&m[835]));
    m[580] = (((~m[137]&~m[234]&~m[836])|(m[137]&m[234]&~m[836]))&BiasedRNG[803])|(((m[137]&~m[234]&~m[836])|(~m[137]&m[234]&m[836]))&~BiasedRNG[803])|((~m[137]&~m[234]&m[836])|(m[137]&~m[234]&m[836])|(m[137]&m[234]&m[836]));
    m[581] = (((~m[137]&~m[250]&~m[837])|(m[137]&m[250]&~m[837]))&BiasedRNG[804])|(((m[137]&~m[250]&~m[837])|(~m[137]&m[250]&m[837]))&~BiasedRNG[804])|((~m[137]&~m[250]&m[837])|(m[137]&~m[250]&m[837])|(m[137]&m[250]&m[837]));
    m[582] = (((~m[137]&~m[266]&~m[838])|(m[137]&m[266]&~m[838]))&BiasedRNG[805])|(((m[137]&~m[266]&~m[838])|(~m[137]&m[266]&m[838]))&~BiasedRNG[805])|((~m[137]&~m[266]&m[838])|(m[137]&~m[266]&m[838])|(m[137]&m[266]&m[838]));
    m[583] = (((~m[137]&~m[282]&~m[839])|(m[137]&m[282]&~m[839]))&BiasedRNG[806])|(((m[137]&~m[282]&~m[839])|(~m[137]&m[282]&m[839]))&~BiasedRNG[806])|((~m[137]&~m[282]&m[839])|(m[137]&~m[282]&m[839])|(m[137]&m[282]&m[839]));
    m[584] = (((~m[138]&~m[298]&~m[840])|(m[138]&m[298]&~m[840]))&BiasedRNG[807])|(((m[138]&~m[298]&~m[840])|(~m[138]&m[298]&m[840]))&~BiasedRNG[807])|((~m[138]&~m[298]&m[840])|(m[138]&~m[298]&m[840])|(m[138]&m[298]&m[840]));
    m[585] = (((~m[138]&~m[314]&~m[841])|(m[138]&m[314]&~m[841]))&BiasedRNG[808])|(((m[138]&~m[314]&~m[841])|(~m[138]&m[314]&m[841]))&~BiasedRNG[808])|((~m[138]&~m[314]&m[841])|(m[138]&~m[314]&m[841])|(m[138]&m[314]&m[841]));
    m[586] = (((~m[138]&~m[330]&~m[842])|(m[138]&m[330]&~m[842]))&BiasedRNG[809])|(((m[138]&~m[330]&~m[842])|(~m[138]&m[330]&m[842]))&~BiasedRNG[809])|((~m[138]&~m[330]&m[842])|(m[138]&~m[330]&m[842])|(m[138]&m[330]&m[842]));
    m[587] = (((~m[138]&~m[346]&~m[843])|(m[138]&m[346]&~m[843]))&BiasedRNG[810])|(((m[138]&~m[346]&~m[843])|(~m[138]&m[346]&m[843]))&~BiasedRNG[810])|((~m[138]&~m[346]&m[843])|(m[138]&~m[346]&m[843])|(m[138]&m[346]&m[843]));
    m[588] = (((~m[139]&~m[362]&~m[844])|(m[139]&m[362]&~m[844]))&BiasedRNG[811])|(((m[139]&~m[362]&~m[844])|(~m[139]&m[362]&m[844]))&~BiasedRNG[811])|((~m[139]&~m[362]&m[844])|(m[139]&~m[362]&m[844])|(m[139]&m[362]&m[844]));
    m[589] = (((~m[139]&~m[378]&~m[845])|(m[139]&m[378]&~m[845]))&BiasedRNG[812])|(((m[139]&~m[378]&~m[845])|(~m[139]&m[378]&m[845]))&~BiasedRNG[812])|((~m[139]&~m[378]&m[845])|(m[139]&~m[378]&m[845])|(m[139]&m[378]&m[845]));
    m[590] = (((~m[139]&~m[394]&~m[846])|(m[139]&m[394]&~m[846]))&BiasedRNG[813])|(((m[139]&~m[394]&~m[846])|(~m[139]&m[394]&m[846]))&~BiasedRNG[813])|((~m[139]&~m[394]&m[846])|(m[139]&~m[394]&m[846])|(m[139]&m[394]&m[846]));
    m[591] = (((~m[139]&~m[410]&~m[847])|(m[139]&m[410]&~m[847]))&BiasedRNG[814])|(((m[139]&~m[410]&~m[847])|(~m[139]&m[410]&m[847]))&~BiasedRNG[814])|((~m[139]&~m[410]&m[847])|(m[139]&~m[410]&m[847])|(m[139]&m[410]&m[847]));
    m[592] = (((~m[140]&~m[171]&~m[848])|(m[140]&m[171]&~m[848]))&BiasedRNG[815])|(((m[140]&~m[171]&~m[848])|(~m[140]&m[171]&m[848]))&~BiasedRNG[815])|((~m[140]&~m[171]&m[848])|(m[140]&~m[171]&m[848])|(m[140]&m[171]&m[848]));
    m[593] = (((~m[140]&~m[187]&~m[849])|(m[140]&m[187]&~m[849]))&BiasedRNG[816])|(((m[140]&~m[187]&~m[849])|(~m[140]&m[187]&m[849]))&~BiasedRNG[816])|((~m[140]&~m[187]&m[849])|(m[140]&~m[187]&m[849])|(m[140]&m[187]&m[849]));
    m[594] = (((~m[140]&~m[203]&~m[850])|(m[140]&m[203]&~m[850]))&BiasedRNG[817])|(((m[140]&~m[203]&~m[850])|(~m[140]&m[203]&m[850]))&~BiasedRNG[817])|((~m[140]&~m[203]&m[850])|(m[140]&~m[203]&m[850])|(m[140]&m[203]&m[850]));
    m[595] = (((~m[140]&~m[219]&~m[851])|(m[140]&m[219]&~m[851]))&BiasedRNG[818])|(((m[140]&~m[219]&~m[851])|(~m[140]&m[219]&m[851]))&~BiasedRNG[818])|((~m[140]&~m[219]&m[851])|(m[140]&~m[219]&m[851])|(m[140]&m[219]&m[851]));
    m[596] = (((~m[141]&~m[235]&~m[852])|(m[141]&m[235]&~m[852]))&BiasedRNG[819])|(((m[141]&~m[235]&~m[852])|(~m[141]&m[235]&m[852]))&~BiasedRNG[819])|((~m[141]&~m[235]&m[852])|(m[141]&~m[235]&m[852])|(m[141]&m[235]&m[852]));
    m[597] = (((~m[141]&~m[251]&~m[853])|(m[141]&m[251]&~m[853]))&BiasedRNG[820])|(((m[141]&~m[251]&~m[853])|(~m[141]&m[251]&m[853]))&~BiasedRNG[820])|((~m[141]&~m[251]&m[853])|(m[141]&~m[251]&m[853])|(m[141]&m[251]&m[853]));
    m[598] = (((~m[141]&~m[267]&~m[854])|(m[141]&m[267]&~m[854]))&BiasedRNG[821])|(((m[141]&~m[267]&~m[854])|(~m[141]&m[267]&m[854]))&~BiasedRNG[821])|((~m[141]&~m[267]&m[854])|(m[141]&~m[267]&m[854])|(m[141]&m[267]&m[854]));
    m[599] = (((~m[141]&~m[283]&~m[855])|(m[141]&m[283]&~m[855]))&BiasedRNG[822])|(((m[141]&~m[283]&~m[855])|(~m[141]&m[283]&m[855]))&~BiasedRNG[822])|((~m[141]&~m[283]&m[855])|(m[141]&~m[283]&m[855])|(m[141]&m[283]&m[855]));
    m[600] = (((~m[142]&~m[299]&~m[856])|(m[142]&m[299]&~m[856]))&BiasedRNG[823])|(((m[142]&~m[299]&~m[856])|(~m[142]&m[299]&m[856]))&~BiasedRNG[823])|((~m[142]&~m[299]&m[856])|(m[142]&~m[299]&m[856])|(m[142]&m[299]&m[856]));
    m[601] = (((~m[142]&~m[315]&~m[857])|(m[142]&m[315]&~m[857]))&BiasedRNG[824])|(((m[142]&~m[315]&~m[857])|(~m[142]&m[315]&m[857]))&~BiasedRNG[824])|((~m[142]&~m[315]&m[857])|(m[142]&~m[315]&m[857])|(m[142]&m[315]&m[857]));
    m[602] = (((~m[142]&~m[331]&~m[858])|(m[142]&m[331]&~m[858]))&BiasedRNG[825])|(((m[142]&~m[331]&~m[858])|(~m[142]&m[331]&m[858]))&~BiasedRNG[825])|((~m[142]&~m[331]&m[858])|(m[142]&~m[331]&m[858])|(m[142]&m[331]&m[858]));
    m[603] = (((~m[142]&~m[347]&~m[859])|(m[142]&m[347]&~m[859]))&BiasedRNG[826])|(((m[142]&~m[347]&~m[859])|(~m[142]&m[347]&m[859]))&~BiasedRNG[826])|((~m[142]&~m[347]&m[859])|(m[142]&~m[347]&m[859])|(m[142]&m[347]&m[859]));
    m[604] = (((~m[143]&~m[363]&~m[860])|(m[143]&m[363]&~m[860]))&BiasedRNG[827])|(((m[143]&~m[363]&~m[860])|(~m[143]&m[363]&m[860]))&~BiasedRNG[827])|((~m[143]&~m[363]&m[860])|(m[143]&~m[363]&m[860])|(m[143]&m[363]&m[860]));
    m[605] = (((~m[143]&~m[379]&~m[861])|(m[143]&m[379]&~m[861]))&BiasedRNG[828])|(((m[143]&~m[379]&~m[861])|(~m[143]&m[379]&m[861]))&~BiasedRNG[828])|((~m[143]&~m[379]&m[861])|(m[143]&~m[379]&m[861])|(m[143]&m[379]&m[861]));
    m[606] = (((~m[143]&~m[395]&~m[862])|(m[143]&m[395]&~m[862]))&BiasedRNG[829])|(((m[143]&~m[395]&~m[862])|(~m[143]&m[395]&m[862]))&~BiasedRNG[829])|((~m[143]&~m[395]&m[862])|(m[143]&~m[395]&m[862])|(m[143]&m[395]&m[862]));
    m[607] = (((~m[143]&~m[411]&~m[863])|(m[143]&m[411]&~m[863]))&BiasedRNG[830])|(((m[143]&~m[411]&~m[863])|(~m[143]&m[411]&m[863]))&~BiasedRNG[830])|((~m[143]&~m[411]&m[863])|(m[143]&~m[411]&m[863])|(m[143]&m[411]&m[863]));
    m[608] = (((~m[144]&~m[172]&~m[864])|(m[144]&m[172]&~m[864]))&BiasedRNG[831])|(((m[144]&~m[172]&~m[864])|(~m[144]&m[172]&m[864]))&~BiasedRNG[831])|((~m[144]&~m[172]&m[864])|(m[144]&~m[172]&m[864])|(m[144]&m[172]&m[864]));
    m[609] = (((~m[144]&~m[188]&~m[865])|(m[144]&m[188]&~m[865]))&BiasedRNG[832])|(((m[144]&~m[188]&~m[865])|(~m[144]&m[188]&m[865]))&~BiasedRNG[832])|((~m[144]&~m[188]&m[865])|(m[144]&~m[188]&m[865])|(m[144]&m[188]&m[865]));
    m[610] = (((~m[144]&~m[204]&~m[866])|(m[144]&m[204]&~m[866]))&BiasedRNG[833])|(((m[144]&~m[204]&~m[866])|(~m[144]&m[204]&m[866]))&~BiasedRNG[833])|((~m[144]&~m[204]&m[866])|(m[144]&~m[204]&m[866])|(m[144]&m[204]&m[866]));
    m[611] = (((~m[144]&~m[220]&~m[867])|(m[144]&m[220]&~m[867]))&BiasedRNG[834])|(((m[144]&~m[220]&~m[867])|(~m[144]&m[220]&m[867]))&~BiasedRNG[834])|((~m[144]&~m[220]&m[867])|(m[144]&~m[220]&m[867])|(m[144]&m[220]&m[867]));
    m[612] = (((~m[145]&~m[236]&~m[868])|(m[145]&m[236]&~m[868]))&BiasedRNG[835])|(((m[145]&~m[236]&~m[868])|(~m[145]&m[236]&m[868]))&~BiasedRNG[835])|((~m[145]&~m[236]&m[868])|(m[145]&~m[236]&m[868])|(m[145]&m[236]&m[868]));
    m[613] = (((~m[145]&~m[252]&~m[869])|(m[145]&m[252]&~m[869]))&BiasedRNG[836])|(((m[145]&~m[252]&~m[869])|(~m[145]&m[252]&m[869]))&~BiasedRNG[836])|((~m[145]&~m[252]&m[869])|(m[145]&~m[252]&m[869])|(m[145]&m[252]&m[869]));
    m[614] = (((~m[145]&~m[268]&~m[870])|(m[145]&m[268]&~m[870]))&BiasedRNG[837])|(((m[145]&~m[268]&~m[870])|(~m[145]&m[268]&m[870]))&~BiasedRNG[837])|((~m[145]&~m[268]&m[870])|(m[145]&~m[268]&m[870])|(m[145]&m[268]&m[870]));
    m[615] = (((~m[145]&~m[284]&~m[871])|(m[145]&m[284]&~m[871]))&BiasedRNG[838])|(((m[145]&~m[284]&~m[871])|(~m[145]&m[284]&m[871]))&~BiasedRNG[838])|((~m[145]&~m[284]&m[871])|(m[145]&~m[284]&m[871])|(m[145]&m[284]&m[871]));
    m[616] = (((~m[146]&~m[300]&~m[872])|(m[146]&m[300]&~m[872]))&BiasedRNG[839])|(((m[146]&~m[300]&~m[872])|(~m[146]&m[300]&m[872]))&~BiasedRNG[839])|((~m[146]&~m[300]&m[872])|(m[146]&~m[300]&m[872])|(m[146]&m[300]&m[872]));
    m[617] = (((~m[146]&~m[316]&~m[873])|(m[146]&m[316]&~m[873]))&BiasedRNG[840])|(((m[146]&~m[316]&~m[873])|(~m[146]&m[316]&m[873]))&~BiasedRNG[840])|((~m[146]&~m[316]&m[873])|(m[146]&~m[316]&m[873])|(m[146]&m[316]&m[873]));
    m[618] = (((~m[146]&~m[332]&~m[874])|(m[146]&m[332]&~m[874]))&BiasedRNG[841])|(((m[146]&~m[332]&~m[874])|(~m[146]&m[332]&m[874]))&~BiasedRNG[841])|((~m[146]&~m[332]&m[874])|(m[146]&~m[332]&m[874])|(m[146]&m[332]&m[874]));
    m[619] = (((~m[146]&~m[348]&~m[875])|(m[146]&m[348]&~m[875]))&BiasedRNG[842])|(((m[146]&~m[348]&~m[875])|(~m[146]&m[348]&m[875]))&~BiasedRNG[842])|((~m[146]&~m[348]&m[875])|(m[146]&~m[348]&m[875])|(m[146]&m[348]&m[875]));
    m[620] = (((~m[147]&~m[364]&~m[876])|(m[147]&m[364]&~m[876]))&BiasedRNG[843])|(((m[147]&~m[364]&~m[876])|(~m[147]&m[364]&m[876]))&~BiasedRNG[843])|((~m[147]&~m[364]&m[876])|(m[147]&~m[364]&m[876])|(m[147]&m[364]&m[876]));
    m[621] = (((~m[147]&~m[380]&~m[877])|(m[147]&m[380]&~m[877]))&BiasedRNG[844])|(((m[147]&~m[380]&~m[877])|(~m[147]&m[380]&m[877]))&~BiasedRNG[844])|((~m[147]&~m[380]&m[877])|(m[147]&~m[380]&m[877])|(m[147]&m[380]&m[877]));
    m[622] = (((~m[147]&~m[396]&~m[878])|(m[147]&m[396]&~m[878]))&BiasedRNG[845])|(((m[147]&~m[396]&~m[878])|(~m[147]&m[396]&m[878]))&~BiasedRNG[845])|((~m[147]&~m[396]&m[878])|(m[147]&~m[396]&m[878])|(m[147]&m[396]&m[878]));
    m[623] = (((~m[147]&~m[412]&~m[879])|(m[147]&m[412]&~m[879]))&BiasedRNG[846])|(((m[147]&~m[412]&~m[879])|(~m[147]&m[412]&m[879]))&~BiasedRNG[846])|((~m[147]&~m[412]&m[879])|(m[147]&~m[412]&m[879])|(m[147]&m[412]&m[879]));
    m[624] = (((~m[148]&~m[173]&~m[880])|(m[148]&m[173]&~m[880]))&BiasedRNG[847])|(((m[148]&~m[173]&~m[880])|(~m[148]&m[173]&m[880]))&~BiasedRNG[847])|((~m[148]&~m[173]&m[880])|(m[148]&~m[173]&m[880])|(m[148]&m[173]&m[880]));
    m[625] = (((~m[148]&~m[189]&~m[881])|(m[148]&m[189]&~m[881]))&BiasedRNG[848])|(((m[148]&~m[189]&~m[881])|(~m[148]&m[189]&m[881]))&~BiasedRNG[848])|((~m[148]&~m[189]&m[881])|(m[148]&~m[189]&m[881])|(m[148]&m[189]&m[881]));
    m[626] = (((~m[148]&~m[205]&~m[882])|(m[148]&m[205]&~m[882]))&BiasedRNG[849])|(((m[148]&~m[205]&~m[882])|(~m[148]&m[205]&m[882]))&~BiasedRNG[849])|((~m[148]&~m[205]&m[882])|(m[148]&~m[205]&m[882])|(m[148]&m[205]&m[882]));
    m[627] = (((~m[148]&~m[221]&~m[883])|(m[148]&m[221]&~m[883]))&BiasedRNG[850])|(((m[148]&~m[221]&~m[883])|(~m[148]&m[221]&m[883]))&~BiasedRNG[850])|((~m[148]&~m[221]&m[883])|(m[148]&~m[221]&m[883])|(m[148]&m[221]&m[883]));
    m[628] = (((~m[149]&~m[237]&~m[884])|(m[149]&m[237]&~m[884]))&BiasedRNG[851])|(((m[149]&~m[237]&~m[884])|(~m[149]&m[237]&m[884]))&~BiasedRNG[851])|((~m[149]&~m[237]&m[884])|(m[149]&~m[237]&m[884])|(m[149]&m[237]&m[884]));
    m[629] = (((~m[149]&~m[253]&~m[885])|(m[149]&m[253]&~m[885]))&BiasedRNG[852])|(((m[149]&~m[253]&~m[885])|(~m[149]&m[253]&m[885]))&~BiasedRNG[852])|((~m[149]&~m[253]&m[885])|(m[149]&~m[253]&m[885])|(m[149]&m[253]&m[885]));
    m[630] = (((~m[149]&~m[269]&~m[886])|(m[149]&m[269]&~m[886]))&BiasedRNG[853])|(((m[149]&~m[269]&~m[886])|(~m[149]&m[269]&m[886]))&~BiasedRNG[853])|((~m[149]&~m[269]&m[886])|(m[149]&~m[269]&m[886])|(m[149]&m[269]&m[886]));
    m[631] = (((~m[149]&~m[285]&~m[887])|(m[149]&m[285]&~m[887]))&BiasedRNG[854])|(((m[149]&~m[285]&~m[887])|(~m[149]&m[285]&m[887]))&~BiasedRNG[854])|((~m[149]&~m[285]&m[887])|(m[149]&~m[285]&m[887])|(m[149]&m[285]&m[887]));
    m[632] = (((~m[150]&~m[301]&~m[888])|(m[150]&m[301]&~m[888]))&BiasedRNG[855])|(((m[150]&~m[301]&~m[888])|(~m[150]&m[301]&m[888]))&~BiasedRNG[855])|((~m[150]&~m[301]&m[888])|(m[150]&~m[301]&m[888])|(m[150]&m[301]&m[888]));
    m[633] = (((~m[150]&~m[317]&~m[889])|(m[150]&m[317]&~m[889]))&BiasedRNG[856])|(((m[150]&~m[317]&~m[889])|(~m[150]&m[317]&m[889]))&~BiasedRNG[856])|((~m[150]&~m[317]&m[889])|(m[150]&~m[317]&m[889])|(m[150]&m[317]&m[889]));
    m[634] = (((~m[150]&~m[333]&~m[890])|(m[150]&m[333]&~m[890]))&BiasedRNG[857])|(((m[150]&~m[333]&~m[890])|(~m[150]&m[333]&m[890]))&~BiasedRNG[857])|((~m[150]&~m[333]&m[890])|(m[150]&~m[333]&m[890])|(m[150]&m[333]&m[890]));
    m[635] = (((~m[150]&~m[349]&~m[891])|(m[150]&m[349]&~m[891]))&BiasedRNG[858])|(((m[150]&~m[349]&~m[891])|(~m[150]&m[349]&m[891]))&~BiasedRNG[858])|((~m[150]&~m[349]&m[891])|(m[150]&~m[349]&m[891])|(m[150]&m[349]&m[891]));
    m[636] = (((~m[151]&~m[365]&~m[892])|(m[151]&m[365]&~m[892]))&BiasedRNG[859])|(((m[151]&~m[365]&~m[892])|(~m[151]&m[365]&m[892]))&~BiasedRNG[859])|((~m[151]&~m[365]&m[892])|(m[151]&~m[365]&m[892])|(m[151]&m[365]&m[892]));
    m[637] = (((~m[151]&~m[381]&~m[893])|(m[151]&m[381]&~m[893]))&BiasedRNG[860])|(((m[151]&~m[381]&~m[893])|(~m[151]&m[381]&m[893]))&~BiasedRNG[860])|((~m[151]&~m[381]&m[893])|(m[151]&~m[381]&m[893])|(m[151]&m[381]&m[893]));
    m[638] = (((~m[151]&~m[397]&~m[894])|(m[151]&m[397]&~m[894]))&BiasedRNG[861])|(((m[151]&~m[397]&~m[894])|(~m[151]&m[397]&m[894]))&~BiasedRNG[861])|((~m[151]&~m[397]&m[894])|(m[151]&~m[397]&m[894])|(m[151]&m[397]&m[894]));
    m[639] = (((~m[151]&~m[413]&~m[895])|(m[151]&m[413]&~m[895]))&BiasedRNG[862])|(((m[151]&~m[413]&~m[895])|(~m[151]&m[413]&m[895]))&~BiasedRNG[862])|((~m[151]&~m[413]&m[895])|(m[151]&~m[413]&m[895])|(m[151]&m[413]&m[895]));
    m[640] = (((~m[152]&~m[174]&~m[896])|(m[152]&m[174]&~m[896]))&BiasedRNG[863])|(((m[152]&~m[174]&~m[896])|(~m[152]&m[174]&m[896]))&~BiasedRNG[863])|((~m[152]&~m[174]&m[896])|(m[152]&~m[174]&m[896])|(m[152]&m[174]&m[896]));
    m[641] = (((~m[152]&~m[190]&~m[897])|(m[152]&m[190]&~m[897]))&BiasedRNG[864])|(((m[152]&~m[190]&~m[897])|(~m[152]&m[190]&m[897]))&~BiasedRNG[864])|((~m[152]&~m[190]&m[897])|(m[152]&~m[190]&m[897])|(m[152]&m[190]&m[897]));
    m[642] = (((~m[152]&~m[206]&~m[898])|(m[152]&m[206]&~m[898]))&BiasedRNG[865])|(((m[152]&~m[206]&~m[898])|(~m[152]&m[206]&m[898]))&~BiasedRNG[865])|((~m[152]&~m[206]&m[898])|(m[152]&~m[206]&m[898])|(m[152]&m[206]&m[898]));
    m[643] = (((~m[152]&~m[222]&~m[899])|(m[152]&m[222]&~m[899]))&BiasedRNG[866])|(((m[152]&~m[222]&~m[899])|(~m[152]&m[222]&m[899]))&~BiasedRNG[866])|((~m[152]&~m[222]&m[899])|(m[152]&~m[222]&m[899])|(m[152]&m[222]&m[899]));
    m[644] = (((~m[153]&~m[238]&~m[900])|(m[153]&m[238]&~m[900]))&BiasedRNG[867])|(((m[153]&~m[238]&~m[900])|(~m[153]&m[238]&m[900]))&~BiasedRNG[867])|((~m[153]&~m[238]&m[900])|(m[153]&~m[238]&m[900])|(m[153]&m[238]&m[900]));
    m[645] = (((~m[153]&~m[254]&~m[901])|(m[153]&m[254]&~m[901]))&BiasedRNG[868])|(((m[153]&~m[254]&~m[901])|(~m[153]&m[254]&m[901]))&~BiasedRNG[868])|((~m[153]&~m[254]&m[901])|(m[153]&~m[254]&m[901])|(m[153]&m[254]&m[901]));
    m[646] = (((~m[153]&~m[270]&~m[902])|(m[153]&m[270]&~m[902]))&BiasedRNG[869])|(((m[153]&~m[270]&~m[902])|(~m[153]&m[270]&m[902]))&~BiasedRNG[869])|((~m[153]&~m[270]&m[902])|(m[153]&~m[270]&m[902])|(m[153]&m[270]&m[902]));
    m[647] = (((~m[153]&~m[286]&~m[903])|(m[153]&m[286]&~m[903]))&BiasedRNG[870])|(((m[153]&~m[286]&~m[903])|(~m[153]&m[286]&m[903]))&~BiasedRNG[870])|((~m[153]&~m[286]&m[903])|(m[153]&~m[286]&m[903])|(m[153]&m[286]&m[903]));
    m[648] = (((~m[154]&~m[302]&~m[904])|(m[154]&m[302]&~m[904]))&BiasedRNG[871])|(((m[154]&~m[302]&~m[904])|(~m[154]&m[302]&m[904]))&~BiasedRNG[871])|((~m[154]&~m[302]&m[904])|(m[154]&~m[302]&m[904])|(m[154]&m[302]&m[904]));
    m[649] = (((~m[154]&~m[318]&~m[905])|(m[154]&m[318]&~m[905]))&BiasedRNG[872])|(((m[154]&~m[318]&~m[905])|(~m[154]&m[318]&m[905]))&~BiasedRNG[872])|((~m[154]&~m[318]&m[905])|(m[154]&~m[318]&m[905])|(m[154]&m[318]&m[905]));
    m[650] = (((~m[154]&~m[334]&~m[906])|(m[154]&m[334]&~m[906]))&BiasedRNG[873])|(((m[154]&~m[334]&~m[906])|(~m[154]&m[334]&m[906]))&~BiasedRNG[873])|((~m[154]&~m[334]&m[906])|(m[154]&~m[334]&m[906])|(m[154]&m[334]&m[906]));
    m[651] = (((~m[154]&~m[350]&~m[907])|(m[154]&m[350]&~m[907]))&BiasedRNG[874])|(((m[154]&~m[350]&~m[907])|(~m[154]&m[350]&m[907]))&~BiasedRNG[874])|((~m[154]&~m[350]&m[907])|(m[154]&~m[350]&m[907])|(m[154]&m[350]&m[907]));
    m[652] = (((~m[155]&~m[366]&~m[908])|(m[155]&m[366]&~m[908]))&BiasedRNG[875])|(((m[155]&~m[366]&~m[908])|(~m[155]&m[366]&m[908]))&~BiasedRNG[875])|((~m[155]&~m[366]&m[908])|(m[155]&~m[366]&m[908])|(m[155]&m[366]&m[908]));
    m[653] = (((~m[155]&~m[382]&~m[909])|(m[155]&m[382]&~m[909]))&BiasedRNG[876])|(((m[155]&~m[382]&~m[909])|(~m[155]&m[382]&m[909]))&~BiasedRNG[876])|((~m[155]&~m[382]&m[909])|(m[155]&~m[382]&m[909])|(m[155]&m[382]&m[909]));
    m[654] = (((~m[155]&~m[398]&~m[910])|(m[155]&m[398]&~m[910]))&BiasedRNG[877])|(((m[155]&~m[398]&~m[910])|(~m[155]&m[398]&m[910]))&~BiasedRNG[877])|((~m[155]&~m[398]&m[910])|(m[155]&~m[398]&m[910])|(m[155]&m[398]&m[910]));
    m[655] = (((~m[155]&~m[414]&~m[911])|(m[155]&m[414]&~m[911]))&BiasedRNG[878])|(((m[155]&~m[414]&~m[911])|(~m[155]&m[414]&m[911]))&~BiasedRNG[878])|((~m[155]&~m[414]&m[911])|(m[155]&~m[414]&m[911])|(m[155]&m[414]&m[911]));
    m[656] = (((~m[156]&~m[175]&~m[912])|(m[156]&m[175]&~m[912]))&BiasedRNG[879])|(((m[156]&~m[175]&~m[912])|(~m[156]&m[175]&m[912]))&~BiasedRNG[879])|((~m[156]&~m[175]&m[912])|(m[156]&~m[175]&m[912])|(m[156]&m[175]&m[912]));
    m[657] = (((~m[156]&~m[191]&~m[913])|(m[156]&m[191]&~m[913]))&BiasedRNG[880])|(((m[156]&~m[191]&~m[913])|(~m[156]&m[191]&m[913]))&~BiasedRNG[880])|((~m[156]&~m[191]&m[913])|(m[156]&~m[191]&m[913])|(m[156]&m[191]&m[913]));
    m[658] = (((~m[156]&~m[207]&~m[914])|(m[156]&m[207]&~m[914]))&BiasedRNG[881])|(((m[156]&~m[207]&~m[914])|(~m[156]&m[207]&m[914]))&~BiasedRNG[881])|((~m[156]&~m[207]&m[914])|(m[156]&~m[207]&m[914])|(m[156]&m[207]&m[914]));
    m[659] = (((~m[156]&~m[223]&~m[915])|(m[156]&m[223]&~m[915]))&BiasedRNG[882])|(((m[156]&~m[223]&~m[915])|(~m[156]&m[223]&m[915]))&~BiasedRNG[882])|((~m[156]&~m[223]&m[915])|(m[156]&~m[223]&m[915])|(m[156]&m[223]&m[915]));
    m[660] = (((~m[157]&~m[239]&~m[916])|(m[157]&m[239]&~m[916]))&BiasedRNG[883])|(((m[157]&~m[239]&~m[916])|(~m[157]&m[239]&m[916]))&~BiasedRNG[883])|((~m[157]&~m[239]&m[916])|(m[157]&~m[239]&m[916])|(m[157]&m[239]&m[916]));
    m[661] = (((~m[157]&~m[255]&~m[917])|(m[157]&m[255]&~m[917]))&BiasedRNG[884])|(((m[157]&~m[255]&~m[917])|(~m[157]&m[255]&m[917]))&~BiasedRNG[884])|((~m[157]&~m[255]&m[917])|(m[157]&~m[255]&m[917])|(m[157]&m[255]&m[917]));
    m[662] = (((~m[157]&~m[271]&~m[918])|(m[157]&m[271]&~m[918]))&BiasedRNG[885])|(((m[157]&~m[271]&~m[918])|(~m[157]&m[271]&m[918]))&~BiasedRNG[885])|((~m[157]&~m[271]&m[918])|(m[157]&~m[271]&m[918])|(m[157]&m[271]&m[918]));
    m[663] = (((~m[157]&~m[287]&~m[919])|(m[157]&m[287]&~m[919]))&BiasedRNG[886])|(((m[157]&~m[287]&~m[919])|(~m[157]&m[287]&m[919]))&~BiasedRNG[886])|((~m[157]&~m[287]&m[919])|(m[157]&~m[287]&m[919])|(m[157]&m[287]&m[919]));
    m[664] = (((~m[158]&~m[303]&~m[920])|(m[158]&m[303]&~m[920]))&BiasedRNG[887])|(((m[158]&~m[303]&~m[920])|(~m[158]&m[303]&m[920]))&~BiasedRNG[887])|((~m[158]&~m[303]&m[920])|(m[158]&~m[303]&m[920])|(m[158]&m[303]&m[920]));
    m[665] = (((~m[158]&~m[319]&~m[921])|(m[158]&m[319]&~m[921]))&BiasedRNG[888])|(((m[158]&~m[319]&~m[921])|(~m[158]&m[319]&m[921]))&~BiasedRNG[888])|((~m[158]&~m[319]&m[921])|(m[158]&~m[319]&m[921])|(m[158]&m[319]&m[921]));
    m[666] = (((~m[158]&~m[335]&~m[922])|(m[158]&m[335]&~m[922]))&BiasedRNG[889])|(((m[158]&~m[335]&~m[922])|(~m[158]&m[335]&m[922]))&~BiasedRNG[889])|((~m[158]&~m[335]&m[922])|(m[158]&~m[335]&m[922])|(m[158]&m[335]&m[922]));
    m[667] = (((~m[158]&~m[351]&~m[923])|(m[158]&m[351]&~m[923]))&BiasedRNG[890])|(((m[158]&~m[351]&~m[923])|(~m[158]&m[351]&m[923]))&~BiasedRNG[890])|((~m[158]&~m[351]&m[923])|(m[158]&~m[351]&m[923])|(m[158]&m[351]&m[923]));
    m[668] = (((~m[159]&~m[367]&~m[924])|(m[159]&m[367]&~m[924]))&BiasedRNG[891])|(((m[159]&~m[367]&~m[924])|(~m[159]&m[367]&m[924]))&~BiasedRNG[891])|((~m[159]&~m[367]&m[924])|(m[159]&~m[367]&m[924])|(m[159]&m[367]&m[924]));
    m[669] = (((~m[159]&~m[383]&~m[925])|(m[159]&m[383]&~m[925]))&BiasedRNG[892])|(((m[159]&~m[383]&~m[925])|(~m[159]&m[383]&m[925]))&~BiasedRNG[892])|((~m[159]&~m[383]&m[925])|(m[159]&~m[383]&m[925])|(m[159]&m[383]&m[925]));
    m[670] = (((~m[159]&~m[399]&~m[926])|(m[159]&m[399]&~m[926]))&BiasedRNG[893])|(((m[159]&~m[399]&~m[926])|(~m[159]&m[399]&m[926]))&~BiasedRNG[893])|((~m[159]&~m[399]&m[926])|(m[159]&~m[399]&m[926])|(m[159]&m[399]&m[926]));
    m[671] = (((~m[159]&~m[415]&~m[927])|(m[159]&m[415]&~m[927]))&BiasedRNG[894])|(((m[159]&~m[415]&~m[927])|(~m[159]&m[415]&m[927]))&~BiasedRNG[894])|((~m[159]&~m[415]&m[927])|(m[159]&~m[415]&m[927])|(m[159]&m[415]&m[927]));
    m[929] = (((m[688]&~m[928]&~m[930]&~m[931]&~m[932])|(~m[688]&~m[928]&~m[930]&m[931]&~m[932])|(m[688]&m[928]&~m[930]&m[931]&~m[932])|(m[688]&~m[928]&m[930]&m[931]&~m[932])|(~m[688]&m[928]&~m[930]&~m[931]&m[932])|(~m[688]&~m[928]&m[930]&~m[931]&m[932])|(m[688]&m[928]&m[930]&~m[931]&m[932])|(~m[688]&m[928]&m[930]&m[931]&m[932]))&UnbiasedRNG[496])|((m[688]&~m[928]&~m[930]&m[931]&~m[932])|(~m[688]&~m[928]&~m[930]&~m[931]&m[932])|(m[688]&~m[928]&~m[930]&~m[931]&m[932])|(m[688]&m[928]&~m[930]&~m[931]&m[932])|(m[688]&~m[928]&m[930]&~m[931]&m[932])|(~m[688]&~m[928]&~m[930]&m[931]&m[932])|(m[688]&~m[928]&~m[930]&m[931]&m[932])|(~m[688]&m[928]&~m[930]&m[931]&m[932])|(m[688]&m[928]&~m[930]&m[931]&m[932])|(~m[688]&~m[928]&m[930]&m[931]&m[932])|(m[688]&~m[928]&m[930]&m[931]&m[932])|(m[688]&m[928]&m[930]&m[931]&m[932]));
    m[934] = (((m[689]&~m[933]&~m[935]&~m[936]&~m[937])|(~m[689]&~m[933]&~m[935]&m[936]&~m[937])|(m[689]&m[933]&~m[935]&m[936]&~m[937])|(m[689]&~m[933]&m[935]&m[936]&~m[937])|(~m[689]&m[933]&~m[935]&~m[936]&m[937])|(~m[689]&~m[933]&m[935]&~m[936]&m[937])|(m[689]&m[933]&m[935]&~m[936]&m[937])|(~m[689]&m[933]&m[935]&m[936]&m[937]))&UnbiasedRNG[497])|((m[689]&~m[933]&~m[935]&m[936]&~m[937])|(~m[689]&~m[933]&~m[935]&~m[936]&m[937])|(m[689]&~m[933]&~m[935]&~m[936]&m[937])|(m[689]&m[933]&~m[935]&~m[936]&m[937])|(m[689]&~m[933]&m[935]&~m[936]&m[937])|(~m[689]&~m[933]&~m[935]&m[936]&m[937])|(m[689]&~m[933]&~m[935]&m[936]&m[937])|(~m[689]&m[933]&~m[935]&m[936]&m[937])|(m[689]&m[933]&~m[935]&m[936]&m[937])|(~m[689]&~m[933]&m[935]&m[936]&m[937])|(m[689]&~m[933]&m[935]&m[936]&m[937])|(m[689]&m[933]&m[935]&m[936]&m[937]));
    m[939] = (((m[704]&~m[938]&~m[940]&~m[941]&~m[942])|(~m[704]&~m[938]&~m[940]&m[941]&~m[942])|(m[704]&m[938]&~m[940]&m[941]&~m[942])|(m[704]&~m[938]&m[940]&m[941]&~m[942])|(~m[704]&m[938]&~m[940]&~m[941]&m[942])|(~m[704]&~m[938]&m[940]&~m[941]&m[942])|(m[704]&m[938]&m[940]&~m[941]&m[942])|(~m[704]&m[938]&m[940]&m[941]&m[942]))&UnbiasedRNG[498])|((m[704]&~m[938]&~m[940]&m[941]&~m[942])|(~m[704]&~m[938]&~m[940]&~m[941]&m[942])|(m[704]&~m[938]&~m[940]&~m[941]&m[942])|(m[704]&m[938]&~m[940]&~m[941]&m[942])|(m[704]&~m[938]&m[940]&~m[941]&m[942])|(~m[704]&~m[938]&~m[940]&m[941]&m[942])|(m[704]&~m[938]&~m[940]&m[941]&m[942])|(~m[704]&m[938]&~m[940]&m[941]&m[942])|(m[704]&m[938]&~m[940]&m[941]&m[942])|(~m[704]&~m[938]&m[940]&m[941]&m[942])|(m[704]&~m[938]&m[940]&m[941]&m[942])|(m[704]&m[938]&m[940]&m[941]&m[942]));
    m[944] = (((m[690]&~m[943]&~m[945]&~m[946]&~m[947])|(~m[690]&~m[943]&~m[945]&m[946]&~m[947])|(m[690]&m[943]&~m[945]&m[946]&~m[947])|(m[690]&~m[943]&m[945]&m[946]&~m[947])|(~m[690]&m[943]&~m[945]&~m[946]&m[947])|(~m[690]&~m[943]&m[945]&~m[946]&m[947])|(m[690]&m[943]&m[945]&~m[946]&m[947])|(~m[690]&m[943]&m[945]&m[946]&m[947]))&UnbiasedRNG[499])|((m[690]&~m[943]&~m[945]&m[946]&~m[947])|(~m[690]&~m[943]&~m[945]&~m[946]&m[947])|(m[690]&~m[943]&~m[945]&~m[946]&m[947])|(m[690]&m[943]&~m[945]&~m[946]&m[947])|(m[690]&~m[943]&m[945]&~m[946]&m[947])|(~m[690]&~m[943]&~m[945]&m[946]&m[947])|(m[690]&~m[943]&~m[945]&m[946]&m[947])|(~m[690]&m[943]&~m[945]&m[946]&m[947])|(m[690]&m[943]&~m[945]&m[946]&m[947])|(~m[690]&~m[943]&m[945]&m[946]&m[947])|(m[690]&~m[943]&m[945]&m[946]&m[947])|(m[690]&m[943]&m[945]&m[946]&m[947]));
    m[949] = (((m[705]&~m[948]&~m[950]&~m[951]&~m[952])|(~m[705]&~m[948]&~m[950]&m[951]&~m[952])|(m[705]&m[948]&~m[950]&m[951]&~m[952])|(m[705]&~m[948]&m[950]&m[951]&~m[952])|(~m[705]&m[948]&~m[950]&~m[951]&m[952])|(~m[705]&~m[948]&m[950]&~m[951]&m[952])|(m[705]&m[948]&m[950]&~m[951]&m[952])|(~m[705]&m[948]&m[950]&m[951]&m[952]))&UnbiasedRNG[500])|((m[705]&~m[948]&~m[950]&m[951]&~m[952])|(~m[705]&~m[948]&~m[950]&~m[951]&m[952])|(m[705]&~m[948]&~m[950]&~m[951]&m[952])|(m[705]&m[948]&~m[950]&~m[951]&m[952])|(m[705]&~m[948]&m[950]&~m[951]&m[952])|(~m[705]&~m[948]&~m[950]&m[951]&m[952])|(m[705]&~m[948]&~m[950]&m[951]&m[952])|(~m[705]&m[948]&~m[950]&m[951]&m[952])|(m[705]&m[948]&~m[950]&m[951]&m[952])|(~m[705]&~m[948]&m[950]&m[951]&m[952])|(m[705]&~m[948]&m[950]&m[951]&m[952])|(m[705]&m[948]&m[950]&m[951]&m[952]));
    m[954] = (((m[720]&~m[953]&~m[955]&~m[956]&~m[957])|(~m[720]&~m[953]&~m[955]&m[956]&~m[957])|(m[720]&m[953]&~m[955]&m[956]&~m[957])|(m[720]&~m[953]&m[955]&m[956]&~m[957])|(~m[720]&m[953]&~m[955]&~m[956]&m[957])|(~m[720]&~m[953]&m[955]&~m[956]&m[957])|(m[720]&m[953]&m[955]&~m[956]&m[957])|(~m[720]&m[953]&m[955]&m[956]&m[957]))&UnbiasedRNG[501])|((m[720]&~m[953]&~m[955]&m[956]&~m[957])|(~m[720]&~m[953]&~m[955]&~m[956]&m[957])|(m[720]&~m[953]&~m[955]&~m[956]&m[957])|(m[720]&m[953]&~m[955]&~m[956]&m[957])|(m[720]&~m[953]&m[955]&~m[956]&m[957])|(~m[720]&~m[953]&~m[955]&m[956]&m[957])|(m[720]&~m[953]&~m[955]&m[956]&m[957])|(~m[720]&m[953]&~m[955]&m[956]&m[957])|(m[720]&m[953]&~m[955]&m[956]&m[957])|(~m[720]&~m[953]&m[955]&m[956]&m[957])|(m[720]&~m[953]&m[955]&m[956]&m[957])|(m[720]&m[953]&m[955]&m[956]&m[957]));
    m[959] = (((m[691]&~m[958]&~m[960]&~m[961]&~m[962])|(~m[691]&~m[958]&~m[960]&m[961]&~m[962])|(m[691]&m[958]&~m[960]&m[961]&~m[962])|(m[691]&~m[958]&m[960]&m[961]&~m[962])|(~m[691]&m[958]&~m[960]&~m[961]&m[962])|(~m[691]&~m[958]&m[960]&~m[961]&m[962])|(m[691]&m[958]&m[960]&~m[961]&m[962])|(~m[691]&m[958]&m[960]&m[961]&m[962]))&UnbiasedRNG[502])|((m[691]&~m[958]&~m[960]&m[961]&~m[962])|(~m[691]&~m[958]&~m[960]&~m[961]&m[962])|(m[691]&~m[958]&~m[960]&~m[961]&m[962])|(m[691]&m[958]&~m[960]&~m[961]&m[962])|(m[691]&~m[958]&m[960]&~m[961]&m[962])|(~m[691]&~m[958]&~m[960]&m[961]&m[962])|(m[691]&~m[958]&~m[960]&m[961]&m[962])|(~m[691]&m[958]&~m[960]&m[961]&m[962])|(m[691]&m[958]&~m[960]&m[961]&m[962])|(~m[691]&~m[958]&m[960]&m[961]&m[962])|(m[691]&~m[958]&m[960]&m[961]&m[962])|(m[691]&m[958]&m[960]&m[961]&m[962]));
    m[964] = (((m[706]&~m[963]&~m[965]&~m[966]&~m[967])|(~m[706]&~m[963]&~m[965]&m[966]&~m[967])|(m[706]&m[963]&~m[965]&m[966]&~m[967])|(m[706]&~m[963]&m[965]&m[966]&~m[967])|(~m[706]&m[963]&~m[965]&~m[966]&m[967])|(~m[706]&~m[963]&m[965]&~m[966]&m[967])|(m[706]&m[963]&m[965]&~m[966]&m[967])|(~m[706]&m[963]&m[965]&m[966]&m[967]))&UnbiasedRNG[503])|((m[706]&~m[963]&~m[965]&m[966]&~m[967])|(~m[706]&~m[963]&~m[965]&~m[966]&m[967])|(m[706]&~m[963]&~m[965]&~m[966]&m[967])|(m[706]&m[963]&~m[965]&~m[966]&m[967])|(m[706]&~m[963]&m[965]&~m[966]&m[967])|(~m[706]&~m[963]&~m[965]&m[966]&m[967])|(m[706]&~m[963]&~m[965]&m[966]&m[967])|(~m[706]&m[963]&~m[965]&m[966]&m[967])|(m[706]&m[963]&~m[965]&m[966]&m[967])|(~m[706]&~m[963]&m[965]&m[966]&m[967])|(m[706]&~m[963]&m[965]&m[966]&m[967])|(m[706]&m[963]&m[965]&m[966]&m[967]));
    m[969] = (((m[721]&~m[968]&~m[970]&~m[971]&~m[972])|(~m[721]&~m[968]&~m[970]&m[971]&~m[972])|(m[721]&m[968]&~m[970]&m[971]&~m[972])|(m[721]&~m[968]&m[970]&m[971]&~m[972])|(~m[721]&m[968]&~m[970]&~m[971]&m[972])|(~m[721]&~m[968]&m[970]&~m[971]&m[972])|(m[721]&m[968]&m[970]&~m[971]&m[972])|(~m[721]&m[968]&m[970]&m[971]&m[972]))&UnbiasedRNG[504])|((m[721]&~m[968]&~m[970]&m[971]&~m[972])|(~m[721]&~m[968]&~m[970]&~m[971]&m[972])|(m[721]&~m[968]&~m[970]&~m[971]&m[972])|(m[721]&m[968]&~m[970]&~m[971]&m[972])|(m[721]&~m[968]&m[970]&~m[971]&m[972])|(~m[721]&~m[968]&~m[970]&m[971]&m[972])|(m[721]&~m[968]&~m[970]&m[971]&m[972])|(~m[721]&m[968]&~m[970]&m[971]&m[972])|(m[721]&m[968]&~m[970]&m[971]&m[972])|(~m[721]&~m[968]&m[970]&m[971]&m[972])|(m[721]&~m[968]&m[970]&m[971]&m[972])|(m[721]&m[968]&m[970]&m[971]&m[972]));
    m[974] = (((m[736]&~m[973]&~m[975]&~m[976]&~m[977])|(~m[736]&~m[973]&~m[975]&m[976]&~m[977])|(m[736]&m[973]&~m[975]&m[976]&~m[977])|(m[736]&~m[973]&m[975]&m[976]&~m[977])|(~m[736]&m[973]&~m[975]&~m[976]&m[977])|(~m[736]&~m[973]&m[975]&~m[976]&m[977])|(m[736]&m[973]&m[975]&~m[976]&m[977])|(~m[736]&m[973]&m[975]&m[976]&m[977]))&UnbiasedRNG[505])|((m[736]&~m[973]&~m[975]&m[976]&~m[977])|(~m[736]&~m[973]&~m[975]&~m[976]&m[977])|(m[736]&~m[973]&~m[975]&~m[976]&m[977])|(m[736]&m[973]&~m[975]&~m[976]&m[977])|(m[736]&~m[973]&m[975]&~m[976]&m[977])|(~m[736]&~m[973]&~m[975]&m[976]&m[977])|(m[736]&~m[973]&~m[975]&m[976]&m[977])|(~m[736]&m[973]&~m[975]&m[976]&m[977])|(m[736]&m[973]&~m[975]&m[976]&m[977])|(~m[736]&~m[973]&m[975]&m[976]&m[977])|(m[736]&~m[973]&m[975]&m[976]&m[977])|(m[736]&m[973]&m[975]&m[976]&m[977]));
    m[979] = (((m[692]&~m[978]&~m[980]&~m[981]&~m[982])|(~m[692]&~m[978]&~m[980]&m[981]&~m[982])|(m[692]&m[978]&~m[980]&m[981]&~m[982])|(m[692]&~m[978]&m[980]&m[981]&~m[982])|(~m[692]&m[978]&~m[980]&~m[981]&m[982])|(~m[692]&~m[978]&m[980]&~m[981]&m[982])|(m[692]&m[978]&m[980]&~m[981]&m[982])|(~m[692]&m[978]&m[980]&m[981]&m[982]))&UnbiasedRNG[506])|((m[692]&~m[978]&~m[980]&m[981]&~m[982])|(~m[692]&~m[978]&~m[980]&~m[981]&m[982])|(m[692]&~m[978]&~m[980]&~m[981]&m[982])|(m[692]&m[978]&~m[980]&~m[981]&m[982])|(m[692]&~m[978]&m[980]&~m[981]&m[982])|(~m[692]&~m[978]&~m[980]&m[981]&m[982])|(m[692]&~m[978]&~m[980]&m[981]&m[982])|(~m[692]&m[978]&~m[980]&m[981]&m[982])|(m[692]&m[978]&~m[980]&m[981]&m[982])|(~m[692]&~m[978]&m[980]&m[981]&m[982])|(m[692]&~m[978]&m[980]&m[981]&m[982])|(m[692]&m[978]&m[980]&m[981]&m[982]));
    m[984] = (((m[707]&~m[983]&~m[985]&~m[986]&~m[987])|(~m[707]&~m[983]&~m[985]&m[986]&~m[987])|(m[707]&m[983]&~m[985]&m[986]&~m[987])|(m[707]&~m[983]&m[985]&m[986]&~m[987])|(~m[707]&m[983]&~m[985]&~m[986]&m[987])|(~m[707]&~m[983]&m[985]&~m[986]&m[987])|(m[707]&m[983]&m[985]&~m[986]&m[987])|(~m[707]&m[983]&m[985]&m[986]&m[987]))&UnbiasedRNG[507])|((m[707]&~m[983]&~m[985]&m[986]&~m[987])|(~m[707]&~m[983]&~m[985]&~m[986]&m[987])|(m[707]&~m[983]&~m[985]&~m[986]&m[987])|(m[707]&m[983]&~m[985]&~m[986]&m[987])|(m[707]&~m[983]&m[985]&~m[986]&m[987])|(~m[707]&~m[983]&~m[985]&m[986]&m[987])|(m[707]&~m[983]&~m[985]&m[986]&m[987])|(~m[707]&m[983]&~m[985]&m[986]&m[987])|(m[707]&m[983]&~m[985]&m[986]&m[987])|(~m[707]&~m[983]&m[985]&m[986]&m[987])|(m[707]&~m[983]&m[985]&m[986]&m[987])|(m[707]&m[983]&m[985]&m[986]&m[987]));
    m[989] = (((m[722]&~m[988]&~m[990]&~m[991]&~m[992])|(~m[722]&~m[988]&~m[990]&m[991]&~m[992])|(m[722]&m[988]&~m[990]&m[991]&~m[992])|(m[722]&~m[988]&m[990]&m[991]&~m[992])|(~m[722]&m[988]&~m[990]&~m[991]&m[992])|(~m[722]&~m[988]&m[990]&~m[991]&m[992])|(m[722]&m[988]&m[990]&~m[991]&m[992])|(~m[722]&m[988]&m[990]&m[991]&m[992]))&UnbiasedRNG[508])|((m[722]&~m[988]&~m[990]&m[991]&~m[992])|(~m[722]&~m[988]&~m[990]&~m[991]&m[992])|(m[722]&~m[988]&~m[990]&~m[991]&m[992])|(m[722]&m[988]&~m[990]&~m[991]&m[992])|(m[722]&~m[988]&m[990]&~m[991]&m[992])|(~m[722]&~m[988]&~m[990]&m[991]&m[992])|(m[722]&~m[988]&~m[990]&m[991]&m[992])|(~m[722]&m[988]&~m[990]&m[991]&m[992])|(m[722]&m[988]&~m[990]&m[991]&m[992])|(~m[722]&~m[988]&m[990]&m[991]&m[992])|(m[722]&~m[988]&m[990]&m[991]&m[992])|(m[722]&m[988]&m[990]&m[991]&m[992]));
    m[994] = (((m[737]&~m[993]&~m[995]&~m[996]&~m[997])|(~m[737]&~m[993]&~m[995]&m[996]&~m[997])|(m[737]&m[993]&~m[995]&m[996]&~m[997])|(m[737]&~m[993]&m[995]&m[996]&~m[997])|(~m[737]&m[993]&~m[995]&~m[996]&m[997])|(~m[737]&~m[993]&m[995]&~m[996]&m[997])|(m[737]&m[993]&m[995]&~m[996]&m[997])|(~m[737]&m[993]&m[995]&m[996]&m[997]))&UnbiasedRNG[509])|((m[737]&~m[993]&~m[995]&m[996]&~m[997])|(~m[737]&~m[993]&~m[995]&~m[996]&m[997])|(m[737]&~m[993]&~m[995]&~m[996]&m[997])|(m[737]&m[993]&~m[995]&~m[996]&m[997])|(m[737]&~m[993]&m[995]&~m[996]&m[997])|(~m[737]&~m[993]&~m[995]&m[996]&m[997])|(m[737]&~m[993]&~m[995]&m[996]&m[997])|(~m[737]&m[993]&~m[995]&m[996]&m[997])|(m[737]&m[993]&~m[995]&m[996]&m[997])|(~m[737]&~m[993]&m[995]&m[996]&m[997])|(m[737]&~m[993]&m[995]&m[996]&m[997])|(m[737]&m[993]&m[995]&m[996]&m[997]));
    m[999] = (((m[752]&~m[998]&~m[1000]&~m[1001]&~m[1002])|(~m[752]&~m[998]&~m[1000]&m[1001]&~m[1002])|(m[752]&m[998]&~m[1000]&m[1001]&~m[1002])|(m[752]&~m[998]&m[1000]&m[1001]&~m[1002])|(~m[752]&m[998]&~m[1000]&~m[1001]&m[1002])|(~m[752]&~m[998]&m[1000]&~m[1001]&m[1002])|(m[752]&m[998]&m[1000]&~m[1001]&m[1002])|(~m[752]&m[998]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[510])|((m[752]&~m[998]&~m[1000]&m[1001]&~m[1002])|(~m[752]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[752]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[752]&m[998]&~m[1000]&~m[1001]&m[1002])|(m[752]&~m[998]&m[1000]&~m[1001]&m[1002])|(~m[752]&~m[998]&~m[1000]&m[1001]&m[1002])|(m[752]&~m[998]&~m[1000]&m[1001]&m[1002])|(~m[752]&m[998]&~m[1000]&m[1001]&m[1002])|(m[752]&m[998]&~m[1000]&m[1001]&m[1002])|(~m[752]&~m[998]&m[1000]&m[1001]&m[1002])|(m[752]&~m[998]&m[1000]&m[1001]&m[1002])|(m[752]&m[998]&m[1000]&m[1001]&m[1002]));
    m[1004] = (((m[693]&~m[1003]&~m[1005]&~m[1006]&~m[1007])|(~m[693]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(m[693]&m[1003]&~m[1005]&m[1006]&~m[1007])|(m[693]&~m[1003]&m[1005]&m[1006]&~m[1007])|(~m[693]&m[1003]&~m[1005]&~m[1006]&m[1007])|(~m[693]&~m[1003]&m[1005]&~m[1006]&m[1007])|(m[693]&m[1003]&m[1005]&~m[1006]&m[1007])|(~m[693]&m[1003]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[511])|((m[693]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(~m[693]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[693]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[693]&m[1003]&~m[1005]&~m[1006]&m[1007])|(m[693]&~m[1003]&m[1005]&~m[1006]&m[1007])|(~m[693]&~m[1003]&~m[1005]&m[1006]&m[1007])|(m[693]&~m[1003]&~m[1005]&m[1006]&m[1007])|(~m[693]&m[1003]&~m[1005]&m[1006]&m[1007])|(m[693]&m[1003]&~m[1005]&m[1006]&m[1007])|(~m[693]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[693]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[693]&m[1003]&m[1005]&m[1006]&m[1007]));
    m[1009] = (((m[708]&~m[1008]&~m[1010]&~m[1011]&~m[1012])|(~m[708]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(m[708]&m[1008]&~m[1010]&m[1011]&~m[1012])|(m[708]&~m[1008]&m[1010]&m[1011]&~m[1012])|(~m[708]&m[1008]&~m[1010]&~m[1011]&m[1012])|(~m[708]&~m[1008]&m[1010]&~m[1011]&m[1012])|(m[708]&m[1008]&m[1010]&~m[1011]&m[1012])|(~m[708]&m[1008]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[512])|((m[708]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(~m[708]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[708]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[708]&m[1008]&~m[1010]&~m[1011]&m[1012])|(m[708]&~m[1008]&m[1010]&~m[1011]&m[1012])|(~m[708]&~m[1008]&~m[1010]&m[1011]&m[1012])|(m[708]&~m[1008]&~m[1010]&m[1011]&m[1012])|(~m[708]&m[1008]&~m[1010]&m[1011]&m[1012])|(m[708]&m[1008]&~m[1010]&m[1011]&m[1012])|(~m[708]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[708]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[708]&m[1008]&m[1010]&m[1011]&m[1012]));
    m[1014] = (((m[723]&~m[1013]&~m[1015]&~m[1016]&~m[1017])|(~m[723]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(m[723]&m[1013]&~m[1015]&m[1016]&~m[1017])|(m[723]&~m[1013]&m[1015]&m[1016]&~m[1017])|(~m[723]&m[1013]&~m[1015]&~m[1016]&m[1017])|(~m[723]&~m[1013]&m[1015]&~m[1016]&m[1017])|(m[723]&m[1013]&m[1015]&~m[1016]&m[1017])|(~m[723]&m[1013]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[513])|((m[723]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(~m[723]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[723]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[723]&m[1013]&~m[1015]&~m[1016]&m[1017])|(m[723]&~m[1013]&m[1015]&~m[1016]&m[1017])|(~m[723]&~m[1013]&~m[1015]&m[1016]&m[1017])|(m[723]&~m[1013]&~m[1015]&m[1016]&m[1017])|(~m[723]&m[1013]&~m[1015]&m[1016]&m[1017])|(m[723]&m[1013]&~m[1015]&m[1016]&m[1017])|(~m[723]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[723]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[723]&m[1013]&m[1015]&m[1016]&m[1017]));
    m[1019] = (((m[738]&~m[1018]&~m[1020]&~m[1021]&~m[1022])|(~m[738]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(m[738]&m[1018]&~m[1020]&m[1021]&~m[1022])|(m[738]&~m[1018]&m[1020]&m[1021]&~m[1022])|(~m[738]&m[1018]&~m[1020]&~m[1021]&m[1022])|(~m[738]&~m[1018]&m[1020]&~m[1021]&m[1022])|(m[738]&m[1018]&m[1020]&~m[1021]&m[1022])|(~m[738]&m[1018]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[514])|((m[738]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(~m[738]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[738]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[738]&m[1018]&~m[1020]&~m[1021]&m[1022])|(m[738]&~m[1018]&m[1020]&~m[1021]&m[1022])|(~m[738]&~m[1018]&~m[1020]&m[1021]&m[1022])|(m[738]&~m[1018]&~m[1020]&m[1021]&m[1022])|(~m[738]&m[1018]&~m[1020]&m[1021]&m[1022])|(m[738]&m[1018]&~m[1020]&m[1021]&m[1022])|(~m[738]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[738]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[738]&m[1018]&m[1020]&m[1021]&m[1022]));
    m[1024] = (((m[753]&~m[1023]&~m[1025]&~m[1026]&~m[1027])|(~m[753]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(m[753]&m[1023]&~m[1025]&m[1026]&~m[1027])|(m[753]&~m[1023]&m[1025]&m[1026]&~m[1027])|(~m[753]&m[1023]&~m[1025]&~m[1026]&m[1027])|(~m[753]&~m[1023]&m[1025]&~m[1026]&m[1027])|(m[753]&m[1023]&m[1025]&~m[1026]&m[1027])|(~m[753]&m[1023]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[515])|((m[753]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(~m[753]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[753]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[753]&m[1023]&~m[1025]&~m[1026]&m[1027])|(m[753]&~m[1023]&m[1025]&~m[1026]&m[1027])|(~m[753]&~m[1023]&~m[1025]&m[1026]&m[1027])|(m[753]&~m[1023]&~m[1025]&m[1026]&m[1027])|(~m[753]&m[1023]&~m[1025]&m[1026]&m[1027])|(m[753]&m[1023]&~m[1025]&m[1026]&m[1027])|(~m[753]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[753]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[753]&m[1023]&m[1025]&m[1026]&m[1027]));
    m[1029] = (((m[768]&~m[1028]&~m[1030]&~m[1031]&~m[1032])|(~m[768]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(m[768]&m[1028]&~m[1030]&m[1031]&~m[1032])|(m[768]&~m[1028]&m[1030]&m[1031]&~m[1032])|(~m[768]&m[1028]&~m[1030]&~m[1031]&m[1032])|(~m[768]&~m[1028]&m[1030]&~m[1031]&m[1032])|(m[768]&m[1028]&m[1030]&~m[1031]&m[1032])|(~m[768]&m[1028]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[516])|((m[768]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(~m[768]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[768]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[768]&m[1028]&~m[1030]&~m[1031]&m[1032])|(m[768]&~m[1028]&m[1030]&~m[1031]&m[1032])|(~m[768]&~m[1028]&~m[1030]&m[1031]&m[1032])|(m[768]&~m[1028]&~m[1030]&m[1031]&m[1032])|(~m[768]&m[1028]&~m[1030]&m[1031]&m[1032])|(m[768]&m[1028]&~m[1030]&m[1031]&m[1032])|(~m[768]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[768]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[768]&m[1028]&m[1030]&m[1031]&m[1032]));
    m[1034] = (((m[694]&~m[1033]&~m[1035]&~m[1036]&~m[1037])|(~m[694]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(m[694]&m[1033]&~m[1035]&m[1036]&~m[1037])|(m[694]&~m[1033]&m[1035]&m[1036]&~m[1037])|(~m[694]&m[1033]&~m[1035]&~m[1036]&m[1037])|(~m[694]&~m[1033]&m[1035]&~m[1036]&m[1037])|(m[694]&m[1033]&m[1035]&~m[1036]&m[1037])|(~m[694]&m[1033]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[517])|((m[694]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(~m[694]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[694]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[694]&m[1033]&~m[1035]&~m[1036]&m[1037])|(m[694]&~m[1033]&m[1035]&~m[1036]&m[1037])|(~m[694]&~m[1033]&~m[1035]&m[1036]&m[1037])|(m[694]&~m[1033]&~m[1035]&m[1036]&m[1037])|(~m[694]&m[1033]&~m[1035]&m[1036]&m[1037])|(m[694]&m[1033]&~m[1035]&m[1036]&m[1037])|(~m[694]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[694]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[694]&m[1033]&m[1035]&m[1036]&m[1037]));
    m[1039] = (((m[709]&~m[1038]&~m[1040]&~m[1041]&~m[1042])|(~m[709]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(m[709]&m[1038]&~m[1040]&m[1041]&~m[1042])|(m[709]&~m[1038]&m[1040]&m[1041]&~m[1042])|(~m[709]&m[1038]&~m[1040]&~m[1041]&m[1042])|(~m[709]&~m[1038]&m[1040]&~m[1041]&m[1042])|(m[709]&m[1038]&m[1040]&~m[1041]&m[1042])|(~m[709]&m[1038]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[518])|((m[709]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(~m[709]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[709]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[709]&m[1038]&~m[1040]&~m[1041]&m[1042])|(m[709]&~m[1038]&m[1040]&~m[1041]&m[1042])|(~m[709]&~m[1038]&~m[1040]&m[1041]&m[1042])|(m[709]&~m[1038]&~m[1040]&m[1041]&m[1042])|(~m[709]&m[1038]&~m[1040]&m[1041]&m[1042])|(m[709]&m[1038]&~m[1040]&m[1041]&m[1042])|(~m[709]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[709]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[709]&m[1038]&m[1040]&m[1041]&m[1042]));
    m[1044] = (((m[724]&~m[1043]&~m[1045]&~m[1046]&~m[1047])|(~m[724]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(m[724]&m[1043]&~m[1045]&m[1046]&~m[1047])|(m[724]&~m[1043]&m[1045]&m[1046]&~m[1047])|(~m[724]&m[1043]&~m[1045]&~m[1046]&m[1047])|(~m[724]&~m[1043]&m[1045]&~m[1046]&m[1047])|(m[724]&m[1043]&m[1045]&~m[1046]&m[1047])|(~m[724]&m[1043]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[519])|((m[724]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(~m[724]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[724]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[724]&m[1043]&~m[1045]&~m[1046]&m[1047])|(m[724]&~m[1043]&m[1045]&~m[1046]&m[1047])|(~m[724]&~m[1043]&~m[1045]&m[1046]&m[1047])|(m[724]&~m[1043]&~m[1045]&m[1046]&m[1047])|(~m[724]&m[1043]&~m[1045]&m[1046]&m[1047])|(m[724]&m[1043]&~m[1045]&m[1046]&m[1047])|(~m[724]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[724]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[724]&m[1043]&m[1045]&m[1046]&m[1047]));
    m[1049] = (((m[739]&~m[1048]&~m[1050]&~m[1051]&~m[1052])|(~m[739]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(m[739]&m[1048]&~m[1050]&m[1051]&~m[1052])|(m[739]&~m[1048]&m[1050]&m[1051]&~m[1052])|(~m[739]&m[1048]&~m[1050]&~m[1051]&m[1052])|(~m[739]&~m[1048]&m[1050]&~m[1051]&m[1052])|(m[739]&m[1048]&m[1050]&~m[1051]&m[1052])|(~m[739]&m[1048]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[520])|((m[739]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(~m[739]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[739]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[739]&m[1048]&~m[1050]&~m[1051]&m[1052])|(m[739]&~m[1048]&m[1050]&~m[1051]&m[1052])|(~m[739]&~m[1048]&~m[1050]&m[1051]&m[1052])|(m[739]&~m[1048]&~m[1050]&m[1051]&m[1052])|(~m[739]&m[1048]&~m[1050]&m[1051]&m[1052])|(m[739]&m[1048]&~m[1050]&m[1051]&m[1052])|(~m[739]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[739]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[739]&m[1048]&m[1050]&m[1051]&m[1052]));
    m[1054] = (((m[754]&~m[1053]&~m[1055]&~m[1056]&~m[1057])|(~m[754]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(m[754]&m[1053]&~m[1055]&m[1056]&~m[1057])|(m[754]&~m[1053]&m[1055]&m[1056]&~m[1057])|(~m[754]&m[1053]&~m[1055]&~m[1056]&m[1057])|(~m[754]&~m[1053]&m[1055]&~m[1056]&m[1057])|(m[754]&m[1053]&m[1055]&~m[1056]&m[1057])|(~m[754]&m[1053]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[521])|((m[754]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(~m[754]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[754]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[754]&m[1053]&~m[1055]&~m[1056]&m[1057])|(m[754]&~m[1053]&m[1055]&~m[1056]&m[1057])|(~m[754]&~m[1053]&~m[1055]&m[1056]&m[1057])|(m[754]&~m[1053]&~m[1055]&m[1056]&m[1057])|(~m[754]&m[1053]&~m[1055]&m[1056]&m[1057])|(m[754]&m[1053]&~m[1055]&m[1056]&m[1057])|(~m[754]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[754]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[754]&m[1053]&m[1055]&m[1056]&m[1057]));
    m[1059] = (((m[769]&~m[1058]&~m[1060]&~m[1061]&~m[1062])|(~m[769]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(m[769]&m[1058]&~m[1060]&m[1061]&~m[1062])|(m[769]&~m[1058]&m[1060]&m[1061]&~m[1062])|(~m[769]&m[1058]&~m[1060]&~m[1061]&m[1062])|(~m[769]&~m[1058]&m[1060]&~m[1061]&m[1062])|(m[769]&m[1058]&m[1060]&~m[1061]&m[1062])|(~m[769]&m[1058]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[522])|((m[769]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(~m[769]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[769]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[769]&m[1058]&~m[1060]&~m[1061]&m[1062])|(m[769]&~m[1058]&m[1060]&~m[1061]&m[1062])|(~m[769]&~m[1058]&~m[1060]&m[1061]&m[1062])|(m[769]&~m[1058]&~m[1060]&m[1061]&m[1062])|(~m[769]&m[1058]&~m[1060]&m[1061]&m[1062])|(m[769]&m[1058]&~m[1060]&m[1061]&m[1062])|(~m[769]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[769]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[769]&m[1058]&m[1060]&m[1061]&m[1062]));
    m[1064] = (((m[784]&~m[1063]&~m[1065]&~m[1066]&~m[1067])|(~m[784]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(m[784]&m[1063]&~m[1065]&m[1066]&~m[1067])|(m[784]&~m[1063]&m[1065]&m[1066]&~m[1067])|(~m[784]&m[1063]&~m[1065]&~m[1066]&m[1067])|(~m[784]&~m[1063]&m[1065]&~m[1066]&m[1067])|(m[784]&m[1063]&m[1065]&~m[1066]&m[1067])|(~m[784]&m[1063]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[523])|((m[784]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(~m[784]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[784]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[784]&m[1063]&~m[1065]&~m[1066]&m[1067])|(m[784]&~m[1063]&m[1065]&~m[1066]&m[1067])|(~m[784]&~m[1063]&~m[1065]&m[1066]&m[1067])|(m[784]&~m[1063]&~m[1065]&m[1066]&m[1067])|(~m[784]&m[1063]&~m[1065]&m[1066]&m[1067])|(m[784]&m[1063]&~m[1065]&m[1066]&m[1067])|(~m[784]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[784]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[784]&m[1063]&m[1065]&m[1066]&m[1067]));
    m[1069] = (((m[695]&~m[1068]&~m[1070]&~m[1071]&~m[1072])|(~m[695]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(m[695]&m[1068]&~m[1070]&m[1071]&~m[1072])|(m[695]&~m[1068]&m[1070]&m[1071]&~m[1072])|(~m[695]&m[1068]&~m[1070]&~m[1071]&m[1072])|(~m[695]&~m[1068]&m[1070]&~m[1071]&m[1072])|(m[695]&m[1068]&m[1070]&~m[1071]&m[1072])|(~m[695]&m[1068]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[524])|((m[695]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(~m[695]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[695]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[695]&m[1068]&~m[1070]&~m[1071]&m[1072])|(m[695]&~m[1068]&m[1070]&~m[1071]&m[1072])|(~m[695]&~m[1068]&~m[1070]&m[1071]&m[1072])|(m[695]&~m[1068]&~m[1070]&m[1071]&m[1072])|(~m[695]&m[1068]&~m[1070]&m[1071]&m[1072])|(m[695]&m[1068]&~m[1070]&m[1071]&m[1072])|(~m[695]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[695]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[695]&m[1068]&m[1070]&m[1071]&m[1072]));
    m[1074] = (((m[710]&~m[1073]&~m[1075]&~m[1076]&~m[1077])|(~m[710]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(m[710]&m[1073]&~m[1075]&m[1076]&~m[1077])|(m[710]&~m[1073]&m[1075]&m[1076]&~m[1077])|(~m[710]&m[1073]&~m[1075]&~m[1076]&m[1077])|(~m[710]&~m[1073]&m[1075]&~m[1076]&m[1077])|(m[710]&m[1073]&m[1075]&~m[1076]&m[1077])|(~m[710]&m[1073]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[525])|((m[710]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(~m[710]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[710]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[710]&m[1073]&~m[1075]&~m[1076]&m[1077])|(m[710]&~m[1073]&m[1075]&~m[1076]&m[1077])|(~m[710]&~m[1073]&~m[1075]&m[1076]&m[1077])|(m[710]&~m[1073]&~m[1075]&m[1076]&m[1077])|(~m[710]&m[1073]&~m[1075]&m[1076]&m[1077])|(m[710]&m[1073]&~m[1075]&m[1076]&m[1077])|(~m[710]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[710]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[710]&m[1073]&m[1075]&m[1076]&m[1077]));
    m[1079] = (((m[725]&~m[1078]&~m[1080]&~m[1081]&~m[1082])|(~m[725]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(m[725]&m[1078]&~m[1080]&m[1081]&~m[1082])|(m[725]&~m[1078]&m[1080]&m[1081]&~m[1082])|(~m[725]&m[1078]&~m[1080]&~m[1081]&m[1082])|(~m[725]&~m[1078]&m[1080]&~m[1081]&m[1082])|(m[725]&m[1078]&m[1080]&~m[1081]&m[1082])|(~m[725]&m[1078]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[526])|((m[725]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(~m[725]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[725]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[725]&m[1078]&~m[1080]&~m[1081]&m[1082])|(m[725]&~m[1078]&m[1080]&~m[1081]&m[1082])|(~m[725]&~m[1078]&~m[1080]&m[1081]&m[1082])|(m[725]&~m[1078]&~m[1080]&m[1081]&m[1082])|(~m[725]&m[1078]&~m[1080]&m[1081]&m[1082])|(m[725]&m[1078]&~m[1080]&m[1081]&m[1082])|(~m[725]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[725]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[725]&m[1078]&m[1080]&m[1081]&m[1082]));
    m[1084] = (((m[740]&~m[1083]&~m[1085]&~m[1086]&~m[1087])|(~m[740]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(m[740]&m[1083]&~m[1085]&m[1086]&~m[1087])|(m[740]&~m[1083]&m[1085]&m[1086]&~m[1087])|(~m[740]&m[1083]&~m[1085]&~m[1086]&m[1087])|(~m[740]&~m[1083]&m[1085]&~m[1086]&m[1087])|(m[740]&m[1083]&m[1085]&~m[1086]&m[1087])|(~m[740]&m[1083]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[527])|((m[740]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(~m[740]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[740]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[740]&m[1083]&~m[1085]&~m[1086]&m[1087])|(m[740]&~m[1083]&m[1085]&~m[1086]&m[1087])|(~m[740]&~m[1083]&~m[1085]&m[1086]&m[1087])|(m[740]&~m[1083]&~m[1085]&m[1086]&m[1087])|(~m[740]&m[1083]&~m[1085]&m[1086]&m[1087])|(m[740]&m[1083]&~m[1085]&m[1086]&m[1087])|(~m[740]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[740]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[740]&m[1083]&m[1085]&m[1086]&m[1087]));
    m[1089] = (((m[755]&~m[1088]&~m[1090]&~m[1091]&~m[1092])|(~m[755]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(m[755]&m[1088]&~m[1090]&m[1091]&~m[1092])|(m[755]&~m[1088]&m[1090]&m[1091]&~m[1092])|(~m[755]&m[1088]&~m[1090]&~m[1091]&m[1092])|(~m[755]&~m[1088]&m[1090]&~m[1091]&m[1092])|(m[755]&m[1088]&m[1090]&~m[1091]&m[1092])|(~m[755]&m[1088]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[528])|((m[755]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(~m[755]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[755]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[755]&m[1088]&~m[1090]&~m[1091]&m[1092])|(m[755]&~m[1088]&m[1090]&~m[1091]&m[1092])|(~m[755]&~m[1088]&~m[1090]&m[1091]&m[1092])|(m[755]&~m[1088]&~m[1090]&m[1091]&m[1092])|(~m[755]&m[1088]&~m[1090]&m[1091]&m[1092])|(m[755]&m[1088]&~m[1090]&m[1091]&m[1092])|(~m[755]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[755]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[755]&m[1088]&m[1090]&m[1091]&m[1092]));
    m[1094] = (((m[770]&~m[1093]&~m[1095]&~m[1096]&~m[1097])|(~m[770]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(m[770]&m[1093]&~m[1095]&m[1096]&~m[1097])|(m[770]&~m[1093]&m[1095]&m[1096]&~m[1097])|(~m[770]&m[1093]&~m[1095]&~m[1096]&m[1097])|(~m[770]&~m[1093]&m[1095]&~m[1096]&m[1097])|(m[770]&m[1093]&m[1095]&~m[1096]&m[1097])|(~m[770]&m[1093]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[529])|((m[770]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(~m[770]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[770]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[770]&m[1093]&~m[1095]&~m[1096]&m[1097])|(m[770]&~m[1093]&m[1095]&~m[1096]&m[1097])|(~m[770]&~m[1093]&~m[1095]&m[1096]&m[1097])|(m[770]&~m[1093]&~m[1095]&m[1096]&m[1097])|(~m[770]&m[1093]&~m[1095]&m[1096]&m[1097])|(m[770]&m[1093]&~m[1095]&m[1096]&m[1097])|(~m[770]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[770]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[770]&m[1093]&m[1095]&m[1096]&m[1097]));
    m[1099] = (((m[785]&~m[1098]&~m[1100]&~m[1101]&~m[1102])|(~m[785]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(m[785]&m[1098]&~m[1100]&m[1101]&~m[1102])|(m[785]&~m[1098]&m[1100]&m[1101]&~m[1102])|(~m[785]&m[1098]&~m[1100]&~m[1101]&m[1102])|(~m[785]&~m[1098]&m[1100]&~m[1101]&m[1102])|(m[785]&m[1098]&m[1100]&~m[1101]&m[1102])|(~m[785]&m[1098]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[530])|((m[785]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(~m[785]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[785]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[785]&m[1098]&~m[1100]&~m[1101]&m[1102])|(m[785]&~m[1098]&m[1100]&~m[1101]&m[1102])|(~m[785]&~m[1098]&~m[1100]&m[1101]&m[1102])|(m[785]&~m[1098]&~m[1100]&m[1101]&m[1102])|(~m[785]&m[1098]&~m[1100]&m[1101]&m[1102])|(m[785]&m[1098]&~m[1100]&m[1101]&m[1102])|(~m[785]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[785]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[785]&m[1098]&m[1100]&m[1101]&m[1102]));
    m[1104] = (((m[800]&~m[1103]&~m[1105]&~m[1106]&~m[1107])|(~m[800]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(m[800]&m[1103]&~m[1105]&m[1106]&~m[1107])|(m[800]&~m[1103]&m[1105]&m[1106]&~m[1107])|(~m[800]&m[1103]&~m[1105]&~m[1106]&m[1107])|(~m[800]&~m[1103]&m[1105]&~m[1106]&m[1107])|(m[800]&m[1103]&m[1105]&~m[1106]&m[1107])|(~m[800]&m[1103]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[531])|((m[800]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(~m[800]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[800]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[800]&m[1103]&~m[1105]&~m[1106]&m[1107])|(m[800]&~m[1103]&m[1105]&~m[1106]&m[1107])|(~m[800]&~m[1103]&~m[1105]&m[1106]&m[1107])|(m[800]&~m[1103]&~m[1105]&m[1106]&m[1107])|(~m[800]&m[1103]&~m[1105]&m[1106]&m[1107])|(m[800]&m[1103]&~m[1105]&m[1106]&m[1107])|(~m[800]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[800]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[800]&m[1103]&m[1105]&m[1106]&m[1107]));
    m[1109] = (((m[696]&~m[1108]&~m[1110]&~m[1111]&~m[1112])|(~m[696]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(m[696]&m[1108]&~m[1110]&m[1111]&~m[1112])|(m[696]&~m[1108]&m[1110]&m[1111]&~m[1112])|(~m[696]&m[1108]&~m[1110]&~m[1111]&m[1112])|(~m[696]&~m[1108]&m[1110]&~m[1111]&m[1112])|(m[696]&m[1108]&m[1110]&~m[1111]&m[1112])|(~m[696]&m[1108]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[532])|((m[696]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(~m[696]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[696]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[696]&m[1108]&~m[1110]&~m[1111]&m[1112])|(m[696]&~m[1108]&m[1110]&~m[1111]&m[1112])|(~m[696]&~m[1108]&~m[1110]&m[1111]&m[1112])|(m[696]&~m[1108]&~m[1110]&m[1111]&m[1112])|(~m[696]&m[1108]&~m[1110]&m[1111]&m[1112])|(m[696]&m[1108]&~m[1110]&m[1111]&m[1112])|(~m[696]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[696]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[696]&m[1108]&m[1110]&m[1111]&m[1112]));
    m[1114] = (((m[711]&~m[1113]&~m[1115]&~m[1116]&~m[1117])|(~m[711]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(m[711]&m[1113]&~m[1115]&m[1116]&~m[1117])|(m[711]&~m[1113]&m[1115]&m[1116]&~m[1117])|(~m[711]&m[1113]&~m[1115]&~m[1116]&m[1117])|(~m[711]&~m[1113]&m[1115]&~m[1116]&m[1117])|(m[711]&m[1113]&m[1115]&~m[1116]&m[1117])|(~m[711]&m[1113]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[533])|((m[711]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(~m[711]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[711]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[711]&m[1113]&~m[1115]&~m[1116]&m[1117])|(m[711]&~m[1113]&m[1115]&~m[1116]&m[1117])|(~m[711]&~m[1113]&~m[1115]&m[1116]&m[1117])|(m[711]&~m[1113]&~m[1115]&m[1116]&m[1117])|(~m[711]&m[1113]&~m[1115]&m[1116]&m[1117])|(m[711]&m[1113]&~m[1115]&m[1116]&m[1117])|(~m[711]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[711]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[711]&m[1113]&m[1115]&m[1116]&m[1117]));
    m[1119] = (((m[726]&~m[1118]&~m[1120]&~m[1121]&~m[1122])|(~m[726]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(m[726]&m[1118]&~m[1120]&m[1121]&~m[1122])|(m[726]&~m[1118]&m[1120]&m[1121]&~m[1122])|(~m[726]&m[1118]&~m[1120]&~m[1121]&m[1122])|(~m[726]&~m[1118]&m[1120]&~m[1121]&m[1122])|(m[726]&m[1118]&m[1120]&~m[1121]&m[1122])|(~m[726]&m[1118]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[534])|((m[726]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(~m[726]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[726]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[726]&m[1118]&~m[1120]&~m[1121]&m[1122])|(m[726]&~m[1118]&m[1120]&~m[1121]&m[1122])|(~m[726]&~m[1118]&~m[1120]&m[1121]&m[1122])|(m[726]&~m[1118]&~m[1120]&m[1121]&m[1122])|(~m[726]&m[1118]&~m[1120]&m[1121]&m[1122])|(m[726]&m[1118]&~m[1120]&m[1121]&m[1122])|(~m[726]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[726]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[726]&m[1118]&m[1120]&m[1121]&m[1122]));
    m[1124] = (((m[741]&~m[1123]&~m[1125]&~m[1126]&~m[1127])|(~m[741]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(m[741]&m[1123]&~m[1125]&m[1126]&~m[1127])|(m[741]&~m[1123]&m[1125]&m[1126]&~m[1127])|(~m[741]&m[1123]&~m[1125]&~m[1126]&m[1127])|(~m[741]&~m[1123]&m[1125]&~m[1126]&m[1127])|(m[741]&m[1123]&m[1125]&~m[1126]&m[1127])|(~m[741]&m[1123]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[535])|((m[741]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(~m[741]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[741]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[741]&m[1123]&~m[1125]&~m[1126]&m[1127])|(m[741]&~m[1123]&m[1125]&~m[1126]&m[1127])|(~m[741]&~m[1123]&~m[1125]&m[1126]&m[1127])|(m[741]&~m[1123]&~m[1125]&m[1126]&m[1127])|(~m[741]&m[1123]&~m[1125]&m[1126]&m[1127])|(m[741]&m[1123]&~m[1125]&m[1126]&m[1127])|(~m[741]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[741]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[741]&m[1123]&m[1125]&m[1126]&m[1127]));
    m[1129] = (((m[756]&~m[1128]&~m[1130]&~m[1131]&~m[1132])|(~m[756]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(m[756]&m[1128]&~m[1130]&m[1131]&~m[1132])|(m[756]&~m[1128]&m[1130]&m[1131]&~m[1132])|(~m[756]&m[1128]&~m[1130]&~m[1131]&m[1132])|(~m[756]&~m[1128]&m[1130]&~m[1131]&m[1132])|(m[756]&m[1128]&m[1130]&~m[1131]&m[1132])|(~m[756]&m[1128]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[536])|((m[756]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(~m[756]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[756]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[756]&m[1128]&~m[1130]&~m[1131]&m[1132])|(m[756]&~m[1128]&m[1130]&~m[1131]&m[1132])|(~m[756]&~m[1128]&~m[1130]&m[1131]&m[1132])|(m[756]&~m[1128]&~m[1130]&m[1131]&m[1132])|(~m[756]&m[1128]&~m[1130]&m[1131]&m[1132])|(m[756]&m[1128]&~m[1130]&m[1131]&m[1132])|(~m[756]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[756]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[756]&m[1128]&m[1130]&m[1131]&m[1132]));
    m[1134] = (((m[771]&~m[1133]&~m[1135]&~m[1136]&~m[1137])|(~m[771]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(m[771]&m[1133]&~m[1135]&m[1136]&~m[1137])|(m[771]&~m[1133]&m[1135]&m[1136]&~m[1137])|(~m[771]&m[1133]&~m[1135]&~m[1136]&m[1137])|(~m[771]&~m[1133]&m[1135]&~m[1136]&m[1137])|(m[771]&m[1133]&m[1135]&~m[1136]&m[1137])|(~m[771]&m[1133]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[537])|((m[771]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(~m[771]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[771]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[771]&m[1133]&~m[1135]&~m[1136]&m[1137])|(m[771]&~m[1133]&m[1135]&~m[1136]&m[1137])|(~m[771]&~m[1133]&~m[1135]&m[1136]&m[1137])|(m[771]&~m[1133]&~m[1135]&m[1136]&m[1137])|(~m[771]&m[1133]&~m[1135]&m[1136]&m[1137])|(m[771]&m[1133]&~m[1135]&m[1136]&m[1137])|(~m[771]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[771]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[771]&m[1133]&m[1135]&m[1136]&m[1137]));
    m[1139] = (((m[786]&~m[1138]&~m[1140]&~m[1141]&~m[1142])|(~m[786]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(m[786]&m[1138]&~m[1140]&m[1141]&~m[1142])|(m[786]&~m[1138]&m[1140]&m[1141]&~m[1142])|(~m[786]&m[1138]&~m[1140]&~m[1141]&m[1142])|(~m[786]&~m[1138]&m[1140]&~m[1141]&m[1142])|(m[786]&m[1138]&m[1140]&~m[1141]&m[1142])|(~m[786]&m[1138]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[538])|((m[786]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(~m[786]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[786]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[786]&m[1138]&~m[1140]&~m[1141]&m[1142])|(m[786]&~m[1138]&m[1140]&~m[1141]&m[1142])|(~m[786]&~m[1138]&~m[1140]&m[1141]&m[1142])|(m[786]&~m[1138]&~m[1140]&m[1141]&m[1142])|(~m[786]&m[1138]&~m[1140]&m[1141]&m[1142])|(m[786]&m[1138]&~m[1140]&m[1141]&m[1142])|(~m[786]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[786]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[786]&m[1138]&m[1140]&m[1141]&m[1142]));
    m[1144] = (((m[801]&~m[1143]&~m[1145]&~m[1146]&~m[1147])|(~m[801]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(m[801]&m[1143]&~m[1145]&m[1146]&~m[1147])|(m[801]&~m[1143]&m[1145]&m[1146]&~m[1147])|(~m[801]&m[1143]&~m[1145]&~m[1146]&m[1147])|(~m[801]&~m[1143]&m[1145]&~m[1146]&m[1147])|(m[801]&m[1143]&m[1145]&~m[1146]&m[1147])|(~m[801]&m[1143]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[539])|((m[801]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(~m[801]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[801]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[801]&m[1143]&~m[1145]&~m[1146]&m[1147])|(m[801]&~m[1143]&m[1145]&~m[1146]&m[1147])|(~m[801]&~m[1143]&~m[1145]&m[1146]&m[1147])|(m[801]&~m[1143]&~m[1145]&m[1146]&m[1147])|(~m[801]&m[1143]&~m[1145]&m[1146]&m[1147])|(m[801]&m[1143]&~m[1145]&m[1146]&m[1147])|(~m[801]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[801]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[801]&m[1143]&m[1145]&m[1146]&m[1147]));
    m[1149] = (((m[816]&~m[1148]&~m[1150]&~m[1151]&~m[1152])|(~m[816]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(m[816]&m[1148]&~m[1150]&m[1151]&~m[1152])|(m[816]&~m[1148]&m[1150]&m[1151]&~m[1152])|(~m[816]&m[1148]&~m[1150]&~m[1151]&m[1152])|(~m[816]&~m[1148]&m[1150]&~m[1151]&m[1152])|(m[816]&m[1148]&m[1150]&~m[1151]&m[1152])|(~m[816]&m[1148]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[540])|((m[816]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(~m[816]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[816]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[816]&m[1148]&~m[1150]&~m[1151]&m[1152])|(m[816]&~m[1148]&m[1150]&~m[1151]&m[1152])|(~m[816]&~m[1148]&~m[1150]&m[1151]&m[1152])|(m[816]&~m[1148]&~m[1150]&m[1151]&m[1152])|(~m[816]&m[1148]&~m[1150]&m[1151]&m[1152])|(m[816]&m[1148]&~m[1150]&m[1151]&m[1152])|(~m[816]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[816]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[816]&m[1148]&m[1150]&m[1151]&m[1152]));
    m[1154] = (((m[697]&~m[1153]&~m[1155]&~m[1156]&~m[1157])|(~m[697]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(m[697]&m[1153]&~m[1155]&m[1156]&~m[1157])|(m[697]&~m[1153]&m[1155]&m[1156]&~m[1157])|(~m[697]&m[1153]&~m[1155]&~m[1156]&m[1157])|(~m[697]&~m[1153]&m[1155]&~m[1156]&m[1157])|(m[697]&m[1153]&m[1155]&~m[1156]&m[1157])|(~m[697]&m[1153]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[541])|((m[697]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(~m[697]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[697]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[697]&m[1153]&~m[1155]&~m[1156]&m[1157])|(m[697]&~m[1153]&m[1155]&~m[1156]&m[1157])|(~m[697]&~m[1153]&~m[1155]&m[1156]&m[1157])|(m[697]&~m[1153]&~m[1155]&m[1156]&m[1157])|(~m[697]&m[1153]&~m[1155]&m[1156]&m[1157])|(m[697]&m[1153]&~m[1155]&m[1156]&m[1157])|(~m[697]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[697]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[697]&m[1153]&m[1155]&m[1156]&m[1157]));
    m[1159] = (((m[712]&~m[1158]&~m[1160]&~m[1161]&~m[1162])|(~m[712]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(m[712]&m[1158]&~m[1160]&m[1161]&~m[1162])|(m[712]&~m[1158]&m[1160]&m[1161]&~m[1162])|(~m[712]&m[1158]&~m[1160]&~m[1161]&m[1162])|(~m[712]&~m[1158]&m[1160]&~m[1161]&m[1162])|(m[712]&m[1158]&m[1160]&~m[1161]&m[1162])|(~m[712]&m[1158]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[542])|((m[712]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(~m[712]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[712]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[712]&m[1158]&~m[1160]&~m[1161]&m[1162])|(m[712]&~m[1158]&m[1160]&~m[1161]&m[1162])|(~m[712]&~m[1158]&~m[1160]&m[1161]&m[1162])|(m[712]&~m[1158]&~m[1160]&m[1161]&m[1162])|(~m[712]&m[1158]&~m[1160]&m[1161]&m[1162])|(m[712]&m[1158]&~m[1160]&m[1161]&m[1162])|(~m[712]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[712]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[712]&m[1158]&m[1160]&m[1161]&m[1162]));
    m[1164] = (((m[727]&~m[1163]&~m[1165]&~m[1166]&~m[1167])|(~m[727]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(m[727]&m[1163]&~m[1165]&m[1166]&~m[1167])|(m[727]&~m[1163]&m[1165]&m[1166]&~m[1167])|(~m[727]&m[1163]&~m[1165]&~m[1166]&m[1167])|(~m[727]&~m[1163]&m[1165]&~m[1166]&m[1167])|(m[727]&m[1163]&m[1165]&~m[1166]&m[1167])|(~m[727]&m[1163]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[543])|((m[727]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(~m[727]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[727]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[727]&m[1163]&~m[1165]&~m[1166]&m[1167])|(m[727]&~m[1163]&m[1165]&~m[1166]&m[1167])|(~m[727]&~m[1163]&~m[1165]&m[1166]&m[1167])|(m[727]&~m[1163]&~m[1165]&m[1166]&m[1167])|(~m[727]&m[1163]&~m[1165]&m[1166]&m[1167])|(m[727]&m[1163]&~m[1165]&m[1166]&m[1167])|(~m[727]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[727]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[727]&m[1163]&m[1165]&m[1166]&m[1167]));
    m[1169] = (((m[742]&~m[1168]&~m[1170]&~m[1171]&~m[1172])|(~m[742]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(m[742]&m[1168]&~m[1170]&m[1171]&~m[1172])|(m[742]&~m[1168]&m[1170]&m[1171]&~m[1172])|(~m[742]&m[1168]&~m[1170]&~m[1171]&m[1172])|(~m[742]&~m[1168]&m[1170]&~m[1171]&m[1172])|(m[742]&m[1168]&m[1170]&~m[1171]&m[1172])|(~m[742]&m[1168]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[544])|((m[742]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(~m[742]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[742]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[742]&m[1168]&~m[1170]&~m[1171]&m[1172])|(m[742]&~m[1168]&m[1170]&~m[1171]&m[1172])|(~m[742]&~m[1168]&~m[1170]&m[1171]&m[1172])|(m[742]&~m[1168]&~m[1170]&m[1171]&m[1172])|(~m[742]&m[1168]&~m[1170]&m[1171]&m[1172])|(m[742]&m[1168]&~m[1170]&m[1171]&m[1172])|(~m[742]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[742]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[742]&m[1168]&m[1170]&m[1171]&m[1172]));
    m[1174] = (((m[757]&~m[1173]&~m[1175]&~m[1176]&~m[1177])|(~m[757]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(m[757]&m[1173]&~m[1175]&m[1176]&~m[1177])|(m[757]&~m[1173]&m[1175]&m[1176]&~m[1177])|(~m[757]&m[1173]&~m[1175]&~m[1176]&m[1177])|(~m[757]&~m[1173]&m[1175]&~m[1176]&m[1177])|(m[757]&m[1173]&m[1175]&~m[1176]&m[1177])|(~m[757]&m[1173]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[545])|((m[757]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(~m[757]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[757]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[757]&m[1173]&~m[1175]&~m[1176]&m[1177])|(m[757]&~m[1173]&m[1175]&~m[1176]&m[1177])|(~m[757]&~m[1173]&~m[1175]&m[1176]&m[1177])|(m[757]&~m[1173]&~m[1175]&m[1176]&m[1177])|(~m[757]&m[1173]&~m[1175]&m[1176]&m[1177])|(m[757]&m[1173]&~m[1175]&m[1176]&m[1177])|(~m[757]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[757]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[757]&m[1173]&m[1175]&m[1176]&m[1177]));
    m[1179] = (((m[772]&~m[1178]&~m[1180]&~m[1181]&~m[1182])|(~m[772]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(m[772]&m[1178]&~m[1180]&m[1181]&~m[1182])|(m[772]&~m[1178]&m[1180]&m[1181]&~m[1182])|(~m[772]&m[1178]&~m[1180]&~m[1181]&m[1182])|(~m[772]&~m[1178]&m[1180]&~m[1181]&m[1182])|(m[772]&m[1178]&m[1180]&~m[1181]&m[1182])|(~m[772]&m[1178]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[546])|((m[772]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(~m[772]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[772]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[772]&m[1178]&~m[1180]&~m[1181]&m[1182])|(m[772]&~m[1178]&m[1180]&~m[1181]&m[1182])|(~m[772]&~m[1178]&~m[1180]&m[1181]&m[1182])|(m[772]&~m[1178]&~m[1180]&m[1181]&m[1182])|(~m[772]&m[1178]&~m[1180]&m[1181]&m[1182])|(m[772]&m[1178]&~m[1180]&m[1181]&m[1182])|(~m[772]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[772]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[772]&m[1178]&m[1180]&m[1181]&m[1182]));
    m[1184] = (((m[787]&~m[1183]&~m[1185]&~m[1186]&~m[1187])|(~m[787]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(m[787]&m[1183]&~m[1185]&m[1186]&~m[1187])|(m[787]&~m[1183]&m[1185]&m[1186]&~m[1187])|(~m[787]&m[1183]&~m[1185]&~m[1186]&m[1187])|(~m[787]&~m[1183]&m[1185]&~m[1186]&m[1187])|(m[787]&m[1183]&m[1185]&~m[1186]&m[1187])|(~m[787]&m[1183]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[547])|((m[787]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(~m[787]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[787]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[787]&m[1183]&~m[1185]&~m[1186]&m[1187])|(m[787]&~m[1183]&m[1185]&~m[1186]&m[1187])|(~m[787]&~m[1183]&~m[1185]&m[1186]&m[1187])|(m[787]&~m[1183]&~m[1185]&m[1186]&m[1187])|(~m[787]&m[1183]&~m[1185]&m[1186]&m[1187])|(m[787]&m[1183]&~m[1185]&m[1186]&m[1187])|(~m[787]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[787]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[787]&m[1183]&m[1185]&m[1186]&m[1187]));
    m[1189] = (((m[802]&~m[1188]&~m[1190]&~m[1191]&~m[1192])|(~m[802]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(m[802]&m[1188]&~m[1190]&m[1191]&~m[1192])|(m[802]&~m[1188]&m[1190]&m[1191]&~m[1192])|(~m[802]&m[1188]&~m[1190]&~m[1191]&m[1192])|(~m[802]&~m[1188]&m[1190]&~m[1191]&m[1192])|(m[802]&m[1188]&m[1190]&~m[1191]&m[1192])|(~m[802]&m[1188]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[548])|((m[802]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(~m[802]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[802]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[802]&m[1188]&~m[1190]&~m[1191]&m[1192])|(m[802]&~m[1188]&m[1190]&~m[1191]&m[1192])|(~m[802]&~m[1188]&~m[1190]&m[1191]&m[1192])|(m[802]&~m[1188]&~m[1190]&m[1191]&m[1192])|(~m[802]&m[1188]&~m[1190]&m[1191]&m[1192])|(m[802]&m[1188]&~m[1190]&m[1191]&m[1192])|(~m[802]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[802]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[802]&m[1188]&m[1190]&m[1191]&m[1192]));
    m[1194] = (((m[817]&~m[1193]&~m[1195]&~m[1196]&~m[1197])|(~m[817]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(m[817]&m[1193]&~m[1195]&m[1196]&~m[1197])|(m[817]&~m[1193]&m[1195]&m[1196]&~m[1197])|(~m[817]&m[1193]&~m[1195]&~m[1196]&m[1197])|(~m[817]&~m[1193]&m[1195]&~m[1196]&m[1197])|(m[817]&m[1193]&m[1195]&~m[1196]&m[1197])|(~m[817]&m[1193]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[549])|((m[817]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(~m[817]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[817]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[817]&m[1193]&~m[1195]&~m[1196]&m[1197])|(m[817]&~m[1193]&m[1195]&~m[1196]&m[1197])|(~m[817]&~m[1193]&~m[1195]&m[1196]&m[1197])|(m[817]&~m[1193]&~m[1195]&m[1196]&m[1197])|(~m[817]&m[1193]&~m[1195]&m[1196]&m[1197])|(m[817]&m[1193]&~m[1195]&m[1196]&m[1197])|(~m[817]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[817]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[817]&m[1193]&m[1195]&m[1196]&m[1197]));
    m[1199] = (((m[832]&~m[1198]&~m[1200]&~m[1201]&~m[1202])|(~m[832]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(m[832]&m[1198]&~m[1200]&m[1201]&~m[1202])|(m[832]&~m[1198]&m[1200]&m[1201]&~m[1202])|(~m[832]&m[1198]&~m[1200]&~m[1201]&m[1202])|(~m[832]&~m[1198]&m[1200]&~m[1201]&m[1202])|(m[832]&m[1198]&m[1200]&~m[1201]&m[1202])|(~m[832]&m[1198]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[550])|((m[832]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(~m[832]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[832]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[832]&m[1198]&~m[1200]&~m[1201]&m[1202])|(m[832]&~m[1198]&m[1200]&~m[1201]&m[1202])|(~m[832]&~m[1198]&~m[1200]&m[1201]&m[1202])|(m[832]&~m[1198]&~m[1200]&m[1201]&m[1202])|(~m[832]&m[1198]&~m[1200]&m[1201]&m[1202])|(m[832]&m[1198]&~m[1200]&m[1201]&m[1202])|(~m[832]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[832]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[832]&m[1198]&m[1200]&m[1201]&m[1202]));
    m[1204] = (((m[698]&~m[1203]&~m[1205]&~m[1206]&~m[1207])|(~m[698]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(m[698]&m[1203]&~m[1205]&m[1206]&~m[1207])|(m[698]&~m[1203]&m[1205]&m[1206]&~m[1207])|(~m[698]&m[1203]&~m[1205]&~m[1206]&m[1207])|(~m[698]&~m[1203]&m[1205]&~m[1206]&m[1207])|(m[698]&m[1203]&m[1205]&~m[1206]&m[1207])|(~m[698]&m[1203]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[551])|((m[698]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(~m[698]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[698]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[698]&m[1203]&~m[1205]&~m[1206]&m[1207])|(m[698]&~m[1203]&m[1205]&~m[1206]&m[1207])|(~m[698]&~m[1203]&~m[1205]&m[1206]&m[1207])|(m[698]&~m[1203]&~m[1205]&m[1206]&m[1207])|(~m[698]&m[1203]&~m[1205]&m[1206]&m[1207])|(m[698]&m[1203]&~m[1205]&m[1206]&m[1207])|(~m[698]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[698]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[698]&m[1203]&m[1205]&m[1206]&m[1207]));
    m[1209] = (((m[713]&~m[1208]&~m[1210]&~m[1211]&~m[1212])|(~m[713]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(m[713]&m[1208]&~m[1210]&m[1211]&~m[1212])|(m[713]&~m[1208]&m[1210]&m[1211]&~m[1212])|(~m[713]&m[1208]&~m[1210]&~m[1211]&m[1212])|(~m[713]&~m[1208]&m[1210]&~m[1211]&m[1212])|(m[713]&m[1208]&m[1210]&~m[1211]&m[1212])|(~m[713]&m[1208]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[552])|((m[713]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(~m[713]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[713]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[713]&m[1208]&~m[1210]&~m[1211]&m[1212])|(m[713]&~m[1208]&m[1210]&~m[1211]&m[1212])|(~m[713]&~m[1208]&~m[1210]&m[1211]&m[1212])|(m[713]&~m[1208]&~m[1210]&m[1211]&m[1212])|(~m[713]&m[1208]&~m[1210]&m[1211]&m[1212])|(m[713]&m[1208]&~m[1210]&m[1211]&m[1212])|(~m[713]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[713]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[713]&m[1208]&m[1210]&m[1211]&m[1212]));
    m[1214] = (((m[728]&~m[1213]&~m[1215]&~m[1216]&~m[1217])|(~m[728]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(m[728]&m[1213]&~m[1215]&m[1216]&~m[1217])|(m[728]&~m[1213]&m[1215]&m[1216]&~m[1217])|(~m[728]&m[1213]&~m[1215]&~m[1216]&m[1217])|(~m[728]&~m[1213]&m[1215]&~m[1216]&m[1217])|(m[728]&m[1213]&m[1215]&~m[1216]&m[1217])|(~m[728]&m[1213]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[553])|((m[728]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(~m[728]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[728]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[728]&m[1213]&~m[1215]&~m[1216]&m[1217])|(m[728]&~m[1213]&m[1215]&~m[1216]&m[1217])|(~m[728]&~m[1213]&~m[1215]&m[1216]&m[1217])|(m[728]&~m[1213]&~m[1215]&m[1216]&m[1217])|(~m[728]&m[1213]&~m[1215]&m[1216]&m[1217])|(m[728]&m[1213]&~m[1215]&m[1216]&m[1217])|(~m[728]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[728]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[728]&m[1213]&m[1215]&m[1216]&m[1217]));
    m[1219] = (((m[743]&~m[1218]&~m[1220]&~m[1221]&~m[1222])|(~m[743]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(m[743]&m[1218]&~m[1220]&m[1221]&~m[1222])|(m[743]&~m[1218]&m[1220]&m[1221]&~m[1222])|(~m[743]&m[1218]&~m[1220]&~m[1221]&m[1222])|(~m[743]&~m[1218]&m[1220]&~m[1221]&m[1222])|(m[743]&m[1218]&m[1220]&~m[1221]&m[1222])|(~m[743]&m[1218]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[554])|((m[743]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(~m[743]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[743]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[743]&m[1218]&~m[1220]&~m[1221]&m[1222])|(m[743]&~m[1218]&m[1220]&~m[1221]&m[1222])|(~m[743]&~m[1218]&~m[1220]&m[1221]&m[1222])|(m[743]&~m[1218]&~m[1220]&m[1221]&m[1222])|(~m[743]&m[1218]&~m[1220]&m[1221]&m[1222])|(m[743]&m[1218]&~m[1220]&m[1221]&m[1222])|(~m[743]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[743]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[743]&m[1218]&m[1220]&m[1221]&m[1222]));
    m[1224] = (((m[758]&~m[1223]&~m[1225]&~m[1226]&~m[1227])|(~m[758]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(m[758]&m[1223]&~m[1225]&m[1226]&~m[1227])|(m[758]&~m[1223]&m[1225]&m[1226]&~m[1227])|(~m[758]&m[1223]&~m[1225]&~m[1226]&m[1227])|(~m[758]&~m[1223]&m[1225]&~m[1226]&m[1227])|(m[758]&m[1223]&m[1225]&~m[1226]&m[1227])|(~m[758]&m[1223]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[555])|((m[758]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(~m[758]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[758]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[758]&m[1223]&~m[1225]&~m[1226]&m[1227])|(m[758]&~m[1223]&m[1225]&~m[1226]&m[1227])|(~m[758]&~m[1223]&~m[1225]&m[1226]&m[1227])|(m[758]&~m[1223]&~m[1225]&m[1226]&m[1227])|(~m[758]&m[1223]&~m[1225]&m[1226]&m[1227])|(m[758]&m[1223]&~m[1225]&m[1226]&m[1227])|(~m[758]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[758]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[758]&m[1223]&m[1225]&m[1226]&m[1227]));
    m[1229] = (((m[773]&~m[1228]&~m[1230]&~m[1231]&~m[1232])|(~m[773]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(m[773]&m[1228]&~m[1230]&m[1231]&~m[1232])|(m[773]&~m[1228]&m[1230]&m[1231]&~m[1232])|(~m[773]&m[1228]&~m[1230]&~m[1231]&m[1232])|(~m[773]&~m[1228]&m[1230]&~m[1231]&m[1232])|(m[773]&m[1228]&m[1230]&~m[1231]&m[1232])|(~m[773]&m[1228]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[556])|((m[773]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(~m[773]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[773]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[773]&m[1228]&~m[1230]&~m[1231]&m[1232])|(m[773]&~m[1228]&m[1230]&~m[1231]&m[1232])|(~m[773]&~m[1228]&~m[1230]&m[1231]&m[1232])|(m[773]&~m[1228]&~m[1230]&m[1231]&m[1232])|(~m[773]&m[1228]&~m[1230]&m[1231]&m[1232])|(m[773]&m[1228]&~m[1230]&m[1231]&m[1232])|(~m[773]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[773]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[773]&m[1228]&m[1230]&m[1231]&m[1232]));
    m[1234] = (((m[788]&~m[1233]&~m[1235]&~m[1236]&~m[1237])|(~m[788]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(m[788]&m[1233]&~m[1235]&m[1236]&~m[1237])|(m[788]&~m[1233]&m[1235]&m[1236]&~m[1237])|(~m[788]&m[1233]&~m[1235]&~m[1236]&m[1237])|(~m[788]&~m[1233]&m[1235]&~m[1236]&m[1237])|(m[788]&m[1233]&m[1235]&~m[1236]&m[1237])|(~m[788]&m[1233]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[557])|((m[788]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(~m[788]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[788]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[788]&m[1233]&~m[1235]&~m[1236]&m[1237])|(m[788]&~m[1233]&m[1235]&~m[1236]&m[1237])|(~m[788]&~m[1233]&~m[1235]&m[1236]&m[1237])|(m[788]&~m[1233]&~m[1235]&m[1236]&m[1237])|(~m[788]&m[1233]&~m[1235]&m[1236]&m[1237])|(m[788]&m[1233]&~m[1235]&m[1236]&m[1237])|(~m[788]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[788]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[788]&m[1233]&m[1235]&m[1236]&m[1237]));
    m[1239] = (((m[803]&~m[1238]&~m[1240]&~m[1241]&~m[1242])|(~m[803]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(m[803]&m[1238]&~m[1240]&m[1241]&~m[1242])|(m[803]&~m[1238]&m[1240]&m[1241]&~m[1242])|(~m[803]&m[1238]&~m[1240]&~m[1241]&m[1242])|(~m[803]&~m[1238]&m[1240]&~m[1241]&m[1242])|(m[803]&m[1238]&m[1240]&~m[1241]&m[1242])|(~m[803]&m[1238]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[558])|((m[803]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(~m[803]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[803]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[803]&m[1238]&~m[1240]&~m[1241]&m[1242])|(m[803]&~m[1238]&m[1240]&~m[1241]&m[1242])|(~m[803]&~m[1238]&~m[1240]&m[1241]&m[1242])|(m[803]&~m[1238]&~m[1240]&m[1241]&m[1242])|(~m[803]&m[1238]&~m[1240]&m[1241]&m[1242])|(m[803]&m[1238]&~m[1240]&m[1241]&m[1242])|(~m[803]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[803]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[803]&m[1238]&m[1240]&m[1241]&m[1242]));
    m[1244] = (((m[818]&~m[1243]&~m[1245]&~m[1246]&~m[1247])|(~m[818]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(m[818]&m[1243]&~m[1245]&m[1246]&~m[1247])|(m[818]&~m[1243]&m[1245]&m[1246]&~m[1247])|(~m[818]&m[1243]&~m[1245]&~m[1246]&m[1247])|(~m[818]&~m[1243]&m[1245]&~m[1246]&m[1247])|(m[818]&m[1243]&m[1245]&~m[1246]&m[1247])|(~m[818]&m[1243]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[559])|((m[818]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(~m[818]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[818]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[818]&m[1243]&~m[1245]&~m[1246]&m[1247])|(m[818]&~m[1243]&m[1245]&~m[1246]&m[1247])|(~m[818]&~m[1243]&~m[1245]&m[1246]&m[1247])|(m[818]&~m[1243]&~m[1245]&m[1246]&m[1247])|(~m[818]&m[1243]&~m[1245]&m[1246]&m[1247])|(m[818]&m[1243]&~m[1245]&m[1246]&m[1247])|(~m[818]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[818]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[818]&m[1243]&m[1245]&m[1246]&m[1247]));
    m[1249] = (((m[833]&~m[1248]&~m[1250]&~m[1251]&~m[1252])|(~m[833]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(m[833]&m[1248]&~m[1250]&m[1251]&~m[1252])|(m[833]&~m[1248]&m[1250]&m[1251]&~m[1252])|(~m[833]&m[1248]&~m[1250]&~m[1251]&m[1252])|(~m[833]&~m[1248]&m[1250]&~m[1251]&m[1252])|(m[833]&m[1248]&m[1250]&~m[1251]&m[1252])|(~m[833]&m[1248]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[560])|((m[833]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(~m[833]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[833]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[833]&m[1248]&~m[1250]&~m[1251]&m[1252])|(m[833]&~m[1248]&m[1250]&~m[1251]&m[1252])|(~m[833]&~m[1248]&~m[1250]&m[1251]&m[1252])|(m[833]&~m[1248]&~m[1250]&m[1251]&m[1252])|(~m[833]&m[1248]&~m[1250]&m[1251]&m[1252])|(m[833]&m[1248]&~m[1250]&m[1251]&m[1252])|(~m[833]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[833]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[833]&m[1248]&m[1250]&m[1251]&m[1252]));
    m[1254] = (((m[848]&~m[1253]&~m[1255]&~m[1256]&~m[1257])|(~m[848]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(m[848]&m[1253]&~m[1255]&m[1256]&~m[1257])|(m[848]&~m[1253]&m[1255]&m[1256]&~m[1257])|(~m[848]&m[1253]&~m[1255]&~m[1256]&m[1257])|(~m[848]&~m[1253]&m[1255]&~m[1256]&m[1257])|(m[848]&m[1253]&m[1255]&~m[1256]&m[1257])|(~m[848]&m[1253]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[561])|((m[848]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(~m[848]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[848]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[848]&m[1253]&~m[1255]&~m[1256]&m[1257])|(m[848]&~m[1253]&m[1255]&~m[1256]&m[1257])|(~m[848]&~m[1253]&~m[1255]&m[1256]&m[1257])|(m[848]&~m[1253]&~m[1255]&m[1256]&m[1257])|(~m[848]&m[1253]&~m[1255]&m[1256]&m[1257])|(m[848]&m[1253]&~m[1255]&m[1256]&m[1257])|(~m[848]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[848]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[848]&m[1253]&m[1255]&m[1256]&m[1257]));
    m[1259] = (((m[699]&~m[1258]&~m[1260]&~m[1261]&~m[1262])|(~m[699]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(m[699]&m[1258]&~m[1260]&m[1261]&~m[1262])|(m[699]&~m[1258]&m[1260]&m[1261]&~m[1262])|(~m[699]&m[1258]&~m[1260]&~m[1261]&m[1262])|(~m[699]&~m[1258]&m[1260]&~m[1261]&m[1262])|(m[699]&m[1258]&m[1260]&~m[1261]&m[1262])|(~m[699]&m[1258]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[562])|((m[699]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(~m[699]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[699]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[699]&m[1258]&~m[1260]&~m[1261]&m[1262])|(m[699]&~m[1258]&m[1260]&~m[1261]&m[1262])|(~m[699]&~m[1258]&~m[1260]&m[1261]&m[1262])|(m[699]&~m[1258]&~m[1260]&m[1261]&m[1262])|(~m[699]&m[1258]&~m[1260]&m[1261]&m[1262])|(m[699]&m[1258]&~m[1260]&m[1261]&m[1262])|(~m[699]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[699]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[699]&m[1258]&m[1260]&m[1261]&m[1262]));
    m[1264] = (((m[714]&~m[1263]&~m[1265]&~m[1266]&~m[1267])|(~m[714]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(m[714]&m[1263]&~m[1265]&m[1266]&~m[1267])|(m[714]&~m[1263]&m[1265]&m[1266]&~m[1267])|(~m[714]&m[1263]&~m[1265]&~m[1266]&m[1267])|(~m[714]&~m[1263]&m[1265]&~m[1266]&m[1267])|(m[714]&m[1263]&m[1265]&~m[1266]&m[1267])|(~m[714]&m[1263]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[563])|((m[714]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(~m[714]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[714]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[714]&m[1263]&~m[1265]&~m[1266]&m[1267])|(m[714]&~m[1263]&m[1265]&~m[1266]&m[1267])|(~m[714]&~m[1263]&~m[1265]&m[1266]&m[1267])|(m[714]&~m[1263]&~m[1265]&m[1266]&m[1267])|(~m[714]&m[1263]&~m[1265]&m[1266]&m[1267])|(m[714]&m[1263]&~m[1265]&m[1266]&m[1267])|(~m[714]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[714]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[714]&m[1263]&m[1265]&m[1266]&m[1267]));
    m[1269] = (((m[729]&~m[1268]&~m[1270]&~m[1271]&~m[1272])|(~m[729]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(m[729]&m[1268]&~m[1270]&m[1271]&~m[1272])|(m[729]&~m[1268]&m[1270]&m[1271]&~m[1272])|(~m[729]&m[1268]&~m[1270]&~m[1271]&m[1272])|(~m[729]&~m[1268]&m[1270]&~m[1271]&m[1272])|(m[729]&m[1268]&m[1270]&~m[1271]&m[1272])|(~m[729]&m[1268]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[564])|((m[729]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(~m[729]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[729]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[729]&m[1268]&~m[1270]&~m[1271]&m[1272])|(m[729]&~m[1268]&m[1270]&~m[1271]&m[1272])|(~m[729]&~m[1268]&~m[1270]&m[1271]&m[1272])|(m[729]&~m[1268]&~m[1270]&m[1271]&m[1272])|(~m[729]&m[1268]&~m[1270]&m[1271]&m[1272])|(m[729]&m[1268]&~m[1270]&m[1271]&m[1272])|(~m[729]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[729]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[729]&m[1268]&m[1270]&m[1271]&m[1272]));
    m[1274] = (((m[744]&~m[1273]&~m[1275]&~m[1276]&~m[1277])|(~m[744]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(m[744]&m[1273]&~m[1275]&m[1276]&~m[1277])|(m[744]&~m[1273]&m[1275]&m[1276]&~m[1277])|(~m[744]&m[1273]&~m[1275]&~m[1276]&m[1277])|(~m[744]&~m[1273]&m[1275]&~m[1276]&m[1277])|(m[744]&m[1273]&m[1275]&~m[1276]&m[1277])|(~m[744]&m[1273]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[565])|((m[744]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(~m[744]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[744]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[744]&m[1273]&~m[1275]&~m[1276]&m[1277])|(m[744]&~m[1273]&m[1275]&~m[1276]&m[1277])|(~m[744]&~m[1273]&~m[1275]&m[1276]&m[1277])|(m[744]&~m[1273]&~m[1275]&m[1276]&m[1277])|(~m[744]&m[1273]&~m[1275]&m[1276]&m[1277])|(m[744]&m[1273]&~m[1275]&m[1276]&m[1277])|(~m[744]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[744]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[744]&m[1273]&m[1275]&m[1276]&m[1277]));
    m[1279] = (((m[759]&~m[1278]&~m[1280]&~m[1281]&~m[1282])|(~m[759]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(m[759]&m[1278]&~m[1280]&m[1281]&~m[1282])|(m[759]&~m[1278]&m[1280]&m[1281]&~m[1282])|(~m[759]&m[1278]&~m[1280]&~m[1281]&m[1282])|(~m[759]&~m[1278]&m[1280]&~m[1281]&m[1282])|(m[759]&m[1278]&m[1280]&~m[1281]&m[1282])|(~m[759]&m[1278]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[566])|((m[759]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(~m[759]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[759]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[759]&m[1278]&~m[1280]&~m[1281]&m[1282])|(m[759]&~m[1278]&m[1280]&~m[1281]&m[1282])|(~m[759]&~m[1278]&~m[1280]&m[1281]&m[1282])|(m[759]&~m[1278]&~m[1280]&m[1281]&m[1282])|(~m[759]&m[1278]&~m[1280]&m[1281]&m[1282])|(m[759]&m[1278]&~m[1280]&m[1281]&m[1282])|(~m[759]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[759]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[759]&m[1278]&m[1280]&m[1281]&m[1282]));
    m[1284] = (((m[774]&~m[1283]&~m[1285]&~m[1286]&~m[1287])|(~m[774]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(m[774]&m[1283]&~m[1285]&m[1286]&~m[1287])|(m[774]&~m[1283]&m[1285]&m[1286]&~m[1287])|(~m[774]&m[1283]&~m[1285]&~m[1286]&m[1287])|(~m[774]&~m[1283]&m[1285]&~m[1286]&m[1287])|(m[774]&m[1283]&m[1285]&~m[1286]&m[1287])|(~m[774]&m[1283]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[567])|((m[774]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(~m[774]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[774]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[774]&m[1283]&~m[1285]&~m[1286]&m[1287])|(m[774]&~m[1283]&m[1285]&~m[1286]&m[1287])|(~m[774]&~m[1283]&~m[1285]&m[1286]&m[1287])|(m[774]&~m[1283]&~m[1285]&m[1286]&m[1287])|(~m[774]&m[1283]&~m[1285]&m[1286]&m[1287])|(m[774]&m[1283]&~m[1285]&m[1286]&m[1287])|(~m[774]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[774]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[774]&m[1283]&m[1285]&m[1286]&m[1287]));
    m[1289] = (((m[789]&~m[1288]&~m[1290]&~m[1291]&~m[1292])|(~m[789]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(m[789]&m[1288]&~m[1290]&m[1291]&~m[1292])|(m[789]&~m[1288]&m[1290]&m[1291]&~m[1292])|(~m[789]&m[1288]&~m[1290]&~m[1291]&m[1292])|(~m[789]&~m[1288]&m[1290]&~m[1291]&m[1292])|(m[789]&m[1288]&m[1290]&~m[1291]&m[1292])|(~m[789]&m[1288]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[568])|((m[789]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(~m[789]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[789]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[789]&m[1288]&~m[1290]&~m[1291]&m[1292])|(m[789]&~m[1288]&m[1290]&~m[1291]&m[1292])|(~m[789]&~m[1288]&~m[1290]&m[1291]&m[1292])|(m[789]&~m[1288]&~m[1290]&m[1291]&m[1292])|(~m[789]&m[1288]&~m[1290]&m[1291]&m[1292])|(m[789]&m[1288]&~m[1290]&m[1291]&m[1292])|(~m[789]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[789]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[789]&m[1288]&m[1290]&m[1291]&m[1292]));
    m[1294] = (((m[804]&~m[1293]&~m[1295]&~m[1296]&~m[1297])|(~m[804]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(m[804]&m[1293]&~m[1295]&m[1296]&~m[1297])|(m[804]&~m[1293]&m[1295]&m[1296]&~m[1297])|(~m[804]&m[1293]&~m[1295]&~m[1296]&m[1297])|(~m[804]&~m[1293]&m[1295]&~m[1296]&m[1297])|(m[804]&m[1293]&m[1295]&~m[1296]&m[1297])|(~m[804]&m[1293]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[569])|((m[804]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(~m[804]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[804]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[804]&m[1293]&~m[1295]&~m[1296]&m[1297])|(m[804]&~m[1293]&m[1295]&~m[1296]&m[1297])|(~m[804]&~m[1293]&~m[1295]&m[1296]&m[1297])|(m[804]&~m[1293]&~m[1295]&m[1296]&m[1297])|(~m[804]&m[1293]&~m[1295]&m[1296]&m[1297])|(m[804]&m[1293]&~m[1295]&m[1296]&m[1297])|(~m[804]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[804]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[804]&m[1293]&m[1295]&m[1296]&m[1297]));
    m[1299] = (((m[819]&~m[1298]&~m[1300]&~m[1301]&~m[1302])|(~m[819]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(m[819]&m[1298]&~m[1300]&m[1301]&~m[1302])|(m[819]&~m[1298]&m[1300]&m[1301]&~m[1302])|(~m[819]&m[1298]&~m[1300]&~m[1301]&m[1302])|(~m[819]&~m[1298]&m[1300]&~m[1301]&m[1302])|(m[819]&m[1298]&m[1300]&~m[1301]&m[1302])|(~m[819]&m[1298]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[570])|((m[819]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(~m[819]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[819]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[819]&m[1298]&~m[1300]&~m[1301]&m[1302])|(m[819]&~m[1298]&m[1300]&~m[1301]&m[1302])|(~m[819]&~m[1298]&~m[1300]&m[1301]&m[1302])|(m[819]&~m[1298]&~m[1300]&m[1301]&m[1302])|(~m[819]&m[1298]&~m[1300]&m[1301]&m[1302])|(m[819]&m[1298]&~m[1300]&m[1301]&m[1302])|(~m[819]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[819]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[819]&m[1298]&m[1300]&m[1301]&m[1302]));
    m[1304] = (((m[834]&~m[1303]&~m[1305]&~m[1306]&~m[1307])|(~m[834]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(m[834]&m[1303]&~m[1305]&m[1306]&~m[1307])|(m[834]&~m[1303]&m[1305]&m[1306]&~m[1307])|(~m[834]&m[1303]&~m[1305]&~m[1306]&m[1307])|(~m[834]&~m[1303]&m[1305]&~m[1306]&m[1307])|(m[834]&m[1303]&m[1305]&~m[1306]&m[1307])|(~m[834]&m[1303]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[571])|((m[834]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(~m[834]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[834]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[834]&m[1303]&~m[1305]&~m[1306]&m[1307])|(m[834]&~m[1303]&m[1305]&~m[1306]&m[1307])|(~m[834]&~m[1303]&~m[1305]&m[1306]&m[1307])|(m[834]&~m[1303]&~m[1305]&m[1306]&m[1307])|(~m[834]&m[1303]&~m[1305]&m[1306]&m[1307])|(m[834]&m[1303]&~m[1305]&m[1306]&m[1307])|(~m[834]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[834]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[834]&m[1303]&m[1305]&m[1306]&m[1307]));
    m[1309] = (((m[849]&~m[1308]&~m[1310]&~m[1311]&~m[1312])|(~m[849]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(m[849]&m[1308]&~m[1310]&m[1311]&~m[1312])|(m[849]&~m[1308]&m[1310]&m[1311]&~m[1312])|(~m[849]&m[1308]&~m[1310]&~m[1311]&m[1312])|(~m[849]&~m[1308]&m[1310]&~m[1311]&m[1312])|(m[849]&m[1308]&m[1310]&~m[1311]&m[1312])|(~m[849]&m[1308]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[572])|((m[849]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(~m[849]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[849]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[849]&m[1308]&~m[1310]&~m[1311]&m[1312])|(m[849]&~m[1308]&m[1310]&~m[1311]&m[1312])|(~m[849]&~m[1308]&~m[1310]&m[1311]&m[1312])|(m[849]&~m[1308]&~m[1310]&m[1311]&m[1312])|(~m[849]&m[1308]&~m[1310]&m[1311]&m[1312])|(m[849]&m[1308]&~m[1310]&m[1311]&m[1312])|(~m[849]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[849]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[849]&m[1308]&m[1310]&m[1311]&m[1312]));
    m[1314] = (((m[864]&~m[1313]&~m[1315]&~m[1316]&~m[1317])|(~m[864]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(m[864]&m[1313]&~m[1315]&m[1316]&~m[1317])|(m[864]&~m[1313]&m[1315]&m[1316]&~m[1317])|(~m[864]&m[1313]&~m[1315]&~m[1316]&m[1317])|(~m[864]&~m[1313]&m[1315]&~m[1316]&m[1317])|(m[864]&m[1313]&m[1315]&~m[1316]&m[1317])|(~m[864]&m[1313]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[573])|((m[864]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(~m[864]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[864]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[864]&m[1313]&~m[1315]&~m[1316]&m[1317])|(m[864]&~m[1313]&m[1315]&~m[1316]&m[1317])|(~m[864]&~m[1313]&~m[1315]&m[1316]&m[1317])|(m[864]&~m[1313]&~m[1315]&m[1316]&m[1317])|(~m[864]&m[1313]&~m[1315]&m[1316]&m[1317])|(m[864]&m[1313]&~m[1315]&m[1316]&m[1317])|(~m[864]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[864]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[864]&m[1313]&m[1315]&m[1316]&m[1317]));
    m[1319] = (((m[700]&~m[1318]&~m[1320]&~m[1321]&~m[1322])|(~m[700]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(m[700]&m[1318]&~m[1320]&m[1321]&~m[1322])|(m[700]&~m[1318]&m[1320]&m[1321]&~m[1322])|(~m[700]&m[1318]&~m[1320]&~m[1321]&m[1322])|(~m[700]&~m[1318]&m[1320]&~m[1321]&m[1322])|(m[700]&m[1318]&m[1320]&~m[1321]&m[1322])|(~m[700]&m[1318]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[574])|((m[700]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(~m[700]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[700]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[700]&m[1318]&~m[1320]&~m[1321]&m[1322])|(m[700]&~m[1318]&m[1320]&~m[1321]&m[1322])|(~m[700]&~m[1318]&~m[1320]&m[1321]&m[1322])|(m[700]&~m[1318]&~m[1320]&m[1321]&m[1322])|(~m[700]&m[1318]&~m[1320]&m[1321]&m[1322])|(m[700]&m[1318]&~m[1320]&m[1321]&m[1322])|(~m[700]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[700]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[700]&m[1318]&m[1320]&m[1321]&m[1322]));
    m[1324] = (((m[715]&~m[1323]&~m[1325]&~m[1326]&~m[1327])|(~m[715]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(m[715]&m[1323]&~m[1325]&m[1326]&~m[1327])|(m[715]&~m[1323]&m[1325]&m[1326]&~m[1327])|(~m[715]&m[1323]&~m[1325]&~m[1326]&m[1327])|(~m[715]&~m[1323]&m[1325]&~m[1326]&m[1327])|(m[715]&m[1323]&m[1325]&~m[1326]&m[1327])|(~m[715]&m[1323]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[575])|((m[715]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(~m[715]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[715]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[715]&m[1323]&~m[1325]&~m[1326]&m[1327])|(m[715]&~m[1323]&m[1325]&~m[1326]&m[1327])|(~m[715]&~m[1323]&~m[1325]&m[1326]&m[1327])|(m[715]&~m[1323]&~m[1325]&m[1326]&m[1327])|(~m[715]&m[1323]&~m[1325]&m[1326]&m[1327])|(m[715]&m[1323]&~m[1325]&m[1326]&m[1327])|(~m[715]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[715]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[715]&m[1323]&m[1325]&m[1326]&m[1327]));
    m[1329] = (((m[730]&~m[1328]&~m[1330]&~m[1331]&~m[1332])|(~m[730]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(m[730]&m[1328]&~m[1330]&m[1331]&~m[1332])|(m[730]&~m[1328]&m[1330]&m[1331]&~m[1332])|(~m[730]&m[1328]&~m[1330]&~m[1331]&m[1332])|(~m[730]&~m[1328]&m[1330]&~m[1331]&m[1332])|(m[730]&m[1328]&m[1330]&~m[1331]&m[1332])|(~m[730]&m[1328]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[576])|((m[730]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(~m[730]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[730]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[730]&m[1328]&~m[1330]&~m[1331]&m[1332])|(m[730]&~m[1328]&m[1330]&~m[1331]&m[1332])|(~m[730]&~m[1328]&~m[1330]&m[1331]&m[1332])|(m[730]&~m[1328]&~m[1330]&m[1331]&m[1332])|(~m[730]&m[1328]&~m[1330]&m[1331]&m[1332])|(m[730]&m[1328]&~m[1330]&m[1331]&m[1332])|(~m[730]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[730]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[730]&m[1328]&m[1330]&m[1331]&m[1332]));
    m[1334] = (((m[745]&~m[1333]&~m[1335]&~m[1336]&~m[1337])|(~m[745]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(m[745]&m[1333]&~m[1335]&m[1336]&~m[1337])|(m[745]&~m[1333]&m[1335]&m[1336]&~m[1337])|(~m[745]&m[1333]&~m[1335]&~m[1336]&m[1337])|(~m[745]&~m[1333]&m[1335]&~m[1336]&m[1337])|(m[745]&m[1333]&m[1335]&~m[1336]&m[1337])|(~m[745]&m[1333]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[577])|((m[745]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(~m[745]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[745]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[745]&m[1333]&~m[1335]&~m[1336]&m[1337])|(m[745]&~m[1333]&m[1335]&~m[1336]&m[1337])|(~m[745]&~m[1333]&~m[1335]&m[1336]&m[1337])|(m[745]&~m[1333]&~m[1335]&m[1336]&m[1337])|(~m[745]&m[1333]&~m[1335]&m[1336]&m[1337])|(m[745]&m[1333]&~m[1335]&m[1336]&m[1337])|(~m[745]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[745]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[745]&m[1333]&m[1335]&m[1336]&m[1337]));
    m[1339] = (((m[760]&~m[1338]&~m[1340]&~m[1341]&~m[1342])|(~m[760]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(m[760]&m[1338]&~m[1340]&m[1341]&~m[1342])|(m[760]&~m[1338]&m[1340]&m[1341]&~m[1342])|(~m[760]&m[1338]&~m[1340]&~m[1341]&m[1342])|(~m[760]&~m[1338]&m[1340]&~m[1341]&m[1342])|(m[760]&m[1338]&m[1340]&~m[1341]&m[1342])|(~m[760]&m[1338]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[578])|((m[760]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(~m[760]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[760]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[760]&m[1338]&~m[1340]&~m[1341]&m[1342])|(m[760]&~m[1338]&m[1340]&~m[1341]&m[1342])|(~m[760]&~m[1338]&~m[1340]&m[1341]&m[1342])|(m[760]&~m[1338]&~m[1340]&m[1341]&m[1342])|(~m[760]&m[1338]&~m[1340]&m[1341]&m[1342])|(m[760]&m[1338]&~m[1340]&m[1341]&m[1342])|(~m[760]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[760]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[760]&m[1338]&m[1340]&m[1341]&m[1342]));
    m[1344] = (((m[775]&~m[1343]&~m[1345]&~m[1346]&~m[1347])|(~m[775]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(m[775]&m[1343]&~m[1345]&m[1346]&~m[1347])|(m[775]&~m[1343]&m[1345]&m[1346]&~m[1347])|(~m[775]&m[1343]&~m[1345]&~m[1346]&m[1347])|(~m[775]&~m[1343]&m[1345]&~m[1346]&m[1347])|(m[775]&m[1343]&m[1345]&~m[1346]&m[1347])|(~m[775]&m[1343]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[579])|((m[775]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(~m[775]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[775]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[775]&m[1343]&~m[1345]&~m[1346]&m[1347])|(m[775]&~m[1343]&m[1345]&~m[1346]&m[1347])|(~m[775]&~m[1343]&~m[1345]&m[1346]&m[1347])|(m[775]&~m[1343]&~m[1345]&m[1346]&m[1347])|(~m[775]&m[1343]&~m[1345]&m[1346]&m[1347])|(m[775]&m[1343]&~m[1345]&m[1346]&m[1347])|(~m[775]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[775]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[775]&m[1343]&m[1345]&m[1346]&m[1347]));
    m[1349] = (((m[790]&~m[1348]&~m[1350]&~m[1351]&~m[1352])|(~m[790]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(m[790]&m[1348]&~m[1350]&m[1351]&~m[1352])|(m[790]&~m[1348]&m[1350]&m[1351]&~m[1352])|(~m[790]&m[1348]&~m[1350]&~m[1351]&m[1352])|(~m[790]&~m[1348]&m[1350]&~m[1351]&m[1352])|(m[790]&m[1348]&m[1350]&~m[1351]&m[1352])|(~m[790]&m[1348]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[580])|((m[790]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(~m[790]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[790]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[790]&m[1348]&~m[1350]&~m[1351]&m[1352])|(m[790]&~m[1348]&m[1350]&~m[1351]&m[1352])|(~m[790]&~m[1348]&~m[1350]&m[1351]&m[1352])|(m[790]&~m[1348]&~m[1350]&m[1351]&m[1352])|(~m[790]&m[1348]&~m[1350]&m[1351]&m[1352])|(m[790]&m[1348]&~m[1350]&m[1351]&m[1352])|(~m[790]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[790]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[790]&m[1348]&m[1350]&m[1351]&m[1352]));
    m[1354] = (((m[805]&~m[1353]&~m[1355]&~m[1356]&~m[1357])|(~m[805]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(m[805]&m[1353]&~m[1355]&m[1356]&~m[1357])|(m[805]&~m[1353]&m[1355]&m[1356]&~m[1357])|(~m[805]&m[1353]&~m[1355]&~m[1356]&m[1357])|(~m[805]&~m[1353]&m[1355]&~m[1356]&m[1357])|(m[805]&m[1353]&m[1355]&~m[1356]&m[1357])|(~m[805]&m[1353]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[581])|((m[805]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(~m[805]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[805]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[805]&m[1353]&~m[1355]&~m[1356]&m[1357])|(m[805]&~m[1353]&m[1355]&~m[1356]&m[1357])|(~m[805]&~m[1353]&~m[1355]&m[1356]&m[1357])|(m[805]&~m[1353]&~m[1355]&m[1356]&m[1357])|(~m[805]&m[1353]&~m[1355]&m[1356]&m[1357])|(m[805]&m[1353]&~m[1355]&m[1356]&m[1357])|(~m[805]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[805]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[805]&m[1353]&m[1355]&m[1356]&m[1357]));
    m[1359] = (((m[820]&~m[1358]&~m[1360]&~m[1361]&~m[1362])|(~m[820]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(m[820]&m[1358]&~m[1360]&m[1361]&~m[1362])|(m[820]&~m[1358]&m[1360]&m[1361]&~m[1362])|(~m[820]&m[1358]&~m[1360]&~m[1361]&m[1362])|(~m[820]&~m[1358]&m[1360]&~m[1361]&m[1362])|(m[820]&m[1358]&m[1360]&~m[1361]&m[1362])|(~m[820]&m[1358]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[582])|((m[820]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(~m[820]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[820]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[820]&m[1358]&~m[1360]&~m[1361]&m[1362])|(m[820]&~m[1358]&m[1360]&~m[1361]&m[1362])|(~m[820]&~m[1358]&~m[1360]&m[1361]&m[1362])|(m[820]&~m[1358]&~m[1360]&m[1361]&m[1362])|(~m[820]&m[1358]&~m[1360]&m[1361]&m[1362])|(m[820]&m[1358]&~m[1360]&m[1361]&m[1362])|(~m[820]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[820]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[820]&m[1358]&m[1360]&m[1361]&m[1362]));
    m[1364] = (((m[835]&~m[1363]&~m[1365]&~m[1366]&~m[1367])|(~m[835]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(m[835]&m[1363]&~m[1365]&m[1366]&~m[1367])|(m[835]&~m[1363]&m[1365]&m[1366]&~m[1367])|(~m[835]&m[1363]&~m[1365]&~m[1366]&m[1367])|(~m[835]&~m[1363]&m[1365]&~m[1366]&m[1367])|(m[835]&m[1363]&m[1365]&~m[1366]&m[1367])|(~m[835]&m[1363]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[583])|((m[835]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(~m[835]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[835]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[835]&m[1363]&~m[1365]&~m[1366]&m[1367])|(m[835]&~m[1363]&m[1365]&~m[1366]&m[1367])|(~m[835]&~m[1363]&~m[1365]&m[1366]&m[1367])|(m[835]&~m[1363]&~m[1365]&m[1366]&m[1367])|(~m[835]&m[1363]&~m[1365]&m[1366]&m[1367])|(m[835]&m[1363]&~m[1365]&m[1366]&m[1367])|(~m[835]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[835]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[835]&m[1363]&m[1365]&m[1366]&m[1367]));
    m[1369] = (((m[850]&~m[1368]&~m[1370]&~m[1371]&~m[1372])|(~m[850]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(m[850]&m[1368]&~m[1370]&m[1371]&~m[1372])|(m[850]&~m[1368]&m[1370]&m[1371]&~m[1372])|(~m[850]&m[1368]&~m[1370]&~m[1371]&m[1372])|(~m[850]&~m[1368]&m[1370]&~m[1371]&m[1372])|(m[850]&m[1368]&m[1370]&~m[1371]&m[1372])|(~m[850]&m[1368]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[584])|((m[850]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(~m[850]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[850]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[850]&m[1368]&~m[1370]&~m[1371]&m[1372])|(m[850]&~m[1368]&m[1370]&~m[1371]&m[1372])|(~m[850]&~m[1368]&~m[1370]&m[1371]&m[1372])|(m[850]&~m[1368]&~m[1370]&m[1371]&m[1372])|(~m[850]&m[1368]&~m[1370]&m[1371]&m[1372])|(m[850]&m[1368]&~m[1370]&m[1371]&m[1372])|(~m[850]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[850]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[850]&m[1368]&m[1370]&m[1371]&m[1372]));
    m[1374] = (((m[865]&~m[1373]&~m[1375]&~m[1376]&~m[1377])|(~m[865]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(m[865]&m[1373]&~m[1375]&m[1376]&~m[1377])|(m[865]&~m[1373]&m[1375]&m[1376]&~m[1377])|(~m[865]&m[1373]&~m[1375]&~m[1376]&m[1377])|(~m[865]&~m[1373]&m[1375]&~m[1376]&m[1377])|(m[865]&m[1373]&m[1375]&~m[1376]&m[1377])|(~m[865]&m[1373]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[585])|((m[865]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(~m[865]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[865]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[865]&m[1373]&~m[1375]&~m[1376]&m[1377])|(m[865]&~m[1373]&m[1375]&~m[1376]&m[1377])|(~m[865]&~m[1373]&~m[1375]&m[1376]&m[1377])|(m[865]&~m[1373]&~m[1375]&m[1376]&m[1377])|(~m[865]&m[1373]&~m[1375]&m[1376]&m[1377])|(m[865]&m[1373]&~m[1375]&m[1376]&m[1377])|(~m[865]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[865]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[865]&m[1373]&m[1375]&m[1376]&m[1377]));
    m[1379] = (((m[880]&~m[1378]&~m[1380]&~m[1381]&~m[1382])|(~m[880]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(m[880]&m[1378]&~m[1380]&m[1381]&~m[1382])|(m[880]&~m[1378]&m[1380]&m[1381]&~m[1382])|(~m[880]&m[1378]&~m[1380]&~m[1381]&m[1382])|(~m[880]&~m[1378]&m[1380]&~m[1381]&m[1382])|(m[880]&m[1378]&m[1380]&~m[1381]&m[1382])|(~m[880]&m[1378]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[586])|((m[880]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(~m[880]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[880]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[880]&m[1378]&~m[1380]&~m[1381]&m[1382])|(m[880]&~m[1378]&m[1380]&~m[1381]&m[1382])|(~m[880]&~m[1378]&~m[1380]&m[1381]&m[1382])|(m[880]&~m[1378]&~m[1380]&m[1381]&m[1382])|(~m[880]&m[1378]&~m[1380]&m[1381]&m[1382])|(m[880]&m[1378]&~m[1380]&m[1381]&m[1382])|(~m[880]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[880]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[880]&m[1378]&m[1380]&m[1381]&m[1382]));
    m[1384] = (((m[701]&~m[1383]&~m[1385]&~m[1386]&~m[1387])|(~m[701]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(m[701]&m[1383]&~m[1385]&m[1386]&~m[1387])|(m[701]&~m[1383]&m[1385]&m[1386]&~m[1387])|(~m[701]&m[1383]&~m[1385]&~m[1386]&m[1387])|(~m[701]&~m[1383]&m[1385]&~m[1386]&m[1387])|(m[701]&m[1383]&m[1385]&~m[1386]&m[1387])|(~m[701]&m[1383]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[587])|((m[701]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(~m[701]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[701]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[701]&m[1383]&~m[1385]&~m[1386]&m[1387])|(m[701]&~m[1383]&m[1385]&~m[1386]&m[1387])|(~m[701]&~m[1383]&~m[1385]&m[1386]&m[1387])|(m[701]&~m[1383]&~m[1385]&m[1386]&m[1387])|(~m[701]&m[1383]&~m[1385]&m[1386]&m[1387])|(m[701]&m[1383]&~m[1385]&m[1386]&m[1387])|(~m[701]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[701]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[701]&m[1383]&m[1385]&m[1386]&m[1387]));
    m[1389] = (((m[716]&~m[1388]&~m[1390]&~m[1391]&~m[1392])|(~m[716]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(m[716]&m[1388]&~m[1390]&m[1391]&~m[1392])|(m[716]&~m[1388]&m[1390]&m[1391]&~m[1392])|(~m[716]&m[1388]&~m[1390]&~m[1391]&m[1392])|(~m[716]&~m[1388]&m[1390]&~m[1391]&m[1392])|(m[716]&m[1388]&m[1390]&~m[1391]&m[1392])|(~m[716]&m[1388]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[588])|((m[716]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(~m[716]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[716]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[716]&m[1388]&~m[1390]&~m[1391]&m[1392])|(m[716]&~m[1388]&m[1390]&~m[1391]&m[1392])|(~m[716]&~m[1388]&~m[1390]&m[1391]&m[1392])|(m[716]&~m[1388]&~m[1390]&m[1391]&m[1392])|(~m[716]&m[1388]&~m[1390]&m[1391]&m[1392])|(m[716]&m[1388]&~m[1390]&m[1391]&m[1392])|(~m[716]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[716]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[716]&m[1388]&m[1390]&m[1391]&m[1392]));
    m[1394] = (((m[731]&~m[1393]&~m[1395]&~m[1396]&~m[1397])|(~m[731]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(m[731]&m[1393]&~m[1395]&m[1396]&~m[1397])|(m[731]&~m[1393]&m[1395]&m[1396]&~m[1397])|(~m[731]&m[1393]&~m[1395]&~m[1396]&m[1397])|(~m[731]&~m[1393]&m[1395]&~m[1396]&m[1397])|(m[731]&m[1393]&m[1395]&~m[1396]&m[1397])|(~m[731]&m[1393]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[589])|((m[731]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(~m[731]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[731]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[731]&m[1393]&~m[1395]&~m[1396]&m[1397])|(m[731]&~m[1393]&m[1395]&~m[1396]&m[1397])|(~m[731]&~m[1393]&~m[1395]&m[1396]&m[1397])|(m[731]&~m[1393]&~m[1395]&m[1396]&m[1397])|(~m[731]&m[1393]&~m[1395]&m[1396]&m[1397])|(m[731]&m[1393]&~m[1395]&m[1396]&m[1397])|(~m[731]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[731]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[731]&m[1393]&m[1395]&m[1396]&m[1397]));
    m[1399] = (((m[746]&~m[1398]&~m[1400]&~m[1401]&~m[1402])|(~m[746]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(m[746]&m[1398]&~m[1400]&m[1401]&~m[1402])|(m[746]&~m[1398]&m[1400]&m[1401]&~m[1402])|(~m[746]&m[1398]&~m[1400]&~m[1401]&m[1402])|(~m[746]&~m[1398]&m[1400]&~m[1401]&m[1402])|(m[746]&m[1398]&m[1400]&~m[1401]&m[1402])|(~m[746]&m[1398]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[590])|((m[746]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(~m[746]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[746]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[746]&m[1398]&~m[1400]&~m[1401]&m[1402])|(m[746]&~m[1398]&m[1400]&~m[1401]&m[1402])|(~m[746]&~m[1398]&~m[1400]&m[1401]&m[1402])|(m[746]&~m[1398]&~m[1400]&m[1401]&m[1402])|(~m[746]&m[1398]&~m[1400]&m[1401]&m[1402])|(m[746]&m[1398]&~m[1400]&m[1401]&m[1402])|(~m[746]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[746]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[746]&m[1398]&m[1400]&m[1401]&m[1402]));
    m[1404] = (((m[761]&~m[1403]&~m[1405]&~m[1406]&~m[1407])|(~m[761]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(m[761]&m[1403]&~m[1405]&m[1406]&~m[1407])|(m[761]&~m[1403]&m[1405]&m[1406]&~m[1407])|(~m[761]&m[1403]&~m[1405]&~m[1406]&m[1407])|(~m[761]&~m[1403]&m[1405]&~m[1406]&m[1407])|(m[761]&m[1403]&m[1405]&~m[1406]&m[1407])|(~m[761]&m[1403]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[591])|((m[761]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(~m[761]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[761]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[761]&m[1403]&~m[1405]&~m[1406]&m[1407])|(m[761]&~m[1403]&m[1405]&~m[1406]&m[1407])|(~m[761]&~m[1403]&~m[1405]&m[1406]&m[1407])|(m[761]&~m[1403]&~m[1405]&m[1406]&m[1407])|(~m[761]&m[1403]&~m[1405]&m[1406]&m[1407])|(m[761]&m[1403]&~m[1405]&m[1406]&m[1407])|(~m[761]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[761]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[761]&m[1403]&m[1405]&m[1406]&m[1407]));
    m[1409] = (((m[776]&~m[1408]&~m[1410]&~m[1411]&~m[1412])|(~m[776]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(m[776]&m[1408]&~m[1410]&m[1411]&~m[1412])|(m[776]&~m[1408]&m[1410]&m[1411]&~m[1412])|(~m[776]&m[1408]&~m[1410]&~m[1411]&m[1412])|(~m[776]&~m[1408]&m[1410]&~m[1411]&m[1412])|(m[776]&m[1408]&m[1410]&~m[1411]&m[1412])|(~m[776]&m[1408]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[592])|((m[776]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(~m[776]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[776]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[776]&m[1408]&~m[1410]&~m[1411]&m[1412])|(m[776]&~m[1408]&m[1410]&~m[1411]&m[1412])|(~m[776]&~m[1408]&~m[1410]&m[1411]&m[1412])|(m[776]&~m[1408]&~m[1410]&m[1411]&m[1412])|(~m[776]&m[1408]&~m[1410]&m[1411]&m[1412])|(m[776]&m[1408]&~m[1410]&m[1411]&m[1412])|(~m[776]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[776]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[776]&m[1408]&m[1410]&m[1411]&m[1412]));
    m[1414] = (((m[791]&~m[1413]&~m[1415]&~m[1416]&~m[1417])|(~m[791]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(m[791]&m[1413]&~m[1415]&m[1416]&~m[1417])|(m[791]&~m[1413]&m[1415]&m[1416]&~m[1417])|(~m[791]&m[1413]&~m[1415]&~m[1416]&m[1417])|(~m[791]&~m[1413]&m[1415]&~m[1416]&m[1417])|(m[791]&m[1413]&m[1415]&~m[1416]&m[1417])|(~m[791]&m[1413]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[593])|((m[791]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(~m[791]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[791]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[791]&m[1413]&~m[1415]&~m[1416]&m[1417])|(m[791]&~m[1413]&m[1415]&~m[1416]&m[1417])|(~m[791]&~m[1413]&~m[1415]&m[1416]&m[1417])|(m[791]&~m[1413]&~m[1415]&m[1416]&m[1417])|(~m[791]&m[1413]&~m[1415]&m[1416]&m[1417])|(m[791]&m[1413]&~m[1415]&m[1416]&m[1417])|(~m[791]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[791]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[791]&m[1413]&m[1415]&m[1416]&m[1417]));
    m[1419] = (((m[806]&~m[1418]&~m[1420]&~m[1421]&~m[1422])|(~m[806]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(m[806]&m[1418]&~m[1420]&m[1421]&~m[1422])|(m[806]&~m[1418]&m[1420]&m[1421]&~m[1422])|(~m[806]&m[1418]&~m[1420]&~m[1421]&m[1422])|(~m[806]&~m[1418]&m[1420]&~m[1421]&m[1422])|(m[806]&m[1418]&m[1420]&~m[1421]&m[1422])|(~m[806]&m[1418]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[594])|((m[806]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(~m[806]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[806]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[806]&m[1418]&~m[1420]&~m[1421]&m[1422])|(m[806]&~m[1418]&m[1420]&~m[1421]&m[1422])|(~m[806]&~m[1418]&~m[1420]&m[1421]&m[1422])|(m[806]&~m[1418]&~m[1420]&m[1421]&m[1422])|(~m[806]&m[1418]&~m[1420]&m[1421]&m[1422])|(m[806]&m[1418]&~m[1420]&m[1421]&m[1422])|(~m[806]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[806]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[806]&m[1418]&m[1420]&m[1421]&m[1422]));
    m[1424] = (((m[821]&~m[1423]&~m[1425]&~m[1426]&~m[1427])|(~m[821]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(m[821]&m[1423]&~m[1425]&m[1426]&~m[1427])|(m[821]&~m[1423]&m[1425]&m[1426]&~m[1427])|(~m[821]&m[1423]&~m[1425]&~m[1426]&m[1427])|(~m[821]&~m[1423]&m[1425]&~m[1426]&m[1427])|(m[821]&m[1423]&m[1425]&~m[1426]&m[1427])|(~m[821]&m[1423]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[595])|((m[821]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(~m[821]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[821]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[821]&m[1423]&~m[1425]&~m[1426]&m[1427])|(m[821]&~m[1423]&m[1425]&~m[1426]&m[1427])|(~m[821]&~m[1423]&~m[1425]&m[1426]&m[1427])|(m[821]&~m[1423]&~m[1425]&m[1426]&m[1427])|(~m[821]&m[1423]&~m[1425]&m[1426]&m[1427])|(m[821]&m[1423]&~m[1425]&m[1426]&m[1427])|(~m[821]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[821]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[821]&m[1423]&m[1425]&m[1426]&m[1427]));
    m[1429] = (((m[836]&~m[1428]&~m[1430]&~m[1431]&~m[1432])|(~m[836]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(m[836]&m[1428]&~m[1430]&m[1431]&~m[1432])|(m[836]&~m[1428]&m[1430]&m[1431]&~m[1432])|(~m[836]&m[1428]&~m[1430]&~m[1431]&m[1432])|(~m[836]&~m[1428]&m[1430]&~m[1431]&m[1432])|(m[836]&m[1428]&m[1430]&~m[1431]&m[1432])|(~m[836]&m[1428]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[596])|((m[836]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(~m[836]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[836]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[836]&m[1428]&~m[1430]&~m[1431]&m[1432])|(m[836]&~m[1428]&m[1430]&~m[1431]&m[1432])|(~m[836]&~m[1428]&~m[1430]&m[1431]&m[1432])|(m[836]&~m[1428]&~m[1430]&m[1431]&m[1432])|(~m[836]&m[1428]&~m[1430]&m[1431]&m[1432])|(m[836]&m[1428]&~m[1430]&m[1431]&m[1432])|(~m[836]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[836]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[836]&m[1428]&m[1430]&m[1431]&m[1432]));
    m[1434] = (((m[851]&~m[1433]&~m[1435]&~m[1436]&~m[1437])|(~m[851]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(m[851]&m[1433]&~m[1435]&m[1436]&~m[1437])|(m[851]&~m[1433]&m[1435]&m[1436]&~m[1437])|(~m[851]&m[1433]&~m[1435]&~m[1436]&m[1437])|(~m[851]&~m[1433]&m[1435]&~m[1436]&m[1437])|(m[851]&m[1433]&m[1435]&~m[1436]&m[1437])|(~m[851]&m[1433]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[597])|((m[851]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(~m[851]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[851]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[851]&m[1433]&~m[1435]&~m[1436]&m[1437])|(m[851]&~m[1433]&m[1435]&~m[1436]&m[1437])|(~m[851]&~m[1433]&~m[1435]&m[1436]&m[1437])|(m[851]&~m[1433]&~m[1435]&m[1436]&m[1437])|(~m[851]&m[1433]&~m[1435]&m[1436]&m[1437])|(m[851]&m[1433]&~m[1435]&m[1436]&m[1437])|(~m[851]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[851]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[851]&m[1433]&m[1435]&m[1436]&m[1437]));
    m[1439] = (((m[866]&~m[1438]&~m[1440]&~m[1441]&~m[1442])|(~m[866]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(m[866]&m[1438]&~m[1440]&m[1441]&~m[1442])|(m[866]&~m[1438]&m[1440]&m[1441]&~m[1442])|(~m[866]&m[1438]&~m[1440]&~m[1441]&m[1442])|(~m[866]&~m[1438]&m[1440]&~m[1441]&m[1442])|(m[866]&m[1438]&m[1440]&~m[1441]&m[1442])|(~m[866]&m[1438]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[598])|((m[866]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(~m[866]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[866]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[866]&m[1438]&~m[1440]&~m[1441]&m[1442])|(m[866]&~m[1438]&m[1440]&~m[1441]&m[1442])|(~m[866]&~m[1438]&~m[1440]&m[1441]&m[1442])|(m[866]&~m[1438]&~m[1440]&m[1441]&m[1442])|(~m[866]&m[1438]&~m[1440]&m[1441]&m[1442])|(m[866]&m[1438]&~m[1440]&m[1441]&m[1442])|(~m[866]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[866]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[866]&m[1438]&m[1440]&m[1441]&m[1442]));
    m[1444] = (((m[881]&~m[1443]&~m[1445]&~m[1446]&~m[1447])|(~m[881]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(m[881]&m[1443]&~m[1445]&m[1446]&~m[1447])|(m[881]&~m[1443]&m[1445]&m[1446]&~m[1447])|(~m[881]&m[1443]&~m[1445]&~m[1446]&m[1447])|(~m[881]&~m[1443]&m[1445]&~m[1446]&m[1447])|(m[881]&m[1443]&m[1445]&~m[1446]&m[1447])|(~m[881]&m[1443]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[599])|((m[881]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(~m[881]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[881]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[881]&m[1443]&~m[1445]&~m[1446]&m[1447])|(m[881]&~m[1443]&m[1445]&~m[1446]&m[1447])|(~m[881]&~m[1443]&~m[1445]&m[1446]&m[1447])|(m[881]&~m[1443]&~m[1445]&m[1446]&m[1447])|(~m[881]&m[1443]&~m[1445]&m[1446]&m[1447])|(m[881]&m[1443]&~m[1445]&m[1446]&m[1447])|(~m[881]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[881]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[881]&m[1443]&m[1445]&m[1446]&m[1447]));
    m[1449] = (((m[896]&~m[1448]&~m[1450]&~m[1451]&~m[1452])|(~m[896]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(m[896]&m[1448]&~m[1450]&m[1451]&~m[1452])|(m[896]&~m[1448]&m[1450]&m[1451]&~m[1452])|(~m[896]&m[1448]&~m[1450]&~m[1451]&m[1452])|(~m[896]&~m[1448]&m[1450]&~m[1451]&m[1452])|(m[896]&m[1448]&m[1450]&~m[1451]&m[1452])|(~m[896]&m[1448]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[600])|((m[896]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(~m[896]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[896]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[896]&m[1448]&~m[1450]&~m[1451]&m[1452])|(m[896]&~m[1448]&m[1450]&~m[1451]&m[1452])|(~m[896]&~m[1448]&~m[1450]&m[1451]&m[1452])|(m[896]&~m[1448]&~m[1450]&m[1451]&m[1452])|(~m[896]&m[1448]&~m[1450]&m[1451]&m[1452])|(m[896]&m[1448]&~m[1450]&m[1451]&m[1452])|(~m[896]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[896]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[896]&m[1448]&m[1450]&m[1451]&m[1452]));
    m[1454] = (((m[702]&~m[1453]&~m[1455]&~m[1456]&~m[1457])|(~m[702]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(m[702]&m[1453]&~m[1455]&m[1456]&~m[1457])|(m[702]&~m[1453]&m[1455]&m[1456]&~m[1457])|(~m[702]&m[1453]&~m[1455]&~m[1456]&m[1457])|(~m[702]&~m[1453]&m[1455]&~m[1456]&m[1457])|(m[702]&m[1453]&m[1455]&~m[1456]&m[1457])|(~m[702]&m[1453]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[601])|((m[702]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(~m[702]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[702]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[702]&m[1453]&~m[1455]&~m[1456]&m[1457])|(m[702]&~m[1453]&m[1455]&~m[1456]&m[1457])|(~m[702]&~m[1453]&~m[1455]&m[1456]&m[1457])|(m[702]&~m[1453]&~m[1455]&m[1456]&m[1457])|(~m[702]&m[1453]&~m[1455]&m[1456]&m[1457])|(m[702]&m[1453]&~m[1455]&m[1456]&m[1457])|(~m[702]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[702]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[702]&m[1453]&m[1455]&m[1456]&m[1457]));
    m[1459] = (((m[717]&~m[1458]&~m[1460]&~m[1461]&~m[1462])|(~m[717]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(m[717]&m[1458]&~m[1460]&m[1461]&~m[1462])|(m[717]&~m[1458]&m[1460]&m[1461]&~m[1462])|(~m[717]&m[1458]&~m[1460]&~m[1461]&m[1462])|(~m[717]&~m[1458]&m[1460]&~m[1461]&m[1462])|(m[717]&m[1458]&m[1460]&~m[1461]&m[1462])|(~m[717]&m[1458]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[602])|((m[717]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(~m[717]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[717]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[717]&m[1458]&~m[1460]&~m[1461]&m[1462])|(m[717]&~m[1458]&m[1460]&~m[1461]&m[1462])|(~m[717]&~m[1458]&~m[1460]&m[1461]&m[1462])|(m[717]&~m[1458]&~m[1460]&m[1461]&m[1462])|(~m[717]&m[1458]&~m[1460]&m[1461]&m[1462])|(m[717]&m[1458]&~m[1460]&m[1461]&m[1462])|(~m[717]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[717]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[717]&m[1458]&m[1460]&m[1461]&m[1462]));
    m[1464] = (((m[732]&~m[1463]&~m[1465]&~m[1466]&~m[1467])|(~m[732]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(m[732]&m[1463]&~m[1465]&m[1466]&~m[1467])|(m[732]&~m[1463]&m[1465]&m[1466]&~m[1467])|(~m[732]&m[1463]&~m[1465]&~m[1466]&m[1467])|(~m[732]&~m[1463]&m[1465]&~m[1466]&m[1467])|(m[732]&m[1463]&m[1465]&~m[1466]&m[1467])|(~m[732]&m[1463]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[603])|((m[732]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(~m[732]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[732]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[732]&m[1463]&~m[1465]&~m[1466]&m[1467])|(m[732]&~m[1463]&m[1465]&~m[1466]&m[1467])|(~m[732]&~m[1463]&~m[1465]&m[1466]&m[1467])|(m[732]&~m[1463]&~m[1465]&m[1466]&m[1467])|(~m[732]&m[1463]&~m[1465]&m[1466]&m[1467])|(m[732]&m[1463]&~m[1465]&m[1466]&m[1467])|(~m[732]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[732]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[732]&m[1463]&m[1465]&m[1466]&m[1467]));
    m[1469] = (((m[747]&~m[1468]&~m[1470]&~m[1471]&~m[1472])|(~m[747]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(m[747]&m[1468]&~m[1470]&m[1471]&~m[1472])|(m[747]&~m[1468]&m[1470]&m[1471]&~m[1472])|(~m[747]&m[1468]&~m[1470]&~m[1471]&m[1472])|(~m[747]&~m[1468]&m[1470]&~m[1471]&m[1472])|(m[747]&m[1468]&m[1470]&~m[1471]&m[1472])|(~m[747]&m[1468]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[604])|((m[747]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(~m[747]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[747]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[747]&m[1468]&~m[1470]&~m[1471]&m[1472])|(m[747]&~m[1468]&m[1470]&~m[1471]&m[1472])|(~m[747]&~m[1468]&~m[1470]&m[1471]&m[1472])|(m[747]&~m[1468]&~m[1470]&m[1471]&m[1472])|(~m[747]&m[1468]&~m[1470]&m[1471]&m[1472])|(m[747]&m[1468]&~m[1470]&m[1471]&m[1472])|(~m[747]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[747]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[747]&m[1468]&m[1470]&m[1471]&m[1472]));
    m[1474] = (((m[762]&~m[1473]&~m[1475]&~m[1476]&~m[1477])|(~m[762]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(m[762]&m[1473]&~m[1475]&m[1476]&~m[1477])|(m[762]&~m[1473]&m[1475]&m[1476]&~m[1477])|(~m[762]&m[1473]&~m[1475]&~m[1476]&m[1477])|(~m[762]&~m[1473]&m[1475]&~m[1476]&m[1477])|(m[762]&m[1473]&m[1475]&~m[1476]&m[1477])|(~m[762]&m[1473]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[605])|((m[762]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(~m[762]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[762]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[762]&m[1473]&~m[1475]&~m[1476]&m[1477])|(m[762]&~m[1473]&m[1475]&~m[1476]&m[1477])|(~m[762]&~m[1473]&~m[1475]&m[1476]&m[1477])|(m[762]&~m[1473]&~m[1475]&m[1476]&m[1477])|(~m[762]&m[1473]&~m[1475]&m[1476]&m[1477])|(m[762]&m[1473]&~m[1475]&m[1476]&m[1477])|(~m[762]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[762]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[762]&m[1473]&m[1475]&m[1476]&m[1477]));
    m[1479] = (((m[777]&~m[1478]&~m[1480]&~m[1481]&~m[1482])|(~m[777]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(m[777]&m[1478]&~m[1480]&m[1481]&~m[1482])|(m[777]&~m[1478]&m[1480]&m[1481]&~m[1482])|(~m[777]&m[1478]&~m[1480]&~m[1481]&m[1482])|(~m[777]&~m[1478]&m[1480]&~m[1481]&m[1482])|(m[777]&m[1478]&m[1480]&~m[1481]&m[1482])|(~m[777]&m[1478]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[606])|((m[777]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(~m[777]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[777]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[777]&m[1478]&~m[1480]&~m[1481]&m[1482])|(m[777]&~m[1478]&m[1480]&~m[1481]&m[1482])|(~m[777]&~m[1478]&~m[1480]&m[1481]&m[1482])|(m[777]&~m[1478]&~m[1480]&m[1481]&m[1482])|(~m[777]&m[1478]&~m[1480]&m[1481]&m[1482])|(m[777]&m[1478]&~m[1480]&m[1481]&m[1482])|(~m[777]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[777]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[777]&m[1478]&m[1480]&m[1481]&m[1482]));
    m[1484] = (((m[792]&~m[1483]&~m[1485]&~m[1486]&~m[1487])|(~m[792]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(m[792]&m[1483]&~m[1485]&m[1486]&~m[1487])|(m[792]&~m[1483]&m[1485]&m[1486]&~m[1487])|(~m[792]&m[1483]&~m[1485]&~m[1486]&m[1487])|(~m[792]&~m[1483]&m[1485]&~m[1486]&m[1487])|(m[792]&m[1483]&m[1485]&~m[1486]&m[1487])|(~m[792]&m[1483]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[607])|((m[792]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(~m[792]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[792]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[792]&m[1483]&~m[1485]&~m[1486]&m[1487])|(m[792]&~m[1483]&m[1485]&~m[1486]&m[1487])|(~m[792]&~m[1483]&~m[1485]&m[1486]&m[1487])|(m[792]&~m[1483]&~m[1485]&m[1486]&m[1487])|(~m[792]&m[1483]&~m[1485]&m[1486]&m[1487])|(m[792]&m[1483]&~m[1485]&m[1486]&m[1487])|(~m[792]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[792]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[792]&m[1483]&m[1485]&m[1486]&m[1487]));
    m[1489] = (((m[807]&~m[1488]&~m[1490]&~m[1491]&~m[1492])|(~m[807]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(m[807]&m[1488]&~m[1490]&m[1491]&~m[1492])|(m[807]&~m[1488]&m[1490]&m[1491]&~m[1492])|(~m[807]&m[1488]&~m[1490]&~m[1491]&m[1492])|(~m[807]&~m[1488]&m[1490]&~m[1491]&m[1492])|(m[807]&m[1488]&m[1490]&~m[1491]&m[1492])|(~m[807]&m[1488]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[608])|((m[807]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(~m[807]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[807]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[807]&m[1488]&~m[1490]&~m[1491]&m[1492])|(m[807]&~m[1488]&m[1490]&~m[1491]&m[1492])|(~m[807]&~m[1488]&~m[1490]&m[1491]&m[1492])|(m[807]&~m[1488]&~m[1490]&m[1491]&m[1492])|(~m[807]&m[1488]&~m[1490]&m[1491]&m[1492])|(m[807]&m[1488]&~m[1490]&m[1491]&m[1492])|(~m[807]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[807]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[807]&m[1488]&m[1490]&m[1491]&m[1492]));
    m[1494] = (((m[822]&~m[1493]&~m[1495]&~m[1496]&~m[1497])|(~m[822]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(m[822]&m[1493]&~m[1495]&m[1496]&~m[1497])|(m[822]&~m[1493]&m[1495]&m[1496]&~m[1497])|(~m[822]&m[1493]&~m[1495]&~m[1496]&m[1497])|(~m[822]&~m[1493]&m[1495]&~m[1496]&m[1497])|(m[822]&m[1493]&m[1495]&~m[1496]&m[1497])|(~m[822]&m[1493]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[609])|((m[822]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(~m[822]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[822]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[822]&m[1493]&~m[1495]&~m[1496]&m[1497])|(m[822]&~m[1493]&m[1495]&~m[1496]&m[1497])|(~m[822]&~m[1493]&~m[1495]&m[1496]&m[1497])|(m[822]&~m[1493]&~m[1495]&m[1496]&m[1497])|(~m[822]&m[1493]&~m[1495]&m[1496]&m[1497])|(m[822]&m[1493]&~m[1495]&m[1496]&m[1497])|(~m[822]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[822]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[822]&m[1493]&m[1495]&m[1496]&m[1497]));
    m[1499] = (((m[837]&~m[1498]&~m[1500]&~m[1501]&~m[1502])|(~m[837]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(m[837]&m[1498]&~m[1500]&m[1501]&~m[1502])|(m[837]&~m[1498]&m[1500]&m[1501]&~m[1502])|(~m[837]&m[1498]&~m[1500]&~m[1501]&m[1502])|(~m[837]&~m[1498]&m[1500]&~m[1501]&m[1502])|(m[837]&m[1498]&m[1500]&~m[1501]&m[1502])|(~m[837]&m[1498]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[610])|((m[837]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(~m[837]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[837]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[837]&m[1498]&~m[1500]&~m[1501]&m[1502])|(m[837]&~m[1498]&m[1500]&~m[1501]&m[1502])|(~m[837]&~m[1498]&~m[1500]&m[1501]&m[1502])|(m[837]&~m[1498]&~m[1500]&m[1501]&m[1502])|(~m[837]&m[1498]&~m[1500]&m[1501]&m[1502])|(m[837]&m[1498]&~m[1500]&m[1501]&m[1502])|(~m[837]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[837]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[837]&m[1498]&m[1500]&m[1501]&m[1502]));
    m[1504] = (((m[852]&~m[1503]&~m[1505]&~m[1506]&~m[1507])|(~m[852]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(m[852]&m[1503]&~m[1505]&m[1506]&~m[1507])|(m[852]&~m[1503]&m[1505]&m[1506]&~m[1507])|(~m[852]&m[1503]&~m[1505]&~m[1506]&m[1507])|(~m[852]&~m[1503]&m[1505]&~m[1506]&m[1507])|(m[852]&m[1503]&m[1505]&~m[1506]&m[1507])|(~m[852]&m[1503]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[611])|((m[852]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(~m[852]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[852]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[852]&m[1503]&~m[1505]&~m[1506]&m[1507])|(m[852]&~m[1503]&m[1505]&~m[1506]&m[1507])|(~m[852]&~m[1503]&~m[1505]&m[1506]&m[1507])|(m[852]&~m[1503]&~m[1505]&m[1506]&m[1507])|(~m[852]&m[1503]&~m[1505]&m[1506]&m[1507])|(m[852]&m[1503]&~m[1505]&m[1506]&m[1507])|(~m[852]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[852]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[852]&m[1503]&m[1505]&m[1506]&m[1507]));
    m[1509] = (((m[867]&~m[1508]&~m[1510]&~m[1511]&~m[1512])|(~m[867]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(m[867]&m[1508]&~m[1510]&m[1511]&~m[1512])|(m[867]&~m[1508]&m[1510]&m[1511]&~m[1512])|(~m[867]&m[1508]&~m[1510]&~m[1511]&m[1512])|(~m[867]&~m[1508]&m[1510]&~m[1511]&m[1512])|(m[867]&m[1508]&m[1510]&~m[1511]&m[1512])|(~m[867]&m[1508]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[612])|((m[867]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(~m[867]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[867]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[867]&m[1508]&~m[1510]&~m[1511]&m[1512])|(m[867]&~m[1508]&m[1510]&~m[1511]&m[1512])|(~m[867]&~m[1508]&~m[1510]&m[1511]&m[1512])|(m[867]&~m[1508]&~m[1510]&m[1511]&m[1512])|(~m[867]&m[1508]&~m[1510]&m[1511]&m[1512])|(m[867]&m[1508]&~m[1510]&m[1511]&m[1512])|(~m[867]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[867]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[867]&m[1508]&m[1510]&m[1511]&m[1512]));
    m[1514] = (((m[882]&~m[1513]&~m[1515]&~m[1516]&~m[1517])|(~m[882]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(m[882]&m[1513]&~m[1515]&m[1516]&~m[1517])|(m[882]&~m[1513]&m[1515]&m[1516]&~m[1517])|(~m[882]&m[1513]&~m[1515]&~m[1516]&m[1517])|(~m[882]&~m[1513]&m[1515]&~m[1516]&m[1517])|(m[882]&m[1513]&m[1515]&~m[1516]&m[1517])|(~m[882]&m[1513]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[613])|((m[882]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(~m[882]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[882]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[882]&m[1513]&~m[1515]&~m[1516]&m[1517])|(m[882]&~m[1513]&m[1515]&~m[1516]&m[1517])|(~m[882]&~m[1513]&~m[1515]&m[1516]&m[1517])|(m[882]&~m[1513]&~m[1515]&m[1516]&m[1517])|(~m[882]&m[1513]&~m[1515]&m[1516]&m[1517])|(m[882]&m[1513]&~m[1515]&m[1516]&m[1517])|(~m[882]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[882]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[882]&m[1513]&m[1515]&m[1516]&m[1517]));
    m[1519] = (((m[897]&~m[1518]&~m[1520]&~m[1521]&~m[1522])|(~m[897]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(m[897]&m[1518]&~m[1520]&m[1521]&~m[1522])|(m[897]&~m[1518]&m[1520]&m[1521]&~m[1522])|(~m[897]&m[1518]&~m[1520]&~m[1521]&m[1522])|(~m[897]&~m[1518]&m[1520]&~m[1521]&m[1522])|(m[897]&m[1518]&m[1520]&~m[1521]&m[1522])|(~m[897]&m[1518]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[614])|((m[897]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(~m[897]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[897]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[897]&m[1518]&~m[1520]&~m[1521]&m[1522])|(m[897]&~m[1518]&m[1520]&~m[1521]&m[1522])|(~m[897]&~m[1518]&~m[1520]&m[1521]&m[1522])|(m[897]&~m[1518]&~m[1520]&m[1521]&m[1522])|(~m[897]&m[1518]&~m[1520]&m[1521]&m[1522])|(m[897]&m[1518]&~m[1520]&m[1521]&m[1522])|(~m[897]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[897]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[897]&m[1518]&m[1520]&m[1521]&m[1522]));
    m[1524] = (((m[912]&~m[1523]&~m[1525]&~m[1526]&~m[1527])|(~m[912]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(m[912]&m[1523]&~m[1525]&m[1526]&~m[1527])|(m[912]&~m[1523]&m[1525]&m[1526]&~m[1527])|(~m[912]&m[1523]&~m[1525]&~m[1526]&m[1527])|(~m[912]&~m[1523]&m[1525]&~m[1526]&m[1527])|(m[912]&m[1523]&m[1525]&~m[1526]&m[1527])|(~m[912]&m[1523]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[615])|((m[912]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(~m[912]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[912]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[912]&m[1523]&~m[1525]&~m[1526]&m[1527])|(m[912]&~m[1523]&m[1525]&~m[1526]&m[1527])|(~m[912]&~m[1523]&~m[1525]&m[1526]&m[1527])|(m[912]&~m[1523]&~m[1525]&m[1526]&m[1527])|(~m[912]&m[1523]&~m[1525]&m[1526]&m[1527])|(m[912]&m[1523]&~m[1525]&m[1526]&m[1527])|(~m[912]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[912]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[912]&m[1523]&m[1525]&m[1526]&m[1527]));
    m[1529] = (((m[703]&~m[1528]&~m[1530]&~m[1531]&~m[1532])|(~m[703]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(m[703]&m[1528]&~m[1530]&m[1531]&~m[1532])|(m[703]&~m[1528]&m[1530]&m[1531]&~m[1532])|(~m[703]&m[1528]&~m[1530]&~m[1531]&m[1532])|(~m[703]&~m[1528]&m[1530]&~m[1531]&m[1532])|(m[703]&m[1528]&m[1530]&~m[1531]&m[1532])|(~m[703]&m[1528]&m[1530]&m[1531]&m[1532]))&UnbiasedRNG[616])|((m[703]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(~m[703]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[703]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[703]&m[1528]&~m[1530]&~m[1531]&m[1532])|(m[703]&~m[1528]&m[1530]&~m[1531]&m[1532])|(~m[703]&~m[1528]&~m[1530]&m[1531]&m[1532])|(m[703]&~m[1528]&~m[1530]&m[1531]&m[1532])|(~m[703]&m[1528]&~m[1530]&m[1531]&m[1532])|(m[703]&m[1528]&~m[1530]&m[1531]&m[1532])|(~m[703]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[703]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[703]&m[1528]&m[1530]&m[1531]&m[1532]));
    m[1534] = (((m[718]&~m[1533]&~m[1535]&~m[1536]&~m[1537])|(~m[718]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(m[718]&m[1533]&~m[1535]&m[1536]&~m[1537])|(m[718]&~m[1533]&m[1535]&m[1536]&~m[1537])|(~m[718]&m[1533]&~m[1535]&~m[1536]&m[1537])|(~m[718]&~m[1533]&m[1535]&~m[1536]&m[1537])|(m[718]&m[1533]&m[1535]&~m[1536]&m[1537])|(~m[718]&m[1533]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[617])|((m[718]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(~m[718]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[718]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[718]&m[1533]&~m[1535]&~m[1536]&m[1537])|(m[718]&~m[1533]&m[1535]&~m[1536]&m[1537])|(~m[718]&~m[1533]&~m[1535]&m[1536]&m[1537])|(m[718]&~m[1533]&~m[1535]&m[1536]&m[1537])|(~m[718]&m[1533]&~m[1535]&m[1536]&m[1537])|(m[718]&m[1533]&~m[1535]&m[1536]&m[1537])|(~m[718]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[718]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[718]&m[1533]&m[1535]&m[1536]&m[1537]));
    m[1539] = (((m[733]&~m[1538]&~m[1540]&~m[1541]&~m[1542])|(~m[733]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(m[733]&m[1538]&~m[1540]&m[1541]&~m[1542])|(m[733]&~m[1538]&m[1540]&m[1541]&~m[1542])|(~m[733]&m[1538]&~m[1540]&~m[1541]&m[1542])|(~m[733]&~m[1538]&m[1540]&~m[1541]&m[1542])|(m[733]&m[1538]&m[1540]&~m[1541]&m[1542])|(~m[733]&m[1538]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[618])|((m[733]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(~m[733]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[733]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[733]&m[1538]&~m[1540]&~m[1541]&m[1542])|(m[733]&~m[1538]&m[1540]&~m[1541]&m[1542])|(~m[733]&~m[1538]&~m[1540]&m[1541]&m[1542])|(m[733]&~m[1538]&~m[1540]&m[1541]&m[1542])|(~m[733]&m[1538]&~m[1540]&m[1541]&m[1542])|(m[733]&m[1538]&~m[1540]&m[1541]&m[1542])|(~m[733]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[733]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[733]&m[1538]&m[1540]&m[1541]&m[1542]));
    m[1544] = (((m[748]&~m[1543]&~m[1545]&~m[1546]&~m[1547])|(~m[748]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(m[748]&m[1543]&~m[1545]&m[1546]&~m[1547])|(m[748]&~m[1543]&m[1545]&m[1546]&~m[1547])|(~m[748]&m[1543]&~m[1545]&~m[1546]&m[1547])|(~m[748]&~m[1543]&m[1545]&~m[1546]&m[1547])|(m[748]&m[1543]&m[1545]&~m[1546]&m[1547])|(~m[748]&m[1543]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[619])|((m[748]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(~m[748]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[748]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[748]&m[1543]&~m[1545]&~m[1546]&m[1547])|(m[748]&~m[1543]&m[1545]&~m[1546]&m[1547])|(~m[748]&~m[1543]&~m[1545]&m[1546]&m[1547])|(m[748]&~m[1543]&~m[1545]&m[1546]&m[1547])|(~m[748]&m[1543]&~m[1545]&m[1546]&m[1547])|(m[748]&m[1543]&~m[1545]&m[1546]&m[1547])|(~m[748]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[748]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[748]&m[1543]&m[1545]&m[1546]&m[1547]));
    m[1549] = (((m[763]&~m[1548]&~m[1550]&~m[1551]&~m[1552])|(~m[763]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(m[763]&m[1548]&~m[1550]&m[1551]&~m[1552])|(m[763]&~m[1548]&m[1550]&m[1551]&~m[1552])|(~m[763]&m[1548]&~m[1550]&~m[1551]&m[1552])|(~m[763]&~m[1548]&m[1550]&~m[1551]&m[1552])|(m[763]&m[1548]&m[1550]&~m[1551]&m[1552])|(~m[763]&m[1548]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[620])|((m[763]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(~m[763]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[763]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[763]&m[1548]&~m[1550]&~m[1551]&m[1552])|(m[763]&~m[1548]&m[1550]&~m[1551]&m[1552])|(~m[763]&~m[1548]&~m[1550]&m[1551]&m[1552])|(m[763]&~m[1548]&~m[1550]&m[1551]&m[1552])|(~m[763]&m[1548]&~m[1550]&m[1551]&m[1552])|(m[763]&m[1548]&~m[1550]&m[1551]&m[1552])|(~m[763]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[763]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[763]&m[1548]&m[1550]&m[1551]&m[1552]));
    m[1554] = (((m[778]&~m[1553]&~m[1555]&~m[1556]&~m[1557])|(~m[778]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(m[778]&m[1553]&~m[1555]&m[1556]&~m[1557])|(m[778]&~m[1553]&m[1555]&m[1556]&~m[1557])|(~m[778]&m[1553]&~m[1555]&~m[1556]&m[1557])|(~m[778]&~m[1553]&m[1555]&~m[1556]&m[1557])|(m[778]&m[1553]&m[1555]&~m[1556]&m[1557])|(~m[778]&m[1553]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[621])|((m[778]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(~m[778]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[778]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[778]&m[1553]&~m[1555]&~m[1556]&m[1557])|(m[778]&~m[1553]&m[1555]&~m[1556]&m[1557])|(~m[778]&~m[1553]&~m[1555]&m[1556]&m[1557])|(m[778]&~m[1553]&~m[1555]&m[1556]&m[1557])|(~m[778]&m[1553]&~m[1555]&m[1556]&m[1557])|(m[778]&m[1553]&~m[1555]&m[1556]&m[1557])|(~m[778]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[778]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[778]&m[1553]&m[1555]&m[1556]&m[1557]));
    m[1559] = (((m[793]&~m[1558]&~m[1560]&~m[1561]&~m[1562])|(~m[793]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(m[793]&m[1558]&~m[1560]&m[1561]&~m[1562])|(m[793]&~m[1558]&m[1560]&m[1561]&~m[1562])|(~m[793]&m[1558]&~m[1560]&~m[1561]&m[1562])|(~m[793]&~m[1558]&m[1560]&~m[1561]&m[1562])|(m[793]&m[1558]&m[1560]&~m[1561]&m[1562])|(~m[793]&m[1558]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[622])|((m[793]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(~m[793]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[793]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[793]&m[1558]&~m[1560]&~m[1561]&m[1562])|(m[793]&~m[1558]&m[1560]&~m[1561]&m[1562])|(~m[793]&~m[1558]&~m[1560]&m[1561]&m[1562])|(m[793]&~m[1558]&~m[1560]&m[1561]&m[1562])|(~m[793]&m[1558]&~m[1560]&m[1561]&m[1562])|(m[793]&m[1558]&~m[1560]&m[1561]&m[1562])|(~m[793]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[793]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[793]&m[1558]&m[1560]&m[1561]&m[1562]));
    m[1564] = (((m[808]&~m[1563]&~m[1565]&~m[1566]&~m[1567])|(~m[808]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(m[808]&m[1563]&~m[1565]&m[1566]&~m[1567])|(m[808]&~m[1563]&m[1565]&m[1566]&~m[1567])|(~m[808]&m[1563]&~m[1565]&~m[1566]&m[1567])|(~m[808]&~m[1563]&m[1565]&~m[1566]&m[1567])|(m[808]&m[1563]&m[1565]&~m[1566]&m[1567])|(~m[808]&m[1563]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[623])|((m[808]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(~m[808]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[808]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[808]&m[1563]&~m[1565]&~m[1566]&m[1567])|(m[808]&~m[1563]&m[1565]&~m[1566]&m[1567])|(~m[808]&~m[1563]&~m[1565]&m[1566]&m[1567])|(m[808]&~m[1563]&~m[1565]&m[1566]&m[1567])|(~m[808]&m[1563]&~m[1565]&m[1566]&m[1567])|(m[808]&m[1563]&~m[1565]&m[1566]&m[1567])|(~m[808]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[808]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[808]&m[1563]&m[1565]&m[1566]&m[1567]));
    m[1569] = (((m[823]&~m[1568]&~m[1570]&~m[1571]&~m[1572])|(~m[823]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(m[823]&m[1568]&~m[1570]&m[1571]&~m[1572])|(m[823]&~m[1568]&m[1570]&m[1571]&~m[1572])|(~m[823]&m[1568]&~m[1570]&~m[1571]&m[1572])|(~m[823]&~m[1568]&m[1570]&~m[1571]&m[1572])|(m[823]&m[1568]&m[1570]&~m[1571]&m[1572])|(~m[823]&m[1568]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[624])|((m[823]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(~m[823]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[823]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[823]&m[1568]&~m[1570]&~m[1571]&m[1572])|(m[823]&~m[1568]&m[1570]&~m[1571]&m[1572])|(~m[823]&~m[1568]&~m[1570]&m[1571]&m[1572])|(m[823]&~m[1568]&~m[1570]&m[1571]&m[1572])|(~m[823]&m[1568]&~m[1570]&m[1571]&m[1572])|(m[823]&m[1568]&~m[1570]&m[1571]&m[1572])|(~m[823]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[823]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[823]&m[1568]&m[1570]&m[1571]&m[1572]));
    m[1574] = (((m[838]&~m[1573]&~m[1575]&~m[1576]&~m[1577])|(~m[838]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(m[838]&m[1573]&~m[1575]&m[1576]&~m[1577])|(m[838]&~m[1573]&m[1575]&m[1576]&~m[1577])|(~m[838]&m[1573]&~m[1575]&~m[1576]&m[1577])|(~m[838]&~m[1573]&m[1575]&~m[1576]&m[1577])|(m[838]&m[1573]&m[1575]&~m[1576]&m[1577])|(~m[838]&m[1573]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[625])|((m[838]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(~m[838]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[838]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[838]&m[1573]&~m[1575]&~m[1576]&m[1577])|(m[838]&~m[1573]&m[1575]&~m[1576]&m[1577])|(~m[838]&~m[1573]&~m[1575]&m[1576]&m[1577])|(m[838]&~m[1573]&~m[1575]&m[1576]&m[1577])|(~m[838]&m[1573]&~m[1575]&m[1576]&m[1577])|(m[838]&m[1573]&~m[1575]&m[1576]&m[1577])|(~m[838]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[838]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[838]&m[1573]&m[1575]&m[1576]&m[1577]));
    m[1579] = (((m[853]&~m[1578]&~m[1580]&~m[1581]&~m[1582])|(~m[853]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(m[853]&m[1578]&~m[1580]&m[1581]&~m[1582])|(m[853]&~m[1578]&m[1580]&m[1581]&~m[1582])|(~m[853]&m[1578]&~m[1580]&~m[1581]&m[1582])|(~m[853]&~m[1578]&m[1580]&~m[1581]&m[1582])|(m[853]&m[1578]&m[1580]&~m[1581]&m[1582])|(~m[853]&m[1578]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[626])|((m[853]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(~m[853]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[853]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[853]&m[1578]&~m[1580]&~m[1581]&m[1582])|(m[853]&~m[1578]&m[1580]&~m[1581]&m[1582])|(~m[853]&~m[1578]&~m[1580]&m[1581]&m[1582])|(m[853]&~m[1578]&~m[1580]&m[1581]&m[1582])|(~m[853]&m[1578]&~m[1580]&m[1581]&m[1582])|(m[853]&m[1578]&~m[1580]&m[1581]&m[1582])|(~m[853]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[853]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[853]&m[1578]&m[1580]&m[1581]&m[1582]));
    m[1584] = (((m[868]&~m[1583]&~m[1585]&~m[1586]&~m[1587])|(~m[868]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(m[868]&m[1583]&~m[1585]&m[1586]&~m[1587])|(m[868]&~m[1583]&m[1585]&m[1586]&~m[1587])|(~m[868]&m[1583]&~m[1585]&~m[1586]&m[1587])|(~m[868]&~m[1583]&m[1585]&~m[1586]&m[1587])|(m[868]&m[1583]&m[1585]&~m[1586]&m[1587])|(~m[868]&m[1583]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[627])|((m[868]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(~m[868]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[868]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[868]&m[1583]&~m[1585]&~m[1586]&m[1587])|(m[868]&~m[1583]&m[1585]&~m[1586]&m[1587])|(~m[868]&~m[1583]&~m[1585]&m[1586]&m[1587])|(m[868]&~m[1583]&~m[1585]&m[1586]&m[1587])|(~m[868]&m[1583]&~m[1585]&m[1586]&m[1587])|(m[868]&m[1583]&~m[1585]&m[1586]&m[1587])|(~m[868]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[868]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[868]&m[1583]&m[1585]&m[1586]&m[1587]));
    m[1589] = (((m[883]&~m[1588]&~m[1590]&~m[1591]&~m[1592])|(~m[883]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(m[883]&m[1588]&~m[1590]&m[1591]&~m[1592])|(m[883]&~m[1588]&m[1590]&m[1591]&~m[1592])|(~m[883]&m[1588]&~m[1590]&~m[1591]&m[1592])|(~m[883]&~m[1588]&m[1590]&~m[1591]&m[1592])|(m[883]&m[1588]&m[1590]&~m[1591]&m[1592])|(~m[883]&m[1588]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[628])|((m[883]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(~m[883]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[883]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[883]&m[1588]&~m[1590]&~m[1591]&m[1592])|(m[883]&~m[1588]&m[1590]&~m[1591]&m[1592])|(~m[883]&~m[1588]&~m[1590]&m[1591]&m[1592])|(m[883]&~m[1588]&~m[1590]&m[1591]&m[1592])|(~m[883]&m[1588]&~m[1590]&m[1591]&m[1592])|(m[883]&m[1588]&~m[1590]&m[1591]&m[1592])|(~m[883]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[883]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[883]&m[1588]&m[1590]&m[1591]&m[1592]));
    m[1594] = (((m[898]&~m[1593]&~m[1595]&~m[1596]&~m[1597])|(~m[898]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(m[898]&m[1593]&~m[1595]&m[1596]&~m[1597])|(m[898]&~m[1593]&m[1595]&m[1596]&~m[1597])|(~m[898]&m[1593]&~m[1595]&~m[1596]&m[1597])|(~m[898]&~m[1593]&m[1595]&~m[1596]&m[1597])|(m[898]&m[1593]&m[1595]&~m[1596]&m[1597])|(~m[898]&m[1593]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[629])|((m[898]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(~m[898]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[898]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[898]&m[1593]&~m[1595]&~m[1596]&m[1597])|(m[898]&~m[1593]&m[1595]&~m[1596]&m[1597])|(~m[898]&~m[1593]&~m[1595]&m[1596]&m[1597])|(m[898]&~m[1593]&~m[1595]&m[1596]&m[1597])|(~m[898]&m[1593]&~m[1595]&m[1596]&m[1597])|(m[898]&m[1593]&~m[1595]&m[1596]&m[1597])|(~m[898]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[898]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[898]&m[1593]&m[1595]&m[1596]&m[1597]));
    m[1599] = (((m[913]&~m[1598]&~m[1600]&~m[1601]&~m[1602])|(~m[913]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(m[913]&m[1598]&~m[1600]&m[1601]&~m[1602])|(m[913]&~m[1598]&m[1600]&m[1601]&~m[1602])|(~m[913]&m[1598]&~m[1600]&~m[1601]&m[1602])|(~m[913]&~m[1598]&m[1600]&~m[1601]&m[1602])|(m[913]&m[1598]&m[1600]&~m[1601]&m[1602])|(~m[913]&m[1598]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[630])|((m[913]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(~m[913]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[913]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[913]&m[1598]&~m[1600]&~m[1601]&m[1602])|(m[913]&~m[1598]&m[1600]&~m[1601]&m[1602])|(~m[913]&~m[1598]&~m[1600]&m[1601]&m[1602])|(m[913]&~m[1598]&~m[1600]&m[1601]&m[1602])|(~m[913]&m[1598]&~m[1600]&m[1601]&m[1602])|(m[913]&m[1598]&~m[1600]&m[1601]&m[1602])|(~m[913]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[913]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[913]&m[1598]&m[1600]&m[1601]&m[1602]));
    m[1604] = (((m[719]&~m[1603]&~m[1605]&~m[1606]&~m[1607])|(~m[719]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(m[719]&m[1603]&~m[1605]&m[1606]&~m[1607])|(m[719]&~m[1603]&m[1605]&m[1606]&~m[1607])|(~m[719]&m[1603]&~m[1605]&~m[1606]&m[1607])|(~m[719]&~m[1603]&m[1605]&~m[1606]&m[1607])|(m[719]&m[1603]&m[1605]&~m[1606]&m[1607])|(~m[719]&m[1603]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[631])|((m[719]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(~m[719]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[719]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[719]&m[1603]&~m[1605]&~m[1606]&m[1607])|(m[719]&~m[1603]&m[1605]&~m[1606]&m[1607])|(~m[719]&~m[1603]&~m[1605]&m[1606]&m[1607])|(m[719]&~m[1603]&~m[1605]&m[1606]&m[1607])|(~m[719]&m[1603]&~m[1605]&m[1606]&m[1607])|(m[719]&m[1603]&~m[1605]&m[1606]&m[1607])|(~m[719]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[719]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[719]&m[1603]&m[1605]&m[1606]&m[1607]));
    m[1609] = (((m[734]&~m[1608]&~m[1610]&~m[1611]&~m[1612])|(~m[734]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(m[734]&m[1608]&~m[1610]&m[1611]&~m[1612])|(m[734]&~m[1608]&m[1610]&m[1611]&~m[1612])|(~m[734]&m[1608]&~m[1610]&~m[1611]&m[1612])|(~m[734]&~m[1608]&m[1610]&~m[1611]&m[1612])|(m[734]&m[1608]&m[1610]&~m[1611]&m[1612])|(~m[734]&m[1608]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[632])|((m[734]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(~m[734]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[734]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[734]&m[1608]&~m[1610]&~m[1611]&m[1612])|(m[734]&~m[1608]&m[1610]&~m[1611]&m[1612])|(~m[734]&~m[1608]&~m[1610]&m[1611]&m[1612])|(m[734]&~m[1608]&~m[1610]&m[1611]&m[1612])|(~m[734]&m[1608]&~m[1610]&m[1611]&m[1612])|(m[734]&m[1608]&~m[1610]&m[1611]&m[1612])|(~m[734]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[734]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[734]&m[1608]&m[1610]&m[1611]&m[1612]));
    m[1614] = (((m[749]&~m[1613]&~m[1615]&~m[1616]&~m[1617])|(~m[749]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(m[749]&m[1613]&~m[1615]&m[1616]&~m[1617])|(m[749]&~m[1613]&m[1615]&m[1616]&~m[1617])|(~m[749]&m[1613]&~m[1615]&~m[1616]&m[1617])|(~m[749]&~m[1613]&m[1615]&~m[1616]&m[1617])|(m[749]&m[1613]&m[1615]&~m[1616]&m[1617])|(~m[749]&m[1613]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[633])|((m[749]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(~m[749]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[749]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[749]&m[1613]&~m[1615]&~m[1616]&m[1617])|(m[749]&~m[1613]&m[1615]&~m[1616]&m[1617])|(~m[749]&~m[1613]&~m[1615]&m[1616]&m[1617])|(m[749]&~m[1613]&~m[1615]&m[1616]&m[1617])|(~m[749]&m[1613]&~m[1615]&m[1616]&m[1617])|(m[749]&m[1613]&~m[1615]&m[1616]&m[1617])|(~m[749]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[749]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[749]&m[1613]&m[1615]&m[1616]&m[1617]));
    m[1619] = (((m[764]&~m[1618]&~m[1620]&~m[1621]&~m[1622])|(~m[764]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(m[764]&m[1618]&~m[1620]&m[1621]&~m[1622])|(m[764]&~m[1618]&m[1620]&m[1621]&~m[1622])|(~m[764]&m[1618]&~m[1620]&~m[1621]&m[1622])|(~m[764]&~m[1618]&m[1620]&~m[1621]&m[1622])|(m[764]&m[1618]&m[1620]&~m[1621]&m[1622])|(~m[764]&m[1618]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[634])|((m[764]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(~m[764]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[764]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[764]&m[1618]&~m[1620]&~m[1621]&m[1622])|(m[764]&~m[1618]&m[1620]&~m[1621]&m[1622])|(~m[764]&~m[1618]&~m[1620]&m[1621]&m[1622])|(m[764]&~m[1618]&~m[1620]&m[1621]&m[1622])|(~m[764]&m[1618]&~m[1620]&m[1621]&m[1622])|(m[764]&m[1618]&~m[1620]&m[1621]&m[1622])|(~m[764]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[764]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[764]&m[1618]&m[1620]&m[1621]&m[1622]));
    m[1624] = (((m[779]&~m[1623]&~m[1625]&~m[1626]&~m[1627])|(~m[779]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(m[779]&m[1623]&~m[1625]&m[1626]&~m[1627])|(m[779]&~m[1623]&m[1625]&m[1626]&~m[1627])|(~m[779]&m[1623]&~m[1625]&~m[1626]&m[1627])|(~m[779]&~m[1623]&m[1625]&~m[1626]&m[1627])|(m[779]&m[1623]&m[1625]&~m[1626]&m[1627])|(~m[779]&m[1623]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[635])|((m[779]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(~m[779]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[779]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[779]&m[1623]&~m[1625]&~m[1626]&m[1627])|(m[779]&~m[1623]&m[1625]&~m[1626]&m[1627])|(~m[779]&~m[1623]&~m[1625]&m[1626]&m[1627])|(m[779]&~m[1623]&~m[1625]&m[1626]&m[1627])|(~m[779]&m[1623]&~m[1625]&m[1626]&m[1627])|(m[779]&m[1623]&~m[1625]&m[1626]&m[1627])|(~m[779]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[779]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[779]&m[1623]&m[1625]&m[1626]&m[1627]));
    m[1629] = (((m[794]&~m[1628]&~m[1630]&~m[1631]&~m[1632])|(~m[794]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(m[794]&m[1628]&~m[1630]&m[1631]&~m[1632])|(m[794]&~m[1628]&m[1630]&m[1631]&~m[1632])|(~m[794]&m[1628]&~m[1630]&~m[1631]&m[1632])|(~m[794]&~m[1628]&m[1630]&~m[1631]&m[1632])|(m[794]&m[1628]&m[1630]&~m[1631]&m[1632])|(~m[794]&m[1628]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[636])|((m[794]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(~m[794]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[794]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[794]&m[1628]&~m[1630]&~m[1631]&m[1632])|(m[794]&~m[1628]&m[1630]&~m[1631]&m[1632])|(~m[794]&~m[1628]&~m[1630]&m[1631]&m[1632])|(m[794]&~m[1628]&~m[1630]&m[1631]&m[1632])|(~m[794]&m[1628]&~m[1630]&m[1631]&m[1632])|(m[794]&m[1628]&~m[1630]&m[1631]&m[1632])|(~m[794]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[794]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[794]&m[1628]&m[1630]&m[1631]&m[1632]));
    m[1634] = (((m[809]&~m[1633]&~m[1635]&~m[1636]&~m[1637])|(~m[809]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(m[809]&m[1633]&~m[1635]&m[1636]&~m[1637])|(m[809]&~m[1633]&m[1635]&m[1636]&~m[1637])|(~m[809]&m[1633]&~m[1635]&~m[1636]&m[1637])|(~m[809]&~m[1633]&m[1635]&~m[1636]&m[1637])|(m[809]&m[1633]&m[1635]&~m[1636]&m[1637])|(~m[809]&m[1633]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[637])|((m[809]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(~m[809]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[809]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[809]&m[1633]&~m[1635]&~m[1636]&m[1637])|(m[809]&~m[1633]&m[1635]&~m[1636]&m[1637])|(~m[809]&~m[1633]&~m[1635]&m[1636]&m[1637])|(m[809]&~m[1633]&~m[1635]&m[1636]&m[1637])|(~m[809]&m[1633]&~m[1635]&m[1636]&m[1637])|(m[809]&m[1633]&~m[1635]&m[1636]&m[1637])|(~m[809]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[809]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[809]&m[1633]&m[1635]&m[1636]&m[1637]));
    m[1639] = (((m[824]&~m[1638]&~m[1640]&~m[1641]&~m[1642])|(~m[824]&~m[1638]&~m[1640]&m[1641]&~m[1642])|(m[824]&m[1638]&~m[1640]&m[1641]&~m[1642])|(m[824]&~m[1638]&m[1640]&m[1641]&~m[1642])|(~m[824]&m[1638]&~m[1640]&~m[1641]&m[1642])|(~m[824]&~m[1638]&m[1640]&~m[1641]&m[1642])|(m[824]&m[1638]&m[1640]&~m[1641]&m[1642])|(~m[824]&m[1638]&m[1640]&m[1641]&m[1642]))&UnbiasedRNG[638])|((m[824]&~m[1638]&~m[1640]&m[1641]&~m[1642])|(~m[824]&~m[1638]&~m[1640]&~m[1641]&m[1642])|(m[824]&~m[1638]&~m[1640]&~m[1641]&m[1642])|(m[824]&m[1638]&~m[1640]&~m[1641]&m[1642])|(m[824]&~m[1638]&m[1640]&~m[1641]&m[1642])|(~m[824]&~m[1638]&~m[1640]&m[1641]&m[1642])|(m[824]&~m[1638]&~m[1640]&m[1641]&m[1642])|(~m[824]&m[1638]&~m[1640]&m[1641]&m[1642])|(m[824]&m[1638]&~m[1640]&m[1641]&m[1642])|(~m[824]&~m[1638]&m[1640]&m[1641]&m[1642])|(m[824]&~m[1638]&m[1640]&m[1641]&m[1642])|(m[824]&m[1638]&m[1640]&m[1641]&m[1642]));
    m[1644] = (((m[839]&~m[1643]&~m[1645]&~m[1646]&~m[1647])|(~m[839]&~m[1643]&~m[1645]&m[1646]&~m[1647])|(m[839]&m[1643]&~m[1645]&m[1646]&~m[1647])|(m[839]&~m[1643]&m[1645]&m[1646]&~m[1647])|(~m[839]&m[1643]&~m[1645]&~m[1646]&m[1647])|(~m[839]&~m[1643]&m[1645]&~m[1646]&m[1647])|(m[839]&m[1643]&m[1645]&~m[1646]&m[1647])|(~m[839]&m[1643]&m[1645]&m[1646]&m[1647]))&UnbiasedRNG[639])|((m[839]&~m[1643]&~m[1645]&m[1646]&~m[1647])|(~m[839]&~m[1643]&~m[1645]&~m[1646]&m[1647])|(m[839]&~m[1643]&~m[1645]&~m[1646]&m[1647])|(m[839]&m[1643]&~m[1645]&~m[1646]&m[1647])|(m[839]&~m[1643]&m[1645]&~m[1646]&m[1647])|(~m[839]&~m[1643]&~m[1645]&m[1646]&m[1647])|(m[839]&~m[1643]&~m[1645]&m[1646]&m[1647])|(~m[839]&m[1643]&~m[1645]&m[1646]&m[1647])|(m[839]&m[1643]&~m[1645]&m[1646]&m[1647])|(~m[839]&~m[1643]&m[1645]&m[1646]&m[1647])|(m[839]&~m[1643]&m[1645]&m[1646]&m[1647])|(m[839]&m[1643]&m[1645]&m[1646]&m[1647]));
    m[1649] = (((m[854]&~m[1648]&~m[1650]&~m[1651]&~m[1652])|(~m[854]&~m[1648]&~m[1650]&m[1651]&~m[1652])|(m[854]&m[1648]&~m[1650]&m[1651]&~m[1652])|(m[854]&~m[1648]&m[1650]&m[1651]&~m[1652])|(~m[854]&m[1648]&~m[1650]&~m[1651]&m[1652])|(~m[854]&~m[1648]&m[1650]&~m[1651]&m[1652])|(m[854]&m[1648]&m[1650]&~m[1651]&m[1652])|(~m[854]&m[1648]&m[1650]&m[1651]&m[1652]))&UnbiasedRNG[640])|((m[854]&~m[1648]&~m[1650]&m[1651]&~m[1652])|(~m[854]&~m[1648]&~m[1650]&~m[1651]&m[1652])|(m[854]&~m[1648]&~m[1650]&~m[1651]&m[1652])|(m[854]&m[1648]&~m[1650]&~m[1651]&m[1652])|(m[854]&~m[1648]&m[1650]&~m[1651]&m[1652])|(~m[854]&~m[1648]&~m[1650]&m[1651]&m[1652])|(m[854]&~m[1648]&~m[1650]&m[1651]&m[1652])|(~m[854]&m[1648]&~m[1650]&m[1651]&m[1652])|(m[854]&m[1648]&~m[1650]&m[1651]&m[1652])|(~m[854]&~m[1648]&m[1650]&m[1651]&m[1652])|(m[854]&~m[1648]&m[1650]&m[1651]&m[1652])|(m[854]&m[1648]&m[1650]&m[1651]&m[1652]));
    m[1654] = (((m[869]&~m[1653]&~m[1655]&~m[1656]&~m[1657])|(~m[869]&~m[1653]&~m[1655]&m[1656]&~m[1657])|(m[869]&m[1653]&~m[1655]&m[1656]&~m[1657])|(m[869]&~m[1653]&m[1655]&m[1656]&~m[1657])|(~m[869]&m[1653]&~m[1655]&~m[1656]&m[1657])|(~m[869]&~m[1653]&m[1655]&~m[1656]&m[1657])|(m[869]&m[1653]&m[1655]&~m[1656]&m[1657])|(~m[869]&m[1653]&m[1655]&m[1656]&m[1657]))&UnbiasedRNG[641])|((m[869]&~m[1653]&~m[1655]&m[1656]&~m[1657])|(~m[869]&~m[1653]&~m[1655]&~m[1656]&m[1657])|(m[869]&~m[1653]&~m[1655]&~m[1656]&m[1657])|(m[869]&m[1653]&~m[1655]&~m[1656]&m[1657])|(m[869]&~m[1653]&m[1655]&~m[1656]&m[1657])|(~m[869]&~m[1653]&~m[1655]&m[1656]&m[1657])|(m[869]&~m[1653]&~m[1655]&m[1656]&m[1657])|(~m[869]&m[1653]&~m[1655]&m[1656]&m[1657])|(m[869]&m[1653]&~m[1655]&m[1656]&m[1657])|(~m[869]&~m[1653]&m[1655]&m[1656]&m[1657])|(m[869]&~m[1653]&m[1655]&m[1656]&m[1657])|(m[869]&m[1653]&m[1655]&m[1656]&m[1657]));
    m[1659] = (((m[884]&~m[1658]&~m[1660]&~m[1661]&~m[1662])|(~m[884]&~m[1658]&~m[1660]&m[1661]&~m[1662])|(m[884]&m[1658]&~m[1660]&m[1661]&~m[1662])|(m[884]&~m[1658]&m[1660]&m[1661]&~m[1662])|(~m[884]&m[1658]&~m[1660]&~m[1661]&m[1662])|(~m[884]&~m[1658]&m[1660]&~m[1661]&m[1662])|(m[884]&m[1658]&m[1660]&~m[1661]&m[1662])|(~m[884]&m[1658]&m[1660]&m[1661]&m[1662]))&UnbiasedRNG[642])|((m[884]&~m[1658]&~m[1660]&m[1661]&~m[1662])|(~m[884]&~m[1658]&~m[1660]&~m[1661]&m[1662])|(m[884]&~m[1658]&~m[1660]&~m[1661]&m[1662])|(m[884]&m[1658]&~m[1660]&~m[1661]&m[1662])|(m[884]&~m[1658]&m[1660]&~m[1661]&m[1662])|(~m[884]&~m[1658]&~m[1660]&m[1661]&m[1662])|(m[884]&~m[1658]&~m[1660]&m[1661]&m[1662])|(~m[884]&m[1658]&~m[1660]&m[1661]&m[1662])|(m[884]&m[1658]&~m[1660]&m[1661]&m[1662])|(~m[884]&~m[1658]&m[1660]&m[1661]&m[1662])|(m[884]&~m[1658]&m[1660]&m[1661]&m[1662])|(m[884]&m[1658]&m[1660]&m[1661]&m[1662]));
    m[1664] = (((m[899]&~m[1663]&~m[1665]&~m[1666]&~m[1667])|(~m[899]&~m[1663]&~m[1665]&m[1666]&~m[1667])|(m[899]&m[1663]&~m[1665]&m[1666]&~m[1667])|(m[899]&~m[1663]&m[1665]&m[1666]&~m[1667])|(~m[899]&m[1663]&~m[1665]&~m[1666]&m[1667])|(~m[899]&~m[1663]&m[1665]&~m[1666]&m[1667])|(m[899]&m[1663]&m[1665]&~m[1666]&m[1667])|(~m[899]&m[1663]&m[1665]&m[1666]&m[1667]))&UnbiasedRNG[643])|((m[899]&~m[1663]&~m[1665]&m[1666]&~m[1667])|(~m[899]&~m[1663]&~m[1665]&~m[1666]&m[1667])|(m[899]&~m[1663]&~m[1665]&~m[1666]&m[1667])|(m[899]&m[1663]&~m[1665]&~m[1666]&m[1667])|(m[899]&~m[1663]&m[1665]&~m[1666]&m[1667])|(~m[899]&~m[1663]&~m[1665]&m[1666]&m[1667])|(m[899]&~m[1663]&~m[1665]&m[1666]&m[1667])|(~m[899]&m[1663]&~m[1665]&m[1666]&m[1667])|(m[899]&m[1663]&~m[1665]&m[1666]&m[1667])|(~m[899]&~m[1663]&m[1665]&m[1666]&m[1667])|(m[899]&~m[1663]&m[1665]&m[1666]&m[1667])|(m[899]&m[1663]&m[1665]&m[1666]&m[1667]));
    m[1669] = (((m[914]&~m[1668]&~m[1670]&~m[1671]&~m[1672])|(~m[914]&~m[1668]&~m[1670]&m[1671]&~m[1672])|(m[914]&m[1668]&~m[1670]&m[1671]&~m[1672])|(m[914]&~m[1668]&m[1670]&m[1671]&~m[1672])|(~m[914]&m[1668]&~m[1670]&~m[1671]&m[1672])|(~m[914]&~m[1668]&m[1670]&~m[1671]&m[1672])|(m[914]&m[1668]&m[1670]&~m[1671]&m[1672])|(~m[914]&m[1668]&m[1670]&m[1671]&m[1672]))&UnbiasedRNG[644])|((m[914]&~m[1668]&~m[1670]&m[1671]&~m[1672])|(~m[914]&~m[1668]&~m[1670]&~m[1671]&m[1672])|(m[914]&~m[1668]&~m[1670]&~m[1671]&m[1672])|(m[914]&m[1668]&~m[1670]&~m[1671]&m[1672])|(m[914]&~m[1668]&m[1670]&~m[1671]&m[1672])|(~m[914]&~m[1668]&~m[1670]&m[1671]&m[1672])|(m[914]&~m[1668]&~m[1670]&m[1671]&m[1672])|(~m[914]&m[1668]&~m[1670]&m[1671]&m[1672])|(m[914]&m[1668]&~m[1670]&m[1671]&m[1672])|(~m[914]&~m[1668]&m[1670]&m[1671]&m[1672])|(m[914]&~m[1668]&m[1670]&m[1671]&m[1672])|(m[914]&m[1668]&m[1670]&m[1671]&m[1672]));
    m[1674] = (((m[735]&~m[1673]&~m[1675]&~m[1676]&~m[1677])|(~m[735]&~m[1673]&~m[1675]&m[1676]&~m[1677])|(m[735]&m[1673]&~m[1675]&m[1676]&~m[1677])|(m[735]&~m[1673]&m[1675]&m[1676]&~m[1677])|(~m[735]&m[1673]&~m[1675]&~m[1676]&m[1677])|(~m[735]&~m[1673]&m[1675]&~m[1676]&m[1677])|(m[735]&m[1673]&m[1675]&~m[1676]&m[1677])|(~m[735]&m[1673]&m[1675]&m[1676]&m[1677]))&UnbiasedRNG[645])|((m[735]&~m[1673]&~m[1675]&m[1676]&~m[1677])|(~m[735]&~m[1673]&~m[1675]&~m[1676]&m[1677])|(m[735]&~m[1673]&~m[1675]&~m[1676]&m[1677])|(m[735]&m[1673]&~m[1675]&~m[1676]&m[1677])|(m[735]&~m[1673]&m[1675]&~m[1676]&m[1677])|(~m[735]&~m[1673]&~m[1675]&m[1676]&m[1677])|(m[735]&~m[1673]&~m[1675]&m[1676]&m[1677])|(~m[735]&m[1673]&~m[1675]&m[1676]&m[1677])|(m[735]&m[1673]&~m[1675]&m[1676]&m[1677])|(~m[735]&~m[1673]&m[1675]&m[1676]&m[1677])|(m[735]&~m[1673]&m[1675]&m[1676]&m[1677])|(m[735]&m[1673]&m[1675]&m[1676]&m[1677]));
    m[1679] = (((m[750]&~m[1678]&~m[1680]&~m[1681]&~m[1682])|(~m[750]&~m[1678]&~m[1680]&m[1681]&~m[1682])|(m[750]&m[1678]&~m[1680]&m[1681]&~m[1682])|(m[750]&~m[1678]&m[1680]&m[1681]&~m[1682])|(~m[750]&m[1678]&~m[1680]&~m[1681]&m[1682])|(~m[750]&~m[1678]&m[1680]&~m[1681]&m[1682])|(m[750]&m[1678]&m[1680]&~m[1681]&m[1682])|(~m[750]&m[1678]&m[1680]&m[1681]&m[1682]))&UnbiasedRNG[646])|((m[750]&~m[1678]&~m[1680]&m[1681]&~m[1682])|(~m[750]&~m[1678]&~m[1680]&~m[1681]&m[1682])|(m[750]&~m[1678]&~m[1680]&~m[1681]&m[1682])|(m[750]&m[1678]&~m[1680]&~m[1681]&m[1682])|(m[750]&~m[1678]&m[1680]&~m[1681]&m[1682])|(~m[750]&~m[1678]&~m[1680]&m[1681]&m[1682])|(m[750]&~m[1678]&~m[1680]&m[1681]&m[1682])|(~m[750]&m[1678]&~m[1680]&m[1681]&m[1682])|(m[750]&m[1678]&~m[1680]&m[1681]&m[1682])|(~m[750]&~m[1678]&m[1680]&m[1681]&m[1682])|(m[750]&~m[1678]&m[1680]&m[1681]&m[1682])|(m[750]&m[1678]&m[1680]&m[1681]&m[1682]));
    m[1684] = (((m[765]&~m[1683]&~m[1685]&~m[1686]&~m[1687])|(~m[765]&~m[1683]&~m[1685]&m[1686]&~m[1687])|(m[765]&m[1683]&~m[1685]&m[1686]&~m[1687])|(m[765]&~m[1683]&m[1685]&m[1686]&~m[1687])|(~m[765]&m[1683]&~m[1685]&~m[1686]&m[1687])|(~m[765]&~m[1683]&m[1685]&~m[1686]&m[1687])|(m[765]&m[1683]&m[1685]&~m[1686]&m[1687])|(~m[765]&m[1683]&m[1685]&m[1686]&m[1687]))&UnbiasedRNG[647])|((m[765]&~m[1683]&~m[1685]&m[1686]&~m[1687])|(~m[765]&~m[1683]&~m[1685]&~m[1686]&m[1687])|(m[765]&~m[1683]&~m[1685]&~m[1686]&m[1687])|(m[765]&m[1683]&~m[1685]&~m[1686]&m[1687])|(m[765]&~m[1683]&m[1685]&~m[1686]&m[1687])|(~m[765]&~m[1683]&~m[1685]&m[1686]&m[1687])|(m[765]&~m[1683]&~m[1685]&m[1686]&m[1687])|(~m[765]&m[1683]&~m[1685]&m[1686]&m[1687])|(m[765]&m[1683]&~m[1685]&m[1686]&m[1687])|(~m[765]&~m[1683]&m[1685]&m[1686]&m[1687])|(m[765]&~m[1683]&m[1685]&m[1686]&m[1687])|(m[765]&m[1683]&m[1685]&m[1686]&m[1687]));
    m[1689] = (((m[780]&~m[1688]&~m[1690]&~m[1691]&~m[1692])|(~m[780]&~m[1688]&~m[1690]&m[1691]&~m[1692])|(m[780]&m[1688]&~m[1690]&m[1691]&~m[1692])|(m[780]&~m[1688]&m[1690]&m[1691]&~m[1692])|(~m[780]&m[1688]&~m[1690]&~m[1691]&m[1692])|(~m[780]&~m[1688]&m[1690]&~m[1691]&m[1692])|(m[780]&m[1688]&m[1690]&~m[1691]&m[1692])|(~m[780]&m[1688]&m[1690]&m[1691]&m[1692]))&UnbiasedRNG[648])|((m[780]&~m[1688]&~m[1690]&m[1691]&~m[1692])|(~m[780]&~m[1688]&~m[1690]&~m[1691]&m[1692])|(m[780]&~m[1688]&~m[1690]&~m[1691]&m[1692])|(m[780]&m[1688]&~m[1690]&~m[1691]&m[1692])|(m[780]&~m[1688]&m[1690]&~m[1691]&m[1692])|(~m[780]&~m[1688]&~m[1690]&m[1691]&m[1692])|(m[780]&~m[1688]&~m[1690]&m[1691]&m[1692])|(~m[780]&m[1688]&~m[1690]&m[1691]&m[1692])|(m[780]&m[1688]&~m[1690]&m[1691]&m[1692])|(~m[780]&~m[1688]&m[1690]&m[1691]&m[1692])|(m[780]&~m[1688]&m[1690]&m[1691]&m[1692])|(m[780]&m[1688]&m[1690]&m[1691]&m[1692]));
    m[1694] = (((m[795]&~m[1693]&~m[1695]&~m[1696]&~m[1697])|(~m[795]&~m[1693]&~m[1695]&m[1696]&~m[1697])|(m[795]&m[1693]&~m[1695]&m[1696]&~m[1697])|(m[795]&~m[1693]&m[1695]&m[1696]&~m[1697])|(~m[795]&m[1693]&~m[1695]&~m[1696]&m[1697])|(~m[795]&~m[1693]&m[1695]&~m[1696]&m[1697])|(m[795]&m[1693]&m[1695]&~m[1696]&m[1697])|(~m[795]&m[1693]&m[1695]&m[1696]&m[1697]))&UnbiasedRNG[649])|((m[795]&~m[1693]&~m[1695]&m[1696]&~m[1697])|(~m[795]&~m[1693]&~m[1695]&~m[1696]&m[1697])|(m[795]&~m[1693]&~m[1695]&~m[1696]&m[1697])|(m[795]&m[1693]&~m[1695]&~m[1696]&m[1697])|(m[795]&~m[1693]&m[1695]&~m[1696]&m[1697])|(~m[795]&~m[1693]&~m[1695]&m[1696]&m[1697])|(m[795]&~m[1693]&~m[1695]&m[1696]&m[1697])|(~m[795]&m[1693]&~m[1695]&m[1696]&m[1697])|(m[795]&m[1693]&~m[1695]&m[1696]&m[1697])|(~m[795]&~m[1693]&m[1695]&m[1696]&m[1697])|(m[795]&~m[1693]&m[1695]&m[1696]&m[1697])|(m[795]&m[1693]&m[1695]&m[1696]&m[1697]));
    m[1699] = (((m[810]&~m[1698]&~m[1700]&~m[1701]&~m[1702])|(~m[810]&~m[1698]&~m[1700]&m[1701]&~m[1702])|(m[810]&m[1698]&~m[1700]&m[1701]&~m[1702])|(m[810]&~m[1698]&m[1700]&m[1701]&~m[1702])|(~m[810]&m[1698]&~m[1700]&~m[1701]&m[1702])|(~m[810]&~m[1698]&m[1700]&~m[1701]&m[1702])|(m[810]&m[1698]&m[1700]&~m[1701]&m[1702])|(~m[810]&m[1698]&m[1700]&m[1701]&m[1702]))&UnbiasedRNG[650])|((m[810]&~m[1698]&~m[1700]&m[1701]&~m[1702])|(~m[810]&~m[1698]&~m[1700]&~m[1701]&m[1702])|(m[810]&~m[1698]&~m[1700]&~m[1701]&m[1702])|(m[810]&m[1698]&~m[1700]&~m[1701]&m[1702])|(m[810]&~m[1698]&m[1700]&~m[1701]&m[1702])|(~m[810]&~m[1698]&~m[1700]&m[1701]&m[1702])|(m[810]&~m[1698]&~m[1700]&m[1701]&m[1702])|(~m[810]&m[1698]&~m[1700]&m[1701]&m[1702])|(m[810]&m[1698]&~m[1700]&m[1701]&m[1702])|(~m[810]&~m[1698]&m[1700]&m[1701]&m[1702])|(m[810]&~m[1698]&m[1700]&m[1701]&m[1702])|(m[810]&m[1698]&m[1700]&m[1701]&m[1702]));
    m[1704] = (((m[825]&~m[1703]&~m[1705]&~m[1706]&~m[1707])|(~m[825]&~m[1703]&~m[1705]&m[1706]&~m[1707])|(m[825]&m[1703]&~m[1705]&m[1706]&~m[1707])|(m[825]&~m[1703]&m[1705]&m[1706]&~m[1707])|(~m[825]&m[1703]&~m[1705]&~m[1706]&m[1707])|(~m[825]&~m[1703]&m[1705]&~m[1706]&m[1707])|(m[825]&m[1703]&m[1705]&~m[1706]&m[1707])|(~m[825]&m[1703]&m[1705]&m[1706]&m[1707]))&UnbiasedRNG[651])|((m[825]&~m[1703]&~m[1705]&m[1706]&~m[1707])|(~m[825]&~m[1703]&~m[1705]&~m[1706]&m[1707])|(m[825]&~m[1703]&~m[1705]&~m[1706]&m[1707])|(m[825]&m[1703]&~m[1705]&~m[1706]&m[1707])|(m[825]&~m[1703]&m[1705]&~m[1706]&m[1707])|(~m[825]&~m[1703]&~m[1705]&m[1706]&m[1707])|(m[825]&~m[1703]&~m[1705]&m[1706]&m[1707])|(~m[825]&m[1703]&~m[1705]&m[1706]&m[1707])|(m[825]&m[1703]&~m[1705]&m[1706]&m[1707])|(~m[825]&~m[1703]&m[1705]&m[1706]&m[1707])|(m[825]&~m[1703]&m[1705]&m[1706]&m[1707])|(m[825]&m[1703]&m[1705]&m[1706]&m[1707]));
    m[1709] = (((m[840]&~m[1708]&~m[1710]&~m[1711]&~m[1712])|(~m[840]&~m[1708]&~m[1710]&m[1711]&~m[1712])|(m[840]&m[1708]&~m[1710]&m[1711]&~m[1712])|(m[840]&~m[1708]&m[1710]&m[1711]&~m[1712])|(~m[840]&m[1708]&~m[1710]&~m[1711]&m[1712])|(~m[840]&~m[1708]&m[1710]&~m[1711]&m[1712])|(m[840]&m[1708]&m[1710]&~m[1711]&m[1712])|(~m[840]&m[1708]&m[1710]&m[1711]&m[1712]))&UnbiasedRNG[652])|((m[840]&~m[1708]&~m[1710]&m[1711]&~m[1712])|(~m[840]&~m[1708]&~m[1710]&~m[1711]&m[1712])|(m[840]&~m[1708]&~m[1710]&~m[1711]&m[1712])|(m[840]&m[1708]&~m[1710]&~m[1711]&m[1712])|(m[840]&~m[1708]&m[1710]&~m[1711]&m[1712])|(~m[840]&~m[1708]&~m[1710]&m[1711]&m[1712])|(m[840]&~m[1708]&~m[1710]&m[1711]&m[1712])|(~m[840]&m[1708]&~m[1710]&m[1711]&m[1712])|(m[840]&m[1708]&~m[1710]&m[1711]&m[1712])|(~m[840]&~m[1708]&m[1710]&m[1711]&m[1712])|(m[840]&~m[1708]&m[1710]&m[1711]&m[1712])|(m[840]&m[1708]&m[1710]&m[1711]&m[1712]));
    m[1714] = (((m[855]&~m[1713]&~m[1715]&~m[1716]&~m[1717])|(~m[855]&~m[1713]&~m[1715]&m[1716]&~m[1717])|(m[855]&m[1713]&~m[1715]&m[1716]&~m[1717])|(m[855]&~m[1713]&m[1715]&m[1716]&~m[1717])|(~m[855]&m[1713]&~m[1715]&~m[1716]&m[1717])|(~m[855]&~m[1713]&m[1715]&~m[1716]&m[1717])|(m[855]&m[1713]&m[1715]&~m[1716]&m[1717])|(~m[855]&m[1713]&m[1715]&m[1716]&m[1717]))&UnbiasedRNG[653])|((m[855]&~m[1713]&~m[1715]&m[1716]&~m[1717])|(~m[855]&~m[1713]&~m[1715]&~m[1716]&m[1717])|(m[855]&~m[1713]&~m[1715]&~m[1716]&m[1717])|(m[855]&m[1713]&~m[1715]&~m[1716]&m[1717])|(m[855]&~m[1713]&m[1715]&~m[1716]&m[1717])|(~m[855]&~m[1713]&~m[1715]&m[1716]&m[1717])|(m[855]&~m[1713]&~m[1715]&m[1716]&m[1717])|(~m[855]&m[1713]&~m[1715]&m[1716]&m[1717])|(m[855]&m[1713]&~m[1715]&m[1716]&m[1717])|(~m[855]&~m[1713]&m[1715]&m[1716]&m[1717])|(m[855]&~m[1713]&m[1715]&m[1716]&m[1717])|(m[855]&m[1713]&m[1715]&m[1716]&m[1717]));
    m[1719] = (((m[870]&~m[1718]&~m[1720]&~m[1721]&~m[1722])|(~m[870]&~m[1718]&~m[1720]&m[1721]&~m[1722])|(m[870]&m[1718]&~m[1720]&m[1721]&~m[1722])|(m[870]&~m[1718]&m[1720]&m[1721]&~m[1722])|(~m[870]&m[1718]&~m[1720]&~m[1721]&m[1722])|(~m[870]&~m[1718]&m[1720]&~m[1721]&m[1722])|(m[870]&m[1718]&m[1720]&~m[1721]&m[1722])|(~m[870]&m[1718]&m[1720]&m[1721]&m[1722]))&UnbiasedRNG[654])|((m[870]&~m[1718]&~m[1720]&m[1721]&~m[1722])|(~m[870]&~m[1718]&~m[1720]&~m[1721]&m[1722])|(m[870]&~m[1718]&~m[1720]&~m[1721]&m[1722])|(m[870]&m[1718]&~m[1720]&~m[1721]&m[1722])|(m[870]&~m[1718]&m[1720]&~m[1721]&m[1722])|(~m[870]&~m[1718]&~m[1720]&m[1721]&m[1722])|(m[870]&~m[1718]&~m[1720]&m[1721]&m[1722])|(~m[870]&m[1718]&~m[1720]&m[1721]&m[1722])|(m[870]&m[1718]&~m[1720]&m[1721]&m[1722])|(~m[870]&~m[1718]&m[1720]&m[1721]&m[1722])|(m[870]&~m[1718]&m[1720]&m[1721]&m[1722])|(m[870]&m[1718]&m[1720]&m[1721]&m[1722]));
    m[1724] = (((m[885]&~m[1723]&~m[1725]&~m[1726]&~m[1727])|(~m[885]&~m[1723]&~m[1725]&m[1726]&~m[1727])|(m[885]&m[1723]&~m[1725]&m[1726]&~m[1727])|(m[885]&~m[1723]&m[1725]&m[1726]&~m[1727])|(~m[885]&m[1723]&~m[1725]&~m[1726]&m[1727])|(~m[885]&~m[1723]&m[1725]&~m[1726]&m[1727])|(m[885]&m[1723]&m[1725]&~m[1726]&m[1727])|(~m[885]&m[1723]&m[1725]&m[1726]&m[1727]))&UnbiasedRNG[655])|((m[885]&~m[1723]&~m[1725]&m[1726]&~m[1727])|(~m[885]&~m[1723]&~m[1725]&~m[1726]&m[1727])|(m[885]&~m[1723]&~m[1725]&~m[1726]&m[1727])|(m[885]&m[1723]&~m[1725]&~m[1726]&m[1727])|(m[885]&~m[1723]&m[1725]&~m[1726]&m[1727])|(~m[885]&~m[1723]&~m[1725]&m[1726]&m[1727])|(m[885]&~m[1723]&~m[1725]&m[1726]&m[1727])|(~m[885]&m[1723]&~m[1725]&m[1726]&m[1727])|(m[885]&m[1723]&~m[1725]&m[1726]&m[1727])|(~m[885]&~m[1723]&m[1725]&m[1726]&m[1727])|(m[885]&~m[1723]&m[1725]&m[1726]&m[1727])|(m[885]&m[1723]&m[1725]&m[1726]&m[1727]));
    m[1729] = (((m[900]&~m[1728]&~m[1730]&~m[1731]&~m[1732])|(~m[900]&~m[1728]&~m[1730]&m[1731]&~m[1732])|(m[900]&m[1728]&~m[1730]&m[1731]&~m[1732])|(m[900]&~m[1728]&m[1730]&m[1731]&~m[1732])|(~m[900]&m[1728]&~m[1730]&~m[1731]&m[1732])|(~m[900]&~m[1728]&m[1730]&~m[1731]&m[1732])|(m[900]&m[1728]&m[1730]&~m[1731]&m[1732])|(~m[900]&m[1728]&m[1730]&m[1731]&m[1732]))&UnbiasedRNG[656])|((m[900]&~m[1728]&~m[1730]&m[1731]&~m[1732])|(~m[900]&~m[1728]&~m[1730]&~m[1731]&m[1732])|(m[900]&~m[1728]&~m[1730]&~m[1731]&m[1732])|(m[900]&m[1728]&~m[1730]&~m[1731]&m[1732])|(m[900]&~m[1728]&m[1730]&~m[1731]&m[1732])|(~m[900]&~m[1728]&~m[1730]&m[1731]&m[1732])|(m[900]&~m[1728]&~m[1730]&m[1731]&m[1732])|(~m[900]&m[1728]&~m[1730]&m[1731]&m[1732])|(m[900]&m[1728]&~m[1730]&m[1731]&m[1732])|(~m[900]&~m[1728]&m[1730]&m[1731]&m[1732])|(m[900]&~m[1728]&m[1730]&m[1731]&m[1732])|(m[900]&m[1728]&m[1730]&m[1731]&m[1732]));
    m[1734] = (((m[915]&~m[1733]&~m[1735]&~m[1736]&~m[1737])|(~m[915]&~m[1733]&~m[1735]&m[1736]&~m[1737])|(m[915]&m[1733]&~m[1735]&m[1736]&~m[1737])|(m[915]&~m[1733]&m[1735]&m[1736]&~m[1737])|(~m[915]&m[1733]&~m[1735]&~m[1736]&m[1737])|(~m[915]&~m[1733]&m[1735]&~m[1736]&m[1737])|(m[915]&m[1733]&m[1735]&~m[1736]&m[1737])|(~m[915]&m[1733]&m[1735]&m[1736]&m[1737]))&UnbiasedRNG[657])|((m[915]&~m[1733]&~m[1735]&m[1736]&~m[1737])|(~m[915]&~m[1733]&~m[1735]&~m[1736]&m[1737])|(m[915]&~m[1733]&~m[1735]&~m[1736]&m[1737])|(m[915]&m[1733]&~m[1735]&~m[1736]&m[1737])|(m[915]&~m[1733]&m[1735]&~m[1736]&m[1737])|(~m[915]&~m[1733]&~m[1735]&m[1736]&m[1737])|(m[915]&~m[1733]&~m[1735]&m[1736]&m[1737])|(~m[915]&m[1733]&~m[1735]&m[1736]&m[1737])|(m[915]&m[1733]&~m[1735]&m[1736]&m[1737])|(~m[915]&~m[1733]&m[1735]&m[1736]&m[1737])|(m[915]&~m[1733]&m[1735]&m[1736]&m[1737])|(m[915]&m[1733]&m[1735]&m[1736]&m[1737]));
    m[1739] = (((m[751]&~m[1738]&~m[1740]&~m[1741]&~m[1742])|(~m[751]&~m[1738]&~m[1740]&m[1741]&~m[1742])|(m[751]&m[1738]&~m[1740]&m[1741]&~m[1742])|(m[751]&~m[1738]&m[1740]&m[1741]&~m[1742])|(~m[751]&m[1738]&~m[1740]&~m[1741]&m[1742])|(~m[751]&~m[1738]&m[1740]&~m[1741]&m[1742])|(m[751]&m[1738]&m[1740]&~m[1741]&m[1742])|(~m[751]&m[1738]&m[1740]&m[1741]&m[1742]))&UnbiasedRNG[658])|((m[751]&~m[1738]&~m[1740]&m[1741]&~m[1742])|(~m[751]&~m[1738]&~m[1740]&~m[1741]&m[1742])|(m[751]&~m[1738]&~m[1740]&~m[1741]&m[1742])|(m[751]&m[1738]&~m[1740]&~m[1741]&m[1742])|(m[751]&~m[1738]&m[1740]&~m[1741]&m[1742])|(~m[751]&~m[1738]&~m[1740]&m[1741]&m[1742])|(m[751]&~m[1738]&~m[1740]&m[1741]&m[1742])|(~m[751]&m[1738]&~m[1740]&m[1741]&m[1742])|(m[751]&m[1738]&~m[1740]&m[1741]&m[1742])|(~m[751]&~m[1738]&m[1740]&m[1741]&m[1742])|(m[751]&~m[1738]&m[1740]&m[1741]&m[1742])|(m[751]&m[1738]&m[1740]&m[1741]&m[1742]));
    m[1744] = (((m[766]&~m[1743]&~m[1745]&~m[1746]&~m[1747])|(~m[766]&~m[1743]&~m[1745]&m[1746]&~m[1747])|(m[766]&m[1743]&~m[1745]&m[1746]&~m[1747])|(m[766]&~m[1743]&m[1745]&m[1746]&~m[1747])|(~m[766]&m[1743]&~m[1745]&~m[1746]&m[1747])|(~m[766]&~m[1743]&m[1745]&~m[1746]&m[1747])|(m[766]&m[1743]&m[1745]&~m[1746]&m[1747])|(~m[766]&m[1743]&m[1745]&m[1746]&m[1747]))&UnbiasedRNG[659])|((m[766]&~m[1743]&~m[1745]&m[1746]&~m[1747])|(~m[766]&~m[1743]&~m[1745]&~m[1746]&m[1747])|(m[766]&~m[1743]&~m[1745]&~m[1746]&m[1747])|(m[766]&m[1743]&~m[1745]&~m[1746]&m[1747])|(m[766]&~m[1743]&m[1745]&~m[1746]&m[1747])|(~m[766]&~m[1743]&~m[1745]&m[1746]&m[1747])|(m[766]&~m[1743]&~m[1745]&m[1746]&m[1747])|(~m[766]&m[1743]&~m[1745]&m[1746]&m[1747])|(m[766]&m[1743]&~m[1745]&m[1746]&m[1747])|(~m[766]&~m[1743]&m[1745]&m[1746]&m[1747])|(m[766]&~m[1743]&m[1745]&m[1746]&m[1747])|(m[766]&m[1743]&m[1745]&m[1746]&m[1747]));
    m[1749] = (((m[781]&~m[1748]&~m[1750]&~m[1751]&~m[1752])|(~m[781]&~m[1748]&~m[1750]&m[1751]&~m[1752])|(m[781]&m[1748]&~m[1750]&m[1751]&~m[1752])|(m[781]&~m[1748]&m[1750]&m[1751]&~m[1752])|(~m[781]&m[1748]&~m[1750]&~m[1751]&m[1752])|(~m[781]&~m[1748]&m[1750]&~m[1751]&m[1752])|(m[781]&m[1748]&m[1750]&~m[1751]&m[1752])|(~m[781]&m[1748]&m[1750]&m[1751]&m[1752]))&UnbiasedRNG[660])|((m[781]&~m[1748]&~m[1750]&m[1751]&~m[1752])|(~m[781]&~m[1748]&~m[1750]&~m[1751]&m[1752])|(m[781]&~m[1748]&~m[1750]&~m[1751]&m[1752])|(m[781]&m[1748]&~m[1750]&~m[1751]&m[1752])|(m[781]&~m[1748]&m[1750]&~m[1751]&m[1752])|(~m[781]&~m[1748]&~m[1750]&m[1751]&m[1752])|(m[781]&~m[1748]&~m[1750]&m[1751]&m[1752])|(~m[781]&m[1748]&~m[1750]&m[1751]&m[1752])|(m[781]&m[1748]&~m[1750]&m[1751]&m[1752])|(~m[781]&~m[1748]&m[1750]&m[1751]&m[1752])|(m[781]&~m[1748]&m[1750]&m[1751]&m[1752])|(m[781]&m[1748]&m[1750]&m[1751]&m[1752]));
    m[1754] = (((m[796]&~m[1753]&~m[1755]&~m[1756]&~m[1757])|(~m[796]&~m[1753]&~m[1755]&m[1756]&~m[1757])|(m[796]&m[1753]&~m[1755]&m[1756]&~m[1757])|(m[796]&~m[1753]&m[1755]&m[1756]&~m[1757])|(~m[796]&m[1753]&~m[1755]&~m[1756]&m[1757])|(~m[796]&~m[1753]&m[1755]&~m[1756]&m[1757])|(m[796]&m[1753]&m[1755]&~m[1756]&m[1757])|(~m[796]&m[1753]&m[1755]&m[1756]&m[1757]))&UnbiasedRNG[661])|((m[796]&~m[1753]&~m[1755]&m[1756]&~m[1757])|(~m[796]&~m[1753]&~m[1755]&~m[1756]&m[1757])|(m[796]&~m[1753]&~m[1755]&~m[1756]&m[1757])|(m[796]&m[1753]&~m[1755]&~m[1756]&m[1757])|(m[796]&~m[1753]&m[1755]&~m[1756]&m[1757])|(~m[796]&~m[1753]&~m[1755]&m[1756]&m[1757])|(m[796]&~m[1753]&~m[1755]&m[1756]&m[1757])|(~m[796]&m[1753]&~m[1755]&m[1756]&m[1757])|(m[796]&m[1753]&~m[1755]&m[1756]&m[1757])|(~m[796]&~m[1753]&m[1755]&m[1756]&m[1757])|(m[796]&~m[1753]&m[1755]&m[1756]&m[1757])|(m[796]&m[1753]&m[1755]&m[1756]&m[1757]));
    m[1759] = (((m[811]&~m[1758]&~m[1760]&~m[1761]&~m[1762])|(~m[811]&~m[1758]&~m[1760]&m[1761]&~m[1762])|(m[811]&m[1758]&~m[1760]&m[1761]&~m[1762])|(m[811]&~m[1758]&m[1760]&m[1761]&~m[1762])|(~m[811]&m[1758]&~m[1760]&~m[1761]&m[1762])|(~m[811]&~m[1758]&m[1760]&~m[1761]&m[1762])|(m[811]&m[1758]&m[1760]&~m[1761]&m[1762])|(~m[811]&m[1758]&m[1760]&m[1761]&m[1762]))&UnbiasedRNG[662])|((m[811]&~m[1758]&~m[1760]&m[1761]&~m[1762])|(~m[811]&~m[1758]&~m[1760]&~m[1761]&m[1762])|(m[811]&~m[1758]&~m[1760]&~m[1761]&m[1762])|(m[811]&m[1758]&~m[1760]&~m[1761]&m[1762])|(m[811]&~m[1758]&m[1760]&~m[1761]&m[1762])|(~m[811]&~m[1758]&~m[1760]&m[1761]&m[1762])|(m[811]&~m[1758]&~m[1760]&m[1761]&m[1762])|(~m[811]&m[1758]&~m[1760]&m[1761]&m[1762])|(m[811]&m[1758]&~m[1760]&m[1761]&m[1762])|(~m[811]&~m[1758]&m[1760]&m[1761]&m[1762])|(m[811]&~m[1758]&m[1760]&m[1761]&m[1762])|(m[811]&m[1758]&m[1760]&m[1761]&m[1762]));
    m[1764] = (((m[826]&~m[1763]&~m[1765]&~m[1766]&~m[1767])|(~m[826]&~m[1763]&~m[1765]&m[1766]&~m[1767])|(m[826]&m[1763]&~m[1765]&m[1766]&~m[1767])|(m[826]&~m[1763]&m[1765]&m[1766]&~m[1767])|(~m[826]&m[1763]&~m[1765]&~m[1766]&m[1767])|(~m[826]&~m[1763]&m[1765]&~m[1766]&m[1767])|(m[826]&m[1763]&m[1765]&~m[1766]&m[1767])|(~m[826]&m[1763]&m[1765]&m[1766]&m[1767]))&UnbiasedRNG[663])|((m[826]&~m[1763]&~m[1765]&m[1766]&~m[1767])|(~m[826]&~m[1763]&~m[1765]&~m[1766]&m[1767])|(m[826]&~m[1763]&~m[1765]&~m[1766]&m[1767])|(m[826]&m[1763]&~m[1765]&~m[1766]&m[1767])|(m[826]&~m[1763]&m[1765]&~m[1766]&m[1767])|(~m[826]&~m[1763]&~m[1765]&m[1766]&m[1767])|(m[826]&~m[1763]&~m[1765]&m[1766]&m[1767])|(~m[826]&m[1763]&~m[1765]&m[1766]&m[1767])|(m[826]&m[1763]&~m[1765]&m[1766]&m[1767])|(~m[826]&~m[1763]&m[1765]&m[1766]&m[1767])|(m[826]&~m[1763]&m[1765]&m[1766]&m[1767])|(m[826]&m[1763]&m[1765]&m[1766]&m[1767]));
    m[1769] = (((m[841]&~m[1768]&~m[1770]&~m[1771]&~m[1772])|(~m[841]&~m[1768]&~m[1770]&m[1771]&~m[1772])|(m[841]&m[1768]&~m[1770]&m[1771]&~m[1772])|(m[841]&~m[1768]&m[1770]&m[1771]&~m[1772])|(~m[841]&m[1768]&~m[1770]&~m[1771]&m[1772])|(~m[841]&~m[1768]&m[1770]&~m[1771]&m[1772])|(m[841]&m[1768]&m[1770]&~m[1771]&m[1772])|(~m[841]&m[1768]&m[1770]&m[1771]&m[1772]))&UnbiasedRNG[664])|((m[841]&~m[1768]&~m[1770]&m[1771]&~m[1772])|(~m[841]&~m[1768]&~m[1770]&~m[1771]&m[1772])|(m[841]&~m[1768]&~m[1770]&~m[1771]&m[1772])|(m[841]&m[1768]&~m[1770]&~m[1771]&m[1772])|(m[841]&~m[1768]&m[1770]&~m[1771]&m[1772])|(~m[841]&~m[1768]&~m[1770]&m[1771]&m[1772])|(m[841]&~m[1768]&~m[1770]&m[1771]&m[1772])|(~m[841]&m[1768]&~m[1770]&m[1771]&m[1772])|(m[841]&m[1768]&~m[1770]&m[1771]&m[1772])|(~m[841]&~m[1768]&m[1770]&m[1771]&m[1772])|(m[841]&~m[1768]&m[1770]&m[1771]&m[1772])|(m[841]&m[1768]&m[1770]&m[1771]&m[1772]));
    m[1774] = (((m[856]&~m[1773]&~m[1775]&~m[1776]&~m[1777])|(~m[856]&~m[1773]&~m[1775]&m[1776]&~m[1777])|(m[856]&m[1773]&~m[1775]&m[1776]&~m[1777])|(m[856]&~m[1773]&m[1775]&m[1776]&~m[1777])|(~m[856]&m[1773]&~m[1775]&~m[1776]&m[1777])|(~m[856]&~m[1773]&m[1775]&~m[1776]&m[1777])|(m[856]&m[1773]&m[1775]&~m[1776]&m[1777])|(~m[856]&m[1773]&m[1775]&m[1776]&m[1777]))&UnbiasedRNG[665])|((m[856]&~m[1773]&~m[1775]&m[1776]&~m[1777])|(~m[856]&~m[1773]&~m[1775]&~m[1776]&m[1777])|(m[856]&~m[1773]&~m[1775]&~m[1776]&m[1777])|(m[856]&m[1773]&~m[1775]&~m[1776]&m[1777])|(m[856]&~m[1773]&m[1775]&~m[1776]&m[1777])|(~m[856]&~m[1773]&~m[1775]&m[1776]&m[1777])|(m[856]&~m[1773]&~m[1775]&m[1776]&m[1777])|(~m[856]&m[1773]&~m[1775]&m[1776]&m[1777])|(m[856]&m[1773]&~m[1775]&m[1776]&m[1777])|(~m[856]&~m[1773]&m[1775]&m[1776]&m[1777])|(m[856]&~m[1773]&m[1775]&m[1776]&m[1777])|(m[856]&m[1773]&m[1775]&m[1776]&m[1777]));
    m[1779] = (((m[871]&~m[1778]&~m[1780]&~m[1781]&~m[1782])|(~m[871]&~m[1778]&~m[1780]&m[1781]&~m[1782])|(m[871]&m[1778]&~m[1780]&m[1781]&~m[1782])|(m[871]&~m[1778]&m[1780]&m[1781]&~m[1782])|(~m[871]&m[1778]&~m[1780]&~m[1781]&m[1782])|(~m[871]&~m[1778]&m[1780]&~m[1781]&m[1782])|(m[871]&m[1778]&m[1780]&~m[1781]&m[1782])|(~m[871]&m[1778]&m[1780]&m[1781]&m[1782]))&UnbiasedRNG[666])|((m[871]&~m[1778]&~m[1780]&m[1781]&~m[1782])|(~m[871]&~m[1778]&~m[1780]&~m[1781]&m[1782])|(m[871]&~m[1778]&~m[1780]&~m[1781]&m[1782])|(m[871]&m[1778]&~m[1780]&~m[1781]&m[1782])|(m[871]&~m[1778]&m[1780]&~m[1781]&m[1782])|(~m[871]&~m[1778]&~m[1780]&m[1781]&m[1782])|(m[871]&~m[1778]&~m[1780]&m[1781]&m[1782])|(~m[871]&m[1778]&~m[1780]&m[1781]&m[1782])|(m[871]&m[1778]&~m[1780]&m[1781]&m[1782])|(~m[871]&~m[1778]&m[1780]&m[1781]&m[1782])|(m[871]&~m[1778]&m[1780]&m[1781]&m[1782])|(m[871]&m[1778]&m[1780]&m[1781]&m[1782]));
    m[1784] = (((m[886]&~m[1783]&~m[1785]&~m[1786]&~m[1787])|(~m[886]&~m[1783]&~m[1785]&m[1786]&~m[1787])|(m[886]&m[1783]&~m[1785]&m[1786]&~m[1787])|(m[886]&~m[1783]&m[1785]&m[1786]&~m[1787])|(~m[886]&m[1783]&~m[1785]&~m[1786]&m[1787])|(~m[886]&~m[1783]&m[1785]&~m[1786]&m[1787])|(m[886]&m[1783]&m[1785]&~m[1786]&m[1787])|(~m[886]&m[1783]&m[1785]&m[1786]&m[1787]))&UnbiasedRNG[667])|((m[886]&~m[1783]&~m[1785]&m[1786]&~m[1787])|(~m[886]&~m[1783]&~m[1785]&~m[1786]&m[1787])|(m[886]&~m[1783]&~m[1785]&~m[1786]&m[1787])|(m[886]&m[1783]&~m[1785]&~m[1786]&m[1787])|(m[886]&~m[1783]&m[1785]&~m[1786]&m[1787])|(~m[886]&~m[1783]&~m[1785]&m[1786]&m[1787])|(m[886]&~m[1783]&~m[1785]&m[1786]&m[1787])|(~m[886]&m[1783]&~m[1785]&m[1786]&m[1787])|(m[886]&m[1783]&~m[1785]&m[1786]&m[1787])|(~m[886]&~m[1783]&m[1785]&m[1786]&m[1787])|(m[886]&~m[1783]&m[1785]&m[1786]&m[1787])|(m[886]&m[1783]&m[1785]&m[1786]&m[1787]));
    m[1789] = (((m[901]&~m[1788]&~m[1790]&~m[1791]&~m[1792])|(~m[901]&~m[1788]&~m[1790]&m[1791]&~m[1792])|(m[901]&m[1788]&~m[1790]&m[1791]&~m[1792])|(m[901]&~m[1788]&m[1790]&m[1791]&~m[1792])|(~m[901]&m[1788]&~m[1790]&~m[1791]&m[1792])|(~m[901]&~m[1788]&m[1790]&~m[1791]&m[1792])|(m[901]&m[1788]&m[1790]&~m[1791]&m[1792])|(~m[901]&m[1788]&m[1790]&m[1791]&m[1792]))&UnbiasedRNG[668])|((m[901]&~m[1788]&~m[1790]&m[1791]&~m[1792])|(~m[901]&~m[1788]&~m[1790]&~m[1791]&m[1792])|(m[901]&~m[1788]&~m[1790]&~m[1791]&m[1792])|(m[901]&m[1788]&~m[1790]&~m[1791]&m[1792])|(m[901]&~m[1788]&m[1790]&~m[1791]&m[1792])|(~m[901]&~m[1788]&~m[1790]&m[1791]&m[1792])|(m[901]&~m[1788]&~m[1790]&m[1791]&m[1792])|(~m[901]&m[1788]&~m[1790]&m[1791]&m[1792])|(m[901]&m[1788]&~m[1790]&m[1791]&m[1792])|(~m[901]&~m[1788]&m[1790]&m[1791]&m[1792])|(m[901]&~m[1788]&m[1790]&m[1791]&m[1792])|(m[901]&m[1788]&m[1790]&m[1791]&m[1792]));
    m[1794] = (((m[916]&~m[1793]&~m[1795]&~m[1796]&~m[1797])|(~m[916]&~m[1793]&~m[1795]&m[1796]&~m[1797])|(m[916]&m[1793]&~m[1795]&m[1796]&~m[1797])|(m[916]&~m[1793]&m[1795]&m[1796]&~m[1797])|(~m[916]&m[1793]&~m[1795]&~m[1796]&m[1797])|(~m[916]&~m[1793]&m[1795]&~m[1796]&m[1797])|(m[916]&m[1793]&m[1795]&~m[1796]&m[1797])|(~m[916]&m[1793]&m[1795]&m[1796]&m[1797]))&UnbiasedRNG[669])|((m[916]&~m[1793]&~m[1795]&m[1796]&~m[1797])|(~m[916]&~m[1793]&~m[1795]&~m[1796]&m[1797])|(m[916]&~m[1793]&~m[1795]&~m[1796]&m[1797])|(m[916]&m[1793]&~m[1795]&~m[1796]&m[1797])|(m[916]&~m[1793]&m[1795]&~m[1796]&m[1797])|(~m[916]&~m[1793]&~m[1795]&m[1796]&m[1797])|(m[916]&~m[1793]&~m[1795]&m[1796]&m[1797])|(~m[916]&m[1793]&~m[1795]&m[1796]&m[1797])|(m[916]&m[1793]&~m[1795]&m[1796]&m[1797])|(~m[916]&~m[1793]&m[1795]&m[1796]&m[1797])|(m[916]&~m[1793]&m[1795]&m[1796]&m[1797])|(m[916]&m[1793]&m[1795]&m[1796]&m[1797]));
    m[1799] = (((m[767]&~m[1798]&~m[1800]&~m[1801]&~m[1802])|(~m[767]&~m[1798]&~m[1800]&m[1801]&~m[1802])|(m[767]&m[1798]&~m[1800]&m[1801]&~m[1802])|(m[767]&~m[1798]&m[1800]&m[1801]&~m[1802])|(~m[767]&m[1798]&~m[1800]&~m[1801]&m[1802])|(~m[767]&~m[1798]&m[1800]&~m[1801]&m[1802])|(m[767]&m[1798]&m[1800]&~m[1801]&m[1802])|(~m[767]&m[1798]&m[1800]&m[1801]&m[1802]))&UnbiasedRNG[670])|((m[767]&~m[1798]&~m[1800]&m[1801]&~m[1802])|(~m[767]&~m[1798]&~m[1800]&~m[1801]&m[1802])|(m[767]&~m[1798]&~m[1800]&~m[1801]&m[1802])|(m[767]&m[1798]&~m[1800]&~m[1801]&m[1802])|(m[767]&~m[1798]&m[1800]&~m[1801]&m[1802])|(~m[767]&~m[1798]&~m[1800]&m[1801]&m[1802])|(m[767]&~m[1798]&~m[1800]&m[1801]&m[1802])|(~m[767]&m[1798]&~m[1800]&m[1801]&m[1802])|(m[767]&m[1798]&~m[1800]&m[1801]&m[1802])|(~m[767]&~m[1798]&m[1800]&m[1801]&m[1802])|(m[767]&~m[1798]&m[1800]&m[1801]&m[1802])|(m[767]&m[1798]&m[1800]&m[1801]&m[1802]));
    m[1804] = (((m[782]&~m[1803]&~m[1805]&~m[1806]&~m[1807])|(~m[782]&~m[1803]&~m[1805]&m[1806]&~m[1807])|(m[782]&m[1803]&~m[1805]&m[1806]&~m[1807])|(m[782]&~m[1803]&m[1805]&m[1806]&~m[1807])|(~m[782]&m[1803]&~m[1805]&~m[1806]&m[1807])|(~m[782]&~m[1803]&m[1805]&~m[1806]&m[1807])|(m[782]&m[1803]&m[1805]&~m[1806]&m[1807])|(~m[782]&m[1803]&m[1805]&m[1806]&m[1807]))&UnbiasedRNG[671])|((m[782]&~m[1803]&~m[1805]&m[1806]&~m[1807])|(~m[782]&~m[1803]&~m[1805]&~m[1806]&m[1807])|(m[782]&~m[1803]&~m[1805]&~m[1806]&m[1807])|(m[782]&m[1803]&~m[1805]&~m[1806]&m[1807])|(m[782]&~m[1803]&m[1805]&~m[1806]&m[1807])|(~m[782]&~m[1803]&~m[1805]&m[1806]&m[1807])|(m[782]&~m[1803]&~m[1805]&m[1806]&m[1807])|(~m[782]&m[1803]&~m[1805]&m[1806]&m[1807])|(m[782]&m[1803]&~m[1805]&m[1806]&m[1807])|(~m[782]&~m[1803]&m[1805]&m[1806]&m[1807])|(m[782]&~m[1803]&m[1805]&m[1806]&m[1807])|(m[782]&m[1803]&m[1805]&m[1806]&m[1807]));
    m[1809] = (((m[797]&~m[1808]&~m[1810]&~m[1811]&~m[1812])|(~m[797]&~m[1808]&~m[1810]&m[1811]&~m[1812])|(m[797]&m[1808]&~m[1810]&m[1811]&~m[1812])|(m[797]&~m[1808]&m[1810]&m[1811]&~m[1812])|(~m[797]&m[1808]&~m[1810]&~m[1811]&m[1812])|(~m[797]&~m[1808]&m[1810]&~m[1811]&m[1812])|(m[797]&m[1808]&m[1810]&~m[1811]&m[1812])|(~m[797]&m[1808]&m[1810]&m[1811]&m[1812]))&UnbiasedRNG[672])|((m[797]&~m[1808]&~m[1810]&m[1811]&~m[1812])|(~m[797]&~m[1808]&~m[1810]&~m[1811]&m[1812])|(m[797]&~m[1808]&~m[1810]&~m[1811]&m[1812])|(m[797]&m[1808]&~m[1810]&~m[1811]&m[1812])|(m[797]&~m[1808]&m[1810]&~m[1811]&m[1812])|(~m[797]&~m[1808]&~m[1810]&m[1811]&m[1812])|(m[797]&~m[1808]&~m[1810]&m[1811]&m[1812])|(~m[797]&m[1808]&~m[1810]&m[1811]&m[1812])|(m[797]&m[1808]&~m[1810]&m[1811]&m[1812])|(~m[797]&~m[1808]&m[1810]&m[1811]&m[1812])|(m[797]&~m[1808]&m[1810]&m[1811]&m[1812])|(m[797]&m[1808]&m[1810]&m[1811]&m[1812]));
    m[1814] = (((m[812]&~m[1813]&~m[1815]&~m[1816]&~m[1817])|(~m[812]&~m[1813]&~m[1815]&m[1816]&~m[1817])|(m[812]&m[1813]&~m[1815]&m[1816]&~m[1817])|(m[812]&~m[1813]&m[1815]&m[1816]&~m[1817])|(~m[812]&m[1813]&~m[1815]&~m[1816]&m[1817])|(~m[812]&~m[1813]&m[1815]&~m[1816]&m[1817])|(m[812]&m[1813]&m[1815]&~m[1816]&m[1817])|(~m[812]&m[1813]&m[1815]&m[1816]&m[1817]))&UnbiasedRNG[673])|((m[812]&~m[1813]&~m[1815]&m[1816]&~m[1817])|(~m[812]&~m[1813]&~m[1815]&~m[1816]&m[1817])|(m[812]&~m[1813]&~m[1815]&~m[1816]&m[1817])|(m[812]&m[1813]&~m[1815]&~m[1816]&m[1817])|(m[812]&~m[1813]&m[1815]&~m[1816]&m[1817])|(~m[812]&~m[1813]&~m[1815]&m[1816]&m[1817])|(m[812]&~m[1813]&~m[1815]&m[1816]&m[1817])|(~m[812]&m[1813]&~m[1815]&m[1816]&m[1817])|(m[812]&m[1813]&~m[1815]&m[1816]&m[1817])|(~m[812]&~m[1813]&m[1815]&m[1816]&m[1817])|(m[812]&~m[1813]&m[1815]&m[1816]&m[1817])|(m[812]&m[1813]&m[1815]&m[1816]&m[1817]));
    m[1819] = (((m[827]&~m[1818]&~m[1820]&~m[1821]&~m[1822])|(~m[827]&~m[1818]&~m[1820]&m[1821]&~m[1822])|(m[827]&m[1818]&~m[1820]&m[1821]&~m[1822])|(m[827]&~m[1818]&m[1820]&m[1821]&~m[1822])|(~m[827]&m[1818]&~m[1820]&~m[1821]&m[1822])|(~m[827]&~m[1818]&m[1820]&~m[1821]&m[1822])|(m[827]&m[1818]&m[1820]&~m[1821]&m[1822])|(~m[827]&m[1818]&m[1820]&m[1821]&m[1822]))&UnbiasedRNG[674])|((m[827]&~m[1818]&~m[1820]&m[1821]&~m[1822])|(~m[827]&~m[1818]&~m[1820]&~m[1821]&m[1822])|(m[827]&~m[1818]&~m[1820]&~m[1821]&m[1822])|(m[827]&m[1818]&~m[1820]&~m[1821]&m[1822])|(m[827]&~m[1818]&m[1820]&~m[1821]&m[1822])|(~m[827]&~m[1818]&~m[1820]&m[1821]&m[1822])|(m[827]&~m[1818]&~m[1820]&m[1821]&m[1822])|(~m[827]&m[1818]&~m[1820]&m[1821]&m[1822])|(m[827]&m[1818]&~m[1820]&m[1821]&m[1822])|(~m[827]&~m[1818]&m[1820]&m[1821]&m[1822])|(m[827]&~m[1818]&m[1820]&m[1821]&m[1822])|(m[827]&m[1818]&m[1820]&m[1821]&m[1822]));
    m[1824] = (((m[842]&~m[1823]&~m[1825]&~m[1826]&~m[1827])|(~m[842]&~m[1823]&~m[1825]&m[1826]&~m[1827])|(m[842]&m[1823]&~m[1825]&m[1826]&~m[1827])|(m[842]&~m[1823]&m[1825]&m[1826]&~m[1827])|(~m[842]&m[1823]&~m[1825]&~m[1826]&m[1827])|(~m[842]&~m[1823]&m[1825]&~m[1826]&m[1827])|(m[842]&m[1823]&m[1825]&~m[1826]&m[1827])|(~m[842]&m[1823]&m[1825]&m[1826]&m[1827]))&UnbiasedRNG[675])|((m[842]&~m[1823]&~m[1825]&m[1826]&~m[1827])|(~m[842]&~m[1823]&~m[1825]&~m[1826]&m[1827])|(m[842]&~m[1823]&~m[1825]&~m[1826]&m[1827])|(m[842]&m[1823]&~m[1825]&~m[1826]&m[1827])|(m[842]&~m[1823]&m[1825]&~m[1826]&m[1827])|(~m[842]&~m[1823]&~m[1825]&m[1826]&m[1827])|(m[842]&~m[1823]&~m[1825]&m[1826]&m[1827])|(~m[842]&m[1823]&~m[1825]&m[1826]&m[1827])|(m[842]&m[1823]&~m[1825]&m[1826]&m[1827])|(~m[842]&~m[1823]&m[1825]&m[1826]&m[1827])|(m[842]&~m[1823]&m[1825]&m[1826]&m[1827])|(m[842]&m[1823]&m[1825]&m[1826]&m[1827]));
    m[1829] = (((m[857]&~m[1828]&~m[1830]&~m[1831]&~m[1832])|(~m[857]&~m[1828]&~m[1830]&m[1831]&~m[1832])|(m[857]&m[1828]&~m[1830]&m[1831]&~m[1832])|(m[857]&~m[1828]&m[1830]&m[1831]&~m[1832])|(~m[857]&m[1828]&~m[1830]&~m[1831]&m[1832])|(~m[857]&~m[1828]&m[1830]&~m[1831]&m[1832])|(m[857]&m[1828]&m[1830]&~m[1831]&m[1832])|(~m[857]&m[1828]&m[1830]&m[1831]&m[1832]))&UnbiasedRNG[676])|((m[857]&~m[1828]&~m[1830]&m[1831]&~m[1832])|(~m[857]&~m[1828]&~m[1830]&~m[1831]&m[1832])|(m[857]&~m[1828]&~m[1830]&~m[1831]&m[1832])|(m[857]&m[1828]&~m[1830]&~m[1831]&m[1832])|(m[857]&~m[1828]&m[1830]&~m[1831]&m[1832])|(~m[857]&~m[1828]&~m[1830]&m[1831]&m[1832])|(m[857]&~m[1828]&~m[1830]&m[1831]&m[1832])|(~m[857]&m[1828]&~m[1830]&m[1831]&m[1832])|(m[857]&m[1828]&~m[1830]&m[1831]&m[1832])|(~m[857]&~m[1828]&m[1830]&m[1831]&m[1832])|(m[857]&~m[1828]&m[1830]&m[1831]&m[1832])|(m[857]&m[1828]&m[1830]&m[1831]&m[1832]));
    m[1834] = (((m[872]&~m[1833]&~m[1835]&~m[1836]&~m[1837])|(~m[872]&~m[1833]&~m[1835]&m[1836]&~m[1837])|(m[872]&m[1833]&~m[1835]&m[1836]&~m[1837])|(m[872]&~m[1833]&m[1835]&m[1836]&~m[1837])|(~m[872]&m[1833]&~m[1835]&~m[1836]&m[1837])|(~m[872]&~m[1833]&m[1835]&~m[1836]&m[1837])|(m[872]&m[1833]&m[1835]&~m[1836]&m[1837])|(~m[872]&m[1833]&m[1835]&m[1836]&m[1837]))&UnbiasedRNG[677])|((m[872]&~m[1833]&~m[1835]&m[1836]&~m[1837])|(~m[872]&~m[1833]&~m[1835]&~m[1836]&m[1837])|(m[872]&~m[1833]&~m[1835]&~m[1836]&m[1837])|(m[872]&m[1833]&~m[1835]&~m[1836]&m[1837])|(m[872]&~m[1833]&m[1835]&~m[1836]&m[1837])|(~m[872]&~m[1833]&~m[1835]&m[1836]&m[1837])|(m[872]&~m[1833]&~m[1835]&m[1836]&m[1837])|(~m[872]&m[1833]&~m[1835]&m[1836]&m[1837])|(m[872]&m[1833]&~m[1835]&m[1836]&m[1837])|(~m[872]&~m[1833]&m[1835]&m[1836]&m[1837])|(m[872]&~m[1833]&m[1835]&m[1836]&m[1837])|(m[872]&m[1833]&m[1835]&m[1836]&m[1837]));
    m[1839] = (((m[887]&~m[1838]&~m[1840]&~m[1841]&~m[1842])|(~m[887]&~m[1838]&~m[1840]&m[1841]&~m[1842])|(m[887]&m[1838]&~m[1840]&m[1841]&~m[1842])|(m[887]&~m[1838]&m[1840]&m[1841]&~m[1842])|(~m[887]&m[1838]&~m[1840]&~m[1841]&m[1842])|(~m[887]&~m[1838]&m[1840]&~m[1841]&m[1842])|(m[887]&m[1838]&m[1840]&~m[1841]&m[1842])|(~m[887]&m[1838]&m[1840]&m[1841]&m[1842]))&UnbiasedRNG[678])|((m[887]&~m[1838]&~m[1840]&m[1841]&~m[1842])|(~m[887]&~m[1838]&~m[1840]&~m[1841]&m[1842])|(m[887]&~m[1838]&~m[1840]&~m[1841]&m[1842])|(m[887]&m[1838]&~m[1840]&~m[1841]&m[1842])|(m[887]&~m[1838]&m[1840]&~m[1841]&m[1842])|(~m[887]&~m[1838]&~m[1840]&m[1841]&m[1842])|(m[887]&~m[1838]&~m[1840]&m[1841]&m[1842])|(~m[887]&m[1838]&~m[1840]&m[1841]&m[1842])|(m[887]&m[1838]&~m[1840]&m[1841]&m[1842])|(~m[887]&~m[1838]&m[1840]&m[1841]&m[1842])|(m[887]&~m[1838]&m[1840]&m[1841]&m[1842])|(m[887]&m[1838]&m[1840]&m[1841]&m[1842]));
    m[1844] = (((m[902]&~m[1843]&~m[1845]&~m[1846]&~m[1847])|(~m[902]&~m[1843]&~m[1845]&m[1846]&~m[1847])|(m[902]&m[1843]&~m[1845]&m[1846]&~m[1847])|(m[902]&~m[1843]&m[1845]&m[1846]&~m[1847])|(~m[902]&m[1843]&~m[1845]&~m[1846]&m[1847])|(~m[902]&~m[1843]&m[1845]&~m[1846]&m[1847])|(m[902]&m[1843]&m[1845]&~m[1846]&m[1847])|(~m[902]&m[1843]&m[1845]&m[1846]&m[1847]))&UnbiasedRNG[679])|((m[902]&~m[1843]&~m[1845]&m[1846]&~m[1847])|(~m[902]&~m[1843]&~m[1845]&~m[1846]&m[1847])|(m[902]&~m[1843]&~m[1845]&~m[1846]&m[1847])|(m[902]&m[1843]&~m[1845]&~m[1846]&m[1847])|(m[902]&~m[1843]&m[1845]&~m[1846]&m[1847])|(~m[902]&~m[1843]&~m[1845]&m[1846]&m[1847])|(m[902]&~m[1843]&~m[1845]&m[1846]&m[1847])|(~m[902]&m[1843]&~m[1845]&m[1846]&m[1847])|(m[902]&m[1843]&~m[1845]&m[1846]&m[1847])|(~m[902]&~m[1843]&m[1845]&m[1846]&m[1847])|(m[902]&~m[1843]&m[1845]&m[1846]&m[1847])|(m[902]&m[1843]&m[1845]&m[1846]&m[1847]));
    m[1849] = (((m[917]&~m[1848]&~m[1850]&~m[1851]&~m[1852])|(~m[917]&~m[1848]&~m[1850]&m[1851]&~m[1852])|(m[917]&m[1848]&~m[1850]&m[1851]&~m[1852])|(m[917]&~m[1848]&m[1850]&m[1851]&~m[1852])|(~m[917]&m[1848]&~m[1850]&~m[1851]&m[1852])|(~m[917]&~m[1848]&m[1850]&~m[1851]&m[1852])|(m[917]&m[1848]&m[1850]&~m[1851]&m[1852])|(~m[917]&m[1848]&m[1850]&m[1851]&m[1852]))&UnbiasedRNG[680])|((m[917]&~m[1848]&~m[1850]&m[1851]&~m[1852])|(~m[917]&~m[1848]&~m[1850]&~m[1851]&m[1852])|(m[917]&~m[1848]&~m[1850]&~m[1851]&m[1852])|(m[917]&m[1848]&~m[1850]&~m[1851]&m[1852])|(m[917]&~m[1848]&m[1850]&~m[1851]&m[1852])|(~m[917]&~m[1848]&~m[1850]&m[1851]&m[1852])|(m[917]&~m[1848]&~m[1850]&m[1851]&m[1852])|(~m[917]&m[1848]&~m[1850]&m[1851]&m[1852])|(m[917]&m[1848]&~m[1850]&m[1851]&m[1852])|(~m[917]&~m[1848]&m[1850]&m[1851]&m[1852])|(m[917]&~m[1848]&m[1850]&m[1851]&m[1852])|(m[917]&m[1848]&m[1850]&m[1851]&m[1852]));
    m[1854] = (((m[783]&~m[1853]&~m[1855]&~m[1856]&~m[1857])|(~m[783]&~m[1853]&~m[1855]&m[1856]&~m[1857])|(m[783]&m[1853]&~m[1855]&m[1856]&~m[1857])|(m[783]&~m[1853]&m[1855]&m[1856]&~m[1857])|(~m[783]&m[1853]&~m[1855]&~m[1856]&m[1857])|(~m[783]&~m[1853]&m[1855]&~m[1856]&m[1857])|(m[783]&m[1853]&m[1855]&~m[1856]&m[1857])|(~m[783]&m[1853]&m[1855]&m[1856]&m[1857]))&UnbiasedRNG[681])|((m[783]&~m[1853]&~m[1855]&m[1856]&~m[1857])|(~m[783]&~m[1853]&~m[1855]&~m[1856]&m[1857])|(m[783]&~m[1853]&~m[1855]&~m[1856]&m[1857])|(m[783]&m[1853]&~m[1855]&~m[1856]&m[1857])|(m[783]&~m[1853]&m[1855]&~m[1856]&m[1857])|(~m[783]&~m[1853]&~m[1855]&m[1856]&m[1857])|(m[783]&~m[1853]&~m[1855]&m[1856]&m[1857])|(~m[783]&m[1853]&~m[1855]&m[1856]&m[1857])|(m[783]&m[1853]&~m[1855]&m[1856]&m[1857])|(~m[783]&~m[1853]&m[1855]&m[1856]&m[1857])|(m[783]&~m[1853]&m[1855]&m[1856]&m[1857])|(m[783]&m[1853]&m[1855]&m[1856]&m[1857]));
    m[1859] = (((m[798]&~m[1858]&~m[1860]&~m[1861]&~m[1862])|(~m[798]&~m[1858]&~m[1860]&m[1861]&~m[1862])|(m[798]&m[1858]&~m[1860]&m[1861]&~m[1862])|(m[798]&~m[1858]&m[1860]&m[1861]&~m[1862])|(~m[798]&m[1858]&~m[1860]&~m[1861]&m[1862])|(~m[798]&~m[1858]&m[1860]&~m[1861]&m[1862])|(m[798]&m[1858]&m[1860]&~m[1861]&m[1862])|(~m[798]&m[1858]&m[1860]&m[1861]&m[1862]))&UnbiasedRNG[682])|((m[798]&~m[1858]&~m[1860]&m[1861]&~m[1862])|(~m[798]&~m[1858]&~m[1860]&~m[1861]&m[1862])|(m[798]&~m[1858]&~m[1860]&~m[1861]&m[1862])|(m[798]&m[1858]&~m[1860]&~m[1861]&m[1862])|(m[798]&~m[1858]&m[1860]&~m[1861]&m[1862])|(~m[798]&~m[1858]&~m[1860]&m[1861]&m[1862])|(m[798]&~m[1858]&~m[1860]&m[1861]&m[1862])|(~m[798]&m[1858]&~m[1860]&m[1861]&m[1862])|(m[798]&m[1858]&~m[1860]&m[1861]&m[1862])|(~m[798]&~m[1858]&m[1860]&m[1861]&m[1862])|(m[798]&~m[1858]&m[1860]&m[1861]&m[1862])|(m[798]&m[1858]&m[1860]&m[1861]&m[1862]));
    m[1864] = (((m[813]&~m[1863]&~m[1865]&~m[1866]&~m[1867])|(~m[813]&~m[1863]&~m[1865]&m[1866]&~m[1867])|(m[813]&m[1863]&~m[1865]&m[1866]&~m[1867])|(m[813]&~m[1863]&m[1865]&m[1866]&~m[1867])|(~m[813]&m[1863]&~m[1865]&~m[1866]&m[1867])|(~m[813]&~m[1863]&m[1865]&~m[1866]&m[1867])|(m[813]&m[1863]&m[1865]&~m[1866]&m[1867])|(~m[813]&m[1863]&m[1865]&m[1866]&m[1867]))&UnbiasedRNG[683])|((m[813]&~m[1863]&~m[1865]&m[1866]&~m[1867])|(~m[813]&~m[1863]&~m[1865]&~m[1866]&m[1867])|(m[813]&~m[1863]&~m[1865]&~m[1866]&m[1867])|(m[813]&m[1863]&~m[1865]&~m[1866]&m[1867])|(m[813]&~m[1863]&m[1865]&~m[1866]&m[1867])|(~m[813]&~m[1863]&~m[1865]&m[1866]&m[1867])|(m[813]&~m[1863]&~m[1865]&m[1866]&m[1867])|(~m[813]&m[1863]&~m[1865]&m[1866]&m[1867])|(m[813]&m[1863]&~m[1865]&m[1866]&m[1867])|(~m[813]&~m[1863]&m[1865]&m[1866]&m[1867])|(m[813]&~m[1863]&m[1865]&m[1866]&m[1867])|(m[813]&m[1863]&m[1865]&m[1866]&m[1867]));
    m[1869] = (((m[828]&~m[1868]&~m[1870]&~m[1871]&~m[1872])|(~m[828]&~m[1868]&~m[1870]&m[1871]&~m[1872])|(m[828]&m[1868]&~m[1870]&m[1871]&~m[1872])|(m[828]&~m[1868]&m[1870]&m[1871]&~m[1872])|(~m[828]&m[1868]&~m[1870]&~m[1871]&m[1872])|(~m[828]&~m[1868]&m[1870]&~m[1871]&m[1872])|(m[828]&m[1868]&m[1870]&~m[1871]&m[1872])|(~m[828]&m[1868]&m[1870]&m[1871]&m[1872]))&UnbiasedRNG[684])|((m[828]&~m[1868]&~m[1870]&m[1871]&~m[1872])|(~m[828]&~m[1868]&~m[1870]&~m[1871]&m[1872])|(m[828]&~m[1868]&~m[1870]&~m[1871]&m[1872])|(m[828]&m[1868]&~m[1870]&~m[1871]&m[1872])|(m[828]&~m[1868]&m[1870]&~m[1871]&m[1872])|(~m[828]&~m[1868]&~m[1870]&m[1871]&m[1872])|(m[828]&~m[1868]&~m[1870]&m[1871]&m[1872])|(~m[828]&m[1868]&~m[1870]&m[1871]&m[1872])|(m[828]&m[1868]&~m[1870]&m[1871]&m[1872])|(~m[828]&~m[1868]&m[1870]&m[1871]&m[1872])|(m[828]&~m[1868]&m[1870]&m[1871]&m[1872])|(m[828]&m[1868]&m[1870]&m[1871]&m[1872]));
    m[1874] = (((m[843]&~m[1873]&~m[1875]&~m[1876]&~m[1877])|(~m[843]&~m[1873]&~m[1875]&m[1876]&~m[1877])|(m[843]&m[1873]&~m[1875]&m[1876]&~m[1877])|(m[843]&~m[1873]&m[1875]&m[1876]&~m[1877])|(~m[843]&m[1873]&~m[1875]&~m[1876]&m[1877])|(~m[843]&~m[1873]&m[1875]&~m[1876]&m[1877])|(m[843]&m[1873]&m[1875]&~m[1876]&m[1877])|(~m[843]&m[1873]&m[1875]&m[1876]&m[1877]))&UnbiasedRNG[685])|((m[843]&~m[1873]&~m[1875]&m[1876]&~m[1877])|(~m[843]&~m[1873]&~m[1875]&~m[1876]&m[1877])|(m[843]&~m[1873]&~m[1875]&~m[1876]&m[1877])|(m[843]&m[1873]&~m[1875]&~m[1876]&m[1877])|(m[843]&~m[1873]&m[1875]&~m[1876]&m[1877])|(~m[843]&~m[1873]&~m[1875]&m[1876]&m[1877])|(m[843]&~m[1873]&~m[1875]&m[1876]&m[1877])|(~m[843]&m[1873]&~m[1875]&m[1876]&m[1877])|(m[843]&m[1873]&~m[1875]&m[1876]&m[1877])|(~m[843]&~m[1873]&m[1875]&m[1876]&m[1877])|(m[843]&~m[1873]&m[1875]&m[1876]&m[1877])|(m[843]&m[1873]&m[1875]&m[1876]&m[1877]));
    m[1879] = (((m[858]&~m[1878]&~m[1880]&~m[1881]&~m[1882])|(~m[858]&~m[1878]&~m[1880]&m[1881]&~m[1882])|(m[858]&m[1878]&~m[1880]&m[1881]&~m[1882])|(m[858]&~m[1878]&m[1880]&m[1881]&~m[1882])|(~m[858]&m[1878]&~m[1880]&~m[1881]&m[1882])|(~m[858]&~m[1878]&m[1880]&~m[1881]&m[1882])|(m[858]&m[1878]&m[1880]&~m[1881]&m[1882])|(~m[858]&m[1878]&m[1880]&m[1881]&m[1882]))&UnbiasedRNG[686])|((m[858]&~m[1878]&~m[1880]&m[1881]&~m[1882])|(~m[858]&~m[1878]&~m[1880]&~m[1881]&m[1882])|(m[858]&~m[1878]&~m[1880]&~m[1881]&m[1882])|(m[858]&m[1878]&~m[1880]&~m[1881]&m[1882])|(m[858]&~m[1878]&m[1880]&~m[1881]&m[1882])|(~m[858]&~m[1878]&~m[1880]&m[1881]&m[1882])|(m[858]&~m[1878]&~m[1880]&m[1881]&m[1882])|(~m[858]&m[1878]&~m[1880]&m[1881]&m[1882])|(m[858]&m[1878]&~m[1880]&m[1881]&m[1882])|(~m[858]&~m[1878]&m[1880]&m[1881]&m[1882])|(m[858]&~m[1878]&m[1880]&m[1881]&m[1882])|(m[858]&m[1878]&m[1880]&m[1881]&m[1882]));
    m[1884] = (((m[873]&~m[1883]&~m[1885]&~m[1886]&~m[1887])|(~m[873]&~m[1883]&~m[1885]&m[1886]&~m[1887])|(m[873]&m[1883]&~m[1885]&m[1886]&~m[1887])|(m[873]&~m[1883]&m[1885]&m[1886]&~m[1887])|(~m[873]&m[1883]&~m[1885]&~m[1886]&m[1887])|(~m[873]&~m[1883]&m[1885]&~m[1886]&m[1887])|(m[873]&m[1883]&m[1885]&~m[1886]&m[1887])|(~m[873]&m[1883]&m[1885]&m[1886]&m[1887]))&UnbiasedRNG[687])|((m[873]&~m[1883]&~m[1885]&m[1886]&~m[1887])|(~m[873]&~m[1883]&~m[1885]&~m[1886]&m[1887])|(m[873]&~m[1883]&~m[1885]&~m[1886]&m[1887])|(m[873]&m[1883]&~m[1885]&~m[1886]&m[1887])|(m[873]&~m[1883]&m[1885]&~m[1886]&m[1887])|(~m[873]&~m[1883]&~m[1885]&m[1886]&m[1887])|(m[873]&~m[1883]&~m[1885]&m[1886]&m[1887])|(~m[873]&m[1883]&~m[1885]&m[1886]&m[1887])|(m[873]&m[1883]&~m[1885]&m[1886]&m[1887])|(~m[873]&~m[1883]&m[1885]&m[1886]&m[1887])|(m[873]&~m[1883]&m[1885]&m[1886]&m[1887])|(m[873]&m[1883]&m[1885]&m[1886]&m[1887]));
    m[1889] = (((m[888]&~m[1888]&~m[1890]&~m[1891]&~m[1892])|(~m[888]&~m[1888]&~m[1890]&m[1891]&~m[1892])|(m[888]&m[1888]&~m[1890]&m[1891]&~m[1892])|(m[888]&~m[1888]&m[1890]&m[1891]&~m[1892])|(~m[888]&m[1888]&~m[1890]&~m[1891]&m[1892])|(~m[888]&~m[1888]&m[1890]&~m[1891]&m[1892])|(m[888]&m[1888]&m[1890]&~m[1891]&m[1892])|(~m[888]&m[1888]&m[1890]&m[1891]&m[1892]))&UnbiasedRNG[688])|((m[888]&~m[1888]&~m[1890]&m[1891]&~m[1892])|(~m[888]&~m[1888]&~m[1890]&~m[1891]&m[1892])|(m[888]&~m[1888]&~m[1890]&~m[1891]&m[1892])|(m[888]&m[1888]&~m[1890]&~m[1891]&m[1892])|(m[888]&~m[1888]&m[1890]&~m[1891]&m[1892])|(~m[888]&~m[1888]&~m[1890]&m[1891]&m[1892])|(m[888]&~m[1888]&~m[1890]&m[1891]&m[1892])|(~m[888]&m[1888]&~m[1890]&m[1891]&m[1892])|(m[888]&m[1888]&~m[1890]&m[1891]&m[1892])|(~m[888]&~m[1888]&m[1890]&m[1891]&m[1892])|(m[888]&~m[1888]&m[1890]&m[1891]&m[1892])|(m[888]&m[1888]&m[1890]&m[1891]&m[1892]));
    m[1894] = (((m[903]&~m[1893]&~m[1895]&~m[1896]&~m[1897])|(~m[903]&~m[1893]&~m[1895]&m[1896]&~m[1897])|(m[903]&m[1893]&~m[1895]&m[1896]&~m[1897])|(m[903]&~m[1893]&m[1895]&m[1896]&~m[1897])|(~m[903]&m[1893]&~m[1895]&~m[1896]&m[1897])|(~m[903]&~m[1893]&m[1895]&~m[1896]&m[1897])|(m[903]&m[1893]&m[1895]&~m[1896]&m[1897])|(~m[903]&m[1893]&m[1895]&m[1896]&m[1897]))&UnbiasedRNG[689])|((m[903]&~m[1893]&~m[1895]&m[1896]&~m[1897])|(~m[903]&~m[1893]&~m[1895]&~m[1896]&m[1897])|(m[903]&~m[1893]&~m[1895]&~m[1896]&m[1897])|(m[903]&m[1893]&~m[1895]&~m[1896]&m[1897])|(m[903]&~m[1893]&m[1895]&~m[1896]&m[1897])|(~m[903]&~m[1893]&~m[1895]&m[1896]&m[1897])|(m[903]&~m[1893]&~m[1895]&m[1896]&m[1897])|(~m[903]&m[1893]&~m[1895]&m[1896]&m[1897])|(m[903]&m[1893]&~m[1895]&m[1896]&m[1897])|(~m[903]&~m[1893]&m[1895]&m[1896]&m[1897])|(m[903]&~m[1893]&m[1895]&m[1896]&m[1897])|(m[903]&m[1893]&m[1895]&m[1896]&m[1897]));
    m[1899] = (((m[918]&~m[1898]&~m[1900]&~m[1901]&~m[1902])|(~m[918]&~m[1898]&~m[1900]&m[1901]&~m[1902])|(m[918]&m[1898]&~m[1900]&m[1901]&~m[1902])|(m[918]&~m[1898]&m[1900]&m[1901]&~m[1902])|(~m[918]&m[1898]&~m[1900]&~m[1901]&m[1902])|(~m[918]&~m[1898]&m[1900]&~m[1901]&m[1902])|(m[918]&m[1898]&m[1900]&~m[1901]&m[1902])|(~m[918]&m[1898]&m[1900]&m[1901]&m[1902]))&UnbiasedRNG[690])|((m[918]&~m[1898]&~m[1900]&m[1901]&~m[1902])|(~m[918]&~m[1898]&~m[1900]&~m[1901]&m[1902])|(m[918]&~m[1898]&~m[1900]&~m[1901]&m[1902])|(m[918]&m[1898]&~m[1900]&~m[1901]&m[1902])|(m[918]&~m[1898]&m[1900]&~m[1901]&m[1902])|(~m[918]&~m[1898]&~m[1900]&m[1901]&m[1902])|(m[918]&~m[1898]&~m[1900]&m[1901]&m[1902])|(~m[918]&m[1898]&~m[1900]&m[1901]&m[1902])|(m[918]&m[1898]&~m[1900]&m[1901]&m[1902])|(~m[918]&~m[1898]&m[1900]&m[1901]&m[1902])|(m[918]&~m[1898]&m[1900]&m[1901]&m[1902])|(m[918]&m[1898]&m[1900]&m[1901]&m[1902]));
    m[1904] = (((m[799]&~m[1903]&~m[1905]&~m[1906]&~m[1907])|(~m[799]&~m[1903]&~m[1905]&m[1906]&~m[1907])|(m[799]&m[1903]&~m[1905]&m[1906]&~m[1907])|(m[799]&~m[1903]&m[1905]&m[1906]&~m[1907])|(~m[799]&m[1903]&~m[1905]&~m[1906]&m[1907])|(~m[799]&~m[1903]&m[1905]&~m[1906]&m[1907])|(m[799]&m[1903]&m[1905]&~m[1906]&m[1907])|(~m[799]&m[1903]&m[1905]&m[1906]&m[1907]))&UnbiasedRNG[691])|((m[799]&~m[1903]&~m[1905]&m[1906]&~m[1907])|(~m[799]&~m[1903]&~m[1905]&~m[1906]&m[1907])|(m[799]&~m[1903]&~m[1905]&~m[1906]&m[1907])|(m[799]&m[1903]&~m[1905]&~m[1906]&m[1907])|(m[799]&~m[1903]&m[1905]&~m[1906]&m[1907])|(~m[799]&~m[1903]&~m[1905]&m[1906]&m[1907])|(m[799]&~m[1903]&~m[1905]&m[1906]&m[1907])|(~m[799]&m[1903]&~m[1905]&m[1906]&m[1907])|(m[799]&m[1903]&~m[1905]&m[1906]&m[1907])|(~m[799]&~m[1903]&m[1905]&m[1906]&m[1907])|(m[799]&~m[1903]&m[1905]&m[1906]&m[1907])|(m[799]&m[1903]&m[1905]&m[1906]&m[1907]));
    m[1909] = (((m[814]&~m[1908]&~m[1910]&~m[1911]&~m[1912])|(~m[814]&~m[1908]&~m[1910]&m[1911]&~m[1912])|(m[814]&m[1908]&~m[1910]&m[1911]&~m[1912])|(m[814]&~m[1908]&m[1910]&m[1911]&~m[1912])|(~m[814]&m[1908]&~m[1910]&~m[1911]&m[1912])|(~m[814]&~m[1908]&m[1910]&~m[1911]&m[1912])|(m[814]&m[1908]&m[1910]&~m[1911]&m[1912])|(~m[814]&m[1908]&m[1910]&m[1911]&m[1912]))&UnbiasedRNG[692])|((m[814]&~m[1908]&~m[1910]&m[1911]&~m[1912])|(~m[814]&~m[1908]&~m[1910]&~m[1911]&m[1912])|(m[814]&~m[1908]&~m[1910]&~m[1911]&m[1912])|(m[814]&m[1908]&~m[1910]&~m[1911]&m[1912])|(m[814]&~m[1908]&m[1910]&~m[1911]&m[1912])|(~m[814]&~m[1908]&~m[1910]&m[1911]&m[1912])|(m[814]&~m[1908]&~m[1910]&m[1911]&m[1912])|(~m[814]&m[1908]&~m[1910]&m[1911]&m[1912])|(m[814]&m[1908]&~m[1910]&m[1911]&m[1912])|(~m[814]&~m[1908]&m[1910]&m[1911]&m[1912])|(m[814]&~m[1908]&m[1910]&m[1911]&m[1912])|(m[814]&m[1908]&m[1910]&m[1911]&m[1912]));
    m[1914] = (((m[829]&~m[1913]&~m[1915]&~m[1916]&~m[1917])|(~m[829]&~m[1913]&~m[1915]&m[1916]&~m[1917])|(m[829]&m[1913]&~m[1915]&m[1916]&~m[1917])|(m[829]&~m[1913]&m[1915]&m[1916]&~m[1917])|(~m[829]&m[1913]&~m[1915]&~m[1916]&m[1917])|(~m[829]&~m[1913]&m[1915]&~m[1916]&m[1917])|(m[829]&m[1913]&m[1915]&~m[1916]&m[1917])|(~m[829]&m[1913]&m[1915]&m[1916]&m[1917]))&UnbiasedRNG[693])|((m[829]&~m[1913]&~m[1915]&m[1916]&~m[1917])|(~m[829]&~m[1913]&~m[1915]&~m[1916]&m[1917])|(m[829]&~m[1913]&~m[1915]&~m[1916]&m[1917])|(m[829]&m[1913]&~m[1915]&~m[1916]&m[1917])|(m[829]&~m[1913]&m[1915]&~m[1916]&m[1917])|(~m[829]&~m[1913]&~m[1915]&m[1916]&m[1917])|(m[829]&~m[1913]&~m[1915]&m[1916]&m[1917])|(~m[829]&m[1913]&~m[1915]&m[1916]&m[1917])|(m[829]&m[1913]&~m[1915]&m[1916]&m[1917])|(~m[829]&~m[1913]&m[1915]&m[1916]&m[1917])|(m[829]&~m[1913]&m[1915]&m[1916]&m[1917])|(m[829]&m[1913]&m[1915]&m[1916]&m[1917]));
    m[1919] = (((m[844]&~m[1918]&~m[1920]&~m[1921]&~m[1922])|(~m[844]&~m[1918]&~m[1920]&m[1921]&~m[1922])|(m[844]&m[1918]&~m[1920]&m[1921]&~m[1922])|(m[844]&~m[1918]&m[1920]&m[1921]&~m[1922])|(~m[844]&m[1918]&~m[1920]&~m[1921]&m[1922])|(~m[844]&~m[1918]&m[1920]&~m[1921]&m[1922])|(m[844]&m[1918]&m[1920]&~m[1921]&m[1922])|(~m[844]&m[1918]&m[1920]&m[1921]&m[1922]))&UnbiasedRNG[694])|((m[844]&~m[1918]&~m[1920]&m[1921]&~m[1922])|(~m[844]&~m[1918]&~m[1920]&~m[1921]&m[1922])|(m[844]&~m[1918]&~m[1920]&~m[1921]&m[1922])|(m[844]&m[1918]&~m[1920]&~m[1921]&m[1922])|(m[844]&~m[1918]&m[1920]&~m[1921]&m[1922])|(~m[844]&~m[1918]&~m[1920]&m[1921]&m[1922])|(m[844]&~m[1918]&~m[1920]&m[1921]&m[1922])|(~m[844]&m[1918]&~m[1920]&m[1921]&m[1922])|(m[844]&m[1918]&~m[1920]&m[1921]&m[1922])|(~m[844]&~m[1918]&m[1920]&m[1921]&m[1922])|(m[844]&~m[1918]&m[1920]&m[1921]&m[1922])|(m[844]&m[1918]&m[1920]&m[1921]&m[1922]));
    m[1924] = (((m[859]&~m[1923]&~m[1925]&~m[1926]&~m[1927])|(~m[859]&~m[1923]&~m[1925]&m[1926]&~m[1927])|(m[859]&m[1923]&~m[1925]&m[1926]&~m[1927])|(m[859]&~m[1923]&m[1925]&m[1926]&~m[1927])|(~m[859]&m[1923]&~m[1925]&~m[1926]&m[1927])|(~m[859]&~m[1923]&m[1925]&~m[1926]&m[1927])|(m[859]&m[1923]&m[1925]&~m[1926]&m[1927])|(~m[859]&m[1923]&m[1925]&m[1926]&m[1927]))&UnbiasedRNG[695])|((m[859]&~m[1923]&~m[1925]&m[1926]&~m[1927])|(~m[859]&~m[1923]&~m[1925]&~m[1926]&m[1927])|(m[859]&~m[1923]&~m[1925]&~m[1926]&m[1927])|(m[859]&m[1923]&~m[1925]&~m[1926]&m[1927])|(m[859]&~m[1923]&m[1925]&~m[1926]&m[1927])|(~m[859]&~m[1923]&~m[1925]&m[1926]&m[1927])|(m[859]&~m[1923]&~m[1925]&m[1926]&m[1927])|(~m[859]&m[1923]&~m[1925]&m[1926]&m[1927])|(m[859]&m[1923]&~m[1925]&m[1926]&m[1927])|(~m[859]&~m[1923]&m[1925]&m[1926]&m[1927])|(m[859]&~m[1923]&m[1925]&m[1926]&m[1927])|(m[859]&m[1923]&m[1925]&m[1926]&m[1927]));
    m[1929] = (((m[874]&~m[1928]&~m[1930]&~m[1931]&~m[1932])|(~m[874]&~m[1928]&~m[1930]&m[1931]&~m[1932])|(m[874]&m[1928]&~m[1930]&m[1931]&~m[1932])|(m[874]&~m[1928]&m[1930]&m[1931]&~m[1932])|(~m[874]&m[1928]&~m[1930]&~m[1931]&m[1932])|(~m[874]&~m[1928]&m[1930]&~m[1931]&m[1932])|(m[874]&m[1928]&m[1930]&~m[1931]&m[1932])|(~m[874]&m[1928]&m[1930]&m[1931]&m[1932]))&UnbiasedRNG[696])|((m[874]&~m[1928]&~m[1930]&m[1931]&~m[1932])|(~m[874]&~m[1928]&~m[1930]&~m[1931]&m[1932])|(m[874]&~m[1928]&~m[1930]&~m[1931]&m[1932])|(m[874]&m[1928]&~m[1930]&~m[1931]&m[1932])|(m[874]&~m[1928]&m[1930]&~m[1931]&m[1932])|(~m[874]&~m[1928]&~m[1930]&m[1931]&m[1932])|(m[874]&~m[1928]&~m[1930]&m[1931]&m[1932])|(~m[874]&m[1928]&~m[1930]&m[1931]&m[1932])|(m[874]&m[1928]&~m[1930]&m[1931]&m[1932])|(~m[874]&~m[1928]&m[1930]&m[1931]&m[1932])|(m[874]&~m[1928]&m[1930]&m[1931]&m[1932])|(m[874]&m[1928]&m[1930]&m[1931]&m[1932]));
    m[1934] = (((m[889]&~m[1933]&~m[1935]&~m[1936]&~m[1937])|(~m[889]&~m[1933]&~m[1935]&m[1936]&~m[1937])|(m[889]&m[1933]&~m[1935]&m[1936]&~m[1937])|(m[889]&~m[1933]&m[1935]&m[1936]&~m[1937])|(~m[889]&m[1933]&~m[1935]&~m[1936]&m[1937])|(~m[889]&~m[1933]&m[1935]&~m[1936]&m[1937])|(m[889]&m[1933]&m[1935]&~m[1936]&m[1937])|(~m[889]&m[1933]&m[1935]&m[1936]&m[1937]))&UnbiasedRNG[697])|((m[889]&~m[1933]&~m[1935]&m[1936]&~m[1937])|(~m[889]&~m[1933]&~m[1935]&~m[1936]&m[1937])|(m[889]&~m[1933]&~m[1935]&~m[1936]&m[1937])|(m[889]&m[1933]&~m[1935]&~m[1936]&m[1937])|(m[889]&~m[1933]&m[1935]&~m[1936]&m[1937])|(~m[889]&~m[1933]&~m[1935]&m[1936]&m[1937])|(m[889]&~m[1933]&~m[1935]&m[1936]&m[1937])|(~m[889]&m[1933]&~m[1935]&m[1936]&m[1937])|(m[889]&m[1933]&~m[1935]&m[1936]&m[1937])|(~m[889]&~m[1933]&m[1935]&m[1936]&m[1937])|(m[889]&~m[1933]&m[1935]&m[1936]&m[1937])|(m[889]&m[1933]&m[1935]&m[1936]&m[1937]));
    m[1939] = (((m[904]&~m[1938]&~m[1940]&~m[1941]&~m[1942])|(~m[904]&~m[1938]&~m[1940]&m[1941]&~m[1942])|(m[904]&m[1938]&~m[1940]&m[1941]&~m[1942])|(m[904]&~m[1938]&m[1940]&m[1941]&~m[1942])|(~m[904]&m[1938]&~m[1940]&~m[1941]&m[1942])|(~m[904]&~m[1938]&m[1940]&~m[1941]&m[1942])|(m[904]&m[1938]&m[1940]&~m[1941]&m[1942])|(~m[904]&m[1938]&m[1940]&m[1941]&m[1942]))&UnbiasedRNG[698])|((m[904]&~m[1938]&~m[1940]&m[1941]&~m[1942])|(~m[904]&~m[1938]&~m[1940]&~m[1941]&m[1942])|(m[904]&~m[1938]&~m[1940]&~m[1941]&m[1942])|(m[904]&m[1938]&~m[1940]&~m[1941]&m[1942])|(m[904]&~m[1938]&m[1940]&~m[1941]&m[1942])|(~m[904]&~m[1938]&~m[1940]&m[1941]&m[1942])|(m[904]&~m[1938]&~m[1940]&m[1941]&m[1942])|(~m[904]&m[1938]&~m[1940]&m[1941]&m[1942])|(m[904]&m[1938]&~m[1940]&m[1941]&m[1942])|(~m[904]&~m[1938]&m[1940]&m[1941]&m[1942])|(m[904]&~m[1938]&m[1940]&m[1941]&m[1942])|(m[904]&m[1938]&m[1940]&m[1941]&m[1942]));
    m[1944] = (((m[919]&~m[1943]&~m[1945]&~m[1946]&~m[1947])|(~m[919]&~m[1943]&~m[1945]&m[1946]&~m[1947])|(m[919]&m[1943]&~m[1945]&m[1946]&~m[1947])|(m[919]&~m[1943]&m[1945]&m[1946]&~m[1947])|(~m[919]&m[1943]&~m[1945]&~m[1946]&m[1947])|(~m[919]&~m[1943]&m[1945]&~m[1946]&m[1947])|(m[919]&m[1943]&m[1945]&~m[1946]&m[1947])|(~m[919]&m[1943]&m[1945]&m[1946]&m[1947]))&UnbiasedRNG[699])|((m[919]&~m[1943]&~m[1945]&m[1946]&~m[1947])|(~m[919]&~m[1943]&~m[1945]&~m[1946]&m[1947])|(m[919]&~m[1943]&~m[1945]&~m[1946]&m[1947])|(m[919]&m[1943]&~m[1945]&~m[1946]&m[1947])|(m[919]&~m[1943]&m[1945]&~m[1946]&m[1947])|(~m[919]&~m[1943]&~m[1945]&m[1946]&m[1947])|(m[919]&~m[1943]&~m[1945]&m[1946]&m[1947])|(~m[919]&m[1943]&~m[1945]&m[1946]&m[1947])|(m[919]&m[1943]&~m[1945]&m[1946]&m[1947])|(~m[919]&~m[1943]&m[1945]&m[1946]&m[1947])|(m[919]&~m[1943]&m[1945]&m[1946]&m[1947])|(m[919]&m[1943]&m[1945]&m[1946]&m[1947]));
    m[1949] = (((m[815]&~m[1948]&~m[1950]&~m[1951]&~m[1952])|(~m[815]&~m[1948]&~m[1950]&m[1951]&~m[1952])|(m[815]&m[1948]&~m[1950]&m[1951]&~m[1952])|(m[815]&~m[1948]&m[1950]&m[1951]&~m[1952])|(~m[815]&m[1948]&~m[1950]&~m[1951]&m[1952])|(~m[815]&~m[1948]&m[1950]&~m[1951]&m[1952])|(m[815]&m[1948]&m[1950]&~m[1951]&m[1952])|(~m[815]&m[1948]&m[1950]&m[1951]&m[1952]))&UnbiasedRNG[700])|((m[815]&~m[1948]&~m[1950]&m[1951]&~m[1952])|(~m[815]&~m[1948]&~m[1950]&~m[1951]&m[1952])|(m[815]&~m[1948]&~m[1950]&~m[1951]&m[1952])|(m[815]&m[1948]&~m[1950]&~m[1951]&m[1952])|(m[815]&~m[1948]&m[1950]&~m[1951]&m[1952])|(~m[815]&~m[1948]&~m[1950]&m[1951]&m[1952])|(m[815]&~m[1948]&~m[1950]&m[1951]&m[1952])|(~m[815]&m[1948]&~m[1950]&m[1951]&m[1952])|(m[815]&m[1948]&~m[1950]&m[1951]&m[1952])|(~m[815]&~m[1948]&m[1950]&m[1951]&m[1952])|(m[815]&~m[1948]&m[1950]&m[1951]&m[1952])|(m[815]&m[1948]&m[1950]&m[1951]&m[1952]));
    m[1954] = (((m[830]&~m[1953]&~m[1955]&~m[1956]&~m[1957])|(~m[830]&~m[1953]&~m[1955]&m[1956]&~m[1957])|(m[830]&m[1953]&~m[1955]&m[1956]&~m[1957])|(m[830]&~m[1953]&m[1955]&m[1956]&~m[1957])|(~m[830]&m[1953]&~m[1955]&~m[1956]&m[1957])|(~m[830]&~m[1953]&m[1955]&~m[1956]&m[1957])|(m[830]&m[1953]&m[1955]&~m[1956]&m[1957])|(~m[830]&m[1953]&m[1955]&m[1956]&m[1957]))&UnbiasedRNG[701])|((m[830]&~m[1953]&~m[1955]&m[1956]&~m[1957])|(~m[830]&~m[1953]&~m[1955]&~m[1956]&m[1957])|(m[830]&~m[1953]&~m[1955]&~m[1956]&m[1957])|(m[830]&m[1953]&~m[1955]&~m[1956]&m[1957])|(m[830]&~m[1953]&m[1955]&~m[1956]&m[1957])|(~m[830]&~m[1953]&~m[1955]&m[1956]&m[1957])|(m[830]&~m[1953]&~m[1955]&m[1956]&m[1957])|(~m[830]&m[1953]&~m[1955]&m[1956]&m[1957])|(m[830]&m[1953]&~m[1955]&m[1956]&m[1957])|(~m[830]&~m[1953]&m[1955]&m[1956]&m[1957])|(m[830]&~m[1953]&m[1955]&m[1956]&m[1957])|(m[830]&m[1953]&m[1955]&m[1956]&m[1957]));
    m[1959] = (((m[845]&~m[1958]&~m[1960]&~m[1961]&~m[1962])|(~m[845]&~m[1958]&~m[1960]&m[1961]&~m[1962])|(m[845]&m[1958]&~m[1960]&m[1961]&~m[1962])|(m[845]&~m[1958]&m[1960]&m[1961]&~m[1962])|(~m[845]&m[1958]&~m[1960]&~m[1961]&m[1962])|(~m[845]&~m[1958]&m[1960]&~m[1961]&m[1962])|(m[845]&m[1958]&m[1960]&~m[1961]&m[1962])|(~m[845]&m[1958]&m[1960]&m[1961]&m[1962]))&UnbiasedRNG[702])|((m[845]&~m[1958]&~m[1960]&m[1961]&~m[1962])|(~m[845]&~m[1958]&~m[1960]&~m[1961]&m[1962])|(m[845]&~m[1958]&~m[1960]&~m[1961]&m[1962])|(m[845]&m[1958]&~m[1960]&~m[1961]&m[1962])|(m[845]&~m[1958]&m[1960]&~m[1961]&m[1962])|(~m[845]&~m[1958]&~m[1960]&m[1961]&m[1962])|(m[845]&~m[1958]&~m[1960]&m[1961]&m[1962])|(~m[845]&m[1958]&~m[1960]&m[1961]&m[1962])|(m[845]&m[1958]&~m[1960]&m[1961]&m[1962])|(~m[845]&~m[1958]&m[1960]&m[1961]&m[1962])|(m[845]&~m[1958]&m[1960]&m[1961]&m[1962])|(m[845]&m[1958]&m[1960]&m[1961]&m[1962]));
    m[1964] = (((m[860]&~m[1963]&~m[1965]&~m[1966]&~m[1967])|(~m[860]&~m[1963]&~m[1965]&m[1966]&~m[1967])|(m[860]&m[1963]&~m[1965]&m[1966]&~m[1967])|(m[860]&~m[1963]&m[1965]&m[1966]&~m[1967])|(~m[860]&m[1963]&~m[1965]&~m[1966]&m[1967])|(~m[860]&~m[1963]&m[1965]&~m[1966]&m[1967])|(m[860]&m[1963]&m[1965]&~m[1966]&m[1967])|(~m[860]&m[1963]&m[1965]&m[1966]&m[1967]))&UnbiasedRNG[703])|((m[860]&~m[1963]&~m[1965]&m[1966]&~m[1967])|(~m[860]&~m[1963]&~m[1965]&~m[1966]&m[1967])|(m[860]&~m[1963]&~m[1965]&~m[1966]&m[1967])|(m[860]&m[1963]&~m[1965]&~m[1966]&m[1967])|(m[860]&~m[1963]&m[1965]&~m[1966]&m[1967])|(~m[860]&~m[1963]&~m[1965]&m[1966]&m[1967])|(m[860]&~m[1963]&~m[1965]&m[1966]&m[1967])|(~m[860]&m[1963]&~m[1965]&m[1966]&m[1967])|(m[860]&m[1963]&~m[1965]&m[1966]&m[1967])|(~m[860]&~m[1963]&m[1965]&m[1966]&m[1967])|(m[860]&~m[1963]&m[1965]&m[1966]&m[1967])|(m[860]&m[1963]&m[1965]&m[1966]&m[1967]));
    m[1969] = (((m[875]&~m[1968]&~m[1970]&~m[1971]&~m[1972])|(~m[875]&~m[1968]&~m[1970]&m[1971]&~m[1972])|(m[875]&m[1968]&~m[1970]&m[1971]&~m[1972])|(m[875]&~m[1968]&m[1970]&m[1971]&~m[1972])|(~m[875]&m[1968]&~m[1970]&~m[1971]&m[1972])|(~m[875]&~m[1968]&m[1970]&~m[1971]&m[1972])|(m[875]&m[1968]&m[1970]&~m[1971]&m[1972])|(~m[875]&m[1968]&m[1970]&m[1971]&m[1972]))&UnbiasedRNG[704])|((m[875]&~m[1968]&~m[1970]&m[1971]&~m[1972])|(~m[875]&~m[1968]&~m[1970]&~m[1971]&m[1972])|(m[875]&~m[1968]&~m[1970]&~m[1971]&m[1972])|(m[875]&m[1968]&~m[1970]&~m[1971]&m[1972])|(m[875]&~m[1968]&m[1970]&~m[1971]&m[1972])|(~m[875]&~m[1968]&~m[1970]&m[1971]&m[1972])|(m[875]&~m[1968]&~m[1970]&m[1971]&m[1972])|(~m[875]&m[1968]&~m[1970]&m[1971]&m[1972])|(m[875]&m[1968]&~m[1970]&m[1971]&m[1972])|(~m[875]&~m[1968]&m[1970]&m[1971]&m[1972])|(m[875]&~m[1968]&m[1970]&m[1971]&m[1972])|(m[875]&m[1968]&m[1970]&m[1971]&m[1972]));
    m[1974] = (((m[890]&~m[1973]&~m[1975]&~m[1976]&~m[1977])|(~m[890]&~m[1973]&~m[1975]&m[1976]&~m[1977])|(m[890]&m[1973]&~m[1975]&m[1976]&~m[1977])|(m[890]&~m[1973]&m[1975]&m[1976]&~m[1977])|(~m[890]&m[1973]&~m[1975]&~m[1976]&m[1977])|(~m[890]&~m[1973]&m[1975]&~m[1976]&m[1977])|(m[890]&m[1973]&m[1975]&~m[1976]&m[1977])|(~m[890]&m[1973]&m[1975]&m[1976]&m[1977]))&UnbiasedRNG[705])|((m[890]&~m[1973]&~m[1975]&m[1976]&~m[1977])|(~m[890]&~m[1973]&~m[1975]&~m[1976]&m[1977])|(m[890]&~m[1973]&~m[1975]&~m[1976]&m[1977])|(m[890]&m[1973]&~m[1975]&~m[1976]&m[1977])|(m[890]&~m[1973]&m[1975]&~m[1976]&m[1977])|(~m[890]&~m[1973]&~m[1975]&m[1976]&m[1977])|(m[890]&~m[1973]&~m[1975]&m[1976]&m[1977])|(~m[890]&m[1973]&~m[1975]&m[1976]&m[1977])|(m[890]&m[1973]&~m[1975]&m[1976]&m[1977])|(~m[890]&~m[1973]&m[1975]&m[1976]&m[1977])|(m[890]&~m[1973]&m[1975]&m[1976]&m[1977])|(m[890]&m[1973]&m[1975]&m[1976]&m[1977]));
    m[1979] = (((m[905]&~m[1978]&~m[1980]&~m[1981]&~m[1982])|(~m[905]&~m[1978]&~m[1980]&m[1981]&~m[1982])|(m[905]&m[1978]&~m[1980]&m[1981]&~m[1982])|(m[905]&~m[1978]&m[1980]&m[1981]&~m[1982])|(~m[905]&m[1978]&~m[1980]&~m[1981]&m[1982])|(~m[905]&~m[1978]&m[1980]&~m[1981]&m[1982])|(m[905]&m[1978]&m[1980]&~m[1981]&m[1982])|(~m[905]&m[1978]&m[1980]&m[1981]&m[1982]))&UnbiasedRNG[706])|((m[905]&~m[1978]&~m[1980]&m[1981]&~m[1982])|(~m[905]&~m[1978]&~m[1980]&~m[1981]&m[1982])|(m[905]&~m[1978]&~m[1980]&~m[1981]&m[1982])|(m[905]&m[1978]&~m[1980]&~m[1981]&m[1982])|(m[905]&~m[1978]&m[1980]&~m[1981]&m[1982])|(~m[905]&~m[1978]&~m[1980]&m[1981]&m[1982])|(m[905]&~m[1978]&~m[1980]&m[1981]&m[1982])|(~m[905]&m[1978]&~m[1980]&m[1981]&m[1982])|(m[905]&m[1978]&~m[1980]&m[1981]&m[1982])|(~m[905]&~m[1978]&m[1980]&m[1981]&m[1982])|(m[905]&~m[1978]&m[1980]&m[1981]&m[1982])|(m[905]&m[1978]&m[1980]&m[1981]&m[1982]));
    m[1984] = (((m[920]&~m[1983]&~m[1985]&~m[1986]&~m[1987])|(~m[920]&~m[1983]&~m[1985]&m[1986]&~m[1987])|(m[920]&m[1983]&~m[1985]&m[1986]&~m[1987])|(m[920]&~m[1983]&m[1985]&m[1986]&~m[1987])|(~m[920]&m[1983]&~m[1985]&~m[1986]&m[1987])|(~m[920]&~m[1983]&m[1985]&~m[1986]&m[1987])|(m[920]&m[1983]&m[1985]&~m[1986]&m[1987])|(~m[920]&m[1983]&m[1985]&m[1986]&m[1987]))&UnbiasedRNG[707])|((m[920]&~m[1983]&~m[1985]&m[1986]&~m[1987])|(~m[920]&~m[1983]&~m[1985]&~m[1986]&m[1987])|(m[920]&~m[1983]&~m[1985]&~m[1986]&m[1987])|(m[920]&m[1983]&~m[1985]&~m[1986]&m[1987])|(m[920]&~m[1983]&m[1985]&~m[1986]&m[1987])|(~m[920]&~m[1983]&~m[1985]&m[1986]&m[1987])|(m[920]&~m[1983]&~m[1985]&m[1986]&m[1987])|(~m[920]&m[1983]&~m[1985]&m[1986]&m[1987])|(m[920]&m[1983]&~m[1985]&m[1986]&m[1987])|(~m[920]&~m[1983]&m[1985]&m[1986]&m[1987])|(m[920]&~m[1983]&m[1985]&m[1986]&m[1987])|(m[920]&m[1983]&m[1985]&m[1986]&m[1987]));
    m[1989] = (((m[831]&~m[1988]&~m[1990]&~m[1991]&~m[1992])|(~m[831]&~m[1988]&~m[1990]&m[1991]&~m[1992])|(m[831]&m[1988]&~m[1990]&m[1991]&~m[1992])|(m[831]&~m[1988]&m[1990]&m[1991]&~m[1992])|(~m[831]&m[1988]&~m[1990]&~m[1991]&m[1992])|(~m[831]&~m[1988]&m[1990]&~m[1991]&m[1992])|(m[831]&m[1988]&m[1990]&~m[1991]&m[1992])|(~m[831]&m[1988]&m[1990]&m[1991]&m[1992]))&UnbiasedRNG[708])|((m[831]&~m[1988]&~m[1990]&m[1991]&~m[1992])|(~m[831]&~m[1988]&~m[1990]&~m[1991]&m[1992])|(m[831]&~m[1988]&~m[1990]&~m[1991]&m[1992])|(m[831]&m[1988]&~m[1990]&~m[1991]&m[1992])|(m[831]&~m[1988]&m[1990]&~m[1991]&m[1992])|(~m[831]&~m[1988]&~m[1990]&m[1991]&m[1992])|(m[831]&~m[1988]&~m[1990]&m[1991]&m[1992])|(~m[831]&m[1988]&~m[1990]&m[1991]&m[1992])|(m[831]&m[1988]&~m[1990]&m[1991]&m[1992])|(~m[831]&~m[1988]&m[1990]&m[1991]&m[1992])|(m[831]&~m[1988]&m[1990]&m[1991]&m[1992])|(m[831]&m[1988]&m[1990]&m[1991]&m[1992]));
    m[1994] = (((m[846]&~m[1993]&~m[1995]&~m[1996]&~m[1997])|(~m[846]&~m[1993]&~m[1995]&m[1996]&~m[1997])|(m[846]&m[1993]&~m[1995]&m[1996]&~m[1997])|(m[846]&~m[1993]&m[1995]&m[1996]&~m[1997])|(~m[846]&m[1993]&~m[1995]&~m[1996]&m[1997])|(~m[846]&~m[1993]&m[1995]&~m[1996]&m[1997])|(m[846]&m[1993]&m[1995]&~m[1996]&m[1997])|(~m[846]&m[1993]&m[1995]&m[1996]&m[1997]))&UnbiasedRNG[709])|((m[846]&~m[1993]&~m[1995]&m[1996]&~m[1997])|(~m[846]&~m[1993]&~m[1995]&~m[1996]&m[1997])|(m[846]&~m[1993]&~m[1995]&~m[1996]&m[1997])|(m[846]&m[1993]&~m[1995]&~m[1996]&m[1997])|(m[846]&~m[1993]&m[1995]&~m[1996]&m[1997])|(~m[846]&~m[1993]&~m[1995]&m[1996]&m[1997])|(m[846]&~m[1993]&~m[1995]&m[1996]&m[1997])|(~m[846]&m[1993]&~m[1995]&m[1996]&m[1997])|(m[846]&m[1993]&~m[1995]&m[1996]&m[1997])|(~m[846]&~m[1993]&m[1995]&m[1996]&m[1997])|(m[846]&~m[1993]&m[1995]&m[1996]&m[1997])|(m[846]&m[1993]&m[1995]&m[1996]&m[1997]));
    m[1999] = (((m[861]&~m[1998]&~m[2000]&~m[2001]&~m[2002])|(~m[861]&~m[1998]&~m[2000]&m[2001]&~m[2002])|(m[861]&m[1998]&~m[2000]&m[2001]&~m[2002])|(m[861]&~m[1998]&m[2000]&m[2001]&~m[2002])|(~m[861]&m[1998]&~m[2000]&~m[2001]&m[2002])|(~m[861]&~m[1998]&m[2000]&~m[2001]&m[2002])|(m[861]&m[1998]&m[2000]&~m[2001]&m[2002])|(~m[861]&m[1998]&m[2000]&m[2001]&m[2002]))&UnbiasedRNG[710])|((m[861]&~m[1998]&~m[2000]&m[2001]&~m[2002])|(~m[861]&~m[1998]&~m[2000]&~m[2001]&m[2002])|(m[861]&~m[1998]&~m[2000]&~m[2001]&m[2002])|(m[861]&m[1998]&~m[2000]&~m[2001]&m[2002])|(m[861]&~m[1998]&m[2000]&~m[2001]&m[2002])|(~m[861]&~m[1998]&~m[2000]&m[2001]&m[2002])|(m[861]&~m[1998]&~m[2000]&m[2001]&m[2002])|(~m[861]&m[1998]&~m[2000]&m[2001]&m[2002])|(m[861]&m[1998]&~m[2000]&m[2001]&m[2002])|(~m[861]&~m[1998]&m[2000]&m[2001]&m[2002])|(m[861]&~m[1998]&m[2000]&m[2001]&m[2002])|(m[861]&m[1998]&m[2000]&m[2001]&m[2002]));
    m[2004] = (((m[876]&~m[2003]&~m[2005]&~m[2006]&~m[2007])|(~m[876]&~m[2003]&~m[2005]&m[2006]&~m[2007])|(m[876]&m[2003]&~m[2005]&m[2006]&~m[2007])|(m[876]&~m[2003]&m[2005]&m[2006]&~m[2007])|(~m[876]&m[2003]&~m[2005]&~m[2006]&m[2007])|(~m[876]&~m[2003]&m[2005]&~m[2006]&m[2007])|(m[876]&m[2003]&m[2005]&~m[2006]&m[2007])|(~m[876]&m[2003]&m[2005]&m[2006]&m[2007]))&UnbiasedRNG[711])|((m[876]&~m[2003]&~m[2005]&m[2006]&~m[2007])|(~m[876]&~m[2003]&~m[2005]&~m[2006]&m[2007])|(m[876]&~m[2003]&~m[2005]&~m[2006]&m[2007])|(m[876]&m[2003]&~m[2005]&~m[2006]&m[2007])|(m[876]&~m[2003]&m[2005]&~m[2006]&m[2007])|(~m[876]&~m[2003]&~m[2005]&m[2006]&m[2007])|(m[876]&~m[2003]&~m[2005]&m[2006]&m[2007])|(~m[876]&m[2003]&~m[2005]&m[2006]&m[2007])|(m[876]&m[2003]&~m[2005]&m[2006]&m[2007])|(~m[876]&~m[2003]&m[2005]&m[2006]&m[2007])|(m[876]&~m[2003]&m[2005]&m[2006]&m[2007])|(m[876]&m[2003]&m[2005]&m[2006]&m[2007]));
    m[2009] = (((m[891]&~m[2008]&~m[2010]&~m[2011]&~m[2012])|(~m[891]&~m[2008]&~m[2010]&m[2011]&~m[2012])|(m[891]&m[2008]&~m[2010]&m[2011]&~m[2012])|(m[891]&~m[2008]&m[2010]&m[2011]&~m[2012])|(~m[891]&m[2008]&~m[2010]&~m[2011]&m[2012])|(~m[891]&~m[2008]&m[2010]&~m[2011]&m[2012])|(m[891]&m[2008]&m[2010]&~m[2011]&m[2012])|(~m[891]&m[2008]&m[2010]&m[2011]&m[2012]))&UnbiasedRNG[712])|((m[891]&~m[2008]&~m[2010]&m[2011]&~m[2012])|(~m[891]&~m[2008]&~m[2010]&~m[2011]&m[2012])|(m[891]&~m[2008]&~m[2010]&~m[2011]&m[2012])|(m[891]&m[2008]&~m[2010]&~m[2011]&m[2012])|(m[891]&~m[2008]&m[2010]&~m[2011]&m[2012])|(~m[891]&~m[2008]&~m[2010]&m[2011]&m[2012])|(m[891]&~m[2008]&~m[2010]&m[2011]&m[2012])|(~m[891]&m[2008]&~m[2010]&m[2011]&m[2012])|(m[891]&m[2008]&~m[2010]&m[2011]&m[2012])|(~m[891]&~m[2008]&m[2010]&m[2011]&m[2012])|(m[891]&~m[2008]&m[2010]&m[2011]&m[2012])|(m[891]&m[2008]&m[2010]&m[2011]&m[2012]));
    m[2014] = (((m[906]&~m[2013]&~m[2015]&~m[2016]&~m[2017])|(~m[906]&~m[2013]&~m[2015]&m[2016]&~m[2017])|(m[906]&m[2013]&~m[2015]&m[2016]&~m[2017])|(m[906]&~m[2013]&m[2015]&m[2016]&~m[2017])|(~m[906]&m[2013]&~m[2015]&~m[2016]&m[2017])|(~m[906]&~m[2013]&m[2015]&~m[2016]&m[2017])|(m[906]&m[2013]&m[2015]&~m[2016]&m[2017])|(~m[906]&m[2013]&m[2015]&m[2016]&m[2017]))&UnbiasedRNG[713])|((m[906]&~m[2013]&~m[2015]&m[2016]&~m[2017])|(~m[906]&~m[2013]&~m[2015]&~m[2016]&m[2017])|(m[906]&~m[2013]&~m[2015]&~m[2016]&m[2017])|(m[906]&m[2013]&~m[2015]&~m[2016]&m[2017])|(m[906]&~m[2013]&m[2015]&~m[2016]&m[2017])|(~m[906]&~m[2013]&~m[2015]&m[2016]&m[2017])|(m[906]&~m[2013]&~m[2015]&m[2016]&m[2017])|(~m[906]&m[2013]&~m[2015]&m[2016]&m[2017])|(m[906]&m[2013]&~m[2015]&m[2016]&m[2017])|(~m[906]&~m[2013]&m[2015]&m[2016]&m[2017])|(m[906]&~m[2013]&m[2015]&m[2016]&m[2017])|(m[906]&m[2013]&m[2015]&m[2016]&m[2017]));
    m[2019] = (((m[921]&~m[2018]&~m[2020]&~m[2021]&~m[2022])|(~m[921]&~m[2018]&~m[2020]&m[2021]&~m[2022])|(m[921]&m[2018]&~m[2020]&m[2021]&~m[2022])|(m[921]&~m[2018]&m[2020]&m[2021]&~m[2022])|(~m[921]&m[2018]&~m[2020]&~m[2021]&m[2022])|(~m[921]&~m[2018]&m[2020]&~m[2021]&m[2022])|(m[921]&m[2018]&m[2020]&~m[2021]&m[2022])|(~m[921]&m[2018]&m[2020]&m[2021]&m[2022]))&UnbiasedRNG[714])|((m[921]&~m[2018]&~m[2020]&m[2021]&~m[2022])|(~m[921]&~m[2018]&~m[2020]&~m[2021]&m[2022])|(m[921]&~m[2018]&~m[2020]&~m[2021]&m[2022])|(m[921]&m[2018]&~m[2020]&~m[2021]&m[2022])|(m[921]&~m[2018]&m[2020]&~m[2021]&m[2022])|(~m[921]&~m[2018]&~m[2020]&m[2021]&m[2022])|(m[921]&~m[2018]&~m[2020]&m[2021]&m[2022])|(~m[921]&m[2018]&~m[2020]&m[2021]&m[2022])|(m[921]&m[2018]&~m[2020]&m[2021]&m[2022])|(~m[921]&~m[2018]&m[2020]&m[2021]&m[2022])|(m[921]&~m[2018]&m[2020]&m[2021]&m[2022])|(m[921]&m[2018]&m[2020]&m[2021]&m[2022]));
    m[2024] = (((m[847]&~m[2023]&~m[2025]&~m[2026]&~m[2027])|(~m[847]&~m[2023]&~m[2025]&m[2026]&~m[2027])|(m[847]&m[2023]&~m[2025]&m[2026]&~m[2027])|(m[847]&~m[2023]&m[2025]&m[2026]&~m[2027])|(~m[847]&m[2023]&~m[2025]&~m[2026]&m[2027])|(~m[847]&~m[2023]&m[2025]&~m[2026]&m[2027])|(m[847]&m[2023]&m[2025]&~m[2026]&m[2027])|(~m[847]&m[2023]&m[2025]&m[2026]&m[2027]))&UnbiasedRNG[715])|((m[847]&~m[2023]&~m[2025]&m[2026]&~m[2027])|(~m[847]&~m[2023]&~m[2025]&~m[2026]&m[2027])|(m[847]&~m[2023]&~m[2025]&~m[2026]&m[2027])|(m[847]&m[2023]&~m[2025]&~m[2026]&m[2027])|(m[847]&~m[2023]&m[2025]&~m[2026]&m[2027])|(~m[847]&~m[2023]&~m[2025]&m[2026]&m[2027])|(m[847]&~m[2023]&~m[2025]&m[2026]&m[2027])|(~m[847]&m[2023]&~m[2025]&m[2026]&m[2027])|(m[847]&m[2023]&~m[2025]&m[2026]&m[2027])|(~m[847]&~m[2023]&m[2025]&m[2026]&m[2027])|(m[847]&~m[2023]&m[2025]&m[2026]&m[2027])|(m[847]&m[2023]&m[2025]&m[2026]&m[2027]));
    m[2029] = (((m[862]&~m[2028]&~m[2030]&~m[2031]&~m[2032])|(~m[862]&~m[2028]&~m[2030]&m[2031]&~m[2032])|(m[862]&m[2028]&~m[2030]&m[2031]&~m[2032])|(m[862]&~m[2028]&m[2030]&m[2031]&~m[2032])|(~m[862]&m[2028]&~m[2030]&~m[2031]&m[2032])|(~m[862]&~m[2028]&m[2030]&~m[2031]&m[2032])|(m[862]&m[2028]&m[2030]&~m[2031]&m[2032])|(~m[862]&m[2028]&m[2030]&m[2031]&m[2032]))&UnbiasedRNG[716])|((m[862]&~m[2028]&~m[2030]&m[2031]&~m[2032])|(~m[862]&~m[2028]&~m[2030]&~m[2031]&m[2032])|(m[862]&~m[2028]&~m[2030]&~m[2031]&m[2032])|(m[862]&m[2028]&~m[2030]&~m[2031]&m[2032])|(m[862]&~m[2028]&m[2030]&~m[2031]&m[2032])|(~m[862]&~m[2028]&~m[2030]&m[2031]&m[2032])|(m[862]&~m[2028]&~m[2030]&m[2031]&m[2032])|(~m[862]&m[2028]&~m[2030]&m[2031]&m[2032])|(m[862]&m[2028]&~m[2030]&m[2031]&m[2032])|(~m[862]&~m[2028]&m[2030]&m[2031]&m[2032])|(m[862]&~m[2028]&m[2030]&m[2031]&m[2032])|(m[862]&m[2028]&m[2030]&m[2031]&m[2032]));
    m[2034] = (((m[877]&~m[2033]&~m[2035]&~m[2036]&~m[2037])|(~m[877]&~m[2033]&~m[2035]&m[2036]&~m[2037])|(m[877]&m[2033]&~m[2035]&m[2036]&~m[2037])|(m[877]&~m[2033]&m[2035]&m[2036]&~m[2037])|(~m[877]&m[2033]&~m[2035]&~m[2036]&m[2037])|(~m[877]&~m[2033]&m[2035]&~m[2036]&m[2037])|(m[877]&m[2033]&m[2035]&~m[2036]&m[2037])|(~m[877]&m[2033]&m[2035]&m[2036]&m[2037]))&UnbiasedRNG[717])|((m[877]&~m[2033]&~m[2035]&m[2036]&~m[2037])|(~m[877]&~m[2033]&~m[2035]&~m[2036]&m[2037])|(m[877]&~m[2033]&~m[2035]&~m[2036]&m[2037])|(m[877]&m[2033]&~m[2035]&~m[2036]&m[2037])|(m[877]&~m[2033]&m[2035]&~m[2036]&m[2037])|(~m[877]&~m[2033]&~m[2035]&m[2036]&m[2037])|(m[877]&~m[2033]&~m[2035]&m[2036]&m[2037])|(~m[877]&m[2033]&~m[2035]&m[2036]&m[2037])|(m[877]&m[2033]&~m[2035]&m[2036]&m[2037])|(~m[877]&~m[2033]&m[2035]&m[2036]&m[2037])|(m[877]&~m[2033]&m[2035]&m[2036]&m[2037])|(m[877]&m[2033]&m[2035]&m[2036]&m[2037]));
    m[2039] = (((m[892]&~m[2038]&~m[2040]&~m[2041]&~m[2042])|(~m[892]&~m[2038]&~m[2040]&m[2041]&~m[2042])|(m[892]&m[2038]&~m[2040]&m[2041]&~m[2042])|(m[892]&~m[2038]&m[2040]&m[2041]&~m[2042])|(~m[892]&m[2038]&~m[2040]&~m[2041]&m[2042])|(~m[892]&~m[2038]&m[2040]&~m[2041]&m[2042])|(m[892]&m[2038]&m[2040]&~m[2041]&m[2042])|(~m[892]&m[2038]&m[2040]&m[2041]&m[2042]))&UnbiasedRNG[718])|((m[892]&~m[2038]&~m[2040]&m[2041]&~m[2042])|(~m[892]&~m[2038]&~m[2040]&~m[2041]&m[2042])|(m[892]&~m[2038]&~m[2040]&~m[2041]&m[2042])|(m[892]&m[2038]&~m[2040]&~m[2041]&m[2042])|(m[892]&~m[2038]&m[2040]&~m[2041]&m[2042])|(~m[892]&~m[2038]&~m[2040]&m[2041]&m[2042])|(m[892]&~m[2038]&~m[2040]&m[2041]&m[2042])|(~m[892]&m[2038]&~m[2040]&m[2041]&m[2042])|(m[892]&m[2038]&~m[2040]&m[2041]&m[2042])|(~m[892]&~m[2038]&m[2040]&m[2041]&m[2042])|(m[892]&~m[2038]&m[2040]&m[2041]&m[2042])|(m[892]&m[2038]&m[2040]&m[2041]&m[2042]));
    m[2044] = (((m[907]&~m[2043]&~m[2045]&~m[2046]&~m[2047])|(~m[907]&~m[2043]&~m[2045]&m[2046]&~m[2047])|(m[907]&m[2043]&~m[2045]&m[2046]&~m[2047])|(m[907]&~m[2043]&m[2045]&m[2046]&~m[2047])|(~m[907]&m[2043]&~m[2045]&~m[2046]&m[2047])|(~m[907]&~m[2043]&m[2045]&~m[2046]&m[2047])|(m[907]&m[2043]&m[2045]&~m[2046]&m[2047])|(~m[907]&m[2043]&m[2045]&m[2046]&m[2047]))&UnbiasedRNG[719])|((m[907]&~m[2043]&~m[2045]&m[2046]&~m[2047])|(~m[907]&~m[2043]&~m[2045]&~m[2046]&m[2047])|(m[907]&~m[2043]&~m[2045]&~m[2046]&m[2047])|(m[907]&m[2043]&~m[2045]&~m[2046]&m[2047])|(m[907]&~m[2043]&m[2045]&~m[2046]&m[2047])|(~m[907]&~m[2043]&~m[2045]&m[2046]&m[2047])|(m[907]&~m[2043]&~m[2045]&m[2046]&m[2047])|(~m[907]&m[2043]&~m[2045]&m[2046]&m[2047])|(m[907]&m[2043]&~m[2045]&m[2046]&m[2047])|(~m[907]&~m[2043]&m[2045]&m[2046]&m[2047])|(m[907]&~m[2043]&m[2045]&m[2046]&m[2047])|(m[907]&m[2043]&m[2045]&m[2046]&m[2047]));
    m[2049] = (((m[922]&~m[2048]&~m[2050]&~m[2051]&~m[2052])|(~m[922]&~m[2048]&~m[2050]&m[2051]&~m[2052])|(m[922]&m[2048]&~m[2050]&m[2051]&~m[2052])|(m[922]&~m[2048]&m[2050]&m[2051]&~m[2052])|(~m[922]&m[2048]&~m[2050]&~m[2051]&m[2052])|(~m[922]&~m[2048]&m[2050]&~m[2051]&m[2052])|(m[922]&m[2048]&m[2050]&~m[2051]&m[2052])|(~m[922]&m[2048]&m[2050]&m[2051]&m[2052]))&UnbiasedRNG[720])|((m[922]&~m[2048]&~m[2050]&m[2051]&~m[2052])|(~m[922]&~m[2048]&~m[2050]&~m[2051]&m[2052])|(m[922]&~m[2048]&~m[2050]&~m[2051]&m[2052])|(m[922]&m[2048]&~m[2050]&~m[2051]&m[2052])|(m[922]&~m[2048]&m[2050]&~m[2051]&m[2052])|(~m[922]&~m[2048]&~m[2050]&m[2051]&m[2052])|(m[922]&~m[2048]&~m[2050]&m[2051]&m[2052])|(~m[922]&m[2048]&~m[2050]&m[2051]&m[2052])|(m[922]&m[2048]&~m[2050]&m[2051]&m[2052])|(~m[922]&~m[2048]&m[2050]&m[2051]&m[2052])|(m[922]&~m[2048]&m[2050]&m[2051]&m[2052])|(m[922]&m[2048]&m[2050]&m[2051]&m[2052]));
    m[2054] = (((m[863]&~m[2053]&~m[2055]&~m[2056]&~m[2057])|(~m[863]&~m[2053]&~m[2055]&m[2056]&~m[2057])|(m[863]&m[2053]&~m[2055]&m[2056]&~m[2057])|(m[863]&~m[2053]&m[2055]&m[2056]&~m[2057])|(~m[863]&m[2053]&~m[2055]&~m[2056]&m[2057])|(~m[863]&~m[2053]&m[2055]&~m[2056]&m[2057])|(m[863]&m[2053]&m[2055]&~m[2056]&m[2057])|(~m[863]&m[2053]&m[2055]&m[2056]&m[2057]))&UnbiasedRNG[721])|((m[863]&~m[2053]&~m[2055]&m[2056]&~m[2057])|(~m[863]&~m[2053]&~m[2055]&~m[2056]&m[2057])|(m[863]&~m[2053]&~m[2055]&~m[2056]&m[2057])|(m[863]&m[2053]&~m[2055]&~m[2056]&m[2057])|(m[863]&~m[2053]&m[2055]&~m[2056]&m[2057])|(~m[863]&~m[2053]&~m[2055]&m[2056]&m[2057])|(m[863]&~m[2053]&~m[2055]&m[2056]&m[2057])|(~m[863]&m[2053]&~m[2055]&m[2056]&m[2057])|(m[863]&m[2053]&~m[2055]&m[2056]&m[2057])|(~m[863]&~m[2053]&m[2055]&m[2056]&m[2057])|(m[863]&~m[2053]&m[2055]&m[2056]&m[2057])|(m[863]&m[2053]&m[2055]&m[2056]&m[2057]));
    m[2059] = (((m[878]&~m[2058]&~m[2060]&~m[2061]&~m[2062])|(~m[878]&~m[2058]&~m[2060]&m[2061]&~m[2062])|(m[878]&m[2058]&~m[2060]&m[2061]&~m[2062])|(m[878]&~m[2058]&m[2060]&m[2061]&~m[2062])|(~m[878]&m[2058]&~m[2060]&~m[2061]&m[2062])|(~m[878]&~m[2058]&m[2060]&~m[2061]&m[2062])|(m[878]&m[2058]&m[2060]&~m[2061]&m[2062])|(~m[878]&m[2058]&m[2060]&m[2061]&m[2062]))&UnbiasedRNG[722])|((m[878]&~m[2058]&~m[2060]&m[2061]&~m[2062])|(~m[878]&~m[2058]&~m[2060]&~m[2061]&m[2062])|(m[878]&~m[2058]&~m[2060]&~m[2061]&m[2062])|(m[878]&m[2058]&~m[2060]&~m[2061]&m[2062])|(m[878]&~m[2058]&m[2060]&~m[2061]&m[2062])|(~m[878]&~m[2058]&~m[2060]&m[2061]&m[2062])|(m[878]&~m[2058]&~m[2060]&m[2061]&m[2062])|(~m[878]&m[2058]&~m[2060]&m[2061]&m[2062])|(m[878]&m[2058]&~m[2060]&m[2061]&m[2062])|(~m[878]&~m[2058]&m[2060]&m[2061]&m[2062])|(m[878]&~m[2058]&m[2060]&m[2061]&m[2062])|(m[878]&m[2058]&m[2060]&m[2061]&m[2062]));
    m[2064] = (((m[893]&~m[2063]&~m[2065]&~m[2066]&~m[2067])|(~m[893]&~m[2063]&~m[2065]&m[2066]&~m[2067])|(m[893]&m[2063]&~m[2065]&m[2066]&~m[2067])|(m[893]&~m[2063]&m[2065]&m[2066]&~m[2067])|(~m[893]&m[2063]&~m[2065]&~m[2066]&m[2067])|(~m[893]&~m[2063]&m[2065]&~m[2066]&m[2067])|(m[893]&m[2063]&m[2065]&~m[2066]&m[2067])|(~m[893]&m[2063]&m[2065]&m[2066]&m[2067]))&UnbiasedRNG[723])|((m[893]&~m[2063]&~m[2065]&m[2066]&~m[2067])|(~m[893]&~m[2063]&~m[2065]&~m[2066]&m[2067])|(m[893]&~m[2063]&~m[2065]&~m[2066]&m[2067])|(m[893]&m[2063]&~m[2065]&~m[2066]&m[2067])|(m[893]&~m[2063]&m[2065]&~m[2066]&m[2067])|(~m[893]&~m[2063]&~m[2065]&m[2066]&m[2067])|(m[893]&~m[2063]&~m[2065]&m[2066]&m[2067])|(~m[893]&m[2063]&~m[2065]&m[2066]&m[2067])|(m[893]&m[2063]&~m[2065]&m[2066]&m[2067])|(~m[893]&~m[2063]&m[2065]&m[2066]&m[2067])|(m[893]&~m[2063]&m[2065]&m[2066]&m[2067])|(m[893]&m[2063]&m[2065]&m[2066]&m[2067]));
    m[2069] = (((m[908]&~m[2068]&~m[2070]&~m[2071]&~m[2072])|(~m[908]&~m[2068]&~m[2070]&m[2071]&~m[2072])|(m[908]&m[2068]&~m[2070]&m[2071]&~m[2072])|(m[908]&~m[2068]&m[2070]&m[2071]&~m[2072])|(~m[908]&m[2068]&~m[2070]&~m[2071]&m[2072])|(~m[908]&~m[2068]&m[2070]&~m[2071]&m[2072])|(m[908]&m[2068]&m[2070]&~m[2071]&m[2072])|(~m[908]&m[2068]&m[2070]&m[2071]&m[2072]))&UnbiasedRNG[724])|((m[908]&~m[2068]&~m[2070]&m[2071]&~m[2072])|(~m[908]&~m[2068]&~m[2070]&~m[2071]&m[2072])|(m[908]&~m[2068]&~m[2070]&~m[2071]&m[2072])|(m[908]&m[2068]&~m[2070]&~m[2071]&m[2072])|(m[908]&~m[2068]&m[2070]&~m[2071]&m[2072])|(~m[908]&~m[2068]&~m[2070]&m[2071]&m[2072])|(m[908]&~m[2068]&~m[2070]&m[2071]&m[2072])|(~m[908]&m[2068]&~m[2070]&m[2071]&m[2072])|(m[908]&m[2068]&~m[2070]&m[2071]&m[2072])|(~m[908]&~m[2068]&m[2070]&m[2071]&m[2072])|(m[908]&~m[2068]&m[2070]&m[2071]&m[2072])|(m[908]&m[2068]&m[2070]&m[2071]&m[2072]));
    m[2074] = (((m[923]&~m[2073]&~m[2075]&~m[2076]&~m[2077])|(~m[923]&~m[2073]&~m[2075]&m[2076]&~m[2077])|(m[923]&m[2073]&~m[2075]&m[2076]&~m[2077])|(m[923]&~m[2073]&m[2075]&m[2076]&~m[2077])|(~m[923]&m[2073]&~m[2075]&~m[2076]&m[2077])|(~m[923]&~m[2073]&m[2075]&~m[2076]&m[2077])|(m[923]&m[2073]&m[2075]&~m[2076]&m[2077])|(~m[923]&m[2073]&m[2075]&m[2076]&m[2077]))&UnbiasedRNG[725])|((m[923]&~m[2073]&~m[2075]&m[2076]&~m[2077])|(~m[923]&~m[2073]&~m[2075]&~m[2076]&m[2077])|(m[923]&~m[2073]&~m[2075]&~m[2076]&m[2077])|(m[923]&m[2073]&~m[2075]&~m[2076]&m[2077])|(m[923]&~m[2073]&m[2075]&~m[2076]&m[2077])|(~m[923]&~m[2073]&~m[2075]&m[2076]&m[2077])|(m[923]&~m[2073]&~m[2075]&m[2076]&m[2077])|(~m[923]&m[2073]&~m[2075]&m[2076]&m[2077])|(m[923]&m[2073]&~m[2075]&m[2076]&m[2077])|(~m[923]&~m[2073]&m[2075]&m[2076]&m[2077])|(m[923]&~m[2073]&m[2075]&m[2076]&m[2077])|(m[923]&m[2073]&m[2075]&m[2076]&m[2077]));
    m[2079] = (((m[879]&~m[2078]&~m[2080]&~m[2081]&~m[2082])|(~m[879]&~m[2078]&~m[2080]&m[2081]&~m[2082])|(m[879]&m[2078]&~m[2080]&m[2081]&~m[2082])|(m[879]&~m[2078]&m[2080]&m[2081]&~m[2082])|(~m[879]&m[2078]&~m[2080]&~m[2081]&m[2082])|(~m[879]&~m[2078]&m[2080]&~m[2081]&m[2082])|(m[879]&m[2078]&m[2080]&~m[2081]&m[2082])|(~m[879]&m[2078]&m[2080]&m[2081]&m[2082]))&UnbiasedRNG[726])|((m[879]&~m[2078]&~m[2080]&m[2081]&~m[2082])|(~m[879]&~m[2078]&~m[2080]&~m[2081]&m[2082])|(m[879]&~m[2078]&~m[2080]&~m[2081]&m[2082])|(m[879]&m[2078]&~m[2080]&~m[2081]&m[2082])|(m[879]&~m[2078]&m[2080]&~m[2081]&m[2082])|(~m[879]&~m[2078]&~m[2080]&m[2081]&m[2082])|(m[879]&~m[2078]&~m[2080]&m[2081]&m[2082])|(~m[879]&m[2078]&~m[2080]&m[2081]&m[2082])|(m[879]&m[2078]&~m[2080]&m[2081]&m[2082])|(~m[879]&~m[2078]&m[2080]&m[2081]&m[2082])|(m[879]&~m[2078]&m[2080]&m[2081]&m[2082])|(m[879]&m[2078]&m[2080]&m[2081]&m[2082]));
    m[2084] = (((m[894]&~m[2083]&~m[2085]&~m[2086]&~m[2087])|(~m[894]&~m[2083]&~m[2085]&m[2086]&~m[2087])|(m[894]&m[2083]&~m[2085]&m[2086]&~m[2087])|(m[894]&~m[2083]&m[2085]&m[2086]&~m[2087])|(~m[894]&m[2083]&~m[2085]&~m[2086]&m[2087])|(~m[894]&~m[2083]&m[2085]&~m[2086]&m[2087])|(m[894]&m[2083]&m[2085]&~m[2086]&m[2087])|(~m[894]&m[2083]&m[2085]&m[2086]&m[2087]))&UnbiasedRNG[727])|((m[894]&~m[2083]&~m[2085]&m[2086]&~m[2087])|(~m[894]&~m[2083]&~m[2085]&~m[2086]&m[2087])|(m[894]&~m[2083]&~m[2085]&~m[2086]&m[2087])|(m[894]&m[2083]&~m[2085]&~m[2086]&m[2087])|(m[894]&~m[2083]&m[2085]&~m[2086]&m[2087])|(~m[894]&~m[2083]&~m[2085]&m[2086]&m[2087])|(m[894]&~m[2083]&~m[2085]&m[2086]&m[2087])|(~m[894]&m[2083]&~m[2085]&m[2086]&m[2087])|(m[894]&m[2083]&~m[2085]&m[2086]&m[2087])|(~m[894]&~m[2083]&m[2085]&m[2086]&m[2087])|(m[894]&~m[2083]&m[2085]&m[2086]&m[2087])|(m[894]&m[2083]&m[2085]&m[2086]&m[2087]));
    m[2089] = (((m[909]&~m[2088]&~m[2090]&~m[2091]&~m[2092])|(~m[909]&~m[2088]&~m[2090]&m[2091]&~m[2092])|(m[909]&m[2088]&~m[2090]&m[2091]&~m[2092])|(m[909]&~m[2088]&m[2090]&m[2091]&~m[2092])|(~m[909]&m[2088]&~m[2090]&~m[2091]&m[2092])|(~m[909]&~m[2088]&m[2090]&~m[2091]&m[2092])|(m[909]&m[2088]&m[2090]&~m[2091]&m[2092])|(~m[909]&m[2088]&m[2090]&m[2091]&m[2092]))&UnbiasedRNG[728])|((m[909]&~m[2088]&~m[2090]&m[2091]&~m[2092])|(~m[909]&~m[2088]&~m[2090]&~m[2091]&m[2092])|(m[909]&~m[2088]&~m[2090]&~m[2091]&m[2092])|(m[909]&m[2088]&~m[2090]&~m[2091]&m[2092])|(m[909]&~m[2088]&m[2090]&~m[2091]&m[2092])|(~m[909]&~m[2088]&~m[2090]&m[2091]&m[2092])|(m[909]&~m[2088]&~m[2090]&m[2091]&m[2092])|(~m[909]&m[2088]&~m[2090]&m[2091]&m[2092])|(m[909]&m[2088]&~m[2090]&m[2091]&m[2092])|(~m[909]&~m[2088]&m[2090]&m[2091]&m[2092])|(m[909]&~m[2088]&m[2090]&m[2091]&m[2092])|(m[909]&m[2088]&m[2090]&m[2091]&m[2092]));
    m[2094] = (((m[924]&~m[2093]&~m[2095]&~m[2096]&~m[2097])|(~m[924]&~m[2093]&~m[2095]&m[2096]&~m[2097])|(m[924]&m[2093]&~m[2095]&m[2096]&~m[2097])|(m[924]&~m[2093]&m[2095]&m[2096]&~m[2097])|(~m[924]&m[2093]&~m[2095]&~m[2096]&m[2097])|(~m[924]&~m[2093]&m[2095]&~m[2096]&m[2097])|(m[924]&m[2093]&m[2095]&~m[2096]&m[2097])|(~m[924]&m[2093]&m[2095]&m[2096]&m[2097]))&UnbiasedRNG[729])|((m[924]&~m[2093]&~m[2095]&m[2096]&~m[2097])|(~m[924]&~m[2093]&~m[2095]&~m[2096]&m[2097])|(m[924]&~m[2093]&~m[2095]&~m[2096]&m[2097])|(m[924]&m[2093]&~m[2095]&~m[2096]&m[2097])|(m[924]&~m[2093]&m[2095]&~m[2096]&m[2097])|(~m[924]&~m[2093]&~m[2095]&m[2096]&m[2097])|(m[924]&~m[2093]&~m[2095]&m[2096]&m[2097])|(~m[924]&m[2093]&~m[2095]&m[2096]&m[2097])|(m[924]&m[2093]&~m[2095]&m[2096]&m[2097])|(~m[924]&~m[2093]&m[2095]&m[2096]&m[2097])|(m[924]&~m[2093]&m[2095]&m[2096]&m[2097])|(m[924]&m[2093]&m[2095]&m[2096]&m[2097]));
    m[2099] = (((m[895]&~m[2098]&~m[2100]&~m[2101]&~m[2102])|(~m[895]&~m[2098]&~m[2100]&m[2101]&~m[2102])|(m[895]&m[2098]&~m[2100]&m[2101]&~m[2102])|(m[895]&~m[2098]&m[2100]&m[2101]&~m[2102])|(~m[895]&m[2098]&~m[2100]&~m[2101]&m[2102])|(~m[895]&~m[2098]&m[2100]&~m[2101]&m[2102])|(m[895]&m[2098]&m[2100]&~m[2101]&m[2102])|(~m[895]&m[2098]&m[2100]&m[2101]&m[2102]))&UnbiasedRNG[730])|((m[895]&~m[2098]&~m[2100]&m[2101]&~m[2102])|(~m[895]&~m[2098]&~m[2100]&~m[2101]&m[2102])|(m[895]&~m[2098]&~m[2100]&~m[2101]&m[2102])|(m[895]&m[2098]&~m[2100]&~m[2101]&m[2102])|(m[895]&~m[2098]&m[2100]&~m[2101]&m[2102])|(~m[895]&~m[2098]&~m[2100]&m[2101]&m[2102])|(m[895]&~m[2098]&~m[2100]&m[2101]&m[2102])|(~m[895]&m[2098]&~m[2100]&m[2101]&m[2102])|(m[895]&m[2098]&~m[2100]&m[2101]&m[2102])|(~m[895]&~m[2098]&m[2100]&m[2101]&m[2102])|(m[895]&~m[2098]&m[2100]&m[2101]&m[2102])|(m[895]&m[2098]&m[2100]&m[2101]&m[2102]));
    m[2104] = (((m[910]&~m[2103]&~m[2105]&~m[2106]&~m[2107])|(~m[910]&~m[2103]&~m[2105]&m[2106]&~m[2107])|(m[910]&m[2103]&~m[2105]&m[2106]&~m[2107])|(m[910]&~m[2103]&m[2105]&m[2106]&~m[2107])|(~m[910]&m[2103]&~m[2105]&~m[2106]&m[2107])|(~m[910]&~m[2103]&m[2105]&~m[2106]&m[2107])|(m[910]&m[2103]&m[2105]&~m[2106]&m[2107])|(~m[910]&m[2103]&m[2105]&m[2106]&m[2107]))&UnbiasedRNG[731])|((m[910]&~m[2103]&~m[2105]&m[2106]&~m[2107])|(~m[910]&~m[2103]&~m[2105]&~m[2106]&m[2107])|(m[910]&~m[2103]&~m[2105]&~m[2106]&m[2107])|(m[910]&m[2103]&~m[2105]&~m[2106]&m[2107])|(m[910]&~m[2103]&m[2105]&~m[2106]&m[2107])|(~m[910]&~m[2103]&~m[2105]&m[2106]&m[2107])|(m[910]&~m[2103]&~m[2105]&m[2106]&m[2107])|(~m[910]&m[2103]&~m[2105]&m[2106]&m[2107])|(m[910]&m[2103]&~m[2105]&m[2106]&m[2107])|(~m[910]&~m[2103]&m[2105]&m[2106]&m[2107])|(m[910]&~m[2103]&m[2105]&m[2106]&m[2107])|(m[910]&m[2103]&m[2105]&m[2106]&m[2107]));
    m[2109] = (((m[925]&~m[2108]&~m[2110]&~m[2111]&~m[2112])|(~m[925]&~m[2108]&~m[2110]&m[2111]&~m[2112])|(m[925]&m[2108]&~m[2110]&m[2111]&~m[2112])|(m[925]&~m[2108]&m[2110]&m[2111]&~m[2112])|(~m[925]&m[2108]&~m[2110]&~m[2111]&m[2112])|(~m[925]&~m[2108]&m[2110]&~m[2111]&m[2112])|(m[925]&m[2108]&m[2110]&~m[2111]&m[2112])|(~m[925]&m[2108]&m[2110]&m[2111]&m[2112]))&UnbiasedRNG[732])|((m[925]&~m[2108]&~m[2110]&m[2111]&~m[2112])|(~m[925]&~m[2108]&~m[2110]&~m[2111]&m[2112])|(m[925]&~m[2108]&~m[2110]&~m[2111]&m[2112])|(m[925]&m[2108]&~m[2110]&~m[2111]&m[2112])|(m[925]&~m[2108]&m[2110]&~m[2111]&m[2112])|(~m[925]&~m[2108]&~m[2110]&m[2111]&m[2112])|(m[925]&~m[2108]&~m[2110]&m[2111]&m[2112])|(~m[925]&m[2108]&~m[2110]&m[2111]&m[2112])|(m[925]&m[2108]&~m[2110]&m[2111]&m[2112])|(~m[925]&~m[2108]&m[2110]&m[2111]&m[2112])|(m[925]&~m[2108]&m[2110]&m[2111]&m[2112])|(m[925]&m[2108]&m[2110]&m[2111]&m[2112]));
    m[2114] = (((m[911]&~m[2113]&~m[2115]&~m[2116]&~m[2117])|(~m[911]&~m[2113]&~m[2115]&m[2116]&~m[2117])|(m[911]&m[2113]&~m[2115]&m[2116]&~m[2117])|(m[911]&~m[2113]&m[2115]&m[2116]&~m[2117])|(~m[911]&m[2113]&~m[2115]&~m[2116]&m[2117])|(~m[911]&~m[2113]&m[2115]&~m[2116]&m[2117])|(m[911]&m[2113]&m[2115]&~m[2116]&m[2117])|(~m[911]&m[2113]&m[2115]&m[2116]&m[2117]))&UnbiasedRNG[733])|((m[911]&~m[2113]&~m[2115]&m[2116]&~m[2117])|(~m[911]&~m[2113]&~m[2115]&~m[2116]&m[2117])|(m[911]&~m[2113]&~m[2115]&~m[2116]&m[2117])|(m[911]&m[2113]&~m[2115]&~m[2116]&m[2117])|(m[911]&~m[2113]&m[2115]&~m[2116]&m[2117])|(~m[911]&~m[2113]&~m[2115]&m[2116]&m[2117])|(m[911]&~m[2113]&~m[2115]&m[2116]&m[2117])|(~m[911]&m[2113]&~m[2115]&m[2116]&m[2117])|(m[911]&m[2113]&~m[2115]&m[2116]&m[2117])|(~m[911]&~m[2113]&m[2115]&m[2116]&m[2117])|(m[911]&~m[2113]&m[2115]&m[2116]&m[2117])|(m[911]&m[2113]&m[2115]&m[2116]&m[2117]));
    m[2119] = (((m[926]&~m[2118]&~m[2120]&~m[2121]&~m[2122])|(~m[926]&~m[2118]&~m[2120]&m[2121]&~m[2122])|(m[926]&m[2118]&~m[2120]&m[2121]&~m[2122])|(m[926]&~m[2118]&m[2120]&m[2121]&~m[2122])|(~m[926]&m[2118]&~m[2120]&~m[2121]&m[2122])|(~m[926]&~m[2118]&m[2120]&~m[2121]&m[2122])|(m[926]&m[2118]&m[2120]&~m[2121]&m[2122])|(~m[926]&m[2118]&m[2120]&m[2121]&m[2122]))&UnbiasedRNG[734])|((m[926]&~m[2118]&~m[2120]&m[2121]&~m[2122])|(~m[926]&~m[2118]&~m[2120]&~m[2121]&m[2122])|(m[926]&~m[2118]&~m[2120]&~m[2121]&m[2122])|(m[926]&m[2118]&~m[2120]&~m[2121]&m[2122])|(m[926]&~m[2118]&m[2120]&~m[2121]&m[2122])|(~m[926]&~m[2118]&~m[2120]&m[2121]&m[2122])|(m[926]&~m[2118]&~m[2120]&m[2121]&m[2122])|(~m[926]&m[2118]&~m[2120]&m[2121]&m[2122])|(m[926]&m[2118]&~m[2120]&m[2121]&m[2122])|(~m[926]&~m[2118]&m[2120]&m[2121]&m[2122])|(m[926]&~m[2118]&m[2120]&m[2121]&m[2122])|(m[926]&m[2118]&m[2120]&m[2121]&m[2122]));
    m[2124] = (((m[927]&~m[2123]&~m[2125]&~m[2126]&~m[2127])|(~m[927]&~m[2123]&~m[2125]&m[2126]&~m[2127])|(m[927]&m[2123]&~m[2125]&m[2126]&~m[2127])|(m[927]&~m[2123]&m[2125]&m[2126]&~m[2127])|(~m[927]&m[2123]&~m[2125]&~m[2126]&m[2127])|(~m[927]&~m[2123]&m[2125]&~m[2126]&m[2127])|(m[927]&m[2123]&m[2125]&~m[2126]&m[2127])|(~m[927]&m[2123]&m[2125]&m[2126]&m[2127]))&UnbiasedRNG[735])|((m[927]&~m[2123]&~m[2125]&m[2126]&~m[2127])|(~m[927]&~m[2123]&~m[2125]&~m[2126]&m[2127])|(m[927]&~m[2123]&~m[2125]&~m[2126]&m[2127])|(m[927]&m[2123]&~m[2125]&~m[2126]&m[2127])|(m[927]&~m[2123]&m[2125]&~m[2126]&m[2127])|(~m[927]&~m[2123]&~m[2125]&m[2126]&m[2127])|(m[927]&~m[2123]&~m[2125]&m[2126]&m[2127])|(~m[927]&m[2123]&~m[2125]&m[2126]&m[2127])|(m[927]&m[2123]&~m[2125]&m[2126]&m[2127])|(~m[927]&~m[2123]&m[2125]&m[2126]&m[2127])|(m[927]&~m[2123]&m[2125]&m[2126]&m[2127])|(m[927]&m[2123]&m[2125]&m[2126]&m[2127]));
end

always @(posedge color3_clk) begin
    m[936] = (((m[933]&~m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&~m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&m[937]&~m[938])|(~m[933]&~m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&m[937]&m[938])|(m[933]&~m[934]&m[935]&m[937]&m[938])|(~m[933]&m[934]&m[935]&m[937]&m[938]))&UnbiasedRNG[736])|((m[933]&m[934]&~m[935]&~m[937]&~m[938])|(m[933]&~m[934]&m[935]&~m[937]&~m[938])|(~m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&~m[934]&~m[935]&~m[937]&m[938])|(~m[933]&m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&~m[937]&m[938])|(~m[933]&~m[934]&m[935]&~m[937]&m[938])|(m[933]&~m[934]&m[935]&~m[937]&m[938])|(~m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&m[937]&m[938]));
    m[946] = (((m[943]&~m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&~m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&m[947]&~m[948])|(~m[943]&~m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&m[947]&m[948])|(m[943]&~m[944]&m[945]&m[947]&m[948])|(~m[943]&m[944]&m[945]&m[947]&m[948]))&UnbiasedRNG[737])|((m[943]&m[944]&~m[945]&~m[947]&~m[948])|(m[943]&~m[944]&m[945]&~m[947]&~m[948])|(~m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&~m[944]&~m[945]&~m[947]&m[948])|(~m[943]&m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&~m[947]&m[948])|(~m[943]&~m[944]&m[945]&~m[947]&m[948])|(m[943]&~m[944]&m[945]&~m[947]&m[948])|(~m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&m[947]&m[948]));
    m[951] = (((m[948]&~m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&~m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&m[952]&~m[953])|(~m[948]&~m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&m[952]&m[953])|(m[948]&~m[949]&m[950]&m[952]&m[953])|(~m[948]&m[949]&m[950]&m[952]&m[953]))&UnbiasedRNG[738])|((m[948]&m[949]&~m[950]&~m[952]&~m[953])|(m[948]&~m[949]&m[950]&~m[952]&~m[953])|(~m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&~m[949]&~m[950]&~m[952]&m[953])|(~m[948]&m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&~m[952]&m[953])|(~m[948]&~m[949]&m[950]&~m[952]&m[953])|(m[948]&~m[949]&m[950]&~m[952]&m[953])|(~m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&m[952]&m[953]));
    m[961] = (((m[958]&~m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&~m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&m[962]&~m[963])|(~m[958]&~m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&m[962]&m[963])|(m[958]&~m[959]&m[960]&m[962]&m[963])|(~m[958]&m[959]&m[960]&m[962]&m[963]))&UnbiasedRNG[739])|((m[958]&m[959]&~m[960]&~m[962]&~m[963])|(m[958]&~m[959]&m[960]&~m[962]&~m[963])|(~m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&~m[959]&~m[960]&~m[962]&m[963])|(~m[958]&m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&~m[962]&m[963])|(~m[958]&~m[959]&m[960]&~m[962]&m[963])|(m[958]&~m[959]&m[960]&~m[962]&m[963])|(~m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&m[962]&m[963]));
    m[966] = (((m[963]&~m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&~m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&m[967]&~m[968])|(~m[963]&~m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&m[967]&m[968])|(m[963]&~m[964]&m[965]&m[967]&m[968])|(~m[963]&m[964]&m[965]&m[967]&m[968]))&UnbiasedRNG[740])|((m[963]&m[964]&~m[965]&~m[967]&~m[968])|(m[963]&~m[964]&m[965]&~m[967]&~m[968])|(~m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&~m[964]&~m[965]&~m[967]&m[968])|(~m[963]&m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&~m[967]&m[968])|(~m[963]&~m[964]&m[965]&~m[967]&m[968])|(m[963]&~m[964]&m[965]&~m[967]&m[968])|(~m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&m[967]&m[968]));
    m[971] = (((m[968]&~m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&~m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&m[972]&~m[973])|(~m[968]&~m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&m[972]&m[973])|(m[968]&~m[969]&m[970]&m[972]&m[973])|(~m[968]&m[969]&m[970]&m[972]&m[973]))&UnbiasedRNG[741])|((m[968]&m[969]&~m[970]&~m[972]&~m[973])|(m[968]&~m[969]&m[970]&~m[972]&~m[973])|(~m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&~m[969]&~m[970]&~m[972]&m[973])|(~m[968]&m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&~m[972]&m[973])|(~m[968]&~m[969]&m[970]&~m[972]&m[973])|(m[968]&~m[969]&m[970]&~m[972]&m[973])|(~m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&m[972]&m[973]));
    m[981] = (((m[978]&~m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&~m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&m[982]&~m[983])|(~m[978]&~m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&m[982]&m[983])|(m[978]&~m[979]&m[980]&m[982]&m[983])|(~m[978]&m[979]&m[980]&m[982]&m[983]))&UnbiasedRNG[742])|((m[978]&m[979]&~m[980]&~m[982]&~m[983])|(m[978]&~m[979]&m[980]&~m[982]&~m[983])|(~m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&~m[979]&~m[980]&~m[982]&m[983])|(~m[978]&m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&~m[982]&m[983])|(~m[978]&~m[979]&m[980]&~m[982]&m[983])|(m[978]&~m[979]&m[980]&~m[982]&m[983])|(~m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&m[982]&m[983]));
    m[986] = (((m[983]&~m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&~m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&m[987]&~m[988])|(~m[983]&~m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&m[987]&m[988])|(m[983]&~m[984]&m[985]&m[987]&m[988])|(~m[983]&m[984]&m[985]&m[987]&m[988]))&UnbiasedRNG[743])|((m[983]&m[984]&~m[985]&~m[987]&~m[988])|(m[983]&~m[984]&m[985]&~m[987]&~m[988])|(~m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&~m[984]&~m[985]&~m[987]&m[988])|(~m[983]&m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&~m[987]&m[988])|(~m[983]&~m[984]&m[985]&~m[987]&m[988])|(m[983]&~m[984]&m[985]&~m[987]&m[988])|(~m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&m[987]&m[988]));
    m[991] = (((m[988]&~m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&~m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&m[992]&~m[993])|(~m[988]&~m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&m[992]&m[993])|(m[988]&~m[989]&m[990]&m[992]&m[993])|(~m[988]&m[989]&m[990]&m[992]&m[993]))&UnbiasedRNG[744])|((m[988]&m[989]&~m[990]&~m[992]&~m[993])|(m[988]&~m[989]&m[990]&~m[992]&~m[993])|(~m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&~m[989]&~m[990]&~m[992]&m[993])|(~m[988]&m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&~m[992]&m[993])|(~m[988]&~m[989]&m[990]&~m[992]&m[993])|(m[988]&~m[989]&m[990]&~m[992]&m[993])|(~m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&m[992]&m[993]));
    m[996] = (((m[993]&~m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&~m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&m[997]&~m[998])|(~m[993]&~m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&m[997]&m[998])|(m[993]&~m[994]&m[995]&m[997]&m[998])|(~m[993]&m[994]&m[995]&m[997]&m[998]))&UnbiasedRNG[745])|((m[993]&m[994]&~m[995]&~m[997]&~m[998])|(m[993]&~m[994]&m[995]&~m[997]&~m[998])|(~m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&~m[994]&~m[995]&~m[997]&m[998])|(~m[993]&m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&~m[997]&m[998])|(~m[993]&~m[994]&m[995]&~m[997]&m[998])|(m[993]&~m[994]&m[995]&~m[997]&m[998])|(~m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&m[997]&m[998]));
    m[1006] = (((m[1003]&~m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&~m[1008])|(~m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&m[1007]&m[1008]))&UnbiasedRNG[746])|((m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&m[1008]));
    m[1011] = (((m[1008]&~m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&~m[1013])|(~m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))&UnbiasedRNG[747])|((m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&m[1013]));
    m[1016] = (((m[1013]&~m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&~m[1018])|(~m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))&UnbiasedRNG[748])|((m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&m[1018]));
    m[1021] = (((m[1018]&~m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&~m[1023])|(~m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))&UnbiasedRNG[749])|((m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&m[1023]));
    m[1026] = (((m[1023]&~m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&~m[1028])|(~m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))&UnbiasedRNG[750])|((m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&m[1028]));
    m[1036] = (((m[1033]&~m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&~m[1038])|(~m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))&UnbiasedRNG[751])|((m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&m[1038]));
    m[1041] = (((m[1038]&~m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&~m[1043])|(~m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))&UnbiasedRNG[752])|((m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&m[1043]));
    m[1046] = (((m[1043]&~m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&~m[1048])|(~m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&m[1047]&m[1048]))&UnbiasedRNG[753])|((m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&m[1048]));
    m[1051] = (((m[1048]&~m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&~m[1053])|(~m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))&UnbiasedRNG[754])|((m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&m[1053]));
    m[1056] = (((m[1053]&~m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&~m[1058])|(~m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&m[1057]&m[1058]))&UnbiasedRNG[755])|((m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&m[1058]));
    m[1061] = (((m[1058]&~m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&~m[1063])|(~m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))&UnbiasedRNG[756])|((m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&m[1063]));
    m[1071] = (((m[1068]&~m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&~m[1073])|(~m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))&UnbiasedRNG[757])|((m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&m[1073]));
    m[1076] = (((m[1073]&~m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&~m[1078])|(~m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))&UnbiasedRNG[758])|((m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&m[1078]));
    m[1081] = (((m[1078]&~m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&~m[1083])|(~m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&m[1082]&m[1083]))&UnbiasedRNG[759])|((m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&m[1083]));
    m[1086] = (((m[1083]&~m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&~m[1088])|(~m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))&UnbiasedRNG[760])|((m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&m[1088]));
    m[1091] = (((m[1088]&~m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&~m[1093])|(~m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))&UnbiasedRNG[761])|((m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&m[1093]));
    m[1096] = (((m[1093]&~m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&~m[1098])|(~m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))&UnbiasedRNG[762])|((m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&m[1098]));
    m[1101] = (((m[1098]&~m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&~m[1103])|(~m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))&UnbiasedRNG[763])|((m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&m[1103]));
    m[1111] = (((m[1108]&~m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&~m[1113])|(~m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&m[1112]&m[1113]))&UnbiasedRNG[764])|((m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&m[1113]));
    m[1116] = (((m[1113]&~m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&~m[1118])|(~m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&m[1117]&m[1118]))&UnbiasedRNG[765])|((m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&m[1118]));
    m[1121] = (((m[1118]&~m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&~m[1123])|(~m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))&UnbiasedRNG[766])|((m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&m[1123]));
    m[1126] = (((m[1123]&~m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&~m[1128])|(~m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))&UnbiasedRNG[767])|((m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&m[1128]));
    m[1131] = (((m[1128]&~m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&~m[1133])|(~m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))&UnbiasedRNG[768])|((m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&m[1133]));
    m[1136] = (((m[1133]&~m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&~m[1138])|(~m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&m[1137]&m[1138]))&UnbiasedRNG[769])|((m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&m[1138]));
    m[1141] = (((m[1138]&~m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&~m[1143])|(~m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))&UnbiasedRNG[770])|((m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&m[1143]));
    m[1146] = (((m[1143]&~m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&~m[1148])|(~m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))&UnbiasedRNG[771])|((m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&m[1148]));
    m[1156] = (((m[1153]&~m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&~m[1158])|(~m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&m[1157]&m[1158]))&UnbiasedRNG[772])|((m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&m[1158]));
    m[1161] = (((m[1158]&~m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&~m[1163])|(~m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))&UnbiasedRNG[773])|((m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&m[1163]));
    m[1166] = (((m[1163]&~m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&~m[1168])|(~m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))&UnbiasedRNG[774])|((m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&m[1168]));
    m[1171] = (((m[1168]&~m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&~m[1173])|(~m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&m[1172]&m[1173]))&UnbiasedRNG[775])|((m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&m[1173]));
    m[1176] = (((m[1173]&~m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&~m[1178])|(~m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))&UnbiasedRNG[776])|((m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&m[1178]));
    m[1181] = (((m[1178]&~m[1179]&~m[1180]&~m[1182]&~m[1183])|(~m[1178]&m[1179]&~m[1180]&~m[1182]&~m[1183])|(~m[1178]&~m[1179]&m[1180]&~m[1182]&~m[1183])|(m[1178]&m[1179]&m[1180]&m[1182]&~m[1183])|(~m[1178]&~m[1179]&~m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&~m[1180]&m[1182]&m[1183])|(m[1178]&~m[1179]&m[1180]&m[1182]&m[1183])|(~m[1178]&m[1179]&m[1180]&m[1182]&m[1183]))&UnbiasedRNG[777])|((m[1178]&m[1179]&~m[1180]&~m[1182]&~m[1183])|(m[1178]&~m[1179]&m[1180]&~m[1182]&~m[1183])|(~m[1178]&m[1179]&m[1180]&~m[1182]&~m[1183])|(m[1178]&m[1179]&m[1180]&~m[1182]&~m[1183])|(m[1178]&~m[1179]&~m[1180]&~m[1182]&m[1183])|(~m[1178]&m[1179]&~m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&~m[1180]&~m[1182]&m[1183])|(~m[1178]&~m[1179]&m[1180]&~m[1182]&m[1183])|(m[1178]&~m[1179]&m[1180]&~m[1182]&m[1183])|(~m[1178]&m[1179]&m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&m[1180]&m[1182]&m[1183]));
    m[1186] = (((m[1183]&~m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&~m[1188])|(~m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&m[1187]&m[1188]))&UnbiasedRNG[778])|((m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&m[1188]));
    m[1191] = (((m[1188]&~m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&~m[1193])|(~m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&m[1192]&m[1193]))&UnbiasedRNG[779])|((m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&m[1193]));
    m[1196] = (((m[1193]&~m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&~m[1198])|(~m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&m[1197]&m[1198]))&UnbiasedRNG[780])|((m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&m[1198]));
    m[1206] = (((m[1203]&~m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&~m[1208])|(~m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&m[1207]&m[1208]))&UnbiasedRNG[781])|((m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&m[1208]));
    m[1211] = (((m[1208]&~m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&~m[1213])|(~m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&m[1212]&m[1213]))&UnbiasedRNG[782])|((m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&m[1213]));
    m[1216] = (((m[1213]&~m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&~m[1218])|(~m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&m[1217]&m[1218]))&UnbiasedRNG[783])|((m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&m[1218]));
    m[1221] = (((m[1218]&~m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&~m[1223])|(~m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&m[1222]&m[1223]))&UnbiasedRNG[784])|((m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&m[1223]));
    m[1226] = (((m[1223]&~m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&~m[1228])|(~m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&m[1227]&m[1228]))&UnbiasedRNG[785])|((m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&m[1228]));
    m[1231] = (((m[1228]&~m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&~m[1233])|(~m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&m[1232]&m[1233]))&UnbiasedRNG[786])|((m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&m[1233]));
    m[1236] = (((m[1233]&~m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&~m[1238])|(~m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&m[1237]&m[1238]))&UnbiasedRNG[787])|((m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&m[1238]));
    m[1241] = (((m[1238]&~m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&~m[1243])|(~m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&m[1242]&m[1243]))&UnbiasedRNG[788])|((m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&m[1243]));
    m[1246] = (((m[1243]&~m[1244]&~m[1245]&~m[1247]&~m[1248])|(~m[1243]&m[1244]&~m[1245]&~m[1247]&~m[1248])|(~m[1243]&~m[1244]&m[1245]&~m[1247]&~m[1248])|(m[1243]&m[1244]&m[1245]&m[1247]&~m[1248])|(~m[1243]&~m[1244]&~m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&~m[1245]&m[1247]&m[1248])|(m[1243]&~m[1244]&m[1245]&m[1247]&m[1248])|(~m[1243]&m[1244]&m[1245]&m[1247]&m[1248]))&UnbiasedRNG[789])|((m[1243]&m[1244]&~m[1245]&~m[1247]&~m[1248])|(m[1243]&~m[1244]&m[1245]&~m[1247]&~m[1248])|(~m[1243]&m[1244]&m[1245]&~m[1247]&~m[1248])|(m[1243]&m[1244]&m[1245]&~m[1247]&~m[1248])|(m[1243]&~m[1244]&~m[1245]&~m[1247]&m[1248])|(~m[1243]&m[1244]&~m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&~m[1245]&~m[1247]&m[1248])|(~m[1243]&~m[1244]&m[1245]&~m[1247]&m[1248])|(m[1243]&~m[1244]&m[1245]&~m[1247]&m[1248])|(~m[1243]&m[1244]&m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&m[1245]&m[1247]&m[1248]));
    m[1251] = (((m[1248]&~m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&~m[1253])|(~m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&m[1252]&m[1253]))&UnbiasedRNG[790])|((m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&m[1253]));
    m[1261] = (((m[1258]&~m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&~m[1263])|(~m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&m[1262]&m[1263]))&UnbiasedRNG[791])|((m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&m[1263]));
    m[1266] = (((m[1263]&~m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&~m[1268])|(~m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&m[1267]&m[1268]))&UnbiasedRNG[792])|((m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&m[1268]));
    m[1271] = (((m[1268]&~m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&~m[1273])|(~m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&m[1272]&m[1273]))&UnbiasedRNG[793])|((m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&m[1273]));
    m[1276] = (((m[1273]&~m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&~m[1278])|(~m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&m[1277]&m[1278]))&UnbiasedRNG[794])|((m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&m[1278]));
    m[1281] = (((m[1278]&~m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&~m[1283])|(~m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&m[1282]&m[1283]))&UnbiasedRNG[795])|((m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&m[1283]));
    m[1286] = (((m[1283]&~m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&~m[1288])|(~m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&m[1287]&m[1288]))&UnbiasedRNG[796])|((m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&m[1288]));
    m[1291] = (((m[1288]&~m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&~m[1293])|(~m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&m[1292]&m[1293]))&UnbiasedRNG[797])|((m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&m[1293]));
    m[1296] = (((m[1293]&~m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&~m[1298])|(~m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&m[1297]&m[1298]))&UnbiasedRNG[798])|((m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&m[1298]));
    m[1301] = (((m[1298]&~m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&~m[1303])|(~m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&m[1302]&m[1303]))&UnbiasedRNG[799])|((m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&m[1303]));
    m[1306] = (((m[1303]&~m[1304]&~m[1305]&~m[1307]&~m[1308])|(~m[1303]&m[1304]&~m[1305]&~m[1307]&~m[1308])|(~m[1303]&~m[1304]&m[1305]&~m[1307]&~m[1308])|(m[1303]&m[1304]&m[1305]&m[1307]&~m[1308])|(~m[1303]&~m[1304]&~m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&~m[1305]&m[1307]&m[1308])|(m[1303]&~m[1304]&m[1305]&m[1307]&m[1308])|(~m[1303]&m[1304]&m[1305]&m[1307]&m[1308]))&UnbiasedRNG[800])|((m[1303]&m[1304]&~m[1305]&~m[1307]&~m[1308])|(m[1303]&~m[1304]&m[1305]&~m[1307]&~m[1308])|(~m[1303]&m[1304]&m[1305]&~m[1307]&~m[1308])|(m[1303]&m[1304]&m[1305]&~m[1307]&~m[1308])|(m[1303]&~m[1304]&~m[1305]&~m[1307]&m[1308])|(~m[1303]&m[1304]&~m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&~m[1305]&~m[1307]&m[1308])|(~m[1303]&~m[1304]&m[1305]&~m[1307]&m[1308])|(m[1303]&~m[1304]&m[1305]&~m[1307]&m[1308])|(~m[1303]&m[1304]&m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&m[1305]&m[1307]&m[1308]));
    m[1311] = (((m[1308]&~m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&~m[1313])|(~m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&m[1312]&m[1313]))&UnbiasedRNG[801])|((m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&m[1313]));
    m[1321] = (((m[1318]&~m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&~m[1323])|(~m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&m[1322]&m[1323]))&UnbiasedRNG[802])|((m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&m[1323]));
    m[1326] = (((m[1323]&~m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&~m[1328])|(~m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&m[1327]&m[1328]))&UnbiasedRNG[803])|((m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&m[1328]));
    m[1331] = (((m[1328]&~m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&~m[1333])|(~m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&m[1332]&m[1333]))&UnbiasedRNG[804])|((m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&m[1333]));
    m[1336] = (((m[1333]&~m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&~m[1338])|(~m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&m[1337]&m[1338]))&UnbiasedRNG[805])|((m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&m[1338]));
    m[1341] = (((m[1338]&~m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&~m[1343])|(~m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&m[1342]&m[1343]))&UnbiasedRNG[806])|((m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&m[1343]));
    m[1346] = (((m[1343]&~m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&~m[1348])|(~m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&m[1347]&m[1348]))&UnbiasedRNG[807])|((m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&m[1348]));
    m[1351] = (((m[1348]&~m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&~m[1353])|(~m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&m[1352]&m[1353]))&UnbiasedRNG[808])|((m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&m[1353]));
    m[1356] = (((m[1353]&~m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&~m[1358])|(~m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&m[1357]&m[1358]))&UnbiasedRNG[809])|((m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&m[1358]));
    m[1361] = (((m[1358]&~m[1359]&~m[1360]&~m[1362]&~m[1363])|(~m[1358]&m[1359]&~m[1360]&~m[1362]&~m[1363])|(~m[1358]&~m[1359]&m[1360]&~m[1362]&~m[1363])|(m[1358]&m[1359]&m[1360]&m[1362]&~m[1363])|(~m[1358]&~m[1359]&~m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&~m[1360]&m[1362]&m[1363])|(m[1358]&~m[1359]&m[1360]&m[1362]&m[1363])|(~m[1358]&m[1359]&m[1360]&m[1362]&m[1363]))&UnbiasedRNG[810])|((m[1358]&m[1359]&~m[1360]&~m[1362]&~m[1363])|(m[1358]&~m[1359]&m[1360]&~m[1362]&~m[1363])|(~m[1358]&m[1359]&m[1360]&~m[1362]&~m[1363])|(m[1358]&m[1359]&m[1360]&~m[1362]&~m[1363])|(m[1358]&~m[1359]&~m[1360]&~m[1362]&m[1363])|(~m[1358]&m[1359]&~m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&~m[1360]&~m[1362]&m[1363])|(~m[1358]&~m[1359]&m[1360]&~m[1362]&m[1363])|(m[1358]&~m[1359]&m[1360]&~m[1362]&m[1363])|(~m[1358]&m[1359]&m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&m[1360]&m[1362]&m[1363]));
    m[1366] = (((m[1363]&~m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&~m[1368])|(~m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&m[1367]&m[1368]))&UnbiasedRNG[811])|((m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&m[1368]));
    m[1371] = (((m[1368]&~m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&~m[1373])|(~m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&m[1372]&m[1373]))&UnbiasedRNG[812])|((m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&m[1373]));
    m[1376] = (((m[1373]&~m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&~m[1378])|(~m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&m[1377]&m[1378]))&UnbiasedRNG[813])|((m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&m[1378]));
    m[1386] = (((m[1383]&~m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&~m[1388])|(~m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&m[1387]&m[1388]))&UnbiasedRNG[814])|((m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&m[1388]));
    m[1391] = (((m[1388]&~m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&~m[1393])|(~m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&m[1392]&m[1393]))&UnbiasedRNG[815])|((m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&m[1393]));
    m[1396] = (((m[1393]&~m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&~m[1398])|(~m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&m[1397]&m[1398]))&UnbiasedRNG[816])|((m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&m[1398]));
    m[1401] = (((m[1398]&~m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&~m[1403])|(~m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&m[1402]&m[1403]))&UnbiasedRNG[817])|((m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&m[1403]));
    m[1406] = (((m[1403]&~m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&~m[1408])|(~m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&m[1407]&m[1408]))&UnbiasedRNG[818])|((m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&m[1408]));
    m[1411] = (((m[1408]&~m[1409]&~m[1410]&~m[1412]&~m[1413])|(~m[1408]&m[1409]&~m[1410]&~m[1412]&~m[1413])|(~m[1408]&~m[1409]&m[1410]&~m[1412]&~m[1413])|(m[1408]&m[1409]&m[1410]&m[1412]&~m[1413])|(~m[1408]&~m[1409]&~m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&~m[1410]&m[1412]&m[1413])|(m[1408]&~m[1409]&m[1410]&m[1412]&m[1413])|(~m[1408]&m[1409]&m[1410]&m[1412]&m[1413]))&UnbiasedRNG[819])|((m[1408]&m[1409]&~m[1410]&~m[1412]&~m[1413])|(m[1408]&~m[1409]&m[1410]&~m[1412]&~m[1413])|(~m[1408]&m[1409]&m[1410]&~m[1412]&~m[1413])|(m[1408]&m[1409]&m[1410]&~m[1412]&~m[1413])|(m[1408]&~m[1409]&~m[1410]&~m[1412]&m[1413])|(~m[1408]&m[1409]&~m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&~m[1410]&~m[1412]&m[1413])|(~m[1408]&~m[1409]&m[1410]&~m[1412]&m[1413])|(m[1408]&~m[1409]&m[1410]&~m[1412]&m[1413])|(~m[1408]&m[1409]&m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&m[1410]&m[1412]&m[1413]));
    m[1416] = (((m[1413]&~m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&~m[1418])|(~m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&m[1417]&m[1418]))&UnbiasedRNG[820])|((m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&m[1418]));
    m[1421] = (((m[1418]&~m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&~m[1423])|(~m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&m[1422]&m[1423]))&UnbiasedRNG[821])|((m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&m[1423]));
    m[1426] = (((m[1423]&~m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&~m[1428])|(~m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&m[1427]&m[1428]))&UnbiasedRNG[822])|((m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&m[1428]));
    m[1431] = (((m[1428]&~m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&~m[1433])|(~m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&m[1432]&m[1433]))&UnbiasedRNG[823])|((m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&m[1433]));
    m[1436] = (((m[1433]&~m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&~m[1438])|(~m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&m[1437]&m[1438]))&UnbiasedRNG[824])|((m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&m[1438]));
    m[1441] = (((m[1438]&~m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&~m[1443])|(~m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&m[1442]&m[1443]))&UnbiasedRNG[825])|((m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&m[1443]));
    m[1446] = (((m[1443]&~m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&~m[1448])|(~m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&m[1447]&m[1448]))&UnbiasedRNG[826])|((m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&m[1448]));
    m[1456] = (((m[1453]&~m[1454]&~m[1455]&~m[1457]&~m[1458])|(~m[1453]&m[1454]&~m[1455]&~m[1457]&~m[1458])|(~m[1453]&~m[1454]&m[1455]&~m[1457]&~m[1458])|(m[1453]&m[1454]&m[1455]&m[1457]&~m[1458])|(~m[1453]&~m[1454]&~m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&~m[1455]&m[1457]&m[1458])|(m[1453]&~m[1454]&m[1455]&m[1457]&m[1458])|(~m[1453]&m[1454]&m[1455]&m[1457]&m[1458]))&UnbiasedRNG[827])|((m[1453]&m[1454]&~m[1455]&~m[1457]&~m[1458])|(m[1453]&~m[1454]&m[1455]&~m[1457]&~m[1458])|(~m[1453]&m[1454]&m[1455]&~m[1457]&~m[1458])|(m[1453]&m[1454]&m[1455]&~m[1457]&~m[1458])|(m[1453]&~m[1454]&~m[1455]&~m[1457]&m[1458])|(~m[1453]&m[1454]&~m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&~m[1455]&~m[1457]&m[1458])|(~m[1453]&~m[1454]&m[1455]&~m[1457]&m[1458])|(m[1453]&~m[1454]&m[1455]&~m[1457]&m[1458])|(~m[1453]&m[1454]&m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&m[1455]&m[1457]&m[1458]));
    m[1461] = (((m[1458]&~m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&~m[1463])|(~m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&m[1462]&m[1463]))&UnbiasedRNG[828])|((m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&m[1463]));
    m[1466] = (((m[1463]&~m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&~m[1468])|(~m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&m[1467]&m[1468]))&UnbiasedRNG[829])|((m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&m[1468]));
    m[1471] = (((m[1468]&~m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&~m[1473])|(~m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&m[1472]&m[1473]))&UnbiasedRNG[830])|((m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&m[1473]));
    m[1476] = (((m[1473]&~m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&~m[1478])|(~m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&m[1477]&m[1478]))&UnbiasedRNG[831])|((m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&m[1478]));
    m[1481] = (((m[1478]&~m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&~m[1483])|(~m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&m[1482]&m[1483]))&UnbiasedRNG[832])|((m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&m[1483]));
    m[1486] = (((m[1483]&~m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&~m[1488])|(~m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&m[1487]&m[1488]))&UnbiasedRNG[833])|((m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&m[1488]));
    m[1491] = (((m[1488]&~m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&~m[1493])|(~m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&m[1492]&m[1493]))&UnbiasedRNG[834])|((m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&m[1493]));
    m[1496] = (((m[1493]&~m[1494]&~m[1495]&~m[1497]&~m[1498])|(~m[1493]&m[1494]&~m[1495]&~m[1497]&~m[1498])|(~m[1493]&~m[1494]&m[1495]&~m[1497]&~m[1498])|(m[1493]&m[1494]&m[1495]&m[1497]&~m[1498])|(~m[1493]&~m[1494]&~m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&~m[1495]&m[1497]&m[1498])|(m[1493]&~m[1494]&m[1495]&m[1497]&m[1498])|(~m[1493]&m[1494]&m[1495]&m[1497]&m[1498]))&UnbiasedRNG[835])|((m[1493]&m[1494]&~m[1495]&~m[1497]&~m[1498])|(m[1493]&~m[1494]&m[1495]&~m[1497]&~m[1498])|(~m[1493]&m[1494]&m[1495]&~m[1497]&~m[1498])|(m[1493]&m[1494]&m[1495]&~m[1497]&~m[1498])|(m[1493]&~m[1494]&~m[1495]&~m[1497]&m[1498])|(~m[1493]&m[1494]&~m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&~m[1495]&~m[1497]&m[1498])|(~m[1493]&~m[1494]&m[1495]&~m[1497]&m[1498])|(m[1493]&~m[1494]&m[1495]&~m[1497]&m[1498])|(~m[1493]&m[1494]&m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&m[1495]&m[1497]&m[1498]));
    m[1501] = (((m[1498]&~m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&~m[1503])|(~m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&m[1502]&m[1503]))&UnbiasedRNG[836])|((m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&m[1503]));
    m[1506] = (((m[1503]&~m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&~m[1508])|(~m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&m[1507]&m[1508]))&UnbiasedRNG[837])|((m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&m[1508]));
    m[1511] = (((m[1508]&~m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&~m[1513])|(~m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&m[1512]&m[1513]))&UnbiasedRNG[838])|((m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&m[1513]));
    m[1516] = (((m[1513]&~m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&~m[1518])|(~m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&m[1517]&m[1518]))&UnbiasedRNG[839])|((m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&m[1518]));
    m[1521] = (((m[1518]&~m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&~m[1523])|(~m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&m[1522]&m[1523]))&UnbiasedRNG[840])|((m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&m[1523]));
    m[1531] = (((m[1528]&~m[1529]&~m[1530]&~m[1532]&~m[1533])|(~m[1528]&m[1529]&~m[1530]&~m[1532]&~m[1533])|(~m[1528]&~m[1529]&m[1530]&~m[1532]&~m[1533])|(m[1528]&m[1529]&m[1530]&m[1532]&~m[1533])|(~m[1528]&~m[1529]&~m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&~m[1530]&m[1532]&m[1533])|(m[1528]&~m[1529]&m[1530]&m[1532]&m[1533])|(~m[1528]&m[1529]&m[1530]&m[1532]&m[1533]))&UnbiasedRNG[841])|((m[1528]&m[1529]&~m[1530]&~m[1532]&~m[1533])|(m[1528]&~m[1529]&m[1530]&~m[1532]&~m[1533])|(~m[1528]&m[1529]&m[1530]&~m[1532]&~m[1533])|(m[1528]&m[1529]&m[1530]&~m[1532]&~m[1533])|(m[1528]&~m[1529]&~m[1530]&~m[1532]&m[1533])|(~m[1528]&m[1529]&~m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&~m[1530]&~m[1532]&m[1533])|(~m[1528]&~m[1529]&m[1530]&~m[1532]&m[1533])|(m[1528]&~m[1529]&m[1530]&~m[1532]&m[1533])|(~m[1528]&m[1529]&m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&m[1530]&m[1532]&m[1533]));
    m[1536] = (((m[1533]&~m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&~m[1538])|(~m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&m[1537]&m[1538]))&UnbiasedRNG[842])|((m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&m[1538]));
    m[1541] = (((m[1538]&~m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&~m[1543])|(~m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&m[1542]&m[1543]))&UnbiasedRNG[843])|((m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&m[1543]));
    m[1546] = (((m[1543]&~m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&~m[1548])|(~m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&m[1547]&m[1548]))&UnbiasedRNG[844])|((m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&m[1548]));
    m[1551] = (((m[1548]&~m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&~m[1553])|(~m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&m[1552]&m[1553]))&UnbiasedRNG[845])|((m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&m[1553]));
    m[1556] = (((m[1553]&~m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&~m[1558])|(~m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&m[1557]&m[1558]))&UnbiasedRNG[846])|((m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&m[1558]));
    m[1561] = (((m[1558]&~m[1559]&~m[1560]&~m[1562]&~m[1563])|(~m[1558]&m[1559]&~m[1560]&~m[1562]&~m[1563])|(~m[1558]&~m[1559]&m[1560]&~m[1562]&~m[1563])|(m[1558]&m[1559]&m[1560]&m[1562]&~m[1563])|(~m[1558]&~m[1559]&~m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&~m[1560]&m[1562]&m[1563])|(m[1558]&~m[1559]&m[1560]&m[1562]&m[1563])|(~m[1558]&m[1559]&m[1560]&m[1562]&m[1563]))&UnbiasedRNG[847])|((m[1558]&m[1559]&~m[1560]&~m[1562]&~m[1563])|(m[1558]&~m[1559]&m[1560]&~m[1562]&~m[1563])|(~m[1558]&m[1559]&m[1560]&~m[1562]&~m[1563])|(m[1558]&m[1559]&m[1560]&~m[1562]&~m[1563])|(m[1558]&~m[1559]&~m[1560]&~m[1562]&m[1563])|(~m[1558]&m[1559]&~m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&~m[1560]&~m[1562]&m[1563])|(~m[1558]&~m[1559]&m[1560]&~m[1562]&m[1563])|(m[1558]&~m[1559]&m[1560]&~m[1562]&m[1563])|(~m[1558]&m[1559]&m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&m[1560]&m[1562]&m[1563]));
    m[1566] = (((m[1563]&~m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&~m[1568])|(~m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&m[1567]&m[1568]))&UnbiasedRNG[848])|((m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&m[1568]));
    m[1571] = (((m[1568]&~m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&~m[1573])|(~m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&m[1572]&m[1573]))&UnbiasedRNG[849])|((m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&m[1573]));
    m[1576] = (((m[1573]&~m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&~m[1578])|(~m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&m[1577]&m[1578]))&UnbiasedRNG[850])|((m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&m[1578]));
    m[1581] = (((m[1578]&~m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&~m[1583])|(~m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&m[1582]&m[1583]))&UnbiasedRNG[851])|((m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&m[1583]));
    m[1586] = (((m[1583]&~m[1584]&~m[1585]&~m[1587]&~m[1588])|(~m[1583]&m[1584]&~m[1585]&~m[1587]&~m[1588])|(~m[1583]&~m[1584]&m[1585]&~m[1587]&~m[1588])|(m[1583]&m[1584]&m[1585]&m[1587]&~m[1588])|(~m[1583]&~m[1584]&~m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&~m[1585]&m[1587]&m[1588])|(m[1583]&~m[1584]&m[1585]&m[1587]&m[1588])|(~m[1583]&m[1584]&m[1585]&m[1587]&m[1588]))&UnbiasedRNG[852])|((m[1583]&m[1584]&~m[1585]&~m[1587]&~m[1588])|(m[1583]&~m[1584]&m[1585]&~m[1587]&~m[1588])|(~m[1583]&m[1584]&m[1585]&~m[1587]&~m[1588])|(m[1583]&m[1584]&m[1585]&~m[1587]&~m[1588])|(m[1583]&~m[1584]&~m[1585]&~m[1587]&m[1588])|(~m[1583]&m[1584]&~m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&~m[1585]&~m[1587]&m[1588])|(~m[1583]&~m[1584]&m[1585]&~m[1587]&m[1588])|(m[1583]&~m[1584]&m[1585]&~m[1587]&m[1588])|(~m[1583]&m[1584]&m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&m[1585]&m[1587]&m[1588]));
    m[1591] = (((m[1588]&~m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&~m[1593])|(~m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&m[1592]&m[1593]))&UnbiasedRNG[853])|((m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&m[1593]));
    m[1596] = (((m[1593]&~m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&~m[1598])|(~m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&m[1597]&m[1598]))&UnbiasedRNG[854])|((m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&m[1598]));
    m[1606] = (((m[1603]&~m[1604]&~m[1605]&~m[1607]&~m[1608])|(~m[1603]&m[1604]&~m[1605]&~m[1607]&~m[1608])|(~m[1603]&~m[1604]&m[1605]&~m[1607]&~m[1608])|(m[1603]&m[1604]&m[1605]&m[1607]&~m[1608])|(~m[1603]&~m[1604]&~m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&~m[1605]&m[1607]&m[1608])|(m[1603]&~m[1604]&m[1605]&m[1607]&m[1608])|(~m[1603]&m[1604]&m[1605]&m[1607]&m[1608]))&UnbiasedRNG[855])|((m[1603]&m[1604]&~m[1605]&~m[1607]&~m[1608])|(m[1603]&~m[1604]&m[1605]&~m[1607]&~m[1608])|(~m[1603]&m[1604]&m[1605]&~m[1607]&~m[1608])|(m[1603]&m[1604]&m[1605]&~m[1607]&~m[1608])|(m[1603]&~m[1604]&~m[1605]&~m[1607]&m[1608])|(~m[1603]&m[1604]&~m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&~m[1605]&~m[1607]&m[1608])|(~m[1603]&~m[1604]&m[1605]&~m[1607]&m[1608])|(m[1603]&~m[1604]&m[1605]&~m[1607]&m[1608])|(~m[1603]&m[1604]&m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&m[1605]&m[1607]&m[1608]));
    m[1611] = (((m[1608]&~m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&~m[1613])|(~m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&m[1612]&m[1613]))&UnbiasedRNG[856])|((m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&m[1613]));
    m[1616] = (((m[1613]&~m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&~m[1618])|(~m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&m[1617]&m[1618]))&UnbiasedRNG[857])|((m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&m[1618]));
    m[1621] = (((m[1618]&~m[1619]&~m[1620]&~m[1622]&~m[1623])|(~m[1618]&m[1619]&~m[1620]&~m[1622]&~m[1623])|(~m[1618]&~m[1619]&m[1620]&~m[1622]&~m[1623])|(m[1618]&m[1619]&m[1620]&m[1622]&~m[1623])|(~m[1618]&~m[1619]&~m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&~m[1620]&m[1622]&m[1623])|(m[1618]&~m[1619]&m[1620]&m[1622]&m[1623])|(~m[1618]&m[1619]&m[1620]&m[1622]&m[1623]))&UnbiasedRNG[858])|((m[1618]&m[1619]&~m[1620]&~m[1622]&~m[1623])|(m[1618]&~m[1619]&m[1620]&~m[1622]&~m[1623])|(~m[1618]&m[1619]&m[1620]&~m[1622]&~m[1623])|(m[1618]&m[1619]&m[1620]&~m[1622]&~m[1623])|(m[1618]&~m[1619]&~m[1620]&~m[1622]&m[1623])|(~m[1618]&m[1619]&~m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&~m[1620]&~m[1622]&m[1623])|(~m[1618]&~m[1619]&m[1620]&~m[1622]&m[1623])|(m[1618]&~m[1619]&m[1620]&~m[1622]&m[1623])|(~m[1618]&m[1619]&m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&m[1620]&m[1622]&m[1623]));
    m[1626] = (((m[1623]&~m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&~m[1628])|(~m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&m[1627]&m[1628]))&UnbiasedRNG[859])|((m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&m[1628]));
    m[1631] = (((m[1628]&~m[1629]&~m[1630]&~m[1632]&~m[1633])|(~m[1628]&m[1629]&~m[1630]&~m[1632]&~m[1633])|(~m[1628]&~m[1629]&m[1630]&~m[1632]&~m[1633])|(m[1628]&m[1629]&m[1630]&m[1632]&~m[1633])|(~m[1628]&~m[1629]&~m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&~m[1630]&m[1632]&m[1633])|(m[1628]&~m[1629]&m[1630]&m[1632]&m[1633])|(~m[1628]&m[1629]&m[1630]&m[1632]&m[1633]))&UnbiasedRNG[860])|((m[1628]&m[1629]&~m[1630]&~m[1632]&~m[1633])|(m[1628]&~m[1629]&m[1630]&~m[1632]&~m[1633])|(~m[1628]&m[1629]&m[1630]&~m[1632]&~m[1633])|(m[1628]&m[1629]&m[1630]&~m[1632]&~m[1633])|(m[1628]&~m[1629]&~m[1630]&~m[1632]&m[1633])|(~m[1628]&m[1629]&~m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&~m[1630]&~m[1632]&m[1633])|(~m[1628]&~m[1629]&m[1630]&~m[1632]&m[1633])|(m[1628]&~m[1629]&m[1630]&~m[1632]&m[1633])|(~m[1628]&m[1629]&m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&m[1630]&m[1632]&m[1633]));
    m[1636] = (((m[1633]&~m[1634]&~m[1635]&~m[1637]&~m[1638])|(~m[1633]&m[1634]&~m[1635]&~m[1637]&~m[1638])|(~m[1633]&~m[1634]&m[1635]&~m[1637]&~m[1638])|(m[1633]&m[1634]&m[1635]&m[1637]&~m[1638])|(~m[1633]&~m[1634]&~m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&~m[1635]&m[1637]&m[1638])|(m[1633]&~m[1634]&m[1635]&m[1637]&m[1638])|(~m[1633]&m[1634]&m[1635]&m[1637]&m[1638]))&UnbiasedRNG[861])|((m[1633]&m[1634]&~m[1635]&~m[1637]&~m[1638])|(m[1633]&~m[1634]&m[1635]&~m[1637]&~m[1638])|(~m[1633]&m[1634]&m[1635]&~m[1637]&~m[1638])|(m[1633]&m[1634]&m[1635]&~m[1637]&~m[1638])|(m[1633]&~m[1634]&~m[1635]&~m[1637]&m[1638])|(~m[1633]&m[1634]&~m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&~m[1635]&~m[1637]&m[1638])|(~m[1633]&~m[1634]&m[1635]&~m[1637]&m[1638])|(m[1633]&~m[1634]&m[1635]&~m[1637]&m[1638])|(~m[1633]&m[1634]&m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&m[1635]&m[1637]&m[1638]));
    m[1641] = (((m[1638]&~m[1639]&~m[1640]&~m[1642]&~m[1643])|(~m[1638]&m[1639]&~m[1640]&~m[1642]&~m[1643])|(~m[1638]&~m[1639]&m[1640]&~m[1642]&~m[1643])|(m[1638]&m[1639]&m[1640]&m[1642]&~m[1643])|(~m[1638]&~m[1639]&~m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&~m[1640]&m[1642]&m[1643])|(m[1638]&~m[1639]&m[1640]&m[1642]&m[1643])|(~m[1638]&m[1639]&m[1640]&m[1642]&m[1643]))&UnbiasedRNG[862])|((m[1638]&m[1639]&~m[1640]&~m[1642]&~m[1643])|(m[1638]&~m[1639]&m[1640]&~m[1642]&~m[1643])|(~m[1638]&m[1639]&m[1640]&~m[1642]&~m[1643])|(m[1638]&m[1639]&m[1640]&~m[1642]&~m[1643])|(m[1638]&~m[1639]&~m[1640]&~m[1642]&m[1643])|(~m[1638]&m[1639]&~m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&~m[1640]&~m[1642]&m[1643])|(~m[1638]&~m[1639]&m[1640]&~m[1642]&m[1643])|(m[1638]&~m[1639]&m[1640]&~m[1642]&m[1643])|(~m[1638]&m[1639]&m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&m[1640]&m[1642]&m[1643]));
    m[1646] = (((m[1643]&~m[1644]&~m[1645]&~m[1647]&~m[1648])|(~m[1643]&m[1644]&~m[1645]&~m[1647]&~m[1648])|(~m[1643]&~m[1644]&m[1645]&~m[1647]&~m[1648])|(m[1643]&m[1644]&m[1645]&m[1647]&~m[1648])|(~m[1643]&~m[1644]&~m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&~m[1645]&m[1647]&m[1648])|(m[1643]&~m[1644]&m[1645]&m[1647]&m[1648])|(~m[1643]&m[1644]&m[1645]&m[1647]&m[1648]))&UnbiasedRNG[863])|((m[1643]&m[1644]&~m[1645]&~m[1647]&~m[1648])|(m[1643]&~m[1644]&m[1645]&~m[1647]&~m[1648])|(~m[1643]&m[1644]&m[1645]&~m[1647]&~m[1648])|(m[1643]&m[1644]&m[1645]&~m[1647]&~m[1648])|(m[1643]&~m[1644]&~m[1645]&~m[1647]&m[1648])|(~m[1643]&m[1644]&~m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&~m[1645]&~m[1647]&m[1648])|(~m[1643]&~m[1644]&m[1645]&~m[1647]&m[1648])|(m[1643]&~m[1644]&m[1645]&~m[1647]&m[1648])|(~m[1643]&m[1644]&m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&m[1645]&m[1647]&m[1648]));
    m[1651] = (((m[1648]&~m[1649]&~m[1650]&~m[1652]&~m[1653])|(~m[1648]&m[1649]&~m[1650]&~m[1652]&~m[1653])|(~m[1648]&~m[1649]&m[1650]&~m[1652]&~m[1653])|(m[1648]&m[1649]&m[1650]&m[1652]&~m[1653])|(~m[1648]&~m[1649]&~m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&~m[1650]&m[1652]&m[1653])|(m[1648]&~m[1649]&m[1650]&m[1652]&m[1653])|(~m[1648]&m[1649]&m[1650]&m[1652]&m[1653]))&UnbiasedRNG[864])|((m[1648]&m[1649]&~m[1650]&~m[1652]&~m[1653])|(m[1648]&~m[1649]&m[1650]&~m[1652]&~m[1653])|(~m[1648]&m[1649]&m[1650]&~m[1652]&~m[1653])|(m[1648]&m[1649]&m[1650]&~m[1652]&~m[1653])|(m[1648]&~m[1649]&~m[1650]&~m[1652]&m[1653])|(~m[1648]&m[1649]&~m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&~m[1650]&~m[1652]&m[1653])|(~m[1648]&~m[1649]&m[1650]&~m[1652]&m[1653])|(m[1648]&~m[1649]&m[1650]&~m[1652]&m[1653])|(~m[1648]&m[1649]&m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&m[1650]&m[1652]&m[1653]));
    m[1656] = (((m[1653]&~m[1654]&~m[1655]&~m[1657]&~m[1658])|(~m[1653]&m[1654]&~m[1655]&~m[1657]&~m[1658])|(~m[1653]&~m[1654]&m[1655]&~m[1657]&~m[1658])|(m[1653]&m[1654]&m[1655]&m[1657]&~m[1658])|(~m[1653]&~m[1654]&~m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&~m[1655]&m[1657]&m[1658])|(m[1653]&~m[1654]&m[1655]&m[1657]&m[1658])|(~m[1653]&m[1654]&m[1655]&m[1657]&m[1658]))&UnbiasedRNG[865])|((m[1653]&m[1654]&~m[1655]&~m[1657]&~m[1658])|(m[1653]&~m[1654]&m[1655]&~m[1657]&~m[1658])|(~m[1653]&m[1654]&m[1655]&~m[1657]&~m[1658])|(m[1653]&m[1654]&m[1655]&~m[1657]&~m[1658])|(m[1653]&~m[1654]&~m[1655]&~m[1657]&m[1658])|(~m[1653]&m[1654]&~m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&~m[1655]&~m[1657]&m[1658])|(~m[1653]&~m[1654]&m[1655]&~m[1657]&m[1658])|(m[1653]&~m[1654]&m[1655]&~m[1657]&m[1658])|(~m[1653]&m[1654]&m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&m[1655]&m[1657]&m[1658]));
    m[1661] = (((m[1658]&~m[1659]&~m[1660]&~m[1662]&~m[1663])|(~m[1658]&m[1659]&~m[1660]&~m[1662]&~m[1663])|(~m[1658]&~m[1659]&m[1660]&~m[1662]&~m[1663])|(m[1658]&m[1659]&m[1660]&m[1662]&~m[1663])|(~m[1658]&~m[1659]&~m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&~m[1660]&m[1662]&m[1663])|(m[1658]&~m[1659]&m[1660]&m[1662]&m[1663])|(~m[1658]&m[1659]&m[1660]&m[1662]&m[1663]))&UnbiasedRNG[866])|((m[1658]&m[1659]&~m[1660]&~m[1662]&~m[1663])|(m[1658]&~m[1659]&m[1660]&~m[1662]&~m[1663])|(~m[1658]&m[1659]&m[1660]&~m[1662]&~m[1663])|(m[1658]&m[1659]&m[1660]&~m[1662]&~m[1663])|(m[1658]&~m[1659]&~m[1660]&~m[1662]&m[1663])|(~m[1658]&m[1659]&~m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&~m[1660]&~m[1662]&m[1663])|(~m[1658]&~m[1659]&m[1660]&~m[1662]&m[1663])|(m[1658]&~m[1659]&m[1660]&~m[1662]&m[1663])|(~m[1658]&m[1659]&m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&m[1660]&m[1662]&m[1663]));
    m[1666] = (((m[1663]&~m[1664]&~m[1665]&~m[1667]&~m[1668])|(~m[1663]&m[1664]&~m[1665]&~m[1667]&~m[1668])|(~m[1663]&~m[1664]&m[1665]&~m[1667]&~m[1668])|(m[1663]&m[1664]&m[1665]&m[1667]&~m[1668])|(~m[1663]&~m[1664]&~m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&~m[1665]&m[1667]&m[1668])|(m[1663]&~m[1664]&m[1665]&m[1667]&m[1668])|(~m[1663]&m[1664]&m[1665]&m[1667]&m[1668]))&UnbiasedRNG[867])|((m[1663]&m[1664]&~m[1665]&~m[1667]&~m[1668])|(m[1663]&~m[1664]&m[1665]&~m[1667]&~m[1668])|(~m[1663]&m[1664]&m[1665]&~m[1667]&~m[1668])|(m[1663]&m[1664]&m[1665]&~m[1667]&~m[1668])|(m[1663]&~m[1664]&~m[1665]&~m[1667]&m[1668])|(~m[1663]&m[1664]&~m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&~m[1665]&~m[1667]&m[1668])|(~m[1663]&~m[1664]&m[1665]&~m[1667]&m[1668])|(m[1663]&~m[1664]&m[1665]&~m[1667]&m[1668])|(~m[1663]&m[1664]&m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&m[1665]&m[1667]&m[1668]));
    m[1676] = (((m[1673]&~m[1674]&~m[1675]&~m[1677]&~m[1678])|(~m[1673]&m[1674]&~m[1675]&~m[1677]&~m[1678])|(~m[1673]&~m[1674]&m[1675]&~m[1677]&~m[1678])|(m[1673]&m[1674]&m[1675]&m[1677]&~m[1678])|(~m[1673]&~m[1674]&~m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&~m[1675]&m[1677]&m[1678])|(m[1673]&~m[1674]&m[1675]&m[1677]&m[1678])|(~m[1673]&m[1674]&m[1675]&m[1677]&m[1678]))&UnbiasedRNG[868])|((m[1673]&m[1674]&~m[1675]&~m[1677]&~m[1678])|(m[1673]&~m[1674]&m[1675]&~m[1677]&~m[1678])|(~m[1673]&m[1674]&m[1675]&~m[1677]&~m[1678])|(m[1673]&m[1674]&m[1675]&~m[1677]&~m[1678])|(m[1673]&~m[1674]&~m[1675]&~m[1677]&m[1678])|(~m[1673]&m[1674]&~m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&~m[1675]&~m[1677]&m[1678])|(~m[1673]&~m[1674]&m[1675]&~m[1677]&m[1678])|(m[1673]&~m[1674]&m[1675]&~m[1677]&m[1678])|(~m[1673]&m[1674]&m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&m[1675]&m[1677]&m[1678]));
    m[1681] = (((m[1678]&~m[1679]&~m[1680]&~m[1682]&~m[1683])|(~m[1678]&m[1679]&~m[1680]&~m[1682]&~m[1683])|(~m[1678]&~m[1679]&m[1680]&~m[1682]&~m[1683])|(m[1678]&m[1679]&m[1680]&m[1682]&~m[1683])|(~m[1678]&~m[1679]&~m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&~m[1680]&m[1682]&m[1683])|(m[1678]&~m[1679]&m[1680]&m[1682]&m[1683])|(~m[1678]&m[1679]&m[1680]&m[1682]&m[1683]))&UnbiasedRNG[869])|((m[1678]&m[1679]&~m[1680]&~m[1682]&~m[1683])|(m[1678]&~m[1679]&m[1680]&~m[1682]&~m[1683])|(~m[1678]&m[1679]&m[1680]&~m[1682]&~m[1683])|(m[1678]&m[1679]&m[1680]&~m[1682]&~m[1683])|(m[1678]&~m[1679]&~m[1680]&~m[1682]&m[1683])|(~m[1678]&m[1679]&~m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&~m[1680]&~m[1682]&m[1683])|(~m[1678]&~m[1679]&m[1680]&~m[1682]&m[1683])|(m[1678]&~m[1679]&m[1680]&~m[1682]&m[1683])|(~m[1678]&m[1679]&m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&m[1680]&m[1682]&m[1683]));
    m[1686] = (((m[1683]&~m[1684]&~m[1685]&~m[1687]&~m[1688])|(~m[1683]&m[1684]&~m[1685]&~m[1687]&~m[1688])|(~m[1683]&~m[1684]&m[1685]&~m[1687]&~m[1688])|(m[1683]&m[1684]&m[1685]&m[1687]&~m[1688])|(~m[1683]&~m[1684]&~m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&~m[1685]&m[1687]&m[1688])|(m[1683]&~m[1684]&m[1685]&m[1687]&m[1688])|(~m[1683]&m[1684]&m[1685]&m[1687]&m[1688]))&UnbiasedRNG[870])|((m[1683]&m[1684]&~m[1685]&~m[1687]&~m[1688])|(m[1683]&~m[1684]&m[1685]&~m[1687]&~m[1688])|(~m[1683]&m[1684]&m[1685]&~m[1687]&~m[1688])|(m[1683]&m[1684]&m[1685]&~m[1687]&~m[1688])|(m[1683]&~m[1684]&~m[1685]&~m[1687]&m[1688])|(~m[1683]&m[1684]&~m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&~m[1685]&~m[1687]&m[1688])|(~m[1683]&~m[1684]&m[1685]&~m[1687]&m[1688])|(m[1683]&~m[1684]&m[1685]&~m[1687]&m[1688])|(~m[1683]&m[1684]&m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&m[1685]&m[1687]&m[1688]));
    m[1691] = (((m[1688]&~m[1689]&~m[1690]&~m[1692]&~m[1693])|(~m[1688]&m[1689]&~m[1690]&~m[1692]&~m[1693])|(~m[1688]&~m[1689]&m[1690]&~m[1692]&~m[1693])|(m[1688]&m[1689]&m[1690]&m[1692]&~m[1693])|(~m[1688]&~m[1689]&~m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&~m[1690]&m[1692]&m[1693])|(m[1688]&~m[1689]&m[1690]&m[1692]&m[1693])|(~m[1688]&m[1689]&m[1690]&m[1692]&m[1693]))&UnbiasedRNG[871])|((m[1688]&m[1689]&~m[1690]&~m[1692]&~m[1693])|(m[1688]&~m[1689]&m[1690]&~m[1692]&~m[1693])|(~m[1688]&m[1689]&m[1690]&~m[1692]&~m[1693])|(m[1688]&m[1689]&m[1690]&~m[1692]&~m[1693])|(m[1688]&~m[1689]&~m[1690]&~m[1692]&m[1693])|(~m[1688]&m[1689]&~m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&~m[1690]&~m[1692]&m[1693])|(~m[1688]&~m[1689]&m[1690]&~m[1692]&m[1693])|(m[1688]&~m[1689]&m[1690]&~m[1692]&m[1693])|(~m[1688]&m[1689]&m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&m[1690]&m[1692]&m[1693]));
    m[1696] = (((m[1693]&~m[1694]&~m[1695]&~m[1697]&~m[1698])|(~m[1693]&m[1694]&~m[1695]&~m[1697]&~m[1698])|(~m[1693]&~m[1694]&m[1695]&~m[1697]&~m[1698])|(m[1693]&m[1694]&m[1695]&m[1697]&~m[1698])|(~m[1693]&~m[1694]&~m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&~m[1695]&m[1697]&m[1698])|(m[1693]&~m[1694]&m[1695]&m[1697]&m[1698])|(~m[1693]&m[1694]&m[1695]&m[1697]&m[1698]))&UnbiasedRNG[872])|((m[1693]&m[1694]&~m[1695]&~m[1697]&~m[1698])|(m[1693]&~m[1694]&m[1695]&~m[1697]&~m[1698])|(~m[1693]&m[1694]&m[1695]&~m[1697]&~m[1698])|(m[1693]&m[1694]&m[1695]&~m[1697]&~m[1698])|(m[1693]&~m[1694]&~m[1695]&~m[1697]&m[1698])|(~m[1693]&m[1694]&~m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&~m[1695]&~m[1697]&m[1698])|(~m[1693]&~m[1694]&m[1695]&~m[1697]&m[1698])|(m[1693]&~m[1694]&m[1695]&~m[1697]&m[1698])|(~m[1693]&m[1694]&m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&m[1695]&m[1697]&m[1698]));
    m[1701] = (((m[1698]&~m[1699]&~m[1700]&~m[1702]&~m[1703])|(~m[1698]&m[1699]&~m[1700]&~m[1702]&~m[1703])|(~m[1698]&~m[1699]&m[1700]&~m[1702]&~m[1703])|(m[1698]&m[1699]&m[1700]&m[1702]&~m[1703])|(~m[1698]&~m[1699]&~m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&~m[1700]&m[1702]&m[1703])|(m[1698]&~m[1699]&m[1700]&m[1702]&m[1703])|(~m[1698]&m[1699]&m[1700]&m[1702]&m[1703]))&UnbiasedRNG[873])|((m[1698]&m[1699]&~m[1700]&~m[1702]&~m[1703])|(m[1698]&~m[1699]&m[1700]&~m[1702]&~m[1703])|(~m[1698]&m[1699]&m[1700]&~m[1702]&~m[1703])|(m[1698]&m[1699]&m[1700]&~m[1702]&~m[1703])|(m[1698]&~m[1699]&~m[1700]&~m[1702]&m[1703])|(~m[1698]&m[1699]&~m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&~m[1700]&~m[1702]&m[1703])|(~m[1698]&~m[1699]&m[1700]&~m[1702]&m[1703])|(m[1698]&~m[1699]&m[1700]&~m[1702]&m[1703])|(~m[1698]&m[1699]&m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&m[1700]&m[1702]&m[1703]));
    m[1706] = (((m[1703]&~m[1704]&~m[1705]&~m[1707]&~m[1708])|(~m[1703]&m[1704]&~m[1705]&~m[1707]&~m[1708])|(~m[1703]&~m[1704]&m[1705]&~m[1707]&~m[1708])|(m[1703]&m[1704]&m[1705]&m[1707]&~m[1708])|(~m[1703]&~m[1704]&~m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&~m[1705]&m[1707]&m[1708])|(m[1703]&~m[1704]&m[1705]&m[1707]&m[1708])|(~m[1703]&m[1704]&m[1705]&m[1707]&m[1708]))&UnbiasedRNG[874])|((m[1703]&m[1704]&~m[1705]&~m[1707]&~m[1708])|(m[1703]&~m[1704]&m[1705]&~m[1707]&~m[1708])|(~m[1703]&m[1704]&m[1705]&~m[1707]&~m[1708])|(m[1703]&m[1704]&m[1705]&~m[1707]&~m[1708])|(m[1703]&~m[1704]&~m[1705]&~m[1707]&m[1708])|(~m[1703]&m[1704]&~m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&~m[1705]&~m[1707]&m[1708])|(~m[1703]&~m[1704]&m[1705]&~m[1707]&m[1708])|(m[1703]&~m[1704]&m[1705]&~m[1707]&m[1708])|(~m[1703]&m[1704]&m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&m[1705]&m[1707]&m[1708]));
    m[1711] = (((m[1708]&~m[1709]&~m[1710]&~m[1712]&~m[1713])|(~m[1708]&m[1709]&~m[1710]&~m[1712]&~m[1713])|(~m[1708]&~m[1709]&m[1710]&~m[1712]&~m[1713])|(m[1708]&m[1709]&m[1710]&m[1712]&~m[1713])|(~m[1708]&~m[1709]&~m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&~m[1710]&m[1712]&m[1713])|(m[1708]&~m[1709]&m[1710]&m[1712]&m[1713])|(~m[1708]&m[1709]&m[1710]&m[1712]&m[1713]))&UnbiasedRNG[875])|((m[1708]&m[1709]&~m[1710]&~m[1712]&~m[1713])|(m[1708]&~m[1709]&m[1710]&~m[1712]&~m[1713])|(~m[1708]&m[1709]&m[1710]&~m[1712]&~m[1713])|(m[1708]&m[1709]&m[1710]&~m[1712]&~m[1713])|(m[1708]&~m[1709]&~m[1710]&~m[1712]&m[1713])|(~m[1708]&m[1709]&~m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&~m[1710]&~m[1712]&m[1713])|(~m[1708]&~m[1709]&m[1710]&~m[1712]&m[1713])|(m[1708]&~m[1709]&m[1710]&~m[1712]&m[1713])|(~m[1708]&m[1709]&m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&m[1710]&m[1712]&m[1713]));
    m[1716] = (((m[1713]&~m[1714]&~m[1715]&~m[1717]&~m[1718])|(~m[1713]&m[1714]&~m[1715]&~m[1717]&~m[1718])|(~m[1713]&~m[1714]&m[1715]&~m[1717]&~m[1718])|(m[1713]&m[1714]&m[1715]&m[1717]&~m[1718])|(~m[1713]&~m[1714]&~m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&~m[1715]&m[1717]&m[1718])|(m[1713]&~m[1714]&m[1715]&m[1717]&m[1718])|(~m[1713]&m[1714]&m[1715]&m[1717]&m[1718]))&UnbiasedRNG[876])|((m[1713]&m[1714]&~m[1715]&~m[1717]&~m[1718])|(m[1713]&~m[1714]&m[1715]&~m[1717]&~m[1718])|(~m[1713]&m[1714]&m[1715]&~m[1717]&~m[1718])|(m[1713]&m[1714]&m[1715]&~m[1717]&~m[1718])|(m[1713]&~m[1714]&~m[1715]&~m[1717]&m[1718])|(~m[1713]&m[1714]&~m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&~m[1715]&~m[1717]&m[1718])|(~m[1713]&~m[1714]&m[1715]&~m[1717]&m[1718])|(m[1713]&~m[1714]&m[1715]&~m[1717]&m[1718])|(~m[1713]&m[1714]&m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&m[1715]&m[1717]&m[1718]));
    m[1721] = (((m[1718]&~m[1719]&~m[1720]&~m[1722]&~m[1723])|(~m[1718]&m[1719]&~m[1720]&~m[1722]&~m[1723])|(~m[1718]&~m[1719]&m[1720]&~m[1722]&~m[1723])|(m[1718]&m[1719]&m[1720]&m[1722]&~m[1723])|(~m[1718]&~m[1719]&~m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&~m[1720]&m[1722]&m[1723])|(m[1718]&~m[1719]&m[1720]&m[1722]&m[1723])|(~m[1718]&m[1719]&m[1720]&m[1722]&m[1723]))&UnbiasedRNG[877])|((m[1718]&m[1719]&~m[1720]&~m[1722]&~m[1723])|(m[1718]&~m[1719]&m[1720]&~m[1722]&~m[1723])|(~m[1718]&m[1719]&m[1720]&~m[1722]&~m[1723])|(m[1718]&m[1719]&m[1720]&~m[1722]&~m[1723])|(m[1718]&~m[1719]&~m[1720]&~m[1722]&m[1723])|(~m[1718]&m[1719]&~m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&~m[1720]&~m[1722]&m[1723])|(~m[1718]&~m[1719]&m[1720]&~m[1722]&m[1723])|(m[1718]&~m[1719]&m[1720]&~m[1722]&m[1723])|(~m[1718]&m[1719]&m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&m[1720]&m[1722]&m[1723]));
    m[1726] = (((m[1723]&~m[1724]&~m[1725]&~m[1727]&~m[1728])|(~m[1723]&m[1724]&~m[1725]&~m[1727]&~m[1728])|(~m[1723]&~m[1724]&m[1725]&~m[1727]&~m[1728])|(m[1723]&m[1724]&m[1725]&m[1727]&~m[1728])|(~m[1723]&~m[1724]&~m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&~m[1725]&m[1727]&m[1728])|(m[1723]&~m[1724]&m[1725]&m[1727]&m[1728])|(~m[1723]&m[1724]&m[1725]&m[1727]&m[1728]))&UnbiasedRNG[878])|((m[1723]&m[1724]&~m[1725]&~m[1727]&~m[1728])|(m[1723]&~m[1724]&m[1725]&~m[1727]&~m[1728])|(~m[1723]&m[1724]&m[1725]&~m[1727]&~m[1728])|(m[1723]&m[1724]&m[1725]&~m[1727]&~m[1728])|(m[1723]&~m[1724]&~m[1725]&~m[1727]&m[1728])|(~m[1723]&m[1724]&~m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&~m[1725]&~m[1727]&m[1728])|(~m[1723]&~m[1724]&m[1725]&~m[1727]&m[1728])|(m[1723]&~m[1724]&m[1725]&~m[1727]&m[1728])|(~m[1723]&m[1724]&m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&m[1725]&m[1727]&m[1728]));
    m[1731] = (((m[1728]&~m[1729]&~m[1730]&~m[1732]&~m[1733])|(~m[1728]&m[1729]&~m[1730]&~m[1732]&~m[1733])|(~m[1728]&~m[1729]&m[1730]&~m[1732]&~m[1733])|(m[1728]&m[1729]&m[1730]&m[1732]&~m[1733])|(~m[1728]&~m[1729]&~m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&~m[1730]&m[1732]&m[1733])|(m[1728]&~m[1729]&m[1730]&m[1732]&m[1733])|(~m[1728]&m[1729]&m[1730]&m[1732]&m[1733]))&UnbiasedRNG[879])|((m[1728]&m[1729]&~m[1730]&~m[1732]&~m[1733])|(m[1728]&~m[1729]&m[1730]&~m[1732]&~m[1733])|(~m[1728]&m[1729]&m[1730]&~m[1732]&~m[1733])|(m[1728]&m[1729]&m[1730]&~m[1732]&~m[1733])|(m[1728]&~m[1729]&~m[1730]&~m[1732]&m[1733])|(~m[1728]&m[1729]&~m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&~m[1730]&~m[1732]&m[1733])|(~m[1728]&~m[1729]&m[1730]&~m[1732]&m[1733])|(m[1728]&~m[1729]&m[1730]&~m[1732]&m[1733])|(~m[1728]&m[1729]&m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&m[1730]&m[1732]&m[1733]));
    m[1741] = (((m[1738]&~m[1739]&~m[1740]&~m[1742]&~m[1743])|(~m[1738]&m[1739]&~m[1740]&~m[1742]&~m[1743])|(~m[1738]&~m[1739]&m[1740]&~m[1742]&~m[1743])|(m[1738]&m[1739]&m[1740]&m[1742]&~m[1743])|(~m[1738]&~m[1739]&~m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&~m[1740]&m[1742]&m[1743])|(m[1738]&~m[1739]&m[1740]&m[1742]&m[1743])|(~m[1738]&m[1739]&m[1740]&m[1742]&m[1743]))&UnbiasedRNG[880])|((m[1738]&m[1739]&~m[1740]&~m[1742]&~m[1743])|(m[1738]&~m[1739]&m[1740]&~m[1742]&~m[1743])|(~m[1738]&m[1739]&m[1740]&~m[1742]&~m[1743])|(m[1738]&m[1739]&m[1740]&~m[1742]&~m[1743])|(m[1738]&~m[1739]&~m[1740]&~m[1742]&m[1743])|(~m[1738]&m[1739]&~m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&~m[1740]&~m[1742]&m[1743])|(~m[1738]&~m[1739]&m[1740]&~m[1742]&m[1743])|(m[1738]&~m[1739]&m[1740]&~m[1742]&m[1743])|(~m[1738]&m[1739]&m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&m[1740]&m[1742]&m[1743]));
    m[1746] = (((m[1743]&~m[1744]&~m[1745]&~m[1747]&~m[1748])|(~m[1743]&m[1744]&~m[1745]&~m[1747]&~m[1748])|(~m[1743]&~m[1744]&m[1745]&~m[1747]&~m[1748])|(m[1743]&m[1744]&m[1745]&m[1747]&~m[1748])|(~m[1743]&~m[1744]&~m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&~m[1745]&m[1747]&m[1748])|(m[1743]&~m[1744]&m[1745]&m[1747]&m[1748])|(~m[1743]&m[1744]&m[1745]&m[1747]&m[1748]))&UnbiasedRNG[881])|((m[1743]&m[1744]&~m[1745]&~m[1747]&~m[1748])|(m[1743]&~m[1744]&m[1745]&~m[1747]&~m[1748])|(~m[1743]&m[1744]&m[1745]&~m[1747]&~m[1748])|(m[1743]&m[1744]&m[1745]&~m[1747]&~m[1748])|(m[1743]&~m[1744]&~m[1745]&~m[1747]&m[1748])|(~m[1743]&m[1744]&~m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&~m[1745]&~m[1747]&m[1748])|(~m[1743]&~m[1744]&m[1745]&~m[1747]&m[1748])|(m[1743]&~m[1744]&m[1745]&~m[1747]&m[1748])|(~m[1743]&m[1744]&m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&m[1745]&m[1747]&m[1748]));
    m[1751] = (((m[1748]&~m[1749]&~m[1750]&~m[1752]&~m[1753])|(~m[1748]&m[1749]&~m[1750]&~m[1752]&~m[1753])|(~m[1748]&~m[1749]&m[1750]&~m[1752]&~m[1753])|(m[1748]&m[1749]&m[1750]&m[1752]&~m[1753])|(~m[1748]&~m[1749]&~m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&~m[1750]&m[1752]&m[1753])|(m[1748]&~m[1749]&m[1750]&m[1752]&m[1753])|(~m[1748]&m[1749]&m[1750]&m[1752]&m[1753]))&UnbiasedRNG[882])|((m[1748]&m[1749]&~m[1750]&~m[1752]&~m[1753])|(m[1748]&~m[1749]&m[1750]&~m[1752]&~m[1753])|(~m[1748]&m[1749]&m[1750]&~m[1752]&~m[1753])|(m[1748]&m[1749]&m[1750]&~m[1752]&~m[1753])|(m[1748]&~m[1749]&~m[1750]&~m[1752]&m[1753])|(~m[1748]&m[1749]&~m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&~m[1750]&~m[1752]&m[1753])|(~m[1748]&~m[1749]&m[1750]&~m[1752]&m[1753])|(m[1748]&~m[1749]&m[1750]&~m[1752]&m[1753])|(~m[1748]&m[1749]&m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&m[1750]&m[1752]&m[1753]));
    m[1756] = (((m[1753]&~m[1754]&~m[1755]&~m[1757]&~m[1758])|(~m[1753]&m[1754]&~m[1755]&~m[1757]&~m[1758])|(~m[1753]&~m[1754]&m[1755]&~m[1757]&~m[1758])|(m[1753]&m[1754]&m[1755]&m[1757]&~m[1758])|(~m[1753]&~m[1754]&~m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&~m[1755]&m[1757]&m[1758])|(m[1753]&~m[1754]&m[1755]&m[1757]&m[1758])|(~m[1753]&m[1754]&m[1755]&m[1757]&m[1758]))&UnbiasedRNG[883])|((m[1753]&m[1754]&~m[1755]&~m[1757]&~m[1758])|(m[1753]&~m[1754]&m[1755]&~m[1757]&~m[1758])|(~m[1753]&m[1754]&m[1755]&~m[1757]&~m[1758])|(m[1753]&m[1754]&m[1755]&~m[1757]&~m[1758])|(m[1753]&~m[1754]&~m[1755]&~m[1757]&m[1758])|(~m[1753]&m[1754]&~m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&~m[1755]&~m[1757]&m[1758])|(~m[1753]&~m[1754]&m[1755]&~m[1757]&m[1758])|(m[1753]&~m[1754]&m[1755]&~m[1757]&m[1758])|(~m[1753]&m[1754]&m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&m[1755]&m[1757]&m[1758]));
    m[1761] = (((m[1758]&~m[1759]&~m[1760]&~m[1762]&~m[1763])|(~m[1758]&m[1759]&~m[1760]&~m[1762]&~m[1763])|(~m[1758]&~m[1759]&m[1760]&~m[1762]&~m[1763])|(m[1758]&m[1759]&m[1760]&m[1762]&~m[1763])|(~m[1758]&~m[1759]&~m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&~m[1760]&m[1762]&m[1763])|(m[1758]&~m[1759]&m[1760]&m[1762]&m[1763])|(~m[1758]&m[1759]&m[1760]&m[1762]&m[1763]))&UnbiasedRNG[884])|((m[1758]&m[1759]&~m[1760]&~m[1762]&~m[1763])|(m[1758]&~m[1759]&m[1760]&~m[1762]&~m[1763])|(~m[1758]&m[1759]&m[1760]&~m[1762]&~m[1763])|(m[1758]&m[1759]&m[1760]&~m[1762]&~m[1763])|(m[1758]&~m[1759]&~m[1760]&~m[1762]&m[1763])|(~m[1758]&m[1759]&~m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&~m[1760]&~m[1762]&m[1763])|(~m[1758]&~m[1759]&m[1760]&~m[1762]&m[1763])|(m[1758]&~m[1759]&m[1760]&~m[1762]&m[1763])|(~m[1758]&m[1759]&m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&m[1760]&m[1762]&m[1763]));
    m[1766] = (((m[1763]&~m[1764]&~m[1765]&~m[1767]&~m[1768])|(~m[1763]&m[1764]&~m[1765]&~m[1767]&~m[1768])|(~m[1763]&~m[1764]&m[1765]&~m[1767]&~m[1768])|(m[1763]&m[1764]&m[1765]&m[1767]&~m[1768])|(~m[1763]&~m[1764]&~m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&~m[1765]&m[1767]&m[1768])|(m[1763]&~m[1764]&m[1765]&m[1767]&m[1768])|(~m[1763]&m[1764]&m[1765]&m[1767]&m[1768]))&UnbiasedRNG[885])|((m[1763]&m[1764]&~m[1765]&~m[1767]&~m[1768])|(m[1763]&~m[1764]&m[1765]&~m[1767]&~m[1768])|(~m[1763]&m[1764]&m[1765]&~m[1767]&~m[1768])|(m[1763]&m[1764]&m[1765]&~m[1767]&~m[1768])|(m[1763]&~m[1764]&~m[1765]&~m[1767]&m[1768])|(~m[1763]&m[1764]&~m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&~m[1765]&~m[1767]&m[1768])|(~m[1763]&~m[1764]&m[1765]&~m[1767]&m[1768])|(m[1763]&~m[1764]&m[1765]&~m[1767]&m[1768])|(~m[1763]&m[1764]&m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&m[1765]&m[1767]&m[1768]));
    m[1771] = (((m[1768]&~m[1769]&~m[1770]&~m[1772]&~m[1773])|(~m[1768]&m[1769]&~m[1770]&~m[1772]&~m[1773])|(~m[1768]&~m[1769]&m[1770]&~m[1772]&~m[1773])|(m[1768]&m[1769]&m[1770]&m[1772]&~m[1773])|(~m[1768]&~m[1769]&~m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&~m[1770]&m[1772]&m[1773])|(m[1768]&~m[1769]&m[1770]&m[1772]&m[1773])|(~m[1768]&m[1769]&m[1770]&m[1772]&m[1773]))&UnbiasedRNG[886])|((m[1768]&m[1769]&~m[1770]&~m[1772]&~m[1773])|(m[1768]&~m[1769]&m[1770]&~m[1772]&~m[1773])|(~m[1768]&m[1769]&m[1770]&~m[1772]&~m[1773])|(m[1768]&m[1769]&m[1770]&~m[1772]&~m[1773])|(m[1768]&~m[1769]&~m[1770]&~m[1772]&m[1773])|(~m[1768]&m[1769]&~m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&~m[1770]&~m[1772]&m[1773])|(~m[1768]&~m[1769]&m[1770]&~m[1772]&m[1773])|(m[1768]&~m[1769]&m[1770]&~m[1772]&m[1773])|(~m[1768]&m[1769]&m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&m[1770]&m[1772]&m[1773]));
    m[1776] = (((m[1773]&~m[1774]&~m[1775]&~m[1777]&~m[1778])|(~m[1773]&m[1774]&~m[1775]&~m[1777]&~m[1778])|(~m[1773]&~m[1774]&m[1775]&~m[1777]&~m[1778])|(m[1773]&m[1774]&m[1775]&m[1777]&~m[1778])|(~m[1773]&~m[1774]&~m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&~m[1775]&m[1777]&m[1778])|(m[1773]&~m[1774]&m[1775]&m[1777]&m[1778])|(~m[1773]&m[1774]&m[1775]&m[1777]&m[1778]))&UnbiasedRNG[887])|((m[1773]&m[1774]&~m[1775]&~m[1777]&~m[1778])|(m[1773]&~m[1774]&m[1775]&~m[1777]&~m[1778])|(~m[1773]&m[1774]&m[1775]&~m[1777]&~m[1778])|(m[1773]&m[1774]&m[1775]&~m[1777]&~m[1778])|(m[1773]&~m[1774]&~m[1775]&~m[1777]&m[1778])|(~m[1773]&m[1774]&~m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&~m[1775]&~m[1777]&m[1778])|(~m[1773]&~m[1774]&m[1775]&~m[1777]&m[1778])|(m[1773]&~m[1774]&m[1775]&~m[1777]&m[1778])|(~m[1773]&m[1774]&m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&m[1775]&m[1777]&m[1778]));
    m[1781] = (((m[1778]&~m[1779]&~m[1780]&~m[1782]&~m[1783])|(~m[1778]&m[1779]&~m[1780]&~m[1782]&~m[1783])|(~m[1778]&~m[1779]&m[1780]&~m[1782]&~m[1783])|(m[1778]&m[1779]&m[1780]&m[1782]&~m[1783])|(~m[1778]&~m[1779]&~m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&~m[1780]&m[1782]&m[1783])|(m[1778]&~m[1779]&m[1780]&m[1782]&m[1783])|(~m[1778]&m[1779]&m[1780]&m[1782]&m[1783]))&UnbiasedRNG[888])|((m[1778]&m[1779]&~m[1780]&~m[1782]&~m[1783])|(m[1778]&~m[1779]&m[1780]&~m[1782]&~m[1783])|(~m[1778]&m[1779]&m[1780]&~m[1782]&~m[1783])|(m[1778]&m[1779]&m[1780]&~m[1782]&~m[1783])|(m[1778]&~m[1779]&~m[1780]&~m[1782]&m[1783])|(~m[1778]&m[1779]&~m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&~m[1780]&~m[1782]&m[1783])|(~m[1778]&~m[1779]&m[1780]&~m[1782]&m[1783])|(m[1778]&~m[1779]&m[1780]&~m[1782]&m[1783])|(~m[1778]&m[1779]&m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&m[1780]&m[1782]&m[1783]));
    m[1786] = (((m[1783]&~m[1784]&~m[1785]&~m[1787]&~m[1788])|(~m[1783]&m[1784]&~m[1785]&~m[1787]&~m[1788])|(~m[1783]&~m[1784]&m[1785]&~m[1787]&~m[1788])|(m[1783]&m[1784]&m[1785]&m[1787]&~m[1788])|(~m[1783]&~m[1784]&~m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&~m[1785]&m[1787]&m[1788])|(m[1783]&~m[1784]&m[1785]&m[1787]&m[1788])|(~m[1783]&m[1784]&m[1785]&m[1787]&m[1788]))&UnbiasedRNG[889])|((m[1783]&m[1784]&~m[1785]&~m[1787]&~m[1788])|(m[1783]&~m[1784]&m[1785]&~m[1787]&~m[1788])|(~m[1783]&m[1784]&m[1785]&~m[1787]&~m[1788])|(m[1783]&m[1784]&m[1785]&~m[1787]&~m[1788])|(m[1783]&~m[1784]&~m[1785]&~m[1787]&m[1788])|(~m[1783]&m[1784]&~m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&~m[1785]&~m[1787]&m[1788])|(~m[1783]&~m[1784]&m[1785]&~m[1787]&m[1788])|(m[1783]&~m[1784]&m[1785]&~m[1787]&m[1788])|(~m[1783]&m[1784]&m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&m[1785]&m[1787]&m[1788]));
    m[1791] = (((m[1788]&~m[1789]&~m[1790]&~m[1792]&~m[1793])|(~m[1788]&m[1789]&~m[1790]&~m[1792]&~m[1793])|(~m[1788]&~m[1789]&m[1790]&~m[1792]&~m[1793])|(m[1788]&m[1789]&m[1790]&m[1792]&~m[1793])|(~m[1788]&~m[1789]&~m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&~m[1790]&m[1792]&m[1793])|(m[1788]&~m[1789]&m[1790]&m[1792]&m[1793])|(~m[1788]&m[1789]&m[1790]&m[1792]&m[1793]))&UnbiasedRNG[890])|((m[1788]&m[1789]&~m[1790]&~m[1792]&~m[1793])|(m[1788]&~m[1789]&m[1790]&~m[1792]&~m[1793])|(~m[1788]&m[1789]&m[1790]&~m[1792]&~m[1793])|(m[1788]&m[1789]&m[1790]&~m[1792]&~m[1793])|(m[1788]&~m[1789]&~m[1790]&~m[1792]&m[1793])|(~m[1788]&m[1789]&~m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&~m[1790]&~m[1792]&m[1793])|(~m[1788]&~m[1789]&m[1790]&~m[1792]&m[1793])|(m[1788]&~m[1789]&m[1790]&~m[1792]&m[1793])|(~m[1788]&m[1789]&m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&m[1790]&m[1792]&m[1793]));
    m[1801] = (((m[1798]&~m[1799]&~m[1800]&~m[1802]&~m[1803])|(~m[1798]&m[1799]&~m[1800]&~m[1802]&~m[1803])|(~m[1798]&~m[1799]&m[1800]&~m[1802]&~m[1803])|(m[1798]&m[1799]&m[1800]&m[1802]&~m[1803])|(~m[1798]&~m[1799]&~m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&~m[1800]&m[1802]&m[1803])|(m[1798]&~m[1799]&m[1800]&m[1802]&m[1803])|(~m[1798]&m[1799]&m[1800]&m[1802]&m[1803]))&UnbiasedRNG[891])|((m[1798]&m[1799]&~m[1800]&~m[1802]&~m[1803])|(m[1798]&~m[1799]&m[1800]&~m[1802]&~m[1803])|(~m[1798]&m[1799]&m[1800]&~m[1802]&~m[1803])|(m[1798]&m[1799]&m[1800]&~m[1802]&~m[1803])|(m[1798]&~m[1799]&~m[1800]&~m[1802]&m[1803])|(~m[1798]&m[1799]&~m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&~m[1800]&~m[1802]&m[1803])|(~m[1798]&~m[1799]&m[1800]&~m[1802]&m[1803])|(m[1798]&~m[1799]&m[1800]&~m[1802]&m[1803])|(~m[1798]&m[1799]&m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&m[1800]&m[1802]&m[1803]));
    m[1806] = (((m[1803]&~m[1804]&~m[1805]&~m[1807]&~m[1808])|(~m[1803]&m[1804]&~m[1805]&~m[1807]&~m[1808])|(~m[1803]&~m[1804]&m[1805]&~m[1807]&~m[1808])|(m[1803]&m[1804]&m[1805]&m[1807]&~m[1808])|(~m[1803]&~m[1804]&~m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&~m[1805]&m[1807]&m[1808])|(m[1803]&~m[1804]&m[1805]&m[1807]&m[1808])|(~m[1803]&m[1804]&m[1805]&m[1807]&m[1808]))&UnbiasedRNG[892])|((m[1803]&m[1804]&~m[1805]&~m[1807]&~m[1808])|(m[1803]&~m[1804]&m[1805]&~m[1807]&~m[1808])|(~m[1803]&m[1804]&m[1805]&~m[1807]&~m[1808])|(m[1803]&m[1804]&m[1805]&~m[1807]&~m[1808])|(m[1803]&~m[1804]&~m[1805]&~m[1807]&m[1808])|(~m[1803]&m[1804]&~m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&~m[1805]&~m[1807]&m[1808])|(~m[1803]&~m[1804]&m[1805]&~m[1807]&m[1808])|(m[1803]&~m[1804]&m[1805]&~m[1807]&m[1808])|(~m[1803]&m[1804]&m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&m[1805]&m[1807]&m[1808]));
    m[1811] = (((m[1808]&~m[1809]&~m[1810]&~m[1812]&~m[1813])|(~m[1808]&m[1809]&~m[1810]&~m[1812]&~m[1813])|(~m[1808]&~m[1809]&m[1810]&~m[1812]&~m[1813])|(m[1808]&m[1809]&m[1810]&m[1812]&~m[1813])|(~m[1808]&~m[1809]&~m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&~m[1810]&m[1812]&m[1813])|(m[1808]&~m[1809]&m[1810]&m[1812]&m[1813])|(~m[1808]&m[1809]&m[1810]&m[1812]&m[1813]))&UnbiasedRNG[893])|((m[1808]&m[1809]&~m[1810]&~m[1812]&~m[1813])|(m[1808]&~m[1809]&m[1810]&~m[1812]&~m[1813])|(~m[1808]&m[1809]&m[1810]&~m[1812]&~m[1813])|(m[1808]&m[1809]&m[1810]&~m[1812]&~m[1813])|(m[1808]&~m[1809]&~m[1810]&~m[1812]&m[1813])|(~m[1808]&m[1809]&~m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&~m[1810]&~m[1812]&m[1813])|(~m[1808]&~m[1809]&m[1810]&~m[1812]&m[1813])|(m[1808]&~m[1809]&m[1810]&~m[1812]&m[1813])|(~m[1808]&m[1809]&m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&m[1810]&m[1812]&m[1813]));
    m[1816] = (((m[1813]&~m[1814]&~m[1815]&~m[1817]&~m[1818])|(~m[1813]&m[1814]&~m[1815]&~m[1817]&~m[1818])|(~m[1813]&~m[1814]&m[1815]&~m[1817]&~m[1818])|(m[1813]&m[1814]&m[1815]&m[1817]&~m[1818])|(~m[1813]&~m[1814]&~m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&~m[1815]&m[1817]&m[1818])|(m[1813]&~m[1814]&m[1815]&m[1817]&m[1818])|(~m[1813]&m[1814]&m[1815]&m[1817]&m[1818]))&UnbiasedRNG[894])|((m[1813]&m[1814]&~m[1815]&~m[1817]&~m[1818])|(m[1813]&~m[1814]&m[1815]&~m[1817]&~m[1818])|(~m[1813]&m[1814]&m[1815]&~m[1817]&~m[1818])|(m[1813]&m[1814]&m[1815]&~m[1817]&~m[1818])|(m[1813]&~m[1814]&~m[1815]&~m[1817]&m[1818])|(~m[1813]&m[1814]&~m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&~m[1815]&~m[1817]&m[1818])|(~m[1813]&~m[1814]&m[1815]&~m[1817]&m[1818])|(m[1813]&~m[1814]&m[1815]&~m[1817]&m[1818])|(~m[1813]&m[1814]&m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&m[1815]&m[1817]&m[1818]));
    m[1821] = (((m[1818]&~m[1819]&~m[1820]&~m[1822]&~m[1823])|(~m[1818]&m[1819]&~m[1820]&~m[1822]&~m[1823])|(~m[1818]&~m[1819]&m[1820]&~m[1822]&~m[1823])|(m[1818]&m[1819]&m[1820]&m[1822]&~m[1823])|(~m[1818]&~m[1819]&~m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&~m[1820]&m[1822]&m[1823])|(m[1818]&~m[1819]&m[1820]&m[1822]&m[1823])|(~m[1818]&m[1819]&m[1820]&m[1822]&m[1823]))&UnbiasedRNG[895])|((m[1818]&m[1819]&~m[1820]&~m[1822]&~m[1823])|(m[1818]&~m[1819]&m[1820]&~m[1822]&~m[1823])|(~m[1818]&m[1819]&m[1820]&~m[1822]&~m[1823])|(m[1818]&m[1819]&m[1820]&~m[1822]&~m[1823])|(m[1818]&~m[1819]&~m[1820]&~m[1822]&m[1823])|(~m[1818]&m[1819]&~m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&~m[1820]&~m[1822]&m[1823])|(~m[1818]&~m[1819]&m[1820]&~m[1822]&m[1823])|(m[1818]&~m[1819]&m[1820]&~m[1822]&m[1823])|(~m[1818]&m[1819]&m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&m[1820]&m[1822]&m[1823]));
    m[1826] = (((m[1823]&~m[1824]&~m[1825]&~m[1827]&~m[1828])|(~m[1823]&m[1824]&~m[1825]&~m[1827]&~m[1828])|(~m[1823]&~m[1824]&m[1825]&~m[1827]&~m[1828])|(m[1823]&m[1824]&m[1825]&m[1827]&~m[1828])|(~m[1823]&~m[1824]&~m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&~m[1825]&m[1827]&m[1828])|(m[1823]&~m[1824]&m[1825]&m[1827]&m[1828])|(~m[1823]&m[1824]&m[1825]&m[1827]&m[1828]))&UnbiasedRNG[896])|((m[1823]&m[1824]&~m[1825]&~m[1827]&~m[1828])|(m[1823]&~m[1824]&m[1825]&~m[1827]&~m[1828])|(~m[1823]&m[1824]&m[1825]&~m[1827]&~m[1828])|(m[1823]&m[1824]&m[1825]&~m[1827]&~m[1828])|(m[1823]&~m[1824]&~m[1825]&~m[1827]&m[1828])|(~m[1823]&m[1824]&~m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&~m[1825]&~m[1827]&m[1828])|(~m[1823]&~m[1824]&m[1825]&~m[1827]&m[1828])|(m[1823]&~m[1824]&m[1825]&~m[1827]&m[1828])|(~m[1823]&m[1824]&m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&m[1825]&m[1827]&m[1828]));
    m[1831] = (((m[1828]&~m[1829]&~m[1830]&~m[1832]&~m[1833])|(~m[1828]&m[1829]&~m[1830]&~m[1832]&~m[1833])|(~m[1828]&~m[1829]&m[1830]&~m[1832]&~m[1833])|(m[1828]&m[1829]&m[1830]&m[1832]&~m[1833])|(~m[1828]&~m[1829]&~m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&~m[1830]&m[1832]&m[1833])|(m[1828]&~m[1829]&m[1830]&m[1832]&m[1833])|(~m[1828]&m[1829]&m[1830]&m[1832]&m[1833]))&UnbiasedRNG[897])|((m[1828]&m[1829]&~m[1830]&~m[1832]&~m[1833])|(m[1828]&~m[1829]&m[1830]&~m[1832]&~m[1833])|(~m[1828]&m[1829]&m[1830]&~m[1832]&~m[1833])|(m[1828]&m[1829]&m[1830]&~m[1832]&~m[1833])|(m[1828]&~m[1829]&~m[1830]&~m[1832]&m[1833])|(~m[1828]&m[1829]&~m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&~m[1830]&~m[1832]&m[1833])|(~m[1828]&~m[1829]&m[1830]&~m[1832]&m[1833])|(m[1828]&~m[1829]&m[1830]&~m[1832]&m[1833])|(~m[1828]&m[1829]&m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&m[1830]&m[1832]&m[1833]));
    m[1836] = (((m[1833]&~m[1834]&~m[1835]&~m[1837]&~m[1838])|(~m[1833]&m[1834]&~m[1835]&~m[1837]&~m[1838])|(~m[1833]&~m[1834]&m[1835]&~m[1837]&~m[1838])|(m[1833]&m[1834]&m[1835]&m[1837]&~m[1838])|(~m[1833]&~m[1834]&~m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&~m[1835]&m[1837]&m[1838])|(m[1833]&~m[1834]&m[1835]&m[1837]&m[1838])|(~m[1833]&m[1834]&m[1835]&m[1837]&m[1838]))&UnbiasedRNG[898])|((m[1833]&m[1834]&~m[1835]&~m[1837]&~m[1838])|(m[1833]&~m[1834]&m[1835]&~m[1837]&~m[1838])|(~m[1833]&m[1834]&m[1835]&~m[1837]&~m[1838])|(m[1833]&m[1834]&m[1835]&~m[1837]&~m[1838])|(m[1833]&~m[1834]&~m[1835]&~m[1837]&m[1838])|(~m[1833]&m[1834]&~m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&~m[1835]&~m[1837]&m[1838])|(~m[1833]&~m[1834]&m[1835]&~m[1837]&m[1838])|(m[1833]&~m[1834]&m[1835]&~m[1837]&m[1838])|(~m[1833]&m[1834]&m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&m[1835]&m[1837]&m[1838]));
    m[1841] = (((m[1838]&~m[1839]&~m[1840]&~m[1842]&~m[1843])|(~m[1838]&m[1839]&~m[1840]&~m[1842]&~m[1843])|(~m[1838]&~m[1839]&m[1840]&~m[1842]&~m[1843])|(m[1838]&m[1839]&m[1840]&m[1842]&~m[1843])|(~m[1838]&~m[1839]&~m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&~m[1840]&m[1842]&m[1843])|(m[1838]&~m[1839]&m[1840]&m[1842]&m[1843])|(~m[1838]&m[1839]&m[1840]&m[1842]&m[1843]))&UnbiasedRNG[899])|((m[1838]&m[1839]&~m[1840]&~m[1842]&~m[1843])|(m[1838]&~m[1839]&m[1840]&~m[1842]&~m[1843])|(~m[1838]&m[1839]&m[1840]&~m[1842]&~m[1843])|(m[1838]&m[1839]&m[1840]&~m[1842]&~m[1843])|(m[1838]&~m[1839]&~m[1840]&~m[1842]&m[1843])|(~m[1838]&m[1839]&~m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&~m[1840]&~m[1842]&m[1843])|(~m[1838]&~m[1839]&m[1840]&~m[1842]&m[1843])|(m[1838]&~m[1839]&m[1840]&~m[1842]&m[1843])|(~m[1838]&m[1839]&m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&m[1840]&m[1842]&m[1843]));
    m[1846] = (((m[1843]&~m[1844]&~m[1845]&~m[1847]&~m[1848])|(~m[1843]&m[1844]&~m[1845]&~m[1847]&~m[1848])|(~m[1843]&~m[1844]&m[1845]&~m[1847]&~m[1848])|(m[1843]&m[1844]&m[1845]&m[1847]&~m[1848])|(~m[1843]&~m[1844]&~m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&~m[1845]&m[1847]&m[1848])|(m[1843]&~m[1844]&m[1845]&m[1847]&m[1848])|(~m[1843]&m[1844]&m[1845]&m[1847]&m[1848]))&UnbiasedRNG[900])|((m[1843]&m[1844]&~m[1845]&~m[1847]&~m[1848])|(m[1843]&~m[1844]&m[1845]&~m[1847]&~m[1848])|(~m[1843]&m[1844]&m[1845]&~m[1847]&~m[1848])|(m[1843]&m[1844]&m[1845]&~m[1847]&~m[1848])|(m[1843]&~m[1844]&~m[1845]&~m[1847]&m[1848])|(~m[1843]&m[1844]&~m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&~m[1845]&~m[1847]&m[1848])|(~m[1843]&~m[1844]&m[1845]&~m[1847]&m[1848])|(m[1843]&~m[1844]&m[1845]&~m[1847]&m[1848])|(~m[1843]&m[1844]&m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&m[1845]&m[1847]&m[1848]));
    m[1856] = (((m[1853]&~m[1854]&~m[1855]&~m[1857]&~m[1858])|(~m[1853]&m[1854]&~m[1855]&~m[1857]&~m[1858])|(~m[1853]&~m[1854]&m[1855]&~m[1857]&~m[1858])|(m[1853]&m[1854]&m[1855]&m[1857]&~m[1858])|(~m[1853]&~m[1854]&~m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&~m[1855]&m[1857]&m[1858])|(m[1853]&~m[1854]&m[1855]&m[1857]&m[1858])|(~m[1853]&m[1854]&m[1855]&m[1857]&m[1858]))&UnbiasedRNG[901])|((m[1853]&m[1854]&~m[1855]&~m[1857]&~m[1858])|(m[1853]&~m[1854]&m[1855]&~m[1857]&~m[1858])|(~m[1853]&m[1854]&m[1855]&~m[1857]&~m[1858])|(m[1853]&m[1854]&m[1855]&~m[1857]&~m[1858])|(m[1853]&~m[1854]&~m[1855]&~m[1857]&m[1858])|(~m[1853]&m[1854]&~m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&~m[1855]&~m[1857]&m[1858])|(~m[1853]&~m[1854]&m[1855]&~m[1857]&m[1858])|(m[1853]&~m[1854]&m[1855]&~m[1857]&m[1858])|(~m[1853]&m[1854]&m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&m[1855]&m[1857]&m[1858]));
    m[1861] = (((m[1858]&~m[1859]&~m[1860]&~m[1862]&~m[1863])|(~m[1858]&m[1859]&~m[1860]&~m[1862]&~m[1863])|(~m[1858]&~m[1859]&m[1860]&~m[1862]&~m[1863])|(m[1858]&m[1859]&m[1860]&m[1862]&~m[1863])|(~m[1858]&~m[1859]&~m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&~m[1860]&m[1862]&m[1863])|(m[1858]&~m[1859]&m[1860]&m[1862]&m[1863])|(~m[1858]&m[1859]&m[1860]&m[1862]&m[1863]))&UnbiasedRNG[902])|((m[1858]&m[1859]&~m[1860]&~m[1862]&~m[1863])|(m[1858]&~m[1859]&m[1860]&~m[1862]&~m[1863])|(~m[1858]&m[1859]&m[1860]&~m[1862]&~m[1863])|(m[1858]&m[1859]&m[1860]&~m[1862]&~m[1863])|(m[1858]&~m[1859]&~m[1860]&~m[1862]&m[1863])|(~m[1858]&m[1859]&~m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&~m[1860]&~m[1862]&m[1863])|(~m[1858]&~m[1859]&m[1860]&~m[1862]&m[1863])|(m[1858]&~m[1859]&m[1860]&~m[1862]&m[1863])|(~m[1858]&m[1859]&m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&m[1860]&m[1862]&m[1863]));
    m[1866] = (((m[1863]&~m[1864]&~m[1865]&~m[1867]&~m[1868])|(~m[1863]&m[1864]&~m[1865]&~m[1867]&~m[1868])|(~m[1863]&~m[1864]&m[1865]&~m[1867]&~m[1868])|(m[1863]&m[1864]&m[1865]&m[1867]&~m[1868])|(~m[1863]&~m[1864]&~m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&~m[1865]&m[1867]&m[1868])|(m[1863]&~m[1864]&m[1865]&m[1867]&m[1868])|(~m[1863]&m[1864]&m[1865]&m[1867]&m[1868]))&UnbiasedRNG[903])|((m[1863]&m[1864]&~m[1865]&~m[1867]&~m[1868])|(m[1863]&~m[1864]&m[1865]&~m[1867]&~m[1868])|(~m[1863]&m[1864]&m[1865]&~m[1867]&~m[1868])|(m[1863]&m[1864]&m[1865]&~m[1867]&~m[1868])|(m[1863]&~m[1864]&~m[1865]&~m[1867]&m[1868])|(~m[1863]&m[1864]&~m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&~m[1865]&~m[1867]&m[1868])|(~m[1863]&~m[1864]&m[1865]&~m[1867]&m[1868])|(m[1863]&~m[1864]&m[1865]&~m[1867]&m[1868])|(~m[1863]&m[1864]&m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&m[1865]&m[1867]&m[1868]));
    m[1871] = (((m[1868]&~m[1869]&~m[1870]&~m[1872]&~m[1873])|(~m[1868]&m[1869]&~m[1870]&~m[1872]&~m[1873])|(~m[1868]&~m[1869]&m[1870]&~m[1872]&~m[1873])|(m[1868]&m[1869]&m[1870]&m[1872]&~m[1873])|(~m[1868]&~m[1869]&~m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&~m[1870]&m[1872]&m[1873])|(m[1868]&~m[1869]&m[1870]&m[1872]&m[1873])|(~m[1868]&m[1869]&m[1870]&m[1872]&m[1873]))&UnbiasedRNG[904])|((m[1868]&m[1869]&~m[1870]&~m[1872]&~m[1873])|(m[1868]&~m[1869]&m[1870]&~m[1872]&~m[1873])|(~m[1868]&m[1869]&m[1870]&~m[1872]&~m[1873])|(m[1868]&m[1869]&m[1870]&~m[1872]&~m[1873])|(m[1868]&~m[1869]&~m[1870]&~m[1872]&m[1873])|(~m[1868]&m[1869]&~m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&~m[1870]&~m[1872]&m[1873])|(~m[1868]&~m[1869]&m[1870]&~m[1872]&m[1873])|(m[1868]&~m[1869]&m[1870]&~m[1872]&m[1873])|(~m[1868]&m[1869]&m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&m[1870]&m[1872]&m[1873]));
    m[1876] = (((m[1873]&~m[1874]&~m[1875]&~m[1877]&~m[1878])|(~m[1873]&m[1874]&~m[1875]&~m[1877]&~m[1878])|(~m[1873]&~m[1874]&m[1875]&~m[1877]&~m[1878])|(m[1873]&m[1874]&m[1875]&m[1877]&~m[1878])|(~m[1873]&~m[1874]&~m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&~m[1875]&m[1877]&m[1878])|(m[1873]&~m[1874]&m[1875]&m[1877]&m[1878])|(~m[1873]&m[1874]&m[1875]&m[1877]&m[1878]))&UnbiasedRNG[905])|((m[1873]&m[1874]&~m[1875]&~m[1877]&~m[1878])|(m[1873]&~m[1874]&m[1875]&~m[1877]&~m[1878])|(~m[1873]&m[1874]&m[1875]&~m[1877]&~m[1878])|(m[1873]&m[1874]&m[1875]&~m[1877]&~m[1878])|(m[1873]&~m[1874]&~m[1875]&~m[1877]&m[1878])|(~m[1873]&m[1874]&~m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&~m[1875]&~m[1877]&m[1878])|(~m[1873]&~m[1874]&m[1875]&~m[1877]&m[1878])|(m[1873]&~m[1874]&m[1875]&~m[1877]&m[1878])|(~m[1873]&m[1874]&m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&m[1875]&m[1877]&m[1878]));
    m[1881] = (((m[1878]&~m[1879]&~m[1880]&~m[1882]&~m[1883])|(~m[1878]&m[1879]&~m[1880]&~m[1882]&~m[1883])|(~m[1878]&~m[1879]&m[1880]&~m[1882]&~m[1883])|(m[1878]&m[1879]&m[1880]&m[1882]&~m[1883])|(~m[1878]&~m[1879]&~m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&~m[1880]&m[1882]&m[1883])|(m[1878]&~m[1879]&m[1880]&m[1882]&m[1883])|(~m[1878]&m[1879]&m[1880]&m[1882]&m[1883]))&UnbiasedRNG[906])|((m[1878]&m[1879]&~m[1880]&~m[1882]&~m[1883])|(m[1878]&~m[1879]&m[1880]&~m[1882]&~m[1883])|(~m[1878]&m[1879]&m[1880]&~m[1882]&~m[1883])|(m[1878]&m[1879]&m[1880]&~m[1882]&~m[1883])|(m[1878]&~m[1879]&~m[1880]&~m[1882]&m[1883])|(~m[1878]&m[1879]&~m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&~m[1880]&~m[1882]&m[1883])|(~m[1878]&~m[1879]&m[1880]&~m[1882]&m[1883])|(m[1878]&~m[1879]&m[1880]&~m[1882]&m[1883])|(~m[1878]&m[1879]&m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&m[1880]&m[1882]&m[1883]));
    m[1886] = (((m[1883]&~m[1884]&~m[1885]&~m[1887]&~m[1888])|(~m[1883]&m[1884]&~m[1885]&~m[1887]&~m[1888])|(~m[1883]&~m[1884]&m[1885]&~m[1887]&~m[1888])|(m[1883]&m[1884]&m[1885]&m[1887]&~m[1888])|(~m[1883]&~m[1884]&~m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&~m[1885]&m[1887]&m[1888])|(m[1883]&~m[1884]&m[1885]&m[1887]&m[1888])|(~m[1883]&m[1884]&m[1885]&m[1887]&m[1888]))&UnbiasedRNG[907])|((m[1883]&m[1884]&~m[1885]&~m[1887]&~m[1888])|(m[1883]&~m[1884]&m[1885]&~m[1887]&~m[1888])|(~m[1883]&m[1884]&m[1885]&~m[1887]&~m[1888])|(m[1883]&m[1884]&m[1885]&~m[1887]&~m[1888])|(m[1883]&~m[1884]&~m[1885]&~m[1887]&m[1888])|(~m[1883]&m[1884]&~m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&~m[1885]&~m[1887]&m[1888])|(~m[1883]&~m[1884]&m[1885]&~m[1887]&m[1888])|(m[1883]&~m[1884]&m[1885]&~m[1887]&m[1888])|(~m[1883]&m[1884]&m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&m[1885]&m[1887]&m[1888]));
    m[1891] = (((m[1888]&~m[1889]&~m[1890]&~m[1892]&~m[1893])|(~m[1888]&m[1889]&~m[1890]&~m[1892]&~m[1893])|(~m[1888]&~m[1889]&m[1890]&~m[1892]&~m[1893])|(m[1888]&m[1889]&m[1890]&m[1892]&~m[1893])|(~m[1888]&~m[1889]&~m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&~m[1890]&m[1892]&m[1893])|(m[1888]&~m[1889]&m[1890]&m[1892]&m[1893])|(~m[1888]&m[1889]&m[1890]&m[1892]&m[1893]))&UnbiasedRNG[908])|((m[1888]&m[1889]&~m[1890]&~m[1892]&~m[1893])|(m[1888]&~m[1889]&m[1890]&~m[1892]&~m[1893])|(~m[1888]&m[1889]&m[1890]&~m[1892]&~m[1893])|(m[1888]&m[1889]&m[1890]&~m[1892]&~m[1893])|(m[1888]&~m[1889]&~m[1890]&~m[1892]&m[1893])|(~m[1888]&m[1889]&~m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&~m[1890]&~m[1892]&m[1893])|(~m[1888]&~m[1889]&m[1890]&~m[1892]&m[1893])|(m[1888]&~m[1889]&m[1890]&~m[1892]&m[1893])|(~m[1888]&m[1889]&m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&m[1890]&m[1892]&m[1893]));
    m[1896] = (((m[1893]&~m[1894]&~m[1895]&~m[1897]&~m[1898])|(~m[1893]&m[1894]&~m[1895]&~m[1897]&~m[1898])|(~m[1893]&~m[1894]&m[1895]&~m[1897]&~m[1898])|(m[1893]&m[1894]&m[1895]&m[1897]&~m[1898])|(~m[1893]&~m[1894]&~m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&~m[1895]&m[1897]&m[1898])|(m[1893]&~m[1894]&m[1895]&m[1897]&m[1898])|(~m[1893]&m[1894]&m[1895]&m[1897]&m[1898]))&UnbiasedRNG[909])|((m[1893]&m[1894]&~m[1895]&~m[1897]&~m[1898])|(m[1893]&~m[1894]&m[1895]&~m[1897]&~m[1898])|(~m[1893]&m[1894]&m[1895]&~m[1897]&~m[1898])|(m[1893]&m[1894]&m[1895]&~m[1897]&~m[1898])|(m[1893]&~m[1894]&~m[1895]&~m[1897]&m[1898])|(~m[1893]&m[1894]&~m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&~m[1895]&~m[1897]&m[1898])|(~m[1893]&~m[1894]&m[1895]&~m[1897]&m[1898])|(m[1893]&~m[1894]&m[1895]&~m[1897]&m[1898])|(~m[1893]&m[1894]&m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&m[1895]&m[1897]&m[1898]));
    m[1906] = (((m[1903]&~m[1904]&~m[1905]&~m[1907]&~m[1908])|(~m[1903]&m[1904]&~m[1905]&~m[1907]&~m[1908])|(~m[1903]&~m[1904]&m[1905]&~m[1907]&~m[1908])|(m[1903]&m[1904]&m[1905]&m[1907]&~m[1908])|(~m[1903]&~m[1904]&~m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&~m[1905]&m[1907]&m[1908])|(m[1903]&~m[1904]&m[1905]&m[1907]&m[1908])|(~m[1903]&m[1904]&m[1905]&m[1907]&m[1908]))&UnbiasedRNG[910])|((m[1903]&m[1904]&~m[1905]&~m[1907]&~m[1908])|(m[1903]&~m[1904]&m[1905]&~m[1907]&~m[1908])|(~m[1903]&m[1904]&m[1905]&~m[1907]&~m[1908])|(m[1903]&m[1904]&m[1905]&~m[1907]&~m[1908])|(m[1903]&~m[1904]&~m[1905]&~m[1907]&m[1908])|(~m[1903]&m[1904]&~m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&~m[1905]&~m[1907]&m[1908])|(~m[1903]&~m[1904]&m[1905]&~m[1907]&m[1908])|(m[1903]&~m[1904]&m[1905]&~m[1907]&m[1908])|(~m[1903]&m[1904]&m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&m[1905]&m[1907]&m[1908]));
    m[1911] = (((m[1908]&~m[1909]&~m[1910]&~m[1912]&~m[1913])|(~m[1908]&m[1909]&~m[1910]&~m[1912]&~m[1913])|(~m[1908]&~m[1909]&m[1910]&~m[1912]&~m[1913])|(m[1908]&m[1909]&m[1910]&m[1912]&~m[1913])|(~m[1908]&~m[1909]&~m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&~m[1910]&m[1912]&m[1913])|(m[1908]&~m[1909]&m[1910]&m[1912]&m[1913])|(~m[1908]&m[1909]&m[1910]&m[1912]&m[1913]))&UnbiasedRNG[911])|((m[1908]&m[1909]&~m[1910]&~m[1912]&~m[1913])|(m[1908]&~m[1909]&m[1910]&~m[1912]&~m[1913])|(~m[1908]&m[1909]&m[1910]&~m[1912]&~m[1913])|(m[1908]&m[1909]&m[1910]&~m[1912]&~m[1913])|(m[1908]&~m[1909]&~m[1910]&~m[1912]&m[1913])|(~m[1908]&m[1909]&~m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&~m[1910]&~m[1912]&m[1913])|(~m[1908]&~m[1909]&m[1910]&~m[1912]&m[1913])|(m[1908]&~m[1909]&m[1910]&~m[1912]&m[1913])|(~m[1908]&m[1909]&m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&m[1910]&m[1912]&m[1913]));
    m[1916] = (((m[1913]&~m[1914]&~m[1915]&~m[1917]&~m[1918])|(~m[1913]&m[1914]&~m[1915]&~m[1917]&~m[1918])|(~m[1913]&~m[1914]&m[1915]&~m[1917]&~m[1918])|(m[1913]&m[1914]&m[1915]&m[1917]&~m[1918])|(~m[1913]&~m[1914]&~m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&~m[1915]&m[1917]&m[1918])|(m[1913]&~m[1914]&m[1915]&m[1917]&m[1918])|(~m[1913]&m[1914]&m[1915]&m[1917]&m[1918]))&UnbiasedRNG[912])|((m[1913]&m[1914]&~m[1915]&~m[1917]&~m[1918])|(m[1913]&~m[1914]&m[1915]&~m[1917]&~m[1918])|(~m[1913]&m[1914]&m[1915]&~m[1917]&~m[1918])|(m[1913]&m[1914]&m[1915]&~m[1917]&~m[1918])|(m[1913]&~m[1914]&~m[1915]&~m[1917]&m[1918])|(~m[1913]&m[1914]&~m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&~m[1915]&~m[1917]&m[1918])|(~m[1913]&~m[1914]&m[1915]&~m[1917]&m[1918])|(m[1913]&~m[1914]&m[1915]&~m[1917]&m[1918])|(~m[1913]&m[1914]&m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&m[1915]&m[1917]&m[1918]));
    m[1921] = (((m[1918]&~m[1919]&~m[1920]&~m[1922]&~m[1923])|(~m[1918]&m[1919]&~m[1920]&~m[1922]&~m[1923])|(~m[1918]&~m[1919]&m[1920]&~m[1922]&~m[1923])|(m[1918]&m[1919]&m[1920]&m[1922]&~m[1923])|(~m[1918]&~m[1919]&~m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&~m[1920]&m[1922]&m[1923])|(m[1918]&~m[1919]&m[1920]&m[1922]&m[1923])|(~m[1918]&m[1919]&m[1920]&m[1922]&m[1923]))&UnbiasedRNG[913])|((m[1918]&m[1919]&~m[1920]&~m[1922]&~m[1923])|(m[1918]&~m[1919]&m[1920]&~m[1922]&~m[1923])|(~m[1918]&m[1919]&m[1920]&~m[1922]&~m[1923])|(m[1918]&m[1919]&m[1920]&~m[1922]&~m[1923])|(m[1918]&~m[1919]&~m[1920]&~m[1922]&m[1923])|(~m[1918]&m[1919]&~m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&~m[1920]&~m[1922]&m[1923])|(~m[1918]&~m[1919]&m[1920]&~m[1922]&m[1923])|(m[1918]&~m[1919]&m[1920]&~m[1922]&m[1923])|(~m[1918]&m[1919]&m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&m[1920]&m[1922]&m[1923]));
    m[1926] = (((m[1923]&~m[1924]&~m[1925]&~m[1927]&~m[1928])|(~m[1923]&m[1924]&~m[1925]&~m[1927]&~m[1928])|(~m[1923]&~m[1924]&m[1925]&~m[1927]&~m[1928])|(m[1923]&m[1924]&m[1925]&m[1927]&~m[1928])|(~m[1923]&~m[1924]&~m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&~m[1925]&m[1927]&m[1928])|(m[1923]&~m[1924]&m[1925]&m[1927]&m[1928])|(~m[1923]&m[1924]&m[1925]&m[1927]&m[1928]))&UnbiasedRNG[914])|((m[1923]&m[1924]&~m[1925]&~m[1927]&~m[1928])|(m[1923]&~m[1924]&m[1925]&~m[1927]&~m[1928])|(~m[1923]&m[1924]&m[1925]&~m[1927]&~m[1928])|(m[1923]&m[1924]&m[1925]&~m[1927]&~m[1928])|(m[1923]&~m[1924]&~m[1925]&~m[1927]&m[1928])|(~m[1923]&m[1924]&~m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&~m[1925]&~m[1927]&m[1928])|(~m[1923]&~m[1924]&m[1925]&~m[1927]&m[1928])|(m[1923]&~m[1924]&m[1925]&~m[1927]&m[1928])|(~m[1923]&m[1924]&m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&m[1925]&m[1927]&m[1928]));
    m[1931] = (((m[1928]&~m[1929]&~m[1930]&~m[1932]&~m[1933])|(~m[1928]&m[1929]&~m[1930]&~m[1932]&~m[1933])|(~m[1928]&~m[1929]&m[1930]&~m[1932]&~m[1933])|(m[1928]&m[1929]&m[1930]&m[1932]&~m[1933])|(~m[1928]&~m[1929]&~m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&~m[1930]&m[1932]&m[1933])|(m[1928]&~m[1929]&m[1930]&m[1932]&m[1933])|(~m[1928]&m[1929]&m[1930]&m[1932]&m[1933]))&UnbiasedRNG[915])|((m[1928]&m[1929]&~m[1930]&~m[1932]&~m[1933])|(m[1928]&~m[1929]&m[1930]&~m[1932]&~m[1933])|(~m[1928]&m[1929]&m[1930]&~m[1932]&~m[1933])|(m[1928]&m[1929]&m[1930]&~m[1932]&~m[1933])|(m[1928]&~m[1929]&~m[1930]&~m[1932]&m[1933])|(~m[1928]&m[1929]&~m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&~m[1930]&~m[1932]&m[1933])|(~m[1928]&~m[1929]&m[1930]&~m[1932]&m[1933])|(m[1928]&~m[1929]&m[1930]&~m[1932]&m[1933])|(~m[1928]&m[1929]&m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&m[1930]&m[1932]&m[1933]));
    m[1936] = (((m[1933]&~m[1934]&~m[1935]&~m[1937]&~m[1938])|(~m[1933]&m[1934]&~m[1935]&~m[1937]&~m[1938])|(~m[1933]&~m[1934]&m[1935]&~m[1937]&~m[1938])|(m[1933]&m[1934]&m[1935]&m[1937]&~m[1938])|(~m[1933]&~m[1934]&~m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&~m[1935]&m[1937]&m[1938])|(m[1933]&~m[1934]&m[1935]&m[1937]&m[1938])|(~m[1933]&m[1934]&m[1935]&m[1937]&m[1938]))&UnbiasedRNG[916])|((m[1933]&m[1934]&~m[1935]&~m[1937]&~m[1938])|(m[1933]&~m[1934]&m[1935]&~m[1937]&~m[1938])|(~m[1933]&m[1934]&m[1935]&~m[1937]&~m[1938])|(m[1933]&m[1934]&m[1935]&~m[1937]&~m[1938])|(m[1933]&~m[1934]&~m[1935]&~m[1937]&m[1938])|(~m[1933]&m[1934]&~m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&~m[1935]&~m[1937]&m[1938])|(~m[1933]&~m[1934]&m[1935]&~m[1937]&m[1938])|(m[1933]&~m[1934]&m[1935]&~m[1937]&m[1938])|(~m[1933]&m[1934]&m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&m[1935]&m[1937]&m[1938]));
    m[1941] = (((m[1938]&~m[1939]&~m[1940]&~m[1942]&~m[1943])|(~m[1938]&m[1939]&~m[1940]&~m[1942]&~m[1943])|(~m[1938]&~m[1939]&m[1940]&~m[1942]&~m[1943])|(m[1938]&m[1939]&m[1940]&m[1942]&~m[1943])|(~m[1938]&~m[1939]&~m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&~m[1940]&m[1942]&m[1943])|(m[1938]&~m[1939]&m[1940]&m[1942]&m[1943])|(~m[1938]&m[1939]&m[1940]&m[1942]&m[1943]))&UnbiasedRNG[917])|((m[1938]&m[1939]&~m[1940]&~m[1942]&~m[1943])|(m[1938]&~m[1939]&m[1940]&~m[1942]&~m[1943])|(~m[1938]&m[1939]&m[1940]&~m[1942]&~m[1943])|(m[1938]&m[1939]&m[1940]&~m[1942]&~m[1943])|(m[1938]&~m[1939]&~m[1940]&~m[1942]&m[1943])|(~m[1938]&m[1939]&~m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&~m[1940]&~m[1942]&m[1943])|(~m[1938]&~m[1939]&m[1940]&~m[1942]&m[1943])|(m[1938]&~m[1939]&m[1940]&~m[1942]&m[1943])|(~m[1938]&m[1939]&m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&m[1940]&m[1942]&m[1943]));
    m[1951] = (((m[1948]&~m[1949]&~m[1950]&~m[1952]&~m[1953])|(~m[1948]&m[1949]&~m[1950]&~m[1952]&~m[1953])|(~m[1948]&~m[1949]&m[1950]&~m[1952]&~m[1953])|(m[1948]&m[1949]&m[1950]&m[1952]&~m[1953])|(~m[1948]&~m[1949]&~m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&~m[1950]&m[1952]&m[1953])|(m[1948]&~m[1949]&m[1950]&m[1952]&m[1953])|(~m[1948]&m[1949]&m[1950]&m[1952]&m[1953]))&UnbiasedRNG[918])|((m[1948]&m[1949]&~m[1950]&~m[1952]&~m[1953])|(m[1948]&~m[1949]&m[1950]&~m[1952]&~m[1953])|(~m[1948]&m[1949]&m[1950]&~m[1952]&~m[1953])|(m[1948]&m[1949]&m[1950]&~m[1952]&~m[1953])|(m[1948]&~m[1949]&~m[1950]&~m[1952]&m[1953])|(~m[1948]&m[1949]&~m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&~m[1950]&~m[1952]&m[1953])|(~m[1948]&~m[1949]&m[1950]&~m[1952]&m[1953])|(m[1948]&~m[1949]&m[1950]&~m[1952]&m[1953])|(~m[1948]&m[1949]&m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&m[1950]&m[1952]&m[1953]));
    m[1956] = (((m[1953]&~m[1954]&~m[1955]&~m[1957]&~m[1958])|(~m[1953]&m[1954]&~m[1955]&~m[1957]&~m[1958])|(~m[1953]&~m[1954]&m[1955]&~m[1957]&~m[1958])|(m[1953]&m[1954]&m[1955]&m[1957]&~m[1958])|(~m[1953]&~m[1954]&~m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&~m[1955]&m[1957]&m[1958])|(m[1953]&~m[1954]&m[1955]&m[1957]&m[1958])|(~m[1953]&m[1954]&m[1955]&m[1957]&m[1958]))&UnbiasedRNG[919])|((m[1953]&m[1954]&~m[1955]&~m[1957]&~m[1958])|(m[1953]&~m[1954]&m[1955]&~m[1957]&~m[1958])|(~m[1953]&m[1954]&m[1955]&~m[1957]&~m[1958])|(m[1953]&m[1954]&m[1955]&~m[1957]&~m[1958])|(m[1953]&~m[1954]&~m[1955]&~m[1957]&m[1958])|(~m[1953]&m[1954]&~m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&~m[1955]&~m[1957]&m[1958])|(~m[1953]&~m[1954]&m[1955]&~m[1957]&m[1958])|(m[1953]&~m[1954]&m[1955]&~m[1957]&m[1958])|(~m[1953]&m[1954]&m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&m[1955]&m[1957]&m[1958]));
    m[1961] = (((m[1958]&~m[1959]&~m[1960]&~m[1962]&~m[1963])|(~m[1958]&m[1959]&~m[1960]&~m[1962]&~m[1963])|(~m[1958]&~m[1959]&m[1960]&~m[1962]&~m[1963])|(m[1958]&m[1959]&m[1960]&m[1962]&~m[1963])|(~m[1958]&~m[1959]&~m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&~m[1960]&m[1962]&m[1963])|(m[1958]&~m[1959]&m[1960]&m[1962]&m[1963])|(~m[1958]&m[1959]&m[1960]&m[1962]&m[1963]))&UnbiasedRNG[920])|((m[1958]&m[1959]&~m[1960]&~m[1962]&~m[1963])|(m[1958]&~m[1959]&m[1960]&~m[1962]&~m[1963])|(~m[1958]&m[1959]&m[1960]&~m[1962]&~m[1963])|(m[1958]&m[1959]&m[1960]&~m[1962]&~m[1963])|(m[1958]&~m[1959]&~m[1960]&~m[1962]&m[1963])|(~m[1958]&m[1959]&~m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&~m[1960]&~m[1962]&m[1963])|(~m[1958]&~m[1959]&m[1960]&~m[1962]&m[1963])|(m[1958]&~m[1959]&m[1960]&~m[1962]&m[1963])|(~m[1958]&m[1959]&m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&m[1960]&m[1962]&m[1963]));
    m[1966] = (((m[1963]&~m[1964]&~m[1965]&~m[1967]&~m[1968])|(~m[1963]&m[1964]&~m[1965]&~m[1967]&~m[1968])|(~m[1963]&~m[1964]&m[1965]&~m[1967]&~m[1968])|(m[1963]&m[1964]&m[1965]&m[1967]&~m[1968])|(~m[1963]&~m[1964]&~m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&~m[1965]&m[1967]&m[1968])|(m[1963]&~m[1964]&m[1965]&m[1967]&m[1968])|(~m[1963]&m[1964]&m[1965]&m[1967]&m[1968]))&UnbiasedRNG[921])|((m[1963]&m[1964]&~m[1965]&~m[1967]&~m[1968])|(m[1963]&~m[1964]&m[1965]&~m[1967]&~m[1968])|(~m[1963]&m[1964]&m[1965]&~m[1967]&~m[1968])|(m[1963]&m[1964]&m[1965]&~m[1967]&~m[1968])|(m[1963]&~m[1964]&~m[1965]&~m[1967]&m[1968])|(~m[1963]&m[1964]&~m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&~m[1965]&~m[1967]&m[1968])|(~m[1963]&~m[1964]&m[1965]&~m[1967]&m[1968])|(m[1963]&~m[1964]&m[1965]&~m[1967]&m[1968])|(~m[1963]&m[1964]&m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&m[1965]&m[1967]&m[1968]));
    m[1971] = (((m[1968]&~m[1969]&~m[1970]&~m[1972]&~m[1973])|(~m[1968]&m[1969]&~m[1970]&~m[1972]&~m[1973])|(~m[1968]&~m[1969]&m[1970]&~m[1972]&~m[1973])|(m[1968]&m[1969]&m[1970]&m[1972]&~m[1973])|(~m[1968]&~m[1969]&~m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&~m[1970]&m[1972]&m[1973])|(m[1968]&~m[1969]&m[1970]&m[1972]&m[1973])|(~m[1968]&m[1969]&m[1970]&m[1972]&m[1973]))&UnbiasedRNG[922])|((m[1968]&m[1969]&~m[1970]&~m[1972]&~m[1973])|(m[1968]&~m[1969]&m[1970]&~m[1972]&~m[1973])|(~m[1968]&m[1969]&m[1970]&~m[1972]&~m[1973])|(m[1968]&m[1969]&m[1970]&~m[1972]&~m[1973])|(m[1968]&~m[1969]&~m[1970]&~m[1972]&m[1973])|(~m[1968]&m[1969]&~m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&~m[1970]&~m[1972]&m[1973])|(~m[1968]&~m[1969]&m[1970]&~m[1972]&m[1973])|(m[1968]&~m[1969]&m[1970]&~m[1972]&m[1973])|(~m[1968]&m[1969]&m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&m[1970]&m[1972]&m[1973]));
    m[1976] = (((m[1973]&~m[1974]&~m[1975]&~m[1977]&~m[1978])|(~m[1973]&m[1974]&~m[1975]&~m[1977]&~m[1978])|(~m[1973]&~m[1974]&m[1975]&~m[1977]&~m[1978])|(m[1973]&m[1974]&m[1975]&m[1977]&~m[1978])|(~m[1973]&~m[1974]&~m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&~m[1975]&m[1977]&m[1978])|(m[1973]&~m[1974]&m[1975]&m[1977]&m[1978])|(~m[1973]&m[1974]&m[1975]&m[1977]&m[1978]))&UnbiasedRNG[923])|((m[1973]&m[1974]&~m[1975]&~m[1977]&~m[1978])|(m[1973]&~m[1974]&m[1975]&~m[1977]&~m[1978])|(~m[1973]&m[1974]&m[1975]&~m[1977]&~m[1978])|(m[1973]&m[1974]&m[1975]&~m[1977]&~m[1978])|(m[1973]&~m[1974]&~m[1975]&~m[1977]&m[1978])|(~m[1973]&m[1974]&~m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&~m[1975]&~m[1977]&m[1978])|(~m[1973]&~m[1974]&m[1975]&~m[1977]&m[1978])|(m[1973]&~m[1974]&m[1975]&~m[1977]&m[1978])|(~m[1973]&m[1974]&m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&m[1975]&m[1977]&m[1978]));
    m[1981] = (((m[1978]&~m[1979]&~m[1980]&~m[1982]&~m[1983])|(~m[1978]&m[1979]&~m[1980]&~m[1982]&~m[1983])|(~m[1978]&~m[1979]&m[1980]&~m[1982]&~m[1983])|(m[1978]&m[1979]&m[1980]&m[1982]&~m[1983])|(~m[1978]&~m[1979]&~m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&~m[1980]&m[1982]&m[1983])|(m[1978]&~m[1979]&m[1980]&m[1982]&m[1983])|(~m[1978]&m[1979]&m[1980]&m[1982]&m[1983]))&UnbiasedRNG[924])|((m[1978]&m[1979]&~m[1980]&~m[1982]&~m[1983])|(m[1978]&~m[1979]&m[1980]&~m[1982]&~m[1983])|(~m[1978]&m[1979]&m[1980]&~m[1982]&~m[1983])|(m[1978]&m[1979]&m[1980]&~m[1982]&~m[1983])|(m[1978]&~m[1979]&~m[1980]&~m[1982]&m[1983])|(~m[1978]&m[1979]&~m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&~m[1980]&~m[1982]&m[1983])|(~m[1978]&~m[1979]&m[1980]&~m[1982]&m[1983])|(m[1978]&~m[1979]&m[1980]&~m[1982]&m[1983])|(~m[1978]&m[1979]&m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&m[1980]&m[1982]&m[1983]));
    m[1991] = (((m[1988]&~m[1989]&~m[1990]&~m[1992]&~m[1993])|(~m[1988]&m[1989]&~m[1990]&~m[1992]&~m[1993])|(~m[1988]&~m[1989]&m[1990]&~m[1992]&~m[1993])|(m[1988]&m[1989]&m[1990]&m[1992]&~m[1993])|(~m[1988]&~m[1989]&~m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&~m[1990]&m[1992]&m[1993])|(m[1988]&~m[1989]&m[1990]&m[1992]&m[1993])|(~m[1988]&m[1989]&m[1990]&m[1992]&m[1993]))&UnbiasedRNG[925])|((m[1988]&m[1989]&~m[1990]&~m[1992]&~m[1993])|(m[1988]&~m[1989]&m[1990]&~m[1992]&~m[1993])|(~m[1988]&m[1989]&m[1990]&~m[1992]&~m[1993])|(m[1988]&m[1989]&m[1990]&~m[1992]&~m[1993])|(m[1988]&~m[1989]&~m[1990]&~m[1992]&m[1993])|(~m[1988]&m[1989]&~m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&~m[1990]&~m[1992]&m[1993])|(~m[1988]&~m[1989]&m[1990]&~m[1992]&m[1993])|(m[1988]&~m[1989]&m[1990]&~m[1992]&m[1993])|(~m[1988]&m[1989]&m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&m[1990]&m[1992]&m[1993]));
    m[1996] = (((m[1993]&~m[1994]&~m[1995]&~m[1997]&~m[1998])|(~m[1993]&m[1994]&~m[1995]&~m[1997]&~m[1998])|(~m[1993]&~m[1994]&m[1995]&~m[1997]&~m[1998])|(m[1993]&m[1994]&m[1995]&m[1997]&~m[1998])|(~m[1993]&~m[1994]&~m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&~m[1995]&m[1997]&m[1998])|(m[1993]&~m[1994]&m[1995]&m[1997]&m[1998])|(~m[1993]&m[1994]&m[1995]&m[1997]&m[1998]))&UnbiasedRNG[926])|((m[1993]&m[1994]&~m[1995]&~m[1997]&~m[1998])|(m[1993]&~m[1994]&m[1995]&~m[1997]&~m[1998])|(~m[1993]&m[1994]&m[1995]&~m[1997]&~m[1998])|(m[1993]&m[1994]&m[1995]&~m[1997]&~m[1998])|(m[1993]&~m[1994]&~m[1995]&~m[1997]&m[1998])|(~m[1993]&m[1994]&~m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&~m[1995]&~m[1997]&m[1998])|(~m[1993]&~m[1994]&m[1995]&~m[1997]&m[1998])|(m[1993]&~m[1994]&m[1995]&~m[1997]&m[1998])|(~m[1993]&m[1994]&m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&m[1995]&m[1997]&m[1998]));
    m[2001] = (((m[1998]&~m[1999]&~m[2000]&~m[2002]&~m[2003])|(~m[1998]&m[1999]&~m[2000]&~m[2002]&~m[2003])|(~m[1998]&~m[1999]&m[2000]&~m[2002]&~m[2003])|(m[1998]&m[1999]&m[2000]&m[2002]&~m[2003])|(~m[1998]&~m[1999]&~m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&~m[2000]&m[2002]&m[2003])|(m[1998]&~m[1999]&m[2000]&m[2002]&m[2003])|(~m[1998]&m[1999]&m[2000]&m[2002]&m[2003]))&UnbiasedRNG[927])|((m[1998]&m[1999]&~m[2000]&~m[2002]&~m[2003])|(m[1998]&~m[1999]&m[2000]&~m[2002]&~m[2003])|(~m[1998]&m[1999]&m[2000]&~m[2002]&~m[2003])|(m[1998]&m[1999]&m[2000]&~m[2002]&~m[2003])|(m[1998]&~m[1999]&~m[2000]&~m[2002]&m[2003])|(~m[1998]&m[1999]&~m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&~m[2000]&~m[2002]&m[2003])|(~m[1998]&~m[1999]&m[2000]&~m[2002]&m[2003])|(m[1998]&~m[1999]&m[2000]&~m[2002]&m[2003])|(~m[1998]&m[1999]&m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&m[2000]&m[2002]&m[2003]));
    m[2006] = (((m[2003]&~m[2004]&~m[2005]&~m[2007]&~m[2008])|(~m[2003]&m[2004]&~m[2005]&~m[2007]&~m[2008])|(~m[2003]&~m[2004]&m[2005]&~m[2007]&~m[2008])|(m[2003]&m[2004]&m[2005]&m[2007]&~m[2008])|(~m[2003]&~m[2004]&~m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&~m[2005]&m[2007]&m[2008])|(m[2003]&~m[2004]&m[2005]&m[2007]&m[2008])|(~m[2003]&m[2004]&m[2005]&m[2007]&m[2008]))&UnbiasedRNG[928])|((m[2003]&m[2004]&~m[2005]&~m[2007]&~m[2008])|(m[2003]&~m[2004]&m[2005]&~m[2007]&~m[2008])|(~m[2003]&m[2004]&m[2005]&~m[2007]&~m[2008])|(m[2003]&m[2004]&m[2005]&~m[2007]&~m[2008])|(m[2003]&~m[2004]&~m[2005]&~m[2007]&m[2008])|(~m[2003]&m[2004]&~m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&~m[2005]&~m[2007]&m[2008])|(~m[2003]&~m[2004]&m[2005]&~m[2007]&m[2008])|(m[2003]&~m[2004]&m[2005]&~m[2007]&m[2008])|(~m[2003]&m[2004]&m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&m[2005]&m[2007]&m[2008]));
    m[2011] = (((m[2008]&~m[2009]&~m[2010]&~m[2012]&~m[2013])|(~m[2008]&m[2009]&~m[2010]&~m[2012]&~m[2013])|(~m[2008]&~m[2009]&m[2010]&~m[2012]&~m[2013])|(m[2008]&m[2009]&m[2010]&m[2012]&~m[2013])|(~m[2008]&~m[2009]&~m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&~m[2010]&m[2012]&m[2013])|(m[2008]&~m[2009]&m[2010]&m[2012]&m[2013])|(~m[2008]&m[2009]&m[2010]&m[2012]&m[2013]))&UnbiasedRNG[929])|((m[2008]&m[2009]&~m[2010]&~m[2012]&~m[2013])|(m[2008]&~m[2009]&m[2010]&~m[2012]&~m[2013])|(~m[2008]&m[2009]&m[2010]&~m[2012]&~m[2013])|(m[2008]&m[2009]&m[2010]&~m[2012]&~m[2013])|(m[2008]&~m[2009]&~m[2010]&~m[2012]&m[2013])|(~m[2008]&m[2009]&~m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&~m[2010]&~m[2012]&m[2013])|(~m[2008]&~m[2009]&m[2010]&~m[2012]&m[2013])|(m[2008]&~m[2009]&m[2010]&~m[2012]&m[2013])|(~m[2008]&m[2009]&m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&m[2010]&m[2012]&m[2013]));
    m[2016] = (((m[2013]&~m[2014]&~m[2015]&~m[2017]&~m[2018])|(~m[2013]&m[2014]&~m[2015]&~m[2017]&~m[2018])|(~m[2013]&~m[2014]&m[2015]&~m[2017]&~m[2018])|(m[2013]&m[2014]&m[2015]&m[2017]&~m[2018])|(~m[2013]&~m[2014]&~m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&~m[2015]&m[2017]&m[2018])|(m[2013]&~m[2014]&m[2015]&m[2017]&m[2018])|(~m[2013]&m[2014]&m[2015]&m[2017]&m[2018]))&UnbiasedRNG[930])|((m[2013]&m[2014]&~m[2015]&~m[2017]&~m[2018])|(m[2013]&~m[2014]&m[2015]&~m[2017]&~m[2018])|(~m[2013]&m[2014]&m[2015]&~m[2017]&~m[2018])|(m[2013]&m[2014]&m[2015]&~m[2017]&~m[2018])|(m[2013]&~m[2014]&~m[2015]&~m[2017]&m[2018])|(~m[2013]&m[2014]&~m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&~m[2015]&~m[2017]&m[2018])|(~m[2013]&~m[2014]&m[2015]&~m[2017]&m[2018])|(m[2013]&~m[2014]&m[2015]&~m[2017]&m[2018])|(~m[2013]&m[2014]&m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&m[2015]&m[2017]&m[2018]));
    m[2026] = (((m[2023]&~m[2024]&~m[2025]&~m[2027]&~m[2028])|(~m[2023]&m[2024]&~m[2025]&~m[2027]&~m[2028])|(~m[2023]&~m[2024]&m[2025]&~m[2027]&~m[2028])|(m[2023]&m[2024]&m[2025]&m[2027]&~m[2028])|(~m[2023]&~m[2024]&~m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&~m[2025]&m[2027]&m[2028])|(m[2023]&~m[2024]&m[2025]&m[2027]&m[2028])|(~m[2023]&m[2024]&m[2025]&m[2027]&m[2028]))&UnbiasedRNG[931])|((m[2023]&m[2024]&~m[2025]&~m[2027]&~m[2028])|(m[2023]&~m[2024]&m[2025]&~m[2027]&~m[2028])|(~m[2023]&m[2024]&m[2025]&~m[2027]&~m[2028])|(m[2023]&m[2024]&m[2025]&~m[2027]&~m[2028])|(m[2023]&~m[2024]&~m[2025]&~m[2027]&m[2028])|(~m[2023]&m[2024]&~m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&~m[2025]&~m[2027]&m[2028])|(~m[2023]&~m[2024]&m[2025]&~m[2027]&m[2028])|(m[2023]&~m[2024]&m[2025]&~m[2027]&m[2028])|(~m[2023]&m[2024]&m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&m[2025]&m[2027]&m[2028]));
    m[2031] = (((m[2028]&~m[2029]&~m[2030]&~m[2032]&~m[2033])|(~m[2028]&m[2029]&~m[2030]&~m[2032]&~m[2033])|(~m[2028]&~m[2029]&m[2030]&~m[2032]&~m[2033])|(m[2028]&m[2029]&m[2030]&m[2032]&~m[2033])|(~m[2028]&~m[2029]&~m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&~m[2030]&m[2032]&m[2033])|(m[2028]&~m[2029]&m[2030]&m[2032]&m[2033])|(~m[2028]&m[2029]&m[2030]&m[2032]&m[2033]))&UnbiasedRNG[932])|((m[2028]&m[2029]&~m[2030]&~m[2032]&~m[2033])|(m[2028]&~m[2029]&m[2030]&~m[2032]&~m[2033])|(~m[2028]&m[2029]&m[2030]&~m[2032]&~m[2033])|(m[2028]&m[2029]&m[2030]&~m[2032]&~m[2033])|(m[2028]&~m[2029]&~m[2030]&~m[2032]&m[2033])|(~m[2028]&m[2029]&~m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&~m[2030]&~m[2032]&m[2033])|(~m[2028]&~m[2029]&m[2030]&~m[2032]&m[2033])|(m[2028]&~m[2029]&m[2030]&~m[2032]&m[2033])|(~m[2028]&m[2029]&m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&m[2030]&m[2032]&m[2033]));
    m[2036] = (((m[2033]&~m[2034]&~m[2035]&~m[2037]&~m[2038])|(~m[2033]&m[2034]&~m[2035]&~m[2037]&~m[2038])|(~m[2033]&~m[2034]&m[2035]&~m[2037]&~m[2038])|(m[2033]&m[2034]&m[2035]&m[2037]&~m[2038])|(~m[2033]&~m[2034]&~m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&~m[2035]&m[2037]&m[2038])|(m[2033]&~m[2034]&m[2035]&m[2037]&m[2038])|(~m[2033]&m[2034]&m[2035]&m[2037]&m[2038]))&UnbiasedRNG[933])|((m[2033]&m[2034]&~m[2035]&~m[2037]&~m[2038])|(m[2033]&~m[2034]&m[2035]&~m[2037]&~m[2038])|(~m[2033]&m[2034]&m[2035]&~m[2037]&~m[2038])|(m[2033]&m[2034]&m[2035]&~m[2037]&~m[2038])|(m[2033]&~m[2034]&~m[2035]&~m[2037]&m[2038])|(~m[2033]&m[2034]&~m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&~m[2035]&~m[2037]&m[2038])|(~m[2033]&~m[2034]&m[2035]&~m[2037]&m[2038])|(m[2033]&~m[2034]&m[2035]&~m[2037]&m[2038])|(~m[2033]&m[2034]&m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&m[2035]&m[2037]&m[2038]));
    m[2041] = (((m[2038]&~m[2039]&~m[2040]&~m[2042]&~m[2043])|(~m[2038]&m[2039]&~m[2040]&~m[2042]&~m[2043])|(~m[2038]&~m[2039]&m[2040]&~m[2042]&~m[2043])|(m[2038]&m[2039]&m[2040]&m[2042]&~m[2043])|(~m[2038]&~m[2039]&~m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&~m[2040]&m[2042]&m[2043])|(m[2038]&~m[2039]&m[2040]&m[2042]&m[2043])|(~m[2038]&m[2039]&m[2040]&m[2042]&m[2043]))&UnbiasedRNG[934])|((m[2038]&m[2039]&~m[2040]&~m[2042]&~m[2043])|(m[2038]&~m[2039]&m[2040]&~m[2042]&~m[2043])|(~m[2038]&m[2039]&m[2040]&~m[2042]&~m[2043])|(m[2038]&m[2039]&m[2040]&~m[2042]&~m[2043])|(m[2038]&~m[2039]&~m[2040]&~m[2042]&m[2043])|(~m[2038]&m[2039]&~m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&~m[2040]&~m[2042]&m[2043])|(~m[2038]&~m[2039]&m[2040]&~m[2042]&m[2043])|(m[2038]&~m[2039]&m[2040]&~m[2042]&m[2043])|(~m[2038]&m[2039]&m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&m[2040]&m[2042]&m[2043]));
    m[2046] = (((m[2043]&~m[2044]&~m[2045]&~m[2047]&~m[2048])|(~m[2043]&m[2044]&~m[2045]&~m[2047]&~m[2048])|(~m[2043]&~m[2044]&m[2045]&~m[2047]&~m[2048])|(m[2043]&m[2044]&m[2045]&m[2047]&~m[2048])|(~m[2043]&~m[2044]&~m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&~m[2045]&m[2047]&m[2048])|(m[2043]&~m[2044]&m[2045]&m[2047]&m[2048])|(~m[2043]&m[2044]&m[2045]&m[2047]&m[2048]))&UnbiasedRNG[935])|((m[2043]&m[2044]&~m[2045]&~m[2047]&~m[2048])|(m[2043]&~m[2044]&m[2045]&~m[2047]&~m[2048])|(~m[2043]&m[2044]&m[2045]&~m[2047]&~m[2048])|(m[2043]&m[2044]&m[2045]&~m[2047]&~m[2048])|(m[2043]&~m[2044]&~m[2045]&~m[2047]&m[2048])|(~m[2043]&m[2044]&~m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&~m[2045]&~m[2047]&m[2048])|(~m[2043]&~m[2044]&m[2045]&~m[2047]&m[2048])|(m[2043]&~m[2044]&m[2045]&~m[2047]&m[2048])|(~m[2043]&m[2044]&m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&m[2045]&m[2047]&m[2048]));
    m[2056] = (((m[2053]&~m[2054]&~m[2055]&~m[2057]&~m[2058])|(~m[2053]&m[2054]&~m[2055]&~m[2057]&~m[2058])|(~m[2053]&~m[2054]&m[2055]&~m[2057]&~m[2058])|(m[2053]&m[2054]&m[2055]&m[2057]&~m[2058])|(~m[2053]&~m[2054]&~m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&~m[2055]&m[2057]&m[2058])|(m[2053]&~m[2054]&m[2055]&m[2057]&m[2058])|(~m[2053]&m[2054]&m[2055]&m[2057]&m[2058]))&UnbiasedRNG[936])|((m[2053]&m[2054]&~m[2055]&~m[2057]&~m[2058])|(m[2053]&~m[2054]&m[2055]&~m[2057]&~m[2058])|(~m[2053]&m[2054]&m[2055]&~m[2057]&~m[2058])|(m[2053]&m[2054]&m[2055]&~m[2057]&~m[2058])|(m[2053]&~m[2054]&~m[2055]&~m[2057]&m[2058])|(~m[2053]&m[2054]&~m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&~m[2055]&~m[2057]&m[2058])|(~m[2053]&~m[2054]&m[2055]&~m[2057]&m[2058])|(m[2053]&~m[2054]&m[2055]&~m[2057]&m[2058])|(~m[2053]&m[2054]&m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&m[2055]&m[2057]&m[2058]));
    m[2061] = (((m[2058]&~m[2059]&~m[2060]&~m[2062]&~m[2063])|(~m[2058]&m[2059]&~m[2060]&~m[2062]&~m[2063])|(~m[2058]&~m[2059]&m[2060]&~m[2062]&~m[2063])|(m[2058]&m[2059]&m[2060]&m[2062]&~m[2063])|(~m[2058]&~m[2059]&~m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&~m[2060]&m[2062]&m[2063])|(m[2058]&~m[2059]&m[2060]&m[2062]&m[2063])|(~m[2058]&m[2059]&m[2060]&m[2062]&m[2063]))&UnbiasedRNG[937])|((m[2058]&m[2059]&~m[2060]&~m[2062]&~m[2063])|(m[2058]&~m[2059]&m[2060]&~m[2062]&~m[2063])|(~m[2058]&m[2059]&m[2060]&~m[2062]&~m[2063])|(m[2058]&m[2059]&m[2060]&~m[2062]&~m[2063])|(m[2058]&~m[2059]&~m[2060]&~m[2062]&m[2063])|(~m[2058]&m[2059]&~m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&~m[2060]&~m[2062]&m[2063])|(~m[2058]&~m[2059]&m[2060]&~m[2062]&m[2063])|(m[2058]&~m[2059]&m[2060]&~m[2062]&m[2063])|(~m[2058]&m[2059]&m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&m[2060]&m[2062]&m[2063]));
    m[2066] = (((m[2063]&~m[2064]&~m[2065]&~m[2067]&~m[2068])|(~m[2063]&m[2064]&~m[2065]&~m[2067]&~m[2068])|(~m[2063]&~m[2064]&m[2065]&~m[2067]&~m[2068])|(m[2063]&m[2064]&m[2065]&m[2067]&~m[2068])|(~m[2063]&~m[2064]&~m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&~m[2065]&m[2067]&m[2068])|(m[2063]&~m[2064]&m[2065]&m[2067]&m[2068])|(~m[2063]&m[2064]&m[2065]&m[2067]&m[2068]))&UnbiasedRNG[938])|((m[2063]&m[2064]&~m[2065]&~m[2067]&~m[2068])|(m[2063]&~m[2064]&m[2065]&~m[2067]&~m[2068])|(~m[2063]&m[2064]&m[2065]&~m[2067]&~m[2068])|(m[2063]&m[2064]&m[2065]&~m[2067]&~m[2068])|(m[2063]&~m[2064]&~m[2065]&~m[2067]&m[2068])|(~m[2063]&m[2064]&~m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&~m[2065]&~m[2067]&m[2068])|(~m[2063]&~m[2064]&m[2065]&~m[2067]&m[2068])|(m[2063]&~m[2064]&m[2065]&~m[2067]&m[2068])|(~m[2063]&m[2064]&m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&m[2065]&m[2067]&m[2068]));
    m[2071] = (((m[2068]&~m[2069]&~m[2070]&~m[2072]&~m[2073])|(~m[2068]&m[2069]&~m[2070]&~m[2072]&~m[2073])|(~m[2068]&~m[2069]&m[2070]&~m[2072]&~m[2073])|(m[2068]&m[2069]&m[2070]&m[2072]&~m[2073])|(~m[2068]&~m[2069]&~m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&~m[2070]&m[2072]&m[2073])|(m[2068]&~m[2069]&m[2070]&m[2072]&m[2073])|(~m[2068]&m[2069]&m[2070]&m[2072]&m[2073]))&UnbiasedRNG[939])|((m[2068]&m[2069]&~m[2070]&~m[2072]&~m[2073])|(m[2068]&~m[2069]&m[2070]&~m[2072]&~m[2073])|(~m[2068]&m[2069]&m[2070]&~m[2072]&~m[2073])|(m[2068]&m[2069]&m[2070]&~m[2072]&~m[2073])|(m[2068]&~m[2069]&~m[2070]&~m[2072]&m[2073])|(~m[2068]&m[2069]&~m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&~m[2070]&~m[2072]&m[2073])|(~m[2068]&~m[2069]&m[2070]&~m[2072]&m[2073])|(m[2068]&~m[2069]&m[2070]&~m[2072]&m[2073])|(~m[2068]&m[2069]&m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&m[2070]&m[2072]&m[2073]));
    m[2081] = (((m[2078]&~m[2079]&~m[2080]&~m[2082]&~m[2083])|(~m[2078]&m[2079]&~m[2080]&~m[2082]&~m[2083])|(~m[2078]&~m[2079]&m[2080]&~m[2082]&~m[2083])|(m[2078]&m[2079]&m[2080]&m[2082]&~m[2083])|(~m[2078]&~m[2079]&~m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&~m[2080]&m[2082]&m[2083])|(m[2078]&~m[2079]&m[2080]&m[2082]&m[2083])|(~m[2078]&m[2079]&m[2080]&m[2082]&m[2083]))&UnbiasedRNG[940])|((m[2078]&m[2079]&~m[2080]&~m[2082]&~m[2083])|(m[2078]&~m[2079]&m[2080]&~m[2082]&~m[2083])|(~m[2078]&m[2079]&m[2080]&~m[2082]&~m[2083])|(m[2078]&m[2079]&m[2080]&~m[2082]&~m[2083])|(m[2078]&~m[2079]&~m[2080]&~m[2082]&m[2083])|(~m[2078]&m[2079]&~m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&~m[2080]&~m[2082]&m[2083])|(~m[2078]&~m[2079]&m[2080]&~m[2082]&m[2083])|(m[2078]&~m[2079]&m[2080]&~m[2082]&m[2083])|(~m[2078]&m[2079]&m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&m[2080]&m[2082]&m[2083]));
    m[2086] = (((m[2083]&~m[2084]&~m[2085]&~m[2087]&~m[2088])|(~m[2083]&m[2084]&~m[2085]&~m[2087]&~m[2088])|(~m[2083]&~m[2084]&m[2085]&~m[2087]&~m[2088])|(m[2083]&m[2084]&m[2085]&m[2087]&~m[2088])|(~m[2083]&~m[2084]&~m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&~m[2085]&m[2087]&m[2088])|(m[2083]&~m[2084]&m[2085]&m[2087]&m[2088])|(~m[2083]&m[2084]&m[2085]&m[2087]&m[2088]))&UnbiasedRNG[941])|((m[2083]&m[2084]&~m[2085]&~m[2087]&~m[2088])|(m[2083]&~m[2084]&m[2085]&~m[2087]&~m[2088])|(~m[2083]&m[2084]&m[2085]&~m[2087]&~m[2088])|(m[2083]&m[2084]&m[2085]&~m[2087]&~m[2088])|(m[2083]&~m[2084]&~m[2085]&~m[2087]&m[2088])|(~m[2083]&m[2084]&~m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&~m[2085]&~m[2087]&m[2088])|(~m[2083]&~m[2084]&m[2085]&~m[2087]&m[2088])|(m[2083]&~m[2084]&m[2085]&~m[2087]&m[2088])|(~m[2083]&m[2084]&m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&m[2085]&m[2087]&m[2088]));
    m[2091] = (((m[2088]&~m[2089]&~m[2090]&~m[2092]&~m[2093])|(~m[2088]&m[2089]&~m[2090]&~m[2092]&~m[2093])|(~m[2088]&~m[2089]&m[2090]&~m[2092]&~m[2093])|(m[2088]&m[2089]&m[2090]&m[2092]&~m[2093])|(~m[2088]&~m[2089]&~m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&~m[2090]&m[2092]&m[2093])|(m[2088]&~m[2089]&m[2090]&m[2092]&m[2093])|(~m[2088]&m[2089]&m[2090]&m[2092]&m[2093]))&UnbiasedRNG[942])|((m[2088]&m[2089]&~m[2090]&~m[2092]&~m[2093])|(m[2088]&~m[2089]&m[2090]&~m[2092]&~m[2093])|(~m[2088]&m[2089]&m[2090]&~m[2092]&~m[2093])|(m[2088]&m[2089]&m[2090]&~m[2092]&~m[2093])|(m[2088]&~m[2089]&~m[2090]&~m[2092]&m[2093])|(~m[2088]&m[2089]&~m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&~m[2090]&~m[2092]&m[2093])|(~m[2088]&~m[2089]&m[2090]&~m[2092]&m[2093])|(m[2088]&~m[2089]&m[2090]&~m[2092]&m[2093])|(~m[2088]&m[2089]&m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&m[2090]&m[2092]&m[2093]));
    m[2101] = (((m[2098]&~m[2099]&~m[2100]&~m[2102]&~m[2103])|(~m[2098]&m[2099]&~m[2100]&~m[2102]&~m[2103])|(~m[2098]&~m[2099]&m[2100]&~m[2102]&~m[2103])|(m[2098]&m[2099]&m[2100]&m[2102]&~m[2103])|(~m[2098]&~m[2099]&~m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&~m[2100]&m[2102]&m[2103])|(m[2098]&~m[2099]&m[2100]&m[2102]&m[2103])|(~m[2098]&m[2099]&m[2100]&m[2102]&m[2103]))&UnbiasedRNG[943])|((m[2098]&m[2099]&~m[2100]&~m[2102]&~m[2103])|(m[2098]&~m[2099]&m[2100]&~m[2102]&~m[2103])|(~m[2098]&m[2099]&m[2100]&~m[2102]&~m[2103])|(m[2098]&m[2099]&m[2100]&~m[2102]&~m[2103])|(m[2098]&~m[2099]&~m[2100]&~m[2102]&m[2103])|(~m[2098]&m[2099]&~m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&~m[2100]&~m[2102]&m[2103])|(~m[2098]&~m[2099]&m[2100]&~m[2102]&m[2103])|(m[2098]&~m[2099]&m[2100]&~m[2102]&m[2103])|(~m[2098]&m[2099]&m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&m[2100]&m[2102]&m[2103]));
    m[2106] = (((m[2103]&~m[2104]&~m[2105]&~m[2107]&~m[2108])|(~m[2103]&m[2104]&~m[2105]&~m[2107]&~m[2108])|(~m[2103]&~m[2104]&m[2105]&~m[2107]&~m[2108])|(m[2103]&m[2104]&m[2105]&m[2107]&~m[2108])|(~m[2103]&~m[2104]&~m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&~m[2105]&m[2107]&m[2108])|(m[2103]&~m[2104]&m[2105]&m[2107]&m[2108])|(~m[2103]&m[2104]&m[2105]&m[2107]&m[2108]))&UnbiasedRNG[944])|((m[2103]&m[2104]&~m[2105]&~m[2107]&~m[2108])|(m[2103]&~m[2104]&m[2105]&~m[2107]&~m[2108])|(~m[2103]&m[2104]&m[2105]&~m[2107]&~m[2108])|(m[2103]&m[2104]&m[2105]&~m[2107]&~m[2108])|(m[2103]&~m[2104]&~m[2105]&~m[2107]&m[2108])|(~m[2103]&m[2104]&~m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&~m[2105]&~m[2107]&m[2108])|(~m[2103]&~m[2104]&m[2105]&~m[2107]&m[2108])|(m[2103]&~m[2104]&m[2105]&~m[2107]&m[2108])|(~m[2103]&m[2104]&m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&m[2105]&m[2107]&m[2108]));
    m[2116] = (((m[2113]&~m[2114]&~m[2115]&~m[2117]&~m[2118])|(~m[2113]&m[2114]&~m[2115]&~m[2117]&~m[2118])|(~m[2113]&~m[2114]&m[2115]&~m[2117]&~m[2118])|(m[2113]&m[2114]&m[2115]&m[2117]&~m[2118])|(~m[2113]&~m[2114]&~m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&~m[2115]&m[2117]&m[2118])|(m[2113]&~m[2114]&m[2115]&m[2117]&m[2118])|(~m[2113]&m[2114]&m[2115]&m[2117]&m[2118]))&UnbiasedRNG[945])|((m[2113]&m[2114]&~m[2115]&~m[2117]&~m[2118])|(m[2113]&~m[2114]&m[2115]&~m[2117]&~m[2118])|(~m[2113]&m[2114]&m[2115]&~m[2117]&~m[2118])|(m[2113]&m[2114]&m[2115]&~m[2117]&~m[2118])|(m[2113]&~m[2114]&~m[2115]&~m[2117]&m[2118])|(~m[2113]&m[2114]&~m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&~m[2115]&~m[2117]&m[2118])|(~m[2113]&~m[2114]&m[2115]&~m[2117]&m[2118])|(m[2113]&~m[2114]&m[2115]&~m[2117]&m[2118])|(~m[2113]&m[2114]&m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&m[2115]&m[2117]&m[2118]));
end

always @(posedge color4_clk) begin
    m[932] = (((m[928]&~m[929]&~m[930]&~m[931]&~m[935])|(~m[928]&m[929]&~m[930]&~m[931]&~m[935])|(~m[928]&~m[929]&m[930]&~m[931]&~m[935])|(m[928]&m[929]&~m[930]&m[931]&~m[935])|(m[928]&~m[929]&m[930]&m[931]&~m[935])|(~m[928]&m[929]&m[930]&m[931]&~m[935]))&BiasedRNG[895])|(((m[928]&~m[929]&~m[930]&~m[931]&m[935])|(~m[928]&m[929]&~m[930]&~m[931]&m[935])|(~m[928]&~m[929]&m[930]&~m[931]&m[935])|(m[928]&m[929]&~m[930]&m[931]&m[935])|(m[928]&~m[929]&m[930]&m[931]&m[935])|(~m[928]&m[929]&m[930]&m[931]&m[935]))&~BiasedRNG[895])|((m[928]&m[929]&~m[930]&~m[931]&~m[935])|(m[928]&~m[929]&m[930]&~m[931]&~m[935])|(~m[928]&m[929]&m[930]&~m[931]&~m[935])|(m[928]&m[929]&m[930]&~m[931]&~m[935])|(m[928]&m[929]&m[930]&m[931]&~m[935])|(m[928]&m[929]&~m[930]&~m[931]&m[935])|(m[928]&~m[929]&m[930]&~m[931]&m[935])|(~m[928]&m[929]&m[930]&~m[931]&m[935])|(m[928]&m[929]&m[930]&~m[931]&m[935])|(m[928]&m[929]&m[930]&m[931]&m[935]));
    m[937] = (((m[933]&~m[934]&~m[935]&~m[936]&~m[945])|(~m[933]&m[934]&~m[935]&~m[936]&~m[945])|(~m[933]&~m[934]&m[935]&~m[936]&~m[945])|(m[933]&m[934]&~m[935]&m[936]&~m[945])|(m[933]&~m[934]&m[935]&m[936]&~m[945])|(~m[933]&m[934]&m[935]&m[936]&~m[945]))&BiasedRNG[896])|(((m[933]&~m[934]&~m[935]&~m[936]&m[945])|(~m[933]&m[934]&~m[935]&~m[936]&m[945])|(~m[933]&~m[934]&m[935]&~m[936]&m[945])|(m[933]&m[934]&~m[935]&m[936]&m[945])|(m[933]&~m[934]&m[935]&m[936]&m[945])|(~m[933]&m[934]&m[935]&m[936]&m[945]))&~BiasedRNG[896])|((m[933]&m[934]&~m[935]&~m[936]&~m[945])|(m[933]&~m[934]&m[935]&~m[936]&~m[945])|(~m[933]&m[934]&m[935]&~m[936]&~m[945])|(m[933]&m[934]&m[935]&~m[936]&~m[945])|(m[933]&m[934]&m[935]&m[936]&~m[945])|(m[933]&m[934]&~m[935]&~m[936]&m[945])|(m[933]&~m[934]&m[935]&~m[936]&m[945])|(~m[933]&m[934]&m[935]&~m[936]&m[945])|(m[933]&m[934]&m[935]&~m[936]&m[945])|(m[933]&m[934]&m[935]&m[936]&m[945]));
    m[942] = (((m[938]&~m[939]&~m[940]&~m[941]&~m[950])|(~m[938]&m[939]&~m[940]&~m[941]&~m[950])|(~m[938]&~m[939]&m[940]&~m[941]&~m[950])|(m[938]&m[939]&~m[940]&m[941]&~m[950])|(m[938]&~m[939]&m[940]&m[941]&~m[950])|(~m[938]&m[939]&m[940]&m[941]&~m[950]))&BiasedRNG[897])|(((m[938]&~m[939]&~m[940]&~m[941]&m[950])|(~m[938]&m[939]&~m[940]&~m[941]&m[950])|(~m[938]&~m[939]&m[940]&~m[941]&m[950])|(m[938]&m[939]&~m[940]&m[941]&m[950])|(m[938]&~m[939]&m[940]&m[941]&m[950])|(~m[938]&m[939]&m[940]&m[941]&m[950]))&~BiasedRNG[897])|((m[938]&m[939]&~m[940]&~m[941]&~m[950])|(m[938]&~m[939]&m[940]&~m[941]&~m[950])|(~m[938]&m[939]&m[940]&~m[941]&~m[950])|(m[938]&m[939]&m[940]&~m[941]&~m[950])|(m[938]&m[939]&m[940]&m[941]&~m[950])|(m[938]&m[939]&~m[940]&~m[941]&m[950])|(m[938]&~m[939]&m[940]&~m[941]&m[950])|(~m[938]&m[939]&m[940]&~m[941]&m[950])|(m[938]&m[939]&m[940]&~m[941]&m[950])|(m[938]&m[939]&m[940]&m[941]&m[950]));
    m[947] = (((m[943]&~m[944]&~m[945]&~m[946]&~m[960])|(~m[943]&m[944]&~m[945]&~m[946]&~m[960])|(~m[943]&~m[944]&m[945]&~m[946]&~m[960])|(m[943]&m[944]&~m[945]&m[946]&~m[960])|(m[943]&~m[944]&m[945]&m[946]&~m[960])|(~m[943]&m[944]&m[945]&m[946]&~m[960]))&BiasedRNG[898])|(((m[943]&~m[944]&~m[945]&~m[946]&m[960])|(~m[943]&m[944]&~m[945]&~m[946]&m[960])|(~m[943]&~m[944]&m[945]&~m[946]&m[960])|(m[943]&m[944]&~m[945]&m[946]&m[960])|(m[943]&~m[944]&m[945]&m[946]&m[960])|(~m[943]&m[944]&m[945]&m[946]&m[960]))&~BiasedRNG[898])|((m[943]&m[944]&~m[945]&~m[946]&~m[960])|(m[943]&~m[944]&m[945]&~m[946]&~m[960])|(~m[943]&m[944]&m[945]&~m[946]&~m[960])|(m[943]&m[944]&m[945]&~m[946]&~m[960])|(m[943]&m[944]&m[945]&m[946]&~m[960])|(m[943]&m[944]&~m[945]&~m[946]&m[960])|(m[943]&~m[944]&m[945]&~m[946]&m[960])|(~m[943]&m[944]&m[945]&~m[946]&m[960])|(m[943]&m[944]&m[945]&~m[946]&m[960])|(m[943]&m[944]&m[945]&m[946]&m[960]));
    m[952] = (((m[948]&~m[949]&~m[950]&~m[951]&~m[965])|(~m[948]&m[949]&~m[950]&~m[951]&~m[965])|(~m[948]&~m[949]&m[950]&~m[951]&~m[965])|(m[948]&m[949]&~m[950]&m[951]&~m[965])|(m[948]&~m[949]&m[950]&m[951]&~m[965])|(~m[948]&m[949]&m[950]&m[951]&~m[965]))&BiasedRNG[899])|(((m[948]&~m[949]&~m[950]&~m[951]&m[965])|(~m[948]&m[949]&~m[950]&~m[951]&m[965])|(~m[948]&~m[949]&m[950]&~m[951]&m[965])|(m[948]&m[949]&~m[950]&m[951]&m[965])|(m[948]&~m[949]&m[950]&m[951]&m[965])|(~m[948]&m[949]&m[950]&m[951]&m[965]))&~BiasedRNG[899])|((m[948]&m[949]&~m[950]&~m[951]&~m[965])|(m[948]&~m[949]&m[950]&~m[951]&~m[965])|(~m[948]&m[949]&m[950]&~m[951]&~m[965])|(m[948]&m[949]&m[950]&~m[951]&~m[965])|(m[948]&m[949]&m[950]&m[951]&~m[965])|(m[948]&m[949]&~m[950]&~m[951]&m[965])|(m[948]&~m[949]&m[950]&~m[951]&m[965])|(~m[948]&m[949]&m[950]&~m[951]&m[965])|(m[948]&m[949]&m[950]&~m[951]&m[965])|(m[948]&m[949]&m[950]&m[951]&m[965]));
    m[957] = (((m[953]&~m[954]&~m[955]&~m[956]&~m[970])|(~m[953]&m[954]&~m[955]&~m[956]&~m[970])|(~m[953]&~m[954]&m[955]&~m[956]&~m[970])|(m[953]&m[954]&~m[955]&m[956]&~m[970])|(m[953]&~m[954]&m[955]&m[956]&~m[970])|(~m[953]&m[954]&m[955]&m[956]&~m[970]))&BiasedRNG[900])|(((m[953]&~m[954]&~m[955]&~m[956]&m[970])|(~m[953]&m[954]&~m[955]&~m[956]&m[970])|(~m[953]&~m[954]&m[955]&~m[956]&m[970])|(m[953]&m[954]&~m[955]&m[956]&m[970])|(m[953]&~m[954]&m[955]&m[956]&m[970])|(~m[953]&m[954]&m[955]&m[956]&m[970]))&~BiasedRNG[900])|((m[953]&m[954]&~m[955]&~m[956]&~m[970])|(m[953]&~m[954]&m[955]&~m[956]&~m[970])|(~m[953]&m[954]&m[955]&~m[956]&~m[970])|(m[953]&m[954]&m[955]&~m[956]&~m[970])|(m[953]&m[954]&m[955]&m[956]&~m[970])|(m[953]&m[954]&~m[955]&~m[956]&m[970])|(m[953]&~m[954]&m[955]&~m[956]&m[970])|(~m[953]&m[954]&m[955]&~m[956]&m[970])|(m[953]&m[954]&m[955]&~m[956]&m[970])|(m[953]&m[954]&m[955]&m[956]&m[970]));
    m[962] = (((m[958]&~m[959]&~m[960]&~m[961]&~m[980])|(~m[958]&m[959]&~m[960]&~m[961]&~m[980])|(~m[958]&~m[959]&m[960]&~m[961]&~m[980])|(m[958]&m[959]&~m[960]&m[961]&~m[980])|(m[958]&~m[959]&m[960]&m[961]&~m[980])|(~m[958]&m[959]&m[960]&m[961]&~m[980]))&BiasedRNG[901])|(((m[958]&~m[959]&~m[960]&~m[961]&m[980])|(~m[958]&m[959]&~m[960]&~m[961]&m[980])|(~m[958]&~m[959]&m[960]&~m[961]&m[980])|(m[958]&m[959]&~m[960]&m[961]&m[980])|(m[958]&~m[959]&m[960]&m[961]&m[980])|(~m[958]&m[959]&m[960]&m[961]&m[980]))&~BiasedRNG[901])|((m[958]&m[959]&~m[960]&~m[961]&~m[980])|(m[958]&~m[959]&m[960]&~m[961]&~m[980])|(~m[958]&m[959]&m[960]&~m[961]&~m[980])|(m[958]&m[959]&m[960]&~m[961]&~m[980])|(m[958]&m[959]&m[960]&m[961]&~m[980])|(m[958]&m[959]&~m[960]&~m[961]&m[980])|(m[958]&~m[959]&m[960]&~m[961]&m[980])|(~m[958]&m[959]&m[960]&~m[961]&m[980])|(m[958]&m[959]&m[960]&~m[961]&m[980])|(m[958]&m[959]&m[960]&m[961]&m[980]));
    m[967] = (((m[963]&~m[964]&~m[965]&~m[966]&~m[985])|(~m[963]&m[964]&~m[965]&~m[966]&~m[985])|(~m[963]&~m[964]&m[965]&~m[966]&~m[985])|(m[963]&m[964]&~m[965]&m[966]&~m[985])|(m[963]&~m[964]&m[965]&m[966]&~m[985])|(~m[963]&m[964]&m[965]&m[966]&~m[985]))&BiasedRNG[902])|(((m[963]&~m[964]&~m[965]&~m[966]&m[985])|(~m[963]&m[964]&~m[965]&~m[966]&m[985])|(~m[963]&~m[964]&m[965]&~m[966]&m[985])|(m[963]&m[964]&~m[965]&m[966]&m[985])|(m[963]&~m[964]&m[965]&m[966]&m[985])|(~m[963]&m[964]&m[965]&m[966]&m[985]))&~BiasedRNG[902])|((m[963]&m[964]&~m[965]&~m[966]&~m[985])|(m[963]&~m[964]&m[965]&~m[966]&~m[985])|(~m[963]&m[964]&m[965]&~m[966]&~m[985])|(m[963]&m[964]&m[965]&~m[966]&~m[985])|(m[963]&m[964]&m[965]&m[966]&~m[985])|(m[963]&m[964]&~m[965]&~m[966]&m[985])|(m[963]&~m[964]&m[965]&~m[966]&m[985])|(~m[963]&m[964]&m[965]&~m[966]&m[985])|(m[963]&m[964]&m[965]&~m[966]&m[985])|(m[963]&m[964]&m[965]&m[966]&m[985]));
    m[972] = (((m[968]&~m[969]&~m[970]&~m[971]&~m[990])|(~m[968]&m[969]&~m[970]&~m[971]&~m[990])|(~m[968]&~m[969]&m[970]&~m[971]&~m[990])|(m[968]&m[969]&~m[970]&m[971]&~m[990])|(m[968]&~m[969]&m[970]&m[971]&~m[990])|(~m[968]&m[969]&m[970]&m[971]&~m[990]))&BiasedRNG[903])|(((m[968]&~m[969]&~m[970]&~m[971]&m[990])|(~m[968]&m[969]&~m[970]&~m[971]&m[990])|(~m[968]&~m[969]&m[970]&~m[971]&m[990])|(m[968]&m[969]&~m[970]&m[971]&m[990])|(m[968]&~m[969]&m[970]&m[971]&m[990])|(~m[968]&m[969]&m[970]&m[971]&m[990]))&~BiasedRNG[903])|((m[968]&m[969]&~m[970]&~m[971]&~m[990])|(m[968]&~m[969]&m[970]&~m[971]&~m[990])|(~m[968]&m[969]&m[970]&~m[971]&~m[990])|(m[968]&m[969]&m[970]&~m[971]&~m[990])|(m[968]&m[969]&m[970]&m[971]&~m[990])|(m[968]&m[969]&~m[970]&~m[971]&m[990])|(m[968]&~m[969]&m[970]&~m[971]&m[990])|(~m[968]&m[969]&m[970]&~m[971]&m[990])|(m[968]&m[969]&m[970]&~m[971]&m[990])|(m[968]&m[969]&m[970]&m[971]&m[990]));
    m[977] = (((m[973]&~m[974]&~m[975]&~m[976]&~m[995])|(~m[973]&m[974]&~m[975]&~m[976]&~m[995])|(~m[973]&~m[974]&m[975]&~m[976]&~m[995])|(m[973]&m[974]&~m[975]&m[976]&~m[995])|(m[973]&~m[974]&m[975]&m[976]&~m[995])|(~m[973]&m[974]&m[975]&m[976]&~m[995]))&BiasedRNG[904])|(((m[973]&~m[974]&~m[975]&~m[976]&m[995])|(~m[973]&m[974]&~m[975]&~m[976]&m[995])|(~m[973]&~m[974]&m[975]&~m[976]&m[995])|(m[973]&m[974]&~m[975]&m[976]&m[995])|(m[973]&~m[974]&m[975]&m[976]&m[995])|(~m[973]&m[974]&m[975]&m[976]&m[995]))&~BiasedRNG[904])|((m[973]&m[974]&~m[975]&~m[976]&~m[995])|(m[973]&~m[974]&m[975]&~m[976]&~m[995])|(~m[973]&m[974]&m[975]&~m[976]&~m[995])|(m[973]&m[974]&m[975]&~m[976]&~m[995])|(m[973]&m[974]&m[975]&m[976]&~m[995])|(m[973]&m[974]&~m[975]&~m[976]&m[995])|(m[973]&~m[974]&m[975]&~m[976]&m[995])|(~m[973]&m[974]&m[975]&~m[976]&m[995])|(m[973]&m[974]&m[975]&~m[976]&m[995])|(m[973]&m[974]&m[975]&m[976]&m[995]));
    m[982] = (((m[978]&~m[979]&~m[980]&~m[981]&~m[1005])|(~m[978]&m[979]&~m[980]&~m[981]&~m[1005])|(~m[978]&~m[979]&m[980]&~m[981]&~m[1005])|(m[978]&m[979]&~m[980]&m[981]&~m[1005])|(m[978]&~m[979]&m[980]&m[981]&~m[1005])|(~m[978]&m[979]&m[980]&m[981]&~m[1005]))&BiasedRNG[905])|(((m[978]&~m[979]&~m[980]&~m[981]&m[1005])|(~m[978]&m[979]&~m[980]&~m[981]&m[1005])|(~m[978]&~m[979]&m[980]&~m[981]&m[1005])|(m[978]&m[979]&~m[980]&m[981]&m[1005])|(m[978]&~m[979]&m[980]&m[981]&m[1005])|(~m[978]&m[979]&m[980]&m[981]&m[1005]))&~BiasedRNG[905])|((m[978]&m[979]&~m[980]&~m[981]&~m[1005])|(m[978]&~m[979]&m[980]&~m[981]&~m[1005])|(~m[978]&m[979]&m[980]&~m[981]&~m[1005])|(m[978]&m[979]&m[980]&~m[981]&~m[1005])|(m[978]&m[979]&m[980]&m[981]&~m[1005])|(m[978]&m[979]&~m[980]&~m[981]&m[1005])|(m[978]&~m[979]&m[980]&~m[981]&m[1005])|(~m[978]&m[979]&m[980]&~m[981]&m[1005])|(m[978]&m[979]&m[980]&~m[981]&m[1005])|(m[978]&m[979]&m[980]&m[981]&m[1005]));
    m[987] = (((m[983]&~m[984]&~m[985]&~m[986]&~m[1010])|(~m[983]&m[984]&~m[985]&~m[986]&~m[1010])|(~m[983]&~m[984]&m[985]&~m[986]&~m[1010])|(m[983]&m[984]&~m[985]&m[986]&~m[1010])|(m[983]&~m[984]&m[985]&m[986]&~m[1010])|(~m[983]&m[984]&m[985]&m[986]&~m[1010]))&BiasedRNG[906])|(((m[983]&~m[984]&~m[985]&~m[986]&m[1010])|(~m[983]&m[984]&~m[985]&~m[986]&m[1010])|(~m[983]&~m[984]&m[985]&~m[986]&m[1010])|(m[983]&m[984]&~m[985]&m[986]&m[1010])|(m[983]&~m[984]&m[985]&m[986]&m[1010])|(~m[983]&m[984]&m[985]&m[986]&m[1010]))&~BiasedRNG[906])|((m[983]&m[984]&~m[985]&~m[986]&~m[1010])|(m[983]&~m[984]&m[985]&~m[986]&~m[1010])|(~m[983]&m[984]&m[985]&~m[986]&~m[1010])|(m[983]&m[984]&m[985]&~m[986]&~m[1010])|(m[983]&m[984]&m[985]&m[986]&~m[1010])|(m[983]&m[984]&~m[985]&~m[986]&m[1010])|(m[983]&~m[984]&m[985]&~m[986]&m[1010])|(~m[983]&m[984]&m[985]&~m[986]&m[1010])|(m[983]&m[984]&m[985]&~m[986]&m[1010])|(m[983]&m[984]&m[985]&m[986]&m[1010]));
    m[992] = (((m[988]&~m[989]&~m[990]&~m[991]&~m[1015])|(~m[988]&m[989]&~m[990]&~m[991]&~m[1015])|(~m[988]&~m[989]&m[990]&~m[991]&~m[1015])|(m[988]&m[989]&~m[990]&m[991]&~m[1015])|(m[988]&~m[989]&m[990]&m[991]&~m[1015])|(~m[988]&m[989]&m[990]&m[991]&~m[1015]))&BiasedRNG[907])|(((m[988]&~m[989]&~m[990]&~m[991]&m[1015])|(~m[988]&m[989]&~m[990]&~m[991]&m[1015])|(~m[988]&~m[989]&m[990]&~m[991]&m[1015])|(m[988]&m[989]&~m[990]&m[991]&m[1015])|(m[988]&~m[989]&m[990]&m[991]&m[1015])|(~m[988]&m[989]&m[990]&m[991]&m[1015]))&~BiasedRNG[907])|((m[988]&m[989]&~m[990]&~m[991]&~m[1015])|(m[988]&~m[989]&m[990]&~m[991]&~m[1015])|(~m[988]&m[989]&m[990]&~m[991]&~m[1015])|(m[988]&m[989]&m[990]&~m[991]&~m[1015])|(m[988]&m[989]&m[990]&m[991]&~m[1015])|(m[988]&m[989]&~m[990]&~m[991]&m[1015])|(m[988]&~m[989]&m[990]&~m[991]&m[1015])|(~m[988]&m[989]&m[990]&~m[991]&m[1015])|(m[988]&m[989]&m[990]&~m[991]&m[1015])|(m[988]&m[989]&m[990]&m[991]&m[1015]));
    m[997] = (((m[993]&~m[994]&~m[995]&~m[996]&~m[1020])|(~m[993]&m[994]&~m[995]&~m[996]&~m[1020])|(~m[993]&~m[994]&m[995]&~m[996]&~m[1020])|(m[993]&m[994]&~m[995]&m[996]&~m[1020])|(m[993]&~m[994]&m[995]&m[996]&~m[1020])|(~m[993]&m[994]&m[995]&m[996]&~m[1020]))&BiasedRNG[908])|(((m[993]&~m[994]&~m[995]&~m[996]&m[1020])|(~m[993]&m[994]&~m[995]&~m[996]&m[1020])|(~m[993]&~m[994]&m[995]&~m[996]&m[1020])|(m[993]&m[994]&~m[995]&m[996]&m[1020])|(m[993]&~m[994]&m[995]&m[996]&m[1020])|(~m[993]&m[994]&m[995]&m[996]&m[1020]))&~BiasedRNG[908])|((m[993]&m[994]&~m[995]&~m[996]&~m[1020])|(m[993]&~m[994]&m[995]&~m[996]&~m[1020])|(~m[993]&m[994]&m[995]&~m[996]&~m[1020])|(m[993]&m[994]&m[995]&~m[996]&~m[1020])|(m[993]&m[994]&m[995]&m[996]&~m[1020])|(m[993]&m[994]&~m[995]&~m[996]&m[1020])|(m[993]&~m[994]&m[995]&~m[996]&m[1020])|(~m[993]&m[994]&m[995]&~m[996]&m[1020])|(m[993]&m[994]&m[995]&~m[996]&m[1020])|(m[993]&m[994]&m[995]&m[996]&m[1020]));
    m[1002] = (((m[998]&~m[999]&~m[1000]&~m[1001]&~m[1025])|(~m[998]&m[999]&~m[1000]&~m[1001]&~m[1025])|(~m[998]&~m[999]&m[1000]&~m[1001]&~m[1025])|(m[998]&m[999]&~m[1000]&m[1001]&~m[1025])|(m[998]&~m[999]&m[1000]&m[1001]&~m[1025])|(~m[998]&m[999]&m[1000]&m[1001]&~m[1025]))&BiasedRNG[909])|(((m[998]&~m[999]&~m[1000]&~m[1001]&m[1025])|(~m[998]&m[999]&~m[1000]&~m[1001]&m[1025])|(~m[998]&~m[999]&m[1000]&~m[1001]&m[1025])|(m[998]&m[999]&~m[1000]&m[1001]&m[1025])|(m[998]&~m[999]&m[1000]&m[1001]&m[1025])|(~m[998]&m[999]&m[1000]&m[1001]&m[1025]))&~BiasedRNG[909])|((m[998]&m[999]&~m[1000]&~m[1001]&~m[1025])|(m[998]&~m[999]&m[1000]&~m[1001]&~m[1025])|(~m[998]&m[999]&m[1000]&~m[1001]&~m[1025])|(m[998]&m[999]&m[1000]&~m[1001]&~m[1025])|(m[998]&m[999]&m[1000]&m[1001]&~m[1025])|(m[998]&m[999]&~m[1000]&~m[1001]&m[1025])|(m[998]&~m[999]&m[1000]&~m[1001]&m[1025])|(~m[998]&m[999]&m[1000]&~m[1001]&m[1025])|(m[998]&m[999]&m[1000]&~m[1001]&m[1025])|(m[998]&m[999]&m[1000]&m[1001]&m[1025]));
    m[1007] = (((m[1003]&~m[1004]&~m[1005]&~m[1006]&~m[1035])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1035])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1035])|(m[1003]&m[1004]&~m[1005]&m[1006]&~m[1035])|(m[1003]&~m[1004]&m[1005]&m[1006]&~m[1035])|(~m[1003]&m[1004]&m[1005]&m[1006]&~m[1035]))&BiasedRNG[910])|(((m[1003]&~m[1004]&~m[1005]&~m[1006]&m[1035])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&m[1035])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&m[1035])|(m[1003]&m[1004]&~m[1005]&m[1006]&m[1035])|(m[1003]&~m[1004]&m[1005]&m[1006]&m[1035])|(~m[1003]&m[1004]&m[1005]&m[1006]&m[1035]))&~BiasedRNG[910])|((m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1035])|(m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1035])|(~m[1003]&m[1004]&m[1005]&~m[1006]&~m[1035])|(m[1003]&m[1004]&m[1005]&~m[1006]&~m[1035])|(m[1003]&m[1004]&m[1005]&m[1006]&~m[1035])|(m[1003]&m[1004]&~m[1005]&~m[1006]&m[1035])|(m[1003]&~m[1004]&m[1005]&~m[1006]&m[1035])|(~m[1003]&m[1004]&m[1005]&~m[1006]&m[1035])|(m[1003]&m[1004]&m[1005]&~m[1006]&m[1035])|(m[1003]&m[1004]&m[1005]&m[1006]&m[1035]));
    m[1012] = (((m[1008]&~m[1009]&~m[1010]&~m[1011]&~m[1040])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1040])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1040])|(m[1008]&m[1009]&~m[1010]&m[1011]&~m[1040])|(m[1008]&~m[1009]&m[1010]&m[1011]&~m[1040])|(~m[1008]&m[1009]&m[1010]&m[1011]&~m[1040]))&BiasedRNG[911])|(((m[1008]&~m[1009]&~m[1010]&~m[1011]&m[1040])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&m[1040])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&m[1040])|(m[1008]&m[1009]&~m[1010]&m[1011]&m[1040])|(m[1008]&~m[1009]&m[1010]&m[1011]&m[1040])|(~m[1008]&m[1009]&m[1010]&m[1011]&m[1040]))&~BiasedRNG[911])|((m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1040])|(m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1040])|(~m[1008]&m[1009]&m[1010]&~m[1011]&~m[1040])|(m[1008]&m[1009]&m[1010]&~m[1011]&~m[1040])|(m[1008]&m[1009]&m[1010]&m[1011]&~m[1040])|(m[1008]&m[1009]&~m[1010]&~m[1011]&m[1040])|(m[1008]&~m[1009]&m[1010]&~m[1011]&m[1040])|(~m[1008]&m[1009]&m[1010]&~m[1011]&m[1040])|(m[1008]&m[1009]&m[1010]&~m[1011]&m[1040])|(m[1008]&m[1009]&m[1010]&m[1011]&m[1040]));
    m[1017] = (((m[1013]&~m[1014]&~m[1015]&~m[1016]&~m[1045])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1045])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1045])|(m[1013]&m[1014]&~m[1015]&m[1016]&~m[1045])|(m[1013]&~m[1014]&m[1015]&m[1016]&~m[1045])|(~m[1013]&m[1014]&m[1015]&m[1016]&~m[1045]))&BiasedRNG[912])|(((m[1013]&~m[1014]&~m[1015]&~m[1016]&m[1045])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&m[1045])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&m[1045])|(m[1013]&m[1014]&~m[1015]&m[1016]&m[1045])|(m[1013]&~m[1014]&m[1015]&m[1016]&m[1045])|(~m[1013]&m[1014]&m[1015]&m[1016]&m[1045]))&~BiasedRNG[912])|((m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1045])|(m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1045])|(~m[1013]&m[1014]&m[1015]&~m[1016]&~m[1045])|(m[1013]&m[1014]&m[1015]&~m[1016]&~m[1045])|(m[1013]&m[1014]&m[1015]&m[1016]&~m[1045])|(m[1013]&m[1014]&~m[1015]&~m[1016]&m[1045])|(m[1013]&~m[1014]&m[1015]&~m[1016]&m[1045])|(~m[1013]&m[1014]&m[1015]&~m[1016]&m[1045])|(m[1013]&m[1014]&m[1015]&~m[1016]&m[1045])|(m[1013]&m[1014]&m[1015]&m[1016]&m[1045]));
    m[1022] = (((m[1018]&~m[1019]&~m[1020]&~m[1021]&~m[1050])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1050])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1050])|(m[1018]&m[1019]&~m[1020]&m[1021]&~m[1050])|(m[1018]&~m[1019]&m[1020]&m[1021]&~m[1050])|(~m[1018]&m[1019]&m[1020]&m[1021]&~m[1050]))&BiasedRNG[913])|(((m[1018]&~m[1019]&~m[1020]&~m[1021]&m[1050])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&m[1050])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&m[1050])|(m[1018]&m[1019]&~m[1020]&m[1021]&m[1050])|(m[1018]&~m[1019]&m[1020]&m[1021]&m[1050])|(~m[1018]&m[1019]&m[1020]&m[1021]&m[1050]))&~BiasedRNG[913])|((m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1050])|(m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1050])|(~m[1018]&m[1019]&m[1020]&~m[1021]&~m[1050])|(m[1018]&m[1019]&m[1020]&~m[1021]&~m[1050])|(m[1018]&m[1019]&m[1020]&m[1021]&~m[1050])|(m[1018]&m[1019]&~m[1020]&~m[1021]&m[1050])|(m[1018]&~m[1019]&m[1020]&~m[1021]&m[1050])|(~m[1018]&m[1019]&m[1020]&~m[1021]&m[1050])|(m[1018]&m[1019]&m[1020]&~m[1021]&m[1050])|(m[1018]&m[1019]&m[1020]&m[1021]&m[1050]));
    m[1027] = (((m[1023]&~m[1024]&~m[1025]&~m[1026]&~m[1055])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1055])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1055])|(m[1023]&m[1024]&~m[1025]&m[1026]&~m[1055])|(m[1023]&~m[1024]&m[1025]&m[1026]&~m[1055])|(~m[1023]&m[1024]&m[1025]&m[1026]&~m[1055]))&BiasedRNG[914])|(((m[1023]&~m[1024]&~m[1025]&~m[1026]&m[1055])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&m[1055])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&m[1055])|(m[1023]&m[1024]&~m[1025]&m[1026]&m[1055])|(m[1023]&~m[1024]&m[1025]&m[1026]&m[1055])|(~m[1023]&m[1024]&m[1025]&m[1026]&m[1055]))&~BiasedRNG[914])|((m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1055])|(m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1055])|(~m[1023]&m[1024]&m[1025]&~m[1026]&~m[1055])|(m[1023]&m[1024]&m[1025]&~m[1026]&~m[1055])|(m[1023]&m[1024]&m[1025]&m[1026]&~m[1055])|(m[1023]&m[1024]&~m[1025]&~m[1026]&m[1055])|(m[1023]&~m[1024]&m[1025]&~m[1026]&m[1055])|(~m[1023]&m[1024]&m[1025]&~m[1026]&m[1055])|(m[1023]&m[1024]&m[1025]&~m[1026]&m[1055])|(m[1023]&m[1024]&m[1025]&m[1026]&m[1055]));
    m[1032] = (((m[1028]&~m[1029]&~m[1030]&~m[1031]&~m[1060])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1060])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1060])|(m[1028]&m[1029]&~m[1030]&m[1031]&~m[1060])|(m[1028]&~m[1029]&m[1030]&m[1031]&~m[1060])|(~m[1028]&m[1029]&m[1030]&m[1031]&~m[1060]))&BiasedRNG[915])|(((m[1028]&~m[1029]&~m[1030]&~m[1031]&m[1060])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&m[1060])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&m[1060])|(m[1028]&m[1029]&~m[1030]&m[1031]&m[1060])|(m[1028]&~m[1029]&m[1030]&m[1031]&m[1060])|(~m[1028]&m[1029]&m[1030]&m[1031]&m[1060]))&~BiasedRNG[915])|((m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1060])|(m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1060])|(~m[1028]&m[1029]&m[1030]&~m[1031]&~m[1060])|(m[1028]&m[1029]&m[1030]&~m[1031]&~m[1060])|(m[1028]&m[1029]&m[1030]&m[1031]&~m[1060])|(m[1028]&m[1029]&~m[1030]&~m[1031]&m[1060])|(m[1028]&~m[1029]&m[1030]&~m[1031]&m[1060])|(~m[1028]&m[1029]&m[1030]&~m[1031]&m[1060])|(m[1028]&m[1029]&m[1030]&~m[1031]&m[1060])|(m[1028]&m[1029]&m[1030]&m[1031]&m[1060]));
    m[1037] = (((m[1033]&~m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&~m[1070]))&BiasedRNG[916])|(((m[1033]&~m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&m[1070]))&~BiasedRNG[916])|((m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&m[1070]));
    m[1042] = (((m[1038]&~m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&~m[1075]))&BiasedRNG[917])|(((m[1038]&~m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&m[1075]))&~BiasedRNG[917])|((m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&m[1075]));
    m[1047] = (((m[1043]&~m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&~m[1080]))&BiasedRNG[918])|(((m[1043]&~m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&m[1080]))&~BiasedRNG[918])|((m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&m[1080]));
    m[1052] = (((m[1048]&~m[1049]&~m[1050]&~m[1051]&~m[1085])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1085])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1085])|(m[1048]&m[1049]&~m[1050]&m[1051]&~m[1085])|(m[1048]&~m[1049]&m[1050]&m[1051]&~m[1085])|(~m[1048]&m[1049]&m[1050]&m[1051]&~m[1085]))&BiasedRNG[919])|(((m[1048]&~m[1049]&~m[1050]&~m[1051]&m[1085])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&m[1085])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&m[1085])|(m[1048]&m[1049]&~m[1050]&m[1051]&m[1085])|(m[1048]&~m[1049]&m[1050]&m[1051]&m[1085])|(~m[1048]&m[1049]&m[1050]&m[1051]&m[1085]))&~BiasedRNG[919])|((m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1085])|(m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1085])|(~m[1048]&m[1049]&m[1050]&~m[1051]&~m[1085])|(m[1048]&m[1049]&m[1050]&~m[1051]&~m[1085])|(m[1048]&m[1049]&m[1050]&m[1051]&~m[1085])|(m[1048]&m[1049]&~m[1050]&~m[1051]&m[1085])|(m[1048]&~m[1049]&m[1050]&~m[1051]&m[1085])|(~m[1048]&m[1049]&m[1050]&~m[1051]&m[1085])|(m[1048]&m[1049]&m[1050]&~m[1051]&m[1085])|(m[1048]&m[1049]&m[1050]&m[1051]&m[1085]));
    m[1057] = (((m[1053]&~m[1054]&~m[1055]&~m[1056]&~m[1090])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1090])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1090])|(m[1053]&m[1054]&~m[1055]&m[1056]&~m[1090])|(m[1053]&~m[1054]&m[1055]&m[1056]&~m[1090])|(~m[1053]&m[1054]&m[1055]&m[1056]&~m[1090]))&BiasedRNG[920])|(((m[1053]&~m[1054]&~m[1055]&~m[1056]&m[1090])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&m[1090])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&m[1090])|(m[1053]&m[1054]&~m[1055]&m[1056]&m[1090])|(m[1053]&~m[1054]&m[1055]&m[1056]&m[1090])|(~m[1053]&m[1054]&m[1055]&m[1056]&m[1090]))&~BiasedRNG[920])|((m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1090])|(m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1090])|(~m[1053]&m[1054]&m[1055]&~m[1056]&~m[1090])|(m[1053]&m[1054]&m[1055]&~m[1056]&~m[1090])|(m[1053]&m[1054]&m[1055]&m[1056]&~m[1090])|(m[1053]&m[1054]&~m[1055]&~m[1056]&m[1090])|(m[1053]&~m[1054]&m[1055]&~m[1056]&m[1090])|(~m[1053]&m[1054]&m[1055]&~m[1056]&m[1090])|(m[1053]&m[1054]&m[1055]&~m[1056]&m[1090])|(m[1053]&m[1054]&m[1055]&m[1056]&m[1090]));
    m[1062] = (((m[1058]&~m[1059]&~m[1060]&~m[1061]&~m[1095])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1095])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1095])|(m[1058]&m[1059]&~m[1060]&m[1061]&~m[1095])|(m[1058]&~m[1059]&m[1060]&m[1061]&~m[1095])|(~m[1058]&m[1059]&m[1060]&m[1061]&~m[1095]))&BiasedRNG[921])|(((m[1058]&~m[1059]&~m[1060]&~m[1061]&m[1095])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&m[1095])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&m[1095])|(m[1058]&m[1059]&~m[1060]&m[1061]&m[1095])|(m[1058]&~m[1059]&m[1060]&m[1061]&m[1095])|(~m[1058]&m[1059]&m[1060]&m[1061]&m[1095]))&~BiasedRNG[921])|((m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1095])|(m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1095])|(~m[1058]&m[1059]&m[1060]&~m[1061]&~m[1095])|(m[1058]&m[1059]&m[1060]&~m[1061]&~m[1095])|(m[1058]&m[1059]&m[1060]&m[1061]&~m[1095])|(m[1058]&m[1059]&~m[1060]&~m[1061]&m[1095])|(m[1058]&~m[1059]&m[1060]&~m[1061]&m[1095])|(~m[1058]&m[1059]&m[1060]&~m[1061]&m[1095])|(m[1058]&m[1059]&m[1060]&~m[1061]&m[1095])|(m[1058]&m[1059]&m[1060]&m[1061]&m[1095]));
    m[1067] = (((m[1063]&~m[1064]&~m[1065]&~m[1066]&~m[1100])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1100])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1100])|(m[1063]&m[1064]&~m[1065]&m[1066]&~m[1100])|(m[1063]&~m[1064]&m[1065]&m[1066]&~m[1100])|(~m[1063]&m[1064]&m[1065]&m[1066]&~m[1100]))&BiasedRNG[922])|(((m[1063]&~m[1064]&~m[1065]&~m[1066]&m[1100])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&m[1100])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&m[1100])|(m[1063]&m[1064]&~m[1065]&m[1066]&m[1100])|(m[1063]&~m[1064]&m[1065]&m[1066]&m[1100])|(~m[1063]&m[1064]&m[1065]&m[1066]&m[1100]))&~BiasedRNG[922])|((m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1100])|(m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1100])|(~m[1063]&m[1064]&m[1065]&~m[1066]&~m[1100])|(m[1063]&m[1064]&m[1065]&~m[1066]&~m[1100])|(m[1063]&m[1064]&m[1065]&m[1066]&~m[1100])|(m[1063]&m[1064]&~m[1065]&~m[1066]&m[1100])|(m[1063]&~m[1064]&m[1065]&~m[1066]&m[1100])|(~m[1063]&m[1064]&m[1065]&~m[1066]&m[1100])|(m[1063]&m[1064]&m[1065]&~m[1066]&m[1100])|(m[1063]&m[1064]&m[1065]&m[1066]&m[1100]));
    m[1072] = (((m[1068]&~m[1069]&~m[1070]&~m[1071]&~m[1110])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1110])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1110])|(m[1068]&m[1069]&~m[1070]&m[1071]&~m[1110])|(m[1068]&~m[1069]&m[1070]&m[1071]&~m[1110])|(~m[1068]&m[1069]&m[1070]&m[1071]&~m[1110]))&BiasedRNG[923])|(((m[1068]&~m[1069]&~m[1070]&~m[1071]&m[1110])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&m[1110])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&m[1110])|(m[1068]&m[1069]&~m[1070]&m[1071]&m[1110])|(m[1068]&~m[1069]&m[1070]&m[1071]&m[1110])|(~m[1068]&m[1069]&m[1070]&m[1071]&m[1110]))&~BiasedRNG[923])|((m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1110])|(m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1110])|(~m[1068]&m[1069]&m[1070]&~m[1071]&~m[1110])|(m[1068]&m[1069]&m[1070]&~m[1071]&~m[1110])|(m[1068]&m[1069]&m[1070]&m[1071]&~m[1110])|(m[1068]&m[1069]&~m[1070]&~m[1071]&m[1110])|(m[1068]&~m[1069]&m[1070]&~m[1071]&m[1110])|(~m[1068]&m[1069]&m[1070]&~m[1071]&m[1110])|(m[1068]&m[1069]&m[1070]&~m[1071]&m[1110])|(m[1068]&m[1069]&m[1070]&m[1071]&m[1110]));
    m[1077] = (((m[1073]&~m[1074]&~m[1075]&~m[1076]&~m[1115])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1115])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1115])|(m[1073]&m[1074]&~m[1075]&m[1076]&~m[1115])|(m[1073]&~m[1074]&m[1075]&m[1076]&~m[1115])|(~m[1073]&m[1074]&m[1075]&m[1076]&~m[1115]))&BiasedRNG[924])|(((m[1073]&~m[1074]&~m[1075]&~m[1076]&m[1115])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&m[1115])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&m[1115])|(m[1073]&m[1074]&~m[1075]&m[1076]&m[1115])|(m[1073]&~m[1074]&m[1075]&m[1076]&m[1115])|(~m[1073]&m[1074]&m[1075]&m[1076]&m[1115]))&~BiasedRNG[924])|((m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1115])|(m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1115])|(~m[1073]&m[1074]&m[1075]&~m[1076]&~m[1115])|(m[1073]&m[1074]&m[1075]&~m[1076]&~m[1115])|(m[1073]&m[1074]&m[1075]&m[1076]&~m[1115])|(m[1073]&m[1074]&~m[1075]&~m[1076]&m[1115])|(m[1073]&~m[1074]&m[1075]&~m[1076]&m[1115])|(~m[1073]&m[1074]&m[1075]&~m[1076]&m[1115])|(m[1073]&m[1074]&m[1075]&~m[1076]&m[1115])|(m[1073]&m[1074]&m[1075]&m[1076]&m[1115]));
    m[1082] = (((m[1078]&~m[1079]&~m[1080]&~m[1081]&~m[1120])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1120])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1120])|(m[1078]&m[1079]&~m[1080]&m[1081]&~m[1120])|(m[1078]&~m[1079]&m[1080]&m[1081]&~m[1120])|(~m[1078]&m[1079]&m[1080]&m[1081]&~m[1120]))&BiasedRNG[925])|(((m[1078]&~m[1079]&~m[1080]&~m[1081]&m[1120])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&m[1120])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&m[1120])|(m[1078]&m[1079]&~m[1080]&m[1081]&m[1120])|(m[1078]&~m[1079]&m[1080]&m[1081]&m[1120])|(~m[1078]&m[1079]&m[1080]&m[1081]&m[1120]))&~BiasedRNG[925])|((m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1120])|(m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1120])|(~m[1078]&m[1079]&m[1080]&~m[1081]&~m[1120])|(m[1078]&m[1079]&m[1080]&~m[1081]&~m[1120])|(m[1078]&m[1079]&m[1080]&m[1081]&~m[1120])|(m[1078]&m[1079]&~m[1080]&~m[1081]&m[1120])|(m[1078]&~m[1079]&m[1080]&~m[1081]&m[1120])|(~m[1078]&m[1079]&m[1080]&~m[1081]&m[1120])|(m[1078]&m[1079]&m[1080]&~m[1081]&m[1120])|(m[1078]&m[1079]&m[1080]&m[1081]&m[1120]));
    m[1087] = (((m[1083]&~m[1084]&~m[1085]&~m[1086]&~m[1125])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1125])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1125])|(m[1083]&m[1084]&~m[1085]&m[1086]&~m[1125])|(m[1083]&~m[1084]&m[1085]&m[1086]&~m[1125])|(~m[1083]&m[1084]&m[1085]&m[1086]&~m[1125]))&BiasedRNG[926])|(((m[1083]&~m[1084]&~m[1085]&~m[1086]&m[1125])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&m[1125])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&m[1125])|(m[1083]&m[1084]&~m[1085]&m[1086]&m[1125])|(m[1083]&~m[1084]&m[1085]&m[1086]&m[1125])|(~m[1083]&m[1084]&m[1085]&m[1086]&m[1125]))&~BiasedRNG[926])|((m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1125])|(m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1125])|(~m[1083]&m[1084]&m[1085]&~m[1086]&~m[1125])|(m[1083]&m[1084]&m[1085]&~m[1086]&~m[1125])|(m[1083]&m[1084]&m[1085]&m[1086]&~m[1125])|(m[1083]&m[1084]&~m[1085]&~m[1086]&m[1125])|(m[1083]&~m[1084]&m[1085]&~m[1086]&m[1125])|(~m[1083]&m[1084]&m[1085]&~m[1086]&m[1125])|(m[1083]&m[1084]&m[1085]&~m[1086]&m[1125])|(m[1083]&m[1084]&m[1085]&m[1086]&m[1125]));
    m[1092] = (((m[1088]&~m[1089]&~m[1090]&~m[1091]&~m[1130])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1130])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1130])|(m[1088]&m[1089]&~m[1090]&m[1091]&~m[1130])|(m[1088]&~m[1089]&m[1090]&m[1091]&~m[1130])|(~m[1088]&m[1089]&m[1090]&m[1091]&~m[1130]))&BiasedRNG[927])|(((m[1088]&~m[1089]&~m[1090]&~m[1091]&m[1130])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&m[1130])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&m[1130])|(m[1088]&m[1089]&~m[1090]&m[1091]&m[1130])|(m[1088]&~m[1089]&m[1090]&m[1091]&m[1130])|(~m[1088]&m[1089]&m[1090]&m[1091]&m[1130]))&~BiasedRNG[927])|((m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1130])|(m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1130])|(~m[1088]&m[1089]&m[1090]&~m[1091]&~m[1130])|(m[1088]&m[1089]&m[1090]&~m[1091]&~m[1130])|(m[1088]&m[1089]&m[1090]&m[1091]&~m[1130])|(m[1088]&m[1089]&~m[1090]&~m[1091]&m[1130])|(m[1088]&~m[1089]&m[1090]&~m[1091]&m[1130])|(~m[1088]&m[1089]&m[1090]&~m[1091]&m[1130])|(m[1088]&m[1089]&m[1090]&~m[1091]&m[1130])|(m[1088]&m[1089]&m[1090]&m[1091]&m[1130]));
    m[1097] = (((m[1093]&~m[1094]&~m[1095]&~m[1096]&~m[1135])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1135])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1135])|(m[1093]&m[1094]&~m[1095]&m[1096]&~m[1135])|(m[1093]&~m[1094]&m[1095]&m[1096]&~m[1135])|(~m[1093]&m[1094]&m[1095]&m[1096]&~m[1135]))&BiasedRNG[928])|(((m[1093]&~m[1094]&~m[1095]&~m[1096]&m[1135])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&m[1135])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&m[1135])|(m[1093]&m[1094]&~m[1095]&m[1096]&m[1135])|(m[1093]&~m[1094]&m[1095]&m[1096]&m[1135])|(~m[1093]&m[1094]&m[1095]&m[1096]&m[1135]))&~BiasedRNG[928])|((m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1135])|(m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1135])|(~m[1093]&m[1094]&m[1095]&~m[1096]&~m[1135])|(m[1093]&m[1094]&m[1095]&~m[1096]&~m[1135])|(m[1093]&m[1094]&m[1095]&m[1096]&~m[1135])|(m[1093]&m[1094]&~m[1095]&~m[1096]&m[1135])|(m[1093]&~m[1094]&m[1095]&~m[1096]&m[1135])|(~m[1093]&m[1094]&m[1095]&~m[1096]&m[1135])|(m[1093]&m[1094]&m[1095]&~m[1096]&m[1135])|(m[1093]&m[1094]&m[1095]&m[1096]&m[1135]));
    m[1102] = (((m[1098]&~m[1099]&~m[1100]&~m[1101]&~m[1140])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1140])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1140])|(m[1098]&m[1099]&~m[1100]&m[1101]&~m[1140])|(m[1098]&~m[1099]&m[1100]&m[1101]&~m[1140])|(~m[1098]&m[1099]&m[1100]&m[1101]&~m[1140]))&BiasedRNG[929])|(((m[1098]&~m[1099]&~m[1100]&~m[1101]&m[1140])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&m[1140])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&m[1140])|(m[1098]&m[1099]&~m[1100]&m[1101]&m[1140])|(m[1098]&~m[1099]&m[1100]&m[1101]&m[1140])|(~m[1098]&m[1099]&m[1100]&m[1101]&m[1140]))&~BiasedRNG[929])|((m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1140])|(m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1140])|(~m[1098]&m[1099]&m[1100]&~m[1101]&~m[1140])|(m[1098]&m[1099]&m[1100]&~m[1101]&~m[1140])|(m[1098]&m[1099]&m[1100]&m[1101]&~m[1140])|(m[1098]&m[1099]&~m[1100]&~m[1101]&m[1140])|(m[1098]&~m[1099]&m[1100]&~m[1101]&m[1140])|(~m[1098]&m[1099]&m[1100]&~m[1101]&m[1140])|(m[1098]&m[1099]&m[1100]&~m[1101]&m[1140])|(m[1098]&m[1099]&m[1100]&m[1101]&m[1140]));
    m[1107] = (((m[1103]&~m[1104]&~m[1105]&~m[1106]&~m[1145])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1145])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1145])|(m[1103]&m[1104]&~m[1105]&m[1106]&~m[1145])|(m[1103]&~m[1104]&m[1105]&m[1106]&~m[1145])|(~m[1103]&m[1104]&m[1105]&m[1106]&~m[1145]))&BiasedRNG[930])|(((m[1103]&~m[1104]&~m[1105]&~m[1106]&m[1145])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&m[1145])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&m[1145])|(m[1103]&m[1104]&~m[1105]&m[1106]&m[1145])|(m[1103]&~m[1104]&m[1105]&m[1106]&m[1145])|(~m[1103]&m[1104]&m[1105]&m[1106]&m[1145]))&~BiasedRNG[930])|((m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1145])|(m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1145])|(~m[1103]&m[1104]&m[1105]&~m[1106]&~m[1145])|(m[1103]&m[1104]&m[1105]&~m[1106]&~m[1145])|(m[1103]&m[1104]&m[1105]&m[1106]&~m[1145])|(m[1103]&m[1104]&~m[1105]&~m[1106]&m[1145])|(m[1103]&~m[1104]&m[1105]&~m[1106]&m[1145])|(~m[1103]&m[1104]&m[1105]&~m[1106]&m[1145])|(m[1103]&m[1104]&m[1105]&~m[1106]&m[1145])|(m[1103]&m[1104]&m[1105]&m[1106]&m[1145]));
    m[1112] = (((m[1108]&~m[1109]&~m[1110]&~m[1111]&~m[1155])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1155])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1155])|(m[1108]&m[1109]&~m[1110]&m[1111]&~m[1155])|(m[1108]&~m[1109]&m[1110]&m[1111]&~m[1155])|(~m[1108]&m[1109]&m[1110]&m[1111]&~m[1155]))&BiasedRNG[931])|(((m[1108]&~m[1109]&~m[1110]&~m[1111]&m[1155])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&m[1155])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&m[1155])|(m[1108]&m[1109]&~m[1110]&m[1111]&m[1155])|(m[1108]&~m[1109]&m[1110]&m[1111]&m[1155])|(~m[1108]&m[1109]&m[1110]&m[1111]&m[1155]))&~BiasedRNG[931])|((m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1155])|(m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1155])|(~m[1108]&m[1109]&m[1110]&~m[1111]&~m[1155])|(m[1108]&m[1109]&m[1110]&~m[1111]&~m[1155])|(m[1108]&m[1109]&m[1110]&m[1111]&~m[1155])|(m[1108]&m[1109]&~m[1110]&~m[1111]&m[1155])|(m[1108]&~m[1109]&m[1110]&~m[1111]&m[1155])|(~m[1108]&m[1109]&m[1110]&~m[1111]&m[1155])|(m[1108]&m[1109]&m[1110]&~m[1111]&m[1155])|(m[1108]&m[1109]&m[1110]&m[1111]&m[1155]));
    m[1117] = (((m[1113]&~m[1114]&~m[1115]&~m[1116]&~m[1160])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1160])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1160])|(m[1113]&m[1114]&~m[1115]&m[1116]&~m[1160])|(m[1113]&~m[1114]&m[1115]&m[1116]&~m[1160])|(~m[1113]&m[1114]&m[1115]&m[1116]&~m[1160]))&BiasedRNG[932])|(((m[1113]&~m[1114]&~m[1115]&~m[1116]&m[1160])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&m[1160])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&m[1160])|(m[1113]&m[1114]&~m[1115]&m[1116]&m[1160])|(m[1113]&~m[1114]&m[1115]&m[1116]&m[1160])|(~m[1113]&m[1114]&m[1115]&m[1116]&m[1160]))&~BiasedRNG[932])|((m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1160])|(m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1160])|(~m[1113]&m[1114]&m[1115]&~m[1116]&~m[1160])|(m[1113]&m[1114]&m[1115]&~m[1116]&~m[1160])|(m[1113]&m[1114]&m[1115]&m[1116]&~m[1160])|(m[1113]&m[1114]&~m[1115]&~m[1116]&m[1160])|(m[1113]&~m[1114]&m[1115]&~m[1116]&m[1160])|(~m[1113]&m[1114]&m[1115]&~m[1116]&m[1160])|(m[1113]&m[1114]&m[1115]&~m[1116]&m[1160])|(m[1113]&m[1114]&m[1115]&m[1116]&m[1160]));
    m[1122] = (((m[1118]&~m[1119]&~m[1120]&~m[1121]&~m[1165])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1165])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1165])|(m[1118]&m[1119]&~m[1120]&m[1121]&~m[1165])|(m[1118]&~m[1119]&m[1120]&m[1121]&~m[1165])|(~m[1118]&m[1119]&m[1120]&m[1121]&~m[1165]))&BiasedRNG[933])|(((m[1118]&~m[1119]&~m[1120]&~m[1121]&m[1165])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&m[1165])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&m[1165])|(m[1118]&m[1119]&~m[1120]&m[1121]&m[1165])|(m[1118]&~m[1119]&m[1120]&m[1121]&m[1165])|(~m[1118]&m[1119]&m[1120]&m[1121]&m[1165]))&~BiasedRNG[933])|((m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1165])|(m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1165])|(~m[1118]&m[1119]&m[1120]&~m[1121]&~m[1165])|(m[1118]&m[1119]&m[1120]&~m[1121]&~m[1165])|(m[1118]&m[1119]&m[1120]&m[1121]&~m[1165])|(m[1118]&m[1119]&~m[1120]&~m[1121]&m[1165])|(m[1118]&~m[1119]&m[1120]&~m[1121]&m[1165])|(~m[1118]&m[1119]&m[1120]&~m[1121]&m[1165])|(m[1118]&m[1119]&m[1120]&~m[1121]&m[1165])|(m[1118]&m[1119]&m[1120]&m[1121]&m[1165]));
    m[1127] = (((m[1123]&~m[1124]&~m[1125]&~m[1126]&~m[1170])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1170])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1170])|(m[1123]&m[1124]&~m[1125]&m[1126]&~m[1170])|(m[1123]&~m[1124]&m[1125]&m[1126]&~m[1170])|(~m[1123]&m[1124]&m[1125]&m[1126]&~m[1170]))&BiasedRNG[934])|(((m[1123]&~m[1124]&~m[1125]&~m[1126]&m[1170])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&m[1170])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&m[1170])|(m[1123]&m[1124]&~m[1125]&m[1126]&m[1170])|(m[1123]&~m[1124]&m[1125]&m[1126]&m[1170])|(~m[1123]&m[1124]&m[1125]&m[1126]&m[1170]))&~BiasedRNG[934])|((m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1170])|(m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1170])|(~m[1123]&m[1124]&m[1125]&~m[1126]&~m[1170])|(m[1123]&m[1124]&m[1125]&~m[1126]&~m[1170])|(m[1123]&m[1124]&m[1125]&m[1126]&~m[1170])|(m[1123]&m[1124]&~m[1125]&~m[1126]&m[1170])|(m[1123]&~m[1124]&m[1125]&~m[1126]&m[1170])|(~m[1123]&m[1124]&m[1125]&~m[1126]&m[1170])|(m[1123]&m[1124]&m[1125]&~m[1126]&m[1170])|(m[1123]&m[1124]&m[1125]&m[1126]&m[1170]));
    m[1132] = (((m[1128]&~m[1129]&~m[1130]&~m[1131]&~m[1175])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1175])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1175])|(m[1128]&m[1129]&~m[1130]&m[1131]&~m[1175])|(m[1128]&~m[1129]&m[1130]&m[1131]&~m[1175])|(~m[1128]&m[1129]&m[1130]&m[1131]&~m[1175]))&BiasedRNG[935])|(((m[1128]&~m[1129]&~m[1130]&~m[1131]&m[1175])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&m[1175])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&m[1175])|(m[1128]&m[1129]&~m[1130]&m[1131]&m[1175])|(m[1128]&~m[1129]&m[1130]&m[1131]&m[1175])|(~m[1128]&m[1129]&m[1130]&m[1131]&m[1175]))&~BiasedRNG[935])|((m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1175])|(m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1175])|(~m[1128]&m[1129]&m[1130]&~m[1131]&~m[1175])|(m[1128]&m[1129]&m[1130]&~m[1131]&~m[1175])|(m[1128]&m[1129]&m[1130]&m[1131]&~m[1175])|(m[1128]&m[1129]&~m[1130]&~m[1131]&m[1175])|(m[1128]&~m[1129]&m[1130]&~m[1131]&m[1175])|(~m[1128]&m[1129]&m[1130]&~m[1131]&m[1175])|(m[1128]&m[1129]&m[1130]&~m[1131]&m[1175])|(m[1128]&m[1129]&m[1130]&m[1131]&m[1175]));
    m[1137] = (((m[1133]&~m[1134]&~m[1135]&~m[1136]&~m[1180])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1180])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1180])|(m[1133]&m[1134]&~m[1135]&m[1136]&~m[1180])|(m[1133]&~m[1134]&m[1135]&m[1136]&~m[1180])|(~m[1133]&m[1134]&m[1135]&m[1136]&~m[1180]))&BiasedRNG[936])|(((m[1133]&~m[1134]&~m[1135]&~m[1136]&m[1180])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&m[1180])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&m[1180])|(m[1133]&m[1134]&~m[1135]&m[1136]&m[1180])|(m[1133]&~m[1134]&m[1135]&m[1136]&m[1180])|(~m[1133]&m[1134]&m[1135]&m[1136]&m[1180]))&~BiasedRNG[936])|((m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1180])|(m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1180])|(~m[1133]&m[1134]&m[1135]&~m[1136]&~m[1180])|(m[1133]&m[1134]&m[1135]&~m[1136]&~m[1180])|(m[1133]&m[1134]&m[1135]&m[1136]&~m[1180])|(m[1133]&m[1134]&~m[1135]&~m[1136]&m[1180])|(m[1133]&~m[1134]&m[1135]&~m[1136]&m[1180])|(~m[1133]&m[1134]&m[1135]&~m[1136]&m[1180])|(m[1133]&m[1134]&m[1135]&~m[1136]&m[1180])|(m[1133]&m[1134]&m[1135]&m[1136]&m[1180]));
    m[1142] = (((m[1138]&~m[1139]&~m[1140]&~m[1141]&~m[1185])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1185])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1185])|(m[1138]&m[1139]&~m[1140]&m[1141]&~m[1185])|(m[1138]&~m[1139]&m[1140]&m[1141]&~m[1185])|(~m[1138]&m[1139]&m[1140]&m[1141]&~m[1185]))&BiasedRNG[937])|(((m[1138]&~m[1139]&~m[1140]&~m[1141]&m[1185])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&m[1185])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&m[1185])|(m[1138]&m[1139]&~m[1140]&m[1141]&m[1185])|(m[1138]&~m[1139]&m[1140]&m[1141]&m[1185])|(~m[1138]&m[1139]&m[1140]&m[1141]&m[1185]))&~BiasedRNG[937])|((m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1185])|(m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1185])|(~m[1138]&m[1139]&m[1140]&~m[1141]&~m[1185])|(m[1138]&m[1139]&m[1140]&~m[1141]&~m[1185])|(m[1138]&m[1139]&m[1140]&m[1141]&~m[1185])|(m[1138]&m[1139]&~m[1140]&~m[1141]&m[1185])|(m[1138]&~m[1139]&m[1140]&~m[1141]&m[1185])|(~m[1138]&m[1139]&m[1140]&~m[1141]&m[1185])|(m[1138]&m[1139]&m[1140]&~m[1141]&m[1185])|(m[1138]&m[1139]&m[1140]&m[1141]&m[1185]));
    m[1147] = (((m[1143]&~m[1144]&~m[1145]&~m[1146]&~m[1190])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1190])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1190])|(m[1143]&m[1144]&~m[1145]&m[1146]&~m[1190])|(m[1143]&~m[1144]&m[1145]&m[1146]&~m[1190])|(~m[1143]&m[1144]&m[1145]&m[1146]&~m[1190]))&BiasedRNG[938])|(((m[1143]&~m[1144]&~m[1145]&~m[1146]&m[1190])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&m[1190])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&m[1190])|(m[1143]&m[1144]&~m[1145]&m[1146]&m[1190])|(m[1143]&~m[1144]&m[1145]&m[1146]&m[1190])|(~m[1143]&m[1144]&m[1145]&m[1146]&m[1190]))&~BiasedRNG[938])|((m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1190])|(m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1190])|(~m[1143]&m[1144]&m[1145]&~m[1146]&~m[1190])|(m[1143]&m[1144]&m[1145]&~m[1146]&~m[1190])|(m[1143]&m[1144]&m[1145]&m[1146]&~m[1190])|(m[1143]&m[1144]&~m[1145]&~m[1146]&m[1190])|(m[1143]&~m[1144]&m[1145]&~m[1146]&m[1190])|(~m[1143]&m[1144]&m[1145]&~m[1146]&m[1190])|(m[1143]&m[1144]&m[1145]&~m[1146]&m[1190])|(m[1143]&m[1144]&m[1145]&m[1146]&m[1190]));
    m[1152] = (((m[1148]&~m[1149]&~m[1150]&~m[1151]&~m[1195])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1195])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1195])|(m[1148]&m[1149]&~m[1150]&m[1151]&~m[1195])|(m[1148]&~m[1149]&m[1150]&m[1151]&~m[1195])|(~m[1148]&m[1149]&m[1150]&m[1151]&~m[1195]))&BiasedRNG[939])|(((m[1148]&~m[1149]&~m[1150]&~m[1151]&m[1195])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&m[1195])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&m[1195])|(m[1148]&m[1149]&~m[1150]&m[1151]&m[1195])|(m[1148]&~m[1149]&m[1150]&m[1151]&m[1195])|(~m[1148]&m[1149]&m[1150]&m[1151]&m[1195]))&~BiasedRNG[939])|((m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1195])|(m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1195])|(~m[1148]&m[1149]&m[1150]&~m[1151]&~m[1195])|(m[1148]&m[1149]&m[1150]&~m[1151]&~m[1195])|(m[1148]&m[1149]&m[1150]&m[1151]&~m[1195])|(m[1148]&m[1149]&~m[1150]&~m[1151]&m[1195])|(m[1148]&~m[1149]&m[1150]&~m[1151]&m[1195])|(~m[1148]&m[1149]&m[1150]&~m[1151]&m[1195])|(m[1148]&m[1149]&m[1150]&~m[1151]&m[1195])|(m[1148]&m[1149]&m[1150]&m[1151]&m[1195]));
    m[1157] = (((m[1153]&~m[1154]&~m[1155]&~m[1156]&~m[1205])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1205])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1205])|(m[1153]&m[1154]&~m[1155]&m[1156]&~m[1205])|(m[1153]&~m[1154]&m[1155]&m[1156]&~m[1205])|(~m[1153]&m[1154]&m[1155]&m[1156]&~m[1205]))&BiasedRNG[940])|(((m[1153]&~m[1154]&~m[1155]&~m[1156]&m[1205])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&m[1205])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&m[1205])|(m[1153]&m[1154]&~m[1155]&m[1156]&m[1205])|(m[1153]&~m[1154]&m[1155]&m[1156]&m[1205])|(~m[1153]&m[1154]&m[1155]&m[1156]&m[1205]))&~BiasedRNG[940])|((m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1205])|(m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1205])|(~m[1153]&m[1154]&m[1155]&~m[1156]&~m[1205])|(m[1153]&m[1154]&m[1155]&~m[1156]&~m[1205])|(m[1153]&m[1154]&m[1155]&m[1156]&~m[1205])|(m[1153]&m[1154]&~m[1155]&~m[1156]&m[1205])|(m[1153]&~m[1154]&m[1155]&~m[1156]&m[1205])|(~m[1153]&m[1154]&m[1155]&~m[1156]&m[1205])|(m[1153]&m[1154]&m[1155]&~m[1156]&m[1205])|(m[1153]&m[1154]&m[1155]&m[1156]&m[1205]));
    m[1162] = (((m[1158]&~m[1159]&~m[1160]&~m[1161]&~m[1210])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1210])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1210])|(m[1158]&m[1159]&~m[1160]&m[1161]&~m[1210])|(m[1158]&~m[1159]&m[1160]&m[1161]&~m[1210])|(~m[1158]&m[1159]&m[1160]&m[1161]&~m[1210]))&BiasedRNG[941])|(((m[1158]&~m[1159]&~m[1160]&~m[1161]&m[1210])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&m[1210])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&m[1210])|(m[1158]&m[1159]&~m[1160]&m[1161]&m[1210])|(m[1158]&~m[1159]&m[1160]&m[1161]&m[1210])|(~m[1158]&m[1159]&m[1160]&m[1161]&m[1210]))&~BiasedRNG[941])|((m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1210])|(m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1210])|(~m[1158]&m[1159]&m[1160]&~m[1161]&~m[1210])|(m[1158]&m[1159]&m[1160]&~m[1161]&~m[1210])|(m[1158]&m[1159]&m[1160]&m[1161]&~m[1210])|(m[1158]&m[1159]&~m[1160]&~m[1161]&m[1210])|(m[1158]&~m[1159]&m[1160]&~m[1161]&m[1210])|(~m[1158]&m[1159]&m[1160]&~m[1161]&m[1210])|(m[1158]&m[1159]&m[1160]&~m[1161]&m[1210])|(m[1158]&m[1159]&m[1160]&m[1161]&m[1210]));
    m[1167] = (((m[1163]&~m[1164]&~m[1165]&~m[1166]&~m[1215])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1215])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1215])|(m[1163]&m[1164]&~m[1165]&m[1166]&~m[1215])|(m[1163]&~m[1164]&m[1165]&m[1166]&~m[1215])|(~m[1163]&m[1164]&m[1165]&m[1166]&~m[1215]))&BiasedRNG[942])|(((m[1163]&~m[1164]&~m[1165]&~m[1166]&m[1215])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&m[1215])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&m[1215])|(m[1163]&m[1164]&~m[1165]&m[1166]&m[1215])|(m[1163]&~m[1164]&m[1165]&m[1166]&m[1215])|(~m[1163]&m[1164]&m[1165]&m[1166]&m[1215]))&~BiasedRNG[942])|((m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1215])|(m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1215])|(~m[1163]&m[1164]&m[1165]&~m[1166]&~m[1215])|(m[1163]&m[1164]&m[1165]&~m[1166]&~m[1215])|(m[1163]&m[1164]&m[1165]&m[1166]&~m[1215])|(m[1163]&m[1164]&~m[1165]&~m[1166]&m[1215])|(m[1163]&~m[1164]&m[1165]&~m[1166]&m[1215])|(~m[1163]&m[1164]&m[1165]&~m[1166]&m[1215])|(m[1163]&m[1164]&m[1165]&~m[1166]&m[1215])|(m[1163]&m[1164]&m[1165]&m[1166]&m[1215]));
    m[1172] = (((m[1168]&~m[1169]&~m[1170]&~m[1171]&~m[1220])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1220])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1220])|(m[1168]&m[1169]&~m[1170]&m[1171]&~m[1220])|(m[1168]&~m[1169]&m[1170]&m[1171]&~m[1220])|(~m[1168]&m[1169]&m[1170]&m[1171]&~m[1220]))&BiasedRNG[943])|(((m[1168]&~m[1169]&~m[1170]&~m[1171]&m[1220])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&m[1220])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&m[1220])|(m[1168]&m[1169]&~m[1170]&m[1171]&m[1220])|(m[1168]&~m[1169]&m[1170]&m[1171]&m[1220])|(~m[1168]&m[1169]&m[1170]&m[1171]&m[1220]))&~BiasedRNG[943])|((m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1220])|(m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1220])|(~m[1168]&m[1169]&m[1170]&~m[1171]&~m[1220])|(m[1168]&m[1169]&m[1170]&~m[1171]&~m[1220])|(m[1168]&m[1169]&m[1170]&m[1171]&~m[1220])|(m[1168]&m[1169]&~m[1170]&~m[1171]&m[1220])|(m[1168]&~m[1169]&m[1170]&~m[1171]&m[1220])|(~m[1168]&m[1169]&m[1170]&~m[1171]&m[1220])|(m[1168]&m[1169]&m[1170]&~m[1171]&m[1220])|(m[1168]&m[1169]&m[1170]&m[1171]&m[1220]));
    m[1177] = (((m[1173]&~m[1174]&~m[1175]&~m[1176]&~m[1225])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1225])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1225])|(m[1173]&m[1174]&~m[1175]&m[1176]&~m[1225])|(m[1173]&~m[1174]&m[1175]&m[1176]&~m[1225])|(~m[1173]&m[1174]&m[1175]&m[1176]&~m[1225]))&BiasedRNG[944])|(((m[1173]&~m[1174]&~m[1175]&~m[1176]&m[1225])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&m[1225])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&m[1225])|(m[1173]&m[1174]&~m[1175]&m[1176]&m[1225])|(m[1173]&~m[1174]&m[1175]&m[1176]&m[1225])|(~m[1173]&m[1174]&m[1175]&m[1176]&m[1225]))&~BiasedRNG[944])|((m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1225])|(m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1225])|(~m[1173]&m[1174]&m[1175]&~m[1176]&~m[1225])|(m[1173]&m[1174]&m[1175]&~m[1176]&~m[1225])|(m[1173]&m[1174]&m[1175]&m[1176]&~m[1225])|(m[1173]&m[1174]&~m[1175]&~m[1176]&m[1225])|(m[1173]&~m[1174]&m[1175]&~m[1176]&m[1225])|(~m[1173]&m[1174]&m[1175]&~m[1176]&m[1225])|(m[1173]&m[1174]&m[1175]&~m[1176]&m[1225])|(m[1173]&m[1174]&m[1175]&m[1176]&m[1225]));
    m[1182] = (((m[1178]&~m[1179]&~m[1180]&~m[1181]&~m[1230])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1230])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1230])|(m[1178]&m[1179]&~m[1180]&m[1181]&~m[1230])|(m[1178]&~m[1179]&m[1180]&m[1181]&~m[1230])|(~m[1178]&m[1179]&m[1180]&m[1181]&~m[1230]))&BiasedRNG[945])|(((m[1178]&~m[1179]&~m[1180]&~m[1181]&m[1230])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&m[1230])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&m[1230])|(m[1178]&m[1179]&~m[1180]&m[1181]&m[1230])|(m[1178]&~m[1179]&m[1180]&m[1181]&m[1230])|(~m[1178]&m[1179]&m[1180]&m[1181]&m[1230]))&~BiasedRNG[945])|((m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1230])|(m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1230])|(~m[1178]&m[1179]&m[1180]&~m[1181]&~m[1230])|(m[1178]&m[1179]&m[1180]&~m[1181]&~m[1230])|(m[1178]&m[1179]&m[1180]&m[1181]&~m[1230])|(m[1178]&m[1179]&~m[1180]&~m[1181]&m[1230])|(m[1178]&~m[1179]&m[1180]&~m[1181]&m[1230])|(~m[1178]&m[1179]&m[1180]&~m[1181]&m[1230])|(m[1178]&m[1179]&m[1180]&~m[1181]&m[1230])|(m[1178]&m[1179]&m[1180]&m[1181]&m[1230]));
    m[1187] = (((m[1183]&~m[1184]&~m[1185]&~m[1186]&~m[1235])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1235])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1235])|(m[1183]&m[1184]&~m[1185]&m[1186]&~m[1235])|(m[1183]&~m[1184]&m[1185]&m[1186]&~m[1235])|(~m[1183]&m[1184]&m[1185]&m[1186]&~m[1235]))&BiasedRNG[946])|(((m[1183]&~m[1184]&~m[1185]&~m[1186]&m[1235])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&m[1235])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&m[1235])|(m[1183]&m[1184]&~m[1185]&m[1186]&m[1235])|(m[1183]&~m[1184]&m[1185]&m[1186]&m[1235])|(~m[1183]&m[1184]&m[1185]&m[1186]&m[1235]))&~BiasedRNG[946])|((m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1235])|(m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1235])|(~m[1183]&m[1184]&m[1185]&~m[1186]&~m[1235])|(m[1183]&m[1184]&m[1185]&~m[1186]&~m[1235])|(m[1183]&m[1184]&m[1185]&m[1186]&~m[1235])|(m[1183]&m[1184]&~m[1185]&~m[1186]&m[1235])|(m[1183]&~m[1184]&m[1185]&~m[1186]&m[1235])|(~m[1183]&m[1184]&m[1185]&~m[1186]&m[1235])|(m[1183]&m[1184]&m[1185]&~m[1186]&m[1235])|(m[1183]&m[1184]&m[1185]&m[1186]&m[1235]));
    m[1192] = (((m[1188]&~m[1189]&~m[1190]&~m[1191]&~m[1240])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1240])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1240])|(m[1188]&m[1189]&~m[1190]&m[1191]&~m[1240])|(m[1188]&~m[1189]&m[1190]&m[1191]&~m[1240])|(~m[1188]&m[1189]&m[1190]&m[1191]&~m[1240]))&BiasedRNG[947])|(((m[1188]&~m[1189]&~m[1190]&~m[1191]&m[1240])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&m[1240])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&m[1240])|(m[1188]&m[1189]&~m[1190]&m[1191]&m[1240])|(m[1188]&~m[1189]&m[1190]&m[1191]&m[1240])|(~m[1188]&m[1189]&m[1190]&m[1191]&m[1240]))&~BiasedRNG[947])|((m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1240])|(m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1240])|(~m[1188]&m[1189]&m[1190]&~m[1191]&~m[1240])|(m[1188]&m[1189]&m[1190]&~m[1191]&~m[1240])|(m[1188]&m[1189]&m[1190]&m[1191]&~m[1240])|(m[1188]&m[1189]&~m[1190]&~m[1191]&m[1240])|(m[1188]&~m[1189]&m[1190]&~m[1191]&m[1240])|(~m[1188]&m[1189]&m[1190]&~m[1191]&m[1240])|(m[1188]&m[1189]&m[1190]&~m[1191]&m[1240])|(m[1188]&m[1189]&m[1190]&m[1191]&m[1240]));
    m[1197] = (((m[1193]&~m[1194]&~m[1195]&~m[1196]&~m[1245])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1245])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1245])|(m[1193]&m[1194]&~m[1195]&m[1196]&~m[1245])|(m[1193]&~m[1194]&m[1195]&m[1196]&~m[1245])|(~m[1193]&m[1194]&m[1195]&m[1196]&~m[1245]))&BiasedRNG[948])|(((m[1193]&~m[1194]&~m[1195]&~m[1196]&m[1245])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&m[1245])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&m[1245])|(m[1193]&m[1194]&~m[1195]&m[1196]&m[1245])|(m[1193]&~m[1194]&m[1195]&m[1196]&m[1245])|(~m[1193]&m[1194]&m[1195]&m[1196]&m[1245]))&~BiasedRNG[948])|((m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1245])|(m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1245])|(~m[1193]&m[1194]&m[1195]&~m[1196]&~m[1245])|(m[1193]&m[1194]&m[1195]&~m[1196]&~m[1245])|(m[1193]&m[1194]&m[1195]&m[1196]&~m[1245])|(m[1193]&m[1194]&~m[1195]&~m[1196]&m[1245])|(m[1193]&~m[1194]&m[1195]&~m[1196]&m[1245])|(~m[1193]&m[1194]&m[1195]&~m[1196]&m[1245])|(m[1193]&m[1194]&m[1195]&~m[1196]&m[1245])|(m[1193]&m[1194]&m[1195]&m[1196]&m[1245]));
    m[1202] = (((m[1198]&~m[1199]&~m[1200]&~m[1201]&~m[1250])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1250])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1250])|(m[1198]&m[1199]&~m[1200]&m[1201]&~m[1250])|(m[1198]&~m[1199]&m[1200]&m[1201]&~m[1250])|(~m[1198]&m[1199]&m[1200]&m[1201]&~m[1250]))&BiasedRNG[949])|(((m[1198]&~m[1199]&~m[1200]&~m[1201]&m[1250])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&m[1250])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&m[1250])|(m[1198]&m[1199]&~m[1200]&m[1201]&m[1250])|(m[1198]&~m[1199]&m[1200]&m[1201]&m[1250])|(~m[1198]&m[1199]&m[1200]&m[1201]&m[1250]))&~BiasedRNG[949])|((m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1250])|(m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1250])|(~m[1198]&m[1199]&m[1200]&~m[1201]&~m[1250])|(m[1198]&m[1199]&m[1200]&~m[1201]&~m[1250])|(m[1198]&m[1199]&m[1200]&m[1201]&~m[1250])|(m[1198]&m[1199]&~m[1200]&~m[1201]&m[1250])|(m[1198]&~m[1199]&m[1200]&~m[1201]&m[1250])|(~m[1198]&m[1199]&m[1200]&~m[1201]&m[1250])|(m[1198]&m[1199]&m[1200]&~m[1201]&m[1250])|(m[1198]&m[1199]&m[1200]&m[1201]&m[1250]));
    m[1207] = (((m[1203]&~m[1204]&~m[1205]&~m[1206]&~m[1260])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1260])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1260])|(m[1203]&m[1204]&~m[1205]&m[1206]&~m[1260])|(m[1203]&~m[1204]&m[1205]&m[1206]&~m[1260])|(~m[1203]&m[1204]&m[1205]&m[1206]&~m[1260]))&BiasedRNG[950])|(((m[1203]&~m[1204]&~m[1205]&~m[1206]&m[1260])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&m[1260])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&m[1260])|(m[1203]&m[1204]&~m[1205]&m[1206]&m[1260])|(m[1203]&~m[1204]&m[1205]&m[1206]&m[1260])|(~m[1203]&m[1204]&m[1205]&m[1206]&m[1260]))&~BiasedRNG[950])|((m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1260])|(m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1260])|(~m[1203]&m[1204]&m[1205]&~m[1206]&~m[1260])|(m[1203]&m[1204]&m[1205]&~m[1206]&~m[1260])|(m[1203]&m[1204]&m[1205]&m[1206]&~m[1260])|(m[1203]&m[1204]&~m[1205]&~m[1206]&m[1260])|(m[1203]&~m[1204]&m[1205]&~m[1206]&m[1260])|(~m[1203]&m[1204]&m[1205]&~m[1206]&m[1260])|(m[1203]&m[1204]&m[1205]&~m[1206]&m[1260])|(m[1203]&m[1204]&m[1205]&m[1206]&m[1260]));
    m[1212] = (((m[1208]&~m[1209]&~m[1210]&~m[1211]&~m[1265])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1265])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1265])|(m[1208]&m[1209]&~m[1210]&m[1211]&~m[1265])|(m[1208]&~m[1209]&m[1210]&m[1211]&~m[1265])|(~m[1208]&m[1209]&m[1210]&m[1211]&~m[1265]))&BiasedRNG[951])|(((m[1208]&~m[1209]&~m[1210]&~m[1211]&m[1265])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&m[1265])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&m[1265])|(m[1208]&m[1209]&~m[1210]&m[1211]&m[1265])|(m[1208]&~m[1209]&m[1210]&m[1211]&m[1265])|(~m[1208]&m[1209]&m[1210]&m[1211]&m[1265]))&~BiasedRNG[951])|((m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1265])|(m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1265])|(~m[1208]&m[1209]&m[1210]&~m[1211]&~m[1265])|(m[1208]&m[1209]&m[1210]&~m[1211]&~m[1265])|(m[1208]&m[1209]&m[1210]&m[1211]&~m[1265])|(m[1208]&m[1209]&~m[1210]&~m[1211]&m[1265])|(m[1208]&~m[1209]&m[1210]&~m[1211]&m[1265])|(~m[1208]&m[1209]&m[1210]&~m[1211]&m[1265])|(m[1208]&m[1209]&m[1210]&~m[1211]&m[1265])|(m[1208]&m[1209]&m[1210]&m[1211]&m[1265]));
    m[1217] = (((m[1213]&~m[1214]&~m[1215]&~m[1216]&~m[1270])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1270])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1270])|(m[1213]&m[1214]&~m[1215]&m[1216]&~m[1270])|(m[1213]&~m[1214]&m[1215]&m[1216]&~m[1270])|(~m[1213]&m[1214]&m[1215]&m[1216]&~m[1270]))&BiasedRNG[952])|(((m[1213]&~m[1214]&~m[1215]&~m[1216]&m[1270])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&m[1270])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&m[1270])|(m[1213]&m[1214]&~m[1215]&m[1216]&m[1270])|(m[1213]&~m[1214]&m[1215]&m[1216]&m[1270])|(~m[1213]&m[1214]&m[1215]&m[1216]&m[1270]))&~BiasedRNG[952])|((m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1270])|(m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1270])|(~m[1213]&m[1214]&m[1215]&~m[1216]&~m[1270])|(m[1213]&m[1214]&m[1215]&~m[1216]&~m[1270])|(m[1213]&m[1214]&m[1215]&m[1216]&~m[1270])|(m[1213]&m[1214]&~m[1215]&~m[1216]&m[1270])|(m[1213]&~m[1214]&m[1215]&~m[1216]&m[1270])|(~m[1213]&m[1214]&m[1215]&~m[1216]&m[1270])|(m[1213]&m[1214]&m[1215]&~m[1216]&m[1270])|(m[1213]&m[1214]&m[1215]&m[1216]&m[1270]));
    m[1222] = (((m[1218]&~m[1219]&~m[1220]&~m[1221]&~m[1275])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1275])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1275])|(m[1218]&m[1219]&~m[1220]&m[1221]&~m[1275])|(m[1218]&~m[1219]&m[1220]&m[1221]&~m[1275])|(~m[1218]&m[1219]&m[1220]&m[1221]&~m[1275]))&BiasedRNG[953])|(((m[1218]&~m[1219]&~m[1220]&~m[1221]&m[1275])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&m[1275])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&m[1275])|(m[1218]&m[1219]&~m[1220]&m[1221]&m[1275])|(m[1218]&~m[1219]&m[1220]&m[1221]&m[1275])|(~m[1218]&m[1219]&m[1220]&m[1221]&m[1275]))&~BiasedRNG[953])|((m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1275])|(m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1275])|(~m[1218]&m[1219]&m[1220]&~m[1221]&~m[1275])|(m[1218]&m[1219]&m[1220]&~m[1221]&~m[1275])|(m[1218]&m[1219]&m[1220]&m[1221]&~m[1275])|(m[1218]&m[1219]&~m[1220]&~m[1221]&m[1275])|(m[1218]&~m[1219]&m[1220]&~m[1221]&m[1275])|(~m[1218]&m[1219]&m[1220]&~m[1221]&m[1275])|(m[1218]&m[1219]&m[1220]&~m[1221]&m[1275])|(m[1218]&m[1219]&m[1220]&m[1221]&m[1275]));
    m[1227] = (((m[1223]&~m[1224]&~m[1225]&~m[1226]&~m[1280])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1280])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1280])|(m[1223]&m[1224]&~m[1225]&m[1226]&~m[1280])|(m[1223]&~m[1224]&m[1225]&m[1226]&~m[1280])|(~m[1223]&m[1224]&m[1225]&m[1226]&~m[1280]))&BiasedRNG[954])|(((m[1223]&~m[1224]&~m[1225]&~m[1226]&m[1280])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&m[1280])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&m[1280])|(m[1223]&m[1224]&~m[1225]&m[1226]&m[1280])|(m[1223]&~m[1224]&m[1225]&m[1226]&m[1280])|(~m[1223]&m[1224]&m[1225]&m[1226]&m[1280]))&~BiasedRNG[954])|((m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1280])|(m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1280])|(~m[1223]&m[1224]&m[1225]&~m[1226]&~m[1280])|(m[1223]&m[1224]&m[1225]&~m[1226]&~m[1280])|(m[1223]&m[1224]&m[1225]&m[1226]&~m[1280])|(m[1223]&m[1224]&~m[1225]&~m[1226]&m[1280])|(m[1223]&~m[1224]&m[1225]&~m[1226]&m[1280])|(~m[1223]&m[1224]&m[1225]&~m[1226]&m[1280])|(m[1223]&m[1224]&m[1225]&~m[1226]&m[1280])|(m[1223]&m[1224]&m[1225]&m[1226]&m[1280]));
    m[1232] = (((m[1228]&~m[1229]&~m[1230]&~m[1231]&~m[1285])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1285])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1285])|(m[1228]&m[1229]&~m[1230]&m[1231]&~m[1285])|(m[1228]&~m[1229]&m[1230]&m[1231]&~m[1285])|(~m[1228]&m[1229]&m[1230]&m[1231]&~m[1285]))&BiasedRNG[955])|(((m[1228]&~m[1229]&~m[1230]&~m[1231]&m[1285])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&m[1285])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&m[1285])|(m[1228]&m[1229]&~m[1230]&m[1231]&m[1285])|(m[1228]&~m[1229]&m[1230]&m[1231]&m[1285])|(~m[1228]&m[1229]&m[1230]&m[1231]&m[1285]))&~BiasedRNG[955])|((m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1285])|(m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1285])|(~m[1228]&m[1229]&m[1230]&~m[1231]&~m[1285])|(m[1228]&m[1229]&m[1230]&~m[1231]&~m[1285])|(m[1228]&m[1229]&m[1230]&m[1231]&~m[1285])|(m[1228]&m[1229]&~m[1230]&~m[1231]&m[1285])|(m[1228]&~m[1229]&m[1230]&~m[1231]&m[1285])|(~m[1228]&m[1229]&m[1230]&~m[1231]&m[1285])|(m[1228]&m[1229]&m[1230]&~m[1231]&m[1285])|(m[1228]&m[1229]&m[1230]&m[1231]&m[1285]));
    m[1237] = (((m[1233]&~m[1234]&~m[1235]&~m[1236]&~m[1290])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1290])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1290])|(m[1233]&m[1234]&~m[1235]&m[1236]&~m[1290])|(m[1233]&~m[1234]&m[1235]&m[1236]&~m[1290])|(~m[1233]&m[1234]&m[1235]&m[1236]&~m[1290]))&BiasedRNG[956])|(((m[1233]&~m[1234]&~m[1235]&~m[1236]&m[1290])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&m[1290])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&m[1290])|(m[1233]&m[1234]&~m[1235]&m[1236]&m[1290])|(m[1233]&~m[1234]&m[1235]&m[1236]&m[1290])|(~m[1233]&m[1234]&m[1235]&m[1236]&m[1290]))&~BiasedRNG[956])|((m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1290])|(m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1290])|(~m[1233]&m[1234]&m[1235]&~m[1236]&~m[1290])|(m[1233]&m[1234]&m[1235]&~m[1236]&~m[1290])|(m[1233]&m[1234]&m[1235]&m[1236]&~m[1290])|(m[1233]&m[1234]&~m[1235]&~m[1236]&m[1290])|(m[1233]&~m[1234]&m[1235]&~m[1236]&m[1290])|(~m[1233]&m[1234]&m[1235]&~m[1236]&m[1290])|(m[1233]&m[1234]&m[1235]&~m[1236]&m[1290])|(m[1233]&m[1234]&m[1235]&m[1236]&m[1290]));
    m[1242] = (((m[1238]&~m[1239]&~m[1240]&~m[1241]&~m[1295])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1295])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1295])|(m[1238]&m[1239]&~m[1240]&m[1241]&~m[1295])|(m[1238]&~m[1239]&m[1240]&m[1241]&~m[1295])|(~m[1238]&m[1239]&m[1240]&m[1241]&~m[1295]))&BiasedRNG[957])|(((m[1238]&~m[1239]&~m[1240]&~m[1241]&m[1295])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&m[1295])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&m[1295])|(m[1238]&m[1239]&~m[1240]&m[1241]&m[1295])|(m[1238]&~m[1239]&m[1240]&m[1241]&m[1295])|(~m[1238]&m[1239]&m[1240]&m[1241]&m[1295]))&~BiasedRNG[957])|((m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1295])|(m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1295])|(~m[1238]&m[1239]&m[1240]&~m[1241]&~m[1295])|(m[1238]&m[1239]&m[1240]&~m[1241]&~m[1295])|(m[1238]&m[1239]&m[1240]&m[1241]&~m[1295])|(m[1238]&m[1239]&~m[1240]&~m[1241]&m[1295])|(m[1238]&~m[1239]&m[1240]&~m[1241]&m[1295])|(~m[1238]&m[1239]&m[1240]&~m[1241]&m[1295])|(m[1238]&m[1239]&m[1240]&~m[1241]&m[1295])|(m[1238]&m[1239]&m[1240]&m[1241]&m[1295]));
    m[1247] = (((m[1243]&~m[1244]&~m[1245]&~m[1246]&~m[1300])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1300])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1300])|(m[1243]&m[1244]&~m[1245]&m[1246]&~m[1300])|(m[1243]&~m[1244]&m[1245]&m[1246]&~m[1300])|(~m[1243]&m[1244]&m[1245]&m[1246]&~m[1300]))&BiasedRNG[958])|(((m[1243]&~m[1244]&~m[1245]&~m[1246]&m[1300])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&m[1300])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&m[1300])|(m[1243]&m[1244]&~m[1245]&m[1246]&m[1300])|(m[1243]&~m[1244]&m[1245]&m[1246]&m[1300])|(~m[1243]&m[1244]&m[1245]&m[1246]&m[1300]))&~BiasedRNG[958])|((m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1300])|(m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1300])|(~m[1243]&m[1244]&m[1245]&~m[1246]&~m[1300])|(m[1243]&m[1244]&m[1245]&~m[1246]&~m[1300])|(m[1243]&m[1244]&m[1245]&m[1246]&~m[1300])|(m[1243]&m[1244]&~m[1245]&~m[1246]&m[1300])|(m[1243]&~m[1244]&m[1245]&~m[1246]&m[1300])|(~m[1243]&m[1244]&m[1245]&~m[1246]&m[1300])|(m[1243]&m[1244]&m[1245]&~m[1246]&m[1300])|(m[1243]&m[1244]&m[1245]&m[1246]&m[1300]));
    m[1252] = (((m[1248]&~m[1249]&~m[1250]&~m[1251]&~m[1305])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1305])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1305])|(m[1248]&m[1249]&~m[1250]&m[1251]&~m[1305])|(m[1248]&~m[1249]&m[1250]&m[1251]&~m[1305])|(~m[1248]&m[1249]&m[1250]&m[1251]&~m[1305]))&BiasedRNG[959])|(((m[1248]&~m[1249]&~m[1250]&~m[1251]&m[1305])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&m[1305])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&m[1305])|(m[1248]&m[1249]&~m[1250]&m[1251]&m[1305])|(m[1248]&~m[1249]&m[1250]&m[1251]&m[1305])|(~m[1248]&m[1249]&m[1250]&m[1251]&m[1305]))&~BiasedRNG[959])|((m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1305])|(m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1305])|(~m[1248]&m[1249]&m[1250]&~m[1251]&~m[1305])|(m[1248]&m[1249]&m[1250]&~m[1251]&~m[1305])|(m[1248]&m[1249]&m[1250]&m[1251]&~m[1305])|(m[1248]&m[1249]&~m[1250]&~m[1251]&m[1305])|(m[1248]&~m[1249]&m[1250]&~m[1251]&m[1305])|(~m[1248]&m[1249]&m[1250]&~m[1251]&m[1305])|(m[1248]&m[1249]&m[1250]&~m[1251]&m[1305])|(m[1248]&m[1249]&m[1250]&m[1251]&m[1305]));
    m[1257] = (((m[1253]&~m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&~m[1310]))&BiasedRNG[960])|(((m[1253]&~m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&m[1310]))&~BiasedRNG[960])|((m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&m[1310]));
    m[1262] = (((m[1258]&~m[1259]&~m[1260]&~m[1261]&~m[1320])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1320])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1320])|(m[1258]&m[1259]&~m[1260]&m[1261]&~m[1320])|(m[1258]&~m[1259]&m[1260]&m[1261]&~m[1320])|(~m[1258]&m[1259]&m[1260]&m[1261]&~m[1320]))&BiasedRNG[961])|(((m[1258]&~m[1259]&~m[1260]&~m[1261]&m[1320])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&m[1320])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&m[1320])|(m[1258]&m[1259]&~m[1260]&m[1261]&m[1320])|(m[1258]&~m[1259]&m[1260]&m[1261]&m[1320])|(~m[1258]&m[1259]&m[1260]&m[1261]&m[1320]))&~BiasedRNG[961])|((m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1320])|(m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1320])|(~m[1258]&m[1259]&m[1260]&~m[1261]&~m[1320])|(m[1258]&m[1259]&m[1260]&~m[1261]&~m[1320])|(m[1258]&m[1259]&m[1260]&m[1261]&~m[1320])|(m[1258]&m[1259]&~m[1260]&~m[1261]&m[1320])|(m[1258]&~m[1259]&m[1260]&~m[1261]&m[1320])|(~m[1258]&m[1259]&m[1260]&~m[1261]&m[1320])|(m[1258]&m[1259]&m[1260]&~m[1261]&m[1320])|(m[1258]&m[1259]&m[1260]&m[1261]&m[1320]));
    m[1267] = (((m[1263]&~m[1264]&~m[1265]&~m[1266]&~m[1325])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1325])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1325])|(m[1263]&m[1264]&~m[1265]&m[1266]&~m[1325])|(m[1263]&~m[1264]&m[1265]&m[1266]&~m[1325])|(~m[1263]&m[1264]&m[1265]&m[1266]&~m[1325]))&BiasedRNG[962])|(((m[1263]&~m[1264]&~m[1265]&~m[1266]&m[1325])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&m[1325])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&m[1325])|(m[1263]&m[1264]&~m[1265]&m[1266]&m[1325])|(m[1263]&~m[1264]&m[1265]&m[1266]&m[1325])|(~m[1263]&m[1264]&m[1265]&m[1266]&m[1325]))&~BiasedRNG[962])|((m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1325])|(m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1325])|(~m[1263]&m[1264]&m[1265]&~m[1266]&~m[1325])|(m[1263]&m[1264]&m[1265]&~m[1266]&~m[1325])|(m[1263]&m[1264]&m[1265]&m[1266]&~m[1325])|(m[1263]&m[1264]&~m[1265]&~m[1266]&m[1325])|(m[1263]&~m[1264]&m[1265]&~m[1266]&m[1325])|(~m[1263]&m[1264]&m[1265]&~m[1266]&m[1325])|(m[1263]&m[1264]&m[1265]&~m[1266]&m[1325])|(m[1263]&m[1264]&m[1265]&m[1266]&m[1325]));
    m[1272] = (((m[1268]&~m[1269]&~m[1270]&~m[1271]&~m[1330])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1330])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1330])|(m[1268]&m[1269]&~m[1270]&m[1271]&~m[1330])|(m[1268]&~m[1269]&m[1270]&m[1271]&~m[1330])|(~m[1268]&m[1269]&m[1270]&m[1271]&~m[1330]))&BiasedRNG[963])|(((m[1268]&~m[1269]&~m[1270]&~m[1271]&m[1330])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&m[1330])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&m[1330])|(m[1268]&m[1269]&~m[1270]&m[1271]&m[1330])|(m[1268]&~m[1269]&m[1270]&m[1271]&m[1330])|(~m[1268]&m[1269]&m[1270]&m[1271]&m[1330]))&~BiasedRNG[963])|((m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1330])|(m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1330])|(~m[1268]&m[1269]&m[1270]&~m[1271]&~m[1330])|(m[1268]&m[1269]&m[1270]&~m[1271]&~m[1330])|(m[1268]&m[1269]&m[1270]&m[1271]&~m[1330])|(m[1268]&m[1269]&~m[1270]&~m[1271]&m[1330])|(m[1268]&~m[1269]&m[1270]&~m[1271]&m[1330])|(~m[1268]&m[1269]&m[1270]&~m[1271]&m[1330])|(m[1268]&m[1269]&m[1270]&~m[1271]&m[1330])|(m[1268]&m[1269]&m[1270]&m[1271]&m[1330]));
    m[1277] = (((m[1273]&~m[1274]&~m[1275]&~m[1276]&~m[1335])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1335])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1335])|(m[1273]&m[1274]&~m[1275]&m[1276]&~m[1335])|(m[1273]&~m[1274]&m[1275]&m[1276]&~m[1335])|(~m[1273]&m[1274]&m[1275]&m[1276]&~m[1335]))&BiasedRNG[964])|(((m[1273]&~m[1274]&~m[1275]&~m[1276]&m[1335])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&m[1335])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&m[1335])|(m[1273]&m[1274]&~m[1275]&m[1276]&m[1335])|(m[1273]&~m[1274]&m[1275]&m[1276]&m[1335])|(~m[1273]&m[1274]&m[1275]&m[1276]&m[1335]))&~BiasedRNG[964])|((m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1335])|(m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1335])|(~m[1273]&m[1274]&m[1275]&~m[1276]&~m[1335])|(m[1273]&m[1274]&m[1275]&~m[1276]&~m[1335])|(m[1273]&m[1274]&m[1275]&m[1276]&~m[1335])|(m[1273]&m[1274]&~m[1275]&~m[1276]&m[1335])|(m[1273]&~m[1274]&m[1275]&~m[1276]&m[1335])|(~m[1273]&m[1274]&m[1275]&~m[1276]&m[1335])|(m[1273]&m[1274]&m[1275]&~m[1276]&m[1335])|(m[1273]&m[1274]&m[1275]&m[1276]&m[1335]));
    m[1282] = (((m[1278]&~m[1279]&~m[1280]&~m[1281]&~m[1340])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1340])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1340])|(m[1278]&m[1279]&~m[1280]&m[1281]&~m[1340])|(m[1278]&~m[1279]&m[1280]&m[1281]&~m[1340])|(~m[1278]&m[1279]&m[1280]&m[1281]&~m[1340]))&BiasedRNG[965])|(((m[1278]&~m[1279]&~m[1280]&~m[1281]&m[1340])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&m[1340])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&m[1340])|(m[1278]&m[1279]&~m[1280]&m[1281]&m[1340])|(m[1278]&~m[1279]&m[1280]&m[1281]&m[1340])|(~m[1278]&m[1279]&m[1280]&m[1281]&m[1340]))&~BiasedRNG[965])|((m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1340])|(m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1340])|(~m[1278]&m[1279]&m[1280]&~m[1281]&~m[1340])|(m[1278]&m[1279]&m[1280]&~m[1281]&~m[1340])|(m[1278]&m[1279]&m[1280]&m[1281]&~m[1340])|(m[1278]&m[1279]&~m[1280]&~m[1281]&m[1340])|(m[1278]&~m[1279]&m[1280]&~m[1281]&m[1340])|(~m[1278]&m[1279]&m[1280]&~m[1281]&m[1340])|(m[1278]&m[1279]&m[1280]&~m[1281]&m[1340])|(m[1278]&m[1279]&m[1280]&m[1281]&m[1340]));
    m[1287] = (((m[1283]&~m[1284]&~m[1285]&~m[1286]&~m[1345])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1345])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1345])|(m[1283]&m[1284]&~m[1285]&m[1286]&~m[1345])|(m[1283]&~m[1284]&m[1285]&m[1286]&~m[1345])|(~m[1283]&m[1284]&m[1285]&m[1286]&~m[1345]))&BiasedRNG[966])|(((m[1283]&~m[1284]&~m[1285]&~m[1286]&m[1345])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&m[1345])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&m[1345])|(m[1283]&m[1284]&~m[1285]&m[1286]&m[1345])|(m[1283]&~m[1284]&m[1285]&m[1286]&m[1345])|(~m[1283]&m[1284]&m[1285]&m[1286]&m[1345]))&~BiasedRNG[966])|((m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1345])|(m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1345])|(~m[1283]&m[1284]&m[1285]&~m[1286]&~m[1345])|(m[1283]&m[1284]&m[1285]&~m[1286]&~m[1345])|(m[1283]&m[1284]&m[1285]&m[1286]&~m[1345])|(m[1283]&m[1284]&~m[1285]&~m[1286]&m[1345])|(m[1283]&~m[1284]&m[1285]&~m[1286]&m[1345])|(~m[1283]&m[1284]&m[1285]&~m[1286]&m[1345])|(m[1283]&m[1284]&m[1285]&~m[1286]&m[1345])|(m[1283]&m[1284]&m[1285]&m[1286]&m[1345]));
    m[1292] = (((m[1288]&~m[1289]&~m[1290]&~m[1291]&~m[1350])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1350])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1350])|(m[1288]&m[1289]&~m[1290]&m[1291]&~m[1350])|(m[1288]&~m[1289]&m[1290]&m[1291]&~m[1350])|(~m[1288]&m[1289]&m[1290]&m[1291]&~m[1350]))&BiasedRNG[967])|(((m[1288]&~m[1289]&~m[1290]&~m[1291]&m[1350])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&m[1350])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&m[1350])|(m[1288]&m[1289]&~m[1290]&m[1291]&m[1350])|(m[1288]&~m[1289]&m[1290]&m[1291]&m[1350])|(~m[1288]&m[1289]&m[1290]&m[1291]&m[1350]))&~BiasedRNG[967])|((m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1350])|(m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1350])|(~m[1288]&m[1289]&m[1290]&~m[1291]&~m[1350])|(m[1288]&m[1289]&m[1290]&~m[1291]&~m[1350])|(m[1288]&m[1289]&m[1290]&m[1291]&~m[1350])|(m[1288]&m[1289]&~m[1290]&~m[1291]&m[1350])|(m[1288]&~m[1289]&m[1290]&~m[1291]&m[1350])|(~m[1288]&m[1289]&m[1290]&~m[1291]&m[1350])|(m[1288]&m[1289]&m[1290]&~m[1291]&m[1350])|(m[1288]&m[1289]&m[1290]&m[1291]&m[1350]));
    m[1297] = (((m[1293]&~m[1294]&~m[1295]&~m[1296]&~m[1355])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1355])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1355])|(m[1293]&m[1294]&~m[1295]&m[1296]&~m[1355])|(m[1293]&~m[1294]&m[1295]&m[1296]&~m[1355])|(~m[1293]&m[1294]&m[1295]&m[1296]&~m[1355]))&BiasedRNG[968])|(((m[1293]&~m[1294]&~m[1295]&~m[1296]&m[1355])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&m[1355])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&m[1355])|(m[1293]&m[1294]&~m[1295]&m[1296]&m[1355])|(m[1293]&~m[1294]&m[1295]&m[1296]&m[1355])|(~m[1293]&m[1294]&m[1295]&m[1296]&m[1355]))&~BiasedRNG[968])|((m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1355])|(m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1355])|(~m[1293]&m[1294]&m[1295]&~m[1296]&~m[1355])|(m[1293]&m[1294]&m[1295]&~m[1296]&~m[1355])|(m[1293]&m[1294]&m[1295]&m[1296]&~m[1355])|(m[1293]&m[1294]&~m[1295]&~m[1296]&m[1355])|(m[1293]&~m[1294]&m[1295]&~m[1296]&m[1355])|(~m[1293]&m[1294]&m[1295]&~m[1296]&m[1355])|(m[1293]&m[1294]&m[1295]&~m[1296]&m[1355])|(m[1293]&m[1294]&m[1295]&m[1296]&m[1355]));
    m[1302] = (((m[1298]&~m[1299]&~m[1300]&~m[1301]&~m[1360])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1360])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1360])|(m[1298]&m[1299]&~m[1300]&m[1301]&~m[1360])|(m[1298]&~m[1299]&m[1300]&m[1301]&~m[1360])|(~m[1298]&m[1299]&m[1300]&m[1301]&~m[1360]))&BiasedRNG[969])|(((m[1298]&~m[1299]&~m[1300]&~m[1301]&m[1360])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&m[1360])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&m[1360])|(m[1298]&m[1299]&~m[1300]&m[1301]&m[1360])|(m[1298]&~m[1299]&m[1300]&m[1301]&m[1360])|(~m[1298]&m[1299]&m[1300]&m[1301]&m[1360]))&~BiasedRNG[969])|((m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1360])|(m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1360])|(~m[1298]&m[1299]&m[1300]&~m[1301]&~m[1360])|(m[1298]&m[1299]&m[1300]&~m[1301]&~m[1360])|(m[1298]&m[1299]&m[1300]&m[1301]&~m[1360])|(m[1298]&m[1299]&~m[1300]&~m[1301]&m[1360])|(m[1298]&~m[1299]&m[1300]&~m[1301]&m[1360])|(~m[1298]&m[1299]&m[1300]&~m[1301]&m[1360])|(m[1298]&m[1299]&m[1300]&~m[1301]&m[1360])|(m[1298]&m[1299]&m[1300]&m[1301]&m[1360]));
    m[1307] = (((m[1303]&~m[1304]&~m[1305]&~m[1306]&~m[1365])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1365])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1365])|(m[1303]&m[1304]&~m[1305]&m[1306]&~m[1365])|(m[1303]&~m[1304]&m[1305]&m[1306]&~m[1365])|(~m[1303]&m[1304]&m[1305]&m[1306]&~m[1365]))&BiasedRNG[970])|(((m[1303]&~m[1304]&~m[1305]&~m[1306]&m[1365])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&m[1365])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&m[1365])|(m[1303]&m[1304]&~m[1305]&m[1306]&m[1365])|(m[1303]&~m[1304]&m[1305]&m[1306]&m[1365])|(~m[1303]&m[1304]&m[1305]&m[1306]&m[1365]))&~BiasedRNG[970])|((m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1365])|(m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1365])|(~m[1303]&m[1304]&m[1305]&~m[1306]&~m[1365])|(m[1303]&m[1304]&m[1305]&~m[1306]&~m[1365])|(m[1303]&m[1304]&m[1305]&m[1306]&~m[1365])|(m[1303]&m[1304]&~m[1305]&~m[1306]&m[1365])|(m[1303]&~m[1304]&m[1305]&~m[1306]&m[1365])|(~m[1303]&m[1304]&m[1305]&~m[1306]&m[1365])|(m[1303]&m[1304]&m[1305]&~m[1306]&m[1365])|(m[1303]&m[1304]&m[1305]&m[1306]&m[1365]));
    m[1312] = (((m[1308]&~m[1309]&~m[1310]&~m[1311]&~m[1370])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1370])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1370])|(m[1308]&m[1309]&~m[1310]&m[1311]&~m[1370])|(m[1308]&~m[1309]&m[1310]&m[1311]&~m[1370])|(~m[1308]&m[1309]&m[1310]&m[1311]&~m[1370]))&BiasedRNG[971])|(((m[1308]&~m[1309]&~m[1310]&~m[1311]&m[1370])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&m[1370])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&m[1370])|(m[1308]&m[1309]&~m[1310]&m[1311]&m[1370])|(m[1308]&~m[1309]&m[1310]&m[1311]&m[1370])|(~m[1308]&m[1309]&m[1310]&m[1311]&m[1370]))&~BiasedRNG[971])|((m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1370])|(m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1370])|(~m[1308]&m[1309]&m[1310]&~m[1311]&~m[1370])|(m[1308]&m[1309]&m[1310]&~m[1311]&~m[1370])|(m[1308]&m[1309]&m[1310]&m[1311]&~m[1370])|(m[1308]&m[1309]&~m[1310]&~m[1311]&m[1370])|(m[1308]&~m[1309]&m[1310]&~m[1311]&m[1370])|(~m[1308]&m[1309]&m[1310]&~m[1311]&m[1370])|(m[1308]&m[1309]&m[1310]&~m[1311]&m[1370])|(m[1308]&m[1309]&m[1310]&m[1311]&m[1370]));
    m[1317] = (((m[1313]&~m[1314]&~m[1315]&~m[1316]&~m[1375])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1375])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1375])|(m[1313]&m[1314]&~m[1315]&m[1316]&~m[1375])|(m[1313]&~m[1314]&m[1315]&m[1316]&~m[1375])|(~m[1313]&m[1314]&m[1315]&m[1316]&~m[1375]))&BiasedRNG[972])|(((m[1313]&~m[1314]&~m[1315]&~m[1316]&m[1375])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&m[1375])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&m[1375])|(m[1313]&m[1314]&~m[1315]&m[1316]&m[1375])|(m[1313]&~m[1314]&m[1315]&m[1316]&m[1375])|(~m[1313]&m[1314]&m[1315]&m[1316]&m[1375]))&~BiasedRNG[972])|((m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1375])|(m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1375])|(~m[1313]&m[1314]&m[1315]&~m[1316]&~m[1375])|(m[1313]&m[1314]&m[1315]&~m[1316]&~m[1375])|(m[1313]&m[1314]&m[1315]&m[1316]&~m[1375])|(m[1313]&m[1314]&~m[1315]&~m[1316]&m[1375])|(m[1313]&~m[1314]&m[1315]&~m[1316]&m[1375])|(~m[1313]&m[1314]&m[1315]&~m[1316]&m[1375])|(m[1313]&m[1314]&m[1315]&~m[1316]&m[1375])|(m[1313]&m[1314]&m[1315]&m[1316]&m[1375]));
    m[1322] = (((m[1318]&~m[1319]&~m[1320]&~m[1321]&~m[1385])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1385])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1385])|(m[1318]&m[1319]&~m[1320]&m[1321]&~m[1385])|(m[1318]&~m[1319]&m[1320]&m[1321]&~m[1385])|(~m[1318]&m[1319]&m[1320]&m[1321]&~m[1385]))&BiasedRNG[973])|(((m[1318]&~m[1319]&~m[1320]&~m[1321]&m[1385])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&m[1385])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&m[1385])|(m[1318]&m[1319]&~m[1320]&m[1321]&m[1385])|(m[1318]&~m[1319]&m[1320]&m[1321]&m[1385])|(~m[1318]&m[1319]&m[1320]&m[1321]&m[1385]))&~BiasedRNG[973])|((m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1385])|(m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1385])|(~m[1318]&m[1319]&m[1320]&~m[1321]&~m[1385])|(m[1318]&m[1319]&m[1320]&~m[1321]&~m[1385])|(m[1318]&m[1319]&m[1320]&m[1321]&~m[1385])|(m[1318]&m[1319]&~m[1320]&~m[1321]&m[1385])|(m[1318]&~m[1319]&m[1320]&~m[1321]&m[1385])|(~m[1318]&m[1319]&m[1320]&~m[1321]&m[1385])|(m[1318]&m[1319]&m[1320]&~m[1321]&m[1385])|(m[1318]&m[1319]&m[1320]&m[1321]&m[1385]));
    m[1327] = (((m[1323]&~m[1324]&~m[1325]&~m[1326]&~m[1390])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1390])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1390])|(m[1323]&m[1324]&~m[1325]&m[1326]&~m[1390])|(m[1323]&~m[1324]&m[1325]&m[1326]&~m[1390])|(~m[1323]&m[1324]&m[1325]&m[1326]&~m[1390]))&BiasedRNG[974])|(((m[1323]&~m[1324]&~m[1325]&~m[1326]&m[1390])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&m[1390])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&m[1390])|(m[1323]&m[1324]&~m[1325]&m[1326]&m[1390])|(m[1323]&~m[1324]&m[1325]&m[1326]&m[1390])|(~m[1323]&m[1324]&m[1325]&m[1326]&m[1390]))&~BiasedRNG[974])|((m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1390])|(m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1390])|(~m[1323]&m[1324]&m[1325]&~m[1326]&~m[1390])|(m[1323]&m[1324]&m[1325]&~m[1326]&~m[1390])|(m[1323]&m[1324]&m[1325]&m[1326]&~m[1390])|(m[1323]&m[1324]&~m[1325]&~m[1326]&m[1390])|(m[1323]&~m[1324]&m[1325]&~m[1326]&m[1390])|(~m[1323]&m[1324]&m[1325]&~m[1326]&m[1390])|(m[1323]&m[1324]&m[1325]&~m[1326]&m[1390])|(m[1323]&m[1324]&m[1325]&m[1326]&m[1390]));
    m[1332] = (((m[1328]&~m[1329]&~m[1330]&~m[1331]&~m[1395])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1395])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1395])|(m[1328]&m[1329]&~m[1330]&m[1331]&~m[1395])|(m[1328]&~m[1329]&m[1330]&m[1331]&~m[1395])|(~m[1328]&m[1329]&m[1330]&m[1331]&~m[1395]))&BiasedRNG[975])|(((m[1328]&~m[1329]&~m[1330]&~m[1331]&m[1395])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&m[1395])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&m[1395])|(m[1328]&m[1329]&~m[1330]&m[1331]&m[1395])|(m[1328]&~m[1329]&m[1330]&m[1331]&m[1395])|(~m[1328]&m[1329]&m[1330]&m[1331]&m[1395]))&~BiasedRNG[975])|((m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1395])|(m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1395])|(~m[1328]&m[1329]&m[1330]&~m[1331]&~m[1395])|(m[1328]&m[1329]&m[1330]&~m[1331]&~m[1395])|(m[1328]&m[1329]&m[1330]&m[1331]&~m[1395])|(m[1328]&m[1329]&~m[1330]&~m[1331]&m[1395])|(m[1328]&~m[1329]&m[1330]&~m[1331]&m[1395])|(~m[1328]&m[1329]&m[1330]&~m[1331]&m[1395])|(m[1328]&m[1329]&m[1330]&~m[1331]&m[1395])|(m[1328]&m[1329]&m[1330]&m[1331]&m[1395]));
    m[1337] = (((m[1333]&~m[1334]&~m[1335]&~m[1336]&~m[1400])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1400])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1400])|(m[1333]&m[1334]&~m[1335]&m[1336]&~m[1400])|(m[1333]&~m[1334]&m[1335]&m[1336]&~m[1400])|(~m[1333]&m[1334]&m[1335]&m[1336]&~m[1400]))&BiasedRNG[976])|(((m[1333]&~m[1334]&~m[1335]&~m[1336]&m[1400])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&m[1400])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&m[1400])|(m[1333]&m[1334]&~m[1335]&m[1336]&m[1400])|(m[1333]&~m[1334]&m[1335]&m[1336]&m[1400])|(~m[1333]&m[1334]&m[1335]&m[1336]&m[1400]))&~BiasedRNG[976])|((m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1400])|(m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1400])|(~m[1333]&m[1334]&m[1335]&~m[1336]&~m[1400])|(m[1333]&m[1334]&m[1335]&~m[1336]&~m[1400])|(m[1333]&m[1334]&m[1335]&m[1336]&~m[1400])|(m[1333]&m[1334]&~m[1335]&~m[1336]&m[1400])|(m[1333]&~m[1334]&m[1335]&~m[1336]&m[1400])|(~m[1333]&m[1334]&m[1335]&~m[1336]&m[1400])|(m[1333]&m[1334]&m[1335]&~m[1336]&m[1400])|(m[1333]&m[1334]&m[1335]&m[1336]&m[1400]));
    m[1342] = (((m[1338]&~m[1339]&~m[1340]&~m[1341]&~m[1405])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1405])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1405])|(m[1338]&m[1339]&~m[1340]&m[1341]&~m[1405])|(m[1338]&~m[1339]&m[1340]&m[1341]&~m[1405])|(~m[1338]&m[1339]&m[1340]&m[1341]&~m[1405]))&BiasedRNG[977])|(((m[1338]&~m[1339]&~m[1340]&~m[1341]&m[1405])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&m[1405])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&m[1405])|(m[1338]&m[1339]&~m[1340]&m[1341]&m[1405])|(m[1338]&~m[1339]&m[1340]&m[1341]&m[1405])|(~m[1338]&m[1339]&m[1340]&m[1341]&m[1405]))&~BiasedRNG[977])|((m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1405])|(m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1405])|(~m[1338]&m[1339]&m[1340]&~m[1341]&~m[1405])|(m[1338]&m[1339]&m[1340]&~m[1341]&~m[1405])|(m[1338]&m[1339]&m[1340]&m[1341]&~m[1405])|(m[1338]&m[1339]&~m[1340]&~m[1341]&m[1405])|(m[1338]&~m[1339]&m[1340]&~m[1341]&m[1405])|(~m[1338]&m[1339]&m[1340]&~m[1341]&m[1405])|(m[1338]&m[1339]&m[1340]&~m[1341]&m[1405])|(m[1338]&m[1339]&m[1340]&m[1341]&m[1405]));
    m[1347] = (((m[1343]&~m[1344]&~m[1345]&~m[1346]&~m[1410])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1410])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1410])|(m[1343]&m[1344]&~m[1345]&m[1346]&~m[1410])|(m[1343]&~m[1344]&m[1345]&m[1346]&~m[1410])|(~m[1343]&m[1344]&m[1345]&m[1346]&~m[1410]))&BiasedRNG[978])|(((m[1343]&~m[1344]&~m[1345]&~m[1346]&m[1410])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&m[1410])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&m[1410])|(m[1343]&m[1344]&~m[1345]&m[1346]&m[1410])|(m[1343]&~m[1344]&m[1345]&m[1346]&m[1410])|(~m[1343]&m[1344]&m[1345]&m[1346]&m[1410]))&~BiasedRNG[978])|((m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1410])|(m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1410])|(~m[1343]&m[1344]&m[1345]&~m[1346]&~m[1410])|(m[1343]&m[1344]&m[1345]&~m[1346]&~m[1410])|(m[1343]&m[1344]&m[1345]&m[1346]&~m[1410])|(m[1343]&m[1344]&~m[1345]&~m[1346]&m[1410])|(m[1343]&~m[1344]&m[1345]&~m[1346]&m[1410])|(~m[1343]&m[1344]&m[1345]&~m[1346]&m[1410])|(m[1343]&m[1344]&m[1345]&~m[1346]&m[1410])|(m[1343]&m[1344]&m[1345]&m[1346]&m[1410]));
    m[1352] = (((m[1348]&~m[1349]&~m[1350]&~m[1351]&~m[1415])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1415])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1415])|(m[1348]&m[1349]&~m[1350]&m[1351]&~m[1415])|(m[1348]&~m[1349]&m[1350]&m[1351]&~m[1415])|(~m[1348]&m[1349]&m[1350]&m[1351]&~m[1415]))&BiasedRNG[979])|(((m[1348]&~m[1349]&~m[1350]&~m[1351]&m[1415])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&m[1415])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&m[1415])|(m[1348]&m[1349]&~m[1350]&m[1351]&m[1415])|(m[1348]&~m[1349]&m[1350]&m[1351]&m[1415])|(~m[1348]&m[1349]&m[1350]&m[1351]&m[1415]))&~BiasedRNG[979])|((m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1415])|(m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1415])|(~m[1348]&m[1349]&m[1350]&~m[1351]&~m[1415])|(m[1348]&m[1349]&m[1350]&~m[1351]&~m[1415])|(m[1348]&m[1349]&m[1350]&m[1351]&~m[1415])|(m[1348]&m[1349]&~m[1350]&~m[1351]&m[1415])|(m[1348]&~m[1349]&m[1350]&~m[1351]&m[1415])|(~m[1348]&m[1349]&m[1350]&~m[1351]&m[1415])|(m[1348]&m[1349]&m[1350]&~m[1351]&m[1415])|(m[1348]&m[1349]&m[1350]&m[1351]&m[1415]));
    m[1357] = (((m[1353]&~m[1354]&~m[1355]&~m[1356]&~m[1420])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1420])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1420])|(m[1353]&m[1354]&~m[1355]&m[1356]&~m[1420])|(m[1353]&~m[1354]&m[1355]&m[1356]&~m[1420])|(~m[1353]&m[1354]&m[1355]&m[1356]&~m[1420]))&BiasedRNG[980])|(((m[1353]&~m[1354]&~m[1355]&~m[1356]&m[1420])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&m[1420])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&m[1420])|(m[1353]&m[1354]&~m[1355]&m[1356]&m[1420])|(m[1353]&~m[1354]&m[1355]&m[1356]&m[1420])|(~m[1353]&m[1354]&m[1355]&m[1356]&m[1420]))&~BiasedRNG[980])|((m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1420])|(m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1420])|(~m[1353]&m[1354]&m[1355]&~m[1356]&~m[1420])|(m[1353]&m[1354]&m[1355]&~m[1356]&~m[1420])|(m[1353]&m[1354]&m[1355]&m[1356]&~m[1420])|(m[1353]&m[1354]&~m[1355]&~m[1356]&m[1420])|(m[1353]&~m[1354]&m[1355]&~m[1356]&m[1420])|(~m[1353]&m[1354]&m[1355]&~m[1356]&m[1420])|(m[1353]&m[1354]&m[1355]&~m[1356]&m[1420])|(m[1353]&m[1354]&m[1355]&m[1356]&m[1420]));
    m[1362] = (((m[1358]&~m[1359]&~m[1360]&~m[1361]&~m[1425])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1425])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1425])|(m[1358]&m[1359]&~m[1360]&m[1361]&~m[1425])|(m[1358]&~m[1359]&m[1360]&m[1361]&~m[1425])|(~m[1358]&m[1359]&m[1360]&m[1361]&~m[1425]))&BiasedRNG[981])|(((m[1358]&~m[1359]&~m[1360]&~m[1361]&m[1425])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&m[1425])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&m[1425])|(m[1358]&m[1359]&~m[1360]&m[1361]&m[1425])|(m[1358]&~m[1359]&m[1360]&m[1361]&m[1425])|(~m[1358]&m[1359]&m[1360]&m[1361]&m[1425]))&~BiasedRNG[981])|((m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1425])|(m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1425])|(~m[1358]&m[1359]&m[1360]&~m[1361]&~m[1425])|(m[1358]&m[1359]&m[1360]&~m[1361]&~m[1425])|(m[1358]&m[1359]&m[1360]&m[1361]&~m[1425])|(m[1358]&m[1359]&~m[1360]&~m[1361]&m[1425])|(m[1358]&~m[1359]&m[1360]&~m[1361]&m[1425])|(~m[1358]&m[1359]&m[1360]&~m[1361]&m[1425])|(m[1358]&m[1359]&m[1360]&~m[1361]&m[1425])|(m[1358]&m[1359]&m[1360]&m[1361]&m[1425]));
    m[1367] = (((m[1363]&~m[1364]&~m[1365]&~m[1366]&~m[1430])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1430])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1430])|(m[1363]&m[1364]&~m[1365]&m[1366]&~m[1430])|(m[1363]&~m[1364]&m[1365]&m[1366]&~m[1430])|(~m[1363]&m[1364]&m[1365]&m[1366]&~m[1430]))&BiasedRNG[982])|(((m[1363]&~m[1364]&~m[1365]&~m[1366]&m[1430])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&m[1430])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&m[1430])|(m[1363]&m[1364]&~m[1365]&m[1366]&m[1430])|(m[1363]&~m[1364]&m[1365]&m[1366]&m[1430])|(~m[1363]&m[1364]&m[1365]&m[1366]&m[1430]))&~BiasedRNG[982])|((m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1430])|(m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1430])|(~m[1363]&m[1364]&m[1365]&~m[1366]&~m[1430])|(m[1363]&m[1364]&m[1365]&~m[1366]&~m[1430])|(m[1363]&m[1364]&m[1365]&m[1366]&~m[1430])|(m[1363]&m[1364]&~m[1365]&~m[1366]&m[1430])|(m[1363]&~m[1364]&m[1365]&~m[1366]&m[1430])|(~m[1363]&m[1364]&m[1365]&~m[1366]&m[1430])|(m[1363]&m[1364]&m[1365]&~m[1366]&m[1430])|(m[1363]&m[1364]&m[1365]&m[1366]&m[1430]));
    m[1372] = (((m[1368]&~m[1369]&~m[1370]&~m[1371]&~m[1435])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1435])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1435])|(m[1368]&m[1369]&~m[1370]&m[1371]&~m[1435])|(m[1368]&~m[1369]&m[1370]&m[1371]&~m[1435])|(~m[1368]&m[1369]&m[1370]&m[1371]&~m[1435]))&BiasedRNG[983])|(((m[1368]&~m[1369]&~m[1370]&~m[1371]&m[1435])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&m[1435])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&m[1435])|(m[1368]&m[1369]&~m[1370]&m[1371]&m[1435])|(m[1368]&~m[1369]&m[1370]&m[1371]&m[1435])|(~m[1368]&m[1369]&m[1370]&m[1371]&m[1435]))&~BiasedRNG[983])|((m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1435])|(m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1435])|(~m[1368]&m[1369]&m[1370]&~m[1371]&~m[1435])|(m[1368]&m[1369]&m[1370]&~m[1371]&~m[1435])|(m[1368]&m[1369]&m[1370]&m[1371]&~m[1435])|(m[1368]&m[1369]&~m[1370]&~m[1371]&m[1435])|(m[1368]&~m[1369]&m[1370]&~m[1371]&m[1435])|(~m[1368]&m[1369]&m[1370]&~m[1371]&m[1435])|(m[1368]&m[1369]&m[1370]&~m[1371]&m[1435])|(m[1368]&m[1369]&m[1370]&m[1371]&m[1435]));
    m[1377] = (((m[1373]&~m[1374]&~m[1375]&~m[1376]&~m[1440])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1440])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1440])|(m[1373]&m[1374]&~m[1375]&m[1376]&~m[1440])|(m[1373]&~m[1374]&m[1375]&m[1376]&~m[1440])|(~m[1373]&m[1374]&m[1375]&m[1376]&~m[1440]))&BiasedRNG[984])|(((m[1373]&~m[1374]&~m[1375]&~m[1376]&m[1440])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&m[1440])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&m[1440])|(m[1373]&m[1374]&~m[1375]&m[1376]&m[1440])|(m[1373]&~m[1374]&m[1375]&m[1376]&m[1440])|(~m[1373]&m[1374]&m[1375]&m[1376]&m[1440]))&~BiasedRNG[984])|((m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1440])|(m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1440])|(~m[1373]&m[1374]&m[1375]&~m[1376]&~m[1440])|(m[1373]&m[1374]&m[1375]&~m[1376]&~m[1440])|(m[1373]&m[1374]&m[1375]&m[1376]&~m[1440])|(m[1373]&m[1374]&~m[1375]&~m[1376]&m[1440])|(m[1373]&~m[1374]&m[1375]&~m[1376]&m[1440])|(~m[1373]&m[1374]&m[1375]&~m[1376]&m[1440])|(m[1373]&m[1374]&m[1375]&~m[1376]&m[1440])|(m[1373]&m[1374]&m[1375]&m[1376]&m[1440]));
    m[1382] = (((m[1378]&~m[1379]&~m[1380]&~m[1381]&~m[1445])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1445])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1445])|(m[1378]&m[1379]&~m[1380]&m[1381]&~m[1445])|(m[1378]&~m[1379]&m[1380]&m[1381]&~m[1445])|(~m[1378]&m[1379]&m[1380]&m[1381]&~m[1445]))&BiasedRNG[985])|(((m[1378]&~m[1379]&~m[1380]&~m[1381]&m[1445])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&m[1445])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&m[1445])|(m[1378]&m[1379]&~m[1380]&m[1381]&m[1445])|(m[1378]&~m[1379]&m[1380]&m[1381]&m[1445])|(~m[1378]&m[1379]&m[1380]&m[1381]&m[1445]))&~BiasedRNG[985])|((m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1445])|(m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1445])|(~m[1378]&m[1379]&m[1380]&~m[1381]&~m[1445])|(m[1378]&m[1379]&m[1380]&~m[1381]&~m[1445])|(m[1378]&m[1379]&m[1380]&m[1381]&~m[1445])|(m[1378]&m[1379]&~m[1380]&~m[1381]&m[1445])|(m[1378]&~m[1379]&m[1380]&~m[1381]&m[1445])|(~m[1378]&m[1379]&m[1380]&~m[1381]&m[1445])|(m[1378]&m[1379]&m[1380]&~m[1381]&m[1445])|(m[1378]&m[1379]&m[1380]&m[1381]&m[1445]));
    m[1387] = (((m[1383]&~m[1384]&~m[1385]&~m[1386]&~m[1455])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1455])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1455])|(m[1383]&m[1384]&~m[1385]&m[1386]&~m[1455])|(m[1383]&~m[1384]&m[1385]&m[1386]&~m[1455])|(~m[1383]&m[1384]&m[1385]&m[1386]&~m[1455]))&BiasedRNG[986])|(((m[1383]&~m[1384]&~m[1385]&~m[1386]&m[1455])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&m[1455])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&m[1455])|(m[1383]&m[1384]&~m[1385]&m[1386]&m[1455])|(m[1383]&~m[1384]&m[1385]&m[1386]&m[1455])|(~m[1383]&m[1384]&m[1385]&m[1386]&m[1455]))&~BiasedRNG[986])|((m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1455])|(m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1455])|(~m[1383]&m[1384]&m[1385]&~m[1386]&~m[1455])|(m[1383]&m[1384]&m[1385]&~m[1386]&~m[1455])|(m[1383]&m[1384]&m[1385]&m[1386]&~m[1455])|(m[1383]&m[1384]&~m[1385]&~m[1386]&m[1455])|(m[1383]&~m[1384]&m[1385]&~m[1386]&m[1455])|(~m[1383]&m[1384]&m[1385]&~m[1386]&m[1455])|(m[1383]&m[1384]&m[1385]&~m[1386]&m[1455])|(m[1383]&m[1384]&m[1385]&m[1386]&m[1455]));
    m[1392] = (((m[1388]&~m[1389]&~m[1390]&~m[1391]&~m[1460])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1460])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1460])|(m[1388]&m[1389]&~m[1390]&m[1391]&~m[1460])|(m[1388]&~m[1389]&m[1390]&m[1391]&~m[1460])|(~m[1388]&m[1389]&m[1390]&m[1391]&~m[1460]))&BiasedRNG[987])|(((m[1388]&~m[1389]&~m[1390]&~m[1391]&m[1460])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&m[1460])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&m[1460])|(m[1388]&m[1389]&~m[1390]&m[1391]&m[1460])|(m[1388]&~m[1389]&m[1390]&m[1391]&m[1460])|(~m[1388]&m[1389]&m[1390]&m[1391]&m[1460]))&~BiasedRNG[987])|((m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1460])|(m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1460])|(~m[1388]&m[1389]&m[1390]&~m[1391]&~m[1460])|(m[1388]&m[1389]&m[1390]&~m[1391]&~m[1460])|(m[1388]&m[1389]&m[1390]&m[1391]&~m[1460])|(m[1388]&m[1389]&~m[1390]&~m[1391]&m[1460])|(m[1388]&~m[1389]&m[1390]&~m[1391]&m[1460])|(~m[1388]&m[1389]&m[1390]&~m[1391]&m[1460])|(m[1388]&m[1389]&m[1390]&~m[1391]&m[1460])|(m[1388]&m[1389]&m[1390]&m[1391]&m[1460]));
    m[1397] = (((m[1393]&~m[1394]&~m[1395]&~m[1396]&~m[1465])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1465])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1465])|(m[1393]&m[1394]&~m[1395]&m[1396]&~m[1465])|(m[1393]&~m[1394]&m[1395]&m[1396]&~m[1465])|(~m[1393]&m[1394]&m[1395]&m[1396]&~m[1465]))&BiasedRNG[988])|(((m[1393]&~m[1394]&~m[1395]&~m[1396]&m[1465])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&m[1465])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&m[1465])|(m[1393]&m[1394]&~m[1395]&m[1396]&m[1465])|(m[1393]&~m[1394]&m[1395]&m[1396]&m[1465])|(~m[1393]&m[1394]&m[1395]&m[1396]&m[1465]))&~BiasedRNG[988])|((m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1465])|(m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1465])|(~m[1393]&m[1394]&m[1395]&~m[1396]&~m[1465])|(m[1393]&m[1394]&m[1395]&~m[1396]&~m[1465])|(m[1393]&m[1394]&m[1395]&m[1396]&~m[1465])|(m[1393]&m[1394]&~m[1395]&~m[1396]&m[1465])|(m[1393]&~m[1394]&m[1395]&~m[1396]&m[1465])|(~m[1393]&m[1394]&m[1395]&~m[1396]&m[1465])|(m[1393]&m[1394]&m[1395]&~m[1396]&m[1465])|(m[1393]&m[1394]&m[1395]&m[1396]&m[1465]));
    m[1402] = (((m[1398]&~m[1399]&~m[1400]&~m[1401]&~m[1470])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1470])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1470])|(m[1398]&m[1399]&~m[1400]&m[1401]&~m[1470])|(m[1398]&~m[1399]&m[1400]&m[1401]&~m[1470])|(~m[1398]&m[1399]&m[1400]&m[1401]&~m[1470]))&BiasedRNG[989])|(((m[1398]&~m[1399]&~m[1400]&~m[1401]&m[1470])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&m[1470])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&m[1470])|(m[1398]&m[1399]&~m[1400]&m[1401]&m[1470])|(m[1398]&~m[1399]&m[1400]&m[1401]&m[1470])|(~m[1398]&m[1399]&m[1400]&m[1401]&m[1470]))&~BiasedRNG[989])|((m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1470])|(m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1470])|(~m[1398]&m[1399]&m[1400]&~m[1401]&~m[1470])|(m[1398]&m[1399]&m[1400]&~m[1401]&~m[1470])|(m[1398]&m[1399]&m[1400]&m[1401]&~m[1470])|(m[1398]&m[1399]&~m[1400]&~m[1401]&m[1470])|(m[1398]&~m[1399]&m[1400]&~m[1401]&m[1470])|(~m[1398]&m[1399]&m[1400]&~m[1401]&m[1470])|(m[1398]&m[1399]&m[1400]&~m[1401]&m[1470])|(m[1398]&m[1399]&m[1400]&m[1401]&m[1470]));
    m[1407] = (((m[1403]&~m[1404]&~m[1405]&~m[1406]&~m[1475])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1475])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1475])|(m[1403]&m[1404]&~m[1405]&m[1406]&~m[1475])|(m[1403]&~m[1404]&m[1405]&m[1406]&~m[1475])|(~m[1403]&m[1404]&m[1405]&m[1406]&~m[1475]))&BiasedRNG[990])|(((m[1403]&~m[1404]&~m[1405]&~m[1406]&m[1475])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&m[1475])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&m[1475])|(m[1403]&m[1404]&~m[1405]&m[1406]&m[1475])|(m[1403]&~m[1404]&m[1405]&m[1406]&m[1475])|(~m[1403]&m[1404]&m[1405]&m[1406]&m[1475]))&~BiasedRNG[990])|((m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1475])|(m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1475])|(~m[1403]&m[1404]&m[1405]&~m[1406]&~m[1475])|(m[1403]&m[1404]&m[1405]&~m[1406]&~m[1475])|(m[1403]&m[1404]&m[1405]&m[1406]&~m[1475])|(m[1403]&m[1404]&~m[1405]&~m[1406]&m[1475])|(m[1403]&~m[1404]&m[1405]&~m[1406]&m[1475])|(~m[1403]&m[1404]&m[1405]&~m[1406]&m[1475])|(m[1403]&m[1404]&m[1405]&~m[1406]&m[1475])|(m[1403]&m[1404]&m[1405]&m[1406]&m[1475]));
    m[1412] = (((m[1408]&~m[1409]&~m[1410]&~m[1411]&~m[1480])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1480])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1480])|(m[1408]&m[1409]&~m[1410]&m[1411]&~m[1480])|(m[1408]&~m[1409]&m[1410]&m[1411]&~m[1480])|(~m[1408]&m[1409]&m[1410]&m[1411]&~m[1480]))&BiasedRNG[991])|(((m[1408]&~m[1409]&~m[1410]&~m[1411]&m[1480])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&m[1480])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&m[1480])|(m[1408]&m[1409]&~m[1410]&m[1411]&m[1480])|(m[1408]&~m[1409]&m[1410]&m[1411]&m[1480])|(~m[1408]&m[1409]&m[1410]&m[1411]&m[1480]))&~BiasedRNG[991])|((m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1480])|(m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1480])|(~m[1408]&m[1409]&m[1410]&~m[1411]&~m[1480])|(m[1408]&m[1409]&m[1410]&~m[1411]&~m[1480])|(m[1408]&m[1409]&m[1410]&m[1411]&~m[1480])|(m[1408]&m[1409]&~m[1410]&~m[1411]&m[1480])|(m[1408]&~m[1409]&m[1410]&~m[1411]&m[1480])|(~m[1408]&m[1409]&m[1410]&~m[1411]&m[1480])|(m[1408]&m[1409]&m[1410]&~m[1411]&m[1480])|(m[1408]&m[1409]&m[1410]&m[1411]&m[1480]));
    m[1417] = (((m[1413]&~m[1414]&~m[1415]&~m[1416]&~m[1485])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1485])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1485])|(m[1413]&m[1414]&~m[1415]&m[1416]&~m[1485])|(m[1413]&~m[1414]&m[1415]&m[1416]&~m[1485])|(~m[1413]&m[1414]&m[1415]&m[1416]&~m[1485]))&BiasedRNG[992])|(((m[1413]&~m[1414]&~m[1415]&~m[1416]&m[1485])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&m[1485])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&m[1485])|(m[1413]&m[1414]&~m[1415]&m[1416]&m[1485])|(m[1413]&~m[1414]&m[1415]&m[1416]&m[1485])|(~m[1413]&m[1414]&m[1415]&m[1416]&m[1485]))&~BiasedRNG[992])|((m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1485])|(m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1485])|(~m[1413]&m[1414]&m[1415]&~m[1416]&~m[1485])|(m[1413]&m[1414]&m[1415]&~m[1416]&~m[1485])|(m[1413]&m[1414]&m[1415]&m[1416]&~m[1485])|(m[1413]&m[1414]&~m[1415]&~m[1416]&m[1485])|(m[1413]&~m[1414]&m[1415]&~m[1416]&m[1485])|(~m[1413]&m[1414]&m[1415]&~m[1416]&m[1485])|(m[1413]&m[1414]&m[1415]&~m[1416]&m[1485])|(m[1413]&m[1414]&m[1415]&m[1416]&m[1485]));
    m[1422] = (((m[1418]&~m[1419]&~m[1420]&~m[1421]&~m[1490])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1490])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1490])|(m[1418]&m[1419]&~m[1420]&m[1421]&~m[1490])|(m[1418]&~m[1419]&m[1420]&m[1421]&~m[1490])|(~m[1418]&m[1419]&m[1420]&m[1421]&~m[1490]))&BiasedRNG[993])|(((m[1418]&~m[1419]&~m[1420]&~m[1421]&m[1490])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&m[1490])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&m[1490])|(m[1418]&m[1419]&~m[1420]&m[1421]&m[1490])|(m[1418]&~m[1419]&m[1420]&m[1421]&m[1490])|(~m[1418]&m[1419]&m[1420]&m[1421]&m[1490]))&~BiasedRNG[993])|((m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1490])|(m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1490])|(~m[1418]&m[1419]&m[1420]&~m[1421]&~m[1490])|(m[1418]&m[1419]&m[1420]&~m[1421]&~m[1490])|(m[1418]&m[1419]&m[1420]&m[1421]&~m[1490])|(m[1418]&m[1419]&~m[1420]&~m[1421]&m[1490])|(m[1418]&~m[1419]&m[1420]&~m[1421]&m[1490])|(~m[1418]&m[1419]&m[1420]&~m[1421]&m[1490])|(m[1418]&m[1419]&m[1420]&~m[1421]&m[1490])|(m[1418]&m[1419]&m[1420]&m[1421]&m[1490]));
    m[1427] = (((m[1423]&~m[1424]&~m[1425]&~m[1426]&~m[1495])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1495])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1495])|(m[1423]&m[1424]&~m[1425]&m[1426]&~m[1495])|(m[1423]&~m[1424]&m[1425]&m[1426]&~m[1495])|(~m[1423]&m[1424]&m[1425]&m[1426]&~m[1495]))&BiasedRNG[994])|(((m[1423]&~m[1424]&~m[1425]&~m[1426]&m[1495])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&m[1495])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&m[1495])|(m[1423]&m[1424]&~m[1425]&m[1426]&m[1495])|(m[1423]&~m[1424]&m[1425]&m[1426]&m[1495])|(~m[1423]&m[1424]&m[1425]&m[1426]&m[1495]))&~BiasedRNG[994])|((m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1495])|(m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1495])|(~m[1423]&m[1424]&m[1425]&~m[1426]&~m[1495])|(m[1423]&m[1424]&m[1425]&~m[1426]&~m[1495])|(m[1423]&m[1424]&m[1425]&m[1426]&~m[1495])|(m[1423]&m[1424]&~m[1425]&~m[1426]&m[1495])|(m[1423]&~m[1424]&m[1425]&~m[1426]&m[1495])|(~m[1423]&m[1424]&m[1425]&~m[1426]&m[1495])|(m[1423]&m[1424]&m[1425]&~m[1426]&m[1495])|(m[1423]&m[1424]&m[1425]&m[1426]&m[1495]));
    m[1432] = (((m[1428]&~m[1429]&~m[1430]&~m[1431]&~m[1500])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1500])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1500])|(m[1428]&m[1429]&~m[1430]&m[1431]&~m[1500])|(m[1428]&~m[1429]&m[1430]&m[1431]&~m[1500])|(~m[1428]&m[1429]&m[1430]&m[1431]&~m[1500]))&BiasedRNG[995])|(((m[1428]&~m[1429]&~m[1430]&~m[1431]&m[1500])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&m[1500])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&m[1500])|(m[1428]&m[1429]&~m[1430]&m[1431]&m[1500])|(m[1428]&~m[1429]&m[1430]&m[1431]&m[1500])|(~m[1428]&m[1429]&m[1430]&m[1431]&m[1500]))&~BiasedRNG[995])|((m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1500])|(m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1500])|(~m[1428]&m[1429]&m[1430]&~m[1431]&~m[1500])|(m[1428]&m[1429]&m[1430]&~m[1431]&~m[1500])|(m[1428]&m[1429]&m[1430]&m[1431]&~m[1500])|(m[1428]&m[1429]&~m[1430]&~m[1431]&m[1500])|(m[1428]&~m[1429]&m[1430]&~m[1431]&m[1500])|(~m[1428]&m[1429]&m[1430]&~m[1431]&m[1500])|(m[1428]&m[1429]&m[1430]&~m[1431]&m[1500])|(m[1428]&m[1429]&m[1430]&m[1431]&m[1500]));
    m[1437] = (((m[1433]&~m[1434]&~m[1435]&~m[1436]&~m[1505])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1505])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1505])|(m[1433]&m[1434]&~m[1435]&m[1436]&~m[1505])|(m[1433]&~m[1434]&m[1435]&m[1436]&~m[1505])|(~m[1433]&m[1434]&m[1435]&m[1436]&~m[1505]))&BiasedRNG[996])|(((m[1433]&~m[1434]&~m[1435]&~m[1436]&m[1505])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&m[1505])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&m[1505])|(m[1433]&m[1434]&~m[1435]&m[1436]&m[1505])|(m[1433]&~m[1434]&m[1435]&m[1436]&m[1505])|(~m[1433]&m[1434]&m[1435]&m[1436]&m[1505]))&~BiasedRNG[996])|((m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1505])|(m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1505])|(~m[1433]&m[1434]&m[1435]&~m[1436]&~m[1505])|(m[1433]&m[1434]&m[1435]&~m[1436]&~m[1505])|(m[1433]&m[1434]&m[1435]&m[1436]&~m[1505])|(m[1433]&m[1434]&~m[1435]&~m[1436]&m[1505])|(m[1433]&~m[1434]&m[1435]&~m[1436]&m[1505])|(~m[1433]&m[1434]&m[1435]&~m[1436]&m[1505])|(m[1433]&m[1434]&m[1435]&~m[1436]&m[1505])|(m[1433]&m[1434]&m[1435]&m[1436]&m[1505]));
    m[1442] = (((m[1438]&~m[1439]&~m[1440]&~m[1441]&~m[1510])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1510])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1510])|(m[1438]&m[1439]&~m[1440]&m[1441]&~m[1510])|(m[1438]&~m[1439]&m[1440]&m[1441]&~m[1510])|(~m[1438]&m[1439]&m[1440]&m[1441]&~m[1510]))&BiasedRNG[997])|(((m[1438]&~m[1439]&~m[1440]&~m[1441]&m[1510])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&m[1510])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&m[1510])|(m[1438]&m[1439]&~m[1440]&m[1441]&m[1510])|(m[1438]&~m[1439]&m[1440]&m[1441]&m[1510])|(~m[1438]&m[1439]&m[1440]&m[1441]&m[1510]))&~BiasedRNG[997])|((m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1510])|(m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1510])|(~m[1438]&m[1439]&m[1440]&~m[1441]&~m[1510])|(m[1438]&m[1439]&m[1440]&~m[1441]&~m[1510])|(m[1438]&m[1439]&m[1440]&m[1441]&~m[1510])|(m[1438]&m[1439]&~m[1440]&~m[1441]&m[1510])|(m[1438]&~m[1439]&m[1440]&~m[1441]&m[1510])|(~m[1438]&m[1439]&m[1440]&~m[1441]&m[1510])|(m[1438]&m[1439]&m[1440]&~m[1441]&m[1510])|(m[1438]&m[1439]&m[1440]&m[1441]&m[1510]));
    m[1447] = (((m[1443]&~m[1444]&~m[1445]&~m[1446]&~m[1515])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1515])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1515])|(m[1443]&m[1444]&~m[1445]&m[1446]&~m[1515])|(m[1443]&~m[1444]&m[1445]&m[1446]&~m[1515])|(~m[1443]&m[1444]&m[1445]&m[1446]&~m[1515]))&BiasedRNG[998])|(((m[1443]&~m[1444]&~m[1445]&~m[1446]&m[1515])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&m[1515])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&m[1515])|(m[1443]&m[1444]&~m[1445]&m[1446]&m[1515])|(m[1443]&~m[1444]&m[1445]&m[1446]&m[1515])|(~m[1443]&m[1444]&m[1445]&m[1446]&m[1515]))&~BiasedRNG[998])|((m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1515])|(m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1515])|(~m[1443]&m[1444]&m[1445]&~m[1446]&~m[1515])|(m[1443]&m[1444]&m[1445]&~m[1446]&~m[1515])|(m[1443]&m[1444]&m[1445]&m[1446]&~m[1515])|(m[1443]&m[1444]&~m[1445]&~m[1446]&m[1515])|(m[1443]&~m[1444]&m[1445]&~m[1446]&m[1515])|(~m[1443]&m[1444]&m[1445]&~m[1446]&m[1515])|(m[1443]&m[1444]&m[1445]&~m[1446]&m[1515])|(m[1443]&m[1444]&m[1445]&m[1446]&m[1515]));
    m[1452] = (((m[1448]&~m[1449]&~m[1450]&~m[1451]&~m[1520])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1520])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1520])|(m[1448]&m[1449]&~m[1450]&m[1451]&~m[1520])|(m[1448]&~m[1449]&m[1450]&m[1451]&~m[1520])|(~m[1448]&m[1449]&m[1450]&m[1451]&~m[1520]))&BiasedRNG[999])|(((m[1448]&~m[1449]&~m[1450]&~m[1451]&m[1520])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&m[1520])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&m[1520])|(m[1448]&m[1449]&~m[1450]&m[1451]&m[1520])|(m[1448]&~m[1449]&m[1450]&m[1451]&m[1520])|(~m[1448]&m[1449]&m[1450]&m[1451]&m[1520]))&~BiasedRNG[999])|((m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1520])|(m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1520])|(~m[1448]&m[1449]&m[1450]&~m[1451]&~m[1520])|(m[1448]&m[1449]&m[1450]&~m[1451]&~m[1520])|(m[1448]&m[1449]&m[1450]&m[1451]&~m[1520])|(m[1448]&m[1449]&~m[1450]&~m[1451]&m[1520])|(m[1448]&~m[1449]&m[1450]&~m[1451]&m[1520])|(~m[1448]&m[1449]&m[1450]&~m[1451]&m[1520])|(m[1448]&m[1449]&m[1450]&~m[1451]&m[1520])|(m[1448]&m[1449]&m[1450]&m[1451]&m[1520]));
    m[1457] = (((m[1453]&~m[1454]&~m[1455]&~m[1456]&~m[1530])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1530])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1530])|(m[1453]&m[1454]&~m[1455]&m[1456]&~m[1530])|(m[1453]&~m[1454]&m[1455]&m[1456]&~m[1530])|(~m[1453]&m[1454]&m[1455]&m[1456]&~m[1530]))&BiasedRNG[1000])|(((m[1453]&~m[1454]&~m[1455]&~m[1456]&m[1530])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&m[1530])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&m[1530])|(m[1453]&m[1454]&~m[1455]&m[1456]&m[1530])|(m[1453]&~m[1454]&m[1455]&m[1456]&m[1530])|(~m[1453]&m[1454]&m[1455]&m[1456]&m[1530]))&~BiasedRNG[1000])|((m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1530])|(m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1530])|(~m[1453]&m[1454]&m[1455]&~m[1456]&~m[1530])|(m[1453]&m[1454]&m[1455]&~m[1456]&~m[1530])|(m[1453]&m[1454]&m[1455]&m[1456]&~m[1530])|(m[1453]&m[1454]&~m[1455]&~m[1456]&m[1530])|(m[1453]&~m[1454]&m[1455]&~m[1456]&m[1530])|(~m[1453]&m[1454]&m[1455]&~m[1456]&m[1530])|(m[1453]&m[1454]&m[1455]&~m[1456]&m[1530])|(m[1453]&m[1454]&m[1455]&m[1456]&m[1530]));
    m[1462] = (((m[1458]&~m[1459]&~m[1460]&~m[1461]&~m[1535])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1535])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1535])|(m[1458]&m[1459]&~m[1460]&m[1461]&~m[1535])|(m[1458]&~m[1459]&m[1460]&m[1461]&~m[1535])|(~m[1458]&m[1459]&m[1460]&m[1461]&~m[1535]))&BiasedRNG[1001])|(((m[1458]&~m[1459]&~m[1460]&~m[1461]&m[1535])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&m[1535])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&m[1535])|(m[1458]&m[1459]&~m[1460]&m[1461]&m[1535])|(m[1458]&~m[1459]&m[1460]&m[1461]&m[1535])|(~m[1458]&m[1459]&m[1460]&m[1461]&m[1535]))&~BiasedRNG[1001])|((m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1535])|(m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1535])|(~m[1458]&m[1459]&m[1460]&~m[1461]&~m[1535])|(m[1458]&m[1459]&m[1460]&~m[1461]&~m[1535])|(m[1458]&m[1459]&m[1460]&m[1461]&~m[1535])|(m[1458]&m[1459]&~m[1460]&~m[1461]&m[1535])|(m[1458]&~m[1459]&m[1460]&~m[1461]&m[1535])|(~m[1458]&m[1459]&m[1460]&~m[1461]&m[1535])|(m[1458]&m[1459]&m[1460]&~m[1461]&m[1535])|(m[1458]&m[1459]&m[1460]&m[1461]&m[1535]));
    m[1467] = (((m[1463]&~m[1464]&~m[1465]&~m[1466]&~m[1540])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1540])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1540])|(m[1463]&m[1464]&~m[1465]&m[1466]&~m[1540])|(m[1463]&~m[1464]&m[1465]&m[1466]&~m[1540])|(~m[1463]&m[1464]&m[1465]&m[1466]&~m[1540]))&BiasedRNG[1002])|(((m[1463]&~m[1464]&~m[1465]&~m[1466]&m[1540])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&m[1540])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&m[1540])|(m[1463]&m[1464]&~m[1465]&m[1466]&m[1540])|(m[1463]&~m[1464]&m[1465]&m[1466]&m[1540])|(~m[1463]&m[1464]&m[1465]&m[1466]&m[1540]))&~BiasedRNG[1002])|((m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1540])|(m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1540])|(~m[1463]&m[1464]&m[1465]&~m[1466]&~m[1540])|(m[1463]&m[1464]&m[1465]&~m[1466]&~m[1540])|(m[1463]&m[1464]&m[1465]&m[1466]&~m[1540])|(m[1463]&m[1464]&~m[1465]&~m[1466]&m[1540])|(m[1463]&~m[1464]&m[1465]&~m[1466]&m[1540])|(~m[1463]&m[1464]&m[1465]&~m[1466]&m[1540])|(m[1463]&m[1464]&m[1465]&~m[1466]&m[1540])|(m[1463]&m[1464]&m[1465]&m[1466]&m[1540]));
    m[1472] = (((m[1468]&~m[1469]&~m[1470]&~m[1471]&~m[1545])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1545])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1545])|(m[1468]&m[1469]&~m[1470]&m[1471]&~m[1545])|(m[1468]&~m[1469]&m[1470]&m[1471]&~m[1545])|(~m[1468]&m[1469]&m[1470]&m[1471]&~m[1545]))&BiasedRNG[1003])|(((m[1468]&~m[1469]&~m[1470]&~m[1471]&m[1545])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&m[1545])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&m[1545])|(m[1468]&m[1469]&~m[1470]&m[1471]&m[1545])|(m[1468]&~m[1469]&m[1470]&m[1471]&m[1545])|(~m[1468]&m[1469]&m[1470]&m[1471]&m[1545]))&~BiasedRNG[1003])|((m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1545])|(m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1545])|(~m[1468]&m[1469]&m[1470]&~m[1471]&~m[1545])|(m[1468]&m[1469]&m[1470]&~m[1471]&~m[1545])|(m[1468]&m[1469]&m[1470]&m[1471]&~m[1545])|(m[1468]&m[1469]&~m[1470]&~m[1471]&m[1545])|(m[1468]&~m[1469]&m[1470]&~m[1471]&m[1545])|(~m[1468]&m[1469]&m[1470]&~m[1471]&m[1545])|(m[1468]&m[1469]&m[1470]&~m[1471]&m[1545])|(m[1468]&m[1469]&m[1470]&m[1471]&m[1545]));
    m[1477] = (((m[1473]&~m[1474]&~m[1475]&~m[1476]&~m[1550])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1550])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1550])|(m[1473]&m[1474]&~m[1475]&m[1476]&~m[1550])|(m[1473]&~m[1474]&m[1475]&m[1476]&~m[1550])|(~m[1473]&m[1474]&m[1475]&m[1476]&~m[1550]))&BiasedRNG[1004])|(((m[1473]&~m[1474]&~m[1475]&~m[1476]&m[1550])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&m[1550])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&m[1550])|(m[1473]&m[1474]&~m[1475]&m[1476]&m[1550])|(m[1473]&~m[1474]&m[1475]&m[1476]&m[1550])|(~m[1473]&m[1474]&m[1475]&m[1476]&m[1550]))&~BiasedRNG[1004])|((m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1550])|(m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1550])|(~m[1473]&m[1474]&m[1475]&~m[1476]&~m[1550])|(m[1473]&m[1474]&m[1475]&~m[1476]&~m[1550])|(m[1473]&m[1474]&m[1475]&m[1476]&~m[1550])|(m[1473]&m[1474]&~m[1475]&~m[1476]&m[1550])|(m[1473]&~m[1474]&m[1475]&~m[1476]&m[1550])|(~m[1473]&m[1474]&m[1475]&~m[1476]&m[1550])|(m[1473]&m[1474]&m[1475]&~m[1476]&m[1550])|(m[1473]&m[1474]&m[1475]&m[1476]&m[1550]));
    m[1482] = (((m[1478]&~m[1479]&~m[1480]&~m[1481]&~m[1555])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1555])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1555])|(m[1478]&m[1479]&~m[1480]&m[1481]&~m[1555])|(m[1478]&~m[1479]&m[1480]&m[1481]&~m[1555])|(~m[1478]&m[1479]&m[1480]&m[1481]&~m[1555]))&BiasedRNG[1005])|(((m[1478]&~m[1479]&~m[1480]&~m[1481]&m[1555])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&m[1555])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&m[1555])|(m[1478]&m[1479]&~m[1480]&m[1481]&m[1555])|(m[1478]&~m[1479]&m[1480]&m[1481]&m[1555])|(~m[1478]&m[1479]&m[1480]&m[1481]&m[1555]))&~BiasedRNG[1005])|((m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1555])|(m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1555])|(~m[1478]&m[1479]&m[1480]&~m[1481]&~m[1555])|(m[1478]&m[1479]&m[1480]&~m[1481]&~m[1555])|(m[1478]&m[1479]&m[1480]&m[1481]&~m[1555])|(m[1478]&m[1479]&~m[1480]&~m[1481]&m[1555])|(m[1478]&~m[1479]&m[1480]&~m[1481]&m[1555])|(~m[1478]&m[1479]&m[1480]&~m[1481]&m[1555])|(m[1478]&m[1479]&m[1480]&~m[1481]&m[1555])|(m[1478]&m[1479]&m[1480]&m[1481]&m[1555]));
    m[1487] = (((m[1483]&~m[1484]&~m[1485]&~m[1486]&~m[1560])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1560])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1560])|(m[1483]&m[1484]&~m[1485]&m[1486]&~m[1560])|(m[1483]&~m[1484]&m[1485]&m[1486]&~m[1560])|(~m[1483]&m[1484]&m[1485]&m[1486]&~m[1560]))&BiasedRNG[1006])|(((m[1483]&~m[1484]&~m[1485]&~m[1486]&m[1560])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&m[1560])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&m[1560])|(m[1483]&m[1484]&~m[1485]&m[1486]&m[1560])|(m[1483]&~m[1484]&m[1485]&m[1486]&m[1560])|(~m[1483]&m[1484]&m[1485]&m[1486]&m[1560]))&~BiasedRNG[1006])|((m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1560])|(m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1560])|(~m[1483]&m[1484]&m[1485]&~m[1486]&~m[1560])|(m[1483]&m[1484]&m[1485]&~m[1486]&~m[1560])|(m[1483]&m[1484]&m[1485]&m[1486]&~m[1560])|(m[1483]&m[1484]&~m[1485]&~m[1486]&m[1560])|(m[1483]&~m[1484]&m[1485]&~m[1486]&m[1560])|(~m[1483]&m[1484]&m[1485]&~m[1486]&m[1560])|(m[1483]&m[1484]&m[1485]&~m[1486]&m[1560])|(m[1483]&m[1484]&m[1485]&m[1486]&m[1560]));
    m[1492] = (((m[1488]&~m[1489]&~m[1490]&~m[1491]&~m[1565])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1565])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1565])|(m[1488]&m[1489]&~m[1490]&m[1491]&~m[1565])|(m[1488]&~m[1489]&m[1490]&m[1491]&~m[1565])|(~m[1488]&m[1489]&m[1490]&m[1491]&~m[1565]))&BiasedRNG[1007])|(((m[1488]&~m[1489]&~m[1490]&~m[1491]&m[1565])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&m[1565])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&m[1565])|(m[1488]&m[1489]&~m[1490]&m[1491]&m[1565])|(m[1488]&~m[1489]&m[1490]&m[1491]&m[1565])|(~m[1488]&m[1489]&m[1490]&m[1491]&m[1565]))&~BiasedRNG[1007])|((m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1565])|(m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1565])|(~m[1488]&m[1489]&m[1490]&~m[1491]&~m[1565])|(m[1488]&m[1489]&m[1490]&~m[1491]&~m[1565])|(m[1488]&m[1489]&m[1490]&m[1491]&~m[1565])|(m[1488]&m[1489]&~m[1490]&~m[1491]&m[1565])|(m[1488]&~m[1489]&m[1490]&~m[1491]&m[1565])|(~m[1488]&m[1489]&m[1490]&~m[1491]&m[1565])|(m[1488]&m[1489]&m[1490]&~m[1491]&m[1565])|(m[1488]&m[1489]&m[1490]&m[1491]&m[1565]));
    m[1497] = (((m[1493]&~m[1494]&~m[1495]&~m[1496]&~m[1570])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1570])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1570])|(m[1493]&m[1494]&~m[1495]&m[1496]&~m[1570])|(m[1493]&~m[1494]&m[1495]&m[1496]&~m[1570])|(~m[1493]&m[1494]&m[1495]&m[1496]&~m[1570]))&BiasedRNG[1008])|(((m[1493]&~m[1494]&~m[1495]&~m[1496]&m[1570])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&m[1570])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&m[1570])|(m[1493]&m[1494]&~m[1495]&m[1496]&m[1570])|(m[1493]&~m[1494]&m[1495]&m[1496]&m[1570])|(~m[1493]&m[1494]&m[1495]&m[1496]&m[1570]))&~BiasedRNG[1008])|((m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1570])|(m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1570])|(~m[1493]&m[1494]&m[1495]&~m[1496]&~m[1570])|(m[1493]&m[1494]&m[1495]&~m[1496]&~m[1570])|(m[1493]&m[1494]&m[1495]&m[1496]&~m[1570])|(m[1493]&m[1494]&~m[1495]&~m[1496]&m[1570])|(m[1493]&~m[1494]&m[1495]&~m[1496]&m[1570])|(~m[1493]&m[1494]&m[1495]&~m[1496]&m[1570])|(m[1493]&m[1494]&m[1495]&~m[1496]&m[1570])|(m[1493]&m[1494]&m[1495]&m[1496]&m[1570]));
    m[1502] = (((m[1498]&~m[1499]&~m[1500]&~m[1501]&~m[1575])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1575])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1575])|(m[1498]&m[1499]&~m[1500]&m[1501]&~m[1575])|(m[1498]&~m[1499]&m[1500]&m[1501]&~m[1575])|(~m[1498]&m[1499]&m[1500]&m[1501]&~m[1575]))&BiasedRNG[1009])|(((m[1498]&~m[1499]&~m[1500]&~m[1501]&m[1575])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&m[1575])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&m[1575])|(m[1498]&m[1499]&~m[1500]&m[1501]&m[1575])|(m[1498]&~m[1499]&m[1500]&m[1501]&m[1575])|(~m[1498]&m[1499]&m[1500]&m[1501]&m[1575]))&~BiasedRNG[1009])|((m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1575])|(m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1575])|(~m[1498]&m[1499]&m[1500]&~m[1501]&~m[1575])|(m[1498]&m[1499]&m[1500]&~m[1501]&~m[1575])|(m[1498]&m[1499]&m[1500]&m[1501]&~m[1575])|(m[1498]&m[1499]&~m[1500]&~m[1501]&m[1575])|(m[1498]&~m[1499]&m[1500]&~m[1501]&m[1575])|(~m[1498]&m[1499]&m[1500]&~m[1501]&m[1575])|(m[1498]&m[1499]&m[1500]&~m[1501]&m[1575])|(m[1498]&m[1499]&m[1500]&m[1501]&m[1575]));
    m[1507] = (((m[1503]&~m[1504]&~m[1505]&~m[1506]&~m[1580])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1580])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1580])|(m[1503]&m[1504]&~m[1505]&m[1506]&~m[1580])|(m[1503]&~m[1504]&m[1505]&m[1506]&~m[1580])|(~m[1503]&m[1504]&m[1505]&m[1506]&~m[1580]))&BiasedRNG[1010])|(((m[1503]&~m[1504]&~m[1505]&~m[1506]&m[1580])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&m[1580])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&m[1580])|(m[1503]&m[1504]&~m[1505]&m[1506]&m[1580])|(m[1503]&~m[1504]&m[1505]&m[1506]&m[1580])|(~m[1503]&m[1504]&m[1505]&m[1506]&m[1580]))&~BiasedRNG[1010])|((m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1580])|(m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1580])|(~m[1503]&m[1504]&m[1505]&~m[1506]&~m[1580])|(m[1503]&m[1504]&m[1505]&~m[1506]&~m[1580])|(m[1503]&m[1504]&m[1505]&m[1506]&~m[1580])|(m[1503]&m[1504]&~m[1505]&~m[1506]&m[1580])|(m[1503]&~m[1504]&m[1505]&~m[1506]&m[1580])|(~m[1503]&m[1504]&m[1505]&~m[1506]&m[1580])|(m[1503]&m[1504]&m[1505]&~m[1506]&m[1580])|(m[1503]&m[1504]&m[1505]&m[1506]&m[1580]));
    m[1512] = (((m[1508]&~m[1509]&~m[1510]&~m[1511]&~m[1585])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1585])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1585])|(m[1508]&m[1509]&~m[1510]&m[1511]&~m[1585])|(m[1508]&~m[1509]&m[1510]&m[1511]&~m[1585])|(~m[1508]&m[1509]&m[1510]&m[1511]&~m[1585]))&BiasedRNG[1011])|(((m[1508]&~m[1509]&~m[1510]&~m[1511]&m[1585])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&m[1585])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&m[1585])|(m[1508]&m[1509]&~m[1510]&m[1511]&m[1585])|(m[1508]&~m[1509]&m[1510]&m[1511]&m[1585])|(~m[1508]&m[1509]&m[1510]&m[1511]&m[1585]))&~BiasedRNG[1011])|((m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1585])|(m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1585])|(~m[1508]&m[1509]&m[1510]&~m[1511]&~m[1585])|(m[1508]&m[1509]&m[1510]&~m[1511]&~m[1585])|(m[1508]&m[1509]&m[1510]&m[1511]&~m[1585])|(m[1508]&m[1509]&~m[1510]&~m[1511]&m[1585])|(m[1508]&~m[1509]&m[1510]&~m[1511]&m[1585])|(~m[1508]&m[1509]&m[1510]&~m[1511]&m[1585])|(m[1508]&m[1509]&m[1510]&~m[1511]&m[1585])|(m[1508]&m[1509]&m[1510]&m[1511]&m[1585]));
    m[1517] = (((m[1513]&~m[1514]&~m[1515]&~m[1516]&~m[1590])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1590])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1590])|(m[1513]&m[1514]&~m[1515]&m[1516]&~m[1590])|(m[1513]&~m[1514]&m[1515]&m[1516]&~m[1590])|(~m[1513]&m[1514]&m[1515]&m[1516]&~m[1590]))&BiasedRNG[1012])|(((m[1513]&~m[1514]&~m[1515]&~m[1516]&m[1590])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&m[1590])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&m[1590])|(m[1513]&m[1514]&~m[1515]&m[1516]&m[1590])|(m[1513]&~m[1514]&m[1515]&m[1516]&m[1590])|(~m[1513]&m[1514]&m[1515]&m[1516]&m[1590]))&~BiasedRNG[1012])|((m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1590])|(m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1590])|(~m[1513]&m[1514]&m[1515]&~m[1516]&~m[1590])|(m[1513]&m[1514]&m[1515]&~m[1516]&~m[1590])|(m[1513]&m[1514]&m[1515]&m[1516]&~m[1590])|(m[1513]&m[1514]&~m[1515]&~m[1516]&m[1590])|(m[1513]&~m[1514]&m[1515]&~m[1516]&m[1590])|(~m[1513]&m[1514]&m[1515]&~m[1516]&m[1590])|(m[1513]&m[1514]&m[1515]&~m[1516]&m[1590])|(m[1513]&m[1514]&m[1515]&m[1516]&m[1590]));
    m[1522] = (((m[1518]&~m[1519]&~m[1520]&~m[1521]&~m[1595])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1595])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1595])|(m[1518]&m[1519]&~m[1520]&m[1521]&~m[1595])|(m[1518]&~m[1519]&m[1520]&m[1521]&~m[1595])|(~m[1518]&m[1519]&m[1520]&m[1521]&~m[1595]))&BiasedRNG[1013])|(((m[1518]&~m[1519]&~m[1520]&~m[1521]&m[1595])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&m[1595])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&m[1595])|(m[1518]&m[1519]&~m[1520]&m[1521]&m[1595])|(m[1518]&~m[1519]&m[1520]&m[1521]&m[1595])|(~m[1518]&m[1519]&m[1520]&m[1521]&m[1595]))&~BiasedRNG[1013])|((m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1595])|(m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1595])|(~m[1518]&m[1519]&m[1520]&~m[1521]&~m[1595])|(m[1518]&m[1519]&m[1520]&~m[1521]&~m[1595])|(m[1518]&m[1519]&m[1520]&m[1521]&~m[1595])|(m[1518]&m[1519]&~m[1520]&~m[1521]&m[1595])|(m[1518]&~m[1519]&m[1520]&~m[1521]&m[1595])|(~m[1518]&m[1519]&m[1520]&~m[1521]&m[1595])|(m[1518]&m[1519]&m[1520]&~m[1521]&m[1595])|(m[1518]&m[1519]&m[1520]&m[1521]&m[1595]));
    m[1527] = (((m[1523]&~m[1524]&~m[1525]&~m[1526]&~m[1600])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1600])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1600])|(m[1523]&m[1524]&~m[1525]&m[1526]&~m[1600])|(m[1523]&~m[1524]&m[1525]&m[1526]&~m[1600])|(~m[1523]&m[1524]&m[1525]&m[1526]&~m[1600]))&BiasedRNG[1014])|(((m[1523]&~m[1524]&~m[1525]&~m[1526]&m[1600])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&m[1600])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&m[1600])|(m[1523]&m[1524]&~m[1525]&m[1526]&m[1600])|(m[1523]&~m[1524]&m[1525]&m[1526]&m[1600])|(~m[1523]&m[1524]&m[1525]&m[1526]&m[1600]))&~BiasedRNG[1014])|((m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1600])|(m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1600])|(~m[1523]&m[1524]&m[1525]&~m[1526]&~m[1600])|(m[1523]&m[1524]&m[1525]&~m[1526]&~m[1600])|(m[1523]&m[1524]&m[1525]&m[1526]&~m[1600])|(m[1523]&m[1524]&~m[1525]&~m[1526]&m[1600])|(m[1523]&~m[1524]&m[1525]&~m[1526]&m[1600])|(~m[1523]&m[1524]&m[1525]&~m[1526]&m[1600])|(m[1523]&m[1524]&m[1525]&~m[1526]&m[1600])|(m[1523]&m[1524]&m[1525]&m[1526]&m[1600]));
    m[1532] = (((m[1528]&~m[1529]&~m[1530]&~m[1531]&~m[1603])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1603])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1603])|(m[1528]&m[1529]&~m[1530]&m[1531]&~m[1603])|(m[1528]&~m[1529]&m[1530]&m[1531]&~m[1603])|(~m[1528]&m[1529]&m[1530]&m[1531]&~m[1603]))&BiasedRNG[1015])|(((m[1528]&~m[1529]&~m[1530]&~m[1531]&m[1603])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&m[1603])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&m[1603])|(m[1528]&m[1529]&~m[1530]&m[1531]&m[1603])|(m[1528]&~m[1529]&m[1530]&m[1531]&m[1603])|(~m[1528]&m[1529]&m[1530]&m[1531]&m[1603]))&~BiasedRNG[1015])|((m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1603])|(m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1603])|(~m[1528]&m[1529]&m[1530]&~m[1531]&~m[1603])|(m[1528]&m[1529]&m[1530]&~m[1531]&~m[1603])|(m[1528]&m[1529]&m[1530]&m[1531]&~m[1603])|(m[1528]&m[1529]&~m[1530]&~m[1531]&m[1603])|(m[1528]&~m[1529]&m[1530]&~m[1531]&m[1603])|(~m[1528]&m[1529]&m[1530]&~m[1531]&m[1603])|(m[1528]&m[1529]&m[1530]&~m[1531]&m[1603])|(m[1528]&m[1529]&m[1530]&m[1531]&m[1603]));
    m[1537] = (((m[1533]&~m[1534]&~m[1535]&~m[1536]&~m[1605])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1605])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1605])|(m[1533]&m[1534]&~m[1535]&m[1536]&~m[1605])|(m[1533]&~m[1534]&m[1535]&m[1536]&~m[1605])|(~m[1533]&m[1534]&m[1535]&m[1536]&~m[1605]))&BiasedRNG[1016])|(((m[1533]&~m[1534]&~m[1535]&~m[1536]&m[1605])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&m[1605])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&m[1605])|(m[1533]&m[1534]&~m[1535]&m[1536]&m[1605])|(m[1533]&~m[1534]&m[1535]&m[1536]&m[1605])|(~m[1533]&m[1534]&m[1535]&m[1536]&m[1605]))&~BiasedRNG[1016])|((m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1605])|(m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1605])|(~m[1533]&m[1534]&m[1535]&~m[1536]&~m[1605])|(m[1533]&m[1534]&m[1535]&~m[1536]&~m[1605])|(m[1533]&m[1534]&m[1535]&m[1536]&~m[1605])|(m[1533]&m[1534]&~m[1535]&~m[1536]&m[1605])|(m[1533]&~m[1534]&m[1535]&~m[1536]&m[1605])|(~m[1533]&m[1534]&m[1535]&~m[1536]&m[1605])|(m[1533]&m[1534]&m[1535]&~m[1536]&m[1605])|(m[1533]&m[1534]&m[1535]&m[1536]&m[1605]));
    m[1542] = (((m[1538]&~m[1539]&~m[1540]&~m[1541]&~m[1610])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1610])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1610])|(m[1538]&m[1539]&~m[1540]&m[1541]&~m[1610])|(m[1538]&~m[1539]&m[1540]&m[1541]&~m[1610])|(~m[1538]&m[1539]&m[1540]&m[1541]&~m[1610]))&BiasedRNG[1017])|(((m[1538]&~m[1539]&~m[1540]&~m[1541]&m[1610])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&m[1610])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&m[1610])|(m[1538]&m[1539]&~m[1540]&m[1541]&m[1610])|(m[1538]&~m[1539]&m[1540]&m[1541]&m[1610])|(~m[1538]&m[1539]&m[1540]&m[1541]&m[1610]))&~BiasedRNG[1017])|((m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1610])|(m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1610])|(~m[1538]&m[1539]&m[1540]&~m[1541]&~m[1610])|(m[1538]&m[1539]&m[1540]&~m[1541]&~m[1610])|(m[1538]&m[1539]&m[1540]&m[1541]&~m[1610])|(m[1538]&m[1539]&~m[1540]&~m[1541]&m[1610])|(m[1538]&~m[1539]&m[1540]&~m[1541]&m[1610])|(~m[1538]&m[1539]&m[1540]&~m[1541]&m[1610])|(m[1538]&m[1539]&m[1540]&~m[1541]&m[1610])|(m[1538]&m[1539]&m[1540]&m[1541]&m[1610]));
    m[1547] = (((m[1543]&~m[1544]&~m[1545]&~m[1546]&~m[1615])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1615])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1615])|(m[1543]&m[1544]&~m[1545]&m[1546]&~m[1615])|(m[1543]&~m[1544]&m[1545]&m[1546]&~m[1615])|(~m[1543]&m[1544]&m[1545]&m[1546]&~m[1615]))&BiasedRNG[1018])|(((m[1543]&~m[1544]&~m[1545]&~m[1546]&m[1615])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&m[1615])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&m[1615])|(m[1543]&m[1544]&~m[1545]&m[1546]&m[1615])|(m[1543]&~m[1544]&m[1545]&m[1546]&m[1615])|(~m[1543]&m[1544]&m[1545]&m[1546]&m[1615]))&~BiasedRNG[1018])|((m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1615])|(m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1615])|(~m[1543]&m[1544]&m[1545]&~m[1546]&~m[1615])|(m[1543]&m[1544]&m[1545]&~m[1546]&~m[1615])|(m[1543]&m[1544]&m[1545]&m[1546]&~m[1615])|(m[1543]&m[1544]&~m[1545]&~m[1546]&m[1615])|(m[1543]&~m[1544]&m[1545]&~m[1546]&m[1615])|(~m[1543]&m[1544]&m[1545]&~m[1546]&m[1615])|(m[1543]&m[1544]&m[1545]&~m[1546]&m[1615])|(m[1543]&m[1544]&m[1545]&m[1546]&m[1615]));
    m[1552] = (((m[1548]&~m[1549]&~m[1550]&~m[1551]&~m[1620])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1620])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1620])|(m[1548]&m[1549]&~m[1550]&m[1551]&~m[1620])|(m[1548]&~m[1549]&m[1550]&m[1551]&~m[1620])|(~m[1548]&m[1549]&m[1550]&m[1551]&~m[1620]))&BiasedRNG[1019])|(((m[1548]&~m[1549]&~m[1550]&~m[1551]&m[1620])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&m[1620])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&m[1620])|(m[1548]&m[1549]&~m[1550]&m[1551]&m[1620])|(m[1548]&~m[1549]&m[1550]&m[1551]&m[1620])|(~m[1548]&m[1549]&m[1550]&m[1551]&m[1620]))&~BiasedRNG[1019])|((m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1620])|(m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1620])|(~m[1548]&m[1549]&m[1550]&~m[1551]&~m[1620])|(m[1548]&m[1549]&m[1550]&~m[1551]&~m[1620])|(m[1548]&m[1549]&m[1550]&m[1551]&~m[1620])|(m[1548]&m[1549]&~m[1550]&~m[1551]&m[1620])|(m[1548]&~m[1549]&m[1550]&~m[1551]&m[1620])|(~m[1548]&m[1549]&m[1550]&~m[1551]&m[1620])|(m[1548]&m[1549]&m[1550]&~m[1551]&m[1620])|(m[1548]&m[1549]&m[1550]&m[1551]&m[1620]));
    m[1557] = (((m[1553]&~m[1554]&~m[1555]&~m[1556]&~m[1625])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1625])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1625])|(m[1553]&m[1554]&~m[1555]&m[1556]&~m[1625])|(m[1553]&~m[1554]&m[1555]&m[1556]&~m[1625])|(~m[1553]&m[1554]&m[1555]&m[1556]&~m[1625]))&BiasedRNG[1020])|(((m[1553]&~m[1554]&~m[1555]&~m[1556]&m[1625])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&m[1625])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&m[1625])|(m[1553]&m[1554]&~m[1555]&m[1556]&m[1625])|(m[1553]&~m[1554]&m[1555]&m[1556]&m[1625])|(~m[1553]&m[1554]&m[1555]&m[1556]&m[1625]))&~BiasedRNG[1020])|((m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1625])|(m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1625])|(~m[1553]&m[1554]&m[1555]&~m[1556]&~m[1625])|(m[1553]&m[1554]&m[1555]&~m[1556]&~m[1625])|(m[1553]&m[1554]&m[1555]&m[1556]&~m[1625])|(m[1553]&m[1554]&~m[1555]&~m[1556]&m[1625])|(m[1553]&~m[1554]&m[1555]&~m[1556]&m[1625])|(~m[1553]&m[1554]&m[1555]&~m[1556]&m[1625])|(m[1553]&m[1554]&m[1555]&~m[1556]&m[1625])|(m[1553]&m[1554]&m[1555]&m[1556]&m[1625]));
    m[1562] = (((m[1558]&~m[1559]&~m[1560]&~m[1561]&~m[1630])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1630])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1630])|(m[1558]&m[1559]&~m[1560]&m[1561]&~m[1630])|(m[1558]&~m[1559]&m[1560]&m[1561]&~m[1630])|(~m[1558]&m[1559]&m[1560]&m[1561]&~m[1630]))&BiasedRNG[1021])|(((m[1558]&~m[1559]&~m[1560]&~m[1561]&m[1630])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&m[1630])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&m[1630])|(m[1558]&m[1559]&~m[1560]&m[1561]&m[1630])|(m[1558]&~m[1559]&m[1560]&m[1561]&m[1630])|(~m[1558]&m[1559]&m[1560]&m[1561]&m[1630]))&~BiasedRNG[1021])|((m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1630])|(m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1630])|(~m[1558]&m[1559]&m[1560]&~m[1561]&~m[1630])|(m[1558]&m[1559]&m[1560]&~m[1561]&~m[1630])|(m[1558]&m[1559]&m[1560]&m[1561]&~m[1630])|(m[1558]&m[1559]&~m[1560]&~m[1561]&m[1630])|(m[1558]&~m[1559]&m[1560]&~m[1561]&m[1630])|(~m[1558]&m[1559]&m[1560]&~m[1561]&m[1630])|(m[1558]&m[1559]&m[1560]&~m[1561]&m[1630])|(m[1558]&m[1559]&m[1560]&m[1561]&m[1630]));
    m[1567] = (((m[1563]&~m[1564]&~m[1565]&~m[1566]&~m[1635])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1635])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1635])|(m[1563]&m[1564]&~m[1565]&m[1566]&~m[1635])|(m[1563]&~m[1564]&m[1565]&m[1566]&~m[1635])|(~m[1563]&m[1564]&m[1565]&m[1566]&~m[1635]))&BiasedRNG[1022])|(((m[1563]&~m[1564]&~m[1565]&~m[1566]&m[1635])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&m[1635])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&m[1635])|(m[1563]&m[1564]&~m[1565]&m[1566]&m[1635])|(m[1563]&~m[1564]&m[1565]&m[1566]&m[1635])|(~m[1563]&m[1564]&m[1565]&m[1566]&m[1635]))&~BiasedRNG[1022])|((m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1635])|(m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1635])|(~m[1563]&m[1564]&m[1565]&~m[1566]&~m[1635])|(m[1563]&m[1564]&m[1565]&~m[1566]&~m[1635])|(m[1563]&m[1564]&m[1565]&m[1566]&~m[1635])|(m[1563]&m[1564]&~m[1565]&~m[1566]&m[1635])|(m[1563]&~m[1564]&m[1565]&~m[1566]&m[1635])|(~m[1563]&m[1564]&m[1565]&~m[1566]&m[1635])|(m[1563]&m[1564]&m[1565]&~m[1566]&m[1635])|(m[1563]&m[1564]&m[1565]&m[1566]&m[1635]));
    m[1572] = (((m[1568]&~m[1569]&~m[1570]&~m[1571]&~m[1640])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1640])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1640])|(m[1568]&m[1569]&~m[1570]&m[1571]&~m[1640])|(m[1568]&~m[1569]&m[1570]&m[1571]&~m[1640])|(~m[1568]&m[1569]&m[1570]&m[1571]&~m[1640]))&BiasedRNG[1023])|(((m[1568]&~m[1569]&~m[1570]&~m[1571]&m[1640])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&m[1640])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&m[1640])|(m[1568]&m[1569]&~m[1570]&m[1571]&m[1640])|(m[1568]&~m[1569]&m[1570]&m[1571]&m[1640])|(~m[1568]&m[1569]&m[1570]&m[1571]&m[1640]))&~BiasedRNG[1023])|((m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1640])|(m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1640])|(~m[1568]&m[1569]&m[1570]&~m[1571]&~m[1640])|(m[1568]&m[1569]&m[1570]&~m[1571]&~m[1640])|(m[1568]&m[1569]&m[1570]&m[1571]&~m[1640])|(m[1568]&m[1569]&~m[1570]&~m[1571]&m[1640])|(m[1568]&~m[1569]&m[1570]&~m[1571]&m[1640])|(~m[1568]&m[1569]&m[1570]&~m[1571]&m[1640])|(m[1568]&m[1569]&m[1570]&~m[1571]&m[1640])|(m[1568]&m[1569]&m[1570]&m[1571]&m[1640]));
    m[1577] = (((m[1573]&~m[1574]&~m[1575]&~m[1576]&~m[1645])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1645])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1645])|(m[1573]&m[1574]&~m[1575]&m[1576]&~m[1645])|(m[1573]&~m[1574]&m[1575]&m[1576]&~m[1645])|(~m[1573]&m[1574]&m[1575]&m[1576]&~m[1645]))&BiasedRNG[1024])|(((m[1573]&~m[1574]&~m[1575]&~m[1576]&m[1645])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&m[1645])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&m[1645])|(m[1573]&m[1574]&~m[1575]&m[1576]&m[1645])|(m[1573]&~m[1574]&m[1575]&m[1576]&m[1645])|(~m[1573]&m[1574]&m[1575]&m[1576]&m[1645]))&~BiasedRNG[1024])|((m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1645])|(m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1645])|(~m[1573]&m[1574]&m[1575]&~m[1576]&~m[1645])|(m[1573]&m[1574]&m[1575]&~m[1576]&~m[1645])|(m[1573]&m[1574]&m[1575]&m[1576]&~m[1645])|(m[1573]&m[1574]&~m[1575]&~m[1576]&m[1645])|(m[1573]&~m[1574]&m[1575]&~m[1576]&m[1645])|(~m[1573]&m[1574]&m[1575]&~m[1576]&m[1645])|(m[1573]&m[1574]&m[1575]&~m[1576]&m[1645])|(m[1573]&m[1574]&m[1575]&m[1576]&m[1645]));
    m[1582] = (((m[1578]&~m[1579]&~m[1580]&~m[1581]&~m[1650])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1650])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1650])|(m[1578]&m[1579]&~m[1580]&m[1581]&~m[1650])|(m[1578]&~m[1579]&m[1580]&m[1581]&~m[1650])|(~m[1578]&m[1579]&m[1580]&m[1581]&~m[1650]))&BiasedRNG[1025])|(((m[1578]&~m[1579]&~m[1580]&~m[1581]&m[1650])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&m[1650])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&m[1650])|(m[1578]&m[1579]&~m[1580]&m[1581]&m[1650])|(m[1578]&~m[1579]&m[1580]&m[1581]&m[1650])|(~m[1578]&m[1579]&m[1580]&m[1581]&m[1650]))&~BiasedRNG[1025])|((m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1650])|(m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1650])|(~m[1578]&m[1579]&m[1580]&~m[1581]&~m[1650])|(m[1578]&m[1579]&m[1580]&~m[1581]&~m[1650])|(m[1578]&m[1579]&m[1580]&m[1581]&~m[1650])|(m[1578]&m[1579]&~m[1580]&~m[1581]&m[1650])|(m[1578]&~m[1579]&m[1580]&~m[1581]&m[1650])|(~m[1578]&m[1579]&m[1580]&~m[1581]&m[1650])|(m[1578]&m[1579]&m[1580]&~m[1581]&m[1650])|(m[1578]&m[1579]&m[1580]&m[1581]&m[1650]));
    m[1587] = (((m[1583]&~m[1584]&~m[1585]&~m[1586]&~m[1655])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1655])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1655])|(m[1583]&m[1584]&~m[1585]&m[1586]&~m[1655])|(m[1583]&~m[1584]&m[1585]&m[1586]&~m[1655])|(~m[1583]&m[1584]&m[1585]&m[1586]&~m[1655]))&BiasedRNG[1026])|(((m[1583]&~m[1584]&~m[1585]&~m[1586]&m[1655])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&m[1655])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&m[1655])|(m[1583]&m[1584]&~m[1585]&m[1586]&m[1655])|(m[1583]&~m[1584]&m[1585]&m[1586]&m[1655])|(~m[1583]&m[1584]&m[1585]&m[1586]&m[1655]))&~BiasedRNG[1026])|((m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1655])|(m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1655])|(~m[1583]&m[1584]&m[1585]&~m[1586]&~m[1655])|(m[1583]&m[1584]&m[1585]&~m[1586]&~m[1655])|(m[1583]&m[1584]&m[1585]&m[1586]&~m[1655])|(m[1583]&m[1584]&~m[1585]&~m[1586]&m[1655])|(m[1583]&~m[1584]&m[1585]&~m[1586]&m[1655])|(~m[1583]&m[1584]&m[1585]&~m[1586]&m[1655])|(m[1583]&m[1584]&m[1585]&~m[1586]&m[1655])|(m[1583]&m[1584]&m[1585]&m[1586]&m[1655]));
    m[1592] = (((m[1588]&~m[1589]&~m[1590]&~m[1591]&~m[1660])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1660])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1660])|(m[1588]&m[1589]&~m[1590]&m[1591]&~m[1660])|(m[1588]&~m[1589]&m[1590]&m[1591]&~m[1660])|(~m[1588]&m[1589]&m[1590]&m[1591]&~m[1660]))&BiasedRNG[1027])|(((m[1588]&~m[1589]&~m[1590]&~m[1591]&m[1660])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&m[1660])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&m[1660])|(m[1588]&m[1589]&~m[1590]&m[1591]&m[1660])|(m[1588]&~m[1589]&m[1590]&m[1591]&m[1660])|(~m[1588]&m[1589]&m[1590]&m[1591]&m[1660]))&~BiasedRNG[1027])|((m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1660])|(m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1660])|(~m[1588]&m[1589]&m[1590]&~m[1591]&~m[1660])|(m[1588]&m[1589]&m[1590]&~m[1591]&~m[1660])|(m[1588]&m[1589]&m[1590]&m[1591]&~m[1660])|(m[1588]&m[1589]&~m[1590]&~m[1591]&m[1660])|(m[1588]&~m[1589]&m[1590]&~m[1591]&m[1660])|(~m[1588]&m[1589]&m[1590]&~m[1591]&m[1660])|(m[1588]&m[1589]&m[1590]&~m[1591]&m[1660])|(m[1588]&m[1589]&m[1590]&m[1591]&m[1660]));
    m[1597] = (((m[1593]&~m[1594]&~m[1595]&~m[1596]&~m[1665])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1665])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1665])|(m[1593]&m[1594]&~m[1595]&m[1596]&~m[1665])|(m[1593]&~m[1594]&m[1595]&m[1596]&~m[1665])|(~m[1593]&m[1594]&m[1595]&m[1596]&~m[1665]))&BiasedRNG[1028])|(((m[1593]&~m[1594]&~m[1595]&~m[1596]&m[1665])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&m[1665])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&m[1665])|(m[1593]&m[1594]&~m[1595]&m[1596]&m[1665])|(m[1593]&~m[1594]&m[1595]&m[1596]&m[1665])|(~m[1593]&m[1594]&m[1595]&m[1596]&m[1665]))&~BiasedRNG[1028])|((m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1665])|(m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1665])|(~m[1593]&m[1594]&m[1595]&~m[1596]&~m[1665])|(m[1593]&m[1594]&m[1595]&~m[1596]&~m[1665])|(m[1593]&m[1594]&m[1595]&m[1596]&~m[1665])|(m[1593]&m[1594]&~m[1595]&~m[1596]&m[1665])|(m[1593]&~m[1594]&m[1595]&~m[1596]&m[1665])|(~m[1593]&m[1594]&m[1595]&~m[1596]&m[1665])|(m[1593]&m[1594]&m[1595]&~m[1596]&m[1665])|(m[1593]&m[1594]&m[1595]&m[1596]&m[1665]));
    m[1602] = (((m[1598]&~m[1599]&~m[1600]&~m[1601]&~m[1670])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1670])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1670])|(m[1598]&m[1599]&~m[1600]&m[1601]&~m[1670])|(m[1598]&~m[1599]&m[1600]&m[1601]&~m[1670])|(~m[1598]&m[1599]&m[1600]&m[1601]&~m[1670]))&BiasedRNG[1029])|(((m[1598]&~m[1599]&~m[1600]&~m[1601]&m[1670])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&m[1670])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&m[1670])|(m[1598]&m[1599]&~m[1600]&m[1601]&m[1670])|(m[1598]&~m[1599]&m[1600]&m[1601]&m[1670])|(~m[1598]&m[1599]&m[1600]&m[1601]&m[1670]))&~BiasedRNG[1029])|((m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1670])|(m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1670])|(~m[1598]&m[1599]&m[1600]&~m[1601]&~m[1670])|(m[1598]&m[1599]&m[1600]&~m[1601]&~m[1670])|(m[1598]&m[1599]&m[1600]&m[1601]&~m[1670])|(m[1598]&m[1599]&~m[1600]&~m[1601]&m[1670])|(m[1598]&~m[1599]&m[1600]&~m[1601]&m[1670])|(~m[1598]&m[1599]&m[1600]&~m[1601]&m[1670])|(m[1598]&m[1599]&m[1600]&~m[1601]&m[1670])|(m[1598]&m[1599]&m[1600]&m[1601]&m[1670]));
    m[1607] = (((m[1603]&~m[1604]&~m[1605]&~m[1606]&~m[1673])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1673])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1673])|(m[1603]&m[1604]&~m[1605]&m[1606]&~m[1673])|(m[1603]&~m[1604]&m[1605]&m[1606]&~m[1673])|(~m[1603]&m[1604]&m[1605]&m[1606]&~m[1673]))&BiasedRNG[1030])|(((m[1603]&~m[1604]&~m[1605]&~m[1606]&m[1673])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&m[1673])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&m[1673])|(m[1603]&m[1604]&~m[1605]&m[1606]&m[1673])|(m[1603]&~m[1604]&m[1605]&m[1606]&m[1673])|(~m[1603]&m[1604]&m[1605]&m[1606]&m[1673]))&~BiasedRNG[1030])|((m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1673])|(m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1673])|(~m[1603]&m[1604]&m[1605]&~m[1606]&~m[1673])|(m[1603]&m[1604]&m[1605]&~m[1606]&~m[1673])|(m[1603]&m[1604]&m[1605]&m[1606]&~m[1673])|(m[1603]&m[1604]&~m[1605]&~m[1606]&m[1673])|(m[1603]&~m[1604]&m[1605]&~m[1606]&m[1673])|(~m[1603]&m[1604]&m[1605]&~m[1606]&m[1673])|(m[1603]&m[1604]&m[1605]&~m[1606]&m[1673])|(m[1603]&m[1604]&m[1605]&m[1606]&m[1673]));
    m[1612] = (((m[1608]&~m[1609]&~m[1610]&~m[1611]&~m[1675])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1675])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1675])|(m[1608]&m[1609]&~m[1610]&m[1611]&~m[1675])|(m[1608]&~m[1609]&m[1610]&m[1611]&~m[1675])|(~m[1608]&m[1609]&m[1610]&m[1611]&~m[1675]))&BiasedRNG[1031])|(((m[1608]&~m[1609]&~m[1610]&~m[1611]&m[1675])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&m[1675])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&m[1675])|(m[1608]&m[1609]&~m[1610]&m[1611]&m[1675])|(m[1608]&~m[1609]&m[1610]&m[1611]&m[1675])|(~m[1608]&m[1609]&m[1610]&m[1611]&m[1675]))&~BiasedRNG[1031])|((m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1675])|(m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1675])|(~m[1608]&m[1609]&m[1610]&~m[1611]&~m[1675])|(m[1608]&m[1609]&m[1610]&~m[1611]&~m[1675])|(m[1608]&m[1609]&m[1610]&m[1611]&~m[1675])|(m[1608]&m[1609]&~m[1610]&~m[1611]&m[1675])|(m[1608]&~m[1609]&m[1610]&~m[1611]&m[1675])|(~m[1608]&m[1609]&m[1610]&~m[1611]&m[1675])|(m[1608]&m[1609]&m[1610]&~m[1611]&m[1675])|(m[1608]&m[1609]&m[1610]&m[1611]&m[1675]));
    m[1617] = (((m[1613]&~m[1614]&~m[1615]&~m[1616]&~m[1680])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1680])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1680])|(m[1613]&m[1614]&~m[1615]&m[1616]&~m[1680])|(m[1613]&~m[1614]&m[1615]&m[1616]&~m[1680])|(~m[1613]&m[1614]&m[1615]&m[1616]&~m[1680]))&BiasedRNG[1032])|(((m[1613]&~m[1614]&~m[1615]&~m[1616]&m[1680])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&m[1680])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&m[1680])|(m[1613]&m[1614]&~m[1615]&m[1616]&m[1680])|(m[1613]&~m[1614]&m[1615]&m[1616]&m[1680])|(~m[1613]&m[1614]&m[1615]&m[1616]&m[1680]))&~BiasedRNG[1032])|((m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1680])|(m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1680])|(~m[1613]&m[1614]&m[1615]&~m[1616]&~m[1680])|(m[1613]&m[1614]&m[1615]&~m[1616]&~m[1680])|(m[1613]&m[1614]&m[1615]&m[1616]&~m[1680])|(m[1613]&m[1614]&~m[1615]&~m[1616]&m[1680])|(m[1613]&~m[1614]&m[1615]&~m[1616]&m[1680])|(~m[1613]&m[1614]&m[1615]&~m[1616]&m[1680])|(m[1613]&m[1614]&m[1615]&~m[1616]&m[1680])|(m[1613]&m[1614]&m[1615]&m[1616]&m[1680]));
    m[1622] = (((m[1618]&~m[1619]&~m[1620]&~m[1621]&~m[1685])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1685])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1685])|(m[1618]&m[1619]&~m[1620]&m[1621]&~m[1685])|(m[1618]&~m[1619]&m[1620]&m[1621]&~m[1685])|(~m[1618]&m[1619]&m[1620]&m[1621]&~m[1685]))&BiasedRNG[1033])|(((m[1618]&~m[1619]&~m[1620]&~m[1621]&m[1685])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&m[1685])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&m[1685])|(m[1618]&m[1619]&~m[1620]&m[1621]&m[1685])|(m[1618]&~m[1619]&m[1620]&m[1621]&m[1685])|(~m[1618]&m[1619]&m[1620]&m[1621]&m[1685]))&~BiasedRNG[1033])|((m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1685])|(m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1685])|(~m[1618]&m[1619]&m[1620]&~m[1621]&~m[1685])|(m[1618]&m[1619]&m[1620]&~m[1621]&~m[1685])|(m[1618]&m[1619]&m[1620]&m[1621]&~m[1685])|(m[1618]&m[1619]&~m[1620]&~m[1621]&m[1685])|(m[1618]&~m[1619]&m[1620]&~m[1621]&m[1685])|(~m[1618]&m[1619]&m[1620]&~m[1621]&m[1685])|(m[1618]&m[1619]&m[1620]&~m[1621]&m[1685])|(m[1618]&m[1619]&m[1620]&m[1621]&m[1685]));
    m[1627] = (((m[1623]&~m[1624]&~m[1625]&~m[1626]&~m[1690])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1690])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1690])|(m[1623]&m[1624]&~m[1625]&m[1626]&~m[1690])|(m[1623]&~m[1624]&m[1625]&m[1626]&~m[1690])|(~m[1623]&m[1624]&m[1625]&m[1626]&~m[1690]))&BiasedRNG[1034])|(((m[1623]&~m[1624]&~m[1625]&~m[1626]&m[1690])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&m[1690])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&m[1690])|(m[1623]&m[1624]&~m[1625]&m[1626]&m[1690])|(m[1623]&~m[1624]&m[1625]&m[1626]&m[1690])|(~m[1623]&m[1624]&m[1625]&m[1626]&m[1690]))&~BiasedRNG[1034])|((m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1690])|(m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1690])|(~m[1623]&m[1624]&m[1625]&~m[1626]&~m[1690])|(m[1623]&m[1624]&m[1625]&~m[1626]&~m[1690])|(m[1623]&m[1624]&m[1625]&m[1626]&~m[1690])|(m[1623]&m[1624]&~m[1625]&~m[1626]&m[1690])|(m[1623]&~m[1624]&m[1625]&~m[1626]&m[1690])|(~m[1623]&m[1624]&m[1625]&~m[1626]&m[1690])|(m[1623]&m[1624]&m[1625]&~m[1626]&m[1690])|(m[1623]&m[1624]&m[1625]&m[1626]&m[1690]));
    m[1632] = (((m[1628]&~m[1629]&~m[1630]&~m[1631]&~m[1695])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1695])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1695])|(m[1628]&m[1629]&~m[1630]&m[1631]&~m[1695])|(m[1628]&~m[1629]&m[1630]&m[1631]&~m[1695])|(~m[1628]&m[1629]&m[1630]&m[1631]&~m[1695]))&BiasedRNG[1035])|(((m[1628]&~m[1629]&~m[1630]&~m[1631]&m[1695])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&m[1695])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&m[1695])|(m[1628]&m[1629]&~m[1630]&m[1631]&m[1695])|(m[1628]&~m[1629]&m[1630]&m[1631]&m[1695])|(~m[1628]&m[1629]&m[1630]&m[1631]&m[1695]))&~BiasedRNG[1035])|((m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1695])|(m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1695])|(~m[1628]&m[1629]&m[1630]&~m[1631]&~m[1695])|(m[1628]&m[1629]&m[1630]&~m[1631]&~m[1695])|(m[1628]&m[1629]&m[1630]&m[1631]&~m[1695])|(m[1628]&m[1629]&~m[1630]&~m[1631]&m[1695])|(m[1628]&~m[1629]&m[1630]&~m[1631]&m[1695])|(~m[1628]&m[1629]&m[1630]&~m[1631]&m[1695])|(m[1628]&m[1629]&m[1630]&~m[1631]&m[1695])|(m[1628]&m[1629]&m[1630]&m[1631]&m[1695]));
    m[1637] = (((m[1633]&~m[1634]&~m[1635]&~m[1636]&~m[1700])|(~m[1633]&m[1634]&~m[1635]&~m[1636]&~m[1700])|(~m[1633]&~m[1634]&m[1635]&~m[1636]&~m[1700])|(m[1633]&m[1634]&~m[1635]&m[1636]&~m[1700])|(m[1633]&~m[1634]&m[1635]&m[1636]&~m[1700])|(~m[1633]&m[1634]&m[1635]&m[1636]&~m[1700]))&BiasedRNG[1036])|(((m[1633]&~m[1634]&~m[1635]&~m[1636]&m[1700])|(~m[1633]&m[1634]&~m[1635]&~m[1636]&m[1700])|(~m[1633]&~m[1634]&m[1635]&~m[1636]&m[1700])|(m[1633]&m[1634]&~m[1635]&m[1636]&m[1700])|(m[1633]&~m[1634]&m[1635]&m[1636]&m[1700])|(~m[1633]&m[1634]&m[1635]&m[1636]&m[1700]))&~BiasedRNG[1036])|((m[1633]&m[1634]&~m[1635]&~m[1636]&~m[1700])|(m[1633]&~m[1634]&m[1635]&~m[1636]&~m[1700])|(~m[1633]&m[1634]&m[1635]&~m[1636]&~m[1700])|(m[1633]&m[1634]&m[1635]&~m[1636]&~m[1700])|(m[1633]&m[1634]&m[1635]&m[1636]&~m[1700])|(m[1633]&m[1634]&~m[1635]&~m[1636]&m[1700])|(m[1633]&~m[1634]&m[1635]&~m[1636]&m[1700])|(~m[1633]&m[1634]&m[1635]&~m[1636]&m[1700])|(m[1633]&m[1634]&m[1635]&~m[1636]&m[1700])|(m[1633]&m[1634]&m[1635]&m[1636]&m[1700]));
    m[1642] = (((m[1638]&~m[1639]&~m[1640]&~m[1641]&~m[1705])|(~m[1638]&m[1639]&~m[1640]&~m[1641]&~m[1705])|(~m[1638]&~m[1639]&m[1640]&~m[1641]&~m[1705])|(m[1638]&m[1639]&~m[1640]&m[1641]&~m[1705])|(m[1638]&~m[1639]&m[1640]&m[1641]&~m[1705])|(~m[1638]&m[1639]&m[1640]&m[1641]&~m[1705]))&BiasedRNG[1037])|(((m[1638]&~m[1639]&~m[1640]&~m[1641]&m[1705])|(~m[1638]&m[1639]&~m[1640]&~m[1641]&m[1705])|(~m[1638]&~m[1639]&m[1640]&~m[1641]&m[1705])|(m[1638]&m[1639]&~m[1640]&m[1641]&m[1705])|(m[1638]&~m[1639]&m[1640]&m[1641]&m[1705])|(~m[1638]&m[1639]&m[1640]&m[1641]&m[1705]))&~BiasedRNG[1037])|((m[1638]&m[1639]&~m[1640]&~m[1641]&~m[1705])|(m[1638]&~m[1639]&m[1640]&~m[1641]&~m[1705])|(~m[1638]&m[1639]&m[1640]&~m[1641]&~m[1705])|(m[1638]&m[1639]&m[1640]&~m[1641]&~m[1705])|(m[1638]&m[1639]&m[1640]&m[1641]&~m[1705])|(m[1638]&m[1639]&~m[1640]&~m[1641]&m[1705])|(m[1638]&~m[1639]&m[1640]&~m[1641]&m[1705])|(~m[1638]&m[1639]&m[1640]&~m[1641]&m[1705])|(m[1638]&m[1639]&m[1640]&~m[1641]&m[1705])|(m[1638]&m[1639]&m[1640]&m[1641]&m[1705]));
    m[1647] = (((m[1643]&~m[1644]&~m[1645]&~m[1646]&~m[1710])|(~m[1643]&m[1644]&~m[1645]&~m[1646]&~m[1710])|(~m[1643]&~m[1644]&m[1645]&~m[1646]&~m[1710])|(m[1643]&m[1644]&~m[1645]&m[1646]&~m[1710])|(m[1643]&~m[1644]&m[1645]&m[1646]&~m[1710])|(~m[1643]&m[1644]&m[1645]&m[1646]&~m[1710]))&BiasedRNG[1038])|(((m[1643]&~m[1644]&~m[1645]&~m[1646]&m[1710])|(~m[1643]&m[1644]&~m[1645]&~m[1646]&m[1710])|(~m[1643]&~m[1644]&m[1645]&~m[1646]&m[1710])|(m[1643]&m[1644]&~m[1645]&m[1646]&m[1710])|(m[1643]&~m[1644]&m[1645]&m[1646]&m[1710])|(~m[1643]&m[1644]&m[1645]&m[1646]&m[1710]))&~BiasedRNG[1038])|((m[1643]&m[1644]&~m[1645]&~m[1646]&~m[1710])|(m[1643]&~m[1644]&m[1645]&~m[1646]&~m[1710])|(~m[1643]&m[1644]&m[1645]&~m[1646]&~m[1710])|(m[1643]&m[1644]&m[1645]&~m[1646]&~m[1710])|(m[1643]&m[1644]&m[1645]&m[1646]&~m[1710])|(m[1643]&m[1644]&~m[1645]&~m[1646]&m[1710])|(m[1643]&~m[1644]&m[1645]&~m[1646]&m[1710])|(~m[1643]&m[1644]&m[1645]&~m[1646]&m[1710])|(m[1643]&m[1644]&m[1645]&~m[1646]&m[1710])|(m[1643]&m[1644]&m[1645]&m[1646]&m[1710]));
    m[1652] = (((m[1648]&~m[1649]&~m[1650]&~m[1651]&~m[1715])|(~m[1648]&m[1649]&~m[1650]&~m[1651]&~m[1715])|(~m[1648]&~m[1649]&m[1650]&~m[1651]&~m[1715])|(m[1648]&m[1649]&~m[1650]&m[1651]&~m[1715])|(m[1648]&~m[1649]&m[1650]&m[1651]&~m[1715])|(~m[1648]&m[1649]&m[1650]&m[1651]&~m[1715]))&BiasedRNG[1039])|(((m[1648]&~m[1649]&~m[1650]&~m[1651]&m[1715])|(~m[1648]&m[1649]&~m[1650]&~m[1651]&m[1715])|(~m[1648]&~m[1649]&m[1650]&~m[1651]&m[1715])|(m[1648]&m[1649]&~m[1650]&m[1651]&m[1715])|(m[1648]&~m[1649]&m[1650]&m[1651]&m[1715])|(~m[1648]&m[1649]&m[1650]&m[1651]&m[1715]))&~BiasedRNG[1039])|((m[1648]&m[1649]&~m[1650]&~m[1651]&~m[1715])|(m[1648]&~m[1649]&m[1650]&~m[1651]&~m[1715])|(~m[1648]&m[1649]&m[1650]&~m[1651]&~m[1715])|(m[1648]&m[1649]&m[1650]&~m[1651]&~m[1715])|(m[1648]&m[1649]&m[1650]&m[1651]&~m[1715])|(m[1648]&m[1649]&~m[1650]&~m[1651]&m[1715])|(m[1648]&~m[1649]&m[1650]&~m[1651]&m[1715])|(~m[1648]&m[1649]&m[1650]&~m[1651]&m[1715])|(m[1648]&m[1649]&m[1650]&~m[1651]&m[1715])|(m[1648]&m[1649]&m[1650]&m[1651]&m[1715]));
    m[1657] = (((m[1653]&~m[1654]&~m[1655]&~m[1656]&~m[1720])|(~m[1653]&m[1654]&~m[1655]&~m[1656]&~m[1720])|(~m[1653]&~m[1654]&m[1655]&~m[1656]&~m[1720])|(m[1653]&m[1654]&~m[1655]&m[1656]&~m[1720])|(m[1653]&~m[1654]&m[1655]&m[1656]&~m[1720])|(~m[1653]&m[1654]&m[1655]&m[1656]&~m[1720]))&BiasedRNG[1040])|(((m[1653]&~m[1654]&~m[1655]&~m[1656]&m[1720])|(~m[1653]&m[1654]&~m[1655]&~m[1656]&m[1720])|(~m[1653]&~m[1654]&m[1655]&~m[1656]&m[1720])|(m[1653]&m[1654]&~m[1655]&m[1656]&m[1720])|(m[1653]&~m[1654]&m[1655]&m[1656]&m[1720])|(~m[1653]&m[1654]&m[1655]&m[1656]&m[1720]))&~BiasedRNG[1040])|((m[1653]&m[1654]&~m[1655]&~m[1656]&~m[1720])|(m[1653]&~m[1654]&m[1655]&~m[1656]&~m[1720])|(~m[1653]&m[1654]&m[1655]&~m[1656]&~m[1720])|(m[1653]&m[1654]&m[1655]&~m[1656]&~m[1720])|(m[1653]&m[1654]&m[1655]&m[1656]&~m[1720])|(m[1653]&m[1654]&~m[1655]&~m[1656]&m[1720])|(m[1653]&~m[1654]&m[1655]&~m[1656]&m[1720])|(~m[1653]&m[1654]&m[1655]&~m[1656]&m[1720])|(m[1653]&m[1654]&m[1655]&~m[1656]&m[1720])|(m[1653]&m[1654]&m[1655]&m[1656]&m[1720]));
    m[1662] = (((m[1658]&~m[1659]&~m[1660]&~m[1661]&~m[1725])|(~m[1658]&m[1659]&~m[1660]&~m[1661]&~m[1725])|(~m[1658]&~m[1659]&m[1660]&~m[1661]&~m[1725])|(m[1658]&m[1659]&~m[1660]&m[1661]&~m[1725])|(m[1658]&~m[1659]&m[1660]&m[1661]&~m[1725])|(~m[1658]&m[1659]&m[1660]&m[1661]&~m[1725]))&BiasedRNG[1041])|(((m[1658]&~m[1659]&~m[1660]&~m[1661]&m[1725])|(~m[1658]&m[1659]&~m[1660]&~m[1661]&m[1725])|(~m[1658]&~m[1659]&m[1660]&~m[1661]&m[1725])|(m[1658]&m[1659]&~m[1660]&m[1661]&m[1725])|(m[1658]&~m[1659]&m[1660]&m[1661]&m[1725])|(~m[1658]&m[1659]&m[1660]&m[1661]&m[1725]))&~BiasedRNG[1041])|((m[1658]&m[1659]&~m[1660]&~m[1661]&~m[1725])|(m[1658]&~m[1659]&m[1660]&~m[1661]&~m[1725])|(~m[1658]&m[1659]&m[1660]&~m[1661]&~m[1725])|(m[1658]&m[1659]&m[1660]&~m[1661]&~m[1725])|(m[1658]&m[1659]&m[1660]&m[1661]&~m[1725])|(m[1658]&m[1659]&~m[1660]&~m[1661]&m[1725])|(m[1658]&~m[1659]&m[1660]&~m[1661]&m[1725])|(~m[1658]&m[1659]&m[1660]&~m[1661]&m[1725])|(m[1658]&m[1659]&m[1660]&~m[1661]&m[1725])|(m[1658]&m[1659]&m[1660]&m[1661]&m[1725]));
    m[1667] = (((m[1663]&~m[1664]&~m[1665]&~m[1666]&~m[1730])|(~m[1663]&m[1664]&~m[1665]&~m[1666]&~m[1730])|(~m[1663]&~m[1664]&m[1665]&~m[1666]&~m[1730])|(m[1663]&m[1664]&~m[1665]&m[1666]&~m[1730])|(m[1663]&~m[1664]&m[1665]&m[1666]&~m[1730])|(~m[1663]&m[1664]&m[1665]&m[1666]&~m[1730]))&BiasedRNG[1042])|(((m[1663]&~m[1664]&~m[1665]&~m[1666]&m[1730])|(~m[1663]&m[1664]&~m[1665]&~m[1666]&m[1730])|(~m[1663]&~m[1664]&m[1665]&~m[1666]&m[1730])|(m[1663]&m[1664]&~m[1665]&m[1666]&m[1730])|(m[1663]&~m[1664]&m[1665]&m[1666]&m[1730])|(~m[1663]&m[1664]&m[1665]&m[1666]&m[1730]))&~BiasedRNG[1042])|((m[1663]&m[1664]&~m[1665]&~m[1666]&~m[1730])|(m[1663]&~m[1664]&m[1665]&~m[1666]&~m[1730])|(~m[1663]&m[1664]&m[1665]&~m[1666]&~m[1730])|(m[1663]&m[1664]&m[1665]&~m[1666]&~m[1730])|(m[1663]&m[1664]&m[1665]&m[1666]&~m[1730])|(m[1663]&m[1664]&~m[1665]&~m[1666]&m[1730])|(m[1663]&~m[1664]&m[1665]&~m[1666]&m[1730])|(~m[1663]&m[1664]&m[1665]&~m[1666]&m[1730])|(m[1663]&m[1664]&m[1665]&~m[1666]&m[1730])|(m[1663]&m[1664]&m[1665]&m[1666]&m[1730]));
    m[1672] = (((m[1668]&~m[1669]&~m[1670]&~m[1671]&~m[1735])|(~m[1668]&m[1669]&~m[1670]&~m[1671]&~m[1735])|(~m[1668]&~m[1669]&m[1670]&~m[1671]&~m[1735])|(m[1668]&m[1669]&~m[1670]&m[1671]&~m[1735])|(m[1668]&~m[1669]&m[1670]&m[1671]&~m[1735])|(~m[1668]&m[1669]&m[1670]&m[1671]&~m[1735]))&BiasedRNG[1043])|(((m[1668]&~m[1669]&~m[1670]&~m[1671]&m[1735])|(~m[1668]&m[1669]&~m[1670]&~m[1671]&m[1735])|(~m[1668]&~m[1669]&m[1670]&~m[1671]&m[1735])|(m[1668]&m[1669]&~m[1670]&m[1671]&m[1735])|(m[1668]&~m[1669]&m[1670]&m[1671]&m[1735])|(~m[1668]&m[1669]&m[1670]&m[1671]&m[1735]))&~BiasedRNG[1043])|((m[1668]&m[1669]&~m[1670]&~m[1671]&~m[1735])|(m[1668]&~m[1669]&m[1670]&~m[1671]&~m[1735])|(~m[1668]&m[1669]&m[1670]&~m[1671]&~m[1735])|(m[1668]&m[1669]&m[1670]&~m[1671]&~m[1735])|(m[1668]&m[1669]&m[1670]&m[1671]&~m[1735])|(m[1668]&m[1669]&~m[1670]&~m[1671]&m[1735])|(m[1668]&~m[1669]&m[1670]&~m[1671]&m[1735])|(~m[1668]&m[1669]&m[1670]&~m[1671]&m[1735])|(m[1668]&m[1669]&m[1670]&~m[1671]&m[1735])|(m[1668]&m[1669]&m[1670]&m[1671]&m[1735]));
    m[1677] = (((m[1673]&~m[1674]&~m[1675]&~m[1676]&~m[1738])|(~m[1673]&m[1674]&~m[1675]&~m[1676]&~m[1738])|(~m[1673]&~m[1674]&m[1675]&~m[1676]&~m[1738])|(m[1673]&m[1674]&~m[1675]&m[1676]&~m[1738])|(m[1673]&~m[1674]&m[1675]&m[1676]&~m[1738])|(~m[1673]&m[1674]&m[1675]&m[1676]&~m[1738]))&BiasedRNG[1044])|(((m[1673]&~m[1674]&~m[1675]&~m[1676]&m[1738])|(~m[1673]&m[1674]&~m[1675]&~m[1676]&m[1738])|(~m[1673]&~m[1674]&m[1675]&~m[1676]&m[1738])|(m[1673]&m[1674]&~m[1675]&m[1676]&m[1738])|(m[1673]&~m[1674]&m[1675]&m[1676]&m[1738])|(~m[1673]&m[1674]&m[1675]&m[1676]&m[1738]))&~BiasedRNG[1044])|((m[1673]&m[1674]&~m[1675]&~m[1676]&~m[1738])|(m[1673]&~m[1674]&m[1675]&~m[1676]&~m[1738])|(~m[1673]&m[1674]&m[1675]&~m[1676]&~m[1738])|(m[1673]&m[1674]&m[1675]&~m[1676]&~m[1738])|(m[1673]&m[1674]&m[1675]&m[1676]&~m[1738])|(m[1673]&m[1674]&~m[1675]&~m[1676]&m[1738])|(m[1673]&~m[1674]&m[1675]&~m[1676]&m[1738])|(~m[1673]&m[1674]&m[1675]&~m[1676]&m[1738])|(m[1673]&m[1674]&m[1675]&~m[1676]&m[1738])|(m[1673]&m[1674]&m[1675]&m[1676]&m[1738]));
    m[1682] = (((m[1678]&~m[1679]&~m[1680]&~m[1681]&~m[1740])|(~m[1678]&m[1679]&~m[1680]&~m[1681]&~m[1740])|(~m[1678]&~m[1679]&m[1680]&~m[1681]&~m[1740])|(m[1678]&m[1679]&~m[1680]&m[1681]&~m[1740])|(m[1678]&~m[1679]&m[1680]&m[1681]&~m[1740])|(~m[1678]&m[1679]&m[1680]&m[1681]&~m[1740]))&BiasedRNG[1045])|(((m[1678]&~m[1679]&~m[1680]&~m[1681]&m[1740])|(~m[1678]&m[1679]&~m[1680]&~m[1681]&m[1740])|(~m[1678]&~m[1679]&m[1680]&~m[1681]&m[1740])|(m[1678]&m[1679]&~m[1680]&m[1681]&m[1740])|(m[1678]&~m[1679]&m[1680]&m[1681]&m[1740])|(~m[1678]&m[1679]&m[1680]&m[1681]&m[1740]))&~BiasedRNG[1045])|((m[1678]&m[1679]&~m[1680]&~m[1681]&~m[1740])|(m[1678]&~m[1679]&m[1680]&~m[1681]&~m[1740])|(~m[1678]&m[1679]&m[1680]&~m[1681]&~m[1740])|(m[1678]&m[1679]&m[1680]&~m[1681]&~m[1740])|(m[1678]&m[1679]&m[1680]&m[1681]&~m[1740])|(m[1678]&m[1679]&~m[1680]&~m[1681]&m[1740])|(m[1678]&~m[1679]&m[1680]&~m[1681]&m[1740])|(~m[1678]&m[1679]&m[1680]&~m[1681]&m[1740])|(m[1678]&m[1679]&m[1680]&~m[1681]&m[1740])|(m[1678]&m[1679]&m[1680]&m[1681]&m[1740]));
    m[1687] = (((m[1683]&~m[1684]&~m[1685]&~m[1686]&~m[1745])|(~m[1683]&m[1684]&~m[1685]&~m[1686]&~m[1745])|(~m[1683]&~m[1684]&m[1685]&~m[1686]&~m[1745])|(m[1683]&m[1684]&~m[1685]&m[1686]&~m[1745])|(m[1683]&~m[1684]&m[1685]&m[1686]&~m[1745])|(~m[1683]&m[1684]&m[1685]&m[1686]&~m[1745]))&BiasedRNG[1046])|(((m[1683]&~m[1684]&~m[1685]&~m[1686]&m[1745])|(~m[1683]&m[1684]&~m[1685]&~m[1686]&m[1745])|(~m[1683]&~m[1684]&m[1685]&~m[1686]&m[1745])|(m[1683]&m[1684]&~m[1685]&m[1686]&m[1745])|(m[1683]&~m[1684]&m[1685]&m[1686]&m[1745])|(~m[1683]&m[1684]&m[1685]&m[1686]&m[1745]))&~BiasedRNG[1046])|((m[1683]&m[1684]&~m[1685]&~m[1686]&~m[1745])|(m[1683]&~m[1684]&m[1685]&~m[1686]&~m[1745])|(~m[1683]&m[1684]&m[1685]&~m[1686]&~m[1745])|(m[1683]&m[1684]&m[1685]&~m[1686]&~m[1745])|(m[1683]&m[1684]&m[1685]&m[1686]&~m[1745])|(m[1683]&m[1684]&~m[1685]&~m[1686]&m[1745])|(m[1683]&~m[1684]&m[1685]&~m[1686]&m[1745])|(~m[1683]&m[1684]&m[1685]&~m[1686]&m[1745])|(m[1683]&m[1684]&m[1685]&~m[1686]&m[1745])|(m[1683]&m[1684]&m[1685]&m[1686]&m[1745]));
    m[1692] = (((m[1688]&~m[1689]&~m[1690]&~m[1691]&~m[1750])|(~m[1688]&m[1689]&~m[1690]&~m[1691]&~m[1750])|(~m[1688]&~m[1689]&m[1690]&~m[1691]&~m[1750])|(m[1688]&m[1689]&~m[1690]&m[1691]&~m[1750])|(m[1688]&~m[1689]&m[1690]&m[1691]&~m[1750])|(~m[1688]&m[1689]&m[1690]&m[1691]&~m[1750]))&BiasedRNG[1047])|(((m[1688]&~m[1689]&~m[1690]&~m[1691]&m[1750])|(~m[1688]&m[1689]&~m[1690]&~m[1691]&m[1750])|(~m[1688]&~m[1689]&m[1690]&~m[1691]&m[1750])|(m[1688]&m[1689]&~m[1690]&m[1691]&m[1750])|(m[1688]&~m[1689]&m[1690]&m[1691]&m[1750])|(~m[1688]&m[1689]&m[1690]&m[1691]&m[1750]))&~BiasedRNG[1047])|((m[1688]&m[1689]&~m[1690]&~m[1691]&~m[1750])|(m[1688]&~m[1689]&m[1690]&~m[1691]&~m[1750])|(~m[1688]&m[1689]&m[1690]&~m[1691]&~m[1750])|(m[1688]&m[1689]&m[1690]&~m[1691]&~m[1750])|(m[1688]&m[1689]&m[1690]&m[1691]&~m[1750])|(m[1688]&m[1689]&~m[1690]&~m[1691]&m[1750])|(m[1688]&~m[1689]&m[1690]&~m[1691]&m[1750])|(~m[1688]&m[1689]&m[1690]&~m[1691]&m[1750])|(m[1688]&m[1689]&m[1690]&~m[1691]&m[1750])|(m[1688]&m[1689]&m[1690]&m[1691]&m[1750]));
    m[1697] = (((m[1693]&~m[1694]&~m[1695]&~m[1696]&~m[1755])|(~m[1693]&m[1694]&~m[1695]&~m[1696]&~m[1755])|(~m[1693]&~m[1694]&m[1695]&~m[1696]&~m[1755])|(m[1693]&m[1694]&~m[1695]&m[1696]&~m[1755])|(m[1693]&~m[1694]&m[1695]&m[1696]&~m[1755])|(~m[1693]&m[1694]&m[1695]&m[1696]&~m[1755]))&BiasedRNG[1048])|(((m[1693]&~m[1694]&~m[1695]&~m[1696]&m[1755])|(~m[1693]&m[1694]&~m[1695]&~m[1696]&m[1755])|(~m[1693]&~m[1694]&m[1695]&~m[1696]&m[1755])|(m[1693]&m[1694]&~m[1695]&m[1696]&m[1755])|(m[1693]&~m[1694]&m[1695]&m[1696]&m[1755])|(~m[1693]&m[1694]&m[1695]&m[1696]&m[1755]))&~BiasedRNG[1048])|((m[1693]&m[1694]&~m[1695]&~m[1696]&~m[1755])|(m[1693]&~m[1694]&m[1695]&~m[1696]&~m[1755])|(~m[1693]&m[1694]&m[1695]&~m[1696]&~m[1755])|(m[1693]&m[1694]&m[1695]&~m[1696]&~m[1755])|(m[1693]&m[1694]&m[1695]&m[1696]&~m[1755])|(m[1693]&m[1694]&~m[1695]&~m[1696]&m[1755])|(m[1693]&~m[1694]&m[1695]&~m[1696]&m[1755])|(~m[1693]&m[1694]&m[1695]&~m[1696]&m[1755])|(m[1693]&m[1694]&m[1695]&~m[1696]&m[1755])|(m[1693]&m[1694]&m[1695]&m[1696]&m[1755]));
    m[1702] = (((m[1698]&~m[1699]&~m[1700]&~m[1701]&~m[1760])|(~m[1698]&m[1699]&~m[1700]&~m[1701]&~m[1760])|(~m[1698]&~m[1699]&m[1700]&~m[1701]&~m[1760])|(m[1698]&m[1699]&~m[1700]&m[1701]&~m[1760])|(m[1698]&~m[1699]&m[1700]&m[1701]&~m[1760])|(~m[1698]&m[1699]&m[1700]&m[1701]&~m[1760]))&BiasedRNG[1049])|(((m[1698]&~m[1699]&~m[1700]&~m[1701]&m[1760])|(~m[1698]&m[1699]&~m[1700]&~m[1701]&m[1760])|(~m[1698]&~m[1699]&m[1700]&~m[1701]&m[1760])|(m[1698]&m[1699]&~m[1700]&m[1701]&m[1760])|(m[1698]&~m[1699]&m[1700]&m[1701]&m[1760])|(~m[1698]&m[1699]&m[1700]&m[1701]&m[1760]))&~BiasedRNG[1049])|((m[1698]&m[1699]&~m[1700]&~m[1701]&~m[1760])|(m[1698]&~m[1699]&m[1700]&~m[1701]&~m[1760])|(~m[1698]&m[1699]&m[1700]&~m[1701]&~m[1760])|(m[1698]&m[1699]&m[1700]&~m[1701]&~m[1760])|(m[1698]&m[1699]&m[1700]&m[1701]&~m[1760])|(m[1698]&m[1699]&~m[1700]&~m[1701]&m[1760])|(m[1698]&~m[1699]&m[1700]&~m[1701]&m[1760])|(~m[1698]&m[1699]&m[1700]&~m[1701]&m[1760])|(m[1698]&m[1699]&m[1700]&~m[1701]&m[1760])|(m[1698]&m[1699]&m[1700]&m[1701]&m[1760]));
    m[1707] = (((m[1703]&~m[1704]&~m[1705]&~m[1706]&~m[1765])|(~m[1703]&m[1704]&~m[1705]&~m[1706]&~m[1765])|(~m[1703]&~m[1704]&m[1705]&~m[1706]&~m[1765])|(m[1703]&m[1704]&~m[1705]&m[1706]&~m[1765])|(m[1703]&~m[1704]&m[1705]&m[1706]&~m[1765])|(~m[1703]&m[1704]&m[1705]&m[1706]&~m[1765]))&BiasedRNG[1050])|(((m[1703]&~m[1704]&~m[1705]&~m[1706]&m[1765])|(~m[1703]&m[1704]&~m[1705]&~m[1706]&m[1765])|(~m[1703]&~m[1704]&m[1705]&~m[1706]&m[1765])|(m[1703]&m[1704]&~m[1705]&m[1706]&m[1765])|(m[1703]&~m[1704]&m[1705]&m[1706]&m[1765])|(~m[1703]&m[1704]&m[1705]&m[1706]&m[1765]))&~BiasedRNG[1050])|((m[1703]&m[1704]&~m[1705]&~m[1706]&~m[1765])|(m[1703]&~m[1704]&m[1705]&~m[1706]&~m[1765])|(~m[1703]&m[1704]&m[1705]&~m[1706]&~m[1765])|(m[1703]&m[1704]&m[1705]&~m[1706]&~m[1765])|(m[1703]&m[1704]&m[1705]&m[1706]&~m[1765])|(m[1703]&m[1704]&~m[1705]&~m[1706]&m[1765])|(m[1703]&~m[1704]&m[1705]&~m[1706]&m[1765])|(~m[1703]&m[1704]&m[1705]&~m[1706]&m[1765])|(m[1703]&m[1704]&m[1705]&~m[1706]&m[1765])|(m[1703]&m[1704]&m[1705]&m[1706]&m[1765]));
    m[1712] = (((m[1708]&~m[1709]&~m[1710]&~m[1711]&~m[1770])|(~m[1708]&m[1709]&~m[1710]&~m[1711]&~m[1770])|(~m[1708]&~m[1709]&m[1710]&~m[1711]&~m[1770])|(m[1708]&m[1709]&~m[1710]&m[1711]&~m[1770])|(m[1708]&~m[1709]&m[1710]&m[1711]&~m[1770])|(~m[1708]&m[1709]&m[1710]&m[1711]&~m[1770]))&BiasedRNG[1051])|(((m[1708]&~m[1709]&~m[1710]&~m[1711]&m[1770])|(~m[1708]&m[1709]&~m[1710]&~m[1711]&m[1770])|(~m[1708]&~m[1709]&m[1710]&~m[1711]&m[1770])|(m[1708]&m[1709]&~m[1710]&m[1711]&m[1770])|(m[1708]&~m[1709]&m[1710]&m[1711]&m[1770])|(~m[1708]&m[1709]&m[1710]&m[1711]&m[1770]))&~BiasedRNG[1051])|((m[1708]&m[1709]&~m[1710]&~m[1711]&~m[1770])|(m[1708]&~m[1709]&m[1710]&~m[1711]&~m[1770])|(~m[1708]&m[1709]&m[1710]&~m[1711]&~m[1770])|(m[1708]&m[1709]&m[1710]&~m[1711]&~m[1770])|(m[1708]&m[1709]&m[1710]&m[1711]&~m[1770])|(m[1708]&m[1709]&~m[1710]&~m[1711]&m[1770])|(m[1708]&~m[1709]&m[1710]&~m[1711]&m[1770])|(~m[1708]&m[1709]&m[1710]&~m[1711]&m[1770])|(m[1708]&m[1709]&m[1710]&~m[1711]&m[1770])|(m[1708]&m[1709]&m[1710]&m[1711]&m[1770]));
    m[1717] = (((m[1713]&~m[1714]&~m[1715]&~m[1716]&~m[1775])|(~m[1713]&m[1714]&~m[1715]&~m[1716]&~m[1775])|(~m[1713]&~m[1714]&m[1715]&~m[1716]&~m[1775])|(m[1713]&m[1714]&~m[1715]&m[1716]&~m[1775])|(m[1713]&~m[1714]&m[1715]&m[1716]&~m[1775])|(~m[1713]&m[1714]&m[1715]&m[1716]&~m[1775]))&BiasedRNG[1052])|(((m[1713]&~m[1714]&~m[1715]&~m[1716]&m[1775])|(~m[1713]&m[1714]&~m[1715]&~m[1716]&m[1775])|(~m[1713]&~m[1714]&m[1715]&~m[1716]&m[1775])|(m[1713]&m[1714]&~m[1715]&m[1716]&m[1775])|(m[1713]&~m[1714]&m[1715]&m[1716]&m[1775])|(~m[1713]&m[1714]&m[1715]&m[1716]&m[1775]))&~BiasedRNG[1052])|((m[1713]&m[1714]&~m[1715]&~m[1716]&~m[1775])|(m[1713]&~m[1714]&m[1715]&~m[1716]&~m[1775])|(~m[1713]&m[1714]&m[1715]&~m[1716]&~m[1775])|(m[1713]&m[1714]&m[1715]&~m[1716]&~m[1775])|(m[1713]&m[1714]&m[1715]&m[1716]&~m[1775])|(m[1713]&m[1714]&~m[1715]&~m[1716]&m[1775])|(m[1713]&~m[1714]&m[1715]&~m[1716]&m[1775])|(~m[1713]&m[1714]&m[1715]&~m[1716]&m[1775])|(m[1713]&m[1714]&m[1715]&~m[1716]&m[1775])|(m[1713]&m[1714]&m[1715]&m[1716]&m[1775]));
    m[1722] = (((m[1718]&~m[1719]&~m[1720]&~m[1721]&~m[1780])|(~m[1718]&m[1719]&~m[1720]&~m[1721]&~m[1780])|(~m[1718]&~m[1719]&m[1720]&~m[1721]&~m[1780])|(m[1718]&m[1719]&~m[1720]&m[1721]&~m[1780])|(m[1718]&~m[1719]&m[1720]&m[1721]&~m[1780])|(~m[1718]&m[1719]&m[1720]&m[1721]&~m[1780]))&BiasedRNG[1053])|(((m[1718]&~m[1719]&~m[1720]&~m[1721]&m[1780])|(~m[1718]&m[1719]&~m[1720]&~m[1721]&m[1780])|(~m[1718]&~m[1719]&m[1720]&~m[1721]&m[1780])|(m[1718]&m[1719]&~m[1720]&m[1721]&m[1780])|(m[1718]&~m[1719]&m[1720]&m[1721]&m[1780])|(~m[1718]&m[1719]&m[1720]&m[1721]&m[1780]))&~BiasedRNG[1053])|((m[1718]&m[1719]&~m[1720]&~m[1721]&~m[1780])|(m[1718]&~m[1719]&m[1720]&~m[1721]&~m[1780])|(~m[1718]&m[1719]&m[1720]&~m[1721]&~m[1780])|(m[1718]&m[1719]&m[1720]&~m[1721]&~m[1780])|(m[1718]&m[1719]&m[1720]&m[1721]&~m[1780])|(m[1718]&m[1719]&~m[1720]&~m[1721]&m[1780])|(m[1718]&~m[1719]&m[1720]&~m[1721]&m[1780])|(~m[1718]&m[1719]&m[1720]&~m[1721]&m[1780])|(m[1718]&m[1719]&m[1720]&~m[1721]&m[1780])|(m[1718]&m[1719]&m[1720]&m[1721]&m[1780]));
    m[1727] = (((m[1723]&~m[1724]&~m[1725]&~m[1726]&~m[1785])|(~m[1723]&m[1724]&~m[1725]&~m[1726]&~m[1785])|(~m[1723]&~m[1724]&m[1725]&~m[1726]&~m[1785])|(m[1723]&m[1724]&~m[1725]&m[1726]&~m[1785])|(m[1723]&~m[1724]&m[1725]&m[1726]&~m[1785])|(~m[1723]&m[1724]&m[1725]&m[1726]&~m[1785]))&BiasedRNG[1054])|(((m[1723]&~m[1724]&~m[1725]&~m[1726]&m[1785])|(~m[1723]&m[1724]&~m[1725]&~m[1726]&m[1785])|(~m[1723]&~m[1724]&m[1725]&~m[1726]&m[1785])|(m[1723]&m[1724]&~m[1725]&m[1726]&m[1785])|(m[1723]&~m[1724]&m[1725]&m[1726]&m[1785])|(~m[1723]&m[1724]&m[1725]&m[1726]&m[1785]))&~BiasedRNG[1054])|((m[1723]&m[1724]&~m[1725]&~m[1726]&~m[1785])|(m[1723]&~m[1724]&m[1725]&~m[1726]&~m[1785])|(~m[1723]&m[1724]&m[1725]&~m[1726]&~m[1785])|(m[1723]&m[1724]&m[1725]&~m[1726]&~m[1785])|(m[1723]&m[1724]&m[1725]&m[1726]&~m[1785])|(m[1723]&m[1724]&~m[1725]&~m[1726]&m[1785])|(m[1723]&~m[1724]&m[1725]&~m[1726]&m[1785])|(~m[1723]&m[1724]&m[1725]&~m[1726]&m[1785])|(m[1723]&m[1724]&m[1725]&~m[1726]&m[1785])|(m[1723]&m[1724]&m[1725]&m[1726]&m[1785]));
    m[1732] = (((m[1728]&~m[1729]&~m[1730]&~m[1731]&~m[1790])|(~m[1728]&m[1729]&~m[1730]&~m[1731]&~m[1790])|(~m[1728]&~m[1729]&m[1730]&~m[1731]&~m[1790])|(m[1728]&m[1729]&~m[1730]&m[1731]&~m[1790])|(m[1728]&~m[1729]&m[1730]&m[1731]&~m[1790])|(~m[1728]&m[1729]&m[1730]&m[1731]&~m[1790]))&BiasedRNG[1055])|(((m[1728]&~m[1729]&~m[1730]&~m[1731]&m[1790])|(~m[1728]&m[1729]&~m[1730]&~m[1731]&m[1790])|(~m[1728]&~m[1729]&m[1730]&~m[1731]&m[1790])|(m[1728]&m[1729]&~m[1730]&m[1731]&m[1790])|(m[1728]&~m[1729]&m[1730]&m[1731]&m[1790])|(~m[1728]&m[1729]&m[1730]&m[1731]&m[1790]))&~BiasedRNG[1055])|((m[1728]&m[1729]&~m[1730]&~m[1731]&~m[1790])|(m[1728]&~m[1729]&m[1730]&~m[1731]&~m[1790])|(~m[1728]&m[1729]&m[1730]&~m[1731]&~m[1790])|(m[1728]&m[1729]&m[1730]&~m[1731]&~m[1790])|(m[1728]&m[1729]&m[1730]&m[1731]&~m[1790])|(m[1728]&m[1729]&~m[1730]&~m[1731]&m[1790])|(m[1728]&~m[1729]&m[1730]&~m[1731]&m[1790])|(~m[1728]&m[1729]&m[1730]&~m[1731]&m[1790])|(m[1728]&m[1729]&m[1730]&~m[1731]&m[1790])|(m[1728]&m[1729]&m[1730]&m[1731]&m[1790]));
    m[1737] = (((m[1733]&~m[1734]&~m[1735]&~m[1736]&~m[1795])|(~m[1733]&m[1734]&~m[1735]&~m[1736]&~m[1795])|(~m[1733]&~m[1734]&m[1735]&~m[1736]&~m[1795])|(m[1733]&m[1734]&~m[1735]&m[1736]&~m[1795])|(m[1733]&~m[1734]&m[1735]&m[1736]&~m[1795])|(~m[1733]&m[1734]&m[1735]&m[1736]&~m[1795]))&BiasedRNG[1056])|(((m[1733]&~m[1734]&~m[1735]&~m[1736]&m[1795])|(~m[1733]&m[1734]&~m[1735]&~m[1736]&m[1795])|(~m[1733]&~m[1734]&m[1735]&~m[1736]&m[1795])|(m[1733]&m[1734]&~m[1735]&m[1736]&m[1795])|(m[1733]&~m[1734]&m[1735]&m[1736]&m[1795])|(~m[1733]&m[1734]&m[1735]&m[1736]&m[1795]))&~BiasedRNG[1056])|((m[1733]&m[1734]&~m[1735]&~m[1736]&~m[1795])|(m[1733]&~m[1734]&m[1735]&~m[1736]&~m[1795])|(~m[1733]&m[1734]&m[1735]&~m[1736]&~m[1795])|(m[1733]&m[1734]&m[1735]&~m[1736]&~m[1795])|(m[1733]&m[1734]&m[1735]&m[1736]&~m[1795])|(m[1733]&m[1734]&~m[1735]&~m[1736]&m[1795])|(m[1733]&~m[1734]&m[1735]&~m[1736]&m[1795])|(~m[1733]&m[1734]&m[1735]&~m[1736]&m[1795])|(m[1733]&m[1734]&m[1735]&~m[1736]&m[1795])|(m[1733]&m[1734]&m[1735]&m[1736]&m[1795]));
    m[1742] = (((m[1738]&~m[1739]&~m[1740]&~m[1741]&~m[1798])|(~m[1738]&m[1739]&~m[1740]&~m[1741]&~m[1798])|(~m[1738]&~m[1739]&m[1740]&~m[1741]&~m[1798])|(m[1738]&m[1739]&~m[1740]&m[1741]&~m[1798])|(m[1738]&~m[1739]&m[1740]&m[1741]&~m[1798])|(~m[1738]&m[1739]&m[1740]&m[1741]&~m[1798]))&BiasedRNG[1057])|(((m[1738]&~m[1739]&~m[1740]&~m[1741]&m[1798])|(~m[1738]&m[1739]&~m[1740]&~m[1741]&m[1798])|(~m[1738]&~m[1739]&m[1740]&~m[1741]&m[1798])|(m[1738]&m[1739]&~m[1740]&m[1741]&m[1798])|(m[1738]&~m[1739]&m[1740]&m[1741]&m[1798])|(~m[1738]&m[1739]&m[1740]&m[1741]&m[1798]))&~BiasedRNG[1057])|((m[1738]&m[1739]&~m[1740]&~m[1741]&~m[1798])|(m[1738]&~m[1739]&m[1740]&~m[1741]&~m[1798])|(~m[1738]&m[1739]&m[1740]&~m[1741]&~m[1798])|(m[1738]&m[1739]&m[1740]&~m[1741]&~m[1798])|(m[1738]&m[1739]&m[1740]&m[1741]&~m[1798])|(m[1738]&m[1739]&~m[1740]&~m[1741]&m[1798])|(m[1738]&~m[1739]&m[1740]&~m[1741]&m[1798])|(~m[1738]&m[1739]&m[1740]&~m[1741]&m[1798])|(m[1738]&m[1739]&m[1740]&~m[1741]&m[1798])|(m[1738]&m[1739]&m[1740]&m[1741]&m[1798]));
    m[1747] = (((m[1743]&~m[1744]&~m[1745]&~m[1746]&~m[1800])|(~m[1743]&m[1744]&~m[1745]&~m[1746]&~m[1800])|(~m[1743]&~m[1744]&m[1745]&~m[1746]&~m[1800])|(m[1743]&m[1744]&~m[1745]&m[1746]&~m[1800])|(m[1743]&~m[1744]&m[1745]&m[1746]&~m[1800])|(~m[1743]&m[1744]&m[1745]&m[1746]&~m[1800]))&BiasedRNG[1058])|(((m[1743]&~m[1744]&~m[1745]&~m[1746]&m[1800])|(~m[1743]&m[1744]&~m[1745]&~m[1746]&m[1800])|(~m[1743]&~m[1744]&m[1745]&~m[1746]&m[1800])|(m[1743]&m[1744]&~m[1745]&m[1746]&m[1800])|(m[1743]&~m[1744]&m[1745]&m[1746]&m[1800])|(~m[1743]&m[1744]&m[1745]&m[1746]&m[1800]))&~BiasedRNG[1058])|((m[1743]&m[1744]&~m[1745]&~m[1746]&~m[1800])|(m[1743]&~m[1744]&m[1745]&~m[1746]&~m[1800])|(~m[1743]&m[1744]&m[1745]&~m[1746]&~m[1800])|(m[1743]&m[1744]&m[1745]&~m[1746]&~m[1800])|(m[1743]&m[1744]&m[1745]&m[1746]&~m[1800])|(m[1743]&m[1744]&~m[1745]&~m[1746]&m[1800])|(m[1743]&~m[1744]&m[1745]&~m[1746]&m[1800])|(~m[1743]&m[1744]&m[1745]&~m[1746]&m[1800])|(m[1743]&m[1744]&m[1745]&~m[1746]&m[1800])|(m[1743]&m[1744]&m[1745]&m[1746]&m[1800]));
    m[1752] = (((m[1748]&~m[1749]&~m[1750]&~m[1751]&~m[1805])|(~m[1748]&m[1749]&~m[1750]&~m[1751]&~m[1805])|(~m[1748]&~m[1749]&m[1750]&~m[1751]&~m[1805])|(m[1748]&m[1749]&~m[1750]&m[1751]&~m[1805])|(m[1748]&~m[1749]&m[1750]&m[1751]&~m[1805])|(~m[1748]&m[1749]&m[1750]&m[1751]&~m[1805]))&BiasedRNG[1059])|(((m[1748]&~m[1749]&~m[1750]&~m[1751]&m[1805])|(~m[1748]&m[1749]&~m[1750]&~m[1751]&m[1805])|(~m[1748]&~m[1749]&m[1750]&~m[1751]&m[1805])|(m[1748]&m[1749]&~m[1750]&m[1751]&m[1805])|(m[1748]&~m[1749]&m[1750]&m[1751]&m[1805])|(~m[1748]&m[1749]&m[1750]&m[1751]&m[1805]))&~BiasedRNG[1059])|((m[1748]&m[1749]&~m[1750]&~m[1751]&~m[1805])|(m[1748]&~m[1749]&m[1750]&~m[1751]&~m[1805])|(~m[1748]&m[1749]&m[1750]&~m[1751]&~m[1805])|(m[1748]&m[1749]&m[1750]&~m[1751]&~m[1805])|(m[1748]&m[1749]&m[1750]&m[1751]&~m[1805])|(m[1748]&m[1749]&~m[1750]&~m[1751]&m[1805])|(m[1748]&~m[1749]&m[1750]&~m[1751]&m[1805])|(~m[1748]&m[1749]&m[1750]&~m[1751]&m[1805])|(m[1748]&m[1749]&m[1750]&~m[1751]&m[1805])|(m[1748]&m[1749]&m[1750]&m[1751]&m[1805]));
    m[1757] = (((m[1753]&~m[1754]&~m[1755]&~m[1756]&~m[1810])|(~m[1753]&m[1754]&~m[1755]&~m[1756]&~m[1810])|(~m[1753]&~m[1754]&m[1755]&~m[1756]&~m[1810])|(m[1753]&m[1754]&~m[1755]&m[1756]&~m[1810])|(m[1753]&~m[1754]&m[1755]&m[1756]&~m[1810])|(~m[1753]&m[1754]&m[1755]&m[1756]&~m[1810]))&BiasedRNG[1060])|(((m[1753]&~m[1754]&~m[1755]&~m[1756]&m[1810])|(~m[1753]&m[1754]&~m[1755]&~m[1756]&m[1810])|(~m[1753]&~m[1754]&m[1755]&~m[1756]&m[1810])|(m[1753]&m[1754]&~m[1755]&m[1756]&m[1810])|(m[1753]&~m[1754]&m[1755]&m[1756]&m[1810])|(~m[1753]&m[1754]&m[1755]&m[1756]&m[1810]))&~BiasedRNG[1060])|((m[1753]&m[1754]&~m[1755]&~m[1756]&~m[1810])|(m[1753]&~m[1754]&m[1755]&~m[1756]&~m[1810])|(~m[1753]&m[1754]&m[1755]&~m[1756]&~m[1810])|(m[1753]&m[1754]&m[1755]&~m[1756]&~m[1810])|(m[1753]&m[1754]&m[1755]&m[1756]&~m[1810])|(m[1753]&m[1754]&~m[1755]&~m[1756]&m[1810])|(m[1753]&~m[1754]&m[1755]&~m[1756]&m[1810])|(~m[1753]&m[1754]&m[1755]&~m[1756]&m[1810])|(m[1753]&m[1754]&m[1755]&~m[1756]&m[1810])|(m[1753]&m[1754]&m[1755]&m[1756]&m[1810]));
    m[1762] = (((m[1758]&~m[1759]&~m[1760]&~m[1761]&~m[1815])|(~m[1758]&m[1759]&~m[1760]&~m[1761]&~m[1815])|(~m[1758]&~m[1759]&m[1760]&~m[1761]&~m[1815])|(m[1758]&m[1759]&~m[1760]&m[1761]&~m[1815])|(m[1758]&~m[1759]&m[1760]&m[1761]&~m[1815])|(~m[1758]&m[1759]&m[1760]&m[1761]&~m[1815]))&BiasedRNG[1061])|(((m[1758]&~m[1759]&~m[1760]&~m[1761]&m[1815])|(~m[1758]&m[1759]&~m[1760]&~m[1761]&m[1815])|(~m[1758]&~m[1759]&m[1760]&~m[1761]&m[1815])|(m[1758]&m[1759]&~m[1760]&m[1761]&m[1815])|(m[1758]&~m[1759]&m[1760]&m[1761]&m[1815])|(~m[1758]&m[1759]&m[1760]&m[1761]&m[1815]))&~BiasedRNG[1061])|((m[1758]&m[1759]&~m[1760]&~m[1761]&~m[1815])|(m[1758]&~m[1759]&m[1760]&~m[1761]&~m[1815])|(~m[1758]&m[1759]&m[1760]&~m[1761]&~m[1815])|(m[1758]&m[1759]&m[1760]&~m[1761]&~m[1815])|(m[1758]&m[1759]&m[1760]&m[1761]&~m[1815])|(m[1758]&m[1759]&~m[1760]&~m[1761]&m[1815])|(m[1758]&~m[1759]&m[1760]&~m[1761]&m[1815])|(~m[1758]&m[1759]&m[1760]&~m[1761]&m[1815])|(m[1758]&m[1759]&m[1760]&~m[1761]&m[1815])|(m[1758]&m[1759]&m[1760]&m[1761]&m[1815]));
    m[1767] = (((m[1763]&~m[1764]&~m[1765]&~m[1766]&~m[1820])|(~m[1763]&m[1764]&~m[1765]&~m[1766]&~m[1820])|(~m[1763]&~m[1764]&m[1765]&~m[1766]&~m[1820])|(m[1763]&m[1764]&~m[1765]&m[1766]&~m[1820])|(m[1763]&~m[1764]&m[1765]&m[1766]&~m[1820])|(~m[1763]&m[1764]&m[1765]&m[1766]&~m[1820]))&BiasedRNG[1062])|(((m[1763]&~m[1764]&~m[1765]&~m[1766]&m[1820])|(~m[1763]&m[1764]&~m[1765]&~m[1766]&m[1820])|(~m[1763]&~m[1764]&m[1765]&~m[1766]&m[1820])|(m[1763]&m[1764]&~m[1765]&m[1766]&m[1820])|(m[1763]&~m[1764]&m[1765]&m[1766]&m[1820])|(~m[1763]&m[1764]&m[1765]&m[1766]&m[1820]))&~BiasedRNG[1062])|((m[1763]&m[1764]&~m[1765]&~m[1766]&~m[1820])|(m[1763]&~m[1764]&m[1765]&~m[1766]&~m[1820])|(~m[1763]&m[1764]&m[1765]&~m[1766]&~m[1820])|(m[1763]&m[1764]&m[1765]&~m[1766]&~m[1820])|(m[1763]&m[1764]&m[1765]&m[1766]&~m[1820])|(m[1763]&m[1764]&~m[1765]&~m[1766]&m[1820])|(m[1763]&~m[1764]&m[1765]&~m[1766]&m[1820])|(~m[1763]&m[1764]&m[1765]&~m[1766]&m[1820])|(m[1763]&m[1764]&m[1765]&~m[1766]&m[1820])|(m[1763]&m[1764]&m[1765]&m[1766]&m[1820]));
    m[1772] = (((m[1768]&~m[1769]&~m[1770]&~m[1771]&~m[1825])|(~m[1768]&m[1769]&~m[1770]&~m[1771]&~m[1825])|(~m[1768]&~m[1769]&m[1770]&~m[1771]&~m[1825])|(m[1768]&m[1769]&~m[1770]&m[1771]&~m[1825])|(m[1768]&~m[1769]&m[1770]&m[1771]&~m[1825])|(~m[1768]&m[1769]&m[1770]&m[1771]&~m[1825]))&BiasedRNG[1063])|(((m[1768]&~m[1769]&~m[1770]&~m[1771]&m[1825])|(~m[1768]&m[1769]&~m[1770]&~m[1771]&m[1825])|(~m[1768]&~m[1769]&m[1770]&~m[1771]&m[1825])|(m[1768]&m[1769]&~m[1770]&m[1771]&m[1825])|(m[1768]&~m[1769]&m[1770]&m[1771]&m[1825])|(~m[1768]&m[1769]&m[1770]&m[1771]&m[1825]))&~BiasedRNG[1063])|((m[1768]&m[1769]&~m[1770]&~m[1771]&~m[1825])|(m[1768]&~m[1769]&m[1770]&~m[1771]&~m[1825])|(~m[1768]&m[1769]&m[1770]&~m[1771]&~m[1825])|(m[1768]&m[1769]&m[1770]&~m[1771]&~m[1825])|(m[1768]&m[1769]&m[1770]&m[1771]&~m[1825])|(m[1768]&m[1769]&~m[1770]&~m[1771]&m[1825])|(m[1768]&~m[1769]&m[1770]&~m[1771]&m[1825])|(~m[1768]&m[1769]&m[1770]&~m[1771]&m[1825])|(m[1768]&m[1769]&m[1770]&~m[1771]&m[1825])|(m[1768]&m[1769]&m[1770]&m[1771]&m[1825]));
    m[1777] = (((m[1773]&~m[1774]&~m[1775]&~m[1776]&~m[1830])|(~m[1773]&m[1774]&~m[1775]&~m[1776]&~m[1830])|(~m[1773]&~m[1774]&m[1775]&~m[1776]&~m[1830])|(m[1773]&m[1774]&~m[1775]&m[1776]&~m[1830])|(m[1773]&~m[1774]&m[1775]&m[1776]&~m[1830])|(~m[1773]&m[1774]&m[1775]&m[1776]&~m[1830]))&BiasedRNG[1064])|(((m[1773]&~m[1774]&~m[1775]&~m[1776]&m[1830])|(~m[1773]&m[1774]&~m[1775]&~m[1776]&m[1830])|(~m[1773]&~m[1774]&m[1775]&~m[1776]&m[1830])|(m[1773]&m[1774]&~m[1775]&m[1776]&m[1830])|(m[1773]&~m[1774]&m[1775]&m[1776]&m[1830])|(~m[1773]&m[1774]&m[1775]&m[1776]&m[1830]))&~BiasedRNG[1064])|((m[1773]&m[1774]&~m[1775]&~m[1776]&~m[1830])|(m[1773]&~m[1774]&m[1775]&~m[1776]&~m[1830])|(~m[1773]&m[1774]&m[1775]&~m[1776]&~m[1830])|(m[1773]&m[1774]&m[1775]&~m[1776]&~m[1830])|(m[1773]&m[1774]&m[1775]&m[1776]&~m[1830])|(m[1773]&m[1774]&~m[1775]&~m[1776]&m[1830])|(m[1773]&~m[1774]&m[1775]&~m[1776]&m[1830])|(~m[1773]&m[1774]&m[1775]&~m[1776]&m[1830])|(m[1773]&m[1774]&m[1775]&~m[1776]&m[1830])|(m[1773]&m[1774]&m[1775]&m[1776]&m[1830]));
    m[1782] = (((m[1778]&~m[1779]&~m[1780]&~m[1781]&~m[1835])|(~m[1778]&m[1779]&~m[1780]&~m[1781]&~m[1835])|(~m[1778]&~m[1779]&m[1780]&~m[1781]&~m[1835])|(m[1778]&m[1779]&~m[1780]&m[1781]&~m[1835])|(m[1778]&~m[1779]&m[1780]&m[1781]&~m[1835])|(~m[1778]&m[1779]&m[1780]&m[1781]&~m[1835]))&BiasedRNG[1065])|(((m[1778]&~m[1779]&~m[1780]&~m[1781]&m[1835])|(~m[1778]&m[1779]&~m[1780]&~m[1781]&m[1835])|(~m[1778]&~m[1779]&m[1780]&~m[1781]&m[1835])|(m[1778]&m[1779]&~m[1780]&m[1781]&m[1835])|(m[1778]&~m[1779]&m[1780]&m[1781]&m[1835])|(~m[1778]&m[1779]&m[1780]&m[1781]&m[1835]))&~BiasedRNG[1065])|((m[1778]&m[1779]&~m[1780]&~m[1781]&~m[1835])|(m[1778]&~m[1779]&m[1780]&~m[1781]&~m[1835])|(~m[1778]&m[1779]&m[1780]&~m[1781]&~m[1835])|(m[1778]&m[1779]&m[1780]&~m[1781]&~m[1835])|(m[1778]&m[1779]&m[1780]&m[1781]&~m[1835])|(m[1778]&m[1779]&~m[1780]&~m[1781]&m[1835])|(m[1778]&~m[1779]&m[1780]&~m[1781]&m[1835])|(~m[1778]&m[1779]&m[1780]&~m[1781]&m[1835])|(m[1778]&m[1779]&m[1780]&~m[1781]&m[1835])|(m[1778]&m[1779]&m[1780]&m[1781]&m[1835]));
    m[1787] = (((m[1783]&~m[1784]&~m[1785]&~m[1786]&~m[1840])|(~m[1783]&m[1784]&~m[1785]&~m[1786]&~m[1840])|(~m[1783]&~m[1784]&m[1785]&~m[1786]&~m[1840])|(m[1783]&m[1784]&~m[1785]&m[1786]&~m[1840])|(m[1783]&~m[1784]&m[1785]&m[1786]&~m[1840])|(~m[1783]&m[1784]&m[1785]&m[1786]&~m[1840]))&BiasedRNG[1066])|(((m[1783]&~m[1784]&~m[1785]&~m[1786]&m[1840])|(~m[1783]&m[1784]&~m[1785]&~m[1786]&m[1840])|(~m[1783]&~m[1784]&m[1785]&~m[1786]&m[1840])|(m[1783]&m[1784]&~m[1785]&m[1786]&m[1840])|(m[1783]&~m[1784]&m[1785]&m[1786]&m[1840])|(~m[1783]&m[1784]&m[1785]&m[1786]&m[1840]))&~BiasedRNG[1066])|((m[1783]&m[1784]&~m[1785]&~m[1786]&~m[1840])|(m[1783]&~m[1784]&m[1785]&~m[1786]&~m[1840])|(~m[1783]&m[1784]&m[1785]&~m[1786]&~m[1840])|(m[1783]&m[1784]&m[1785]&~m[1786]&~m[1840])|(m[1783]&m[1784]&m[1785]&m[1786]&~m[1840])|(m[1783]&m[1784]&~m[1785]&~m[1786]&m[1840])|(m[1783]&~m[1784]&m[1785]&~m[1786]&m[1840])|(~m[1783]&m[1784]&m[1785]&~m[1786]&m[1840])|(m[1783]&m[1784]&m[1785]&~m[1786]&m[1840])|(m[1783]&m[1784]&m[1785]&m[1786]&m[1840]));
    m[1792] = (((m[1788]&~m[1789]&~m[1790]&~m[1791]&~m[1845])|(~m[1788]&m[1789]&~m[1790]&~m[1791]&~m[1845])|(~m[1788]&~m[1789]&m[1790]&~m[1791]&~m[1845])|(m[1788]&m[1789]&~m[1790]&m[1791]&~m[1845])|(m[1788]&~m[1789]&m[1790]&m[1791]&~m[1845])|(~m[1788]&m[1789]&m[1790]&m[1791]&~m[1845]))&BiasedRNG[1067])|(((m[1788]&~m[1789]&~m[1790]&~m[1791]&m[1845])|(~m[1788]&m[1789]&~m[1790]&~m[1791]&m[1845])|(~m[1788]&~m[1789]&m[1790]&~m[1791]&m[1845])|(m[1788]&m[1789]&~m[1790]&m[1791]&m[1845])|(m[1788]&~m[1789]&m[1790]&m[1791]&m[1845])|(~m[1788]&m[1789]&m[1790]&m[1791]&m[1845]))&~BiasedRNG[1067])|((m[1788]&m[1789]&~m[1790]&~m[1791]&~m[1845])|(m[1788]&~m[1789]&m[1790]&~m[1791]&~m[1845])|(~m[1788]&m[1789]&m[1790]&~m[1791]&~m[1845])|(m[1788]&m[1789]&m[1790]&~m[1791]&~m[1845])|(m[1788]&m[1789]&m[1790]&m[1791]&~m[1845])|(m[1788]&m[1789]&~m[1790]&~m[1791]&m[1845])|(m[1788]&~m[1789]&m[1790]&~m[1791]&m[1845])|(~m[1788]&m[1789]&m[1790]&~m[1791]&m[1845])|(m[1788]&m[1789]&m[1790]&~m[1791]&m[1845])|(m[1788]&m[1789]&m[1790]&m[1791]&m[1845]));
    m[1797] = (((m[1793]&~m[1794]&~m[1795]&~m[1796]&~m[1850])|(~m[1793]&m[1794]&~m[1795]&~m[1796]&~m[1850])|(~m[1793]&~m[1794]&m[1795]&~m[1796]&~m[1850])|(m[1793]&m[1794]&~m[1795]&m[1796]&~m[1850])|(m[1793]&~m[1794]&m[1795]&m[1796]&~m[1850])|(~m[1793]&m[1794]&m[1795]&m[1796]&~m[1850]))&BiasedRNG[1068])|(((m[1793]&~m[1794]&~m[1795]&~m[1796]&m[1850])|(~m[1793]&m[1794]&~m[1795]&~m[1796]&m[1850])|(~m[1793]&~m[1794]&m[1795]&~m[1796]&m[1850])|(m[1793]&m[1794]&~m[1795]&m[1796]&m[1850])|(m[1793]&~m[1794]&m[1795]&m[1796]&m[1850])|(~m[1793]&m[1794]&m[1795]&m[1796]&m[1850]))&~BiasedRNG[1068])|((m[1793]&m[1794]&~m[1795]&~m[1796]&~m[1850])|(m[1793]&~m[1794]&m[1795]&~m[1796]&~m[1850])|(~m[1793]&m[1794]&m[1795]&~m[1796]&~m[1850])|(m[1793]&m[1794]&m[1795]&~m[1796]&~m[1850])|(m[1793]&m[1794]&m[1795]&m[1796]&~m[1850])|(m[1793]&m[1794]&~m[1795]&~m[1796]&m[1850])|(m[1793]&~m[1794]&m[1795]&~m[1796]&m[1850])|(~m[1793]&m[1794]&m[1795]&~m[1796]&m[1850])|(m[1793]&m[1794]&m[1795]&~m[1796]&m[1850])|(m[1793]&m[1794]&m[1795]&m[1796]&m[1850]));
    m[1802] = (((m[1798]&~m[1799]&~m[1800]&~m[1801]&~m[1853])|(~m[1798]&m[1799]&~m[1800]&~m[1801]&~m[1853])|(~m[1798]&~m[1799]&m[1800]&~m[1801]&~m[1853])|(m[1798]&m[1799]&~m[1800]&m[1801]&~m[1853])|(m[1798]&~m[1799]&m[1800]&m[1801]&~m[1853])|(~m[1798]&m[1799]&m[1800]&m[1801]&~m[1853]))&BiasedRNG[1069])|(((m[1798]&~m[1799]&~m[1800]&~m[1801]&m[1853])|(~m[1798]&m[1799]&~m[1800]&~m[1801]&m[1853])|(~m[1798]&~m[1799]&m[1800]&~m[1801]&m[1853])|(m[1798]&m[1799]&~m[1800]&m[1801]&m[1853])|(m[1798]&~m[1799]&m[1800]&m[1801]&m[1853])|(~m[1798]&m[1799]&m[1800]&m[1801]&m[1853]))&~BiasedRNG[1069])|((m[1798]&m[1799]&~m[1800]&~m[1801]&~m[1853])|(m[1798]&~m[1799]&m[1800]&~m[1801]&~m[1853])|(~m[1798]&m[1799]&m[1800]&~m[1801]&~m[1853])|(m[1798]&m[1799]&m[1800]&~m[1801]&~m[1853])|(m[1798]&m[1799]&m[1800]&m[1801]&~m[1853])|(m[1798]&m[1799]&~m[1800]&~m[1801]&m[1853])|(m[1798]&~m[1799]&m[1800]&~m[1801]&m[1853])|(~m[1798]&m[1799]&m[1800]&~m[1801]&m[1853])|(m[1798]&m[1799]&m[1800]&~m[1801]&m[1853])|(m[1798]&m[1799]&m[1800]&m[1801]&m[1853]));
    m[1807] = (((m[1803]&~m[1804]&~m[1805]&~m[1806]&~m[1855])|(~m[1803]&m[1804]&~m[1805]&~m[1806]&~m[1855])|(~m[1803]&~m[1804]&m[1805]&~m[1806]&~m[1855])|(m[1803]&m[1804]&~m[1805]&m[1806]&~m[1855])|(m[1803]&~m[1804]&m[1805]&m[1806]&~m[1855])|(~m[1803]&m[1804]&m[1805]&m[1806]&~m[1855]))&BiasedRNG[1070])|(((m[1803]&~m[1804]&~m[1805]&~m[1806]&m[1855])|(~m[1803]&m[1804]&~m[1805]&~m[1806]&m[1855])|(~m[1803]&~m[1804]&m[1805]&~m[1806]&m[1855])|(m[1803]&m[1804]&~m[1805]&m[1806]&m[1855])|(m[1803]&~m[1804]&m[1805]&m[1806]&m[1855])|(~m[1803]&m[1804]&m[1805]&m[1806]&m[1855]))&~BiasedRNG[1070])|((m[1803]&m[1804]&~m[1805]&~m[1806]&~m[1855])|(m[1803]&~m[1804]&m[1805]&~m[1806]&~m[1855])|(~m[1803]&m[1804]&m[1805]&~m[1806]&~m[1855])|(m[1803]&m[1804]&m[1805]&~m[1806]&~m[1855])|(m[1803]&m[1804]&m[1805]&m[1806]&~m[1855])|(m[1803]&m[1804]&~m[1805]&~m[1806]&m[1855])|(m[1803]&~m[1804]&m[1805]&~m[1806]&m[1855])|(~m[1803]&m[1804]&m[1805]&~m[1806]&m[1855])|(m[1803]&m[1804]&m[1805]&~m[1806]&m[1855])|(m[1803]&m[1804]&m[1805]&m[1806]&m[1855]));
    m[1812] = (((m[1808]&~m[1809]&~m[1810]&~m[1811]&~m[1860])|(~m[1808]&m[1809]&~m[1810]&~m[1811]&~m[1860])|(~m[1808]&~m[1809]&m[1810]&~m[1811]&~m[1860])|(m[1808]&m[1809]&~m[1810]&m[1811]&~m[1860])|(m[1808]&~m[1809]&m[1810]&m[1811]&~m[1860])|(~m[1808]&m[1809]&m[1810]&m[1811]&~m[1860]))&BiasedRNG[1071])|(((m[1808]&~m[1809]&~m[1810]&~m[1811]&m[1860])|(~m[1808]&m[1809]&~m[1810]&~m[1811]&m[1860])|(~m[1808]&~m[1809]&m[1810]&~m[1811]&m[1860])|(m[1808]&m[1809]&~m[1810]&m[1811]&m[1860])|(m[1808]&~m[1809]&m[1810]&m[1811]&m[1860])|(~m[1808]&m[1809]&m[1810]&m[1811]&m[1860]))&~BiasedRNG[1071])|((m[1808]&m[1809]&~m[1810]&~m[1811]&~m[1860])|(m[1808]&~m[1809]&m[1810]&~m[1811]&~m[1860])|(~m[1808]&m[1809]&m[1810]&~m[1811]&~m[1860])|(m[1808]&m[1809]&m[1810]&~m[1811]&~m[1860])|(m[1808]&m[1809]&m[1810]&m[1811]&~m[1860])|(m[1808]&m[1809]&~m[1810]&~m[1811]&m[1860])|(m[1808]&~m[1809]&m[1810]&~m[1811]&m[1860])|(~m[1808]&m[1809]&m[1810]&~m[1811]&m[1860])|(m[1808]&m[1809]&m[1810]&~m[1811]&m[1860])|(m[1808]&m[1809]&m[1810]&m[1811]&m[1860]));
    m[1817] = (((m[1813]&~m[1814]&~m[1815]&~m[1816]&~m[1865])|(~m[1813]&m[1814]&~m[1815]&~m[1816]&~m[1865])|(~m[1813]&~m[1814]&m[1815]&~m[1816]&~m[1865])|(m[1813]&m[1814]&~m[1815]&m[1816]&~m[1865])|(m[1813]&~m[1814]&m[1815]&m[1816]&~m[1865])|(~m[1813]&m[1814]&m[1815]&m[1816]&~m[1865]))&BiasedRNG[1072])|(((m[1813]&~m[1814]&~m[1815]&~m[1816]&m[1865])|(~m[1813]&m[1814]&~m[1815]&~m[1816]&m[1865])|(~m[1813]&~m[1814]&m[1815]&~m[1816]&m[1865])|(m[1813]&m[1814]&~m[1815]&m[1816]&m[1865])|(m[1813]&~m[1814]&m[1815]&m[1816]&m[1865])|(~m[1813]&m[1814]&m[1815]&m[1816]&m[1865]))&~BiasedRNG[1072])|((m[1813]&m[1814]&~m[1815]&~m[1816]&~m[1865])|(m[1813]&~m[1814]&m[1815]&~m[1816]&~m[1865])|(~m[1813]&m[1814]&m[1815]&~m[1816]&~m[1865])|(m[1813]&m[1814]&m[1815]&~m[1816]&~m[1865])|(m[1813]&m[1814]&m[1815]&m[1816]&~m[1865])|(m[1813]&m[1814]&~m[1815]&~m[1816]&m[1865])|(m[1813]&~m[1814]&m[1815]&~m[1816]&m[1865])|(~m[1813]&m[1814]&m[1815]&~m[1816]&m[1865])|(m[1813]&m[1814]&m[1815]&~m[1816]&m[1865])|(m[1813]&m[1814]&m[1815]&m[1816]&m[1865]));
    m[1822] = (((m[1818]&~m[1819]&~m[1820]&~m[1821]&~m[1870])|(~m[1818]&m[1819]&~m[1820]&~m[1821]&~m[1870])|(~m[1818]&~m[1819]&m[1820]&~m[1821]&~m[1870])|(m[1818]&m[1819]&~m[1820]&m[1821]&~m[1870])|(m[1818]&~m[1819]&m[1820]&m[1821]&~m[1870])|(~m[1818]&m[1819]&m[1820]&m[1821]&~m[1870]))&BiasedRNG[1073])|(((m[1818]&~m[1819]&~m[1820]&~m[1821]&m[1870])|(~m[1818]&m[1819]&~m[1820]&~m[1821]&m[1870])|(~m[1818]&~m[1819]&m[1820]&~m[1821]&m[1870])|(m[1818]&m[1819]&~m[1820]&m[1821]&m[1870])|(m[1818]&~m[1819]&m[1820]&m[1821]&m[1870])|(~m[1818]&m[1819]&m[1820]&m[1821]&m[1870]))&~BiasedRNG[1073])|((m[1818]&m[1819]&~m[1820]&~m[1821]&~m[1870])|(m[1818]&~m[1819]&m[1820]&~m[1821]&~m[1870])|(~m[1818]&m[1819]&m[1820]&~m[1821]&~m[1870])|(m[1818]&m[1819]&m[1820]&~m[1821]&~m[1870])|(m[1818]&m[1819]&m[1820]&m[1821]&~m[1870])|(m[1818]&m[1819]&~m[1820]&~m[1821]&m[1870])|(m[1818]&~m[1819]&m[1820]&~m[1821]&m[1870])|(~m[1818]&m[1819]&m[1820]&~m[1821]&m[1870])|(m[1818]&m[1819]&m[1820]&~m[1821]&m[1870])|(m[1818]&m[1819]&m[1820]&m[1821]&m[1870]));
    m[1827] = (((m[1823]&~m[1824]&~m[1825]&~m[1826]&~m[1875])|(~m[1823]&m[1824]&~m[1825]&~m[1826]&~m[1875])|(~m[1823]&~m[1824]&m[1825]&~m[1826]&~m[1875])|(m[1823]&m[1824]&~m[1825]&m[1826]&~m[1875])|(m[1823]&~m[1824]&m[1825]&m[1826]&~m[1875])|(~m[1823]&m[1824]&m[1825]&m[1826]&~m[1875]))&BiasedRNG[1074])|(((m[1823]&~m[1824]&~m[1825]&~m[1826]&m[1875])|(~m[1823]&m[1824]&~m[1825]&~m[1826]&m[1875])|(~m[1823]&~m[1824]&m[1825]&~m[1826]&m[1875])|(m[1823]&m[1824]&~m[1825]&m[1826]&m[1875])|(m[1823]&~m[1824]&m[1825]&m[1826]&m[1875])|(~m[1823]&m[1824]&m[1825]&m[1826]&m[1875]))&~BiasedRNG[1074])|((m[1823]&m[1824]&~m[1825]&~m[1826]&~m[1875])|(m[1823]&~m[1824]&m[1825]&~m[1826]&~m[1875])|(~m[1823]&m[1824]&m[1825]&~m[1826]&~m[1875])|(m[1823]&m[1824]&m[1825]&~m[1826]&~m[1875])|(m[1823]&m[1824]&m[1825]&m[1826]&~m[1875])|(m[1823]&m[1824]&~m[1825]&~m[1826]&m[1875])|(m[1823]&~m[1824]&m[1825]&~m[1826]&m[1875])|(~m[1823]&m[1824]&m[1825]&~m[1826]&m[1875])|(m[1823]&m[1824]&m[1825]&~m[1826]&m[1875])|(m[1823]&m[1824]&m[1825]&m[1826]&m[1875]));
    m[1832] = (((m[1828]&~m[1829]&~m[1830]&~m[1831]&~m[1880])|(~m[1828]&m[1829]&~m[1830]&~m[1831]&~m[1880])|(~m[1828]&~m[1829]&m[1830]&~m[1831]&~m[1880])|(m[1828]&m[1829]&~m[1830]&m[1831]&~m[1880])|(m[1828]&~m[1829]&m[1830]&m[1831]&~m[1880])|(~m[1828]&m[1829]&m[1830]&m[1831]&~m[1880]))&BiasedRNG[1075])|(((m[1828]&~m[1829]&~m[1830]&~m[1831]&m[1880])|(~m[1828]&m[1829]&~m[1830]&~m[1831]&m[1880])|(~m[1828]&~m[1829]&m[1830]&~m[1831]&m[1880])|(m[1828]&m[1829]&~m[1830]&m[1831]&m[1880])|(m[1828]&~m[1829]&m[1830]&m[1831]&m[1880])|(~m[1828]&m[1829]&m[1830]&m[1831]&m[1880]))&~BiasedRNG[1075])|((m[1828]&m[1829]&~m[1830]&~m[1831]&~m[1880])|(m[1828]&~m[1829]&m[1830]&~m[1831]&~m[1880])|(~m[1828]&m[1829]&m[1830]&~m[1831]&~m[1880])|(m[1828]&m[1829]&m[1830]&~m[1831]&~m[1880])|(m[1828]&m[1829]&m[1830]&m[1831]&~m[1880])|(m[1828]&m[1829]&~m[1830]&~m[1831]&m[1880])|(m[1828]&~m[1829]&m[1830]&~m[1831]&m[1880])|(~m[1828]&m[1829]&m[1830]&~m[1831]&m[1880])|(m[1828]&m[1829]&m[1830]&~m[1831]&m[1880])|(m[1828]&m[1829]&m[1830]&m[1831]&m[1880]));
    m[1837] = (((m[1833]&~m[1834]&~m[1835]&~m[1836]&~m[1885])|(~m[1833]&m[1834]&~m[1835]&~m[1836]&~m[1885])|(~m[1833]&~m[1834]&m[1835]&~m[1836]&~m[1885])|(m[1833]&m[1834]&~m[1835]&m[1836]&~m[1885])|(m[1833]&~m[1834]&m[1835]&m[1836]&~m[1885])|(~m[1833]&m[1834]&m[1835]&m[1836]&~m[1885]))&BiasedRNG[1076])|(((m[1833]&~m[1834]&~m[1835]&~m[1836]&m[1885])|(~m[1833]&m[1834]&~m[1835]&~m[1836]&m[1885])|(~m[1833]&~m[1834]&m[1835]&~m[1836]&m[1885])|(m[1833]&m[1834]&~m[1835]&m[1836]&m[1885])|(m[1833]&~m[1834]&m[1835]&m[1836]&m[1885])|(~m[1833]&m[1834]&m[1835]&m[1836]&m[1885]))&~BiasedRNG[1076])|((m[1833]&m[1834]&~m[1835]&~m[1836]&~m[1885])|(m[1833]&~m[1834]&m[1835]&~m[1836]&~m[1885])|(~m[1833]&m[1834]&m[1835]&~m[1836]&~m[1885])|(m[1833]&m[1834]&m[1835]&~m[1836]&~m[1885])|(m[1833]&m[1834]&m[1835]&m[1836]&~m[1885])|(m[1833]&m[1834]&~m[1835]&~m[1836]&m[1885])|(m[1833]&~m[1834]&m[1835]&~m[1836]&m[1885])|(~m[1833]&m[1834]&m[1835]&~m[1836]&m[1885])|(m[1833]&m[1834]&m[1835]&~m[1836]&m[1885])|(m[1833]&m[1834]&m[1835]&m[1836]&m[1885]));
    m[1842] = (((m[1838]&~m[1839]&~m[1840]&~m[1841]&~m[1890])|(~m[1838]&m[1839]&~m[1840]&~m[1841]&~m[1890])|(~m[1838]&~m[1839]&m[1840]&~m[1841]&~m[1890])|(m[1838]&m[1839]&~m[1840]&m[1841]&~m[1890])|(m[1838]&~m[1839]&m[1840]&m[1841]&~m[1890])|(~m[1838]&m[1839]&m[1840]&m[1841]&~m[1890]))&BiasedRNG[1077])|(((m[1838]&~m[1839]&~m[1840]&~m[1841]&m[1890])|(~m[1838]&m[1839]&~m[1840]&~m[1841]&m[1890])|(~m[1838]&~m[1839]&m[1840]&~m[1841]&m[1890])|(m[1838]&m[1839]&~m[1840]&m[1841]&m[1890])|(m[1838]&~m[1839]&m[1840]&m[1841]&m[1890])|(~m[1838]&m[1839]&m[1840]&m[1841]&m[1890]))&~BiasedRNG[1077])|((m[1838]&m[1839]&~m[1840]&~m[1841]&~m[1890])|(m[1838]&~m[1839]&m[1840]&~m[1841]&~m[1890])|(~m[1838]&m[1839]&m[1840]&~m[1841]&~m[1890])|(m[1838]&m[1839]&m[1840]&~m[1841]&~m[1890])|(m[1838]&m[1839]&m[1840]&m[1841]&~m[1890])|(m[1838]&m[1839]&~m[1840]&~m[1841]&m[1890])|(m[1838]&~m[1839]&m[1840]&~m[1841]&m[1890])|(~m[1838]&m[1839]&m[1840]&~m[1841]&m[1890])|(m[1838]&m[1839]&m[1840]&~m[1841]&m[1890])|(m[1838]&m[1839]&m[1840]&m[1841]&m[1890]));
    m[1847] = (((m[1843]&~m[1844]&~m[1845]&~m[1846]&~m[1895])|(~m[1843]&m[1844]&~m[1845]&~m[1846]&~m[1895])|(~m[1843]&~m[1844]&m[1845]&~m[1846]&~m[1895])|(m[1843]&m[1844]&~m[1845]&m[1846]&~m[1895])|(m[1843]&~m[1844]&m[1845]&m[1846]&~m[1895])|(~m[1843]&m[1844]&m[1845]&m[1846]&~m[1895]))&BiasedRNG[1078])|(((m[1843]&~m[1844]&~m[1845]&~m[1846]&m[1895])|(~m[1843]&m[1844]&~m[1845]&~m[1846]&m[1895])|(~m[1843]&~m[1844]&m[1845]&~m[1846]&m[1895])|(m[1843]&m[1844]&~m[1845]&m[1846]&m[1895])|(m[1843]&~m[1844]&m[1845]&m[1846]&m[1895])|(~m[1843]&m[1844]&m[1845]&m[1846]&m[1895]))&~BiasedRNG[1078])|((m[1843]&m[1844]&~m[1845]&~m[1846]&~m[1895])|(m[1843]&~m[1844]&m[1845]&~m[1846]&~m[1895])|(~m[1843]&m[1844]&m[1845]&~m[1846]&~m[1895])|(m[1843]&m[1844]&m[1845]&~m[1846]&~m[1895])|(m[1843]&m[1844]&m[1845]&m[1846]&~m[1895])|(m[1843]&m[1844]&~m[1845]&~m[1846]&m[1895])|(m[1843]&~m[1844]&m[1845]&~m[1846]&m[1895])|(~m[1843]&m[1844]&m[1845]&~m[1846]&m[1895])|(m[1843]&m[1844]&m[1845]&~m[1846]&m[1895])|(m[1843]&m[1844]&m[1845]&m[1846]&m[1895]));
    m[1852] = (((m[1848]&~m[1849]&~m[1850]&~m[1851]&~m[1900])|(~m[1848]&m[1849]&~m[1850]&~m[1851]&~m[1900])|(~m[1848]&~m[1849]&m[1850]&~m[1851]&~m[1900])|(m[1848]&m[1849]&~m[1850]&m[1851]&~m[1900])|(m[1848]&~m[1849]&m[1850]&m[1851]&~m[1900])|(~m[1848]&m[1849]&m[1850]&m[1851]&~m[1900]))&BiasedRNG[1079])|(((m[1848]&~m[1849]&~m[1850]&~m[1851]&m[1900])|(~m[1848]&m[1849]&~m[1850]&~m[1851]&m[1900])|(~m[1848]&~m[1849]&m[1850]&~m[1851]&m[1900])|(m[1848]&m[1849]&~m[1850]&m[1851]&m[1900])|(m[1848]&~m[1849]&m[1850]&m[1851]&m[1900])|(~m[1848]&m[1849]&m[1850]&m[1851]&m[1900]))&~BiasedRNG[1079])|((m[1848]&m[1849]&~m[1850]&~m[1851]&~m[1900])|(m[1848]&~m[1849]&m[1850]&~m[1851]&~m[1900])|(~m[1848]&m[1849]&m[1850]&~m[1851]&~m[1900])|(m[1848]&m[1849]&m[1850]&~m[1851]&~m[1900])|(m[1848]&m[1849]&m[1850]&m[1851]&~m[1900])|(m[1848]&m[1849]&~m[1850]&~m[1851]&m[1900])|(m[1848]&~m[1849]&m[1850]&~m[1851]&m[1900])|(~m[1848]&m[1849]&m[1850]&~m[1851]&m[1900])|(m[1848]&m[1849]&m[1850]&~m[1851]&m[1900])|(m[1848]&m[1849]&m[1850]&m[1851]&m[1900]));
    m[1857] = (((m[1853]&~m[1854]&~m[1855]&~m[1856]&~m[1903])|(~m[1853]&m[1854]&~m[1855]&~m[1856]&~m[1903])|(~m[1853]&~m[1854]&m[1855]&~m[1856]&~m[1903])|(m[1853]&m[1854]&~m[1855]&m[1856]&~m[1903])|(m[1853]&~m[1854]&m[1855]&m[1856]&~m[1903])|(~m[1853]&m[1854]&m[1855]&m[1856]&~m[1903]))&BiasedRNG[1080])|(((m[1853]&~m[1854]&~m[1855]&~m[1856]&m[1903])|(~m[1853]&m[1854]&~m[1855]&~m[1856]&m[1903])|(~m[1853]&~m[1854]&m[1855]&~m[1856]&m[1903])|(m[1853]&m[1854]&~m[1855]&m[1856]&m[1903])|(m[1853]&~m[1854]&m[1855]&m[1856]&m[1903])|(~m[1853]&m[1854]&m[1855]&m[1856]&m[1903]))&~BiasedRNG[1080])|((m[1853]&m[1854]&~m[1855]&~m[1856]&~m[1903])|(m[1853]&~m[1854]&m[1855]&~m[1856]&~m[1903])|(~m[1853]&m[1854]&m[1855]&~m[1856]&~m[1903])|(m[1853]&m[1854]&m[1855]&~m[1856]&~m[1903])|(m[1853]&m[1854]&m[1855]&m[1856]&~m[1903])|(m[1853]&m[1854]&~m[1855]&~m[1856]&m[1903])|(m[1853]&~m[1854]&m[1855]&~m[1856]&m[1903])|(~m[1853]&m[1854]&m[1855]&~m[1856]&m[1903])|(m[1853]&m[1854]&m[1855]&~m[1856]&m[1903])|(m[1853]&m[1854]&m[1855]&m[1856]&m[1903]));
    m[1862] = (((m[1858]&~m[1859]&~m[1860]&~m[1861]&~m[1905])|(~m[1858]&m[1859]&~m[1860]&~m[1861]&~m[1905])|(~m[1858]&~m[1859]&m[1860]&~m[1861]&~m[1905])|(m[1858]&m[1859]&~m[1860]&m[1861]&~m[1905])|(m[1858]&~m[1859]&m[1860]&m[1861]&~m[1905])|(~m[1858]&m[1859]&m[1860]&m[1861]&~m[1905]))&BiasedRNG[1081])|(((m[1858]&~m[1859]&~m[1860]&~m[1861]&m[1905])|(~m[1858]&m[1859]&~m[1860]&~m[1861]&m[1905])|(~m[1858]&~m[1859]&m[1860]&~m[1861]&m[1905])|(m[1858]&m[1859]&~m[1860]&m[1861]&m[1905])|(m[1858]&~m[1859]&m[1860]&m[1861]&m[1905])|(~m[1858]&m[1859]&m[1860]&m[1861]&m[1905]))&~BiasedRNG[1081])|((m[1858]&m[1859]&~m[1860]&~m[1861]&~m[1905])|(m[1858]&~m[1859]&m[1860]&~m[1861]&~m[1905])|(~m[1858]&m[1859]&m[1860]&~m[1861]&~m[1905])|(m[1858]&m[1859]&m[1860]&~m[1861]&~m[1905])|(m[1858]&m[1859]&m[1860]&m[1861]&~m[1905])|(m[1858]&m[1859]&~m[1860]&~m[1861]&m[1905])|(m[1858]&~m[1859]&m[1860]&~m[1861]&m[1905])|(~m[1858]&m[1859]&m[1860]&~m[1861]&m[1905])|(m[1858]&m[1859]&m[1860]&~m[1861]&m[1905])|(m[1858]&m[1859]&m[1860]&m[1861]&m[1905]));
    m[1867] = (((m[1863]&~m[1864]&~m[1865]&~m[1866]&~m[1910])|(~m[1863]&m[1864]&~m[1865]&~m[1866]&~m[1910])|(~m[1863]&~m[1864]&m[1865]&~m[1866]&~m[1910])|(m[1863]&m[1864]&~m[1865]&m[1866]&~m[1910])|(m[1863]&~m[1864]&m[1865]&m[1866]&~m[1910])|(~m[1863]&m[1864]&m[1865]&m[1866]&~m[1910]))&BiasedRNG[1082])|(((m[1863]&~m[1864]&~m[1865]&~m[1866]&m[1910])|(~m[1863]&m[1864]&~m[1865]&~m[1866]&m[1910])|(~m[1863]&~m[1864]&m[1865]&~m[1866]&m[1910])|(m[1863]&m[1864]&~m[1865]&m[1866]&m[1910])|(m[1863]&~m[1864]&m[1865]&m[1866]&m[1910])|(~m[1863]&m[1864]&m[1865]&m[1866]&m[1910]))&~BiasedRNG[1082])|((m[1863]&m[1864]&~m[1865]&~m[1866]&~m[1910])|(m[1863]&~m[1864]&m[1865]&~m[1866]&~m[1910])|(~m[1863]&m[1864]&m[1865]&~m[1866]&~m[1910])|(m[1863]&m[1864]&m[1865]&~m[1866]&~m[1910])|(m[1863]&m[1864]&m[1865]&m[1866]&~m[1910])|(m[1863]&m[1864]&~m[1865]&~m[1866]&m[1910])|(m[1863]&~m[1864]&m[1865]&~m[1866]&m[1910])|(~m[1863]&m[1864]&m[1865]&~m[1866]&m[1910])|(m[1863]&m[1864]&m[1865]&~m[1866]&m[1910])|(m[1863]&m[1864]&m[1865]&m[1866]&m[1910]));
    m[1872] = (((m[1868]&~m[1869]&~m[1870]&~m[1871]&~m[1915])|(~m[1868]&m[1869]&~m[1870]&~m[1871]&~m[1915])|(~m[1868]&~m[1869]&m[1870]&~m[1871]&~m[1915])|(m[1868]&m[1869]&~m[1870]&m[1871]&~m[1915])|(m[1868]&~m[1869]&m[1870]&m[1871]&~m[1915])|(~m[1868]&m[1869]&m[1870]&m[1871]&~m[1915]))&BiasedRNG[1083])|(((m[1868]&~m[1869]&~m[1870]&~m[1871]&m[1915])|(~m[1868]&m[1869]&~m[1870]&~m[1871]&m[1915])|(~m[1868]&~m[1869]&m[1870]&~m[1871]&m[1915])|(m[1868]&m[1869]&~m[1870]&m[1871]&m[1915])|(m[1868]&~m[1869]&m[1870]&m[1871]&m[1915])|(~m[1868]&m[1869]&m[1870]&m[1871]&m[1915]))&~BiasedRNG[1083])|((m[1868]&m[1869]&~m[1870]&~m[1871]&~m[1915])|(m[1868]&~m[1869]&m[1870]&~m[1871]&~m[1915])|(~m[1868]&m[1869]&m[1870]&~m[1871]&~m[1915])|(m[1868]&m[1869]&m[1870]&~m[1871]&~m[1915])|(m[1868]&m[1869]&m[1870]&m[1871]&~m[1915])|(m[1868]&m[1869]&~m[1870]&~m[1871]&m[1915])|(m[1868]&~m[1869]&m[1870]&~m[1871]&m[1915])|(~m[1868]&m[1869]&m[1870]&~m[1871]&m[1915])|(m[1868]&m[1869]&m[1870]&~m[1871]&m[1915])|(m[1868]&m[1869]&m[1870]&m[1871]&m[1915]));
    m[1877] = (((m[1873]&~m[1874]&~m[1875]&~m[1876]&~m[1920])|(~m[1873]&m[1874]&~m[1875]&~m[1876]&~m[1920])|(~m[1873]&~m[1874]&m[1875]&~m[1876]&~m[1920])|(m[1873]&m[1874]&~m[1875]&m[1876]&~m[1920])|(m[1873]&~m[1874]&m[1875]&m[1876]&~m[1920])|(~m[1873]&m[1874]&m[1875]&m[1876]&~m[1920]))&BiasedRNG[1084])|(((m[1873]&~m[1874]&~m[1875]&~m[1876]&m[1920])|(~m[1873]&m[1874]&~m[1875]&~m[1876]&m[1920])|(~m[1873]&~m[1874]&m[1875]&~m[1876]&m[1920])|(m[1873]&m[1874]&~m[1875]&m[1876]&m[1920])|(m[1873]&~m[1874]&m[1875]&m[1876]&m[1920])|(~m[1873]&m[1874]&m[1875]&m[1876]&m[1920]))&~BiasedRNG[1084])|((m[1873]&m[1874]&~m[1875]&~m[1876]&~m[1920])|(m[1873]&~m[1874]&m[1875]&~m[1876]&~m[1920])|(~m[1873]&m[1874]&m[1875]&~m[1876]&~m[1920])|(m[1873]&m[1874]&m[1875]&~m[1876]&~m[1920])|(m[1873]&m[1874]&m[1875]&m[1876]&~m[1920])|(m[1873]&m[1874]&~m[1875]&~m[1876]&m[1920])|(m[1873]&~m[1874]&m[1875]&~m[1876]&m[1920])|(~m[1873]&m[1874]&m[1875]&~m[1876]&m[1920])|(m[1873]&m[1874]&m[1875]&~m[1876]&m[1920])|(m[1873]&m[1874]&m[1875]&m[1876]&m[1920]));
    m[1882] = (((m[1878]&~m[1879]&~m[1880]&~m[1881]&~m[1925])|(~m[1878]&m[1879]&~m[1880]&~m[1881]&~m[1925])|(~m[1878]&~m[1879]&m[1880]&~m[1881]&~m[1925])|(m[1878]&m[1879]&~m[1880]&m[1881]&~m[1925])|(m[1878]&~m[1879]&m[1880]&m[1881]&~m[1925])|(~m[1878]&m[1879]&m[1880]&m[1881]&~m[1925]))&BiasedRNG[1085])|(((m[1878]&~m[1879]&~m[1880]&~m[1881]&m[1925])|(~m[1878]&m[1879]&~m[1880]&~m[1881]&m[1925])|(~m[1878]&~m[1879]&m[1880]&~m[1881]&m[1925])|(m[1878]&m[1879]&~m[1880]&m[1881]&m[1925])|(m[1878]&~m[1879]&m[1880]&m[1881]&m[1925])|(~m[1878]&m[1879]&m[1880]&m[1881]&m[1925]))&~BiasedRNG[1085])|((m[1878]&m[1879]&~m[1880]&~m[1881]&~m[1925])|(m[1878]&~m[1879]&m[1880]&~m[1881]&~m[1925])|(~m[1878]&m[1879]&m[1880]&~m[1881]&~m[1925])|(m[1878]&m[1879]&m[1880]&~m[1881]&~m[1925])|(m[1878]&m[1879]&m[1880]&m[1881]&~m[1925])|(m[1878]&m[1879]&~m[1880]&~m[1881]&m[1925])|(m[1878]&~m[1879]&m[1880]&~m[1881]&m[1925])|(~m[1878]&m[1879]&m[1880]&~m[1881]&m[1925])|(m[1878]&m[1879]&m[1880]&~m[1881]&m[1925])|(m[1878]&m[1879]&m[1880]&m[1881]&m[1925]));
    m[1887] = (((m[1883]&~m[1884]&~m[1885]&~m[1886]&~m[1930])|(~m[1883]&m[1884]&~m[1885]&~m[1886]&~m[1930])|(~m[1883]&~m[1884]&m[1885]&~m[1886]&~m[1930])|(m[1883]&m[1884]&~m[1885]&m[1886]&~m[1930])|(m[1883]&~m[1884]&m[1885]&m[1886]&~m[1930])|(~m[1883]&m[1884]&m[1885]&m[1886]&~m[1930]))&BiasedRNG[1086])|(((m[1883]&~m[1884]&~m[1885]&~m[1886]&m[1930])|(~m[1883]&m[1884]&~m[1885]&~m[1886]&m[1930])|(~m[1883]&~m[1884]&m[1885]&~m[1886]&m[1930])|(m[1883]&m[1884]&~m[1885]&m[1886]&m[1930])|(m[1883]&~m[1884]&m[1885]&m[1886]&m[1930])|(~m[1883]&m[1884]&m[1885]&m[1886]&m[1930]))&~BiasedRNG[1086])|((m[1883]&m[1884]&~m[1885]&~m[1886]&~m[1930])|(m[1883]&~m[1884]&m[1885]&~m[1886]&~m[1930])|(~m[1883]&m[1884]&m[1885]&~m[1886]&~m[1930])|(m[1883]&m[1884]&m[1885]&~m[1886]&~m[1930])|(m[1883]&m[1884]&m[1885]&m[1886]&~m[1930])|(m[1883]&m[1884]&~m[1885]&~m[1886]&m[1930])|(m[1883]&~m[1884]&m[1885]&~m[1886]&m[1930])|(~m[1883]&m[1884]&m[1885]&~m[1886]&m[1930])|(m[1883]&m[1884]&m[1885]&~m[1886]&m[1930])|(m[1883]&m[1884]&m[1885]&m[1886]&m[1930]));
    m[1892] = (((m[1888]&~m[1889]&~m[1890]&~m[1891]&~m[1935])|(~m[1888]&m[1889]&~m[1890]&~m[1891]&~m[1935])|(~m[1888]&~m[1889]&m[1890]&~m[1891]&~m[1935])|(m[1888]&m[1889]&~m[1890]&m[1891]&~m[1935])|(m[1888]&~m[1889]&m[1890]&m[1891]&~m[1935])|(~m[1888]&m[1889]&m[1890]&m[1891]&~m[1935]))&BiasedRNG[1087])|(((m[1888]&~m[1889]&~m[1890]&~m[1891]&m[1935])|(~m[1888]&m[1889]&~m[1890]&~m[1891]&m[1935])|(~m[1888]&~m[1889]&m[1890]&~m[1891]&m[1935])|(m[1888]&m[1889]&~m[1890]&m[1891]&m[1935])|(m[1888]&~m[1889]&m[1890]&m[1891]&m[1935])|(~m[1888]&m[1889]&m[1890]&m[1891]&m[1935]))&~BiasedRNG[1087])|((m[1888]&m[1889]&~m[1890]&~m[1891]&~m[1935])|(m[1888]&~m[1889]&m[1890]&~m[1891]&~m[1935])|(~m[1888]&m[1889]&m[1890]&~m[1891]&~m[1935])|(m[1888]&m[1889]&m[1890]&~m[1891]&~m[1935])|(m[1888]&m[1889]&m[1890]&m[1891]&~m[1935])|(m[1888]&m[1889]&~m[1890]&~m[1891]&m[1935])|(m[1888]&~m[1889]&m[1890]&~m[1891]&m[1935])|(~m[1888]&m[1889]&m[1890]&~m[1891]&m[1935])|(m[1888]&m[1889]&m[1890]&~m[1891]&m[1935])|(m[1888]&m[1889]&m[1890]&m[1891]&m[1935]));
    m[1897] = (((m[1893]&~m[1894]&~m[1895]&~m[1896]&~m[1940])|(~m[1893]&m[1894]&~m[1895]&~m[1896]&~m[1940])|(~m[1893]&~m[1894]&m[1895]&~m[1896]&~m[1940])|(m[1893]&m[1894]&~m[1895]&m[1896]&~m[1940])|(m[1893]&~m[1894]&m[1895]&m[1896]&~m[1940])|(~m[1893]&m[1894]&m[1895]&m[1896]&~m[1940]))&BiasedRNG[1088])|(((m[1893]&~m[1894]&~m[1895]&~m[1896]&m[1940])|(~m[1893]&m[1894]&~m[1895]&~m[1896]&m[1940])|(~m[1893]&~m[1894]&m[1895]&~m[1896]&m[1940])|(m[1893]&m[1894]&~m[1895]&m[1896]&m[1940])|(m[1893]&~m[1894]&m[1895]&m[1896]&m[1940])|(~m[1893]&m[1894]&m[1895]&m[1896]&m[1940]))&~BiasedRNG[1088])|((m[1893]&m[1894]&~m[1895]&~m[1896]&~m[1940])|(m[1893]&~m[1894]&m[1895]&~m[1896]&~m[1940])|(~m[1893]&m[1894]&m[1895]&~m[1896]&~m[1940])|(m[1893]&m[1894]&m[1895]&~m[1896]&~m[1940])|(m[1893]&m[1894]&m[1895]&m[1896]&~m[1940])|(m[1893]&m[1894]&~m[1895]&~m[1896]&m[1940])|(m[1893]&~m[1894]&m[1895]&~m[1896]&m[1940])|(~m[1893]&m[1894]&m[1895]&~m[1896]&m[1940])|(m[1893]&m[1894]&m[1895]&~m[1896]&m[1940])|(m[1893]&m[1894]&m[1895]&m[1896]&m[1940]));
    m[1902] = (((m[1898]&~m[1899]&~m[1900]&~m[1901]&~m[1945])|(~m[1898]&m[1899]&~m[1900]&~m[1901]&~m[1945])|(~m[1898]&~m[1899]&m[1900]&~m[1901]&~m[1945])|(m[1898]&m[1899]&~m[1900]&m[1901]&~m[1945])|(m[1898]&~m[1899]&m[1900]&m[1901]&~m[1945])|(~m[1898]&m[1899]&m[1900]&m[1901]&~m[1945]))&BiasedRNG[1089])|(((m[1898]&~m[1899]&~m[1900]&~m[1901]&m[1945])|(~m[1898]&m[1899]&~m[1900]&~m[1901]&m[1945])|(~m[1898]&~m[1899]&m[1900]&~m[1901]&m[1945])|(m[1898]&m[1899]&~m[1900]&m[1901]&m[1945])|(m[1898]&~m[1899]&m[1900]&m[1901]&m[1945])|(~m[1898]&m[1899]&m[1900]&m[1901]&m[1945]))&~BiasedRNG[1089])|((m[1898]&m[1899]&~m[1900]&~m[1901]&~m[1945])|(m[1898]&~m[1899]&m[1900]&~m[1901]&~m[1945])|(~m[1898]&m[1899]&m[1900]&~m[1901]&~m[1945])|(m[1898]&m[1899]&m[1900]&~m[1901]&~m[1945])|(m[1898]&m[1899]&m[1900]&m[1901]&~m[1945])|(m[1898]&m[1899]&~m[1900]&~m[1901]&m[1945])|(m[1898]&~m[1899]&m[1900]&~m[1901]&m[1945])|(~m[1898]&m[1899]&m[1900]&~m[1901]&m[1945])|(m[1898]&m[1899]&m[1900]&~m[1901]&m[1945])|(m[1898]&m[1899]&m[1900]&m[1901]&m[1945]));
    m[1907] = (((m[1903]&~m[1904]&~m[1905]&~m[1906]&~m[1948])|(~m[1903]&m[1904]&~m[1905]&~m[1906]&~m[1948])|(~m[1903]&~m[1904]&m[1905]&~m[1906]&~m[1948])|(m[1903]&m[1904]&~m[1905]&m[1906]&~m[1948])|(m[1903]&~m[1904]&m[1905]&m[1906]&~m[1948])|(~m[1903]&m[1904]&m[1905]&m[1906]&~m[1948]))&BiasedRNG[1090])|(((m[1903]&~m[1904]&~m[1905]&~m[1906]&m[1948])|(~m[1903]&m[1904]&~m[1905]&~m[1906]&m[1948])|(~m[1903]&~m[1904]&m[1905]&~m[1906]&m[1948])|(m[1903]&m[1904]&~m[1905]&m[1906]&m[1948])|(m[1903]&~m[1904]&m[1905]&m[1906]&m[1948])|(~m[1903]&m[1904]&m[1905]&m[1906]&m[1948]))&~BiasedRNG[1090])|((m[1903]&m[1904]&~m[1905]&~m[1906]&~m[1948])|(m[1903]&~m[1904]&m[1905]&~m[1906]&~m[1948])|(~m[1903]&m[1904]&m[1905]&~m[1906]&~m[1948])|(m[1903]&m[1904]&m[1905]&~m[1906]&~m[1948])|(m[1903]&m[1904]&m[1905]&m[1906]&~m[1948])|(m[1903]&m[1904]&~m[1905]&~m[1906]&m[1948])|(m[1903]&~m[1904]&m[1905]&~m[1906]&m[1948])|(~m[1903]&m[1904]&m[1905]&~m[1906]&m[1948])|(m[1903]&m[1904]&m[1905]&~m[1906]&m[1948])|(m[1903]&m[1904]&m[1905]&m[1906]&m[1948]));
    m[1912] = (((m[1908]&~m[1909]&~m[1910]&~m[1911]&~m[1950])|(~m[1908]&m[1909]&~m[1910]&~m[1911]&~m[1950])|(~m[1908]&~m[1909]&m[1910]&~m[1911]&~m[1950])|(m[1908]&m[1909]&~m[1910]&m[1911]&~m[1950])|(m[1908]&~m[1909]&m[1910]&m[1911]&~m[1950])|(~m[1908]&m[1909]&m[1910]&m[1911]&~m[1950]))&BiasedRNG[1091])|(((m[1908]&~m[1909]&~m[1910]&~m[1911]&m[1950])|(~m[1908]&m[1909]&~m[1910]&~m[1911]&m[1950])|(~m[1908]&~m[1909]&m[1910]&~m[1911]&m[1950])|(m[1908]&m[1909]&~m[1910]&m[1911]&m[1950])|(m[1908]&~m[1909]&m[1910]&m[1911]&m[1950])|(~m[1908]&m[1909]&m[1910]&m[1911]&m[1950]))&~BiasedRNG[1091])|((m[1908]&m[1909]&~m[1910]&~m[1911]&~m[1950])|(m[1908]&~m[1909]&m[1910]&~m[1911]&~m[1950])|(~m[1908]&m[1909]&m[1910]&~m[1911]&~m[1950])|(m[1908]&m[1909]&m[1910]&~m[1911]&~m[1950])|(m[1908]&m[1909]&m[1910]&m[1911]&~m[1950])|(m[1908]&m[1909]&~m[1910]&~m[1911]&m[1950])|(m[1908]&~m[1909]&m[1910]&~m[1911]&m[1950])|(~m[1908]&m[1909]&m[1910]&~m[1911]&m[1950])|(m[1908]&m[1909]&m[1910]&~m[1911]&m[1950])|(m[1908]&m[1909]&m[1910]&m[1911]&m[1950]));
    m[1917] = (((m[1913]&~m[1914]&~m[1915]&~m[1916]&~m[1955])|(~m[1913]&m[1914]&~m[1915]&~m[1916]&~m[1955])|(~m[1913]&~m[1914]&m[1915]&~m[1916]&~m[1955])|(m[1913]&m[1914]&~m[1915]&m[1916]&~m[1955])|(m[1913]&~m[1914]&m[1915]&m[1916]&~m[1955])|(~m[1913]&m[1914]&m[1915]&m[1916]&~m[1955]))&BiasedRNG[1092])|(((m[1913]&~m[1914]&~m[1915]&~m[1916]&m[1955])|(~m[1913]&m[1914]&~m[1915]&~m[1916]&m[1955])|(~m[1913]&~m[1914]&m[1915]&~m[1916]&m[1955])|(m[1913]&m[1914]&~m[1915]&m[1916]&m[1955])|(m[1913]&~m[1914]&m[1915]&m[1916]&m[1955])|(~m[1913]&m[1914]&m[1915]&m[1916]&m[1955]))&~BiasedRNG[1092])|((m[1913]&m[1914]&~m[1915]&~m[1916]&~m[1955])|(m[1913]&~m[1914]&m[1915]&~m[1916]&~m[1955])|(~m[1913]&m[1914]&m[1915]&~m[1916]&~m[1955])|(m[1913]&m[1914]&m[1915]&~m[1916]&~m[1955])|(m[1913]&m[1914]&m[1915]&m[1916]&~m[1955])|(m[1913]&m[1914]&~m[1915]&~m[1916]&m[1955])|(m[1913]&~m[1914]&m[1915]&~m[1916]&m[1955])|(~m[1913]&m[1914]&m[1915]&~m[1916]&m[1955])|(m[1913]&m[1914]&m[1915]&~m[1916]&m[1955])|(m[1913]&m[1914]&m[1915]&m[1916]&m[1955]));
    m[1922] = (((m[1918]&~m[1919]&~m[1920]&~m[1921]&~m[1960])|(~m[1918]&m[1919]&~m[1920]&~m[1921]&~m[1960])|(~m[1918]&~m[1919]&m[1920]&~m[1921]&~m[1960])|(m[1918]&m[1919]&~m[1920]&m[1921]&~m[1960])|(m[1918]&~m[1919]&m[1920]&m[1921]&~m[1960])|(~m[1918]&m[1919]&m[1920]&m[1921]&~m[1960]))&BiasedRNG[1093])|(((m[1918]&~m[1919]&~m[1920]&~m[1921]&m[1960])|(~m[1918]&m[1919]&~m[1920]&~m[1921]&m[1960])|(~m[1918]&~m[1919]&m[1920]&~m[1921]&m[1960])|(m[1918]&m[1919]&~m[1920]&m[1921]&m[1960])|(m[1918]&~m[1919]&m[1920]&m[1921]&m[1960])|(~m[1918]&m[1919]&m[1920]&m[1921]&m[1960]))&~BiasedRNG[1093])|((m[1918]&m[1919]&~m[1920]&~m[1921]&~m[1960])|(m[1918]&~m[1919]&m[1920]&~m[1921]&~m[1960])|(~m[1918]&m[1919]&m[1920]&~m[1921]&~m[1960])|(m[1918]&m[1919]&m[1920]&~m[1921]&~m[1960])|(m[1918]&m[1919]&m[1920]&m[1921]&~m[1960])|(m[1918]&m[1919]&~m[1920]&~m[1921]&m[1960])|(m[1918]&~m[1919]&m[1920]&~m[1921]&m[1960])|(~m[1918]&m[1919]&m[1920]&~m[1921]&m[1960])|(m[1918]&m[1919]&m[1920]&~m[1921]&m[1960])|(m[1918]&m[1919]&m[1920]&m[1921]&m[1960]));
    m[1927] = (((m[1923]&~m[1924]&~m[1925]&~m[1926]&~m[1965])|(~m[1923]&m[1924]&~m[1925]&~m[1926]&~m[1965])|(~m[1923]&~m[1924]&m[1925]&~m[1926]&~m[1965])|(m[1923]&m[1924]&~m[1925]&m[1926]&~m[1965])|(m[1923]&~m[1924]&m[1925]&m[1926]&~m[1965])|(~m[1923]&m[1924]&m[1925]&m[1926]&~m[1965]))&BiasedRNG[1094])|(((m[1923]&~m[1924]&~m[1925]&~m[1926]&m[1965])|(~m[1923]&m[1924]&~m[1925]&~m[1926]&m[1965])|(~m[1923]&~m[1924]&m[1925]&~m[1926]&m[1965])|(m[1923]&m[1924]&~m[1925]&m[1926]&m[1965])|(m[1923]&~m[1924]&m[1925]&m[1926]&m[1965])|(~m[1923]&m[1924]&m[1925]&m[1926]&m[1965]))&~BiasedRNG[1094])|((m[1923]&m[1924]&~m[1925]&~m[1926]&~m[1965])|(m[1923]&~m[1924]&m[1925]&~m[1926]&~m[1965])|(~m[1923]&m[1924]&m[1925]&~m[1926]&~m[1965])|(m[1923]&m[1924]&m[1925]&~m[1926]&~m[1965])|(m[1923]&m[1924]&m[1925]&m[1926]&~m[1965])|(m[1923]&m[1924]&~m[1925]&~m[1926]&m[1965])|(m[1923]&~m[1924]&m[1925]&~m[1926]&m[1965])|(~m[1923]&m[1924]&m[1925]&~m[1926]&m[1965])|(m[1923]&m[1924]&m[1925]&~m[1926]&m[1965])|(m[1923]&m[1924]&m[1925]&m[1926]&m[1965]));
    m[1932] = (((m[1928]&~m[1929]&~m[1930]&~m[1931]&~m[1970])|(~m[1928]&m[1929]&~m[1930]&~m[1931]&~m[1970])|(~m[1928]&~m[1929]&m[1930]&~m[1931]&~m[1970])|(m[1928]&m[1929]&~m[1930]&m[1931]&~m[1970])|(m[1928]&~m[1929]&m[1930]&m[1931]&~m[1970])|(~m[1928]&m[1929]&m[1930]&m[1931]&~m[1970]))&BiasedRNG[1095])|(((m[1928]&~m[1929]&~m[1930]&~m[1931]&m[1970])|(~m[1928]&m[1929]&~m[1930]&~m[1931]&m[1970])|(~m[1928]&~m[1929]&m[1930]&~m[1931]&m[1970])|(m[1928]&m[1929]&~m[1930]&m[1931]&m[1970])|(m[1928]&~m[1929]&m[1930]&m[1931]&m[1970])|(~m[1928]&m[1929]&m[1930]&m[1931]&m[1970]))&~BiasedRNG[1095])|((m[1928]&m[1929]&~m[1930]&~m[1931]&~m[1970])|(m[1928]&~m[1929]&m[1930]&~m[1931]&~m[1970])|(~m[1928]&m[1929]&m[1930]&~m[1931]&~m[1970])|(m[1928]&m[1929]&m[1930]&~m[1931]&~m[1970])|(m[1928]&m[1929]&m[1930]&m[1931]&~m[1970])|(m[1928]&m[1929]&~m[1930]&~m[1931]&m[1970])|(m[1928]&~m[1929]&m[1930]&~m[1931]&m[1970])|(~m[1928]&m[1929]&m[1930]&~m[1931]&m[1970])|(m[1928]&m[1929]&m[1930]&~m[1931]&m[1970])|(m[1928]&m[1929]&m[1930]&m[1931]&m[1970]));
    m[1937] = (((m[1933]&~m[1934]&~m[1935]&~m[1936]&~m[1975])|(~m[1933]&m[1934]&~m[1935]&~m[1936]&~m[1975])|(~m[1933]&~m[1934]&m[1935]&~m[1936]&~m[1975])|(m[1933]&m[1934]&~m[1935]&m[1936]&~m[1975])|(m[1933]&~m[1934]&m[1935]&m[1936]&~m[1975])|(~m[1933]&m[1934]&m[1935]&m[1936]&~m[1975]))&BiasedRNG[1096])|(((m[1933]&~m[1934]&~m[1935]&~m[1936]&m[1975])|(~m[1933]&m[1934]&~m[1935]&~m[1936]&m[1975])|(~m[1933]&~m[1934]&m[1935]&~m[1936]&m[1975])|(m[1933]&m[1934]&~m[1935]&m[1936]&m[1975])|(m[1933]&~m[1934]&m[1935]&m[1936]&m[1975])|(~m[1933]&m[1934]&m[1935]&m[1936]&m[1975]))&~BiasedRNG[1096])|((m[1933]&m[1934]&~m[1935]&~m[1936]&~m[1975])|(m[1933]&~m[1934]&m[1935]&~m[1936]&~m[1975])|(~m[1933]&m[1934]&m[1935]&~m[1936]&~m[1975])|(m[1933]&m[1934]&m[1935]&~m[1936]&~m[1975])|(m[1933]&m[1934]&m[1935]&m[1936]&~m[1975])|(m[1933]&m[1934]&~m[1935]&~m[1936]&m[1975])|(m[1933]&~m[1934]&m[1935]&~m[1936]&m[1975])|(~m[1933]&m[1934]&m[1935]&~m[1936]&m[1975])|(m[1933]&m[1934]&m[1935]&~m[1936]&m[1975])|(m[1933]&m[1934]&m[1935]&m[1936]&m[1975]));
    m[1942] = (((m[1938]&~m[1939]&~m[1940]&~m[1941]&~m[1980])|(~m[1938]&m[1939]&~m[1940]&~m[1941]&~m[1980])|(~m[1938]&~m[1939]&m[1940]&~m[1941]&~m[1980])|(m[1938]&m[1939]&~m[1940]&m[1941]&~m[1980])|(m[1938]&~m[1939]&m[1940]&m[1941]&~m[1980])|(~m[1938]&m[1939]&m[1940]&m[1941]&~m[1980]))&BiasedRNG[1097])|(((m[1938]&~m[1939]&~m[1940]&~m[1941]&m[1980])|(~m[1938]&m[1939]&~m[1940]&~m[1941]&m[1980])|(~m[1938]&~m[1939]&m[1940]&~m[1941]&m[1980])|(m[1938]&m[1939]&~m[1940]&m[1941]&m[1980])|(m[1938]&~m[1939]&m[1940]&m[1941]&m[1980])|(~m[1938]&m[1939]&m[1940]&m[1941]&m[1980]))&~BiasedRNG[1097])|((m[1938]&m[1939]&~m[1940]&~m[1941]&~m[1980])|(m[1938]&~m[1939]&m[1940]&~m[1941]&~m[1980])|(~m[1938]&m[1939]&m[1940]&~m[1941]&~m[1980])|(m[1938]&m[1939]&m[1940]&~m[1941]&~m[1980])|(m[1938]&m[1939]&m[1940]&m[1941]&~m[1980])|(m[1938]&m[1939]&~m[1940]&~m[1941]&m[1980])|(m[1938]&~m[1939]&m[1940]&~m[1941]&m[1980])|(~m[1938]&m[1939]&m[1940]&~m[1941]&m[1980])|(m[1938]&m[1939]&m[1940]&~m[1941]&m[1980])|(m[1938]&m[1939]&m[1940]&m[1941]&m[1980]));
    m[1947] = (((m[1943]&~m[1944]&~m[1945]&~m[1946]&~m[1985])|(~m[1943]&m[1944]&~m[1945]&~m[1946]&~m[1985])|(~m[1943]&~m[1944]&m[1945]&~m[1946]&~m[1985])|(m[1943]&m[1944]&~m[1945]&m[1946]&~m[1985])|(m[1943]&~m[1944]&m[1945]&m[1946]&~m[1985])|(~m[1943]&m[1944]&m[1945]&m[1946]&~m[1985]))&BiasedRNG[1098])|(((m[1943]&~m[1944]&~m[1945]&~m[1946]&m[1985])|(~m[1943]&m[1944]&~m[1945]&~m[1946]&m[1985])|(~m[1943]&~m[1944]&m[1945]&~m[1946]&m[1985])|(m[1943]&m[1944]&~m[1945]&m[1946]&m[1985])|(m[1943]&~m[1944]&m[1945]&m[1946]&m[1985])|(~m[1943]&m[1944]&m[1945]&m[1946]&m[1985]))&~BiasedRNG[1098])|((m[1943]&m[1944]&~m[1945]&~m[1946]&~m[1985])|(m[1943]&~m[1944]&m[1945]&~m[1946]&~m[1985])|(~m[1943]&m[1944]&m[1945]&~m[1946]&~m[1985])|(m[1943]&m[1944]&m[1945]&~m[1946]&~m[1985])|(m[1943]&m[1944]&m[1945]&m[1946]&~m[1985])|(m[1943]&m[1944]&~m[1945]&~m[1946]&m[1985])|(m[1943]&~m[1944]&m[1945]&~m[1946]&m[1985])|(~m[1943]&m[1944]&m[1945]&~m[1946]&m[1985])|(m[1943]&m[1944]&m[1945]&~m[1946]&m[1985])|(m[1943]&m[1944]&m[1945]&m[1946]&m[1985]));
    m[1952] = (((m[1948]&~m[1949]&~m[1950]&~m[1951]&~m[1988])|(~m[1948]&m[1949]&~m[1950]&~m[1951]&~m[1988])|(~m[1948]&~m[1949]&m[1950]&~m[1951]&~m[1988])|(m[1948]&m[1949]&~m[1950]&m[1951]&~m[1988])|(m[1948]&~m[1949]&m[1950]&m[1951]&~m[1988])|(~m[1948]&m[1949]&m[1950]&m[1951]&~m[1988]))&BiasedRNG[1099])|(((m[1948]&~m[1949]&~m[1950]&~m[1951]&m[1988])|(~m[1948]&m[1949]&~m[1950]&~m[1951]&m[1988])|(~m[1948]&~m[1949]&m[1950]&~m[1951]&m[1988])|(m[1948]&m[1949]&~m[1950]&m[1951]&m[1988])|(m[1948]&~m[1949]&m[1950]&m[1951]&m[1988])|(~m[1948]&m[1949]&m[1950]&m[1951]&m[1988]))&~BiasedRNG[1099])|((m[1948]&m[1949]&~m[1950]&~m[1951]&~m[1988])|(m[1948]&~m[1949]&m[1950]&~m[1951]&~m[1988])|(~m[1948]&m[1949]&m[1950]&~m[1951]&~m[1988])|(m[1948]&m[1949]&m[1950]&~m[1951]&~m[1988])|(m[1948]&m[1949]&m[1950]&m[1951]&~m[1988])|(m[1948]&m[1949]&~m[1950]&~m[1951]&m[1988])|(m[1948]&~m[1949]&m[1950]&~m[1951]&m[1988])|(~m[1948]&m[1949]&m[1950]&~m[1951]&m[1988])|(m[1948]&m[1949]&m[1950]&~m[1951]&m[1988])|(m[1948]&m[1949]&m[1950]&m[1951]&m[1988]));
    m[1957] = (((m[1953]&~m[1954]&~m[1955]&~m[1956]&~m[1990])|(~m[1953]&m[1954]&~m[1955]&~m[1956]&~m[1990])|(~m[1953]&~m[1954]&m[1955]&~m[1956]&~m[1990])|(m[1953]&m[1954]&~m[1955]&m[1956]&~m[1990])|(m[1953]&~m[1954]&m[1955]&m[1956]&~m[1990])|(~m[1953]&m[1954]&m[1955]&m[1956]&~m[1990]))&BiasedRNG[1100])|(((m[1953]&~m[1954]&~m[1955]&~m[1956]&m[1990])|(~m[1953]&m[1954]&~m[1955]&~m[1956]&m[1990])|(~m[1953]&~m[1954]&m[1955]&~m[1956]&m[1990])|(m[1953]&m[1954]&~m[1955]&m[1956]&m[1990])|(m[1953]&~m[1954]&m[1955]&m[1956]&m[1990])|(~m[1953]&m[1954]&m[1955]&m[1956]&m[1990]))&~BiasedRNG[1100])|((m[1953]&m[1954]&~m[1955]&~m[1956]&~m[1990])|(m[1953]&~m[1954]&m[1955]&~m[1956]&~m[1990])|(~m[1953]&m[1954]&m[1955]&~m[1956]&~m[1990])|(m[1953]&m[1954]&m[1955]&~m[1956]&~m[1990])|(m[1953]&m[1954]&m[1955]&m[1956]&~m[1990])|(m[1953]&m[1954]&~m[1955]&~m[1956]&m[1990])|(m[1953]&~m[1954]&m[1955]&~m[1956]&m[1990])|(~m[1953]&m[1954]&m[1955]&~m[1956]&m[1990])|(m[1953]&m[1954]&m[1955]&~m[1956]&m[1990])|(m[1953]&m[1954]&m[1955]&m[1956]&m[1990]));
    m[1962] = (((m[1958]&~m[1959]&~m[1960]&~m[1961]&~m[1995])|(~m[1958]&m[1959]&~m[1960]&~m[1961]&~m[1995])|(~m[1958]&~m[1959]&m[1960]&~m[1961]&~m[1995])|(m[1958]&m[1959]&~m[1960]&m[1961]&~m[1995])|(m[1958]&~m[1959]&m[1960]&m[1961]&~m[1995])|(~m[1958]&m[1959]&m[1960]&m[1961]&~m[1995]))&BiasedRNG[1101])|(((m[1958]&~m[1959]&~m[1960]&~m[1961]&m[1995])|(~m[1958]&m[1959]&~m[1960]&~m[1961]&m[1995])|(~m[1958]&~m[1959]&m[1960]&~m[1961]&m[1995])|(m[1958]&m[1959]&~m[1960]&m[1961]&m[1995])|(m[1958]&~m[1959]&m[1960]&m[1961]&m[1995])|(~m[1958]&m[1959]&m[1960]&m[1961]&m[1995]))&~BiasedRNG[1101])|((m[1958]&m[1959]&~m[1960]&~m[1961]&~m[1995])|(m[1958]&~m[1959]&m[1960]&~m[1961]&~m[1995])|(~m[1958]&m[1959]&m[1960]&~m[1961]&~m[1995])|(m[1958]&m[1959]&m[1960]&~m[1961]&~m[1995])|(m[1958]&m[1959]&m[1960]&m[1961]&~m[1995])|(m[1958]&m[1959]&~m[1960]&~m[1961]&m[1995])|(m[1958]&~m[1959]&m[1960]&~m[1961]&m[1995])|(~m[1958]&m[1959]&m[1960]&~m[1961]&m[1995])|(m[1958]&m[1959]&m[1960]&~m[1961]&m[1995])|(m[1958]&m[1959]&m[1960]&m[1961]&m[1995]));
    m[1967] = (((m[1963]&~m[1964]&~m[1965]&~m[1966]&~m[2000])|(~m[1963]&m[1964]&~m[1965]&~m[1966]&~m[2000])|(~m[1963]&~m[1964]&m[1965]&~m[1966]&~m[2000])|(m[1963]&m[1964]&~m[1965]&m[1966]&~m[2000])|(m[1963]&~m[1964]&m[1965]&m[1966]&~m[2000])|(~m[1963]&m[1964]&m[1965]&m[1966]&~m[2000]))&BiasedRNG[1102])|(((m[1963]&~m[1964]&~m[1965]&~m[1966]&m[2000])|(~m[1963]&m[1964]&~m[1965]&~m[1966]&m[2000])|(~m[1963]&~m[1964]&m[1965]&~m[1966]&m[2000])|(m[1963]&m[1964]&~m[1965]&m[1966]&m[2000])|(m[1963]&~m[1964]&m[1965]&m[1966]&m[2000])|(~m[1963]&m[1964]&m[1965]&m[1966]&m[2000]))&~BiasedRNG[1102])|((m[1963]&m[1964]&~m[1965]&~m[1966]&~m[2000])|(m[1963]&~m[1964]&m[1965]&~m[1966]&~m[2000])|(~m[1963]&m[1964]&m[1965]&~m[1966]&~m[2000])|(m[1963]&m[1964]&m[1965]&~m[1966]&~m[2000])|(m[1963]&m[1964]&m[1965]&m[1966]&~m[2000])|(m[1963]&m[1964]&~m[1965]&~m[1966]&m[2000])|(m[1963]&~m[1964]&m[1965]&~m[1966]&m[2000])|(~m[1963]&m[1964]&m[1965]&~m[1966]&m[2000])|(m[1963]&m[1964]&m[1965]&~m[1966]&m[2000])|(m[1963]&m[1964]&m[1965]&m[1966]&m[2000]));
    m[1972] = (((m[1968]&~m[1969]&~m[1970]&~m[1971]&~m[2005])|(~m[1968]&m[1969]&~m[1970]&~m[1971]&~m[2005])|(~m[1968]&~m[1969]&m[1970]&~m[1971]&~m[2005])|(m[1968]&m[1969]&~m[1970]&m[1971]&~m[2005])|(m[1968]&~m[1969]&m[1970]&m[1971]&~m[2005])|(~m[1968]&m[1969]&m[1970]&m[1971]&~m[2005]))&BiasedRNG[1103])|(((m[1968]&~m[1969]&~m[1970]&~m[1971]&m[2005])|(~m[1968]&m[1969]&~m[1970]&~m[1971]&m[2005])|(~m[1968]&~m[1969]&m[1970]&~m[1971]&m[2005])|(m[1968]&m[1969]&~m[1970]&m[1971]&m[2005])|(m[1968]&~m[1969]&m[1970]&m[1971]&m[2005])|(~m[1968]&m[1969]&m[1970]&m[1971]&m[2005]))&~BiasedRNG[1103])|((m[1968]&m[1969]&~m[1970]&~m[1971]&~m[2005])|(m[1968]&~m[1969]&m[1970]&~m[1971]&~m[2005])|(~m[1968]&m[1969]&m[1970]&~m[1971]&~m[2005])|(m[1968]&m[1969]&m[1970]&~m[1971]&~m[2005])|(m[1968]&m[1969]&m[1970]&m[1971]&~m[2005])|(m[1968]&m[1969]&~m[1970]&~m[1971]&m[2005])|(m[1968]&~m[1969]&m[1970]&~m[1971]&m[2005])|(~m[1968]&m[1969]&m[1970]&~m[1971]&m[2005])|(m[1968]&m[1969]&m[1970]&~m[1971]&m[2005])|(m[1968]&m[1969]&m[1970]&m[1971]&m[2005]));
    m[1977] = (((m[1973]&~m[1974]&~m[1975]&~m[1976]&~m[2010])|(~m[1973]&m[1974]&~m[1975]&~m[1976]&~m[2010])|(~m[1973]&~m[1974]&m[1975]&~m[1976]&~m[2010])|(m[1973]&m[1974]&~m[1975]&m[1976]&~m[2010])|(m[1973]&~m[1974]&m[1975]&m[1976]&~m[2010])|(~m[1973]&m[1974]&m[1975]&m[1976]&~m[2010]))&BiasedRNG[1104])|(((m[1973]&~m[1974]&~m[1975]&~m[1976]&m[2010])|(~m[1973]&m[1974]&~m[1975]&~m[1976]&m[2010])|(~m[1973]&~m[1974]&m[1975]&~m[1976]&m[2010])|(m[1973]&m[1974]&~m[1975]&m[1976]&m[2010])|(m[1973]&~m[1974]&m[1975]&m[1976]&m[2010])|(~m[1973]&m[1974]&m[1975]&m[1976]&m[2010]))&~BiasedRNG[1104])|((m[1973]&m[1974]&~m[1975]&~m[1976]&~m[2010])|(m[1973]&~m[1974]&m[1975]&~m[1976]&~m[2010])|(~m[1973]&m[1974]&m[1975]&~m[1976]&~m[2010])|(m[1973]&m[1974]&m[1975]&~m[1976]&~m[2010])|(m[1973]&m[1974]&m[1975]&m[1976]&~m[2010])|(m[1973]&m[1974]&~m[1975]&~m[1976]&m[2010])|(m[1973]&~m[1974]&m[1975]&~m[1976]&m[2010])|(~m[1973]&m[1974]&m[1975]&~m[1976]&m[2010])|(m[1973]&m[1974]&m[1975]&~m[1976]&m[2010])|(m[1973]&m[1974]&m[1975]&m[1976]&m[2010]));
    m[1982] = (((m[1978]&~m[1979]&~m[1980]&~m[1981]&~m[2015])|(~m[1978]&m[1979]&~m[1980]&~m[1981]&~m[2015])|(~m[1978]&~m[1979]&m[1980]&~m[1981]&~m[2015])|(m[1978]&m[1979]&~m[1980]&m[1981]&~m[2015])|(m[1978]&~m[1979]&m[1980]&m[1981]&~m[2015])|(~m[1978]&m[1979]&m[1980]&m[1981]&~m[2015]))&BiasedRNG[1105])|(((m[1978]&~m[1979]&~m[1980]&~m[1981]&m[2015])|(~m[1978]&m[1979]&~m[1980]&~m[1981]&m[2015])|(~m[1978]&~m[1979]&m[1980]&~m[1981]&m[2015])|(m[1978]&m[1979]&~m[1980]&m[1981]&m[2015])|(m[1978]&~m[1979]&m[1980]&m[1981]&m[2015])|(~m[1978]&m[1979]&m[1980]&m[1981]&m[2015]))&~BiasedRNG[1105])|((m[1978]&m[1979]&~m[1980]&~m[1981]&~m[2015])|(m[1978]&~m[1979]&m[1980]&~m[1981]&~m[2015])|(~m[1978]&m[1979]&m[1980]&~m[1981]&~m[2015])|(m[1978]&m[1979]&m[1980]&~m[1981]&~m[2015])|(m[1978]&m[1979]&m[1980]&m[1981]&~m[2015])|(m[1978]&m[1979]&~m[1980]&~m[1981]&m[2015])|(m[1978]&~m[1979]&m[1980]&~m[1981]&m[2015])|(~m[1978]&m[1979]&m[1980]&~m[1981]&m[2015])|(m[1978]&m[1979]&m[1980]&~m[1981]&m[2015])|(m[1978]&m[1979]&m[1980]&m[1981]&m[2015]));
    m[1987] = (((m[1983]&~m[1984]&~m[1985]&~m[1986]&~m[2020])|(~m[1983]&m[1984]&~m[1985]&~m[1986]&~m[2020])|(~m[1983]&~m[1984]&m[1985]&~m[1986]&~m[2020])|(m[1983]&m[1984]&~m[1985]&m[1986]&~m[2020])|(m[1983]&~m[1984]&m[1985]&m[1986]&~m[2020])|(~m[1983]&m[1984]&m[1985]&m[1986]&~m[2020]))&BiasedRNG[1106])|(((m[1983]&~m[1984]&~m[1985]&~m[1986]&m[2020])|(~m[1983]&m[1984]&~m[1985]&~m[1986]&m[2020])|(~m[1983]&~m[1984]&m[1985]&~m[1986]&m[2020])|(m[1983]&m[1984]&~m[1985]&m[1986]&m[2020])|(m[1983]&~m[1984]&m[1985]&m[1986]&m[2020])|(~m[1983]&m[1984]&m[1985]&m[1986]&m[2020]))&~BiasedRNG[1106])|((m[1983]&m[1984]&~m[1985]&~m[1986]&~m[2020])|(m[1983]&~m[1984]&m[1985]&~m[1986]&~m[2020])|(~m[1983]&m[1984]&m[1985]&~m[1986]&~m[2020])|(m[1983]&m[1984]&m[1985]&~m[1986]&~m[2020])|(m[1983]&m[1984]&m[1985]&m[1986]&~m[2020])|(m[1983]&m[1984]&~m[1985]&~m[1986]&m[2020])|(m[1983]&~m[1984]&m[1985]&~m[1986]&m[2020])|(~m[1983]&m[1984]&m[1985]&~m[1986]&m[2020])|(m[1983]&m[1984]&m[1985]&~m[1986]&m[2020])|(m[1983]&m[1984]&m[1985]&m[1986]&m[2020]));
    m[1992] = (((m[1988]&~m[1989]&~m[1990]&~m[1991]&~m[2023])|(~m[1988]&m[1989]&~m[1990]&~m[1991]&~m[2023])|(~m[1988]&~m[1989]&m[1990]&~m[1991]&~m[2023])|(m[1988]&m[1989]&~m[1990]&m[1991]&~m[2023])|(m[1988]&~m[1989]&m[1990]&m[1991]&~m[2023])|(~m[1988]&m[1989]&m[1990]&m[1991]&~m[2023]))&BiasedRNG[1107])|(((m[1988]&~m[1989]&~m[1990]&~m[1991]&m[2023])|(~m[1988]&m[1989]&~m[1990]&~m[1991]&m[2023])|(~m[1988]&~m[1989]&m[1990]&~m[1991]&m[2023])|(m[1988]&m[1989]&~m[1990]&m[1991]&m[2023])|(m[1988]&~m[1989]&m[1990]&m[1991]&m[2023])|(~m[1988]&m[1989]&m[1990]&m[1991]&m[2023]))&~BiasedRNG[1107])|((m[1988]&m[1989]&~m[1990]&~m[1991]&~m[2023])|(m[1988]&~m[1989]&m[1990]&~m[1991]&~m[2023])|(~m[1988]&m[1989]&m[1990]&~m[1991]&~m[2023])|(m[1988]&m[1989]&m[1990]&~m[1991]&~m[2023])|(m[1988]&m[1989]&m[1990]&m[1991]&~m[2023])|(m[1988]&m[1989]&~m[1990]&~m[1991]&m[2023])|(m[1988]&~m[1989]&m[1990]&~m[1991]&m[2023])|(~m[1988]&m[1989]&m[1990]&~m[1991]&m[2023])|(m[1988]&m[1989]&m[1990]&~m[1991]&m[2023])|(m[1988]&m[1989]&m[1990]&m[1991]&m[2023]));
    m[1997] = (((m[1993]&~m[1994]&~m[1995]&~m[1996]&~m[2025])|(~m[1993]&m[1994]&~m[1995]&~m[1996]&~m[2025])|(~m[1993]&~m[1994]&m[1995]&~m[1996]&~m[2025])|(m[1993]&m[1994]&~m[1995]&m[1996]&~m[2025])|(m[1993]&~m[1994]&m[1995]&m[1996]&~m[2025])|(~m[1993]&m[1994]&m[1995]&m[1996]&~m[2025]))&BiasedRNG[1108])|(((m[1993]&~m[1994]&~m[1995]&~m[1996]&m[2025])|(~m[1993]&m[1994]&~m[1995]&~m[1996]&m[2025])|(~m[1993]&~m[1994]&m[1995]&~m[1996]&m[2025])|(m[1993]&m[1994]&~m[1995]&m[1996]&m[2025])|(m[1993]&~m[1994]&m[1995]&m[1996]&m[2025])|(~m[1993]&m[1994]&m[1995]&m[1996]&m[2025]))&~BiasedRNG[1108])|((m[1993]&m[1994]&~m[1995]&~m[1996]&~m[2025])|(m[1993]&~m[1994]&m[1995]&~m[1996]&~m[2025])|(~m[1993]&m[1994]&m[1995]&~m[1996]&~m[2025])|(m[1993]&m[1994]&m[1995]&~m[1996]&~m[2025])|(m[1993]&m[1994]&m[1995]&m[1996]&~m[2025])|(m[1993]&m[1994]&~m[1995]&~m[1996]&m[2025])|(m[1993]&~m[1994]&m[1995]&~m[1996]&m[2025])|(~m[1993]&m[1994]&m[1995]&~m[1996]&m[2025])|(m[1993]&m[1994]&m[1995]&~m[1996]&m[2025])|(m[1993]&m[1994]&m[1995]&m[1996]&m[2025]));
    m[2002] = (((m[1998]&~m[1999]&~m[2000]&~m[2001]&~m[2030])|(~m[1998]&m[1999]&~m[2000]&~m[2001]&~m[2030])|(~m[1998]&~m[1999]&m[2000]&~m[2001]&~m[2030])|(m[1998]&m[1999]&~m[2000]&m[2001]&~m[2030])|(m[1998]&~m[1999]&m[2000]&m[2001]&~m[2030])|(~m[1998]&m[1999]&m[2000]&m[2001]&~m[2030]))&BiasedRNG[1109])|(((m[1998]&~m[1999]&~m[2000]&~m[2001]&m[2030])|(~m[1998]&m[1999]&~m[2000]&~m[2001]&m[2030])|(~m[1998]&~m[1999]&m[2000]&~m[2001]&m[2030])|(m[1998]&m[1999]&~m[2000]&m[2001]&m[2030])|(m[1998]&~m[1999]&m[2000]&m[2001]&m[2030])|(~m[1998]&m[1999]&m[2000]&m[2001]&m[2030]))&~BiasedRNG[1109])|((m[1998]&m[1999]&~m[2000]&~m[2001]&~m[2030])|(m[1998]&~m[1999]&m[2000]&~m[2001]&~m[2030])|(~m[1998]&m[1999]&m[2000]&~m[2001]&~m[2030])|(m[1998]&m[1999]&m[2000]&~m[2001]&~m[2030])|(m[1998]&m[1999]&m[2000]&m[2001]&~m[2030])|(m[1998]&m[1999]&~m[2000]&~m[2001]&m[2030])|(m[1998]&~m[1999]&m[2000]&~m[2001]&m[2030])|(~m[1998]&m[1999]&m[2000]&~m[2001]&m[2030])|(m[1998]&m[1999]&m[2000]&~m[2001]&m[2030])|(m[1998]&m[1999]&m[2000]&m[2001]&m[2030]));
    m[2007] = (((m[2003]&~m[2004]&~m[2005]&~m[2006]&~m[2035])|(~m[2003]&m[2004]&~m[2005]&~m[2006]&~m[2035])|(~m[2003]&~m[2004]&m[2005]&~m[2006]&~m[2035])|(m[2003]&m[2004]&~m[2005]&m[2006]&~m[2035])|(m[2003]&~m[2004]&m[2005]&m[2006]&~m[2035])|(~m[2003]&m[2004]&m[2005]&m[2006]&~m[2035]))&BiasedRNG[1110])|(((m[2003]&~m[2004]&~m[2005]&~m[2006]&m[2035])|(~m[2003]&m[2004]&~m[2005]&~m[2006]&m[2035])|(~m[2003]&~m[2004]&m[2005]&~m[2006]&m[2035])|(m[2003]&m[2004]&~m[2005]&m[2006]&m[2035])|(m[2003]&~m[2004]&m[2005]&m[2006]&m[2035])|(~m[2003]&m[2004]&m[2005]&m[2006]&m[2035]))&~BiasedRNG[1110])|((m[2003]&m[2004]&~m[2005]&~m[2006]&~m[2035])|(m[2003]&~m[2004]&m[2005]&~m[2006]&~m[2035])|(~m[2003]&m[2004]&m[2005]&~m[2006]&~m[2035])|(m[2003]&m[2004]&m[2005]&~m[2006]&~m[2035])|(m[2003]&m[2004]&m[2005]&m[2006]&~m[2035])|(m[2003]&m[2004]&~m[2005]&~m[2006]&m[2035])|(m[2003]&~m[2004]&m[2005]&~m[2006]&m[2035])|(~m[2003]&m[2004]&m[2005]&~m[2006]&m[2035])|(m[2003]&m[2004]&m[2005]&~m[2006]&m[2035])|(m[2003]&m[2004]&m[2005]&m[2006]&m[2035]));
    m[2012] = (((m[2008]&~m[2009]&~m[2010]&~m[2011]&~m[2040])|(~m[2008]&m[2009]&~m[2010]&~m[2011]&~m[2040])|(~m[2008]&~m[2009]&m[2010]&~m[2011]&~m[2040])|(m[2008]&m[2009]&~m[2010]&m[2011]&~m[2040])|(m[2008]&~m[2009]&m[2010]&m[2011]&~m[2040])|(~m[2008]&m[2009]&m[2010]&m[2011]&~m[2040]))&BiasedRNG[1111])|(((m[2008]&~m[2009]&~m[2010]&~m[2011]&m[2040])|(~m[2008]&m[2009]&~m[2010]&~m[2011]&m[2040])|(~m[2008]&~m[2009]&m[2010]&~m[2011]&m[2040])|(m[2008]&m[2009]&~m[2010]&m[2011]&m[2040])|(m[2008]&~m[2009]&m[2010]&m[2011]&m[2040])|(~m[2008]&m[2009]&m[2010]&m[2011]&m[2040]))&~BiasedRNG[1111])|((m[2008]&m[2009]&~m[2010]&~m[2011]&~m[2040])|(m[2008]&~m[2009]&m[2010]&~m[2011]&~m[2040])|(~m[2008]&m[2009]&m[2010]&~m[2011]&~m[2040])|(m[2008]&m[2009]&m[2010]&~m[2011]&~m[2040])|(m[2008]&m[2009]&m[2010]&m[2011]&~m[2040])|(m[2008]&m[2009]&~m[2010]&~m[2011]&m[2040])|(m[2008]&~m[2009]&m[2010]&~m[2011]&m[2040])|(~m[2008]&m[2009]&m[2010]&~m[2011]&m[2040])|(m[2008]&m[2009]&m[2010]&~m[2011]&m[2040])|(m[2008]&m[2009]&m[2010]&m[2011]&m[2040]));
    m[2017] = (((m[2013]&~m[2014]&~m[2015]&~m[2016]&~m[2045])|(~m[2013]&m[2014]&~m[2015]&~m[2016]&~m[2045])|(~m[2013]&~m[2014]&m[2015]&~m[2016]&~m[2045])|(m[2013]&m[2014]&~m[2015]&m[2016]&~m[2045])|(m[2013]&~m[2014]&m[2015]&m[2016]&~m[2045])|(~m[2013]&m[2014]&m[2015]&m[2016]&~m[2045]))&BiasedRNG[1112])|(((m[2013]&~m[2014]&~m[2015]&~m[2016]&m[2045])|(~m[2013]&m[2014]&~m[2015]&~m[2016]&m[2045])|(~m[2013]&~m[2014]&m[2015]&~m[2016]&m[2045])|(m[2013]&m[2014]&~m[2015]&m[2016]&m[2045])|(m[2013]&~m[2014]&m[2015]&m[2016]&m[2045])|(~m[2013]&m[2014]&m[2015]&m[2016]&m[2045]))&~BiasedRNG[1112])|((m[2013]&m[2014]&~m[2015]&~m[2016]&~m[2045])|(m[2013]&~m[2014]&m[2015]&~m[2016]&~m[2045])|(~m[2013]&m[2014]&m[2015]&~m[2016]&~m[2045])|(m[2013]&m[2014]&m[2015]&~m[2016]&~m[2045])|(m[2013]&m[2014]&m[2015]&m[2016]&~m[2045])|(m[2013]&m[2014]&~m[2015]&~m[2016]&m[2045])|(m[2013]&~m[2014]&m[2015]&~m[2016]&m[2045])|(~m[2013]&m[2014]&m[2015]&~m[2016]&m[2045])|(m[2013]&m[2014]&m[2015]&~m[2016]&m[2045])|(m[2013]&m[2014]&m[2015]&m[2016]&m[2045]));
    m[2022] = (((m[2018]&~m[2019]&~m[2020]&~m[2021]&~m[2050])|(~m[2018]&m[2019]&~m[2020]&~m[2021]&~m[2050])|(~m[2018]&~m[2019]&m[2020]&~m[2021]&~m[2050])|(m[2018]&m[2019]&~m[2020]&m[2021]&~m[2050])|(m[2018]&~m[2019]&m[2020]&m[2021]&~m[2050])|(~m[2018]&m[2019]&m[2020]&m[2021]&~m[2050]))&BiasedRNG[1113])|(((m[2018]&~m[2019]&~m[2020]&~m[2021]&m[2050])|(~m[2018]&m[2019]&~m[2020]&~m[2021]&m[2050])|(~m[2018]&~m[2019]&m[2020]&~m[2021]&m[2050])|(m[2018]&m[2019]&~m[2020]&m[2021]&m[2050])|(m[2018]&~m[2019]&m[2020]&m[2021]&m[2050])|(~m[2018]&m[2019]&m[2020]&m[2021]&m[2050]))&~BiasedRNG[1113])|((m[2018]&m[2019]&~m[2020]&~m[2021]&~m[2050])|(m[2018]&~m[2019]&m[2020]&~m[2021]&~m[2050])|(~m[2018]&m[2019]&m[2020]&~m[2021]&~m[2050])|(m[2018]&m[2019]&m[2020]&~m[2021]&~m[2050])|(m[2018]&m[2019]&m[2020]&m[2021]&~m[2050])|(m[2018]&m[2019]&~m[2020]&~m[2021]&m[2050])|(m[2018]&~m[2019]&m[2020]&~m[2021]&m[2050])|(~m[2018]&m[2019]&m[2020]&~m[2021]&m[2050])|(m[2018]&m[2019]&m[2020]&~m[2021]&m[2050])|(m[2018]&m[2019]&m[2020]&m[2021]&m[2050]));
    m[2027] = (((m[2023]&~m[2024]&~m[2025]&~m[2026]&~m[2053])|(~m[2023]&m[2024]&~m[2025]&~m[2026]&~m[2053])|(~m[2023]&~m[2024]&m[2025]&~m[2026]&~m[2053])|(m[2023]&m[2024]&~m[2025]&m[2026]&~m[2053])|(m[2023]&~m[2024]&m[2025]&m[2026]&~m[2053])|(~m[2023]&m[2024]&m[2025]&m[2026]&~m[2053]))&BiasedRNG[1114])|(((m[2023]&~m[2024]&~m[2025]&~m[2026]&m[2053])|(~m[2023]&m[2024]&~m[2025]&~m[2026]&m[2053])|(~m[2023]&~m[2024]&m[2025]&~m[2026]&m[2053])|(m[2023]&m[2024]&~m[2025]&m[2026]&m[2053])|(m[2023]&~m[2024]&m[2025]&m[2026]&m[2053])|(~m[2023]&m[2024]&m[2025]&m[2026]&m[2053]))&~BiasedRNG[1114])|((m[2023]&m[2024]&~m[2025]&~m[2026]&~m[2053])|(m[2023]&~m[2024]&m[2025]&~m[2026]&~m[2053])|(~m[2023]&m[2024]&m[2025]&~m[2026]&~m[2053])|(m[2023]&m[2024]&m[2025]&~m[2026]&~m[2053])|(m[2023]&m[2024]&m[2025]&m[2026]&~m[2053])|(m[2023]&m[2024]&~m[2025]&~m[2026]&m[2053])|(m[2023]&~m[2024]&m[2025]&~m[2026]&m[2053])|(~m[2023]&m[2024]&m[2025]&~m[2026]&m[2053])|(m[2023]&m[2024]&m[2025]&~m[2026]&m[2053])|(m[2023]&m[2024]&m[2025]&m[2026]&m[2053]));
    m[2032] = (((m[2028]&~m[2029]&~m[2030]&~m[2031]&~m[2055])|(~m[2028]&m[2029]&~m[2030]&~m[2031]&~m[2055])|(~m[2028]&~m[2029]&m[2030]&~m[2031]&~m[2055])|(m[2028]&m[2029]&~m[2030]&m[2031]&~m[2055])|(m[2028]&~m[2029]&m[2030]&m[2031]&~m[2055])|(~m[2028]&m[2029]&m[2030]&m[2031]&~m[2055]))&BiasedRNG[1115])|(((m[2028]&~m[2029]&~m[2030]&~m[2031]&m[2055])|(~m[2028]&m[2029]&~m[2030]&~m[2031]&m[2055])|(~m[2028]&~m[2029]&m[2030]&~m[2031]&m[2055])|(m[2028]&m[2029]&~m[2030]&m[2031]&m[2055])|(m[2028]&~m[2029]&m[2030]&m[2031]&m[2055])|(~m[2028]&m[2029]&m[2030]&m[2031]&m[2055]))&~BiasedRNG[1115])|((m[2028]&m[2029]&~m[2030]&~m[2031]&~m[2055])|(m[2028]&~m[2029]&m[2030]&~m[2031]&~m[2055])|(~m[2028]&m[2029]&m[2030]&~m[2031]&~m[2055])|(m[2028]&m[2029]&m[2030]&~m[2031]&~m[2055])|(m[2028]&m[2029]&m[2030]&m[2031]&~m[2055])|(m[2028]&m[2029]&~m[2030]&~m[2031]&m[2055])|(m[2028]&~m[2029]&m[2030]&~m[2031]&m[2055])|(~m[2028]&m[2029]&m[2030]&~m[2031]&m[2055])|(m[2028]&m[2029]&m[2030]&~m[2031]&m[2055])|(m[2028]&m[2029]&m[2030]&m[2031]&m[2055]));
    m[2037] = (((m[2033]&~m[2034]&~m[2035]&~m[2036]&~m[2060])|(~m[2033]&m[2034]&~m[2035]&~m[2036]&~m[2060])|(~m[2033]&~m[2034]&m[2035]&~m[2036]&~m[2060])|(m[2033]&m[2034]&~m[2035]&m[2036]&~m[2060])|(m[2033]&~m[2034]&m[2035]&m[2036]&~m[2060])|(~m[2033]&m[2034]&m[2035]&m[2036]&~m[2060]))&BiasedRNG[1116])|(((m[2033]&~m[2034]&~m[2035]&~m[2036]&m[2060])|(~m[2033]&m[2034]&~m[2035]&~m[2036]&m[2060])|(~m[2033]&~m[2034]&m[2035]&~m[2036]&m[2060])|(m[2033]&m[2034]&~m[2035]&m[2036]&m[2060])|(m[2033]&~m[2034]&m[2035]&m[2036]&m[2060])|(~m[2033]&m[2034]&m[2035]&m[2036]&m[2060]))&~BiasedRNG[1116])|((m[2033]&m[2034]&~m[2035]&~m[2036]&~m[2060])|(m[2033]&~m[2034]&m[2035]&~m[2036]&~m[2060])|(~m[2033]&m[2034]&m[2035]&~m[2036]&~m[2060])|(m[2033]&m[2034]&m[2035]&~m[2036]&~m[2060])|(m[2033]&m[2034]&m[2035]&m[2036]&~m[2060])|(m[2033]&m[2034]&~m[2035]&~m[2036]&m[2060])|(m[2033]&~m[2034]&m[2035]&~m[2036]&m[2060])|(~m[2033]&m[2034]&m[2035]&~m[2036]&m[2060])|(m[2033]&m[2034]&m[2035]&~m[2036]&m[2060])|(m[2033]&m[2034]&m[2035]&m[2036]&m[2060]));
    m[2042] = (((m[2038]&~m[2039]&~m[2040]&~m[2041]&~m[2065])|(~m[2038]&m[2039]&~m[2040]&~m[2041]&~m[2065])|(~m[2038]&~m[2039]&m[2040]&~m[2041]&~m[2065])|(m[2038]&m[2039]&~m[2040]&m[2041]&~m[2065])|(m[2038]&~m[2039]&m[2040]&m[2041]&~m[2065])|(~m[2038]&m[2039]&m[2040]&m[2041]&~m[2065]))&BiasedRNG[1117])|(((m[2038]&~m[2039]&~m[2040]&~m[2041]&m[2065])|(~m[2038]&m[2039]&~m[2040]&~m[2041]&m[2065])|(~m[2038]&~m[2039]&m[2040]&~m[2041]&m[2065])|(m[2038]&m[2039]&~m[2040]&m[2041]&m[2065])|(m[2038]&~m[2039]&m[2040]&m[2041]&m[2065])|(~m[2038]&m[2039]&m[2040]&m[2041]&m[2065]))&~BiasedRNG[1117])|((m[2038]&m[2039]&~m[2040]&~m[2041]&~m[2065])|(m[2038]&~m[2039]&m[2040]&~m[2041]&~m[2065])|(~m[2038]&m[2039]&m[2040]&~m[2041]&~m[2065])|(m[2038]&m[2039]&m[2040]&~m[2041]&~m[2065])|(m[2038]&m[2039]&m[2040]&m[2041]&~m[2065])|(m[2038]&m[2039]&~m[2040]&~m[2041]&m[2065])|(m[2038]&~m[2039]&m[2040]&~m[2041]&m[2065])|(~m[2038]&m[2039]&m[2040]&~m[2041]&m[2065])|(m[2038]&m[2039]&m[2040]&~m[2041]&m[2065])|(m[2038]&m[2039]&m[2040]&m[2041]&m[2065]));
    m[2047] = (((m[2043]&~m[2044]&~m[2045]&~m[2046]&~m[2070])|(~m[2043]&m[2044]&~m[2045]&~m[2046]&~m[2070])|(~m[2043]&~m[2044]&m[2045]&~m[2046]&~m[2070])|(m[2043]&m[2044]&~m[2045]&m[2046]&~m[2070])|(m[2043]&~m[2044]&m[2045]&m[2046]&~m[2070])|(~m[2043]&m[2044]&m[2045]&m[2046]&~m[2070]))&BiasedRNG[1118])|(((m[2043]&~m[2044]&~m[2045]&~m[2046]&m[2070])|(~m[2043]&m[2044]&~m[2045]&~m[2046]&m[2070])|(~m[2043]&~m[2044]&m[2045]&~m[2046]&m[2070])|(m[2043]&m[2044]&~m[2045]&m[2046]&m[2070])|(m[2043]&~m[2044]&m[2045]&m[2046]&m[2070])|(~m[2043]&m[2044]&m[2045]&m[2046]&m[2070]))&~BiasedRNG[1118])|((m[2043]&m[2044]&~m[2045]&~m[2046]&~m[2070])|(m[2043]&~m[2044]&m[2045]&~m[2046]&~m[2070])|(~m[2043]&m[2044]&m[2045]&~m[2046]&~m[2070])|(m[2043]&m[2044]&m[2045]&~m[2046]&~m[2070])|(m[2043]&m[2044]&m[2045]&m[2046]&~m[2070])|(m[2043]&m[2044]&~m[2045]&~m[2046]&m[2070])|(m[2043]&~m[2044]&m[2045]&~m[2046]&m[2070])|(~m[2043]&m[2044]&m[2045]&~m[2046]&m[2070])|(m[2043]&m[2044]&m[2045]&~m[2046]&m[2070])|(m[2043]&m[2044]&m[2045]&m[2046]&m[2070]));
    m[2052] = (((m[2048]&~m[2049]&~m[2050]&~m[2051]&~m[2075])|(~m[2048]&m[2049]&~m[2050]&~m[2051]&~m[2075])|(~m[2048]&~m[2049]&m[2050]&~m[2051]&~m[2075])|(m[2048]&m[2049]&~m[2050]&m[2051]&~m[2075])|(m[2048]&~m[2049]&m[2050]&m[2051]&~m[2075])|(~m[2048]&m[2049]&m[2050]&m[2051]&~m[2075]))&BiasedRNG[1119])|(((m[2048]&~m[2049]&~m[2050]&~m[2051]&m[2075])|(~m[2048]&m[2049]&~m[2050]&~m[2051]&m[2075])|(~m[2048]&~m[2049]&m[2050]&~m[2051]&m[2075])|(m[2048]&m[2049]&~m[2050]&m[2051]&m[2075])|(m[2048]&~m[2049]&m[2050]&m[2051]&m[2075])|(~m[2048]&m[2049]&m[2050]&m[2051]&m[2075]))&~BiasedRNG[1119])|((m[2048]&m[2049]&~m[2050]&~m[2051]&~m[2075])|(m[2048]&~m[2049]&m[2050]&~m[2051]&~m[2075])|(~m[2048]&m[2049]&m[2050]&~m[2051]&~m[2075])|(m[2048]&m[2049]&m[2050]&~m[2051]&~m[2075])|(m[2048]&m[2049]&m[2050]&m[2051]&~m[2075])|(m[2048]&m[2049]&~m[2050]&~m[2051]&m[2075])|(m[2048]&~m[2049]&m[2050]&~m[2051]&m[2075])|(~m[2048]&m[2049]&m[2050]&~m[2051]&m[2075])|(m[2048]&m[2049]&m[2050]&~m[2051]&m[2075])|(m[2048]&m[2049]&m[2050]&m[2051]&m[2075]));
    m[2057] = (((m[2053]&~m[2054]&~m[2055]&~m[2056]&~m[2078])|(~m[2053]&m[2054]&~m[2055]&~m[2056]&~m[2078])|(~m[2053]&~m[2054]&m[2055]&~m[2056]&~m[2078])|(m[2053]&m[2054]&~m[2055]&m[2056]&~m[2078])|(m[2053]&~m[2054]&m[2055]&m[2056]&~m[2078])|(~m[2053]&m[2054]&m[2055]&m[2056]&~m[2078]))&BiasedRNG[1120])|(((m[2053]&~m[2054]&~m[2055]&~m[2056]&m[2078])|(~m[2053]&m[2054]&~m[2055]&~m[2056]&m[2078])|(~m[2053]&~m[2054]&m[2055]&~m[2056]&m[2078])|(m[2053]&m[2054]&~m[2055]&m[2056]&m[2078])|(m[2053]&~m[2054]&m[2055]&m[2056]&m[2078])|(~m[2053]&m[2054]&m[2055]&m[2056]&m[2078]))&~BiasedRNG[1120])|((m[2053]&m[2054]&~m[2055]&~m[2056]&~m[2078])|(m[2053]&~m[2054]&m[2055]&~m[2056]&~m[2078])|(~m[2053]&m[2054]&m[2055]&~m[2056]&~m[2078])|(m[2053]&m[2054]&m[2055]&~m[2056]&~m[2078])|(m[2053]&m[2054]&m[2055]&m[2056]&~m[2078])|(m[2053]&m[2054]&~m[2055]&~m[2056]&m[2078])|(m[2053]&~m[2054]&m[2055]&~m[2056]&m[2078])|(~m[2053]&m[2054]&m[2055]&~m[2056]&m[2078])|(m[2053]&m[2054]&m[2055]&~m[2056]&m[2078])|(m[2053]&m[2054]&m[2055]&m[2056]&m[2078]));
    m[2062] = (((m[2058]&~m[2059]&~m[2060]&~m[2061]&~m[2080])|(~m[2058]&m[2059]&~m[2060]&~m[2061]&~m[2080])|(~m[2058]&~m[2059]&m[2060]&~m[2061]&~m[2080])|(m[2058]&m[2059]&~m[2060]&m[2061]&~m[2080])|(m[2058]&~m[2059]&m[2060]&m[2061]&~m[2080])|(~m[2058]&m[2059]&m[2060]&m[2061]&~m[2080]))&BiasedRNG[1121])|(((m[2058]&~m[2059]&~m[2060]&~m[2061]&m[2080])|(~m[2058]&m[2059]&~m[2060]&~m[2061]&m[2080])|(~m[2058]&~m[2059]&m[2060]&~m[2061]&m[2080])|(m[2058]&m[2059]&~m[2060]&m[2061]&m[2080])|(m[2058]&~m[2059]&m[2060]&m[2061]&m[2080])|(~m[2058]&m[2059]&m[2060]&m[2061]&m[2080]))&~BiasedRNG[1121])|((m[2058]&m[2059]&~m[2060]&~m[2061]&~m[2080])|(m[2058]&~m[2059]&m[2060]&~m[2061]&~m[2080])|(~m[2058]&m[2059]&m[2060]&~m[2061]&~m[2080])|(m[2058]&m[2059]&m[2060]&~m[2061]&~m[2080])|(m[2058]&m[2059]&m[2060]&m[2061]&~m[2080])|(m[2058]&m[2059]&~m[2060]&~m[2061]&m[2080])|(m[2058]&~m[2059]&m[2060]&~m[2061]&m[2080])|(~m[2058]&m[2059]&m[2060]&~m[2061]&m[2080])|(m[2058]&m[2059]&m[2060]&~m[2061]&m[2080])|(m[2058]&m[2059]&m[2060]&m[2061]&m[2080]));
    m[2067] = (((m[2063]&~m[2064]&~m[2065]&~m[2066]&~m[2085])|(~m[2063]&m[2064]&~m[2065]&~m[2066]&~m[2085])|(~m[2063]&~m[2064]&m[2065]&~m[2066]&~m[2085])|(m[2063]&m[2064]&~m[2065]&m[2066]&~m[2085])|(m[2063]&~m[2064]&m[2065]&m[2066]&~m[2085])|(~m[2063]&m[2064]&m[2065]&m[2066]&~m[2085]))&BiasedRNG[1122])|(((m[2063]&~m[2064]&~m[2065]&~m[2066]&m[2085])|(~m[2063]&m[2064]&~m[2065]&~m[2066]&m[2085])|(~m[2063]&~m[2064]&m[2065]&~m[2066]&m[2085])|(m[2063]&m[2064]&~m[2065]&m[2066]&m[2085])|(m[2063]&~m[2064]&m[2065]&m[2066]&m[2085])|(~m[2063]&m[2064]&m[2065]&m[2066]&m[2085]))&~BiasedRNG[1122])|((m[2063]&m[2064]&~m[2065]&~m[2066]&~m[2085])|(m[2063]&~m[2064]&m[2065]&~m[2066]&~m[2085])|(~m[2063]&m[2064]&m[2065]&~m[2066]&~m[2085])|(m[2063]&m[2064]&m[2065]&~m[2066]&~m[2085])|(m[2063]&m[2064]&m[2065]&m[2066]&~m[2085])|(m[2063]&m[2064]&~m[2065]&~m[2066]&m[2085])|(m[2063]&~m[2064]&m[2065]&~m[2066]&m[2085])|(~m[2063]&m[2064]&m[2065]&~m[2066]&m[2085])|(m[2063]&m[2064]&m[2065]&~m[2066]&m[2085])|(m[2063]&m[2064]&m[2065]&m[2066]&m[2085]));
    m[2072] = (((m[2068]&~m[2069]&~m[2070]&~m[2071]&~m[2090])|(~m[2068]&m[2069]&~m[2070]&~m[2071]&~m[2090])|(~m[2068]&~m[2069]&m[2070]&~m[2071]&~m[2090])|(m[2068]&m[2069]&~m[2070]&m[2071]&~m[2090])|(m[2068]&~m[2069]&m[2070]&m[2071]&~m[2090])|(~m[2068]&m[2069]&m[2070]&m[2071]&~m[2090]))&BiasedRNG[1123])|(((m[2068]&~m[2069]&~m[2070]&~m[2071]&m[2090])|(~m[2068]&m[2069]&~m[2070]&~m[2071]&m[2090])|(~m[2068]&~m[2069]&m[2070]&~m[2071]&m[2090])|(m[2068]&m[2069]&~m[2070]&m[2071]&m[2090])|(m[2068]&~m[2069]&m[2070]&m[2071]&m[2090])|(~m[2068]&m[2069]&m[2070]&m[2071]&m[2090]))&~BiasedRNG[1123])|((m[2068]&m[2069]&~m[2070]&~m[2071]&~m[2090])|(m[2068]&~m[2069]&m[2070]&~m[2071]&~m[2090])|(~m[2068]&m[2069]&m[2070]&~m[2071]&~m[2090])|(m[2068]&m[2069]&m[2070]&~m[2071]&~m[2090])|(m[2068]&m[2069]&m[2070]&m[2071]&~m[2090])|(m[2068]&m[2069]&~m[2070]&~m[2071]&m[2090])|(m[2068]&~m[2069]&m[2070]&~m[2071]&m[2090])|(~m[2068]&m[2069]&m[2070]&~m[2071]&m[2090])|(m[2068]&m[2069]&m[2070]&~m[2071]&m[2090])|(m[2068]&m[2069]&m[2070]&m[2071]&m[2090]));
    m[2077] = (((m[2073]&~m[2074]&~m[2075]&~m[2076]&~m[2095])|(~m[2073]&m[2074]&~m[2075]&~m[2076]&~m[2095])|(~m[2073]&~m[2074]&m[2075]&~m[2076]&~m[2095])|(m[2073]&m[2074]&~m[2075]&m[2076]&~m[2095])|(m[2073]&~m[2074]&m[2075]&m[2076]&~m[2095])|(~m[2073]&m[2074]&m[2075]&m[2076]&~m[2095]))&BiasedRNG[1124])|(((m[2073]&~m[2074]&~m[2075]&~m[2076]&m[2095])|(~m[2073]&m[2074]&~m[2075]&~m[2076]&m[2095])|(~m[2073]&~m[2074]&m[2075]&~m[2076]&m[2095])|(m[2073]&m[2074]&~m[2075]&m[2076]&m[2095])|(m[2073]&~m[2074]&m[2075]&m[2076]&m[2095])|(~m[2073]&m[2074]&m[2075]&m[2076]&m[2095]))&~BiasedRNG[1124])|((m[2073]&m[2074]&~m[2075]&~m[2076]&~m[2095])|(m[2073]&~m[2074]&m[2075]&~m[2076]&~m[2095])|(~m[2073]&m[2074]&m[2075]&~m[2076]&~m[2095])|(m[2073]&m[2074]&m[2075]&~m[2076]&~m[2095])|(m[2073]&m[2074]&m[2075]&m[2076]&~m[2095])|(m[2073]&m[2074]&~m[2075]&~m[2076]&m[2095])|(m[2073]&~m[2074]&m[2075]&~m[2076]&m[2095])|(~m[2073]&m[2074]&m[2075]&~m[2076]&m[2095])|(m[2073]&m[2074]&m[2075]&~m[2076]&m[2095])|(m[2073]&m[2074]&m[2075]&m[2076]&m[2095]));
    m[2082] = (((m[2078]&~m[2079]&~m[2080]&~m[2081]&~m[2098])|(~m[2078]&m[2079]&~m[2080]&~m[2081]&~m[2098])|(~m[2078]&~m[2079]&m[2080]&~m[2081]&~m[2098])|(m[2078]&m[2079]&~m[2080]&m[2081]&~m[2098])|(m[2078]&~m[2079]&m[2080]&m[2081]&~m[2098])|(~m[2078]&m[2079]&m[2080]&m[2081]&~m[2098]))&BiasedRNG[1125])|(((m[2078]&~m[2079]&~m[2080]&~m[2081]&m[2098])|(~m[2078]&m[2079]&~m[2080]&~m[2081]&m[2098])|(~m[2078]&~m[2079]&m[2080]&~m[2081]&m[2098])|(m[2078]&m[2079]&~m[2080]&m[2081]&m[2098])|(m[2078]&~m[2079]&m[2080]&m[2081]&m[2098])|(~m[2078]&m[2079]&m[2080]&m[2081]&m[2098]))&~BiasedRNG[1125])|((m[2078]&m[2079]&~m[2080]&~m[2081]&~m[2098])|(m[2078]&~m[2079]&m[2080]&~m[2081]&~m[2098])|(~m[2078]&m[2079]&m[2080]&~m[2081]&~m[2098])|(m[2078]&m[2079]&m[2080]&~m[2081]&~m[2098])|(m[2078]&m[2079]&m[2080]&m[2081]&~m[2098])|(m[2078]&m[2079]&~m[2080]&~m[2081]&m[2098])|(m[2078]&~m[2079]&m[2080]&~m[2081]&m[2098])|(~m[2078]&m[2079]&m[2080]&~m[2081]&m[2098])|(m[2078]&m[2079]&m[2080]&~m[2081]&m[2098])|(m[2078]&m[2079]&m[2080]&m[2081]&m[2098]));
    m[2087] = (((m[2083]&~m[2084]&~m[2085]&~m[2086]&~m[2100])|(~m[2083]&m[2084]&~m[2085]&~m[2086]&~m[2100])|(~m[2083]&~m[2084]&m[2085]&~m[2086]&~m[2100])|(m[2083]&m[2084]&~m[2085]&m[2086]&~m[2100])|(m[2083]&~m[2084]&m[2085]&m[2086]&~m[2100])|(~m[2083]&m[2084]&m[2085]&m[2086]&~m[2100]))&BiasedRNG[1126])|(((m[2083]&~m[2084]&~m[2085]&~m[2086]&m[2100])|(~m[2083]&m[2084]&~m[2085]&~m[2086]&m[2100])|(~m[2083]&~m[2084]&m[2085]&~m[2086]&m[2100])|(m[2083]&m[2084]&~m[2085]&m[2086]&m[2100])|(m[2083]&~m[2084]&m[2085]&m[2086]&m[2100])|(~m[2083]&m[2084]&m[2085]&m[2086]&m[2100]))&~BiasedRNG[1126])|((m[2083]&m[2084]&~m[2085]&~m[2086]&~m[2100])|(m[2083]&~m[2084]&m[2085]&~m[2086]&~m[2100])|(~m[2083]&m[2084]&m[2085]&~m[2086]&~m[2100])|(m[2083]&m[2084]&m[2085]&~m[2086]&~m[2100])|(m[2083]&m[2084]&m[2085]&m[2086]&~m[2100])|(m[2083]&m[2084]&~m[2085]&~m[2086]&m[2100])|(m[2083]&~m[2084]&m[2085]&~m[2086]&m[2100])|(~m[2083]&m[2084]&m[2085]&~m[2086]&m[2100])|(m[2083]&m[2084]&m[2085]&~m[2086]&m[2100])|(m[2083]&m[2084]&m[2085]&m[2086]&m[2100]));
    m[2092] = (((m[2088]&~m[2089]&~m[2090]&~m[2091]&~m[2105])|(~m[2088]&m[2089]&~m[2090]&~m[2091]&~m[2105])|(~m[2088]&~m[2089]&m[2090]&~m[2091]&~m[2105])|(m[2088]&m[2089]&~m[2090]&m[2091]&~m[2105])|(m[2088]&~m[2089]&m[2090]&m[2091]&~m[2105])|(~m[2088]&m[2089]&m[2090]&m[2091]&~m[2105]))&BiasedRNG[1127])|(((m[2088]&~m[2089]&~m[2090]&~m[2091]&m[2105])|(~m[2088]&m[2089]&~m[2090]&~m[2091]&m[2105])|(~m[2088]&~m[2089]&m[2090]&~m[2091]&m[2105])|(m[2088]&m[2089]&~m[2090]&m[2091]&m[2105])|(m[2088]&~m[2089]&m[2090]&m[2091]&m[2105])|(~m[2088]&m[2089]&m[2090]&m[2091]&m[2105]))&~BiasedRNG[1127])|((m[2088]&m[2089]&~m[2090]&~m[2091]&~m[2105])|(m[2088]&~m[2089]&m[2090]&~m[2091]&~m[2105])|(~m[2088]&m[2089]&m[2090]&~m[2091]&~m[2105])|(m[2088]&m[2089]&m[2090]&~m[2091]&~m[2105])|(m[2088]&m[2089]&m[2090]&m[2091]&~m[2105])|(m[2088]&m[2089]&~m[2090]&~m[2091]&m[2105])|(m[2088]&~m[2089]&m[2090]&~m[2091]&m[2105])|(~m[2088]&m[2089]&m[2090]&~m[2091]&m[2105])|(m[2088]&m[2089]&m[2090]&~m[2091]&m[2105])|(m[2088]&m[2089]&m[2090]&m[2091]&m[2105]));
    m[2097] = (((m[2093]&~m[2094]&~m[2095]&~m[2096]&~m[2110])|(~m[2093]&m[2094]&~m[2095]&~m[2096]&~m[2110])|(~m[2093]&~m[2094]&m[2095]&~m[2096]&~m[2110])|(m[2093]&m[2094]&~m[2095]&m[2096]&~m[2110])|(m[2093]&~m[2094]&m[2095]&m[2096]&~m[2110])|(~m[2093]&m[2094]&m[2095]&m[2096]&~m[2110]))&BiasedRNG[1128])|(((m[2093]&~m[2094]&~m[2095]&~m[2096]&m[2110])|(~m[2093]&m[2094]&~m[2095]&~m[2096]&m[2110])|(~m[2093]&~m[2094]&m[2095]&~m[2096]&m[2110])|(m[2093]&m[2094]&~m[2095]&m[2096]&m[2110])|(m[2093]&~m[2094]&m[2095]&m[2096]&m[2110])|(~m[2093]&m[2094]&m[2095]&m[2096]&m[2110]))&~BiasedRNG[1128])|((m[2093]&m[2094]&~m[2095]&~m[2096]&~m[2110])|(m[2093]&~m[2094]&m[2095]&~m[2096]&~m[2110])|(~m[2093]&m[2094]&m[2095]&~m[2096]&~m[2110])|(m[2093]&m[2094]&m[2095]&~m[2096]&~m[2110])|(m[2093]&m[2094]&m[2095]&m[2096]&~m[2110])|(m[2093]&m[2094]&~m[2095]&~m[2096]&m[2110])|(m[2093]&~m[2094]&m[2095]&~m[2096]&m[2110])|(~m[2093]&m[2094]&m[2095]&~m[2096]&m[2110])|(m[2093]&m[2094]&m[2095]&~m[2096]&m[2110])|(m[2093]&m[2094]&m[2095]&m[2096]&m[2110]));
    m[2102] = (((m[2098]&~m[2099]&~m[2100]&~m[2101]&~m[2113])|(~m[2098]&m[2099]&~m[2100]&~m[2101]&~m[2113])|(~m[2098]&~m[2099]&m[2100]&~m[2101]&~m[2113])|(m[2098]&m[2099]&~m[2100]&m[2101]&~m[2113])|(m[2098]&~m[2099]&m[2100]&m[2101]&~m[2113])|(~m[2098]&m[2099]&m[2100]&m[2101]&~m[2113]))&BiasedRNG[1129])|(((m[2098]&~m[2099]&~m[2100]&~m[2101]&m[2113])|(~m[2098]&m[2099]&~m[2100]&~m[2101]&m[2113])|(~m[2098]&~m[2099]&m[2100]&~m[2101]&m[2113])|(m[2098]&m[2099]&~m[2100]&m[2101]&m[2113])|(m[2098]&~m[2099]&m[2100]&m[2101]&m[2113])|(~m[2098]&m[2099]&m[2100]&m[2101]&m[2113]))&~BiasedRNG[1129])|((m[2098]&m[2099]&~m[2100]&~m[2101]&~m[2113])|(m[2098]&~m[2099]&m[2100]&~m[2101]&~m[2113])|(~m[2098]&m[2099]&m[2100]&~m[2101]&~m[2113])|(m[2098]&m[2099]&m[2100]&~m[2101]&~m[2113])|(m[2098]&m[2099]&m[2100]&m[2101]&~m[2113])|(m[2098]&m[2099]&~m[2100]&~m[2101]&m[2113])|(m[2098]&~m[2099]&m[2100]&~m[2101]&m[2113])|(~m[2098]&m[2099]&m[2100]&~m[2101]&m[2113])|(m[2098]&m[2099]&m[2100]&~m[2101]&m[2113])|(m[2098]&m[2099]&m[2100]&m[2101]&m[2113]));
    m[2107] = (((m[2103]&~m[2104]&~m[2105]&~m[2106]&~m[2115])|(~m[2103]&m[2104]&~m[2105]&~m[2106]&~m[2115])|(~m[2103]&~m[2104]&m[2105]&~m[2106]&~m[2115])|(m[2103]&m[2104]&~m[2105]&m[2106]&~m[2115])|(m[2103]&~m[2104]&m[2105]&m[2106]&~m[2115])|(~m[2103]&m[2104]&m[2105]&m[2106]&~m[2115]))&BiasedRNG[1130])|(((m[2103]&~m[2104]&~m[2105]&~m[2106]&m[2115])|(~m[2103]&m[2104]&~m[2105]&~m[2106]&m[2115])|(~m[2103]&~m[2104]&m[2105]&~m[2106]&m[2115])|(m[2103]&m[2104]&~m[2105]&m[2106]&m[2115])|(m[2103]&~m[2104]&m[2105]&m[2106]&m[2115])|(~m[2103]&m[2104]&m[2105]&m[2106]&m[2115]))&~BiasedRNG[1130])|((m[2103]&m[2104]&~m[2105]&~m[2106]&~m[2115])|(m[2103]&~m[2104]&m[2105]&~m[2106]&~m[2115])|(~m[2103]&m[2104]&m[2105]&~m[2106]&~m[2115])|(m[2103]&m[2104]&m[2105]&~m[2106]&~m[2115])|(m[2103]&m[2104]&m[2105]&m[2106]&~m[2115])|(m[2103]&m[2104]&~m[2105]&~m[2106]&m[2115])|(m[2103]&~m[2104]&m[2105]&~m[2106]&m[2115])|(~m[2103]&m[2104]&m[2105]&~m[2106]&m[2115])|(m[2103]&m[2104]&m[2105]&~m[2106]&m[2115])|(m[2103]&m[2104]&m[2105]&m[2106]&m[2115]));
    m[2112] = (((m[2108]&~m[2109]&~m[2110]&~m[2111]&~m[2120])|(~m[2108]&m[2109]&~m[2110]&~m[2111]&~m[2120])|(~m[2108]&~m[2109]&m[2110]&~m[2111]&~m[2120])|(m[2108]&m[2109]&~m[2110]&m[2111]&~m[2120])|(m[2108]&~m[2109]&m[2110]&m[2111]&~m[2120])|(~m[2108]&m[2109]&m[2110]&m[2111]&~m[2120]))&BiasedRNG[1131])|(((m[2108]&~m[2109]&~m[2110]&~m[2111]&m[2120])|(~m[2108]&m[2109]&~m[2110]&~m[2111]&m[2120])|(~m[2108]&~m[2109]&m[2110]&~m[2111]&m[2120])|(m[2108]&m[2109]&~m[2110]&m[2111]&m[2120])|(m[2108]&~m[2109]&m[2110]&m[2111]&m[2120])|(~m[2108]&m[2109]&m[2110]&m[2111]&m[2120]))&~BiasedRNG[1131])|((m[2108]&m[2109]&~m[2110]&~m[2111]&~m[2120])|(m[2108]&~m[2109]&m[2110]&~m[2111]&~m[2120])|(~m[2108]&m[2109]&m[2110]&~m[2111]&~m[2120])|(m[2108]&m[2109]&m[2110]&~m[2111]&~m[2120])|(m[2108]&m[2109]&m[2110]&m[2111]&~m[2120])|(m[2108]&m[2109]&~m[2110]&~m[2111]&m[2120])|(m[2108]&~m[2109]&m[2110]&~m[2111]&m[2120])|(~m[2108]&m[2109]&m[2110]&~m[2111]&m[2120])|(m[2108]&m[2109]&m[2110]&~m[2111]&m[2120])|(m[2108]&m[2109]&m[2110]&m[2111]&m[2120]));
    m[2117] = (((m[2113]&~m[2114]&~m[2115]&~m[2116]&~m[2123])|(~m[2113]&m[2114]&~m[2115]&~m[2116]&~m[2123])|(~m[2113]&~m[2114]&m[2115]&~m[2116]&~m[2123])|(m[2113]&m[2114]&~m[2115]&m[2116]&~m[2123])|(m[2113]&~m[2114]&m[2115]&m[2116]&~m[2123])|(~m[2113]&m[2114]&m[2115]&m[2116]&~m[2123]))&BiasedRNG[1132])|(((m[2113]&~m[2114]&~m[2115]&~m[2116]&m[2123])|(~m[2113]&m[2114]&~m[2115]&~m[2116]&m[2123])|(~m[2113]&~m[2114]&m[2115]&~m[2116]&m[2123])|(m[2113]&m[2114]&~m[2115]&m[2116]&m[2123])|(m[2113]&~m[2114]&m[2115]&m[2116]&m[2123])|(~m[2113]&m[2114]&m[2115]&m[2116]&m[2123]))&~BiasedRNG[1132])|((m[2113]&m[2114]&~m[2115]&~m[2116]&~m[2123])|(m[2113]&~m[2114]&m[2115]&~m[2116]&~m[2123])|(~m[2113]&m[2114]&m[2115]&~m[2116]&~m[2123])|(m[2113]&m[2114]&m[2115]&~m[2116]&~m[2123])|(m[2113]&m[2114]&m[2115]&m[2116]&~m[2123])|(m[2113]&m[2114]&~m[2115]&~m[2116]&m[2123])|(m[2113]&~m[2114]&m[2115]&~m[2116]&m[2123])|(~m[2113]&m[2114]&m[2115]&~m[2116]&m[2123])|(m[2113]&m[2114]&m[2115]&~m[2116]&m[2123])|(m[2113]&m[2114]&m[2115]&m[2116]&m[2123]));
    m[2122] = (((m[2118]&~m[2119]&~m[2120]&~m[2121]&~m[2125])|(~m[2118]&m[2119]&~m[2120]&~m[2121]&~m[2125])|(~m[2118]&~m[2119]&m[2120]&~m[2121]&~m[2125])|(m[2118]&m[2119]&~m[2120]&m[2121]&~m[2125])|(m[2118]&~m[2119]&m[2120]&m[2121]&~m[2125])|(~m[2118]&m[2119]&m[2120]&m[2121]&~m[2125]))&BiasedRNG[1133])|(((m[2118]&~m[2119]&~m[2120]&~m[2121]&m[2125])|(~m[2118]&m[2119]&~m[2120]&~m[2121]&m[2125])|(~m[2118]&~m[2119]&m[2120]&~m[2121]&m[2125])|(m[2118]&m[2119]&~m[2120]&m[2121]&m[2125])|(m[2118]&~m[2119]&m[2120]&m[2121]&m[2125])|(~m[2118]&m[2119]&m[2120]&m[2121]&m[2125]))&~BiasedRNG[1133])|((m[2118]&m[2119]&~m[2120]&~m[2121]&~m[2125])|(m[2118]&~m[2119]&m[2120]&~m[2121]&~m[2125])|(~m[2118]&m[2119]&m[2120]&~m[2121]&~m[2125])|(m[2118]&m[2119]&m[2120]&~m[2121]&~m[2125])|(m[2118]&m[2119]&m[2120]&m[2121]&~m[2125])|(m[2118]&m[2119]&~m[2120]&~m[2121]&m[2125])|(m[2118]&~m[2119]&m[2120]&~m[2121]&m[2125])|(~m[2118]&m[2119]&m[2120]&~m[2121]&m[2125])|(m[2118]&m[2119]&m[2120]&~m[2121]&m[2125])|(m[2118]&m[2119]&m[2120]&m[2121]&m[2125]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[975]&LFSRcolor0[1243]&LFSRcolor0[496]&LFSRcolor0[409]);
    BiasedRNG[1] = (LFSRcolor0[1093]&LFSRcolor0[68]&LFSRcolor0[568]&LFSRcolor0[334]);
    BiasedRNG[2] = (LFSRcolor0[47]&LFSRcolor0[146]&LFSRcolor0[11]&LFSRcolor0[885]);
    BiasedRNG[3] = (LFSRcolor0[700]&LFSRcolor0[260]&LFSRcolor0[359]&LFSRcolor0[346]);
    BiasedRNG[4] = (LFSRcolor0[1059]&LFSRcolor0[755]&LFSRcolor0[464]&LFSRcolor0[775]);
    BiasedRNG[5] = (LFSRcolor0[522]&LFSRcolor0[353]&LFSRcolor0[321]&LFSRcolor0[1207]);
    BiasedRNG[6] = (LFSRcolor0[113]&LFSRcolor0[80]&LFSRcolor0[1128]&LFSRcolor0[1293]);
    BiasedRNG[7] = (LFSRcolor0[258]&LFSRcolor0[363]&LFSRcolor0[1053]&LFSRcolor0[724]);
    BiasedRNG[8] = (LFSRcolor0[355]&LFSRcolor0[750]&LFSRcolor0[770]&LFSRcolor0[671]);
    BiasedRNG[9] = (LFSRcolor0[666]&LFSRcolor0[962]&LFSRcolor0[783]&LFSRcolor0[1068]);
    BiasedRNG[10] = (LFSRcolor0[874]&LFSRcolor0[497]&LFSRcolor0[1130]&LFSRcolor0[858]);
    BiasedRNG[11] = (LFSRcolor0[1186]&LFSRcolor0[92]&LFSRcolor0[212]&LFSRcolor0[259]);
    BiasedRNG[12] = (LFSRcolor0[112]&LFSRcolor0[276]&LFSRcolor0[907]&LFSRcolor0[797]);
    BiasedRNG[13] = (LFSRcolor0[661]&LFSRcolor0[0]&LFSRcolor0[746]&LFSRcolor0[658]);
    BiasedRNG[14] = (LFSRcolor0[896]&LFSRcolor0[1064]&LFSRcolor0[761]&LFSRcolor0[1137]);
    BiasedRNG[15] = (LFSRcolor0[237]&LFSRcolor0[160]&LFSRcolor0[829]&LFSRcolor0[233]);
    BiasedRNG[16] = (LFSRcolor0[304]&LFSRcolor0[517]&LFSRcolor0[422]&LFSRcolor0[1256]);
    BiasedRNG[17] = (LFSRcolor0[45]&LFSRcolor0[850]&LFSRcolor0[544]&LFSRcolor0[728]);
    BiasedRNG[18] = (LFSRcolor0[966]&LFSRcolor0[734]&LFSRcolor0[570]&LFSRcolor0[295]);
    BiasedRNG[19] = (LFSRcolor0[478]&LFSRcolor0[191]&LFSRcolor0[876]&LFSRcolor0[1094]);
    BiasedRNG[20] = (LFSRcolor0[504]&LFSRcolor0[401]&LFSRcolor0[34]&LFSRcolor0[602]);
    BiasedRNG[21] = (LFSRcolor0[832]&LFSRcolor0[837]&LFSRcolor0[1028]&LFSRcolor0[733]);
    BiasedRNG[22] = (LFSRcolor0[1300]&LFSRcolor0[703]&LFSRcolor0[208]&LFSRcolor0[1277]);
    BiasedRNG[23] = (LFSRcolor0[803]&LFSRcolor0[609]&LFSRcolor0[1272]&LFSRcolor0[83]);
    BiasedRNG[24] = (LFSRcolor0[668]&LFSRcolor0[1124]&LFSRcolor0[1139]&LFSRcolor0[1126]);
    BiasedRNG[25] = (LFSRcolor0[615]&LFSRcolor0[109]&LFSRcolor0[434]&LFSRcolor0[732]);
    BiasedRNG[26] = (LFSRcolor0[238]&LFSRcolor0[808]&LFSRcolor0[373]&LFSRcolor0[78]);
    BiasedRNG[27] = (LFSRcolor0[784]&LFSRcolor0[788]&LFSRcolor0[690]&LFSRcolor0[210]);
    BiasedRNG[28] = (LFSRcolor0[1180]&LFSRcolor0[33]&LFSRcolor0[252]&LFSRcolor0[991]);
    BiasedRNG[29] = (LFSRcolor0[2]&LFSRcolor0[860]&LFSRcolor0[394]&LFSRcolor0[667]);
    BiasedRNG[30] = (LFSRcolor0[339]&LFSRcolor0[1141]&LFSRcolor0[1212]&LFSRcolor0[1257]);
    BiasedRNG[31] = (LFSRcolor0[121]&LFSRcolor0[799]&LFSRcolor0[1072]&LFSRcolor0[1190]);
    BiasedRNG[32] = (LFSRcolor0[681]&LFSRcolor0[763]&LFSRcolor0[777]&LFSRcolor0[593]);
    BiasedRNG[33] = (LFSRcolor0[696]&LFSRcolor0[220]&LFSRcolor0[941]&LFSRcolor0[391]);
    BiasedRNG[34] = (LFSRcolor0[999]&LFSRcolor0[1001]&LFSRcolor0[389]&LFSRcolor0[582]);
    BiasedRNG[35] = (LFSRcolor0[145]&LFSRcolor0[133]&LFSRcolor0[764]&LFSRcolor0[126]);
    BiasedRNG[36] = (LFSRcolor0[688]&LFSRcolor0[1177]&LFSRcolor0[1062]&LFSRcolor0[66]);
    BiasedRNG[37] = (LFSRcolor0[1118]&LFSRcolor0[580]&LFSRcolor0[30]&LFSRcolor0[123]);
    BiasedRNG[38] = (LFSRcolor0[108]&LFSRcolor0[936]&LFSRcolor0[909]&LFSRcolor0[919]);
    BiasedRNG[39] = (LFSRcolor0[1058]&LFSRcolor0[228]&LFSRcolor0[125]&LFSRcolor0[82]);
    BiasedRNG[40] = (LFSRcolor0[959]&LFSRcolor0[342]&LFSRcolor0[807]&LFSRcolor0[1239]);
    BiasedRNG[41] = (LFSRcolor0[1101]&LFSRcolor0[617]&LFSRcolor0[794]&LFSRcolor0[531]);
    BiasedRNG[42] = (LFSRcolor0[217]&LFSRcolor0[597]&LFSRcolor0[51]&LFSRcolor0[1333]);
    BiasedRNG[43] = (LFSRcolor0[815]&LFSRcolor0[542]&LFSRcolor0[347]&LFSRcolor0[1060]);
    BiasedRNG[44] = (LFSRcolor0[157]&LFSRcolor0[447]&LFSRcolor0[49]&LFSRcolor0[287]);
    BiasedRNG[45] = (LFSRcolor0[891]&LFSRcolor0[935]&LFSRcolor0[1013]&LFSRcolor0[350]);
    BiasedRNG[46] = (LFSRcolor0[1092]&LFSRcolor0[1329]&LFSRcolor0[1229]&LFSRcolor0[1275]);
    BiasedRNG[47] = (LFSRcolor0[611]&LFSRcolor0[336]&LFSRcolor0[281]&LFSRcolor0[972]);
    BiasedRNG[48] = (LFSRcolor0[69]&LFSRcolor0[620]&LFSRcolor0[767]&LFSRcolor0[599]);
    BiasedRNG[49] = (LFSRcolor0[296]&LFSRcolor0[664]&LFSRcolor0[1230]&LFSRcolor0[171]);
    BiasedRNG[50] = (LFSRcolor0[902]&LFSRcolor0[326]&LFSRcolor0[247]&LFSRcolor0[152]);
    BiasedRNG[51] = (LFSRcolor0[453]&LFSRcolor0[984]&LFSRcolor0[562]&LFSRcolor0[1081]);
    BiasedRNG[52] = (LFSRcolor0[1220]&LFSRcolor0[1318]&LFSRcolor0[132]&LFSRcolor0[234]);
    BiasedRNG[53] = (LFSRcolor0[44]&LFSRcolor0[1269]&LFSRcolor0[134]&LFSRcolor0[718]);
    BiasedRNG[54] = (LFSRcolor0[94]&LFSRcolor0[1222]&LFSRcolor0[705]&LFSRcolor0[560]);
    BiasedRNG[55] = (LFSRcolor0[1145]&LFSRcolor0[563]&LFSRcolor0[1122]&LFSRcolor0[840]);
    BiasedRNG[56] = (LFSRcolor0[880]&LFSRcolor0[1245]&LFSRcolor0[1163]&LFSRcolor0[120]);
    BiasedRNG[57] = (LFSRcolor0[50]&LFSRcolor0[1106]&LFSRcolor0[614]&LFSRcolor0[298]);
    BiasedRNG[58] = (LFSRcolor0[766]&LFSRcolor0[381]&LFSRcolor0[987]&LFSRcolor0[692]);
    BiasedRNG[59] = (LFSRcolor0[1078]&LFSRcolor0[140]&LFSRcolor0[56]&LFSRcolor0[1255]);
    BiasedRNG[60] = (LFSRcolor0[1317]&LFSRcolor0[40]&LFSRcolor0[595]&LFSRcolor0[214]);
    BiasedRNG[61] = (LFSRcolor0[1276]&LFSRcolor0[370]&LFSRcolor0[236]&LFSRcolor0[1291]);
    BiasedRNG[62] = (LFSRcolor0[1085]&LFSRcolor0[149]&LFSRcolor0[424]&LFSRcolor0[185]);
    BiasedRNG[63] = (LFSRcolor0[933]&LFSRcolor0[616]&LFSRcolor0[1202]&LFSRcolor0[1018]);
    BiasedRNG[64] = (LFSRcolor0[632]&LFSRcolor0[806]&LFSRcolor0[871]&LFSRcolor0[795]);
    BiasedRNG[65] = (LFSRcolor0[556]&LFSRcolor0[195]&LFSRcolor0[813]&LFSRcolor0[1054]);
    BiasedRNG[66] = (LFSRcolor0[1017]&LFSRcolor0[1065]&LFSRcolor0[1203]&LFSRcolor0[899]);
    BiasedRNG[67] = (LFSRcolor0[659]&LFSRcolor0[357]&LFSRcolor0[589]&LFSRcolor0[629]);
    BiasedRNG[68] = (LFSRcolor0[787]&LFSRcolor0[1007]&LFSRcolor0[340]&LFSRcolor0[20]);
    BiasedRNG[69] = (LFSRcolor0[303]&LFSRcolor0[317]&LFSRcolor0[141]&LFSRcolor0[253]);
    BiasedRNG[70] = (LFSRcolor0[1042]&LFSRcolor0[172]&LFSRcolor0[178]&LFSRcolor0[992]);
    BiasedRNG[71] = (LFSRcolor0[205]&LFSRcolor0[1200]&LFSRcolor0[385]&LFSRcolor0[757]);
    BiasedRNG[72] = (LFSRcolor0[493]&LFSRcolor0[79]&LFSRcolor0[331]&LFSRcolor0[436]);
    BiasedRNG[73] = (LFSRcolor0[390]&LFSRcolor0[367]&LFSRcolor0[491]&LFSRcolor0[285]);
    BiasedRNG[74] = (LFSRcolor0[1161]&LFSRcolor0[868]&LFSRcolor0[515]&LFSRcolor0[546]);
    BiasedRNG[75] = (LFSRcolor0[519]&LFSRcolor0[279]&LFSRcolor0[442]&LFSRcolor0[882]);
    BiasedRNG[76] = (LFSRcolor0[360]&LFSRcolor0[159]&LFSRcolor0[914]&LFSRcolor0[313]);
    BiasedRNG[77] = (LFSRcolor0[1216]&LFSRcolor0[366]&LFSRcolor0[811]&LFSRcolor0[356]);
    BiasedRNG[78] = (LFSRcolor0[1132]&LFSRcolor0[384]&LFSRcolor0[571]&LFSRcolor0[19]);
    BiasedRNG[79] = (LFSRcolor0[84]&LFSRcolor0[219]&LFSRcolor0[1008]&LFSRcolor0[168]);
    BiasedRNG[80] = (LFSRcolor0[1250]&LFSRcolor0[1172]&LFSRcolor0[1321]&LFSRcolor0[549]);
    BiasedRNG[81] = (LFSRcolor0[679]&LFSRcolor0[1160]&LFSRcolor0[328]&LFSRcolor0[721]);
    BiasedRNG[82] = (LFSRcolor0[1103]&LFSRcolor0[392]&LFSRcolor0[1020]&LFSRcolor0[894]);
    BiasedRNG[83] = (LFSRcolor0[680]&LFSRcolor0[583]&LFSRcolor0[793]&LFSRcolor0[470]);
    BiasedRNG[84] = (LFSRcolor0[165]&LFSRcolor0[1148]&LFSRcolor0[1181]&LFSRcolor0[268]);
    BiasedRNG[85] = (LFSRcolor0[1284]&LFSRcolor0[812]&LFSRcolor0[1251]&LFSRcolor0[849]);
    BiasedRNG[86] = (LFSRcolor0[820]&LFSRcolor0[708]&LFSRcolor0[456]&LFSRcolor0[591]);
    BiasedRNG[87] = (LFSRcolor0[1098]&LFSRcolor0[1120]&LFSRcolor0[1090]&LFSRcolor0[254]);
    BiasedRNG[88] = (LFSRcolor0[1082]&LFSRcolor0[978]&LFSRcolor0[62]&LFSRcolor0[600]);
    BiasedRNG[89] = (LFSRcolor0[528]&LFSRcolor0[1301]&LFSRcolor0[1119]&LFSRcolor0[809]);
    BiasedRNG[90] = (LFSRcolor0[652]&LFSRcolor0[476]&LFSRcolor0[1114]&LFSRcolor0[378]);
    BiasedRNG[91] = (LFSRcolor0[156]&LFSRcolor0[506]&LFSRcolor0[908]&LFSRcolor0[854]);
    BiasedRNG[92] = (LFSRcolor0[691]&LFSRcolor0[1012]&LFSRcolor0[230]&LFSRcolor0[1158]);
    BiasedRNG[93] = (LFSRcolor0[1194]&LFSRcolor0[1112]&LFSRcolor0[877]&LFSRcolor0[663]);
    BiasedRNG[94] = (LFSRcolor0[744]&LFSRcolor0[869]&LFSRcolor0[1070]&LFSRcolor0[547]);
    BiasedRNG[95] = (LFSRcolor0[830]&LFSRcolor0[558]&LFSRcolor0[895]&LFSRcolor0[118]);
    BiasedRNG[96] = (LFSRcolor0[557]&LFSRcolor0[417]&LFSRcolor0[1156]&LFSRcolor0[459]);
    BiasedRNG[97] = (LFSRcolor0[1288]&LFSRcolor0[527]&LFSRcolor0[1253]&LFSRcolor0[512]);
    BiasedRNG[98] = (LFSRcolor0[364]&LFSRcolor0[211]&LFSRcolor0[315]&LFSRcolor0[225]);
    BiasedRNG[99] = (LFSRcolor0[818]&LFSRcolor0[129]&LFSRcolor0[1049]&LFSRcolor0[400]);
    BiasedRNG[100] = (LFSRcolor0[596]&LFSRcolor0[1170]&LFSRcolor0[628]&LFSRcolor0[17]);
    BiasedRNG[101] = (LFSRcolor0[535]&LFSRcolor0[1208]&LFSRcolor0[741]&LFSRcolor0[10]);
    BiasedRNG[102] = (LFSRcolor0[525]&LFSRcolor0[748]&LFSRcolor0[606]&LFSRcolor0[248]);
    BiasedRNG[103] = (LFSRcolor0[727]&LFSRcolor0[202]&LFSRcolor0[1209]&LFSRcolor0[102]);
    BiasedRNG[104] = (LFSRcolor0[856]&LFSRcolor0[939]&LFSRcolor0[46]&LFSRcolor0[1285]);
    BiasedRNG[105] = (LFSRcolor0[408]&LFSRcolor0[1066]&LFSRcolor0[779]&LFSRcolor0[1009]);
    BiasedRNG[106] = (LFSRcolor0[301]&LFSRcolor0[627]&LFSRcolor0[87]&LFSRcolor0[1313]);
    BiasedRNG[107] = (LFSRcolor0[587]&LFSRcolor0[857]&LFSRcolor0[901]&LFSRcolor0[601]);
    BiasedRNG[108] = (LFSRcolor0[119]&LFSRcolor0[404]&LFSRcolor0[98]&LFSRcolor0[906]);
    BiasedRNG[109] = (LFSRcolor0[451]&LFSRcolor0[1004]&LFSRcolor0[6]&LFSRcolor0[865]);
    BiasedRNG[110] = (LFSRcolor0[760]&LFSRcolor0[1029]&LFSRcolor0[1149]&LFSRcolor0[863]);
    BiasedRNG[111] = (LFSRcolor0[508]&LFSRcolor0[416]&LFSRcolor0[1270]&LFSRcolor0[709]);
    BiasedRNG[112] = (LFSRcolor0[977]&LFSRcolor0[270]&LFSRcolor0[501]&LFSRcolor0[673]);
    BiasedRNG[113] = (LFSRcolor0[1109]&LFSRcolor0[1296]&LFSRcolor0[433]&LFSRcolor0[244]);
    BiasedRNG[114] = (LFSRcolor0[1314]&LFSRcolor0[930]&LFSRcolor0[1290]&LFSRcolor0[32]);
    BiasedRNG[115] = (LFSRcolor0[26]&LFSRcolor0[484]&LFSRcolor0[280]&LFSRcolor0[153]);
    BiasedRNG[116] = (LFSRcolor0[100]&LFSRcolor0[621]&LFSRcolor0[675]&LFSRcolor0[550]);
    BiasedRNG[117] = (LFSRcolor0[1030]&LFSRcolor0[1011]&LFSRcolor0[655]&LFSRcolor0[1217]);
    BiasedRNG[118] = (LFSRcolor0[27]&LFSRcolor0[1278]&LFSRcolor0[561]&LFSRcolor0[25]);
    BiasedRNG[119] = (LFSRcolor0[862]&LFSRcolor0[931]&LFSRcolor0[1038]&LFSRcolor0[695]);
    BiasedRNG[120] = (LFSRcolor0[740]&LFSRcolor0[1297]&LFSRcolor0[272]&LFSRcolor0[574]);
    BiasedRNG[121] = (LFSRcolor0[643]&LFSRcolor0[911]&LFSRcolor0[239]&LFSRcolor0[81]);
    BiasedRNG[122] = (LFSRcolor0[576]&LFSRcolor0[492]&LFSRcolor0[866]&LFSRcolor0[1302]);
    BiasedRNG[123] = (LFSRcolor0[1240]&LFSRcolor0[1056]&LFSRcolor0[624]&LFSRcolor0[241]);
    BiasedRNG[124] = (LFSRcolor0[175]&LFSRcolor0[870]&LFSRcolor0[289]&LFSRcolor0[853]);
    BiasedRNG[125] = (LFSRcolor0[1043]&LFSRcolor0[878]&LFSRcolor0[1281]&LFSRcolor0[101]);
    BiasedRNG[126] = (LFSRcolor0[67]&LFSRcolor0[1136]&LFSRcolor0[686]&LFSRcolor0[828]);
    BiasedRNG[127] = (LFSRcolor0[1260]&LFSRcolor0[534]&LFSRcolor0[640]&LFSRcolor0[349]);
    BiasedRNG[128] = (LFSRcolor0[509]&LFSRcolor0[946]&LFSRcolor0[91]&LFSRcolor0[224]);
    BiasedRNG[129] = (LFSRcolor0[312]&LFSRcolor0[1330]&LFSRcolor0[440]&LFSRcolor0[754]);
    BiasedRNG[130] = (LFSRcolor0[1002]&LFSRcolor0[446]&LFSRcolor0[405]&LFSRcolor0[330]);
    BiasedRNG[131] = (LFSRcolor0[1283]&LFSRcolor0[927]&LFSRcolor0[1005]&LFSRcolor0[213]);
    BiasedRNG[132] = (LFSRcolor0[1102]&LFSRcolor0[677]&LFSRcolor0[720]&LFSRcolor0[368]);
    BiasedRNG[133] = (LFSRcolor0[541]&LFSRcolor0[533]&LFSRcolor0[308]&LFSRcolor0[299]);
    BiasedRNG[134] = (LFSRcolor0[827]&LFSRcolor0[204]&LFSRcolor0[462]&LFSRcolor0[318]);
    BiasedRNG[135] = (LFSRcolor0[64]&LFSRcolor0[277]&LFSRcolor0[106]&LFSRcolor0[465]);
    BiasedRNG[136] = (LFSRcolor0[1211]&LFSRcolor0[35]&LFSRcolor0[415]&LFSRcolor0[848]);
    BiasedRNG[137] = (LFSRcolor0[431]&LFSRcolor0[993]&LFSRcolor0[1201]&LFSRcolor0[1228]);
    BiasedRNG[138] = (LFSRcolor0[618]&LFSRcolor0[193]&LFSRcolor0[324]&LFSRcolor0[316]);
    BiasedRNG[139] = (LFSRcolor0[89]&LFSRcolor0[28]&LFSRcolor0[58]&LFSRcolor0[524]);
    BiasedRNG[140] = (LFSRcolor0[425]&LFSRcolor0[472]&LFSRcolor0[539]&LFSRcolor0[1238]);
    BiasedRNG[141] = (LFSRcolor0[957]&LFSRcolor0[791]&LFSRcolor0[973]&LFSRcolor0[575]);
    BiasedRNG[142] = (LFSRcolor0[735]&LFSRcolor0[707]&LFSRcolor0[545]&LFSRcolor0[262]);
    BiasedRNG[143] = (LFSRcolor0[521]&LFSRcolor0[598]&LFSRcolor0[76]&LFSRcolor0[179]);
    BiasedRNG[144] = (LFSRcolor0[960]&LFSRcolor0[771]&LFSRcolor0[685]&LFSRcolor0[1069]);
    BiasedRNG[145] = (LFSRcolor0[1178]&LFSRcolor0[590]&LFSRcolor0[1032]&LFSRcolor0[608]);
    BiasedRNG[146] = (LFSRcolor0[971]&LFSRcolor0[768]&LFSRcolor0[834]&LFSRcolor0[762]);
    BiasedRNG[147] = (LFSRcolor0[31]&LFSRcolor0[790]&LFSRcolor0[698]&LFSRcolor0[485]);
    BiasedRNG[148] = (LFSRcolor0[699]&LFSRcolor0[294]&LFSRcolor0[243]&LFSRcolor0[581]);
    BiasedRNG[149] = (LFSRcolor0[482]&LFSRcolor0[42]&LFSRcolor0[1045]&LFSRcolor0[1117]);
    BiasedRNG[150] = (LFSRcolor0[271]&LFSRcolor0[293]&LFSRcolor0[1096]&LFSRcolor0[921]);
    BiasedRNG[151] = (LFSRcolor0[753]&LFSRcolor0[1021]&LFSRcolor0[898]&LFSRcolor0[619]);
    BiasedRNG[152] = (LFSRcolor0[148]&LFSRcolor0[578]&LFSRcolor0[189]&LFSRcolor0[73]);
    BiasedRNG[153] = (LFSRcolor0[256]&LFSRcolor0[523]&LFSRcolor0[170]&LFSRcolor0[1057]);
    BiasedRNG[154] = (LFSRcolor0[432]&LFSRcolor0[955]&LFSRcolor0[418]&LFSRcolor0[477]);
    BiasedRNG[155] = (LFSRcolor0[1127]&LFSRcolor0[839]&LFSRcolor0[713]&LFSRcolor0[88]);
    BiasedRNG[156] = (LFSRcolor0[502]&LFSRcolor0[825]&LFSRcolor0[518]&LFSRcolor0[116]);
    BiasedRNG[157] = (LFSRcolor0[197]&LFSRcolor0[1031]&LFSRcolor0[1048]&LFSRcolor0[65]);
    BiasedRNG[158] = (LFSRcolor0[372]&LFSRcolor0[607]&LFSRcolor0[1155]&LFSRcolor0[448]);
    BiasedRNG[159] = (LFSRcolor0[333]&LFSRcolor0[36]&LFSRcolor0[507]&LFSRcolor0[22]);
    BiasedRNG[160] = (LFSRcolor0[752]&LFSRcolor0[1306]&LFSRcolor0[466]&LFSRcolor0[449]);
    BiasedRNG[161] = (LFSRcolor0[943]&LFSRcolor0[1295]&LFSRcolor0[500]&LFSRcolor0[57]);
    BiasedRNG[162] = (LFSRcolor0[613]&LFSRcolor0[1328]&LFSRcolor0[1184]&LFSRcolor0[351]);
    BiasedRNG[163] = (LFSRcolor0[631]&LFSRcolor0[879]&LFSRcolor0[892]&LFSRcolor0[352]);
    BiasedRNG[164] = (LFSRcolor0[128]&LFSRcolor0[1135]&LFSRcolor0[1263]&LFSRcolor0[814]);
    BiasedRNG[165] = (LFSRcolor0[445]&LFSRcolor0[1324]&LFSRcolor0[437]&LFSRcolor0[520]);
    BiasedRNG[166] = (LFSRcolor0[1322]&LFSRcolor0[647]&LFSRcolor0[639]&LFSRcolor0[41]);
    BiasedRNG[167] = (LFSRcolor0[60]&LFSRcolor0[24]&LFSRcolor0[945]&LFSRcolor0[846]);
    BiasedRNG[168] = (LFSRcolor0[325]&LFSRcolor0[656]&LFSRcolor0[444]&LFSRcolor0[1192]);
    BiasedRNG[169] = (LFSRcolor0[1041]&LFSRcolor0[824]&LFSRcolor0[864]&LFSRcolor0[963]);
    BiasedRNG[170] = (LFSRcolor0[124]&LFSRcolor0[747]&LFSRcolor0[105]&LFSRcolor0[940]);
    BiasedRNG[171] = (LFSRcolor0[1143]&LFSRcolor0[821]&LFSRcolor0[9]&LFSRcolor0[851]);
    BiasedRNG[172] = (LFSRcolor0[458]&LFSRcolor0[805]&LFSRcolor0[884]&LFSRcolor0[242]);
    BiasedRNG[173] = (LFSRcolor0[1168]&LFSRcolor0[548]&LFSRcolor0[1129]&LFSRcolor0[934]);
    BiasedRNG[174] = (LFSRcolor0[756]&LFSRcolor0[1280]&LFSRcolor0[457]&LFSRcolor0[274]);
    BiasedRNG[175] = (LFSRcolor0[1016]&LFSRcolor0[1022]&LFSRcolor0[786]&LFSRcolor0[798]);
    BiasedRNG[176] = (LFSRcolor0[883]&LFSRcolor0[142]&LFSRcolor0[209]&LFSRcolor0[637]);
    BiasedRNG[177] = (LFSRcolor0[54]&LFSRcolor0[111]&LFSRcolor0[1188]&LFSRcolor0[956]);
    BiasedRNG[178] = (LFSRcolor0[947]&LFSRcolor0[785]&LFSRcolor0[14]&LFSRcolor0[226]);
    BiasedRNG[179] = (LFSRcolor0[166]&LFSRcolor0[1121]&LFSRcolor0[246]&LFSRcolor0[642]);
    BiasedRNG[180] = (LFSRcolor0[93]&LFSRcolor0[1182]&LFSRcolor0[1036]&LFSRcolor0[1311]);
    BiasedRNG[181] = (LFSRcolor0[345]&LFSRcolor0[710]&LFSRcolor0[1171]&LFSRcolor0[486]);
    BiasedRNG[182] = (LFSRcolor0[207]&LFSRcolor0[950]&LFSRcolor0[650]&LFSRcolor0[537]);
    BiasedRNG[183] = (LFSRcolor0[1100]&LFSRcolor0[499]&LFSRcolor0[739]&LFSRcolor0[269]);
    BiasedRNG[184] = (LFSRcolor0[490]&LFSRcolor0[1206]&LFSRcolor0[1153]&LFSRcolor0[1046]);
    BiasedRNG[185] = (LFSRcolor0[130]&LFSRcolor0[920]&LFSRcolor0[173]&LFSRcolor0[396]);
    BiasedRNG[186] = (LFSRcolor0[605]&LFSRcolor0[264]&LFSRcolor0[634]&LFSRcolor0[654]);
    BiasedRNG[187] = (LFSRcolor0[18]&LFSRcolor0[665]&LFSRcolor0[1232]&LFSRcolor0[1286]);
    BiasedRNG[188] = (LFSRcolor0[1292]&LFSRcolor0[90]&LFSRcolor0[354]&LFSRcolor0[163]);
    BiasedRNG[189] = (LFSRcolor0[473]&LFSRcolor0[131]&LFSRcolor0[375]&LFSRcolor0[1165]);
    BiasedRNG[190] = (LFSRcolor0[398]&LFSRcolor0[1264]&LFSRcolor0[223]&LFSRcolor0[822]);
    BiasedRNG[191] = (LFSRcolor0[592]&LFSRcolor0[180]&LFSRcolor0[1144]&LFSRcolor0[722]);
    BiasedRNG[192] = (LFSRcolor0[684]&LFSRcolor0[672]&LFSRcolor0[630]&LFSRcolor0[660]);
    BiasedRNG[193] = (LFSRcolor0[538]&LFSRcolor0[320]&LFSRcolor0[1089]&LFSRcolor0[923]);
    BiasedRNG[194] = (LFSRcolor0[104]&LFSRcolor0[831]&LFSRcolor0[693]&LFSRcolor0[471]);
    BiasedRNG[195] = (LFSRcolor0[701]&LFSRcolor0[998]&LFSRcolor0[689]&LFSRcolor0[964]);
    BiasedRNG[196] = (LFSRcolor0[670]&LFSRcolor0[1010]&LFSRcolor0[1254]&LFSRcolor0[1095]);
    BiasedRNG[197] = (LFSRcolor0[913]&LFSRcolor0[71]&LFSRcolor0[139]&LFSRcolor0[737]);
    BiasedRNG[198] = (LFSRcolor0[994]&LFSRcolor0[21]&LFSRcolor0[719]&LFSRcolor0[1104]);
    BiasedRNG[199] = (LFSRcolor0[96]&LFSRcolor0[887]&LFSRcolor0[644]&LFSRcolor0[203]);
    BiasedRNG[200] = (LFSRcolor0[1258]&LFSRcolor0[751]&LFSRcolor0[604]&LFSRcolor0[855]);
    BiasedRNG[201] = (LFSRcolor0[989]&LFSRcolor0[74]&LFSRcolor0[439]&LFSRcolor0[161]);
    BiasedRNG[202] = (LFSRcolor0[335]&LFSRcolor0[199]&LFSRcolor0[1227]&LFSRcolor0[711]);
    BiasedRNG[203] = (LFSRcolor0[1074]&LFSRcolor0[1076]&LFSRcolor0[286]&LFSRcolor0[1086]);
    BiasedRNG[204] = (LFSRcolor0[1193]&LFSRcolor0[1003]&LFSRcolor0[377]&LFSRcolor0[844]);
    BiasedRNG[205] = (LFSRcolor0[1]&LFSRcolor0[968]&LFSRcolor0[469]&LFSRcolor0[441]);
    BiasedRNG[206] = (LFSRcolor0[625]&LFSRcolor0[266]&LFSRcolor0[97]&LFSRcolor0[261]);
    BiasedRNG[207] = (LFSRcolor0[986]&LFSRcolor0[122]&LFSRcolor0[291]&LFSRcolor0[974]);
    BiasedRNG[208] = (LFSRcolor0[1214]&LFSRcolor0[454]&LFSRcolor0[382]&LFSRcolor0[817]);
    BiasedRNG[209] = (LFSRcolor0[183]&LFSRcolor0[781]&LFSRcolor0[1271]&LFSRcolor0[3]);
    BiasedRNG[210] = (LFSRcolor0[323]&LFSRcolor0[988]&LFSRcolor0[383]&LFSRcolor0[1235]);
    BiasedRNG[211] = (LFSRcolor0[1267]&LFSRcolor0[192]&LFSRcolor0[15]&LFSRcolor0[1289]);
    BiasedRNG[212] = (LFSRcolor0[765]&LFSRcolor0[951]&LFSRcolor0[420]&LFSRcolor0[85]);
    BiasedRNG[213] = (LFSRcolor0[1331]&LFSRcolor0[358]&LFSRcolor0[704]&LFSRcolor0[626]);
    BiasedRNG[214] = (LFSRcolor0[958]&LFSRcolor0[529]&LFSRcolor0[263]&LFSRcolor0[1261]);
    BiasedRNG[215] = (LFSRcolor0[218]&LFSRcolor0[343]&LFSRcolor0[635]&LFSRcolor0[310]);
    BiasedRNG[216] = (LFSRcolor0[553]&LFSRcolor0[1294]&LFSRcolor0[1248]&LFSRcolor0[715]);
    BiasedRNG[217] = (LFSRcolor0[1304]&LFSRcolor0[344]&LFSRcolor0[136]&LFSRcolor0[1325]);
    BiasedRNG[218] = (LFSRcolor0[567]&LFSRcolor0[1199]&LFSRcolor0[769]&LFSRcolor0[657]);
    BiasedRNG[219] = (LFSRcolor0[1195]&LFSRcolor0[7]&LFSRcolor0[290]&LFSRcolor0[683]);
    BiasedRNG[220] = (LFSRcolor0[184]&LFSRcolor0[526]&LFSRcolor0[1252]&LFSRcolor0[479]);
    BiasedRNG[221] = (LFSRcolor0[905]&LFSRcolor0[1219]&LFSRcolor0[1279]&LFSRcolor0[886]);
    BiasedRNG[222] = (LFSRcolor0[603]&LFSRcolor0[435]&LFSRcolor0[990]&LFSRcolor0[669]);
    BiasedRNG[223] = (LFSRcolor0[115]&LFSRcolor0[16]&LFSRcolor0[970]&LFSRcolor0[151]);
    BiasedRNG[224] = (LFSRcolor0[1115]&LFSRcolor0[1191]&LFSRcolor0[810]&LFSRcolor0[155]);
    BiasedRNG[225] = (LFSRcolor0[778]&LFSRcolor0[726]&LFSRcolor0[421]&LFSRcolor0[1047]);
    BiasedRNG[226] = (LFSRcolor0[206]&LFSRcolor0[443]&LFSRcolor0[949]&LFSRcolor0[841]);
    BiasedRNG[227] = (LFSRcolor0[468]&LFSRcolor0[1088]&LFSRcolor0[1034]&LFSRcolor0[284]);
    BiasedRNG[228] = (LFSRcolor0[379]&LFSRcolor0[414]&LFSRcolor0[198]&LFSRcolor0[1298]);
    BiasedRNG[229] = (LFSRcolor0[588]&LFSRcolor0[835]&LFSRcolor0[1308]&LFSRcolor0[43]);
    BiasedRNG[230] = (LFSRcolor0[932]&LFSRcolor0[399]&LFSRcolor0[229]&LFSRcolor0[1175]);
    BiasedRNG[231] = (LFSRcolor0[1262]&LFSRcolor0[337]&LFSRcolor0[1079]&LFSRcolor0[221]);
    BiasedRNG[232] = (LFSRcolor0[1146]&LFSRcolor0[127]&LFSRcolor0[1242]&LFSRcolor0[257]);
    BiasedRNG[233] = (LFSRcolor0[283]&LFSRcolor0[427]&LFSRcolor0[633]&LFSRcolor0[843]);
    BiasedRNG[234] = (LFSRcolor0[965]&LFSRcolor0[742]&LFSRcolor0[338]&LFSRcolor0[413]);
    BiasedRNG[235] = (LFSRcolor0[926]&LFSRcolor0[1315]&LFSRcolor0[1223]&LFSRcolor0[1097]);
    BiasedRNG[236] = (LFSRcolor0[980]&LFSRcolor0[403]&LFSRcolor0[369]&LFSRcolor0[516]);
    BiasedRNG[237] = (LFSRcolor0[1080]&LFSRcolor0[460]&LFSRcolor0[103]&LFSRcolor0[232]);
    BiasedRNG[238] = (LFSRcolor0[873]&LFSRcolor0[376]&LFSRcolor0[307]&LFSRcolor0[532]);
    BiasedRNG[239] = (LFSRcolor0[474]&LFSRcolor0[1015]&LFSRcolor0[386]&LFSRcolor0[407]);
    BiasedRNG[240] = (LFSRcolor0[961]&LFSRcolor0[952]&LFSRcolor0[985]&LFSRcolor0[1234]);
    BiasedRNG[241] = (LFSRcolor0[543]&LFSRcolor0[245]&LFSRcolor0[99]&LFSRcolor0[530]);
    BiasedRNG[242] = (LFSRcolor0[428]&LFSRcolor0[1237]&LFSRcolor0[847]&LFSRcolor0[72]);
    BiasedRNG[243] = (LFSRcolor0[1187]&LFSRcolor0[678]&LFSRcolor0[774]&LFSRcolor0[967]);
    BiasedRNG[244] = (LFSRcolor0[1332]&LFSRcolor0[37]&LFSRcolor0[503]&LFSRcolor0[1326]);
    BiasedRNG[245] = (LFSRcolor0[86]&LFSRcolor0[181]&LFSRcolor0[826]&LFSRcolor0[942]);
    BiasedRNG[246] = (LFSRcolor0[1159]&LFSRcolor0[297]&LFSRcolor0[694]&LFSRcolor0[1152]);
    BiasedRNG[247] = (LFSRcolor0[572]&LFSRcolor0[1309]&LFSRcolor0[566]&LFSRcolor0[1108]);
    BiasedRNG[248] = (LFSRcolor0[893]&LFSRcolor0[8]&LFSRcolor0[1044]&LFSRcolor0[314]);
    BiasedRNG[249] = (LFSRcolor0[1131]&LFSRcolor0[182]&LFSRcolor0[75]&LFSRcolor0[59]);
    BiasedRNG[250] = (LFSRcolor0[1083]&LFSRcolor0[641]&LFSRcolor0[897]&LFSRcolor0[107]);
    BiasedRNG[251] = (LFSRcolor0[687]&LFSRcolor0[743]&LFSRcolor0[1169]&LFSRcolor0[610]);
    BiasedRNG[252] = (LFSRcolor0[1259]&LFSRcolor0[61]&LFSRcolor0[676]&LFSRcolor0[1224]);
    BiasedRNG[253] = (LFSRcolor0[514]&LFSRcolor0[995]&LFSRcolor0[481]&LFSRcolor0[1173]);
    BiasedRNG[254] = (LFSRcolor0[1307]&LFSRcolor0[915]&LFSRcolor0[565]&LFSRcolor0[475]);
    BiasedRNG[255] = (LFSRcolor0[937]&LFSRcolor0[309]&LFSRcolor0[1204]&LFSRcolor0[410]);
    UnbiasedRNG[0] = LFSRcolor0[586];
    UnbiasedRNG[1] = LFSRcolor0[282];
    UnbiasedRNG[2] = LFSRcolor0[861];
    UnbiasedRNG[3] = LFSRcolor0[1166];
    UnbiasedRNG[4] = LFSRcolor0[1084];
    UnbiasedRNG[5] = LFSRcolor0[215];
    UnbiasedRNG[6] = LFSRcolor0[265];
    UnbiasedRNG[7] = LFSRcolor0[143];
    UnbiasedRNG[8] = LFSRcolor0[1150];
    UnbiasedRNG[9] = LFSRcolor0[55];
    UnbiasedRNG[10] = LFSRcolor0[1215];
    UnbiasedRNG[11] = LFSRcolor0[1000];
    UnbiasedRNG[12] = LFSRcolor0[216];
    UnbiasedRNG[13] = LFSRcolor0[196];
    UnbiasedRNG[14] = LFSRcolor0[833];
    UnbiasedRNG[15] = LFSRcolor0[725];
    UnbiasedRNG[16] = LFSRcolor0[736];
    UnbiasedRNG[17] = LFSRcolor0[1073];
    UnbiasedRNG[18] = LFSRcolor0[564];
    UnbiasedRNG[19] = LFSRcolor0[300];
    UnbiasedRNG[20] = LFSRcolor0[1035];
    UnbiasedRNG[21] = LFSRcolor0[510];
    UnbiasedRNG[22] = LFSRcolor0[622];
    UnbiasedRNG[23] = LFSRcolor0[1310];
    UnbiasedRNG[24] = LFSRcolor0[387];
    UnbiasedRNG[25] = LFSRcolor0[227];
    UnbiasedRNG[26] = LFSRcolor0[1320];
    UnbiasedRNG[27] = LFSRcolor0[1205];
    UnbiasedRNG[28] = LFSRcolor0[979];
    UnbiasedRNG[29] = LFSRcolor0[1316];
    UnbiasedRNG[30] = LFSRcolor0[922];
    UnbiasedRNG[31] = LFSRcolor0[1125];
    UnbiasedRNG[32] = LFSRcolor0[1312];
    UnbiasedRNG[33] = LFSRcolor0[306];
    UnbiasedRNG[34] = LFSRcolor0[200];
    UnbiasedRNG[35] = LFSRcolor0[682];
    UnbiasedRNG[36] = LFSRcolor0[1266];
    UnbiasedRNG[37] = LFSRcolor0[483];
    UnbiasedRNG[38] = LFSRcolor0[39];
    UnbiasedRNG[39] = LFSRcolor0[1189];
    UnbiasedRNG[40] = LFSRcolor0[190];
    UnbiasedRNG[41] = LFSRcolor0[1327];
    UnbiasedRNG[42] = LFSRcolor0[1183];
    UnbiasedRNG[43] = LFSRcolor0[362];
    UnbiasedRNG[44] = LFSRcolor0[1147];
    UnbiasedRNG[45] = LFSRcolor0[1138];
    UnbiasedRNG[46] = LFSRcolor0[406];
    UnbiasedRNG[47] = LFSRcolor0[1176];
    UnbiasedRNG[48] = LFSRcolor0[154];
    UnbiasedRNG[49] = LFSRcolor0[801];
    UnbiasedRNG[50] = LFSRcolor0[249];
    UnbiasedRNG[51] = LFSRcolor0[646];
    UnbiasedRNG[52] = LFSRcolor0[1105];
    UnbiasedRNG[53] = LFSRcolor0[585];
    UnbiasedRNG[54] = LFSRcolor0[1196];
    UnbiasedRNG[55] = LFSRcolor0[996];
    UnbiasedRNG[56] = LFSRcolor0[1055];
    UnbiasedRNG[57] = LFSRcolor0[186];
    UnbiasedRNG[58] = LFSRcolor0[759];
    UnbiasedRNG[59] = LFSRcolor0[1063];
    UnbiasedRNG[60] = LFSRcolor0[1123];
    UnbiasedRNG[61] = LFSRcolor0[823];
    UnbiasedRNG[62] = LFSRcolor0[4];
    UnbiasedRNG[63] = LFSRcolor0[1026];
    UnbiasedRNG[64] = LFSRcolor0[1218];
    UnbiasedRNG[65] = LFSRcolor0[250];
    UnbiasedRNG[66] = LFSRcolor0[928];
    UnbiasedRNG[67] = LFSRcolor0[240];
    UnbiasedRNG[68] = LFSRcolor0[53];
    UnbiasedRNG[69] = LFSRcolor0[1157];
    UnbiasedRNG[70] = LFSRcolor0[1244];
    UnbiasedRNG[71] = LFSRcolor0[114];
    UnbiasedRNG[72] = LFSRcolor0[487];
    UnbiasedRNG[73] = LFSRcolor0[780];
    UnbiasedRNG[74] = LFSRcolor0[397];
    UnbiasedRNG[75] = LFSRcolor0[278];
    UnbiasedRNG[76] = LFSRcolor0[135];
    UnbiasedRNG[77] = LFSRcolor0[329];
    UnbiasedRNG[78] = LFSRcolor0[1221];
    UnbiasedRNG[79] = LFSRcolor0[38];
    UnbiasedRNG[80] = LFSRcolor0[636];
    UnbiasedRNG[81] = LFSRcolor0[222];
    UnbiasedRNG[82] = LFSRcolor0[395];
    UnbiasedRNG[83] = LFSRcolor0[981];
    UnbiasedRNG[84] = LFSRcolor0[137];
    UnbiasedRNG[85] = LFSRcolor0[900];
    UnbiasedRNG[86] = LFSRcolor0[1140];
    UnbiasedRNG[87] = LFSRcolor0[380];
    UnbiasedRNG[88] = LFSRcolor0[292];
    UnbiasedRNG[89] = LFSRcolor0[1142];
    UnbiasedRNG[90] = LFSRcolor0[938];
    UnbiasedRNG[91] = LFSRcolor0[5];
    UnbiasedRNG[92] = LFSRcolor0[662];
    UnbiasedRNG[93] = LFSRcolor0[374];
    UnbiasedRNG[94] = LFSRcolor0[953];
    UnbiasedRNG[95] = LFSRcolor0[569];
    UnbiasedRNG[96] = LFSRcolor0[1268];
    UnbiasedRNG[97] = LFSRcolor0[1197];
    UnbiasedRNG[98] = LFSRcolor0[789];
    UnbiasedRNG[99] = LFSRcolor0[1033];
    UnbiasedRNG[100] = LFSRcolor0[1052];
    UnbiasedRNG[101] = LFSRcolor0[463];
    UnbiasedRNG[102] = LFSRcolor0[467];
    UnbiasedRNG[103] = LFSRcolor0[231];
    UnbiasedRNG[104] = LFSRcolor0[623];
    UnbiasedRNG[105] = LFSRcolor0[792];
    UnbiasedRNG[106] = LFSRcolor0[776];
    UnbiasedRNG[107] = LFSRcolor0[273];
    UnbiasedRNG[108] = LFSRcolor0[917];
    UnbiasedRNG[109] = LFSRcolor0[174];
    UnbiasedRNG[110] = LFSRcolor0[1179];
    UnbiasedRNG[111] = LFSRcolor0[1303];
    UnbiasedRNG[112] = LFSRcolor0[1241];
    UnbiasedRNG[113] = LFSRcolor0[144];
    UnbiasedRNG[114] = LFSRcolor0[559];
    UnbiasedRNG[115] = LFSRcolor0[536];
    UnbiasedRNG[116] = LFSRcolor0[881];
    UnbiasedRNG[117] = LFSRcolor0[697];
    UnbiasedRNG[118] = LFSRcolor0[1287];
    UnbiasedRNG[119] = LFSRcolor0[361];
    UnbiasedRNG[120] = LFSRcolor0[716];
    UnbiasedRNG[121] = LFSRcolor0[461];
    UnbiasedRNG[122] = LFSRcolor0[888];
    UnbiasedRNG[123] = LFSRcolor0[912];
    UnbiasedRNG[124] = LFSRcolor0[852];
    UnbiasedRNG[125] = LFSRcolor0[1133];
    UnbiasedRNG[126] = LFSRcolor0[579];
    UnbiasedRNG[127] = LFSRcolor0[177];
    UnbiasedRNG[128] = LFSRcolor0[275];
    UnbiasedRNG[129] = LFSRcolor0[1265];
    UnbiasedRNG[130] = LFSRcolor0[505];
    UnbiasedRNG[131] = LFSRcolor0[1006];
    UnbiasedRNG[132] = LFSRcolor0[12];
    UnbiasedRNG[133] = LFSRcolor0[1249];
    UnbiasedRNG[134] = LFSRcolor0[48];
    UnbiasedRNG[135] = LFSRcolor0[311];
    UnbiasedRNG[136] = LFSRcolor0[138];
    UnbiasedRNG[137] = LFSRcolor0[944];
    UnbiasedRNG[138] = LFSRcolor0[819];
    UnbiasedRNG[139] = LFSRcolor0[1305];
    UnbiasedRNG[140] = LFSRcolor0[430];
    UnbiasedRNG[141] = LFSRcolor0[573];
    UnbiasedRNG[142] = LFSRcolor0[1282];
    UnbiasedRNG[143] = LFSRcolor0[1226];
    UnbiasedRNG[144] = LFSRcolor0[1134];
    UnbiasedRNG[145] = LFSRcolor0[554];
    UnbiasedRNG[146] = LFSRcolor0[706];
    UnbiasedRNG[147] = LFSRcolor0[674];
    UnbiasedRNG[148] = LFSRcolor0[194];
    UnbiasedRNG[149] = LFSRcolor0[1273];
    UnbiasedRNG[150] = LFSRcolor0[859];
    UnbiasedRNG[151] = LFSRcolor0[745];
    UnbiasedRNG[152] = LFSRcolor0[717];
    UnbiasedRNG[153] = LFSRcolor0[1061];
    UnbiasedRNG[154] = LFSRcolor0[782];
    UnbiasedRNG[155] = LFSRcolor0[904];
    UnbiasedRNG[156] = LFSRcolor0[651];
    UnbiasedRNG[157] = LFSRcolor0[816];
    UnbiasedRNG[158] = LFSRcolor0[1091];
    UnbiasedRNG[159] = LFSRcolor0[1039];
    UnbiasedRNG[160] = LFSRcolor0[969];
    UnbiasedRNG[161] = LFSRcolor0[1174];
    UnbiasedRNG[162] = LFSRcolor0[201];
    UnbiasedRNG[163] = LFSRcolor0[1323];
    UnbiasedRNG[164] = LFSRcolor0[924];
    UnbiasedRNG[165] = LFSRcolor0[890];
    UnbiasedRNG[166] = LFSRcolor0[1051];
    UnbiasedRNG[167] = LFSRcolor0[423];
    UnbiasedRNG[168] = LFSRcolor0[842];
    UnbiasedRNG[169] = LFSRcolor0[302];
    UnbiasedRNG[170] = LFSRcolor0[162];
    UnbiasedRNG[171] = LFSRcolor0[875];
    UnbiasedRNG[172] = LFSRcolor0[796];
    UnbiasedRNG[173] = LFSRcolor0[872];
    UnbiasedRNG[174] = LFSRcolor0[23];
    UnbiasedRNG[175] = LFSRcolor0[1110];
    UnbiasedRNG[176] = LFSRcolor0[1299];
    UnbiasedRNG[177] = LFSRcolor0[649];
    UnbiasedRNG[178] = LFSRcolor0[169];
    UnbiasedRNG[179] = LFSRcolor0[552];
    UnbiasedRNG[180] = LFSRcolor0[729];
    UnbiasedRNG[181] = LFSRcolor0[1037];
    UnbiasedRNG[182] = LFSRcolor0[1210];
    UnbiasedRNG[183] = LFSRcolor0[1024];
    UnbiasedRNG[184] = LFSRcolor0[712];
    UnbiasedRNG[185] = LFSRcolor0[702];
    UnbiasedRNG[186] = LFSRcolor0[63];
    UnbiasedRNG[187] = LFSRcolor0[867];
    UnbiasedRNG[188] = LFSRcolor0[645];
    UnbiasedRNG[189] = LFSRcolor0[480];
    UnbiasedRNG[190] = LFSRcolor0[929];
    UnbiasedRNG[191] = LFSRcolor0[1198];
    UnbiasedRNG[192] = LFSRcolor0[251];
    UnbiasedRNG[193] = LFSRcolor0[714];
    UnbiasedRNG[194] = LFSRcolor0[1319];
    UnbiasedRNG[195] = LFSRcolor0[1213];
    UnbiasedRNG[196] = LFSRcolor0[117];
    UnbiasedRNG[197] = LFSRcolor0[836];
    UnbiasedRNG[198] = LFSRcolor0[540];
    UnbiasedRNG[199] = LFSRcolor0[577];
    UnbiasedRNG[200] = LFSRcolor0[164];
    UnbiasedRNG[201] = LFSRcolor0[412];
    UnbiasedRNG[202] = LFSRcolor0[1019];
    UnbiasedRNG[203] = LFSRcolor0[838];
    UnbiasedRNG[204] = LFSRcolor0[371];
    UnbiasedRNG[205] = LFSRcolor0[730];
    UnbiasedRNG[206] = LFSRcolor0[1151];
    UnbiasedRNG[207] = LFSRcolor0[1040];
    UnbiasedRNG[208] = LFSRcolor0[1107];
    UnbiasedRNG[209] = LFSRcolor0[1071];
    UnbiasedRNG[210] = LFSRcolor0[1087];
    UnbiasedRNG[211] = LFSRcolor0[365];
    UnbiasedRNG[212] = LFSRcolor0[738];
    UnbiasedRNG[213] = LFSRcolor0[150];
    UnbiasedRNG[214] = LFSRcolor0[954];
    UnbiasedRNG[215] = LFSRcolor0[1075];
    UnbiasedRNG[216] = LFSRcolor0[267];
    UnbiasedRNG[217] = LFSRcolor0[1231];
    UnbiasedRNG[218] = LFSRcolor0[513];
    UnbiasedRNG[219] = LFSRcolor0[29];
    UnbiasedRNG[220] = LFSRcolor0[1077];
    UnbiasedRNG[221] = LFSRcolor0[1050];
    UnbiasedRNG[222] = LFSRcolor0[77];
    UnbiasedRNG[223] = LFSRcolor0[1116];
    UnbiasedRNG[224] = LFSRcolor0[158];
    UnbiasedRNG[225] = LFSRcolor0[52];
    UnbiasedRNG[226] = LFSRcolor0[653];
    UnbiasedRNG[227] = LFSRcolor0[723];
    UnbiasedRNG[228] = LFSRcolor0[1014];
    UnbiasedRNG[229] = LFSRcolor0[976];
    UnbiasedRNG[230] = LFSRcolor0[167];
    UnbiasedRNG[231] = LFSRcolor0[341];
    UnbiasedRNG[232] = LFSRcolor0[419];
    UnbiasedRNG[233] = LFSRcolor0[511];
    UnbiasedRNG[234] = LFSRcolor0[176];
    UnbiasedRNG[235] = LFSRcolor0[997];
    UnbiasedRNG[236] = LFSRcolor0[903];
    UnbiasedRNG[237] = LFSRcolor0[1167];
    UnbiasedRNG[238] = LFSRcolor0[731];
    UnbiasedRNG[239] = LFSRcolor0[1025];
    UnbiasedRNG[240] = LFSRcolor0[916];
    UnbiasedRNG[241] = LFSRcolor0[322];
    UnbiasedRNG[242] = LFSRcolor0[426];
    UnbiasedRNG[243] = LFSRcolor0[1113];
    UnbiasedRNG[244] = LFSRcolor0[332];
    UnbiasedRNG[245] = LFSRcolor0[1099];
    UnbiasedRNG[246] = LFSRcolor0[495];
    UnbiasedRNG[247] = LFSRcolor0[638];
    UnbiasedRNG[248] = LFSRcolor0[188];
    UnbiasedRNG[249] = LFSRcolor0[1246];
    UnbiasedRNG[250] = LFSRcolor0[13];
    UnbiasedRNG[251] = LFSRcolor0[1233];
    UnbiasedRNG[252] = LFSRcolor0[910];
    UnbiasedRNG[253] = LFSRcolor0[402];
    UnbiasedRNG[254] = LFSRcolor0[348];
    UnbiasedRNG[255] = LFSRcolor0[773];
    UnbiasedRNG[256] = LFSRcolor0[1023];
    UnbiasedRNG[257] = LFSRcolor0[804];
    UnbiasedRNG[258] = LFSRcolor0[305];
    UnbiasedRNG[259] = LFSRcolor0[1236];
    UnbiasedRNG[260] = LFSRcolor0[1274];
    UnbiasedRNG[261] = LFSRcolor0[749];
    UnbiasedRNG[262] = LFSRcolor0[845];
    UnbiasedRNG[263] = LFSRcolor0[772];
    UnbiasedRNG[264] = LFSRcolor0[455];
    UnbiasedRNG[265] = LFSRcolor0[1111];
    UnbiasedRNG[266] = LFSRcolor0[327];
    UnbiasedRNG[267] = LFSRcolor0[235];
    UnbiasedRNG[268] = LFSRcolor0[648];
    UnbiasedRNG[269] = LFSRcolor0[555];
    UnbiasedRNG[270] = LFSRcolor0[288];
end

always @(posedge color0_clk) begin
    BiasedRNG[256] = (LFSRcolor1[265]&LFSRcolor1[1438]&LFSRcolor1[1081]&LFSRcolor1[1640]);
    BiasedRNG[257] = (LFSRcolor1[1124]&LFSRcolor1[1689]&LFSRcolor1[4]&LFSRcolor1[208]);
    BiasedRNG[258] = (LFSRcolor1[602]&LFSRcolor1[1696]&LFSRcolor1[1574]&LFSRcolor1[447]);
    BiasedRNG[259] = (LFSRcolor1[1773]&LFSRcolor1[1615]&LFSRcolor1[745]&LFSRcolor1[1333]);
    BiasedRNG[260] = (LFSRcolor1[1616]&LFSRcolor1[1493]&LFSRcolor1[327]&LFSRcolor1[234]);
    BiasedRNG[261] = (LFSRcolor1[1722]&LFSRcolor1[860]&LFSRcolor1[1406]&LFSRcolor1[1661]);
    BiasedRNG[262] = (LFSRcolor1[459]&LFSRcolor1[1684]&LFSRcolor1[674]&LFSRcolor1[686]);
    BiasedRNG[263] = (LFSRcolor1[1112]&LFSRcolor1[1668]&LFSRcolor1[1035]&LFSRcolor1[71]);
    BiasedRNG[264] = (LFSRcolor1[2]&LFSRcolor1[1259]&LFSRcolor1[1651]&LFSRcolor1[954]);
    BiasedRNG[265] = (LFSRcolor1[730]&LFSRcolor1[1290]&LFSRcolor1[1256]&LFSRcolor1[1061]);
    BiasedRNG[266] = (LFSRcolor1[1404]&LFSRcolor1[1146]&LFSRcolor1[256]&LFSRcolor1[1449]);
    BiasedRNG[267] = (LFSRcolor1[1141]&LFSRcolor1[717]&LFSRcolor1[165]&LFSRcolor1[1709]);
    BiasedRNG[268] = (LFSRcolor1[98]&LFSRcolor1[1046]&LFSRcolor1[1360]&LFSRcolor1[123]);
    BiasedRNG[269] = (LFSRcolor1[1350]&LFSRcolor1[758]&LFSRcolor1[461]&LFSRcolor1[1136]);
    BiasedRNG[270] = (LFSRcolor1[1443]&LFSRcolor1[693]&LFSRcolor1[400]&LFSRcolor1[689]);
    BiasedRNG[271] = (LFSRcolor1[205]&LFSRcolor1[1174]&LFSRcolor1[403]&LFSRcolor1[1473]);
    BiasedRNG[272] = (LFSRcolor1[470]&LFSRcolor1[1636]&LFSRcolor1[247]&LFSRcolor1[1535]);
    BiasedRNG[273] = (LFSRcolor1[785]&LFSRcolor1[856]&LFSRcolor1[985]&LFSRcolor1[539]);
    BiasedRNG[274] = (LFSRcolor1[1508]&LFSRcolor1[1400]&LFSRcolor1[1422]&LFSRcolor1[8]);
    BiasedRNG[275] = (LFSRcolor1[616]&LFSRcolor1[24]&LFSRcolor1[775]&LFSRcolor1[408]);
    BiasedRNG[276] = (LFSRcolor1[1056]&LFSRcolor1[570]&LFSRcolor1[1240]&LFSRcolor1[1315]);
    BiasedRNG[277] = (LFSRcolor1[1392]&LFSRcolor1[527]&LFSRcolor1[336]&LFSRcolor1[1424]);
    BiasedRNG[278] = (LFSRcolor1[1247]&LFSRcolor1[1733]&LFSRcolor1[1526]&LFSRcolor1[1725]);
    BiasedRNG[279] = (LFSRcolor1[1691]&LFSRcolor1[473]&LFSRcolor1[1243]&LFSRcolor1[180]);
    BiasedRNG[280] = (LFSRcolor1[706]&LFSRcolor1[101]&LFSRcolor1[1569]&LFSRcolor1[436]);
    BiasedRNG[281] = (LFSRcolor1[409]&LFSRcolor1[680]&LFSRcolor1[608]&LFSRcolor1[1450]);
    BiasedRNG[282] = (LFSRcolor1[574]&LFSRcolor1[1425]&LFSRcolor1[1628]&LFSRcolor1[115]);
    BiasedRNG[283] = (LFSRcolor1[892]&LFSRcolor1[1102]&LFSRcolor1[1657]&LFSRcolor1[57]);
    BiasedRNG[284] = (LFSRcolor1[543]&LFSRcolor1[1228]&LFSRcolor1[827]&LFSRcolor1[1652]);
    BiasedRNG[285] = (LFSRcolor1[232]&LFSRcolor1[1180]&LFSRcolor1[1492]&LFSRcolor1[586]);
    BiasedRNG[286] = (LFSRcolor1[688]&LFSRcolor1[261]&LFSRcolor1[972]&LFSRcolor1[545]);
    BiasedRNG[287] = (LFSRcolor1[924]&LFSRcolor1[1052]&LFSRcolor1[139]&LFSRcolor1[503]);
    BiasedRNG[288] = (LFSRcolor1[1607]&LFSRcolor1[1195]&LFSRcolor1[1674]&LFSRcolor1[1059]);
    BiasedRNG[289] = (LFSRcolor1[1557]&LFSRcolor1[1467]&LFSRcolor1[1591]&LFSRcolor1[1504]);
    BiasedRNG[290] = (LFSRcolor1[508]&LFSRcolor1[561]&LFSRcolor1[429]&LFSRcolor1[1008]);
    BiasedRNG[291] = (LFSRcolor1[1369]&LFSRcolor1[1731]&LFSRcolor1[1030]&LFSRcolor1[1118]);
    BiasedRNG[292] = (LFSRcolor1[721]&LFSRcolor1[1439]&LFSRcolor1[460]&LFSRcolor1[1649]);
    BiasedRNG[293] = (LFSRcolor1[83]&LFSRcolor1[1673]&LFSRcolor1[883]&LFSRcolor1[1074]);
    BiasedRNG[294] = (LFSRcolor1[536]&LFSRcolor1[1643]&LFSRcolor1[1749]&LFSRcolor1[264]);
    BiasedRNG[295] = (LFSRcolor1[908]&LFSRcolor1[426]&LFSRcolor1[1275]&LFSRcolor1[1561]);
    BiasedRNG[296] = (LFSRcolor1[450]&LFSRcolor1[1343]&LFSRcolor1[1476]&LFSRcolor1[1381]);
    BiasedRNG[297] = (LFSRcolor1[238]&LFSRcolor1[287]&LFSRcolor1[798]&LFSRcolor1[214]);
    BiasedRNG[298] = (LFSRcolor1[1599]&LFSRcolor1[1262]&LFSRcolor1[431]&LFSRcolor1[19]);
    BiasedRNG[299] = (LFSRcolor1[1325]&LFSRcolor1[1051]&LFSRcolor1[476]&LFSRcolor1[617]);
    BiasedRNG[300] = (LFSRcolor1[366]&LFSRcolor1[1276]&LFSRcolor1[913]&LFSRcolor1[834]);
    BiasedRNG[301] = (LFSRcolor1[1700]&LFSRcolor1[812]&LFSRcolor1[184]&LFSRcolor1[458]);
    BiasedRNG[302] = (LFSRcolor1[1190]&LFSRcolor1[1341]&LFSRcolor1[1328]&LFSRcolor1[41]);
    BiasedRNG[303] = (LFSRcolor1[708]&LFSRcolor1[696]&LFSRcolor1[894]&LFSRcolor1[504]);
    BiasedRNG[304] = (LFSRcolor1[289]&LFSRcolor1[1172]&LFSRcolor1[505]&LFSRcolor1[992]);
    BiasedRNG[305] = (LFSRcolor1[500]&LFSRcolor1[278]&LFSRcolor1[67]&LFSRcolor1[1274]);
    BiasedRNG[306] = (LFSRcolor1[698]&LFSRcolor1[765]&LFSRcolor1[229]&LFSRcolor1[1047]);
    BiasedRNG[307] = (LFSRcolor1[1025]&LFSRcolor1[750]&LFSRcolor1[1735]&LFSRcolor1[1101]);
    BiasedRNG[308] = (LFSRcolor1[420]&LFSRcolor1[286]&LFSRcolor1[653]&LFSRcolor1[1017]);
    BiasedRNG[309] = (LFSRcolor1[1223]&LFSRcolor1[1384]&LFSRcolor1[89]&LFSRcolor1[1241]);
    BiasedRNG[310] = (LFSRcolor1[726]&LFSRcolor1[1265]&LFSRcolor1[112]&LFSRcolor1[1553]);
    BiasedRNG[311] = (LFSRcolor1[1785]&LFSRcolor1[915]&LFSRcolor1[874]&LFSRcolor1[996]);
    BiasedRNG[312] = (LFSRcolor1[1686]&LFSRcolor1[725]&LFSRcolor1[1612]&LFSRcolor1[937]);
    BiasedRNG[313] = (LFSRcolor1[890]&LFSRcolor1[227]&LFSRcolor1[772]&LFSRcolor1[660]);
    BiasedRNG[314] = (LFSRcolor1[490]&LFSRcolor1[948]&LFSRcolor1[18]&LFSRcolor1[567]);
    BiasedRNG[315] = (LFSRcolor1[451]&LFSRcolor1[1373]&LFSRcolor1[1159]&LFSRcolor1[1489]);
    BiasedRNG[316] = (LFSRcolor1[957]&LFSRcolor1[1513]&LFSRcolor1[442]&LFSRcolor1[899]);
    BiasedRNG[317] = (LFSRcolor1[242]&LFSRcolor1[26]&LFSRcolor1[559]&LFSRcolor1[1533]);
    BiasedRNG[318] = (LFSRcolor1[789]&LFSRcolor1[170]&LFSRcolor1[1723]&LFSRcolor1[585]);
    BiasedRNG[319] = (LFSRcolor1[111]&LFSRcolor1[1710]&LFSRcolor1[484]&LFSRcolor1[638]);
    BiasedRNG[320] = (LFSRcolor1[353]&LFSRcolor1[1342]&LFSRcolor1[1311]&LFSRcolor1[72]);
    BiasedRNG[321] = (LFSRcolor1[1405]&LFSRcolor1[842]&LFSRcolor1[879]&LFSRcolor1[1633]);
    BiasedRNG[322] = (LFSRcolor1[1745]&LFSRcolor1[1507]&LFSRcolor1[1349]&LFSRcolor1[1625]);
    BiasedRNG[323] = (LFSRcolor1[1585]&LFSRcolor1[1165]&LFSRcolor1[1481]&LFSRcolor1[1727]);
    BiasedRNG[324] = (LFSRcolor1[99]&LFSRcolor1[1642]&LFSRcolor1[0]&LFSRcolor1[393]);
    BiasedRNG[325] = (LFSRcolor1[1483]&LFSRcolor1[747]&LFSRcolor1[1445]&LFSRcolor1[671]);
    BiasedRNG[326] = (LFSRcolor1[1544]&LFSRcolor1[1637]&LFSRcolor1[42]&LFSRcolor1[1313]);
    BiasedRNG[327] = (LFSRcolor1[813]&LFSRcolor1[1293]&LFSRcolor1[91]&LFSRcolor1[969]);
    BiasedRNG[328] = (LFSRcolor1[1041]&LFSRcolor1[1221]&LFSRcolor1[1094]&LFSRcolor1[627]);
    BiasedRNG[329] = (LFSRcolor1[368]&LFSRcolor1[603]&LFSRcolor1[1435]&LFSRcolor1[299]);
    BiasedRNG[330] = (LFSRcolor1[667]&LFSRcolor1[1344]&LFSRcolor1[923]&LFSRcolor1[498]);
    BiasedRNG[331] = (LFSRcolor1[774]&LFSRcolor1[1635]&LFSRcolor1[938]&LFSRcolor1[1188]);
    BiasedRNG[332] = (LFSRcolor1[802]&LFSRcolor1[1609]&LFSRcolor1[1494]&LFSRcolor1[1181]);
    BiasedRNG[333] = (LFSRcolor1[1656]&LFSRcolor1[1237]&LFSRcolor1[1490]&LFSRcolor1[1429]);
    BiasedRNG[334] = (LFSRcolor1[1571]&LFSRcolor1[358]&LFSRcolor1[11]&LFSRcolor1[791]);
    BiasedRNG[335] = (LFSRcolor1[421]&LFSRcolor1[554]&LFSRcolor1[77]&LFSRcolor1[347]);
    BiasedRNG[336] = (LFSRcolor1[1132]&LFSRcolor1[1289]&LFSRcolor1[1464]&LFSRcolor1[1201]);
    BiasedRNG[337] = (LFSRcolor1[1552]&LFSRcolor1[649]&LFSRcolor1[676]&LFSRcolor1[869]);
    BiasedRNG[338] = (LFSRcolor1[998]&LFSRcolor1[1442]&LFSRcolor1[1430]&LFSRcolor1[413]);
    BiasedRNG[339] = (LFSRcolor1[404]&LFSRcolor1[886]&LFSRcolor1[1354]&LFSRcolor1[1732]);
    BiasedRNG[340] = (LFSRcolor1[1724]&LFSRcolor1[1194]&LFSRcolor1[63]&LFSRcolor1[532]);
    BiasedRNG[341] = (LFSRcolor1[795]&LFSRcolor1[257]&LFSRcolor1[1002]&LFSRcolor1[1261]);
    BiasedRNG[342] = (LFSRcolor1[794]&LFSRcolor1[97]&LFSRcolor1[1152]&LFSRcolor1[1126]);
    BiasedRNG[343] = (LFSRcolor1[632]&LFSRcolor1[968]&LFSRcolor1[1522]&LFSRcolor1[132]);
    BiasedRNG[344] = (LFSRcolor1[22]&LFSRcolor1[878]&LFSRcolor1[1095]&LFSRcolor1[663]);
    BiasedRNG[345] = (LFSRcolor1[1378]&LFSRcolor1[204]&LFSRcolor1[399]&LFSRcolor1[583]);
    BiasedRNG[346] = (LFSRcolor1[1418]&LFSRcolor1[131]&LFSRcolor1[1768]&LFSRcolor1[1231]);
    BiasedRNG[347] = (LFSRcolor1[1060]&LFSRcolor1[613]&LFSRcolor1[1570]&LFSRcolor1[1695]);
    BiasedRNG[348] = (LFSRcolor1[363]&LFSRcolor1[32]&LFSRcolor1[321]&LFSRcolor1[736]);
    BiasedRNG[349] = (LFSRcolor1[96]&LFSRcolor1[1245]&LFSRcolor1[1119]&LFSRcolor1[876]);
    BiasedRNG[350] = (LFSRcolor1[1189]&LFSRcolor1[1105]&LFSRcolor1[1138]&LFSRcolor1[926]);
    BiasedRNG[351] = (LFSRcolor1[1605]&LFSRcolor1[1776]&LFSRcolor1[323]&LFSRcolor1[658]);
    BiasedRNG[352] = (LFSRcolor1[1516]&LFSRcolor1[1206]&LFSRcolor1[704]&LFSRcolor1[974]);
    BiasedRNG[353] = (LFSRcolor1[1498]&LFSRcolor1[1220]&LFSRcolor1[1394]&LFSRcolor1[1252]);
    BiasedRNG[354] = (LFSRcolor1[1239]&LFSRcolor1[1414]&LFSRcolor1[1639]&LFSRcolor1[1721]);
    BiasedRNG[355] = (LFSRcolor1[1043]&LFSRcolor1[1110]&LFSRcolor1[448]&LFSRcolor1[1023]);
    BiasedRNG[356] = (LFSRcolor1[1235]&LFSRcolor1[1715]&LFSRcolor1[1428]&LFSRcolor1[1743]);
    BiasedRNG[357] = (LFSRcolor1[994]&LFSRcolor1[501]&LFSRcolor1[1753]&LFSRcolor1[953]);
    BiasedRNG[358] = (LFSRcolor1[1198]&LFSRcolor1[455]&LFSRcolor1[64]&LFSRcolor1[1362]);
    BiasedRNG[359] = (LFSRcolor1[1559]&LFSRcolor1[292]&LFSRcolor1[1737]&LFSRcolor1[906]);
    BiasedRNG[360] = (LFSRcolor1[845]&LFSRcolor1[1249]&LFSRcolor1[1368]&LFSRcolor1[433]);
    BiasedRNG[361] = (LFSRcolor1[499]&LFSRcolor1[17]&LFSRcolor1[304]&LFSRcolor1[997]);
    BiasedRNG[362] = (LFSRcolor1[650]&LFSRcolor1[1408]&LFSRcolor1[1789]&LFSRcolor1[140]);
    BiasedRNG[363] = (LFSRcolor1[138]&LFSRcolor1[1560]&LFSRcolor1[1558]&LFSRcolor1[916]);
    BiasedRNG[364] = (LFSRcolor1[907]&LFSRcolor1[691]&LFSRcolor1[762]&LFSRcolor1[1326]);
    BiasedRNG[365] = (LFSRcolor1[1212]&LFSRcolor1[701]&LFSRcolor1[58]&LFSRcolor1[1503]);
    BiasedRNG[366] = (LFSRcolor1[855]&LFSRcolor1[437]&LFSRcolor1[1086]&LFSRcolor1[1312]);
    BiasedRNG[367] = (LFSRcolor1[1543]&LFSRcolor1[1401]&LFSRcolor1[1683]&LFSRcolor1[526]);
    BiasedRNG[368] = (LFSRcolor1[1462]&LFSRcolor1[237]&LFSRcolor1[578]&LFSRcolor1[777]);
    BiasedRNG[369] = (LFSRcolor1[183]&LFSRcolor1[1200]&LFSRcolor1[1440]&LFSRcolor1[1042]);
    BiasedRNG[370] = (LFSRcolor1[666]&LFSRcolor1[300]&LFSRcolor1[1109]&LFSRcolor1[1088]);
    BiasedRNG[371] = (LFSRcolor1[843]&LFSRcolor1[1031]&LFSRcolor1[1524]&LFSRcolor1[697]);
    BiasedRNG[372] = (LFSRcolor1[298]&LFSRcolor1[1143]&LFSRcolor1[1171]&LFSRcolor1[1161]);
    BiasedRNG[373] = (LFSRcolor1[1793]&LFSRcolor1[75]&LFSRcolor1[415]&LFSRcolor1[823]);
    BiasedRNG[374] = (LFSRcolor1[1595]&LFSRcolor1[418]&LFSRcolor1[528]&LFSRcolor1[659]);
    BiasedRNG[375] = (LFSRcolor1[86]&LFSRcolor1[1374]&LFSRcolor1[253]&LFSRcolor1[1011]);
    BiasedRNG[376] = (LFSRcolor1[1336]&LFSRcolor1[1741]&LFSRcolor1[565]&LFSRcolor1[607]);
    BiasedRNG[377] = (LFSRcolor1[1331]&LFSRcolor1[778]&LFSRcolor1[861]&LFSRcolor1[1775]);
    BiasedRNG[378] = (LFSRcolor1[1549]&LFSRcolor1[1216]&LFSRcolor1[40]&LFSRcolor1[1075]);
    BiasedRNG[379] = (LFSRcolor1[1679]&LFSRcolor1[695]&LFSRcolor1[702]&LFSRcolor1[1254]);
    BiasedRNG[380] = (LFSRcolor1[308]&LFSRcolor1[944]&LFSRcolor1[1644]&LFSRcolor1[322]);
    BiasedRNG[381] = (LFSRcolor1[362]&LFSRcolor1[1510]&LFSRcolor1[1012]&LFSRcolor1[1663]);
    BiasedRNG[382] = (LFSRcolor1[853]&LFSRcolor1[984]&LFSRcolor1[82]&LFSRcolor1[831]);
    BiasedRNG[383] = (LFSRcolor1[349]&LFSRcolor1[1078]&LFSRcolor1[1779]&LFSRcolor1[457]);
    BiasedRNG[384] = (LFSRcolor1[1787]&LFSRcolor1[1055]&LFSRcolor1[1505]&LFSRcolor1[942]);
    BiasedRNG[385] = (LFSRcolor1[50]&LFSRcolor1[1547]&LFSRcolor1[35]&LFSRcolor1[1566]);
    BiasedRNG[386] = (LFSRcolor1[1366]&LFSRcolor1[93]&LFSRcolor1[623]&LFSRcolor1[48]);
    BiasedRNG[387] = (LFSRcolor1[1379]&LFSRcolor1[754]&LFSRcolor1[1626]&LFSRcolor1[85]);
    BiasedRNG[388] = (LFSRcolor1[748]&LFSRcolor1[84]&LFSRcolor1[880]&LFSRcolor1[637]);
    BiasedRNG[389] = (LFSRcolor1[1104]&LFSRcolor1[562]&LFSRcolor1[1458]&LFSRcolor1[866]);
    BiasedRNG[390] = (LFSRcolor1[1415]&LFSRcolor1[1213]&LFSRcolor1[673]&LFSRcolor1[120]);
    BiasedRNG[391] = (LFSRcolor1[474]&LFSRcolor1[918]&LFSRcolor1[177]&LFSRcolor1[1608]);
    BiasedRNG[392] = (LFSRcolor1[1281]&LFSRcolor1[144]&LFSRcolor1[192]&LFSRcolor1[714]);
    BiasedRNG[393] = (LFSRcolor1[446]&LFSRcolor1[1089]&LFSRcolor1[266]&LFSRcolor1[44]);
    BiasedRNG[394] = (LFSRcolor1[328]&LFSRcolor1[864]&LFSRcolor1[276]&LFSRcolor1[49]);
    BiasedRNG[395] = (LFSRcolor1[711]&LFSRcolor1[424]&LFSRcolor1[575]&LFSRcolor1[639]);
    BiasedRNG[396] = (LFSRcolor1[1085]&LFSRcolor1[206]&LFSRcolor1[255]&LFSRcolor1[146]);
    BiasedRNG[397] = (LFSRcolor1[1209]&LFSRcolor1[1226]&LFSRcolor1[518]&LFSRcolor1[482]);
    BiasedRNG[398] = (LFSRcolor1[1752]&LFSRcolor1[194]&LFSRcolor1[764]&LFSRcolor1[1116]);
    BiasedRNG[399] = (LFSRcolor1[1665]&LFSRcolor1[1092]&LFSRcolor1[1764]&LFSRcolor1[30]);
    BiasedRNG[400] = (LFSRcolor1[579]&LFSRcolor1[181]&LFSRcolor1[1769]&LFSRcolor1[1766]);
    BiasedRNG[401] = (LFSRcolor1[1199]&LFSRcolor1[382]&LFSRcolor1[423]&LFSRcolor1[1371]);
    BiasedRNG[402] = (LFSRcolor1[912]&LFSRcolor1[312]&LFSRcolor1[1627]&LFSRcolor1[1598]);
    BiasedRNG[403] = (LFSRcolor1[1246]&LFSRcolor1[1495]&LFSRcolor1[1520]&LFSRcolor1[381]);
    BiasedRNG[404] = (LFSRcolor1[1039]&LFSRcolor1[510]&LFSRcolor1[236]&LFSRcolor1[116]);
    BiasedRNG[405] = (LFSRcolor1[1087]&LFSRcolor1[1361]&LFSRcolor1[844]&LFSRcolor1[1417]);
    BiasedRNG[406] = (LFSRcolor1[1630]&LFSRcolor1[1407]&LFSRcolor1[1001]&LFSRcolor1[635]);
    BiasedRNG[407] = (LFSRcolor1[1168]&LFSRcolor1[468]&LFSRcolor1[820]&LFSRcolor1[746]);
    BiasedRNG[408] = (LFSRcolor1[491]&LFSRcolor1[884]&LFSRcolor1[515]&LFSRcolor1[1277]);
    BiasedRNG[409] = (LFSRcolor1[1703]&LFSRcolor1[272]&LFSRcolor1[1077]&LFSRcolor1[963]);
    BiasedRNG[410] = (LFSRcolor1[512]&LFSRcolor1[1090]&LFSRcolor1[1714]&LFSRcolor1[231]);
    BiasedRNG[411] = (LFSRcolor1[857]&LFSRcolor1[1478]&LFSRcolor1[788]&LFSRcolor1[1150]);
    BiasedRNG[412] = (LFSRcolor1[212]&LFSRcolor1[1066]&LFSRcolor1[151]&LFSRcolor1[502]);
    BiasedRNG[413] = (LFSRcolor1[118]&LFSRcolor1[1217]&LFSRcolor1[621]&LFSRcolor1[1049]);
    BiasedRNG[414] = (LFSRcolor1[402]&LFSRcolor1[1063]&LFSRcolor1[525]&LFSRcolor1[369]);
    BiasedRNG[415] = (LFSRcolor1[1113]&LFSRcolor1[1355]&LFSRcolor1[1071]&LFSRcolor1[867]);
    BiasedRNG[416] = (LFSRcolor1[530]&LFSRcolor1[540]&LFSRcolor1[338]&LFSRcolor1[1134]);
    BiasedRNG[417] = (LFSRcolor1[670]&LFSRcolor1[207]&LFSRcolor1[1786]&LFSRcolor1[932]);
    BiasedRNG[418] = (LFSRcolor1[1460]&LFSRcolor1[830]&LFSRcolor1[495]&LFSRcolor1[365]);
    BiasedRNG[419] = (LFSRcolor1[770]&LFSRcolor1[1676]&LFSRcolor1[958]&LFSRcolor1[771]);
    BiasedRNG[420] = (LFSRcolor1[801]&LFSRcolor1[839]&LFSRcolor1[955]&LFSRcolor1[1567]);
    BiasedRNG[421] = (LFSRcolor1[187]&LFSRcolor1[51]&LFSRcolor1[76]&LFSRcolor1[1748]);
    BiasedRNG[422] = (LFSRcolor1[202]&LFSRcolor1[1666]&LFSRcolor1[519]&LFSRcolor1[1632]);
    BiasedRNG[423] = (LFSRcolor1[1704]&LFSRcolor1[1659]&LFSRcolor1[521]&LFSRcolor1[211]);
    BiasedRNG[424] = (LFSRcolor1[1419]&LFSRcolor1[1413]&LFSRcolor1[1057]&LFSRcolor1[462]);
    BiasedRNG[425] = (LFSRcolor1[444]&LFSRcolor1[74]&LFSRcolor1[1365]&LFSRcolor1[376]);
    BiasedRNG[426] = (LFSRcolor1[281]&LFSRcolor1[1534]&LFSRcolor1[563]&LFSRcolor1[95]);
    BiasedRNG[427] = (LFSRcolor1[682]&LFSRcolor1[1781]&LFSRcolor1[69]&LFSRcolor1[1015]);
    BiasedRNG[428] = (LFSRcolor1[1573]&LFSRcolor1[1214]&LFSRcolor1[103]&LFSRcolor1[1203]);
    BiasedRNG[429] = (LFSRcolor1[150]&LFSRcolor1[334]&LFSRcolor1[1587]&LFSRcolor1[1487]);
    BiasedRNG[430] = (LFSRcolor1[43]&LFSRcolor1[1594]&LFSRcolor1[104]&LFSRcolor1[125]);
    BiasedRNG[431] = (LFSRcolor1[590]&LFSRcolor1[117]&LFSRcolor1[29]&LFSRcolor1[1197]);
    BiasedRNG[432] = (LFSRcolor1[1230]&LFSRcolor1[727]&LFSRcolor1[910]&LFSRcolor1[1022]);
    BiasedRNG[433] = (LFSRcolor1[1572]&LFSRcolor1[190]&LFSRcolor1[9]&LFSRcolor1[1701]);
    BiasedRNG[434] = (LFSRcolor1[1515]&LFSRcolor1[854]&LFSRcolor1[1207]&LFSRcolor1[1291]);
    BiasedRNG[435] = (LFSRcolor1[875]&LFSRcolor1[648]&LFSRcolor1[1638]&LFSRcolor1[1588]);
    BiasedRNG[436] = (LFSRcolor1[1028]&LFSRcolor1[1144]&LFSRcolor1[1525]&LFSRcolor1[245]);
    BiasedRNG[437] = (LFSRcolor1[1193]&LFSRcolor1[39]&LFSRcolor1[705]&LFSRcolor1[367]);
    BiasedRNG[438] = (LFSRcolor1[713]&LFSRcolor1[306]&LFSRcolor1[1339]&LFSRcolor1[1211]);
    BiasedRNG[439] = (LFSRcolor1[529]&LFSRcolor1[816]&LFSRcolor1[1]&LFSRcolor1[732]);
    BiasedRNG[440] = (LFSRcolor1[1215]&LFSRcolor1[252]&LFSRcolor1[258]&LFSRcolor1[989]);
    BiasedRNG[441] = (LFSRcolor1[645]&LFSRcolor1[723]&LFSRcolor1[1667]&LFSRcolor1[160]);
    BiasedRNG[442] = (LFSRcolor1[233]&LFSRcolor1[20]&LFSRcolor1[1681]&LFSRcolor1[66]);
    BiasedRNG[443] = (LFSRcolor1[1155]&LFSRcolor1[1114]&LFSRcolor1[1738]&LFSRcolor1[1335]);
    BiasedRNG[444] = (LFSRcolor1[1356]&LFSRcolor1[1634]&LFSRcolor1[1182]&LFSRcolor1[847]);
    BiasedRNG[445] = (LFSRcolor1[153]&LFSRcolor1[1754]&LFSRcolor1[1271]&LFSRcolor1[893]);
    BiasedRNG[446] = (LFSRcolor1[1740]&LFSRcolor1[1772]&LFSRcolor1[269]&LFSRcolor1[925]);
    BiasedRNG[447] = (LFSRcolor1[1660]&LFSRcolor1[1183]&LFSRcolor1[416]&LFSRcolor1[1304]);
    BiasedRNG[448] = (LFSRcolor1[124]&LFSRcolor1[1372]&LFSRcolor1[1530]&LFSRcolor1[136]);
    BiasedRNG[449] = (LFSRcolor1[828]&LFSRcolor1[1387]&LFSRcolor1[1545]&LFSRcolor1[249]);
    BiasedRNG[450] = (LFSRcolor1[55]&LFSRcolor1[589]&LFSRcolor1[1316]&LFSRcolor1[166]);
    BiasedRNG[451] = (LFSRcolor1[1410]&LFSRcolor1[1421]&LFSRcolor1[405]&LFSRcolor1[511]);
    BiasedRNG[452] = (LFSRcolor1[819]&LFSRcolor1[439]&LFSRcolor1[930]&LFSRcolor1[449]);
    BiasedRNG[453] = (LFSRcolor1[1003]&LFSRcolor1[243]&LFSRcolor1[1096]&LFSRcolor1[1208]);
    BiasedRNG[454] = (LFSRcolor1[235]&LFSRcolor1[288]&LFSRcolor1[1184]&LFSRcolor1[414]);
    BiasedRNG[455] = (LFSRcolor1[1034]&LFSRcolor1[401]&LFSRcolor1[1680]&LFSRcolor1[1500]);
    BiasedRNG[456] = (LFSRcolor1[241]&LFSRcolor1[224]&LFSRcolor1[975]&LFSRcolor1[513]);
    BiasedRNG[457] = (LFSRcolor1[1556]&LFSRcolor1[546]&LFSRcolor1[709]&LFSRcolor1[1238]);
    BiasedRNG[458] = (LFSRcolor1[542]&LFSRcolor1[216]&LFSRcolor1[901]&LFSRcolor1[1348]);
    BiasedRNG[459] = (LFSRcolor1[13]&LFSRcolor1[392]&LFSRcolor1[881]&LFSRcolor1[1771]);
    BiasedRNG[460] = (LFSRcolor1[419]&LFSRcolor1[940]&LFSRcolor1[991]&LFSRcolor1[980]);
    BiasedRNG[461] = (LFSRcolor1[1229]&LFSRcolor1[427]&LFSRcolor1[1502]&LFSRcolor1[538]);
    BiasedRNG[462] = (LFSRcolor1[710]&LFSRcolor1[100]&LFSRcolor1[262]&LFSRcolor1[1029]);
    BiasedRNG[463] = (LFSRcolor1[580]&LFSRcolor1[1314]&LFSRcolor1[1353]&LFSRcolor1[496]);
    BiasedRNG[464] = (LFSRcolor1[1248]&LFSRcolor1[412]&LFSRcolor1[1330]&LFSRcolor1[1431]);
    BiasedRNG[465] = (LFSRcolor1[152]&LFSRcolor1[1364]&LFSRcolor1[331]&LFSRcolor1[1582]);
    BiasedRNG[466] = (LFSRcolor1[641]&LFSRcolor1[161]&LFSRcolor1[1453]&LFSRcolor1[1286]);
    BiasedRNG[467] = (LFSRcolor1[897]&LFSRcolor1[220]&LFSRcolor1[1045]&LFSRcolor1[1363]);
    BiasedRNG[468] = (LFSRcolor1[887]&LFSRcolor1[1338]&LFSRcolor1[1367]&LFSRcolor1[397]);
    BiasedRNG[469] = (LFSRcolor1[572]&LFSRcolor1[1603]&LFSRcolor1[230]&LFSRcolor1[1411]);
    BiasedRNG[470] = (LFSRcolor1[986]&LFSRcolor1[1447]&LFSRcolor1[773]&LFSRcolor1[284]);
    BiasedRNG[471] = (LFSRcolor1[1514]&LFSRcolor1[1084]&LFSRcolor1[62]&LFSRcolor1[1337]);
    BiasedRNG[472] = (LFSRcolor1[1670]&LFSRcolor1[1537]&LFSRcolor1[517]&LFSRcolor1[1162]);
    BiasedRNG[473] = (LFSRcolor1[268]&LFSRcolor1[489]&LFSRcolor1[1597]&LFSRcolor1[352]);
    BiasedRNG[474] = (LFSRcolor1[1050]&LFSRcolor1[1299]&LFSRcolor1[990]&LFSRcolor1[1153]);
    BiasedRNG[475] = (LFSRcolor1[1488]&LFSRcolor1[1370]&LFSRcolor1[805]&LFSRcolor1[279]);
    BiasedRNG[476] = (LFSRcolor1[961]&LFSRcolor1[657]&LFSRcolor1[1541]&LFSRcolor1[1347]);
    BiasedRNG[477] = (LFSRcolor1[1512]&LFSRcolor1[425]&LFSRcolor1[781]&LFSRcolor1[612]);
    BiasedRNG[478] = (LFSRcolor1[1076]&LFSRcolor1[1466]&LFSRcolor1[1279]&LFSRcolor1[840]);
    BiasedRNG[479] = (LFSRcolor1[625]&LFSRcolor1[1164]&LFSRcolor1[552]&LFSRcolor1[1523]);
    BiasedRNG[480] = (LFSRcolor1[1376]&LFSRcolor1[1690]&LFSRcolor1[598]&LFSRcolor1[463]);
    BiasedRNG[481] = (LFSRcolor1[154]&LFSRcolor1[1497]&LFSRcolor1[1222]&LFSRcolor1[1482]);
    BiasedRNG[482] = (LFSRcolor1[1589]&LFSRcolor1[1033]&LFSRcolor1[1079]&LFSRcolor1[178]);
    BiasedRNG[483] = (LFSRcolor1[1619]&LFSRcolor1[1474]&LFSRcolor1[939]&LFSRcolor1[1359]);
    BiasedRNG[484] = (LFSRcolor1[1321]&LFSRcolor1[1485]&LFSRcolor1[1097]&LFSRcolor1[295]);
    BiasedRNG[485] = (LFSRcolor1[56]&LFSRcolor1[868]&LFSRcolor1[587]&LFSRcolor1[1380]);
    BiasedRNG[486] = (LFSRcolor1[1306]&LFSRcolor1[1436]&LFSRcolor1[922]&LFSRcolor1[228]);
    BiasedRNG[487] = (LFSRcolor1[1307]&LFSRcolor1[949]&LFSRcolor1[556]&LFSRcolor1[927]);
    BiasedRNG[488] = (LFSRcolor1[335]&LFSRcolor1[445]&LFSRcolor1[1602]&LFSRcolor1[933]);
    BiasedRNG[489] = (LFSRcolor1[768]&LFSRcolor1[655]&LFSRcolor1[1053]&LFSRcolor1[1219]);
    BiasedRNG[490] = (LFSRcolor1[620]&LFSRcolor1[1151]&LFSRcolor1[804]&LFSRcolor1[1593]);
    BiasedRNG[491] = (LFSRcolor1[1726]&LFSRcolor1[1565]&LFSRcolor1[776]&LFSRcolor1[950]);
    BiasedRNG[492] = (LFSRcolor1[379]&LFSRcolor1[1528]&LFSRcolor1[685]&LFSRcolor1[604]);
    BiasedRNG[493] = (LFSRcolor1[1020]&LFSRcolor1[1302]&LFSRcolor1[1391]&LFSRcolor1[25]);
    BiasedRNG[494] = (LFSRcolor1[430]&LFSRcolor1[553]&LFSRcolor1[81]&LFSRcolor1[1461]);
    BiasedRNG[495] = (LFSRcolor1[600]&LFSRcolor1[21]&LFSRcolor1[800]&LFSRcolor1[201]);
    BiasedRNG[496] = (LFSRcolor1[825]&LFSRcolor1[905]&LFSRcolor1[1122]&LFSRcolor1[157]);
    BiasedRNG[497] = (LFSRcolor1[1527]&LFSRcolor1[549]&LFSRcolor1[1728]&LFSRcolor1[756]);
    BiasedRNG[498] = (LFSRcolor1[320]&LFSRcolor1[387]&LFSRcolor1[1128]&LFSRcolor1[977]);
    BiasedRNG[499] = (LFSRcolor1[438]&LFSRcolor1[1613]&LFSRcolor1[122]&LFSRcolor1[1285]);
    BiasedRNG[500] = (LFSRcolor1[1098]&LFSRcolor1[485]&LFSRcolor1[1499]&LFSRcolor1[707]);
    BiasedRNG[501] = (LFSRcolor1[339]&LFSRcolor1[1253]&LFSRcolor1[715]&LFSRcolor1[176]);
    BiasedRNG[502] = (LFSRcolor1[1133]&LFSRcolor1[53]&LFSRcolor1[1539]&LFSRcolor1[1434]);
    BiasedRNG[503] = (LFSRcolor1[80]&LFSRcolor1[456]&LFSRcolor1[631]&LFSRcolor1[226]);
    BiasedRNG[504] = (LFSRcolor1[143]&LFSRcolor1[1121]&LFSRcolor1[1068]&LFSRcolor1[656]);
    BiasedRNG[505] = (LFSRcolor1[718]&LFSRcolor1[740]&LFSRcolor1[469]&LFSRcolor1[1037]);
    BiasedRNG[506] = (LFSRcolor1[987]&LFSRcolor1[615]&LFSRcolor1[1270]&LFSRcolor1[838]);
    BiasedRNG[507] = (LFSRcolor1[1480]&LFSRcolor1[1324]&LFSRcolor1[10]&LFSRcolor1[999]);
    BiasedRNG[508] = (LFSRcolor1[668]&LFSRcolor1[640]&LFSRcolor1[751]&LFSRcolor1[1352]);
    BiasedRNG[509] = (LFSRcolor1[163]&LFSRcolor1[629]&LFSRcolor1[1019]&LFSRcolor1[1519]);
    BiasedRNG[510] = (LFSRcolor1[162]&LFSRcolor1[1191]&LFSRcolor1[330]&LFSRcolor1[642]);
    BiasedRNG[511] = (LFSRcolor1[135]&LFSRcolor1[1268]&LFSRcolor1[1554]&LFSRcolor1[646]);
    BiasedRNG[512] = (LFSRcolor1[946]&LFSRcolor1[675]&LFSRcolor1[1083]&LFSRcolor1[179]);
    BiasedRNG[513] = (LFSRcolor1[1170]&LFSRcolor1[1210]&LFSRcolor1[1529]&LFSRcolor1[889]);
    BiasedRNG[514] = (LFSRcolor1[951]&LFSRcolor1[46]&LFSRcolor1[12]&LFSRcolor1[142]);
    BiasedRNG[515] = (LFSRcolor1[829]&LFSRcolor1[1386]&LFSRcolor1[1318]&LFSRcolor1[1303]);
    BiasedRNG[516] = (LFSRcolor1[564]&LFSRcolor1[597]&LFSRcolor1[1496]&LFSRcolor1[681]);
    BiasedRNG[517] = (LFSRcolor1[1662]&LFSRcolor1[282]&LFSRcolor1[581]&LFSRcolor1[846]);
    BiasedRNG[518] = (LFSRcolor1[1009]&LFSRcolor1[863]&LFSRcolor1[983]&LFSRcolor1[1763]);
    BiasedRNG[519] = (LFSRcolor1[683]&LFSRcolor1[584]&LFSRcolor1[652]&LFSRcolor1[1024]);
    BiasedRNG[520] = (LFSRcolor1[622]&LFSRcolor1[1777]&LFSRcolor1[1131]&LFSRcolor1[1036]);
    BiasedRNG[521] = (LFSRcolor1[222]&LFSRcolor1[1111]&LFSRcolor1[1156]&LFSRcolor1[716]);
    BiasedRNG[522] = (LFSRcolor1[1654]&LFSRcolor1[73]&LFSRcolor1[341]&LFSRcolor1[1575]);
    BiasedRNG[523] = (LFSRcolor1[1308]&LFSRcolor1[630]&LFSRcolor1[1760]&LFSRcolor1[848]);
    BiasedRNG[524] = (LFSRcolor1[1402]&LFSRcolor1[1007]&LFSRcolor1[1677]&LFSRcolor1[885]);
    BiasedRNG[525] = (LFSRcolor1[221]&LFSRcolor1[767]&LFSRcolor1[475]&LFSRcolor1[70]);
    BiasedRNG[526] = (LFSRcolor1[687]&LFSRcolor1[199]&LFSRcolor1[147]&LFSRcolor1[1295]);
    BiasedRNG[527] = (LFSRcolor1[354]&LFSRcolor1[1175]&LFSRcolor1[1106]&LFSRcolor1[1396]);
    BiasedRNG[528] = (LFSRcolor1[728]&LFSRcolor1[815]&LFSRcolor1[441]&LFSRcolor1[859]);
    BiasedRNG[529] = (LFSRcolor1[760]&LFSRcolor1[88]&LFSRcolor1[210]&LFSRcolor1[1655]);
    BiasedRNG[530] = (LFSRcolor1[375]&LFSRcolor1[1581]&LFSRcolor1[1576]&LFSRcolor1[315]);
    BiasedRNG[531] = (LFSRcolor1[1621]&LFSRcolor1[1300]&LFSRcolor1[1255]&LFSRcolor1[836]);
    BiasedRNG[532] = (LFSRcolor1[1296]&LFSRcolor1[669]&LFSRcolor1[193]&LFSRcolor1[1491]);
    BiasedRNG[533] = (LFSRcolor1[1005]&LFSRcolor1[1334]&LFSRcolor1[248]&LFSRcolor1[1389]);
    BiasedRNG[534] = (LFSRcolor1[1166]&LFSRcolor1[601]&LFSRcolor1[1579]&LFSRcolor1[1123]);
    BiasedRNG[535] = (LFSRcolor1[1412]&LFSRcolor1[1399]&LFSRcolor1[593]&LFSRcolor1[1179]);
    BiasedRNG[536] = (LFSRcolor1[1454]&LFSRcolor1[664]&LFSRcolor1[137]&LFSRcolor1[428]);
    BiasedRNG[537] = (LFSRcolor1[763]&LFSRcolor1[127]&LFSRcolor1[1590]&LFSRcolor1[394]);
    BiasedRNG[538] = (LFSRcolor1[558]&LFSRcolor1[1236]&LFSRcolor1[1205]&LFSRcolor1[1471]);
    BiasedRNG[539] = (LFSRcolor1[599]&LFSRcolor1[1192]&LFSRcolor1[1000]&LFSRcolor1[1457]);
    BiasedRNG[540] = (LFSRcolor1[824]&LFSRcolor1[285]&LFSRcolor1[821]&LFSRcolor1[1287]);
    BiasedRNG[541] = (LFSRcolor1[1158]&LFSRcolor1[1301]&LFSRcolor1[1173]&LFSRcolor1[121]);
    BiasedRNG[542] = (LFSRcolor1[865]&LFSRcolor1[1792]&LFSRcolor1[1073]&LFSRcolor1[544]);
    BiasedRNG[543] = (LFSRcolor1[1778]&LFSRcolor1[724]&LFSRcolor1[1697]&LFSRcolor1[38]);
    BiasedRNG[544] = (LFSRcolor1[5]&LFSRcolor1[1108]&LFSRcolor1[1509]&LFSRcolor1[309]);
    BiasedRNG[545] = (LFSRcolor1[722]&LFSRcolor1[891]&LFSRcolor1[36]&LFSRcolor1[509]);
    BiasedRNG[546] = (LFSRcolor1[1294]&LFSRcolor1[168]&LFSRcolor1[167]&LFSRcolor1[743]);
    BiasedRNG[547] = (LFSRcolor1[595]&LFSRcolor1[411]&LFSRcolor1[793]&LFSRcolor1[275]);
    BiasedRNG[548] = (LFSRcolor1[1218]&LFSRcolor1[114]&LFSRcolor1[296]&LFSRcolor1[873]);
    BiasedRNG[549] = (LFSRcolor1[1604]&LFSRcolor1[1169]&LFSRcolor1[129]&LFSRcolor1[377]);
    BiasedRNG[550] = (LFSRcolor1[102]&LFSRcolor1[311]&LFSRcolor1[332]&LFSRcolor1[934]);
    BiasedRNG[551] = (LFSRcolor1[197]&LFSRcolor1[1671]&LFSRcolor1[407]&LFSRcolor1[1742]);
    BiasedRNG[552] = (LFSRcolor1[23]&LFSRcolor1[1583]&LFSRcolor1[1375]&LFSRcolor1[303]);
    BiasedRNG[553] = (LFSRcolor1[246]&LFSRcolor1[935]&LFSRcolor1[684]&LFSRcolor1[1322]);
    BiasedRNG[554] = (LFSRcolor1[779]&LFSRcolor1[921]&LFSRcolor1[270]&LFSRcolor1[1472]);
    BiasedRNG[555] = (LFSRcolor1[1140]&LFSRcolor1[752]&LFSRcolor1[1761]&LFSRcolor1[1641]);
    BiasedRNG[556] = (LFSRcolor1[1720]&LFSRcolor1[592]&LFSRcolor1[171]&LFSRcolor1[223]);
    BiasedRNG[557] = (LFSRcolor1[810]&LFSRcolor1[472]&LFSRcolor1[1791]&LFSRcolor1[1160]);
    BiasedRNG[558] = (LFSRcolor1[60]&LFSRcolor1[52]&LFSRcolor1[1459]&LFSRcolor1[1377]);
    BiasedRNG[559] = (LFSRcolor1[1427]&LFSRcolor1[550]&LFSRcolor1[355]&LFSRcolor1[1708]);
    BiasedRNG[560] = (LFSRcolor1[1264]&LFSRcolor1[1780]&LFSRcolor1[628]&LFSRcolor1[920]);
    BiasedRNG[561] = (LFSRcolor1[1251]&LFSRcolor1[719]&LFSRcolor1[1517]&LFSRcolor1[149]);
    BiasedRNG[562] = (LFSRcolor1[218]&LFSRcolor1[33]&LFSRcolor1[342]&LFSRcolor1[766]);
    BiasedRNG[563] = (LFSRcolor1[516]&LFSRcolor1[1451]&LFSRcolor1[280]&LFSRcolor1[1091]);
    BiasedRNG[564] = (LFSRcolor1[1163]&LFSRcolor1[158]&LFSRcolor1[172]&LFSRcolor1[654]);
    BiasedRNG[565] = (LFSRcolor1[1358]&LFSRcolor1[734]&LFSRcolor1[1135]&LFSRcolor1[1601]);
    BiasedRNG[566] = (LFSRcolor1[551]&LFSRcolor1[965]&LFSRcolor1[643]&LFSRcolor1[488]);
    BiasedRNG[567] = (LFSRcolor1[110]&LFSRcolor1[440]&LFSRcolor1[979]&LFSRcolor1[1719]);
    BiasedRNG[568] = (LFSRcolor1[398]&LFSRcolor1[1606]&LFSRcolor1[466]&LFSRcolor1[1196]);
    BiasedRNG[569] = (LFSRcolor1[555]&LFSRcolor1[943]&LFSRcolor1[931]&LFSRcolor1[1319]);
    BiasedRNG[570] = (LFSRcolor1[1790]&LFSRcolor1[318]&LFSRcolor1[982]&LFSRcolor1[1388]);
    BiasedRNG[571] = (LFSRcolor1[960]&LFSRcolor1[1137]&LFSRcolor1[454]&LFSRcolor1[164]);
    BiasedRNG[572] = (LFSRcolor1[1617]&LFSRcolor1[1225]&LFSRcolor1[271]&LFSRcolor1[811]);
    BiasedRNG[573] = (LFSRcolor1[267]&LFSRcolor1[31]&LFSRcolor1[1687]&LFSRcolor1[699]);
    BiasedRNG[574] = (LFSRcolor1[28]&LFSRcolor1[1538]&LFSRcolor1[514]&LFSRcolor1[945]);
    BiasedRNG[575] = (LFSRcolor1[560]&LFSRcolor1[333]&LFSRcolor1[735]&LFSRcolor1[385]);
    BiasedRNG[576] = (LFSRcolor1[786]&LFSRcolor1[1139]&LFSRcolor1[1062]&LFSRcolor1[822]);
    BiasedRNG[577] = (LFSRcolor1[1455]&LFSRcolor1[967]&LFSRcolor1[1469]&LFSRcolor1[557]);
    BiasedRNG[578] = (LFSRcolor1[471]&LFSRcolor1[1395]&LFSRcolor1[16]&LFSRcolor1[105]);
    BiasedRNG[579] = (LFSRcolor1[119]&LFSRcolor1[250]&LFSRcolor1[1755]&LFSRcolor1[213]);
    BiasedRNG[580] = (LFSRcolor1[345]&LFSRcolor1[1624]&LFSRcolor1[290]&LFSRcolor1[1272]);
    BiasedRNG[581] = (LFSRcolor1[959]&LFSRcolor1[1320]&LFSRcolor1[1759]&LFSRcolor1[919]);
    BiasedRNG[582] = (LFSRcolor1[1645]&LFSRcolor1[283]&LFSRcolor1[1653]&LFSRcolor1[1346]);
    BiasedRNG[583] = (LFSRcolor1[1044]&LFSRcolor1[483]&LFSRcolor1[217]&LFSRcolor1[742]);
    BiasedRNG[584] = (LFSRcolor1[1712]&LFSRcolor1[1563]&LFSRcolor1[1309]&LFSRcolor1[1784]);
    BiasedRNG[585] = (LFSRcolor1[1646]&LFSRcolor1[494]&LFSRcolor1[1650]&LFSRcolor1[1729]);
    BiasedRNG[586] = (LFSRcolor1[1578]&LFSRcolor1[1470]&LFSRcolor1[1016]&LFSRcolor1[406]);
    BiasedRNG[587] = (LFSRcolor1[1692]&LFSRcolor1[314]&LFSRcolor1[350]&LFSRcolor1[1204]);
    BiasedRNG[588] = (LFSRcolor1[537]&LFSRcolor1[782]&LFSRcolor1[941]&LFSRcolor1[87]);
    BiasedRNG[589] = (LFSRcolor1[479]&LFSRcolor1[898]&LFSRcolor1[1546]&LFSRcolor1[1278]);
    BiasedRNG[590] = (LFSRcolor1[1475]&LFSRcolor1[310]&LFSRcolor1[329]&LFSRcolor1[1682]);
    BiasedRNG[591] = (LFSRcolor1[1623]&LFSRcolor1[594]&LFSRcolor1[850]&LFSRcolor1[1069]);
    BiasedRNG[592] = (LFSRcolor1[1477]&LFSRcolor1[523]&LFSRcolor1[305]&LFSRcolor1[1532]);
    BiasedRNG[593] = (LFSRcolor1[259]&LFSRcolor1[1718]&LFSRcolor1[1664]&LFSRcolor1[759]);
    BiasedRNG[594] = (LFSRcolor1[477]&LFSRcolor1[79]&LFSRcolor1[1048]&LFSRcolor1[611]);
    BiasedRNG[595] = (LFSRcolor1[1397]&LFSRcolor1[548]&LFSRcolor1[818]&LFSRcolor1[1332]);
    BiasedRNG[596] = (LFSRcolor1[1040]&LFSRcolor1[636]&LFSRcolor1[978]&LFSRcolor1[534]);
    BiasedRNG[597] = (LFSRcolor1[524]&LFSRcolor1[988]&LFSRcolor1[1224]&LFSRcolor1[107]);
    BiasedRNG[598] = (LFSRcolor1[1305]&LFSRcolor1[1064]&LFSRcolor1[173]&LFSRcolor1[835]);
    BiasedRNG[599] = (LFSRcolor1[148]&LFSRcolor1[364]&LFSRcolor1[753]&LFSRcolor1[324]);
    BiasedRNG[600] = (LFSRcolor1[852]&LFSRcolor1[1774]&LFSRcolor1[1021]&LFSRcolor1[966]);
    BiasedRNG[601] = (LFSRcolor1[956]&LFSRcolor1[92]&LFSRcolor1[749]&LFSRcolor1[1187]);
    BiasedRNG[602] = (LFSRcolor1[1486]&LFSRcolor1[1711]&LFSRcolor1[738]&LFSRcolor1[1568]);
    BiasedRNG[603] = (LFSRcolor1[45]&LFSRcolor1[435]&LFSRcolor1[1584]&LFSRcolor1[113]);
    BiasedRNG[604] = (LFSRcolor1[1297]&LFSRcolor1[263]&LFSRcolor1[464]&LFSRcolor1[1054]);
    BiasedRNG[605] = (LFSRcolor1[384]&LFSRcolor1[582]&LFSRcolor1[337]&LFSRcolor1[1058]);
    BiasedRNG[606] = (LFSRcolor1[344]&LFSRcolor1[134]&LFSRcolor1[273]&LFSRcolor1[1250]);
    BiasedRNG[607] = (LFSRcolor1[1107]&LFSRcolor1[1283]&LFSRcolor1[1284]&LFSRcolor1[1027]);
    BiasedRNG[608] = (LFSRcolor1[1511]&LFSRcolor1[796]&LFSRcolor1[361]&LFSRcolor1[1260]);
    BiasedRNG[609] = (LFSRcolor1[378]&LFSRcolor1[340]&LFSRcolor1[126]&LFSRcolor1[573]);
    BiasedRNG[610] = (LFSRcolor1[535]&LFSRcolor1[928]&LFSRcolor1[301]&LFSRcolor1[1178]);
    BiasedRNG[611] = (LFSRcolor1[260]&LFSRcolor1[1327]&LFSRcolor1[174]&LFSRcolor1[1032]);
    BiasedRNG[612] = (LFSRcolor1[1080]&LFSRcolor1[1648]&LFSRcolor1[877]&LFSRcolor1[870]);
    BiasedRNG[613] = (LFSRcolor1[588]&LFSRcolor1[467]&LFSRcolor1[90]&LFSRcolor1[1018]);
    BiasedRNG[614] = (LFSRcolor1[453]&LFSRcolor1[1072]&LFSRcolor1[1734]&LFSRcolor1[976]);
    BiasedRNG[615] = (LFSRcolor1[1550]&LFSRcolor1[896]&LFSRcolor1[739]&LFSRcolor1[251]);
    BiasedRNG[616] = (LFSRcolor1[373]&LFSRcolor1[1357]&LFSRcolor1[319]&LFSRcolor1[1167]);
    BiasedRNG[617] = (LFSRcolor1[799]&LFSRcolor1[1592]&LFSRcolor1[14]&LFSRcolor1[1065]);
    BiasedRNG[618] = (LFSRcolor1[200]&LFSRcolor1[1577]&LFSRcolor1[240]&LFSRcolor1[478]);
    BiasedRNG[619] = (LFSRcolor1[1117]&LFSRcolor1[909]&LFSRcolor1[1770]&LFSRcolor1[175]);
    BiasedRNG[620] = (LFSRcolor1[1329]&LFSRcolor1[571]&LFSRcolor1[215]&LFSRcolor1[1610]);
    BiasedRNG[621] = (LFSRcolor1[452]&LFSRcolor1[1756]&LFSRcolor1[480]&LFSRcolor1[647]);
    BiasedRNG[622] = (LFSRcolor1[947]&LFSRcolor1[94]&LFSRcolor1[1484]&LFSRcolor1[1783]);
    BiasedRNG[623] = (LFSRcolor1[343]&LFSRcolor1[203]&LFSRcolor1[254]&LFSRcolor1[520]);
    BiasedRNG[624] = (LFSRcolor1[790]&LFSRcolor1[1383]&LFSRcolor1[888]&LFSRcolor1[1416]);
    BiasedRNG[625] = (LFSRcolor1[809]&LFSRcolor1[522]&LFSRcolor1[814]&LFSRcolor1[422]);
    BiasedRNG[626] = (LFSRcolor1[481]&LFSRcolor1[1014]&LFSRcolor1[895]&LFSRcolor1[677]);
    BiasedRNG[627] = (LFSRcolor1[614]&LFSRcolor1[109]&LFSRcolor1[1747]&LFSRcolor1[145]);
    BiasedRNG[628] = (LFSRcolor1[1317]&LFSRcolor1[372]&LFSRcolor1[1658]&LFSRcolor1[1468]);
    BiasedRNG[629] = (LFSRcolor1[1393]&LFSRcolor1[317]&LFSRcolor1[487]&LFSRcolor1[1234]);
    BiasedRNG[630] = (LFSRcolor1[690]&LFSRcolor1[325]&LFSRcolor1[493]&LFSRcolor1[1675]);
    BiasedRNG[631] = (LFSRcolor1[1154]&LFSRcolor1[851]&LFSRcolor1[307]&LFSRcolor1[1004]);
    BiasedRNG[632] = (LFSRcolor1[1611]&LFSRcolor1[61]&LFSRcolor1[1157]&LFSRcolor1[1698]);
    BiasedRNG[633] = (LFSRcolor1[1762]&LFSRcolor1[1441]&LFSRcolor1[59]&LFSRcolor1[1600]);
    BiasedRNG[634] = (LFSRcolor1[1120]&LFSRcolor1[106]&LFSRcolor1[626]&LFSRcolor1[1596]);
    BiasedRNG[635] = (LFSRcolor1[196]&LFSRcolor1[1267]&LFSRcolor1[1310]&LFSRcolor1[239]);
    BiasedRNG[636] = (LFSRcolor1[182]&LFSRcolor1[1298]&LFSRcolor1[1551]&LFSRcolor1[1115]);
    BiasedRNG[637] = (LFSRcolor1[541]&LFSRcolor1[858]&LFSRcolor1[1437]&LFSRcolor1[973]);
    BiasedRNG[638] = (LFSRcolor1[507]&LFSRcolor1[294]&LFSRcolor1[389]&LFSRcolor1[929]);
    UnbiasedRNG[271] = LFSRcolor1[1521];
    UnbiasedRNG[272] = LFSRcolor1[130];
    UnbiasedRNG[273] = LFSRcolor1[1147];
    UnbiasedRNG[274] = LFSRcolor1[1244];
    UnbiasedRNG[275] = LFSRcolor1[610];
    UnbiasedRNG[276] = LFSRcolor1[744];
    UnbiasedRNG[277] = LFSRcolor1[302];
    UnbiasedRNG[278] = LFSRcolor1[609];
    UnbiasedRNG[279] = LFSRcolor1[817];
    UnbiasedRNG[280] = LFSRcolor1[692];
    UnbiasedRNG[281] = LFSRcolor1[1026];
    UnbiasedRNG[282] = LFSRcolor1[1351];
    UnbiasedRNG[283] = LFSRcolor1[1233];
    UnbiasedRNG[284] = LFSRcolor1[1531];
    UnbiasedRNG[285] = LFSRcolor1[729];
    UnbiasedRNG[286] = LFSRcolor1[195];
    UnbiasedRNG[287] = LFSRcolor1[6];
    UnbiasedRNG[288] = LFSRcolor1[506];
    UnbiasedRNG[289] = LFSRcolor1[841];
    UnbiasedRNG[290] = LFSRcolor1[807];
    UnbiasedRNG[291] = LFSRcolor1[1390];
    UnbiasedRNG[292] = LFSRcolor1[971];
    UnbiasedRNG[293] = LFSRcolor1[169];
    UnbiasedRNG[294] = LFSRcolor1[7];
    UnbiasedRNG[295] = LFSRcolor1[1432];
    UnbiasedRNG[296] = LFSRcolor1[962];
    UnbiasedRNG[297] = LFSRcolor1[1757];
    UnbiasedRNG[298] = LFSRcolor1[712];
    UnbiasedRNG[299] = LFSRcolor1[1142];
    UnbiasedRNG[300] = LFSRcolor1[1730];
    UnbiasedRNG[301] = LFSRcolor1[391];
    UnbiasedRNG[302] = LFSRcolor1[1788];
    UnbiasedRNG[303] = LFSRcolor1[1750];
    UnbiasedRNG[304] = LFSRcolor1[356];
    UnbiasedRNG[305] = LFSRcolor1[1694];
    UnbiasedRNG[306] = LFSRcolor1[1765];
    UnbiasedRNG[307] = LFSRcolor1[497];
    UnbiasedRNG[308] = LFSRcolor1[15];
    UnbiasedRNG[309] = LFSRcolor1[591];
    UnbiasedRNG[310] = LFSRcolor1[797];
    UnbiasedRNG[311] = LFSRcolor1[902];
    UnbiasedRNG[312] = LFSRcolor1[1536];
    UnbiasedRNG[313] = LFSRcolor1[761];
    UnbiasedRNG[314] = LFSRcolor1[914];
    UnbiasedRNG[315] = LFSRcolor1[787];
    UnbiasedRNG[316] = LFSRcolor1[1707];
    UnbiasedRNG[317] = LFSRcolor1[1282];
    UnbiasedRNG[318] = LFSRcolor1[1614];
    UnbiasedRNG[319] = LFSRcolor1[326];
    UnbiasedRNG[320] = LFSRcolor1[1631];
    UnbiasedRNG[321] = LFSRcolor1[1093];
    UnbiasedRNG[322] = LFSRcolor1[970];
    UnbiasedRNG[323] = LFSRcolor1[911];
    UnbiasedRNG[324] = LFSRcolor1[1564];
    UnbiasedRNG[325] = LFSRcolor1[1288];
    UnbiasedRNG[326] = LFSRcolor1[189];
    UnbiasedRNG[327] = LFSRcolor1[1744];
    UnbiasedRNG[328] = LFSRcolor1[1070];
    UnbiasedRNG[329] = LFSRcolor1[1463];
    UnbiasedRNG[330] = LFSRcolor1[1423];
    UnbiasedRNG[331] = LFSRcolor1[1693];
    UnbiasedRNG[332] = LFSRcolor1[679];
    UnbiasedRNG[333] = LFSRcolor1[661];
    UnbiasedRNG[334] = LFSRcolor1[434];
    UnbiasedRNG[335] = LFSRcolor1[1713];
    UnbiasedRNG[336] = LFSRcolor1[1100];
    UnbiasedRNG[337] = LFSRcolor1[191];
    UnbiasedRNG[338] = LFSRcolor1[443];
    UnbiasedRNG[339] = LFSRcolor1[936];
    UnbiasedRNG[340] = LFSRcolor1[792];
    UnbiasedRNG[341] = LFSRcolor1[1340];
    UnbiasedRNG[342] = LFSRcolor1[1678];
    UnbiasedRNG[343] = LFSRcolor1[755];
    UnbiasedRNG[344] = LFSRcolor1[1629];
    UnbiasedRNG[345] = LFSRcolor1[903];
    UnbiasedRNG[346] = LFSRcolor1[386];
    UnbiasedRNG[347] = LFSRcolor1[1420];
    UnbiasedRNG[348] = LFSRcolor1[27];
    UnbiasedRNG[349] = LFSRcolor1[1403];
    UnbiasedRNG[350] = LFSRcolor1[624];
    UnbiasedRNG[351] = LFSRcolor1[374];
    UnbiasedRNG[352] = LFSRcolor1[54];
    UnbiasedRNG[353] = LFSRcolor1[1186];
    UnbiasedRNG[354] = LFSRcolor1[1622];
    UnbiasedRNG[355] = LFSRcolor1[1398];
    UnbiasedRNG[356] = LFSRcolor1[291];
    UnbiasedRNG[357] = LFSRcolor1[1148];
    UnbiasedRNG[358] = LFSRcolor1[316];
    UnbiasedRNG[359] = LFSRcolor1[128];
    UnbiasedRNG[360] = LFSRcolor1[806];
    UnbiasedRNG[361] = LFSRcolor1[68];
    UnbiasedRNG[362] = LFSRcolor1[159];
    UnbiasedRNG[363] = LFSRcolor1[1706];
    UnbiasedRNG[364] = LFSRcolor1[995];
    UnbiasedRNG[365] = LFSRcolor1[1038];
    UnbiasedRNG[366] = LFSRcolor1[108];
    UnbiasedRNG[367] = LFSRcolor1[1185];
    UnbiasedRNG[368] = LFSRcolor1[156];
    UnbiasedRNG[369] = LFSRcolor1[741];
    UnbiasedRNG[370] = LFSRcolor1[1542];
    UnbiasedRNG[371] = LFSRcolor1[808];
    UnbiasedRNG[372] = LFSRcolor1[1555];
    UnbiasedRNG[373] = LFSRcolor1[733];
    UnbiasedRNG[374] = LFSRcolor1[665];
    UnbiasedRNG[375] = LFSRcolor1[872];
    UnbiasedRNG[376] = LFSRcolor1[348];
    UnbiasedRNG[377] = LFSRcolor1[1280];
    UnbiasedRNG[378] = LFSRcolor1[633];
    UnbiasedRNG[379] = LFSRcolor1[1716];
    UnbiasedRNG[380] = LFSRcolor1[244];
    UnbiasedRNG[381] = LFSRcolor1[917];
    UnbiasedRNG[382] = LFSRcolor1[225];
    UnbiasedRNG[383] = LFSRcolor1[651];
    UnbiasedRNG[384] = LFSRcolor1[1618];
    UnbiasedRNG[385] = LFSRcolor1[274];
    UnbiasedRNG[386] = LFSRcolor1[1227];
    UnbiasedRNG[387] = LFSRcolor1[1149];
    UnbiasedRNG[388] = LFSRcolor1[694];
    UnbiasedRNG[389] = LFSRcolor1[141];
    UnbiasedRNG[390] = LFSRcolor1[1127];
    UnbiasedRNG[391] = LFSRcolor1[531];
    UnbiasedRNG[392] = LFSRcolor1[1647];
    UnbiasedRNG[393] = LFSRcolor1[1257];
    UnbiasedRNG[394] = LFSRcolor1[849];
    UnbiasedRNG[395] = LFSRcolor1[1345];
    UnbiasedRNG[396] = LFSRcolor1[1699];
    UnbiasedRNG[397] = LFSRcolor1[198];
    UnbiasedRNG[398] = LFSRcolor1[1540];
    UnbiasedRNG[399] = LFSRcolor1[832];
    UnbiasedRNG[400] = LFSRcolor1[1232];
    UnbiasedRNG[401] = LFSRcolor1[981];
    UnbiasedRNG[402] = LFSRcolor1[1273];
    UnbiasedRNG[403] = LFSRcolor1[568];
    UnbiasedRNG[404] = LFSRcolor1[351];
    UnbiasedRNG[405] = LFSRcolor1[1669];
    UnbiasedRNG[406] = LFSRcolor1[731];
    UnbiasedRNG[407] = LFSRcolor1[1688];
    UnbiasedRNG[408] = LFSRcolor1[1082];
    UnbiasedRNG[409] = LFSRcolor1[371];
    UnbiasedRNG[410] = LFSRcolor1[871];
    UnbiasedRNG[411] = LFSRcolor1[186];
    UnbiasedRNG[412] = LFSRcolor1[904];
    UnbiasedRNG[413] = LFSRcolor1[3];
    UnbiasedRNG[414] = LFSRcolor1[720];
    UnbiasedRNG[415] = LFSRcolor1[644];
    UnbiasedRNG[416] = LFSRcolor1[1586];
    UnbiasedRNG[417] = LFSRcolor1[577];
    UnbiasedRNG[418] = LFSRcolor1[1465];
    UnbiasedRNG[419] = LFSRcolor1[634];
    UnbiasedRNG[420] = LFSRcolor1[1263];
    UnbiasedRNG[421] = LFSRcolor1[533];
    UnbiasedRNG[422] = LFSRcolor1[1705];
    UnbiasedRNG[423] = LFSRcolor1[188];
    UnbiasedRNG[424] = LFSRcolor1[619];
    UnbiasedRNG[425] = LFSRcolor1[313];
    UnbiasedRNG[426] = LFSRcolor1[672];
    UnbiasedRNG[427] = LFSRcolor1[900];
    UnbiasedRNG[428] = LFSRcolor1[1006];
    UnbiasedRNG[429] = LFSRcolor1[492];
    UnbiasedRNG[430] = LFSRcolor1[1518];
    UnbiasedRNG[431] = LFSRcolor1[357];
    UnbiasedRNG[432] = LFSRcolor1[1202];
    UnbiasedRNG[433] = LFSRcolor1[1746];
    UnbiasedRNG[434] = LFSRcolor1[1242];
    UnbiasedRNG[435] = LFSRcolor1[1323];
    UnbiasedRNG[436] = LFSRcolor1[155];
    UnbiasedRNG[437] = LFSRcolor1[47];
    UnbiasedRNG[438] = LFSRcolor1[1129];
    UnbiasedRNG[439] = LFSRcolor1[862];
    UnbiasedRNG[440] = LFSRcolor1[833];
    UnbiasedRNG[441] = LFSRcolor1[1409];
    UnbiasedRNG[442] = LFSRcolor1[1292];
    UnbiasedRNG[443] = LFSRcolor1[1782];
    UnbiasedRNG[444] = LFSRcolor1[606];
    UnbiasedRNG[445] = LFSRcolor1[380];
    UnbiasedRNG[446] = LFSRcolor1[1446];
    UnbiasedRNG[447] = LFSRcolor1[65];
    UnbiasedRNG[448] = LFSRcolor1[1506];
    UnbiasedRNG[449] = LFSRcolor1[780];
    UnbiasedRNG[450] = LFSRcolor1[1767];
    UnbiasedRNG[451] = LFSRcolor1[662];
    UnbiasedRNG[452] = LFSRcolor1[1501];
    UnbiasedRNG[453] = LFSRcolor1[1258];
    UnbiasedRNG[454] = LFSRcolor1[1717];
    UnbiasedRNG[455] = LFSRcolor1[882];
    UnbiasedRNG[456] = LFSRcolor1[1433];
    UnbiasedRNG[457] = LFSRcolor1[277];
    UnbiasedRNG[458] = LFSRcolor1[465];
    UnbiasedRNG[459] = LFSRcolor1[1269];
    UnbiasedRNG[460] = LFSRcolor1[1685];
    UnbiasedRNG[461] = LFSRcolor1[1562];
    UnbiasedRNG[462] = LFSRcolor1[1672];
    UnbiasedRNG[463] = LFSRcolor1[605];
    UnbiasedRNG[464] = LFSRcolor1[1580];
    UnbiasedRNG[465] = LFSRcolor1[1479];
    UnbiasedRNG[466] = LFSRcolor1[826];
    UnbiasedRNG[467] = LFSRcolor1[569];
    UnbiasedRNG[468] = LFSRcolor1[1013];
    UnbiasedRNG[469] = LFSRcolor1[576];
    UnbiasedRNG[470] = LFSRcolor1[803];
    UnbiasedRNG[471] = LFSRcolor1[1382];
    UnbiasedRNG[472] = LFSRcolor1[1130];
    UnbiasedRNG[473] = LFSRcolor1[1758];
    UnbiasedRNG[474] = LFSRcolor1[784];
    UnbiasedRNG[475] = LFSRcolor1[547];
    UnbiasedRNG[476] = LFSRcolor1[410];
    UnbiasedRNG[477] = LFSRcolor1[133];
    UnbiasedRNG[478] = LFSRcolor1[78];
    UnbiasedRNG[479] = LFSRcolor1[359];
    UnbiasedRNG[480] = LFSRcolor1[1426];
    UnbiasedRNG[481] = LFSRcolor1[700];
    UnbiasedRNG[482] = LFSRcolor1[757];
    UnbiasedRNG[483] = LFSRcolor1[395];
    UnbiasedRNG[484] = LFSRcolor1[293];
    UnbiasedRNG[485] = LFSRcolor1[783];
    UnbiasedRNG[486] = LFSRcolor1[678];
    UnbiasedRNG[487] = LFSRcolor1[219];
    UnbiasedRNG[488] = LFSRcolor1[1444];
    UnbiasedRNG[489] = LFSRcolor1[432];
    UnbiasedRNG[490] = LFSRcolor1[837];
    UnbiasedRNG[491] = LFSRcolor1[1702];
    UnbiasedRNG[492] = LFSRcolor1[1177];
    UnbiasedRNG[493] = LFSRcolor1[486];
    UnbiasedRNG[494] = LFSRcolor1[1103];
    UnbiasedRNG[495] = LFSRcolor1[390];
end

always @(posedge color1_clk) begin
    BiasedRNG[639] = (LFSRcolor2[1263]&LFSRcolor2[668]&LFSRcolor2[1088]&LFSRcolor2[530]);
    BiasedRNG[640] = (LFSRcolor2[29]&LFSRcolor2[474]&LFSRcolor2[793]&LFSRcolor2[707]);
    BiasedRNG[641] = (LFSRcolor2[1272]&LFSRcolor2[508]&LFSRcolor2[828]&LFSRcolor2[451]);
    BiasedRNG[642] = (LFSRcolor2[999]&LFSRcolor2[1145]&LFSRcolor2[1062]&LFSRcolor2[3]);
    BiasedRNG[643] = (LFSRcolor2[354]&LFSRcolor2[475]&LFSRcolor2[1044]&LFSRcolor2[157]);
    BiasedRNG[644] = (LFSRcolor2[19]&LFSRcolor2[889]&LFSRcolor2[533]&LFSRcolor2[928]);
    BiasedRNG[645] = (LFSRcolor2[102]&LFSRcolor2[346]&LFSRcolor2[972]&LFSRcolor2[796]);
    BiasedRNG[646] = (LFSRcolor2[446]&LFSRcolor2[995]&LFSRcolor2[761]&LFSRcolor2[1205]);
    BiasedRNG[647] = (LFSRcolor2[421]&LFSRcolor2[1011]&LFSRcolor2[612]&LFSRcolor2[1220]);
    BiasedRNG[648] = (LFSRcolor2[142]&LFSRcolor2[914]&LFSRcolor2[265]&LFSRcolor2[223]);
    BiasedRNG[649] = (LFSRcolor2[602]&LFSRcolor2[1214]&LFSRcolor2[1253]&LFSRcolor2[450]);
    BiasedRNG[650] = (LFSRcolor2[731]&LFSRcolor2[1041]&LFSRcolor2[231]&LFSRcolor2[639]);
    BiasedRNG[651] = (LFSRcolor2[589]&LFSRcolor2[100]&LFSRcolor2[94]&LFSRcolor2[273]);
    BiasedRNG[652] = (LFSRcolor2[1071]&LFSRcolor2[815]&LFSRcolor2[6]&LFSRcolor2[314]);
    BiasedRNG[653] = (LFSRcolor2[1069]&LFSRcolor2[746]&LFSRcolor2[578]&LFSRcolor2[1188]);
    BiasedRNG[654] = (LFSRcolor2[30]&LFSRcolor2[859]&LFSRcolor2[1147]&LFSRcolor2[232]);
    BiasedRNG[655] = (LFSRcolor2[74]&LFSRcolor2[374]&LFSRcolor2[194]&LFSRcolor2[950]);
    BiasedRNG[656] = (LFSRcolor2[1081]&LFSRcolor2[55]&LFSRcolor2[717]&LFSRcolor2[247]);
    BiasedRNG[657] = (LFSRcolor2[593]&LFSRcolor2[1240]&LFSRcolor2[515]&LFSRcolor2[197]);
    BiasedRNG[658] = (LFSRcolor2[177]&LFSRcolor2[316]&LFSRcolor2[33]&LFSRcolor2[483]);
    BiasedRNG[659] = (LFSRcolor2[1164]&LFSRcolor2[188]&LFSRcolor2[1207]&LFSRcolor2[460]);
    BiasedRNG[660] = (LFSRcolor2[583]&LFSRcolor2[1166]&LFSRcolor2[923]&LFSRcolor2[736]);
    BiasedRNG[661] = (LFSRcolor2[62]&LFSRcolor2[866]&LFSRcolor2[686]&LFSRcolor2[820]);
    BiasedRNG[662] = (LFSRcolor2[153]&LFSRcolor2[1172]&LFSRcolor2[1236]&LFSRcolor2[375]);
    BiasedRNG[663] = (LFSRcolor2[766]&LFSRcolor2[581]&LFSRcolor2[984]&LFSRcolor2[468]);
    BiasedRNG[664] = (LFSRcolor2[1268]&LFSRcolor2[149]&LFSRcolor2[242]&LFSRcolor2[559]);
    BiasedRNG[665] = (LFSRcolor2[634]&LFSRcolor2[1130]&LFSRcolor2[66]&LFSRcolor2[814]);
    BiasedRNG[666] = (LFSRcolor2[401]&LFSRcolor2[136]&LFSRcolor2[509]&LFSRcolor2[418]);
    BiasedRNG[667] = (LFSRcolor2[20]&LFSRcolor2[938]&LFSRcolor2[1157]&LFSRcolor2[58]);
    BiasedRNG[668] = (LFSRcolor2[447]&LFSRcolor2[675]&LFSRcolor2[817]&LFSRcolor2[1136]);
    BiasedRNG[669] = (LFSRcolor2[255]&LFSRcolor2[881]&LFSRcolor2[235]&LFSRcolor2[737]);
    BiasedRNG[670] = (LFSRcolor2[1007]&LFSRcolor2[1061]&LFSRcolor2[396]&LFSRcolor2[229]);
    BiasedRNG[671] = (LFSRcolor2[270]&LFSRcolor2[1042]&LFSRcolor2[751]&LFSRcolor2[1196]);
    BiasedRNG[672] = (LFSRcolor2[1161]&LFSRcolor2[37]&LFSRcolor2[558]&LFSRcolor2[308]);
    BiasedRNG[673] = (LFSRcolor2[63]&LFSRcolor2[464]&LFSRcolor2[549]&LFSRcolor2[579]);
    BiasedRNG[674] = (LFSRcolor2[1216]&LFSRcolor2[544]&LFSRcolor2[1075]&LFSRcolor2[221]);
    BiasedRNG[675] = (LFSRcolor2[321]&LFSRcolor2[115]&LFSRcolor2[516]&LFSRcolor2[688]);
    BiasedRNG[676] = (LFSRcolor2[754]&LFSRcolor2[669]&LFSRcolor2[1057]&LFSRcolor2[327]);
    BiasedRNG[677] = (LFSRcolor2[1107]&LFSRcolor2[905]&LFSRcolor2[384]&LFSRcolor2[279]);
    BiasedRNG[678] = (LFSRcolor2[1090]&LFSRcolor2[876]&LFSRcolor2[1143]&LFSRcolor2[187]);
    BiasedRNG[679] = (LFSRcolor2[1033]&LFSRcolor2[1036]&LFSRcolor2[1050]&LFSRcolor2[543]);
    BiasedRNG[680] = (LFSRcolor2[159]&LFSRcolor2[986]&LFSRcolor2[35]&LFSRcolor2[1177]);
    BiasedRNG[681] = (LFSRcolor2[910]&LFSRcolor2[47]&LFSRcolor2[249]&LFSRcolor2[363]);
    BiasedRNG[682] = (LFSRcolor2[1219]&LFSRcolor2[722]&LFSRcolor2[302]&LFSRcolor2[933]);
    BiasedRNG[683] = (LFSRcolor2[880]&LFSRcolor2[521]&LFSRcolor2[1278]&LFSRcolor2[745]);
    BiasedRNG[684] = (LFSRcolor2[811]&LFSRcolor2[156]&LFSRcolor2[61]&LFSRcolor2[858]);
    BiasedRNG[685] = (LFSRcolor2[609]&LFSRcolor2[104]&LFSRcolor2[266]&LFSRcolor2[1001]);
    BiasedRNG[686] = (LFSRcolor2[777]&LFSRcolor2[762]&LFSRcolor2[1258]&LFSRcolor2[69]);
    BiasedRNG[687] = (LFSRcolor2[1048]&LFSRcolor2[961]&LFSRcolor2[1248]&LFSRcolor2[729]);
    BiasedRNG[688] = (LFSRcolor2[903]&LFSRcolor2[584]&LFSRcolor2[598]&LFSRcolor2[196]);
    BiasedRNG[689] = (LFSRcolor2[629]&LFSRcolor2[994]&LFSRcolor2[1068]&LFSRcolor2[288]);
    BiasedRNG[690] = (LFSRcolor2[1101]&LFSRcolor2[476]&LFSRcolor2[46]&LFSRcolor2[503]);
    BiasedRNG[691] = (LFSRcolor2[1226]&LFSRcolor2[730]&LFSRcolor2[224]&LFSRcolor2[806]);
    BiasedRNG[692] = (LFSRcolor2[1039]&LFSRcolor2[748]&LFSRcolor2[1091]&LFSRcolor2[109]);
    BiasedRNG[693] = (LFSRcolor2[840]&LFSRcolor2[304]&LFSRcolor2[630]&LFSRcolor2[557]);
    BiasedRNG[694] = (LFSRcolor2[671]&LFSRcolor2[1179]&LFSRcolor2[932]&LFSRcolor2[172]);
    BiasedRNG[695] = (LFSRcolor2[538]&LFSRcolor2[676]&LFSRcolor2[1189]&LFSRcolor2[871]);
    BiasedRNG[696] = (LFSRcolor2[107]&LFSRcolor2[580]&LFSRcolor2[661]&LFSRcolor2[254]);
    BiasedRNG[697] = (LFSRcolor2[438]&LFSRcolor2[361]&LFSRcolor2[1265]&LFSRcolor2[1133]);
    BiasedRNG[698] = (LFSRcolor2[267]&LFSRcolor2[1000]&LFSRcolor2[114]&LFSRcolor2[642]);
    BiasedRNG[699] = (LFSRcolor2[443]&LFSRcolor2[939]&LFSRcolor2[146]&LFSRcolor2[40]);
    BiasedRNG[700] = (LFSRcolor2[1051]&LFSRcolor2[556]&LFSRcolor2[1217]&LFSRcolor2[1016]);
    BiasedRNG[701] = (LFSRcolor2[162]&LFSRcolor2[43]&LFSRcolor2[175]&LFSRcolor2[1246]);
    BiasedRNG[702] = (LFSRcolor2[1089]&LFSRcolor2[597]&LFSRcolor2[127]&LFSRcolor2[1054]);
    BiasedRNG[703] = (LFSRcolor2[442]&LFSRcolor2[383]&LFSRcolor2[1203]&LFSRcolor2[621]);
    BiasedRNG[704] = (LFSRcolor2[457]&LFSRcolor2[329]&LFSRcolor2[779]&LFSRcolor2[1080]);
    BiasedRNG[705] = (LFSRcolor2[407]&LFSRcolor2[484]&LFSRcolor2[763]&LFSRcolor2[957]);
    BiasedRNG[706] = (LFSRcolor2[497]&LFSRcolor2[571]&LFSRcolor2[1031]&LFSRcolor2[1002]);
    BiasedRNG[707] = (LFSRcolor2[555]&LFSRcolor2[572]&LFSRcolor2[1021]&LFSRcolor2[241]);
    BiasedRNG[708] = (LFSRcolor2[341]&LFSRcolor2[560]&LFSRcolor2[334]&LFSRcolor2[546]);
    BiasedRNG[709] = (LFSRcolor2[121]&LFSRcolor2[166]&LFSRcolor2[394]&LFSRcolor2[253]);
    BiasedRNG[710] = (LFSRcolor2[582]&LFSRcolor2[927]&LFSRcolor2[295]&LFSRcolor2[90]);
    BiasedRNG[711] = (LFSRcolor2[816]&LFSRcolor2[216]&LFSRcolor2[332]&LFSRcolor2[622]);
    BiasedRNG[712] = (LFSRcolor2[168]&LFSRcolor2[171]&LFSRcolor2[1029]&LFSRcolor2[452]);
    BiasedRNG[713] = (LFSRcolor2[1167]&LFSRcolor2[1117]&LFSRcolor2[1153]&LFSRcolor2[207]);
    BiasedRNG[714] = (LFSRcolor2[528]&LFSRcolor2[896]&LFSRcolor2[495]&LFSRcolor2[217]);
    BiasedRNG[715] = (LFSRcolor2[431]&LFSRcolor2[710]&LFSRcolor2[853]&LFSRcolor2[651]);
    BiasedRNG[716] = (LFSRcolor2[1023]&LFSRcolor2[26]&LFSRcolor2[390]&LFSRcolor2[141]);
    BiasedRNG[717] = (LFSRcolor2[1247]&LFSRcolor2[805]&LFSRcolor2[500]&LFSRcolor2[850]);
    BiasedRNG[718] = (LFSRcolor2[1025]&LFSRcolor2[603]&LFSRcolor2[918]&LFSRcolor2[728]);
    BiasedRNG[719] = (LFSRcolor2[1168]&LFSRcolor2[181]&LFSRcolor2[861]&LFSRcolor2[656]);
    BiasedRNG[720] = (LFSRcolor2[381]&LFSRcolor2[420]&LFSRcolor2[548]&LFSRcolor2[883]);
    BiasedRNG[721] = (LFSRcolor2[1221]&LFSRcolor2[236]&LFSRcolor2[764]&LFSRcolor2[1015]);
    BiasedRNG[722] = (LFSRcolor2[1019]&LFSRcolor2[971]&LFSRcolor2[262]&LFSRcolor2[339]);
    BiasedRNG[723] = (LFSRcolor2[1202]&LFSRcolor2[898]&LFSRcolor2[49]&LFSRcolor2[692]);
    BiasedRNG[724] = (LFSRcolor2[180]&LFSRcolor2[203]&LFSRcolor2[1104]&LFSRcolor2[365]);
    BiasedRNG[725] = (LFSRcolor2[264]&LFSRcolor2[344]&LFSRcolor2[313]&LFSRcolor2[818]);
    BiasedRNG[726] = (LFSRcolor2[1077]&LFSRcolor2[887]&LFSRcolor2[380]&LFSRcolor2[408]);
    BiasedRNG[727] = (LFSRcolor2[849]&LFSRcolor2[563]&LFSRcolor2[931]&LFSRcolor2[890]);
    BiasedRNG[728] = (LFSRcolor2[1280]&LFSRcolor2[997]&LFSRcolor2[1200]&LFSRcolor2[623]);
    BiasedRNG[729] = (LFSRcolor2[192]&LFSRcolor2[373]&LFSRcolor2[205]&LFSRcolor2[1178]);
    BiasedRNG[730] = (LFSRcolor2[1225]&LFSRcolor2[1230]&LFSRcolor2[988]&LFSRcolor2[429]);
    BiasedRNG[731] = (LFSRcolor2[195]&LFSRcolor2[1195]&LFSRcolor2[113]&LFSRcolor2[499]);
    BiasedRNG[732] = (LFSRcolor2[1149]&LFSRcolor2[38]&LFSRcolor2[386]&LFSRcolor2[741]);
    BiasedRNG[733] = (LFSRcolor2[1154]&LFSRcolor2[869]&LFSRcolor2[286]&LFSRcolor2[1087]);
    BiasedRNG[734] = (LFSRcolor2[1204]&LFSRcolor2[713]&LFSRcolor2[190]&LFSRcolor2[1233]);
    BiasedRNG[735] = (LFSRcolor2[1274]&LFSRcolor2[1187]&LFSRcolor2[1284]&LFSRcolor2[691]);
    BiasedRNG[736] = (LFSRcolor2[160]&LFSRcolor2[1037]&LFSRcolor2[591]&LFSRcolor2[738]);
    BiasedRNG[737] = (LFSRcolor2[716]&LFSRcolor2[326]&LFSRcolor2[222]&LFSRcolor2[899]);
    BiasedRNG[738] = (LFSRcolor2[1063]&LFSRcolor2[554]&LFSRcolor2[1171]&LFSRcolor2[54]);
    BiasedRNG[739] = (LFSRcolor2[16]&LFSRcolor2[366]&LFSRcolor2[21]&LFSRcolor2[1234]);
    BiasedRNG[740] = (LFSRcolor2[888]&LFSRcolor2[309]&LFSRcolor2[632]&LFSRcolor2[740]);
    BiasedRNG[741] = (LFSRcolor2[864]&LFSRcolor2[263]&LFSRcolor2[574]&LFSRcolor2[935]);
    BiasedRNG[742] = (LFSRcolor2[1218]&LFSRcolor2[570]&LFSRcolor2[228]&LFSRcolor2[960]);
    BiasedRNG[743] = (LFSRcolor2[488]&LFSRcolor2[893]&LFSRcolor2[1201]&LFSRcolor2[300]);
    BiasedRNG[744] = (LFSRcolor2[310]&LFSRcolor2[750]&LFSRcolor2[1120]&LFSRcolor2[809]);
    BiasedRNG[745] = (LFSRcolor2[610]&LFSRcolor2[836]&LFSRcolor2[536]&LFSRcolor2[683]);
    BiasedRNG[746] = (LFSRcolor2[182]&LFSRcolor2[993]&LFSRcolor2[347]&LFSRcolor2[425]);
    BiasedRNG[747] = (LFSRcolor2[826]&LFSRcolor2[714]&LFSRcolor2[250]&LFSRcolor2[117]);
    BiasedRNG[748] = (LFSRcolor2[542]&LFSRcolor2[130]&LFSRcolor2[1093]&LFSRcolor2[727]);
    BiasedRNG[749] = (LFSRcolor2[246]&LFSRcolor2[1140]&LFSRcolor2[843]&LFSRcolor2[284]);
    BiasedRNG[750] = (LFSRcolor2[440]&LFSRcolor2[1275]&LFSRcolor2[1215]&LFSRcolor2[204]);
    BiasedRNG[751] = (LFSRcolor2[448]&LFSRcolor2[1123]&LFSRcolor2[645]&LFSRcolor2[59]);
    BiasedRNG[752] = (LFSRcolor2[875]&LFSRcolor2[663]&LFSRcolor2[919]&LFSRcolor2[70]);
    BiasedRNG[753] = (LFSRcolor2[522]&LFSRcolor2[834]&LFSRcolor2[916]&LFSRcolor2[813]);
    BiasedRNG[754] = (LFSRcolor2[118]&LFSRcolor2[776]&LFSRcolor2[1092]&LFSRcolor2[77]);
    BiasedRNG[755] = (LFSRcolor2[787]&LFSRcolor2[1102]&LFSRcolor2[930]&LFSRcolor2[439]);
    BiasedRNG[756] = (LFSRcolor2[409]&LFSRcolor2[564]&LFSRcolor2[998]&LFSRcolor2[650]);
    BiasedRNG[757] = (LFSRcolor2[747]&LFSRcolor2[28]&LFSRcolor2[703]&LFSRcolor2[1199]);
    BiasedRNG[758] = (LFSRcolor2[342]&LFSRcolor2[27]&LFSRcolor2[87]&LFSRcolor2[856]);
    BiasedRNG[759] = (LFSRcolor2[230]&LFSRcolor2[1010]&LFSRcolor2[699]&LFSRcolor2[1059]);
    BiasedRNG[760] = (LFSRcolor2[356]&LFSRcolor2[783]&LFSRcolor2[897]&LFSRcolor2[1251]);
    BiasedRNG[761] = (LFSRcolor2[406]&LFSRcolor2[139]&LFSRcolor2[592]&LFSRcolor2[274]);
    BiasedRNG[762] = (LFSRcolor2[1232]&LFSRcolor2[937]&LFSRcolor2[1222]&LFSRcolor2[167]);
    BiasedRNG[763] = (LFSRcolor2[1116]&LFSRcolor2[292]&LFSRcolor2[307]&LFSRcolor2[257]);
    BiasedRNG[764] = (LFSRcolor2[635]&LFSRcolor2[1262]&LFSRcolor2[507]&LFSRcolor2[531]);
    BiasedRNG[765] = (LFSRcolor2[912]&LFSRcolor2[336]&LFSRcolor2[98]&LFSRcolor2[36]);
    BiasedRNG[766] = (LFSRcolor2[185]&LFSRcolor2[48]&LFSRcolor2[1198]&LFSRcolor2[1245]);
    BiasedRNG[767] = (LFSRcolor2[872]&LFSRcolor2[788]&LFSRcolor2[165]&LFSRcolor2[289]);
    BiasedRNG[768] = (LFSRcolor2[1254]&LFSRcolor2[829]&LFSRcolor2[99]&LFSRcolor2[470]);
    BiasedRNG[769] = (LFSRcolor2[1127]&LFSRcolor2[970]&LFSRcolor2[697]&LFSRcolor2[744]);
    BiasedRNG[770] = (LFSRcolor2[1257]&LFSRcolor2[680]&LFSRcolor2[1279]&LFSRcolor2[12]);
    BiasedRNG[771] = (LFSRcolor2[311]&LFSRcolor2[1122]&LFSRcolor2[989]&LFSRcolor2[477]);
    BiasedRNG[772] = (LFSRcolor2[1197]&LFSRcolor2[135]&LFSRcolor2[44]&LFSRcolor2[124]);
    BiasedRNG[773] = (LFSRcolor2[298]&LFSRcolor2[550]&LFSRcolor2[68]&LFSRcolor2[1238]);
    BiasedRNG[774] = (LFSRcolor2[403]&LFSRcolor2[322]&LFSRcolor2[388]&LFSRcolor2[371]);
    BiasedRNG[775] = (LFSRcolor2[333]&LFSRcolor2[891]&LFSRcolor2[693]&LFSRcolor2[1287]);
    BiasedRNG[776] = (LFSRcolor2[22]&LFSRcolor2[791]&LFSRcolor2[832]&LFSRcolor2[1260]);
    BiasedRNG[777] = (LFSRcolor2[367]&LFSRcolor2[116]&LFSRcolor2[218]&LFSRcolor2[337]);
    BiasedRNG[778] = (LFSRcolor2[143]&LFSRcolor2[1106]&LFSRcolor2[379]&LFSRcolor2[189]);
    BiasedRNG[779] = (LFSRcolor2[1073]&LFSRcolor2[1244]&LFSRcolor2[773]&LFSRcolor2[1128]);
    BiasedRNG[780] = (LFSRcolor2[5]&LFSRcolor2[353]&LFSRcolor2[924]&LFSRcolor2[473]);
    BiasedRNG[781] = (LFSRcolor2[15]&LFSRcolor2[535]&LFSRcolor2[966]&LFSRcolor2[681]);
    BiasedRNG[782] = (LFSRcolor2[79]&LFSRcolor2[462]&LFSRcolor2[990]&LFSRcolor2[1005]);
    BiasedRNG[783] = (LFSRcolor2[870]&LFSRcolor2[616]&LFSRcolor2[774]&LFSRcolor2[441]);
    BiasedRNG[784] = (LFSRcolor2[282]&LFSRcolor2[677]&LFSRcolor2[9]&LFSRcolor2[186]);
    BiasedRNG[785] = (LFSRcolor2[845]&LFSRcolor2[552]&LFSRcolor2[1270]&LFSRcolor2[1065]);
    BiasedRNG[786] = (LFSRcolor2[387]&LFSRcolor2[934]&LFSRcolor2[414]&LFSRcolor2[112]);
    BiasedRNG[787] = (LFSRcolor2[493]&LFSRcolor2[674]&LFSRcolor2[31]&LFSRcolor2[349]);
    BiasedRNG[788] = (LFSRcolor2[1121]&LFSRcolor2[637]&LFSRcolor2[726]&LFSRcolor2[921]);
    BiasedRNG[789] = (LFSRcolor2[678]&LFSRcolor2[83]&LFSRcolor2[660]&LFSRcolor2[296]);
    BiasedRNG[790] = (LFSRcolor2[780]&LFSRcolor2[513]&LFSRcolor2[444]&LFSRcolor2[163]);
    BiasedRNG[791] = (LFSRcolor2[41]&LFSRcolor2[1129]&LFSRcolor2[733]&LFSRcolor2[665]);
    BiasedRNG[792] = (LFSRcolor2[753]&LFSRcolor2[1035]&LFSRcolor2[734]&LFSRcolor2[906]);
    BiasedRNG[793] = (LFSRcolor2[633]&LFSRcolor2[641]&LFSRcolor2[215]&LFSRcolor2[640]);
    BiasedRNG[794] = (LFSRcolor2[237]&LFSRcolor2[1227]&LFSRcolor2[985]&LFSRcolor2[857]);
    BiasedRNG[795] = (LFSRcolor2[398]&LFSRcolor2[757]&LFSRcolor2[743]&LFSRcolor2[106]);
    BiasedRNG[796] = (LFSRcolor2[1052]&LFSRcolor2[594]&LFSRcolor2[489]&LFSRcolor2[700]);
    BiasedRNG[797] = (LFSRcolor2[1212]&LFSRcolor2[715]&LFSRcolor2[1028]&LFSRcolor2[132]);
    BiasedRNG[798] = (LFSRcolor2[652]&LFSRcolor2[1003]&LFSRcolor2[244]&LFSRcolor2[649]);
    BiasedRNG[799] = (LFSRcolor2[1249]&LFSRcolor2[917]&LFSRcolor2[144]&LFSRcolor2[278]);
    BiasedRNG[800] = (LFSRcolor2[362]&LFSRcolor2[1040]&LFSRcolor2[23]&LFSRcolor2[963]);
    BiasedRNG[801] = (LFSRcolor2[644]&LFSRcolor2[525]&LFSRcolor2[285]&LFSRcolor2[147]);
    BiasedRNG[802] = (LFSRcolor2[682]&LFSRcolor2[1126]&LFSRcolor2[430]&LFSRcolor2[1017]);
    BiasedRNG[803] = (LFSRcolor2[785]&LFSRcolor2[1027]&LFSRcolor2[1229]&LFSRcolor2[614]);
    BiasedRNG[804] = (LFSRcolor2[608]&LFSRcolor2[812]&LFSRcolor2[752]&LFSRcolor2[611]);
    BiasedRNG[805] = (LFSRcolor2[838]&LFSRcolor2[239]&LFSRcolor2[1]&LFSRcolor2[877]);
    BiasedRNG[806] = (LFSRcolor2[1209]&LFSRcolor2[976]&LFSRcolor2[397]&LFSRcolor2[73]);
    BiasedRNG[807] = (LFSRcolor2[725]&LFSRcolor2[32]&LFSRcolor2[706]&LFSRcolor2[1165]);
    BiasedRNG[808] = (LFSRcolor2[666]&LFSRcolor2[685]&LFSRcolor2[945]&LFSRcolor2[718]);
    BiasedRNG[809] = (LFSRcolor2[86]&LFSRcolor2[490]&LFSRcolor2[758]&LFSRcolor2[494]);
    BiasedRNG[810] = (LFSRcolor2[1185]&LFSRcolor2[323]&LFSRcolor2[479]&LFSRcolor2[306]);
    BiasedRNG[811] = (LFSRcolor2[372]&LFSRcolor2[404]&LFSRcolor2[517]&LFSRcolor2[294]);
    BiasedRNG[812] = (LFSRcolor2[835]&LFSRcolor2[1119]&LFSRcolor2[982]&LFSRcolor2[617]);
    BiasedRNG[813] = (LFSRcolor2[359]&LFSRcolor2[895]&LFSRcolor2[1267]&LFSRcolor2[624]);
    BiasedRNG[814] = (LFSRcolor2[673]&LFSRcolor2[1163]&LFSRcolor2[413]&LFSRcolor2[862]);
    BiasedRNG[815] = (LFSRcolor2[213]&LFSRcolor2[170]&LFSRcolor2[1060]&LFSRcolor2[959]);
    BiasedRNG[816] = (LFSRcolor2[654]&LFSRcolor2[291]&LFSRcolor2[695]&LFSRcolor2[281]);
    BiasedRNG[817] = (LFSRcolor2[133]&LFSRcolor2[925]&LFSRcolor2[1241]&LFSRcolor2[863]);
    BiasedRNG[818] = (LFSRcolor2[211]&LFSRcolor2[57]&LFSRcolor2[193]&LFSRcolor2[75]);
    BiasedRNG[819] = (LFSRcolor2[434]&LFSRcolor2[576]&LFSRcolor2[679]&LFSRcolor2[1144]);
    BiasedRNG[820] = (LFSRcolor2[659]&LFSRcolor2[17]&LFSRcolor2[501]&LFSRcolor2[330]);
    BiasedRNG[821] = (LFSRcolor2[1286]&LFSRcolor2[364]&LFSRcolor2[65]&LFSRcolor2[885]);
    BiasedRNG[822] = (LFSRcolor2[11]&LFSRcolor2[1206]&LFSRcolor2[996]&LFSRcolor2[1058]);
    BiasedRNG[823] = (LFSRcolor2[214]&LFSRcolor2[335]&LFSRcolor2[368]&LFSRcolor2[1210]);
    BiasedRNG[824] = (LFSRcolor2[967]&LFSRcolor2[690]&LFSRcolor2[1024]&LFSRcolor2[148]);
    BiasedRNG[825] = (LFSRcolor2[1056]&LFSRcolor2[619]&LFSRcolor2[56]&LFSRcolor2[604]);
    BiasedRNG[826] = (LFSRcolor2[613]&LFSRcolor2[803]&LFSRcolor2[855]&LFSRcolor2[868]);
    BiasedRNG[827] = (LFSRcolor2[944]&LFSRcolor2[245]&LFSRcolor2[1114]&LFSRcolor2[790]);
    BiasedRNG[828] = (LFSRcolor2[91]&LFSRcolor2[472]&LFSRcolor2[759]&LFSRcolor2[689]);
    BiasedRNG[829] = (LFSRcolor2[378]&LFSRcolor2[52]&LFSRcolor2[648]&LFSRcolor2[909]);
    BiasedRNG[830] = (LFSRcolor2[514]&LFSRcolor2[882]&LFSRcolor2[4]&LFSRcolor2[471]);
    BiasedRNG[831] = (LFSRcolor2[878]&LFSRcolor2[1067]&LFSRcolor2[225]&LFSRcolor2[607]);
    BiasedRNG[832] = (LFSRcolor2[784]&LFSRcolor2[88]&LFSRcolor2[687]&LFSRcolor2[1170]);
    BiasedRNG[833] = (LFSRcolor2[423]&LFSRcolor2[71]&LFSRcolor2[569]&LFSRcolor2[271]);
    BiasedRNG[834] = (LFSRcolor2[1277]&LFSRcolor2[82]&LFSRcolor2[978]&LFSRcolor2[980]);
    BiasedRNG[835] = (LFSRcolor2[318]&LFSRcolor2[393]&LFSRcolor2[1252]&LFSRcolor2[325]);
    BiasedRNG[836] = (LFSRcolor2[1014]&LFSRcolor2[951]&LFSRcolor2[1098]&LFSRcolor2[481]);
    BiasedRNG[837] = (LFSRcolor2[103]&LFSRcolor2[251]&LFSRcolor2[210]&LFSRcolor2[467]);
    BiasedRNG[838] = (LFSRcolor2[831]&LFSRcolor2[428]&LFSRcolor2[865]&LFSRcolor2[426]);
    BiasedRNG[839] = (LFSRcolor2[1142]&LFSRcolor2[164]&LFSRcolor2[174]&LFSRcolor2[1281]);
    BiasedRNG[840] = (LFSRcolor2[510]&LFSRcolor2[987]&LFSRcolor2[125]&LFSRcolor2[915]);
    BiasedRNG[841] = (LFSRcolor2[1066]&LFSRcolor2[1175]&LFSRcolor2[176]&LFSRcolor2[105]);
    BiasedRNG[842] = (LFSRcolor2[566]&LFSRcolor2[498]&LFSRcolor2[799]&LFSRcolor2[80]);
    BiasedRNG[843] = (LFSRcolor2[1034]&LFSRcolor2[1103]&LFSRcolor2[672]&LFSRcolor2[599]);
    BiasedRNG[844] = (LFSRcolor2[1231]&LFSRcolor2[860]&LFSRcolor2[1176]&LFSRcolor2[537]);
    BiasedRNG[845] = (LFSRcolor2[395]&LFSRcolor2[453]&LFSRcolor2[590]&LFSRcolor2[756]);
    BiasedRNG[846] = (LFSRcolor2[417]&LFSRcolor2[568]&LFSRcolor2[1158]&LFSRcolor2[1183]);
    BiasedRNG[847] = (LFSRcolor2[1097]&LFSRcolor2[606]&LFSRcolor2[14]&LFSRcolor2[64]);
    BiasedRNG[848] = (LFSRcolor2[502]&LFSRcolor2[586]&LFSRcolor2[702]&LFSRcolor2[258]);
    BiasedRNG[849] = (LFSRcolor2[1174]&LFSRcolor2[436]&LFSRcolor2[601]&LFSRcolor2[600]);
    BiasedRNG[850] = (LFSRcolor2[2]&LFSRcolor2[1155]&LFSRcolor2[1156]&LFSRcolor2[704]);
    BiasedRNG[851] = (LFSRcolor2[772]&LFSRcolor2[385]&LFSRcolor2[810]&LFSRcolor2[34]);
    BiasedRNG[852] = (LFSRcolor2[191]&LFSRcolor2[775]&LFSRcolor2[389]&LFSRcolor2[76]);
    BiasedRNG[853] = (LFSRcolor2[721]&LFSRcolor2[50]&LFSRcolor2[819]&LFSRcolor2[1109]);
    BiasedRNG[854] = (LFSRcolor2[698]&LFSRcolor2[324]&LFSRcolor2[965]&LFSRcolor2[454]);
    BiasedRNG[855] = (LFSRcolor2[527]&LFSRcolor2[220]&LFSRcolor2[7]&LFSRcolor2[991]);
    BiasedRNG[856] = (LFSRcolor2[466]&LFSRcolor2[42]&LFSRcolor2[958]&LFSRcolor2[1182]);
    BiasedRNG[857] = (LFSRcolor2[711]&LFSRcolor2[940]&LFSRcolor2[122]&LFSRcolor2[427]);
    BiasedRNG[858] = (LFSRcolor2[1152]&LFSRcolor2[348]&LFSRcolor2[39]&LFSRcolor2[701]);
    BiasedRNG[859] = (LFSRcolor2[823]&LFSRcolor2[0]&LFSRcolor2[1085]&LFSRcolor2[1193]);
    BiasedRNG[860] = (LFSRcolor2[620]&LFSRcolor2[742]&LFSRcolor2[60]&LFSRcolor2[199]);
    BiasedRNG[861] = (LFSRcolor2[781]&LFSRcolor2[605]&LFSRcolor2[360]&LFSRcolor2[907]);
    BiasedRNG[862] = (LFSRcolor2[1173]&LFSRcolor2[948]&LFSRcolor2[767]&LFSRcolor2[827]);
    BiasedRNG[863] = (LFSRcolor2[485]&LFSRcolor2[646]&LFSRcolor2[1264]&LFSRcolor2[1137]);
    BiasedRNG[864] = (LFSRcolor2[206]&LFSRcolor2[227]&LFSRcolor2[432]&LFSRcolor2[854]);
    BiasedRNG[865] = (LFSRcolor2[1045]&LFSRcolor2[496]&LFSRcolor2[252]&LFSRcolor2[873]);
    BiasedRNG[866] = (LFSRcolor2[1184]&LFSRcolor2[708]&LFSRcolor2[248]&LFSRcolor2[801]);
    BiasedRNG[867] = (LFSRcolor2[667]&LFSRcolor2[575]&LFSRcolor2[280]&LFSRcolor2[1111]);
    BiasedRNG[868] = (LFSRcolor2[1115]&LFSRcolor2[400]&LFSRcolor2[901]&LFSRcolor2[1180]);
    BiasedRNG[869] = (LFSRcolor2[786]&LFSRcolor2[627]&LFSRcolor2[1086]&LFSRcolor2[647]);
    BiasedRNG[870] = (LFSRcolor2[769]&LFSRcolor2[1020]&LFSRcolor2[1026]&LFSRcolor2[276]);
    BiasedRNG[871] = (LFSRcolor2[942]&LFSRcolor2[1094]&LFSRcolor2[134]&LFSRcolor2[523]);
    BiasedRNG[872] = (LFSRcolor2[299]&LFSRcolor2[84]&LFSRcolor2[511]&LFSRcolor2[1190]);
    BiasedRNG[873] = (LFSRcolor2[1009]&LFSRcolor2[1273]&LFSRcolor2[1013]&LFSRcolor2[789]);
    BiasedRNG[874] = (LFSRcolor2[119]&LFSRcolor2[1283]&LFSRcolor2[419]&LFSRcolor2[1064]);
    BiasedRNG[875] = (LFSRcolor2[1038]&LFSRcolor2[657]&LFSRcolor2[947]&LFSRcolor2[545]);
    BiasedRNG[876] = (LFSRcolor2[975]&LFSRcolor2[129]&LFSRcolor2[422]&LFSRcolor2[376]);
    BiasedRNG[877] = (LFSRcolor2[969]&LFSRcolor2[705]&LFSRcolor2[145]&LFSRcolor2[184]);
    BiasedRNG[878] = (LFSRcolor2[89]&LFSRcolor2[664]&LFSRcolor2[392]&LFSRcolor2[618]);
    BiasedRNG[879] = (LFSRcolor2[1112]&LFSRcolor2[1186]&LFSRcolor2[92]&LFSRcolor2[760]);
    BiasedRNG[880] = (LFSRcolor2[137]&LFSRcolor2[140]&LFSRcolor2[662]&LFSRcolor2[128]);
    BiasedRNG[881] = (LFSRcolor2[983]&LFSRcolor2[238]&LFSRcolor2[411]&LFSRcolor2[350]);
    BiasedRNG[882] = (LFSRcolor2[256]&LFSRcolor2[540]&LFSRcolor2[1194]&LFSRcolor2[981]);
    BiasedRNG[883] = (LFSRcolor2[93]&LFSRcolor2[268]&LFSRcolor2[908]&LFSRcolor2[259]);
    BiasedRNG[884] = (LFSRcolor2[1030]&LFSRcolor2[67]&LFSRcolor2[410]&LFSRcolor2[377]);
    BiasedRNG[885] = (LFSRcolor2[962]&LFSRcolor2[1055]&LFSRcolor2[964]&LFSRcolor2[491]);
    BiasedRNG[886] = (LFSRcolor2[351]&LFSRcolor2[97]&LFSRcolor2[839]&LFSRcolor2[312]);
    BiasedRNG[887] = (LFSRcolor2[841]&LFSRcolor2[1138]&LFSRcolor2[161]&LFSRcolor2[732]);
    BiasedRNG[888] = (LFSRcolor2[847]&LFSRcolor2[275]&LFSRcolor2[1213]&LFSRcolor2[825]);
    BiasedRNG[889] = (LFSRcolor2[461]&LFSRcolor2[625]&LFSRcolor2[72]&LFSRcolor2[804]);
    BiasedRNG[890] = (LFSRcolor2[110]&LFSRcolor2[486]&LFSRcolor2[1160]&LFSRcolor2[340]);
    BiasedRNG[891] = (LFSRcolor2[1237]&LFSRcolor2[492]&LFSRcolor2[169]&LFSRcolor2[1047]);
    BiasedRNG[892] = (LFSRcolor2[770]&LFSRcolor2[269]&LFSRcolor2[636]&LFSRcolor2[562]);
    BiasedRNG[893] = (LFSRcolor2[1255]&LFSRcolor2[973]&LFSRcolor2[1235]&LFSRcolor2[830]);
    BiasedRNG[894] = (LFSRcolor2[643]&LFSRcolor2[1012]&LFSRcolor2[587]&LFSRcolor2[178]);
    UnbiasedRNG[496] = LFSRcolor2[1242];
    UnbiasedRNG[497] = LFSRcolor2[1243];
    UnbiasedRNG[498] = LFSRcolor2[886];
    UnbiasedRNG[499] = LFSRcolor2[449];
    UnbiasedRNG[500] = LFSRcolor2[1271];
    UnbiasedRNG[501] = LFSRcolor2[1124];
    UnbiasedRNG[502] = LFSRcolor2[720];
    UnbiasedRNG[503] = LFSRcolor2[290];
    UnbiasedRNG[504] = LFSRcolor2[463];
    UnbiasedRNG[505] = LFSRcolor2[1228];
    UnbiasedRNG[506] = LFSRcolor2[1018];
    UnbiasedRNG[507] = LFSRcolor2[433];
    UnbiasedRNG[508] = LFSRcolor2[913];
    UnbiasedRNG[509] = LFSRcolor2[524];
    UnbiasedRNG[510] = LFSRcolor2[469];
    UnbiasedRNG[511] = LFSRcolor2[807];
    UnbiasedRNG[512] = LFSRcolor2[719];
    UnbiasedRNG[513] = LFSRcolor2[301];
    UnbiasedRNG[514] = LFSRcolor2[151];
    UnbiasedRNG[515] = LFSRcolor2[892];
    UnbiasedRNG[516] = LFSRcolor2[723];
    UnbiasedRNG[517] = LFSRcolor2[233];
    UnbiasedRNG[518] = LFSRcolor2[771];
    UnbiasedRNG[519] = LFSRcolor2[108];
    UnbiasedRNG[520] = LFSRcolor2[25];
    UnbiasedRNG[521] = LFSRcolor2[240];
    UnbiasedRNG[522] = LFSRcolor2[694];
    UnbiasedRNG[523] = LFSRcolor2[846];
    UnbiasedRNG[524] = LFSRcolor2[1006];
    UnbiasedRNG[525] = LFSRcolor2[1282];
    UnbiasedRNG[526] = LFSRcolor2[1118];
    UnbiasedRNG[527] = LFSRcolor2[1108];
    UnbiasedRNG[528] = LFSRcolor2[504];
    UnbiasedRNG[529] = LFSRcolor2[1072];
    UnbiasedRNG[530] = LFSRcolor2[415];
    UnbiasedRNG[531] = LFSRcolor2[1150];
    UnbiasedRNG[532] = LFSRcolor2[551];
    UnbiasedRNG[533] = LFSRcolor2[1131];
    UnbiasedRNG[534] = LFSRcolor2[272];
    UnbiasedRNG[535] = LFSRcolor2[684];
    UnbiasedRNG[536] = LFSRcolor2[155];
    UnbiasedRNG[537] = LFSRcolor2[200];
    UnbiasedRNG[538] = LFSRcolor2[1132];
    UnbiasedRNG[539] = LFSRcolor2[879];
    UnbiasedRNG[540] = LFSRcolor2[658];
    UnbiasedRNG[541] = LFSRcolor2[529];
    UnbiasedRNG[542] = LFSRcolor2[1223];
    UnbiasedRNG[543] = LFSRcolor2[595];
    UnbiasedRNG[544] = LFSRcolor2[85];
    UnbiasedRNG[545] = LFSRcolor2[655];
    UnbiasedRNG[546] = LFSRcolor2[158];
    UnbiasedRNG[547] = LFSRcolor2[929];
    UnbiasedRNG[548] = LFSRcolor2[596];
    UnbiasedRNG[549] = LFSRcolor2[8];
    UnbiasedRNG[550] = LFSRcolor2[111];
    UnbiasedRNG[551] = LFSRcolor2[974];
    UnbiasedRNG[552] = LFSRcolor2[874];
    UnbiasedRNG[553] = LFSRcolor2[512];
    UnbiasedRNG[554] = LFSRcolor2[357];
    UnbiasedRNG[555] = LFSRcolor2[735];
    UnbiasedRNG[556] = LFSRcolor2[956];
    UnbiasedRNG[557] = LFSRcolor2[391];
    UnbiasedRNG[558] = LFSRcolor2[183];
    UnbiasedRNG[559] = LFSRcolor2[260];
    UnbiasedRNG[560] = LFSRcolor2[317];
    UnbiasedRNG[561] = LFSRcolor2[1099];
    UnbiasedRNG[562] = LFSRcolor2[1134];
    UnbiasedRNG[563] = LFSRcolor2[370];
    UnbiasedRNG[564] = LFSRcolor2[953];
    UnbiasedRNG[565] = LFSRcolor2[81];
    UnbiasedRNG[566] = LFSRcolor2[465];
    UnbiasedRNG[567] = LFSRcolor2[1125];
    UnbiasedRNG[568] = LFSRcolor2[585];
    UnbiasedRNG[569] = LFSRcolor2[1261];
    UnbiasedRNG[570] = LFSRcolor2[541];
    UnbiasedRNG[571] = LFSRcolor2[518];
    UnbiasedRNG[572] = LFSRcolor2[261];
    UnbiasedRNG[573] = LFSRcolor2[628];
    UnbiasedRNG[574] = LFSRcolor2[749];
    UnbiasedRNG[575] = LFSRcolor2[884];
    UnbiasedRNG[576] = LFSRcolor2[808];
    UnbiasedRNG[577] = LFSRcolor2[303];
    UnbiasedRNG[578] = LFSRcolor2[954];
    UnbiasedRNG[579] = LFSRcolor2[459];
    UnbiasedRNG[580] = LFSRcolor2[297];
    UnbiasedRNG[581] = LFSRcolor2[96];
    UnbiasedRNG[582] = LFSRcolor2[638];
    UnbiasedRNG[583] = LFSRcolor2[101];
    UnbiasedRNG[584] = LFSRcolor2[123];
    UnbiasedRNG[585] = LFSRcolor2[1208];
    UnbiasedRNG[586] = LFSRcolor2[24];
    UnbiasedRNG[587] = LFSRcolor2[1053];
    UnbiasedRNG[588] = LFSRcolor2[352];
    UnbiasedRNG[589] = LFSRcolor2[505];
    UnbiasedRNG[590] = LFSRcolor2[567];
    UnbiasedRNG[591] = LFSRcolor2[315];
    UnbiasedRNG[592] = LFSRcolor2[1169];
    UnbiasedRNG[593] = LFSRcolor2[402];
    UnbiasedRNG[594] = LFSRcolor2[755];
    UnbiasedRNG[595] = LFSRcolor2[416];
    UnbiasedRNG[596] = LFSRcolor2[95];
    UnbiasedRNG[597] = LFSRcolor2[822];
    UnbiasedRNG[598] = LFSRcolor2[437];
    UnbiasedRNG[599] = LFSRcolor2[724];
    UnbiasedRNG[600] = LFSRcolor2[792];
    UnbiasedRNG[601] = LFSRcolor2[1224];
    UnbiasedRNG[602] = LFSRcolor2[53];
    UnbiasedRNG[603] = LFSRcolor2[709];
    UnbiasedRNG[604] = LFSRcolor2[911];
    UnbiasedRNG[605] = LFSRcolor2[1008];
    UnbiasedRNG[606] = LFSRcolor2[1269];
    UnbiasedRNG[607] = LFSRcolor2[837];
    UnbiasedRNG[608] = LFSRcolor2[1082];
    UnbiasedRNG[609] = LFSRcolor2[1070];
    UnbiasedRNG[610] = LFSRcolor2[209];
    UnbiasedRNG[611] = LFSRcolor2[1135];
    UnbiasedRNG[612] = LFSRcolor2[287];
    UnbiasedRNG[613] = LFSRcolor2[1211];
    UnbiasedRNG[614] = LFSRcolor2[487];
    UnbiasedRNG[615] = LFSRcolor2[778];
    UnbiasedRNG[616] = LFSRcolor2[1049];
    UnbiasedRNG[617] = LFSRcolor2[798];
    UnbiasedRNG[618] = LFSRcolor2[320];
    UnbiasedRNG[619] = LFSRcolor2[615];
    UnbiasedRNG[620] = LFSRcolor2[154];
    UnbiasedRNG[621] = LFSRcolor2[941];
    UnbiasedRNG[622] = LFSRcolor2[900];
    UnbiasedRNG[623] = LFSRcolor2[138];
    UnbiasedRNG[624] = LFSRcolor2[198];
    UnbiasedRNG[625] = LFSRcolor2[1191];
    UnbiasedRNG[626] = LFSRcolor2[358];
    UnbiasedRNG[627] = LFSRcolor2[1276];
    UnbiasedRNG[628] = LFSRcolor2[712];
    UnbiasedRNG[629] = LFSRcolor2[1078];
    UnbiasedRNG[630] = LFSRcolor2[369];
    UnbiasedRNG[631] = LFSRcolor2[631];
    UnbiasedRNG[632] = LFSRcolor2[794];
    UnbiasedRNG[633] = LFSRcolor2[78];
    UnbiasedRNG[634] = LFSRcolor2[179];
    UnbiasedRNG[635] = LFSRcolor2[10];
    UnbiasedRNG[636] = LFSRcolor2[506];
    UnbiasedRNG[637] = LFSRcolor2[842];
    UnbiasedRNG[638] = LFSRcolor2[922];
    UnbiasedRNG[639] = LFSRcolor2[979];
    UnbiasedRNG[640] = LFSRcolor2[1148];
    UnbiasedRNG[641] = LFSRcolor2[573];
    UnbiasedRNG[642] = LFSRcolor2[943];
    UnbiasedRNG[643] = LFSRcolor2[782];
    UnbiasedRNG[644] = LFSRcolor2[1266];
    UnbiasedRNG[645] = LFSRcolor2[867];
    UnbiasedRNG[646] = LFSRcolor2[1004];
    UnbiasedRNG[647] = LFSRcolor2[561];
    UnbiasedRNG[648] = LFSRcolor2[382];
    UnbiasedRNG[649] = LFSRcolor2[1250];
    UnbiasedRNG[650] = LFSRcolor2[208];
    UnbiasedRNG[651] = LFSRcolor2[152];
    UnbiasedRNG[652] = LFSRcolor2[926];
    UnbiasedRNG[653] = LFSRcolor2[283];
    UnbiasedRNG[654] = LFSRcolor2[445];
    UnbiasedRNG[655] = LFSRcolor2[553];
    UnbiasedRNG[656] = LFSRcolor2[435];
    UnbiasedRNG[657] = LFSRcolor2[1139];
    UnbiasedRNG[658] = LFSRcolor2[1159];
    UnbiasedRNG[659] = LFSRcolor2[1079];
    UnbiasedRNG[660] = LFSRcolor2[405];
    UnbiasedRNG[661] = LFSRcolor2[1032];
    UnbiasedRNG[662] = LFSRcolor2[45];
    UnbiasedRNG[663] = LFSRcolor2[202];
    UnbiasedRNG[664] = LFSRcolor2[765];
    UnbiasedRNG[665] = LFSRcolor2[670];
    UnbiasedRNG[666] = LFSRcolor2[946];
    UnbiasedRNG[667] = LFSRcolor2[626];
    UnbiasedRNG[668] = LFSRcolor2[150];
    UnbiasedRNG[669] = LFSRcolor2[1076];
    UnbiasedRNG[670] = LFSRcolor2[653];
    UnbiasedRNG[671] = LFSRcolor2[1096];
    UnbiasedRNG[672] = LFSRcolor2[458];
    UnbiasedRNG[673] = LFSRcolor2[920];
    UnbiasedRNG[674] = LFSRcolor2[821];
    UnbiasedRNG[675] = LFSRcolor2[343];
    UnbiasedRNG[676] = LFSRcolor2[1259];
    UnbiasedRNG[677] = LFSRcolor2[131];
    UnbiasedRNG[678] = LFSRcolor2[1110];
    UnbiasedRNG[679] = LFSRcolor2[768];
    UnbiasedRNG[680] = LFSRcolor2[848];
    UnbiasedRNG[681] = LFSRcolor2[455];
    UnbiasedRNG[682] = LFSRcolor2[345];
    UnbiasedRNG[683] = LFSRcolor2[1285];
    UnbiasedRNG[684] = LFSRcolor2[532];
    UnbiasedRNG[685] = LFSRcolor2[800];
    UnbiasedRNG[686] = LFSRcolor2[1141];
    UnbiasedRNG[687] = LFSRcolor2[894];
    UnbiasedRNG[688] = LFSRcolor2[277];
    UnbiasedRNG[689] = LFSRcolor2[1239];
    UnbiasedRNG[690] = LFSRcolor2[1043];
    UnbiasedRNG[691] = LFSRcolor2[1192];
    UnbiasedRNG[692] = LFSRcolor2[226];
    UnbiasedRNG[693] = LFSRcolor2[519];
    UnbiasedRNG[694] = LFSRcolor2[844];
    UnbiasedRNG[695] = LFSRcolor2[456];
    UnbiasedRNG[696] = LFSRcolor2[1146];
    UnbiasedRNG[697] = LFSRcolor2[1162];
    UnbiasedRNG[698] = LFSRcolor2[802];
    UnbiasedRNG[699] = LFSRcolor2[1113];
    UnbiasedRNG[700] = LFSRcolor2[305];
    UnbiasedRNG[701] = LFSRcolor2[338];
    UnbiasedRNG[702] = LFSRcolor2[482];
    UnbiasedRNG[703] = LFSRcolor2[952];
    UnbiasedRNG[704] = LFSRcolor2[851];
    UnbiasedRNG[705] = LFSRcolor2[526];
    UnbiasedRNG[706] = LFSRcolor2[234];
    UnbiasedRNG[707] = LFSRcolor2[795];
    UnbiasedRNG[708] = LFSRcolor2[173];
    UnbiasedRNG[709] = LFSRcolor2[293];
    UnbiasedRNG[710] = LFSRcolor2[539];
    UnbiasedRNG[711] = LFSRcolor2[547];
    UnbiasedRNG[712] = LFSRcolor2[1083];
    UnbiasedRNG[713] = LFSRcolor2[534];
    UnbiasedRNG[714] = LFSRcolor2[478];
    UnbiasedRNG[715] = LFSRcolor2[824];
    UnbiasedRNG[716] = LFSRcolor2[13];
    UnbiasedRNG[717] = LFSRcolor2[1022];
    UnbiasedRNG[718] = LFSRcolor2[852];
    UnbiasedRNG[719] = LFSRcolor2[1181];
    UnbiasedRNG[720] = LFSRcolor2[1105];
    UnbiasedRNG[721] = LFSRcolor2[319];
    UnbiasedRNG[722] = LFSRcolor2[412];
    UnbiasedRNG[723] = LFSRcolor2[1074];
    UnbiasedRNG[724] = LFSRcolor2[243];
    UnbiasedRNG[725] = LFSRcolor2[1256];
    UnbiasedRNG[726] = LFSRcolor2[201];
    UnbiasedRNG[727] = LFSRcolor2[219];
    UnbiasedRNG[728] = LFSRcolor2[1100];
    UnbiasedRNG[729] = LFSRcolor2[968];
    UnbiasedRNG[730] = LFSRcolor2[424];
    UnbiasedRNG[731] = LFSRcolor2[520];
    UnbiasedRNG[732] = LFSRcolor2[955];
    UnbiasedRNG[733] = LFSRcolor2[1095];
    UnbiasedRNG[734] = LFSRcolor2[399];
    UnbiasedRNG[735] = LFSRcolor2[902];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[736] = LFSRcolor3[98];
    UnbiasedRNG[737] = LFSRcolor3[222];
    UnbiasedRNG[738] = LFSRcolor3[136];
    UnbiasedRNG[739] = LFSRcolor3[227];
    UnbiasedRNG[740] = LFSRcolor3[213];
    UnbiasedRNG[741] = LFSRcolor3[78];
    UnbiasedRNG[742] = LFSRcolor3[65];
    UnbiasedRNG[743] = LFSRcolor3[7];
    UnbiasedRNG[744] = LFSRcolor3[101];
    UnbiasedRNG[745] = LFSRcolor3[191];
    UnbiasedRNG[746] = LFSRcolor3[148];
    UnbiasedRNG[747] = LFSRcolor3[87];
    UnbiasedRNG[748] = LFSRcolor3[44];
    UnbiasedRNG[749] = LFSRcolor3[119];
    UnbiasedRNG[750] = LFSRcolor3[114];
    UnbiasedRNG[751] = LFSRcolor3[153];
    UnbiasedRNG[752] = LFSRcolor3[107];
    UnbiasedRNG[753] = LFSRcolor3[167];
    UnbiasedRNG[754] = LFSRcolor3[219];
    UnbiasedRNG[755] = LFSRcolor3[59];
    UnbiasedRNG[756] = LFSRcolor3[58];
    UnbiasedRNG[757] = LFSRcolor3[46];
    UnbiasedRNG[758] = LFSRcolor3[109];
    UnbiasedRNG[759] = LFSRcolor3[174];
    UnbiasedRNG[760] = LFSRcolor3[193];
    UnbiasedRNG[761] = LFSRcolor3[125];
    UnbiasedRNG[762] = LFSRcolor3[57];
    UnbiasedRNG[763] = LFSRcolor3[75];
    UnbiasedRNG[764] = LFSRcolor3[223];
    UnbiasedRNG[765] = LFSRcolor3[34];
    UnbiasedRNG[766] = LFSRcolor3[228];
    UnbiasedRNG[767] = LFSRcolor3[175];
    UnbiasedRNG[768] = LFSRcolor3[38];
    UnbiasedRNG[769] = LFSRcolor3[16];
    UnbiasedRNG[770] = LFSRcolor3[37];
    UnbiasedRNG[771] = LFSRcolor3[19];
    UnbiasedRNG[772] = LFSRcolor3[189];
    UnbiasedRNG[773] = LFSRcolor3[50];
    UnbiasedRNG[774] = LFSRcolor3[200];
    UnbiasedRNG[775] = LFSRcolor3[225];
    UnbiasedRNG[776] = LFSRcolor3[195];
    UnbiasedRNG[777] = LFSRcolor3[212];
    UnbiasedRNG[778] = LFSRcolor3[90];
    UnbiasedRNG[779] = LFSRcolor3[72];
    UnbiasedRNG[780] = LFSRcolor3[33];
    UnbiasedRNG[781] = LFSRcolor3[24];
    UnbiasedRNG[782] = LFSRcolor3[204];
    UnbiasedRNG[783] = LFSRcolor3[207];
    UnbiasedRNG[784] = LFSRcolor3[142];
    UnbiasedRNG[785] = LFSRcolor3[91];
    UnbiasedRNG[786] = LFSRcolor3[10];
    UnbiasedRNG[787] = LFSRcolor3[56];
    UnbiasedRNG[788] = LFSRcolor3[187];
    UnbiasedRNG[789] = LFSRcolor3[66];
    UnbiasedRNG[790] = LFSRcolor3[103];
    UnbiasedRNG[791] = LFSRcolor3[42];
    UnbiasedRNG[792] = LFSRcolor3[181];
    UnbiasedRNG[793] = LFSRcolor3[12];
    UnbiasedRNG[794] = LFSRcolor3[81];
    UnbiasedRNG[795] = LFSRcolor3[94];
    UnbiasedRNG[796] = LFSRcolor3[144];
    UnbiasedRNG[797] = LFSRcolor3[76];
    UnbiasedRNG[798] = LFSRcolor3[89];
    UnbiasedRNG[799] = LFSRcolor3[128];
    UnbiasedRNG[800] = LFSRcolor3[179];
    UnbiasedRNG[801] = LFSRcolor3[102];
    UnbiasedRNG[802] = LFSRcolor3[84];
    UnbiasedRNG[803] = LFSRcolor3[220];
    UnbiasedRNG[804] = LFSRcolor3[45];
    UnbiasedRNG[805] = LFSRcolor3[40];
    UnbiasedRNG[806] = LFSRcolor3[5];
    UnbiasedRNG[807] = LFSRcolor3[202];
    UnbiasedRNG[808] = LFSRcolor3[18];
    UnbiasedRNG[809] = LFSRcolor3[192];
    UnbiasedRNG[810] = LFSRcolor3[216];
    UnbiasedRNG[811] = LFSRcolor3[182];
    UnbiasedRNG[812] = LFSRcolor3[173];
    UnbiasedRNG[813] = LFSRcolor3[218];
    UnbiasedRNG[814] = LFSRcolor3[158];
    UnbiasedRNG[815] = LFSRcolor3[138];
    UnbiasedRNG[816] = LFSRcolor3[29];
    UnbiasedRNG[817] = LFSRcolor3[137];
    UnbiasedRNG[818] = LFSRcolor3[100];
    UnbiasedRNG[819] = LFSRcolor3[20];
    UnbiasedRNG[820] = LFSRcolor3[130];
    UnbiasedRNG[821] = LFSRcolor3[77];
    UnbiasedRNG[822] = LFSRcolor3[74];
    UnbiasedRNG[823] = LFSRcolor3[224];
    UnbiasedRNG[824] = LFSRcolor3[31];
    UnbiasedRNG[825] = LFSRcolor3[147];
    UnbiasedRNG[826] = LFSRcolor3[118];
    UnbiasedRNG[827] = LFSRcolor3[39];
    UnbiasedRNG[828] = LFSRcolor3[104];
    UnbiasedRNG[829] = LFSRcolor3[61];
    UnbiasedRNG[830] = LFSRcolor3[55];
    UnbiasedRNG[831] = LFSRcolor3[53];
    UnbiasedRNG[832] = LFSRcolor3[30];
    UnbiasedRNG[833] = LFSRcolor3[140];
    UnbiasedRNG[834] = LFSRcolor3[126];
    UnbiasedRNG[835] = LFSRcolor3[154];
    UnbiasedRNG[836] = LFSRcolor3[83];
    UnbiasedRNG[837] = LFSRcolor3[47];
    UnbiasedRNG[838] = LFSRcolor3[35];
    UnbiasedRNG[839] = LFSRcolor3[95];
    UnbiasedRNG[840] = LFSRcolor3[96];
    UnbiasedRNG[841] = LFSRcolor3[129];
    UnbiasedRNG[842] = LFSRcolor3[68];
    UnbiasedRNG[843] = LFSRcolor3[106];
    UnbiasedRNG[844] = LFSRcolor3[1];
    UnbiasedRNG[845] = LFSRcolor3[141];
    UnbiasedRNG[846] = LFSRcolor3[97];
    UnbiasedRNG[847] = LFSRcolor3[64];
    UnbiasedRNG[848] = LFSRcolor3[26];
    UnbiasedRNG[849] = LFSRcolor3[215];
    UnbiasedRNG[850] = LFSRcolor3[111];
    UnbiasedRNG[851] = LFSRcolor3[14];
    UnbiasedRNG[852] = LFSRcolor3[2];
    UnbiasedRNG[853] = LFSRcolor3[197];
    UnbiasedRNG[854] = LFSRcolor3[124];
    UnbiasedRNG[855] = LFSRcolor3[199];
    UnbiasedRNG[856] = LFSRcolor3[188];
    UnbiasedRNG[857] = LFSRcolor3[110];
    UnbiasedRNG[858] = LFSRcolor3[108];
    UnbiasedRNG[859] = LFSRcolor3[41];
    UnbiasedRNG[860] = LFSRcolor3[152];
    UnbiasedRNG[861] = LFSRcolor3[22];
    UnbiasedRNG[862] = LFSRcolor3[205];
    UnbiasedRNG[863] = LFSRcolor3[25];
    UnbiasedRNG[864] = LFSRcolor3[122];
    UnbiasedRNG[865] = LFSRcolor3[11];
    UnbiasedRNG[866] = LFSRcolor3[162];
    UnbiasedRNG[867] = LFSRcolor3[209];
    UnbiasedRNG[868] = LFSRcolor3[139];
    UnbiasedRNG[869] = LFSRcolor3[121];
    UnbiasedRNG[870] = LFSRcolor3[120];
    UnbiasedRNG[871] = LFSRcolor3[0];
    UnbiasedRNG[872] = LFSRcolor3[36];
    UnbiasedRNG[873] = LFSRcolor3[171];
    UnbiasedRNG[874] = LFSRcolor3[164];
    UnbiasedRNG[875] = LFSRcolor3[166];
    UnbiasedRNG[876] = LFSRcolor3[113];
    UnbiasedRNG[877] = LFSRcolor3[79];
    UnbiasedRNG[878] = LFSRcolor3[105];
    UnbiasedRNG[879] = LFSRcolor3[85];
    UnbiasedRNG[880] = LFSRcolor3[229];
    UnbiasedRNG[881] = LFSRcolor3[63];
    UnbiasedRNG[882] = LFSRcolor3[206];
    UnbiasedRNG[883] = LFSRcolor3[211];
    UnbiasedRNG[884] = LFSRcolor3[3];
    UnbiasedRNG[885] = LFSRcolor3[214];
    UnbiasedRNG[886] = LFSRcolor3[184];
    UnbiasedRNG[887] = LFSRcolor3[201];
    UnbiasedRNG[888] = LFSRcolor3[17];
    UnbiasedRNG[889] = LFSRcolor3[9];
    UnbiasedRNG[890] = LFSRcolor3[69];
    UnbiasedRNG[891] = LFSRcolor3[92];
    UnbiasedRNG[892] = LFSRcolor3[132];
    UnbiasedRNG[893] = LFSRcolor3[198];
    UnbiasedRNG[894] = LFSRcolor3[135];
    UnbiasedRNG[895] = LFSRcolor3[80];
    UnbiasedRNG[896] = LFSRcolor3[60];
    UnbiasedRNG[897] = LFSRcolor3[51];
    UnbiasedRNG[898] = LFSRcolor3[62];
    UnbiasedRNG[899] = LFSRcolor3[86];
    UnbiasedRNG[900] = LFSRcolor3[13];
    UnbiasedRNG[901] = LFSRcolor3[226];
    UnbiasedRNG[902] = LFSRcolor3[71];
    UnbiasedRNG[903] = LFSRcolor3[208];
    UnbiasedRNG[904] = LFSRcolor3[177];
    UnbiasedRNG[905] = LFSRcolor3[165];
    UnbiasedRNG[906] = LFSRcolor3[159];
    UnbiasedRNG[907] = LFSRcolor3[49];
    UnbiasedRNG[908] = LFSRcolor3[67];
    UnbiasedRNG[909] = LFSRcolor3[196];
    UnbiasedRNG[910] = LFSRcolor3[190];
    UnbiasedRNG[911] = LFSRcolor3[99];
    UnbiasedRNG[912] = LFSRcolor3[169];
    UnbiasedRNG[913] = LFSRcolor3[28];
    UnbiasedRNG[914] = LFSRcolor3[210];
    UnbiasedRNG[915] = LFSRcolor3[117];
    UnbiasedRNG[916] = LFSRcolor3[134];
    UnbiasedRNG[917] = LFSRcolor3[43];
    UnbiasedRNG[918] = LFSRcolor3[163];
    UnbiasedRNG[919] = LFSRcolor3[143];
    UnbiasedRNG[920] = LFSRcolor3[4];
    UnbiasedRNG[921] = LFSRcolor3[203];
    UnbiasedRNG[922] = LFSRcolor3[23];
    UnbiasedRNG[923] = LFSRcolor3[185];
    UnbiasedRNG[924] = LFSRcolor3[32];
    UnbiasedRNG[925] = LFSRcolor3[168];
    UnbiasedRNG[926] = LFSRcolor3[70];
    UnbiasedRNG[927] = LFSRcolor3[172];
    UnbiasedRNG[928] = LFSRcolor3[127];
    UnbiasedRNG[929] = LFSRcolor3[21];
    UnbiasedRNG[930] = LFSRcolor3[123];
    UnbiasedRNG[931] = LFSRcolor3[112];
    UnbiasedRNG[932] = LFSRcolor3[160];
    UnbiasedRNG[933] = LFSRcolor3[157];
    UnbiasedRNG[934] = LFSRcolor3[27];
    UnbiasedRNG[935] = LFSRcolor3[48];
    UnbiasedRNG[936] = LFSRcolor3[115];
    UnbiasedRNG[937] = LFSRcolor3[93];
    UnbiasedRNG[938] = LFSRcolor3[131];
    UnbiasedRNG[939] = LFSRcolor3[221];
    UnbiasedRNG[940] = LFSRcolor3[161];
    UnbiasedRNG[941] = LFSRcolor3[73];
    UnbiasedRNG[942] = LFSRcolor3[133];
    UnbiasedRNG[943] = LFSRcolor3[149];
    UnbiasedRNG[944] = LFSRcolor3[52];
    UnbiasedRNG[945] = LFSRcolor3[155];
end

always @(posedge color3_clk) begin
    BiasedRNG[895] = (LFSRcolor4[947]&LFSRcolor4[390]&LFSRcolor4[395]&LFSRcolor4[463]);
    BiasedRNG[896] = (LFSRcolor4[937]&LFSRcolor4[832]&LFSRcolor4[10]&LFSRcolor4[870]);
    BiasedRNG[897] = (LFSRcolor4[956]&LFSRcolor4[730]&LFSRcolor4[111]&LFSRcolor4[479]);
    BiasedRNG[898] = (LFSRcolor4[914]&LFSRcolor4[411]&LFSRcolor4[223]&LFSRcolor4[170]);
    BiasedRNG[899] = (LFSRcolor4[360]&LFSRcolor4[639]&LFSRcolor4[873]&LFSRcolor4[869]);
    BiasedRNG[900] = (LFSRcolor4[810]&LFSRcolor4[322]&LFSRcolor4[534]&LFSRcolor4[9]);
    BiasedRNG[901] = (LFSRcolor4[341]&LFSRcolor4[568]&LFSRcolor4[650]&LFSRcolor4[835]);
    BiasedRNG[902] = (LFSRcolor4[583]&LFSRcolor4[124]&LFSRcolor4[63]&LFSRcolor4[321]);
    BiasedRNG[903] = (LFSRcolor4[110]&LFSRcolor4[228]&LFSRcolor4[447]&LFSRcolor4[156]);
    BiasedRNG[904] = (LFSRcolor4[216]&LFSRcolor4[830]&LFSRcolor4[964]&LFSRcolor4[824]);
    BiasedRNG[905] = (LFSRcolor4[593]&LFSRcolor4[30]&LFSRcolor4[191]&LFSRcolor4[459]);
    BiasedRNG[906] = (LFSRcolor4[405]&LFSRcolor4[95]&LFSRcolor4[582]&LFSRcolor4[726]);
    BiasedRNG[907] = (LFSRcolor4[940]&LFSRcolor4[22]&LFSRcolor4[893]&LFSRcolor4[843]);
    BiasedRNG[908] = (LFSRcolor4[778]&LFSRcolor4[508]&LFSRcolor4[884]&LFSRcolor4[437]);
    BiasedRNG[909] = (LFSRcolor4[712]&LFSRcolor4[241]&LFSRcolor4[762]&LFSRcolor4[190]);
    BiasedRNG[910] = (LFSRcolor4[883]&LFSRcolor4[701]&LFSRcolor4[81]&LFSRcolor4[755]);
    BiasedRNG[911] = (LFSRcolor4[444]&LFSRcolor4[649]&LFSRcolor4[692]&LFSRcolor4[652]);
    BiasedRNG[912] = (LFSRcolor4[496]&LFSRcolor4[517]&LFSRcolor4[441]&LFSRcolor4[26]);
    BiasedRNG[913] = (LFSRcolor4[916]&LFSRcolor4[330]&LFSRcolor4[92]&LFSRcolor4[436]);
    BiasedRNG[914] = (LFSRcolor4[754]&LFSRcolor4[766]&LFSRcolor4[244]&LFSRcolor4[335]);
    BiasedRNG[915] = (LFSRcolor4[901]&LFSRcolor4[167]&LFSRcolor4[954]&LFSRcolor4[4]);
    BiasedRNG[916] = (LFSRcolor4[691]&LFSRcolor4[570]&LFSRcolor4[20]&LFSRcolor4[263]);
    BiasedRNG[917] = (LFSRcolor4[819]&LFSRcolor4[461]&LFSRcolor4[779]&LFSRcolor4[688]);
    BiasedRNG[918] = (LFSRcolor4[122]&LFSRcolor4[165]&LFSRcolor4[681]&LFSRcolor4[262]);
    BiasedRNG[919] = (LFSRcolor4[56]&LFSRcolor4[732]&LFSRcolor4[818]&LFSRcolor4[806]);
    BiasedRNG[920] = (LFSRcolor4[229]&LFSRcolor4[339]&LFSRcolor4[47]&LFSRcolor4[592]);
    BiasedRNG[921] = (LFSRcolor4[708]&LFSRcolor4[101]&LFSRcolor4[860]&LFSRcolor4[952]);
    BiasedRNG[922] = (LFSRcolor4[604]&LFSRcolor4[224]&LFSRcolor4[199]&LFSRcolor4[453]);
    BiasedRNG[923] = (LFSRcolor4[451]&LFSRcolor4[38]&LFSRcolor4[306]&LFSRcolor4[72]);
    BiasedRNG[924] = (LFSRcolor4[717]&LFSRcolor4[389]&LFSRcolor4[939]&LFSRcolor4[410]);
    BiasedRNG[925] = (LFSRcolor4[157]&LFSRcolor4[827]&LFSRcolor4[369]&LFSRcolor4[162]);
    BiasedRNG[926] = (LFSRcolor4[529]&LFSRcolor4[15]&LFSRcolor4[235]&LFSRcolor4[640]);
    BiasedRNG[927] = (LFSRcolor4[497]&LFSRcolor4[115]&LFSRcolor4[474]&LFSRcolor4[426]);
    BiasedRNG[928] = (LFSRcolor4[696]&LFSRcolor4[924]&LFSRcolor4[678]&LFSRcolor4[349]);
    BiasedRNG[929] = (LFSRcolor4[23]&LFSRcolor4[19]&LFSRcolor4[350]&LFSRcolor4[328]);
    BiasedRNG[930] = (LFSRcolor4[288]&LFSRcolor4[268]&LFSRcolor4[527]&LFSRcolor4[138]);
    BiasedRNG[931] = (LFSRcolor4[176]&LFSRcolor4[886]&LFSRcolor4[67]&LFSRcolor4[377]);
    BiasedRNG[932] = (LFSRcolor4[14]&LFSRcolor4[599]&LFSRcolor4[727]&LFSRcolor4[890]);
    BiasedRNG[933] = (LFSRcolor4[514]&LFSRcolor4[951]&LFSRcolor4[336]&LFSRcolor4[368]);
    BiasedRNG[934] = (LFSRcolor4[233]&LFSRcolor4[928]&LFSRcolor4[273]&LFSRcolor4[129]);
    BiasedRNG[935] = (LFSRcolor4[710]&LFSRcolor4[677]&LFSRcolor4[629]&LFSRcolor4[292]);
    BiasedRNG[936] = (LFSRcolor4[251]&LFSRcolor4[934]&LFSRcolor4[442]&LFSRcolor4[865]);
    BiasedRNG[937] = (LFSRcolor4[892]&LFSRcolor4[948]&LFSRcolor4[551]&LFSRcolor4[910]);
    BiasedRNG[938] = (LFSRcolor4[185]&LFSRcolor4[700]&LFSRcolor4[345]&LFSRcolor4[329]);
    BiasedRNG[939] = (LFSRcolor4[443]&LFSRcolor4[800]&LFSRcolor4[499]&LFSRcolor4[55]);
    BiasedRNG[940] = (LFSRcolor4[254]&LFSRcolor4[707]&LFSRcolor4[607]&LFSRcolor4[379]);
    BiasedRNG[941] = (LFSRcolor4[135]&LFSRcolor4[693]&LFSRcolor4[638]&LFSRcolor4[378]);
    BiasedRNG[942] = (LFSRcolor4[62]&LFSRcolor4[366]&LFSRcolor4[417]&LFSRcolor4[673]);
    BiasedRNG[943] = (LFSRcolor4[32]&LFSRcolor4[46]&LFSRcolor4[470]&LFSRcolor4[658]);
    BiasedRNG[944] = (LFSRcolor4[578]&LFSRcolor4[687]&LFSRcolor4[187]&LFSRcolor4[724]);
    BiasedRNG[945] = (LFSRcolor4[194]&LFSRcolor4[36]&LFSRcolor4[58]&LFSRcolor4[746]);
    BiasedRNG[946] = (LFSRcolor4[793]&LFSRcolor4[276]&LFSRcolor4[838]&LFSRcolor4[207]);
    BiasedRNG[947] = (LFSRcolor4[949]&LFSRcolor4[872]&LFSRcolor4[236]&LFSRcolor4[795]);
    BiasedRNG[948] = (LFSRcolor4[822]&LFSRcolor4[857]&LFSRcolor4[507]&LFSRcolor4[396]);
    BiasedRNG[949] = (LFSRcolor4[408]&LFSRcolor4[772]&LFSRcolor4[927]&LFSRcolor4[154]);
    BiasedRNG[950] = (LFSRcolor4[178]&LFSRcolor4[504]&LFSRcolor4[622]&LFSRcolor4[674]);
    BiasedRNG[951] = (LFSRcolor4[941]&LFSRcolor4[680]&LFSRcolor4[68]&LFSRcolor4[13]);
    BiasedRNG[952] = (LFSRcolor4[114]&LFSRcolor4[439]&LFSRcolor4[850]&LFSRcolor4[909]);
    BiasedRNG[953] = (LFSRcolor4[289]&LFSRcolor4[773]&LFSRcolor4[323]&LFSRcolor4[149]);
    BiasedRNG[954] = (LFSRcolor4[340]&LFSRcolor4[433]&LFSRcolor4[158]&LFSRcolor4[8]);
    BiasedRNG[955] = (LFSRcolor4[749]&LFSRcolor4[455]&LFSRcolor4[888]&LFSRcolor4[581]);
    BiasedRNG[956] = (LFSRcolor4[509]&LFSRcolor4[282]&LFSRcolor4[896]&LFSRcolor4[719]);
    BiasedRNG[957] = (LFSRcolor4[225]&LFSRcolor4[70]&LFSRcolor4[342]&LFSRcolor4[478]);
    BiasedRNG[958] = (LFSRcolor4[816]&LFSRcolor4[356]&LFSRcolor4[89]&LFSRcolor4[334]);
    BiasedRNG[959] = (LFSRcolor4[314]&LFSRcolor4[57]&LFSRcolor4[351]&LFSRcolor4[784]);
    BiasedRNG[960] = (LFSRcolor4[663]&LFSRcolor4[78]&LFSRcolor4[936]&LFSRcolor4[143]);
    BiasedRNG[961] = (LFSRcolor4[204]&LFSRcolor4[249]&LFSRcolor4[257]&LFSRcolor4[12]);
    BiasedRNG[962] = (LFSRcolor4[813]&LFSRcolor4[697]&LFSRcolor4[247]&LFSRcolor4[875]);
    BiasedRNG[963] = (LFSRcolor4[905]&LFSRcolor4[938]&LFSRcolor4[614]&LFSRcolor4[840]);
    BiasedRNG[964] = (LFSRcolor4[293]&LFSRcolor4[16]&LFSRcolor4[132]&LFSRcolor4[41]);
    BiasedRNG[965] = (LFSRcolor4[213]&LFSRcolor4[29]&LFSRcolor4[242]&LFSRcolor4[182]);
    BiasedRNG[966] = (LFSRcolor4[112]&LFSRcolor4[108]&LFSRcolor4[370]&LFSRcolor4[373]);
    BiasedRNG[967] = (LFSRcolor4[703]&LFSRcolor4[344]&LFSRcolor4[298]&LFSRcolor4[831]);
    BiasedRNG[968] = (LFSRcolor4[105]&LFSRcolor4[492]&LFSRcolor4[706]&LFSRcolor4[828]);
    BiasedRNG[969] = (LFSRcolor4[98]&LFSRcolor4[829]&LFSRcolor4[610]&LFSRcolor4[926]);
    BiasedRNG[970] = (LFSRcolor4[522]&LFSRcolor4[902]&LFSRcolor4[502]&LFSRcolor4[577]);
    BiasedRNG[971] = (LFSRcolor4[222]&LFSRcolor4[300]&LFSRcolor4[603]&LFSRcolor4[163]);
    BiasedRNG[972] = (LFSRcolor4[761]&LFSRcolor4[372]&LFSRcolor4[595]&LFSRcolor4[611]);
    BiasedRNG[973] = (LFSRcolor4[716]&LFSRcolor4[523]&LFSRcolor4[33]&LFSRcolor4[343]);
    BiasedRNG[974] = (LFSRcolor4[547]&LFSRcolor4[807]&LFSRcolor4[31]&LFSRcolor4[432]);
    BiasedRNG[975] = (LFSRcolor4[375]&LFSRcolor4[51]&LFSRcolor4[747]&LFSRcolor4[598]);
    BiasedRNG[976] = (LFSRcolor4[123]&LFSRcolor4[711]&LFSRcolor4[179]&LFSRcolor4[383]);
    BiasedRNG[977] = (LFSRcolor4[572]&LFSRcolor4[198]&LFSRcolor4[933]&LFSRcolor4[615]);
    BiasedRNG[978] = (LFSRcolor4[554]&LFSRcolor4[34]&LFSRcolor4[450]&LFSRcolor4[590]);
    BiasedRNG[979] = (LFSRcolor4[296]&LFSRcolor4[963]&LFSRcolor4[695]&LFSRcolor4[799]);
    BiasedRNG[980] = (LFSRcolor4[161]&LFSRcolor4[391]&LFSRcolor4[906]&LFSRcolor4[526]);
    BiasedRNG[981] = (LFSRcolor4[208]&LFSRcolor4[17]&LFSRcolor4[260]&LFSRcolor4[454]);
    BiasedRNG[982] = (LFSRcolor4[671]&LFSRcolor4[295]&LFSRcolor4[155]&LFSRcolor4[505]);
    BiasedRNG[983] = (LFSRcolor4[218]&LFSRcolor4[69]&LFSRcolor4[291]&LFSRcolor4[768]);
    BiasedRNG[984] = (LFSRcolor4[102]&LFSRcolor4[586]&LFSRcolor4[601]&LFSRcolor4[558]);
    BiasedRNG[985] = (LFSRcolor4[355]&LFSRcolor4[550]&LFSRcolor4[548]&LFSRcolor4[180]);
    BiasedRNG[986] = (LFSRcolor4[245]&LFSRcolor4[929]&LFSRcolor4[43]&LFSRcolor4[556]);
    BiasedRNG[987] = (LFSRcolor4[414]&LFSRcolor4[608]&LFSRcolor4[283]&LFSRcolor4[209]);
    BiasedRNG[988] = (LFSRcolor4[944]&LFSRcolor4[729]&LFSRcolor4[777]&LFSRcolor4[641]);
    BiasedRNG[989] = (LFSRcolor4[506]&LFSRcolor4[6]&LFSRcolor4[647]&LFSRcolor4[636]);
    BiasedRNG[990] = (LFSRcolor4[643]&LFSRcolor4[513]&LFSRcolor4[3]&LFSRcolor4[214]);
    BiasedRNG[991] = (LFSRcolor4[915]&LFSRcolor4[753]&LFSRcolor4[393]&LFSRcolor4[862]);
    BiasedRNG[992] = (LFSRcolor4[544]&LFSRcolor4[400]&LFSRcolor4[965]&LFSRcolor4[859]);
    BiasedRNG[993] = (LFSRcolor4[270]&LFSRcolor4[718]&LFSRcolor4[304]&LFSRcolor4[955]);
    BiasedRNG[994] = (LFSRcolor4[620]&LFSRcolor4[256]&LFSRcolor4[798]&LFSRcolor4[305]);
    BiasedRNG[995] = (LFSRcolor4[169]&LFSRcolor4[477]&LFSRcolor4[734]&LFSRcolor4[324]);
    BiasedRNG[996] = (LFSRcolor4[467]&LFSRcolor4[855]&LFSRcolor4[142]&LFSRcolor4[694]);
    BiasedRNG[997] = (LFSRcolor4[634]&LFSRcolor4[174]&LFSRcolor4[175]&LFSRcolor4[679]);
    BiasedRNG[998] = (LFSRcolor4[488]&LFSRcolor4[404]&LFSRcolor4[118]&LFSRcolor4[460]);
    BiasedRNG[999] = (LFSRcolor4[381]&LFSRcolor4[486]&LFSRcolor4[531]&LFSRcolor4[667]);
    BiasedRNG[1000] = (LFSRcolor4[532]&LFSRcolor4[957]&LFSRcolor4[637]&LFSRcolor4[520]);
    BiasedRNG[1001] = (LFSRcolor4[656]&LFSRcolor4[672]&LFSRcolor4[2]&LFSRcolor4[243]);
    BiasedRNG[1002] = (LFSRcolor4[325]&LFSRcolor4[481]&LFSRcolor4[670]&LFSRcolor4[212]);
    BiasedRNG[1003] = (LFSRcolor4[406]&LFSRcolor4[74]&LFSRcolor4[277]&LFSRcolor4[589]);
    BiasedRNG[1004] = (LFSRcolor4[219]&LFSRcolor4[485]&LFSRcolor4[518]&LFSRcolor4[200]);
    BiasedRNG[1005] = (LFSRcolor4[401]&LFSRcolor4[125]&LFSRcolor4[53]&LFSRcolor4[958]);
    BiasedRNG[1006] = (LFSRcolor4[37]&LFSRcolor4[736]&LFSRcolor4[299]&LFSRcolor4[146]);
    BiasedRNG[1007] = (LFSRcolor4[713]&LFSRcolor4[269]&LFSRcolor4[895]&LFSRcolor4[327]);
    BiasedRNG[1008] = (LFSRcolor4[87]&LFSRcolor4[274]&LFSRcolor4[794]&LFSRcolor4[600]);
    BiasedRNG[1009] = (LFSRcolor4[445]&LFSRcolor4[184]&LFSRcolor4[782]&LFSRcolor4[817]);
    BiasedRNG[1010] = (LFSRcolor4[261]&LFSRcolor4[99]&LFSRcolor4[85]&LFSRcolor4[743]);
    BiasedRNG[1011] = (LFSRcolor4[606]&LFSRcolor4[624]&LFSRcolor4[494]&LFSRcolor4[424]);
    BiasedRNG[1012] = (LFSRcolor4[452]&LFSRcolor4[503]&LFSRcolor4[684]&LFSRcolor4[538]);
    BiasedRNG[1013] = (LFSRcolor4[921]&LFSRcolor4[448]&LFSRcolor4[318]&LFSRcolor4[868]);
    BiasedRNG[1014] = (LFSRcolor4[846]&LFSRcolor4[894]&LFSRcolor4[833]&LFSRcolor4[919]);
    BiasedRNG[1015] = (LFSRcolor4[358]&LFSRcolor4[484]&LFSRcolor4[286]&LFSRcolor4[382]);
    BiasedRNG[1016] = (LFSRcolor4[310]&LFSRcolor4[685]&LFSRcolor4[430]&LFSRcolor4[533]);
    BiasedRNG[1017] = (LFSRcolor4[466]&LFSRcolor4[230]&LFSRcolor4[899]&LFSRcolor4[758]);
    BiasedRNG[1018] = (LFSRcolor4[246]&LFSRcolor4[0]&LFSRcolor4[177]&LFSRcolor4[765]);
    BiasedRNG[1019] = (LFSRcolor4[648]&LFSRcolor4[252]&LFSRcolor4[315]&LFSRcolor4[723]);
    BiasedRNG[1020] = (LFSRcolor4[75]&LFSRcolor4[848]&LFSRcolor4[745]&LFSRcolor4[932]);
    BiasedRNG[1021] = (LFSRcolor4[585]&LFSRcolor4[646]&LFSRcolor4[472]&LFSRcolor4[837]);
    BiasedRNG[1022] = (LFSRcolor4[258]&LFSRcolor4[618]&LFSRcolor4[561]&LFSRcolor4[740]);
    BiasedRNG[1023] = (LFSRcolor4[419]&LFSRcolor4[853]&LFSRcolor4[669]&LFSRcolor4[211]);
    BiasedRNG[1024] = (LFSRcolor4[801]&LFSRcolor4[97]&LFSRcolor4[804]&LFSRcolor4[387]);
    BiasedRNG[1025] = (LFSRcolor4[565]&LFSRcolor4[930]&LFSRcolor4[71]&LFSRcolor4[704]);
    BiasedRNG[1026] = (LFSRcolor4[642]&LFSRcolor4[823]&LFSRcolor4[130]&LFSRcolor4[312]);
    BiasedRNG[1027] = (LFSRcolor4[374]&LFSRcolor4[352]&LFSRcolor4[197]&LFSRcolor4[491]);
    BiasedRNG[1028] = (LFSRcolor4[202]&LFSRcolor4[519]&LFSRcolor4[21]&LFSRcolor4[844]);
    BiasedRNG[1029] = (LFSRcolor4[525]&LFSRcolor4[280]&LFSRcolor4[420]&LFSRcolor4[511]);
    BiasedRNG[1030] = (LFSRcolor4[465]&LFSRcolor4[221]&LFSRcolor4[512]&LFSRcolor4[172]);
    BiasedRNG[1031] = (LFSRcolor4[597]&LFSRcolor4[756]&LFSRcolor4[449]&LFSRcolor4[297]);
    BiasedRNG[1032] = (LFSRcolor4[540]&LFSRcolor4[675]&LFSRcolor4[912]&LFSRcolor4[398]);
    BiasedRNG[1033] = (LFSRcolor4[521]&LFSRcolor4[866]&LFSRcolor4[690]&LFSRcolor4[171]);
    BiasedRNG[1034] = (LFSRcolor4[215]&LFSRcolor4[423]&LFSRcolor4[836]&LFSRcolor4[66]);
    BiasedRNG[1035] = (LFSRcolor4[7]&LFSRcolor4[279]&LFSRcolor4[845]&LFSRcolor4[84]);
    BiasedRNG[1036] = (LFSRcolor4[594]&LFSRcolor4[127]&LFSRcolor4[148]&LFSRcolor4[962]);
    BiasedRNG[1037] = (LFSRcolor4[752]&LFSRcolor4[841]&LFSRcolor4[537]&LFSRcolor4[490]);
    BiasedRNG[1038] = (LFSRcolor4[421]&LFSRcolor4[76]&LFSRcolor4[588]&LFSRcolor4[90]);
    BiasedRNG[1039] = (LFSRcolor4[319]&LFSRcolor4[546]&LFSRcolor4[337]&LFSRcolor4[316]);
    BiasedRNG[1040] = (LFSRcolor4[116]&LFSRcolor4[210]&LFSRcolor4[741]&LFSRcolor4[495]);
    BiasedRNG[1041] = (LFSRcolor4[126]&LFSRcolor4[721]&LFSRcolor4[560]&LFSRcolor4[945]);
    BiasedRNG[1042] = (LFSRcolor4[591]&LFSRcolor4[120]&LFSRcolor4[168]&LFSRcolor4[635]);
    BiasedRNG[1043] = (LFSRcolor4[192]&LFSRcolor4[498]&LFSRcolor4[767]&LFSRcolor4[134]);
    BiasedRNG[1044] = (LFSRcolor4[418]&LFSRcolor4[602]&LFSRcolor4[294]&LFSRcolor4[307]);
    BiasedRNG[1045] = (LFSRcolor4[931]&LFSRcolor4[737]&LFSRcolor4[891]&LFSRcolor4[858]);
    BiasedRNG[1046] = (LFSRcolor4[5]&LFSRcolor4[259]&LFSRcolor4[774]&LFSRcolor4[771]);
    BiasedRNG[1047] = (LFSRcolor4[666]&LFSRcolor4[240]&LFSRcolor4[808]&LFSRcolor4[960]);
    BiasedRNG[1048] = (LFSRcolor4[365]&LFSRcolor4[619]&LFSRcolor4[141]&LFSRcolor4[332]);
    BiasedRNG[1049] = (LFSRcolor4[877]&LFSRcolor4[173]&LFSRcolor4[882]&LFSRcolor4[186]);
    BiasedRNG[1050] = (LFSRcolor4[482]&LFSRcolor4[409]&LFSRcolor4[922]&LFSRcolor4[128]);
    BiasedRNG[1051] = (LFSRcolor4[535]&LFSRcolor4[117]&LFSRcolor4[119]&LFSRcolor4[789]);
    BiasedRNG[1052] = (LFSRcolor4[248]&LFSRcolor4[796]&LFSRcolor4[867]&LFSRcolor4[907]);
    BiasedRNG[1053] = (LFSRcolor4[109]&LFSRcolor4[338]&LFSRcolor4[317]&LFSRcolor4[787]);
    BiasedRNG[1054] = (LFSRcolor4[255]&LFSRcolor4[415]&LFSRcolor4[407]&LFSRcolor4[303]);
    BiasedRNG[1055] = (LFSRcolor4[399]&LFSRcolor4[275]&LFSRcolor4[786]&LFSRcolor4[348]);
    BiasedRNG[1056] = (LFSRcolor4[744]&LFSRcolor4[476]&LFSRcolor4[660]&LFSRcolor4[264]);
    BiasedRNG[1057] = (LFSRcolor4[530]&LFSRcolor4[549]&LFSRcolor4[480]&LFSRcolor4[86]);
    BiasedRNG[1058] = (LFSRcolor4[133]&LFSRcolor4[959]&LFSRcolor4[61]&LFSRcolor4[52]);
    BiasedRNG[1059] = (LFSRcolor4[854]&LFSRcolor4[290]&LFSRcolor4[628]&LFSRcolor4[543]);
    BiasedRNG[1060] = (LFSRcolor4[623]&LFSRcolor4[885]&LFSRcolor4[385]&LFSRcolor4[471]);
    BiasedRNG[1061] = (LFSRcolor4[770]&LFSRcolor4[633]&LFSRcolor4[435]&LFSRcolor4[239]);
    BiasedRNG[1062] = (LFSRcolor4[493]&LFSRcolor4[842]&LFSRcolor4[428]&LFSRcolor4[783]);
    BiasedRNG[1063] = (LFSRcolor4[39]&LFSRcolor4[371]&LFSRcolor4[564]&LFSRcolor4[50]);
    BiasedRNG[1064] = (LFSRcolor4[686]&LFSRcolor4[25]&LFSRcolor4[524]&LFSRcolor4[131]);
    BiasedRNG[1065] = (LFSRcolor4[898]&LFSRcolor4[429]&LFSRcolor4[267]&LFSRcolor4[113]);
    BiasedRNG[1066] = (LFSRcolor4[566]&LFSRcolor4[281]&LFSRcolor4[91]&LFSRcolor4[630]);
    BiasedRNG[1067] = (LFSRcolor4[237]&LFSRcolor4[738]&LFSRcolor4[576]&LFSRcolor4[571]);
    BiasedRNG[1068] = (LFSRcolor4[923]&LFSRcolor4[763]&LFSRcolor4[689]&LFSRcolor4[359]);
    BiasedRNG[1069] = (LFSRcolor4[402]&LFSRcolor4[425]&LFSRcolor4[107]&LFSRcolor4[820]);
    BiasedRNG[1070] = (LFSRcolor4[596]&LFSRcolor4[82]&LFSRcolor4[863]&LFSRcolor4[153]);
    BiasedRNG[1071] = (LFSRcolor4[715]&LFSRcolor4[722]&LFSRcolor4[616]&LFSRcolor4[151]);
    BiasedRNG[1072] = (LFSRcolor4[876]&LFSRcolor4[809]&LFSRcolor4[80]&LFSRcolor4[644]);
    BiasedRNG[1073] = (LFSRcolor4[769]&LFSRcolor4[748]&LFSRcolor4[709]&LFSRcolor4[655]);
    BiasedRNG[1074] = (LFSRcolor4[516]&LFSRcolor4[311]&LFSRcolor4[265]&LFSRcolor4[284]);
    BiasedRNG[1075] = (LFSRcolor4[422]&LFSRcolor4[613]&LFSRcolor4[301]&LFSRcolor4[791]);
    BiasedRNG[1076] = (LFSRcolor4[683]&LFSRcolor4[150]&LFSRcolor4[364]&LFSRcolor4[852]);
    BiasedRNG[1077] = (LFSRcolor4[879]&LFSRcolor4[880]&LFSRcolor4[812]&LFSRcolor4[464]);
    BiasedRNG[1078] = (LFSRcolor4[104]&LFSRcolor4[559]&LFSRcolor4[434]&LFSRcolor4[733]);
    BiasedRNG[1079] = (LFSRcolor4[775]&LFSRcolor4[562]&LFSRcolor4[331]&LFSRcolor4[195]);
    BiasedRNG[1080] = (LFSRcolor4[805]&LFSRcolor4[889]&LFSRcolor4[609]&LFSRcolor4[48]);
    BiasedRNG[1081] = (LFSRcolor4[785]&LFSRcolor4[856]&LFSRcolor4[545]&LFSRcolor4[946]);
    BiasedRNG[1082] = (LFSRcolor4[826]&LFSRcolor4[950]&LFSRcolor4[65]&LFSRcolor4[462]);
    BiasedRNG[1083] = (LFSRcolor4[475]&LFSRcolor4[326]&LFSRcolor4[392]&LFSRcolor4[28]);
    BiasedRNG[1084] = (LFSRcolor4[911]&LFSRcolor4[139]&LFSRcolor4[106]&LFSRcolor4[205]);
    BiasedRNG[1085] = (LFSRcolor4[166]&LFSRcolor4[751]&LFSRcolor4[44]&LFSRcolor4[1]);
    BiasedRNG[1086] = (LFSRcolor4[515]&LFSRcolor4[668]&LFSRcolor4[302]&LFSRcolor4[847]);
    BiasedRNG[1087] = (LFSRcolor4[45]&LFSRcolor4[226]&LFSRcolor4[11]&LFSRcolor4[183]);
    BiasedRNG[1088] = (LFSRcolor4[201]&LFSRcolor4[750]&LFSRcolor4[501]&LFSRcolor4[416]);
    BiasedRNG[1089] = (LFSRcolor4[555]&LFSRcolor4[792]&LFSRcolor4[227]&LFSRcolor4[539]);
    BiasedRNG[1090] = (LFSRcolor4[705]&LFSRcolor4[136]&LFSRcolor4[232]&LFSRcolor4[625]);
    BiasedRNG[1091] = (LFSRcolor4[363]&LFSRcolor4[457]&LFSRcolor4[24]&LFSRcolor4[627]);
    BiasedRNG[1092] = (LFSRcolor4[79]&LFSRcolor4[815]&LFSRcolor4[580]&LFSRcolor4[573]);
    BiasedRNG[1093] = (LFSRcolor4[93]&LFSRcolor4[621]&LFSRcolor4[569]&LFSRcolor4[121]);
    BiasedRNG[1094] = (LFSRcolor4[266]&LFSRcolor4[720]&LFSRcolor4[788]&LFSRcolor4[500]);
    BiasedRNG[1095] = (LFSRcolor4[308]&LFSRcolor4[676]&LFSRcolor4[645]&LFSRcolor4[864]);
    BiasedRNG[1096] = (LFSRcolor4[725]&LFSRcolor4[542]&LFSRcolor4[887]&LFSRcolor4[152]);
    BiasedRNG[1097] = (LFSRcolor4[759]&LFSRcolor4[900]&LFSRcolor4[575]&LFSRcolor4[665]);
    BiasedRNG[1098] = (LFSRcolor4[96]&LFSRcolor4[59]&LFSRcolor4[661]&LFSRcolor4[347]);
    BiasedRNG[1099] = (LFSRcolor4[386]&LFSRcolor4[874]&LFSRcolor4[278]&LFSRcolor4[362]);
    BiasedRNG[1100] = (LFSRcolor4[654]&LFSRcolor4[394]&LFSRcolor4[272]&LFSRcolor4[64]);
    BiasedRNG[1101] = (LFSRcolor4[431]&LFSRcolor4[380]&LFSRcolor4[137]&LFSRcolor4[438]);
    BiasedRNG[1102] = (LFSRcolor4[361]&LFSRcolor4[953]&LFSRcolor4[925]&LFSRcolor4[760]);
    BiasedRNG[1103] = (LFSRcolor4[458]&LFSRcolor4[563]&LFSRcolor4[384]&LFSRcolor4[376]);
    BiasedRNG[1104] = (LFSRcolor4[903]&LFSRcolor4[164]&LFSRcolor4[346]&LFSRcolor4[702]);
    BiasedRNG[1105] = (LFSRcolor4[541]&LFSRcolor4[917]&LFSRcolor4[42]&LFSRcolor4[234]);
    BiasedRNG[1106] = (LFSRcolor4[632]&LFSRcolor4[367]&LFSRcolor4[220]&LFSRcolor4[587]);
    BiasedRNG[1107] = (LFSRcolor4[217]&LFSRcolor4[354]&LFSRcolor4[35]&LFSRcolor4[662]);
    BiasedRNG[1108] = (LFSRcolor4[468]&LFSRcolor4[181]&LFSRcolor4[821]&LFSRcolor4[943]);
    BiasedRNG[1109] = (LFSRcolor4[631]&LFSRcolor4[728]&LFSRcolor4[552]&LFSRcolor4[897]);
    BiasedRNG[1110] = (LFSRcolor4[206]&LFSRcolor4[653]&LFSRcolor4[473]&LFSRcolor4[913]);
    BiasedRNG[1111] = (LFSRcolor4[77]&LFSRcolor4[483]&LFSRcolor4[797]&LFSRcolor4[790]);
    BiasedRNG[1112] = (LFSRcolor4[657]&LFSRcolor4[553]&LFSRcolor4[469]&LFSRcolor4[203]);
    BiasedRNG[1113] = (LFSRcolor4[651]&LFSRcolor4[446]&LFSRcolor4[579]&LFSRcolor4[739]);
    BiasedRNG[1114] = (LFSRcolor4[731]&LFSRcolor4[626]&LFSRcolor4[942]&LFSRcolor4[333]);
    BiasedRNG[1115] = (LFSRcolor4[487]&LFSRcolor4[664]&LFSRcolor4[764]&LFSRcolor4[189]);
    BiasedRNG[1116] = (LFSRcolor4[456]&LFSRcolor4[803]&LFSRcolor4[612]&LFSRcolor4[742]);
    BiasedRNG[1117] = (LFSRcolor4[188]&LFSRcolor4[861]&LFSRcolor4[54]&LFSRcolor4[839]);
    BiasedRNG[1118] = (LFSRcolor4[617]&LFSRcolor4[536]&LFSRcolor4[40]&LFSRcolor4[682]);
    BiasedRNG[1119] = (LFSRcolor4[193]&LFSRcolor4[605]&LFSRcolor4[781]&LFSRcolor4[698]);
    BiasedRNG[1120] = (LFSRcolor4[735]&LFSRcolor4[440]&LFSRcolor4[103]&LFSRcolor4[825]);
    BiasedRNG[1121] = (LFSRcolor4[814]&LFSRcolor4[88]&LFSRcolor4[238]&LFSRcolor4[271]);
    BiasedRNG[1122] = (LFSRcolor4[780]&LFSRcolor4[714]&LFSRcolor4[851]&LFSRcolor4[397]);
    BiasedRNG[1123] = (LFSRcolor4[231]&LFSRcolor4[73]&LFSRcolor4[878]&LFSRcolor4[918]);
    BiasedRNG[1124] = (LFSRcolor4[388]&LFSRcolor4[908]&LFSRcolor4[510]&LFSRcolor4[27]);
    BiasedRNG[1125] = (LFSRcolor4[412]&LFSRcolor4[357]&LFSRcolor4[145]&LFSRcolor4[904]);
    BiasedRNG[1126] = (LFSRcolor4[699]&LFSRcolor4[584]&LFSRcolor4[834]&LFSRcolor4[18]);
    BiasedRNG[1127] = (LFSRcolor4[757]&LFSRcolor4[250]&LFSRcolor4[920]&LFSRcolor4[196]);
    BiasedRNG[1128] = (LFSRcolor4[881]&LFSRcolor4[528]&LFSRcolor4[160]&LFSRcolor4[320]);
    BiasedRNG[1129] = (LFSRcolor4[49]&LFSRcolor4[83]&LFSRcolor4[849]&LFSRcolor4[159]);
    BiasedRNG[1130] = (LFSRcolor4[353]&LFSRcolor4[60]&LFSRcolor4[776]&LFSRcolor4[659]);
    BiasedRNG[1131] = (LFSRcolor4[147]&LFSRcolor4[961]&LFSRcolor4[802]&LFSRcolor4[574]);
    BiasedRNG[1132] = (LFSRcolor4[253]&LFSRcolor4[811]&LFSRcolor4[935]&LFSRcolor4[557]);
    BiasedRNG[1133] = (LFSRcolor4[403]&LFSRcolor4[94]&LFSRcolor4[287]&LFSRcolor4[309]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule