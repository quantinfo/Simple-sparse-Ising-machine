//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [37:0] counter;
initial counter = 38'b0;
reg [23:0] solution;
reg [23:0] solution_check;
wire [23:0] solution_set;
initial solution_check = 24'b111111000010001011111101;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
reg [0:1151] InitCond;
reg run;
wire [643:0] LFSRcolor0;
wire [781:0] LFSRcolor1;
wire [597:0] LFSRcolor2;
wire [137:0] LFSRcolor3;
wire [413:0] LFSRcolor4;
reg [657:0] BiasedRNG;       //For I=+/-1 cases
reg [493:0] UnbiasedRNG;   //For I=0 cases
reg [0:1187] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[384] = 1'b1;
initial m[531] = 1'b0;
initial m[541] = 1'b1;
initial m[556] = 1'b1;
initial m[576] = 1'b1;
initial m[601] = 1'b1;
initial m[631] = 1'b1;
initial m[666] = 1'b1;
initial m[706] = 1'b0;
initial m[751] = 1'b1;
initial m[801] = 1'b0;
initial m[856] = 1'b0;
initial m[911] = 1'b0;
initial m[961] = 1'b1;
initial m[1006] = 1'b0;
initial m[1046] = 1'b0;
initial m[1081] = 1'b0;
initial m[1111] = 1'b0;
initial m[1136] = 1'b1;
initial m[1156] = 1'b1;
initial m[1171] = 1'b1;
initial m[1181] = 1'b1;
initial m[1186] = 1'b1;
initial m[1187] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[530] = 1'b0;
initial m[540] = 1'b0;
initial m[555] = 1'b0;
initial m[575] = 1'b0;
initial m[600] = 1'b0;
initial m[630] = 1'b0;
initial m[665] = 1'b0;
initial m[705] = 1'b0;
initial m[750] = 1'b0;
initial m[800] = 1'b0;
initial m[855] = 1'b0;
initial m[858] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR0_11(.LFSRregister(LFSRcolor0[551:506]),.clk(sample_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR0_12(.LFSRregister(LFSRcolor0[597:552]),.clk(sample_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR0_13(.LFSRregister(LFSRcolor0[643:598]),.clk(sample_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR1_15(.LFSRregister(LFSRcolor1[735:690]),.clk(color0_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR1_16(.LFSRregister(LFSRcolor1[781:736]),.clk(color0_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR2_11(.LFSRregister(LFSRcolor2[551:506]),.clk(color1_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR2_12(.LFSRregister(LFSRcolor2[597:552]),.clk(color1_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR3_2(.LFSRregister(LFSRcolor3[137:92]),.clk(color2_clk));
lfsr #(.seed(46'b0011001000010001001111001110101111011111000110)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b0101000110100000010101001000010000101101100110)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1110011010010011001010111010100101111111100000)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b1001111000010100100001100010110000001111101011)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b0011101001111100110111000000010000101100111110)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b1010111010001100001100010110010011100100101100)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b1101010000110001000001011010110100010000110101)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b0111111000001001010001100011001110110101101001)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));
lfsr #(.seed(46'b0111011110101100100001111000001001111001010010)) LFSR4_8(.LFSRregister(LFSRcolor4[413:368]),.clk(color3_clk));
//To control whether the system runs or resets using VIO and counter:
always @(posedge sample_clk) begin
    if (reset) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 24'b0;
        failure = 1'b0;
        solution_check = solution_set;
        m[384] = solution_set[0];
        m[531] = solution_set[1];
        m[541] = solution_set[2];
        m[556] = solution_set[3];
        m[576] = solution_set[4];
        m[601] = solution_set[5];
        m[631] = solution_set[6];
        m[666] = solution_set[7];
        m[706] = solution_set[8];
        m[751] = solution_set[9];
        m[801] = solution_set[10];
        m[856] = solution_set[11];
        m[911] = solution_set[12];
        m[961] = solution_set[13];
        m[1006] = solution_set[14];
        m[1046] = solution_set[15];
        m[1081] = solution_set[16];
        m[1111] = solution_set[17];
        m[1136] = solution_set[18];
        m[1156] = solution_set[19];
        m[1171] = solution_set[20];
        m[1181] = solution_set[21];
        m[1186] = solution_set[22];
        m[1187] = solution_set[23];
    end else if (solution_flag) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 24'b0;
        failure = 1'b0;
    end else if (counter < 38'b11111111111111111111111111111111111111) begin
        if (counter == 1) begin
            InitCond[0] = UnbiasedRNG[0];
            InitCond[1] = UnbiasedRNG[1];
            InitCond[2] = UnbiasedRNG[2];
            InitCond[3] = UnbiasedRNG[3];
            InitCond[4] = UnbiasedRNG[4];
            InitCond[5] = UnbiasedRNG[5];
            InitCond[6] = UnbiasedRNG[6];
            InitCond[7] = UnbiasedRNG[7];
            InitCond[8] = UnbiasedRNG[8];
            InitCond[9] = UnbiasedRNG[9];
            InitCond[10] = UnbiasedRNG[10];
            InitCond[11] = UnbiasedRNG[11];
            InitCond[12] = UnbiasedRNG[12];
            InitCond[13] = UnbiasedRNG[13];
            InitCond[14] = UnbiasedRNG[14];
            InitCond[15] = UnbiasedRNG[15];
            InitCond[16] = UnbiasedRNG[16];
            InitCond[17] = UnbiasedRNG[17];
            InitCond[18] = UnbiasedRNG[18];
            InitCond[19] = UnbiasedRNG[19];
            InitCond[20] = UnbiasedRNG[20];
            InitCond[21] = UnbiasedRNG[21];
            InitCond[22] = UnbiasedRNG[22];
            InitCond[23] = UnbiasedRNG[23];
            InitCond[24] = UnbiasedRNG[24];
            InitCond[25] = UnbiasedRNG[25];
            InitCond[26] = UnbiasedRNG[26];
            InitCond[27] = UnbiasedRNG[27];
            InitCond[28] = UnbiasedRNG[28];
            InitCond[29] = UnbiasedRNG[29];
            InitCond[30] = UnbiasedRNG[30];
            InitCond[31] = UnbiasedRNG[31];
            InitCond[32] = UnbiasedRNG[32];
            InitCond[33] = UnbiasedRNG[33];
            InitCond[34] = UnbiasedRNG[34];
            InitCond[35] = UnbiasedRNG[35];
            InitCond[36] = UnbiasedRNG[36];
            InitCond[37] = UnbiasedRNG[37];
            InitCond[38] = UnbiasedRNG[38];
            InitCond[39] = UnbiasedRNG[39];
            InitCond[40] = UnbiasedRNG[40];
            InitCond[41] = UnbiasedRNG[41];
            InitCond[42] = UnbiasedRNG[42];
            InitCond[43] = UnbiasedRNG[43];
            InitCond[44] = UnbiasedRNG[44];
            InitCond[45] = UnbiasedRNG[45];
            InitCond[46] = UnbiasedRNG[46];
            InitCond[47] = UnbiasedRNG[47];
            InitCond[48] = UnbiasedRNG[48];
            InitCond[49] = UnbiasedRNG[49];
            InitCond[50] = UnbiasedRNG[50];
            InitCond[51] = UnbiasedRNG[51];
            InitCond[52] = UnbiasedRNG[52];
            InitCond[53] = UnbiasedRNG[53];
            InitCond[54] = UnbiasedRNG[54];
            InitCond[55] = UnbiasedRNG[55];
            InitCond[56] = UnbiasedRNG[56];
            InitCond[57] = UnbiasedRNG[57];
            InitCond[58] = UnbiasedRNG[58];
            InitCond[59] = UnbiasedRNG[59];
            InitCond[60] = UnbiasedRNG[60];
            InitCond[61] = UnbiasedRNG[61];
            InitCond[62] = UnbiasedRNG[62];
            InitCond[63] = UnbiasedRNG[63];
            InitCond[64] = UnbiasedRNG[64];
            InitCond[65] = UnbiasedRNG[65];
            InitCond[66] = UnbiasedRNG[66];
            InitCond[67] = UnbiasedRNG[67];
            InitCond[68] = UnbiasedRNG[68];
            InitCond[69] = UnbiasedRNG[69];
            InitCond[70] = UnbiasedRNG[70];
            InitCond[71] = UnbiasedRNG[71];
            InitCond[72] = UnbiasedRNG[72];
            InitCond[73] = UnbiasedRNG[73];
            InitCond[74] = UnbiasedRNG[74];
            InitCond[75] = UnbiasedRNG[75];
            InitCond[76] = UnbiasedRNG[76];
            InitCond[77] = UnbiasedRNG[77];
            InitCond[78] = UnbiasedRNG[78];
            InitCond[79] = UnbiasedRNG[79];
            InitCond[80] = UnbiasedRNG[80];
            InitCond[81] = UnbiasedRNG[81];
            InitCond[82] = UnbiasedRNG[82];
            InitCond[83] = UnbiasedRNG[83];
            InitCond[84] = UnbiasedRNG[84];
            InitCond[85] = UnbiasedRNG[85];
            InitCond[86] = UnbiasedRNG[86];
            InitCond[87] = UnbiasedRNG[87];
            InitCond[88] = UnbiasedRNG[88];
            InitCond[89] = UnbiasedRNG[89];
            InitCond[90] = UnbiasedRNG[90];
            InitCond[91] = UnbiasedRNG[91];
            InitCond[92] = UnbiasedRNG[92];
            InitCond[93] = UnbiasedRNG[93];
            InitCond[94] = UnbiasedRNG[94];
            InitCond[95] = UnbiasedRNG[95];
            InitCond[96] = UnbiasedRNG[96];
            InitCond[97] = UnbiasedRNG[97];
            InitCond[98] = UnbiasedRNG[98];
            InitCond[99] = UnbiasedRNG[99];
            InitCond[100] = UnbiasedRNG[100];
            InitCond[101] = UnbiasedRNG[101];
            InitCond[102] = UnbiasedRNG[102];
            InitCond[103] = UnbiasedRNG[103];
            InitCond[104] = UnbiasedRNG[104];
            InitCond[105] = UnbiasedRNG[105];
            InitCond[106] = UnbiasedRNG[106];
            InitCond[107] = UnbiasedRNG[107];
            InitCond[108] = UnbiasedRNG[108];
            InitCond[109] = UnbiasedRNG[109];
            InitCond[110] = UnbiasedRNG[110];
            InitCond[111] = UnbiasedRNG[111];
            InitCond[112] = UnbiasedRNG[112];
            InitCond[113] = UnbiasedRNG[113];
            InitCond[114] = UnbiasedRNG[114];
            InitCond[115] = UnbiasedRNG[115];
            InitCond[116] = UnbiasedRNG[116];
            InitCond[117] = UnbiasedRNG[117];
            InitCond[118] = UnbiasedRNG[118];
            InitCond[119] = UnbiasedRNG[119];
            InitCond[120] = UnbiasedRNG[120];
            InitCond[121] = UnbiasedRNG[121];
            InitCond[122] = UnbiasedRNG[122];
            InitCond[123] = UnbiasedRNG[123];
            InitCond[124] = UnbiasedRNG[124];
            InitCond[125] = UnbiasedRNG[125];
            InitCond[126] = UnbiasedRNG[126];
            InitCond[127] = UnbiasedRNG[127];
            InitCond[128] = UnbiasedRNG[128];
            InitCond[129] = UnbiasedRNG[129];
            InitCond[130] = UnbiasedRNG[130];
            InitCond[131] = UnbiasedRNG[131];
            InitCond[132] = UnbiasedRNG[132];
            InitCond[133] = UnbiasedRNG[133];
            InitCond[134] = UnbiasedRNG[134];
            InitCond[135] = UnbiasedRNG[135];
            InitCond[136] = UnbiasedRNG[136];
            InitCond[137] = UnbiasedRNG[137];
            InitCond[138] = UnbiasedRNG[138];
            InitCond[139] = UnbiasedRNG[139];
            InitCond[140] = UnbiasedRNG[140];
            InitCond[141] = UnbiasedRNG[141];
            InitCond[142] = UnbiasedRNG[142];
            InitCond[143] = UnbiasedRNG[143];
            InitCond[144] = UnbiasedRNG[144];
            InitCond[145] = UnbiasedRNG[145];
            InitCond[146] = UnbiasedRNG[146];
            InitCond[147] = UnbiasedRNG[147];
            InitCond[148] = UnbiasedRNG[148];
            InitCond[149] = UnbiasedRNG[149];
            InitCond[150] = UnbiasedRNG[150];
            InitCond[151] = UnbiasedRNG[151];
            InitCond[152] = UnbiasedRNG[152];
            InitCond[153] = UnbiasedRNG[153];
            InitCond[154] = UnbiasedRNG[154];
            InitCond[155] = UnbiasedRNG[155];
            InitCond[156] = UnbiasedRNG[156];
            InitCond[157] = UnbiasedRNG[157];
            InitCond[158] = UnbiasedRNG[158];
            InitCond[159] = UnbiasedRNG[159];
            InitCond[160] = UnbiasedRNG[160];
            InitCond[161] = UnbiasedRNG[161];
            InitCond[162] = UnbiasedRNG[162];
            InitCond[163] = UnbiasedRNG[163];
            InitCond[164] = UnbiasedRNG[164];
            InitCond[165] = UnbiasedRNG[165];
            InitCond[166] = UnbiasedRNG[166];
            InitCond[167] = UnbiasedRNG[167];
            InitCond[168] = UnbiasedRNG[168];
            InitCond[169] = UnbiasedRNG[169];
            InitCond[170] = UnbiasedRNG[170];
            InitCond[171] = UnbiasedRNG[171];
            InitCond[172] = UnbiasedRNG[172];
            InitCond[173] = UnbiasedRNG[173];
            InitCond[174] = UnbiasedRNG[174];
            InitCond[175] = UnbiasedRNG[175];
            InitCond[176] = UnbiasedRNG[176];
            InitCond[177] = UnbiasedRNG[177];
            InitCond[178] = UnbiasedRNG[178];
            InitCond[179] = UnbiasedRNG[179];
            InitCond[180] = UnbiasedRNG[180];
            InitCond[181] = UnbiasedRNG[181];
            InitCond[182] = UnbiasedRNG[182];
            InitCond[183] = UnbiasedRNG[183];
            InitCond[184] = UnbiasedRNG[184];
            InitCond[185] = UnbiasedRNG[185];
            InitCond[186] = UnbiasedRNG[186];
            InitCond[187] = UnbiasedRNG[187];
            InitCond[188] = UnbiasedRNG[188];
            InitCond[189] = UnbiasedRNG[189];
            InitCond[190] = UnbiasedRNG[190];
            InitCond[191] = UnbiasedRNG[191];
            InitCond[192] = UnbiasedRNG[192];
            InitCond[193] = UnbiasedRNG[193];
            InitCond[194] = UnbiasedRNG[194];
            InitCond[195] = UnbiasedRNG[195];
            InitCond[196] = UnbiasedRNG[196];
            InitCond[197] = UnbiasedRNG[197];
            InitCond[198] = UnbiasedRNG[198];
            InitCond[199] = UnbiasedRNG[199];
            InitCond[200] = UnbiasedRNG[200];
            InitCond[201] = UnbiasedRNG[201];
            InitCond[202] = UnbiasedRNG[202];
            InitCond[203] = UnbiasedRNG[203];
            InitCond[204] = UnbiasedRNG[204];
            InitCond[205] = UnbiasedRNG[205];
            InitCond[206] = UnbiasedRNG[206];
            InitCond[207] = UnbiasedRNG[207];
            InitCond[208] = UnbiasedRNG[208];
            InitCond[209] = UnbiasedRNG[209];
            InitCond[210] = UnbiasedRNG[210];
            InitCond[211] = UnbiasedRNG[211];
            InitCond[212] = UnbiasedRNG[212];
            InitCond[213] = UnbiasedRNG[213];
            InitCond[214] = UnbiasedRNG[214];
            InitCond[215] = UnbiasedRNG[215];
            InitCond[216] = UnbiasedRNG[216];
            InitCond[217] = UnbiasedRNG[217];
            InitCond[218] = UnbiasedRNG[218];
            InitCond[219] = UnbiasedRNG[219];
            InitCond[220] = UnbiasedRNG[220];
            InitCond[221] = UnbiasedRNG[221];
            InitCond[222] = UnbiasedRNG[222];
            InitCond[223] = UnbiasedRNG[223];
            InitCond[224] = UnbiasedRNG[224];
            InitCond[225] = UnbiasedRNG[225];
            InitCond[226] = UnbiasedRNG[226];
            InitCond[227] = UnbiasedRNG[227];
            InitCond[228] = UnbiasedRNG[228];
            InitCond[229] = UnbiasedRNG[229];
            InitCond[230] = UnbiasedRNG[230];
            InitCond[231] = UnbiasedRNG[231];
            InitCond[232] = UnbiasedRNG[232];
            InitCond[233] = UnbiasedRNG[233];
            InitCond[234] = UnbiasedRNG[234];
            InitCond[235] = UnbiasedRNG[235];
            InitCond[236] = UnbiasedRNG[236];
            InitCond[237] = UnbiasedRNG[237];
            InitCond[238] = UnbiasedRNG[238];
            InitCond[239] = UnbiasedRNG[239];
            InitCond[240] = UnbiasedRNG[240];
            InitCond[241] = UnbiasedRNG[241];
            InitCond[242] = UnbiasedRNG[242];
            InitCond[243] = UnbiasedRNG[243];
            InitCond[244] = UnbiasedRNG[244];
            InitCond[245] = UnbiasedRNG[245];
            InitCond[246] = UnbiasedRNG[246];
            InitCond[247] = UnbiasedRNG[247];
            InitCond[248] = UnbiasedRNG[248];
            InitCond[249] = UnbiasedRNG[249];
            InitCond[250] = UnbiasedRNG[250];
            InitCond[251] = UnbiasedRNG[251];
            InitCond[252] = UnbiasedRNG[252];
            InitCond[253] = UnbiasedRNG[253];
            InitCond[254] = UnbiasedRNG[254];
            InitCond[255] = UnbiasedRNG[255];
            InitCond[256] = UnbiasedRNG[256];
            InitCond[257] = UnbiasedRNG[257];
            InitCond[258] = UnbiasedRNG[258];
            InitCond[259] = UnbiasedRNG[259];
            InitCond[260] = UnbiasedRNG[260];
            InitCond[261] = UnbiasedRNG[261];
            InitCond[262] = UnbiasedRNG[262];
            InitCond[263] = UnbiasedRNG[263];
            InitCond[264] = UnbiasedRNG[264];
            InitCond[265] = UnbiasedRNG[265];
            InitCond[266] = UnbiasedRNG[266];
            InitCond[267] = UnbiasedRNG[267];
            InitCond[268] = UnbiasedRNG[268];
            InitCond[269] = UnbiasedRNG[269];
            InitCond[270] = UnbiasedRNG[270];
            InitCond[271] = UnbiasedRNG[271];
            InitCond[272] = UnbiasedRNG[272];
            InitCond[273] = UnbiasedRNG[273];
            InitCond[274] = UnbiasedRNG[274];
            InitCond[275] = UnbiasedRNG[275];
            InitCond[276] = UnbiasedRNG[276];
            InitCond[277] = UnbiasedRNG[277];
            InitCond[278] = UnbiasedRNG[278];
            InitCond[279] = UnbiasedRNG[279];
            InitCond[280] = UnbiasedRNG[280];
            InitCond[281] = UnbiasedRNG[281];
            InitCond[282] = UnbiasedRNG[282];
            InitCond[283] = UnbiasedRNG[283];
            InitCond[284] = UnbiasedRNG[284];
            InitCond[285] = UnbiasedRNG[285];
            InitCond[286] = UnbiasedRNG[286];
            InitCond[287] = UnbiasedRNG[287];
            InitCond[288] = UnbiasedRNG[288];
            InitCond[289] = UnbiasedRNG[289];
            InitCond[290] = UnbiasedRNG[290];
            InitCond[291] = UnbiasedRNG[291];
            InitCond[292] = UnbiasedRNG[292];
            InitCond[293] = UnbiasedRNG[293];
            InitCond[294] = UnbiasedRNG[294];
            InitCond[295] = UnbiasedRNG[295];
            InitCond[296] = UnbiasedRNG[296];
            InitCond[297] = UnbiasedRNG[297];
            InitCond[298] = UnbiasedRNG[298];
            InitCond[299] = UnbiasedRNG[299];
            InitCond[300] = UnbiasedRNG[300];
            InitCond[301] = UnbiasedRNG[301];
            InitCond[302] = UnbiasedRNG[302];
            InitCond[303] = UnbiasedRNG[303];
            InitCond[304] = UnbiasedRNG[304];
            InitCond[305] = UnbiasedRNG[305];
            InitCond[306] = UnbiasedRNG[306];
            InitCond[307] = UnbiasedRNG[307];
            InitCond[308] = UnbiasedRNG[308];
            InitCond[309] = UnbiasedRNG[309];
            InitCond[310] = UnbiasedRNG[310];
            InitCond[311] = UnbiasedRNG[311];
            InitCond[312] = UnbiasedRNG[312];
            InitCond[313] = UnbiasedRNG[313];
            InitCond[314] = UnbiasedRNG[314];
            InitCond[315] = UnbiasedRNG[315];
            InitCond[316] = UnbiasedRNG[316];
            InitCond[317] = UnbiasedRNG[317];
            InitCond[318] = UnbiasedRNG[318];
            InitCond[319] = UnbiasedRNG[319];
            InitCond[320] = UnbiasedRNG[320];
            InitCond[321] = UnbiasedRNG[321];
            InitCond[322] = UnbiasedRNG[322];
            InitCond[323] = UnbiasedRNG[323];
            InitCond[324] = UnbiasedRNG[324];
            InitCond[325] = UnbiasedRNG[325];
            InitCond[326] = UnbiasedRNG[326];
            InitCond[327] = UnbiasedRNG[327];
            InitCond[328] = UnbiasedRNG[328];
            InitCond[329] = UnbiasedRNG[329];
            InitCond[330] = UnbiasedRNG[330];
            InitCond[331] = UnbiasedRNG[331];
            InitCond[332] = UnbiasedRNG[332];
            InitCond[333] = UnbiasedRNG[333];
            InitCond[334] = UnbiasedRNG[334];
            InitCond[335] = UnbiasedRNG[335];
            InitCond[336] = UnbiasedRNG[336];
            InitCond[337] = UnbiasedRNG[337];
            InitCond[338] = UnbiasedRNG[338];
            InitCond[339] = UnbiasedRNG[339];
            InitCond[340] = UnbiasedRNG[340];
            InitCond[341] = UnbiasedRNG[341];
            InitCond[342] = UnbiasedRNG[342];
            InitCond[343] = UnbiasedRNG[343];
            InitCond[344] = UnbiasedRNG[344];
            InitCond[345] = UnbiasedRNG[345];
            InitCond[346] = UnbiasedRNG[346];
            InitCond[347] = UnbiasedRNG[347];
            InitCond[348] = UnbiasedRNG[348];
            InitCond[349] = UnbiasedRNG[349];
            InitCond[350] = UnbiasedRNG[350];
            InitCond[351] = UnbiasedRNG[351];
            InitCond[352] = UnbiasedRNG[352];
            InitCond[353] = UnbiasedRNG[353];
            InitCond[354] = UnbiasedRNG[354];
            InitCond[355] = UnbiasedRNG[355];
            InitCond[356] = UnbiasedRNG[356];
            InitCond[357] = UnbiasedRNG[357];
            InitCond[358] = UnbiasedRNG[358];
            InitCond[359] = UnbiasedRNG[359];
            InitCond[360] = UnbiasedRNG[360];
            InitCond[361] = UnbiasedRNG[361];
            InitCond[362] = UnbiasedRNG[362];
            InitCond[363] = UnbiasedRNG[363];
            InitCond[364] = UnbiasedRNG[364];
            InitCond[365] = UnbiasedRNG[365];
            InitCond[366] = UnbiasedRNG[366];
            InitCond[367] = UnbiasedRNG[367];
            InitCond[368] = UnbiasedRNG[368];
            InitCond[369] = UnbiasedRNG[369];
            InitCond[370] = UnbiasedRNG[370];
            InitCond[371] = UnbiasedRNG[371];
            InitCond[372] = UnbiasedRNG[372];
            InitCond[373] = UnbiasedRNG[373];
            InitCond[374] = UnbiasedRNG[374];
            InitCond[375] = UnbiasedRNG[375];
            InitCond[376] = UnbiasedRNG[376];
            InitCond[377] = UnbiasedRNG[377];
            InitCond[378] = UnbiasedRNG[378];
            InitCond[379] = UnbiasedRNG[379];
            InitCond[380] = UnbiasedRNG[380];
            InitCond[381] = UnbiasedRNG[381];
            InitCond[382] = UnbiasedRNG[382];
            InitCond[383] = UnbiasedRNG[383];
            InitCond[384] = UnbiasedRNG[384];
            InitCond[385] = UnbiasedRNG[385];
            InitCond[386] = UnbiasedRNG[386];
            InitCond[387] = UnbiasedRNG[387];
            InitCond[388] = UnbiasedRNG[388];
            InitCond[389] = UnbiasedRNG[389];
            InitCond[390] = UnbiasedRNG[390];
            InitCond[391] = UnbiasedRNG[391];
            InitCond[392] = UnbiasedRNG[392];
            InitCond[393] = UnbiasedRNG[393];
            InitCond[394] = UnbiasedRNG[394];
            InitCond[395] = UnbiasedRNG[395];
            InitCond[396] = UnbiasedRNG[396];
            InitCond[397] = UnbiasedRNG[397];
            InitCond[398] = UnbiasedRNG[398];
            InitCond[399] = UnbiasedRNG[399];
            InitCond[400] = UnbiasedRNG[400];
            InitCond[401] = UnbiasedRNG[401];
            InitCond[402] = UnbiasedRNG[402];
            InitCond[403] = UnbiasedRNG[403];
            InitCond[404] = UnbiasedRNG[404];
            InitCond[405] = UnbiasedRNG[405];
            InitCond[406] = UnbiasedRNG[406];
            InitCond[407] = UnbiasedRNG[407];
            InitCond[408] = UnbiasedRNG[408];
            InitCond[409] = UnbiasedRNG[409];
            InitCond[410] = UnbiasedRNG[410];
            InitCond[411] = UnbiasedRNG[411];
            InitCond[412] = UnbiasedRNG[412];
            InitCond[413] = UnbiasedRNG[413];
            InitCond[414] = UnbiasedRNG[414];
            InitCond[415] = UnbiasedRNG[415];
            InitCond[416] = UnbiasedRNG[416];
            InitCond[417] = UnbiasedRNG[417];
            InitCond[418] = UnbiasedRNG[418];
            InitCond[419] = UnbiasedRNG[419];
            InitCond[420] = UnbiasedRNG[420];
            InitCond[421] = UnbiasedRNG[421];
            InitCond[422] = UnbiasedRNG[422];
            InitCond[423] = UnbiasedRNG[423];
            InitCond[424] = UnbiasedRNG[424];
            InitCond[425] = UnbiasedRNG[425];
            InitCond[426] = UnbiasedRNG[426];
            InitCond[427] = UnbiasedRNG[427];
            InitCond[428] = UnbiasedRNG[428];
            InitCond[429] = UnbiasedRNG[429];
            InitCond[430] = UnbiasedRNG[430];
            InitCond[431] = UnbiasedRNG[431];
            InitCond[432] = UnbiasedRNG[432];
            InitCond[433] = UnbiasedRNG[433];
            InitCond[434] = UnbiasedRNG[434];
            InitCond[435] = UnbiasedRNG[435];
            InitCond[436] = UnbiasedRNG[436];
            InitCond[437] = UnbiasedRNG[437];
            InitCond[438] = UnbiasedRNG[438];
            InitCond[439] = UnbiasedRNG[439];
            InitCond[440] = UnbiasedRNG[440];
            InitCond[441] = UnbiasedRNG[441];
            InitCond[442] = UnbiasedRNG[442];
            InitCond[443] = UnbiasedRNG[443];
            InitCond[444] = UnbiasedRNG[444];
            InitCond[445] = UnbiasedRNG[445];
            InitCond[446] = UnbiasedRNG[446];
            InitCond[447] = UnbiasedRNG[447];
            InitCond[448] = UnbiasedRNG[448];
            InitCond[449] = UnbiasedRNG[449];
            InitCond[450] = UnbiasedRNG[450];
            InitCond[451] = UnbiasedRNG[451];
            InitCond[452] = UnbiasedRNG[452];
            InitCond[453] = UnbiasedRNG[453];
            InitCond[454] = UnbiasedRNG[454];
            InitCond[455] = UnbiasedRNG[455];
            InitCond[456] = UnbiasedRNG[456];
            InitCond[457] = UnbiasedRNG[457];
            InitCond[458] = UnbiasedRNG[458];
            InitCond[459] = UnbiasedRNG[459];
            InitCond[460] = UnbiasedRNG[460];
            InitCond[461] = UnbiasedRNG[461];
            InitCond[462] = UnbiasedRNG[462];
            InitCond[463] = UnbiasedRNG[463];
            InitCond[464] = UnbiasedRNG[464];
            InitCond[465] = UnbiasedRNG[465];
            InitCond[466] = UnbiasedRNG[466];
            InitCond[467] = UnbiasedRNG[467];
            InitCond[468] = UnbiasedRNG[468];
            InitCond[469] = UnbiasedRNG[469];
            InitCond[470] = UnbiasedRNG[470];
            InitCond[471] = UnbiasedRNG[471];
            InitCond[472] = UnbiasedRNG[472];
            InitCond[473] = UnbiasedRNG[473];
            InitCond[474] = UnbiasedRNG[474];
            InitCond[475] = UnbiasedRNG[475];
            InitCond[476] = UnbiasedRNG[476];
            InitCond[477] = UnbiasedRNG[477];
            InitCond[478] = UnbiasedRNG[478];
            InitCond[479] = UnbiasedRNG[479];
            InitCond[480] = UnbiasedRNG[480];
            InitCond[481] = UnbiasedRNG[481];
            InitCond[482] = UnbiasedRNG[482];
            InitCond[483] = UnbiasedRNG[483];
            InitCond[484] = UnbiasedRNG[484];
            InitCond[485] = UnbiasedRNG[485];
            InitCond[486] = UnbiasedRNG[486];
            InitCond[487] = UnbiasedRNG[487];
            InitCond[488] = UnbiasedRNG[488];
            InitCond[489] = UnbiasedRNG[489];
            InitCond[490] = UnbiasedRNG[490];
            InitCond[491] = UnbiasedRNG[491];
            InitCond[492] = UnbiasedRNG[492];
            InitCond[493] = UnbiasedRNG[493];
        end
        else if (counter == 2) begin
            InitCond[494] = UnbiasedRNG[0];
            InitCond[495] = UnbiasedRNG[1];
            InitCond[496] = UnbiasedRNG[2];
            InitCond[497] = UnbiasedRNG[3];
            InitCond[498] = UnbiasedRNG[4];
            InitCond[499] = UnbiasedRNG[5];
            InitCond[500] = UnbiasedRNG[6];
            InitCond[501] = UnbiasedRNG[7];
            InitCond[502] = UnbiasedRNG[8];
            InitCond[503] = UnbiasedRNG[9];
            InitCond[504] = UnbiasedRNG[10];
            InitCond[505] = UnbiasedRNG[11];
            InitCond[506] = UnbiasedRNG[12];
            InitCond[507] = UnbiasedRNG[13];
            InitCond[508] = UnbiasedRNG[14];
            InitCond[509] = UnbiasedRNG[15];
            InitCond[510] = UnbiasedRNG[16];
            InitCond[511] = UnbiasedRNG[17];
            InitCond[512] = UnbiasedRNG[18];
            InitCond[513] = UnbiasedRNG[19];
            InitCond[514] = UnbiasedRNG[20];
            InitCond[515] = UnbiasedRNG[21];
            InitCond[516] = UnbiasedRNG[22];
            InitCond[517] = UnbiasedRNG[23];
            InitCond[518] = UnbiasedRNG[24];
            InitCond[519] = UnbiasedRNG[25];
            InitCond[520] = UnbiasedRNG[26];
            InitCond[521] = UnbiasedRNG[27];
            InitCond[522] = UnbiasedRNG[28];
            InitCond[523] = UnbiasedRNG[29];
            InitCond[524] = UnbiasedRNG[30];
            InitCond[525] = UnbiasedRNG[31];
            InitCond[526] = UnbiasedRNG[32];
            InitCond[527] = UnbiasedRNG[33];
            InitCond[528] = UnbiasedRNG[34];
            InitCond[529] = UnbiasedRNG[35];
            InitCond[530] = UnbiasedRNG[36];
            InitCond[531] = UnbiasedRNG[37];
            InitCond[532] = UnbiasedRNG[38];
            InitCond[533] = UnbiasedRNG[39];
            InitCond[534] = UnbiasedRNG[40];
            InitCond[535] = UnbiasedRNG[41];
            InitCond[536] = UnbiasedRNG[42];
            InitCond[537] = UnbiasedRNG[43];
            InitCond[538] = UnbiasedRNG[44];
            InitCond[539] = UnbiasedRNG[45];
            InitCond[540] = UnbiasedRNG[46];
            InitCond[541] = UnbiasedRNG[47];
            InitCond[542] = UnbiasedRNG[48];
            InitCond[543] = UnbiasedRNG[49];
            InitCond[544] = UnbiasedRNG[50];
            InitCond[545] = UnbiasedRNG[51];
            InitCond[546] = UnbiasedRNG[52];
            InitCond[547] = UnbiasedRNG[53];
            InitCond[548] = UnbiasedRNG[54];
            InitCond[549] = UnbiasedRNG[55];
            InitCond[550] = UnbiasedRNG[56];
            InitCond[551] = UnbiasedRNG[57];
            InitCond[552] = UnbiasedRNG[58];
            InitCond[553] = UnbiasedRNG[59];
            InitCond[554] = UnbiasedRNG[60];
            InitCond[555] = UnbiasedRNG[61];
            InitCond[556] = UnbiasedRNG[62];
            InitCond[557] = UnbiasedRNG[63];
            InitCond[558] = UnbiasedRNG[64];
            InitCond[559] = UnbiasedRNG[65];
            InitCond[560] = UnbiasedRNG[66];
            InitCond[561] = UnbiasedRNG[67];
            InitCond[562] = UnbiasedRNG[68];
            InitCond[563] = UnbiasedRNG[69];
            InitCond[564] = UnbiasedRNG[70];
            InitCond[565] = UnbiasedRNG[71];
            InitCond[566] = UnbiasedRNG[72];
            InitCond[567] = UnbiasedRNG[73];
            InitCond[568] = UnbiasedRNG[74];
            InitCond[569] = UnbiasedRNG[75];
            InitCond[570] = UnbiasedRNG[76];
            InitCond[571] = UnbiasedRNG[77];
            InitCond[572] = UnbiasedRNG[78];
            InitCond[573] = UnbiasedRNG[79];
            InitCond[574] = UnbiasedRNG[80];
            InitCond[575] = UnbiasedRNG[81];
            InitCond[576] = UnbiasedRNG[82];
            InitCond[577] = UnbiasedRNG[83];
            InitCond[578] = UnbiasedRNG[84];
            InitCond[579] = UnbiasedRNG[85];
            InitCond[580] = UnbiasedRNG[86];
            InitCond[581] = UnbiasedRNG[87];
            InitCond[582] = UnbiasedRNG[88];
            InitCond[583] = UnbiasedRNG[89];
            InitCond[584] = UnbiasedRNG[90];
            InitCond[585] = UnbiasedRNG[91];
            InitCond[586] = UnbiasedRNG[92];
            InitCond[587] = UnbiasedRNG[93];
            InitCond[588] = UnbiasedRNG[94];
            InitCond[589] = UnbiasedRNG[95];
            InitCond[590] = UnbiasedRNG[96];
            InitCond[591] = UnbiasedRNG[97];
            InitCond[592] = UnbiasedRNG[98];
            InitCond[593] = UnbiasedRNG[99];
            InitCond[594] = UnbiasedRNG[100];
            InitCond[595] = UnbiasedRNG[101];
            InitCond[596] = UnbiasedRNG[102];
            InitCond[597] = UnbiasedRNG[103];
            InitCond[598] = UnbiasedRNG[104];
            InitCond[599] = UnbiasedRNG[105];
            InitCond[600] = UnbiasedRNG[106];
            InitCond[601] = UnbiasedRNG[107];
            InitCond[602] = UnbiasedRNG[108];
            InitCond[603] = UnbiasedRNG[109];
            InitCond[604] = UnbiasedRNG[110];
            InitCond[605] = UnbiasedRNG[111];
            InitCond[606] = UnbiasedRNG[112];
            InitCond[607] = UnbiasedRNG[113];
            InitCond[608] = UnbiasedRNG[114];
            InitCond[609] = UnbiasedRNG[115];
            InitCond[610] = UnbiasedRNG[116];
            InitCond[611] = UnbiasedRNG[117];
            InitCond[612] = UnbiasedRNG[118];
            InitCond[613] = UnbiasedRNG[119];
            InitCond[614] = UnbiasedRNG[120];
            InitCond[615] = UnbiasedRNG[121];
            InitCond[616] = UnbiasedRNG[122];
            InitCond[617] = UnbiasedRNG[123];
            InitCond[618] = UnbiasedRNG[124];
            InitCond[619] = UnbiasedRNG[125];
            InitCond[620] = UnbiasedRNG[126];
            InitCond[621] = UnbiasedRNG[127];
            InitCond[622] = UnbiasedRNG[128];
            InitCond[623] = UnbiasedRNG[129];
            InitCond[624] = UnbiasedRNG[130];
            InitCond[625] = UnbiasedRNG[131];
            InitCond[626] = UnbiasedRNG[132];
            InitCond[627] = UnbiasedRNG[133];
            InitCond[628] = UnbiasedRNG[134];
            InitCond[629] = UnbiasedRNG[135];
            InitCond[630] = UnbiasedRNG[136];
            InitCond[631] = UnbiasedRNG[137];
            InitCond[632] = UnbiasedRNG[138];
            InitCond[633] = UnbiasedRNG[139];
            InitCond[634] = UnbiasedRNG[140];
            InitCond[635] = UnbiasedRNG[141];
            InitCond[636] = UnbiasedRNG[142];
            InitCond[637] = UnbiasedRNG[143];
            InitCond[638] = UnbiasedRNG[144];
            InitCond[639] = UnbiasedRNG[145];
            InitCond[640] = UnbiasedRNG[146];
            InitCond[641] = UnbiasedRNG[147];
            InitCond[642] = UnbiasedRNG[148];
            InitCond[643] = UnbiasedRNG[149];
            InitCond[644] = UnbiasedRNG[150];
            InitCond[645] = UnbiasedRNG[151];
            InitCond[646] = UnbiasedRNG[152];
            InitCond[647] = UnbiasedRNG[153];
            InitCond[648] = UnbiasedRNG[154];
            InitCond[649] = UnbiasedRNG[155];
            InitCond[650] = UnbiasedRNG[156];
            InitCond[651] = UnbiasedRNG[157];
            InitCond[652] = UnbiasedRNG[158];
            InitCond[653] = UnbiasedRNG[159];
            InitCond[654] = UnbiasedRNG[160];
            InitCond[655] = UnbiasedRNG[161];
            InitCond[656] = UnbiasedRNG[162];
            InitCond[657] = UnbiasedRNG[163];
            InitCond[658] = UnbiasedRNG[164];
            InitCond[659] = UnbiasedRNG[165];
            InitCond[660] = UnbiasedRNG[166];
            InitCond[661] = UnbiasedRNG[167];
            InitCond[662] = UnbiasedRNG[168];
            InitCond[663] = UnbiasedRNG[169];
            InitCond[664] = UnbiasedRNG[170];
            InitCond[665] = UnbiasedRNG[171];
            InitCond[666] = UnbiasedRNG[172];
            InitCond[667] = UnbiasedRNG[173];
            InitCond[668] = UnbiasedRNG[174];
            InitCond[669] = UnbiasedRNG[175];
            InitCond[670] = UnbiasedRNG[176];
            InitCond[671] = UnbiasedRNG[177];
            InitCond[672] = UnbiasedRNG[178];
            InitCond[673] = UnbiasedRNG[179];
            InitCond[674] = UnbiasedRNG[180];
            InitCond[675] = UnbiasedRNG[181];
            InitCond[676] = UnbiasedRNG[182];
            InitCond[677] = UnbiasedRNG[183];
            InitCond[678] = UnbiasedRNG[184];
            InitCond[679] = UnbiasedRNG[185];
            InitCond[680] = UnbiasedRNG[186];
            InitCond[681] = UnbiasedRNG[187];
            InitCond[682] = UnbiasedRNG[188];
            InitCond[683] = UnbiasedRNG[189];
            InitCond[684] = UnbiasedRNG[190];
            InitCond[685] = UnbiasedRNG[191];
            InitCond[686] = UnbiasedRNG[192];
            InitCond[687] = UnbiasedRNG[193];
            InitCond[688] = UnbiasedRNG[194];
            InitCond[689] = UnbiasedRNG[195];
            InitCond[690] = UnbiasedRNG[196];
            InitCond[691] = UnbiasedRNG[197];
            InitCond[692] = UnbiasedRNG[198];
            InitCond[693] = UnbiasedRNG[199];
            InitCond[694] = UnbiasedRNG[200];
            InitCond[695] = UnbiasedRNG[201];
            InitCond[696] = UnbiasedRNG[202];
            InitCond[697] = UnbiasedRNG[203];
            InitCond[698] = UnbiasedRNG[204];
            InitCond[699] = UnbiasedRNG[205];
            InitCond[700] = UnbiasedRNG[206];
            InitCond[701] = UnbiasedRNG[207];
            InitCond[702] = UnbiasedRNG[208];
            InitCond[703] = UnbiasedRNG[209];
            InitCond[704] = UnbiasedRNG[210];
            InitCond[705] = UnbiasedRNG[211];
            InitCond[706] = UnbiasedRNG[212];
            InitCond[707] = UnbiasedRNG[213];
            InitCond[708] = UnbiasedRNG[214];
            InitCond[709] = UnbiasedRNG[215];
            InitCond[710] = UnbiasedRNG[216];
            InitCond[711] = UnbiasedRNG[217];
            InitCond[712] = UnbiasedRNG[218];
            InitCond[713] = UnbiasedRNG[219];
            InitCond[714] = UnbiasedRNG[220];
            InitCond[715] = UnbiasedRNG[221];
            InitCond[716] = UnbiasedRNG[222];
            InitCond[717] = UnbiasedRNG[223];
            InitCond[718] = UnbiasedRNG[224];
            InitCond[719] = UnbiasedRNG[225];
            InitCond[720] = UnbiasedRNG[226];
            InitCond[721] = UnbiasedRNG[227];
            InitCond[722] = UnbiasedRNG[228];
            InitCond[723] = UnbiasedRNG[229];
            InitCond[724] = UnbiasedRNG[230];
            InitCond[725] = UnbiasedRNG[231];
            InitCond[726] = UnbiasedRNG[232];
            InitCond[727] = UnbiasedRNG[233];
            InitCond[728] = UnbiasedRNG[234];
            InitCond[729] = UnbiasedRNG[235];
            InitCond[730] = UnbiasedRNG[236];
            InitCond[731] = UnbiasedRNG[237];
            InitCond[732] = UnbiasedRNG[238];
            InitCond[733] = UnbiasedRNG[239];
            InitCond[734] = UnbiasedRNG[240];
            InitCond[735] = UnbiasedRNG[241];
            InitCond[736] = UnbiasedRNG[242];
            InitCond[737] = UnbiasedRNG[243];
            InitCond[738] = UnbiasedRNG[244];
            InitCond[739] = UnbiasedRNG[245];
            InitCond[740] = UnbiasedRNG[246];
            InitCond[741] = UnbiasedRNG[247];
            InitCond[742] = UnbiasedRNG[248];
            InitCond[743] = UnbiasedRNG[249];
            InitCond[744] = UnbiasedRNG[250];
            InitCond[745] = UnbiasedRNG[251];
            InitCond[746] = UnbiasedRNG[252];
            InitCond[747] = UnbiasedRNG[253];
            InitCond[748] = UnbiasedRNG[254];
            InitCond[749] = UnbiasedRNG[255];
            InitCond[750] = UnbiasedRNG[256];
            InitCond[751] = UnbiasedRNG[257];
            InitCond[752] = UnbiasedRNG[258];
            InitCond[753] = UnbiasedRNG[259];
            InitCond[754] = UnbiasedRNG[260];
            InitCond[755] = UnbiasedRNG[261];
            InitCond[756] = UnbiasedRNG[262];
            InitCond[757] = UnbiasedRNG[263];
            InitCond[758] = UnbiasedRNG[264];
            InitCond[759] = UnbiasedRNG[265];
            InitCond[760] = UnbiasedRNG[266];
            InitCond[761] = UnbiasedRNG[267];
            InitCond[762] = UnbiasedRNG[268];
            InitCond[763] = UnbiasedRNG[269];
            InitCond[764] = UnbiasedRNG[270];
            InitCond[765] = UnbiasedRNG[271];
            InitCond[766] = UnbiasedRNG[272];
            InitCond[767] = UnbiasedRNG[273];
            InitCond[768] = UnbiasedRNG[274];
            InitCond[769] = UnbiasedRNG[275];
            InitCond[770] = UnbiasedRNG[276];
            InitCond[771] = UnbiasedRNG[277];
            InitCond[772] = UnbiasedRNG[278];
            InitCond[773] = UnbiasedRNG[279];
            InitCond[774] = UnbiasedRNG[280];
            InitCond[775] = UnbiasedRNG[281];
            InitCond[776] = UnbiasedRNG[282];
            InitCond[777] = UnbiasedRNG[283];
            InitCond[778] = UnbiasedRNG[284];
            InitCond[779] = UnbiasedRNG[285];
            InitCond[780] = UnbiasedRNG[286];
            InitCond[781] = UnbiasedRNG[287];
            InitCond[782] = UnbiasedRNG[288];
            InitCond[783] = UnbiasedRNG[289];
            InitCond[784] = UnbiasedRNG[290];
            InitCond[785] = UnbiasedRNG[291];
            InitCond[786] = UnbiasedRNG[292];
            InitCond[787] = UnbiasedRNG[293];
            InitCond[788] = UnbiasedRNG[294];
            InitCond[789] = UnbiasedRNG[295];
            InitCond[790] = UnbiasedRNG[296];
            InitCond[791] = UnbiasedRNG[297];
            InitCond[792] = UnbiasedRNG[298];
            InitCond[793] = UnbiasedRNG[299];
            InitCond[794] = UnbiasedRNG[300];
            InitCond[795] = UnbiasedRNG[301];
            InitCond[796] = UnbiasedRNG[302];
            InitCond[797] = UnbiasedRNG[303];
            InitCond[798] = UnbiasedRNG[304];
            InitCond[799] = UnbiasedRNG[305];
            InitCond[800] = UnbiasedRNG[306];
            InitCond[801] = UnbiasedRNG[307];
            InitCond[802] = UnbiasedRNG[308];
            InitCond[803] = UnbiasedRNG[309];
            InitCond[804] = UnbiasedRNG[310];
            InitCond[805] = UnbiasedRNG[311];
            InitCond[806] = UnbiasedRNG[312];
            InitCond[807] = UnbiasedRNG[313];
            InitCond[808] = UnbiasedRNG[314];
            InitCond[809] = UnbiasedRNG[315];
            InitCond[810] = UnbiasedRNG[316];
            InitCond[811] = UnbiasedRNG[317];
            InitCond[812] = UnbiasedRNG[318];
            InitCond[813] = UnbiasedRNG[319];
            InitCond[814] = UnbiasedRNG[320];
            InitCond[815] = UnbiasedRNG[321];
            InitCond[816] = UnbiasedRNG[322];
            InitCond[817] = UnbiasedRNG[323];
            InitCond[818] = UnbiasedRNG[324];
            InitCond[819] = UnbiasedRNG[325];
            InitCond[820] = UnbiasedRNG[326];
            InitCond[821] = UnbiasedRNG[327];
            InitCond[822] = UnbiasedRNG[328];
            InitCond[823] = UnbiasedRNG[329];
            InitCond[824] = UnbiasedRNG[330];
            InitCond[825] = UnbiasedRNG[331];
            InitCond[826] = UnbiasedRNG[332];
            InitCond[827] = UnbiasedRNG[333];
            InitCond[828] = UnbiasedRNG[334];
            InitCond[829] = UnbiasedRNG[335];
            InitCond[830] = UnbiasedRNG[336];
            InitCond[831] = UnbiasedRNG[337];
            InitCond[832] = UnbiasedRNG[338];
            InitCond[833] = UnbiasedRNG[339];
            InitCond[834] = UnbiasedRNG[340];
            InitCond[835] = UnbiasedRNG[341];
            InitCond[836] = UnbiasedRNG[342];
            InitCond[837] = UnbiasedRNG[343];
            InitCond[838] = UnbiasedRNG[344];
            InitCond[839] = UnbiasedRNG[345];
            InitCond[840] = UnbiasedRNG[346];
            InitCond[841] = UnbiasedRNG[347];
            InitCond[842] = UnbiasedRNG[348];
            InitCond[843] = UnbiasedRNG[349];
            InitCond[844] = UnbiasedRNG[350];
            InitCond[845] = UnbiasedRNG[351];
            InitCond[846] = UnbiasedRNG[352];
            InitCond[847] = UnbiasedRNG[353];
            InitCond[848] = UnbiasedRNG[354];
            InitCond[849] = UnbiasedRNG[355];
            InitCond[850] = UnbiasedRNG[356];
            InitCond[851] = UnbiasedRNG[357];
            InitCond[852] = UnbiasedRNG[358];
            InitCond[853] = UnbiasedRNG[359];
            InitCond[854] = UnbiasedRNG[360];
            InitCond[855] = UnbiasedRNG[361];
            InitCond[856] = UnbiasedRNG[362];
            InitCond[857] = UnbiasedRNG[363];
            InitCond[858] = UnbiasedRNG[364];
            InitCond[859] = UnbiasedRNG[365];
            InitCond[860] = UnbiasedRNG[366];
            InitCond[861] = UnbiasedRNG[367];
            InitCond[862] = UnbiasedRNG[368];
            InitCond[863] = UnbiasedRNG[369];
            InitCond[864] = UnbiasedRNG[370];
            InitCond[865] = UnbiasedRNG[371];
            InitCond[866] = UnbiasedRNG[372];
            InitCond[867] = UnbiasedRNG[373];
            InitCond[868] = UnbiasedRNG[374];
            InitCond[869] = UnbiasedRNG[375];
            InitCond[870] = UnbiasedRNG[376];
            InitCond[871] = UnbiasedRNG[377];
            InitCond[872] = UnbiasedRNG[378];
            InitCond[873] = UnbiasedRNG[379];
            InitCond[874] = UnbiasedRNG[380];
            InitCond[875] = UnbiasedRNG[381];
            InitCond[876] = UnbiasedRNG[382];
            InitCond[877] = UnbiasedRNG[383];
            InitCond[878] = UnbiasedRNG[384];
            InitCond[879] = UnbiasedRNG[385];
            InitCond[880] = UnbiasedRNG[386];
            InitCond[881] = UnbiasedRNG[387];
            InitCond[882] = UnbiasedRNG[388];
            InitCond[883] = UnbiasedRNG[389];
            InitCond[884] = UnbiasedRNG[390];
            InitCond[885] = UnbiasedRNG[391];
            InitCond[886] = UnbiasedRNG[392];
            InitCond[887] = UnbiasedRNG[393];
            InitCond[888] = UnbiasedRNG[394];
            InitCond[889] = UnbiasedRNG[395];
            InitCond[890] = UnbiasedRNG[396];
            InitCond[891] = UnbiasedRNG[397];
            InitCond[892] = UnbiasedRNG[398];
            InitCond[893] = UnbiasedRNG[399];
            InitCond[894] = UnbiasedRNG[400];
            InitCond[895] = UnbiasedRNG[401];
            InitCond[896] = UnbiasedRNG[402];
            InitCond[897] = UnbiasedRNG[403];
            InitCond[898] = UnbiasedRNG[404];
            InitCond[899] = UnbiasedRNG[405];
            InitCond[900] = UnbiasedRNG[406];
            InitCond[901] = UnbiasedRNG[407];
            InitCond[902] = UnbiasedRNG[408];
            InitCond[903] = UnbiasedRNG[409];
            InitCond[904] = UnbiasedRNG[410];
            InitCond[905] = UnbiasedRNG[411];
            InitCond[906] = UnbiasedRNG[412];
            InitCond[907] = UnbiasedRNG[413];
            InitCond[908] = UnbiasedRNG[414];
            InitCond[909] = UnbiasedRNG[415];
            InitCond[910] = UnbiasedRNG[416];
            InitCond[911] = UnbiasedRNG[417];
            InitCond[912] = UnbiasedRNG[418];
            InitCond[913] = UnbiasedRNG[419];
            InitCond[914] = UnbiasedRNG[420];
            InitCond[915] = UnbiasedRNG[421];
            InitCond[916] = UnbiasedRNG[422];
            InitCond[917] = UnbiasedRNG[423];
            InitCond[918] = UnbiasedRNG[424];
            InitCond[919] = UnbiasedRNG[425];
            InitCond[920] = UnbiasedRNG[426];
            InitCond[921] = UnbiasedRNG[427];
            InitCond[922] = UnbiasedRNG[428];
            InitCond[923] = UnbiasedRNG[429];
            InitCond[924] = UnbiasedRNG[430];
            InitCond[925] = UnbiasedRNG[431];
            InitCond[926] = UnbiasedRNG[432];
            InitCond[927] = UnbiasedRNG[433];
            InitCond[928] = UnbiasedRNG[434];
            InitCond[929] = UnbiasedRNG[435];
            InitCond[930] = UnbiasedRNG[436];
            InitCond[931] = UnbiasedRNG[437];
            InitCond[932] = UnbiasedRNG[438];
            InitCond[933] = UnbiasedRNG[439];
            InitCond[934] = UnbiasedRNG[440];
            InitCond[935] = UnbiasedRNG[441];
            InitCond[936] = UnbiasedRNG[442];
            InitCond[937] = UnbiasedRNG[443];
            InitCond[938] = UnbiasedRNG[444];
            InitCond[939] = UnbiasedRNG[445];
            InitCond[940] = UnbiasedRNG[446];
            InitCond[941] = UnbiasedRNG[447];
            InitCond[942] = UnbiasedRNG[448];
            InitCond[943] = UnbiasedRNG[449];
            InitCond[944] = UnbiasedRNG[450];
            InitCond[945] = UnbiasedRNG[451];
            InitCond[946] = UnbiasedRNG[452];
            InitCond[947] = UnbiasedRNG[453];
            InitCond[948] = UnbiasedRNG[454];
            InitCond[949] = UnbiasedRNG[455];
            InitCond[950] = UnbiasedRNG[456];
            InitCond[951] = UnbiasedRNG[457];
            InitCond[952] = UnbiasedRNG[458];
            InitCond[953] = UnbiasedRNG[459];
            InitCond[954] = UnbiasedRNG[460];
            InitCond[955] = UnbiasedRNG[461];
            InitCond[956] = UnbiasedRNG[462];
            InitCond[957] = UnbiasedRNG[463];
            InitCond[958] = UnbiasedRNG[464];
            InitCond[959] = UnbiasedRNG[465];
            InitCond[960] = UnbiasedRNG[466];
            InitCond[961] = UnbiasedRNG[467];
            InitCond[962] = UnbiasedRNG[468];
            InitCond[963] = UnbiasedRNG[469];
            InitCond[964] = UnbiasedRNG[470];
            InitCond[965] = UnbiasedRNG[471];
            InitCond[966] = UnbiasedRNG[472];
            InitCond[967] = UnbiasedRNG[473];
            InitCond[968] = UnbiasedRNG[474];
            InitCond[969] = UnbiasedRNG[475];
            InitCond[970] = UnbiasedRNG[476];
            InitCond[971] = UnbiasedRNG[477];
            InitCond[972] = UnbiasedRNG[478];
            InitCond[973] = UnbiasedRNG[479];
            InitCond[974] = UnbiasedRNG[480];
            InitCond[975] = UnbiasedRNG[481];
            InitCond[976] = UnbiasedRNG[482];
            InitCond[977] = UnbiasedRNG[483];
            InitCond[978] = UnbiasedRNG[484];
            InitCond[979] = UnbiasedRNG[485];
            InitCond[980] = UnbiasedRNG[486];
            InitCond[981] = UnbiasedRNG[487];
            InitCond[982] = UnbiasedRNG[488];
            InitCond[983] = UnbiasedRNG[489];
            InitCond[984] = UnbiasedRNG[490];
            InitCond[985] = UnbiasedRNG[491];
            InitCond[986] = UnbiasedRNG[492];
            InitCond[987] = UnbiasedRNG[493];
        end
        else if (counter == 3) begin
            InitCond[988] = UnbiasedRNG[0];
            InitCond[989] = UnbiasedRNG[1];
            InitCond[990] = UnbiasedRNG[2];
            InitCond[991] = UnbiasedRNG[3];
            InitCond[992] = UnbiasedRNG[4];
            InitCond[993] = UnbiasedRNG[5];
            InitCond[994] = UnbiasedRNG[6];
            InitCond[995] = UnbiasedRNG[7];
            InitCond[996] = UnbiasedRNG[8];
            InitCond[997] = UnbiasedRNG[9];
            InitCond[998] = UnbiasedRNG[10];
            InitCond[999] = UnbiasedRNG[11];
            InitCond[1000] = UnbiasedRNG[12];
            InitCond[1001] = UnbiasedRNG[13];
            InitCond[1002] = UnbiasedRNG[14];
            InitCond[1003] = UnbiasedRNG[15];
            InitCond[1004] = UnbiasedRNG[16];
            InitCond[1005] = UnbiasedRNG[17];
            InitCond[1006] = UnbiasedRNG[18];
            InitCond[1007] = UnbiasedRNG[19];
            InitCond[1008] = UnbiasedRNG[20];
            InitCond[1009] = UnbiasedRNG[21];
            InitCond[1010] = UnbiasedRNG[22];
            InitCond[1011] = UnbiasedRNG[23];
            InitCond[1012] = UnbiasedRNG[24];
            InitCond[1013] = UnbiasedRNG[25];
            InitCond[1014] = UnbiasedRNG[26];
            InitCond[1015] = UnbiasedRNG[27];
            InitCond[1016] = UnbiasedRNG[28];
            InitCond[1017] = UnbiasedRNG[29];
            InitCond[1018] = UnbiasedRNG[30];
            InitCond[1019] = UnbiasedRNG[31];
            InitCond[1020] = UnbiasedRNG[32];
            InitCond[1021] = UnbiasedRNG[33];
            InitCond[1022] = UnbiasedRNG[34];
            InitCond[1023] = UnbiasedRNG[35];
            InitCond[1024] = UnbiasedRNG[36];
            InitCond[1025] = UnbiasedRNG[37];
            InitCond[1026] = UnbiasedRNG[38];
            InitCond[1027] = UnbiasedRNG[39];
            InitCond[1028] = UnbiasedRNG[40];
            InitCond[1029] = UnbiasedRNG[41];
            InitCond[1030] = UnbiasedRNG[42];
            InitCond[1031] = UnbiasedRNG[43];
            InitCond[1032] = UnbiasedRNG[44];
            InitCond[1033] = UnbiasedRNG[45];
            InitCond[1034] = UnbiasedRNG[46];
            InitCond[1035] = UnbiasedRNG[47];
            InitCond[1036] = UnbiasedRNG[48];
            InitCond[1037] = UnbiasedRNG[49];
            InitCond[1038] = UnbiasedRNG[50];
            InitCond[1039] = UnbiasedRNG[51];
            InitCond[1040] = UnbiasedRNG[52];
            InitCond[1041] = UnbiasedRNG[53];
            InitCond[1042] = UnbiasedRNG[54];
            InitCond[1043] = UnbiasedRNG[55];
            InitCond[1044] = UnbiasedRNG[56];
            InitCond[1045] = UnbiasedRNG[57];
            InitCond[1046] = UnbiasedRNG[58];
            InitCond[1047] = UnbiasedRNG[59];
            InitCond[1048] = UnbiasedRNG[60];
            InitCond[1049] = UnbiasedRNG[61];
            InitCond[1050] = UnbiasedRNG[62];
            InitCond[1051] = UnbiasedRNG[63];
            InitCond[1052] = UnbiasedRNG[64];
            InitCond[1053] = UnbiasedRNG[65];
            InitCond[1054] = UnbiasedRNG[66];
            InitCond[1055] = UnbiasedRNG[67];
            InitCond[1056] = UnbiasedRNG[68];
            InitCond[1057] = UnbiasedRNG[69];
            InitCond[1058] = UnbiasedRNG[70];
            InitCond[1059] = UnbiasedRNG[71];
            InitCond[1060] = UnbiasedRNG[72];
            InitCond[1061] = UnbiasedRNG[73];
            InitCond[1062] = UnbiasedRNG[74];
            InitCond[1063] = UnbiasedRNG[75];
            InitCond[1064] = UnbiasedRNG[76];
            InitCond[1065] = UnbiasedRNG[77];
            InitCond[1066] = UnbiasedRNG[78];
            InitCond[1067] = UnbiasedRNG[79];
            InitCond[1068] = UnbiasedRNG[80];
            InitCond[1069] = UnbiasedRNG[81];
            InitCond[1070] = UnbiasedRNG[82];
            InitCond[1071] = UnbiasedRNG[83];
            InitCond[1072] = UnbiasedRNG[84];
            InitCond[1073] = UnbiasedRNG[85];
            InitCond[1074] = UnbiasedRNG[86];
            InitCond[1075] = UnbiasedRNG[87];
            InitCond[1076] = UnbiasedRNG[88];
            InitCond[1077] = UnbiasedRNG[89];
            InitCond[1078] = UnbiasedRNG[90];
            InitCond[1079] = UnbiasedRNG[91];
            InitCond[1080] = UnbiasedRNG[92];
            InitCond[1081] = UnbiasedRNG[93];
            InitCond[1082] = UnbiasedRNG[94];
            InitCond[1083] = UnbiasedRNG[95];
            InitCond[1084] = UnbiasedRNG[96];
            InitCond[1085] = UnbiasedRNG[97];
            InitCond[1086] = UnbiasedRNG[98];
            InitCond[1087] = UnbiasedRNG[99];
            InitCond[1088] = UnbiasedRNG[100];
            InitCond[1089] = UnbiasedRNG[101];
            InitCond[1090] = UnbiasedRNG[102];
            InitCond[1091] = UnbiasedRNG[103];
            InitCond[1092] = UnbiasedRNG[104];
            InitCond[1093] = UnbiasedRNG[105];
            InitCond[1094] = UnbiasedRNG[106];
            InitCond[1095] = UnbiasedRNG[107];
            InitCond[1096] = UnbiasedRNG[108];
            InitCond[1097] = UnbiasedRNG[109];
            InitCond[1098] = UnbiasedRNG[110];
            InitCond[1099] = UnbiasedRNG[111];
            InitCond[1100] = UnbiasedRNG[112];
            InitCond[1101] = UnbiasedRNG[113];
            InitCond[1102] = UnbiasedRNG[114];
            InitCond[1103] = UnbiasedRNG[115];
            InitCond[1104] = UnbiasedRNG[116];
            InitCond[1105] = UnbiasedRNG[117];
            InitCond[1106] = UnbiasedRNG[118];
            InitCond[1107] = UnbiasedRNG[119];
            InitCond[1108] = UnbiasedRNG[120];
            InitCond[1109] = UnbiasedRNG[121];
            InitCond[1110] = UnbiasedRNG[122];
            InitCond[1111] = UnbiasedRNG[123];
            InitCond[1112] = UnbiasedRNG[124];
            InitCond[1113] = UnbiasedRNG[125];
            InitCond[1114] = UnbiasedRNG[126];
            InitCond[1115] = UnbiasedRNG[127];
            InitCond[1116] = UnbiasedRNG[128];
            InitCond[1117] = UnbiasedRNG[129];
            InitCond[1118] = UnbiasedRNG[130];
            InitCond[1119] = UnbiasedRNG[131];
            InitCond[1120] = UnbiasedRNG[132];
            InitCond[1121] = UnbiasedRNG[133];
            InitCond[1122] = UnbiasedRNG[134];
            InitCond[1123] = UnbiasedRNG[135];
            InitCond[1124] = UnbiasedRNG[136];
            InitCond[1125] = UnbiasedRNG[137];
            InitCond[1126] = UnbiasedRNG[138];
            InitCond[1127] = UnbiasedRNG[139];
            InitCond[1128] = UnbiasedRNG[140];
            InitCond[1129] = UnbiasedRNG[141];
            InitCond[1130] = UnbiasedRNG[142];
            InitCond[1131] = UnbiasedRNG[143];
            InitCond[1132] = UnbiasedRNG[144];
            InitCond[1133] = UnbiasedRNG[145];
            InitCond[1134] = UnbiasedRNG[146];
            InitCond[1135] = UnbiasedRNG[147];
            InitCond[1136] = UnbiasedRNG[148];
            InitCond[1137] = UnbiasedRNG[149];
            InitCond[1138] = UnbiasedRNG[150];
            InitCond[1139] = UnbiasedRNG[151];
            InitCond[1140] = UnbiasedRNG[152];
            InitCond[1141] = UnbiasedRNG[153];
            InitCond[1142] = UnbiasedRNG[154];
            InitCond[1143] = UnbiasedRNG[155];
            InitCond[1144] = UnbiasedRNG[156];
            InitCond[1145] = UnbiasedRNG[157];
            InitCond[1146] = UnbiasedRNG[158];
            InitCond[1147] = UnbiasedRNG[159];
            InitCond[1148] = UnbiasedRNG[160];
            InitCond[1149] = UnbiasedRNG[161];
            InitCond[1150] = UnbiasedRNG[162];
            InitCond[1151] = UnbiasedRNG[163];
        end
        else if (counter==5)
            run = 1'b1;
        counter = counter+38'b1;
        solution = {m[11],m[10],m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[23],m[22],m[21],m[20],m[19],m[18],m[17],m[16],m[15],m[14],m[13],m[12]};
    end else begin 
        counter = 38'b0;
        failure = 1'b1;
        run = 1'b0;
    end
end

//To measure on only the last step using ILA:
always @(negedge sample_clk) begin
    if (solution_flag)
        solution_flag = 1'b0;
    else if ((run & (solution == solution_check)) | failure)
        solution_flag = 1'b1;
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = run?((((m[24]&~m[25]&~m[26])|(~m[24]&m[25]&~m[26])|(~m[24]&~m[25]&m[26]))&BiasedRNG[0])|(((m[24]&m[25]&~m[26])|(m[24]&~m[25]&m[26])|(~m[24]&m[25]&m[26]))&~BiasedRNG[0])|((m[24]&m[25]&m[26]))):InitCond[0];
    m[1] = run?((((m[27]&~m[28]&~m[29])|(~m[27]&m[28]&~m[29])|(~m[27]&~m[28]&m[29]))&BiasedRNG[1])|(((m[27]&m[28]&~m[29])|(m[27]&~m[28]&m[29])|(~m[27]&m[28]&m[29]))&~BiasedRNG[1])|((m[27]&m[28]&m[29]))):InitCond[1];
    m[2] = run?((((m[30]&~m[31]&~m[32])|(~m[30]&m[31]&~m[32])|(~m[30]&~m[31]&m[32]))&BiasedRNG[2])|(((m[30]&m[31]&~m[32])|(m[30]&~m[31]&m[32])|(~m[30]&m[31]&m[32]))&~BiasedRNG[2])|((m[30]&m[31]&m[32]))):InitCond[2];
    m[3] = run?((((m[33]&~m[34]&~m[35])|(~m[33]&m[34]&~m[35])|(~m[33]&~m[34]&m[35]))&BiasedRNG[3])|(((m[33]&m[34]&~m[35])|(m[33]&~m[34]&m[35])|(~m[33]&m[34]&m[35]))&~BiasedRNG[3])|((m[33]&m[34]&m[35]))):InitCond[3];
    m[4] = run?((((m[36]&~m[37]&~m[38])|(~m[36]&m[37]&~m[38])|(~m[36]&~m[37]&m[38]))&BiasedRNG[4])|(((m[36]&m[37]&~m[38])|(m[36]&~m[37]&m[38])|(~m[36]&m[37]&m[38]))&~BiasedRNG[4])|((m[36]&m[37]&m[38]))):InitCond[4];
    m[5] = run?((((m[39]&~m[40]&~m[41])|(~m[39]&m[40]&~m[41])|(~m[39]&~m[40]&m[41]))&BiasedRNG[5])|(((m[39]&m[40]&~m[41])|(m[39]&~m[40]&m[41])|(~m[39]&m[40]&m[41]))&~BiasedRNG[5])|((m[39]&m[40]&m[41]))):InitCond[5];
    m[6] = run?((((m[42]&~m[43]&~m[44])|(~m[42]&m[43]&~m[44])|(~m[42]&~m[43]&m[44]))&BiasedRNG[6])|(((m[42]&m[43]&~m[44])|(m[42]&~m[43]&m[44])|(~m[42]&m[43]&m[44]))&~BiasedRNG[6])|((m[42]&m[43]&m[44]))):InitCond[6];
    m[7] = run?((((m[45]&~m[46]&~m[47])|(~m[45]&m[46]&~m[47])|(~m[45]&~m[46]&m[47]))&BiasedRNG[7])|(((m[45]&m[46]&~m[47])|(m[45]&~m[46]&m[47])|(~m[45]&m[46]&m[47]))&~BiasedRNG[7])|((m[45]&m[46]&m[47]))):InitCond[7];
    m[8] = run?((((m[48]&~m[49]&~m[50])|(~m[48]&m[49]&~m[50])|(~m[48]&~m[49]&m[50]))&BiasedRNG[8])|(((m[48]&m[49]&~m[50])|(m[48]&~m[49]&m[50])|(~m[48]&m[49]&m[50]))&~BiasedRNG[8])|((m[48]&m[49]&m[50]))):InitCond[8];
    m[9] = run?((((m[51]&~m[52]&~m[53])|(~m[51]&m[52]&~m[53])|(~m[51]&~m[52]&m[53]))&BiasedRNG[9])|(((m[51]&m[52]&~m[53])|(m[51]&~m[52]&m[53])|(~m[51]&m[52]&m[53]))&~BiasedRNG[9])|((m[51]&m[52]&m[53]))):InitCond[9];
    m[10] = run?((((m[54]&~m[55]&~m[56])|(~m[54]&m[55]&~m[56])|(~m[54]&~m[55]&m[56]))&BiasedRNG[10])|(((m[54]&m[55]&~m[56])|(m[54]&~m[55]&m[56])|(~m[54]&m[55]&m[56]))&~BiasedRNG[10])|((m[54]&m[55]&m[56]))):InitCond[10];
    m[11] = run?((((m[57]&~m[58]&~m[59])|(~m[57]&m[58]&~m[59])|(~m[57]&~m[58]&m[59]))&BiasedRNG[11])|(((m[57]&m[58]&~m[59])|(m[57]&~m[58]&m[59])|(~m[57]&m[58]&m[59]))&~BiasedRNG[11])|((m[57]&m[58]&m[59]))):InitCond[11];
    m[12] = run?((((m[60]&~m[61]&~m[62])|(~m[60]&m[61]&~m[62])|(~m[60]&~m[61]&m[62]))&BiasedRNG[12])|(((m[60]&m[61]&~m[62])|(m[60]&~m[61]&m[62])|(~m[60]&m[61]&m[62]))&~BiasedRNG[12])|((m[60]&m[61]&m[62]))):InitCond[12];
    m[13] = run?((((m[63]&~m[64]&~m[65])|(~m[63]&m[64]&~m[65])|(~m[63]&~m[64]&m[65]))&BiasedRNG[13])|(((m[63]&m[64]&~m[65])|(m[63]&~m[64]&m[65])|(~m[63]&m[64]&m[65]))&~BiasedRNG[13])|((m[63]&m[64]&m[65]))):InitCond[13];
    m[14] = run?((((m[66]&~m[67]&~m[68])|(~m[66]&m[67]&~m[68])|(~m[66]&~m[67]&m[68]))&BiasedRNG[14])|(((m[66]&m[67]&~m[68])|(m[66]&~m[67]&m[68])|(~m[66]&m[67]&m[68]))&~BiasedRNG[14])|((m[66]&m[67]&m[68]))):InitCond[14];
    m[15] = run?((((m[69]&~m[70]&~m[71])|(~m[69]&m[70]&~m[71])|(~m[69]&~m[70]&m[71]))&BiasedRNG[15])|(((m[69]&m[70]&~m[71])|(m[69]&~m[70]&m[71])|(~m[69]&m[70]&m[71]))&~BiasedRNG[15])|((m[69]&m[70]&m[71]))):InitCond[15];
    m[16] = run?((((m[72]&~m[73]&~m[74])|(~m[72]&m[73]&~m[74])|(~m[72]&~m[73]&m[74]))&BiasedRNG[16])|(((m[72]&m[73]&~m[74])|(m[72]&~m[73]&m[74])|(~m[72]&m[73]&m[74]))&~BiasedRNG[16])|((m[72]&m[73]&m[74]))):InitCond[16];
    m[17] = run?((((m[75]&~m[76]&~m[77])|(~m[75]&m[76]&~m[77])|(~m[75]&~m[76]&m[77]))&BiasedRNG[17])|(((m[75]&m[76]&~m[77])|(m[75]&~m[76]&m[77])|(~m[75]&m[76]&m[77]))&~BiasedRNG[17])|((m[75]&m[76]&m[77]))):InitCond[17];
    m[18] = run?((((m[78]&~m[79]&~m[80])|(~m[78]&m[79]&~m[80])|(~m[78]&~m[79]&m[80]))&BiasedRNG[18])|(((m[78]&m[79]&~m[80])|(m[78]&~m[79]&m[80])|(~m[78]&m[79]&m[80]))&~BiasedRNG[18])|((m[78]&m[79]&m[80]))):InitCond[18];
    m[19] = run?((((m[81]&~m[82]&~m[83])|(~m[81]&m[82]&~m[83])|(~m[81]&~m[82]&m[83]))&BiasedRNG[19])|(((m[81]&m[82]&~m[83])|(m[81]&~m[82]&m[83])|(~m[81]&m[82]&m[83]))&~BiasedRNG[19])|((m[81]&m[82]&m[83]))):InitCond[19];
    m[20] = run?((((m[84]&~m[85]&~m[86])|(~m[84]&m[85]&~m[86])|(~m[84]&~m[85]&m[86]))&BiasedRNG[20])|(((m[84]&m[85]&~m[86])|(m[84]&~m[85]&m[86])|(~m[84]&m[85]&m[86]))&~BiasedRNG[20])|((m[84]&m[85]&m[86]))):InitCond[20];
    m[21] = run?((((m[87]&~m[88]&~m[89])|(~m[87]&m[88]&~m[89])|(~m[87]&~m[88]&m[89]))&BiasedRNG[21])|(((m[87]&m[88]&~m[89])|(m[87]&~m[88]&m[89])|(~m[87]&m[88]&m[89]))&~BiasedRNG[21])|((m[87]&m[88]&m[89]))):InitCond[21];
    m[22] = run?((((m[90]&~m[91]&~m[92])|(~m[90]&m[91]&~m[92])|(~m[90]&~m[91]&m[92]))&BiasedRNG[22])|(((m[90]&m[91]&~m[92])|(m[90]&~m[91]&m[92])|(~m[90]&m[91]&m[92]))&~BiasedRNG[22])|((m[90]&m[91]&m[92]))):InitCond[22];
    m[23] = run?((((m[93]&~m[94]&~m[95])|(~m[93]&m[94]&~m[95])|(~m[93]&~m[94]&m[95]))&BiasedRNG[23])|(((m[93]&m[94]&~m[95])|(m[93]&~m[94]&m[95])|(~m[93]&m[94]&m[95]))&~BiasedRNG[23])|((m[93]&m[94]&m[95]))):InitCond[23];
    m[96] = run?((((~m[24]&~m[240]&~m[384])|(m[24]&m[240]&~m[384]))&BiasedRNG[24])|(((m[24]&~m[240]&~m[384])|(~m[24]&m[240]&m[384]))&~BiasedRNG[24])|((~m[24]&~m[240]&m[384])|(m[24]&~m[240]&m[384])|(m[24]&m[240]&m[384]))):InitCond[24];
    m[97] = run?((((~m[24]&~m[252]&~m[396])|(m[24]&m[252]&~m[396]))&BiasedRNG[25])|(((m[24]&~m[252]&~m[396])|(~m[24]&m[252]&m[396]))&~BiasedRNG[25])|((~m[24]&~m[252]&m[396])|(m[24]&~m[252]&m[396])|(m[24]&m[252]&m[396]))):InitCond[25];
    m[98] = run?((((~m[24]&~m[264]&~m[408])|(m[24]&m[264]&~m[408]))&BiasedRNG[26])|(((m[24]&~m[264]&~m[408])|(~m[24]&m[264]&m[408]))&~BiasedRNG[26])|((~m[24]&~m[264]&m[408])|(m[24]&~m[264]&m[408])|(m[24]&m[264]&m[408]))):InitCond[26];
    m[99] = run?((((~m[24]&~m[276]&~m[420])|(m[24]&m[276]&~m[420]))&BiasedRNG[27])|(((m[24]&~m[276]&~m[420])|(~m[24]&m[276]&m[420]))&~BiasedRNG[27])|((~m[24]&~m[276]&m[420])|(m[24]&~m[276]&m[420])|(m[24]&m[276]&m[420]))):InitCond[27];
    m[100] = run?((((~m[25]&~m[288]&~m[432])|(m[25]&m[288]&~m[432]))&BiasedRNG[28])|(((m[25]&~m[288]&~m[432])|(~m[25]&m[288]&m[432]))&~BiasedRNG[28])|((~m[25]&~m[288]&m[432])|(m[25]&~m[288]&m[432])|(m[25]&m[288]&m[432]))):InitCond[28];
    m[101] = run?((((~m[25]&~m[300]&~m[444])|(m[25]&m[300]&~m[444]))&BiasedRNG[29])|(((m[25]&~m[300]&~m[444])|(~m[25]&m[300]&m[444]))&~BiasedRNG[29])|((~m[25]&~m[300]&m[444])|(m[25]&~m[300]&m[444])|(m[25]&m[300]&m[444]))):InitCond[29];
    m[102] = run?((((~m[25]&~m[312]&~m[456])|(m[25]&m[312]&~m[456]))&BiasedRNG[30])|(((m[25]&~m[312]&~m[456])|(~m[25]&m[312]&m[456]))&~BiasedRNG[30])|((~m[25]&~m[312]&m[456])|(m[25]&~m[312]&m[456])|(m[25]&m[312]&m[456]))):InitCond[30];
    m[103] = run?((((~m[25]&~m[324]&~m[468])|(m[25]&m[324]&~m[468]))&BiasedRNG[31])|(((m[25]&~m[324]&~m[468])|(~m[25]&m[324]&m[468]))&~BiasedRNG[31])|((~m[25]&~m[324]&m[468])|(m[25]&~m[324]&m[468])|(m[25]&m[324]&m[468]))):InitCond[31];
    m[104] = run?((((~m[26]&~m[336]&~m[480])|(m[26]&m[336]&~m[480]))&BiasedRNG[32])|(((m[26]&~m[336]&~m[480])|(~m[26]&m[336]&m[480]))&~BiasedRNG[32])|((~m[26]&~m[336]&m[480])|(m[26]&~m[336]&m[480])|(m[26]&m[336]&m[480]))):InitCond[32];
    m[105] = run?((((~m[26]&~m[348]&~m[492])|(m[26]&m[348]&~m[492]))&BiasedRNG[33])|(((m[26]&~m[348]&~m[492])|(~m[26]&m[348]&m[492]))&~BiasedRNG[33])|((~m[26]&~m[348]&m[492])|(m[26]&~m[348]&m[492])|(m[26]&m[348]&m[492]))):InitCond[33];
    m[106] = run?((((~m[26]&~m[360]&~m[504])|(m[26]&m[360]&~m[504]))&BiasedRNG[34])|(((m[26]&~m[360]&~m[504])|(~m[26]&m[360]&m[504]))&~BiasedRNG[34])|((~m[26]&~m[360]&m[504])|(m[26]&~m[360]&m[504])|(m[26]&m[360]&m[504]))):InitCond[34];
    m[107] = run?((((~m[26]&~m[372]&~m[516])|(m[26]&m[372]&~m[516]))&BiasedRNG[35])|(((m[26]&~m[372]&~m[516])|(~m[26]&m[372]&m[516]))&~BiasedRNG[35])|((~m[26]&~m[372]&m[516])|(m[26]&~m[372]&m[516])|(m[26]&m[372]&m[516]))):InitCond[35];
    m[108] = run?((((~m[27]&~m[241]&~m[385])|(m[27]&m[241]&~m[385]))&BiasedRNG[36])|(((m[27]&~m[241]&~m[385])|(~m[27]&m[241]&m[385]))&~BiasedRNG[36])|((~m[27]&~m[241]&m[385])|(m[27]&~m[241]&m[385])|(m[27]&m[241]&m[385]))):InitCond[36];
    m[109] = run?((((~m[27]&~m[253]&~m[397])|(m[27]&m[253]&~m[397]))&BiasedRNG[37])|(((m[27]&~m[253]&~m[397])|(~m[27]&m[253]&m[397]))&~BiasedRNG[37])|((~m[27]&~m[253]&m[397])|(m[27]&~m[253]&m[397])|(m[27]&m[253]&m[397]))):InitCond[37];
    m[110] = run?((((~m[27]&~m[265]&~m[409])|(m[27]&m[265]&~m[409]))&BiasedRNG[38])|(((m[27]&~m[265]&~m[409])|(~m[27]&m[265]&m[409]))&~BiasedRNG[38])|((~m[27]&~m[265]&m[409])|(m[27]&~m[265]&m[409])|(m[27]&m[265]&m[409]))):InitCond[38];
    m[111] = run?((((~m[27]&~m[277]&~m[421])|(m[27]&m[277]&~m[421]))&BiasedRNG[39])|(((m[27]&~m[277]&~m[421])|(~m[27]&m[277]&m[421]))&~BiasedRNG[39])|((~m[27]&~m[277]&m[421])|(m[27]&~m[277]&m[421])|(m[27]&m[277]&m[421]))):InitCond[39];
    m[112] = run?((((~m[28]&~m[289]&~m[433])|(m[28]&m[289]&~m[433]))&BiasedRNG[40])|(((m[28]&~m[289]&~m[433])|(~m[28]&m[289]&m[433]))&~BiasedRNG[40])|((~m[28]&~m[289]&m[433])|(m[28]&~m[289]&m[433])|(m[28]&m[289]&m[433]))):InitCond[40];
    m[113] = run?((((~m[28]&~m[301]&~m[445])|(m[28]&m[301]&~m[445]))&BiasedRNG[41])|(((m[28]&~m[301]&~m[445])|(~m[28]&m[301]&m[445]))&~BiasedRNG[41])|((~m[28]&~m[301]&m[445])|(m[28]&~m[301]&m[445])|(m[28]&m[301]&m[445]))):InitCond[41];
    m[114] = run?((((~m[28]&~m[313]&~m[457])|(m[28]&m[313]&~m[457]))&BiasedRNG[42])|(((m[28]&~m[313]&~m[457])|(~m[28]&m[313]&m[457]))&~BiasedRNG[42])|((~m[28]&~m[313]&m[457])|(m[28]&~m[313]&m[457])|(m[28]&m[313]&m[457]))):InitCond[42];
    m[115] = run?((((~m[28]&~m[325]&~m[469])|(m[28]&m[325]&~m[469]))&BiasedRNG[43])|(((m[28]&~m[325]&~m[469])|(~m[28]&m[325]&m[469]))&~BiasedRNG[43])|((~m[28]&~m[325]&m[469])|(m[28]&~m[325]&m[469])|(m[28]&m[325]&m[469]))):InitCond[43];
    m[116] = run?((((~m[29]&~m[337]&~m[481])|(m[29]&m[337]&~m[481]))&BiasedRNG[44])|(((m[29]&~m[337]&~m[481])|(~m[29]&m[337]&m[481]))&~BiasedRNG[44])|((~m[29]&~m[337]&m[481])|(m[29]&~m[337]&m[481])|(m[29]&m[337]&m[481]))):InitCond[44];
    m[117] = run?((((~m[29]&~m[349]&~m[493])|(m[29]&m[349]&~m[493]))&BiasedRNG[45])|(((m[29]&~m[349]&~m[493])|(~m[29]&m[349]&m[493]))&~BiasedRNG[45])|((~m[29]&~m[349]&m[493])|(m[29]&~m[349]&m[493])|(m[29]&m[349]&m[493]))):InitCond[45];
    m[118] = run?((((~m[29]&~m[361]&~m[505])|(m[29]&m[361]&~m[505]))&BiasedRNG[46])|(((m[29]&~m[361]&~m[505])|(~m[29]&m[361]&m[505]))&~BiasedRNG[46])|((~m[29]&~m[361]&m[505])|(m[29]&~m[361]&m[505])|(m[29]&m[361]&m[505]))):InitCond[46];
    m[119] = run?((((~m[29]&~m[373]&~m[517])|(m[29]&m[373]&~m[517]))&BiasedRNG[47])|(((m[29]&~m[373]&~m[517])|(~m[29]&m[373]&m[517]))&~BiasedRNG[47])|((~m[29]&~m[373]&m[517])|(m[29]&~m[373]&m[517])|(m[29]&m[373]&m[517]))):InitCond[47];
    m[120] = run?((((~m[30]&~m[242]&~m[386])|(m[30]&m[242]&~m[386]))&BiasedRNG[48])|(((m[30]&~m[242]&~m[386])|(~m[30]&m[242]&m[386]))&~BiasedRNG[48])|((~m[30]&~m[242]&m[386])|(m[30]&~m[242]&m[386])|(m[30]&m[242]&m[386]))):InitCond[48];
    m[121] = run?((((~m[30]&~m[254]&~m[398])|(m[30]&m[254]&~m[398]))&BiasedRNG[49])|(((m[30]&~m[254]&~m[398])|(~m[30]&m[254]&m[398]))&~BiasedRNG[49])|((~m[30]&~m[254]&m[398])|(m[30]&~m[254]&m[398])|(m[30]&m[254]&m[398]))):InitCond[49];
    m[122] = run?((((~m[30]&~m[266]&~m[410])|(m[30]&m[266]&~m[410]))&BiasedRNG[50])|(((m[30]&~m[266]&~m[410])|(~m[30]&m[266]&m[410]))&~BiasedRNG[50])|((~m[30]&~m[266]&m[410])|(m[30]&~m[266]&m[410])|(m[30]&m[266]&m[410]))):InitCond[50];
    m[123] = run?((((~m[30]&~m[278]&~m[422])|(m[30]&m[278]&~m[422]))&BiasedRNG[51])|(((m[30]&~m[278]&~m[422])|(~m[30]&m[278]&m[422]))&~BiasedRNG[51])|((~m[30]&~m[278]&m[422])|(m[30]&~m[278]&m[422])|(m[30]&m[278]&m[422]))):InitCond[51];
    m[124] = run?((((~m[31]&~m[290]&~m[434])|(m[31]&m[290]&~m[434]))&BiasedRNG[52])|(((m[31]&~m[290]&~m[434])|(~m[31]&m[290]&m[434]))&~BiasedRNG[52])|((~m[31]&~m[290]&m[434])|(m[31]&~m[290]&m[434])|(m[31]&m[290]&m[434]))):InitCond[52];
    m[125] = run?((((~m[31]&~m[302]&~m[446])|(m[31]&m[302]&~m[446]))&BiasedRNG[53])|(((m[31]&~m[302]&~m[446])|(~m[31]&m[302]&m[446]))&~BiasedRNG[53])|((~m[31]&~m[302]&m[446])|(m[31]&~m[302]&m[446])|(m[31]&m[302]&m[446]))):InitCond[53];
    m[126] = run?((((~m[31]&~m[314]&~m[458])|(m[31]&m[314]&~m[458]))&BiasedRNG[54])|(((m[31]&~m[314]&~m[458])|(~m[31]&m[314]&m[458]))&~BiasedRNG[54])|((~m[31]&~m[314]&m[458])|(m[31]&~m[314]&m[458])|(m[31]&m[314]&m[458]))):InitCond[54];
    m[127] = run?((((~m[31]&~m[326]&~m[470])|(m[31]&m[326]&~m[470]))&BiasedRNG[55])|(((m[31]&~m[326]&~m[470])|(~m[31]&m[326]&m[470]))&~BiasedRNG[55])|((~m[31]&~m[326]&m[470])|(m[31]&~m[326]&m[470])|(m[31]&m[326]&m[470]))):InitCond[55];
    m[128] = run?((((~m[32]&~m[338]&~m[482])|(m[32]&m[338]&~m[482]))&BiasedRNG[56])|(((m[32]&~m[338]&~m[482])|(~m[32]&m[338]&m[482]))&~BiasedRNG[56])|((~m[32]&~m[338]&m[482])|(m[32]&~m[338]&m[482])|(m[32]&m[338]&m[482]))):InitCond[56];
    m[129] = run?((((~m[32]&~m[350]&~m[494])|(m[32]&m[350]&~m[494]))&BiasedRNG[57])|(((m[32]&~m[350]&~m[494])|(~m[32]&m[350]&m[494]))&~BiasedRNG[57])|((~m[32]&~m[350]&m[494])|(m[32]&~m[350]&m[494])|(m[32]&m[350]&m[494]))):InitCond[57];
    m[130] = run?((((~m[32]&~m[362]&~m[506])|(m[32]&m[362]&~m[506]))&BiasedRNG[58])|(((m[32]&~m[362]&~m[506])|(~m[32]&m[362]&m[506]))&~BiasedRNG[58])|((~m[32]&~m[362]&m[506])|(m[32]&~m[362]&m[506])|(m[32]&m[362]&m[506]))):InitCond[58];
    m[131] = run?((((~m[32]&~m[374]&~m[518])|(m[32]&m[374]&~m[518]))&BiasedRNG[59])|(((m[32]&~m[374]&~m[518])|(~m[32]&m[374]&m[518]))&~BiasedRNG[59])|((~m[32]&~m[374]&m[518])|(m[32]&~m[374]&m[518])|(m[32]&m[374]&m[518]))):InitCond[59];
    m[132] = run?((((~m[33]&~m[243]&~m[387])|(m[33]&m[243]&~m[387]))&BiasedRNG[60])|(((m[33]&~m[243]&~m[387])|(~m[33]&m[243]&m[387]))&~BiasedRNG[60])|((~m[33]&~m[243]&m[387])|(m[33]&~m[243]&m[387])|(m[33]&m[243]&m[387]))):InitCond[60];
    m[133] = run?((((~m[33]&~m[255]&~m[399])|(m[33]&m[255]&~m[399]))&BiasedRNG[61])|(((m[33]&~m[255]&~m[399])|(~m[33]&m[255]&m[399]))&~BiasedRNG[61])|((~m[33]&~m[255]&m[399])|(m[33]&~m[255]&m[399])|(m[33]&m[255]&m[399]))):InitCond[61];
    m[134] = run?((((~m[33]&~m[267]&~m[411])|(m[33]&m[267]&~m[411]))&BiasedRNG[62])|(((m[33]&~m[267]&~m[411])|(~m[33]&m[267]&m[411]))&~BiasedRNG[62])|((~m[33]&~m[267]&m[411])|(m[33]&~m[267]&m[411])|(m[33]&m[267]&m[411]))):InitCond[62];
    m[135] = run?((((~m[33]&~m[279]&~m[423])|(m[33]&m[279]&~m[423]))&BiasedRNG[63])|(((m[33]&~m[279]&~m[423])|(~m[33]&m[279]&m[423]))&~BiasedRNG[63])|((~m[33]&~m[279]&m[423])|(m[33]&~m[279]&m[423])|(m[33]&m[279]&m[423]))):InitCond[63];
    m[136] = run?((((~m[34]&~m[291]&~m[435])|(m[34]&m[291]&~m[435]))&BiasedRNG[64])|(((m[34]&~m[291]&~m[435])|(~m[34]&m[291]&m[435]))&~BiasedRNG[64])|((~m[34]&~m[291]&m[435])|(m[34]&~m[291]&m[435])|(m[34]&m[291]&m[435]))):InitCond[64];
    m[137] = run?((((~m[34]&~m[303]&~m[447])|(m[34]&m[303]&~m[447]))&BiasedRNG[65])|(((m[34]&~m[303]&~m[447])|(~m[34]&m[303]&m[447]))&~BiasedRNG[65])|((~m[34]&~m[303]&m[447])|(m[34]&~m[303]&m[447])|(m[34]&m[303]&m[447]))):InitCond[65];
    m[138] = run?((((~m[34]&~m[315]&~m[459])|(m[34]&m[315]&~m[459]))&BiasedRNG[66])|(((m[34]&~m[315]&~m[459])|(~m[34]&m[315]&m[459]))&~BiasedRNG[66])|((~m[34]&~m[315]&m[459])|(m[34]&~m[315]&m[459])|(m[34]&m[315]&m[459]))):InitCond[66];
    m[139] = run?((((~m[34]&~m[327]&~m[471])|(m[34]&m[327]&~m[471]))&BiasedRNG[67])|(((m[34]&~m[327]&~m[471])|(~m[34]&m[327]&m[471]))&~BiasedRNG[67])|((~m[34]&~m[327]&m[471])|(m[34]&~m[327]&m[471])|(m[34]&m[327]&m[471]))):InitCond[67];
    m[140] = run?((((~m[35]&~m[339]&~m[483])|(m[35]&m[339]&~m[483]))&BiasedRNG[68])|(((m[35]&~m[339]&~m[483])|(~m[35]&m[339]&m[483]))&~BiasedRNG[68])|((~m[35]&~m[339]&m[483])|(m[35]&~m[339]&m[483])|(m[35]&m[339]&m[483]))):InitCond[68];
    m[141] = run?((((~m[35]&~m[351]&~m[495])|(m[35]&m[351]&~m[495]))&BiasedRNG[69])|(((m[35]&~m[351]&~m[495])|(~m[35]&m[351]&m[495]))&~BiasedRNG[69])|((~m[35]&~m[351]&m[495])|(m[35]&~m[351]&m[495])|(m[35]&m[351]&m[495]))):InitCond[69];
    m[142] = run?((((~m[35]&~m[363]&~m[507])|(m[35]&m[363]&~m[507]))&BiasedRNG[70])|(((m[35]&~m[363]&~m[507])|(~m[35]&m[363]&m[507]))&~BiasedRNG[70])|((~m[35]&~m[363]&m[507])|(m[35]&~m[363]&m[507])|(m[35]&m[363]&m[507]))):InitCond[70];
    m[143] = run?((((~m[35]&~m[375]&~m[519])|(m[35]&m[375]&~m[519]))&BiasedRNG[71])|(((m[35]&~m[375]&~m[519])|(~m[35]&m[375]&m[519]))&~BiasedRNG[71])|((~m[35]&~m[375]&m[519])|(m[35]&~m[375]&m[519])|(m[35]&m[375]&m[519]))):InitCond[71];
    m[144] = run?((((~m[36]&~m[244]&~m[388])|(m[36]&m[244]&~m[388]))&BiasedRNG[72])|(((m[36]&~m[244]&~m[388])|(~m[36]&m[244]&m[388]))&~BiasedRNG[72])|((~m[36]&~m[244]&m[388])|(m[36]&~m[244]&m[388])|(m[36]&m[244]&m[388]))):InitCond[72];
    m[145] = run?((((~m[36]&~m[256]&~m[400])|(m[36]&m[256]&~m[400]))&BiasedRNG[73])|(((m[36]&~m[256]&~m[400])|(~m[36]&m[256]&m[400]))&~BiasedRNG[73])|((~m[36]&~m[256]&m[400])|(m[36]&~m[256]&m[400])|(m[36]&m[256]&m[400]))):InitCond[73];
    m[146] = run?((((~m[36]&~m[268]&~m[412])|(m[36]&m[268]&~m[412]))&BiasedRNG[74])|(((m[36]&~m[268]&~m[412])|(~m[36]&m[268]&m[412]))&~BiasedRNG[74])|((~m[36]&~m[268]&m[412])|(m[36]&~m[268]&m[412])|(m[36]&m[268]&m[412]))):InitCond[74];
    m[147] = run?((((~m[36]&~m[280]&~m[424])|(m[36]&m[280]&~m[424]))&BiasedRNG[75])|(((m[36]&~m[280]&~m[424])|(~m[36]&m[280]&m[424]))&~BiasedRNG[75])|((~m[36]&~m[280]&m[424])|(m[36]&~m[280]&m[424])|(m[36]&m[280]&m[424]))):InitCond[75];
    m[148] = run?((((~m[37]&~m[292]&~m[436])|(m[37]&m[292]&~m[436]))&BiasedRNG[76])|(((m[37]&~m[292]&~m[436])|(~m[37]&m[292]&m[436]))&~BiasedRNG[76])|((~m[37]&~m[292]&m[436])|(m[37]&~m[292]&m[436])|(m[37]&m[292]&m[436]))):InitCond[76];
    m[149] = run?((((~m[37]&~m[304]&~m[448])|(m[37]&m[304]&~m[448]))&BiasedRNG[77])|(((m[37]&~m[304]&~m[448])|(~m[37]&m[304]&m[448]))&~BiasedRNG[77])|((~m[37]&~m[304]&m[448])|(m[37]&~m[304]&m[448])|(m[37]&m[304]&m[448]))):InitCond[77];
    m[150] = run?((((~m[37]&~m[316]&~m[460])|(m[37]&m[316]&~m[460]))&BiasedRNG[78])|(((m[37]&~m[316]&~m[460])|(~m[37]&m[316]&m[460]))&~BiasedRNG[78])|((~m[37]&~m[316]&m[460])|(m[37]&~m[316]&m[460])|(m[37]&m[316]&m[460]))):InitCond[78];
    m[151] = run?((((~m[37]&~m[328]&~m[472])|(m[37]&m[328]&~m[472]))&BiasedRNG[79])|(((m[37]&~m[328]&~m[472])|(~m[37]&m[328]&m[472]))&~BiasedRNG[79])|((~m[37]&~m[328]&m[472])|(m[37]&~m[328]&m[472])|(m[37]&m[328]&m[472]))):InitCond[79];
    m[152] = run?((((~m[38]&~m[340]&~m[484])|(m[38]&m[340]&~m[484]))&BiasedRNG[80])|(((m[38]&~m[340]&~m[484])|(~m[38]&m[340]&m[484]))&~BiasedRNG[80])|((~m[38]&~m[340]&m[484])|(m[38]&~m[340]&m[484])|(m[38]&m[340]&m[484]))):InitCond[80];
    m[153] = run?((((~m[38]&~m[352]&~m[496])|(m[38]&m[352]&~m[496]))&BiasedRNG[81])|(((m[38]&~m[352]&~m[496])|(~m[38]&m[352]&m[496]))&~BiasedRNG[81])|((~m[38]&~m[352]&m[496])|(m[38]&~m[352]&m[496])|(m[38]&m[352]&m[496]))):InitCond[81];
    m[154] = run?((((~m[38]&~m[364]&~m[508])|(m[38]&m[364]&~m[508]))&BiasedRNG[82])|(((m[38]&~m[364]&~m[508])|(~m[38]&m[364]&m[508]))&~BiasedRNG[82])|((~m[38]&~m[364]&m[508])|(m[38]&~m[364]&m[508])|(m[38]&m[364]&m[508]))):InitCond[82];
    m[155] = run?((((~m[38]&~m[376]&~m[520])|(m[38]&m[376]&~m[520]))&BiasedRNG[83])|(((m[38]&~m[376]&~m[520])|(~m[38]&m[376]&m[520]))&~BiasedRNG[83])|((~m[38]&~m[376]&m[520])|(m[38]&~m[376]&m[520])|(m[38]&m[376]&m[520]))):InitCond[83];
    m[156] = run?((((~m[39]&~m[245]&~m[389])|(m[39]&m[245]&~m[389]))&BiasedRNG[84])|(((m[39]&~m[245]&~m[389])|(~m[39]&m[245]&m[389]))&~BiasedRNG[84])|((~m[39]&~m[245]&m[389])|(m[39]&~m[245]&m[389])|(m[39]&m[245]&m[389]))):InitCond[84];
    m[157] = run?((((~m[39]&~m[257]&~m[401])|(m[39]&m[257]&~m[401]))&BiasedRNG[85])|(((m[39]&~m[257]&~m[401])|(~m[39]&m[257]&m[401]))&~BiasedRNG[85])|((~m[39]&~m[257]&m[401])|(m[39]&~m[257]&m[401])|(m[39]&m[257]&m[401]))):InitCond[85];
    m[158] = run?((((~m[39]&~m[269]&~m[413])|(m[39]&m[269]&~m[413]))&BiasedRNG[86])|(((m[39]&~m[269]&~m[413])|(~m[39]&m[269]&m[413]))&~BiasedRNG[86])|((~m[39]&~m[269]&m[413])|(m[39]&~m[269]&m[413])|(m[39]&m[269]&m[413]))):InitCond[86];
    m[159] = run?((((~m[39]&~m[281]&~m[425])|(m[39]&m[281]&~m[425]))&BiasedRNG[87])|(((m[39]&~m[281]&~m[425])|(~m[39]&m[281]&m[425]))&~BiasedRNG[87])|((~m[39]&~m[281]&m[425])|(m[39]&~m[281]&m[425])|(m[39]&m[281]&m[425]))):InitCond[87];
    m[160] = run?((((~m[40]&~m[293]&~m[437])|(m[40]&m[293]&~m[437]))&BiasedRNG[88])|(((m[40]&~m[293]&~m[437])|(~m[40]&m[293]&m[437]))&~BiasedRNG[88])|((~m[40]&~m[293]&m[437])|(m[40]&~m[293]&m[437])|(m[40]&m[293]&m[437]))):InitCond[88];
    m[161] = run?((((~m[40]&~m[305]&~m[449])|(m[40]&m[305]&~m[449]))&BiasedRNG[89])|(((m[40]&~m[305]&~m[449])|(~m[40]&m[305]&m[449]))&~BiasedRNG[89])|((~m[40]&~m[305]&m[449])|(m[40]&~m[305]&m[449])|(m[40]&m[305]&m[449]))):InitCond[89];
    m[162] = run?((((~m[40]&~m[317]&~m[461])|(m[40]&m[317]&~m[461]))&BiasedRNG[90])|(((m[40]&~m[317]&~m[461])|(~m[40]&m[317]&m[461]))&~BiasedRNG[90])|((~m[40]&~m[317]&m[461])|(m[40]&~m[317]&m[461])|(m[40]&m[317]&m[461]))):InitCond[90];
    m[163] = run?((((~m[40]&~m[329]&~m[473])|(m[40]&m[329]&~m[473]))&BiasedRNG[91])|(((m[40]&~m[329]&~m[473])|(~m[40]&m[329]&m[473]))&~BiasedRNG[91])|((~m[40]&~m[329]&m[473])|(m[40]&~m[329]&m[473])|(m[40]&m[329]&m[473]))):InitCond[91];
    m[164] = run?((((~m[41]&~m[341]&~m[485])|(m[41]&m[341]&~m[485]))&BiasedRNG[92])|(((m[41]&~m[341]&~m[485])|(~m[41]&m[341]&m[485]))&~BiasedRNG[92])|((~m[41]&~m[341]&m[485])|(m[41]&~m[341]&m[485])|(m[41]&m[341]&m[485]))):InitCond[92];
    m[165] = run?((((~m[41]&~m[353]&~m[497])|(m[41]&m[353]&~m[497]))&BiasedRNG[93])|(((m[41]&~m[353]&~m[497])|(~m[41]&m[353]&m[497]))&~BiasedRNG[93])|((~m[41]&~m[353]&m[497])|(m[41]&~m[353]&m[497])|(m[41]&m[353]&m[497]))):InitCond[93];
    m[166] = run?((((~m[41]&~m[365]&~m[509])|(m[41]&m[365]&~m[509]))&BiasedRNG[94])|(((m[41]&~m[365]&~m[509])|(~m[41]&m[365]&m[509]))&~BiasedRNG[94])|((~m[41]&~m[365]&m[509])|(m[41]&~m[365]&m[509])|(m[41]&m[365]&m[509]))):InitCond[94];
    m[167] = run?((((~m[41]&~m[377]&~m[521])|(m[41]&m[377]&~m[521]))&BiasedRNG[95])|(((m[41]&~m[377]&~m[521])|(~m[41]&m[377]&m[521]))&~BiasedRNG[95])|((~m[41]&~m[377]&m[521])|(m[41]&~m[377]&m[521])|(m[41]&m[377]&m[521]))):InitCond[95];
    m[168] = run?((((~m[42]&~m[246]&~m[390])|(m[42]&m[246]&~m[390]))&BiasedRNG[96])|(((m[42]&~m[246]&~m[390])|(~m[42]&m[246]&m[390]))&~BiasedRNG[96])|((~m[42]&~m[246]&m[390])|(m[42]&~m[246]&m[390])|(m[42]&m[246]&m[390]))):InitCond[96];
    m[169] = run?((((~m[42]&~m[258]&~m[402])|(m[42]&m[258]&~m[402]))&BiasedRNG[97])|(((m[42]&~m[258]&~m[402])|(~m[42]&m[258]&m[402]))&~BiasedRNG[97])|((~m[42]&~m[258]&m[402])|(m[42]&~m[258]&m[402])|(m[42]&m[258]&m[402]))):InitCond[97];
    m[170] = run?((((~m[42]&~m[270]&~m[414])|(m[42]&m[270]&~m[414]))&BiasedRNG[98])|(((m[42]&~m[270]&~m[414])|(~m[42]&m[270]&m[414]))&~BiasedRNG[98])|((~m[42]&~m[270]&m[414])|(m[42]&~m[270]&m[414])|(m[42]&m[270]&m[414]))):InitCond[98];
    m[171] = run?((((~m[42]&~m[282]&~m[426])|(m[42]&m[282]&~m[426]))&BiasedRNG[99])|(((m[42]&~m[282]&~m[426])|(~m[42]&m[282]&m[426]))&~BiasedRNG[99])|((~m[42]&~m[282]&m[426])|(m[42]&~m[282]&m[426])|(m[42]&m[282]&m[426]))):InitCond[99];
    m[172] = run?((((~m[43]&~m[294]&~m[438])|(m[43]&m[294]&~m[438]))&BiasedRNG[100])|(((m[43]&~m[294]&~m[438])|(~m[43]&m[294]&m[438]))&~BiasedRNG[100])|((~m[43]&~m[294]&m[438])|(m[43]&~m[294]&m[438])|(m[43]&m[294]&m[438]))):InitCond[100];
    m[173] = run?((((~m[43]&~m[306]&~m[450])|(m[43]&m[306]&~m[450]))&BiasedRNG[101])|(((m[43]&~m[306]&~m[450])|(~m[43]&m[306]&m[450]))&~BiasedRNG[101])|((~m[43]&~m[306]&m[450])|(m[43]&~m[306]&m[450])|(m[43]&m[306]&m[450]))):InitCond[101];
    m[174] = run?((((~m[43]&~m[318]&~m[462])|(m[43]&m[318]&~m[462]))&BiasedRNG[102])|(((m[43]&~m[318]&~m[462])|(~m[43]&m[318]&m[462]))&~BiasedRNG[102])|((~m[43]&~m[318]&m[462])|(m[43]&~m[318]&m[462])|(m[43]&m[318]&m[462]))):InitCond[102];
    m[175] = run?((((~m[43]&~m[330]&~m[474])|(m[43]&m[330]&~m[474]))&BiasedRNG[103])|(((m[43]&~m[330]&~m[474])|(~m[43]&m[330]&m[474]))&~BiasedRNG[103])|((~m[43]&~m[330]&m[474])|(m[43]&~m[330]&m[474])|(m[43]&m[330]&m[474]))):InitCond[103];
    m[176] = run?((((~m[44]&~m[342]&~m[486])|(m[44]&m[342]&~m[486]))&BiasedRNG[104])|(((m[44]&~m[342]&~m[486])|(~m[44]&m[342]&m[486]))&~BiasedRNG[104])|((~m[44]&~m[342]&m[486])|(m[44]&~m[342]&m[486])|(m[44]&m[342]&m[486]))):InitCond[104];
    m[177] = run?((((~m[44]&~m[354]&~m[498])|(m[44]&m[354]&~m[498]))&BiasedRNG[105])|(((m[44]&~m[354]&~m[498])|(~m[44]&m[354]&m[498]))&~BiasedRNG[105])|((~m[44]&~m[354]&m[498])|(m[44]&~m[354]&m[498])|(m[44]&m[354]&m[498]))):InitCond[105];
    m[178] = run?((((~m[44]&~m[366]&~m[510])|(m[44]&m[366]&~m[510]))&BiasedRNG[106])|(((m[44]&~m[366]&~m[510])|(~m[44]&m[366]&m[510]))&~BiasedRNG[106])|((~m[44]&~m[366]&m[510])|(m[44]&~m[366]&m[510])|(m[44]&m[366]&m[510]))):InitCond[106];
    m[179] = run?((((~m[44]&~m[378]&~m[522])|(m[44]&m[378]&~m[522]))&BiasedRNG[107])|(((m[44]&~m[378]&~m[522])|(~m[44]&m[378]&m[522]))&~BiasedRNG[107])|((~m[44]&~m[378]&m[522])|(m[44]&~m[378]&m[522])|(m[44]&m[378]&m[522]))):InitCond[107];
    m[180] = run?((((~m[45]&~m[247]&~m[391])|(m[45]&m[247]&~m[391]))&BiasedRNG[108])|(((m[45]&~m[247]&~m[391])|(~m[45]&m[247]&m[391]))&~BiasedRNG[108])|((~m[45]&~m[247]&m[391])|(m[45]&~m[247]&m[391])|(m[45]&m[247]&m[391]))):InitCond[108];
    m[181] = run?((((~m[45]&~m[259]&~m[403])|(m[45]&m[259]&~m[403]))&BiasedRNG[109])|(((m[45]&~m[259]&~m[403])|(~m[45]&m[259]&m[403]))&~BiasedRNG[109])|((~m[45]&~m[259]&m[403])|(m[45]&~m[259]&m[403])|(m[45]&m[259]&m[403]))):InitCond[109];
    m[182] = run?((((~m[45]&~m[271]&~m[415])|(m[45]&m[271]&~m[415]))&BiasedRNG[110])|(((m[45]&~m[271]&~m[415])|(~m[45]&m[271]&m[415]))&~BiasedRNG[110])|((~m[45]&~m[271]&m[415])|(m[45]&~m[271]&m[415])|(m[45]&m[271]&m[415]))):InitCond[110];
    m[183] = run?((((~m[45]&~m[283]&~m[427])|(m[45]&m[283]&~m[427]))&BiasedRNG[111])|(((m[45]&~m[283]&~m[427])|(~m[45]&m[283]&m[427]))&~BiasedRNG[111])|((~m[45]&~m[283]&m[427])|(m[45]&~m[283]&m[427])|(m[45]&m[283]&m[427]))):InitCond[111];
    m[184] = run?((((~m[46]&~m[295]&~m[439])|(m[46]&m[295]&~m[439]))&BiasedRNG[112])|(((m[46]&~m[295]&~m[439])|(~m[46]&m[295]&m[439]))&~BiasedRNG[112])|((~m[46]&~m[295]&m[439])|(m[46]&~m[295]&m[439])|(m[46]&m[295]&m[439]))):InitCond[112];
    m[185] = run?((((~m[46]&~m[307]&~m[451])|(m[46]&m[307]&~m[451]))&BiasedRNG[113])|(((m[46]&~m[307]&~m[451])|(~m[46]&m[307]&m[451]))&~BiasedRNG[113])|((~m[46]&~m[307]&m[451])|(m[46]&~m[307]&m[451])|(m[46]&m[307]&m[451]))):InitCond[113];
    m[186] = run?((((~m[46]&~m[319]&~m[463])|(m[46]&m[319]&~m[463]))&BiasedRNG[114])|(((m[46]&~m[319]&~m[463])|(~m[46]&m[319]&m[463]))&~BiasedRNG[114])|((~m[46]&~m[319]&m[463])|(m[46]&~m[319]&m[463])|(m[46]&m[319]&m[463]))):InitCond[114];
    m[187] = run?((((~m[46]&~m[331]&~m[475])|(m[46]&m[331]&~m[475]))&BiasedRNG[115])|(((m[46]&~m[331]&~m[475])|(~m[46]&m[331]&m[475]))&~BiasedRNG[115])|((~m[46]&~m[331]&m[475])|(m[46]&~m[331]&m[475])|(m[46]&m[331]&m[475]))):InitCond[115];
    m[188] = run?((((~m[47]&~m[343]&~m[487])|(m[47]&m[343]&~m[487]))&BiasedRNG[116])|(((m[47]&~m[343]&~m[487])|(~m[47]&m[343]&m[487]))&~BiasedRNG[116])|((~m[47]&~m[343]&m[487])|(m[47]&~m[343]&m[487])|(m[47]&m[343]&m[487]))):InitCond[116];
    m[189] = run?((((~m[47]&~m[355]&~m[499])|(m[47]&m[355]&~m[499]))&BiasedRNG[117])|(((m[47]&~m[355]&~m[499])|(~m[47]&m[355]&m[499]))&~BiasedRNG[117])|((~m[47]&~m[355]&m[499])|(m[47]&~m[355]&m[499])|(m[47]&m[355]&m[499]))):InitCond[117];
    m[190] = run?((((~m[47]&~m[367]&~m[511])|(m[47]&m[367]&~m[511]))&BiasedRNG[118])|(((m[47]&~m[367]&~m[511])|(~m[47]&m[367]&m[511]))&~BiasedRNG[118])|((~m[47]&~m[367]&m[511])|(m[47]&~m[367]&m[511])|(m[47]&m[367]&m[511]))):InitCond[118];
    m[191] = run?((((~m[47]&~m[379]&~m[523])|(m[47]&m[379]&~m[523]))&BiasedRNG[119])|(((m[47]&~m[379]&~m[523])|(~m[47]&m[379]&m[523]))&~BiasedRNG[119])|((~m[47]&~m[379]&m[523])|(m[47]&~m[379]&m[523])|(m[47]&m[379]&m[523]))):InitCond[119];
    m[192] = run?((((~m[48]&~m[248]&~m[392])|(m[48]&m[248]&~m[392]))&BiasedRNG[120])|(((m[48]&~m[248]&~m[392])|(~m[48]&m[248]&m[392]))&~BiasedRNG[120])|((~m[48]&~m[248]&m[392])|(m[48]&~m[248]&m[392])|(m[48]&m[248]&m[392]))):InitCond[120];
    m[193] = run?((((~m[48]&~m[260]&~m[404])|(m[48]&m[260]&~m[404]))&BiasedRNG[121])|(((m[48]&~m[260]&~m[404])|(~m[48]&m[260]&m[404]))&~BiasedRNG[121])|((~m[48]&~m[260]&m[404])|(m[48]&~m[260]&m[404])|(m[48]&m[260]&m[404]))):InitCond[121];
    m[194] = run?((((~m[48]&~m[272]&~m[416])|(m[48]&m[272]&~m[416]))&BiasedRNG[122])|(((m[48]&~m[272]&~m[416])|(~m[48]&m[272]&m[416]))&~BiasedRNG[122])|((~m[48]&~m[272]&m[416])|(m[48]&~m[272]&m[416])|(m[48]&m[272]&m[416]))):InitCond[122];
    m[195] = run?((((~m[48]&~m[284]&~m[428])|(m[48]&m[284]&~m[428]))&BiasedRNG[123])|(((m[48]&~m[284]&~m[428])|(~m[48]&m[284]&m[428]))&~BiasedRNG[123])|((~m[48]&~m[284]&m[428])|(m[48]&~m[284]&m[428])|(m[48]&m[284]&m[428]))):InitCond[123];
    m[196] = run?((((~m[49]&~m[296]&~m[440])|(m[49]&m[296]&~m[440]))&BiasedRNG[124])|(((m[49]&~m[296]&~m[440])|(~m[49]&m[296]&m[440]))&~BiasedRNG[124])|((~m[49]&~m[296]&m[440])|(m[49]&~m[296]&m[440])|(m[49]&m[296]&m[440]))):InitCond[124];
    m[197] = run?((((~m[49]&~m[308]&~m[452])|(m[49]&m[308]&~m[452]))&BiasedRNG[125])|(((m[49]&~m[308]&~m[452])|(~m[49]&m[308]&m[452]))&~BiasedRNG[125])|((~m[49]&~m[308]&m[452])|(m[49]&~m[308]&m[452])|(m[49]&m[308]&m[452]))):InitCond[125];
    m[198] = run?((((~m[49]&~m[320]&~m[464])|(m[49]&m[320]&~m[464]))&BiasedRNG[126])|(((m[49]&~m[320]&~m[464])|(~m[49]&m[320]&m[464]))&~BiasedRNG[126])|((~m[49]&~m[320]&m[464])|(m[49]&~m[320]&m[464])|(m[49]&m[320]&m[464]))):InitCond[126];
    m[199] = run?((((~m[49]&~m[332]&~m[476])|(m[49]&m[332]&~m[476]))&BiasedRNG[127])|(((m[49]&~m[332]&~m[476])|(~m[49]&m[332]&m[476]))&~BiasedRNG[127])|((~m[49]&~m[332]&m[476])|(m[49]&~m[332]&m[476])|(m[49]&m[332]&m[476]))):InitCond[127];
    m[200] = run?((((~m[50]&~m[344]&~m[488])|(m[50]&m[344]&~m[488]))&BiasedRNG[128])|(((m[50]&~m[344]&~m[488])|(~m[50]&m[344]&m[488]))&~BiasedRNG[128])|((~m[50]&~m[344]&m[488])|(m[50]&~m[344]&m[488])|(m[50]&m[344]&m[488]))):InitCond[128];
    m[201] = run?((((~m[50]&~m[356]&~m[500])|(m[50]&m[356]&~m[500]))&BiasedRNG[129])|(((m[50]&~m[356]&~m[500])|(~m[50]&m[356]&m[500]))&~BiasedRNG[129])|((~m[50]&~m[356]&m[500])|(m[50]&~m[356]&m[500])|(m[50]&m[356]&m[500]))):InitCond[129];
    m[202] = run?((((~m[50]&~m[368]&~m[512])|(m[50]&m[368]&~m[512]))&BiasedRNG[130])|(((m[50]&~m[368]&~m[512])|(~m[50]&m[368]&m[512]))&~BiasedRNG[130])|((~m[50]&~m[368]&m[512])|(m[50]&~m[368]&m[512])|(m[50]&m[368]&m[512]))):InitCond[130];
    m[203] = run?((((~m[50]&~m[380]&~m[524])|(m[50]&m[380]&~m[524]))&BiasedRNG[131])|(((m[50]&~m[380]&~m[524])|(~m[50]&m[380]&m[524]))&~BiasedRNG[131])|((~m[50]&~m[380]&m[524])|(m[50]&~m[380]&m[524])|(m[50]&m[380]&m[524]))):InitCond[131];
    m[204] = run?((((~m[51]&~m[249]&~m[393])|(m[51]&m[249]&~m[393]))&BiasedRNG[132])|(((m[51]&~m[249]&~m[393])|(~m[51]&m[249]&m[393]))&~BiasedRNG[132])|((~m[51]&~m[249]&m[393])|(m[51]&~m[249]&m[393])|(m[51]&m[249]&m[393]))):InitCond[132];
    m[205] = run?((((~m[51]&~m[261]&~m[405])|(m[51]&m[261]&~m[405]))&BiasedRNG[133])|(((m[51]&~m[261]&~m[405])|(~m[51]&m[261]&m[405]))&~BiasedRNG[133])|((~m[51]&~m[261]&m[405])|(m[51]&~m[261]&m[405])|(m[51]&m[261]&m[405]))):InitCond[133];
    m[206] = run?((((~m[51]&~m[273]&~m[417])|(m[51]&m[273]&~m[417]))&BiasedRNG[134])|(((m[51]&~m[273]&~m[417])|(~m[51]&m[273]&m[417]))&~BiasedRNG[134])|((~m[51]&~m[273]&m[417])|(m[51]&~m[273]&m[417])|(m[51]&m[273]&m[417]))):InitCond[134];
    m[207] = run?((((~m[51]&~m[285]&~m[429])|(m[51]&m[285]&~m[429]))&BiasedRNG[135])|(((m[51]&~m[285]&~m[429])|(~m[51]&m[285]&m[429]))&~BiasedRNG[135])|((~m[51]&~m[285]&m[429])|(m[51]&~m[285]&m[429])|(m[51]&m[285]&m[429]))):InitCond[135];
    m[208] = run?((((~m[52]&~m[297]&~m[441])|(m[52]&m[297]&~m[441]))&BiasedRNG[136])|(((m[52]&~m[297]&~m[441])|(~m[52]&m[297]&m[441]))&~BiasedRNG[136])|((~m[52]&~m[297]&m[441])|(m[52]&~m[297]&m[441])|(m[52]&m[297]&m[441]))):InitCond[136];
    m[209] = run?((((~m[52]&~m[309]&~m[453])|(m[52]&m[309]&~m[453]))&BiasedRNG[137])|(((m[52]&~m[309]&~m[453])|(~m[52]&m[309]&m[453]))&~BiasedRNG[137])|((~m[52]&~m[309]&m[453])|(m[52]&~m[309]&m[453])|(m[52]&m[309]&m[453]))):InitCond[137];
    m[210] = run?((((~m[52]&~m[321]&~m[465])|(m[52]&m[321]&~m[465]))&BiasedRNG[138])|(((m[52]&~m[321]&~m[465])|(~m[52]&m[321]&m[465]))&~BiasedRNG[138])|((~m[52]&~m[321]&m[465])|(m[52]&~m[321]&m[465])|(m[52]&m[321]&m[465]))):InitCond[138];
    m[211] = run?((((~m[52]&~m[333]&~m[477])|(m[52]&m[333]&~m[477]))&BiasedRNG[139])|(((m[52]&~m[333]&~m[477])|(~m[52]&m[333]&m[477]))&~BiasedRNG[139])|((~m[52]&~m[333]&m[477])|(m[52]&~m[333]&m[477])|(m[52]&m[333]&m[477]))):InitCond[139];
    m[212] = run?((((~m[53]&~m[345]&~m[489])|(m[53]&m[345]&~m[489]))&BiasedRNG[140])|(((m[53]&~m[345]&~m[489])|(~m[53]&m[345]&m[489]))&~BiasedRNG[140])|((~m[53]&~m[345]&m[489])|(m[53]&~m[345]&m[489])|(m[53]&m[345]&m[489]))):InitCond[140];
    m[213] = run?((((~m[53]&~m[357]&~m[501])|(m[53]&m[357]&~m[501]))&BiasedRNG[141])|(((m[53]&~m[357]&~m[501])|(~m[53]&m[357]&m[501]))&~BiasedRNG[141])|((~m[53]&~m[357]&m[501])|(m[53]&~m[357]&m[501])|(m[53]&m[357]&m[501]))):InitCond[141];
    m[214] = run?((((~m[53]&~m[369]&~m[513])|(m[53]&m[369]&~m[513]))&BiasedRNG[142])|(((m[53]&~m[369]&~m[513])|(~m[53]&m[369]&m[513]))&~BiasedRNG[142])|((~m[53]&~m[369]&m[513])|(m[53]&~m[369]&m[513])|(m[53]&m[369]&m[513]))):InitCond[142];
    m[215] = run?((((~m[53]&~m[381]&~m[525])|(m[53]&m[381]&~m[525]))&BiasedRNG[143])|(((m[53]&~m[381]&~m[525])|(~m[53]&m[381]&m[525]))&~BiasedRNG[143])|((~m[53]&~m[381]&m[525])|(m[53]&~m[381]&m[525])|(m[53]&m[381]&m[525]))):InitCond[143];
    m[216] = run?((((~m[54]&~m[250]&~m[394])|(m[54]&m[250]&~m[394]))&BiasedRNG[144])|(((m[54]&~m[250]&~m[394])|(~m[54]&m[250]&m[394]))&~BiasedRNG[144])|((~m[54]&~m[250]&m[394])|(m[54]&~m[250]&m[394])|(m[54]&m[250]&m[394]))):InitCond[144];
    m[217] = run?((((~m[54]&~m[262]&~m[406])|(m[54]&m[262]&~m[406]))&BiasedRNG[145])|(((m[54]&~m[262]&~m[406])|(~m[54]&m[262]&m[406]))&~BiasedRNG[145])|((~m[54]&~m[262]&m[406])|(m[54]&~m[262]&m[406])|(m[54]&m[262]&m[406]))):InitCond[145];
    m[218] = run?((((~m[54]&~m[274]&~m[418])|(m[54]&m[274]&~m[418]))&BiasedRNG[146])|(((m[54]&~m[274]&~m[418])|(~m[54]&m[274]&m[418]))&~BiasedRNG[146])|((~m[54]&~m[274]&m[418])|(m[54]&~m[274]&m[418])|(m[54]&m[274]&m[418]))):InitCond[146];
    m[219] = run?((((~m[54]&~m[286]&~m[430])|(m[54]&m[286]&~m[430]))&BiasedRNG[147])|(((m[54]&~m[286]&~m[430])|(~m[54]&m[286]&m[430]))&~BiasedRNG[147])|((~m[54]&~m[286]&m[430])|(m[54]&~m[286]&m[430])|(m[54]&m[286]&m[430]))):InitCond[147];
    m[220] = run?((((~m[55]&~m[298]&~m[442])|(m[55]&m[298]&~m[442]))&BiasedRNG[148])|(((m[55]&~m[298]&~m[442])|(~m[55]&m[298]&m[442]))&~BiasedRNG[148])|((~m[55]&~m[298]&m[442])|(m[55]&~m[298]&m[442])|(m[55]&m[298]&m[442]))):InitCond[148];
    m[221] = run?((((~m[55]&~m[310]&~m[454])|(m[55]&m[310]&~m[454]))&BiasedRNG[149])|(((m[55]&~m[310]&~m[454])|(~m[55]&m[310]&m[454]))&~BiasedRNG[149])|((~m[55]&~m[310]&m[454])|(m[55]&~m[310]&m[454])|(m[55]&m[310]&m[454]))):InitCond[149];
    m[222] = run?((((~m[55]&~m[322]&~m[466])|(m[55]&m[322]&~m[466]))&BiasedRNG[150])|(((m[55]&~m[322]&~m[466])|(~m[55]&m[322]&m[466]))&~BiasedRNG[150])|((~m[55]&~m[322]&m[466])|(m[55]&~m[322]&m[466])|(m[55]&m[322]&m[466]))):InitCond[150];
    m[223] = run?((((~m[55]&~m[334]&~m[478])|(m[55]&m[334]&~m[478]))&BiasedRNG[151])|(((m[55]&~m[334]&~m[478])|(~m[55]&m[334]&m[478]))&~BiasedRNG[151])|((~m[55]&~m[334]&m[478])|(m[55]&~m[334]&m[478])|(m[55]&m[334]&m[478]))):InitCond[151];
    m[224] = run?((((~m[56]&~m[346]&~m[490])|(m[56]&m[346]&~m[490]))&BiasedRNG[152])|(((m[56]&~m[346]&~m[490])|(~m[56]&m[346]&m[490]))&~BiasedRNG[152])|((~m[56]&~m[346]&m[490])|(m[56]&~m[346]&m[490])|(m[56]&m[346]&m[490]))):InitCond[152];
    m[225] = run?((((~m[56]&~m[358]&~m[502])|(m[56]&m[358]&~m[502]))&BiasedRNG[153])|(((m[56]&~m[358]&~m[502])|(~m[56]&m[358]&m[502]))&~BiasedRNG[153])|((~m[56]&~m[358]&m[502])|(m[56]&~m[358]&m[502])|(m[56]&m[358]&m[502]))):InitCond[153];
    m[226] = run?((((~m[56]&~m[370]&~m[514])|(m[56]&m[370]&~m[514]))&BiasedRNG[154])|(((m[56]&~m[370]&~m[514])|(~m[56]&m[370]&m[514]))&~BiasedRNG[154])|((~m[56]&~m[370]&m[514])|(m[56]&~m[370]&m[514])|(m[56]&m[370]&m[514]))):InitCond[154];
    m[227] = run?((((~m[56]&~m[382]&~m[526])|(m[56]&m[382]&~m[526]))&BiasedRNG[155])|(((m[56]&~m[382]&~m[526])|(~m[56]&m[382]&m[526]))&~BiasedRNG[155])|((~m[56]&~m[382]&m[526])|(m[56]&~m[382]&m[526])|(m[56]&m[382]&m[526]))):InitCond[155];
    m[228] = run?((((~m[57]&~m[251]&~m[395])|(m[57]&m[251]&~m[395]))&BiasedRNG[156])|(((m[57]&~m[251]&~m[395])|(~m[57]&m[251]&m[395]))&~BiasedRNG[156])|((~m[57]&~m[251]&m[395])|(m[57]&~m[251]&m[395])|(m[57]&m[251]&m[395]))):InitCond[156];
    m[229] = run?((((~m[57]&~m[263]&~m[407])|(m[57]&m[263]&~m[407]))&BiasedRNG[157])|(((m[57]&~m[263]&~m[407])|(~m[57]&m[263]&m[407]))&~BiasedRNG[157])|((~m[57]&~m[263]&m[407])|(m[57]&~m[263]&m[407])|(m[57]&m[263]&m[407]))):InitCond[157];
    m[230] = run?((((~m[57]&~m[275]&~m[419])|(m[57]&m[275]&~m[419]))&BiasedRNG[158])|(((m[57]&~m[275]&~m[419])|(~m[57]&m[275]&m[419]))&~BiasedRNG[158])|((~m[57]&~m[275]&m[419])|(m[57]&~m[275]&m[419])|(m[57]&m[275]&m[419]))):InitCond[158];
    m[231] = run?((((~m[57]&~m[287]&~m[431])|(m[57]&m[287]&~m[431]))&BiasedRNG[159])|(((m[57]&~m[287]&~m[431])|(~m[57]&m[287]&m[431]))&~BiasedRNG[159])|((~m[57]&~m[287]&m[431])|(m[57]&~m[287]&m[431])|(m[57]&m[287]&m[431]))):InitCond[159];
    m[232] = run?((((~m[58]&~m[299]&~m[443])|(m[58]&m[299]&~m[443]))&BiasedRNG[160])|(((m[58]&~m[299]&~m[443])|(~m[58]&m[299]&m[443]))&~BiasedRNG[160])|((~m[58]&~m[299]&m[443])|(m[58]&~m[299]&m[443])|(m[58]&m[299]&m[443]))):InitCond[160];
    m[233] = run?((((~m[58]&~m[311]&~m[455])|(m[58]&m[311]&~m[455]))&BiasedRNG[161])|(((m[58]&~m[311]&~m[455])|(~m[58]&m[311]&m[455]))&~BiasedRNG[161])|((~m[58]&~m[311]&m[455])|(m[58]&~m[311]&m[455])|(m[58]&m[311]&m[455]))):InitCond[161];
    m[234] = run?((((~m[58]&~m[323]&~m[467])|(m[58]&m[323]&~m[467]))&BiasedRNG[162])|(((m[58]&~m[323]&~m[467])|(~m[58]&m[323]&m[467]))&~BiasedRNG[162])|((~m[58]&~m[323]&m[467])|(m[58]&~m[323]&m[467])|(m[58]&m[323]&m[467]))):InitCond[162];
    m[235] = run?((((~m[58]&~m[335]&~m[479])|(m[58]&m[335]&~m[479]))&BiasedRNG[163])|(((m[58]&~m[335]&~m[479])|(~m[58]&m[335]&m[479]))&~BiasedRNG[163])|((~m[58]&~m[335]&m[479])|(m[58]&~m[335]&m[479])|(m[58]&m[335]&m[479]))):InitCond[163];
    m[236] = run?((((~m[59]&~m[347]&~m[491])|(m[59]&m[347]&~m[491]))&BiasedRNG[164])|(((m[59]&~m[347]&~m[491])|(~m[59]&m[347]&m[491]))&~BiasedRNG[164])|((~m[59]&~m[347]&m[491])|(m[59]&~m[347]&m[491])|(m[59]&m[347]&m[491]))):InitCond[164];
    m[237] = run?((((~m[59]&~m[359]&~m[503])|(m[59]&m[359]&~m[503]))&BiasedRNG[165])|(((m[59]&~m[359]&~m[503])|(~m[59]&m[359]&m[503]))&~BiasedRNG[165])|((~m[59]&~m[359]&m[503])|(m[59]&~m[359]&m[503])|(m[59]&m[359]&m[503]))):InitCond[165];
    m[238] = run?((((~m[59]&~m[371]&~m[515])|(m[59]&m[371]&~m[515]))&BiasedRNG[166])|(((m[59]&~m[371]&~m[515])|(~m[59]&m[371]&m[515]))&~BiasedRNG[166])|((~m[59]&~m[371]&m[515])|(m[59]&~m[371]&m[515])|(m[59]&m[371]&m[515]))):InitCond[166];
    m[239] = run?((((~m[59]&~m[383]&~m[527])|(m[59]&m[383]&~m[527]))&BiasedRNG[167])|(((m[59]&~m[383]&~m[527])|(~m[59]&m[383]&m[527]))&~BiasedRNG[167])|((~m[59]&~m[383]&m[527])|(m[59]&~m[383]&m[527])|(m[59]&m[383]&m[527]))):InitCond[167];
    m[528] = run?((((m[385]&~m[529]&~m[530]&~m[531]&~m[532])|(~m[385]&~m[529]&~m[530]&m[531]&~m[532])|(m[385]&m[529]&~m[530]&m[531]&~m[532])|(m[385]&~m[529]&m[530]&m[531]&~m[532])|(~m[385]&m[529]&~m[530]&~m[531]&m[532])|(~m[385]&~m[529]&m[530]&~m[531]&m[532])|(m[385]&m[529]&m[530]&~m[531]&m[532])|(~m[385]&m[529]&m[530]&m[531]&m[532]))&UnbiasedRNG[0])|((m[385]&~m[529]&~m[530]&m[531]&~m[532])|(~m[385]&~m[529]&~m[530]&~m[531]&m[532])|(m[385]&~m[529]&~m[530]&~m[531]&m[532])|(m[385]&m[529]&~m[530]&~m[531]&m[532])|(m[385]&~m[529]&m[530]&~m[531]&m[532])|(~m[385]&~m[529]&~m[530]&m[531]&m[532])|(m[385]&~m[529]&~m[530]&m[531]&m[532])|(~m[385]&m[529]&~m[530]&m[531]&m[532])|(m[385]&m[529]&~m[530]&m[531]&m[532])|(~m[385]&~m[529]&m[530]&m[531]&m[532])|(m[385]&~m[529]&m[530]&m[531]&m[532])|(m[385]&m[529]&m[530]&m[531]&m[532]))):InitCond[168];
    m[533] = run?((((m[386]&~m[534]&~m[535]&~m[536]&~m[537])|(~m[386]&~m[534]&~m[535]&m[536]&~m[537])|(m[386]&m[534]&~m[535]&m[536]&~m[537])|(m[386]&~m[534]&m[535]&m[536]&~m[537])|(~m[386]&m[534]&~m[535]&~m[536]&m[537])|(~m[386]&~m[534]&m[535]&~m[536]&m[537])|(m[386]&m[534]&m[535]&~m[536]&m[537])|(~m[386]&m[534]&m[535]&m[536]&m[537]))&UnbiasedRNG[1])|((m[386]&~m[534]&~m[535]&m[536]&~m[537])|(~m[386]&~m[534]&~m[535]&~m[536]&m[537])|(m[386]&~m[534]&~m[535]&~m[536]&m[537])|(m[386]&m[534]&~m[535]&~m[536]&m[537])|(m[386]&~m[534]&m[535]&~m[536]&m[537])|(~m[386]&~m[534]&~m[535]&m[536]&m[537])|(m[386]&~m[534]&~m[535]&m[536]&m[537])|(~m[386]&m[534]&~m[535]&m[536]&m[537])|(m[386]&m[534]&~m[535]&m[536]&m[537])|(~m[386]&~m[534]&m[535]&m[536]&m[537])|(m[386]&~m[534]&m[535]&m[536]&m[537])|(m[386]&m[534]&m[535]&m[536]&m[537]))):InitCond[169];
    m[538] = run?((((m[536]&~m[539]&~m[540]&~m[541]&~m[542])|(~m[536]&~m[539]&~m[540]&m[541]&~m[542])|(m[536]&m[539]&~m[540]&m[541]&~m[542])|(m[536]&~m[539]&m[540]&m[541]&~m[542])|(~m[536]&m[539]&~m[540]&~m[541]&m[542])|(~m[536]&~m[539]&m[540]&~m[541]&m[542])|(m[536]&m[539]&m[540]&~m[541]&m[542])|(~m[536]&m[539]&m[540]&m[541]&m[542]))&UnbiasedRNG[2])|((m[536]&~m[539]&~m[540]&m[541]&~m[542])|(~m[536]&~m[539]&~m[540]&~m[541]&m[542])|(m[536]&~m[539]&~m[540]&~m[541]&m[542])|(m[536]&m[539]&~m[540]&~m[541]&m[542])|(m[536]&~m[539]&m[540]&~m[541]&m[542])|(~m[536]&~m[539]&~m[540]&m[541]&m[542])|(m[536]&~m[539]&~m[540]&m[541]&m[542])|(~m[536]&m[539]&~m[540]&m[541]&m[542])|(m[536]&m[539]&~m[540]&m[541]&m[542])|(~m[536]&~m[539]&m[540]&m[541]&m[542])|(m[536]&~m[539]&m[540]&m[541]&m[542])|(m[536]&m[539]&m[540]&m[541]&m[542]))):InitCond[170];
    m[543] = run?((((m[387]&~m[544]&~m[545]&~m[546]&~m[547])|(~m[387]&~m[544]&~m[545]&m[546]&~m[547])|(m[387]&m[544]&~m[545]&m[546]&~m[547])|(m[387]&~m[544]&m[545]&m[546]&~m[547])|(~m[387]&m[544]&~m[545]&~m[546]&m[547])|(~m[387]&~m[544]&m[545]&~m[546]&m[547])|(m[387]&m[544]&m[545]&~m[546]&m[547])|(~m[387]&m[544]&m[545]&m[546]&m[547]))&UnbiasedRNG[3])|((m[387]&~m[544]&~m[545]&m[546]&~m[547])|(~m[387]&~m[544]&~m[545]&~m[546]&m[547])|(m[387]&~m[544]&~m[545]&~m[546]&m[547])|(m[387]&m[544]&~m[545]&~m[546]&m[547])|(m[387]&~m[544]&m[545]&~m[546]&m[547])|(~m[387]&~m[544]&~m[545]&m[546]&m[547])|(m[387]&~m[544]&~m[545]&m[546]&m[547])|(~m[387]&m[544]&~m[545]&m[546]&m[547])|(m[387]&m[544]&~m[545]&m[546]&m[547])|(~m[387]&~m[544]&m[545]&m[546]&m[547])|(m[387]&~m[544]&m[545]&m[546]&m[547])|(m[387]&m[544]&m[545]&m[546]&m[547]))):InitCond[171];
    m[548] = run?((((m[546]&~m[549]&~m[550]&~m[551]&~m[552])|(~m[546]&~m[549]&~m[550]&m[551]&~m[552])|(m[546]&m[549]&~m[550]&m[551]&~m[552])|(m[546]&~m[549]&m[550]&m[551]&~m[552])|(~m[546]&m[549]&~m[550]&~m[551]&m[552])|(~m[546]&~m[549]&m[550]&~m[551]&m[552])|(m[546]&m[549]&m[550]&~m[551]&m[552])|(~m[546]&m[549]&m[550]&m[551]&m[552]))&UnbiasedRNG[4])|((m[546]&~m[549]&~m[550]&m[551]&~m[552])|(~m[546]&~m[549]&~m[550]&~m[551]&m[552])|(m[546]&~m[549]&~m[550]&~m[551]&m[552])|(m[546]&m[549]&~m[550]&~m[551]&m[552])|(m[546]&~m[549]&m[550]&~m[551]&m[552])|(~m[546]&~m[549]&~m[550]&m[551]&m[552])|(m[546]&~m[549]&~m[550]&m[551]&m[552])|(~m[546]&m[549]&~m[550]&m[551]&m[552])|(m[546]&m[549]&~m[550]&m[551]&m[552])|(~m[546]&~m[549]&m[550]&m[551]&m[552])|(m[546]&~m[549]&m[550]&m[551]&m[552])|(m[546]&m[549]&m[550]&m[551]&m[552]))):InitCond[172];
    m[553] = run?((((m[551]&~m[554]&~m[555]&~m[556]&~m[557])|(~m[551]&~m[554]&~m[555]&m[556]&~m[557])|(m[551]&m[554]&~m[555]&m[556]&~m[557])|(m[551]&~m[554]&m[555]&m[556]&~m[557])|(~m[551]&m[554]&~m[555]&~m[556]&m[557])|(~m[551]&~m[554]&m[555]&~m[556]&m[557])|(m[551]&m[554]&m[555]&~m[556]&m[557])|(~m[551]&m[554]&m[555]&m[556]&m[557]))&UnbiasedRNG[5])|((m[551]&~m[554]&~m[555]&m[556]&~m[557])|(~m[551]&~m[554]&~m[555]&~m[556]&m[557])|(m[551]&~m[554]&~m[555]&~m[556]&m[557])|(m[551]&m[554]&~m[555]&~m[556]&m[557])|(m[551]&~m[554]&m[555]&~m[556]&m[557])|(~m[551]&~m[554]&~m[555]&m[556]&m[557])|(m[551]&~m[554]&~m[555]&m[556]&m[557])|(~m[551]&m[554]&~m[555]&m[556]&m[557])|(m[551]&m[554]&~m[555]&m[556]&m[557])|(~m[551]&~m[554]&m[555]&m[556]&m[557])|(m[551]&~m[554]&m[555]&m[556]&m[557])|(m[551]&m[554]&m[555]&m[556]&m[557]))):InitCond[173];
    m[558] = run?((((m[388]&~m[559]&~m[560]&~m[561]&~m[562])|(~m[388]&~m[559]&~m[560]&m[561]&~m[562])|(m[388]&m[559]&~m[560]&m[561]&~m[562])|(m[388]&~m[559]&m[560]&m[561]&~m[562])|(~m[388]&m[559]&~m[560]&~m[561]&m[562])|(~m[388]&~m[559]&m[560]&~m[561]&m[562])|(m[388]&m[559]&m[560]&~m[561]&m[562])|(~m[388]&m[559]&m[560]&m[561]&m[562]))&UnbiasedRNG[6])|((m[388]&~m[559]&~m[560]&m[561]&~m[562])|(~m[388]&~m[559]&~m[560]&~m[561]&m[562])|(m[388]&~m[559]&~m[560]&~m[561]&m[562])|(m[388]&m[559]&~m[560]&~m[561]&m[562])|(m[388]&~m[559]&m[560]&~m[561]&m[562])|(~m[388]&~m[559]&~m[560]&m[561]&m[562])|(m[388]&~m[559]&~m[560]&m[561]&m[562])|(~m[388]&m[559]&~m[560]&m[561]&m[562])|(m[388]&m[559]&~m[560]&m[561]&m[562])|(~m[388]&~m[559]&m[560]&m[561]&m[562])|(m[388]&~m[559]&m[560]&m[561]&m[562])|(m[388]&m[559]&m[560]&m[561]&m[562]))):InitCond[174];
    m[563] = run?((((m[561]&~m[564]&~m[565]&~m[566]&~m[567])|(~m[561]&~m[564]&~m[565]&m[566]&~m[567])|(m[561]&m[564]&~m[565]&m[566]&~m[567])|(m[561]&~m[564]&m[565]&m[566]&~m[567])|(~m[561]&m[564]&~m[565]&~m[566]&m[567])|(~m[561]&~m[564]&m[565]&~m[566]&m[567])|(m[561]&m[564]&m[565]&~m[566]&m[567])|(~m[561]&m[564]&m[565]&m[566]&m[567]))&UnbiasedRNG[7])|((m[561]&~m[564]&~m[565]&m[566]&~m[567])|(~m[561]&~m[564]&~m[565]&~m[566]&m[567])|(m[561]&~m[564]&~m[565]&~m[566]&m[567])|(m[561]&m[564]&~m[565]&~m[566]&m[567])|(m[561]&~m[564]&m[565]&~m[566]&m[567])|(~m[561]&~m[564]&~m[565]&m[566]&m[567])|(m[561]&~m[564]&~m[565]&m[566]&m[567])|(~m[561]&m[564]&~m[565]&m[566]&m[567])|(m[561]&m[564]&~m[565]&m[566]&m[567])|(~m[561]&~m[564]&m[565]&m[566]&m[567])|(m[561]&~m[564]&m[565]&m[566]&m[567])|(m[561]&m[564]&m[565]&m[566]&m[567]))):InitCond[175];
    m[568] = run?((((m[566]&~m[569]&~m[570]&~m[571]&~m[572])|(~m[566]&~m[569]&~m[570]&m[571]&~m[572])|(m[566]&m[569]&~m[570]&m[571]&~m[572])|(m[566]&~m[569]&m[570]&m[571]&~m[572])|(~m[566]&m[569]&~m[570]&~m[571]&m[572])|(~m[566]&~m[569]&m[570]&~m[571]&m[572])|(m[566]&m[569]&m[570]&~m[571]&m[572])|(~m[566]&m[569]&m[570]&m[571]&m[572]))&UnbiasedRNG[8])|((m[566]&~m[569]&~m[570]&m[571]&~m[572])|(~m[566]&~m[569]&~m[570]&~m[571]&m[572])|(m[566]&~m[569]&~m[570]&~m[571]&m[572])|(m[566]&m[569]&~m[570]&~m[571]&m[572])|(m[566]&~m[569]&m[570]&~m[571]&m[572])|(~m[566]&~m[569]&~m[570]&m[571]&m[572])|(m[566]&~m[569]&~m[570]&m[571]&m[572])|(~m[566]&m[569]&~m[570]&m[571]&m[572])|(m[566]&m[569]&~m[570]&m[571]&m[572])|(~m[566]&~m[569]&m[570]&m[571]&m[572])|(m[566]&~m[569]&m[570]&m[571]&m[572])|(m[566]&m[569]&m[570]&m[571]&m[572]))):InitCond[176];
    m[573] = run?((((m[571]&~m[574]&~m[575]&~m[576]&~m[577])|(~m[571]&~m[574]&~m[575]&m[576]&~m[577])|(m[571]&m[574]&~m[575]&m[576]&~m[577])|(m[571]&~m[574]&m[575]&m[576]&~m[577])|(~m[571]&m[574]&~m[575]&~m[576]&m[577])|(~m[571]&~m[574]&m[575]&~m[576]&m[577])|(m[571]&m[574]&m[575]&~m[576]&m[577])|(~m[571]&m[574]&m[575]&m[576]&m[577]))&UnbiasedRNG[9])|((m[571]&~m[574]&~m[575]&m[576]&~m[577])|(~m[571]&~m[574]&~m[575]&~m[576]&m[577])|(m[571]&~m[574]&~m[575]&~m[576]&m[577])|(m[571]&m[574]&~m[575]&~m[576]&m[577])|(m[571]&~m[574]&m[575]&~m[576]&m[577])|(~m[571]&~m[574]&~m[575]&m[576]&m[577])|(m[571]&~m[574]&~m[575]&m[576]&m[577])|(~m[571]&m[574]&~m[575]&m[576]&m[577])|(m[571]&m[574]&~m[575]&m[576]&m[577])|(~m[571]&~m[574]&m[575]&m[576]&m[577])|(m[571]&~m[574]&m[575]&m[576]&m[577])|(m[571]&m[574]&m[575]&m[576]&m[577]))):InitCond[177];
    m[578] = run?((((m[389]&~m[579]&~m[580]&~m[581]&~m[582])|(~m[389]&~m[579]&~m[580]&m[581]&~m[582])|(m[389]&m[579]&~m[580]&m[581]&~m[582])|(m[389]&~m[579]&m[580]&m[581]&~m[582])|(~m[389]&m[579]&~m[580]&~m[581]&m[582])|(~m[389]&~m[579]&m[580]&~m[581]&m[582])|(m[389]&m[579]&m[580]&~m[581]&m[582])|(~m[389]&m[579]&m[580]&m[581]&m[582]))&UnbiasedRNG[10])|((m[389]&~m[579]&~m[580]&m[581]&~m[582])|(~m[389]&~m[579]&~m[580]&~m[581]&m[582])|(m[389]&~m[579]&~m[580]&~m[581]&m[582])|(m[389]&m[579]&~m[580]&~m[581]&m[582])|(m[389]&~m[579]&m[580]&~m[581]&m[582])|(~m[389]&~m[579]&~m[580]&m[581]&m[582])|(m[389]&~m[579]&~m[580]&m[581]&m[582])|(~m[389]&m[579]&~m[580]&m[581]&m[582])|(m[389]&m[579]&~m[580]&m[581]&m[582])|(~m[389]&~m[579]&m[580]&m[581]&m[582])|(m[389]&~m[579]&m[580]&m[581]&m[582])|(m[389]&m[579]&m[580]&m[581]&m[582]))):InitCond[178];
    m[583] = run?((((m[581]&~m[584]&~m[585]&~m[586]&~m[587])|(~m[581]&~m[584]&~m[585]&m[586]&~m[587])|(m[581]&m[584]&~m[585]&m[586]&~m[587])|(m[581]&~m[584]&m[585]&m[586]&~m[587])|(~m[581]&m[584]&~m[585]&~m[586]&m[587])|(~m[581]&~m[584]&m[585]&~m[586]&m[587])|(m[581]&m[584]&m[585]&~m[586]&m[587])|(~m[581]&m[584]&m[585]&m[586]&m[587]))&UnbiasedRNG[11])|((m[581]&~m[584]&~m[585]&m[586]&~m[587])|(~m[581]&~m[584]&~m[585]&~m[586]&m[587])|(m[581]&~m[584]&~m[585]&~m[586]&m[587])|(m[581]&m[584]&~m[585]&~m[586]&m[587])|(m[581]&~m[584]&m[585]&~m[586]&m[587])|(~m[581]&~m[584]&~m[585]&m[586]&m[587])|(m[581]&~m[584]&~m[585]&m[586]&m[587])|(~m[581]&m[584]&~m[585]&m[586]&m[587])|(m[581]&m[584]&~m[585]&m[586]&m[587])|(~m[581]&~m[584]&m[585]&m[586]&m[587])|(m[581]&~m[584]&m[585]&m[586]&m[587])|(m[581]&m[584]&m[585]&m[586]&m[587]))):InitCond[179];
    m[588] = run?((((m[586]&~m[589]&~m[590]&~m[591]&~m[592])|(~m[586]&~m[589]&~m[590]&m[591]&~m[592])|(m[586]&m[589]&~m[590]&m[591]&~m[592])|(m[586]&~m[589]&m[590]&m[591]&~m[592])|(~m[586]&m[589]&~m[590]&~m[591]&m[592])|(~m[586]&~m[589]&m[590]&~m[591]&m[592])|(m[586]&m[589]&m[590]&~m[591]&m[592])|(~m[586]&m[589]&m[590]&m[591]&m[592]))&UnbiasedRNG[12])|((m[586]&~m[589]&~m[590]&m[591]&~m[592])|(~m[586]&~m[589]&~m[590]&~m[591]&m[592])|(m[586]&~m[589]&~m[590]&~m[591]&m[592])|(m[586]&m[589]&~m[590]&~m[591]&m[592])|(m[586]&~m[589]&m[590]&~m[591]&m[592])|(~m[586]&~m[589]&~m[590]&m[591]&m[592])|(m[586]&~m[589]&~m[590]&m[591]&m[592])|(~m[586]&m[589]&~m[590]&m[591]&m[592])|(m[586]&m[589]&~m[590]&m[591]&m[592])|(~m[586]&~m[589]&m[590]&m[591]&m[592])|(m[586]&~m[589]&m[590]&m[591]&m[592])|(m[586]&m[589]&m[590]&m[591]&m[592]))):InitCond[180];
    m[593] = run?((((m[591]&~m[594]&~m[595]&~m[596]&~m[597])|(~m[591]&~m[594]&~m[595]&m[596]&~m[597])|(m[591]&m[594]&~m[595]&m[596]&~m[597])|(m[591]&~m[594]&m[595]&m[596]&~m[597])|(~m[591]&m[594]&~m[595]&~m[596]&m[597])|(~m[591]&~m[594]&m[595]&~m[596]&m[597])|(m[591]&m[594]&m[595]&~m[596]&m[597])|(~m[591]&m[594]&m[595]&m[596]&m[597]))&UnbiasedRNG[13])|((m[591]&~m[594]&~m[595]&m[596]&~m[597])|(~m[591]&~m[594]&~m[595]&~m[596]&m[597])|(m[591]&~m[594]&~m[595]&~m[596]&m[597])|(m[591]&m[594]&~m[595]&~m[596]&m[597])|(m[591]&~m[594]&m[595]&~m[596]&m[597])|(~m[591]&~m[594]&~m[595]&m[596]&m[597])|(m[591]&~m[594]&~m[595]&m[596]&m[597])|(~m[591]&m[594]&~m[595]&m[596]&m[597])|(m[591]&m[594]&~m[595]&m[596]&m[597])|(~m[591]&~m[594]&m[595]&m[596]&m[597])|(m[591]&~m[594]&m[595]&m[596]&m[597])|(m[591]&m[594]&m[595]&m[596]&m[597]))):InitCond[181];
    m[598] = run?((((m[596]&~m[599]&~m[600]&~m[601]&~m[602])|(~m[596]&~m[599]&~m[600]&m[601]&~m[602])|(m[596]&m[599]&~m[600]&m[601]&~m[602])|(m[596]&~m[599]&m[600]&m[601]&~m[602])|(~m[596]&m[599]&~m[600]&~m[601]&m[602])|(~m[596]&~m[599]&m[600]&~m[601]&m[602])|(m[596]&m[599]&m[600]&~m[601]&m[602])|(~m[596]&m[599]&m[600]&m[601]&m[602]))&UnbiasedRNG[14])|((m[596]&~m[599]&~m[600]&m[601]&~m[602])|(~m[596]&~m[599]&~m[600]&~m[601]&m[602])|(m[596]&~m[599]&~m[600]&~m[601]&m[602])|(m[596]&m[599]&~m[600]&~m[601]&m[602])|(m[596]&~m[599]&m[600]&~m[601]&m[602])|(~m[596]&~m[599]&~m[600]&m[601]&m[602])|(m[596]&~m[599]&~m[600]&m[601]&m[602])|(~m[596]&m[599]&~m[600]&m[601]&m[602])|(m[596]&m[599]&~m[600]&m[601]&m[602])|(~m[596]&~m[599]&m[600]&m[601]&m[602])|(m[596]&~m[599]&m[600]&m[601]&m[602])|(m[596]&m[599]&m[600]&m[601]&m[602]))):InitCond[182];
    m[603] = run?((((m[390]&~m[604]&~m[605]&~m[606]&~m[607])|(~m[390]&~m[604]&~m[605]&m[606]&~m[607])|(m[390]&m[604]&~m[605]&m[606]&~m[607])|(m[390]&~m[604]&m[605]&m[606]&~m[607])|(~m[390]&m[604]&~m[605]&~m[606]&m[607])|(~m[390]&~m[604]&m[605]&~m[606]&m[607])|(m[390]&m[604]&m[605]&~m[606]&m[607])|(~m[390]&m[604]&m[605]&m[606]&m[607]))&UnbiasedRNG[15])|((m[390]&~m[604]&~m[605]&m[606]&~m[607])|(~m[390]&~m[604]&~m[605]&~m[606]&m[607])|(m[390]&~m[604]&~m[605]&~m[606]&m[607])|(m[390]&m[604]&~m[605]&~m[606]&m[607])|(m[390]&~m[604]&m[605]&~m[606]&m[607])|(~m[390]&~m[604]&~m[605]&m[606]&m[607])|(m[390]&~m[604]&~m[605]&m[606]&m[607])|(~m[390]&m[604]&~m[605]&m[606]&m[607])|(m[390]&m[604]&~m[605]&m[606]&m[607])|(~m[390]&~m[604]&m[605]&m[606]&m[607])|(m[390]&~m[604]&m[605]&m[606]&m[607])|(m[390]&m[604]&m[605]&m[606]&m[607]))):InitCond[183];
    m[608] = run?((((m[606]&~m[609]&~m[610]&~m[611]&~m[612])|(~m[606]&~m[609]&~m[610]&m[611]&~m[612])|(m[606]&m[609]&~m[610]&m[611]&~m[612])|(m[606]&~m[609]&m[610]&m[611]&~m[612])|(~m[606]&m[609]&~m[610]&~m[611]&m[612])|(~m[606]&~m[609]&m[610]&~m[611]&m[612])|(m[606]&m[609]&m[610]&~m[611]&m[612])|(~m[606]&m[609]&m[610]&m[611]&m[612]))&UnbiasedRNG[16])|((m[606]&~m[609]&~m[610]&m[611]&~m[612])|(~m[606]&~m[609]&~m[610]&~m[611]&m[612])|(m[606]&~m[609]&~m[610]&~m[611]&m[612])|(m[606]&m[609]&~m[610]&~m[611]&m[612])|(m[606]&~m[609]&m[610]&~m[611]&m[612])|(~m[606]&~m[609]&~m[610]&m[611]&m[612])|(m[606]&~m[609]&~m[610]&m[611]&m[612])|(~m[606]&m[609]&~m[610]&m[611]&m[612])|(m[606]&m[609]&~m[610]&m[611]&m[612])|(~m[606]&~m[609]&m[610]&m[611]&m[612])|(m[606]&~m[609]&m[610]&m[611]&m[612])|(m[606]&m[609]&m[610]&m[611]&m[612]))):InitCond[184];
    m[613] = run?((((m[611]&~m[614]&~m[615]&~m[616]&~m[617])|(~m[611]&~m[614]&~m[615]&m[616]&~m[617])|(m[611]&m[614]&~m[615]&m[616]&~m[617])|(m[611]&~m[614]&m[615]&m[616]&~m[617])|(~m[611]&m[614]&~m[615]&~m[616]&m[617])|(~m[611]&~m[614]&m[615]&~m[616]&m[617])|(m[611]&m[614]&m[615]&~m[616]&m[617])|(~m[611]&m[614]&m[615]&m[616]&m[617]))&UnbiasedRNG[17])|((m[611]&~m[614]&~m[615]&m[616]&~m[617])|(~m[611]&~m[614]&~m[615]&~m[616]&m[617])|(m[611]&~m[614]&~m[615]&~m[616]&m[617])|(m[611]&m[614]&~m[615]&~m[616]&m[617])|(m[611]&~m[614]&m[615]&~m[616]&m[617])|(~m[611]&~m[614]&~m[615]&m[616]&m[617])|(m[611]&~m[614]&~m[615]&m[616]&m[617])|(~m[611]&m[614]&~m[615]&m[616]&m[617])|(m[611]&m[614]&~m[615]&m[616]&m[617])|(~m[611]&~m[614]&m[615]&m[616]&m[617])|(m[611]&~m[614]&m[615]&m[616]&m[617])|(m[611]&m[614]&m[615]&m[616]&m[617]))):InitCond[185];
    m[618] = run?((((m[616]&~m[619]&~m[620]&~m[621]&~m[622])|(~m[616]&~m[619]&~m[620]&m[621]&~m[622])|(m[616]&m[619]&~m[620]&m[621]&~m[622])|(m[616]&~m[619]&m[620]&m[621]&~m[622])|(~m[616]&m[619]&~m[620]&~m[621]&m[622])|(~m[616]&~m[619]&m[620]&~m[621]&m[622])|(m[616]&m[619]&m[620]&~m[621]&m[622])|(~m[616]&m[619]&m[620]&m[621]&m[622]))&UnbiasedRNG[18])|((m[616]&~m[619]&~m[620]&m[621]&~m[622])|(~m[616]&~m[619]&~m[620]&~m[621]&m[622])|(m[616]&~m[619]&~m[620]&~m[621]&m[622])|(m[616]&m[619]&~m[620]&~m[621]&m[622])|(m[616]&~m[619]&m[620]&~m[621]&m[622])|(~m[616]&~m[619]&~m[620]&m[621]&m[622])|(m[616]&~m[619]&~m[620]&m[621]&m[622])|(~m[616]&m[619]&~m[620]&m[621]&m[622])|(m[616]&m[619]&~m[620]&m[621]&m[622])|(~m[616]&~m[619]&m[620]&m[621]&m[622])|(m[616]&~m[619]&m[620]&m[621]&m[622])|(m[616]&m[619]&m[620]&m[621]&m[622]))):InitCond[186];
    m[623] = run?((((m[621]&~m[624]&~m[625]&~m[626]&~m[627])|(~m[621]&~m[624]&~m[625]&m[626]&~m[627])|(m[621]&m[624]&~m[625]&m[626]&~m[627])|(m[621]&~m[624]&m[625]&m[626]&~m[627])|(~m[621]&m[624]&~m[625]&~m[626]&m[627])|(~m[621]&~m[624]&m[625]&~m[626]&m[627])|(m[621]&m[624]&m[625]&~m[626]&m[627])|(~m[621]&m[624]&m[625]&m[626]&m[627]))&UnbiasedRNG[19])|((m[621]&~m[624]&~m[625]&m[626]&~m[627])|(~m[621]&~m[624]&~m[625]&~m[626]&m[627])|(m[621]&~m[624]&~m[625]&~m[626]&m[627])|(m[621]&m[624]&~m[625]&~m[626]&m[627])|(m[621]&~m[624]&m[625]&~m[626]&m[627])|(~m[621]&~m[624]&~m[625]&m[626]&m[627])|(m[621]&~m[624]&~m[625]&m[626]&m[627])|(~m[621]&m[624]&~m[625]&m[626]&m[627])|(m[621]&m[624]&~m[625]&m[626]&m[627])|(~m[621]&~m[624]&m[625]&m[626]&m[627])|(m[621]&~m[624]&m[625]&m[626]&m[627])|(m[621]&m[624]&m[625]&m[626]&m[627]))):InitCond[187];
    m[628] = run?((((m[626]&~m[629]&~m[630]&~m[631]&~m[632])|(~m[626]&~m[629]&~m[630]&m[631]&~m[632])|(m[626]&m[629]&~m[630]&m[631]&~m[632])|(m[626]&~m[629]&m[630]&m[631]&~m[632])|(~m[626]&m[629]&~m[630]&~m[631]&m[632])|(~m[626]&~m[629]&m[630]&~m[631]&m[632])|(m[626]&m[629]&m[630]&~m[631]&m[632])|(~m[626]&m[629]&m[630]&m[631]&m[632]))&UnbiasedRNG[20])|((m[626]&~m[629]&~m[630]&m[631]&~m[632])|(~m[626]&~m[629]&~m[630]&~m[631]&m[632])|(m[626]&~m[629]&~m[630]&~m[631]&m[632])|(m[626]&m[629]&~m[630]&~m[631]&m[632])|(m[626]&~m[629]&m[630]&~m[631]&m[632])|(~m[626]&~m[629]&~m[630]&m[631]&m[632])|(m[626]&~m[629]&~m[630]&m[631]&m[632])|(~m[626]&m[629]&~m[630]&m[631]&m[632])|(m[626]&m[629]&~m[630]&m[631]&m[632])|(~m[626]&~m[629]&m[630]&m[631]&m[632])|(m[626]&~m[629]&m[630]&m[631]&m[632])|(m[626]&m[629]&m[630]&m[631]&m[632]))):InitCond[188];
    m[633] = run?((((m[391]&~m[634]&~m[635]&~m[636]&~m[637])|(~m[391]&~m[634]&~m[635]&m[636]&~m[637])|(m[391]&m[634]&~m[635]&m[636]&~m[637])|(m[391]&~m[634]&m[635]&m[636]&~m[637])|(~m[391]&m[634]&~m[635]&~m[636]&m[637])|(~m[391]&~m[634]&m[635]&~m[636]&m[637])|(m[391]&m[634]&m[635]&~m[636]&m[637])|(~m[391]&m[634]&m[635]&m[636]&m[637]))&UnbiasedRNG[21])|((m[391]&~m[634]&~m[635]&m[636]&~m[637])|(~m[391]&~m[634]&~m[635]&~m[636]&m[637])|(m[391]&~m[634]&~m[635]&~m[636]&m[637])|(m[391]&m[634]&~m[635]&~m[636]&m[637])|(m[391]&~m[634]&m[635]&~m[636]&m[637])|(~m[391]&~m[634]&~m[635]&m[636]&m[637])|(m[391]&~m[634]&~m[635]&m[636]&m[637])|(~m[391]&m[634]&~m[635]&m[636]&m[637])|(m[391]&m[634]&~m[635]&m[636]&m[637])|(~m[391]&~m[634]&m[635]&m[636]&m[637])|(m[391]&~m[634]&m[635]&m[636]&m[637])|(m[391]&m[634]&m[635]&m[636]&m[637]))):InitCond[189];
    m[638] = run?((((m[636]&~m[639]&~m[640]&~m[641]&~m[642])|(~m[636]&~m[639]&~m[640]&m[641]&~m[642])|(m[636]&m[639]&~m[640]&m[641]&~m[642])|(m[636]&~m[639]&m[640]&m[641]&~m[642])|(~m[636]&m[639]&~m[640]&~m[641]&m[642])|(~m[636]&~m[639]&m[640]&~m[641]&m[642])|(m[636]&m[639]&m[640]&~m[641]&m[642])|(~m[636]&m[639]&m[640]&m[641]&m[642]))&UnbiasedRNG[22])|((m[636]&~m[639]&~m[640]&m[641]&~m[642])|(~m[636]&~m[639]&~m[640]&~m[641]&m[642])|(m[636]&~m[639]&~m[640]&~m[641]&m[642])|(m[636]&m[639]&~m[640]&~m[641]&m[642])|(m[636]&~m[639]&m[640]&~m[641]&m[642])|(~m[636]&~m[639]&~m[640]&m[641]&m[642])|(m[636]&~m[639]&~m[640]&m[641]&m[642])|(~m[636]&m[639]&~m[640]&m[641]&m[642])|(m[636]&m[639]&~m[640]&m[641]&m[642])|(~m[636]&~m[639]&m[640]&m[641]&m[642])|(m[636]&~m[639]&m[640]&m[641]&m[642])|(m[636]&m[639]&m[640]&m[641]&m[642]))):InitCond[190];
    m[643] = run?((((m[641]&~m[644]&~m[645]&~m[646]&~m[647])|(~m[641]&~m[644]&~m[645]&m[646]&~m[647])|(m[641]&m[644]&~m[645]&m[646]&~m[647])|(m[641]&~m[644]&m[645]&m[646]&~m[647])|(~m[641]&m[644]&~m[645]&~m[646]&m[647])|(~m[641]&~m[644]&m[645]&~m[646]&m[647])|(m[641]&m[644]&m[645]&~m[646]&m[647])|(~m[641]&m[644]&m[645]&m[646]&m[647]))&UnbiasedRNG[23])|((m[641]&~m[644]&~m[645]&m[646]&~m[647])|(~m[641]&~m[644]&~m[645]&~m[646]&m[647])|(m[641]&~m[644]&~m[645]&~m[646]&m[647])|(m[641]&m[644]&~m[645]&~m[646]&m[647])|(m[641]&~m[644]&m[645]&~m[646]&m[647])|(~m[641]&~m[644]&~m[645]&m[646]&m[647])|(m[641]&~m[644]&~m[645]&m[646]&m[647])|(~m[641]&m[644]&~m[645]&m[646]&m[647])|(m[641]&m[644]&~m[645]&m[646]&m[647])|(~m[641]&~m[644]&m[645]&m[646]&m[647])|(m[641]&~m[644]&m[645]&m[646]&m[647])|(m[641]&m[644]&m[645]&m[646]&m[647]))):InitCond[191];
    m[648] = run?((((m[646]&~m[649]&~m[650]&~m[651]&~m[652])|(~m[646]&~m[649]&~m[650]&m[651]&~m[652])|(m[646]&m[649]&~m[650]&m[651]&~m[652])|(m[646]&~m[649]&m[650]&m[651]&~m[652])|(~m[646]&m[649]&~m[650]&~m[651]&m[652])|(~m[646]&~m[649]&m[650]&~m[651]&m[652])|(m[646]&m[649]&m[650]&~m[651]&m[652])|(~m[646]&m[649]&m[650]&m[651]&m[652]))&UnbiasedRNG[24])|((m[646]&~m[649]&~m[650]&m[651]&~m[652])|(~m[646]&~m[649]&~m[650]&~m[651]&m[652])|(m[646]&~m[649]&~m[650]&~m[651]&m[652])|(m[646]&m[649]&~m[650]&~m[651]&m[652])|(m[646]&~m[649]&m[650]&~m[651]&m[652])|(~m[646]&~m[649]&~m[650]&m[651]&m[652])|(m[646]&~m[649]&~m[650]&m[651]&m[652])|(~m[646]&m[649]&~m[650]&m[651]&m[652])|(m[646]&m[649]&~m[650]&m[651]&m[652])|(~m[646]&~m[649]&m[650]&m[651]&m[652])|(m[646]&~m[649]&m[650]&m[651]&m[652])|(m[646]&m[649]&m[650]&m[651]&m[652]))):InitCond[192];
    m[653] = run?((((m[651]&~m[654]&~m[655]&~m[656]&~m[657])|(~m[651]&~m[654]&~m[655]&m[656]&~m[657])|(m[651]&m[654]&~m[655]&m[656]&~m[657])|(m[651]&~m[654]&m[655]&m[656]&~m[657])|(~m[651]&m[654]&~m[655]&~m[656]&m[657])|(~m[651]&~m[654]&m[655]&~m[656]&m[657])|(m[651]&m[654]&m[655]&~m[656]&m[657])|(~m[651]&m[654]&m[655]&m[656]&m[657]))&UnbiasedRNG[25])|((m[651]&~m[654]&~m[655]&m[656]&~m[657])|(~m[651]&~m[654]&~m[655]&~m[656]&m[657])|(m[651]&~m[654]&~m[655]&~m[656]&m[657])|(m[651]&m[654]&~m[655]&~m[656]&m[657])|(m[651]&~m[654]&m[655]&~m[656]&m[657])|(~m[651]&~m[654]&~m[655]&m[656]&m[657])|(m[651]&~m[654]&~m[655]&m[656]&m[657])|(~m[651]&m[654]&~m[655]&m[656]&m[657])|(m[651]&m[654]&~m[655]&m[656]&m[657])|(~m[651]&~m[654]&m[655]&m[656]&m[657])|(m[651]&~m[654]&m[655]&m[656]&m[657])|(m[651]&m[654]&m[655]&m[656]&m[657]))):InitCond[193];
    m[658] = run?((((m[656]&~m[659]&~m[660]&~m[661]&~m[662])|(~m[656]&~m[659]&~m[660]&m[661]&~m[662])|(m[656]&m[659]&~m[660]&m[661]&~m[662])|(m[656]&~m[659]&m[660]&m[661]&~m[662])|(~m[656]&m[659]&~m[660]&~m[661]&m[662])|(~m[656]&~m[659]&m[660]&~m[661]&m[662])|(m[656]&m[659]&m[660]&~m[661]&m[662])|(~m[656]&m[659]&m[660]&m[661]&m[662]))&UnbiasedRNG[26])|((m[656]&~m[659]&~m[660]&m[661]&~m[662])|(~m[656]&~m[659]&~m[660]&~m[661]&m[662])|(m[656]&~m[659]&~m[660]&~m[661]&m[662])|(m[656]&m[659]&~m[660]&~m[661]&m[662])|(m[656]&~m[659]&m[660]&~m[661]&m[662])|(~m[656]&~m[659]&~m[660]&m[661]&m[662])|(m[656]&~m[659]&~m[660]&m[661]&m[662])|(~m[656]&m[659]&~m[660]&m[661]&m[662])|(m[656]&m[659]&~m[660]&m[661]&m[662])|(~m[656]&~m[659]&m[660]&m[661]&m[662])|(m[656]&~m[659]&m[660]&m[661]&m[662])|(m[656]&m[659]&m[660]&m[661]&m[662]))):InitCond[194];
    m[663] = run?((((m[661]&~m[664]&~m[665]&~m[666]&~m[667])|(~m[661]&~m[664]&~m[665]&m[666]&~m[667])|(m[661]&m[664]&~m[665]&m[666]&~m[667])|(m[661]&~m[664]&m[665]&m[666]&~m[667])|(~m[661]&m[664]&~m[665]&~m[666]&m[667])|(~m[661]&~m[664]&m[665]&~m[666]&m[667])|(m[661]&m[664]&m[665]&~m[666]&m[667])|(~m[661]&m[664]&m[665]&m[666]&m[667]))&UnbiasedRNG[27])|((m[661]&~m[664]&~m[665]&m[666]&~m[667])|(~m[661]&~m[664]&~m[665]&~m[666]&m[667])|(m[661]&~m[664]&~m[665]&~m[666]&m[667])|(m[661]&m[664]&~m[665]&~m[666]&m[667])|(m[661]&~m[664]&m[665]&~m[666]&m[667])|(~m[661]&~m[664]&~m[665]&m[666]&m[667])|(m[661]&~m[664]&~m[665]&m[666]&m[667])|(~m[661]&m[664]&~m[665]&m[666]&m[667])|(m[661]&m[664]&~m[665]&m[666]&m[667])|(~m[661]&~m[664]&m[665]&m[666]&m[667])|(m[661]&~m[664]&m[665]&m[666]&m[667])|(m[661]&m[664]&m[665]&m[666]&m[667]))):InitCond[195];
    m[668] = run?((((m[392]&~m[669]&~m[670]&~m[671]&~m[672])|(~m[392]&~m[669]&~m[670]&m[671]&~m[672])|(m[392]&m[669]&~m[670]&m[671]&~m[672])|(m[392]&~m[669]&m[670]&m[671]&~m[672])|(~m[392]&m[669]&~m[670]&~m[671]&m[672])|(~m[392]&~m[669]&m[670]&~m[671]&m[672])|(m[392]&m[669]&m[670]&~m[671]&m[672])|(~m[392]&m[669]&m[670]&m[671]&m[672]))&UnbiasedRNG[28])|((m[392]&~m[669]&~m[670]&m[671]&~m[672])|(~m[392]&~m[669]&~m[670]&~m[671]&m[672])|(m[392]&~m[669]&~m[670]&~m[671]&m[672])|(m[392]&m[669]&~m[670]&~m[671]&m[672])|(m[392]&~m[669]&m[670]&~m[671]&m[672])|(~m[392]&~m[669]&~m[670]&m[671]&m[672])|(m[392]&~m[669]&~m[670]&m[671]&m[672])|(~m[392]&m[669]&~m[670]&m[671]&m[672])|(m[392]&m[669]&~m[670]&m[671]&m[672])|(~m[392]&~m[669]&m[670]&m[671]&m[672])|(m[392]&~m[669]&m[670]&m[671]&m[672])|(m[392]&m[669]&m[670]&m[671]&m[672]))):InitCond[196];
    m[673] = run?((((m[671]&~m[674]&~m[675]&~m[676]&~m[677])|(~m[671]&~m[674]&~m[675]&m[676]&~m[677])|(m[671]&m[674]&~m[675]&m[676]&~m[677])|(m[671]&~m[674]&m[675]&m[676]&~m[677])|(~m[671]&m[674]&~m[675]&~m[676]&m[677])|(~m[671]&~m[674]&m[675]&~m[676]&m[677])|(m[671]&m[674]&m[675]&~m[676]&m[677])|(~m[671]&m[674]&m[675]&m[676]&m[677]))&UnbiasedRNG[29])|((m[671]&~m[674]&~m[675]&m[676]&~m[677])|(~m[671]&~m[674]&~m[675]&~m[676]&m[677])|(m[671]&~m[674]&~m[675]&~m[676]&m[677])|(m[671]&m[674]&~m[675]&~m[676]&m[677])|(m[671]&~m[674]&m[675]&~m[676]&m[677])|(~m[671]&~m[674]&~m[675]&m[676]&m[677])|(m[671]&~m[674]&~m[675]&m[676]&m[677])|(~m[671]&m[674]&~m[675]&m[676]&m[677])|(m[671]&m[674]&~m[675]&m[676]&m[677])|(~m[671]&~m[674]&m[675]&m[676]&m[677])|(m[671]&~m[674]&m[675]&m[676]&m[677])|(m[671]&m[674]&m[675]&m[676]&m[677]))):InitCond[197];
    m[678] = run?((((m[676]&~m[679]&~m[680]&~m[681]&~m[682])|(~m[676]&~m[679]&~m[680]&m[681]&~m[682])|(m[676]&m[679]&~m[680]&m[681]&~m[682])|(m[676]&~m[679]&m[680]&m[681]&~m[682])|(~m[676]&m[679]&~m[680]&~m[681]&m[682])|(~m[676]&~m[679]&m[680]&~m[681]&m[682])|(m[676]&m[679]&m[680]&~m[681]&m[682])|(~m[676]&m[679]&m[680]&m[681]&m[682]))&UnbiasedRNG[30])|((m[676]&~m[679]&~m[680]&m[681]&~m[682])|(~m[676]&~m[679]&~m[680]&~m[681]&m[682])|(m[676]&~m[679]&~m[680]&~m[681]&m[682])|(m[676]&m[679]&~m[680]&~m[681]&m[682])|(m[676]&~m[679]&m[680]&~m[681]&m[682])|(~m[676]&~m[679]&~m[680]&m[681]&m[682])|(m[676]&~m[679]&~m[680]&m[681]&m[682])|(~m[676]&m[679]&~m[680]&m[681]&m[682])|(m[676]&m[679]&~m[680]&m[681]&m[682])|(~m[676]&~m[679]&m[680]&m[681]&m[682])|(m[676]&~m[679]&m[680]&m[681]&m[682])|(m[676]&m[679]&m[680]&m[681]&m[682]))):InitCond[198];
    m[683] = run?((((m[681]&~m[684]&~m[685]&~m[686]&~m[687])|(~m[681]&~m[684]&~m[685]&m[686]&~m[687])|(m[681]&m[684]&~m[685]&m[686]&~m[687])|(m[681]&~m[684]&m[685]&m[686]&~m[687])|(~m[681]&m[684]&~m[685]&~m[686]&m[687])|(~m[681]&~m[684]&m[685]&~m[686]&m[687])|(m[681]&m[684]&m[685]&~m[686]&m[687])|(~m[681]&m[684]&m[685]&m[686]&m[687]))&UnbiasedRNG[31])|((m[681]&~m[684]&~m[685]&m[686]&~m[687])|(~m[681]&~m[684]&~m[685]&~m[686]&m[687])|(m[681]&~m[684]&~m[685]&~m[686]&m[687])|(m[681]&m[684]&~m[685]&~m[686]&m[687])|(m[681]&~m[684]&m[685]&~m[686]&m[687])|(~m[681]&~m[684]&~m[685]&m[686]&m[687])|(m[681]&~m[684]&~m[685]&m[686]&m[687])|(~m[681]&m[684]&~m[685]&m[686]&m[687])|(m[681]&m[684]&~m[685]&m[686]&m[687])|(~m[681]&~m[684]&m[685]&m[686]&m[687])|(m[681]&~m[684]&m[685]&m[686]&m[687])|(m[681]&m[684]&m[685]&m[686]&m[687]))):InitCond[199];
    m[688] = run?((((m[686]&~m[689]&~m[690]&~m[691]&~m[692])|(~m[686]&~m[689]&~m[690]&m[691]&~m[692])|(m[686]&m[689]&~m[690]&m[691]&~m[692])|(m[686]&~m[689]&m[690]&m[691]&~m[692])|(~m[686]&m[689]&~m[690]&~m[691]&m[692])|(~m[686]&~m[689]&m[690]&~m[691]&m[692])|(m[686]&m[689]&m[690]&~m[691]&m[692])|(~m[686]&m[689]&m[690]&m[691]&m[692]))&UnbiasedRNG[32])|((m[686]&~m[689]&~m[690]&m[691]&~m[692])|(~m[686]&~m[689]&~m[690]&~m[691]&m[692])|(m[686]&~m[689]&~m[690]&~m[691]&m[692])|(m[686]&m[689]&~m[690]&~m[691]&m[692])|(m[686]&~m[689]&m[690]&~m[691]&m[692])|(~m[686]&~m[689]&~m[690]&m[691]&m[692])|(m[686]&~m[689]&~m[690]&m[691]&m[692])|(~m[686]&m[689]&~m[690]&m[691]&m[692])|(m[686]&m[689]&~m[690]&m[691]&m[692])|(~m[686]&~m[689]&m[690]&m[691]&m[692])|(m[686]&~m[689]&m[690]&m[691]&m[692])|(m[686]&m[689]&m[690]&m[691]&m[692]))):InitCond[200];
    m[693] = run?((((m[691]&~m[694]&~m[695]&~m[696]&~m[697])|(~m[691]&~m[694]&~m[695]&m[696]&~m[697])|(m[691]&m[694]&~m[695]&m[696]&~m[697])|(m[691]&~m[694]&m[695]&m[696]&~m[697])|(~m[691]&m[694]&~m[695]&~m[696]&m[697])|(~m[691]&~m[694]&m[695]&~m[696]&m[697])|(m[691]&m[694]&m[695]&~m[696]&m[697])|(~m[691]&m[694]&m[695]&m[696]&m[697]))&UnbiasedRNG[33])|((m[691]&~m[694]&~m[695]&m[696]&~m[697])|(~m[691]&~m[694]&~m[695]&~m[696]&m[697])|(m[691]&~m[694]&~m[695]&~m[696]&m[697])|(m[691]&m[694]&~m[695]&~m[696]&m[697])|(m[691]&~m[694]&m[695]&~m[696]&m[697])|(~m[691]&~m[694]&~m[695]&m[696]&m[697])|(m[691]&~m[694]&~m[695]&m[696]&m[697])|(~m[691]&m[694]&~m[695]&m[696]&m[697])|(m[691]&m[694]&~m[695]&m[696]&m[697])|(~m[691]&~m[694]&m[695]&m[696]&m[697])|(m[691]&~m[694]&m[695]&m[696]&m[697])|(m[691]&m[694]&m[695]&m[696]&m[697]))):InitCond[201];
    m[698] = run?((((m[696]&~m[699]&~m[700]&~m[701]&~m[702])|(~m[696]&~m[699]&~m[700]&m[701]&~m[702])|(m[696]&m[699]&~m[700]&m[701]&~m[702])|(m[696]&~m[699]&m[700]&m[701]&~m[702])|(~m[696]&m[699]&~m[700]&~m[701]&m[702])|(~m[696]&~m[699]&m[700]&~m[701]&m[702])|(m[696]&m[699]&m[700]&~m[701]&m[702])|(~m[696]&m[699]&m[700]&m[701]&m[702]))&UnbiasedRNG[34])|((m[696]&~m[699]&~m[700]&m[701]&~m[702])|(~m[696]&~m[699]&~m[700]&~m[701]&m[702])|(m[696]&~m[699]&~m[700]&~m[701]&m[702])|(m[696]&m[699]&~m[700]&~m[701]&m[702])|(m[696]&~m[699]&m[700]&~m[701]&m[702])|(~m[696]&~m[699]&~m[700]&m[701]&m[702])|(m[696]&~m[699]&~m[700]&m[701]&m[702])|(~m[696]&m[699]&~m[700]&m[701]&m[702])|(m[696]&m[699]&~m[700]&m[701]&m[702])|(~m[696]&~m[699]&m[700]&m[701]&m[702])|(m[696]&~m[699]&m[700]&m[701]&m[702])|(m[696]&m[699]&m[700]&m[701]&m[702]))):InitCond[202];
    m[703] = run?((((m[701]&~m[704]&~m[705]&~m[706]&~m[707])|(~m[701]&~m[704]&~m[705]&m[706]&~m[707])|(m[701]&m[704]&~m[705]&m[706]&~m[707])|(m[701]&~m[704]&m[705]&m[706]&~m[707])|(~m[701]&m[704]&~m[705]&~m[706]&m[707])|(~m[701]&~m[704]&m[705]&~m[706]&m[707])|(m[701]&m[704]&m[705]&~m[706]&m[707])|(~m[701]&m[704]&m[705]&m[706]&m[707]))&UnbiasedRNG[35])|((m[701]&~m[704]&~m[705]&m[706]&~m[707])|(~m[701]&~m[704]&~m[705]&~m[706]&m[707])|(m[701]&~m[704]&~m[705]&~m[706]&m[707])|(m[701]&m[704]&~m[705]&~m[706]&m[707])|(m[701]&~m[704]&m[705]&~m[706]&m[707])|(~m[701]&~m[704]&~m[705]&m[706]&m[707])|(m[701]&~m[704]&~m[705]&m[706]&m[707])|(~m[701]&m[704]&~m[705]&m[706]&m[707])|(m[701]&m[704]&~m[705]&m[706]&m[707])|(~m[701]&~m[704]&m[705]&m[706]&m[707])|(m[701]&~m[704]&m[705]&m[706]&m[707])|(m[701]&m[704]&m[705]&m[706]&m[707]))):InitCond[203];
    m[708] = run?((((m[393]&~m[709]&~m[710]&~m[711]&~m[712])|(~m[393]&~m[709]&~m[710]&m[711]&~m[712])|(m[393]&m[709]&~m[710]&m[711]&~m[712])|(m[393]&~m[709]&m[710]&m[711]&~m[712])|(~m[393]&m[709]&~m[710]&~m[711]&m[712])|(~m[393]&~m[709]&m[710]&~m[711]&m[712])|(m[393]&m[709]&m[710]&~m[711]&m[712])|(~m[393]&m[709]&m[710]&m[711]&m[712]))&UnbiasedRNG[36])|((m[393]&~m[709]&~m[710]&m[711]&~m[712])|(~m[393]&~m[709]&~m[710]&~m[711]&m[712])|(m[393]&~m[709]&~m[710]&~m[711]&m[712])|(m[393]&m[709]&~m[710]&~m[711]&m[712])|(m[393]&~m[709]&m[710]&~m[711]&m[712])|(~m[393]&~m[709]&~m[710]&m[711]&m[712])|(m[393]&~m[709]&~m[710]&m[711]&m[712])|(~m[393]&m[709]&~m[710]&m[711]&m[712])|(m[393]&m[709]&~m[710]&m[711]&m[712])|(~m[393]&~m[709]&m[710]&m[711]&m[712])|(m[393]&~m[709]&m[710]&m[711]&m[712])|(m[393]&m[709]&m[710]&m[711]&m[712]))):InitCond[204];
    m[713] = run?((((m[711]&~m[714]&~m[715]&~m[716]&~m[717])|(~m[711]&~m[714]&~m[715]&m[716]&~m[717])|(m[711]&m[714]&~m[715]&m[716]&~m[717])|(m[711]&~m[714]&m[715]&m[716]&~m[717])|(~m[711]&m[714]&~m[715]&~m[716]&m[717])|(~m[711]&~m[714]&m[715]&~m[716]&m[717])|(m[711]&m[714]&m[715]&~m[716]&m[717])|(~m[711]&m[714]&m[715]&m[716]&m[717]))&UnbiasedRNG[37])|((m[711]&~m[714]&~m[715]&m[716]&~m[717])|(~m[711]&~m[714]&~m[715]&~m[716]&m[717])|(m[711]&~m[714]&~m[715]&~m[716]&m[717])|(m[711]&m[714]&~m[715]&~m[716]&m[717])|(m[711]&~m[714]&m[715]&~m[716]&m[717])|(~m[711]&~m[714]&~m[715]&m[716]&m[717])|(m[711]&~m[714]&~m[715]&m[716]&m[717])|(~m[711]&m[714]&~m[715]&m[716]&m[717])|(m[711]&m[714]&~m[715]&m[716]&m[717])|(~m[711]&~m[714]&m[715]&m[716]&m[717])|(m[711]&~m[714]&m[715]&m[716]&m[717])|(m[711]&m[714]&m[715]&m[716]&m[717]))):InitCond[205];
    m[718] = run?((((m[716]&~m[719]&~m[720]&~m[721]&~m[722])|(~m[716]&~m[719]&~m[720]&m[721]&~m[722])|(m[716]&m[719]&~m[720]&m[721]&~m[722])|(m[716]&~m[719]&m[720]&m[721]&~m[722])|(~m[716]&m[719]&~m[720]&~m[721]&m[722])|(~m[716]&~m[719]&m[720]&~m[721]&m[722])|(m[716]&m[719]&m[720]&~m[721]&m[722])|(~m[716]&m[719]&m[720]&m[721]&m[722]))&UnbiasedRNG[38])|((m[716]&~m[719]&~m[720]&m[721]&~m[722])|(~m[716]&~m[719]&~m[720]&~m[721]&m[722])|(m[716]&~m[719]&~m[720]&~m[721]&m[722])|(m[716]&m[719]&~m[720]&~m[721]&m[722])|(m[716]&~m[719]&m[720]&~m[721]&m[722])|(~m[716]&~m[719]&~m[720]&m[721]&m[722])|(m[716]&~m[719]&~m[720]&m[721]&m[722])|(~m[716]&m[719]&~m[720]&m[721]&m[722])|(m[716]&m[719]&~m[720]&m[721]&m[722])|(~m[716]&~m[719]&m[720]&m[721]&m[722])|(m[716]&~m[719]&m[720]&m[721]&m[722])|(m[716]&m[719]&m[720]&m[721]&m[722]))):InitCond[206];
    m[723] = run?((((m[721]&~m[724]&~m[725]&~m[726]&~m[727])|(~m[721]&~m[724]&~m[725]&m[726]&~m[727])|(m[721]&m[724]&~m[725]&m[726]&~m[727])|(m[721]&~m[724]&m[725]&m[726]&~m[727])|(~m[721]&m[724]&~m[725]&~m[726]&m[727])|(~m[721]&~m[724]&m[725]&~m[726]&m[727])|(m[721]&m[724]&m[725]&~m[726]&m[727])|(~m[721]&m[724]&m[725]&m[726]&m[727]))&UnbiasedRNG[39])|((m[721]&~m[724]&~m[725]&m[726]&~m[727])|(~m[721]&~m[724]&~m[725]&~m[726]&m[727])|(m[721]&~m[724]&~m[725]&~m[726]&m[727])|(m[721]&m[724]&~m[725]&~m[726]&m[727])|(m[721]&~m[724]&m[725]&~m[726]&m[727])|(~m[721]&~m[724]&~m[725]&m[726]&m[727])|(m[721]&~m[724]&~m[725]&m[726]&m[727])|(~m[721]&m[724]&~m[725]&m[726]&m[727])|(m[721]&m[724]&~m[725]&m[726]&m[727])|(~m[721]&~m[724]&m[725]&m[726]&m[727])|(m[721]&~m[724]&m[725]&m[726]&m[727])|(m[721]&m[724]&m[725]&m[726]&m[727]))):InitCond[207];
    m[728] = run?((((m[726]&~m[729]&~m[730]&~m[731]&~m[732])|(~m[726]&~m[729]&~m[730]&m[731]&~m[732])|(m[726]&m[729]&~m[730]&m[731]&~m[732])|(m[726]&~m[729]&m[730]&m[731]&~m[732])|(~m[726]&m[729]&~m[730]&~m[731]&m[732])|(~m[726]&~m[729]&m[730]&~m[731]&m[732])|(m[726]&m[729]&m[730]&~m[731]&m[732])|(~m[726]&m[729]&m[730]&m[731]&m[732]))&UnbiasedRNG[40])|((m[726]&~m[729]&~m[730]&m[731]&~m[732])|(~m[726]&~m[729]&~m[730]&~m[731]&m[732])|(m[726]&~m[729]&~m[730]&~m[731]&m[732])|(m[726]&m[729]&~m[730]&~m[731]&m[732])|(m[726]&~m[729]&m[730]&~m[731]&m[732])|(~m[726]&~m[729]&~m[730]&m[731]&m[732])|(m[726]&~m[729]&~m[730]&m[731]&m[732])|(~m[726]&m[729]&~m[730]&m[731]&m[732])|(m[726]&m[729]&~m[730]&m[731]&m[732])|(~m[726]&~m[729]&m[730]&m[731]&m[732])|(m[726]&~m[729]&m[730]&m[731]&m[732])|(m[726]&m[729]&m[730]&m[731]&m[732]))):InitCond[208];
    m[733] = run?((((m[731]&~m[734]&~m[735]&~m[736]&~m[737])|(~m[731]&~m[734]&~m[735]&m[736]&~m[737])|(m[731]&m[734]&~m[735]&m[736]&~m[737])|(m[731]&~m[734]&m[735]&m[736]&~m[737])|(~m[731]&m[734]&~m[735]&~m[736]&m[737])|(~m[731]&~m[734]&m[735]&~m[736]&m[737])|(m[731]&m[734]&m[735]&~m[736]&m[737])|(~m[731]&m[734]&m[735]&m[736]&m[737]))&UnbiasedRNG[41])|((m[731]&~m[734]&~m[735]&m[736]&~m[737])|(~m[731]&~m[734]&~m[735]&~m[736]&m[737])|(m[731]&~m[734]&~m[735]&~m[736]&m[737])|(m[731]&m[734]&~m[735]&~m[736]&m[737])|(m[731]&~m[734]&m[735]&~m[736]&m[737])|(~m[731]&~m[734]&~m[735]&m[736]&m[737])|(m[731]&~m[734]&~m[735]&m[736]&m[737])|(~m[731]&m[734]&~m[735]&m[736]&m[737])|(m[731]&m[734]&~m[735]&m[736]&m[737])|(~m[731]&~m[734]&m[735]&m[736]&m[737])|(m[731]&~m[734]&m[735]&m[736]&m[737])|(m[731]&m[734]&m[735]&m[736]&m[737]))):InitCond[209];
    m[738] = run?((((m[736]&~m[739]&~m[740]&~m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&m[741]&~m[742])|(m[736]&m[739]&~m[740]&m[741]&~m[742])|(m[736]&~m[739]&m[740]&m[741]&~m[742])|(~m[736]&m[739]&~m[740]&~m[741]&m[742])|(~m[736]&~m[739]&m[740]&~m[741]&m[742])|(m[736]&m[739]&m[740]&~m[741]&m[742])|(~m[736]&m[739]&m[740]&m[741]&m[742]))&UnbiasedRNG[42])|((m[736]&~m[739]&~m[740]&m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&m[740]&~m[741]&m[742])|(~m[736]&~m[739]&~m[740]&m[741]&m[742])|(m[736]&~m[739]&~m[740]&m[741]&m[742])|(~m[736]&m[739]&~m[740]&m[741]&m[742])|(m[736]&m[739]&~m[740]&m[741]&m[742])|(~m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&m[739]&m[740]&m[741]&m[742]))):InitCond[210];
    m[743] = run?((((m[741]&~m[744]&~m[745]&~m[746]&~m[747])|(~m[741]&~m[744]&~m[745]&m[746]&~m[747])|(m[741]&m[744]&~m[745]&m[746]&~m[747])|(m[741]&~m[744]&m[745]&m[746]&~m[747])|(~m[741]&m[744]&~m[745]&~m[746]&m[747])|(~m[741]&~m[744]&m[745]&~m[746]&m[747])|(m[741]&m[744]&m[745]&~m[746]&m[747])|(~m[741]&m[744]&m[745]&m[746]&m[747]))&UnbiasedRNG[43])|((m[741]&~m[744]&~m[745]&m[746]&~m[747])|(~m[741]&~m[744]&~m[745]&~m[746]&m[747])|(m[741]&~m[744]&~m[745]&~m[746]&m[747])|(m[741]&m[744]&~m[745]&~m[746]&m[747])|(m[741]&~m[744]&m[745]&~m[746]&m[747])|(~m[741]&~m[744]&~m[745]&m[746]&m[747])|(m[741]&~m[744]&~m[745]&m[746]&m[747])|(~m[741]&m[744]&~m[745]&m[746]&m[747])|(m[741]&m[744]&~m[745]&m[746]&m[747])|(~m[741]&~m[744]&m[745]&m[746]&m[747])|(m[741]&~m[744]&m[745]&m[746]&m[747])|(m[741]&m[744]&m[745]&m[746]&m[747]))):InitCond[211];
    m[748] = run?((((m[746]&~m[749]&~m[750]&~m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&m[751]&~m[752])|(m[746]&m[749]&~m[750]&m[751]&~m[752])|(m[746]&~m[749]&m[750]&m[751]&~m[752])|(~m[746]&m[749]&~m[750]&~m[751]&m[752])|(~m[746]&~m[749]&m[750]&~m[751]&m[752])|(m[746]&m[749]&m[750]&~m[751]&m[752])|(~m[746]&m[749]&m[750]&m[751]&m[752]))&UnbiasedRNG[44])|((m[746]&~m[749]&~m[750]&m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&m[750]&~m[751]&m[752])|(~m[746]&~m[749]&~m[750]&m[751]&m[752])|(m[746]&~m[749]&~m[750]&m[751]&m[752])|(~m[746]&m[749]&~m[750]&m[751]&m[752])|(m[746]&m[749]&~m[750]&m[751]&m[752])|(~m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&m[749]&m[750]&m[751]&m[752]))):InitCond[212];
    m[753] = run?((((m[394]&~m[754]&~m[755]&~m[756]&~m[757])|(~m[394]&~m[754]&~m[755]&m[756]&~m[757])|(m[394]&m[754]&~m[755]&m[756]&~m[757])|(m[394]&~m[754]&m[755]&m[756]&~m[757])|(~m[394]&m[754]&~m[755]&~m[756]&m[757])|(~m[394]&~m[754]&m[755]&~m[756]&m[757])|(m[394]&m[754]&m[755]&~m[756]&m[757])|(~m[394]&m[754]&m[755]&m[756]&m[757]))&UnbiasedRNG[45])|((m[394]&~m[754]&~m[755]&m[756]&~m[757])|(~m[394]&~m[754]&~m[755]&~m[756]&m[757])|(m[394]&~m[754]&~m[755]&~m[756]&m[757])|(m[394]&m[754]&~m[755]&~m[756]&m[757])|(m[394]&~m[754]&m[755]&~m[756]&m[757])|(~m[394]&~m[754]&~m[755]&m[756]&m[757])|(m[394]&~m[754]&~m[755]&m[756]&m[757])|(~m[394]&m[754]&~m[755]&m[756]&m[757])|(m[394]&m[754]&~m[755]&m[756]&m[757])|(~m[394]&~m[754]&m[755]&m[756]&m[757])|(m[394]&~m[754]&m[755]&m[756]&m[757])|(m[394]&m[754]&m[755]&m[756]&m[757]))):InitCond[213];
    m[758] = run?((((m[756]&~m[759]&~m[760]&~m[761]&~m[762])|(~m[756]&~m[759]&~m[760]&m[761]&~m[762])|(m[756]&m[759]&~m[760]&m[761]&~m[762])|(m[756]&~m[759]&m[760]&m[761]&~m[762])|(~m[756]&m[759]&~m[760]&~m[761]&m[762])|(~m[756]&~m[759]&m[760]&~m[761]&m[762])|(m[756]&m[759]&m[760]&~m[761]&m[762])|(~m[756]&m[759]&m[760]&m[761]&m[762]))&UnbiasedRNG[46])|((m[756]&~m[759]&~m[760]&m[761]&~m[762])|(~m[756]&~m[759]&~m[760]&~m[761]&m[762])|(m[756]&~m[759]&~m[760]&~m[761]&m[762])|(m[756]&m[759]&~m[760]&~m[761]&m[762])|(m[756]&~m[759]&m[760]&~m[761]&m[762])|(~m[756]&~m[759]&~m[760]&m[761]&m[762])|(m[756]&~m[759]&~m[760]&m[761]&m[762])|(~m[756]&m[759]&~m[760]&m[761]&m[762])|(m[756]&m[759]&~m[760]&m[761]&m[762])|(~m[756]&~m[759]&m[760]&m[761]&m[762])|(m[756]&~m[759]&m[760]&m[761]&m[762])|(m[756]&m[759]&m[760]&m[761]&m[762]))):InitCond[214];
    m[763] = run?((((m[761]&~m[764]&~m[765]&~m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&m[766]&~m[767])|(m[761]&m[764]&~m[765]&m[766]&~m[767])|(m[761]&~m[764]&m[765]&m[766]&~m[767])|(~m[761]&m[764]&~m[765]&~m[766]&m[767])|(~m[761]&~m[764]&m[765]&~m[766]&m[767])|(m[761]&m[764]&m[765]&~m[766]&m[767])|(~m[761]&m[764]&m[765]&m[766]&m[767]))&UnbiasedRNG[47])|((m[761]&~m[764]&~m[765]&m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&m[765]&~m[766]&m[767])|(~m[761]&~m[764]&~m[765]&m[766]&m[767])|(m[761]&~m[764]&~m[765]&m[766]&m[767])|(~m[761]&m[764]&~m[765]&m[766]&m[767])|(m[761]&m[764]&~m[765]&m[766]&m[767])|(~m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&m[764]&m[765]&m[766]&m[767]))):InitCond[215];
    m[768] = run?((((m[766]&~m[769]&~m[770]&~m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&m[771]&~m[772])|(m[766]&m[769]&~m[770]&m[771]&~m[772])|(m[766]&~m[769]&m[770]&m[771]&~m[772])|(~m[766]&m[769]&~m[770]&~m[771]&m[772])|(~m[766]&~m[769]&m[770]&~m[771]&m[772])|(m[766]&m[769]&m[770]&~m[771]&m[772])|(~m[766]&m[769]&m[770]&m[771]&m[772]))&UnbiasedRNG[48])|((m[766]&~m[769]&~m[770]&m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&m[770]&~m[771]&m[772])|(~m[766]&~m[769]&~m[770]&m[771]&m[772])|(m[766]&~m[769]&~m[770]&m[771]&m[772])|(~m[766]&m[769]&~m[770]&m[771]&m[772])|(m[766]&m[769]&~m[770]&m[771]&m[772])|(~m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&m[769]&m[770]&m[771]&m[772]))):InitCond[216];
    m[773] = run?((((m[771]&~m[774]&~m[775]&~m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&m[776]&~m[777])|(m[771]&m[774]&~m[775]&m[776]&~m[777])|(m[771]&~m[774]&m[775]&m[776]&~m[777])|(~m[771]&m[774]&~m[775]&~m[776]&m[777])|(~m[771]&~m[774]&m[775]&~m[776]&m[777])|(m[771]&m[774]&m[775]&~m[776]&m[777])|(~m[771]&m[774]&m[775]&m[776]&m[777]))&UnbiasedRNG[49])|((m[771]&~m[774]&~m[775]&m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&m[775]&~m[776]&m[777])|(~m[771]&~m[774]&~m[775]&m[776]&m[777])|(m[771]&~m[774]&~m[775]&m[776]&m[777])|(~m[771]&m[774]&~m[775]&m[776]&m[777])|(m[771]&m[774]&~m[775]&m[776]&m[777])|(~m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&m[774]&m[775]&m[776]&m[777]))):InitCond[217];
    m[778] = run?((((m[776]&~m[779]&~m[780]&~m[781]&~m[782])|(~m[776]&~m[779]&~m[780]&m[781]&~m[782])|(m[776]&m[779]&~m[780]&m[781]&~m[782])|(m[776]&~m[779]&m[780]&m[781]&~m[782])|(~m[776]&m[779]&~m[780]&~m[781]&m[782])|(~m[776]&~m[779]&m[780]&~m[781]&m[782])|(m[776]&m[779]&m[780]&~m[781]&m[782])|(~m[776]&m[779]&m[780]&m[781]&m[782]))&UnbiasedRNG[50])|((m[776]&~m[779]&~m[780]&m[781]&~m[782])|(~m[776]&~m[779]&~m[780]&~m[781]&m[782])|(m[776]&~m[779]&~m[780]&~m[781]&m[782])|(m[776]&m[779]&~m[780]&~m[781]&m[782])|(m[776]&~m[779]&m[780]&~m[781]&m[782])|(~m[776]&~m[779]&~m[780]&m[781]&m[782])|(m[776]&~m[779]&~m[780]&m[781]&m[782])|(~m[776]&m[779]&~m[780]&m[781]&m[782])|(m[776]&m[779]&~m[780]&m[781]&m[782])|(~m[776]&~m[779]&m[780]&m[781]&m[782])|(m[776]&~m[779]&m[780]&m[781]&m[782])|(m[776]&m[779]&m[780]&m[781]&m[782]))):InitCond[218];
    m[783] = run?((((m[781]&~m[784]&~m[785]&~m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&m[786]&~m[787])|(m[781]&m[784]&~m[785]&m[786]&~m[787])|(m[781]&~m[784]&m[785]&m[786]&~m[787])|(~m[781]&m[784]&~m[785]&~m[786]&m[787])|(~m[781]&~m[784]&m[785]&~m[786]&m[787])|(m[781]&m[784]&m[785]&~m[786]&m[787])|(~m[781]&m[784]&m[785]&m[786]&m[787]))&UnbiasedRNG[51])|((m[781]&~m[784]&~m[785]&m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&m[785]&~m[786]&m[787])|(~m[781]&~m[784]&~m[785]&m[786]&m[787])|(m[781]&~m[784]&~m[785]&m[786]&m[787])|(~m[781]&m[784]&~m[785]&m[786]&m[787])|(m[781]&m[784]&~m[785]&m[786]&m[787])|(~m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&m[784]&m[785]&m[786]&m[787]))):InitCond[219];
    m[788] = run?((((m[786]&~m[789]&~m[790]&~m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&m[791]&~m[792])|(m[786]&m[789]&~m[790]&m[791]&~m[792])|(m[786]&~m[789]&m[790]&m[791]&~m[792])|(~m[786]&m[789]&~m[790]&~m[791]&m[792])|(~m[786]&~m[789]&m[790]&~m[791]&m[792])|(m[786]&m[789]&m[790]&~m[791]&m[792])|(~m[786]&m[789]&m[790]&m[791]&m[792]))&UnbiasedRNG[52])|((m[786]&~m[789]&~m[790]&m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&m[790]&~m[791]&m[792])|(~m[786]&~m[789]&~m[790]&m[791]&m[792])|(m[786]&~m[789]&~m[790]&m[791]&m[792])|(~m[786]&m[789]&~m[790]&m[791]&m[792])|(m[786]&m[789]&~m[790]&m[791]&m[792])|(~m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&m[789]&m[790]&m[791]&m[792]))):InitCond[220];
    m[793] = run?((((m[791]&~m[794]&~m[795]&~m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&m[796]&~m[797])|(m[791]&m[794]&~m[795]&m[796]&~m[797])|(m[791]&~m[794]&m[795]&m[796]&~m[797])|(~m[791]&m[794]&~m[795]&~m[796]&m[797])|(~m[791]&~m[794]&m[795]&~m[796]&m[797])|(m[791]&m[794]&m[795]&~m[796]&m[797])|(~m[791]&m[794]&m[795]&m[796]&m[797]))&UnbiasedRNG[53])|((m[791]&~m[794]&~m[795]&m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&m[795]&~m[796]&m[797])|(~m[791]&~m[794]&~m[795]&m[796]&m[797])|(m[791]&~m[794]&~m[795]&m[796]&m[797])|(~m[791]&m[794]&~m[795]&m[796]&m[797])|(m[791]&m[794]&~m[795]&m[796]&m[797])|(~m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&m[794]&m[795]&m[796]&m[797]))):InitCond[221];
    m[798] = run?((((m[796]&~m[799]&~m[800]&~m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&m[801]&~m[802])|(m[796]&m[799]&~m[800]&m[801]&~m[802])|(m[796]&~m[799]&m[800]&m[801]&~m[802])|(~m[796]&m[799]&~m[800]&~m[801]&m[802])|(~m[796]&~m[799]&m[800]&~m[801]&m[802])|(m[796]&m[799]&m[800]&~m[801]&m[802])|(~m[796]&m[799]&m[800]&m[801]&m[802]))&UnbiasedRNG[54])|((m[796]&~m[799]&~m[800]&m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&m[800]&~m[801]&m[802])|(~m[796]&~m[799]&~m[800]&m[801]&m[802])|(m[796]&~m[799]&~m[800]&m[801]&m[802])|(~m[796]&m[799]&~m[800]&m[801]&m[802])|(m[796]&m[799]&~m[800]&m[801]&m[802])|(~m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&m[799]&m[800]&m[801]&m[802]))):InitCond[222];
    m[803] = run?((((m[395]&~m[804]&~m[805]&~m[806]&~m[807])|(~m[395]&~m[804]&~m[805]&m[806]&~m[807])|(m[395]&m[804]&~m[805]&m[806]&~m[807])|(m[395]&~m[804]&m[805]&m[806]&~m[807])|(~m[395]&m[804]&~m[805]&~m[806]&m[807])|(~m[395]&~m[804]&m[805]&~m[806]&m[807])|(m[395]&m[804]&m[805]&~m[806]&m[807])|(~m[395]&m[804]&m[805]&m[806]&m[807]))&UnbiasedRNG[55])|((m[395]&~m[804]&~m[805]&m[806]&~m[807])|(~m[395]&~m[804]&~m[805]&~m[806]&m[807])|(m[395]&~m[804]&~m[805]&~m[806]&m[807])|(m[395]&m[804]&~m[805]&~m[806]&m[807])|(m[395]&~m[804]&m[805]&~m[806]&m[807])|(~m[395]&~m[804]&~m[805]&m[806]&m[807])|(m[395]&~m[804]&~m[805]&m[806]&m[807])|(~m[395]&m[804]&~m[805]&m[806]&m[807])|(m[395]&m[804]&~m[805]&m[806]&m[807])|(~m[395]&~m[804]&m[805]&m[806]&m[807])|(m[395]&~m[804]&m[805]&m[806]&m[807])|(m[395]&m[804]&m[805]&m[806]&m[807]))):InitCond[223];
    m[808] = run?((((m[806]&~m[809]&~m[810]&~m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&m[811]&~m[812])|(m[806]&m[809]&~m[810]&m[811]&~m[812])|(m[806]&~m[809]&m[810]&m[811]&~m[812])|(~m[806]&m[809]&~m[810]&~m[811]&m[812])|(~m[806]&~m[809]&m[810]&~m[811]&m[812])|(m[806]&m[809]&m[810]&~m[811]&m[812])|(~m[806]&m[809]&m[810]&m[811]&m[812]))&UnbiasedRNG[56])|((m[806]&~m[809]&~m[810]&m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&m[810]&~m[811]&m[812])|(~m[806]&~m[809]&~m[810]&m[811]&m[812])|(m[806]&~m[809]&~m[810]&m[811]&m[812])|(~m[806]&m[809]&~m[810]&m[811]&m[812])|(m[806]&m[809]&~m[810]&m[811]&m[812])|(~m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&m[809]&m[810]&m[811]&m[812]))):InitCond[224];
    m[813] = run?((((m[811]&~m[814]&~m[815]&~m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&m[816]&~m[817])|(m[811]&m[814]&~m[815]&m[816]&~m[817])|(m[811]&~m[814]&m[815]&m[816]&~m[817])|(~m[811]&m[814]&~m[815]&~m[816]&m[817])|(~m[811]&~m[814]&m[815]&~m[816]&m[817])|(m[811]&m[814]&m[815]&~m[816]&m[817])|(~m[811]&m[814]&m[815]&m[816]&m[817]))&UnbiasedRNG[57])|((m[811]&~m[814]&~m[815]&m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&m[815]&~m[816]&m[817])|(~m[811]&~m[814]&~m[815]&m[816]&m[817])|(m[811]&~m[814]&~m[815]&m[816]&m[817])|(~m[811]&m[814]&~m[815]&m[816]&m[817])|(m[811]&m[814]&~m[815]&m[816]&m[817])|(~m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&m[814]&m[815]&m[816]&m[817]))):InitCond[225];
    m[818] = run?((((m[816]&~m[819]&~m[820]&~m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&m[821]&~m[822])|(m[816]&m[819]&~m[820]&m[821]&~m[822])|(m[816]&~m[819]&m[820]&m[821]&~m[822])|(~m[816]&m[819]&~m[820]&~m[821]&m[822])|(~m[816]&~m[819]&m[820]&~m[821]&m[822])|(m[816]&m[819]&m[820]&~m[821]&m[822])|(~m[816]&m[819]&m[820]&m[821]&m[822]))&UnbiasedRNG[58])|((m[816]&~m[819]&~m[820]&m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&m[820]&~m[821]&m[822])|(~m[816]&~m[819]&~m[820]&m[821]&m[822])|(m[816]&~m[819]&~m[820]&m[821]&m[822])|(~m[816]&m[819]&~m[820]&m[821]&m[822])|(m[816]&m[819]&~m[820]&m[821]&m[822])|(~m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&m[819]&m[820]&m[821]&m[822]))):InitCond[226];
    m[823] = run?((((m[821]&~m[824]&~m[825]&~m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&m[826]&~m[827])|(m[821]&m[824]&~m[825]&m[826]&~m[827])|(m[821]&~m[824]&m[825]&m[826]&~m[827])|(~m[821]&m[824]&~m[825]&~m[826]&m[827])|(~m[821]&~m[824]&m[825]&~m[826]&m[827])|(m[821]&m[824]&m[825]&~m[826]&m[827])|(~m[821]&m[824]&m[825]&m[826]&m[827]))&UnbiasedRNG[59])|((m[821]&~m[824]&~m[825]&m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&m[825]&~m[826]&m[827])|(~m[821]&~m[824]&~m[825]&m[826]&m[827])|(m[821]&~m[824]&~m[825]&m[826]&m[827])|(~m[821]&m[824]&~m[825]&m[826]&m[827])|(m[821]&m[824]&~m[825]&m[826]&m[827])|(~m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&m[824]&m[825]&m[826]&m[827]))):InitCond[227];
    m[828] = run?((((m[826]&~m[829]&~m[830]&~m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&m[831]&~m[832])|(m[826]&m[829]&~m[830]&m[831]&~m[832])|(m[826]&~m[829]&m[830]&m[831]&~m[832])|(~m[826]&m[829]&~m[830]&~m[831]&m[832])|(~m[826]&~m[829]&m[830]&~m[831]&m[832])|(m[826]&m[829]&m[830]&~m[831]&m[832])|(~m[826]&m[829]&m[830]&m[831]&m[832]))&UnbiasedRNG[60])|((m[826]&~m[829]&~m[830]&m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&m[830]&~m[831]&m[832])|(~m[826]&~m[829]&~m[830]&m[831]&m[832])|(m[826]&~m[829]&~m[830]&m[831]&m[832])|(~m[826]&m[829]&~m[830]&m[831]&m[832])|(m[826]&m[829]&~m[830]&m[831]&m[832])|(~m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&m[829]&m[830]&m[831]&m[832]))):InitCond[228];
    m[833] = run?((((m[831]&~m[834]&~m[835]&~m[836]&~m[837])|(~m[831]&~m[834]&~m[835]&m[836]&~m[837])|(m[831]&m[834]&~m[835]&m[836]&~m[837])|(m[831]&~m[834]&m[835]&m[836]&~m[837])|(~m[831]&m[834]&~m[835]&~m[836]&m[837])|(~m[831]&~m[834]&m[835]&~m[836]&m[837])|(m[831]&m[834]&m[835]&~m[836]&m[837])|(~m[831]&m[834]&m[835]&m[836]&m[837]))&UnbiasedRNG[61])|((m[831]&~m[834]&~m[835]&m[836]&~m[837])|(~m[831]&~m[834]&~m[835]&~m[836]&m[837])|(m[831]&~m[834]&~m[835]&~m[836]&m[837])|(m[831]&m[834]&~m[835]&~m[836]&m[837])|(m[831]&~m[834]&m[835]&~m[836]&m[837])|(~m[831]&~m[834]&~m[835]&m[836]&m[837])|(m[831]&~m[834]&~m[835]&m[836]&m[837])|(~m[831]&m[834]&~m[835]&m[836]&m[837])|(m[831]&m[834]&~m[835]&m[836]&m[837])|(~m[831]&~m[834]&m[835]&m[836]&m[837])|(m[831]&~m[834]&m[835]&m[836]&m[837])|(m[831]&m[834]&m[835]&m[836]&m[837]))):InitCond[229];
    m[838] = run?((((m[836]&~m[839]&~m[840]&~m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&m[841]&~m[842])|(m[836]&m[839]&~m[840]&m[841]&~m[842])|(m[836]&~m[839]&m[840]&m[841]&~m[842])|(~m[836]&m[839]&~m[840]&~m[841]&m[842])|(~m[836]&~m[839]&m[840]&~m[841]&m[842])|(m[836]&m[839]&m[840]&~m[841]&m[842])|(~m[836]&m[839]&m[840]&m[841]&m[842]))&UnbiasedRNG[62])|((m[836]&~m[839]&~m[840]&m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&m[840]&~m[841]&m[842])|(~m[836]&~m[839]&~m[840]&m[841]&m[842])|(m[836]&~m[839]&~m[840]&m[841]&m[842])|(~m[836]&m[839]&~m[840]&m[841]&m[842])|(m[836]&m[839]&~m[840]&m[841]&m[842])|(~m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&m[839]&m[840]&m[841]&m[842]))):InitCond[230];
    m[843] = run?((((m[841]&~m[844]&~m[845]&~m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&m[846]&~m[847])|(m[841]&m[844]&~m[845]&m[846]&~m[847])|(m[841]&~m[844]&m[845]&m[846]&~m[847])|(~m[841]&m[844]&~m[845]&~m[846]&m[847])|(~m[841]&~m[844]&m[845]&~m[846]&m[847])|(m[841]&m[844]&m[845]&~m[846]&m[847])|(~m[841]&m[844]&m[845]&m[846]&m[847]))&UnbiasedRNG[63])|((m[841]&~m[844]&~m[845]&m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&m[845]&~m[846]&m[847])|(~m[841]&~m[844]&~m[845]&m[846]&m[847])|(m[841]&~m[844]&~m[845]&m[846]&m[847])|(~m[841]&m[844]&~m[845]&m[846]&m[847])|(m[841]&m[844]&~m[845]&m[846]&m[847])|(~m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&m[844]&m[845]&m[846]&m[847]))):InitCond[231];
    m[848] = run?((((m[846]&~m[849]&~m[850]&~m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&m[851]&~m[852])|(m[846]&m[849]&~m[850]&m[851]&~m[852])|(m[846]&~m[849]&m[850]&m[851]&~m[852])|(~m[846]&m[849]&~m[850]&~m[851]&m[852])|(~m[846]&~m[849]&m[850]&~m[851]&m[852])|(m[846]&m[849]&m[850]&~m[851]&m[852])|(~m[846]&m[849]&m[850]&m[851]&m[852]))&UnbiasedRNG[64])|((m[846]&~m[849]&~m[850]&m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&m[850]&~m[851]&m[852])|(~m[846]&~m[849]&~m[850]&m[851]&m[852])|(m[846]&~m[849]&~m[850]&m[851]&m[852])|(~m[846]&m[849]&~m[850]&m[851]&m[852])|(m[846]&m[849]&~m[850]&m[851]&m[852])|(~m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&m[849]&m[850]&m[851]&m[852]))):InitCond[232];
    m[853] = run?((((m[851]&~m[854]&~m[855]&~m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&m[856]&~m[857])|(m[851]&m[854]&~m[855]&m[856]&~m[857])|(m[851]&~m[854]&m[855]&m[856]&~m[857])|(~m[851]&m[854]&~m[855]&~m[856]&m[857])|(~m[851]&~m[854]&m[855]&~m[856]&m[857])|(m[851]&m[854]&m[855]&~m[856]&m[857])|(~m[851]&m[854]&m[855]&m[856]&m[857]))&UnbiasedRNG[65])|((m[851]&~m[854]&~m[855]&m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&m[855]&~m[856]&m[857])|(~m[851]&~m[854]&~m[855]&m[856]&m[857])|(m[851]&~m[854]&~m[855]&m[856]&m[857])|(~m[851]&m[854]&~m[855]&m[856]&m[857])|(m[851]&m[854]&~m[855]&m[856]&m[857])|(~m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&m[854]&m[855]&m[856]&m[857]))):InitCond[233];
    m[863] = run?((((m[861]&~m[864]&~m[865]&~m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&m[866]&~m[867])|(m[861]&m[864]&~m[865]&m[866]&~m[867])|(m[861]&~m[864]&m[865]&m[866]&~m[867])|(~m[861]&m[864]&~m[865]&~m[866]&m[867])|(~m[861]&~m[864]&m[865]&~m[866]&m[867])|(m[861]&m[864]&m[865]&~m[866]&m[867])|(~m[861]&m[864]&m[865]&m[866]&m[867]))&UnbiasedRNG[66])|((m[861]&~m[864]&~m[865]&m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&m[865]&~m[866]&m[867])|(~m[861]&~m[864]&~m[865]&m[866]&m[867])|(m[861]&~m[864]&~m[865]&m[866]&m[867])|(~m[861]&m[864]&~m[865]&m[866]&m[867])|(m[861]&m[864]&~m[865]&m[866]&m[867])|(~m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&m[864]&m[865]&m[866]&m[867]))):InitCond[234];
    m[868] = run?((((m[866]&~m[869]&~m[870]&~m[871]&~m[872])|(~m[866]&~m[869]&~m[870]&m[871]&~m[872])|(m[866]&m[869]&~m[870]&m[871]&~m[872])|(m[866]&~m[869]&m[870]&m[871]&~m[872])|(~m[866]&m[869]&~m[870]&~m[871]&m[872])|(~m[866]&~m[869]&m[870]&~m[871]&m[872])|(m[866]&m[869]&m[870]&~m[871]&m[872])|(~m[866]&m[869]&m[870]&m[871]&m[872]))&UnbiasedRNG[67])|((m[866]&~m[869]&~m[870]&m[871]&~m[872])|(~m[866]&~m[869]&~m[870]&~m[871]&m[872])|(m[866]&~m[869]&~m[870]&~m[871]&m[872])|(m[866]&m[869]&~m[870]&~m[871]&m[872])|(m[866]&~m[869]&m[870]&~m[871]&m[872])|(~m[866]&~m[869]&~m[870]&m[871]&m[872])|(m[866]&~m[869]&~m[870]&m[871]&m[872])|(~m[866]&m[869]&~m[870]&m[871]&m[872])|(m[866]&m[869]&~m[870]&m[871]&m[872])|(~m[866]&~m[869]&m[870]&m[871]&m[872])|(m[866]&~m[869]&m[870]&m[871]&m[872])|(m[866]&m[869]&m[870]&m[871]&m[872]))):InitCond[235];
    m[873] = run?((((m[871]&~m[874]&~m[875]&~m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&m[876]&~m[877])|(m[871]&m[874]&~m[875]&m[876]&~m[877])|(m[871]&~m[874]&m[875]&m[876]&~m[877])|(~m[871]&m[874]&~m[875]&~m[876]&m[877])|(~m[871]&~m[874]&m[875]&~m[876]&m[877])|(m[871]&m[874]&m[875]&~m[876]&m[877])|(~m[871]&m[874]&m[875]&m[876]&m[877]))&UnbiasedRNG[68])|((m[871]&~m[874]&~m[875]&m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&m[875]&~m[876]&m[877])|(~m[871]&~m[874]&~m[875]&m[876]&m[877])|(m[871]&~m[874]&~m[875]&m[876]&m[877])|(~m[871]&m[874]&~m[875]&m[876]&m[877])|(m[871]&m[874]&~m[875]&m[876]&m[877])|(~m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&m[874]&m[875]&m[876]&m[877]))):InitCond[236];
    m[878] = run?((((m[876]&~m[879]&~m[880]&~m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&m[881]&~m[882])|(m[876]&m[879]&~m[880]&m[881]&~m[882])|(m[876]&~m[879]&m[880]&m[881]&~m[882])|(~m[876]&m[879]&~m[880]&~m[881]&m[882])|(~m[876]&~m[879]&m[880]&~m[881]&m[882])|(m[876]&m[879]&m[880]&~m[881]&m[882])|(~m[876]&m[879]&m[880]&m[881]&m[882]))&UnbiasedRNG[69])|((m[876]&~m[879]&~m[880]&m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&m[880]&~m[881]&m[882])|(~m[876]&~m[879]&~m[880]&m[881]&m[882])|(m[876]&~m[879]&~m[880]&m[881]&m[882])|(~m[876]&m[879]&~m[880]&m[881]&m[882])|(m[876]&m[879]&~m[880]&m[881]&m[882])|(~m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&m[879]&m[880]&m[881]&m[882]))):InitCond[237];
    m[883] = run?((((m[881]&~m[884]&~m[885]&~m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&m[886]&~m[887])|(m[881]&m[884]&~m[885]&m[886]&~m[887])|(m[881]&~m[884]&m[885]&m[886]&~m[887])|(~m[881]&m[884]&~m[885]&~m[886]&m[887])|(~m[881]&~m[884]&m[885]&~m[886]&m[887])|(m[881]&m[884]&m[885]&~m[886]&m[887])|(~m[881]&m[884]&m[885]&m[886]&m[887]))&UnbiasedRNG[70])|((m[881]&~m[884]&~m[885]&m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&m[885]&~m[886]&m[887])|(~m[881]&~m[884]&~m[885]&m[886]&m[887])|(m[881]&~m[884]&~m[885]&m[886]&m[887])|(~m[881]&m[884]&~m[885]&m[886]&m[887])|(m[881]&m[884]&~m[885]&m[886]&m[887])|(~m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&m[884]&m[885]&m[886]&m[887]))):InitCond[238];
    m[888] = run?((((m[886]&~m[889]&~m[890]&~m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&m[891]&~m[892])|(m[886]&m[889]&~m[890]&m[891]&~m[892])|(m[886]&~m[889]&m[890]&m[891]&~m[892])|(~m[886]&m[889]&~m[890]&~m[891]&m[892])|(~m[886]&~m[889]&m[890]&~m[891]&m[892])|(m[886]&m[889]&m[890]&~m[891]&m[892])|(~m[886]&m[889]&m[890]&m[891]&m[892]))&UnbiasedRNG[71])|((m[886]&~m[889]&~m[890]&m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&m[890]&~m[891]&m[892])|(~m[886]&~m[889]&~m[890]&m[891]&m[892])|(m[886]&~m[889]&~m[890]&m[891]&m[892])|(~m[886]&m[889]&~m[890]&m[891]&m[892])|(m[886]&m[889]&~m[890]&m[891]&m[892])|(~m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&m[889]&m[890]&m[891]&m[892]))):InitCond[239];
    m[893] = run?((((m[891]&~m[894]&~m[895]&~m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&m[896]&~m[897])|(m[891]&m[894]&~m[895]&m[896]&~m[897])|(m[891]&~m[894]&m[895]&m[896]&~m[897])|(~m[891]&m[894]&~m[895]&~m[896]&m[897])|(~m[891]&~m[894]&m[895]&~m[896]&m[897])|(m[891]&m[894]&m[895]&~m[896]&m[897])|(~m[891]&m[894]&m[895]&m[896]&m[897]))&UnbiasedRNG[72])|((m[891]&~m[894]&~m[895]&m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&m[895]&~m[896]&m[897])|(~m[891]&~m[894]&~m[895]&m[896]&m[897])|(m[891]&~m[894]&~m[895]&m[896]&m[897])|(~m[891]&m[894]&~m[895]&m[896]&m[897])|(m[891]&m[894]&~m[895]&m[896]&m[897])|(~m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&m[894]&m[895]&m[896]&m[897]))):InitCond[240];
    m[898] = run?((((m[896]&~m[899]&~m[900]&~m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&m[901]&~m[902])|(m[896]&m[899]&~m[900]&m[901]&~m[902])|(m[896]&~m[899]&m[900]&m[901]&~m[902])|(~m[896]&m[899]&~m[900]&~m[901]&m[902])|(~m[896]&~m[899]&m[900]&~m[901]&m[902])|(m[896]&m[899]&m[900]&~m[901]&m[902])|(~m[896]&m[899]&m[900]&m[901]&m[902]))&UnbiasedRNG[73])|((m[896]&~m[899]&~m[900]&m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&m[900]&~m[901]&m[902])|(~m[896]&~m[899]&~m[900]&m[901]&m[902])|(m[896]&~m[899]&~m[900]&m[901]&m[902])|(~m[896]&m[899]&~m[900]&m[901]&m[902])|(m[896]&m[899]&~m[900]&m[901]&m[902])|(~m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&m[899]&m[900]&m[901]&m[902]))):InitCond[241];
    m[903] = run?((((m[901]&~m[904]&~m[905]&~m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&m[906]&~m[907])|(m[901]&m[904]&~m[905]&m[906]&~m[907])|(m[901]&~m[904]&m[905]&m[906]&~m[907])|(~m[901]&m[904]&~m[905]&~m[906]&m[907])|(~m[901]&~m[904]&m[905]&~m[906]&m[907])|(m[901]&m[904]&m[905]&~m[906]&m[907])|(~m[901]&m[904]&m[905]&m[906]&m[907]))&UnbiasedRNG[74])|((m[901]&~m[904]&~m[905]&m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&m[905]&~m[906]&m[907])|(~m[901]&~m[904]&~m[905]&m[906]&m[907])|(m[901]&~m[904]&~m[905]&m[906]&m[907])|(~m[901]&m[904]&~m[905]&m[906]&m[907])|(m[901]&m[904]&~m[905]&m[906]&m[907])|(~m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&m[904]&m[905]&m[906]&m[907]))):InitCond[242];
    m[908] = run?((((m[906]&~m[909]&~m[910]&~m[911]&~m[912])|(~m[906]&~m[909]&~m[910]&m[911]&~m[912])|(m[906]&m[909]&~m[910]&m[911]&~m[912])|(m[906]&~m[909]&m[910]&m[911]&~m[912])|(~m[906]&m[909]&~m[910]&~m[911]&m[912])|(~m[906]&~m[909]&m[910]&~m[911]&m[912])|(m[906]&m[909]&m[910]&~m[911]&m[912])|(~m[906]&m[909]&m[910]&m[911]&m[912]))&UnbiasedRNG[75])|((m[906]&~m[909]&~m[910]&m[911]&~m[912])|(~m[906]&~m[909]&~m[910]&~m[911]&m[912])|(m[906]&~m[909]&~m[910]&~m[911]&m[912])|(m[906]&m[909]&~m[910]&~m[911]&m[912])|(m[906]&~m[909]&m[910]&~m[911]&m[912])|(~m[906]&~m[909]&~m[910]&m[911]&m[912])|(m[906]&~m[909]&~m[910]&m[911]&m[912])|(~m[906]&m[909]&~m[910]&m[911]&m[912])|(m[906]&m[909]&~m[910]&m[911]&m[912])|(~m[906]&~m[909]&m[910]&m[911]&m[912])|(m[906]&~m[909]&m[910]&m[911]&m[912])|(m[906]&m[909]&m[910]&m[911]&m[912]))):InitCond[243];
    m[913] = run?((((m[862]&~m[914]&~m[915]&~m[916]&~m[917])|(~m[862]&~m[914]&~m[915]&m[916]&~m[917])|(m[862]&m[914]&~m[915]&m[916]&~m[917])|(m[862]&~m[914]&m[915]&m[916]&~m[917])|(~m[862]&m[914]&~m[915]&~m[916]&m[917])|(~m[862]&~m[914]&m[915]&~m[916]&m[917])|(m[862]&m[914]&m[915]&~m[916]&m[917])|(~m[862]&m[914]&m[915]&m[916]&m[917]))&UnbiasedRNG[76])|((m[862]&~m[914]&~m[915]&m[916]&~m[917])|(~m[862]&~m[914]&~m[915]&~m[916]&m[917])|(m[862]&~m[914]&~m[915]&~m[916]&m[917])|(m[862]&m[914]&~m[915]&~m[916]&m[917])|(m[862]&~m[914]&m[915]&~m[916]&m[917])|(~m[862]&~m[914]&~m[915]&m[916]&m[917])|(m[862]&~m[914]&~m[915]&m[916]&m[917])|(~m[862]&m[914]&~m[915]&m[916]&m[917])|(m[862]&m[914]&~m[915]&m[916]&m[917])|(~m[862]&~m[914]&m[915]&m[916]&m[917])|(m[862]&~m[914]&m[915]&m[916]&m[917])|(m[862]&m[914]&m[915]&m[916]&m[917]))):InitCond[244];
    m[918] = run?((((m[916]&~m[919]&~m[920]&~m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&m[921]&~m[922])|(m[916]&m[919]&~m[920]&m[921]&~m[922])|(m[916]&~m[919]&m[920]&m[921]&~m[922])|(~m[916]&m[919]&~m[920]&~m[921]&m[922])|(~m[916]&~m[919]&m[920]&~m[921]&m[922])|(m[916]&m[919]&m[920]&~m[921]&m[922])|(~m[916]&m[919]&m[920]&m[921]&m[922]))&UnbiasedRNG[77])|((m[916]&~m[919]&~m[920]&m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&m[920]&~m[921]&m[922])|(~m[916]&~m[919]&~m[920]&m[921]&m[922])|(m[916]&~m[919]&~m[920]&m[921]&m[922])|(~m[916]&m[919]&~m[920]&m[921]&m[922])|(m[916]&m[919]&~m[920]&m[921]&m[922])|(~m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&m[919]&m[920]&m[921]&m[922]))):InitCond[245];
    m[923] = run?((((m[921]&~m[924]&~m[925]&~m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&m[926]&~m[927])|(m[921]&m[924]&~m[925]&m[926]&~m[927])|(m[921]&~m[924]&m[925]&m[926]&~m[927])|(~m[921]&m[924]&~m[925]&~m[926]&m[927])|(~m[921]&~m[924]&m[925]&~m[926]&m[927])|(m[921]&m[924]&m[925]&~m[926]&m[927])|(~m[921]&m[924]&m[925]&m[926]&m[927]))&UnbiasedRNG[78])|((m[921]&~m[924]&~m[925]&m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&m[925]&~m[926]&m[927])|(~m[921]&~m[924]&~m[925]&m[926]&m[927])|(m[921]&~m[924]&~m[925]&m[926]&m[927])|(~m[921]&m[924]&~m[925]&m[926]&m[927])|(m[921]&m[924]&~m[925]&m[926]&m[927])|(~m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&m[924]&m[925]&m[926]&m[927]))):InitCond[246];
    m[928] = run?((((m[926]&~m[929]&~m[930]&~m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&m[931]&~m[932])|(m[926]&m[929]&~m[930]&m[931]&~m[932])|(m[926]&~m[929]&m[930]&m[931]&~m[932])|(~m[926]&m[929]&~m[930]&~m[931]&m[932])|(~m[926]&~m[929]&m[930]&~m[931]&m[932])|(m[926]&m[929]&m[930]&~m[931]&m[932])|(~m[926]&m[929]&m[930]&m[931]&m[932]))&UnbiasedRNG[79])|((m[926]&~m[929]&~m[930]&m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&m[930]&~m[931]&m[932])|(~m[926]&~m[929]&~m[930]&m[931]&m[932])|(m[926]&~m[929]&~m[930]&m[931]&m[932])|(~m[926]&m[929]&~m[930]&m[931]&m[932])|(m[926]&m[929]&~m[930]&m[931]&m[932])|(~m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&m[929]&m[930]&m[931]&m[932]))):InitCond[247];
    m[933] = run?((((m[931]&~m[934]&~m[935]&~m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&m[936]&~m[937])|(m[931]&m[934]&~m[935]&m[936]&~m[937])|(m[931]&~m[934]&m[935]&m[936]&~m[937])|(~m[931]&m[934]&~m[935]&~m[936]&m[937])|(~m[931]&~m[934]&m[935]&~m[936]&m[937])|(m[931]&m[934]&m[935]&~m[936]&m[937])|(~m[931]&m[934]&m[935]&m[936]&m[937]))&UnbiasedRNG[80])|((m[931]&~m[934]&~m[935]&m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&m[935]&~m[936]&m[937])|(~m[931]&~m[934]&~m[935]&m[936]&m[937])|(m[931]&~m[934]&~m[935]&m[936]&m[937])|(~m[931]&m[934]&~m[935]&m[936]&m[937])|(m[931]&m[934]&~m[935]&m[936]&m[937])|(~m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&m[934]&m[935]&m[936]&m[937]))):InitCond[248];
    m[938] = run?((((m[936]&~m[939]&~m[940]&~m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&m[941]&~m[942])|(m[936]&m[939]&~m[940]&m[941]&~m[942])|(m[936]&~m[939]&m[940]&m[941]&~m[942])|(~m[936]&m[939]&~m[940]&~m[941]&m[942])|(~m[936]&~m[939]&m[940]&~m[941]&m[942])|(m[936]&m[939]&m[940]&~m[941]&m[942])|(~m[936]&m[939]&m[940]&m[941]&m[942]))&UnbiasedRNG[81])|((m[936]&~m[939]&~m[940]&m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&m[940]&~m[941]&m[942])|(~m[936]&~m[939]&~m[940]&m[941]&m[942])|(m[936]&~m[939]&~m[940]&m[941]&m[942])|(~m[936]&m[939]&~m[940]&m[941]&m[942])|(m[936]&m[939]&~m[940]&m[941]&m[942])|(~m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&m[939]&m[940]&m[941]&m[942]))):InitCond[249];
    m[943] = run?((((m[941]&~m[944]&~m[945]&~m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&m[946]&~m[947])|(m[941]&m[944]&~m[945]&m[946]&~m[947])|(m[941]&~m[944]&m[945]&m[946]&~m[947])|(~m[941]&m[944]&~m[945]&~m[946]&m[947])|(~m[941]&~m[944]&m[945]&~m[946]&m[947])|(m[941]&m[944]&m[945]&~m[946]&m[947])|(~m[941]&m[944]&m[945]&m[946]&m[947]))&UnbiasedRNG[82])|((m[941]&~m[944]&~m[945]&m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&m[945]&~m[946]&m[947])|(~m[941]&~m[944]&~m[945]&m[946]&m[947])|(m[941]&~m[944]&~m[945]&m[946]&m[947])|(~m[941]&m[944]&~m[945]&m[946]&m[947])|(m[941]&m[944]&~m[945]&m[946]&m[947])|(~m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&m[944]&m[945]&m[946]&m[947]))):InitCond[250];
    m[948] = run?((((m[946]&~m[949]&~m[950]&~m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&m[951]&~m[952])|(m[946]&m[949]&~m[950]&m[951]&~m[952])|(m[946]&~m[949]&m[950]&m[951]&~m[952])|(~m[946]&m[949]&~m[950]&~m[951]&m[952])|(~m[946]&~m[949]&m[950]&~m[951]&m[952])|(m[946]&m[949]&m[950]&~m[951]&m[952])|(~m[946]&m[949]&m[950]&m[951]&m[952]))&UnbiasedRNG[83])|((m[946]&~m[949]&~m[950]&m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&m[950]&~m[951]&m[952])|(~m[946]&~m[949]&~m[950]&m[951]&m[952])|(m[946]&~m[949]&~m[950]&m[951]&m[952])|(~m[946]&m[949]&~m[950]&m[951]&m[952])|(m[946]&m[949]&~m[950]&m[951]&m[952])|(~m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&m[949]&m[950]&m[951]&m[952]))):InitCond[251];
    m[953] = run?((((m[951]&~m[954]&~m[955]&~m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&m[956]&~m[957])|(m[951]&m[954]&~m[955]&m[956]&~m[957])|(m[951]&~m[954]&m[955]&m[956]&~m[957])|(~m[951]&m[954]&~m[955]&~m[956]&m[957])|(~m[951]&~m[954]&m[955]&~m[956]&m[957])|(m[951]&m[954]&m[955]&~m[956]&m[957])|(~m[951]&m[954]&m[955]&m[956]&m[957]))&UnbiasedRNG[84])|((m[951]&~m[954]&~m[955]&m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&m[955]&~m[956]&m[957])|(~m[951]&~m[954]&~m[955]&m[956]&m[957])|(m[951]&~m[954]&~m[955]&m[956]&m[957])|(~m[951]&m[954]&~m[955]&m[956]&m[957])|(m[951]&m[954]&~m[955]&m[956]&m[957])|(~m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&m[954]&m[955]&m[956]&m[957]))):InitCond[252];
    m[958] = run?((((m[956]&~m[959]&~m[960]&~m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&m[961]&~m[962])|(m[956]&m[959]&~m[960]&m[961]&~m[962])|(m[956]&~m[959]&m[960]&m[961]&~m[962])|(~m[956]&m[959]&~m[960]&~m[961]&m[962])|(~m[956]&~m[959]&m[960]&~m[961]&m[962])|(m[956]&m[959]&m[960]&~m[961]&m[962])|(~m[956]&m[959]&m[960]&m[961]&m[962]))&UnbiasedRNG[85])|((m[956]&~m[959]&~m[960]&m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&m[960]&~m[961]&m[962])|(~m[956]&~m[959]&~m[960]&m[961]&m[962])|(m[956]&~m[959]&~m[960]&m[961]&m[962])|(~m[956]&m[959]&~m[960]&m[961]&m[962])|(m[956]&m[959]&~m[960]&m[961]&m[962])|(~m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&m[959]&m[960]&m[961]&m[962]))):InitCond[253];
    m[963] = run?((((m[917]&~m[964]&~m[965]&~m[966]&~m[967])|(~m[917]&~m[964]&~m[965]&m[966]&~m[967])|(m[917]&m[964]&~m[965]&m[966]&~m[967])|(m[917]&~m[964]&m[965]&m[966]&~m[967])|(~m[917]&m[964]&~m[965]&~m[966]&m[967])|(~m[917]&~m[964]&m[965]&~m[966]&m[967])|(m[917]&m[964]&m[965]&~m[966]&m[967])|(~m[917]&m[964]&m[965]&m[966]&m[967]))&UnbiasedRNG[86])|((m[917]&~m[964]&~m[965]&m[966]&~m[967])|(~m[917]&~m[964]&~m[965]&~m[966]&m[967])|(m[917]&~m[964]&~m[965]&~m[966]&m[967])|(m[917]&m[964]&~m[965]&~m[966]&m[967])|(m[917]&~m[964]&m[965]&~m[966]&m[967])|(~m[917]&~m[964]&~m[965]&m[966]&m[967])|(m[917]&~m[964]&~m[965]&m[966]&m[967])|(~m[917]&m[964]&~m[965]&m[966]&m[967])|(m[917]&m[964]&~m[965]&m[966]&m[967])|(~m[917]&~m[964]&m[965]&m[966]&m[967])|(m[917]&~m[964]&m[965]&m[966]&m[967])|(m[917]&m[964]&m[965]&m[966]&m[967]))):InitCond[254];
    m[968] = run?((((m[966]&~m[969]&~m[970]&~m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&m[971]&~m[972])|(m[966]&m[969]&~m[970]&m[971]&~m[972])|(m[966]&~m[969]&m[970]&m[971]&~m[972])|(~m[966]&m[969]&~m[970]&~m[971]&m[972])|(~m[966]&~m[969]&m[970]&~m[971]&m[972])|(m[966]&m[969]&m[970]&~m[971]&m[972])|(~m[966]&m[969]&m[970]&m[971]&m[972]))&UnbiasedRNG[87])|((m[966]&~m[969]&~m[970]&m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&m[970]&~m[971]&m[972])|(~m[966]&~m[969]&~m[970]&m[971]&m[972])|(m[966]&~m[969]&~m[970]&m[971]&m[972])|(~m[966]&m[969]&~m[970]&m[971]&m[972])|(m[966]&m[969]&~m[970]&m[971]&m[972])|(~m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&m[969]&m[970]&m[971]&m[972]))):InitCond[255];
    m[973] = run?((((m[971]&~m[974]&~m[975]&~m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&m[976]&~m[977])|(m[971]&m[974]&~m[975]&m[976]&~m[977])|(m[971]&~m[974]&m[975]&m[976]&~m[977])|(~m[971]&m[974]&~m[975]&~m[976]&m[977])|(~m[971]&~m[974]&m[975]&~m[976]&m[977])|(m[971]&m[974]&m[975]&~m[976]&m[977])|(~m[971]&m[974]&m[975]&m[976]&m[977]))&UnbiasedRNG[88])|((m[971]&~m[974]&~m[975]&m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&m[975]&~m[976]&m[977])|(~m[971]&~m[974]&~m[975]&m[976]&m[977])|(m[971]&~m[974]&~m[975]&m[976]&m[977])|(~m[971]&m[974]&~m[975]&m[976]&m[977])|(m[971]&m[974]&~m[975]&m[976]&m[977])|(~m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&m[974]&m[975]&m[976]&m[977]))):InitCond[256];
    m[978] = run?((((m[976]&~m[979]&~m[980]&~m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&m[981]&~m[982])|(m[976]&m[979]&~m[980]&m[981]&~m[982])|(m[976]&~m[979]&m[980]&m[981]&~m[982])|(~m[976]&m[979]&~m[980]&~m[981]&m[982])|(~m[976]&~m[979]&m[980]&~m[981]&m[982])|(m[976]&m[979]&m[980]&~m[981]&m[982])|(~m[976]&m[979]&m[980]&m[981]&m[982]))&UnbiasedRNG[89])|((m[976]&~m[979]&~m[980]&m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&m[980]&~m[981]&m[982])|(~m[976]&~m[979]&~m[980]&m[981]&m[982])|(m[976]&~m[979]&~m[980]&m[981]&m[982])|(~m[976]&m[979]&~m[980]&m[981]&m[982])|(m[976]&m[979]&~m[980]&m[981]&m[982])|(~m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&m[979]&m[980]&m[981]&m[982]))):InitCond[257];
    m[983] = run?((((m[981]&~m[984]&~m[985]&~m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&m[986]&~m[987])|(m[981]&m[984]&~m[985]&m[986]&~m[987])|(m[981]&~m[984]&m[985]&m[986]&~m[987])|(~m[981]&m[984]&~m[985]&~m[986]&m[987])|(~m[981]&~m[984]&m[985]&~m[986]&m[987])|(m[981]&m[984]&m[985]&~m[986]&m[987])|(~m[981]&m[984]&m[985]&m[986]&m[987]))&UnbiasedRNG[90])|((m[981]&~m[984]&~m[985]&m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&m[985]&~m[986]&m[987])|(~m[981]&~m[984]&~m[985]&m[986]&m[987])|(m[981]&~m[984]&~m[985]&m[986]&m[987])|(~m[981]&m[984]&~m[985]&m[986]&m[987])|(m[981]&m[984]&~m[985]&m[986]&m[987])|(~m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&m[984]&m[985]&m[986]&m[987]))):InitCond[258];
    m[988] = run?((((m[986]&~m[989]&~m[990]&~m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&m[991]&~m[992])|(m[986]&m[989]&~m[990]&m[991]&~m[992])|(m[986]&~m[989]&m[990]&m[991]&~m[992])|(~m[986]&m[989]&~m[990]&~m[991]&m[992])|(~m[986]&~m[989]&m[990]&~m[991]&m[992])|(m[986]&m[989]&m[990]&~m[991]&m[992])|(~m[986]&m[989]&m[990]&m[991]&m[992]))&UnbiasedRNG[91])|((m[986]&~m[989]&~m[990]&m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&m[990]&~m[991]&m[992])|(~m[986]&~m[989]&~m[990]&m[991]&m[992])|(m[986]&~m[989]&~m[990]&m[991]&m[992])|(~m[986]&m[989]&~m[990]&m[991]&m[992])|(m[986]&m[989]&~m[990]&m[991]&m[992])|(~m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&m[989]&m[990]&m[991]&m[992]))):InitCond[259];
    m[993] = run?((((m[991]&~m[994]&~m[995]&~m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&m[996]&~m[997])|(m[991]&m[994]&~m[995]&m[996]&~m[997])|(m[991]&~m[994]&m[995]&m[996]&~m[997])|(~m[991]&m[994]&~m[995]&~m[996]&m[997])|(~m[991]&~m[994]&m[995]&~m[996]&m[997])|(m[991]&m[994]&m[995]&~m[996]&m[997])|(~m[991]&m[994]&m[995]&m[996]&m[997]))&UnbiasedRNG[92])|((m[991]&~m[994]&~m[995]&m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&m[995]&~m[996]&m[997])|(~m[991]&~m[994]&~m[995]&m[996]&m[997])|(m[991]&~m[994]&~m[995]&m[996]&m[997])|(~m[991]&m[994]&~m[995]&m[996]&m[997])|(m[991]&m[994]&~m[995]&m[996]&m[997])|(~m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&m[994]&m[995]&m[996]&m[997]))):InitCond[260];
    m[998] = run?((((m[996]&~m[999]&~m[1000]&~m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&~m[1002])|(~m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&m[999]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[93])|((m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&m[999]&m[1000]&m[1001]&m[1002]))):InitCond[261];
    m[1003] = run?((((m[1001]&~m[1004]&~m[1005]&~m[1006]&~m[1007])|(~m[1001]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(m[1001]&m[1004]&~m[1005]&m[1006]&~m[1007])|(m[1001]&~m[1004]&m[1005]&m[1006]&~m[1007])|(~m[1001]&m[1004]&~m[1005]&~m[1006]&m[1007])|(~m[1001]&~m[1004]&m[1005]&~m[1006]&m[1007])|(m[1001]&m[1004]&m[1005]&~m[1006]&m[1007])|(~m[1001]&m[1004]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[94])|((m[1001]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(~m[1001]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[1001]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[1001]&m[1004]&~m[1005]&~m[1006]&m[1007])|(m[1001]&~m[1004]&m[1005]&~m[1006]&m[1007])|(~m[1001]&~m[1004]&~m[1005]&m[1006]&m[1007])|(m[1001]&~m[1004]&~m[1005]&m[1006]&m[1007])|(~m[1001]&m[1004]&~m[1005]&m[1006]&m[1007])|(m[1001]&m[1004]&~m[1005]&m[1006]&m[1007])|(~m[1001]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[1001]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[1001]&m[1004]&m[1005]&m[1006]&m[1007]))):InitCond[262];
    m[1008] = run?((((m[967]&~m[1009]&~m[1010]&~m[1011]&~m[1012])|(~m[967]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(m[967]&m[1009]&~m[1010]&m[1011]&~m[1012])|(m[967]&~m[1009]&m[1010]&m[1011]&~m[1012])|(~m[967]&m[1009]&~m[1010]&~m[1011]&m[1012])|(~m[967]&~m[1009]&m[1010]&~m[1011]&m[1012])|(m[967]&m[1009]&m[1010]&~m[1011]&m[1012])|(~m[967]&m[1009]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[95])|((m[967]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(~m[967]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[967]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[967]&m[1009]&~m[1010]&~m[1011]&m[1012])|(m[967]&~m[1009]&m[1010]&~m[1011]&m[1012])|(~m[967]&~m[1009]&~m[1010]&m[1011]&m[1012])|(m[967]&~m[1009]&~m[1010]&m[1011]&m[1012])|(~m[967]&m[1009]&~m[1010]&m[1011]&m[1012])|(m[967]&m[1009]&~m[1010]&m[1011]&m[1012])|(~m[967]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[967]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[967]&m[1009]&m[1010]&m[1011]&m[1012]))):InitCond[263];
    m[1013] = run?((((m[1011]&~m[1014]&~m[1015]&~m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&~m[1017])|(~m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[96])|((m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))):InitCond[264];
    m[1018] = run?((((m[1016]&~m[1019]&~m[1020]&~m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&~m[1022])|(~m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[97])|((m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))):InitCond[265];
    m[1023] = run?((((m[1021]&~m[1024]&~m[1025]&~m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&~m[1027])|(~m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[98])|((m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))):InitCond[266];
    m[1028] = run?((((m[1026]&~m[1029]&~m[1030]&~m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&~m[1032])|(~m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[99])|((m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))):InitCond[267];
    m[1033] = run?((((m[1031]&~m[1034]&~m[1035]&~m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&~m[1037])|(~m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&m[1034]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[100])|((m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&m[1036]&m[1037]))):InitCond[268];
    m[1038] = run?((((m[1036]&~m[1039]&~m[1040]&~m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&~m[1042])|(~m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[101])|((m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))):InitCond[269];
    m[1043] = run?((((m[1041]&~m[1044]&~m[1045]&~m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&~m[1047])|(~m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[102])|((m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))):InitCond[270];
    m[1048] = run?((((m[1012]&~m[1049]&~m[1050]&~m[1051]&~m[1052])|(~m[1012]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1012]&m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1012]&~m[1049]&m[1050]&m[1051]&~m[1052])|(~m[1012]&m[1049]&~m[1050]&~m[1051]&m[1052])|(~m[1012]&~m[1049]&m[1050]&~m[1051]&m[1052])|(m[1012]&m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1012]&m[1049]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[103])|((m[1012]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(~m[1012]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1012]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1012]&m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1012]&~m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1012]&~m[1049]&~m[1050]&m[1051]&m[1052])|(m[1012]&~m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1012]&m[1049]&~m[1050]&m[1051]&m[1052])|(m[1012]&m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1012]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1012]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1012]&m[1049]&m[1050]&m[1051]&m[1052]))):InitCond[271];
    m[1053] = run?((((m[1051]&~m[1054]&~m[1055]&~m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&~m[1057])|(~m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[104])|((m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))):InitCond[272];
    m[1058] = run?((((m[1056]&~m[1059]&~m[1060]&~m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&~m[1062])|(~m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&m[1059]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[105])|((m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&m[1061]&m[1062]))):InitCond[273];
    m[1063] = run?((((m[1061]&~m[1064]&~m[1065]&~m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&~m[1067])|(~m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[106])|((m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))):InitCond[274];
    m[1068] = run?((((m[1066]&~m[1069]&~m[1070]&~m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&~m[1072])|(~m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&m[1069]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[107])|((m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&m[1071]&m[1072]))):InitCond[275];
    m[1073] = run?((((m[1071]&~m[1074]&~m[1075]&~m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&~m[1077])|(~m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[108])|((m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))):InitCond[276];
    m[1078] = run?((((m[1076]&~m[1079]&~m[1080]&~m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&~m[1082])|(~m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[109])|((m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))):InitCond[277];
    m[1083] = run?((((m[1052]&~m[1084]&~m[1085]&~m[1086]&~m[1087])|(~m[1052]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1052]&m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1052]&~m[1084]&m[1085]&m[1086]&~m[1087])|(~m[1052]&m[1084]&~m[1085]&~m[1086]&m[1087])|(~m[1052]&~m[1084]&m[1085]&~m[1086]&m[1087])|(m[1052]&m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1052]&m[1084]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[110])|((m[1052]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(~m[1052]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1052]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1052]&m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1052]&~m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1052]&~m[1084]&~m[1085]&m[1086]&m[1087])|(m[1052]&~m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1052]&m[1084]&~m[1085]&m[1086]&m[1087])|(m[1052]&m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1052]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1052]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1052]&m[1084]&m[1085]&m[1086]&m[1087]))):InitCond[278];
    m[1088] = run?((((m[1086]&~m[1089]&~m[1090]&~m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&~m[1092])|(~m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[111])|((m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))):InitCond[279];
    m[1093] = run?((((m[1091]&~m[1094]&~m[1095]&~m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&~m[1097])|(~m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[112])|((m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))):InitCond[280];
    m[1098] = run?((((m[1096]&~m[1099]&~m[1100]&~m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&~m[1102])|(~m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[113])|((m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))):InitCond[281];
    m[1103] = run?((((m[1101]&~m[1104]&~m[1105]&~m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&~m[1107])|(~m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[114])|((m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))):InitCond[282];
    m[1108] = run?((((m[1106]&~m[1109]&~m[1110]&~m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&~m[1112])|(~m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&m[1109]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[115])|((m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&m[1111]&m[1112]))):InitCond[283];
    m[1113] = run?((((m[1087]&~m[1114]&~m[1115]&~m[1116]&~m[1117])|(~m[1087]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1087]&m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1087]&~m[1114]&m[1115]&m[1116]&~m[1117])|(~m[1087]&m[1114]&~m[1115]&~m[1116]&m[1117])|(~m[1087]&~m[1114]&m[1115]&~m[1116]&m[1117])|(m[1087]&m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1087]&m[1114]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[116])|((m[1087]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(~m[1087]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1087]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1087]&m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1087]&~m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1087]&~m[1114]&~m[1115]&m[1116]&m[1117])|(m[1087]&~m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1087]&m[1114]&~m[1115]&m[1116]&m[1117])|(m[1087]&m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1087]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1087]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1087]&m[1114]&m[1115]&m[1116]&m[1117]))):InitCond[284];
    m[1118] = run?((((m[1116]&~m[1119]&~m[1120]&~m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&~m[1122])|(~m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&m[1119]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[117])|((m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&m[1121]&m[1122]))):InitCond[285];
    m[1123] = run?((((m[1121]&~m[1124]&~m[1125]&~m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&~m[1127])|(~m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[118])|((m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))):InitCond[286];
    m[1128] = run?((((m[1126]&~m[1129]&~m[1130]&~m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&~m[1132])|(~m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[119])|((m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))):InitCond[287];
    m[1133] = run?((((m[1131]&~m[1134]&~m[1135]&~m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&~m[1137])|(~m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[120])|((m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))):InitCond[288];
    m[1138] = run?((((m[1117]&~m[1139]&~m[1140]&~m[1141]&~m[1142])|(~m[1117]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1117]&m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1117]&~m[1139]&m[1140]&m[1141]&~m[1142])|(~m[1117]&m[1139]&~m[1140]&~m[1141]&m[1142])|(~m[1117]&~m[1139]&m[1140]&~m[1141]&m[1142])|(m[1117]&m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1117]&m[1139]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[121])|((m[1117]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(~m[1117]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1117]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1117]&m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1117]&~m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1117]&~m[1139]&~m[1140]&m[1141]&m[1142])|(m[1117]&~m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1117]&m[1139]&~m[1140]&m[1141]&m[1142])|(m[1117]&m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1117]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1117]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1117]&m[1139]&m[1140]&m[1141]&m[1142]))):InitCond[289];
    m[1143] = run?((((m[1141]&~m[1144]&~m[1145]&~m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&~m[1147])|(~m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[122])|((m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))):InitCond[290];
    m[1148] = run?((((m[1146]&~m[1149]&~m[1150]&~m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&~m[1152])|(~m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[123])|((m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))):InitCond[291];
    m[1153] = run?((((m[1151]&~m[1154]&~m[1155]&~m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&~m[1157])|(~m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&m[1154]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[124])|((m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&m[1156]&m[1157]))):InitCond[292];
    m[1158] = run?((((m[1142]&~m[1159]&~m[1160]&~m[1161]&~m[1162])|(~m[1142]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1142]&m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1142]&~m[1159]&m[1160]&m[1161]&~m[1162])|(~m[1142]&m[1159]&~m[1160]&~m[1161]&m[1162])|(~m[1142]&~m[1159]&m[1160]&~m[1161]&m[1162])|(m[1142]&m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1142]&m[1159]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[125])|((m[1142]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(~m[1142]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1142]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1142]&m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1142]&~m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1142]&~m[1159]&~m[1160]&m[1161]&m[1162])|(m[1142]&~m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1142]&m[1159]&~m[1160]&m[1161]&m[1162])|(m[1142]&m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1142]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1142]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1142]&m[1159]&m[1160]&m[1161]&m[1162]))):InitCond[293];
    m[1163] = run?((((m[1161]&~m[1164]&~m[1165]&~m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&~m[1167])|(~m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[126])|((m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))):InitCond[294];
    m[1168] = run?((((m[1166]&~m[1169]&~m[1170]&~m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&~m[1172])|(~m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[127])|((m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))):InitCond[295];
    m[1173] = run?((((m[1162]&~m[1174]&~m[1175]&~m[1176]&~m[1177])|(~m[1162]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1162]&m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1162]&~m[1174]&m[1175]&m[1176]&~m[1177])|(~m[1162]&m[1174]&~m[1175]&~m[1176]&m[1177])|(~m[1162]&~m[1174]&m[1175]&~m[1176]&m[1177])|(m[1162]&m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1162]&m[1174]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[128])|((m[1162]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(~m[1162]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1162]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1162]&m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1162]&~m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1162]&~m[1174]&~m[1175]&m[1176]&m[1177])|(m[1162]&~m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1162]&m[1174]&~m[1175]&m[1176]&m[1177])|(m[1162]&m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1162]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1162]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1162]&m[1174]&m[1175]&m[1176]&m[1177]))):InitCond[296];
    m[1178] = run?((((m[1176]&~m[1179]&~m[1180]&~m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&~m[1182])|(~m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[129])|((m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))):InitCond[297];
    m[1183] = run?((((m[1177]&~m[1184]&~m[1185]&~m[1186]&~m[1187])|(~m[1177]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1177]&m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1177]&~m[1184]&m[1185]&m[1186]&~m[1187])|(~m[1177]&m[1184]&~m[1185]&~m[1186]&m[1187])|(~m[1177]&~m[1184]&m[1185]&~m[1186]&m[1187])|(m[1177]&m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1177]&m[1184]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[130])|((m[1177]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(~m[1177]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1177]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1177]&m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1177]&~m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1177]&~m[1184]&~m[1185]&m[1186]&m[1187])|(m[1177]&~m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1177]&m[1184]&~m[1185]&m[1186]&m[1187])|(m[1177]&m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1177]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1177]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1177]&m[1184]&m[1185]&m[1186]&m[1187]))):InitCond[298];
end

always @(posedge color1_clk) begin
    m[24] = run?((((m[0]&m[96]&~m[97]&~m[98]&~m[99])|(m[0]&~m[96]&m[97]&~m[98]&~m[99])|(~m[0]&m[96]&m[97]&~m[98]&~m[99])|(m[0]&~m[96]&~m[97]&m[98]&~m[99])|(~m[0]&m[96]&~m[97]&m[98]&~m[99])|(~m[0]&~m[96]&m[97]&m[98]&~m[99])|(m[0]&~m[96]&~m[97]&~m[98]&m[99])|(~m[0]&m[96]&~m[97]&~m[98]&m[99])|(~m[0]&~m[96]&m[97]&~m[98]&m[99])|(~m[0]&~m[96]&~m[97]&m[98]&m[99]))&BiasedRNG[168])|(((m[0]&m[96]&m[97]&~m[98]&~m[99])|(m[0]&m[96]&~m[97]&m[98]&~m[99])|(m[0]&~m[96]&m[97]&m[98]&~m[99])|(~m[0]&m[96]&m[97]&m[98]&~m[99])|(m[0]&m[96]&~m[97]&~m[98]&m[99])|(m[0]&~m[96]&m[97]&~m[98]&m[99])|(~m[0]&m[96]&m[97]&~m[98]&m[99])|(m[0]&~m[96]&~m[97]&m[98]&m[99])|(~m[0]&m[96]&~m[97]&m[98]&m[99])|(~m[0]&~m[96]&m[97]&m[98]&m[99]))&~BiasedRNG[168])|((m[0]&m[96]&m[97]&m[98]&~m[99])|(m[0]&m[96]&m[97]&~m[98]&m[99])|(m[0]&m[96]&~m[97]&m[98]&m[99])|(m[0]&~m[96]&m[97]&m[98]&m[99])|(~m[0]&m[96]&m[97]&m[98]&m[99])|(m[0]&m[96]&m[97]&m[98]&m[99]))):InitCond[299];
    m[25] = run?((((m[0]&m[100]&~m[101]&~m[102]&~m[103])|(m[0]&~m[100]&m[101]&~m[102]&~m[103])|(~m[0]&m[100]&m[101]&~m[102]&~m[103])|(m[0]&~m[100]&~m[101]&m[102]&~m[103])|(~m[0]&m[100]&~m[101]&m[102]&~m[103])|(~m[0]&~m[100]&m[101]&m[102]&~m[103])|(m[0]&~m[100]&~m[101]&~m[102]&m[103])|(~m[0]&m[100]&~m[101]&~m[102]&m[103])|(~m[0]&~m[100]&m[101]&~m[102]&m[103])|(~m[0]&~m[100]&~m[101]&m[102]&m[103]))&BiasedRNG[169])|(((m[0]&m[100]&m[101]&~m[102]&~m[103])|(m[0]&m[100]&~m[101]&m[102]&~m[103])|(m[0]&~m[100]&m[101]&m[102]&~m[103])|(~m[0]&m[100]&m[101]&m[102]&~m[103])|(m[0]&m[100]&~m[101]&~m[102]&m[103])|(m[0]&~m[100]&m[101]&~m[102]&m[103])|(~m[0]&m[100]&m[101]&~m[102]&m[103])|(m[0]&~m[100]&~m[101]&m[102]&m[103])|(~m[0]&m[100]&~m[101]&m[102]&m[103])|(~m[0]&~m[100]&m[101]&m[102]&m[103]))&~BiasedRNG[169])|((m[0]&m[100]&m[101]&m[102]&~m[103])|(m[0]&m[100]&m[101]&~m[102]&m[103])|(m[0]&m[100]&~m[101]&m[102]&m[103])|(m[0]&~m[100]&m[101]&m[102]&m[103])|(~m[0]&m[100]&m[101]&m[102]&m[103])|(m[0]&m[100]&m[101]&m[102]&m[103]))):InitCond[300];
    m[26] = run?((((m[0]&m[104]&~m[105]&~m[106]&~m[107])|(m[0]&~m[104]&m[105]&~m[106]&~m[107])|(~m[0]&m[104]&m[105]&~m[106]&~m[107])|(m[0]&~m[104]&~m[105]&m[106]&~m[107])|(~m[0]&m[104]&~m[105]&m[106]&~m[107])|(~m[0]&~m[104]&m[105]&m[106]&~m[107])|(m[0]&~m[104]&~m[105]&~m[106]&m[107])|(~m[0]&m[104]&~m[105]&~m[106]&m[107])|(~m[0]&~m[104]&m[105]&~m[106]&m[107])|(~m[0]&~m[104]&~m[105]&m[106]&m[107]))&BiasedRNG[170])|(((m[0]&m[104]&m[105]&~m[106]&~m[107])|(m[0]&m[104]&~m[105]&m[106]&~m[107])|(m[0]&~m[104]&m[105]&m[106]&~m[107])|(~m[0]&m[104]&m[105]&m[106]&~m[107])|(m[0]&m[104]&~m[105]&~m[106]&m[107])|(m[0]&~m[104]&m[105]&~m[106]&m[107])|(~m[0]&m[104]&m[105]&~m[106]&m[107])|(m[0]&~m[104]&~m[105]&m[106]&m[107])|(~m[0]&m[104]&~m[105]&m[106]&m[107])|(~m[0]&~m[104]&m[105]&m[106]&m[107]))&~BiasedRNG[170])|((m[0]&m[104]&m[105]&m[106]&~m[107])|(m[0]&m[104]&m[105]&~m[106]&m[107])|(m[0]&m[104]&~m[105]&m[106]&m[107])|(m[0]&~m[104]&m[105]&m[106]&m[107])|(~m[0]&m[104]&m[105]&m[106]&m[107])|(m[0]&m[104]&m[105]&m[106]&m[107]))):InitCond[301];
    m[27] = run?((((m[1]&m[108]&~m[109]&~m[110]&~m[111])|(m[1]&~m[108]&m[109]&~m[110]&~m[111])|(~m[1]&m[108]&m[109]&~m[110]&~m[111])|(m[1]&~m[108]&~m[109]&m[110]&~m[111])|(~m[1]&m[108]&~m[109]&m[110]&~m[111])|(~m[1]&~m[108]&m[109]&m[110]&~m[111])|(m[1]&~m[108]&~m[109]&~m[110]&m[111])|(~m[1]&m[108]&~m[109]&~m[110]&m[111])|(~m[1]&~m[108]&m[109]&~m[110]&m[111])|(~m[1]&~m[108]&~m[109]&m[110]&m[111]))&BiasedRNG[171])|(((m[1]&m[108]&m[109]&~m[110]&~m[111])|(m[1]&m[108]&~m[109]&m[110]&~m[111])|(m[1]&~m[108]&m[109]&m[110]&~m[111])|(~m[1]&m[108]&m[109]&m[110]&~m[111])|(m[1]&m[108]&~m[109]&~m[110]&m[111])|(m[1]&~m[108]&m[109]&~m[110]&m[111])|(~m[1]&m[108]&m[109]&~m[110]&m[111])|(m[1]&~m[108]&~m[109]&m[110]&m[111])|(~m[1]&m[108]&~m[109]&m[110]&m[111])|(~m[1]&~m[108]&m[109]&m[110]&m[111]))&~BiasedRNG[171])|((m[1]&m[108]&m[109]&m[110]&~m[111])|(m[1]&m[108]&m[109]&~m[110]&m[111])|(m[1]&m[108]&~m[109]&m[110]&m[111])|(m[1]&~m[108]&m[109]&m[110]&m[111])|(~m[1]&m[108]&m[109]&m[110]&m[111])|(m[1]&m[108]&m[109]&m[110]&m[111]))):InitCond[302];
    m[28] = run?((((m[1]&m[112]&~m[113]&~m[114]&~m[115])|(m[1]&~m[112]&m[113]&~m[114]&~m[115])|(~m[1]&m[112]&m[113]&~m[114]&~m[115])|(m[1]&~m[112]&~m[113]&m[114]&~m[115])|(~m[1]&m[112]&~m[113]&m[114]&~m[115])|(~m[1]&~m[112]&m[113]&m[114]&~m[115])|(m[1]&~m[112]&~m[113]&~m[114]&m[115])|(~m[1]&m[112]&~m[113]&~m[114]&m[115])|(~m[1]&~m[112]&m[113]&~m[114]&m[115])|(~m[1]&~m[112]&~m[113]&m[114]&m[115]))&BiasedRNG[172])|(((m[1]&m[112]&m[113]&~m[114]&~m[115])|(m[1]&m[112]&~m[113]&m[114]&~m[115])|(m[1]&~m[112]&m[113]&m[114]&~m[115])|(~m[1]&m[112]&m[113]&m[114]&~m[115])|(m[1]&m[112]&~m[113]&~m[114]&m[115])|(m[1]&~m[112]&m[113]&~m[114]&m[115])|(~m[1]&m[112]&m[113]&~m[114]&m[115])|(m[1]&~m[112]&~m[113]&m[114]&m[115])|(~m[1]&m[112]&~m[113]&m[114]&m[115])|(~m[1]&~m[112]&m[113]&m[114]&m[115]))&~BiasedRNG[172])|((m[1]&m[112]&m[113]&m[114]&~m[115])|(m[1]&m[112]&m[113]&~m[114]&m[115])|(m[1]&m[112]&~m[113]&m[114]&m[115])|(m[1]&~m[112]&m[113]&m[114]&m[115])|(~m[1]&m[112]&m[113]&m[114]&m[115])|(m[1]&m[112]&m[113]&m[114]&m[115]))):InitCond[303];
    m[29] = run?((((m[1]&m[116]&~m[117]&~m[118]&~m[119])|(m[1]&~m[116]&m[117]&~m[118]&~m[119])|(~m[1]&m[116]&m[117]&~m[118]&~m[119])|(m[1]&~m[116]&~m[117]&m[118]&~m[119])|(~m[1]&m[116]&~m[117]&m[118]&~m[119])|(~m[1]&~m[116]&m[117]&m[118]&~m[119])|(m[1]&~m[116]&~m[117]&~m[118]&m[119])|(~m[1]&m[116]&~m[117]&~m[118]&m[119])|(~m[1]&~m[116]&m[117]&~m[118]&m[119])|(~m[1]&~m[116]&~m[117]&m[118]&m[119]))&BiasedRNG[173])|(((m[1]&m[116]&m[117]&~m[118]&~m[119])|(m[1]&m[116]&~m[117]&m[118]&~m[119])|(m[1]&~m[116]&m[117]&m[118]&~m[119])|(~m[1]&m[116]&m[117]&m[118]&~m[119])|(m[1]&m[116]&~m[117]&~m[118]&m[119])|(m[1]&~m[116]&m[117]&~m[118]&m[119])|(~m[1]&m[116]&m[117]&~m[118]&m[119])|(m[1]&~m[116]&~m[117]&m[118]&m[119])|(~m[1]&m[116]&~m[117]&m[118]&m[119])|(~m[1]&~m[116]&m[117]&m[118]&m[119]))&~BiasedRNG[173])|((m[1]&m[116]&m[117]&m[118]&~m[119])|(m[1]&m[116]&m[117]&~m[118]&m[119])|(m[1]&m[116]&~m[117]&m[118]&m[119])|(m[1]&~m[116]&m[117]&m[118]&m[119])|(~m[1]&m[116]&m[117]&m[118]&m[119])|(m[1]&m[116]&m[117]&m[118]&m[119]))):InitCond[304];
    m[30] = run?((((m[2]&m[120]&~m[121]&~m[122]&~m[123])|(m[2]&~m[120]&m[121]&~m[122]&~m[123])|(~m[2]&m[120]&m[121]&~m[122]&~m[123])|(m[2]&~m[120]&~m[121]&m[122]&~m[123])|(~m[2]&m[120]&~m[121]&m[122]&~m[123])|(~m[2]&~m[120]&m[121]&m[122]&~m[123])|(m[2]&~m[120]&~m[121]&~m[122]&m[123])|(~m[2]&m[120]&~m[121]&~m[122]&m[123])|(~m[2]&~m[120]&m[121]&~m[122]&m[123])|(~m[2]&~m[120]&~m[121]&m[122]&m[123]))&BiasedRNG[174])|(((m[2]&m[120]&m[121]&~m[122]&~m[123])|(m[2]&m[120]&~m[121]&m[122]&~m[123])|(m[2]&~m[120]&m[121]&m[122]&~m[123])|(~m[2]&m[120]&m[121]&m[122]&~m[123])|(m[2]&m[120]&~m[121]&~m[122]&m[123])|(m[2]&~m[120]&m[121]&~m[122]&m[123])|(~m[2]&m[120]&m[121]&~m[122]&m[123])|(m[2]&~m[120]&~m[121]&m[122]&m[123])|(~m[2]&m[120]&~m[121]&m[122]&m[123])|(~m[2]&~m[120]&m[121]&m[122]&m[123]))&~BiasedRNG[174])|((m[2]&m[120]&m[121]&m[122]&~m[123])|(m[2]&m[120]&m[121]&~m[122]&m[123])|(m[2]&m[120]&~m[121]&m[122]&m[123])|(m[2]&~m[120]&m[121]&m[122]&m[123])|(~m[2]&m[120]&m[121]&m[122]&m[123])|(m[2]&m[120]&m[121]&m[122]&m[123]))):InitCond[305];
    m[31] = run?((((m[2]&m[124]&~m[125]&~m[126]&~m[127])|(m[2]&~m[124]&m[125]&~m[126]&~m[127])|(~m[2]&m[124]&m[125]&~m[126]&~m[127])|(m[2]&~m[124]&~m[125]&m[126]&~m[127])|(~m[2]&m[124]&~m[125]&m[126]&~m[127])|(~m[2]&~m[124]&m[125]&m[126]&~m[127])|(m[2]&~m[124]&~m[125]&~m[126]&m[127])|(~m[2]&m[124]&~m[125]&~m[126]&m[127])|(~m[2]&~m[124]&m[125]&~m[126]&m[127])|(~m[2]&~m[124]&~m[125]&m[126]&m[127]))&BiasedRNG[175])|(((m[2]&m[124]&m[125]&~m[126]&~m[127])|(m[2]&m[124]&~m[125]&m[126]&~m[127])|(m[2]&~m[124]&m[125]&m[126]&~m[127])|(~m[2]&m[124]&m[125]&m[126]&~m[127])|(m[2]&m[124]&~m[125]&~m[126]&m[127])|(m[2]&~m[124]&m[125]&~m[126]&m[127])|(~m[2]&m[124]&m[125]&~m[126]&m[127])|(m[2]&~m[124]&~m[125]&m[126]&m[127])|(~m[2]&m[124]&~m[125]&m[126]&m[127])|(~m[2]&~m[124]&m[125]&m[126]&m[127]))&~BiasedRNG[175])|((m[2]&m[124]&m[125]&m[126]&~m[127])|(m[2]&m[124]&m[125]&~m[126]&m[127])|(m[2]&m[124]&~m[125]&m[126]&m[127])|(m[2]&~m[124]&m[125]&m[126]&m[127])|(~m[2]&m[124]&m[125]&m[126]&m[127])|(m[2]&m[124]&m[125]&m[126]&m[127]))):InitCond[306];
    m[32] = run?((((m[2]&m[128]&~m[129]&~m[130]&~m[131])|(m[2]&~m[128]&m[129]&~m[130]&~m[131])|(~m[2]&m[128]&m[129]&~m[130]&~m[131])|(m[2]&~m[128]&~m[129]&m[130]&~m[131])|(~m[2]&m[128]&~m[129]&m[130]&~m[131])|(~m[2]&~m[128]&m[129]&m[130]&~m[131])|(m[2]&~m[128]&~m[129]&~m[130]&m[131])|(~m[2]&m[128]&~m[129]&~m[130]&m[131])|(~m[2]&~m[128]&m[129]&~m[130]&m[131])|(~m[2]&~m[128]&~m[129]&m[130]&m[131]))&BiasedRNG[176])|(((m[2]&m[128]&m[129]&~m[130]&~m[131])|(m[2]&m[128]&~m[129]&m[130]&~m[131])|(m[2]&~m[128]&m[129]&m[130]&~m[131])|(~m[2]&m[128]&m[129]&m[130]&~m[131])|(m[2]&m[128]&~m[129]&~m[130]&m[131])|(m[2]&~m[128]&m[129]&~m[130]&m[131])|(~m[2]&m[128]&m[129]&~m[130]&m[131])|(m[2]&~m[128]&~m[129]&m[130]&m[131])|(~m[2]&m[128]&~m[129]&m[130]&m[131])|(~m[2]&~m[128]&m[129]&m[130]&m[131]))&~BiasedRNG[176])|((m[2]&m[128]&m[129]&m[130]&~m[131])|(m[2]&m[128]&m[129]&~m[130]&m[131])|(m[2]&m[128]&~m[129]&m[130]&m[131])|(m[2]&~m[128]&m[129]&m[130]&m[131])|(~m[2]&m[128]&m[129]&m[130]&m[131])|(m[2]&m[128]&m[129]&m[130]&m[131]))):InitCond[307];
    m[33] = run?((((m[3]&m[132]&~m[133]&~m[134]&~m[135])|(m[3]&~m[132]&m[133]&~m[134]&~m[135])|(~m[3]&m[132]&m[133]&~m[134]&~m[135])|(m[3]&~m[132]&~m[133]&m[134]&~m[135])|(~m[3]&m[132]&~m[133]&m[134]&~m[135])|(~m[3]&~m[132]&m[133]&m[134]&~m[135])|(m[3]&~m[132]&~m[133]&~m[134]&m[135])|(~m[3]&m[132]&~m[133]&~m[134]&m[135])|(~m[3]&~m[132]&m[133]&~m[134]&m[135])|(~m[3]&~m[132]&~m[133]&m[134]&m[135]))&BiasedRNG[177])|(((m[3]&m[132]&m[133]&~m[134]&~m[135])|(m[3]&m[132]&~m[133]&m[134]&~m[135])|(m[3]&~m[132]&m[133]&m[134]&~m[135])|(~m[3]&m[132]&m[133]&m[134]&~m[135])|(m[3]&m[132]&~m[133]&~m[134]&m[135])|(m[3]&~m[132]&m[133]&~m[134]&m[135])|(~m[3]&m[132]&m[133]&~m[134]&m[135])|(m[3]&~m[132]&~m[133]&m[134]&m[135])|(~m[3]&m[132]&~m[133]&m[134]&m[135])|(~m[3]&~m[132]&m[133]&m[134]&m[135]))&~BiasedRNG[177])|((m[3]&m[132]&m[133]&m[134]&~m[135])|(m[3]&m[132]&m[133]&~m[134]&m[135])|(m[3]&m[132]&~m[133]&m[134]&m[135])|(m[3]&~m[132]&m[133]&m[134]&m[135])|(~m[3]&m[132]&m[133]&m[134]&m[135])|(m[3]&m[132]&m[133]&m[134]&m[135]))):InitCond[308];
    m[34] = run?((((m[3]&m[136]&~m[137]&~m[138]&~m[139])|(m[3]&~m[136]&m[137]&~m[138]&~m[139])|(~m[3]&m[136]&m[137]&~m[138]&~m[139])|(m[3]&~m[136]&~m[137]&m[138]&~m[139])|(~m[3]&m[136]&~m[137]&m[138]&~m[139])|(~m[3]&~m[136]&m[137]&m[138]&~m[139])|(m[3]&~m[136]&~m[137]&~m[138]&m[139])|(~m[3]&m[136]&~m[137]&~m[138]&m[139])|(~m[3]&~m[136]&m[137]&~m[138]&m[139])|(~m[3]&~m[136]&~m[137]&m[138]&m[139]))&BiasedRNG[178])|(((m[3]&m[136]&m[137]&~m[138]&~m[139])|(m[3]&m[136]&~m[137]&m[138]&~m[139])|(m[3]&~m[136]&m[137]&m[138]&~m[139])|(~m[3]&m[136]&m[137]&m[138]&~m[139])|(m[3]&m[136]&~m[137]&~m[138]&m[139])|(m[3]&~m[136]&m[137]&~m[138]&m[139])|(~m[3]&m[136]&m[137]&~m[138]&m[139])|(m[3]&~m[136]&~m[137]&m[138]&m[139])|(~m[3]&m[136]&~m[137]&m[138]&m[139])|(~m[3]&~m[136]&m[137]&m[138]&m[139]))&~BiasedRNG[178])|((m[3]&m[136]&m[137]&m[138]&~m[139])|(m[3]&m[136]&m[137]&~m[138]&m[139])|(m[3]&m[136]&~m[137]&m[138]&m[139])|(m[3]&~m[136]&m[137]&m[138]&m[139])|(~m[3]&m[136]&m[137]&m[138]&m[139])|(m[3]&m[136]&m[137]&m[138]&m[139]))):InitCond[309];
    m[35] = run?((((m[3]&m[140]&~m[141]&~m[142]&~m[143])|(m[3]&~m[140]&m[141]&~m[142]&~m[143])|(~m[3]&m[140]&m[141]&~m[142]&~m[143])|(m[3]&~m[140]&~m[141]&m[142]&~m[143])|(~m[3]&m[140]&~m[141]&m[142]&~m[143])|(~m[3]&~m[140]&m[141]&m[142]&~m[143])|(m[3]&~m[140]&~m[141]&~m[142]&m[143])|(~m[3]&m[140]&~m[141]&~m[142]&m[143])|(~m[3]&~m[140]&m[141]&~m[142]&m[143])|(~m[3]&~m[140]&~m[141]&m[142]&m[143]))&BiasedRNG[179])|(((m[3]&m[140]&m[141]&~m[142]&~m[143])|(m[3]&m[140]&~m[141]&m[142]&~m[143])|(m[3]&~m[140]&m[141]&m[142]&~m[143])|(~m[3]&m[140]&m[141]&m[142]&~m[143])|(m[3]&m[140]&~m[141]&~m[142]&m[143])|(m[3]&~m[140]&m[141]&~m[142]&m[143])|(~m[3]&m[140]&m[141]&~m[142]&m[143])|(m[3]&~m[140]&~m[141]&m[142]&m[143])|(~m[3]&m[140]&~m[141]&m[142]&m[143])|(~m[3]&~m[140]&m[141]&m[142]&m[143]))&~BiasedRNG[179])|((m[3]&m[140]&m[141]&m[142]&~m[143])|(m[3]&m[140]&m[141]&~m[142]&m[143])|(m[3]&m[140]&~m[141]&m[142]&m[143])|(m[3]&~m[140]&m[141]&m[142]&m[143])|(~m[3]&m[140]&m[141]&m[142]&m[143])|(m[3]&m[140]&m[141]&m[142]&m[143]))):InitCond[310];
    m[36] = run?((((m[4]&m[144]&~m[145]&~m[146]&~m[147])|(m[4]&~m[144]&m[145]&~m[146]&~m[147])|(~m[4]&m[144]&m[145]&~m[146]&~m[147])|(m[4]&~m[144]&~m[145]&m[146]&~m[147])|(~m[4]&m[144]&~m[145]&m[146]&~m[147])|(~m[4]&~m[144]&m[145]&m[146]&~m[147])|(m[4]&~m[144]&~m[145]&~m[146]&m[147])|(~m[4]&m[144]&~m[145]&~m[146]&m[147])|(~m[4]&~m[144]&m[145]&~m[146]&m[147])|(~m[4]&~m[144]&~m[145]&m[146]&m[147]))&BiasedRNG[180])|(((m[4]&m[144]&m[145]&~m[146]&~m[147])|(m[4]&m[144]&~m[145]&m[146]&~m[147])|(m[4]&~m[144]&m[145]&m[146]&~m[147])|(~m[4]&m[144]&m[145]&m[146]&~m[147])|(m[4]&m[144]&~m[145]&~m[146]&m[147])|(m[4]&~m[144]&m[145]&~m[146]&m[147])|(~m[4]&m[144]&m[145]&~m[146]&m[147])|(m[4]&~m[144]&~m[145]&m[146]&m[147])|(~m[4]&m[144]&~m[145]&m[146]&m[147])|(~m[4]&~m[144]&m[145]&m[146]&m[147]))&~BiasedRNG[180])|((m[4]&m[144]&m[145]&m[146]&~m[147])|(m[4]&m[144]&m[145]&~m[146]&m[147])|(m[4]&m[144]&~m[145]&m[146]&m[147])|(m[4]&~m[144]&m[145]&m[146]&m[147])|(~m[4]&m[144]&m[145]&m[146]&m[147])|(m[4]&m[144]&m[145]&m[146]&m[147]))):InitCond[311];
    m[37] = run?((((m[4]&m[148]&~m[149]&~m[150]&~m[151])|(m[4]&~m[148]&m[149]&~m[150]&~m[151])|(~m[4]&m[148]&m[149]&~m[150]&~m[151])|(m[4]&~m[148]&~m[149]&m[150]&~m[151])|(~m[4]&m[148]&~m[149]&m[150]&~m[151])|(~m[4]&~m[148]&m[149]&m[150]&~m[151])|(m[4]&~m[148]&~m[149]&~m[150]&m[151])|(~m[4]&m[148]&~m[149]&~m[150]&m[151])|(~m[4]&~m[148]&m[149]&~m[150]&m[151])|(~m[4]&~m[148]&~m[149]&m[150]&m[151]))&BiasedRNG[181])|(((m[4]&m[148]&m[149]&~m[150]&~m[151])|(m[4]&m[148]&~m[149]&m[150]&~m[151])|(m[4]&~m[148]&m[149]&m[150]&~m[151])|(~m[4]&m[148]&m[149]&m[150]&~m[151])|(m[4]&m[148]&~m[149]&~m[150]&m[151])|(m[4]&~m[148]&m[149]&~m[150]&m[151])|(~m[4]&m[148]&m[149]&~m[150]&m[151])|(m[4]&~m[148]&~m[149]&m[150]&m[151])|(~m[4]&m[148]&~m[149]&m[150]&m[151])|(~m[4]&~m[148]&m[149]&m[150]&m[151]))&~BiasedRNG[181])|((m[4]&m[148]&m[149]&m[150]&~m[151])|(m[4]&m[148]&m[149]&~m[150]&m[151])|(m[4]&m[148]&~m[149]&m[150]&m[151])|(m[4]&~m[148]&m[149]&m[150]&m[151])|(~m[4]&m[148]&m[149]&m[150]&m[151])|(m[4]&m[148]&m[149]&m[150]&m[151]))):InitCond[312];
    m[38] = run?((((m[4]&m[152]&~m[153]&~m[154]&~m[155])|(m[4]&~m[152]&m[153]&~m[154]&~m[155])|(~m[4]&m[152]&m[153]&~m[154]&~m[155])|(m[4]&~m[152]&~m[153]&m[154]&~m[155])|(~m[4]&m[152]&~m[153]&m[154]&~m[155])|(~m[4]&~m[152]&m[153]&m[154]&~m[155])|(m[4]&~m[152]&~m[153]&~m[154]&m[155])|(~m[4]&m[152]&~m[153]&~m[154]&m[155])|(~m[4]&~m[152]&m[153]&~m[154]&m[155])|(~m[4]&~m[152]&~m[153]&m[154]&m[155]))&BiasedRNG[182])|(((m[4]&m[152]&m[153]&~m[154]&~m[155])|(m[4]&m[152]&~m[153]&m[154]&~m[155])|(m[4]&~m[152]&m[153]&m[154]&~m[155])|(~m[4]&m[152]&m[153]&m[154]&~m[155])|(m[4]&m[152]&~m[153]&~m[154]&m[155])|(m[4]&~m[152]&m[153]&~m[154]&m[155])|(~m[4]&m[152]&m[153]&~m[154]&m[155])|(m[4]&~m[152]&~m[153]&m[154]&m[155])|(~m[4]&m[152]&~m[153]&m[154]&m[155])|(~m[4]&~m[152]&m[153]&m[154]&m[155]))&~BiasedRNG[182])|((m[4]&m[152]&m[153]&m[154]&~m[155])|(m[4]&m[152]&m[153]&~m[154]&m[155])|(m[4]&m[152]&~m[153]&m[154]&m[155])|(m[4]&~m[152]&m[153]&m[154]&m[155])|(~m[4]&m[152]&m[153]&m[154]&m[155])|(m[4]&m[152]&m[153]&m[154]&m[155]))):InitCond[313];
    m[39] = run?((((m[5]&m[156]&~m[157]&~m[158]&~m[159])|(m[5]&~m[156]&m[157]&~m[158]&~m[159])|(~m[5]&m[156]&m[157]&~m[158]&~m[159])|(m[5]&~m[156]&~m[157]&m[158]&~m[159])|(~m[5]&m[156]&~m[157]&m[158]&~m[159])|(~m[5]&~m[156]&m[157]&m[158]&~m[159])|(m[5]&~m[156]&~m[157]&~m[158]&m[159])|(~m[5]&m[156]&~m[157]&~m[158]&m[159])|(~m[5]&~m[156]&m[157]&~m[158]&m[159])|(~m[5]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[183])|(((m[5]&m[156]&m[157]&~m[158]&~m[159])|(m[5]&m[156]&~m[157]&m[158]&~m[159])|(m[5]&~m[156]&m[157]&m[158]&~m[159])|(~m[5]&m[156]&m[157]&m[158]&~m[159])|(m[5]&m[156]&~m[157]&~m[158]&m[159])|(m[5]&~m[156]&m[157]&~m[158]&m[159])|(~m[5]&m[156]&m[157]&~m[158]&m[159])|(m[5]&~m[156]&~m[157]&m[158]&m[159])|(~m[5]&m[156]&~m[157]&m[158]&m[159])|(~m[5]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[183])|((m[5]&m[156]&m[157]&m[158]&~m[159])|(m[5]&m[156]&m[157]&~m[158]&m[159])|(m[5]&m[156]&~m[157]&m[158]&m[159])|(m[5]&~m[156]&m[157]&m[158]&m[159])|(~m[5]&m[156]&m[157]&m[158]&m[159])|(m[5]&m[156]&m[157]&m[158]&m[159]))):InitCond[314];
    m[40] = run?((((m[5]&m[160]&~m[161]&~m[162]&~m[163])|(m[5]&~m[160]&m[161]&~m[162]&~m[163])|(~m[5]&m[160]&m[161]&~m[162]&~m[163])|(m[5]&~m[160]&~m[161]&m[162]&~m[163])|(~m[5]&m[160]&~m[161]&m[162]&~m[163])|(~m[5]&~m[160]&m[161]&m[162]&~m[163])|(m[5]&~m[160]&~m[161]&~m[162]&m[163])|(~m[5]&m[160]&~m[161]&~m[162]&m[163])|(~m[5]&~m[160]&m[161]&~m[162]&m[163])|(~m[5]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[184])|(((m[5]&m[160]&m[161]&~m[162]&~m[163])|(m[5]&m[160]&~m[161]&m[162]&~m[163])|(m[5]&~m[160]&m[161]&m[162]&~m[163])|(~m[5]&m[160]&m[161]&m[162]&~m[163])|(m[5]&m[160]&~m[161]&~m[162]&m[163])|(m[5]&~m[160]&m[161]&~m[162]&m[163])|(~m[5]&m[160]&m[161]&~m[162]&m[163])|(m[5]&~m[160]&~m[161]&m[162]&m[163])|(~m[5]&m[160]&~m[161]&m[162]&m[163])|(~m[5]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[184])|((m[5]&m[160]&m[161]&m[162]&~m[163])|(m[5]&m[160]&m[161]&~m[162]&m[163])|(m[5]&m[160]&~m[161]&m[162]&m[163])|(m[5]&~m[160]&m[161]&m[162]&m[163])|(~m[5]&m[160]&m[161]&m[162]&m[163])|(m[5]&m[160]&m[161]&m[162]&m[163]))):InitCond[315];
    m[41] = run?((((m[5]&m[164]&~m[165]&~m[166]&~m[167])|(m[5]&~m[164]&m[165]&~m[166]&~m[167])|(~m[5]&m[164]&m[165]&~m[166]&~m[167])|(m[5]&~m[164]&~m[165]&m[166]&~m[167])|(~m[5]&m[164]&~m[165]&m[166]&~m[167])|(~m[5]&~m[164]&m[165]&m[166]&~m[167])|(m[5]&~m[164]&~m[165]&~m[166]&m[167])|(~m[5]&m[164]&~m[165]&~m[166]&m[167])|(~m[5]&~m[164]&m[165]&~m[166]&m[167])|(~m[5]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[185])|(((m[5]&m[164]&m[165]&~m[166]&~m[167])|(m[5]&m[164]&~m[165]&m[166]&~m[167])|(m[5]&~m[164]&m[165]&m[166]&~m[167])|(~m[5]&m[164]&m[165]&m[166]&~m[167])|(m[5]&m[164]&~m[165]&~m[166]&m[167])|(m[5]&~m[164]&m[165]&~m[166]&m[167])|(~m[5]&m[164]&m[165]&~m[166]&m[167])|(m[5]&~m[164]&~m[165]&m[166]&m[167])|(~m[5]&m[164]&~m[165]&m[166]&m[167])|(~m[5]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[185])|((m[5]&m[164]&m[165]&m[166]&~m[167])|(m[5]&m[164]&m[165]&~m[166]&m[167])|(m[5]&m[164]&~m[165]&m[166]&m[167])|(m[5]&~m[164]&m[165]&m[166]&m[167])|(~m[5]&m[164]&m[165]&m[166]&m[167])|(m[5]&m[164]&m[165]&m[166]&m[167]))):InitCond[316];
    m[42] = run?((((m[6]&m[168]&~m[169]&~m[170]&~m[171])|(m[6]&~m[168]&m[169]&~m[170]&~m[171])|(~m[6]&m[168]&m[169]&~m[170]&~m[171])|(m[6]&~m[168]&~m[169]&m[170]&~m[171])|(~m[6]&m[168]&~m[169]&m[170]&~m[171])|(~m[6]&~m[168]&m[169]&m[170]&~m[171])|(m[6]&~m[168]&~m[169]&~m[170]&m[171])|(~m[6]&m[168]&~m[169]&~m[170]&m[171])|(~m[6]&~m[168]&m[169]&~m[170]&m[171])|(~m[6]&~m[168]&~m[169]&m[170]&m[171]))&BiasedRNG[186])|(((m[6]&m[168]&m[169]&~m[170]&~m[171])|(m[6]&m[168]&~m[169]&m[170]&~m[171])|(m[6]&~m[168]&m[169]&m[170]&~m[171])|(~m[6]&m[168]&m[169]&m[170]&~m[171])|(m[6]&m[168]&~m[169]&~m[170]&m[171])|(m[6]&~m[168]&m[169]&~m[170]&m[171])|(~m[6]&m[168]&m[169]&~m[170]&m[171])|(m[6]&~m[168]&~m[169]&m[170]&m[171])|(~m[6]&m[168]&~m[169]&m[170]&m[171])|(~m[6]&~m[168]&m[169]&m[170]&m[171]))&~BiasedRNG[186])|((m[6]&m[168]&m[169]&m[170]&~m[171])|(m[6]&m[168]&m[169]&~m[170]&m[171])|(m[6]&m[168]&~m[169]&m[170]&m[171])|(m[6]&~m[168]&m[169]&m[170]&m[171])|(~m[6]&m[168]&m[169]&m[170]&m[171])|(m[6]&m[168]&m[169]&m[170]&m[171]))):InitCond[317];
    m[43] = run?((((m[6]&m[172]&~m[173]&~m[174]&~m[175])|(m[6]&~m[172]&m[173]&~m[174]&~m[175])|(~m[6]&m[172]&m[173]&~m[174]&~m[175])|(m[6]&~m[172]&~m[173]&m[174]&~m[175])|(~m[6]&m[172]&~m[173]&m[174]&~m[175])|(~m[6]&~m[172]&m[173]&m[174]&~m[175])|(m[6]&~m[172]&~m[173]&~m[174]&m[175])|(~m[6]&m[172]&~m[173]&~m[174]&m[175])|(~m[6]&~m[172]&m[173]&~m[174]&m[175])|(~m[6]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[187])|(((m[6]&m[172]&m[173]&~m[174]&~m[175])|(m[6]&m[172]&~m[173]&m[174]&~m[175])|(m[6]&~m[172]&m[173]&m[174]&~m[175])|(~m[6]&m[172]&m[173]&m[174]&~m[175])|(m[6]&m[172]&~m[173]&~m[174]&m[175])|(m[6]&~m[172]&m[173]&~m[174]&m[175])|(~m[6]&m[172]&m[173]&~m[174]&m[175])|(m[6]&~m[172]&~m[173]&m[174]&m[175])|(~m[6]&m[172]&~m[173]&m[174]&m[175])|(~m[6]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[187])|((m[6]&m[172]&m[173]&m[174]&~m[175])|(m[6]&m[172]&m[173]&~m[174]&m[175])|(m[6]&m[172]&~m[173]&m[174]&m[175])|(m[6]&~m[172]&m[173]&m[174]&m[175])|(~m[6]&m[172]&m[173]&m[174]&m[175])|(m[6]&m[172]&m[173]&m[174]&m[175]))):InitCond[318];
    m[44] = run?((((m[6]&m[176]&~m[177]&~m[178]&~m[179])|(m[6]&~m[176]&m[177]&~m[178]&~m[179])|(~m[6]&m[176]&m[177]&~m[178]&~m[179])|(m[6]&~m[176]&~m[177]&m[178]&~m[179])|(~m[6]&m[176]&~m[177]&m[178]&~m[179])|(~m[6]&~m[176]&m[177]&m[178]&~m[179])|(m[6]&~m[176]&~m[177]&~m[178]&m[179])|(~m[6]&m[176]&~m[177]&~m[178]&m[179])|(~m[6]&~m[176]&m[177]&~m[178]&m[179])|(~m[6]&~m[176]&~m[177]&m[178]&m[179]))&BiasedRNG[188])|(((m[6]&m[176]&m[177]&~m[178]&~m[179])|(m[6]&m[176]&~m[177]&m[178]&~m[179])|(m[6]&~m[176]&m[177]&m[178]&~m[179])|(~m[6]&m[176]&m[177]&m[178]&~m[179])|(m[6]&m[176]&~m[177]&~m[178]&m[179])|(m[6]&~m[176]&m[177]&~m[178]&m[179])|(~m[6]&m[176]&m[177]&~m[178]&m[179])|(m[6]&~m[176]&~m[177]&m[178]&m[179])|(~m[6]&m[176]&~m[177]&m[178]&m[179])|(~m[6]&~m[176]&m[177]&m[178]&m[179]))&~BiasedRNG[188])|((m[6]&m[176]&m[177]&m[178]&~m[179])|(m[6]&m[176]&m[177]&~m[178]&m[179])|(m[6]&m[176]&~m[177]&m[178]&m[179])|(m[6]&~m[176]&m[177]&m[178]&m[179])|(~m[6]&m[176]&m[177]&m[178]&m[179])|(m[6]&m[176]&m[177]&m[178]&m[179]))):InitCond[319];
    m[45] = run?((((m[7]&m[180]&~m[181]&~m[182]&~m[183])|(m[7]&~m[180]&m[181]&~m[182]&~m[183])|(~m[7]&m[180]&m[181]&~m[182]&~m[183])|(m[7]&~m[180]&~m[181]&m[182]&~m[183])|(~m[7]&m[180]&~m[181]&m[182]&~m[183])|(~m[7]&~m[180]&m[181]&m[182]&~m[183])|(m[7]&~m[180]&~m[181]&~m[182]&m[183])|(~m[7]&m[180]&~m[181]&~m[182]&m[183])|(~m[7]&~m[180]&m[181]&~m[182]&m[183])|(~m[7]&~m[180]&~m[181]&m[182]&m[183]))&BiasedRNG[189])|(((m[7]&m[180]&m[181]&~m[182]&~m[183])|(m[7]&m[180]&~m[181]&m[182]&~m[183])|(m[7]&~m[180]&m[181]&m[182]&~m[183])|(~m[7]&m[180]&m[181]&m[182]&~m[183])|(m[7]&m[180]&~m[181]&~m[182]&m[183])|(m[7]&~m[180]&m[181]&~m[182]&m[183])|(~m[7]&m[180]&m[181]&~m[182]&m[183])|(m[7]&~m[180]&~m[181]&m[182]&m[183])|(~m[7]&m[180]&~m[181]&m[182]&m[183])|(~m[7]&~m[180]&m[181]&m[182]&m[183]))&~BiasedRNG[189])|((m[7]&m[180]&m[181]&m[182]&~m[183])|(m[7]&m[180]&m[181]&~m[182]&m[183])|(m[7]&m[180]&~m[181]&m[182]&m[183])|(m[7]&~m[180]&m[181]&m[182]&m[183])|(~m[7]&m[180]&m[181]&m[182]&m[183])|(m[7]&m[180]&m[181]&m[182]&m[183]))):InitCond[320];
    m[46] = run?((((m[7]&m[184]&~m[185]&~m[186]&~m[187])|(m[7]&~m[184]&m[185]&~m[186]&~m[187])|(~m[7]&m[184]&m[185]&~m[186]&~m[187])|(m[7]&~m[184]&~m[185]&m[186]&~m[187])|(~m[7]&m[184]&~m[185]&m[186]&~m[187])|(~m[7]&~m[184]&m[185]&m[186]&~m[187])|(m[7]&~m[184]&~m[185]&~m[186]&m[187])|(~m[7]&m[184]&~m[185]&~m[186]&m[187])|(~m[7]&~m[184]&m[185]&~m[186]&m[187])|(~m[7]&~m[184]&~m[185]&m[186]&m[187]))&BiasedRNG[190])|(((m[7]&m[184]&m[185]&~m[186]&~m[187])|(m[7]&m[184]&~m[185]&m[186]&~m[187])|(m[7]&~m[184]&m[185]&m[186]&~m[187])|(~m[7]&m[184]&m[185]&m[186]&~m[187])|(m[7]&m[184]&~m[185]&~m[186]&m[187])|(m[7]&~m[184]&m[185]&~m[186]&m[187])|(~m[7]&m[184]&m[185]&~m[186]&m[187])|(m[7]&~m[184]&~m[185]&m[186]&m[187])|(~m[7]&m[184]&~m[185]&m[186]&m[187])|(~m[7]&~m[184]&m[185]&m[186]&m[187]))&~BiasedRNG[190])|((m[7]&m[184]&m[185]&m[186]&~m[187])|(m[7]&m[184]&m[185]&~m[186]&m[187])|(m[7]&m[184]&~m[185]&m[186]&m[187])|(m[7]&~m[184]&m[185]&m[186]&m[187])|(~m[7]&m[184]&m[185]&m[186]&m[187])|(m[7]&m[184]&m[185]&m[186]&m[187]))):InitCond[321];
    m[47] = run?((((m[7]&m[188]&~m[189]&~m[190]&~m[191])|(m[7]&~m[188]&m[189]&~m[190]&~m[191])|(~m[7]&m[188]&m[189]&~m[190]&~m[191])|(m[7]&~m[188]&~m[189]&m[190]&~m[191])|(~m[7]&m[188]&~m[189]&m[190]&~m[191])|(~m[7]&~m[188]&m[189]&m[190]&~m[191])|(m[7]&~m[188]&~m[189]&~m[190]&m[191])|(~m[7]&m[188]&~m[189]&~m[190]&m[191])|(~m[7]&~m[188]&m[189]&~m[190]&m[191])|(~m[7]&~m[188]&~m[189]&m[190]&m[191]))&BiasedRNG[191])|(((m[7]&m[188]&m[189]&~m[190]&~m[191])|(m[7]&m[188]&~m[189]&m[190]&~m[191])|(m[7]&~m[188]&m[189]&m[190]&~m[191])|(~m[7]&m[188]&m[189]&m[190]&~m[191])|(m[7]&m[188]&~m[189]&~m[190]&m[191])|(m[7]&~m[188]&m[189]&~m[190]&m[191])|(~m[7]&m[188]&m[189]&~m[190]&m[191])|(m[7]&~m[188]&~m[189]&m[190]&m[191])|(~m[7]&m[188]&~m[189]&m[190]&m[191])|(~m[7]&~m[188]&m[189]&m[190]&m[191]))&~BiasedRNG[191])|((m[7]&m[188]&m[189]&m[190]&~m[191])|(m[7]&m[188]&m[189]&~m[190]&m[191])|(m[7]&m[188]&~m[189]&m[190]&m[191])|(m[7]&~m[188]&m[189]&m[190]&m[191])|(~m[7]&m[188]&m[189]&m[190]&m[191])|(m[7]&m[188]&m[189]&m[190]&m[191]))):InitCond[322];
    m[48] = run?((((m[8]&m[192]&~m[193]&~m[194]&~m[195])|(m[8]&~m[192]&m[193]&~m[194]&~m[195])|(~m[8]&m[192]&m[193]&~m[194]&~m[195])|(m[8]&~m[192]&~m[193]&m[194]&~m[195])|(~m[8]&m[192]&~m[193]&m[194]&~m[195])|(~m[8]&~m[192]&m[193]&m[194]&~m[195])|(m[8]&~m[192]&~m[193]&~m[194]&m[195])|(~m[8]&m[192]&~m[193]&~m[194]&m[195])|(~m[8]&~m[192]&m[193]&~m[194]&m[195])|(~m[8]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[192])|(((m[8]&m[192]&m[193]&~m[194]&~m[195])|(m[8]&m[192]&~m[193]&m[194]&~m[195])|(m[8]&~m[192]&m[193]&m[194]&~m[195])|(~m[8]&m[192]&m[193]&m[194]&~m[195])|(m[8]&m[192]&~m[193]&~m[194]&m[195])|(m[8]&~m[192]&m[193]&~m[194]&m[195])|(~m[8]&m[192]&m[193]&~m[194]&m[195])|(m[8]&~m[192]&~m[193]&m[194]&m[195])|(~m[8]&m[192]&~m[193]&m[194]&m[195])|(~m[8]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[192])|((m[8]&m[192]&m[193]&m[194]&~m[195])|(m[8]&m[192]&m[193]&~m[194]&m[195])|(m[8]&m[192]&~m[193]&m[194]&m[195])|(m[8]&~m[192]&m[193]&m[194]&m[195])|(~m[8]&m[192]&m[193]&m[194]&m[195])|(m[8]&m[192]&m[193]&m[194]&m[195]))):InitCond[323];
    m[49] = run?((((m[8]&m[196]&~m[197]&~m[198]&~m[199])|(m[8]&~m[196]&m[197]&~m[198]&~m[199])|(~m[8]&m[196]&m[197]&~m[198]&~m[199])|(m[8]&~m[196]&~m[197]&m[198]&~m[199])|(~m[8]&m[196]&~m[197]&m[198]&~m[199])|(~m[8]&~m[196]&m[197]&m[198]&~m[199])|(m[8]&~m[196]&~m[197]&~m[198]&m[199])|(~m[8]&m[196]&~m[197]&~m[198]&m[199])|(~m[8]&~m[196]&m[197]&~m[198]&m[199])|(~m[8]&~m[196]&~m[197]&m[198]&m[199]))&BiasedRNG[193])|(((m[8]&m[196]&m[197]&~m[198]&~m[199])|(m[8]&m[196]&~m[197]&m[198]&~m[199])|(m[8]&~m[196]&m[197]&m[198]&~m[199])|(~m[8]&m[196]&m[197]&m[198]&~m[199])|(m[8]&m[196]&~m[197]&~m[198]&m[199])|(m[8]&~m[196]&m[197]&~m[198]&m[199])|(~m[8]&m[196]&m[197]&~m[198]&m[199])|(m[8]&~m[196]&~m[197]&m[198]&m[199])|(~m[8]&m[196]&~m[197]&m[198]&m[199])|(~m[8]&~m[196]&m[197]&m[198]&m[199]))&~BiasedRNG[193])|((m[8]&m[196]&m[197]&m[198]&~m[199])|(m[8]&m[196]&m[197]&~m[198]&m[199])|(m[8]&m[196]&~m[197]&m[198]&m[199])|(m[8]&~m[196]&m[197]&m[198]&m[199])|(~m[8]&m[196]&m[197]&m[198]&m[199])|(m[8]&m[196]&m[197]&m[198]&m[199]))):InitCond[324];
    m[50] = run?((((m[8]&m[200]&~m[201]&~m[202]&~m[203])|(m[8]&~m[200]&m[201]&~m[202]&~m[203])|(~m[8]&m[200]&m[201]&~m[202]&~m[203])|(m[8]&~m[200]&~m[201]&m[202]&~m[203])|(~m[8]&m[200]&~m[201]&m[202]&~m[203])|(~m[8]&~m[200]&m[201]&m[202]&~m[203])|(m[8]&~m[200]&~m[201]&~m[202]&m[203])|(~m[8]&m[200]&~m[201]&~m[202]&m[203])|(~m[8]&~m[200]&m[201]&~m[202]&m[203])|(~m[8]&~m[200]&~m[201]&m[202]&m[203]))&BiasedRNG[194])|(((m[8]&m[200]&m[201]&~m[202]&~m[203])|(m[8]&m[200]&~m[201]&m[202]&~m[203])|(m[8]&~m[200]&m[201]&m[202]&~m[203])|(~m[8]&m[200]&m[201]&m[202]&~m[203])|(m[8]&m[200]&~m[201]&~m[202]&m[203])|(m[8]&~m[200]&m[201]&~m[202]&m[203])|(~m[8]&m[200]&m[201]&~m[202]&m[203])|(m[8]&~m[200]&~m[201]&m[202]&m[203])|(~m[8]&m[200]&~m[201]&m[202]&m[203])|(~m[8]&~m[200]&m[201]&m[202]&m[203]))&~BiasedRNG[194])|((m[8]&m[200]&m[201]&m[202]&~m[203])|(m[8]&m[200]&m[201]&~m[202]&m[203])|(m[8]&m[200]&~m[201]&m[202]&m[203])|(m[8]&~m[200]&m[201]&m[202]&m[203])|(~m[8]&m[200]&m[201]&m[202]&m[203])|(m[8]&m[200]&m[201]&m[202]&m[203]))):InitCond[325];
    m[51] = run?((((m[9]&m[204]&~m[205]&~m[206]&~m[207])|(m[9]&~m[204]&m[205]&~m[206]&~m[207])|(~m[9]&m[204]&m[205]&~m[206]&~m[207])|(m[9]&~m[204]&~m[205]&m[206]&~m[207])|(~m[9]&m[204]&~m[205]&m[206]&~m[207])|(~m[9]&~m[204]&m[205]&m[206]&~m[207])|(m[9]&~m[204]&~m[205]&~m[206]&m[207])|(~m[9]&m[204]&~m[205]&~m[206]&m[207])|(~m[9]&~m[204]&m[205]&~m[206]&m[207])|(~m[9]&~m[204]&~m[205]&m[206]&m[207]))&BiasedRNG[195])|(((m[9]&m[204]&m[205]&~m[206]&~m[207])|(m[9]&m[204]&~m[205]&m[206]&~m[207])|(m[9]&~m[204]&m[205]&m[206]&~m[207])|(~m[9]&m[204]&m[205]&m[206]&~m[207])|(m[9]&m[204]&~m[205]&~m[206]&m[207])|(m[9]&~m[204]&m[205]&~m[206]&m[207])|(~m[9]&m[204]&m[205]&~m[206]&m[207])|(m[9]&~m[204]&~m[205]&m[206]&m[207])|(~m[9]&m[204]&~m[205]&m[206]&m[207])|(~m[9]&~m[204]&m[205]&m[206]&m[207]))&~BiasedRNG[195])|((m[9]&m[204]&m[205]&m[206]&~m[207])|(m[9]&m[204]&m[205]&~m[206]&m[207])|(m[9]&m[204]&~m[205]&m[206]&m[207])|(m[9]&~m[204]&m[205]&m[206]&m[207])|(~m[9]&m[204]&m[205]&m[206]&m[207])|(m[9]&m[204]&m[205]&m[206]&m[207]))):InitCond[326];
    m[52] = run?((((m[9]&m[208]&~m[209]&~m[210]&~m[211])|(m[9]&~m[208]&m[209]&~m[210]&~m[211])|(~m[9]&m[208]&m[209]&~m[210]&~m[211])|(m[9]&~m[208]&~m[209]&m[210]&~m[211])|(~m[9]&m[208]&~m[209]&m[210]&~m[211])|(~m[9]&~m[208]&m[209]&m[210]&~m[211])|(m[9]&~m[208]&~m[209]&~m[210]&m[211])|(~m[9]&m[208]&~m[209]&~m[210]&m[211])|(~m[9]&~m[208]&m[209]&~m[210]&m[211])|(~m[9]&~m[208]&~m[209]&m[210]&m[211]))&BiasedRNG[196])|(((m[9]&m[208]&m[209]&~m[210]&~m[211])|(m[9]&m[208]&~m[209]&m[210]&~m[211])|(m[9]&~m[208]&m[209]&m[210]&~m[211])|(~m[9]&m[208]&m[209]&m[210]&~m[211])|(m[9]&m[208]&~m[209]&~m[210]&m[211])|(m[9]&~m[208]&m[209]&~m[210]&m[211])|(~m[9]&m[208]&m[209]&~m[210]&m[211])|(m[9]&~m[208]&~m[209]&m[210]&m[211])|(~m[9]&m[208]&~m[209]&m[210]&m[211])|(~m[9]&~m[208]&m[209]&m[210]&m[211]))&~BiasedRNG[196])|((m[9]&m[208]&m[209]&m[210]&~m[211])|(m[9]&m[208]&m[209]&~m[210]&m[211])|(m[9]&m[208]&~m[209]&m[210]&m[211])|(m[9]&~m[208]&m[209]&m[210]&m[211])|(~m[9]&m[208]&m[209]&m[210]&m[211])|(m[9]&m[208]&m[209]&m[210]&m[211]))):InitCond[327];
    m[53] = run?((((m[9]&m[212]&~m[213]&~m[214]&~m[215])|(m[9]&~m[212]&m[213]&~m[214]&~m[215])|(~m[9]&m[212]&m[213]&~m[214]&~m[215])|(m[9]&~m[212]&~m[213]&m[214]&~m[215])|(~m[9]&m[212]&~m[213]&m[214]&~m[215])|(~m[9]&~m[212]&m[213]&m[214]&~m[215])|(m[9]&~m[212]&~m[213]&~m[214]&m[215])|(~m[9]&m[212]&~m[213]&~m[214]&m[215])|(~m[9]&~m[212]&m[213]&~m[214]&m[215])|(~m[9]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[197])|(((m[9]&m[212]&m[213]&~m[214]&~m[215])|(m[9]&m[212]&~m[213]&m[214]&~m[215])|(m[9]&~m[212]&m[213]&m[214]&~m[215])|(~m[9]&m[212]&m[213]&m[214]&~m[215])|(m[9]&m[212]&~m[213]&~m[214]&m[215])|(m[9]&~m[212]&m[213]&~m[214]&m[215])|(~m[9]&m[212]&m[213]&~m[214]&m[215])|(m[9]&~m[212]&~m[213]&m[214]&m[215])|(~m[9]&m[212]&~m[213]&m[214]&m[215])|(~m[9]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[197])|((m[9]&m[212]&m[213]&m[214]&~m[215])|(m[9]&m[212]&m[213]&~m[214]&m[215])|(m[9]&m[212]&~m[213]&m[214]&m[215])|(m[9]&~m[212]&m[213]&m[214]&m[215])|(~m[9]&m[212]&m[213]&m[214]&m[215])|(m[9]&m[212]&m[213]&m[214]&m[215]))):InitCond[328];
    m[54] = run?((((m[10]&m[216]&~m[217]&~m[218]&~m[219])|(m[10]&~m[216]&m[217]&~m[218]&~m[219])|(~m[10]&m[216]&m[217]&~m[218]&~m[219])|(m[10]&~m[216]&~m[217]&m[218]&~m[219])|(~m[10]&m[216]&~m[217]&m[218]&~m[219])|(~m[10]&~m[216]&m[217]&m[218]&~m[219])|(m[10]&~m[216]&~m[217]&~m[218]&m[219])|(~m[10]&m[216]&~m[217]&~m[218]&m[219])|(~m[10]&~m[216]&m[217]&~m[218]&m[219])|(~m[10]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[198])|(((m[10]&m[216]&m[217]&~m[218]&~m[219])|(m[10]&m[216]&~m[217]&m[218]&~m[219])|(m[10]&~m[216]&m[217]&m[218]&~m[219])|(~m[10]&m[216]&m[217]&m[218]&~m[219])|(m[10]&m[216]&~m[217]&~m[218]&m[219])|(m[10]&~m[216]&m[217]&~m[218]&m[219])|(~m[10]&m[216]&m[217]&~m[218]&m[219])|(m[10]&~m[216]&~m[217]&m[218]&m[219])|(~m[10]&m[216]&~m[217]&m[218]&m[219])|(~m[10]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[198])|((m[10]&m[216]&m[217]&m[218]&~m[219])|(m[10]&m[216]&m[217]&~m[218]&m[219])|(m[10]&m[216]&~m[217]&m[218]&m[219])|(m[10]&~m[216]&m[217]&m[218]&m[219])|(~m[10]&m[216]&m[217]&m[218]&m[219])|(m[10]&m[216]&m[217]&m[218]&m[219]))):InitCond[329];
    m[55] = run?((((m[10]&m[220]&~m[221]&~m[222]&~m[223])|(m[10]&~m[220]&m[221]&~m[222]&~m[223])|(~m[10]&m[220]&m[221]&~m[222]&~m[223])|(m[10]&~m[220]&~m[221]&m[222]&~m[223])|(~m[10]&m[220]&~m[221]&m[222]&~m[223])|(~m[10]&~m[220]&m[221]&m[222]&~m[223])|(m[10]&~m[220]&~m[221]&~m[222]&m[223])|(~m[10]&m[220]&~m[221]&~m[222]&m[223])|(~m[10]&~m[220]&m[221]&~m[222]&m[223])|(~m[10]&~m[220]&~m[221]&m[222]&m[223]))&BiasedRNG[199])|(((m[10]&m[220]&m[221]&~m[222]&~m[223])|(m[10]&m[220]&~m[221]&m[222]&~m[223])|(m[10]&~m[220]&m[221]&m[222]&~m[223])|(~m[10]&m[220]&m[221]&m[222]&~m[223])|(m[10]&m[220]&~m[221]&~m[222]&m[223])|(m[10]&~m[220]&m[221]&~m[222]&m[223])|(~m[10]&m[220]&m[221]&~m[222]&m[223])|(m[10]&~m[220]&~m[221]&m[222]&m[223])|(~m[10]&m[220]&~m[221]&m[222]&m[223])|(~m[10]&~m[220]&m[221]&m[222]&m[223]))&~BiasedRNG[199])|((m[10]&m[220]&m[221]&m[222]&~m[223])|(m[10]&m[220]&m[221]&~m[222]&m[223])|(m[10]&m[220]&~m[221]&m[222]&m[223])|(m[10]&~m[220]&m[221]&m[222]&m[223])|(~m[10]&m[220]&m[221]&m[222]&m[223])|(m[10]&m[220]&m[221]&m[222]&m[223]))):InitCond[330];
    m[56] = run?((((m[10]&m[224]&~m[225]&~m[226]&~m[227])|(m[10]&~m[224]&m[225]&~m[226]&~m[227])|(~m[10]&m[224]&m[225]&~m[226]&~m[227])|(m[10]&~m[224]&~m[225]&m[226]&~m[227])|(~m[10]&m[224]&~m[225]&m[226]&~m[227])|(~m[10]&~m[224]&m[225]&m[226]&~m[227])|(m[10]&~m[224]&~m[225]&~m[226]&m[227])|(~m[10]&m[224]&~m[225]&~m[226]&m[227])|(~m[10]&~m[224]&m[225]&~m[226]&m[227])|(~m[10]&~m[224]&~m[225]&m[226]&m[227]))&BiasedRNG[200])|(((m[10]&m[224]&m[225]&~m[226]&~m[227])|(m[10]&m[224]&~m[225]&m[226]&~m[227])|(m[10]&~m[224]&m[225]&m[226]&~m[227])|(~m[10]&m[224]&m[225]&m[226]&~m[227])|(m[10]&m[224]&~m[225]&~m[226]&m[227])|(m[10]&~m[224]&m[225]&~m[226]&m[227])|(~m[10]&m[224]&m[225]&~m[226]&m[227])|(m[10]&~m[224]&~m[225]&m[226]&m[227])|(~m[10]&m[224]&~m[225]&m[226]&m[227])|(~m[10]&~m[224]&m[225]&m[226]&m[227]))&~BiasedRNG[200])|((m[10]&m[224]&m[225]&m[226]&~m[227])|(m[10]&m[224]&m[225]&~m[226]&m[227])|(m[10]&m[224]&~m[225]&m[226]&m[227])|(m[10]&~m[224]&m[225]&m[226]&m[227])|(~m[10]&m[224]&m[225]&m[226]&m[227])|(m[10]&m[224]&m[225]&m[226]&m[227]))):InitCond[331];
    m[57] = run?((((m[11]&m[228]&~m[229]&~m[230]&~m[231])|(m[11]&~m[228]&m[229]&~m[230]&~m[231])|(~m[11]&m[228]&m[229]&~m[230]&~m[231])|(m[11]&~m[228]&~m[229]&m[230]&~m[231])|(~m[11]&m[228]&~m[229]&m[230]&~m[231])|(~m[11]&~m[228]&m[229]&m[230]&~m[231])|(m[11]&~m[228]&~m[229]&~m[230]&m[231])|(~m[11]&m[228]&~m[229]&~m[230]&m[231])|(~m[11]&~m[228]&m[229]&~m[230]&m[231])|(~m[11]&~m[228]&~m[229]&m[230]&m[231]))&BiasedRNG[201])|(((m[11]&m[228]&m[229]&~m[230]&~m[231])|(m[11]&m[228]&~m[229]&m[230]&~m[231])|(m[11]&~m[228]&m[229]&m[230]&~m[231])|(~m[11]&m[228]&m[229]&m[230]&~m[231])|(m[11]&m[228]&~m[229]&~m[230]&m[231])|(m[11]&~m[228]&m[229]&~m[230]&m[231])|(~m[11]&m[228]&m[229]&~m[230]&m[231])|(m[11]&~m[228]&~m[229]&m[230]&m[231])|(~m[11]&m[228]&~m[229]&m[230]&m[231])|(~m[11]&~m[228]&m[229]&m[230]&m[231]))&~BiasedRNG[201])|((m[11]&m[228]&m[229]&m[230]&~m[231])|(m[11]&m[228]&m[229]&~m[230]&m[231])|(m[11]&m[228]&~m[229]&m[230]&m[231])|(m[11]&~m[228]&m[229]&m[230]&m[231])|(~m[11]&m[228]&m[229]&m[230]&m[231])|(m[11]&m[228]&m[229]&m[230]&m[231]))):InitCond[332];
    m[58] = run?((((m[11]&m[232]&~m[233]&~m[234]&~m[235])|(m[11]&~m[232]&m[233]&~m[234]&~m[235])|(~m[11]&m[232]&m[233]&~m[234]&~m[235])|(m[11]&~m[232]&~m[233]&m[234]&~m[235])|(~m[11]&m[232]&~m[233]&m[234]&~m[235])|(~m[11]&~m[232]&m[233]&m[234]&~m[235])|(m[11]&~m[232]&~m[233]&~m[234]&m[235])|(~m[11]&m[232]&~m[233]&~m[234]&m[235])|(~m[11]&~m[232]&m[233]&~m[234]&m[235])|(~m[11]&~m[232]&~m[233]&m[234]&m[235]))&BiasedRNG[202])|(((m[11]&m[232]&m[233]&~m[234]&~m[235])|(m[11]&m[232]&~m[233]&m[234]&~m[235])|(m[11]&~m[232]&m[233]&m[234]&~m[235])|(~m[11]&m[232]&m[233]&m[234]&~m[235])|(m[11]&m[232]&~m[233]&~m[234]&m[235])|(m[11]&~m[232]&m[233]&~m[234]&m[235])|(~m[11]&m[232]&m[233]&~m[234]&m[235])|(m[11]&~m[232]&~m[233]&m[234]&m[235])|(~m[11]&m[232]&~m[233]&m[234]&m[235])|(~m[11]&~m[232]&m[233]&m[234]&m[235]))&~BiasedRNG[202])|((m[11]&m[232]&m[233]&m[234]&~m[235])|(m[11]&m[232]&m[233]&~m[234]&m[235])|(m[11]&m[232]&~m[233]&m[234]&m[235])|(m[11]&~m[232]&m[233]&m[234]&m[235])|(~m[11]&m[232]&m[233]&m[234]&m[235])|(m[11]&m[232]&m[233]&m[234]&m[235]))):InitCond[333];
    m[59] = run?((((m[11]&m[236]&~m[237]&~m[238]&~m[239])|(m[11]&~m[236]&m[237]&~m[238]&~m[239])|(~m[11]&m[236]&m[237]&~m[238]&~m[239])|(m[11]&~m[236]&~m[237]&m[238]&~m[239])|(~m[11]&m[236]&~m[237]&m[238]&~m[239])|(~m[11]&~m[236]&m[237]&m[238]&~m[239])|(m[11]&~m[236]&~m[237]&~m[238]&m[239])|(~m[11]&m[236]&~m[237]&~m[238]&m[239])|(~m[11]&~m[236]&m[237]&~m[238]&m[239])|(~m[11]&~m[236]&~m[237]&m[238]&m[239]))&BiasedRNG[203])|(((m[11]&m[236]&m[237]&~m[238]&~m[239])|(m[11]&m[236]&~m[237]&m[238]&~m[239])|(m[11]&~m[236]&m[237]&m[238]&~m[239])|(~m[11]&m[236]&m[237]&m[238]&~m[239])|(m[11]&m[236]&~m[237]&~m[238]&m[239])|(m[11]&~m[236]&m[237]&~m[238]&m[239])|(~m[11]&m[236]&m[237]&~m[238]&m[239])|(m[11]&~m[236]&~m[237]&m[238]&m[239])|(~m[11]&m[236]&~m[237]&m[238]&m[239])|(~m[11]&~m[236]&m[237]&m[238]&m[239]))&~BiasedRNG[203])|((m[11]&m[236]&m[237]&m[238]&~m[239])|(m[11]&m[236]&m[237]&~m[238]&m[239])|(m[11]&m[236]&~m[237]&m[238]&m[239])|(m[11]&~m[236]&m[237]&m[238]&m[239])|(~m[11]&m[236]&m[237]&m[238]&m[239])|(m[11]&m[236]&m[237]&m[238]&m[239]))):InitCond[334];
    m[60] = run?((((m[12]&m[240]&~m[241]&~m[242]&~m[243])|(m[12]&~m[240]&m[241]&~m[242]&~m[243])|(~m[12]&m[240]&m[241]&~m[242]&~m[243])|(m[12]&~m[240]&~m[241]&m[242]&~m[243])|(~m[12]&m[240]&~m[241]&m[242]&~m[243])|(~m[12]&~m[240]&m[241]&m[242]&~m[243])|(m[12]&~m[240]&~m[241]&~m[242]&m[243])|(~m[12]&m[240]&~m[241]&~m[242]&m[243])|(~m[12]&~m[240]&m[241]&~m[242]&m[243])|(~m[12]&~m[240]&~m[241]&m[242]&m[243]))&BiasedRNG[204])|(((m[12]&m[240]&m[241]&~m[242]&~m[243])|(m[12]&m[240]&~m[241]&m[242]&~m[243])|(m[12]&~m[240]&m[241]&m[242]&~m[243])|(~m[12]&m[240]&m[241]&m[242]&~m[243])|(m[12]&m[240]&~m[241]&~m[242]&m[243])|(m[12]&~m[240]&m[241]&~m[242]&m[243])|(~m[12]&m[240]&m[241]&~m[242]&m[243])|(m[12]&~m[240]&~m[241]&m[242]&m[243])|(~m[12]&m[240]&~m[241]&m[242]&m[243])|(~m[12]&~m[240]&m[241]&m[242]&m[243]))&~BiasedRNG[204])|((m[12]&m[240]&m[241]&m[242]&~m[243])|(m[12]&m[240]&m[241]&~m[242]&m[243])|(m[12]&m[240]&~m[241]&m[242]&m[243])|(m[12]&~m[240]&m[241]&m[242]&m[243])|(~m[12]&m[240]&m[241]&m[242]&m[243])|(m[12]&m[240]&m[241]&m[242]&m[243]))):InitCond[335];
    m[61] = run?((((m[12]&m[244]&~m[245]&~m[246]&~m[247])|(m[12]&~m[244]&m[245]&~m[246]&~m[247])|(~m[12]&m[244]&m[245]&~m[246]&~m[247])|(m[12]&~m[244]&~m[245]&m[246]&~m[247])|(~m[12]&m[244]&~m[245]&m[246]&~m[247])|(~m[12]&~m[244]&m[245]&m[246]&~m[247])|(m[12]&~m[244]&~m[245]&~m[246]&m[247])|(~m[12]&m[244]&~m[245]&~m[246]&m[247])|(~m[12]&~m[244]&m[245]&~m[246]&m[247])|(~m[12]&~m[244]&~m[245]&m[246]&m[247]))&BiasedRNG[205])|(((m[12]&m[244]&m[245]&~m[246]&~m[247])|(m[12]&m[244]&~m[245]&m[246]&~m[247])|(m[12]&~m[244]&m[245]&m[246]&~m[247])|(~m[12]&m[244]&m[245]&m[246]&~m[247])|(m[12]&m[244]&~m[245]&~m[246]&m[247])|(m[12]&~m[244]&m[245]&~m[246]&m[247])|(~m[12]&m[244]&m[245]&~m[246]&m[247])|(m[12]&~m[244]&~m[245]&m[246]&m[247])|(~m[12]&m[244]&~m[245]&m[246]&m[247])|(~m[12]&~m[244]&m[245]&m[246]&m[247]))&~BiasedRNG[205])|((m[12]&m[244]&m[245]&m[246]&~m[247])|(m[12]&m[244]&m[245]&~m[246]&m[247])|(m[12]&m[244]&~m[245]&m[246]&m[247])|(m[12]&~m[244]&m[245]&m[246]&m[247])|(~m[12]&m[244]&m[245]&m[246]&m[247])|(m[12]&m[244]&m[245]&m[246]&m[247]))):InitCond[336];
    m[62] = run?((((m[12]&m[248]&~m[249]&~m[250]&~m[251])|(m[12]&~m[248]&m[249]&~m[250]&~m[251])|(~m[12]&m[248]&m[249]&~m[250]&~m[251])|(m[12]&~m[248]&~m[249]&m[250]&~m[251])|(~m[12]&m[248]&~m[249]&m[250]&~m[251])|(~m[12]&~m[248]&m[249]&m[250]&~m[251])|(m[12]&~m[248]&~m[249]&~m[250]&m[251])|(~m[12]&m[248]&~m[249]&~m[250]&m[251])|(~m[12]&~m[248]&m[249]&~m[250]&m[251])|(~m[12]&~m[248]&~m[249]&m[250]&m[251]))&BiasedRNG[206])|(((m[12]&m[248]&m[249]&~m[250]&~m[251])|(m[12]&m[248]&~m[249]&m[250]&~m[251])|(m[12]&~m[248]&m[249]&m[250]&~m[251])|(~m[12]&m[248]&m[249]&m[250]&~m[251])|(m[12]&m[248]&~m[249]&~m[250]&m[251])|(m[12]&~m[248]&m[249]&~m[250]&m[251])|(~m[12]&m[248]&m[249]&~m[250]&m[251])|(m[12]&~m[248]&~m[249]&m[250]&m[251])|(~m[12]&m[248]&~m[249]&m[250]&m[251])|(~m[12]&~m[248]&m[249]&m[250]&m[251]))&~BiasedRNG[206])|((m[12]&m[248]&m[249]&m[250]&~m[251])|(m[12]&m[248]&m[249]&~m[250]&m[251])|(m[12]&m[248]&~m[249]&m[250]&m[251])|(m[12]&~m[248]&m[249]&m[250]&m[251])|(~m[12]&m[248]&m[249]&m[250]&m[251])|(m[12]&m[248]&m[249]&m[250]&m[251]))):InitCond[337];
    m[63] = run?((((m[13]&m[252]&~m[253]&~m[254]&~m[255])|(m[13]&~m[252]&m[253]&~m[254]&~m[255])|(~m[13]&m[252]&m[253]&~m[254]&~m[255])|(m[13]&~m[252]&~m[253]&m[254]&~m[255])|(~m[13]&m[252]&~m[253]&m[254]&~m[255])|(~m[13]&~m[252]&m[253]&m[254]&~m[255])|(m[13]&~m[252]&~m[253]&~m[254]&m[255])|(~m[13]&m[252]&~m[253]&~m[254]&m[255])|(~m[13]&~m[252]&m[253]&~m[254]&m[255])|(~m[13]&~m[252]&~m[253]&m[254]&m[255]))&BiasedRNG[207])|(((m[13]&m[252]&m[253]&~m[254]&~m[255])|(m[13]&m[252]&~m[253]&m[254]&~m[255])|(m[13]&~m[252]&m[253]&m[254]&~m[255])|(~m[13]&m[252]&m[253]&m[254]&~m[255])|(m[13]&m[252]&~m[253]&~m[254]&m[255])|(m[13]&~m[252]&m[253]&~m[254]&m[255])|(~m[13]&m[252]&m[253]&~m[254]&m[255])|(m[13]&~m[252]&~m[253]&m[254]&m[255])|(~m[13]&m[252]&~m[253]&m[254]&m[255])|(~m[13]&~m[252]&m[253]&m[254]&m[255]))&~BiasedRNG[207])|((m[13]&m[252]&m[253]&m[254]&~m[255])|(m[13]&m[252]&m[253]&~m[254]&m[255])|(m[13]&m[252]&~m[253]&m[254]&m[255])|(m[13]&~m[252]&m[253]&m[254]&m[255])|(~m[13]&m[252]&m[253]&m[254]&m[255])|(m[13]&m[252]&m[253]&m[254]&m[255]))):InitCond[338];
    m[64] = run?((((m[13]&m[256]&~m[257]&~m[258]&~m[259])|(m[13]&~m[256]&m[257]&~m[258]&~m[259])|(~m[13]&m[256]&m[257]&~m[258]&~m[259])|(m[13]&~m[256]&~m[257]&m[258]&~m[259])|(~m[13]&m[256]&~m[257]&m[258]&~m[259])|(~m[13]&~m[256]&m[257]&m[258]&~m[259])|(m[13]&~m[256]&~m[257]&~m[258]&m[259])|(~m[13]&m[256]&~m[257]&~m[258]&m[259])|(~m[13]&~m[256]&m[257]&~m[258]&m[259])|(~m[13]&~m[256]&~m[257]&m[258]&m[259]))&BiasedRNG[208])|(((m[13]&m[256]&m[257]&~m[258]&~m[259])|(m[13]&m[256]&~m[257]&m[258]&~m[259])|(m[13]&~m[256]&m[257]&m[258]&~m[259])|(~m[13]&m[256]&m[257]&m[258]&~m[259])|(m[13]&m[256]&~m[257]&~m[258]&m[259])|(m[13]&~m[256]&m[257]&~m[258]&m[259])|(~m[13]&m[256]&m[257]&~m[258]&m[259])|(m[13]&~m[256]&~m[257]&m[258]&m[259])|(~m[13]&m[256]&~m[257]&m[258]&m[259])|(~m[13]&~m[256]&m[257]&m[258]&m[259]))&~BiasedRNG[208])|((m[13]&m[256]&m[257]&m[258]&~m[259])|(m[13]&m[256]&m[257]&~m[258]&m[259])|(m[13]&m[256]&~m[257]&m[258]&m[259])|(m[13]&~m[256]&m[257]&m[258]&m[259])|(~m[13]&m[256]&m[257]&m[258]&m[259])|(m[13]&m[256]&m[257]&m[258]&m[259]))):InitCond[339];
    m[65] = run?((((m[13]&m[260]&~m[261]&~m[262]&~m[263])|(m[13]&~m[260]&m[261]&~m[262]&~m[263])|(~m[13]&m[260]&m[261]&~m[262]&~m[263])|(m[13]&~m[260]&~m[261]&m[262]&~m[263])|(~m[13]&m[260]&~m[261]&m[262]&~m[263])|(~m[13]&~m[260]&m[261]&m[262]&~m[263])|(m[13]&~m[260]&~m[261]&~m[262]&m[263])|(~m[13]&m[260]&~m[261]&~m[262]&m[263])|(~m[13]&~m[260]&m[261]&~m[262]&m[263])|(~m[13]&~m[260]&~m[261]&m[262]&m[263]))&BiasedRNG[209])|(((m[13]&m[260]&m[261]&~m[262]&~m[263])|(m[13]&m[260]&~m[261]&m[262]&~m[263])|(m[13]&~m[260]&m[261]&m[262]&~m[263])|(~m[13]&m[260]&m[261]&m[262]&~m[263])|(m[13]&m[260]&~m[261]&~m[262]&m[263])|(m[13]&~m[260]&m[261]&~m[262]&m[263])|(~m[13]&m[260]&m[261]&~m[262]&m[263])|(m[13]&~m[260]&~m[261]&m[262]&m[263])|(~m[13]&m[260]&~m[261]&m[262]&m[263])|(~m[13]&~m[260]&m[261]&m[262]&m[263]))&~BiasedRNG[209])|((m[13]&m[260]&m[261]&m[262]&~m[263])|(m[13]&m[260]&m[261]&~m[262]&m[263])|(m[13]&m[260]&~m[261]&m[262]&m[263])|(m[13]&~m[260]&m[261]&m[262]&m[263])|(~m[13]&m[260]&m[261]&m[262]&m[263])|(m[13]&m[260]&m[261]&m[262]&m[263]))):InitCond[340];
    m[66] = run?((((m[14]&m[264]&~m[265]&~m[266]&~m[267])|(m[14]&~m[264]&m[265]&~m[266]&~m[267])|(~m[14]&m[264]&m[265]&~m[266]&~m[267])|(m[14]&~m[264]&~m[265]&m[266]&~m[267])|(~m[14]&m[264]&~m[265]&m[266]&~m[267])|(~m[14]&~m[264]&m[265]&m[266]&~m[267])|(m[14]&~m[264]&~m[265]&~m[266]&m[267])|(~m[14]&m[264]&~m[265]&~m[266]&m[267])|(~m[14]&~m[264]&m[265]&~m[266]&m[267])|(~m[14]&~m[264]&~m[265]&m[266]&m[267]))&BiasedRNG[210])|(((m[14]&m[264]&m[265]&~m[266]&~m[267])|(m[14]&m[264]&~m[265]&m[266]&~m[267])|(m[14]&~m[264]&m[265]&m[266]&~m[267])|(~m[14]&m[264]&m[265]&m[266]&~m[267])|(m[14]&m[264]&~m[265]&~m[266]&m[267])|(m[14]&~m[264]&m[265]&~m[266]&m[267])|(~m[14]&m[264]&m[265]&~m[266]&m[267])|(m[14]&~m[264]&~m[265]&m[266]&m[267])|(~m[14]&m[264]&~m[265]&m[266]&m[267])|(~m[14]&~m[264]&m[265]&m[266]&m[267]))&~BiasedRNG[210])|((m[14]&m[264]&m[265]&m[266]&~m[267])|(m[14]&m[264]&m[265]&~m[266]&m[267])|(m[14]&m[264]&~m[265]&m[266]&m[267])|(m[14]&~m[264]&m[265]&m[266]&m[267])|(~m[14]&m[264]&m[265]&m[266]&m[267])|(m[14]&m[264]&m[265]&m[266]&m[267]))):InitCond[341];
    m[67] = run?((((m[14]&m[268]&~m[269]&~m[270]&~m[271])|(m[14]&~m[268]&m[269]&~m[270]&~m[271])|(~m[14]&m[268]&m[269]&~m[270]&~m[271])|(m[14]&~m[268]&~m[269]&m[270]&~m[271])|(~m[14]&m[268]&~m[269]&m[270]&~m[271])|(~m[14]&~m[268]&m[269]&m[270]&~m[271])|(m[14]&~m[268]&~m[269]&~m[270]&m[271])|(~m[14]&m[268]&~m[269]&~m[270]&m[271])|(~m[14]&~m[268]&m[269]&~m[270]&m[271])|(~m[14]&~m[268]&~m[269]&m[270]&m[271]))&BiasedRNG[211])|(((m[14]&m[268]&m[269]&~m[270]&~m[271])|(m[14]&m[268]&~m[269]&m[270]&~m[271])|(m[14]&~m[268]&m[269]&m[270]&~m[271])|(~m[14]&m[268]&m[269]&m[270]&~m[271])|(m[14]&m[268]&~m[269]&~m[270]&m[271])|(m[14]&~m[268]&m[269]&~m[270]&m[271])|(~m[14]&m[268]&m[269]&~m[270]&m[271])|(m[14]&~m[268]&~m[269]&m[270]&m[271])|(~m[14]&m[268]&~m[269]&m[270]&m[271])|(~m[14]&~m[268]&m[269]&m[270]&m[271]))&~BiasedRNG[211])|((m[14]&m[268]&m[269]&m[270]&~m[271])|(m[14]&m[268]&m[269]&~m[270]&m[271])|(m[14]&m[268]&~m[269]&m[270]&m[271])|(m[14]&~m[268]&m[269]&m[270]&m[271])|(~m[14]&m[268]&m[269]&m[270]&m[271])|(m[14]&m[268]&m[269]&m[270]&m[271]))):InitCond[342];
    m[68] = run?((((m[14]&m[272]&~m[273]&~m[274]&~m[275])|(m[14]&~m[272]&m[273]&~m[274]&~m[275])|(~m[14]&m[272]&m[273]&~m[274]&~m[275])|(m[14]&~m[272]&~m[273]&m[274]&~m[275])|(~m[14]&m[272]&~m[273]&m[274]&~m[275])|(~m[14]&~m[272]&m[273]&m[274]&~m[275])|(m[14]&~m[272]&~m[273]&~m[274]&m[275])|(~m[14]&m[272]&~m[273]&~m[274]&m[275])|(~m[14]&~m[272]&m[273]&~m[274]&m[275])|(~m[14]&~m[272]&~m[273]&m[274]&m[275]))&BiasedRNG[212])|(((m[14]&m[272]&m[273]&~m[274]&~m[275])|(m[14]&m[272]&~m[273]&m[274]&~m[275])|(m[14]&~m[272]&m[273]&m[274]&~m[275])|(~m[14]&m[272]&m[273]&m[274]&~m[275])|(m[14]&m[272]&~m[273]&~m[274]&m[275])|(m[14]&~m[272]&m[273]&~m[274]&m[275])|(~m[14]&m[272]&m[273]&~m[274]&m[275])|(m[14]&~m[272]&~m[273]&m[274]&m[275])|(~m[14]&m[272]&~m[273]&m[274]&m[275])|(~m[14]&~m[272]&m[273]&m[274]&m[275]))&~BiasedRNG[212])|((m[14]&m[272]&m[273]&m[274]&~m[275])|(m[14]&m[272]&m[273]&~m[274]&m[275])|(m[14]&m[272]&~m[273]&m[274]&m[275])|(m[14]&~m[272]&m[273]&m[274]&m[275])|(~m[14]&m[272]&m[273]&m[274]&m[275])|(m[14]&m[272]&m[273]&m[274]&m[275]))):InitCond[343];
    m[69] = run?((((m[15]&m[276]&~m[277]&~m[278]&~m[279])|(m[15]&~m[276]&m[277]&~m[278]&~m[279])|(~m[15]&m[276]&m[277]&~m[278]&~m[279])|(m[15]&~m[276]&~m[277]&m[278]&~m[279])|(~m[15]&m[276]&~m[277]&m[278]&~m[279])|(~m[15]&~m[276]&m[277]&m[278]&~m[279])|(m[15]&~m[276]&~m[277]&~m[278]&m[279])|(~m[15]&m[276]&~m[277]&~m[278]&m[279])|(~m[15]&~m[276]&m[277]&~m[278]&m[279])|(~m[15]&~m[276]&~m[277]&m[278]&m[279]))&BiasedRNG[213])|(((m[15]&m[276]&m[277]&~m[278]&~m[279])|(m[15]&m[276]&~m[277]&m[278]&~m[279])|(m[15]&~m[276]&m[277]&m[278]&~m[279])|(~m[15]&m[276]&m[277]&m[278]&~m[279])|(m[15]&m[276]&~m[277]&~m[278]&m[279])|(m[15]&~m[276]&m[277]&~m[278]&m[279])|(~m[15]&m[276]&m[277]&~m[278]&m[279])|(m[15]&~m[276]&~m[277]&m[278]&m[279])|(~m[15]&m[276]&~m[277]&m[278]&m[279])|(~m[15]&~m[276]&m[277]&m[278]&m[279]))&~BiasedRNG[213])|((m[15]&m[276]&m[277]&m[278]&~m[279])|(m[15]&m[276]&m[277]&~m[278]&m[279])|(m[15]&m[276]&~m[277]&m[278]&m[279])|(m[15]&~m[276]&m[277]&m[278]&m[279])|(~m[15]&m[276]&m[277]&m[278]&m[279])|(m[15]&m[276]&m[277]&m[278]&m[279]))):InitCond[344];
    m[70] = run?((((m[15]&m[280]&~m[281]&~m[282]&~m[283])|(m[15]&~m[280]&m[281]&~m[282]&~m[283])|(~m[15]&m[280]&m[281]&~m[282]&~m[283])|(m[15]&~m[280]&~m[281]&m[282]&~m[283])|(~m[15]&m[280]&~m[281]&m[282]&~m[283])|(~m[15]&~m[280]&m[281]&m[282]&~m[283])|(m[15]&~m[280]&~m[281]&~m[282]&m[283])|(~m[15]&m[280]&~m[281]&~m[282]&m[283])|(~m[15]&~m[280]&m[281]&~m[282]&m[283])|(~m[15]&~m[280]&~m[281]&m[282]&m[283]))&BiasedRNG[214])|(((m[15]&m[280]&m[281]&~m[282]&~m[283])|(m[15]&m[280]&~m[281]&m[282]&~m[283])|(m[15]&~m[280]&m[281]&m[282]&~m[283])|(~m[15]&m[280]&m[281]&m[282]&~m[283])|(m[15]&m[280]&~m[281]&~m[282]&m[283])|(m[15]&~m[280]&m[281]&~m[282]&m[283])|(~m[15]&m[280]&m[281]&~m[282]&m[283])|(m[15]&~m[280]&~m[281]&m[282]&m[283])|(~m[15]&m[280]&~m[281]&m[282]&m[283])|(~m[15]&~m[280]&m[281]&m[282]&m[283]))&~BiasedRNG[214])|((m[15]&m[280]&m[281]&m[282]&~m[283])|(m[15]&m[280]&m[281]&~m[282]&m[283])|(m[15]&m[280]&~m[281]&m[282]&m[283])|(m[15]&~m[280]&m[281]&m[282]&m[283])|(~m[15]&m[280]&m[281]&m[282]&m[283])|(m[15]&m[280]&m[281]&m[282]&m[283]))):InitCond[345];
    m[71] = run?((((m[15]&m[284]&~m[285]&~m[286]&~m[287])|(m[15]&~m[284]&m[285]&~m[286]&~m[287])|(~m[15]&m[284]&m[285]&~m[286]&~m[287])|(m[15]&~m[284]&~m[285]&m[286]&~m[287])|(~m[15]&m[284]&~m[285]&m[286]&~m[287])|(~m[15]&~m[284]&m[285]&m[286]&~m[287])|(m[15]&~m[284]&~m[285]&~m[286]&m[287])|(~m[15]&m[284]&~m[285]&~m[286]&m[287])|(~m[15]&~m[284]&m[285]&~m[286]&m[287])|(~m[15]&~m[284]&~m[285]&m[286]&m[287]))&BiasedRNG[215])|(((m[15]&m[284]&m[285]&~m[286]&~m[287])|(m[15]&m[284]&~m[285]&m[286]&~m[287])|(m[15]&~m[284]&m[285]&m[286]&~m[287])|(~m[15]&m[284]&m[285]&m[286]&~m[287])|(m[15]&m[284]&~m[285]&~m[286]&m[287])|(m[15]&~m[284]&m[285]&~m[286]&m[287])|(~m[15]&m[284]&m[285]&~m[286]&m[287])|(m[15]&~m[284]&~m[285]&m[286]&m[287])|(~m[15]&m[284]&~m[285]&m[286]&m[287])|(~m[15]&~m[284]&m[285]&m[286]&m[287]))&~BiasedRNG[215])|((m[15]&m[284]&m[285]&m[286]&~m[287])|(m[15]&m[284]&m[285]&~m[286]&m[287])|(m[15]&m[284]&~m[285]&m[286]&m[287])|(m[15]&~m[284]&m[285]&m[286]&m[287])|(~m[15]&m[284]&m[285]&m[286]&m[287])|(m[15]&m[284]&m[285]&m[286]&m[287]))):InitCond[346];
    m[72] = run?((((m[16]&m[288]&~m[289]&~m[290]&~m[291])|(m[16]&~m[288]&m[289]&~m[290]&~m[291])|(~m[16]&m[288]&m[289]&~m[290]&~m[291])|(m[16]&~m[288]&~m[289]&m[290]&~m[291])|(~m[16]&m[288]&~m[289]&m[290]&~m[291])|(~m[16]&~m[288]&m[289]&m[290]&~m[291])|(m[16]&~m[288]&~m[289]&~m[290]&m[291])|(~m[16]&m[288]&~m[289]&~m[290]&m[291])|(~m[16]&~m[288]&m[289]&~m[290]&m[291])|(~m[16]&~m[288]&~m[289]&m[290]&m[291]))&BiasedRNG[216])|(((m[16]&m[288]&m[289]&~m[290]&~m[291])|(m[16]&m[288]&~m[289]&m[290]&~m[291])|(m[16]&~m[288]&m[289]&m[290]&~m[291])|(~m[16]&m[288]&m[289]&m[290]&~m[291])|(m[16]&m[288]&~m[289]&~m[290]&m[291])|(m[16]&~m[288]&m[289]&~m[290]&m[291])|(~m[16]&m[288]&m[289]&~m[290]&m[291])|(m[16]&~m[288]&~m[289]&m[290]&m[291])|(~m[16]&m[288]&~m[289]&m[290]&m[291])|(~m[16]&~m[288]&m[289]&m[290]&m[291]))&~BiasedRNG[216])|((m[16]&m[288]&m[289]&m[290]&~m[291])|(m[16]&m[288]&m[289]&~m[290]&m[291])|(m[16]&m[288]&~m[289]&m[290]&m[291])|(m[16]&~m[288]&m[289]&m[290]&m[291])|(~m[16]&m[288]&m[289]&m[290]&m[291])|(m[16]&m[288]&m[289]&m[290]&m[291]))):InitCond[347];
    m[73] = run?((((m[16]&m[292]&~m[293]&~m[294]&~m[295])|(m[16]&~m[292]&m[293]&~m[294]&~m[295])|(~m[16]&m[292]&m[293]&~m[294]&~m[295])|(m[16]&~m[292]&~m[293]&m[294]&~m[295])|(~m[16]&m[292]&~m[293]&m[294]&~m[295])|(~m[16]&~m[292]&m[293]&m[294]&~m[295])|(m[16]&~m[292]&~m[293]&~m[294]&m[295])|(~m[16]&m[292]&~m[293]&~m[294]&m[295])|(~m[16]&~m[292]&m[293]&~m[294]&m[295])|(~m[16]&~m[292]&~m[293]&m[294]&m[295]))&BiasedRNG[217])|(((m[16]&m[292]&m[293]&~m[294]&~m[295])|(m[16]&m[292]&~m[293]&m[294]&~m[295])|(m[16]&~m[292]&m[293]&m[294]&~m[295])|(~m[16]&m[292]&m[293]&m[294]&~m[295])|(m[16]&m[292]&~m[293]&~m[294]&m[295])|(m[16]&~m[292]&m[293]&~m[294]&m[295])|(~m[16]&m[292]&m[293]&~m[294]&m[295])|(m[16]&~m[292]&~m[293]&m[294]&m[295])|(~m[16]&m[292]&~m[293]&m[294]&m[295])|(~m[16]&~m[292]&m[293]&m[294]&m[295]))&~BiasedRNG[217])|((m[16]&m[292]&m[293]&m[294]&~m[295])|(m[16]&m[292]&m[293]&~m[294]&m[295])|(m[16]&m[292]&~m[293]&m[294]&m[295])|(m[16]&~m[292]&m[293]&m[294]&m[295])|(~m[16]&m[292]&m[293]&m[294]&m[295])|(m[16]&m[292]&m[293]&m[294]&m[295]))):InitCond[348];
    m[74] = run?((((m[16]&m[296]&~m[297]&~m[298]&~m[299])|(m[16]&~m[296]&m[297]&~m[298]&~m[299])|(~m[16]&m[296]&m[297]&~m[298]&~m[299])|(m[16]&~m[296]&~m[297]&m[298]&~m[299])|(~m[16]&m[296]&~m[297]&m[298]&~m[299])|(~m[16]&~m[296]&m[297]&m[298]&~m[299])|(m[16]&~m[296]&~m[297]&~m[298]&m[299])|(~m[16]&m[296]&~m[297]&~m[298]&m[299])|(~m[16]&~m[296]&m[297]&~m[298]&m[299])|(~m[16]&~m[296]&~m[297]&m[298]&m[299]))&BiasedRNG[218])|(((m[16]&m[296]&m[297]&~m[298]&~m[299])|(m[16]&m[296]&~m[297]&m[298]&~m[299])|(m[16]&~m[296]&m[297]&m[298]&~m[299])|(~m[16]&m[296]&m[297]&m[298]&~m[299])|(m[16]&m[296]&~m[297]&~m[298]&m[299])|(m[16]&~m[296]&m[297]&~m[298]&m[299])|(~m[16]&m[296]&m[297]&~m[298]&m[299])|(m[16]&~m[296]&~m[297]&m[298]&m[299])|(~m[16]&m[296]&~m[297]&m[298]&m[299])|(~m[16]&~m[296]&m[297]&m[298]&m[299]))&~BiasedRNG[218])|((m[16]&m[296]&m[297]&m[298]&~m[299])|(m[16]&m[296]&m[297]&~m[298]&m[299])|(m[16]&m[296]&~m[297]&m[298]&m[299])|(m[16]&~m[296]&m[297]&m[298]&m[299])|(~m[16]&m[296]&m[297]&m[298]&m[299])|(m[16]&m[296]&m[297]&m[298]&m[299]))):InitCond[349];
    m[75] = run?((((m[17]&m[300]&~m[301]&~m[302]&~m[303])|(m[17]&~m[300]&m[301]&~m[302]&~m[303])|(~m[17]&m[300]&m[301]&~m[302]&~m[303])|(m[17]&~m[300]&~m[301]&m[302]&~m[303])|(~m[17]&m[300]&~m[301]&m[302]&~m[303])|(~m[17]&~m[300]&m[301]&m[302]&~m[303])|(m[17]&~m[300]&~m[301]&~m[302]&m[303])|(~m[17]&m[300]&~m[301]&~m[302]&m[303])|(~m[17]&~m[300]&m[301]&~m[302]&m[303])|(~m[17]&~m[300]&~m[301]&m[302]&m[303]))&BiasedRNG[219])|(((m[17]&m[300]&m[301]&~m[302]&~m[303])|(m[17]&m[300]&~m[301]&m[302]&~m[303])|(m[17]&~m[300]&m[301]&m[302]&~m[303])|(~m[17]&m[300]&m[301]&m[302]&~m[303])|(m[17]&m[300]&~m[301]&~m[302]&m[303])|(m[17]&~m[300]&m[301]&~m[302]&m[303])|(~m[17]&m[300]&m[301]&~m[302]&m[303])|(m[17]&~m[300]&~m[301]&m[302]&m[303])|(~m[17]&m[300]&~m[301]&m[302]&m[303])|(~m[17]&~m[300]&m[301]&m[302]&m[303]))&~BiasedRNG[219])|((m[17]&m[300]&m[301]&m[302]&~m[303])|(m[17]&m[300]&m[301]&~m[302]&m[303])|(m[17]&m[300]&~m[301]&m[302]&m[303])|(m[17]&~m[300]&m[301]&m[302]&m[303])|(~m[17]&m[300]&m[301]&m[302]&m[303])|(m[17]&m[300]&m[301]&m[302]&m[303]))):InitCond[350];
    m[76] = run?((((m[17]&m[304]&~m[305]&~m[306]&~m[307])|(m[17]&~m[304]&m[305]&~m[306]&~m[307])|(~m[17]&m[304]&m[305]&~m[306]&~m[307])|(m[17]&~m[304]&~m[305]&m[306]&~m[307])|(~m[17]&m[304]&~m[305]&m[306]&~m[307])|(~m[17]&~m[304]&m[305]&m[306]&~m[307])|(m[17]&~m[304]&~m[305]&~m[306]&m[307])|(~m[17]&m[304]&~m[305]&~m[306]&m[307])|(~m[17]&~m[304]&m[305]&~m[306]&m[307])|(~m[17]&~m[304]&~m[305]&m[306]&m[307]))&BiasedRNG[220])|(((m[17]&m[304]&m[305]&~m[306]&~m[307])|(m[17]&m[304]&~m[305]&m[306]&~m[307])|(m[17]&~m[304]&m[305]&m[306]&~m[307])|(~m[17]&m[304]&m[305]&m[306]&~m[307])|(m[17]&m[304]&~m[305]&~m[306]&m[307])|(m[17]&~m[304]&m[305]&~m[306]&m[307])|(~m[17]&m[304]&m[305]&~m[306]&m[307])|(m[17]&~m[304]&~m[305]&m[306]&m[307])|(~m[17]&m[304]&~m[305]&m[306]&m[307])|(~m[17]&~m[304]&m[305]&m[306]&m[307]))&~BiasedRNG[220])|((m[17]&m[304]&m[305]&m[306]&~m[307])|(m[17]&m[304]&m[305]&~m[306]&m[307])|(m[17]&m[304]&~m[305]&m[306]&m[307])|(m[17]&~m[304]&m[305]&m[306]&m[307])|(~m[17]&m[304]&m[305]&m[306]&m[307])|(m[17]&m[304]&m[305]&m[306]&m[307]))):InitCond[351];
    m[77] = run?((((m[17]&m[308]&~m[309]&~m[310]&~m[311])|(m[17]&~m[308]&m[309]&~m[310]&~m[311])|(~m[17]&m[308]&m[309]&~m[310]&~m[311])|(m[17]&~m[308]&~m[309]&m[310]&~m[311])|(~m[17]&m[308]&~m[309]&m[310]&~m[311])|(~m[17]&~m[308]&m[309]&m[310]&~m[311])|(m[17]&~m[308]&~m[309]&~m[310]&m[311])|(~m[17]&m[308]&~m[309]&~m[310]&m[311])|(~m[17]&~m[308]&m[309]&~m[310]&m[311])|(~m[17]&~m[308]&~m[309]&m[310]&m[311]))&BiasedRNG[221])|(((m[17]&m[308]&m[309]&~m[310]&~m[311])|(m[17]&m[308]&~m[309]&m[310]&~m[311])|(m[17]&~m[308]&m[309]&m[310]&~m[311])|(~m[17]&m[308]&m[309]&m[310]&~m[311])|(m[17]&m[308]&~m[309]&~m[310]&m[311])|(m[17]&~m[308]&m[309]&~m[310]&m[311])|(~m[17]&m[308]&m[309]&~m[310]&m[311])|(m[17]&~m[308]&~m[309]&m[310]&m[311])|(~m[17]&m[308]&~m[309]&m[310]&m[311])|(~m[17]&~m[308]&m[309]&m[310]&m[311]))&~BiasedRNG[221])|((m[17]&m[308]&m[309]&m[310]&~m[311])|(m[17]&m[308]&m[309]&~m[310]&m[311])|(m[17]&m[308]&~m[309]&m[310]&m[311])|(m[17]&~m[308]&m[309]&m[310]&m[311])|(~m[17]&m[308]&m[309]&m[310]&m[311])|(m[17]&m[308]&m[309]&m[310]&m[311]))):InitCond[352];
    m[78] = run?((((m[18]&m[312]&~m[313]&~m[314]&~m[315])|(m[18]&~m[312]&m[313]&~m[314]&~m[315])|(~m[18]&m[312]&m[313]&~m[314]&~m[315])|(m[18]&~m[312]&~m[313]&m[314]&~m[315])|(~m[18]&m[312]&~m[313]&m[314]&~m[315])|(~m[18]&~m[312]&m[313]&m[314]&~m[315])|(m[18]&~m[312]&~m[313]&~m[314]&m[315])|(~m[18]&m[312]&~m[313]&~m[314]&m[315])|(~m[18]&~m[312]&m[313]&~m[314]&m[315])|(~m[18]&~m[312]&~m[313]&m[314]&m[315]))&BiasedRNG[222])|(((m[18]&m[312]&m[313]&~m[314]&~m[315])|(m[18]&m[312]&~m[313]&m[314]&~m[315])|(m[18]&~m[312]&m[313]&m[314]&~m[315])|(~m[18]&m[312]&m[313]&m[314]&~m[315])|(m[18]&m[312]&~m[313]&~m[314]&m[315])|(m[18]&~m[312]&m[313]&~m[314]&m[315])|(~m[18]&m[312]&m[313]&~m[314]&m[315])|(m[18]&~m[312]&~m[313]&m[314]&m[315])|(~m[18]&m[312]&~m[313]&m[314]&m[315])|(~m[18]&~m[312]&m[313]&m[314]&m[315]))&~BiasedRNG[222])|((m[18]&m[312]&m[313]&m[314]&~m[315])|(m[18]&m[312]&m[313]&~m[314]&m[315])|(m[18]&m[312]&~m[313]&m[314]&m[315])|(m[18]&~m[312]&m[313]&m[314]&m[315])|(~m[18]&m[312]&m[313]&m[314]&m[315])|(m[18]&m[312]&m[313]&m[314]&m[315]))):InitCond[353];
    m[79] = run?((((m[18]&m[316]&~m[317]&~m[318]&~m[319])|(m[18]&~m[316]&m[317]&~m[318]&~m[319])|(~m[18]&m[316]&m[317]&~m[318]&~m[319])|(m[18]&~m[316]&~m[317]&m[318]&~m[319])|(~m[18]&m[316]&~m[317]&m[318]&~m[319])|(~m[18]&~m[316]&m[317]&m[318]&~m[319])|(m[18]&~m[316]&~m[317]&~m[318]&m[319])|(~m[18]&m[316]&~m[317]&~m[318]&m[319])|(~m[18]&~m[316]&m[317]&~m[318]&m[319])|(~m[18]&~m[316]&~m[317]&m[318]&m[319]))&BiasedRNG[223])|(((m[18]&m[316]&m[317]&~m[318]&~m[319])|(m[18]&m[316]&~m[317]&m[318]&~m[319])|(m[18]&~m[316]&m[317]&m[318]&~m[319])|(~m[18]&m[316]&m[317]&m[318]&~m[319])|(m[18]&m[316]&~m[317]&~m[318]&m[319])|(m[18]&~m[316]&m[317]&~m[318]&m[319])|(~m[18]&m[316]&m[317]&~m[318]&m[319])|(m[18]&~m[316]&~m[317]&m[318]&m[319])|(~m[18]&m[316]&~m[317]&m[318]&m[319])|(~m[18]&~m[316]&m[317]&m[318]&m[319]))&~BiasedRNG[223])|((m[18]&m[316]&m[317]&m[318]&~m[319])|(m[18]&m[316]&m[317]&~m[318]&m[319])|(m[18]&m[316]&~m[317]&m[318]&m[319])|(m[18]&~m[316]&m[317]&m[318]&m[319])|(~m[18]&m[316]&m[317]&m[318]&m[319])|(m[18]&m[316]&m[317]&m[318]&m[319]))):InitCond[354];
    m[80] = run?((((m[18]&m[320]&~m[321]&~m[322]&~m[323])|(m[18]&~m[320]&m[321]&~m[322]&~m[323])|(~m[18]&m[320]&m[321]&~m[322]&~m[323])|(m[18]&~m[320]&~m[321]&m[322]&~m[323])|(~m[18]&m[320]&~m[321]&m[322]&~m[323])|(~m[18]&~m[320]&m[321]&m[322]&~m[323])|(m[18]&~m[320]&~m[321]&~m[322]&m[323])|(~m[18]&m[320]&~m[321]&~m[322]&m[323])|(~m[18]&~m[320]&m[321]&~m[322]&m[323])|(~m[18]&~m[320]&~m[321]&m[322]&m[323]))&BiasedRNG[224])|(((m[18]&m[320]&m[321]&~m[322]&~m[323])|(m[18]&m[320]&~m[321]&m[322]&~m[323])|(m[18]&~m[320]&m[321]&m[322]&~m[323])|(~m[18]&m[320]&m[321]&m[322]&~m[323])|(m[18]&m[320]&~m[321]&~m[322]&m[323])|(m[18]&~m[320]&m[321]&~m[322]&m[323])|(~m[18]&m[320]&m[321]&~m[322]&m[323])|(m[18]&~m[320]&~m[321]&m[322]&m[323])|(~m[18]&m[320]&~m[321]&m[322]&m[323])|(~m[18]&~m[320]&m[321]&m[322]&m[323]))&~BiasedRNG[224])|((m[18]&m[320]&m[321]&m[322]&~m[323])|(m[18]&m[320]&m[321]&~m[322]&m[323])|(m[18]&m[320]&~m[321]&m[322]&m[323])|(m[18]&~m[320]&m[321]&m[322]&m[323])|(~m[18]&m[320]&m[321]&m[322]&m[323])|(m[18]&m[320]&m[321]&m[322]&m[323]))):InitCond[355];
    m[81] = run?((((m[19]&m[324]&~m[325]&~m[326]&~m[327])|(m[19]&~m[324]&m[325]&~m[326]&~m[327])|(~m[19]&m[324]&m[325]&~m[326]&~m[327])|(m[19]&~m[324]&~m[325]&m[326]&~m[327])|(~m[19]&m[324]&~m[325]&m[326]&~m[327])|(~m[19]&~m[324]&m[325]&m[326]&~m[327])|(m[19]&~m[324]&~m[325]&~m[326]&m[327])|(~m[19]&m[324]&~m[325]&~m[326]&m[327])|(~m[19]&~m[324]&m[325]&~m[326]&m[327])|(~m[19]&~m[324]&~m[325]&m[326]&m[327]))&BiasedRNG[225])|(((m[19]&m[324]&m[325]&~m[326]&~m[327])|(m[19]&m[324]&~m[325]&m[326]&~m[327])|(m[19]&~m[324]&m[325]&m[326]&~m[327])|(~m[19]&m[324]&m[325]&m[326]&~m[327])|(m[19]&m[324]&~m[325]&~m[326]&m[327])|(m[19]&~m[324]&m[325]&~m[326]&m[327])|(~m[19]&m[324]&m[325]&~m[326]&m[327])|(m[19]&~m[324]&~m[325]&m[326]&m[327])|(~m[19]&m[324]&~m[325]&m[326]&m[327])|(~m[19]&~m[324]&m[325]&m[326]&m[327]))&~BiasedRNG[225])|((m[19]&m[324]&m[325]&m[326]&~m[327])|(m[19]&m[324]&m[325]&~m[326]&m[327])|(m[19]&m[324]&~m[325]&m[326]&m[327])|(m[19]&~m[324]&m[325]&m[326]&m[327])|(~m[19]&m[324]&m[325]&m[326]&m[327])|(m[19]&m[324]&m[325]&m[326]&m[327]))):InitCond[356];
    m[82] = run?((((m[19]&m[328]&~m[329]&~m[330]&~m[331])|(m[19]&~m[328]&m[329]&~m[330]&~m[331])|(~m[19]&m[328]&m[329]&~m[330]&~m[331])|(m[19]&~m[328]&~m[329]&m[330]&~m[331])|(~m[19]&m[328]&~m[329]&m[330]&~m[331])|(~m[19]&~m[328]&m[329]&m[330]&~m[331])|(m[19]&~m[328]&~m[329]&~m[330]&m[331])|(~m[19]&m[328]&~m[329]&~m[330]&m[331])|(~m[19]&~m[328]&m[329]&~m[330]&m[331])|(~m[19]&~m[328]&~m[329]&m[330]&m[331]))&BiasedRNG[226])|(((m[19]&m[328]&m[329]&~m[330]&~m[331])|(m[19]&m[328]&~m[329]&m[330]&~m[331])|(m[19]&~m[328]&m[329]&m[330]&~m[331])|(~m[19]&m[328]&m[329]&m[330]&~m[331])|(m[19]&m[328]&~m[329]&~m[330]&m[331])|(m[19]&~m[328]&m[329]&~m[330]&m[331])|(~m[19]&m[328]&m[329]&~m[330]&m[331])|(m[19]&~m[328]&~m[329]&m[330]&m[331])|(~m[19]&m[328]&~m[329]&m[330]&m[331])|(~m[19]&~m[328]&m[329]&m[330]&m[331]))&~BiasedRNG[226])|((m[19]&m[328]&m[329]&m[330]&~m[331])|(m[19]&m[328]&m[329]&~m[330]&m[331])|(m[19]&m[328]&~m[329]&m[330]&m[331])|(m[19]&~m[328]&m[329]&m[330]&m[331])|(~m[19]&m[328]&m[329]&m[330]&m[331])|(m[19]&m[328]&m[329]&m[330]&m[331]))):InitCond[357];
    m[83] = run?((((m[19]&m[332]&~m[333]&~m[334]&~m[335])|(m[19]&~m[332]&m[333]&~m[334]&~m[335])|(~m[19]&m[332]&m[333]&~m[334]&~m[335])|(m[19]&~m[332]&~m[333]&m[334]&~m[335])|(~m[19]&m[332]&~m[333]&m[334]&~m[335])|(~m[19]&~m[332]&m[333]&m[334]&~m[335])|(m[19]&~m[332]&~m[333]&~m[334]&m[335])|(~m[19]&m[332]&~m[333]&~m[334]&m[335])|(~m[19]&~m[332]&m[333]&~m[334]&m[335])|(~m[19]&~m[332]&~m[333]&m[334]&m[335]))&BiasedRNG[227])|(((m[19]&m[332]&m[333]&~m[334]&~m[335])|(m[19]&m[332]&~m[333]&m[334]&~m[335])|(m[19]&~m[332]&m[333]&m[334]&~m[335])|(~m[19]&m[332]&m[333]&m[334]&~m[335])|(m[19]&m[332]&~m[333]&~m[334]&m[335])|(m[19]&~m[332]&m[333]&~m[334]&m[335])|(~m[19]&m[332]&m[333]&~m[334]&m[335])|(m[19]&~m[332]&~m[333]&m[334]&m[335])|(~m[19]&m[332]&~m[333]&m[334]&m[335])|(~m[19]&~m[332]&m[333]&m[334]&m[335]))&~BiasedRNG[227])|((m[19]&m[332]&m[333]&m[334]&~m[335])|(m[19]&m[332]&m[333]&~m[334]&m[335])|(m[19]&m[332]&~m[333]&m[334]&m[335])|(m[19]&~m[332]&m[333]&m[334]&m[335])|(~m[19]&m[332]&m[333]&m[334]&m[335])|(m[19]&m[332]&m[333]&m[334]&m[335]))):InitCond[358];
    m[84] = run?((((m[20]&m[336]&~m[337]&~m[338]&~m[339])|(m[20]&~m[336]&m[337]&~m[338]&~m[339])|(~m[20]&m[336]&m[337]&~m[338]&~m[339])|(m[20]&~m[336]&~m[337]&m[338]&~m[339])|(~m[20]&m[336]&~m[337]&m[338]&~m[339])|(~m[20]&~m[336]&m[337]&m[338]&~m[339])|(m[20]&~m[336]&~m[337]&~m[338]&m[339])|(~m[20]&m[336]&~m[337]&~m[338]&m[339])|(~m[20]&~m[336]&m[337]&~m[338]&m[339])|(~m[20]&~m[336]&~m[337]&m[338]&m[339]))&BiasedRNG[228])|(((m[20]&m[336]&m[337]&~m[338]&~m[339])|(m[20]&m[336]&~m[337]&m[338]&~m[339])|(m[20]&~m[336]&m[337]&m[338]&~m[339])|(~m[20]&m[336]&m[337]&m[338]&~m[339])|(m[20]&m[336]&~m[337]&~m[338]&m[339])|(m[20]&~m[336]&m[337]&~m[338]&m[339])|(~m[20]&m[336]&m[337]&~m[338]&m[339])|(m[20]&~m[336]&~m[337]&m[338]&m[339])|(~m[20]&m[336]&~m[337]&m[338]&m[339])|(~m[20]&~m[336]&m[337]&m[338]&m[339]))&~BiasedRNG[228])|((m[20]&m[336]&m[337]&m[338]&~m[339])|(m[20]&m[336]&m[337]&~m[338]&m[339])|(m[20]&m[336]&~m[337]&m[338]&m[339])|(m[20]&~m[336]&m[337]&m[338]&m[339])|(~m[20]&m[336]&m[337]&m[338]&m[339])|(m[20]&m[336]&m[337]&m[338]&m[339]))):InitCond[359];
    m[85] = run?((((m[20]&m[340]&~m[341]&~m[342]&~m[343])|(m[20]&~m[340]&m[341]&~m[342]&~m[343])|(~m[20]&m[340]&m[341]&~m[342]&~m[343])|(m[20]&~m[340]&~m[341]&m[342]&~m[343])|(~m[20]&m[340]&~m[341]&m[342]&~m[343])|(~m[20]&~m[340]&m[341]&m[342]&~m[343])|(m[20]&~m[340]&~m[341]&~m[342]&m[343])|(~m[20]&m[340]&~m[341]&~m[342]&m[343])|(~m[20]&~m[340]&m[341]&~m[342]&m[343])|(~m[20]&~m[340]&~m[341]&m[342]&m[343]))&BiasedRNG[229])|(((m[20]&m[340]&m[341]&~m[342]&~m[343])|(m[20]&m[340]&~m[341]&m[342]&~m[343])|(m[20]&~m[340]&m[341]&m[342]&~m[343])|(~m[20]&m[340]&m[341]&m[342]&~m[343])|(m[20]&m[340]&~m[341]&~m[342]&m[343])|(m[20]&~m[340]&m[341]&~m[342]&m[343])|(~m[20]&m[340]&m[341]&~m[342]&m[343])|(m[20]&~m[340]&~m[341]&m[342]&m[343])|(~m[20]&m[340]&~m[341]&m[342]&m[343])|(~m[20]&~m[340]&m[341]&m[342]&m[343]))&~BiasedRNG[229])|((m[20]&m[340]&m[341]&m[342]&~m[343])|(m[20]&m[340]&m[341]&~m[342]&m[343])|(m[20]&m[340]&~m[341]&m[342]&m[343])|(m[20]&~m[340]&m[341]&m[342]&m[343])|(~m[20]&m[340]&m[341]&m[342]&m[343])|(m[20]&m[340]&m[341]&m[342]&m[343]))):InitCond[360];
    m[86] = run?((((m[20]&m[344]&~m[345]&~m[346]&~m[347])|(m[20]&~m[344]&m[345]&~m[346]&~m[347])|(~m[20]&m[344]&m[345]&~m[346]&~m[347])|(m[20]&~m[344]&~m[345]&m[346]&~m[347])|(~m[20]&m[344]&~m[345]&m[346]&~m[347])|(~m[20]&~m[344]&m[345]&m[346]&~m[347])|(m[20]&~m[344]&~m[345]&~m[346]&m[347])|(~m[20]&m[344]&~m[345]&~m[346]&m[347])|(~m[20]&~m[344]&m[345]&~m[346]&m[347])|(~m[20]&~m[344]&~m[345]&m[346]&m[347]))&BiasedRNG[230])|(((m[20]&m[344]&m[345]&~m[346]&~m[347])|(m[20]&m[344]&~m[345]&m[346]&~m[347])|(m[20]&~m[344]&m[345]&m[346]&~m[347])|(~m[20]&m[344]&m[345]&m[346]&~m[347])|(m[20]&m[344]&~m[345]&~m[346]&m[347])|(m[20]&~m[344]&m[345]&~m[346]&m[347])|(~m[20]&m[344]&m[345]&~m[346]&m[347])|(m[20]&~m[344]&~m[345]&m[346]&m[347])|(~m[20]&m[344]&~m[345]&m[346]&m[347])|(~m[20]&~m[344]&m[345]&m[346]&m[347]))&~BiasedRNG[230])|((m[20]&m[344]&m[345]&m[346]&~m[347])|(m[20]&m[344]&m[345]&~m[346]&m[347])|(m[20]&m[344]&~m[345]&m[346]&m[347])|(m[20]&~m[344]&m[345]&m[346]&m[347])|(~m[20]&m[344]&m[345]&m[346]&m[347])|(m[20]&m[344]&m[345]&m[346]&m[347]))):InitCond[361];
    m[87] = run?((((m[21]&m[348]&~m[349]&~m[350]&~m[351])|(m[21]&~m[348]&m[349]&~m[350]&~m[351])|(~m[21]&m[348]&m[349]&~m[350]&~m[351])|(m[21]&~m[348]&~m[349]&m[350]&~m[351])|(~m[21]&m[348]&~m[349]&m[350]&~m[351])|(~m[21]&~m[348]&m[349]&m[350]&~m[351])|(m[21]&~m[348]&~m[349]&~m[350]&m[351])|(~m[21]&m[348]&~m[349]&~m[350]&m[351])|(~m[21]&~m[348]&m[349]&~m[350]&m[351])|(~m[21]&~m[348]&~m[349]&m[350]&m[351]))&BiasedRNG[231])|(((m[21]&m[348]&m[349]&~m[350]&~m[351])|(m[21]&m[348]&~m[349]&m[350]&~m[351])|(m[21]&~m[348]&m[349]&m[350]&~m[351])|(~m[21]&m[348]&m[349]&m[350]&~m[351])|(m[21]&m[348]&~m[349]&~m[350]&m[351])|(m[21]&~m[348]&m[349]&~m[350]&m[351])|(~m[21]&m[348]&m[349]&~m[350]&m[351])|(m[21]&~m[348]&~m[349]&m[350]&m[351])|(~m[21]&m[348]&~m[349]&m[350]&m[351])|(~m[21]&~m[348]&m[349]&m[350]&m[351]))&~BiasedRNG[231])|((m[21]&m[348]&m[349]&m[350]&~m[351])|(m[21]&m[348]&m[349]&~m[350]&m[351])|(m[21]&m[348]&~m[349]&m[350]&m[351])|(m[21]&~m[348]&m[349]&m[350]&m[351])|(~m[21]&m[348]&m[349]&m[350]&m[351])|(m[21]&m[348]&m[349]&m[350]&m[351]))):InitCond[362];
    m[88] = run?((((m[21]&m[352]&~m[353]&~m[354]&~m[355])|(m[21]&~m[352]&m[353]&~m[354]&~m[355])|(~m[21]&m[352]&m[353]&~m[354]&~m[355])|(m[21]&~m[352]&~m[353]&m[354]&~m[355])|(~m[21]&m[352]&~m[353]&m[354]&~m[355])|(~m[21]&~m[352]&m[353]&m[354]&~m[355])|(m[21]&~m[352]&~m[353]&~m[354]&m[355])|(~m[21]&m[352]&~m[353]&~m[354]&m[355])|(~m[21]&~m[352]&m[353]&~m[354]&m[355])|(~m[21]&~m[352]&~m[353]&m[354]&m[355]))&BiasedRNG[232])|(((m[21]&m[352]&m[353]&~m[354]&~m[355])|(m[21]&m[352]&~m[353]&m[354]&~m[355])|(m[21]&~m[352]&m[353]&m[354]&~m[355])|(~m[21]&m[352]&m[353]&m[354]&~m[355])|(m[21]&m[352]&~m[353]&~m[354]&m[355])|(m[21]&~m[352]&m[353]&~m[354]&m[355])|(~m[21]&m[352]&m[353]&~m[354]&m[355])|(m[21]&~m[352]&~m[353]&m[354]&m[355])|(~m[21]&m[352]&~m[353]&m[354]&m[355])|(~m[21]&~m[352]&m[353]&m[354]&m[355]))&~BiasedRNG[232])|((m[21]&m[352]&m[353]&m[354]&~m[355])|(m[21]&m[352]&m[353]&~m[354]&m[355])|(m[21]&m[352]&~m[353]&m[354]&m[355])|(m[21]&~m[352]&m[353]&m[354]&m[355])|(~m[21]&m[352]&m[353]&m[354]&m[355])|(m[21]&m[352]&m[353]&m[354]&m[355]))):InitCond[363];
    m[89] = run?((((m[21]&m[356]&~m[357]&~m[358]&~m[359])|(m[21]&~m[356]&m[357]&~m[358]&~m[359])|(~m[21]&m[356]&m[357]&~m[358]&~m[359])|(m[21]&~m[356]&~m[357]&m[358]&~m[359])|(~m[21]&m[356]&~m[357]&m[358]&~m[359])|(~m[21]&~m[356]&m[357]&m[358]&~m[359])|(m[21]&~m[356]&~m[357]&~m[358]&m[359])|(~m[21]&m[356]&~m[357]&~m[358]&m[359])|(~m[21]&~m[356]&m[357]&~m[358]&m[359])|(~m[21]&~m[356]&~m[357]&m[358]&m[359]))&BiasedRNG[233])|(((m[21]&m[356]&m[357]&~m[358]&~m[359])|(m[21]&m[356]&~m[357]&m[358]&~m[359])|(m[21]&~m[356]&m[357]&m[358]&~m[359])|(~m[21]&m[356]&m[357]&m[358]&~m[359])|(m[21]&m[356]&~m[357]&~m[358]&m[359])|(m[21]&~m[356]&m[357]&~m[358]&m[359])|(~m[21]&m[356]&m[357]&~m[358]&m[359])|(m[21]&~m[356]&~m[357]&m[358]&m[359])|(~m[21]&m[356]&~m[357]&m[358]&m[359])|(~m[21]&~m[356]&m[357]&m[358]&m[359]))&~BiasedRNG[233])|((m[21]&m[356]&m[357]&m[358]&~m[359])|(m[21]&m[356]&m[357]&~m[358]&m[359])|(m[21]&m[356]&~m[357]&m[358]&m[359])|(m[21]&~m[356]&m[357]&m[358]&m[359])|(~m[21]&m[356]&m[357]&m[358]&m[359])|(m[21]&m[356]&m[357]&m[358]&m[359]))):InitCond[364];
    m[90] = run?((((m[22]&m[360]&~m[361]&~m[362]&~m[363])|(m[22]&~m[360]&m[361]&~m[362]&~m[363])|(~m[22]&m[360]&m[361]&~m[362]&~m[363])|(m[22]&~m[360]&~m[361]&m[362]&~m[363])|(~m[22]&m[360]&~m[361]&m[362]&~m[363])|(~m[22]&~m[360]&m[361]&m[362]&~m[363])|(m[22]&~m[360]&~m[361]&~m[362]&m[363])|(~m[22]&m[360]&~m[361]&~m[362]&m[363])|(~m[22]&~m[360]&m[361]&~m[362]&m[363])|(~m[22]&~m[360]&~m[361]&m[362]&m[363]))&BiasedRNG[234])|(((m[22]&m[360]&m[361]&~m[362]&~m[363])|(m[22]&m[360]&~m[361]&m[362]&~m[363])|(m[22]&~m[360]&m[361]&m[362]&~m[363])|(~m[22]&m[360]&m[361]&m[362]&~m[363])|(m[22]&m[360]&~m[361]&~m[362]&m[363])|(m[22]&~m[360]&m[361]&~m[362]&m[363])|(~m[22]&m[360]&m[361]&~m[362]&m[363])|(m[22]&~m[360]&~m[361]&m[362]&m[363])|(~m[22]&m[360]&~m[361]&m[362]&m[363])|(~m[22]&~m[360]&m[361]&m[362]&m[363]))&~BiasedRNG[234])|((m[22]&m[360]&m[361]&m[362]&~m[363])|(m[22]&m[360]&m[361]&~m[362]&m[363])|(m[22]&m[360]&~m[361]&m[362]&m[363])|(m[22]&~m[360]&m[361]&m[362]&m[363])|(~m[22]&m[360]&m[361]&m[362]&m[363])|(m[22]&m[360]&m[361]&m[362]&m[363]))):InitCond[365];
    m[91] = run?((((m[22]&m[364]&~m[365]&~m[366]&~m[367])|(m[22]&~m[364]&m[365]&~m[366]&~m[367])|(~m[22]&m[364]&m[365]&~m[366]&~m[367])|(m[22]&~m[364]&~m[365]&m[366]&~m[367])|(~m[22]&m[364]&~m[365]&m[366]&~m[367])|(~m[22]&~m[364]&m[365]&m[366]&~m[367])|(m[22]&~m[364]&~m[365]&~m[366]&m[367])|(~m[22]&m[364]&~m[365]&~m[366]&m[367])|(~m[22]&~m[364]&m[365]&~m[366]&m[367])|(~m[22]&~m[364]&~m[365]&m[366]&m[367]))&BiasedRNG[235])|(((m[22]&m[364]&m[365]&~m[366]&~m[367])|(m[22]&m[364]&~m[365]&m[366]&~m[367])|(m[22]&~m[364]&m[365]&m[366]&~m[367])|(~m[22]&m[364]&m[365]&m[366]&~m[367])|(m[22]&m[364]&~m[365]&~m[366]&m[367])|(m[22]&~m[364]&m[365]&~m[366]&m[367])|(~m[22]&m[364]&m[365]&~m[366]&m[367])|(m[22]&~m[364]&~m[365]&m[366]&m[367])|(~m[22]&m[364]&~m[365]&m[366]&m[367])|(~m[22]&~m[364]&m[365]&m[366]&m[367]))&~BiasedRNG[235])|((m[22]&m[364]&m[365]&m[366]&~m[367])|(m[22]&m[364]&m[365]&~m[366]&m[367])|(m[22]&m[364]&~m[365]&m[366]&m[367])|(m[22]&~m[364]&m[365]&m[366]&m[367])|(~m[22]&m[364]&m[365]&m[366]&m[367])|(m[22]&m[364]&m[365]&m[366]&m[367]))):InitCond[366];
    m[92] = run?((((m[22]&m[368]&~m[369]&~m[370]&~m[371])|(m[22]&~m[368]&m[369]&~m[370]&~m[371])|(~m[22]&m[368]&m[369]&~m[370]&~m[371])|(m[22]&~m[368]&~m[369]&m[370]&~m[371])|(~m[22]&m[368]&~m[369]&m[370]&~m[371])|(~m[22]&~m[368]&m[369]&m[370]&~m[371])|(m[22]&~m[368]&~m[369]&~m[370]&m[371])|(~m[22]&m[368]&~m[369]&~m[370]&m[371])|(~m[22]&~m[368]&m[369]&~m[370]&m[371])|(~m[22]&~m[368]&~m[369]&m[370]&m[371]))&BiasedRNG[236])|(((m[22]&m[368]&m[369]&~m[370]&~m[371])|(m[22]&m[368]&~m[369]&m[370]&~m[371])|(m[22]&~m[368]&m[369]&m[370]&~m[371])|(~m[22]&m[368]&m[369]&m[370]&~m[371])|(m[22]&m[368]&~m[369]&~m[370]&m[371])|(m[22]&~m[368]&m[369]&~m[370]&m[371])|(~m[22]&m[368]&m[369]&~m[370]&m[371])|(m[22]&~m[368]&~m[369]&m[370]&m[371])|(~m[22]&m[368]&~m[369]&m[370]&m[371])|(~m[22]&~m[368]&m[369]&m[370]&m[371]))&~BiasedRNG[236])|((m[22]&m[368]&m[369]&m[370]&~m[371])|(m[22]&m[368]&m[369]&~m[370]&m[371])|(m[22]&m[368]&~m[369]&m[370]&m[371])|(m[22]&~m[368]&m[369]&m[370]&m[371])|(~m[22]&m[368]&m[369]&m[370]&m[371])|(m[22]&m[368]&m[369]&m[370]&m[371]))):InitCond[367];
    m[93] = run?((((m[23]&m[372]&~m[373]&~m[374]&~m[375])|(m[23]&~m[372]&m[373]&~m[374]&~m[375])|(~m[23]&m[372]&m[373]&~m[374]&~m[375])|(m[23]&~m[372]&~m[373]&m[374]&~m[375])|(~m[23]&m[372]&~m[373]&m[374]&~m[375])|(~m[23]&~m[372]&m[373]&m[374]&~m[375])|(m[23]&~m[372]&~m[373]&~m[374]&m[375])|(~m[23]&m[372]&~m[373]&~m[374]&m[375])|(~m[23]&~m[372]&m[373]&~m[374]&m[375])|(~m[23]&~m[372]&~m[373]&m[374]&m[375]))&BiasedRNG[237])|(((m[23]&m[372]&m[373]&~m[374]&~m[375])|(m[23]&m[372]&~m[373]&m[374]&~m[375])|(m[23]&~m[372]&m[373]&m[374]&~m[375])|(~m[23]&m[372]&m[373]&m[374]&~m[375])|(m[23]&m[372]&~m[373]&~m[374]&m[375])|(m[23]&~m[372]&m[373]&~m[374]&m[375])|(~m[23]&m[372]&m[373]&~m[374]&m[375])|(m[23]&~m[372]&~m[373]&m[374]&m[375])|(~m[23]&m[372]&~m[373]&m[374]&m[375])|(~m[23]&~m[372]&m[373]&m[374]&m[375]))&~BiasedRNG[237])|((m[23]&m[372]&m[373]&m[374]&~m[375])|(m[23]&m[372]&m[373]&~m[374]&m[375])|(m[23]&m[372]&~m[373]&m[374]&m[375])|(m[23]&~m[372]&m[373]&m[374]&m[375])|(~m[23]&m[372]&m[373]&m[374]&m[375])|(m[23]&m[372]&m[373]&m[374]&m[375]))):InitCond[368];
    m[94] = run?((((m[23]&m[376]&~m[377]&~m[378]&~m[379])|(m[23]&~m[376]&m[377]&~m[378]&~m[379])|(~m[23]&m[376]&m[377]&~m[378]&~m[379])|(m[23]&~m[376]&~m[377]&m[378]&~m[379])|(~m[23]&m[376]&~m[377]&m[378]&~m[379])|(~m[23]&~m[376]&m[377]&m[378]&~m[379])|(m[23]&~m[376]&~m[377]&~m[378]&m[379])|(~m[23]&m[376]&~m[377]&~m[378]&m[379])|(~m[23]&~m[376]&m[377]&~m[378]&m[379])|(~m[23]&~m[376]&~m[377]&m[378]&m[379]))&BiasedRNG[238])|(((m[23]&m[376]&m[377]&~m[378]&~m[379])|(m[23]&m[376]&~m[377]&m[378]&~m[379])|(m[23]&~m[376]&m[377]&m[378]&~m[379])|(~m[23]&m[376]&m[377]&m[378]&~m[379])|(m[23]&m[376]&~m[377]&~m[378]&m[379])|(m[23]&~m[376]&m[377]&~m[378]&m[379])|(~m[23]&m[376]&m[377]&~m[378]&m[379])|(m[23]&~m[376]&~m[377]&m[378]&m[379])|(~m[23]&m[376]&~m[377]&m[378]&m[379])|(~m[23]&~m[376]&m[377]&m[378]&m[379]))&~BiasedRNG[238])|((m[23]&m[376]&m[377]&m[378]&~m[379])|(m[23]&m[376]&m[377]&~m[378]&m[379])|(m[23]&m[376]&~m[377]&m[378]&m[379])|(m[23]&~m[376]&m[377]&m[378]&m[379])|(~m[23]&m[376]&m[377]&m[378]&m[379])|(m[23]&m[376]&m[377]&m[378]&m[379]))):InitCond[369];
    m[95] = run?((((m[23]&m[380]&~m[381]&~m[382]&~m[383])|(m[23]&~m[380]&m[381]&~m[382]&~m[383])|(~m[23]&m[380]&m[381]&~m[382]&~m[383])|(m[23]&~m[380]&~m[381]&m[382]&~m[383])|(~m[23]&m[380]&~m[381]&m[382]&~m[383])|(~m[23]&~m[380]&m[381]&m[382]&~m[383])|(m[23]&~m[380]&~m[381]&~m[382]&m[383])|(~m[23]&m[380]&~m[381]&~m[382]&m[383])|(~m[23]&~m[380]&m[381]&~m[382]&m[383])|(~m[23]&~m[380]&~m[381]&m[382]&m[383]))&BiasedRNG[239])|(((m[23]&m[380]&m[381]&~m[382]&~m[383])|(m[23]&m[380]&~m[381]&m[382]&~m[383])|(m[23]&~m[380]&m[381]&m[382]&~m[383])|(~m[23]&m[380]&m[381]&m[382]&~m[383])|(m[23]&m[380]&~m[381]&~m[382]&m[383])|(m[23]&~m[380]&m[381]&~m[382]&m[383])|(~m[23]&m[380]&m[381]&~m[382]&m[383])|(m[23]&~m[380]&~m[381]&m[382]&m[383])|(~m[23]&m[380]&~m[381]&m[382]&m[383])|(~m[23]&~m[380]&m[381]&m[382]&m[383]))&~BiasedRNG[239])|((m[23]&m[380]&m[381]&m[382]&~m[383])|(m[23]&m[380]&m[381]&~m[382]&m[383])|(m[23]&m[380]&~m[381]&m[382]&m[383])|(m[23]&~m[380]&m[381]&m[382]&m[383])|(~m[23]&m[380]&m[381]&m[382]&m[383])|(m[23]&m[380]&m[381]&m[382]&m[383]))):InitCond[370];
    m[385] = run?((((m[108]&~m[241]&m[528])|(~m[108]&m[241]&m[528]))&BiasedRNG[240])|(((m[108]&m[241]&~m[528]))&~BiasedRNG[240])|((m[108]&m[241]&m[528]))):InitCond[371];
    m[386] = run?((((m[120]&~m[242]&m[533])|(~m[120]&m[242]&m[533]))&BiasedRNG[241])|(((m[120]&m[242]&~m[533]))&~BiasedRNG[241])|((m[120]&m[242]&m[533]))):InitCond[372];
    m[387] = run?((((m[132]&~m[243]&m[543])|(~m[132]&m[243]&m[543]))&BiasedRNG[242])|(((m[132]&m[243]&~m[543]))&~BiasedRNG[242])|((m[132]&m[243]&m[543]))):InitCond[373];
    m[388] = run?((((m[144]&~m[244]&m[558])|(~m[144]&m[244]&m[558]))&BiasedRNG[243])|(((m[144]&m[244]&~m[558]))&~BiasedRNG[243])|((m[144]&m[244]&m[558]))):InitCond[374];
    m[389] = run?((((m[156]&~m[245]&m[578])|(~m[156]&m[245]&m[578]))&BiasedRNG[244])|(((m[156]&m[245]&~m[578]))&~BiasedRNG[244])|((m[156]&m[245]&m[578]))):InitCond[375];
    m[390] = run?((((m[168]&~m[246]&m[603])|(~m[168]&m[246]&m[603]))&BiasedRNG[245])|(((m[168]&m[246]&~m[603]))&~BiasedRNG[245])|((m[168]&m[246]&m[603]))):InitCond[376];
    m[391] = run?((((m[180]&~m[247]&m[633])|(~m[180]&m[247]&m[633]))&BiasedRNG[246])|(((m[180]&m[247]&~m[633]))&~BiasedRNG[246])|((m[180]&m[247]&m[633]))):InitCond[377];
    m[392] = run?((((m[192]&~m[248]&m[668])|(~m[192]&m[248]&m[668]))&BiasedRNG[247])|(((m[192]&m[248]&~m[668]))&~BiasedRNG[247])|((m[192]&m[248]&m[668]))):InitCond[378];
    m[393] = run?((((m[204]&~m[249]&m[708])|(~m[204]&m[249]&m[708]))&BiasedRNG[248])|(((m[204]&m[249]&~m[708]))&~BiasedRNG[248])|((m[204]&m[249]&m[708]))):InitCond[379];
    m[394] = run?((((m[216]&~m[250]&m[753])|(~m[216]&m[250]&m[753]))&BiasedRNG[249])|(((m[216]&m[250]&~m[753]))&~BiasedRNG[249])|((m[216]&m[250]&m[753]))):InitCond[380];
    m[395] = run?((((m[228]&~m[251]&m[803])|(~m[228]&m[251]&m[803]))&BiasedRNG[250])|(((m[228]&m[251]&~m[803]))&~BiasedRNG[250])|((m[228]&m[251]&m[803]))):InitCond[381];
    m[396] = run?((((m[97]&~m[252]&m[529])|(~m[97]&m[252]&m[529]))&BiasedRNG[251])|(((m[97]&m[252]&~m[529]))&~BiasedRNG[251])|((m[97]&m[252]&m[529]))):InitCond[382];
    m[397] = run?((((m[109]&~m[253]&m[534])|(~m[109]&m[253]&m[534]))&BiasedRNG[252])|(((m[109]&m[253]&~m[534]))&~BiasedRNG[252])|((m[109]&m[253]&m[534]))):InitCond[383];
    m[398] = run?((((m[121]&~m[254]&m[544])|(~m[121]&m[254]&m[544]))&BiasedRNG[253])|(((m[121]&m[254]&~m[544]))&~BiasedRNG[253])|((m[121]&m[254]&m[544]))):InitCond[384];
    m[399] = run?((((m[133]&~m[255]&m[559])|(~m[133]&m[255]&m[559]))&BiasedRNG[254])|(((m[133]&m[255]&~m[559]))&~BiasedRNG[254])|((m[133]&m[255]&m[559]))):InitCond[385];
    m[400] = run?((((m[145]&~m[256]&m[579])|(~m[145]&m[256]&m[579]))&BiasedRNG[255])|(((m[145]&m[256]&~m[579]))&~BiasedRNG[255])|((m[145]&m[256]&m[579]))):InitCond[386];
    m[401] = run?((((m[157]&~m[257]&m[604])|(~m[157]&m[257]&m[604]))&BiasedRNG[256])|(((m[157]&m[257]&~m[604]))&~BiasedRNG[256])|((m[157]&m[257]&m[604]))):InitCond[387];
    m[402] = run?((((m[169]&~m[258]&m[634])|(~m[169]&m[258]&m[634]))&BiasedRNG[257])|(((m[169]&m[258]&~m[634]))&~BiasedRNG[257])|((m[169]&m[258]&m[634]))):InitCond[388];
    m[403] = run?((((m[181]&~m[259]&m[669])|(~m[181]&m[259]&m[669]))&BiasedRNG[258])|(((m[181]&m[259]&~m[669]))&~BiasedRNG[258])|((m[181]&m[259]&m[669]))):InitCond[389];
    m[404] = run?((((m[193]&~m[260]&m[709])|(~m[193]&m[260]&m[709]))&BiasedRNG[259])|(((m[193]&m[260]&~m[709]))&~BiasedRNG[259])|((m[193]&m[260]&m[709]))):InitCond[390];
    m[405] = run?((((m[205]&~m[261]&m[754])|(~m[205]&m[261]&m[754]))&BiasedRNG[260])|(((m[205]&m[261]&~m[754]))&~BiasedRNG[260])|((m[205]&m[261]&m[754]))):InitCond[391];
    m[406] = run?((((m[217]&~m[262]&m[804])|(~m[217]&m[262]&m[804]))&BiasedRNG[261])|(((m[217]&m[262]&~m[804]))&~BiasedRNG[261])|((m[217]&m[262]&m[804]))):InitCond[392];
    m[407] = run?((((m[229]&~m[263]&m[859])|(~m[229]&m[263]&m[859]))&BiasedRNG[262])|(((m[229]&m[263]&~m[859]))&~BiasedRNG[262])|((m[229]&m[263]&m[859]))):InitCond[393];
    m[408] = run?((((m[98]&~m[264]&m[539])|(~m[98]&m[264]&m[539]))&BiasedRNG[263])|(((m[98]&m[264]&~m[539]))&~BiasedRNG[263])|((m[98]&m[264]&m[539]))):InitCond[394];
    m[409] = run?((((m[110]&~m[265]&m[549])|(~m[110]&m[265]&m[549]))&BiasedRNG[264])|(((m[110]&m[265]&~m[549]))&~BiasedRNG[264])|((m[110]&m[265]&m[549]))):InitCond[395];
    m[410] = run?((((m[122]&~m[266]&m[564])|(~m[122]&m[266]&m[564]))&BiasedRNG[265])|(((m[122]&m[266]&~m[564]))&~BiasedRNG[265])|((m[122]&m[266]&m[564]))):InitCond[396];
    m[411] = run?((((m[134]&~m[267]&m[584])|(~m[134]&m[267]&m[584]))&BiasedRNG[266])|(((m[134]&m[267]&~m[584]))&~BiasedRNG[266])|((m[134]&m[267]&m[584]))):InitCond[397];
    m[412] = run?((((m[146]&~m[268]&m[609])|(~m[146]&m[268]&m[609]))&BiasedRNG[267])|(((m[146]&m[268]&~m[609]))&~BiasedRNG[267])|((m[146]&m[268]&m[609]))):InitCond[398];
    m[413] = run?((((m[158]&~m[269]&m[639])|(~m[158]&m[269]&m[639]))&BiasedRNG[268])|(((m[158]&m[269]&~m[639]))&~BiasedRNG[268])|((m[158]&m[269]&m[639]))):InitCond[399];
    m[414] = run?((((m[170]&~m[270]&m[674])|(~m[170]&m[270]&m[674]))&BiasedRNG[269])|(((m[170]&m[270]&~m[674]))&~BiasedRNG[269])|((m[170]&m[270]&m[674]))):InitCond[400];
    m[415] = run?((((m[182]&~m[271]&m[714])|(~m[182]&m[271]&m[714]))&BiasedRNG[270])|(((m[182]&m[271]&~m[714]))&~BiasedRNG[270])|((m[182]&m[271]&m[714]))):InitCond[401];
    m[416] = run?((((m[194]&~m[272]&m[759])|(~m[194]&m[272]&m[759]))&BiasedRNG[271])|(((m[194]&m[272]&~m[759]))&~BiasedRNG[271])|((m[194]&m[272]&m[759]))):InitCond[402];
    m[417] = run?((((m[206]&~m[273]&m[809])|(~m[206]&m[273]&m[809]))&BiasedRNG[272])|(((m[206]&m[273]&~m[809]))&~BiasedRNG[272])|((m[206]&m[273]&m[809]))):InitCond[403];
    m[418] = run?((((m[218]&~m[274]&m[864])|(~m[218]&m[274]&m[864]))&BiasedRNG[273])|(((m[218]&m[274]&~m[864]))&~BiasedRNG[273])|((m[218]&m[274]&m[864]))):InitCond[404];
    m[419] = run?((((m[230]&~m[275]&m[914])|(~m[230]&m[275]&m[914]))&BiasedRNG[274])|(((m[230]&m[275]&~m[914]))&~BiasedRNG[274])|((m[230]&m[275]&m[914]))):InitCond[405];
    m[420] = run?((((m[99]&~m[276]&m[554])|(~m[99]&m[276]&m[554]))&BiasedRNG[275])|(((m[99]&m[276]&~m[554]))&~BiasedRNG[275])|((m[99]&m[276]&m[554]))):InitCond[406];
    m[421] = run?((((m[111]&~m[277]&m[569])|(~m[111]&m[277]&m[569]))&BiasedRNG[276])|(((m[111]&m[277]&~m[569]))&~BiasedRNG[276])|((m[111]&m[277]&m[569]))):InitCond[407];
    m[422] = run?((((m[123]&~m[278]&m[589])|(~m[123]&m[278]&m[589]))&BiasedRNG[277])|(((m[123]&m[278]&~m[589]))&~BiasedRNG[277])|((m[123]&m[278]&m[589]))):InitCond[408];
    m[423] = run?((((m[135]&~m[279]&m[614])|(~m[135]&m[279]&m[614]))&BiasedRNG[278])|(((m[135]&m[279]&~m[614]))&~BiasedRNG[278])|((m[135]&m[279]&m[614]))):InitCond[409];
    m[424] = run?((((m[147]&~m[280]&m[644])|(~m[147]&m[280]&m[644]))&BiasedRNG[279])|(((m[147]&m[280]&~m[644]))&~BiasedRNG[279])|((m[147]&m[280]&m[644]))):InitCond[410];
    m[425] = run?((((m[159]&~m[281]&m[679])|(~m[159]&m[281]&m[679]))&BiasedRNG[280])|(((m[159]&m[281]&~m[679]))&~BiasedRNG[280])|((m[159]&m[281]&m[679]))):InitCond[411];
    m[426] = run?((((m[171]&~m[282]&m[719])|(~m[171]&m[282]&m[719]))&BiasedRNG[281])|(((m[171]&m[282]&~m[719]))&~BiasedRNG[281])|((m[171]&m[282]&m[719]))):InitCond[412];
    m[427] = run?((((m[183]&~m[283]&m[764])|(~m[183]&m[283]&m[764]))&BiasedRNG[282])|(((m[183]&m[283]&~m[764]))&~BiasedRNG[282])|((m[183]&m[283]&m[764]))):InitCond[413];
    m[428] = run?((((m[195]&~m[284]&m[814])|(~m[195]&m[284]&m[814]))&BiasedRNG[283])|(((m[195]&m[284]&~m[814]))&~BiasedRNG[283])|((m[195]&m[284]&m[814]))):InitCond[414];
    m[429] = run?((((m[207]&~m[285]&m[869])|(~m[207]&m[285]&m[869]))&BiasedRNG[284])|(((m[207]&m[285]&~m[869]))&~BiasedRNG[284])|((m[207]&m[285]&m[869]))):InitCond[415];
    m[430] = run?((((m[219]&~m[286]&m[919])|(~m[219]&m[286]&m[919]))&BiasedRNG[285])|(((m[219]&m[286]&~m[919]))&~BiasedRNG[285])|((m[219]&m[286]&m[919]))):InitCond[416];
    m[431] = run?((((m[231]&~m[287]&m[964])|(~m[231]&m[287]&m[964]))&BiasedRNG[286])|(((m[231]&m[287]&~m[964]))&~BiasedRNG[286])|((m[231]&m[287]&m[964]))):InitCond[417];
    m[432] = run?((((m[100]&~m[288]&m[574])|(~m[100]&m[288]&m[574]))&BiasedRNG[287])|(((m[100]&m[288]&~m[574]))&~BiasedRNG[287])|((m[100]&m[288]&m[574]))):InitCond[418];
    m[433] = run?((((m[112]&~m[289]&m[594])|(~m[112]&m[289]&m[594]))&BiasedRNG[288])|(((m[112]&m[289]&~m[594]))&~BiasedRNG[288])|((m[112]&m[289]&m[594]))):InitCond[419];
    m[434] = run?((((m[124]&~m[290]&m[619])|(~m[124]&m[290]&m[619]))&BiasedRNG[289])|(((m[124]&m[290]&~m[619]))&~BiasedRNG[289])|((m[124]&m[290]&m[619]))):InitCond[420];
    m[435] = run?((((m[136]&~m[291]&m[649])|(~m[136]&m[291]&m[649]))&BiasedRNG[290])|(((m[136]&m[291]&~m[649]))&~BiasedRNG[290])|((m[136]&m[291]&m[649]))):InitCond[421];
    m[436] = run?((((m[148]&~m[292]&m[684])|(~m[148]&m[292]&m[684]))&BiasedRNG[291])|(((m[148]&m[292]&~m[684]))&~BiasedRNG[291])|((m[148]&m[292]&m[684]))):InitCond[422];
    m[437] = run?((((m[160]&~m[293]&m[724])|(~m[160]&m[293]&m[724]))&BiasedRNG[292])|(((m[160]&m[293]&~m[724]))&~BiasedRNG[292])|((m[160]&m[293]&m[724]))):InitCond[423];
    m[438] = run?((((m[172]&~m[294]&m[769])|(~m[172]&m[294]&m[769]))&BiasedRNG[293])|(((m[172]&m[294]&~m[769]))&~BiasedRNG[293])|((m[172]&m[294]&m[769]))):InitCond[424];
    m[439] = run?((((m[184]&~m[295]&m[819])|(~m[184]&m[295]&m[819]))&BiasedRNG[294])|(((m[184]&m[295]&~m[819]))&~BiasedRNG[294])|((m[184]&m[295]&m[819]))):InitCond[425];
    m[440] = run?((((m[196]&~m[296]&m[874])|(~m[196]&m[296]&m[874]))&BiasedRNG[295])|(((m[196]&m[296]&~m[874]))&~BiasedRNG[295])|((m[196]&m[296]&m[874]))):InitCond[426];
    m[441] = run?((((m[208]&~m[297]&m[924])|(~m[208]&m[297]&m[924]))&BiasedRNG[296])|(((m[208]&m[297]&~m[924]))&~BiasedRNG[296])|((m[208]&m[297]&m[924]))):InitCond[427];
    m[442] = run?((((m[220]&~m[298]&m[969])|(~m[220]&m[298]&m[969]))&BiasedRNG[297])|(((m[220]&m[298]&~m[969]))&~BiasedRNG[297])|((m[220]&m[298]&m[969]))):InitCond[428];
    m[443] = run?((((m[232]&~m[299]&m[1009])|(~m[232]&m[299]&m[1009]))&BiasedRNG[298])|(((m[232]&m[299]&~m[1009]))&~BiasedRNG[298])|((m[232]&m[299]&m[1009]))):InitCond[429];
    m[444] = run?((((m[101]&~m[300]&m[599])|(~m[101]&m[300]&m[599]))&BiasedRNG[299])|(((m[101]&m[300]&~m[599]))&~BiasedRNG[299])|((m[101]&m[300]&m[599]))):InitCond[430];
    m[445] = run?((((m[113]&~m[301]&m[624])|(~m[113]&m[301]&m[624]))&BiasedRNG[300])|(((m[113]&m[301]&~m[624]))&~BiasedRNG[300])|((m[113]&m[301]&m[624]))):InitCond[431];
    m[446] = run?((((m[125]&~m[302]&m[654])|(~m[125]&m[302]&m[654]))&BiasedRNG[301])|(((m[125]&m[302]&~m[654]))&~BiasedRNG[301])|((m[125]&m[302]&m[654]))):InitCond[432];
    m[447] = run?((((m[137]&~m[303]&m[689])|(~m[137]&m[303]&m[689]))&BiasedRNG[302])|(((m[137]&m[303]&~m[689]))&~BiasedRNG[302])|((m[137]&m[303]&m[689]))):InitCond[433];
    m[448] = run?((((m[149]&~m[304]&m[729])|(~m[149]&m[304]&m[729]))&BiasedRNG[303])|(((m[149]&m[304]&~m[729]))&~BiasedRNG[303])|((m[149]&m[304]&m[729]))):InitCond[434];
    m[449] = run?((((m[161]&~m[305]&m[774])|(~m[161]&m[305]&m[774]))&BiasedRNG[304])|(((m[161]&m[305]&~m[774]))&~BiasedRNG[304])|((m[161]&m[305]&m[774]))):InitCond[435];
    m[450] = run?((((m[173]&~m[306]&m[824])|(~m[173]&m[306]&m[824]))&BiasedRNG[305])|(((m[173]&m[306]&~m[824]))&~BiasedRNG[305])|((m[173]&m[306]&m[824]))):InitCond[436];
    m[451] = run?((((m[185]&~m[307]&m[879])|(~m[185]&m[307]&m[879]))&BiasedRNG[306])|(((m[185]&m[307]&~m[879]))&~BiasedRNG[306])|((m[185]&m[307]&m[879]))):InitCond[437];
    m[452] = run?((((m[197]&~m[308]&m[929])|(~m[197]&m[308]&m[929]))&BiasedRNG[307])|(((m[197]&m[308]&~m[929]))&~BiasedRNG[307])|((m[197]&m[308]&m[929]))):InitCond[438];
    m[453] = run?((((m[209]&~m[309]&m[974])|(~m[209]&m[309]&m[974]))&BiasedRNG[308])|(((m[209]&m[309]&~m[974]))&~BiasedRNG[308])|((m[209]&m[309]&m[974]))):InitCond[439];
    m[454] = run?((((m[221]&~m[310]&m[1014])|(~m[221]&m[310]&m[1014]))&BiasedRNG[309])|(((m[221]&m[310]&~m[1014]))&~BiasedRNG[309])|((m[221]&m[310]&m[1014]))):InitCond[440];
    m[455] = run?((((m[233]&~m[311]&m[1049])|(~m[233]&m[311]&m[1049]))&BiasedRNG[310])|(((m[233]&m[311]&~m[1049]))&~BiasedRNG[310])|((m[233]&m[311]&m[1049]))):InitCond[441];
    m[456] = run?((((m[102]&~m[312]&m[629])|(~m[102]&m[312]&m[629]))&BiasedRNG[311])|(((m[102]&m[312]&~m[629]))&~BiasedRNG[311])|((m[102]&m[312]&m[629]))):InitCond[442];
    m[457] = run?((((m[114]&~m[313]&m[659])|(~m[114]&m[313]&m[659]))&BiasedRNG[312])|(((m[114]&m[313]&~m[659]))&~BiasedRNG[312])|((m[114]&m[313]&m[659]))):InitCond[443];
    m[458] = run?((((m[126]&~m[314]&m[694])|(~m[126]&m[314]&m[694]))&BiasedRNG[313])|(((m[126]&m[314]&~m[694]))&~BiasedRNG[313])|((m[126]&m[314]&m[694]))):InitCond[444];
    m[459] = run?((((m[138]&~m[315]&m[734])|(~m[138]&m[315]&m[734]))&BiasedRNG[314])|(((m[138]&m[315]&~m[734]))&~BiasedRNG[314])|((m[138]&m[315]&m[734]))):InitCond[445];
    m[460] = run?((((m[150]&~m[316]&m[779])|(~m[150]&m[316]&m[779]))&BiasedRNG[315])|(((m[150]&m[316]&~m[779]))&~BiasedRNG[315])|((m[150]&m[316]&m[779]))):InitCond[446];
    m[461] = run?((((m[162]&~m[317]&m[829])|(~m[162]&m[317]&m[829]))&BiasedRNG[316])|(((m[162]&m[317]&~m[829]))&~BiasedRNG[316])|((m[162]&m[317]&m[829]))):InitCond[447];
    m[462] = run?((((m[174]&~m[318]&m[884])|(~m[174]&m[318]&m[884]))&BiasedRNG[317])|(((m[174]&m[318]&~m[884]))&~BiasedRNG[317])|((m[174]&m[318]&m[884]))):InitCond[448];
    m[463] = run?((((m[186]&~m[319]&m[934])|(~m[186]&m[319]&m[934]))&BiasedRNG[318])|(((m[186]&m[319]&~m[934]))&~BiasedRNG[318])|((m[186]&m[319]&m[934]))):InitCond[449];
    m[464] = run?((((m[198]&~m[320]&m[979])|(~m[198]&m[320]&m[979]))&BiasedRNG[319])|(((m[198]&m[320]&~m[979]))&~BiasedRNG[319])|((m[198]&m[320]&m[979]))):InitCond[450];
    m[465] = run?((((m[210]&~m[321]&m[1019])|(~m[210]&m[321]&m[1019]))&BiasedRNG[320])|(((m[210]&m[321]&~m[1019]))&~BiasedRNG[320])|((m[210]&m[321]&m[1019]))):InitCond[451];
    m[466] = run?((((m[222]&~m[322]&m[1054])|(~m[222]&m[322]&m[1054]))&BiasedRNG[321])|(((m[222]&m[322]&~m[1054]))&~BiasedRNG[321])|((m[222]&m[322]&m[1054]))):InitCond[452];
    m[467] = run?((((m[234]&~m[323]&m[1084])|(~m[234]&m[323]&m[1084]))&BiasedRNG[322])|(((m[234]&m[323]&~m[1084]))&~BiasedRNG[322])|((m[234]&m[323]&m[1084]))):InitCond[453];
    m[468] = run?((((m[103]&~m[324]&m[664])|(~m[103]&m[324]&m[664]))&BiasedRNG[323])|(((m[103]&m[324]&~m[664]))&~BiasedRNG[323])|((m[103]&m[324]&m[664]))):InitCond[454];
    m[469] = run?((((m[115]&~m[325]&m[699])|(~m[115]&m[325]&m[699]))&BiasedRNG[324])|(((m[115]&m[325]&~m[699]))&~BiasedRNG[324])|((m[115]&m[325]&m[699]))):InitCond[455];
    m[470] = run?((((m[127]&~m[326]&m[739])|(~m[127]&m[326]&m[739]))&BiasedRNG[325])|(((m[127]&m[326]&~m[739]))&~BiasedRNG[325])|((m[127]&m[326]&m[739]))):InitCond[456];
    m[471] = run?((((m[139]&~m[327]&m[784])|(~m[139]&m[327]&m[784]))&BiasedRNG[326])|(((m[139]&m[327]&~m[784]))&~BiasedRNG[326])|((m[139]&m[327]&m[784]))):InitCond[457];
    m[472] = run?((((m[151]&~m[328]&m[834])|(~m[151]&m[328]&m[834]))&BiasedRNG[327])|(((m[151]&m[328]&~m[834]))&~BiasedRNG[327])|((m[151]&m[328]&m[834]))):InitCond[458];
    m[473] = run?((((m[163]&~m[329]&m[889])|(~m[163]&m[329]&m[889]))&BiasedRNG[328])|(((m[163]&m[329]&~m[889]))&~BiasedRNG[328])|((m[163]&m[329]&m[889]))):InitCond[459];
    m[474] = run?((((m[175]&~m[330]&m[939])|(~m[175]&m[330]&m[939]))&BiasedRNG[329])|(((m[175]&m[330]&~m[939]))&~BiasedRNG[329])|((m[175]&m[330]&m[939]))):InitCond[460];
    m[475] = run?((((m[187]&~m[331]&m[984])|(~m[187]&m[331]&m[984]))&BiasedRNG[330])|(((m[187]&m[331]&~m[984]))&~BiasedRNG[330])|((m[187]&m[331]&m[984]))):InitCond[461];
    m[476] = run?((((m[199]&~m[332]&m[1024])|(~m[199]&m[332]&m[1024]))&BiasedRNG[331])|(((m[199]&m[332]&~m[1024]))&~BiasedRNG[331])|((m[199]&m[332]&m[1024]))):InitCond[462];
    m[477] = run?((((m[211]&~m[333]&m[1059])|(~m[211]&m[333]&m[1059]))&BiasedRNG[332])|(((m[211]&m[333]&~m[1059]))&~BiasedRNG[332])|((m[211]&m[333]&m[1059]))):InitCond[463];
    m[478] = run?((((m[223]&~m[334]&m[1089])|(~m[223]&m[334]&m[1089]))&BiasedRNG[333])|(((m[223]&m[334]&~m[1089]))&~BiasedRNG[333])|((m[223]&m[334]&m[1089]))):InitCond[464];
    m[479] = run?((((m[235]&~m[335]&m[1114])|(~m[235]&m[335]&m[1114]))&BiasedRNG[334])|(((m[235]&m[335]&~m[1114]))&~BiasedRNG[334])|((m[235]&m[335]&m[1114]))):InitCond[465];
    m[480] = run?((((m[104]&~m[336]&m[704])|(~m[104]&m[336]&m[704]))&BiasedRNG[335])|(((m[104]&m[336]&~m[704]))&~BiasedRNG[335])|((m[104]&m[336]&m[704]))):InitCond[466];
    m[481] = run?((((m[116]&~m[337]&m[744])|(~m[116]&m[337]&m[744]))&BiasedRNG[336])|(((m[116]&m[337]&~m[744]))&~BiasedRNG[336])|((m[116]&m[337]&m[744]))):InitCond[467];
    m[482] = run?((((m[128]&~m[338]&m[789])|(~m[128]&m[338]&m[789]))&BiasedRNG[337])|(((m[128]&m[338]&~m[789]))&~BiasedRNG[337])|((m[128]&m[338]&m[789]))):InitCond[468];
    m[483] = run?((((m[140]&~m[339]&m[839])|(~m[140]&m[339]&m[839]))&BiasedRNG[338])|(((m[140]&m[339]&~m[839]))&~BiasedRNG[338])|((m[140]&m[339]&m[839]))):InitCond[469];
    m[484] = run?((((m[152]&~m[340]&m[894])|(~m[152]&m[340]&m[894]))&BiasedRNG[339])|(((m[152]&m[340]&~m[894]))&~BiasedRNG[339])|((m[152]&m[340]&m[894]))):InitCond[470];
    m[485] = run?((((m[164]&~m[341]&m[944])|(~m[164]&m[341]&m[944]))&BiasedRNG[340])|(((m[164]&m[341]&~m[944]))&~BiasedRNG[340])|((m[164]&m[341]&m[944]))):InitCond[471];
    m[486] = run?((((m[176]&~m[342]&m[989])|(~m[176]&m[342]&m[989]))&BiasedRNG[341])|(((m[176]&m[342]&~m[989]))&~BiasedRNG[341])|((m[176]&m[342]&m[989]))):InitCond[472];
    m[487] = run?((((m[188]&~m[343]&m[1029])|(~m[188]&m[343]&m[1029]))&BiasedRNG[342])|(((m[188]&m[343]&~m[1029]))&~BiasedRNG[342])|((m[188]&m[343]&m[1029]))):InitCond[473];
    m[488] = run?((((m[200]&~m[344]&m[1064])|(~m[200]&m[344]&m[1064]))&BiasedRNG[343])|(((m[200]&m[344]&~m[1064]))&~BiasedRNG[343])|((m[200]&m[344]&m[1064]))):InitCond[474];
    m[489] = run?((((m[212]&~m[345]&m[1094])|(~m[212]&m[345]&m[1094]))&BiasedRNG[344])|(((m[212]&m[345]&~m[1094]))&~BiasedRNG[344])|((m[212]&m[345]&m[1094]))):InitCond[475];
    m[490] = run?((((m[224]&~m[346]&m[1119])|(~m[224]&m[346]&m[1119]))&BiasedRNG[345])|(((m[224]&m[346]&~m[1119]))&~BiasedRNG[345])|((m[224]&m[346]&m[1119]))):InitCond[476];
    m[491] = run?((((m[236]&~m[347]&m[1139])|(~m[236]&m[347]&m[1139]))&BiasedRNG[346])|(((m[236]&m[347]&~m[1139]))&~BiasedRNG[346])|((m[236]&m[347]&m[1139]))):InitCond[477];
    m[492] = run?((((m[105]&~m[348]&m[749])|(~m[105]&m[348]&m[749]))&BiasedRNG[347])|(((m[105]&m[348]&~m[749]))&~BiasedRNG[347])|((m[105]&m[348]&m[749]))):InitCond[478];
    m[493] = run?((((m[117]&~m[349]&m[794])|(~m[117]&m[349]&m[794]))&BiasedRNG[348])|(((m[117]&m[349]&~m[794]))&~BiasedRNG[348])|((m[117]&m[349]&m[794]))):InitCond[479];
    m[494] = run?((((m[129]&~m[350]&m[844])|(~m[129]&m[350]&m[844]))&BiasedRNG[349])|(((m[129]&m[350]&~m[844]))&~BiasedRNG[349])|((m[129]&m[350]&m[844]))):InitCond[480];
    m[495] = run?((((m[141]&~m[351]&m[899])|(~m[141]&m[351]&m[899]))&BiasedRNG[350])|(((m[141]&m[351]&~m[899]))&~BiasedRNG[350])|((m[141]&m[351]&m[899]))):InitCond[481];
    m[496] = run?((((m[153]&~m[352]&m[949])|(~m[153]&m[352]&m[949]))&BiasedRNG[351])|(((m[153]&m[352]&~m[949]))&~BiasedRNG[351])|((m[153]&m[352]&m[949]))):InitCond[482];
    m[497] = run?((((m[165]&~m[353]&m[994])|(~m[165]&m[353]&m[994]))&BiasedRNG[352])|(((m[165]&m[353]&~m[994]))&~BiasedRNG[352])|((m[165]&m[353]&m[994]))):InitCond[483];
    m[498] = run?((((m[177]&~m[354]&m[1034])|(~m[177]&m[354]&m[1034]))&BiasedRNG[353])|(((m[177]&m[354]&~m[1034]))&~BiasedRNG[353])|((m[177]&m[354]&m[1034]))):InitCond[484];
    m[499] = run?((((m[189]&~m[355]&m[1069])|(~m[189]&m[355]&m[1069]))&BiasedRNG[354])|(((m[189]&m[355]&~m[1069]))&~BiasedRNG[354])|((m[189]&m[355]&m[1069]))):InitCond[485];
    m[500] = run?((((m[201]&~m[356]&m[1099])|(~m[201]&m[356]&m[1099]))&BiasedRNG[355])|(((m[201]&m[356]&~m[1099]))&~BiasedRNG[355])|((m[201]&m[356]&m[1099]))):InitCond[486];
    m[501] = run?((((m[213]&~m[357]&m[1124])|(~m[213]&m[357]&m[1124]))&BiasedRNG[356])|(((m[213]&m[357]&~m[1124]))&~BiasedRNG[356])|((m[213]&m[357]&m[1124]))):InitCond[487];
    m[502] = run?((((m[225]&~m[358]&m[1144])|(~m[225]&m[358]&m[1144]))&BiasedRNG[357])|(((m[225]&m[358]&~m[1144]))&~BiasedRNG[357])|((m[225]&m[358]&m[1144]))):InitCond[488];
    m[503] = run?((((m[237]&~m[359]&m[1159])|(~m[237]&m[359]&m[1159]))&BiasedRNG[358])|(((m[237]&m[359]&~m[1159]))&~BiasedRNG[358])|((m[237]&m[359]&m[1159]))):InitCond[489];
    m[504] = run?((((m[106]&~m[360]&m[799])|(~m[106]&m[360]&m[799]))&BiasedRNG[359])|(((m[106]&m[360]&~m[799]))&~BiasedRNG[359])|((m[106]&m[360]&m[799]))):InitCond[490];
    m[505] = run?((((m[118]&~m[361]&m[849])|(~m[118]&m[361]&m[849]))&BiasedRNG[360])|(((m[118]&m[361]&~m[849]))&~BiasedRNG[360])|((m[118]&m[361]&m[849]))):InitCond[491];
    m[506] = run?((((m[130]&~m[362]&m[904])|(~m[130]&m[362]&m[904]))&BiasedRNG[361])|(((m[130]&m[362]&~m[904]))&~BiasedRNG[361])|((m[130]&m[362]&m[904]))):InitCond[492];
    m[507] = run?((((m[142]&~m[363]&m[954])|(~m[142]&m[363]&m[954]))&BiasedRNG[362])|(((m[142]&m[363]&~m[954]))&~BiasedRNG[362])|((m[142]&m[363]&m[954]))):InitCond[493];
    m[508] = run?((((m[154]&~m[364]&m[999])|(~m[154]&m[364]&m[999]))&BiasedRNG[363])|(((m[154]&m[364]&~m[999]))&~BiasedRNG[363])|((m[154]&m[364]&m[999]))):InitCond[494];
    m[509] = run?((((m[166]&~m[365]&m[1039])|(~m[166]&m[365]&m[1039]))&BiasedRNG[364])|(((m[166]&m[365]&~m[1039]))&~BiasedRNG[364])|((m[166]&m[365]&m[1039]))):InitCond[495];
    m[510] = run?((((m[178]&~m[366]&m[1074])|(~m[178]&m[366]&m[1074]))&BiasedRNG[365])|(((m[178]&m[366]&~m[1074]))&~BiasedRNG[365])|((m[178]&m[366]&m[1074]))):InitCond[496];
    m[511] = run?((((m[190]&~m[367]&m[1104])|(~m[190]&m[367]&m[1104]))&BiasedRNG[366])|(((m[190]&m[367]&~m[1104]))&~BiasedRNG[366])|((m[190]&m[367]&m[1104]))):InitCond[497];
    m[512] = run?((((m[202]&~m[368]&m[1129])|(~m[202]&m[368]&m[1129]))&BiasedRNG[367])|(((m[202]&m[368]&~m[1129]))&~BiasedRNG[367])|((m[202]&m[368]&m[1129]))):InitCond[498];
    m[513] = run?((((m[214]&~m[369]&m[1149])|(~m[214]&m[369]&m[1149]))&BiasedRNG[368])|(((m[214]&m[369]&~m[1149]))&~BiasedRNG[368])|((m[214]&m[369]&m[1149]))):InitCond[499];
    m[514] = run?((((m[226]&~m[370]&m[1164])|(~m[226]&m[370]&m[1164]))&BiasedRNG[369])|(((m[226]&m[370]&~m[1164]))&~BiasedRNG[369])|((m[226]&m[370]&m[1164]))):InitCond[500];
    m[515] = run?((((m[238]&~m[371]&m[1174])|(~m[238]&m[371]&m[1174]))&BiasedRNG[370])|(((m[238]&m[371]&~m[1174]))&~BiasedRNG[370])|((m[238]&m[371]&m[1174]))):InitCond[501];
    m[516] = run?((((m[107]&~m[372]&m[854])|(~m[107]&m[372]&m[854]))&BiasedRNG[371])|(((m[107]&m[372]&~m[854]))&~BiasedRNG[371])|((m[107]&m[372]&m[854]))):InitCond[502];
    m[517] = run?((((m[119]&~m[373]&m[909])|(~m[119]&m[373]&m[909]))&BiasedRNG[372])|(((m[119]&m[373]&~m[909]))&~BiasedRNG[372])|((m[119]&m[373]&m[909]))):InitCond[503];
    m[518] = run?((((m[131]&~m[374]&m[959])|(~m[131]&m[374]&m[959]))&BiasedRNG[373])|(((m[131]&m[374]&~m[959]))&~BiasedRNG[373])|((m[131]&m[374]&m[959]))):InitCond[504];
    m[519] = run?((((m[143]&~m[375]&m[1004])|(~m[143]&m[375]&m[1004]))&BiasedRNG[374])|(((m[143]&m[375]&~m[1004]))&~BiasedRNG[374])|((m[143]&m[375]&m[1004]))):InitCond[505];
    m[520] = run?((((m[155]&~m[376]&m[1044])|(~m[155]&m[376]&m[1044]))&BiasedRNG[375])|(((m[155]&m[376]&~m[1044]))&~BiasedRNG[375])|((m[155]&m[376]&m[1044]))):InitCond[506];
    m[521] = run?((((m[167]&~m[377]&m[1079])|(~m[167]&m[377]&m[1079]))&BiasedRNG[376])|(((m[167]&m[377]&~m[1079]))&~BiasedRNG[376])|((m[167]&m[377]&m[1079]))):InitCond[507];
    m[522] = run?((((m[179]&~m[378]&m[1109])|(~m[179]&m[378]&m[1109]))&BiasedRNG[377])|(((m[179]&m[378]&~m[1109]))&~BiasedRNG[377])|((m[179]&m[378]&m[1109]))):InitCond[508];
    m[523] = run?((((m[191]&~m[379]&m[1134])|(~m[191]&m[379]&m[1134]))&BiasedRNG[378])|(((m[191]&m[379]&~m[1134]))&~BiasedRNG[378])|((m[191]&m[379]&m[1134]))):InitCond[509];
    m[524] = run?((((m[203]&~m[380]&m[1154])|(~m[203]&m[380]&m[1154]))&BiasedRNG[379])|(((m[203]&m[380]&~m[1154]))&~BiasedRNG[379])|((m[203]&m[380]&m[1154]))):InitCond[510];
    m[525] = run?((((m[215]&~m[381]&m[1169])|(~m[215]&m[381]&m[1169]))&BiasedRNG[380])|(((m[215]&m[381]&~m[1169]))&~BiasedRNG[380])|((m[215]&m[381]&m[1169]))):InitCond[511];
    m[526] = run?((((m[227]&~m[382]&m[1179])|(~m[227]&m[382]&m[1179]))&BiasedRNG[381])|(((m[227]&m[382]&~m[1179]))&~BiasedRNG[381])|((m[227]&m[382]&m[1179]))):InitCond[512];
    m[527] = run?((((m[239]&~m[383]&m[1184])|(~m[239]&m[383]&m[1184]))&BiasedRNG[382])|(((m[239]&m[383]&~m[1184]))&~BiasedRNG[382])|((m[239]&m[383]&m[1184]))):InitCond[513];
    m[535] = run?((((m[532]&~m[533]&~m[534]&~m[536]&~m[537])|(~m[532]&~m[533]&~m[534]&m[536]&~m[537])|(m[532]&m[533]&~m[534]&m[536]&~m[537])|(m[532]&~m[533]&m[534]&m[536]&~m[537])|(~m[532]&m[533]&~m[534]&~m[536]&m[537])|(~m[532]&~m[533]&m[534]&~m[536]&m[537])|(m[532]&m[533]&m[534]&~m[536]&m[537])|(~m[532]&m[533]&m[534]&m[536]&m[537]))&UnbiasedRNG[131])|((m[532]&~m[533]&~m[534]&m[536]&~m[537])|(~m[532]&~m[533]&~m[534]&~m[536]&m[537])|(m[532]&~m[533]&~m[534]&~m[536]&m[537])|(m[532]&m[533]&~m[534]&~m[536]&m[537])|(m[532]&~m[533]&m[534]&~m[536]&m[537])|(~m[532]&~m[533]&~m[534]&m[536]&m[537])|(m[532]&~m[533]&~m[534]&m[536]&m[537])|(~m[532]&m[533]&~m[534]&m[536]&m[537])|(m[532]&m[533]&~m[534]&m[536]&m[537])|(~m[532]&~m[533]&m[534]&m[536]&m[537])|(m[532]&~m[533]&m[534]&m[536]&m[537])|(m[532]&m[533]&m[534]&m[536]&m[537]))):InitCond[514];
    m[545] = run?((((m[537]&~m[543]&~m[544]&~m[546]&~m[547])|(~m[537]&~m[543]&~m[544]&m[546]&~m[547])|(m[537]&m[543]&~m[544]&m[546]&~m[547])|(m[537]&~m[543]&m[544]&m[546]&~m[547])|(~m[537]&m[543]&~m[544]&~m[546]&m[547])|(~m[537]&~m[543]&m[544]&~m[546]&m[547])|(m[537]&m[543]&m[544]&~m[546]&m[547])|(~m[537]&m[543]&m[544]&m[546]&m[547]))&UnbiasedRNG[132])|((m[537]&~m[543]&~m[544]&m[546]&~m[547])|(~m[537]&~m[543]&~m[544]&~m[546]&m[547])|(m[537]&~m[543]&~m[544]&~m[546]&m[547])|(m[537]&m[543]&~m[544]&~m[546]&m[547])|(m[537]&~m[543]&m[544]&~m[546]&m[547])|(~m[537]&~m[543]&~m[544]&m[546]&m[547])|(m[537]&~m[543]&~m[544]&m[546]&m[547])|(~m[537]&m[543]&~m[544]&m[546]&m[547])|(m[537]&m[543]&~m[544]&m[546]&m[547])|(~m[537]&~m[543]&m[544]&m[546]&m[547])|(m[537]&~m[543]&m[544]&m[546]&m[547])|(m[537]&m[543]&m[544]&m[546]&m[547]))):InitCond[515];
    m[550] = run?((((m[542]&~m[548]&~m[549]&~m[551]&~m[552])|(~m[542]&~m[548]&~m[549]&m[551]&~m[552])|(m[542]&m[548]&~m[549]&m[551]&~m[552])|(m[542]&~m[548]&m[549]&m[551]&~m[552])|(~m[542]&m[548]&~m[549]&~m[551]&m[552])|(~m[542]&~m[548]&m[549]&~m[551]&m[552])|(m[542]&m[548]&m[549]&~m[551]&m[552])|(~m[542]&m[548]&m[549]&m[551]&m[552]))&UnbiasedRNG[133])|((m[542]&~m[548]&~m[549]&m[551]&~m[552])|(~m[542]&~m[548]&~m[549]&~m[551]&m[552])|(m[542]&~m[548]&~m[549]&~m[551]&m[552])|(m[542]&m[548]&~m[549]&~m[551]&m[552])|(m[542]&~m[548]&m[549]&~m[551]&m[552])|(~m[542]&~m[548]&~m[549]&m[551]&m[552])|(m[542]&~m[548]&~m[549]&m[551]&m[552])|(~m[542]&m[548]&~m[549]&m[551]&m[552])|(m[542]&m[548]&~m[549]&m[551]&m[552])|(~m[542]&~m[548]&m[549]&m[551]&m[552])|(m[542]&~m[548]&m[549]&m[551]&m[552])|(m[542]&m[548]&m[549]&m[551]&m[552]))):InitCond[516];
    m[560] = run?((((m[547]&~m[558]&~m[559]&~m[561]&~m[562])|(~m[547]&~m[558]&~m[559]&m[561]&~m[562])|(m[547]&m[558]&~m[559]&m[561]&~m[562])|(m[547]&~m[558]&m[559]&m[561]&~m[562])|(~m[547]&m[558]&~m[559]&~m[561]&m[562])|(~m[547]&~m[558]&m[559]&~m[561]&m[562])|(m[547]&m[558]&m[559]&~m[561]&m[562])|(~m[547]&m[558]&m[559]&m[561]&m[562]))&UnbiasedRNG[134])|((m[547]&~m[558]&~m[559]&m[561]&~m[562])|(~m[547]&~m[558]&~m[559]&~m[561]&m[562])|(m[547]&~m[558]&~m[559]&~m[561]&m[562])|(m[547]&m[558]&~m[559]&~m[561]&m[562])|(m[547]&~m[558]&m[559]&~m[561]&m[562])|(~m[547]&~m[558]&~m[559]&m[561]&m[562])|(m[547]&~m[558]&~m[559]&m[561]&m[562])|(~m[547]&m[558]&~m[559]&m[561]&m[562])|(m[547]&m[558]&~m[559]&m[561]&m[562])|(~m[547]&~m[558]&m[559]&m[561]&m[562])|(m[547]&~m[558]&m[559]&m[561]&m[562])|(m[547]&m[558]&m[559]&m[561]&m[562]))):InitCond[517];
    m[565] = run?((((m[552]&~m[563]&~m[564]&~m[566]&~m[567])|(~m[552]&~m[563]&~m[564]&m[566]&~m[567])|(m[552]&m[563]&~m[564]&m[566]&~m[567])|(m[552]&~m[563]&m[564]&m[566]&~m[567])|(~m[552]&m[563]&~m[564]&~m[566]&m[567])|(~m[552]&~m[563]&m[564]&~m[566]&m[567])|(m[552]&m[563]&m[564]&~m[566]&m[567])|(~m[552]&m[563]&m[564]&m[566]&m[567]))&UnbiasedRNG[135])|((m[552]&~m[563]&~m[564]&m[566]&~m[567])|(~m[552]&~m[563]&~m[564]&~m[566]&m[567])|(m[552]&~m[563]&~m[564]&~m[566]&m[567])|(m[552]&m[563]&~m[564]&~m[566]&m[567])|(m[552]&~m[563]&m[564]&~m[566]&m[567])|(~m[552]&~m[563]&~m[564]&m[566]&m[567])|(m[552]&~m[563]&~m[564]&m[566]&m[567])|(~m[552]&m[563]&~m[564]&m[566]&m[567])|(m[552]&m[563]&~m[564]&m[566]&m[567])|(~m[552]&~m[563]&m[564]&m[566]&m[567])|(m[552]&~m[563]&m[564]&m[566]&m[567])|(m[552]&m[563]&m[564]&m[566]&m[567]))):InitCond[518];
    m[570] = run?((((m[557]&~m[568]&~m[569]&~m[571]&~m[572])|(~m[557]&~m[568]&~m[569]&m[571]&~m[572])|(m[557]&m[568]&~m[569]&m[571]&~m[572])|(m[557]&~m[568]&m[569]&m[571]&~m[572])|(~m[557]&m[568]&~m[569]&~m[571]&m[572])|(~m[557]&~m[568]&m[569]&~m[571]&m[572])|(m[557]&m[568]&m[569]&~m[571]&m[572])|(~m[557]&m[568]&m[569]&m[571]&m[572]))&UnbiasedRNG[136])|((m[557]&~m[568]&~m[569]&m[571]&~m[572])|(~m[557]&~m[568]&~m[569]&~m[571]&m[572])|(m[557]&~m[568]&~m[569]&~m[571]&m[572])|(m[557]&m[568]&~m[569]&~m[571]&m[572])|(m[557]&~m[568]&m[569]&~m[571]&m[572])|(~m[557]&~m[568]&~m[569]&m[571]&m[572])|(m[557]&~m[568]&~m[569]&m[571]&m[572])|(~m[557]&m[568]&~m[569]&m[571]&m[572])|(m[557]&m[568]&~m[569]&m[571]&m[572])|(~m[557]&~m[568]&m[569]&m[571]&m[572])|(m[557]&~m[568]&m[569]&m[571]&m[572])|(m[557]&m[568]&m[569]&m[571]&m[572]))):InitCond[519];
    m[580] = run?((((m[562]&~m[578]&~m[579]&~m[581]&~m[582])|(~m[562]&~m[578]&~m[579]&m[581]&~m[582])|(m[562]&m[578]&~m[579]&m[581]&~m[582])|(m[562]&~m[578]&m[579]&m[581]&~m[582])|(~m[562]&m[578]&~m[579]&~m[581]&m[582])|(~m[562]&~m[578]&m[579]&~m[581]&m[582])|(m[562]&m[578]&m[579]&~m[581]&m[582])|(~m[562]&m[578]&m[579]&m[581]&m[582]))&UnbiasedRNG[137])|((m[562]&~m[578]&~m[579]&m[581]&~m[582])|(~m[562]&~m[578]&~m[579]&~m[581]&m[582])|(m[562]&~m[578]&~m[579]&~m[581]&m[582])|(m[562]&m[578]&~m[579]&~m[581]&m[582])|(m[562]&~m[578]&m[579]&~m[581]&m[582])|(~m[562]&~m[578]&~m[579]&m[581]&m[582])|(m[562]&~m[578]&~m[579]&m[581]&m[582])|(~m[562]&m[578]&~m[579]&m[581]&m[582])|(m[562]&m[578]&~m[579]&m[581]&m[582])|(~m[562]&~m[578]&m[579]&m[581]&m[582])|(m[562]&~m[578]&m[579]&m[581]&m[582])|(m[562]&m[578]&m[579]&m[581]&m[582]))):InitCond[520];
    m[585] = run?((((m[567]&~m[583]&~m[584]&~m[586]&~m[587])|(~m[567]&~m[583]&~m[584]&m[586]&~m[587])|(m[567]&m[583]&~m[584]&m[586]&~m[587])|(m[567]&~m[583]&m[584]&m[586]&~m[587])|(~m[567]&m[583]&~m[584]&~m[586]&m[587])|(~m[567]&~m[583]&m[584]&~m[586]&m[587])|(m[567]&m[583]&m[584]&~m[586]&m[587])|(~m[567]&m[583]&m[584]&m[586]&m[587]))&UnbiasedRNG[138])|((m[567]&~m[583]&~m[584]&m[586]&~m[587])|(~m[567]&~m[583]&~m[584]&~m[586]&m[587])|(m[567]&~m[583]&~m[584]&~m[586]&m[587])|(m[567]&m[583]&~m[584]&~m[586]&m[587])|(m[567]&~m[583]&m[584]&~m[586]&m[587])|(~m[567]&~m[583]&~m[584]&m[586]&m[587])|(m[567]&~m[583]&~m[584]&m[586]&m[587])|(~m[567]&m[583]&~m[584]&m[586]&m[587])|(m[567]&m[583]&~m[584]&m[586]&m[587])|(~m[567]&~m[583]&m[584]&m[586]&m[587])|(m[567]&~m[583]&m[584]&m[586]&m[587])|(m[567]&m[583]&m[584]&m[586]&m[587]))):InitCond[521];
    m[590] = run?((((m[572]&~m[588]&~m[589]&~m[591]&~m[592])|(~m[572]&~m[588]&~m[589]&m[591]&~m[592])|(m[572]&m[588]&~m[589]&m[591]&~m[592])|(m[572]&~m[588]&m[589]&m[591]&~m[592])|(~m[572]&m[588]&~m[589]&~m[591]&m[592])|(~m[572]&~m[588]&m[589]&~m[591]&m[592])|(m[572]&m[588]&m[589]&~m[591]&m[592])|(~m[572]&m[588]&m[589]&m[591]&m[592]))&UnbiasedRNG[139])|((m[572]&~m[588]&~m[589]&m[591]&~m[592])|(~m[572]&~m[588]&~m[589]&~m[591]&m[592])|(m[572]&~m[588]&~m[589]&~m[591]&m[592])|(m[572]&m[588]&~m[589]&~m[591]&m[592])|(m[572]&~m[588]&m[589]&~m[591]&m[592])|(~m[572]&~m[588]&~m[589]&m[591]&m[592])|(m[572]&~m[588]&~m[589]&m[591]&m[592])|(~m[572]&m[588]&~m[589]&m[591]&m[592])|(m[572]&m[588]&~m[589]&m[591]&m[592])|(~m[572]&~m[588]&m[589]&m[591]&m[592])|(m[572]&~m[588]&m[589]&m[591]&m[592])|(m[572]&m[588]&m[589]&m[591]&m[592]))):InitCond[522];
    m[595] = run?((((m[577]&~m[593]&~m[594]&~m[596]&~m[597])|(~m[577]&~m[593]&~m[594]&m[596]&~m[597])|(m[577]&m[593]&~m[594]&m[596]&~m[597])|(m[577]&~m[593]&m[594]&m[596]&~m[597])|(~m[577]&m[593]&~m[594]&~m[596]&m[597])|(~m[577]&~m[593]&m[594]&~m[596]&m[597])|(m[577]&m[593]&m[594]&~m[596]&m[597])|(~m[577]&m[593]&m[594]&m[596]&m[597]))&UnbiasedRNG[140])|((m[577]&~m[593]&~m[594]&m[596]&~m[597])|(~m[577]&~m[593]&~m[594]&~m[596]&m[597])|(m[577]&~m[593]&~m[594]&~m[596]&m[597])|(m[577]&m[593]&~m[594]&~m[596]&m[597])|(m[577]&~m[593]&m[594]&~m[596]&m[597])|(~m[577]&~m[593]&~m[594]&m[596]&m[597])|(m[577]&~m[593]&~m[594]&m[596]&m[597])|(~m[577]&m[593]&~m[594]&m[596]&m[597])|(m[577]&m[593]&~m[594]&m[596]&m[597])|(~m[577]&~m[593]&m[594]&m[596]&m[597])|(m[577]&~m[593]&m[594]&m[596]&m[597])|(m[577]&m[593]&m[594]&m[596]&m[597]))):InitCond[523];
    m[605] = run?((((m[582]&~m[603]&~m[604]&~m[606]&~m[607])|(~m[582]&~m[603]&~m[604]&m[606]&~m[607])|(m[582]&m[603]&~m[604]&m[606]&~m[607])|(m[582]&~m[603]&m[604]&m[606]&~m[607])|(~m[582]&m[603]&~m[604]&~m[606]&m[607])|(~m[582]&~m[603]&m[604]&~m[606]&m[607])|(m[582]&m[603]&m[604]&~m[606]&m[607])|(~m[582]&m[603]&m[604]&m[606]&m[607]))&UnbiasedRNG[141])|((m[582]&~m[603]&~m[604]&m[606]&~m[607])|(~m[582]&~m[603]&~m[604]&~m[606]&m[607])|(m[582]&~m[603]&~m[604]&~m[606]&m[607])|(m[582]&m[603]&~m[604]&~m[606]&m[607])|(m[582]&~m[603]&m[604]&~m[606]&m[607])|(~m[582]&~m[603]&~m[604]&m[606]&m[607])|(m[582]&~m[603]&~m[604]&m[606]&m[607])|(~m[582]&m[603]&~m[604]&m[606]&m[607])|(m[582]&m[603]&~m[604]&m[606]&m[607])|(~m[582]&~m[603]&m[604]&m[606]&m[607])|(m[582]&~m[603]&m[604]&m[606]&m[607])|(m[582]&m[603]&m[604]&m[606]&m[607]))):InitCond[524];
    m[610] = run?((((m[587]&~m[608]&~m[609]&~m[611]&~m[612])|(~m[587]&~m[608]&~m[609]&m[611]&~m[612])|(m[587]&m[608]&~m[609]&m[611]&~m[612])|(m[587]&~m[608]&m[609]&m[611]&~m[612])|(~m[587]&m[608]&~m[609]&~m[611]&m[612])|(~m[587]&~m[608]&m[609]&~m[611]&m[612])|(m[587]&m[608]&m[609]&~m[611]&m[612])|(~m[587]&m[608]&m[609]&m[611]&m[612]))&UnbiasedRNG[142])|((m[587]&~m[608]&~m[609]&m[611]&~m[612])|(~m[587]&~m[608]&~m[609]&~m[611]&m[612])|(m[587]&~m[608]&~m[609]&~m[611]&m[612])|(m[587]&m[608]&~m[609]&~m[611]&m[612])|(m[587]&~m[608]&m[609]&~m[611]&m[612])|(~m[587]&~m[608]&~m[609]&m[611]&m[612])|(m[587]&~m[608]&~m[609]&m[611]&m[612])|(~m[587]&m[608]&~m[609]&m[611]&m[612])|(m[587]&m[608]&~m[609]&m[611]&m[612])|(~m[587]&~m[608]&m[609]&m[611]&m[612])|(m[587]&~m[608]&m[609]&m[611]&m[612])|(m[587]&m[608]&m[609]&m[611]&m[612]))):InitCond[525];
    m[615] = run?((((m[592]&~m[613]&~m[614]&~m[616]&~m[617])|(~m[592]&~m[613]&~m[614]&m[616]&~m[617])|(m[592]&m[613]&~m[614]&m[616]&~m[617])|(m[592]&~m[613]&m[614]&m[616]&~m[617])|(~m[592]&m[613]&~m[614]&~m[616]&m[617])|(~m[592]&~m[613]&m[614]&~m[616]&m[617])|(m[592]&m[613]&m[614]&~m[616]&m[617])|(~m[592]&m[613]&m[614]&m[616]&m[617]))&UnbiasedRNG[143])|((m[592]&~m[613]&~m[614]&m[616]&~m[617])|(~m[592]&~m[613]&~m[614]&~m[616]&m[617])|(m[592]&~m[613]&~m[614]&~m[616]&m[617])|(m[592]&m[613]&~m[614]&~m[616]&m[617])|(m[592]&~m[613]&m[614]&~m[616]&m[617])|(~m[592]&~m[613]&~m[614]&m[616]&m[617])|(m[592]&~m[613]&~m[614]&m[616]&m[617])|(~m[592]&m[613]&~m[614]&m[616]&m[617])|(m[592]&m[613]&~m[614]&m[616]&m[617])|(~m[592]&~m[613]&m[614]&m[616]&m[617])|(m[592]&~m[613]&m[614]&m[616]&m[617])|(m[592]&m[613]&m[614]&m[616]&m[617]))):InitCond[526];
    m[620] = run?((((m[597]&~m[618]&~m[619]&~m[621]&~m[622])|(~m[597]&~m[618]&~m[619]&m[621]&~m[622])|(m[597]&m[618]&~m[619]&m[621]&~m[622])|(m[597]&~m[618]&m[619]&m[621]&~m[622])|(~m[597]&m[618]&~m[619]&~m[621]&m[622])|(~m[597]&~m[618]&m[619]&~m[621]&m[622])|(m[597]&m[618]&m[619]&~m[621]&m[622])|(~m[597]&m[618]&m[619]&m[621]&m[622]))&UnbiasedRNG[144])|((m[597]&~m[618]&~m[619]&m[621]&~m[622])|(~m[597]&~m[618]&~m[619]&~m[621]&m[622])|(m[597]&~m[618]&~m[619]&~m[621]&m[622])|(m[597]&m[618]&~m[619]&~m[621]&m[622])|(m[597]&~m[618]&m[619]&~m[621]&m[622])|(~m[597]&~m[618]&~m[619]&m[621]&m[622])|(m[597]&~m[618]&~m[619]&m[621]&m[622])|(~m[597]&m[618]&~m[619]&m[621]&m[622])|(m[597]&m[618]&~m[619]&m[621]&m[622])|(~m[597]&~m[618]&m[619]&m[621]&m[622])|(m[597]&~m[618]&m[619]&m[621]&m[622])|(m[597]&m[618]&m[619]&m[621]&m[622]))):InitCond[527];
    m[625] = run?((((m[602]&~m[623]&~m[624]&~m[626]&~m[627])|(~m[602]&~m[623]&~m[624]&m[626]&~m[627])|(m[602]&m[623]&~m[624]&m[626]&~m[627])|(m[602]&~m[623]&m[624]&m[626]&~m[627])|(~m[602]&m[623]&~m[624]&~m[626]&m[627])|(~m[602]&~m[623]&m[624]&~m[626]&m[627])|(m[602]&m[623]&m[624]&~m[626]&m[627])|(~m[602]&m[623]&m[624]&m[626]&m[627]))&UnbiasedRNG[145])|((m[602]&~m[623]&~m[624]&m[626]&~m[627])|(~m[602]&~m[623]&~m[624]&~m[626]&m[627])|(m[602]&~m[623]&~m[624]&~m[626]&m[627])|(m[602]&m[623]&~m[624]&~m[626]&m[627])|(m[602]&~m[623]&m[624]&~m[626]&m[627])|(~m[602]&~m[623]&~m[624]&m[626]&m[627])|(m[602]&~m[623]&~m[624]&m[626]&m[627])|(~m[602]&m[623]&~m[624]&m[626]&m[627])|(m[602]&m[623]&~m[624]&m[626]&m[627])|(~m[602]&~m[623]&m[624]&m[626]&m[627])|(m[602]&~m[623]&m[624]&m[626]&m[627])|(m[602]&m[623]&m[624]&m[626]&m[627]))):InitCond[528];
    m[635] = run?((((m[607]&~m[633]&~m[634]&~m[636]&~m[637])|(~m[607]&~m[633]&~m[634]&m[636]&~m[637])|(m[607]&m[633]&~m[634]&m[636]&~m[637])|(m[607]&~m[633]&m[634]&m[636]&~m[637])|(~m[607]&m[633]&~m[634]&~m[636]&m[637])|(~m[607]&~m[633]&m[634]&~m[636]&m[637])|(m[607]&m[633]&m[634]&~m[636]&m[637])|(~m[607]&m[633]&m[634]&m[636]&m[637]))&UnbiasedRNG[146])|((m[607]&~m[633]&~m[634]&m[636]&~m[637])|(~m[607]&~m[633]&~m[634]&~m[636]&m[637])|(m[607]&~m[633]&~m[634]&~m[636]&m[637])|(m[607]&m[633]&~m[634]&~m[636]&m[637])|(m[607]&~m[633]&m[634]&~m[636]&m[637])|(~m[607]&~m[633]&~m[634]&m[636]&m[637])|(m[607]&~m[633]&~m[634]&m[636]&m[637])|(~m[607]&m[633]&~m[634]&m[636]&m[637])|(m[607]&m[633]&~m[634]&m[636]&m[637])|(~m[607]&~m[633]&m[634]&m[636]&m[637])|(m[607]&~m[633]&m[634]&m[636]&m[637])|(m[607]&m[633]&m[634]&m[636]&m[637]))):InitCond[529];
    m[640] = run?((((m[612]&~m[638]&~m[639]&~m[641]&~m[642])|(~m[612]&~m[638]&~m[639]&m[641]&~m[642])|(m[612]&m[638]&~m[639]&m[641]&~m[642])|(m[612]&~m[638]&m[639]&m[641]&~m[642])|(~m[612]&m[638]&~m[639]&~m[641]&m[642])|(~m[612]&~m[638]&m[639]&~m[641]&m[642])|(m[612]&m[638]&m[639]&~m[641]&m[642])|(~m[612]&m[638]&m[639]&m[641]&m[642]))&UnbiasedRNG[147])|((m[612]&~m[638]&~m[639]&m[641]&~m[642])|(~m[612]&~m[638]&~m[639]&~m[641]&m[642])|(m[612]&~m[638]&~m[639]&~m[641]&m[642])|(m[612]&m[638]&~m[639]&~m[641]&m[642])|(m[612]&~m[638]&m[639]&~m[641]&m[642])|(~m[612]&~m[638]&~m[639]&m[641]&m[642])|(m[612]&~m[638]&~m[639]&m[641]&m[642])|(~m[612]&m[638]&~m[639]&m[641]&m[642])|(m[612]&m[638]&~m[639]&m[641]&m[642])|(~m[612]&~m[638]&m[639]&m[641]&m[642])|(m[612]&~m[638]&m[639]&m[641]&m[642])|(m[612]&m[638]&m[639]&m[641]&m[642]))):InitCond[530];
    m[645] = run?((((m[617]&~m[643]&~m[644]&~m[646]&~m[647])|(~m[617]&~m[643]&~m[644]&m[646]&~m[647])|(m[617]&m[643]&~m[644]&m[646]&~m[647])|(m[617]&~m[643]&m[644]&m[646]&~m[647])|(~m[617]&m[643]&~m[644]&~m[646]&m[647])|(~m[617]&~m[643]&m[644]&~m[646]&m[647])|(m[617]&m[643]&m[644]&~m[646]&m[647])|(~m[617]&m[643]&m[644]&m[646]&m[647]))&UnbiasedRNG[148])|((m[617]&~m[643]&~m[644]&m[646]&~m[647])|(~m[617]&~m[643]&~m[644]&~m[646]&m[647])|(m[617]&~m[643]&~m[644]&~m[646]&m[647])|(m[617]&m[643]&~m[644]&~m[646]&m[647])|(m[617]&~m[643]&m[644]&~m[646]&m[647])|(~m[617]&~m[643]&~m[644]&m[646]&m[647])|(m[617]&~m[643]&~m[644]&m[646]&m[647])|(~m[617]&m[643]&~m[644]&m[646]&m[647])|(m[617]&m[643]&~m[644]&m[646]&m[647])|(~m[617]&~m[643]&m[644]&m[646]&m[647])|(m[617]&~m[643]&m[644]&m[646]&m[647])|(m[617]&m[643]&m[644]&m[646]&m[647]))):InitCond[531];
    m[650] = run?((((m[622]&~m[648]&~m[649]&~m[651]&~m[652])|(~m[622]&~m[648]&~m[649]&m[651]&~m[652])|(m[622]&m[648]&~m[649]&m[651]&~m[652])|(m[622]&~m[648]&m[649]&m[651]&~m[652])|(~m[622]&m[648]&~m[649]&~m[651]&m[652])|(~m[622]&~m[648]&m[649]&~m[651]&m[652])|(m[622]&m[648]&m[649]&~m[651]&m[652])|(~m[622]&m[648]&m[649]&m[651]&m[652]))&UnbiasedRNG[149])|((m[622]&~m[648]&~m[649]&m[651]&~m[652])|(~m[622]&~m[648]&~m[649]&~m[651]&m[652])|(m[622]&~m[648]&~m[649]&~m[651]&m[652])|(m[622]&m[648]&~m[649]&~m[651]&m[652])|(m[622]&~m[648]&m[649]&~m[651]&m[652])|(~m[622]&~m[648]&~m[649]&m[651]&m[652])|(m[622]&~m[648]&~m[649]&m[651]&m[652])|(~m[622]&m[648]&~m[649]&m[651]&m[652])|(m[622]&m[648]&~m[649]&m[651]&m[652])|(~m[622]&~m[648]&m[649]&m[651]&m[652])|(m[622]&~m[648]&m[649]&m[651]&m[652])|(m[622]&m[648]&m[649]&m[651]&m[652]))):InitCond[532];
    m[655] = run?((((m[627]&~m[653]&~m[654]&~m[656]&~m[657])|(~m[627]&~m[653]&~m[654]&m[656]&~m[657])|(m[627]&m[653]&~m[654]&m[656]&~m[657])|(m[627]&~m[653]&m[654]&m[656]&~m[657])|(~m[627]&m[653]&~m[654]&~m[656]&m[657])|(~m[627]&~m[653]&m[654]&~m[656]&m[657])|(m[627]&m[653]&m[654]&~m[656]&m[657])|(~m[627]&m[653]&m[654]&m[656]&m[657]))&UnbiasedRNG[150])|((m[627]&~m[653]&~m[654]&m[656]&~m[657])|(~m[627]&~m[653]&~m[654]&~m[656]&m[657])|(m[627]&~m[653]&~m[654]&~m[656]&m[657])|(m[627]&m[653]&~m[654]&~m[656]&m[657])|(m[627]&~m[653]&m[654]&~m[656]&m[657])|(~m[627]&~m[653]&~m[654]&m[656]&m[657])|(m[627]&~m[653]&~m[654]&m[656]&m[657])|(~m[627]&m[653]&~m[654]&m[656]&m[657])|(m[627]&m[653]&~m[654]&m[656]&m[657])|(~m[627]&~m[653]&m[654]&m[656]&m[657])|(m[627]&~m[653]&m[654]&m[656]&m[657])|(m[627]&m[653]&m[654]&m[656]&m[657]))):InitCond[533];
    m[660] = run?((((m[632]&~m[658]&~m[659]&~m[661]&~m[662])|(~m[632]&~m[658]&~m[659]&m[661]&~m[662])|(m[632]&m[658]&~m[659]&m[661]&~m[662])|(m[632]&~m[658]&m[659]&m[661]&~m[662])|(~m[632]&m[658]&~m[659]&~m[661]&m[662])|(~m[632]&~m[658]&m[659]&~m[661]&m[662])|(m[632]&m[658]&m[659]&~m[661]&m[662])|(~m[632]&m[658]&m[659]&m[661]&m[662]))&UnbiasedRNG[151])|((m[632]&~m[658]&~m[659]&m[661]&~m[662])|(~m[632]&~m[658]&~m[659]&~m[661]&m[662])|(m[632]&~m[658]&~m[659]&~m[661]&m[662])|(m[632]&m[658]&~m[659]&~m[661]&m[662])|(m[632]&~m[658]&m[659]&~m[661]&m[662])|(~m[632]&~m[658]&~m[659]&m[661]&m[662])|(m[632]&~m[658]&~m[659]&m[661]&m[662])|(~m[632]&m[658]&~m[659]&m[661]&m[662])|(m[632]&m[658]&~m[659]&m[661]&m[662])|(~m[632]&~m[658]&m[659]&m[661]&m[662])|(m[632]&~m[658]&m[659]&m[661]&m[662])|(m[632]&m[658]&m[659]&m[661]&m[662]))):InitCond[534];
    m[670] = run?((((m[637]&~m[668]&~m[669]&~m[671]&~m[672])|(~m[637]&~m[668]&~m[669]&m[671]&~m[672])|(m[637]&m[668]&~m[669]&m[671]&~m[672])|(m[637]&~m[668]&m[669]&m[671]&~m[672])|(~m[637]&m[668]&~m[669]&~m[671]&m[672])|(~m[637]&~m[668]&m[669]&~m[671]&m[672])|(m[637]&m[668]&m[669]&~m[671]&m[672])|(~m[637]&m[668]&m[669]&m[671]&m[672]))&UnbiasedRNG[152])|((m[637]&~m[668]&~m[669]&m[671]&~m[672])|(~m[637]&~m[668]&~m[669]&~m[671]&m[672])|(m[637]&~m[668]&~m[669]&~m[671]&m[672])|(m[637]&m[668]&~m[669]&~m[671]&m[672])|(m[637]&~m[668]&m[669]&~m[671]&m[672])|(~m[637]&~m[668]&~m[669]&m[671]&m[672])|(m[637]&~m[668]&~m[669]&m[671]&m[672])|(~m[637]&m[668]&~m[669]&m[671]&m[672])|(m[637]&m[668]&~m[669]&m[671]&m[672])|(~m[637]&~m[668]&m[669]&m[671]&m[672])|(m[637]&~m[668]&m[669]&m[671]&m[672])|(m[637]&m[668]&m[669]&m[671]&m[672]))):InitCond[535];
    m[675] = run?((((m[642]&~m[673]&~m[674]&~m[676]&~m[677])|(~m[642]&~m[673]&~m[674]&m[676]&~m[677])|(m[642]&m[673]&~m[674]&m[676]&~m[677])|(m[642]&~m[673]&m[674]&m[676]&~m[677])|(~m[642]&m[673]&~m[674]&~m[676]&m[677])|(~m[642]&~m[673]&m[674]&~m[676]&m[677])|(m[642]&m[673]&m[674]&~m[676]&m[677])|(~m[642]&m[673]&m[674]&m[676]&m[677]))&UnbiasedRNG[153])|((m[642]&~m[673]&~m[674]&m[676]&~m[677])|(~m[642]&~m[673]&~m[674]&~m[676]&m[677])|(m[642]&~m[673]&~m[674]&~m[676]&m[677])|(m[642]&m[673]&~m[674]&~m[676]&m[677])|(m[642]&~m[673]&m[674]&~m[676]&m[677])|(~m[642]&~m[673]&~m[674]&m[676]&m[677])|(m[642]&~m[673]&~m[674]&m[676]&m[677])|(~m[642]&m[673]&~m[674]&m[676]&m[677])|(m[642]&m[673]&~m[674]&m[676]&m[677])|(~m[642]&~m[673]&m[674]&m[676]&m[677])|(m[642]&~m[673]&m[674]&m[676]&m[677])|(m[642]&m[673]&m[674]&m[676]&m[677]))):InitCond[536];
    m[680] = run?((((m[647]&~m[678]&~m[679]&~m[681]&~m[682])|(~m[647]&~m[678]&~m[679]&m[681]&~m[682])|(m[647]&m[678]&~m[679]&m[681]&~m[682])|(m[647]&~m[678]&m[679]&m[681]&~m[682])|(~m[647]&m[678]&~m[679]&~m[681]&m[682])|(~m[647]&~m[678]&m[679]&~m[681]&m[682])|(m[647]&m[678]&m[679]&~m[681]&m[682])|(~m[647]&m[678]&m[679]&m[681]&m[682]))&UnbiasedRNG[154])|((m[647]&~m[678]&~m[679]&m[681]&~m[682])|(~m[647]&~m[678]&~m[679]&~m[681]&m[682])|(m[647]&~m[678]&~m[679]&~m[681]&m[682])|(m[647]&m[678]&~m[679]&~m[681]&m[682])|(m[647]&~m[678]&m[679]&~m[681]&m[682])|(~m[647]&~m[678]&~m[679]&m[681]&m[682])|(m[647]&~m[678]&~m[679]&m[681]&m[682])|(~m[647]&m[678]&~m[679]&m[681]&m[682])|(m[647]&m[678]&~m[679]&m[681]&m[682])|(~m[647]&~m[678]&m[679]&m[681]&m[682])|(m[647]&~m[678]&m[679]&m[681]&m[682])|(m[647]&m[678]&m[679]&m[681]&m[682]))):InitCond[537];
    m[685] = run?((((m[652]&~m[683]&~m[684]&~m[686]&~m[687])|(~m[652]&~m[683]&~m[684]&m[686]&~m[687])|(m[652]&m[683]&~m[684]&m[686]&~m[687])|(m[652]&~m[683]&m[684]&m[686]&~m[687])|(~m[652]&m[683]&~m[684]&~m[686]&m[687])|(~m[652]&~m[683]&m[684]&~m[686]&m[687])|(m[652]&m[683]&m[684]&~m[686]&m[687])|(~m[652]&m[683]&m[684]&m[686]&m[687]))&UnbiasedRNG[155])|((m[652]&~m[683]&~m[684]&m[686]&~m[687])|(~m[652]&~m[683]&~m[684]&~m[686]&m[687])|(m[652]&~m[683]&~m[684]&~m[686]&m[687])|(m[652]&m[683]&~m[684]&~m[686]&m[687])|(m[652]&~m[683]&m[684]&~m[686]&m[687])|(~m[652]&~m[683]&~m[684]&m[686]&m[687])|(m[652]&~m[683]&~m[684]&m[686]&m[687])|(~m[652]&m[683]&~m[684]&m[686]&m[687])|(m[652]&m[683]&~m[684]&m[686]&m[687])|(~m[652]&~m[683]&m[684]&m[686]&m[687])|(m[652]&~m[683]&m[684]&m[686]&m[687])|(m[652]&m[683]&m[684]&m[686]&m[687]))):InitCond[538];
    m[690] = run?((((m[657]&~m[688]&~m[689]&~m[691]&~m[692])|(~m[657]&~m[688]&~m[689]&m[691]&~m[692])|(m[657]&m[688]&~m[689]&m[691]&~m[692])|(m[657]&~m[688]&m[689]&m[691]&~m[692])|(~m[657]&m[688]&~m[689]&~m[691]&m[692])|(~m[657]&~m[688]&m[689]&~m[691]&m[692])|(m[657]&m[688]&m[689]&~m[691]&m[692])|(~m[657]&m[688]&m[689]&m[691]&m[692]))&UnbiasedRNG[156])|((m[657]&~m[688]&~m[689]&m[691]&~m[692])|(~m[657]&~m[688]&~m[689]&~m[691]&m[692])|(m[657]&~m[688]&~m[689]&~m[691]&m[692])|(m[657]&m[688]&~m[689]&~m[691]&m[692])|(m[657]&~m[688]&m[689]&~m[691]&m[692])|(~m[657]&~m[688]&~m[689]&m[691]&m[692])|(m[657]&~m[688]&~m[689]&m[691]&m[692])|(~m[657]&m[688]&~m[689]&m[691]&m[692])|(m[657]&m[688]&~m[689]&m[691]&m[692])|(~m[657]&~m[688]&m[689]&m[691]&m[692])|(m[657]&~m[688]&m[689]&m[691]&m[692])|(m[657]&m[688]&m[689]&m[691]&m[692]))):InitCond[539];
    m[695] = run?((((m[662]&~m[693]&~m[694]&~m[696]&~m[697])|(~m[662]&~m[693]&~m[694]&m[696]&~m[697])|(m[662]&m[693]&~m[694]&m[696]&~m[697])|(m[662]&~m[693]&m[694]&m[696]&~m[697])|(~m[662]&m[693]&~m[694]&~m[696]&m[697])|(~m[662]&~m[693]&m[694]&~m[696]&m[697])|(m[662]&m[693]&m[694]&~m[696]&m[697])|(~m[662]&m[693]&m[694]&m[696]&m[697]))&UnbiasedRNG[157])|((m[662]&~m[693]&~m[694]&m[696]&~m[697])|(~m[662]&~m[693]&~m[694]&~m[696]&m[697])|(m[662]&~m[693]&~m[694]&~m[696]&m[697])|(m[662]&m[693]&~m[694]&~m[696]&m[697])|(m[662]&~m[693]&m[694]&~m[696]&m[697])|(~m[662]&~m[693]&~m[694]&m[696]&m[697])|(m[662]&~m[693]&~m[694]&m[696]&m[697])|(~m[662]&m[693]&~m[694]&m[696]&m[697])|(m[662]&m[693]&~m[694]&m[696]&m[697])|(~m[662]&~m[693]&m[694]&m[696]&m[697])|(m[662]&~m[693]&m[694]&m[696]&m[697])|(m[662]&m[693]&m[694]&m[696]&m[697]))):InitCond[540];
    m[700] = run?((((m[667]&~m[698]&~m[699]&~m[701]&~m[702])|(~m[667]&~m[698]&~m[699]&m[701]&~m[702])|(m[667]&m[698]&~m[699]&m[701]&~m[702])|(m[667]&~m[698]&m[699]&m[701]&~m[702])|(~m[667]&m[698]&~m[699]&~m[701]&m[702])|(~m[667]&~m[698]&m[699]&~m[701]&m[702])|(m[667]&m[698]&m[699]&~m[701]&m[702])|(~m[667]&m[698]&m[699]&m[701]&m[702]))&UnbiasedRNG[158])|((m[667]&~m[698]&~m[699]&m[701]&~m[702])|(~m[667]&~m[698]&~m[699]&~m[701]&m[702])|(m[667]&~m[698]&~m[699]&~m[701]&m[702])|(m[667]&m[698]&~m[699]&~m[701]&m[702])|(m[667]&~m[698]&m[699]&~m[701]&m[702])|(~m[667]&~m[698]&~m[699]&m[701]&m[702])|(m[667]&~m[698]&~m[699]&m[701]&m[702])|(~m[667]&m[698]&~m[699]&m[701]&m[702])|(m[667]&m[698]&~m[699]&m[701]&m[702])|(~m[667]&~m[698]&m[699]&m[701]&m[702])|(m[667]&~m[698]&m[699]&m[701]&m[702])|(m[667]&m[698]&m[699]&m[701]&m[702]))):InitCond[541];
    m[710] = run?((((m[672]&~m[708]&~m[709]&~m[711]&~m[712])|(~m[672]&~m[708]&~m[709]&m[711]&~m[712])|(m[672]&m[708]&~m[709]&m[711]&~m[712])|(m[672]&~m[708]&m[709]&m[711]&~m[712])|(~m[672]&m[708]&~m[709]&~m[711]&m[712])|(~m[672]&~m[708]&m[709]&~m[711]&m[712])|(m[672]&m[708]&m[709]&~m[711]&m[712])|(~m[672]&m[708]&m[709]&m[711]&m[712]))&UnbiasedRNG[159])|((m[672]&~m[708]&~m[709]&m[711]&~m[712])|(~m[672]&~m[708]&~m[709]&~m[711]&m[712])|(m[672]&~m[708]&~m[709]&~m[711]&m[712])|(m[672]&m[708]&~m[709]&~m[711]&m[712])|(m[672]&~m[708]&m[709]&~m[711]&m[712])|(~m[672]&~m[708]&~m[709]&m[711]&m[712])|(m[672]&~m[708]&~m[709]&m[711]&m[712])|(~m[672]&m[708]&~m[709]&m[711]&m[712])|(m[672]&m[708]&~m[709]&m[711]&m[712])|(~m[672]&~m[708]&m[709]&m[711]&m[712])|(m[672]&~m[708]&m[709]&m[711]&m[712])|(m[672]&m[708]&m[709]&m[711]&m[712]))):InitCond[542];
    m[715] = run?((((m[677]&~m[713]&~m[714]&~m[716]&~m[717])|(~m[677]&~m[713]&~m[714]&m[716]&~m[717])|(m[677]&m[713]&~m[714]&m[716]&~m[717])|(m[677]&~m[713]&m[714]&m[716]&~m[717])|(~m[677]&m[713]&~m[714]&~m[716]&m[717])|(~m[677]&~m[713]&m[714]&~m[716]&m[717])|(m[677]&m[713]&m[714]&~m[716]&m[717])|(~m[677]&m[713]&m[714]&m[716]&m[717]))&UnbiasedRNG[160])|((m[677]&~m[713]&~m[714]&m[716]&~m[717])|(~m[677]&~m[713]&~m[714]&~m[716]&m[717])|(m[677]&~m[713]&~m[714]&~m[716]&m[717])|(m[677]&m[713]&~m[714]&~m[716]&m[717])|(m[677]&~m[713]&m[714]&~m[716]&m[717])|(~m[677]&~m[713]&~m[714]&m[716]&m[717])|(m[677]&~m[713]&~m[714]&m[716]&m[717])|(~m[677]&m[713]&~m[714]&m[716]&m[717])|(m[677]&m[713]&~m[714]&m[716]&m[717])|(~m[677]&~m[713]&m[714]&m[716]&m[717])|(m[677]&~m[713]&m[714]&m[716]&m[717])|(m[677]&m[713]&m[714]&m[716]&m[717]))):InitCond[543];
    m[720] = run?((((m[682]&~m[718]&~m[719]&~m[721]&~m[722])|(~m[682]&~m[718]&~m[719]&m[721]&~m[722])|(m[682]&m[718]&~m[719]&m[721]&~m[722])|(m[682]&~m[718]&m[719]&m[721]&~m[722])|(~m[682]&m[718]&~m[719]&~m[721]&m[722])|(~m[682]&~m[718]&m[719]&~m[721]&m[722])|(m[682]&m[718]&m[719]&~m[721]&m[722])|(~m[682]&m[718]&m[719]&m[721]&m[722]))&UnbiasedRNG[161])|((m[682]&~m[718]&~m[719]&m[721]&~m[722])|(~m[682]&~m[718]&~m[719]&~m[721]&m[722])|(m[682]&~m[718]&~m[719]&~m[721]&m[722])|(m[682]&m[718]&~m[719]&~m[721]&m[722])|(m[682]&~m[718]&m[719]&~m[721]&m[722])|(~m[682]&~m[718]&~m[719]&m[721]&m[722])|(m[682]&~m[718]&~m[719]&m[721]&m[722])|(~m[682]&m[718]&~m[719]&m[721]&m[722])|(m[682]&m[718]&~m[719]&m[721]&m[722])|(~m[682]&~m[718]&m[719]&m[721]&m[722])|(m[682]&~m[718]&m[719]&m[721]&m[722])|(m[682]&m[718]&m[719]&m[721]&m[722]))):InitCond[544];
    m[725] = run?((((m[687]&~m[723]&~m[724]&~m[726]&~m[727])|(~m[687]&~m[723]&~m[724]&m[726]&~m[727])|(m[687]&m[723]&~m[724]&m[726]&~m[727])|(m[687]&~m[723]&m[724]&m[726]&~m[727])|(~m[687]&m[723]&~m[724]&~m[726]&m[727])|(~m[687]&~m[723]&m[724]&~m[726]&m[727])|(m[687]&m[723]&m[724]&~m[726]&m[727])|(~m[687]&m[723]&m[724]&m[726]&m[727]))&UnbiasedRNG[162])|((m[687]&~m[723]&~m[724]&m[726]&~m[727])|(~m[687]&~m[723]&~m[724]&~m[726]&m[727])|(m[687]&~m[723]&~m[724]&~m[726]&m[727])|(m[687]&m[723]&~m[724]&~m[726]&m[727])|(m[687]&~m[723]&m[724]&~m[726]&m[727])|(~m[687]&~m[723]&~m[724]&m[726]&m[727])|(m[687]&~m[723]&~m[724]&m[726]&m[727])|(~m[687]&m[723]&~m[724]&m[726]&m[727])|(m[687]&m[723]&~m[724]&m[726]&m[727])|(~m[687]&~m[723]&m[724]&m[726]&m[727])|(m[687]&~m[723]&m[724]&m[726]&m[727])|(m[687]&m[723]&m[724]&m[726]&m[727]))):InitCond[545];
    m[730] = run?((((m[692]&~m[728]&~m[729]&~m[731]&~m[732])|(~m[692]&~m[728]&~m[729]&m[731]&~m[732])|(m[692]&m[728]&~m[729]&m[731]&~m[732])|(m[692]&~m[728]&m[729]&m[731]&~m[732])|(~m[692]&m[728]&~m[729]&~m[731]&m[732])|(~m[692]&~m[728]&m[729]&~m[731]&m[732])|(m[692]&m[728]&m[729]&~m[731]&m[732])|(~m[692]&m[728]&m[729]&m[731]&m[732]))&UnbiasedRNG[163])|((m[692]&~m[728]&~m[729]&m[731]&~m[732])|(~m[692]&~m[728]&~m[729]&~m[731]&m[732])|(m[692]&~m[728]&~m[729]&~m[731]&m[732])|(m[692]&m[728]&~m[729]&~m[731]&m[732])|(m[692]&~m[728]&m[729]&~m[731]&m[732])|(~m[692]&~m[728]&~m[729]&m[731]&m[732])|(m[692]&~m[728]&~m[729]&m[731]&m[732])|(~m[692]&m[728]&~m[729]&m[731]&m[732])|(m[692]&m[728]&~m[729]&m[731]&m[732])|(~m[692]&~m[728]&m[729]&m[731]&m[732])|(m[692]&~m[728]&m[729]&m[731]&m[732])|(m[692]&m[728]&m[729]&m[731]&m[732]))):InitCond[546];
    m[735] = run?((((m[697]&~m[733]&~m[734]&~m[736]&~m[737])|(~m[697]&~m[733]&~m[734]&m[736]&~m[737])|(m[697]&m[733]&~m[734]&m[736]&~m[737])|(m[697]&~m[733]&m[734]&m[736]&~m[737])|(~m[697]&m[733]&~m[734]&~m[736]&m[737])|(~m[697]&~m[733]&m[734]&~m[736]&m[737])|(m[697]&m[733]&m[734]&~m[736]&m[737])|(~m[697]&m[733]&m[734]&m[736]&m[737]))&UnbiasedRNG[164])|((m[697]&~m[733]&~m[734]&m[736]&~m[737])|(~m[697]&~m[733]&~m[734]&~m[736]&m[737])|(m[697]&~m[733]&~m[734]&~m[736]&m[737])|(m[697]&m[733]&~m[734]&~m[736]&m[737])|(m[697]&~m[733]&m[734]&~m[736]&m[737])|(~m[697]&~m[733]&~m[734]&m[736]&m[737])|(m[697]&~m[733]&~m[734]&m[736]&m[737])|(~m[697]&m[733]&~m[734]&m[736]&m[737])|(m[697]&m[733]&~m[734]&m[736]&m[737])|(~m[697]&~m[733]&m[734]&m[736]&m[737])|(m[697]&~m[733]&m[734]&m[736]&m[737])|(m[697]&m[733]&m[734]&m[736]&m[737]))):InitCond[547];
    m[740] = run?((((m[702]&~m[738]&~m[739]&~m[741]&~m[742])|(~m[702]&~m[738]&~m[739]&m[741]&~m[742])|(m[702]&m[738]&~m[739]&m[741]&~m[742])|(m[702]&~m[738]&m[739]&m[741]&~m[742])|(~m[702]&m[738]&~m[739]&~m[741]&m[742])|(~m[702]&~m[738]&m[739]&~m[741]&m[742])|(m[702]&m[738]&m[739]&~m[741]&m[742])|(~m[702]&m[738]&m[739]&m[741]&m[742]))&UnbiasedRNG[165])|((m[702]&~m[738]&~m[739]&m[741]&~m[742])|(~m[702]&~m[738]&~m[739]&~m[741]&m[742])|(m[702]&~m[738]&~m[739]&~m[741]&m[742])|(m[702]&m[738]&~m[739]&~m[741]&m[742])|(m[702]&~m[738]&m[739]&~m[741]&m[742])|(~m[702]&~m[738]&~m[739]&m[741]&m[742])|(m[702]&~m[738]&~m[739]&m[741]&m[742])|(~m[702]&m[738]&~m[739]&m[741]&m[742])|(m[702]&m[738]&~m[739]&m[741]&m[742])|(~m[702]&~m[738]&m[739]&m[741]&m[742])|(m[702]&~m[738]&m[739]&m[741]&m[742])|(m[702]&m[738]&m[739]&m[741]&m[742]))):InitCond[548];
    m[745] = run?((((m[707]&~m[743]&~m[744]&~m[746]&~m[747])|(~m[707]&~m[743]&~m[744]&m[746]&~m[747])|(m[707]&m[743]&~m[744]&m[746]&~m[747])|(m[707]&~m[743]&m[744]&m[746]&~m[747])|(~m[707]&m[743]&~m[744]&~m[746]&m[747])|(~m[707]&~m[743]&m[744]&~m[746]&m[747])|(m[707]&m[743]&m[744]&~m[746]&m[747])|(~m[707]&m[743]&m[744]&m[746]&m[747]))&UnbiasedRNG[166])|((m[707]&~m[743]&~m[744]&m[746]&~m[747])|(~m[707]&~m[743]&~m[744]&~m[746]&m[747])|(m[707]&~m[743]&~m[744]&~m[746]&m[747])|(m[707]&m[743]&~m[744]&~m[746]&m[747])|(m[707]&~m[743]&m[744]&~m[746]&m[747])|(~m[707]&~m[743]&~m[744]&m[746]&m[747])|(m[707]&~m[743]&~m[744]&m[746]&m[747])|(~m[707]&m[743]&~m[744]&m[746]&m[747])|(m[707]&m[743]&~m[744]&m[746]&m[747])|(~m[707]&~m[743]&m[744]&m[746]&m[747])|(m[707]&~m[743]&m[744]&m[746]&m[747])|(m[707]&m[743]&m[744]&m[746]&m[747]))):InitCond[549];
    m[755] = run?((((m[712]&~m[753]&~m[754]&~m[756]&~m[757])|(~m[712]&~m[753]&~m[754]&m[756]&~m[757])|(m[712]&m[753]&~m[754]&m[756]&~m[757])|(m[712]&~m[753]&m[754]&m[756]&~m[757])|(~m[712]&m[753]&~m[754]&~m[756]&m[757])|(~m[712]&~m[753]&m[754]&~m[756]&m[757])|(m[712]&m[753]&m[754]&~m[756]&m[757])|(~m[712]&m[753]&m[754]&m[756]&m[757]))&UnbiasedRNG[167])|((m[712]&~m[753]&~m[754]&m[756]&~m[757])|(~m[712]&~m[753]&~m[754]&~m[756]&m[757])|(m[712]&~m[753]&~m[754]&~m[756]&m[757])|(m[712]&m[753]&~m[754]&~m[756]&m[757])|(m[712]&~m[753]&m[754]&~m[756]&m[757])|(~m[712]&~m[753]&~m[754]&m[756]&m[757])|(m[712]&~m[753]&~m[754]&m[756]&m[757])|(~m[712]&m[753]&~m[754]&m[756]&m[757])|(m[712]&m[753]&~m[754]&m[756]&m[757])|(~m[712]&~m[753]&m[754]&m[756]&m[757])|(m[712]&~m[753]&m[754]&m[756]&m[757])|(m[712]&m[753]&m[754]&m[756]&m[757]))):InitCond[550];
    m[760] = run?((((m[717]&~m[758]&~m[759]&~m[761]&~m[762])|(~m[717]&~m[758]&~m[759]&m[761]&~m[762])|(m[717]&m[758]&~m[759]&m[761]&~m[762])|(m[717]&~m[758]&m[759]&m[761]&~m[762])|(~m[717]&m[758]&~m[759]&~m[761]&m[762])|(~m[717]&~m[758]&m[759]&~m[761]&m[762])|(m[717]&m[758]&m[759]&~m[761]&m[762])|(~m[717]&m[758]&m[759]&m[761]&m[762]))&UnbiasedRNG[168])|((m[717]&~m[758]&~m[759]&m[761]&~m[762])|(~m[717]&~m[758]&~m[759]&~m[761]&m[762])|(m[717]&~m[758]&~m[759]&~m[761]&m[762])|(m[717]&m[758]&~m[759]&~m[761]&m[762])|(m[717]&~m[758]&m[759]&~m[761]&m[762])|(~m[717]&~m[758]&~m[759]&m[761]&m[762])|(m[717]&~m[758]&~m[759]&m[761]&m[762])|(~m[717]&m[758]&~m[759]&m[761]&m[762])|(m[717]&m[758]&~m[759]&m[761]&m[762])|(~m[717]&~m[758]&m[759]&m[761]&m[762])|(m[717]&~m[758]&m[759]&m[761]&m[762])|(m[717]&m[758]&m[759]&m[761]&m[762]))):InitCond[551];
    m[765] = run?((((m[722]&~m[763]&~m[764]&~m[766]&~m[767])|(~m[722]&~m[763]&~m[764]&m[766]&~m[767])|(m[722]&m[763]&~m[764]&m[766]&~m[767])|(m[722]&~m[763]&m[764]&m[766]&~m[767])|(~m[722]&m[763]&~m[764]&~m[766]&m[767])|(~m[722]&~m[763]&m[764]&~m[766]&m[767])|(m[722]&m[763]&m[764]&~m[766]&m[767])|(~m[722]&m[763]&m[764]&m[766]&m[767]))&UnbiasedRNG[169])|((m[722]&~m[763]&~m[764]&m[766]&~m[767])|(~m[722]&~m[763]&~m[764]&~m[766]&m[767])|(m[722]&~m[763]&~m[764]&~m[766]&m[767])|(m[722]&m[763]&~m[764]&~m[766]&m[767])|(m[722]&~m[763]&m[764]&~m[766]&m[767])|(~m[722]&~m[763]&~m[764]&m[766]&m[767])|(m[722]&~m[763]&~m[764]&m[766]&m[767])|(~m[722]&m[763]&~m[764]&m[766]&m[767])|(m[722]&m[763]&~m[764]&m[766]&m[767])|(~m[722]&~m[763]&m[764]&m[766]&m[767])|(m[722]&~m[763]&m[764]&m[766]&m[767])|(m[722]&m[763]&m[764]&m[766]&m[767]))):InitCond[552];
    m[770] = run?((((m[727]&~m[768]&~m[769]&~m[771]&~m[772])|(~m[727]&~m[768]&~m[769]&m[771]&~m[772])|(m[727]&m[768]&~m[769]&m[771]&~m[772])|(m[727]&~m[768]&m[769]&m[771]&~m[772])|(~m[727]&m[768]&~m[769]&~m[771]&m[772])|(~m[727]&~m[768]&m[769]&~m[771]&m[772])|(m[727]&m[768]&m[769]&~m[771]&m[772])|(~m[727]&m[768]&m[769]&m[771]&m[772]))&UnbiasedRNG[170])|((m[727]&~m[768]&~m[769]&m[771]&~m[772])|(~m[727]&~m[768]&~m[769]&~m[771]&m[772])|(m[727]&~m[768]&~m[769]&~m[771]&m[772])|(m[727]&m[768]&~m[769]&~m[771]&m[772])|(m[727]&~m[768]&m[769]&~m[771]&m[772])|(~m[727]&~m[768]&~m[769]&m[771]&m[772])|(m[727]&~m[768]&~m[769]&m[771]&m[772])|(~m[727]&m[768]&~m[769]&m[771]&m[772])|(m[727]&m[768]&~m[769]&m[771]&m[772])|(~m[727]&~m[768]&m[769]&m[771]&m[772])|(m[727]&~m[768]&m[769]&m[771]&m[772])|(m[727]&m[768]&m[769]&m[771]&m[772]))):InitCond[553];
    m[775] = run?((((m[732]&~m[773]&~m[774]&~m[776]&~m[777])|(~m[732]&~m[773]&~m[774]&m[776]&~m[777])|(m[732]&m[773]&~m[774]&m[776]&~m[777])|(m[732]&~m[773]&m[774]&m[776]&~m[777])|(~m[732]&m[773]&~m[774]&~m[776]&m[777])|(~m[732]&~m[773]&m[774]&~m[776]&m[777])|(m[732]&m[773]&m[774]&~m[776]&m[777])|(~m[732]&m[773]&m[774]&m[776]&m[777]))&UnbiasedRNG[171])|((m[732]&~m[773]&~m[774]&m[776]&~m[777])|(~m[732]&~m[773]&~m[774]&~m[776]&m[777])|(m[732]&~m[773]&~m[774]&~m[776]&m[777])|(m[732]&m[773]&~m[774]&~m[776]&m[777])|(m[732]&~m[773]&m[774]&~m[776]&m[777])|(~m[732]&~m[773]&~m[774]&m[776]&m[777])|(m[732]&~m[773]&~m[774]&m[776]&m[777])|(~m[732]&m[773]&~m[774]&m[776]&m[777])|(m[732]&m[773]&~m[774]&m[776]&m[777])|(~m[732]&~m[773]&m[774]&m[776]&m[777])|(m[732]&~m[773]&m[774]&m[776]&m[777])|(m[732]&m[773]&m[774]&m[776]&m[777]))):InitCond[554];
    m[780] = run?((((m[737]&~m[778]&~m[779]&~m[781]&~m[782])|(~m[737]&~m[778]&~m[779]&m[781]&~m[782])|(m[737]&m[778]&~m[779]&m[781]&~m[782])|(m[737]&~m[778]&m[779]&m[781]&~m[782])|(~m[737]&m[778]&~m[779]&~m[781]&m[782])|(~m[737]&~m[778]&m[779]&~m[781]&m[782])|(m[737]&m[778]&m[779]&~m[781]&m[782])|(~m[737]&m[778]&m[779]&m[781]&m[782]))&UnbiasedRNG[172])|((m[737]&~m[778]&~m[779]&m[781]&~m[782])|(~m[737]&~m[778]&~m[779]&~m[781]&m[782])|(m[737]&~m[778]&~m[779]&~m[781]&m[782])|(m[737]&m[778]&~m[779]&~m[781]&m[782])|(m[737]&~m[778]&m[779]&~m[781]&m[782])|(~m[737]&~m[778]&~m[779]&m[781]&m[782])|(m[737]&~m[778]&~m[779]&m[781]&m[782])|(~m[737]&m[778]&~m[779]&m[781]&m[782])|(m[737]&m[778]&~m[779]&m[781]&m[782])|(~m[737]&~m[778]&m[779]&m[781]&m[782])|(m[737]&~m[778]&m[779]&m[781]&m[782])|(m[737]&m[778]&m[779]&m[781]&m[782]))):InitCond[555];
    m[785] = run?((((m[742]&~m[783]&~m[784]&~m[786]&~m[787])|(~m[742]&~m[783]&~m[784]&m[786]&~m[787])|(m[742]&m[783]&~m[784]&m[786]&~m[787])|(m[742]&~m[783]&m[784]&m[786]&~m[787])|(~m[742]&m[783]&~m[784]&~m[786]&m[787])|(~m[742]&~m[783]&m[784]&~m[786]&m[787])|(m[742]&m[783]&m[784]&~m[786]&m[787])|(~m[742]&m[783]&m[784]&m[786]&m[787]))&UnbiasedRNG[173])|((m[742]&~m[783]&~m[784]&m[786]&~m[787])|(~m[742]&~m[783]&~m[784]&~m[786]&m[787])|(m[742]&~m[783]&~m[784]&~m[786]&m[787])|(m[742]&m[783]&~m[784]&~m[786]&m[787])|(m[742]&~m[783]&m[784]&~m[786]&m[787])|(~m[742]&~m[783]&~m[784]&m[786]&m[787])|(m[742]&~m[783]&~m[784]&m[786]&m[787])|(~m[742]&m[783]&~m[784]&m[786]&m[787])|(m[742]&m[783]&~m[784]&m[786]&m[787])|(~m[742]&~m[783]&m[784]&m[786]&m[787])|(m[742]&~m[783]&m[784]&m[786]&m[787])|(m[742]&m[783]&m[784]&m[786]&m[787]))):InitCond[556];
    m[790] = run?((((m[747]&~m[788]&~m[789]&~m[791]&~m[792])|(~m[747]&~m[788]&~m[789]&m[791]&~m[792])|(m[747]&m[788]&~m[789]&m[791]&~m[792])|(m[747]&~m[788]&m[789]&m[791]&~m[792])|(~m[747]&m[788]&~m[789]&~m[791]&m[792])|(~m[747]&~m[788]&m[789]&~m[791]&m[792])|(m[747]&m[788]&m[789]&~m[791]&m[792])|(~m[747]&m[788]&m[789]&m[791]&m[792]))&UnbiasedRNG[174])|((m[747]&~m[788]&~m[789]&m[791]&~m[792])|(~m[747]&~m[788]&~m[789]&~m[791]&m[792])|(m[747]&~m[788]&~m[789]&~m[791]&m[792])|(m[747]&m[788]&~m[789]&~m[791]&m[792])|(m[747]&~m[788]&m[789]&~m[791]&m[792])|(~m[747]&~m[788]&~m[789]&m[791]&m[792])|(m[747]&~m[788]&~m[789]&m[791]&m[792])|(~m[747]&m[788]&~m[789]&m[791]&m[792])|(m[747]&m[788]&~m[789]&m[791]&m[792])|(~m[747]&~m[788]&m[789]&m[791]&m[792])|(m[747]&~m[788]&m[789]&m[791]&m[792])|(m[747]&m[788]&m[789]&m[791]&m[792]))):InitCond[557];
    m[795] = run?((((m[752]&~m[793]&~m[794]&~m[796]&~m[797])|(~m[752]&~m[793]&~m[794]&m[796]&~m[797])|(m[752]&m[793]&~m[794]&m[796]&~m[797])|(m[752]&~m[793]&m[794]&m[796]&~m[797])|(~m[752]&m[793]&~m[794]&~m[796]&m[797])|(~m[752]&~m[793]&m[794]&~m[796]&m[797])|(m[752]&m[793]&m[794]&~m[796]&m[797])|(~m[752]&m[793]&m[794]&m[796]&m[797]))&UnbiasedRNG[175])|((m[752]&~m[793]&~m[794]&m[796]&~m[797])|(~m[752]&~m[793]&~m[794]&~m[796]&m[797])|(m[752]&~m[793]&~m[794]&~m[796]&m[797])|(m[752]&m[793]&~m[794]&~m[796]&m[797])|(m[752]&~m[793]&m[794]&~m[796]&m[797])|(~m[752]&~m[793]&~m[794]&m[796]&m[797])|(m[752]&~m[793]&~m[794]&m[796]&m[797])|(~m[752]&m[793]&~m[794]&m[796]&m[797])|(m[752]&m[793]&~m[794]&m[796]&m[797])|(~m[752]&~m[793]&m[794]&m[796]&m[797])|(m[752]&~m[793]&m[794]&m[796]&m[797])|(m[752]&m[793]&m[794]&m[796]&m[797]))):InitCond[558];
    m[805] = run?((((m[757]&~m[803]&~m[804]&~m[806]&~m[807])|(~m[757]&~m[803]&~m[804]&m[806]&~m[807])|(m[757]&m[803]&~m[804]&m[806]&~m[807])|(m[757]&~m[803]&m[804]&m[806]&~m[807])|(~m[757]&m[803]&~m[804]&~m[806]&m[807])|(~m[757]&~m[803]&m[804]&~m[806]&m[807])|(m[757]&m[803]&m[804]&~m[806]&m[807])|(~m[757]&m[803]&m[804]&m[806]&m[807]))&UnbiasedRNG[176])|((m[757]&~m[803]&~m[804]&m[806]&~m[807])|(~m[757]&~m[803]&~m[804]&~m[806]&m[807])|(m[757]&~m[803]&~m[804]&~m[806]&m[807])|(m[757]&m[803]&~m[804]&~m[806]&m[807])|(m[757]&~m[803]&m[804]&~m[806]&m[807])|(~m[757]&~m[803]&~m[804]&m[806]&m[807])|(m[757]&~m[803]&~m[804]&m[806]&m[807])|(~m[757]&m[803]&~m[804]&m[806]&m[807])|(m[757]&m[803]&~m[804]&m[806]&m[807])|(~m[757]&~m[803]&m[804]&m[806]&m[807])|(m[757]&~m[803]&m[804]&m[806]&m[807])|(m[757]&m[803]&m[804]&m[806]&m[807]))):InitCond[559];
    m[810] = run?((((m[762]&~m[808]&~m[809]&~m[811]&~m[812])|(~m[762]&~m[808]&~m[809]&m[811]&~m[812])|(m[762]&m[808]&~m[809]&m[811]&~m[812])|(m[762]&~m[808]&m[809]&m[811]&~m[812])|(~m[762]&m[808]&~m[809]&~m[811]&m[812])|(~m[762]&~m[808]&m[809]&~m[811]&m[812])|(m[762]&m[808]&m[809]&~m[811]&m[812])|(~m[762]&m[808]&m[809]&m[811]&m[812]))&UnbiasedRNG[177])|((m[762]&~m[808]&~m[809]&m[811]&~m[812])|(~m[762]&~m[808]&~m[809]&~m[811]&m[812])|(m[762]&~m[808]&~m[809]&~m[811]&m[812])|(m[762]&m[808]&~m[809]&~m[811]&m[812])|(m[762]&~m[808]&m[809]&~m[811]&m[812])|(~m[762]&~m[808]&~m[809]&m[811]&m[812])|(m[762]&~m[808]&~m[809]&m[811]&m[812])|(~m[762]&m[808]&~m[809]&m[811]&m[812])|(m[762]&m[808]&~m[809]&m[811]&m[812])|(~m[762]&~m[808]&m[809]&m[811]&m[812])|(m[762]&~m[808]&m[809]&m[811]&m[812])|(m[762]&m[808]&m[809]&m[811]&m[812]))):InitCond[560];
    m[815] = run?((((m[767]&~m[813]&~m[814]&~m[816]&~m[817])|(~m[767]&~m[813]&~m[814]&m[816]&~m[817])|(m[767]&m[813]&~m[814]&m[816]&~m[817])|(m[767]&~m[813]&m[814]&m[816]&~m[817])|(~m[767]&m[813]&~m[814]&~m[816]&m[817])|(~m[767]&~m[813]&m[814]&~m[816]&m[817])|(m[767]&m[813]&m[814]&~m[816]&m[817])|(~m[767]&m[813]&m[814]&m[816]&m[817]))&UnbiasedRNG[178])|((m[767]&~m[813]&~m[814]&m[816]&~m[817])|(~m[767]&~m[813]&~m[814]&~m[816]&m[817])|(m[767]&~m[813]&~m[814]&~m[816]&m[817])|(m[767]&m[813]&~m[814]&~m[816]&m[817])|(m[767]&~m[813]&m[814]&~m[816]&m[817])|(~m[767]&~m[813]&~m[814]&m[816]&m[817])|(m[767]&~m[813]&~m[814]&m[816]&m[817])|(~m[767]&m[813]&~m[814]&m[816]&m[817])|(m[767]&m[813]&~m[814]&m[816]&m[817])|(~m[767]&~m[813]&m[814]&m[816]&m[817])|(m[767]&~m[813]&m[814]&m[816]&m[817])|(m[767]&m[813]&m[814]&m[816]&m[817]))):InitCond[561];
    m[820] = run?((((m[772]&~m[818]&~m[819]&~m[821]&~m[822])|(~m[772]&~m[818]&~m[819]&m[821]&~m[822])|(m[772]&m[818]&~m[819]&m[821]&~m[822])|(m[772]&~m[818]&m[819]&m[821]&~m[822])|(~m[772]&m[818]&~m[819]&~m[821]&m[822])|(~m[772]&~m[818]&m[819]&~m[821]&m[822])|(m[772]&m[818]&m[819]&~m[821]&m[822])|(~m[772]&m[818]&m[819]&m[821]&m[822]))&UnbiasedRNG[179])|((m[772]&~m[818]&~m[819]&m[821]&~m[822])|(~m[772]&~m[818]&~m[819]&~m[821]&m[822])|(m[772]&~m[818]&~m[819]&~m[821]&m[822])|(m[772]&m[818]&~m[819]&~m[821]&m[822])|(m[772]&~m[818]&m[819]&~m[821]&m[822])|(~m[772]&~m[818]&~m[819]&m[821]&m[822])|(m[772]&~m[818]&~m[819]&m[821]&m[822])|(~m[772]&m[818]&~m[819]&m[821]&m[822])|(m[772]&m[818]&~m[819]&m[821]&m[822])|(~m[772]&~m[818]&m[819]&m[821]&m[822])|(m[772]&~m[818]&m[819]&m[821]&m[822])|(m[772]&m[818]&m[819]&m[821]&m[822]))):InitCond[562];
    m[825] = run?((((m[777]&~m[823]&~m[824]&~m[826]&~m[827])|(~m[777]&~m[823]&~m[824]&m[826]&~m[827])|(m[777]&m[823]&~m[824]&m[826]&~m[827])|(m[777]&~m[823]&m[824]&m[826]&~m[827])|(~m[777]&m[823]&~m[824]&~m[826]&m[827])|(~m[777]&~m[823]&m[824]&~m[826]&m[827])|(m[777]&m[823]&m[824]&~m[826]&m[827])|(~m[777]&m[823]&m[824]&m[826]&m[827]))&UnbiasedRNG[180])|((m[777]&~m[823]&~m[824]&m[826]&~m[827])|(~m[777]&~m[823]&~m[824]&~m[826]&m[827])|(m[777]&~m[823]&~m[824]&~m[826]&m[827])|(m[777]&m[823]&~m[824]&~m[826]&m[827])|(m[777]&~m[823]&m[824]&~m[826]&m[827])|(~m[777]&~m[823]&~m[824]&m[826]&m[827])|(m[777]&~m[823]&~m[824]&m[826]&m[827])|(~m[777]&m[823]&~m[824]&m[826]&m[827])|(m[777]&m[823]&~m[824]&m[826]&m[827])|(~m[777]&~m[823]&m[824]&m[826]&m[827])|(m[777]&~m[823]&m[824]&m[826]&m[827])|(m[777]&m[823]&m[824]&m[826]&m[827]))):InitCond[563];
    m[830] = run?((((m[782]&~m[828]&~m[829]&~m[831]&~m[832])|(~m[782]&~m[828]&~m[829]&m[831]&~m[832])|(m[782]&m[828]&~m[829]&m[831]&~m[832])|(m[782]&~m[828]&m[829]&m[831]&~m[832])|(~m[782]&m[828]&~m[829]&~m[831]&m[832])|(~m[782]&~m[828]&m[829]&~m[831]&m[832])|(m[782]&m[828]&m[829]&~m[831]&m[832])|(~m[782]&m[828]&m[829]&m[831]&m[832]))&UnbiasedRNG[181])|((m[782]&~m[828]&~m[829]&m[831]&~m[832])|(~m[782]&~m[828]&~m[829]&~m[831]&m[832])|(m[782]&~m[828]&~m[829]&~m[831]&m[832])|(m[782]&m[828]&~m[829]&~m[831]&m[832])|(m[782]&~m[828]&m[829]&~m[831]&m[832])|(~m[782]&~m[828]&~m[829]&m[831]&m[832])|(m[782]&~m[828]&~m[829]&m[831]&m[832])|(~m[782]&m[828]&~m[829]&m[831]&m[832])|(m[782]&m[828]&~m[829]&m[831]&m[832])|(~m[782]&~m[828]&m[829]&m[831]&m[832])|(m[782]&~m[828]&m[829]&m[831]&m[832])|(m[782]&m[828]&m[829]&m[831]&m[832]))):InitCond[564];
    m[835] = run?((((m[787]&~m[833]&~m[834]&~m[836]&~m[837])|(~m[787]&~m[833]&~m[834]&m[836]&~m[837])|(m[787]&m[833]&~m[834]&m[836]&~m[837])|(m[787]&~m[833]&m[834]&m[836]&~m[837])|(~m[787]&m[833]&~m[834]&~m[836]&m[837])|(~m[787]&~m[833]&m[834]&~m[836]&m[837])|(m[787]&m[833]&m[834]&~m[836]&m[837])|(~m[787]&m[833]&m[834]&m[836]&m[837]))&UnbiasedRNG[182])|((m[787]&~m[833]&~m[834]&m[836]&~m[837])|(~m[787]&~m[833]&~m[834]&~m[836]&m[837])|(m[787]&~m[833]&~m[834]&~m[836]&m[837])|(m[787]&m[833]&~m[834]&~m[836]&m[837])|(m[787]&~m[833]&m[834]&~m[836]&m[837])|(~m[787]&~m[833]&~m[834]&m[836]&m[837])|(m[787]&~m[833]&~m[834]&m[836]&m[837])|(~m[787]&m[833]&~m[834]&m[836]&m[837])|(m[787]&m[833]&~m[834]&m[836]&m[837])|(~m[787]&~m[833]&m[834]&m[836]&m[837])|(m[787]&~m[833]&m[834]&m[836]&m[837])|(m[787]&m[833]&m[834]&m[836]&m[837]))):InitCond[565];
    m[840] = run?((((m[792]&~m[838]&~m[839]&~m[841]&~m[842])|(~m[792]&~m[838]&~m[839]&m[841]&~m[842])|(m[792]&m[838]&~m[839]&m[841]&~m[842])|(m[792]&~m[838]&m[839]&m[841]&~m[842])|(~m[792]&m[838]&~m[839]&~m[841]&m[842])|(~m[792]&~m[838]&m[839]&~m[841]&m[842])|(m[792]&m[838]&m[839]&~m[841]&m[842])|(~m[792]&m[838]&m[839]&m[841]&m[842]))&UnbiasedRNG[183])|((m[792]&~m[838]&~m[839]&m[841]&~m[842])|(~m[792]&~m[838]&~m[839]&~m[841]&m[842])|(m[792]&~m[838]&~m[839]&~m[841]&m[842])|(m[792]&m[838]&~m[839]&~m[841]&m[842])|(m[792]&~m[838]&m[839]&~m[841]&m[842])|(~m[792]&~m[838]&~m[839]&m[841]&m[842])|(m[792]&~m[838]&~m[839]&m[841]&m[842])|(~m[792]&m[838]&~m[839]&m[841]&m[842])|(m[792]&m[838]&~m[839]&m[841]&m[842])|(~m[792]&~m[838]&m[839]&m[841]&m[842])|(m[792]&~m[838]&m[839]&m[841]&m[842])|(m[792]&m[838]&m[839]&m[841]&m[842]))):InitCond[566];
    m[845] = run?((((m[797]&~m[843]&~m[844]&~m[846]&~m[847])|(~m[797]&~m[843]&~m[844]&m[846]&~m[847])|(m[797]&m[843]&~m[844]&m[846]&~m[847])|(m[797]&~m[843]&m[844]&m[846]&~m[847])|(~m[797]&m[843]&~m[844]&~m[846]&m[847])|(~m[797]&~m[843]&m[844]&~m[846]&m[847])|(m[797]&m[843]&m[844]&~m[846]&m[847])|(~m[797]&m[843]&m[844]&m[846]&m[847]))&UnbiasedRNG[184])|((m[797]&~m[843]&~m[844]&m[846]&~m[847])|(~m[797]&~m[843]&~m[844]&~m[846]&m[847])|(m[797]&~m[843]&~m[844]&~m[846]&m[847])|(m[797]&m[843]&~m[844]&~m[846]&m[847])|(m[797]&~m[843]&m[844]&~m[846]&m[847])|(~m[797]&~m[843]&~m[844]&m[846]&m[847])|(m[797]&~m[843]&~m[844]&m[846]&m[847])|(~m[797]&m[843]&~m[844]&m[846]&m[847])|(m[797]&m[843]&~m[844]&m[846]&m[847])|(~m[797]&~m[843]&m[844]&m[846]&m[847])|(m[797]&~m[843]&m[844]&m[846]&m[847])|(m[797]&m[843]&m[844]&m[846]&m[847]))):InitCond[567];
    m[850] = run?((((m[802]&~m[848]&~m[849]&~m[851]&~m[852])|(~m[802]&~m[848]&~m[849]&m[851]&~m[852])|(m[802]&m[848]&~m[849]&m[851]&~m[852])|(m[802]&~m[848]&m[849]&m[851]&~m[852])|(~m[802]&m[848]&~m[849]&~m[851]&m[852])|(~m[802]&~m[848]&m[849]&~m[851]&m[852])|(m[802]&m[848]&m[849]&~m[851]&m[852])|(~m[802]&m[848]&m[849]&m[851]&m[852]))&UnbiasedRNG[185])|((m[802]&~m[848]&~m[849]&m[851]&~m[852])|(~m[802]&~m[848]&~m[849]&~m[851]&m[852])|(m[802]&~m[848]&~m[849]&~m[851]&m[852])|(m[802]&m[848]&~m[849]&~m[851]&m[852])|(m[802]&~m[848]&m[849]&~m[851]&m[852])|(~m[802]&~m[848]&~m[849]&m[851]&m[852])|(m[802]&~m[848]&~m[849]&m[851]&m[852])|(~m[802]&m[848]&~m[849]&m[851]&m[852])|(m[802]&m[848]&~m[849]&m[851]&m[852])|(~m[802]&~m[848]&m[849]&m[851]&m[852])|(m[802]&~m[848]&m[849]&m[851]&m[852])|(m[802]&m[848]&m[849]&m[851]&m[852]))):InitCond[568];
    m[860] = run?((((m[807]&~m[858]&~m[859]&~m[861]&~m[862])|(~m[807]&~m[858]&~m[859]&m[861]&~m[862])|(m[807]&m[858]&~m[859]&m[861]&~m[862])|(m[807]&~m[858]&m[859]&m[861]&~m[862])|(~m[807]&m[858]&~m[859]&~m[861]&m[862])|(~m[807]&~m[858]&m[859]&~m[861]&m[862])|(m[807]&m[858]&m[859]&~m[861]&m[862])|(~m[807]&m[858]&m[859]&m[861]&m[862]))&UnbiasedRNG[186])|((m[807]&~m[858]&~m[859]&m[861]&~m[862])|(~m[807]&~m[858]&~m[859]&~m[861]&m[862])|(m[807]&~m[858]&~m[859]&~m[861]&m[862])|(m[807]&m[858]&~m[859]&~m[861]&m[862])|(m[807]&~m[858]&m[859]&~m[861]&m[862])|(~m[807]&~m[858]&~m[859]&m[861]&m[862])|(m[807]&~m[858]&~m[859]&m[861]&m[862])|(~m[807]&m[858]&~m[859]&m[861]&m[862])|(m[807]&m[858]&~m[859]&m[861]&m[862])|(~m[807]&~m[858]&m[859]&m[861]&m[862])|(m[807]&~m[858]&m[859]&m[861]&m[862])|(m[807]&m[858]&m[859]&m[861]&m[862]))):InitCond[569];
    m[865] = run?((((m[812]&~m[863]&~m[864]&~m[866]&~m[867])|(~m[812]&~m[863]&~m[864]&m[866]&~m[867])|(m[812]&m[863]&~m[864]&m[866]&~m[867])|(m[812]&~m[863]&m[864]&m[866]&~m[867])|(~m[812]&m[863]&~m[864]&~m[866]&m[867])|(~m[812]&~m[863]&m[864]&~m[866]&m[867])|(m[812]&m[863]&m[864]&~m[866]&m[867])|(~m[812]&m[863]&m[864]&m[866]&m[867]))&UnbiasedRNG[187])|((m[812]&~m[863]&~m[864]&m[866]&~m[867])|(~m[812]&~m[863]&~m[864]&~m[866]&m[867])|(m[812]&~m[863]&~m[864]&~m[866]&m[867])|(m[812]&m[863]&~m[864]&~m[866]&m[867])|(m[812]&~m[863]&m[864]&~m[866]&m[867])|(~m[812]&~m[863]&~m[864]&m[866]&m[867])|(m[812]&~m[863]&~m[864]&m[866]&m[867])|(~m[812]&m[863]&~m[864]&m[866]&m[867])|(m[812]&m[863]&~m[864]&m[866]&m[867])|(~m[812]&~m[863]&m[864]&m[866]&m[867])|(m[812]&~m[863]&m[864]&m[866]&m[867])|(m[812]&m[863]&m[864]&m[866]&m[867]))):InitCond[570];
    m[870] = run?((((m[817]&~m[868]&~m[869]&~m[871]&~m[872])|(~m[817]&~m[868]&~m[869]&m[871]&~m[872])|(m[817]&m[868]&~m[869]&m[871]&~m[872])|(m[817]&~m[868]&m[869]&m[871]&~m[872])|(~m[817]&m[868]&~m[869]&~m[871]&m[872])|(~m[817]&~m[868]&m[869]&~m[871]&m[872])|(m[817]&m[868]&m[869]&~m[871]&m[872])|(~m[817]&m[868]&m[869]&m[871]&m[872]))&UnbiasedRNG[188])|((m[817]&~m[868]&~m[869]&m[871]&~m[872])|(~m[817]&~m[868]&~m[869]&~m[871]&m[872])|(m[817]&~m[868]&~m[869]&~m[871]&m[872])|(m[817]&m[868]&~m[869]&~m[871]&m[872])|(m[817]&~m[868]&m[869]&~m[871]&m[872])|(~m[817]&~m[868]&~m[869]&m[871]&m[872])|(m[817]&~m[868]&~m[869]&m[871]&m[872])|(~m[817]&m[868]&~m[869]&m[871]&m[872])|(m[817]&m[868]&~m[869]&m[871]&m[872])|(~m[817]&~m[868]&m[869]&m[871]&m[872])|(m[817]&~m[868]&m[869]&m[871]&m[872])|(m[817]&m[868]&m[869]&m[871]&m[872]))):InitCond[571];
    m[875] = run?((((m[822]&~m[873]&~m[874]&~m[876]&~m[877])|(~m[822]&~m[873]&~m[874]&m[876]&~m[877])|(m[822]&m[873]&~m[874]&m[876]&~m[877])|(m[822]&~m[873]&m[874]&m[876]&~m[877])|(~m[822]&m[873]&~m[874]&~m[876]&m[877])|(~m[822]&~m[873]&m[874]&~m[876]&m[877])|(m[822]&m[873]&m[874]&~m[876]&m[877])|(~m[822]&m[873]&m[874]&m[876]&m[877]))&UnbiasedRNG[189])|((m[822]&~m[873]&~m[874]&m[876]&~m[877])|(~m[822]&~m[873]&~m[874]&~m[876]&m[877])|(m[822]&~m[873]&~m[874]&~m[876]&m[877])|(m[822]&m[873]&~m[874]&~m[876]&m[877])|(m[822]&~m[873]&m[874]&~m[876]&m[877])|(~m[822]&~m[873]&~m[874]&m[876]&m[877])|(m[822]&~m[873]&~m[874]&m[876]&m[877])|(~m[822]&m[873]&~m[874]&m[876]&m[877])|(m[822]&m[873]&~m[874]&m[876]&m[877])|(~m[822]&~m[873]&m[874]&m[876]&m[877])|(m[822]&~m[873]&m[874]&m[876]&m[877])|(m[822]&m[873]&m[874]&m[876]&m[877]))):InitCond[572];
    m[880] = run?((((m[827]&~m[878]&~m[879]&~m[881]&~m[882])|(~m[827]&~m[878]&~m[879]&m[881]&~m[882])|(m[827]&m[878]&~m[879]&m[881]&~m[882])|(m[827]&~m[878]&m[879]&m[881]&~m[882])|(~m[827]&m[878]&~m[879]&~m[881]&m[882])|(~m[827]&~m[878]&m[879]&~m[881]&m[882])|(m[827]&m[878]&m[879]&~m[881]&m[882])|(~m[827]&m[878]&m[879]&m[881]&m[882]))&UnbiasedRNG[190])|((m[827]&~m[878]&~m[879]&m[881]&~m[882])|(~m[827]&~m[878]&~m[879]&~m[881]&m[882])|(m[827]&~m[878]&~m[879]&~m[881]&m[882])|(m[827]&m[878]&~m[879]&~m[881]&m[882])|(m[827]&~m[878]&m[879]&~m[881]&m[882])|(~m[827]&~m[878]&~m[879]&m[881]&m[882])|(m[827]&~m[878]&~m[879]&m[881]&m[882])|(~m[827]&m[878]&~m[879]&m[881]&m[882])|(m[827]&m[878]&~m[879]&m[881]&m[882])|(~m[827]&~m[878]&m[879]&m[881]&m[882])|(m[827]&~m[878]&m[879]&m[881]&m[882])|(m[827]&m[878]&m[879]&m[881]&m[882]))):InitCond[573];
    m[885] = run?((((m[832]&~m[883]&~m[884]&~m[886]&~m[887])|(~m[832]&~m[883]&~m[884]&m[886]&~m[887])|(m[832]&m[883]&~m[884]&m[886]&~m[887])|(m[832]&~m[883]&m[884]&m[886]&~m[887])|(~m[832]&m[883]&~m[884]&~m[886]&m[887])|(~m[832]&~m[883]&m[884]&~m[886]&m[887])|(m[832]&m[883]&m[884]&~m[886]&m[887])|(~m[832]&m[883]&m[884]&m[886]&m[887]))&UnbiasedRNG[191])|((m[832]&~m[883]&~m[884]&m[886]&~m[887])|(~m[832]&~m[883]&~m[884]&~m[886]&m[887])|(m[832]&~m[883]&~m[884]&~m[886]&m[887])|(m[832]&m[883]&~m[884]&~m[886]&m[887])|(m[832]&~m[883]&m[884]&~m[886]&m[887])|(~m[832]&~m[883]&~m[884]&m[886]&m[887])|(m[832]&~m[883]&~m[884]&m[886]&m[887])|(~m[832]&m[883]&~m[884]&m[886]&m[887])|(m[832]&m[883]&~m[884]&m[886]&m[887])|(~m[832]&~m[883]&m[884]&m[886]&m[887])|(m[832]&~m[883]&m[884]&m[886]&m[887])|(m[832]&m[883]&m[884]&m[886]&m[887]))):InitCond[574];
    m[890] = run?((((m[837]&~m[888]&~m[889]&~m[891]&~m[892])|(~m[837]&~m[888]&~m[889]&m[891]&~m[892])|(m[837]&m[888]&~m[889]&m[891]&~m[892])|(m[837]&~m[888]&m[889]&m[891]&~m[892])|(~m[837]&m[888]&~m[889]&~m[891]&m[892])|(~m[837]&~m[888]&m[889]&~m[891]&m[892])|(m[837]&m[888]&m[889]&~m[891]&m[892])|(~m[837]&m[888]&m[889]&m[891]&m[892]))&UnbiasedRNG[192])|((m[837]&~m[888]&~m[889]&m[891]&~m[892])|(~m[837]&~m[888]&~m[889]&~m[891]&m[892])|(m[837]&~m[888]&~m[889]&~m[891]&m[892])|(m[837]&m[888]&~m[889]&~m[891]&m[892])|(m[837]&~m[888]&m[889]&~m[891]&m[892])|(~m[837]&~m[888]&~m[889]&m[891]&m[892])|(m[837]&~m[888]&~m[889]&m[891]&m[892])|(~m[837]&m[888]&~m[889]&m[891]&m[892])|(m[837]&m[888]&~m[889]&m[891]&m[892])|(~m[837]&~m[888]&m[889]&m[891]&m[892])|(m[837]&~m[888]&m[889]&m[891]&m[892])|(m[837]&m[888]&m[889]&m[891]&m[892]))):InitCond[575];
    m[895] = run?((((m[842]&~m[893]&~m[894]&~m[896]&~m[897])|(~m[842]&~m[893]&~m[894]&m[896]&~m[897])|(m[842]&m[893]&~m[894]&m[896]&~m[897])|(m[842]&~m[893]&m[894]&m[896]&~m[897])|(~m[842]&m[893]&~m[894]&~m[896]&m[897])|(~m[842]&~m[893]&m[894]&~m[896]&m[897])|(m[842]&m[893]&m[894]&~m[896]&m[897])|(~m[842]&m[893]&m[894]&m[896]&m[897]))&UnbiasedRNG[193])|((m[842]&~m[893]&~m[894]&m[896]&~m[897])|(~m[842]&~m[893]&~m[894]&~m[896]&m[897])|(m[842]&~m[893]&~m[894]&~m[896]&m[897])|(m[842]&m[893]&~m[894]&~m[896]&m[897])|(m[842]&~m[893]&m[894]&~m[896]&m[897])|(~m[842]&~m[893]&~m[894]&m[896]&m[897])|(m[842]&~m[893]&~m[894]&m[896]&m[897])|(~m[842]&m[893]&~m[894]&m[896]&m[897])|(m[842]&m[893]&~m[894]&m[896]&m[897])|(~m[842]&~m[893]&m[894]&m[896]&m[897])|(m[842]&~m[893]&m[894]&m[896]&m[897])|(m[842]&m[893]&m[894]&m[896]&m[897]))):InitCond[576];
    m[900] = run?((((m[847]&~m[898]&~m[899]&~m[901]&~m[902])|(~m[847]&~m[898]&~m[899]&m[901]&~m[902])|(m[847]&m[898]&~m[899]&m[901]&~m[902])|(m[847]&~m[898]&m[899]&m[901]&~m[902])|(~m[847]&m[898]&~m[899]&~m[901]&m[902])|(~m[847]&~m[898]&m[899]&~m[901]&m[902])|(m[847]&m[898]&m[899]&~m[901]&m[902])|(~m[847]&m[898]&m[899]&m[901]&m[902]))&UnbiasedRNG[194])|((m[847]&~m[898]&~m[899]&m[901]&~m[902])|(~m[847]&~m[898]&~m[899]&~m[901]&m[902])|(m[847]&~m[898]&~m[899]&~m[901]&m[902])|(m[847]&m[898]&~m[899]&~m[901]&m[902])|(m[847]&~m[898]&m[899]&~m[901]&m[902])|(~m[847]&~m[898]&~m[899]&m[901]&m[902])|(m[847]&~m[898]&~m[899]&m[901]&m[902])|(~m[847]&m[898]&~m[899]&m[901]&m[902])|(m[847]&m[898]&~m[899]&m[901]&m[902])|(~m[847]&~m[898]&m[899]&m[901]&m[902])|(m[847]&~m[898]&m[899]&m[901]&m[902])|(m[847]&m[898]&m[899]&m[901]&m[902]))):InitCond[577];
    m[905] = run?((((m[852]&~m[903]&~m[904]&~m[906]&~m[907])|(~m[852]&~m[903]&~m[904]&m[906]&~m[907])|(m[852]&m[903]&~m[904]&m[906]&~m[907])|(m[852]&~m[903]&m[904]&m[906]&~m[907])|(~m[852]&m[903]&~m[904]&~m[906]&m[907])|(~m[852]&~m[903]&m[904]&~m[906]&m[907])|(m[852]&m[903]&m[904]&~m[906]&m[907])|(~m[852]&m[903]&m[904]&m[906]&m[907]))&UnbiasedRNG[195])|((m[852]&~m[903]&~m[904]&m[906]&~m[907])|(~m[852]&~m[903]&~m[904]&~m[906]&m[907])|(m[852]&~m[903]&~m[904]&~m[906]&m[907])|(m[852]&m[903]&~m[904]&~m[906]&m[907])|(m[852]&~m[903]&m[904]&~m[906]&m[907])|(~m[852]&~m[903]&~m[904]&m[906]&m[907])|(m[852]&~m[903]&~m[904]&m[906]&m[907])|(~m[852]&m[903]&~m[904]&m[906]&m[907])|(m[852]&m[903]&~m[904]&m[906]&m[907])|(~m[852]&~m[903]&m[904]&m[906]&m[907])|(m[852]&~m[903]&m[904]&m[906]&m[907])|(m[852]&m[903]&m[904]&m[906]&m[907]))):InitCond[578];
    m[910] = run?((((m[857]&~m[908]&~m[909]&~m[911]&~m[912])|(~m[857]&~m[908]&~m[909]&m[911]&~m[912])|(m[857]&m[908]&~m[909]&m[911]&~m[912])|(m[857]&~m[908]&m[909]&m[911]&~m[912])|(~m[857]&m[908]&~m[909]&~m[911]&m[912])|(~m[857]&~m[908]&m[909]&~m[911]&m[912])|(m[857]&m[908]&m[909]&~m[911]&m[912])|(~m[857]&m[908]&m[909]&m[911]&m[912]))&UnbiasedRNG[196])|((m[857]&~m[908]&~m[909]&m[911]&~m[912])|(~m[857]&~m[908]&~m[909]&~m[911]&m[912])|(m[857]&~m[908]&~m[909]&~m[911]&m[912])|(m[857]&m[908]&~m[909]&~m[911]&m[912])|(m[857]&~m[908]&m[909]&~m[911]&m[912])|(~m[857]&~m[908]&~m[909]&m[911]&m[912])|(m[857]&~m[908]&~m[909]&m[911]&m[912])|(~m[857]&m[908]&~m[909]&m[911]&m[912])|(m[857]&m[908]&~m[909]&m[911]&m[912])|(~m[857]&~m[908]&m[909]&m[911]&m[912])|(m[857]&~m[908]&m[909]&m[911]&m[912])|(m[857]&m[908]&m[909]&m[911]&m[912]))):InitCond[579];
    m[915] = run?((((m[867]&~m[913]&~m[914]&~m[916]&~m[917])|(~m[867]&~m[913]&~m[914]&m[916]&~m[917])|(m[867]&m[913]&~m[914]&m[916]&~m[917])|(m[867]&~m[913]&m[914]&m[916]&~m[917])|(~m[867]&m[913]&~m[914]&~m[916]&m[917])|(~m[867]&~m[913]&m[914]&~m[916]&m[917])|(m[867]&m[913]&m[914]&~m[916]&m[917])|(~m[867]&m[913]&m[914]&m[916]&m[917]))&UnbiasedRNG[197])|((m[867]&~m[913]&~m[914]&m[916]&~m[917])|(~m[867]&~m[913]&~m[914]&~m[916]&m[917])|(m[867]&~m[913]&~m[914]&~m[916]&m[917])|(m[867]&m[913]&~m[914]&~m[916]&m[917])|(m[867]&~m[913]&m[914]&~m[916]&m[917])|(~m[867]&~m[913]&~m[914]&m[916]&m[917])|(m[867]&~m[913]&~m[914]&m[916]&m[917])|(~m[867]&m[913]&~m[914]&m[916]&m[917])|(m[867]&m[913]&~m[914]&m[916]&m[917])|(~m[867]&~m[913]&m[914]&m[916]&m[917])|(m[867]&~m[913]&m[914]&m[916]&m[917])|(m[867]&m[913]&m[914]&m[916]&m[917]))):InitCond[580];
    m[920] = run?((((m[872]&~m[918]&~m[919]&~m[921]&~m[922])|(~m[872]&~m[918]&~m[919]&m[921]&~m[922])|(m[872]&m[918]&~m[919]&m[921]&~m[922])|(m[872]&~m[918]&m[919]&m[921]&~m[922])|(~m[872]&m[918]&~m[919]&~m[921]&m[922])|(~m[872]&~m[918]&m[919]&~m[921]&m[922])|(m[872]&m[918]&m[919]&~m[921]&m[922])|(~m[872]&m[918]&m[919]&m[921]&m[922]))&UnbiasedRNG[198])|((m[872]&~m[918]&~m[919]&m[921]&~m[922])|(~m[872]&~m[918]&~m[919]&~m[921]&m[922])|(m[872]&~m[918]&~m[919]&~m[921]&m[922])|(m[872]&m[918]&~m[919]&~m[921]&m[922])|(m[872]&~m[918]&m[919]&~m[921]&m[922])|(~m[872]&~m[918]&~m[919]&m[921]&m[922])|(m[872]&~m[918]&~m[919]&m[921]&m[922])|(~m[872]&m[918]&~m[919]&m[921]&m[922])|(m[872]&m[918]&~m[919]&m[921]&m[922])|(~m[872]&~m[918]&m[919]&m[921]&m[922])|(m[872]&~m[918]&m[919]&m[921]&m[922])|(m[872]&m[918]&m[919]&m[921]&m[922]))):InitCond[581];
    m[925] = run?((((m[877]&~m[923]&~m[924]&~m[926]&~m[927])|(~m[877]&~m[923]&~m[924]&m[926]&~m[927])|(m[877]&m[923]&~m[924]&m[926]&~m[927])|(m[877]&~m[923]&m[924]&m[926]&~m[927])|(~m[877]&m[923]&~m[924]&~m[926]&m[927])|(~m[877]&~m[923]&m[924]&~m[926]&m[927])|(m[877]&m[923]&m[924]&~m[926]&m[927])|(~m[877]&m[923]&m[924]&m[926]&m[927]))&UnbiasedRNG[199])|((m[877]&~m[923]&~m[924]&m[926]&~m[927])|(~m[877]&~m[923]&~m[924]&~m[926]&m[927])|(m[877]&~m[923]&~m[924]&~m[926]&m[927])|(m[877]&m[923]&~m[924]&~m[926]&m[927])|(m[877]&~m[923]&m[924]&~m[926]&m[927])|(~m[877]&~m[923]&~m[924]&m[926]&m[927])|(m[877]&~m[923]&~m[924]&m[926]&m[927])|(~m[877]&m[923]&~m[924]&m[926]&m[927])|(m[877]&m[923]&~m[924]&m[926]&m[927])|(~m[877]&~m[923]&m[924]&m[926]&m[927])|(m[877]&~m[923]&m[924]&m[926]&m[927])|(m[877]&m[923]&m[924]&m[926]&m[927]))):InitCond[582];
    m[930] = run?((((m[882]&~m[928]&~m[929]&~m[931]&~m[932])|(~m[882]&~m[928]&~m[929]&m[931]&~m[932])|(m[882]&m[928]&~m[929]&m[931]&~m[932])|(m[882]&~m[928]&m[929]&m[931]&~m[932])|(~m[882]&m[928]&~m[929]&~m[931]&m[932])|(~m[882]&~m[928]&m[929]&~m[931]&m[932])|(m[882]&m[928]&m[929]&~m[931]&m[932])|(~m[882]&m[928]&m[929]&m[931]&m[932]))&UnbiasedRNG[200])|((m[882]&~m[928]&~m[929]&m[931]&~m[932])|(~m[882]&~m[928]&~m[929]&~m[931]&m[932])|(m[882]&~m[928]&~m[929]&~m[931]&m[932])|(m[882]&m[928]&~m[929]&~m[931]&m[932])|(m[882]&~m[928]&m[929]&~m[931]&m[932])|(~m[882]&~m[928]&~m[929]&m[931]&m[932])|(m[882]&~m[928]&~m[929]&m[931]&m[932])|(~m[882]&m[928]&~m[929]&m[931]&m[932])|(m[882]&m[928]&~m[929]&m[931]&m[932])|(~m[882]&~m[928]&m[929]&m[931]&m[932])|(m[882]&~m[928]&m[929]&m[931]&m[932])|(m[882]&m[928]&m[929]&m[931]&m[932]))):InitCond[583];
    m[935] = run?((((m[887]&~m[933]&~m[934]&~m[936]&~m[937])|(~m[887]&~m[933]&~m[934]&m[936]&~m[937])|(m[887]&m[933]&~m[934]&m[936]&~m[937])|(m[887]&~m[933]&m[934]&m[936]&~m[937])|(~m[887]&m[933]&~m[934]&~m[936]&m[937])|(~m[887]&~m[933]&m[934]&~m[936]&m[937])|(m[887]&m[933]&m[934]&~m[936]&m[937])|(~m[887]&m[933]&m[934]&m[936]&m[937]))&UnbiasedRNG[201])|((m[887]&~m[933]&~m[934]&m[936]&~m[937])|(~m[887]&~m[933]&~m[934]&~m[936]&m[937])|(m[887]&~m[933]&~m[934]&~m[936]&m[937])|(m[887]&m[933]&~m[934]&~m[936]&m[937])|(m[887]&~m[933]&m[934]&~m[936]&m[937])|(~m[887]&~m[933]&~m[934]&m[936]&m[937])|(m[887]&~m[933]&~m[934]&m[936]&m[937])|(~m[887]&m[933]&~m[934]&m[936]&m[937])|(m[887]&m[933]&~m[934]&m[936]&m[937])|(~m[887]&~m[933]&m[934]&m[936]&m[937])|(m[887]&~m[933]&m[934]&m[936]&m[937])|(m[887]&m[933]&m[934]&m[936]&m[937]))):InitCond[584];
    m[940] = run?((((m[892]&~m[938]&~m[939]&~m[941]&~m[942])|(~m[892]&~m[938]&~m[939]&m[941]&~m[942])|(m[892]&m[938]&~m[939]&m[941]&~m[942])|(m[892]&~m[938]&m[939]&m[941]&~m[942])|(~m[892]&m[938]&~m[939]&~m[941]&m[942])|(~m[892]&~m[938]&m[939]&~m[941]&m[942])|(m[892]&m[938]&m[939]&~m[941]&m[942])|(~m[892]&m[938]&m[939]&m[941]&m[942]))&UnbiasedRNG[202])|((m[892]&~m[938]&~m[939]&m[941]&~m[942])|(~m[892]&~m[938]&~m[939]&~m[941]&m[942])|(m[892]&~m[938]&~m[939]&~m[941]&m[942])|(m[892]&m[938]&~m[939]&~m[941]&m[942])|(m[892]&~m[938]&m[939]&~m[941]&m[942])|(~m[892]&~m[938]&~m[939]&m[941]&m[942])|(m[892]&~m[938]&~m[939]&m[941]&m[942])|(~m[892]&m[938]&~m[939]&m[941]&m[942])|(m[892]&m[938]&~m[939]&m[941]&m[942])|(~m[892]&~m[938]&m[939]&m[941]&m[942])|(m[892]&~m[938]&m[939]&m[941]&m[942])|(m[892]&m[938]&m[939]&m[941]&m[942]))):InitCond[585];
    m[945] = run?((((m[897]&~m[943]&~m[944]&~m[946]&~m[947])|(~m[897]&~m[943]&~m[944]&m[946]&~m[947])|(m[897]&m[943]&~m[944]&m[946]&~m[947])|(m[897]&~m[943]&m[944]&m[946]&~m[947])|(~m[897]&m[943]&~m[944]&~m[946]&m[947])|(~m[897]&~m[943]&m[944]&~m[946]&m[947])|(m[897]&m[943]&m[944]&~m[946]&m[947])|(~m[897]&m[943]&m[944]&m[946]&m[947]))&UnbiasedRNG[203])|((m[897]&~m[943]&~m[944]&m[946]&~m[947])|(~m[897]&~m[943]&~m[944]&~m[946]&m[947])|(m[897]&~m[943]&~m[944]&~m[946]&m[947])|(m[897]&m[943]&~m[944]&~m[946]&m[947])|(m[897]&~m[943]&m[944]&~m[946]&m[947])|(~m[897]&~m[943]&~m[944]&m[946]&m[947])|(m[897]&~m[943]&~m[944]&m[946]&m[947])|(~m[897]&m[943]&~m[944]&m[946]&m[947])|(m[897]&m[943]&~m[944]&m[946]&m[947])|(~m[897]&~m[943]&m[944]&m[946]&m[947])|(m[897]&~m[943]&m[944]&m[946]&m[947])|(m[897]&m[943]&m[944]&m[946]&m[947]))):InitCond[586];
    m[950] = run?((((m[902]&~m[948]&~m[949]&~m[951]&~m[952])|(~m[902]&~m[948]&~m[949]&m[951]&~m[952])|(m[902]&m[948]&~m[949]&m[951]&~m[952])|(m[902]&~m[948]&m[949]&m[951]&~m[952])|(~m[902]&m[948]&~m[949]&~m[951]&m[952])|(~m[902]&~m[948]&m[949]&~m[951]&m[952])|(m[902]&m[948]&m[949]&~m[951]&m[952])|(~m[902]&m[948]&m[949]&m[951]&m[952]))&UnbiasedRNG[204])|((m[902]&~m[948]&~m[949]&m[951]&~m[952])|(~m[902]&~m[948]&~m[949]&~m[951]&m[952])|(m[902]&~m[948]&~m[949]&~m[951]&m[952])|(m[902]&m[948]&~m[949]&~m[951]&m[952])|(m[902]&~m[948]&m[949]&~m[951]&m[952])|(~m[902]&~m[948]&~m[949]&m[951]&m[952])|(m[902]&~m[948]&~m[949]&m[951]&m[952])|(~m[902]&m[948]&~m[949]&m[951]&m[952])|(m[902]&m[948]&~m[949]&m[951]&m[952])|(~m[902]&~m[948]&m[949]&m[951]&m[952])|(m[902]&~m[948]&m[949]&m[951]&m[952])|(m[902]&m[948]&m[949]&m[951]&m[952]))):InitCond[587];
    m[955] = run?((((m[907]&~m[953]&~m[954]&~m[956]&~m[957])|(~m[907]&~m[953]&~m[954]&m[956]&~m[957])|(m[907]&m[953]&~m[954]&m[956]&~m[957])|(m[907]&~m[953]&m[954]&m[956]&~m[957])|(~m[907]&m[953]&~m[954]&~m[956]&m[957])|(~m[907]&~m[953]&m[954]&~m[956]&m[957])|(m[907]&m[953]&m[954]&~m[956]&m[957])|(~m[907]&m[953]&m[954]&m[956]&m[957]))&UnbiasedRNG[205])|((m[907]&~m[953]&~m[954]&m[956]&~m[957])|(~m[907]&~m[953]&~m[954]&~m[956]&m[957])|(m[907]&~m[953]&~m[954]&~m[956]&m[957])|(m[907]&m[953]&~m[954]&~m[956]&m[957])|(m[907]&~m[953]&m[954]&~m[956]&m[957])|(~m[907]&~m[953]&~m[954]&m[956]&m[957])|(m[907]&~m[953]&~m[954]&m[956]&m[957])|(~m[907]&m[953]&~m[954]&m[956]&m[957])|(m[907]&m[953]&~m[954]&m[956]&m[957])|(~m[907]&~m[953]&m[954]&m[956]&m[957])|(m[907]&~m[953]&m[954]&m[956]&m[957])|(m[907]&m[953]&m[954]&m[956]&m[957]))):InitCond[588];
    m[960] = run?((((m[912]&~m[958]&~m[959]&~m[961]&~m[962])|(~m[912]&~m[958]&~m[959]&m[961]&~m[962])|(m[912]&m[958]&~m[959]&m[961]&~m[962])|(m[912]&~m[958]&m[959]&m[961]&~m[962])|(~m[912]&m[958]&~m[959]&~m[961]&m[962])|(~m[912]&~m[958]&m[959]&~m[961]&m[962])|(m[912]&m[958]&m[959]&~m[961]&m[962])|(~m[912]&m[958]&m[959]&m[961]&m[962]))&UnbiasedRNG[206])|((m[912]&~m[958]&~m[959]&m[961]&~m[962])|(~m[912]&~m[958]&~m[959]&~m[961]&m[962])|(m[912]&~m[958]&~m[959]&~m[961]&m[962])|(m[912]&m[958]&~m[959]&~m[961]&m[962])|(m[912]&~m[958]&m[959]&~m[961]&m[962])|(~m[912]&~m[958]&~m[959]&m[961]&m[962])|(m[912]&~m[958]&~m[959]&m[961]&m[962])|(~m[912]&m[958]&~m[959]&m[961]&m[962])|(m[912]&m[958]&~m[959]&m[961]&m[962])|(~m[912]&~m[958]&m[959]&m[961]&m[962])|(m[912]&~m[958]&m[959]&m[961]&m[962])|(m[912]&m[958]&m[959]&m[961]&m[962]))):InitCond[589];
    m[965] = run?((((m[922]&~m[963]&~m[964]&~m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&m[966]&~m[967])|(m[922]&m[963]&~m[964]&m[966]&~m[967])|(m[922]&~m[963]&m[964]&m[966]&~m[967])|(~m[922]&m[963]&~m[964]&~m[966]&m[967])|(~m[922]&~m[963]&m[964]&~m[966]&m[967])|(m[922]&m[963]&m[964]&~m[966]&m[967])|(~m[922]&m[963]&m[964]&m[966]&m[967]))&UnbiasedRNG[207])|((m[922]&~m[963]&~m[964]&m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&m[964]&~m[966]&m[967])|(~m[922]&~m[963]&~m[964]&m[966]&m[967])|(m[922]&~m[963]&~m[964]&m[966]&m[967])|(~m[922]&m[963]&~m[964]&m[966]&m[967])|(m[922]&m[963]&~m[964]&m[966]&m[967])|(~m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&m[963]&m[964]&m[966]&m[967]))):InitCond[590];
    m[970] = run?((((m[927]&~m[968]&~m[969]&~m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&m[971]&~m[972])|(m[927]&m[968]&~m[969]&m[971]&~m[972])|(m[927]&~m[968]&m[969]&m[971]&~m[972])|(~m[927]&m[968]&~m[969]&~m[971]&m[972])|(~m[927]&~m[968]&m[969]&~m[971]&m[972])|(m[927]&m[968]&m[969]&~m[971]&m[972])|(~m[927]&m[968]&m[969]&m[971]&m[972]))&UnbiasedRNG[208])|((m[927]&~m[968]&~m[969]&m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&m[969]&~m[971]&m[972])|(~m[927]&~m[968]&~m[969]&m[971]&m[972])|(m[927]&~m[968]&~m[969]&m[971]&m[972])|(~m[927]&m[968]&~m[969]&m[971]&m[972])|(m[927]&m[968]&~m[969]&m[971]&m[972])|(~m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&m[968]&m[969]&m[971]&m[972]))):InitCond[591];
    m[975] = run?((((m[932]&~m[973]&~m[974]&~m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&m[976]&~m[977])|(m[932]&m[973]&~m[974]&m[976]&~m[977])|(m[932]&~m[973]&m[974]&m[976]&~m[977])|(~m[932]&m[973]&~m[974]&~m[976]&m[977])|(~m[932]&~m[973]&m[974]&~m[976]&m[977])|(m[932]&m[973]&m[974]&~m[976]&m[977])|(~m[932]&m[973]&m[974]&m[976]&m[977]))&UnbiasedRNG[209])|((m[932]&~m[973]&~m[974]&m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&m[974]&~m[976]&m[977])|(~m[932]&~m[973]&~m[974]&m[976]&m[977])|(m[932]&~m[973]&~m[974]&m[976]&m[977])|(~m[932]&m[973]&~m[974]&m[976]&m[977])|(m[932]&m[973]&~m[974]&m[976]&m[977])|(~m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&m[973]&m[974]&m[976]&m[977]))):InitCond[592];
    m[980] = run?((((m[937]&~m[978]&~m[979]&~m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&m[981]&~m[982])|(m[937]&m[978]&~m[979]&m[981]&~m[982])|(m[937]&~m[978]&m[979]&m[981]&~m[982])|(~m[937]&m[978]&~m[979]&~m[981]&m[982])|(~m[937]&~m[978]&m[979]&~m[981]&m[982])|(m[937]&m[978]&m[979]&~m[981]&m[982])|(~m[937]&m[978]&m[979]&m[981]&m[982]))&UnbiasedRNG[210])|((m[937]&~m[978]&~m[979]&m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&m[979]&~m[981]&m[982])|(~m[937]&~m[978]&~m[979]&m[981]&m[982])|(m[937]&~m[978]&~m[979]&m[981]&m[982])|(~m[937]&m[978]&~m[979]&m[981]&m[982])|(m[937]&m[978]&~m[979]&m[981]&m[982])|(~m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&m[978]&m[979]&m[981]&m[982]))):InitCond[593];
    m[985] = run?((((m[942]&~m[983]&~m[984]&~m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&m[986]&~m[987])|(m[942]&m[983]&~m[984]&m[986]&~m[987])|(m[942]&~m[983]&m[984]&m[986]&~m[987])|(~m[942]&m[983]&~m[984]&~m[986]&m[987])|(~m[942]&~m[983]&m[984]&~m[986]&m[987])|(m[942]&m[983]&m[984]&~m[986]&m[987])|(~m[942]&m[983]&m[984]&m[986]&m[987]))&UnbiasedRNG[211])|((m[942]&~m[983]&~m[984]&m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&m[984]&~m[986]&m[987])|(~m[942]&~m[983]&~m[984]&m[986]&m[987])|(m[942]&~m[983]&~m[984]&m[986]&m[987])|(~m[942]&m[983]&~m[984]&m[986]&m[987])|(m[942]&m[983]&~m[984]&m[986]&m[987])|(~m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&m[983]&m[984]&m[986]&m[987]))):InitCond[594];
    m[990] = run?((((m[947]&~m[988]&~m[989]&~m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&m[991]&~m[992])|(m[947]&m[988]&~m[989]&m[991]&~m[992])|(m[947]&~m[988]&m[989]&m[991]&~m[992])|(~m[947]&m[988]&~m[989]&~m[991]&m[992])|(~m[947]&~m[988]&m[989]&~m[991]&m[992])|(m[947]&m[988]&m[989]&~m[991]&m[992])|(~m[947]&m[988]&m[989]&m[991]&m[992]))&UnbiasedRNG[212])|((m[947]&~m[988]&~m[989]&m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&m[989]&~m[991]&m[992])|(~m[947]&~m[988]&~m[989]&m[991]&m[992])|(m[947]&~m[988]&~m[989]&m[991]&m[992])|(~m[947]&m[988]&~m[989]&m[991]&m[992])|(m[947]&m[988]&~m[989]&m[991]&m[992])|(~m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&m[988]&m[989]&m[991]&m[992]))):InitCond[595];
    m[995] = run?((((m[952]&~m[993]&~m[994]&~m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&m[996]&~m[997])|(m[952]&m[993]&~m[994]&m[996]&~m[997])|(m[952]&~m[993]&m[994]&m[996]&~m[997])|(~m[952]&m[993]&~m[994]&~m[996]&m[997])|(~m[952]&~m[993]&m[994]&~m[996]&m[997])|(m[952]&m[993]&m[994]&~m[996]&m[997])|(~m[952]&m[993]&m[994]&m[996]&m[997]))&UnbiasedRNG[213])|((m[952]&~m[993]&~m[994]&m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&m[994]&~m[996]&m[997])|(~m[952]&~m[993]&~m[994]&m[996]&m[997])|(m[952]&~m[993]&~m[994]&m[996]&m[997])|(~m[952]&m[993]&~m[994]&m[996]&m[997])|(m[952]&m[993]&~m[994]&m[996]&m[997])|(~m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&m[993]&m[994]&m[996]&m[997]))):InitCond[596];
    m[1000] = run?((((m[957]&~m[998]&~m[999]&~m[1001]&~m[1002])|(~m[957]&~m[998]&~m[999]&m[1001]&~m[1002])|(m[957]&m[998]&~m[999]&m[1001]&~m[1002])|(m[957]&~m[998]&m[999]&m[1001]&~m[1002])|(~m[957]&m[998]&~m[999]&~m[1001]&m[1002])|(~m[957]&~m[998]&m[999]&~m[1001]&m[1002])|(m[957]&m[998]&m[999]&~m[1001]&m[1002])|(~m[957]&m[998]&m[999]&m[1001]&m[1002]))&UnbiasedRNG[214])|((m[957]&~m[998]&~m[999]&m[1001]&~m[1002])|(~m[957]&~m[998]&~m[999]&~m[1001]&m[1002])|(m[957]&~m[998]&~m[999]&~m[1001]&m[1002])|(m[957]&m[998]&~m[999]&~m[1001]&m[1002])|(m[957]&~m[998]&m[999]&~m[1001]&m[1002])|(~m[957]&~m[998]&~m[999]&m[1001]&m[1002])|(m[957]&~m[998]&~m[999]&m[1001]&m[1002])|(~m[957]&m[998]&~m[999]&m[1001]&m[1002])|(m[957]&m[998]&~m[999]&m[1001]&m[1002])|(~m[957]&~m[998]&m[999]&m[1001]&m[1002])|(m[957]&~m[998]&m[999]&m[1001]&m[1002])|(m[957]&m[998]&m[999]&m[1001]&m[1002]))):InitCond[597];
    m[1005] = run?((((m[962]&~m[1003]&~m[1004]&~m[1006]&~m[1007])|(~m[962]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(m[962]&m[1003]&~m[1004]&m[1006]&~m[1007])|(m[962]&~m[1003]&m[1004]&m[1006]&~m[1007])|(~m[962]&m[1003]&~m[1004]&~m[1006]&m[1007])|(~m[962]&~m[1003]&m[1004]&~m[1006]&m[1007])|(m[962]&m[1003]&m[1004]&~m[1006]&m[1007])|(~m[962]&m[1003]&m[1004]&m[1006]&m[1007]))&UnbiasedRNG[215])|((m[962]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(~m[962]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[962]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[962]&m[1003]&~m[1004]&~m[1006]&m[1007])|(m[962]&~m[1003]&m[1004]&~m[1006]&m[1007])|(~m[962]&~m[1003]&~m[1004]&m[1006]&m[1007])|(m[962]&~m[1003]&~m[1004]&m[1006]&m[1007])|(~m[962]&m[1003]&~m[1004]&m[1006]&m[1007])|(m[962]&m[1003]&~m[1004]&m[1006]&m[1007])|(~m[962]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[962]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[962]&m[1003]&m[1004]&m[1006]&m[1007]))):InitCond[598];
    m[1010] = run?((((m[972]&~m[1008]&~m[1009]&~m[1011]&~m[1012])|(~m[972]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(m[972]&m[1008]&~m[1009]&m[1011]&~m[1012])|(m[972]&~m[1008]&m[1009]&m[1011]&~m[1012])|(~m[972]&m[1008]&~m[1009]&~m[1011]&m[1012])|(~m[972]&~m[1008]&m[1009]&~m[1011]&m[1012])|(m[972]&m[1008]&m[1009]&~m[1011]&m[1012])|(~m[972]&m[1008]&m[1009]&m[1011]&m[1012]))&UnbiasedRNG[216])|((m[972]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(~m[972]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[972]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[972]&m[1008]&~m[1009]&~m[1011]&m[1012])|(m[972]&~m[1008]&m[1009]&~m[1011]&m[1012])|(~m[972]&~m[1008]&~m[1009]&m[1011]&m[1012])|(m[972]&~m[1008]&~m[1009]&m[1011]&m[1012])|(~m[972]&m[1008]&~m[1009]&m[1011]&m[1012])|(m[972]&m[1008]&~m[1009]&m[1011]&m[1012])|(~m[972]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[972]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[972]&m[1008]&m[1009]&m[1011]&m[1012]))):InitCond[599];
    m[1015] = run?((((m[977]&~m[1013]&~m[1014]&~m[1016]&~m[1017])|(~m[977]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(m[977]&m[1013]&~m[1014]&m[1016]&~m[1017])|(m[977]&~m[1013]&m[1014]&m[1016]&~m[1017])|(~m[977]&m[1013]&~m[1014]&~m[1016]&m[1017])|(~m[977]&~m[1013]&m[1014]&~m[1016]&m[1017])|(m[977]&m[1013]&m[1014]&~m[1016]&m[1017])|(~m[977]&m[1013]&m[1014]&m[1016]&m[1017]))&UnbiasedRNG[217])|((m[977]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(~m[977]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[977]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[977]&m[1013]&~m[1014]&~m[1016]&m[1017])|(m[977]&~m[1013]&m[1014]&~m[1016]&m[1017])|(~m[977]&~m[1013]&~m[1014]&m[1016]&m[1017])|(m[977]&~m[1013]&~m[1014]&m[1016]&m[1017])|(~m[977]&m[1013]&~m[1014]&m[1016]&m[1017])|(m[977]&m[1013]&~m[1014]&m[1016]&m[1017])|(~m[977]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[977]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[977]&m[1013]&m[1014]&m[1016]&m[1017]))):InitCond[600];
    m[1020] = run?((((m[982]&~m[1018]&~m[1019]&~m[1021]&~m[1022])|(~m[982]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(m[982]&m[1018]&~m[1019]&m[1021]&~m[1022])|(m[982]&~m[1018]&m[1019]&m[1021]&~m[1022])|(~m[982]&m[1018]&~m[1019]&~m[1021]&m[1022])|(~m[982]&~m[1018]&m[1019]&~m[1021]&m[1022])|(m[982]&m[1018]&m[1019]&~m[1021]&m[1022])|(~m[982]&m[1018]&m[1019]&m[1021]&m[1022]))&UnbiasedRNG[218])|((m[982]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(~m[982]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[982]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[982]&m[1018]&~m[1019]&~m[1021]&m[1022])|(m[982]&~m[1018]&m[1019]&~m[1021]&m[1022])|(~m[982]&~m[1018]&~m[1019]&m[1021]&m[1022])|(m[982]&~m[1018]&~m[1019]&m[1021]&m[1022])|(~m[982]&m[1018]&~m[1019]&m[1021]&m[1022])|(m[982]&m[1018]&~m[1019]&m[1021]&m[1022])|(~m[982]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[982]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[982]&m[1018]&m[1019]&m[1021]&m[1022]))):InitCond[601];
    m[1025] = run?((((m[987]&~m[1023]&~m[1024]&~m[1026]&~m[1027])|(~m[987]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(m[987]&m[1023]&~m[1024]&m[1026]&~m[1027])|(m[987]&~m[1023]&m[1024]&m[1026]&~m[1027])|(~m[987]&m[1023]&~m[1024]&~m[1026]&m[1027])|(~m[987]&~m[1023]&m[1024]&~m[1026]&m[1027])|(m[987]&m[1023]&m[1024]&~m[1026]&m[1027])|(~m[987]&m[1023]&m[1024]&m[1026]&m[1027]))&UnbiasedRNG[219])|((m[987]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(~m[987]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[987]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[987]&m[1023]&~m[1024]&~m[1026]&m[1027])|(m[987]&~m[1023]&m[1024]&~m[1026]&m[1027])|(~m[987]&~m[1023]&~m[1024]&m[1026]&m[1027])|(m[987]&~m[1023]&~m[1024]&m[1026]&m[1027])|(~m[987]&m[1023]&~m[1024]&m[1026]&m[1027])|(m[987]&m[1023]&~m[1024]&m[1026]&m[1027])|(~m[987]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[987]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[987]&m[1023]&m[1024]&m[1026]&m[1027]))):InitCond[602];
    m[1030] = run?((((m[992]&~m[1028]&~m[1029]&~m[1031]&~m[1032])|(~m[992]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(m[992]&m[1028]&~m[1029]&m[1031]&~m[1032])|(m[992]&~m[1028]&m[1029]&m[1031]&~m[1032])|(~m[992]&m[1028]&~m[1029]&~m[1031]&m[1032])|(~m[992]&~m[1028]&m[1029]&~m[1031]&m[1032])|(m[992]&m[1028]&m[1029]&~m[1031]&m[1032])|(~m[992]&m[1028]&m[1029]&m[1031]&m[1032]))&UnbiasedRNG[220])|((m[992]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(~m[992]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[992]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[992]&m[1028]&~m[1029]&~m[1031]&m[1032])|(m[992]&~m[1028]&m[1029]&~m[1031]&m[1032])|(~m[992]&~m[1028]&~m[1029]&m[1031]&m[1032])|(m[992]&~m[1028]&~m[1029]&m[1031]&m[1032])|(~m[992]&m[1028]&~m[1029]&m[1031]&m[1032])|(m[992]&m[1028]&~m[1029]&m[1031]&m[1032])|(~m[992]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[992]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[992]&m[1028]&m[1029]&m[1031]&m[1032]))):InitCond[603];
    m[1035] = run?((((m[997]&~m[1033]&~m[1034]&~m[1036]&~m[1037])|(~m[997]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(m[997]&m[1033]&~m[1034]&m[1036]&~m[1037])|(m[997]&~m[1033]&m[1034]&m[1036]&~m[1037])|(~m[997]&m[1033]&~m[1034]&~m[1036]&m[1037])|(~m[997]&~m[1033]&m[1034]&~m[1036]&m[1037])|(m[997]&m[1033]&m[1034]&~m[1036]&m[1037])|(~m[997]&m[1033]&m[1034]&m[1036]&m[1037]))&UnbiasedRNG[221])|((m[997]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(~m[997]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[997]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[997]&m[1033]&~m[1034]&~m[1036]&m[1037])|(m[997]&~m[1033]&m[1034]&~m[1036]&m[1037])|(~m[997]&~m[1033]&~m[1034]&m[1036]&m[1037])|(m[997]&~m[1033]&~m[1034]&m[1036]&m[1037])|(~m[997]&m[1033]&~m[1034]&m[1036]&m[1037])|(m[997]&m[1033]&~m[1034]&m[1036]&m[1037])|(~m[997]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[997]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[997]&m[1033]&m[1034]&m[1036]&m[1037]))):InitCond[604];
    m[1040] = run?((((m[1002]&~m[1038]&~m[1039]&~m[1041]&~m[1042])|(~m[1002]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1002]&m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1002]&~m[1038]&m[1039]&m[1041]&~m[1042])|(~m[1002]&m[1038]&~m[1039]&~m[1041]&m[1042])|(~m[1002]&~m[1038]&m[1039]&~m[1041]&m[1042])|(m[1002]&m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1002]&m[1038]&m[1039]&m[1041]&m[1042]))&UnbiasedRNG[222])|((m[1002]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(~m[1002]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1002]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1002]&m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1002]&~m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1002]&~m[1038]&~m[1039]&m[1041]&m[1042])|(m[1002]&~m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1002]&m[1038]&~m[1039]&m[1041]&m[1042])|(m[1002]&m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1002]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1002]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1002]&m[1038]&m[1039]&m[1041]&m[1042]))):InitCond[605];
    m[1045] = run?((((m[1007]&~m[1043]&~m[1044]&~m[1046]&~m[1047])|(~m[1007]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1007]&m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1007]&~m[1043]&m[1044]&m[1046]&~m[1047])|(~m[1007]&m[1043]&~m[1044]&~m[1046]&m[1047])|(~m[1007]&~m[1043]&m[1044]&~m[1046]&m[1047])|(m[1007]&m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1007]&m[1043]&m[1044]&m[1046]&m[1047]))&UnbiasedRNG[223])|((m[1007]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(~m[1007]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1007]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1007]&m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1007]&~m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1007]&~m[1043]&~m[1044]&m[1046]&m[1047])|(m[1007]&~m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1007]&m[1043]&~m[1044]&m[1046]&m[1047])|(m[1007]&m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1007]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1007]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1007]&m[1043]&m[1044]&m[1046]&m[1047]))):InitCond[606];
    m[1050] = run?((((m[1017]&~m[1048]&~m[1049]&~m[1051]&~m[1052])|(~m[1017]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1017]&m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1017]&~m[1048]&m[1049]&m[1051]&~m[1052])|(~m[1017]&m[1048]&~m[1049]&~m[1051]&m[1052])|(~m[1017]&~m[1048]&m[1049]&~m[1051]&m[1052])|(m[1017]&m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1017]&m[1048]&m[1049]&m[1051]&m[1052]))&UnbiasedRNG[224])|((m[1017]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(~m[1017]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1017]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1017]&m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1017]&~m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1017]&~m[1048]&~m[1049]&m[1051]&m[1052])|(m[1017]&~m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1017]&m[1048]&~m[1049]&m[1051]&m[1052])|(m[1017]&m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1017]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1017]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1017]&m[1048]&m[1049]&m[1051]&m[1052]))):InitCond[607];
    m[1055] = run?((((m[1022]&~m[1053]&~m[1054]&~m[1056]&~m[1057])|(~m[1022]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1022]&m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1022]&~m[1053]&m[1054]&m[1056]&~m[1057])|(~m[1022]&m[1053]&~m[1054]&~m[1056]&m[1057])|(~m[1022]&~m[1053]&m[1054]&~m[1056]&m[1057])|(m[1022]&m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1022]&m[1053]&m[1054]&m[1056]&m[1057]))&UnbiasedRNG[225])|((m[1022]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(~m[1022]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1022]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1022]&m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1022]&~m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1022]&~m[1053]&~m[1054]&m[1056]&m[1057])|(m[1022]&~m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1022]&m[1053]&~m[1054]&m[1056]&m[1057])|(m[1022]&m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1022]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1022]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1022]&m[1053]&m[1054]&m[1056]&m[1057]))):InitCond[608];
    m[1060] = run?((((m[1027]&~m[1058]&~m[1059]&~m[1061]&~m[1062])|(~m[1027]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1027]&m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1027]&~m[1058]&m[1059]&m[1061]&~m[1062])|(~m[1027]&m[1058]&~m[1059]&~m[1061]&m[1062])|(~m[1027]&~m[1058]&m[1059]&~m[1061]&m[1062])|(m[1027]&m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1027]&m[1058]&m[1059]&m[1061]&m[1062]))&UnbiasedRNG[226])|((m[1027]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(~m[1027]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1027]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1027]&m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1027]&~m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1027]&~m[1058]&~m[1059]&m[1061]&m[1062])|(m[1027]&~m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1027]&m[1058]&~m[1059]&m[1061]&m[1062])|(m[1027]&m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1027]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1027]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1027]&m[1058]&m[1059]&m[1061]&m[1062]))):InitCond[609];
    m[1065] = run?((((m[1032]&~m[1063]&~m[1064]&~m[1066]&~m[1067])|(~m[1032]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1032]&m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1032]&~m[1063]&m[1064]&m[1066]&~m[1067])|(~m[1032]&m[1063]&~m[1064]&~m[1066]&m[1067])|(~m[1032]&~m[1063]&m[1064]&~m[1066]&m[1067])|(m[1032]&m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1032]&m[1063]&m[1064]&m[1066]&m[1067]))&UnbiasedRNG[227])|((m[1032]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(~m[1032]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1032]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1032]&m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1032]&~m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1032]&~m[1063]&~m[1064]&m[1066]&m[1067])|(m[1032]&~m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1032]&m[1063]&~m[1064]&m[1066]&m[1067])|(m[1032]&m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1032]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1032]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1032]&m[1063]&m[1064]&m[1066]&m[1067]))):InitCond[610];
    m[1070] = run?((((m[1037]&~m[1068]&~m[1069]&~m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&~m[1072])|(~m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&m[1068]&m[1069]&m[1071]&m[1072]))&UnbiasedRNG[228])|((m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&m[1071]&m[1072]))):InitCond[611];
    m[1075] = run?((((m[1042]&~m[1073]&~m[1074]&~m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&~m[1077])|(~m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&m[1073]&m[1074]&m[1076]&m[1077]))&UnbiasedRNG[229])|((m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&m[1076]&m[1077]))):InitCond[612];
    m[1080] = run?((((m[1047]&~m[1078]&~m[1079]&~m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&~m[1082])|(~m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&m[1078]&m[1079]&m[1081]&m[1082]))&UnbiasedRNG[230])|((m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&m[1081]&m[1082]))):InitCond[613];
    m[1085] = run?((((m[1057]&~m[1083]&~m[1084]&~m[1086]&~m[1087])|(~m[1057]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1057]&m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1057]&~m[1083]&m[1084]&m[1086]&~m[1087])|(~m[1057]&m[1083]&~m[1084]&~m[1086]&m[1087])|(~m[1057]&~m[1083]&m[1084]&~m[1086]&m[1087])|(m[1057]&m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1057]&m[1083]&m[1084]&m[1086]&m[1087]))&UnbiasedRNG[231])|((m[1057]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(~m[1057]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1057]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1057]&m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1057]&~m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1057]&~m[1083]&~m[1084]&m[1086]&m[1087])|(m[1057]&~m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1057]&m[1083]&~m[1084]&m[1086]&m[1087])|(m[1057]&m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1057]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1057]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1057]&m[1083]&m[1084]&m[1086]&m[1087]))):InitCond[614];
    m[1090] = run?((((m[1062]&~m[1088]&~m[1089]&~m[1091]&~m[1092])|(~m[1062]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1062]&m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1062]&~m[1088]&m[1089]&m[1091]&~m[1092])|(~m[1062]&m[1088]&~m[1089]&~m[1091]&m[1092])|(~m[1062]&~m[1088]&m[1089]&~m[1091]&m[1092])|(m[1062]&m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1062]&m[1088]&m[1089]&m[1091]&m[1092]))&UnbiasedRNG[232])|((m[1062]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(~m[1062]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1062]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1062]&m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1062]&~m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1062]&~m[1088]&~m[1089]&m[1091]&m[1092])|(m[1062]&~m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1062]&m[1088]&~m[1089]&m[1091]&m[1092])|(m[1062]&m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1062]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1062]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1062]&m[1088]&m[1089]&m[1091]&m[1092]))):InitCond[615];
    m[1095] = run?((((m[1067]&~m[1093]&~m[1094]&~m[1096]&~m[1097])|(~m[1067]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1067]&m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1067]&~m[1093]&m[1094]&m[1096]&~m[1097])|(~m[1067]&m[1093]&~m[1094]&~m[1096]&m[1097])|(~m[1067]&~m[1093]&m[1094]&~m[1096]&m[1097])|(m[1067]&m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1067]&m[1093]&m[1094]&m[1096]&m[1097]))&UnbiasedRNG[233])|((m[1067]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(~m[1067]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1067]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1067]&m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1067]&~m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1067]&~m[1093]&~m[1094]&m[1096]&m[1097])|(m[1067]&~m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1067]&m[1093]&~m[1094]&m[1096]&m[1097])|(m[1067]&m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1067]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1067]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1067]&m[1093]&m[1094]&m[1096]&m[1097]))):InitCond[616];
    m[1100] = run?((((m[1072]&~m[1098]&~m[1099]&~m[1101]&~m[1102])|(~m[1072]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1072]&m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1072]&~m[1098]&m[1099]&m[1101]&~m[1102])|(~m[1072]&m[1098]&~m[1099]&~m[1101]&m[1102])|(~m[1072]&~m[1098]&m[1099]&~m[1101]&m[1102])|(m[1072]&m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1072]&m[1098]&m[1099]&m[1101]&m[1102]))&UnbiasedRNG[234])|((m[1072]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(~m[1072]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1072]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1072]&m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1072]&~m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1072]&~m[1098]&~m[1099]&m[1101]&m[1102])|(m[1072]&~m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1072]&m[1098]&~m[1099]&m[1101]&m[1102])|(m[1072]&m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1072]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1072]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1072]&m[1098]&m[1099]&m[1101]&m[1102]))):InitCond[617];
    m[1105] = run?((((m[1077]&~m[1103]&~m[1104]&~m[1106]&~m[1107])|(~m[1077]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1077]&m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1077]&~m[1103]&m[1104]&m[1106]&~m[1107])|(~m[1077]&m[1103]&~m[1104]&~m[1106]&m[1107])|(~m[1077]&~m[1103]&m[1104]&~m[1106]&m[1107])|(m[1077]&m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1077]&m[1103]&m[1104]&m[1106]&m[1107]))&UnbiasedRNG[235])|((m[1077]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(~m[1077]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1077]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1077]&m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1077]&~m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1077]&~m[1103]&~m[1104]&m[1106]&m[1107])|(m[1077]&~m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1077]&m[1103]&~m[1104]&m[1106]&m[1107])|(m[1077]&m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1077]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1077]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1077]&m[1103]&m[1104]&m[1106]&m[1107]))):InitCond[618];
    m[1110] = run?((((m[1082]&~m[1108]&~m[1109]&~m[1111]&~m[1112])|(~m[1082]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1082]&m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1082]&~m[1108]&m[1109]&m[1111]&~m[1112])|(~m[1082]&m[1108]&~m[1109]&~m[1111]&m[1112])|(~m[1082]&~m[1108]&m[1109]&~m[1111]&m[1112])|(m[1082]&m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1082]&m[1108]&m[1109]&m[1111]&m[1112]))&UnbiasedRNG[236])|((m[1082]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(~m[1082]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1082]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1082]&m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1082]&~m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1082]&~m[1108]&~m[1109]&m[1111]&m[1112])|(m[1082]&~m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1082]&m[1108]&~m[1109]&m[1111]&m[1112])|(m[1082]&m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1082]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1082]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1082]&m[1108]&m[1109]&m[1111]&m[1112]))):InitCond[619];
    m[1115] = run?((((m[1092]&~m[1113]&~m[1114]&~m[1116]&~m[1117])|(~m[1092]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1092]&m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1092]&~m[1113]&m[1114]&m[1116]&~m[1117])|(~m[1092]&m[1113]&~m[1114]&~m[1116]&m[1117])|(~m[1092]&~m[1113]&m[1114]&~m[1116]&m[1117])|(m[1092]&m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1092]&m[1113]&m[1114]&m[1116]&m[1117]))&UnbiasedRNG[237])|((m[1092]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(~m[1092]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1092]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1092]&m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1092]&~m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1092]&~m[1113]&~m[1114]&m[1116]&m[1117])|(m[1092]&~m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1092]&m[1113]&~m[1114]&m[1116]&m[1117])|(m[1092]&m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1092]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1092]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1092]&m[1113]&m[1114]&m[1116]&m[1117]))):InitCond[620];
    m[1120] = run?((((m[1097]&~m[1118]&~m[1119]&~m[1121]&~m[1122])|(~m[1097]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1097]&m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1097]&~m[1118]&m[1119]&m[1121]&~m[1122])|(~m[1097]&m[1118]&~m[1119]&~m[1121]&m[1122])|(~m[1097]&~m[1118]&m[1119]&~m[1121]&m[1122])|(m[1097]&m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1097]&m[1118]&m[1119]&m[1121]&m[1122]))&UnbiasedRNG[238])|((m[1097]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(~m[1097]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1097]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1097]&m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1097]&~m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1097]&~m[1118]&~m[1119]&m[1121]&m[1122])|(m[1097]&~m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1097]&m[1118]&~m[1119]&m[1121]&m[1122])|(m[1097]&m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1097]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1097]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1097]&m[1118]&m[1119]&m[1121]&m[1122]))):InitCond[621];
    m[1125] = run?((((m[1102]&~m[1123]&~m[1124]&~m[1126]&~m[1127])|(~m[1102]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1102]&m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1102]&~m[1123]&m[1124]&m[1126]&~m[1127])|(~m[1102]&m[1123]&~m[1124]&~m[1126]&m[1127])|(~m[1102]&~m[1123]&m[1124]&~m[1126]&m[1127])|(m[1102]&m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1102]&m[1123]&m[1124]&m[1126]&m[1127]))&UnbiasedRNG[239])|((m[1102]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(~m[1102]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1102]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1102]&m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1102]&~m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1102]&~m[1123]&~m[1124]&m[1126]&m[1127])|(m[1102]&~m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1102]&m[1123]&~m[1124]&m[1126]&m[1127])|(m[1102]&m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1102]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1102]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1102]&m[1123]&m[1124]&m[1126]&m[1127]))):InitCond[622];
    m[1130] = run?((((m[1107]&~m[1128]&~m[1129]&~m[1131]&~m[1132])|(~m[1107]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1107]&m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1107]&~m[1128]&m[1129]&m[1131]&~m[1132])|(~m[1107]&m[1128]&~m[1129]&~m[1131]&m[1132])|(~m[1107]&~m[1128]&m[1129]&~m[1131]&m[1132])|(m[1107]&m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1107]&m[1128]&m[1129]&m[1131]&m[1132]))&UnbiasedRNG[240])|((m[1107]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(~m[1107]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1107]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1107]&m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1107]&~m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1107]&~m[1128]&~m[1129]&m[1131]&m[1132])|(m[1107]&~m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1107]&m[1128]&~m[1129]&m[1131]&m[1132])|(m[1107]&m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1107]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1107]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1107]&m[1128]&m[1129]&m[1131]&m[1132]))):InitCond[623];
    m[1135] = run?((((m[1112]&~m[1133]&~m[1134]&~m[1136]&~m[1137])|(~m[1112]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1112]&m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1112]&~m[1133]&m[1134]&m[1136]&~m[1137])|(~m[1112]&m[1133]&~m[1134]&~m[1136]&m[1137])|(~m[1112]&~m[1133]&m[1134]&~m[1136]&m[1137])|(m[1112]&m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1112]&m[1133]&m[1134]&m[1136]&m[1137]))&UnbiasedRNG[241])|((m[1112]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(~m[1112]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1112]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1112]&m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1112]&~m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1112]&~m[1133]&~m[1134]&m[1136]&m[1137])|(m[1112]&~m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1112]&m[1133]&~m[1134]&m[1136]&m[1137])|(m[1112]&m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1112]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1112]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1112]&m[1133]&m[1134]&m[1136]&m[1137]))):InitCond[624];
    m[1140] = run?((((m[1122]&~m[1138]&~m[1139]&~m[1141]&~m[1142])|(~m[1122]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1122]&m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1122]&~m[1138]&m[1139]&m[1141]&~m[1142])|(~m[1122]&m[1138]&~m[1139]&~m[1141]&m[1142])|(~m[1122]&~m[1138]&m[1139]&~m[1141]&m[1142])|(m[1122]&m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1122]&m[1138]&m[1139]&m[1141]&m[1142]))&UnbiasedRNG[242])|((m[1122]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(~m[1122]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1122]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1122]&m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1122]&~m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1122]&~m[1138]&~m[1139]&m[1141]&m[1142])|(m[1122]&~m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1122]&m[1138]&~m[1139]&m[1141]&m[1142])|(m[1122]&m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1122]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1122]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1122]&m[1138]&m[1139]&m[1141]&m[1142]))):InitCond[625];
    m[1145] = run?((((m[1127]&~m[1143]&~m[1144]&~m[1146]&~m[1147])|(~m[1127]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1127]&m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1127]&~m[1143]&m[1144]&m[1146]&~m[1147])|(~m[1127]&m[1143]&~m[1144]&~m[1146]&m[1147])|(~m[1127]&~m[1143]&m[1144]&~m[1146]&m[1147])|(m[1127]&m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1127]&m[1143]&m[1144]&m[1146]&m[1147]))&UnbiasedRNG[243])|((m[1127]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(~m[1127]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1127]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1127]&m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1127]&~m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1127]&~m[1143]&~m[1144]&m[1146]&m[1147])|(m[1127]&~m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1127]&m[1143]&~m[1144]&m[1146]&m[1147])|(m[1127]&m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1127]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1127]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1127]&m[1143]&m[1144]&m[1146]&m[1147]))):InitCond[626];
    m[1150] = run?((((m[1132]&~m[1148]&~m[1149]&~m[1151]&~m[1152])|(~m[1132]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1132]&m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1132]&~m[1148]&m[1149]&m[1151]&~m[1152])|(~m[1132]&m[1148]&~m[1149]&~m[1151]&m[1152])|(~m[1132]&~m[1148]&m[1149]&~m[1151]&m[1152])|(m[1132]&m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1132]&m[1148]&m[1149]&m[1151]&m[1152]))&UnbiasedRNG[244])|((m[1132]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(~m[1132]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1132]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1132]&m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1132]&~m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1132]&~m[1148]&~m[1149]&m[1151]&m[1152])|(m[1132]&~m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1132]&m[1148]&~m[1149]&m[1151]&m[1152])|(m[1132]&m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1132]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1132]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1132]&m[1148]&m[1149]&m[1151]&m[1152]))):InitCond[627];
    m[1155] = run?((((m[1137]&~m[1153]&~m[1154]&~m[1156]&~m[1157])|(~m[1137]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1137]&m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1137]&~m[1153]&m[1154]&m[1156]&~m[1157])|(~m[1137]&m[1153]&~m[1154]&~m[1156]&m[1157])|(~m[1137]&~m[1153]&m[1154]&~m[1156]&m[1157])|(m[1137]&m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1137]&m[1153]&m[1154]&m[1156]&m[1157]))&UnbiasedRNG[245])|((m[1137]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(~m[1137]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1137]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1137]&m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1137]&~m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1137]&~m[1153]&~m[1154]&m[1156]&m[1157])|(m[1137]&~m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1137]&m[1153]&~m[1154]&m[1156]&m[1157])|(m[1137]&m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1137]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1137]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1137]&m[1153]&m[1154]&m[1156]&m[1157]))):InitCond[628];
    m[1160] = run?((((m[1147]&~m[1158]&~m[1159]&~m[1161]&~m[1162])|(~m[1147]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1147]&m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1147]&~m[1158]&m[1159]&m[1161]&~m[1162])|(~m[1147]&m[1158]&~m[1159]&~m[1161]&m[1162])|(~m[1147]&~m[1158]&m[1159]&~m[1161]&m[1162])|(m[1147]&m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1147]&m[1158]&m[1159]&m[1161]&m[1162]))&UnbiasedRNG[246])|((m[1147]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(~m[1147]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1147]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1147]&m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1147]&~m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1147]&~m[1158]&~m[1159]&m[1161]&m[1162])|(m[1147]&~m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1147]&m[1158]&~m[1159]&m[1161]&m[1162])|(m[1147]&m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1147]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1147]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1147]&m[1158]&m[1159]&m[1161]&m[1162]))):InitCond[629];
    m[1165] = run?((((m[1152]&~m[1163]&~m[1164]&~m[1166]&~m[1167])|(~m[1152]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1152]&m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1152]&~m[1163]&m[1164]&m[1166]&~m[1167])|(~m[1152]&m[1163]&~m[1164]&~m[1166]&m[1167])|(~m[1152]&~m[1163]&m[1164]&~m[1166]&m[1167])|(m[1152]&m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1152]&m[1163]&m[1164]&m[1166]&m[1167]))&UnbiasedRNG[247])|((m[1152]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(~m[1152]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1152]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1152]&m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1152]&~m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1152]&~m[1163]&~m[1164]&m[1166]&m[1167])|(m[1152]&~m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1152]&m[1163]&~m[1164]&m[1166]&m[1167])|(m[1152]&m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1152]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1152]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1152]&m[1163]&m[1164]&m[1166]&m[1167]))):InitCond[630];
    m[1170] = run?((((m[1157]&~m[1168]&~m[1169]&~m[1171]&~m[1172])|(~m[1157]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1157]&m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1157]&~m[1168]&m[1169]&m[1171]&~m[1172])|(~m[1157]&m[1168]&~m[1169]&~m[1171]&m[1172])|(~m[1157]&~m[1168]&m[1169]&~m[1171]&m[1172])|(m[1157]&m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1157]&m[1168]&m[1169]&m[1171]&m[1172]))&UnbiasedRNG[248])|((m[1157]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(~m[1157]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1157]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1157]&m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1157]&~m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1157]&~m[1168]&~m[1169]&m[1171]&m[1172])|(m[1157]&~m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1157]&m[1168]&~m[1169]&m[1171]&m[1172])|(m[1157]&m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1157]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1157]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1157]&m[1168]&m[1169]&m[1171]&m[1172]))):InitCond[631];
    m[1175] = run?((((m[1167]&~m[1173]&~m[1174]&~m[1176]&~m[1177])|(~m[1167]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1167]&m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1167]&~m[1173]&m[1174]&m[1176]&~m[1177])|(~m[1167]&m[1173]&~m[1174]&~m[1176]&m[1177])|(~m[1167]&~m[1173]&m[1174]&~m[1176]&m[1177])|(m[1167]&m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1167]&m[1173]&m[1174]&m[1176]&m[1177]))&UnbiasedRNG[249])|((m[1167]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(~m[1167]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1167]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1167]&m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1167]&~m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1167]&~m[1173]&~m[1174]&m[1176]&m[1177])|(m[1167]&~m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1167]&m[1173]&~m[1174]&m[1176]&m[1177])|(m[1167]&m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1167]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1167]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1167]&m[1173]&m[1174]&m[1176]&m[1177]))):InitCond[632];
    m[1180] = run?((((m[1172]&~m[1178]&~m[1179]&~m[1181]&~m[1182])|(~m[1172]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1172]&m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1172]&~m[1178]&m[1179]&m[1181]&~m[1182])|(~m[1172]&m[1178]&~m[1179]&~m[1181]&m[1182])|(~m[1172]&~m[1178]&m[1179]&~m[1181]&m[1182])|(m[1172]&m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1172]&m[1178]&m[1179]&m[1181]&m[1182]))&UnbiasedRNG[250])|((m[1172]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(~m[1172]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1172]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1172]&m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1172]&~m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1172]&~m[1178]&~m[1179]&m[1181]&m[1182])|(m[1172]&~m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1172]&m[1178]&~m[1179]&m[1181]&m[1182])|(m[1172]&m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1172]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1172]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1172]&m[1178]&m[1179]&m[1181]&m[1182]))):InitCond[633];
    m[1185] = run?((((m[1182]&~m[1183]&~m[1184]&~m[1186]&~m[1187])|(~m[1182]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1182]&m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1182]&~m[1183]&m[1184]&m[1186]&~m[1187])|(~m[1182]&m[1183]&~m[1184]&~m[1186]&m[1187])|(~m[1182]&~m[1183]&m[1184]&~m[1186]&m[1187])|(m[1182]&m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1182]&m[1183]&m[1184]&m[1186]&m[1187]))&UnbiasedRNG[251])|((m[1182]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(~m[1182]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1182]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1182]&m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1182]&~m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1182]&~m[1183]&~m[1184]&m[1186]&m[1187])|(m[1182]&~m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1182]&m[1183]&~m[1184]&m[1186]&m[1187])|(m[1182]&m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1182]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1182]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1182]&m[1183]&m[1184]&m[1186]&m[1187]))):InitCond[634];
end

always @(posedge color2_clk) begin
    m[240] = run?((((~m[60]&~m[96]&~m[384])|(m[60]&m[96]&~m[384]))&BiasedRNG[383])|(((m[60]&~m[96]&~m[384])|(~m[60]&m[96]&m[384]))&~BiasedRNG[383])|((~m[60]&~m[96]&m[384])|(m[60]&~m[96]&m[384])|(m[60]&m[96]&m[384]))):InitCond[635];
    m[241] = run?((((~m[60]&~m[108]&~m[385])|(m[60]&m[108]&~m[385]))&BiasedRNG[384])|(((m[60]&~m[108]&~m[385])|(~m[60]&m[108]&m[385]))&~BiasedRNG[384])|((~m[60]&~m[108]&m[385])|(m[60]&~m[108]&m[385])|(m[60]&m[108]&m[385]))):InitCond[636];
    m[242] = run?((((~m[60]&~m[120]&~m[386])|(m[60]&m[120]&~m[386]))&BiasedRNG[385])|(((m[60]&~m[120]&~m[386])|(~m[60]&m[120]&m[386]))&~BiasedRNG[385])|((~m[60]&~m[120]&m[386])|(m[60]&~m[120]&m[386])|(m[60]&m[120]&m[386]))):InitCond[637];
    m[243] = run?((((~m[60]&~m[132]&~m[387])|(m[60]&m[132]&~m[387]))&BiasedRNG[386])|(((m[60]&~m[132]&~m[387])|(~m[60]&m[132]&m[387]))&~BiasedRNG[386])|((~m[60]&~m[132]&m[387])|(m[60]&~m[132]&m[387])|(m[60]&m[132]&m[387]))):InitCond[638];
    m[244] = run?((((~m[61]&~m[144]&~m[388])|(m[61]&m[144]&~m[388]))&BiasedRNG[387])|(((m[61]&~m[144]&~m[388])|(~m[61]&m[144]&m[388]))&~BiasedRNG[387])|((~m[61]&~m[144]&m[388])|(m[61]&~m[144]&m[388])|(m[61]&m[144]&m[388]))):InitCond[639];
    m[245] = run?((((~m[61]&~m[156]&~m[389])|(m[61]&m[156]&~m[389]))&BiasedRNG[388])|(((m[61]&~m[156]&~m[389])|(~m[61]&m[156]&m[389]))&~BiasedRNG[388])|((~m[61]&~m[156]&m[389])|(m[61]&~m[156]&m[389])|(m[61]&m[156]&m[389]))):InitCond[640];
    m[246] = run?((((~m[61]&~m[168]&~m[390])|(m[61]&m[168]&~m[390]))&BiasedRNG[389])|(((m[61]&~m[168]&~m[390])|(~m[61]&m[168]&m[390]))&~BiasedRNG[389])|((~m[61]&~m[168]&m[390])|(m[61]&~m[168]&m[390])|(m[61]&m[168]&m[390]))):InitCond[641];
    m[247] = run?((((~m[61]&~m[180]&~m[391])|(m[61]&m[180]&~m[391]))&BiasedRNG[390])|(((m[61]&~m[180]&~m[391])|(~m[61]&m[180]&m[391]))&~BiasedRNG[390])|((~m[61]&~m[180]&m[391])|(m[61]&~m[180]&m[391])|(m[61]&m[180]&m[391]))):InitCond[642];
    m[248] = run?((((~m[62]&~m[192]&~m[392])|(m[62]&m[192]&~m[392]))&BiasedRNG[391])|(((m[62]&~m[192]&~m[392])|(~m[62]&m[192]&m[392]))&~BiasedRNG[391])|((~m[62]&~m[192]&m[392])|(m[62]&~m[192]&m[392])|(m[62]&m[192]&m[392]))):InitCond[643];
    m[249] = run?((((~m[62]&~m[204]&~m[393])|(m[62]&m[204]&~m[393]))&BiasedRNG[392])|(((m[62]&~m[204]&~m[393])|(~m[62]&m[204]&m[393]))&~BiasedRNG[392])|((~m[62]&~m[204]&m[393])|(m[62]&~m[204]&m[393])|(m[62]&m[204]&m[393]))):InitCond[644];
    m[250] = run?((((~m[62]&~m[216]&~m[394])|(m[62]&m[216]&~m[394]))&BiasedRNG[393])|(((m[62]&~m[216]&~m[394])|(~m[62]&m[216]&m[394]))&~BiasedRNG[393])|((~m[62]&~m[216]&m[394])|(m[62]&~m[216]&m[394])|(m[62]&m[216]&m[394]))):InitCond[645];
    m[251] = run?((((~m[62]&~m[228]&~m[395])|(m[62]&m[228]&~m[395]))&BiasedRNG[394])|(((m[62]&~m[228]&~m[395])|(~m[62]&m[228]&m[395]))&~BiasedRNG[394])|((~m[62]&~m[228]&m[395])|(m[62]&~m[228]&m[395])|(m[62]&m[228]&m[395]))):InitCond[646];
    m[252] = run?((((~m[63]&~m[97]&~m[396])|(m[63]&m[97]&~m[396]))&BiasedRNG[395])|(((m[63]&~m[97]&~m[396])|(~m[63]&m[97]&m[396]))&~BiasedRNG[395])|((~m[63]&~m[97]&m[396])|(m[63]&~m[97]&m[396])|(m[63]&m[97]&m[396]))):InitCond[647];
    m[253] = run?((((~m[63]&~m[109]&~m[397])|(m[63]&m[109]&~m[397]))&BiasedRNG[396])|(((m[63]&~m[109]&~m[397])|(~m[63]&m[109]&m[397]))&~BiasedRNG[396])|((~m[63]&~m[109]&m[397])|(m[63]&~m[109]&m[397])|(m[63]&m[109]&m[397]))):InitCond[648];
    m[254] = run?((((~m[63]&~m[121]&~m[398])|(m[63]&m[121]&~m[398]))&BiasedRNG[397])|(((m[63]&~m[121]&~m[398])|(~m[63]&m[121]&m[398]))&~BiasedRNG[397])|((~m[63]&~m[121]&m[398])|(m[63]&~m[121]&m[398])|(m[63]&m[121]&m[398]))):InitCond[649];
    m[255] = run?((((~m[63]&~m[133]&~m[399])|(m[63]&m[133]&~m[399]))&BiasedRNG[398])|(((m[63]&~m[133]&~m[399])|(~m[63]&m[133]&m[399]))&~BiasedRNG[398])|((~m[63]&~m[133]&m[399])|(m[63]&~m[133]&m[399])|(m[63]&m[133]&m[399]))):InitCond[650];
    m[256] = run?((((~m[64]&~m[145]&~m[400])|(m[64]&m[145]&~m[400]))&BiasedRNG[399])|(((m[64]&~m[145]&~m[400])|(~m[64]&m[145]&m[400]))&~BiasedRNG[399])|((~m[64]&~m[145]&m[400])|(m[64]&~m[145]&m[400])|(m[64]&m[145]&m[400]))):InitCond[651];
    m[257] = run?((((~m[64]&~m[157]&~m[401])|(m[64]&m[157]&~m[401]))&BiasedRNG[400])|(((m[64]&~m[157]&~m[401])|(~m[64]&m[157]&m[401]))&~BiasedRNG[400])|((~m[64]&~m[157]&m[401])|(m[64]&~m[157]&m[401])|(m[64]&m[157]&m[401]))):InitCond[652];
    m[258] = run?((((~m[64]&~m[169]&~m[402])|(m[64]&m[169]&~m[402]))&BiasedRNG[401])|(((m[64]&~m[169]&~m[402])|(~m[64]&m[169]&m[402]))&~BiasedRNG[401])|((~m[64]&~m[169]&m[402])|(m[64]&~m[169]&m[402])|(m[64]&m[169]&m[402]))):InitCond[653];
    m[259] = run?((((~m[64]&~m[181]&~m[403])|(m[64]&m[181]&~m[403]))&BiasedRNG[402])|(((m[64]&~m[181]&~m[403])|(~m[64]&m[181]&m[403]))&~BiasedRNG[402])|((~m[64]&~m[181]&m[403])|(m[64]&~m[181]&m[403])|(m[64]&m[181]&m[403]))):InitCond[654];
    m[260] = run?((((~m[65]&~m[193]&~m[404])|(m[65]&m[193]&~m[404]))&BiasedRNG[403])|(((m[65]&~m[193]&~m[404])|(~m[65]&m[193]&m[404]))&~BiasedRNG[403])|((~m[65]&~m[193]&m[404])|(m[65]&~m[193]&m[404])|(m[65]&m[193]&m[404]))):InitCond[655];
    m[261] = run?((((~m[65]&~m[205]&~m[405])|(m[65]&m[205]&~m[405]))&BiasedRNG[404])|(((m[65]&~m[205]&~m[405])|(~m[65]&m[205]&m[405]))&~BiasedRNG[404])|((~m[65]&~m[205]&m[405])|(m[65]&~m[205]&m[405])|(m[65]&m[205]&m[405]))):InitCond[656];
    m[262] = run?((((~m[65]&~m[217]&~m[406])|(m[65]&m[217]&~m[406]))&BiasedRNG[405])|(((m[65]&~m[217]&~m[406])|(~m[65]&m[217]&m[406]))&~BiasedRNG[405])|((~m[65]&~m[217]&m[406])|(m[65]&~m[217]&m[406])|(m[65]&m[217]&m[406]))):InitCond[657];
    m[263] = run?((((~m[65]&~m[229]&~m[407])|(m[65]&m[229]&~m[407]))&BiasedRNG[406])|(((m[65]&~m[229]&~m[407])|(~m[65]&m[229]&m[407]))&~BiasedRNG[406])|((~m[65]&~m[229]&m[407])|(m[65]&~m[229]&m[407])|(m[65]&m[229]&m[407]))):InitCond[658];
    m[264] = run?((((~m[66]&~m[98]&~m[408])|(m[66]&m[98]&~m[408]))&BiasedRNG[407])|(((m[66]&~m[98]&~m[408])|(~m[66]&m[98]&m[408]))&~BiasedRNG[407])|((~m[66]&~m[98]&m[408])|(m[66]&~m[98]&m[408])|(m[66]&m[98]&m[408]))):InitCond[659];
    m[265] = run?((((~m[66]&~m[110]&~m[409])|(m[66]&m[110]&~m[409]))&BiasedRNG[408])|(((m[66]&~m[110]&~m[409])|(~m[66]&m[110]&m[409]))&~BiasedRNG[408])|((~m[66]&~m[110]&m[409])|(m[66]&~m[110]&m[409])|(m[66]&m[110]&m[409]))):InitCond[660];
    m[266] = run?((((~m[66]&~m[122]&~m[410])|(m[66]&m[122]&~m[410]))&BiasedRNG[409])|(((m[66]&~m[122]&~m[410])|(~m[66]&m[122]&m[410]))&~BiasedRNG[409])|((~m[66]&~m[122]&m[410])|(m[66]&~m[122]&m[410])|(m[66]&m[122]&m[410]))):InitCond[661];
    m[267] = run?((((~m[66]&~m[134]&~m[411])|(m[66]&m[134]&~m[411]))&BiasedRNG[410])|(((m[66]&~m[134]&~m[411])|(~m[66]&m[134]&m[411]))&~BiasedRNG[410])|((~m[66]&~m[134]&m[411])|(m[66]&~m[134]&m[411])|(m[66]&m[134]&m[411]))):InitCond[662];
    m[268] = run?((((~m[67]&~m[146]&~m[412])|(m[67]&m[146]&~m[412]))&BiasedRNG[411])|(((m[67]&~m[146]&~m[412])|(~m[67]&m[146]&m[412]))&~BiasedRNG[411])|((~m[67]&~m[146]&m[412])|(m[67]&~m[146]&m[412])|(m[67]&m[146]&m[412]))):InitCond[663];
    m[269] = run?((((~m[67]&~m[158]&~m[413])|(m[67]&m[158]&~m[413]))&BiasedRNG[412])|(((m[67]&~m[158]&~m[413])|(~m[67]&m[158]&m[413]))&~BiasedRNG[412])|((~m[67]&~m[158]&m[413])|(m[67]&~m[158]&m[413])|(m[67]&m[158]&m[413]))):InitCond[664];
    m[270] = run?((((~m[67]&~m[170]&~m[414])|(m[67]&m[170]&~m[414]))&BiasedRNG[413])|(((m[67]&~m[170]&~m[414])|(~m[67]&m[170]&m[414]))&~BiasedRNG[413])|((~m[67]&~m[170]&m[414])|(m[67]&~m[170]&m[414])|(m[67]&m[170]&m[414]))):InitCond[665];
    m[271] = run?((((~m[67]&~m[182]&~m[415])|(m[67]&m[182]&~m[415]))&BiasedRNG[414])|(((m[67]&~m[182]&~m[415])|(~m[67]&m[182]&m[415]))&~BiasedRNG[414])|((~m[67]&~m[182]&m[415])|(m[67]&~m[182]&m[415])|(m[67]&m[182]&m[415]))):InitCond[666];
    m[272] = run?((((~m[68]&~m[194]&~m[416])|(m[68]&m[194]&~m[416]))&BiasedRNG[415])|(((m[68]&~m[194]&~m[416])|(~m[68]&m[194]&m[416]))&~BiasedRNG[415])|((~m[68]&~m[194]&m[416])|(m[68]&~m[194]&m[416])|(m[68]&m[194]&m[416]))):InitCond[667];
    m[273] = run?((((~m[68]&~m[206]&~m[417])|(m[68]&m[206]&~m[417]))&BiasedRNG[416])|(((m[68]&~m[206]&~m[417])|(~m[68]&m[206]&m[417]))&~BiasedRNG[416])|((~m[68]&~m[206]&m[417])|(m[68]&~m[206]&m[417])|(m[68]&m[206]&m[417]))):InitCond[668];
    m[274] = run?((((~m[68]&~m[218]&~m[418])|(m[68]&m[218]&~m[418]))&BiasedRNG[417])|(((m[68]&~m[218]&~m[418])|(~m[68]&m[218]&m[418]))&~BiasedRNG[417])|((~m[68]&~m[218]&m[418])|(m[68]&~m[218]&m[418])|(m[68]&m[218]&m[418]))):InitCond[669];
    m[275] = run?((((~m[68]&~m[230]&~m[419])|(m[68]&m[230]&~m[419]))&BiasedRNG[418])|(((m[68]&~m[230]&~m[419])|(~m[68]&m[230]&m[419]))&~BiasedRNG[418])|((~m[68]&~m[230]&m[419])|(m[68]&~m[230]&m[419])|(m[68]&m[230]&m[419]))):InitCond[670];
    m[276] = run?((((~m[69]&~m[99]&~m[420])|(m[69]&m[99]&~m[420]))&BiasedRNG[419])|(((m[69]&~m[99]&~m[420])|(~m[69]&m[99]&m[420]))&~BiasedRNG[419])|((~m[69]&~m[99]&m[420])|(m[69]&~m[99]&m[420])|(m[69]&m[99]&m[420]))):InitCond[671];
    m[277] = run?((((~m[69]&~m[111]&~m[421])|(m[69]&m[111]&~m[421]))&BiasedRNG[420])|(((m[69]&~m[111]&~m[421])|(~m[69]&m[111]&m[421]))&~BiasedRNG[420])|((~m[69]&~m[111]&m[421])|(m[69]&~m[111]&m[421])|(m[69]&m[111]&m[421]))):InitCond[672];
    m[278] = run?((((~m[69]&~m[123]&~m[422])|(m[69]&m[123]&~m[422]))&BiasedRNG[421])|(((m[69]&~m[123]&~m[422])|(~m[69]&m[123]&m[422]))&~BiasedRNG[421])|((~m[69]&~m[123]&m[422])|(m[69]&~m[123]&m[422])|(m[69]&m[123]&m[422]))):InitCond[673];
    m[279] = run?((((~m[69]&~m[135]&~m[423])|(m[69]&m[135]&~m[423]))&BiasedRNG[422])|(((m[69]&~m[135]&~m[423])|(~m[69]&m[135]&m[423]))&~BiasedRNG[422])|((~m[69]&~m[135]&m[423])|(m[69]&~m[135]&m[423])|(m[69]&m[135]&m[423]))):InitCond[674];
    m[280] = run?((((~m[70]&~m[147]&~m[424])|(m[70]&m[147]&~m[424]))&BiasedRNG[423])|(((m[70]&~m[147]&~m[424])|(~m[70]&m[147]&m[424]))&~BiasedRNG[423])|((~m[70]&~m[147]&m[424])|(m[70]&~m[147]&m[424])|(m[70]&m[147]&m[424]))):InitCond[675];
    m[281] = run?((((~m[70]&~m[159]&~m[425])|(m[70]&m[159]&~m[425]))&BiasedRNG[424])|(((m[70]&~m[159]&~m[425])|(~m[70]&m[159]&m[425]))&~BiasedRNG[424])|((~m[70]&~m[159]&m[425])|(m[70]&~m[159]&m[425])|(m[70]&m[159]&m[425]))):InitCond[676];
    m[282] = run?((((~m[70]&~m[171]&~m[426])|(m[70]&m[171]&~m[426]))&BiasedRNG[425])|(((m[70]&~m[171]&~m[426])|(~m[70]&m[171]&m[426]))&~BiasedRNG[425])|((~m[70]&~m[171]&m[426])|(m[70]&~m[171]&m[426])|(m[70]&m[171]&m[426]))):InitCond[677];
    m[283] = run?((((~m[70]&~m[183]&~m[427])|(m[70]&m[183]&~m[427]))&BiasedRNG[426])|(((m[70]&~m[183]&~m[427])|(~m[70]&m[183]&m[427]))&~BiasedRNG[426])|((~m[70]&~m[183]&m[427])|(m[70]&~m[183]&m[427])|(m[70]&m[183]&m[427]))):InitCond[678];
    m[284] = run?((((~m[71]&~m[195]&~m[428])|(m[71]&m[195]&~m[428]))&BiasedRNG[427])|(((m[71]&~m[195]&~m[428])|(~m[71]&m[195]&m[428]))&~BiasedRNG[427])|((~m[71]&~m[195]&m[428])|(m[71]&~m[195]&m[428])|(m[71]&m[195]&m[428]))):InitCond[679];
    m[285] = run?((((~m[71]&~m[207]&~m[429])|(m[71]&m[207]&~m[429]))&BiasedRNG[428])|(((m[71]&~m[207]&~m[429])|(~m[71]&m[207]&m[429]))&~BiasedRNG[428])|((~m[71]&~m[207]&m[429])|(m[71]&~m[207]&m[429])|(m[71]&m[207]&m[429]))):InitCond[680];
    m[286] = run?((((~m[71]&~m[219]&~m[430])|(m[71]&m[219]&~m[430]))&BiasedRNG[429])|(((m[71]&~m[219]&~m[430])|(~m[71]&m[219]&m[430]))&~BiasedRNG[429])|((~m[71]&~m[219]&m[430])|(m[71]&~m[219]&m[430])|(m[71]&m[219]&m[430]))):InitCond[681];
    m[287] = run?((((~m[71]&~m[231]&~m[431])|(m[71]&m[231]&~m[431]))&BiasedRNG[430])|(((m[71]&~m[231]&~m[431])|(~m[71]&m[231]&m[431]))&~BiasedRNG[430])|((~m[71]&~m[231]&m[431])|(m[71]&~m[231]&m[431])|(m[71]&m[231]&m[431]))):InitCond[682];
    m[288] = run?((((~m[72]&~m[100]&~m[432])|(m[72]&m[100]&~m[432]))&BiasedRNG[431])|(((m[72]&~m[100]&~m[432])|(~m[72]&m[100]&m[432]))&~BiasedRNG[431])|((~m[72]&~m[100]&m[432])|(m[72]&~m[100]&m[432])|(m[72]&m[100]&m[432]))):InitCond[683];
    m[289] = run?((((~m[72]&~m[112]&~m[433])|(m[72]&m[112]&~m[433]))&BiasedRNG[432])|(((m[72]&~m[112]&~m[433])|(~m[72]&m[112]&m[433]))&~BiasedRNG[432])|((~m[72]&~m[112]&m[433])|(m[72]&~m[112]&m[433])|(m[72]&m[112]&m[433]))):InitCond[684];
    m[290] = run?((((~m[72]&~m[124]&~m[434])|(m[72]&m[124]&~m[434]))&BiasedRNG[433])|(((m[72]&~m[124]&~m[434])|(~m[72]&m[124]&m[434]))&~BiasedRNG[433])|((~m[72]&~m[124]&m[434])|(m[72]&~m[124]&m[434])|(m[72]&m[124]&m[434]))):InitCond[685];
    m[291] = run?((((~m[72]&~m[136]&~m[435])|(m[72]&m[136]&~m[435]))&BiasedRNG[434])|(((m[72]&~m[136]&~m[435])|(~m[72]&m[136]&m[435]))&~BiasedRNG[434])|((~m[72]&~m[136]&m[435])|(m[72]&~m[136]&m[435])|(m[72]&m[136]&m[435]))):InitCond[686];
    m[292] = run?((((~m[73]&~m[148]&~m[436])|(m[73]&m[148]&~m[436]))&BiasedRNG[435])|(((m[73]&~m[148]&~m[436])|(~m[73]&m[148]&m[436]))&~BiasedRNG[435])|((~m[73]&~m[148]&m[436])|(m[73]&~m[148]&m[436])|(m[73]&m[148]&m[436]))):InitCond[687];
    m[293] = run?((((~m[73]&~m[160]&~m[437])|(m[73]&m[160]&~m[437]))&BiasedRNG[436])|(((m[73]&~m[160]&~m[437])|(~m[73]&m[160]&m[437]))&~BiasedRNG[436])|((~m[73]&~m[160]&m[437])|(m[73]&~m[160]&m[437])|(m[73]&m[160]&m[437]))):InitCond[688];
    m[294] = run?((((~m[73]&~m[172]&~m[438])|(m[73]&m[172]&~m[438]))&BiasedRNG[437])|(((m[73]&~m[172]&~m[438])|(~m[73]&m[172]&m[438]))&~BiasedRNG[437])|((~m[73]&~m[172]&m[438])|(m[73]&~m[172]&m[438])|(m[73]&m[172]&m[438]))):InitCond[689];
    m[295] = run?((((~m[73]&~m[184]&~m[439])|(m[73]&m[184]&~m[439]))&BiasedRNG[438])|(((m[73]&~m[184]&~m[439])|(~m[73]&m[184]&m[439]))&~BiasedRNG[438])|((~m[73]&~m[184]&m[439])|(m[73]&~m[184]&m[439])|(m[73]&m[184]&m[439]))):InitCond[690];
    m[296] = run?((((~m[74]&~m[196]&~m[440])|(m[74]&m[196]&~m[440]))&BiasedRNG[439])|(((m[74]&~m[196]&~m[440])|(~m[74]&m[196]&m[440]))&~BiasedRNG[439])|((~m[74]&~m[196]&m[440])|(m[74]&~m[196]&m[440])|(m[74]&m[196]&m[440]))):InitCond[691];
    m[297] = run?((((~m[74]&~m[208]&~m[441])|(m[74]&m[208]&~m[441]))&BiasedRNG[440])|(((m[74]&~m[208]&~m[441])|(~m[74]&m[208]&m[441]))&~BiasedRNG[440])|((~m[74]&~m[208]&m[441])|(m[74]&~m[208]&m[441])|(m[74]&m[208]&m[441]))):InitCond[692];
    m[298] = run?((((~m[74]&~m[220]&~m[442])|(m[74]&m[220]&~m[442]))&BiasedRNG[441])|(((m[74]&~m[220]&~m[442])|(~m[74]&m[220]&m[442]))&~BiasedRNG[441])|((~m[74]&~m[220]&m[442])|(m[74]&~m[220]&m[442])|(m[74]&m[220]&m[442]))):InitCond[693];
    m[299] = run?((((~m[74]&~m[232]&~m[443])|(m[74]&m[232]&~m[443]))&BiasedRNG[442])|(((m[74]&~m[232]&~m[443])|(~m[74]&m[232]&m[443]))&~BiasedRNG[442])|((~m[74]&~m[232]&m[443])|(m[74]&~m[232]&m[443])|(m[74]&m[232]&m[443]))):InitCond[694];
    m[300] = run?((((~m[75]&~m[101]&~m[444])|(m[75]&m[101]&~m[444]))&BiasedRNG[443])|(((m[75]&~m[101]&~m[444])|(~m[75]&m[101]&m[444]))&~BiasedRNG[443])|((~m[75]&~m[101]&m[444])|(m[75]&~m[101]&m[444])|(m[75]&m[101]&m[444]))):InitCond[695];
    m[301] = run?((((~m[75]&~m[113]&~m[445])|(m[75]&m[113]&~m[445]))&BiasedRNG[444])|(((m[75]&~m[113]&~m[445])|(~m[75]&m[113]&m[445]))&~BiasedRNG[444])|((~m[75]&~m[113]&m[445])|(m[75]&~m[113]&m[445])|(m[75]&m[113]&m[445]))):InitCond[696];
    m[302] = run?((((~m[75]&~m[125]&~m[446])|(m[75]&m[125]&~m[446]))&BiasedRNG[445])|(((m[75]&~m[125]&~m[446])|(~m[75]&m[125]&m[446]))&~BiasedRNG[445])|((~m[75]&~m[125]&m[446])|(m[75]&~m[125]&m[446])|(m[75]&m[125]&m[446]))):InitCond[697];
    m[303] = run?((((~m[75]&~m[137]&~m[447])|(m[75]&m[137]&~m[447]))&BiasedRNG[446])|(((m[75]&~m[137]&~m[447])|(~m[75]&m[137]&m[447]))&~BiasedRNG[446])|((~m[75]&~m[137]&m[447])|(m[75]&~m[137]&m[447])|(m[75]&m[137]&m[447]))):InitCond[698];
    m[304] = run?((((~m[76]&~m[149]&~m[448])|(m[76]&m[149]&~m[448]))&BiasedRNG[447])|(((m[76]&~m[149]&~m[448])|(~m[76]&m[149]&m[448]))&~BiasedRNG[447])|((~m[76]&~m[149]&m[448])|(m[76]&~m[149]&m[448])|(m[76]&m[149]&m[448]))):InitCond[699];
    m[305] = run?((((~m[76]&~m[161]&~m[449])|(m[76]&m[161]&~m[449]))&BiasedRNG[448])|(((m[76]&~m[161]&~m[449])|(~m[76]&m[161]&m[449]))&~BiasedRNG[448])|((~m[76]&~m[161]&m[449])|(m[76]&~m[161]&m[449])|(m[76]&m[161]&m[449]))):InitCond[700];
    m[306] = run?((((~m[76]&~m[173]&~m[450])|(m[76]&m[173]&~m[450]))&BiasedRNG[449])|(((m[76]&~m[173]&~m[450])|(~m[76]&m[173]&m[450]))&~BiasedRNG[449])|((~m[76]&~m[173]&m[450])|(m[76]&~m[173]&m[450])|(m[76]&m[173]&m[450]))):InitCond[701];
    m[307] = run?((((~m[76]&~m[185]&~m[451])|(m[76]&m[185]&~m[451]))&BiasedRNG[450])|(((m[76]&~m[185]&~m[451])|(~m[76]&m[185]&m[451]))&~BiasedRNG[450])|((~m[76]&~m[185]&m[451])|(m[76]&~m[185]&m[451])|(m[76]&m[185]&m[451]))):InitCond[702];
    m[308] = run?((((~m[77]&~m[197]&~m[452])|(m[77]&m[197]&~m[452]))&BiasedRNG[451])|(((m[77]&~m[197]&~m[452])|(~m[77]&m[197]&m[452]))&~BiasedRNG[451])|((~m[77]&~m[197]&m[452])|(m[77]&~m[197]&m[452])|(m[77]&m[197]&m[452]))):InitCond[703];
    m[309] = run?((((~m[77]&~m[209]&~m[453])|(m[77]&m[209]&~m[453]))&BiasedRNG[452])|(((m[77]&~m[209]&~m[453])|(~m[77]&m[209]&m[453]))&~BiasedRNG[452])|((~m[77]&~m[209]&m[453])|(m[77]&~m[209]&m[453])|(m[77]&m[209]&m[453]))):InitCond[704];
    m[310] = run?((((~m[77]&~m[221]&~m[454])|(m[77]&m[221]&~m[454]))&BiasedRNG[453])|(((m[77]&~m[221]&~m[454])|(~m[77]&m[221]&m[454]))&~BiasedRNG[453])|((~m[77]&~m[221]&m[454])|(m[77]&~m[221]&m[454])|(m[77]&m[221]&m[454]))):InitCond[705];
    m[311] = run?((((~m[77]&~m[233]&~m[455])|(m[77]&m[233]&~m[455]))&BiasedRNG[454])|(((m[77]&~m[233]&~m[455])|(~m[77]&m[233]&m[455]))&~BiasedRNG[454])|((~m[77]&~m[233]&m[455])|(m[77]&~m[233]&m[455])|(m[77]&m[233]&m[455]))):InitCond[706];
    m[312] = run?((((~m[78]&~m[102]&~m[456])|(m[78]&m[102]&~m[456]))&BiasedRNG[455])|(((m[78]&~m[102]&~m[456])|(~m[78]&m[102]&m[456]))&~BiasedRNG[455])|((~m[78]&~m[102]&m[456])|(m[78]&~m[102]&m[456])|(m[78]&m[102]&m[456]))):InitCond[707];
    m[313] = run?((((~m[78]&~m[114]&~m[457])|(m[78]&m[114]&~m[457]))&BiasedRNG[456])|(((m[78]&~m[114]&~m[457])|(~m[78]&m[114]&m[457]))&~BiasedRNG[456])|((~m[78]&~m[114]&m[457])|(m[78]&~m[114]&m[457])|(m[78]&m[114]&m[457]))):InitCond[708];
    m[314] = run?((((~m[78]&~m[126]&~m[458])|(m[78]&m[126]&~m[458]))&BiasedRNG[457])|(((m[78]&~m[126]&~m[458])|(~m[78]&m[126]&m[458]))&~BiasedRNG[457])|((~m[78]&~m[126]&m[458])|(m[78]&~m[126]&m[458])|(m[78]&m[126]&m[458]))):InitCond[709];
    m[315] = run?((((~m[78]&~m[138]&~m[459])|(m[78]&m[138]&~m[459]))&BiasedRNG[458])|(((m[78]&~m[138]&~m[459])|(~m[78]&m[138]&m[459]))&~BiasedRNG[458])|((~m[78]&~m[138]&m[459])|(m[78]&~m[138]&m[459])|(m[78]&m[138]&m[459]))):InitCond[710];
    m[316] = run?((((~m[79]&~m[150]&~m[460])|(m[79]&m[150]&~m[460]))&BiasedRNG[459])|(((m[79]&~m[150]&~m[460])|(~m[79]&m[150]&m[460]))&~BiasedRNG[459])|((~m[79]&~m[150]&m[460])|(m[79]&~m[150]&m[460])|(m[79]&m[150]&m[460]))):InitCond[711];
    m[317] = run?((((~m[79]&~m[162]&~m[461])|(m[79]&m[162]&~m[461]))&BiasedRNG[460])|(((m[79]&~m[162]&~m[461])|(~m[79]&m[162]&m[461]))&~BiasedRNG[460])|((~m[79]&~m[162]&m[461])|(m[79]&~m[162]&m[461])|(m[79]&m[162]&m[461]))):InitCond[712];
    m[318] = run?((((~m[79]&~m[174]&~m[462])|(m[79]&m[174]&~m[462]))&BiasedRNG[461])|(((m[79]&~m[174]&~m[462])|(~m[79]&m[174]&m[462]))&~BiasedRNG[461])|((~m[79]&~m[174]&m[462])|(m[79]&~m[174]&m[462])|(m[79]&m[174]&m[462]))):InitCond[713];
    m[319] = run?((((~m[79]&~m[186]&~m[463])|(m[79]&m[186]&~m[463]))&BiasedRNG[462])|(((m[79]&~m[186]&~m[463])|(~m[79]&m[186]&m[463]))&~BiasedRNG[462])|((~m[79]&~m[186]&m[463])|(m[79]&~m[186]&m[463])|(m[79]&m[186]&m[463]))):InitCond[714];
    m[320] = run?((((~m[80]&~m[198]&~m[464])|(m[80]&m[198]&~m[464]))&BiasedRNG[463])|(((m[80]&~m[198]&~m[464])|(~m[80]&m[198]&m[464]))&~BiasedRNG[463])|((~m[80]&~m[198]&m[464])|(m[80]&~m[198]&m[464])|(m[80]&m[198]&m[464]))):InitCond[715];
    m[321] = run?((((~m[80]&~m[210]&~m[465])|(m[80]&m[210]&~m[465]))&BiasedRNG[464])|(((m[80]&~m[210]&~m[465])|(~m[80]&m[210]&m[465]))&~BiasedRNG[464])|((~m[80]&~m[210]&m[465])|(m[80]&~m[210]&m[465])|(m[80]&m[210]&m[465]))):InitCond[716];
    m[322] = run?((((~m[80]&~m[222]&~m[466])|(m[80]&m[222]&~m[466]))&BiasedRNG[465])|(((m[80]&~m[222]&~m[466])|(~m[80]&m[222]&m[466]))&~BiasedRNG[465])|((~m[80]&~m[222]&m[466])|(m[80]&~m[222]&m[466])|(m[80]&m[222]&m[466]))):InitCond[717];
    m[323] = run?((((~m[80]&~m[234]&~m[467])|(m[80]&m[234]&~m[467]))&BiasedRNG[466])|(((m[80]&~m[234]&~m[467])|(~m[80]&m[234]&m[467]))&~BiasedRNG[466])|((~m[80]&~m[234]&m[467])|(m[80]&~m[234]&m[467])|(m[80]&m[234]&m[467]))):InitCond[718];
    m[324] = run?((((~m[81]&~m[103]&~m[468])|(m[81]&m[103]&~m[468]))&BiasedRNG[467])|(((m[81]&~m[103]&~m[468])|(~m[81]&m[103]&m[468]))&~BiasedRNG[467])|((~m[81]&~m[103]&m[468])|(m[81]&~m[103]&m[468])|(m[81]&m[103]&m[468]))):InitCond[719];
    m[325] = run?((((~m[81]&~m[115]&~m[469])|(m[81]&m[115]&~m[469]))&BiasedRNG[468])|(((m[81]&~m[115]&~m[469])|(~m[81]&m[115]&m[469]))&~BiasedRNG[468])|((~m[81]&~m[115]&m[469])|(m[81]&~m[115]&m[469])|(m[81]&m[115]&m[469]))):InitCond[720];
    m[326] = run?((((~m[81]&~m[127]&~m[470])|(m[81]&m[127]&~m[470]))&BiasedRNG[469])|(((m[81]&~m[127]&~m[470])|(~m[81]&m[127]&m[470]))&~BiasedRNG[469])|((~m[81]&~m[127]&m[470])|(m[81]&~m[127]&m[470])|(m[81]&m[127]&m[470]))):InitCond[721];
    m[327] = run?((((~m[81]&~m[139]&~m[471])|(m[81]&m[139]&~m[471]))&BiasedRNG[470])|(((m[81]&~m[139]&~m[471])|(~m[81]&m[139]&m[471]))&~BiasedRNG[470])|((~m[81]&~m[139]&m[471])|(m[81]&~m[139]&m[471])|(m[81]&m[139]&m[471]))):InitCond[722];
    m[328] = run?((((~m[82]&~m[151]&~m[472])|(m[82]&m[151]&~m[472]))&BiasedRNG[471])|(((m[82]&~m[151]&~m[472])|(~m[82]&m[151]&m[472]))&~BiasedRNG[471])|((~m[82]&~m[151]&m[472])|(m[82]&~m[151]&m[472])|(m[82]&m[151]&m[472]))):InitCond[723];
    m[329] = run?((((~m[82]&~m[163]&~m[473])|(m[82]&m[163]&~m[473]))&BiasedRNG[472])|(((m[82]&~m[163]&~m[473])|(~m[82]&m[163]&m[473]))&~BiasedRNG[472])|((~m[82]&~m[163]&m[473])|(m[82]&~m[163]&m[473])|(m[82]&m[163]&m[473]))):InitCond[724];
    m[330] = run?((((~m[82]&~m[175]&~m[474])|(m[82]&m[175]&~m[474]))&BiasedRNG[473])|(((m[82]&~m[175]&~m[474])|(~m[82]&m[175]&m[474]))&~BiasedRNG[473])|((~m[82]&~m[175]&m[474])|(m[82]&~m[175]&m[474])|(m[82]&m[175]&m[474]))):InitCond[725];
    m[331] = run?((((~m[82]&~m[187]&~m[475])|(m[82]&m[187]&~m[475]))&BiasedRNG[474])|(((m[82]&~m[187]&~m[475])|(~m[82]&m[187]&m[475]))&~BiasedRNG[474])|((~m[82]&~m[187]&m[475])|(m[82]&~m[187]&m[475])|(m[82]&m[187]&m[475]))):InitCond[726];
    m[332] = run?((((~m[83]&~m[199]&~m[476])|(m[83]&m[199]&~m[476]))&BiasedRNG[475])|(((m[83]&~m[199]&~m[476])|(~m[83]&m[199]&m[476]))&~BiasedRNG[475])|((~m[83]&~m[199]&m[476])|(m[83]&~m[199]&m[476])|(m[83]&m[199]&m[476]))):InitCond[727];
    m[333] = run?((((~m[83]&~m[211]&~m[477])|(m[83]&m[211]&~m[477]))&BiasedRNG[476])|(((m[83]&~m[211]&~m[477])|(~m[83]&m[211]&m[477]))&~BiasedRNG[476])|((~m[83]&~m[211]&m[477])|(m[83]&~m[211]&m[477])|(m[83]&m[211]&m[477]))):InitCond[728];
    m[334] = run?((((~m[83]&~m[223]&~m[478])|(m[83]&m[223]&~m[478]))&BiasedRNG[477])|(((m[83]&~m[223]&~m[478])|(~m[83]&m[223]&m[478]))&~BiasedRNG[477])|((~m[83]&~m[223]&m[478])|(m[83]&~m[223]&m[478])|(m[83]&m[223]&m[478]))):InitCond[729];
    m[335] = run?((((~m[83]&~m[235]&~m[479])|(m[83]&m[235]&~m[479]))&BiasedRNG[478])|(((m[83]&~m[235]&~m[479])|(~m[83]&m[235]&m[479]))&~BiasedRNG[478])|((~m[83]&~m[235]&m[479])|(m[83]&~m[235]&m[479])|(m[83]&m[235]&m[479]))):InitCond[730];
    m[336] = run?((((~m[84]&~m[104]&~m[480])|(m[84]&m[104]&~m[480]))&BiasedRNG[479])|(((m[84]&~m[104]&~m[480])|(~m[84]&m[104]&m[480]))&~BiasedRNG[479])|((~m[84]&~m[104]&m[480])|(m[84]&~m[104]&m[480])|(m[84]&m[104]&m[480]))):InitCond[731];
    m[337] = run?((((~m[84]&~m[116]&~m[481])|(m[84]&m[116]&~m[481]))&BiasedRNG[480])|(((m[84]&~m[116]&~m[481])|(~m[84]&m[116]&m[481]))&~BiasedRNG[480])|((~m[84]&~m[116]&m[481])|(m[84]&~m[116]&m[481])|(m[84]&m[116]&m[481]))):InitCond[732];
    m[338] = run?((((~m[84]&~m[128]&~m[482])|(m[84]&m[128]&~m[482]))&BiasedRNG[481])|(((m[84]&~m[128]&~m[482])|(~m[84]&m[128]&m[482]))&~BiasedRNG[481])|((~m[84]&~m[128]&m[482])|(m[84]&~m[128]&m[482])|(m[84]&m[128]&m[482]))):InitCond[733];
    m[339] = run?((((~m[84]&~m[140]&~m[483])|(m[84]&m[140]&~m[483]))&BiasedRNG[482])|(((m[84]&~m[140]&~m[483])|(~m[84]&m[140]&m[483]))&~BiasedRNG[482])|((~m[84]&~m[140]&m[483])|(m[84]&~m[140]&m[483])|(m[84]&m[140]&m[483]))):InitCond[734];
    m[340] = run?((((~m[85]&~m[152]&~m[484])|(m[85]&m[152]&~m[484]))&BiasedRNG[483])|(((m[85]&~m[152]&~m[484])|(~m[85]&m[152]&m[484]))&~BiasedRNG[483])|((~m[85]&~m[152]&m[484])|(m[85]&~m[152]&m[484])|(m[85]&m[152]&m[484]))):InitCond[735];
    m[341] = run?((((~m[85]&~m[164]&~m[485])|(m[85]&m[164]&~m[485]))&BiasedRNG[484])|(((m[85]&~m[164]&~m[485])|(~m[85]&m[164]&m[485]))&~BiasedRNG[484])|((~m[85]&~m[164]&m[485])|(m[85]&~m[164]&m[485])|(m[85]&m[164]&m[485]))):InitCond[736];
    m[342] = run?((((~m[85]&~m[176]&~m[486])|(m[85]&m[176]&~m[486]))&BiasedRNG[485])|(((m[85]&~m[176]&~m[486])|(~m[85]&m[176]&m[486]))&~BiasedRNG[485])|((~m[85]&~m[176]&m[486])|(m[85]&~m[176]&m[486])|(m[85]&m[176]&m[486]))):InitCond[737];
    m[343] = run?((((~m[85]&~m[188]&~m[487])|(m[85]&m[188]&~m[487]))&BiasedRNG[486])|(((m[85]&~m[188]&~m[487])|(~m[85]&m[188]&m[487]))&~BiasedRNG[486])|((~m[85]&~m[188]&m[487])|(m[85]&~m[188]&m[487])|(m[85]&m[188]&m[487]))):InitCond[738];
    m[344] = run?((((~m[86]&~m[200]&~m[488])|(m[86]&m[200]&~m[488]))&BiasedRNG[487])|(((m[86]&~m[200]&~m[488])|(~m[86]&m[200]&m[488]))&~BiasedRNG[487])|((~m[86]&~m[200]&m[488])|(m[86]&~m[200]&m[488])|(m[86]&m[200]&m[488]))):InitCond[739];
    m[345] = run?((((~m[86]&~m[212]&~m[489])|(m[86]&m[212]&~m[489]))&BiasedRNG[488])|(((m[86]&~m[212]&~m[489])|(~m[86]&m[212]&m[489]))&~BiasedRNG[488])|((~m[86]&~m[212]&m[489])|(m[86]&~m[212]&m[489])|(m[86]&m[212]&m[489]))):InitCond[740];
    m[346] = run?((((~m[86]&~m[224]&~m[490])|(m[86]&m[224]&~m[490]))&BiasedRNG[489])|(((m[86]&~m[224]&~m[490])|(~m[86]&m[224]&m[490]))&~BiasedRNG[489])|((~m[86]&~m[224]&m[490])|(m[86]&~m[224]&m[490])|(m[86]&m[224]&m[490]))):InitCond[741];
    m[347] = run?((((~m[86]&~m[236]&~m[491])|(m[86]&m[236]&~m[491]))&BiasedRNG[490])|(((m[86]&~m[236]&~m[491])|(~m[86]&m[236]&m[491]))&~BiasedRNG[490])|((~m[86]&~m[236]&m[491])|(m[86]&~m[236]&m[491])|(m[86]&m[236]&m[491]))):InitCond[742];
    m[348] = run?((((~m[87]&~m[105]&~m[492])|(m[87]&m[105]&~m[492]))&BiasedRNG[491])|(((m[87]&~m[105]&~m[492])|(~m[87]&m[105]&m[492]))&~BiasedRNG[491])|((~m[87]&~m[105]&m[492])|(m[87]&~m[105]&m[492])|(m[87]&m[105]&m[492]))):InitCond[743];
    m[349] = run?((((~m[87]&~m[117]&~m[493])|(m[87]&m[117]&~m[493]))&BiasedRNG[492])|(((m[87]&~m[117]&~m[493])|(~m[87]&m[117]&m[493]))&~BiasedRNG[492])|((~m[87]&~m[117]&m[493])|(m[87]&~m[117]&m[493])|(m[87]&m[117]&m[493]))):InitCond[744];
    m[350] = run?((((~m[87]&~m[129]&~m[494])|(m[87]&m[129]&~m[494]))&BiasedRNG[493])|(((m[87]&~m[129]&~m[494])|(~m[87]&m[129]&m[494]))&~BiasedRNG[493])|((~m[87]&~m[129]&m[494])|(m[87]&~m[129]&m[494])|(m[87]&m[129]&m[494]))):InitCond[745];
    m[351] = run?((((~m[87]&~m[141]&~m[495])|(m[87]&m[141]&~m[495]))&BiasedRNG[494])|(((m[87]&~m[141]&~m[495])|(~m[87]&m[141]&m[495]))&~BiasedRNG[494])|((~m[87]&~m[141]&m[495])|(m[87]&~m[141]&m[495])|(m[87]&m[141]&m[495]))):InitCond[746];
    m[352] = run?((((~m[88]&~m[153]&~m[496])|(m[88]&m[153]&~m[496]))&BiasedRNG[495])|(((m[88]&~m[153]&~m[496])|(~m[88]&m[153]&m[496]))&~BiasedRNG[495])|((~m[88]&~m[153]&m[496])|(m[88]&~m[153]&m[496])|(m[88]&m[153]&m[496]))):InitCond[747];
    m[353] = run?((((~m[88]&~m[165]&~m[497])|(m[88]&m[165]&~m[497]))&BiasedRNG[496])|(((m[88]&~m[165]&~m[497])|(~m[88]&m[165]&m[497]))&~BiasedRNG[496])|((~m[88]&~m[165]&m[497])|(m[88]&~m[165]&m[497])|(m[88]&m[165]&m[497]))):InitCond[748];
    m[354] = run?((((~m[88]&~m[177]&~m[498])|(m[88]&m[177]&~m[498]))&BiasedRNG[497])|(((m[88]&~m[177]&~m[498])|(~m[88]&m[177]&m[498]))&~BiasedRNG[497])|((~m[88]&~m[177]&m[498])|(m[88]&~m[177]&m[498])|(m[88]&m[177]&m[498]))):InitCond[749];
    m[355] = run?((((~m[88]&~m[189]&~m[499])|(m[88]&m[189]&~m[499]))&BiasedRNG[498])|(((m[88]&~m[189]&~m[499])|(~m[88]&m[189]&m[499]))&~BiasedRNG[498])|((~m[88]&~m[189]&m[499])|(m[88]&~m[189]&m[499])|(m[88]&m[189]&m[499]))):InitCond[750];
    m[356] = run?((((~m[89]&~m[201]&~m[500])|(m[89]&m[201]&~m[500]))&BiasedRNG[499])|(((m[89]&~m[201]&~m[500])|(~m[89]&m[201]&m[500]))&~BiasedRNG[499])|((~m[89]&~m[201]&m[500])|(m[89]&~m[201]&m[500])|(m[89]&m[201]&m[500]))):InitCond[751];
    m[357] = run?((((~m[89]&~m[213]&~m[501])|(m[89]&m[213]&~m[501]))&BiasedRNG[500])|(((m[89]&~m[213]&~m[501])|(~m[89]&m[213]&m[501]))&~BiasedRNG[500])|((~m[89]&~m[213]&m[501])|(m[89]&~m[213]&m[501])|(m[89]&m[213]&m[501]))):InitCond[752];
    m[358] = run?((((~m[89]&~m[225]&~m[502])|(m[89]&m[225]&~m[502]))&BiasedRNG[501])|(((m[89]&~m[225]&~m[502])|(~m[89]&m[225]&m[502]))&~BiasedRNG[501])|((~m[89]&~m[225]&m[502])|(m[89]&~m[225]&m[502])|(m[89]&m[225]&m[502]))):InitCond[753];
    m[359] = run?((((~m[89]&~m[237]&~m[503])|(m[89]&m[237]&~m[503]))&BiasedRNG[502])|(((m[89]&~m[237]&~m[503])|(~m[89]&m[237]&m[503]))&~BiasedRNG[502])|((~m[89]&~m[237]&m[503])|(m[89]&~m[237]&m[503])|(m[89]&m[237]&m[503]))):InitCond[754];
    m[360] = run?((((~m[90]&~m[106]&~m[504])|(m[90]&m[106]&~m[504]))&BiasedRNG[503])|(((m[90]&~m[106]&~m[504])|(~m[90]&m[106]&m[504]))&~BiasedRNG[503])|((~m[90]&~m[106]&m[504])|(m[90]&~m[106]&m[504])|(m[90]&m[106]&m[504]))):InitCond[755];
    m[361] = run?((((~m[90]&~m[118]&~m[505])|(m[90]&m[118]&~m[505]))&BiasedRNG[504])|(((m[90]&~m[118]&~m[505])|(~m[90]&m[118]&m[505]))&~BiasedRNG[504])|((~m[90]&~m[118]&m[505])|(m[90]&~m[118]&m[505])|(m[90]&m[118]&m[505]))):InitCond[756];
    m[362] = run?((((~m[90]&~m[130]&~m[506])|(m[90]&m[130]&~m[506]))&BiasedRNG[505])|(((m[90]&~m[130]&~m[506])|(~m[90]&m[130]&m[506]))&~BiasedRNG[505])|((~m[90]&~m[130]&m[506])|(m[90]&~m[130]&m[506])|(m[90]&m[130]&m[506]))):InitCond[757];
    m[363] = run?((((~m[90]&~m[142]&~m[507])|(m[90]&m[142]&~m[507]))&BiasedRNG[506])|(((m[90]&~m[142]&~m[507])|(~m[90]&m[142]&m[507]))&~BiasedRNG[506])|((~m[90]&~m[142]&m[507])|(m[90]&~m[142]&m[507])|(m[90]&m[142]&m[507]))):InitCond[758];
    m[364] = run?((((~m[91]&~m[154]&~m[508])|(m[91]&m[154]&~m[508]))&BiasedRNG[507])|(((m[91]&~m[154]&~m[508])|(~m[91]&m[154]&m[508]))&~BiasedRNG[507])|((~m[91]&~m[154]&m[508])|(m[91]&~m[154]&m[508])|(m[91]&m[154]&m[508]))):InitCond[759];
    m[365] = run?((((~m[91]&~m[166]&~m[509])|(m[91]&m[166]&~m[509]))&BiasedRNG[508])|(((m[91]&~m[166]&~m[509])|(~m[91]&m[166]&m[509]))&~BiasedRNG[508])|((~m[91]&~m[166]&m[509])|(m[91]&~m[166]&m[509])|(m[91]&m[166]&m[509]))):InitCond[760];
    m[366] = run?((((~m[91]&~m[178]&~m[510])|(m[91]&m[178]&~m[510]))&BiasedRNG[509])|(((m[91]&~m[178]&~m[510])|(~m[91]&m[178]&m[510]))&~BiasedRNG[509])|((~m[91]&~m[178]&m[510])|(m[91]&~m[178]&m[510])|(m[91]&m[178]&m[510]))):InitCond[761];
    m[367] = run?((((~m[91]&~m[190]&~m[511])|(m[91]&m[190]&~m[511]))&BiasedRNG[510])|(((m[91]&~m[190]&~m[511])|(~m[91]&m[190]&m[511]))&~BiasedRNG[510])|((~m[91]&~m[190]&m[511])|(m[91]&~m[190]&m[511])|(m[91]&m[190]&m[511]))):InitCond[762];
    m[368] = run?((((~m[92]&~m[202]&~m[512])|(m[92]&m[202]&~m[512]))&BiasedRNG[511])|(((m[92]&~m[202]&~m[512])|(~m[92]&m[202]&m[512]))&~BiasedRNG[511])|((~m[92]&~m[202]&m[512])|(m[92]&~m[202]&m[512])|(m[92]&m[202]&m[512]))):InitCond[763];
    m[369] = run?((((~m[92]&~m[214]&~m[513])|(m[92]&m[214]&~m[513]))&BiasedRNG[512])|(((m[92]&~m[214]&~m[513])|(~m[92]&m[214]&m[513]))&~BiasedRNG[512])|((~m[92]&~m[214]&m[513])|(m[92]&~m[214]&m[513])|(m[92]&m[214]&m[513]))):InitCond[764];
    m[370] = run?((((~m[92]&~m[226]&~m[514])|(m[92]&m[226]&~m[514]))&BiasedRNG[513])|(((m[92]&~m[226]&~m[514])|(~m[92]&m[226]&m[514]))&~BiasedRNG[513])|((~m[92]&~m[226]&m[514])|(m[92]&~m[226]&m[514])|(m[92]&m[226]&m[514]))):InitCond[765];
    m[371] = run?((((~m[92]&~m[238]&~m[515])|(m[92]&m[238]&~m[515]))&BiasedRNG[514])|(((m[92]&~m[238]&~m[515])|(~m[92]&m[238]&m[515]))&~BiasedRNG[514])|((~m[92]&~m[238]&m[515])|(m[92]&~m[238]&m[515])|(m[92]&m[238]&m[515]))):InitCond[766];
    m[372] = run?((((~m[93]&~m[107]&~m[516])|(m[93]&m[107]&~m[516]))&BiasedRNG[515])|(((m[93]&~m[107]&~m[516])|(~m[93]&m[107]&m[516]))&~BiasedRNG[515])|((~m[93]&~m[107]&m[516])|(m[93]&~m[107]&m[516])|(m[93]&m[107]&m[516]))):InitCond[767];
    m[373] = run?((((~m[93]&~m[119]&~m[517])|(m[93]&m[119]&~m[517]))&BiasedRNG[516])|(((m[93]&~m[119]&~m[517])|(~m[93]&m[119]&m[517]))&~BiasedRNG[516])|((~m[93]&~m[119]&m[517])|(m[93]&~m[119]&m[517])|(m[93]&m[119]&m[517]))):InitCond[768];
    m[374] = run?((((~m[93]&~m[131]&~m[518])|(m[93]&m[131]&~m[518]))&BiasedRNG[517])|(((m[93]&~m[131]&~m[518])|(~m[93]&m[131]&m[518]))&~BiasedRNG[517])|((~m[93]&~m[131]&m[518])|(m[93]&~m[131]&m[518])|(m[93]&m[131]&m[518]))):InitCond[769];
    m[375] = run?((((~m[93]&~m[143]&~m[519])|(m[93]&m[143]&~m[519]))&BiasedRNG[518])|(((m[93]&~m[143]&~m[519])|(~m[93]&m[143]&m[519]))&~BiasedRNG[518])|((~m[93]&~m[143]&m[519])|(m[93]&~m[143]&m[519])|(m[93]&m[143]&m[519]))):InitCond[770];
    m[376] = run?((((~m[94]&~m[155]&~m[520])|(m[94]&m[155]&~m[520]))&BiasedRNG[519])|(((m[94]&~m[155]&~m[520])|(~m[94]&m[155]&m[520]))&~BiasedRNG[519])|((~m[94]&~m[155]&m[520])|(m[94]&~m[155]&m[520])|(m[94]&m[155]&m[520]))):InitCond[771];
    m[377] = run?((((~m[94]&~m[167]&~m[521])|(m[94]&m[167]&~m[521]))&BiasedRNG[520])|(((m[94]&~m[167]&~m[521])|(~m[94]&m[167]&m[521]))&~BiasedRNG[520])|((~m[94]&~m[167]&m[521])|(m[94]&~m[167]&m[521])|(m[94]&m[167]&m[521]))):InitCond[772];
    m[378] = run?((((~m[94]&~m[179]&~m[522])|(m[94]&m[179]&~m[522]))&BiasedRNG[521])|(((m[94]&~m[179]&~m[522])|(~m[94]&m[179]&m[522]))&~BiasedRNG[521])|((~m[94]&~m[179]&m[522])|(m[94]&~m[179]&m[522])|(m[94]&m[179]&m[522]))):InitCond[773];
    m[379] = run?((((~m[94]&~m[191]&~m[523])|(m[94]&m[191]&~m[523]))&BiasedRNG[522])|(((m[94]&~m[191]&~m[523])|(~m[94]&m[191]&m[523]))&~BiasedRNG[522])|((~m[94]&~m[191]&m[523])|(m[94]&~m[191]&m[523])|(m[94]&m[191]&m[523]))):InitCond[774];
    m[380] = run?((((~m[95]&~m[203]&~m[524])|(m[95]&m[203]&~m[524]))&BiasedRNG[523])|(((m[95]&~m[203]&~m[524])|(~m[95]&m[203]&m[524]))&~BiasedRNG[523])|((~m[95]&~m[203]&m[524])|(m[95]&~m[203]&m[524])|(m[95]&m[203]&m[524]))):InitCond[775];
    m[381] = run?((((~m[95]&~m[215]&~m[525])|(m[95]&m[215]&~m[525]))&BiasedRNG[524])|(((m[95]&~m[215]&~m[525])|(~m[95]&m[215]&m[525]))&~BiasedRNG[524])|((~m[95]&~m[215]&m[525])|(m[95]&~m[215]&m[525])|(m[95]&m[215]&m[525]))):InitCond[776];
    m[382] = run?((((~m[95]&~m[227]&~m[526])|(m[95]&m[227]&~m[526]))&BiasedRNG[525])|(((m[95]&~m[227]&~m[526])|(~m[95]&m[227]&m[526]))&~BiasedRNG[525])|((~m[95]&~m[227]&m[526])|(m[95]&~m[227]&m[526])|(m[95]&m[227]&m[526]))):InitCond[777];
    m[383] = run?((((~m[95]&~m[239]&~m[527])|(m[95]&m[239]&~m[527]))&BiasedRNG[526])|(((m[95]&~m[239]&~m[527])|(~m[95]&m[239]&m[527]))&~BiasedRNG[526])|((~m[95]&~m[239]&m[527])|(m[95]&~m[239]&m[527])|(m[95]&m[239]&m[527]))):InitCond[778];
    m[529] = run?((((m[396]&~m[528]&~m[530]&~m[531]&~m[532])|(~m[396]&~m[528]&~m[530]&m[531]&~m[532])|(m[396]&m[528]&~m[530]&m[531]&~m[532])|(m[396]&~m[528]&m[530]&m[531]&~m[532])|(~m[396]&m[528]&~m[530]&~m[531]&m[532])|(~m[396]&~m[528]&m[530]&~m[531]&m[532])|(m[396]&m[528]&m[530]&~m[531]&m[532])|(~m[396]&m[528]&m[530]&m[531]&m[532]))&UnbiasedRNG[252])|((m[396]&~m[528]&~m[530]&m[531]&~m[532])|(~m[396]&~m[528]&~m[530]&~m[531]&m[532])|(m[396]&~m[528]&~m[530]&~m[531]&m[532])|(m[396]&m[528]&~m[530]&~m[531]&m[532])|(m[396]&~m[528]&m[530]&~m[531]&m[532])|(~m[396]&~m[528]&~m[530]&m[531]&m[532])|(m[396]&~m[528]&~m[530]&m[531]&m[532])|(~m[396]&m[528]&~m[530]&m[531]&m[532])|(m[396]&m[528]&~m[530]&m[531]&m[532])|(~m[396]&~m[528]&m[530]&m[531]&m[532])|(m[396]&~m[528]&m[530]&m[531]&m[532])|(m[396]&m[528]&m[530]&m[531]&m[532]))):InitCond[779];
    m[534] = run?((((m[397]&~m[533]&~m[535]&~m[536]&~m[537])|(~m[397]&~m[533]&~m[535]&m[536]&~m[537])|(m[397]&m[533]&~m[535]&m[536]&~m[537])|(m[397]&~m[533]&m[535]&m[536]&~m[537])|(~m[397]&m[533]&~m[535]&~m[536]&m[537])|(~m[397]&~m[533]&m[535]&~m[536]&m[537])|(m[397]&m[533]&m[535]&~m[536]&m[537])|(~m[397]&m[533]&m[535]&m[536]&m[537]))&UnbiasedRNG[253])|((m[397]&~m[533]&~m[535]&m[536]&~m[537])|(~m[397]&~m[533]&~m[535]&~m[536]&m[537])|(m[397]&~m[533]&~m[535]&~m[536]&m[537])|(m[397]&m[533]&~m[535]&~m[536]&m[537])|(m[397]&~m[533]&m[535]&~m[536]&m[537])|(~m[397]&~m[533]&~m[535]&m[536]&m[537])|(m[397]&~m[533]&~m[535]&m[536]&m[537])|(~m[397]&m[533]&~m[535]&m[536]&m[537])|(m[397]&m[533]&~m[535]&m[536]&m[537])|(~m[397]&~m[533]&m[535]&m[536]&m[537])|(m[397]&~m[533]&m[535]&m[536]&m[537])|(m[397]&m[533]&m[535]&m[536]&m[537]))):InitCond[780];
    m[539] = run?((((m[408]&~m[538]&~m[540]&~m[541]&~m[542])|(~m[408]&~m[538]&~m[540]&m[541]&~m[542])|(m[408]&m[538]&~m[540]&m[541]&~m[542])|(m[408]&~m[538]&m[540]&m[541]&~m[542])|(~m[408]&m[538]&~m[540]&~m[541]&m[542])|(~m[408]&~m[538]&m[540]&~m[541]&m[542])|(m[408]&m[538]&m[540]&~m[541]&m[542])|(~m[408]&m[538]&m[540]&m[541]&m[542]))&UnbiasedRNG[254])|((m[408]&~m[538]&~m[540]&m[541]&~m[542])|(~m[408]&~m[538]&~m[540]&~m[541]&m[542])|(m[408]&~m[538]&~m[540]&~m[541]&m[542])|(m[408]&m[538]&~m[540]&~m[541]&m[542])|(m[408]&~m[538]&m[540]&~m[541]&m[542])|(~m[408]&~m[538]&~m[540]&m[541]&m[542])|(m[408]&~m[538]&~m[540]&m[541]&m[542])|(~m[408]&m[538]&~m[540]&m[541]&m[542])|(m[408]&m[538]&~m[540]&m[541]&m[542])|(~m[408]&~m[538]&m[540]&m[541]&m[542])|(m[408]&~m[538]&m[540]&m[541]&m[542])|(m[408]&m[538]&m[540]&m[541]&m[542]))):InitCond[781];
    m[544] = run?((((m[398]&~m[543]&~m[545]&~m[546]&~m[547])|(~m[398]&~m[543]&~m[545]&m[546]&~m[547])|(m[398]&m[543]&~m[545]&m[546]&~m[547])|(m[398]&~m[543]&m[545]&m[546]&~m[547])|(~m[398]&m[543]&~m[545]&~m[546]&m[547])|(~m[398]&~m[543]&m[545]&~m[546]&m[547])|(m[398]&m[543]&m[545]&~m[546]&m[547])|(~m[398]&m[543]&m[545]&m[546]&m[547]))&UnbiasedRNG[255])|((m[398]&~m[543]&~m[545]&m[546]&~m[547])|(~m[398]&~m[543]&~m[545]&~m[546]&m[547])|(m[398]&~m[543]&~m[545]&~m[546]&m[547])|(m[398]&m[543]&~m[545]&~m[546]&m[547])|(m[398]&~m[543]&m[545]&~m[546]&m[547])|(~m[398]&~m[543]&~m[545]&m[546]&m[547])|(m[398]&~m[543]&~m[545]&m[546]&m[547])|(~m[398]&m[543]&~m[545]&m[546]&m[547])|(m[398]&m[543]&~m[545]&m[546]&m[547])|(~m[398]&~m[543]&m[545]&m[546]&m[547])|(m[398]&~m[543]&m[545]&m[546]&m[547])|(m[398]&m[543]&m[545]&m[546]&m[547]))):InitCond[782];
    m[549] = run?((((m[409]&~m[548]&~m[550]&~m[551]&~m[552])|(~m[409]&~m[548]&~m[550]&m[551]&~m[552])|(m[409]&m[548]&~m[550]&m[551]&~m[552])|(m[409]&~m[548]&m[550]&m[551]&~m[552])|(~m[409]&m[548]&~m[550]&~m[551]&m[552])|(~m[409]&~m[548]&m[550]&~m[551]&m[552])|(m[409]&m[548]&m[550]&~m[551]&m[552])|(~m[409]&m[548]&m[550]&m[551]&m[552]))&UnbiasedRNG[256])|((m[409]&~m[548]&~m[550]&m[551]&~m[552])|(~m[409]&~m[548]&~m[550]&~m[551]&m[552])|(m[409]&~m[548]&~m[550]&~m[551]&m[552])|(m[409]&m[548]&~m[550]&~m[551]&m[552])|(m[409]&~m[548]&m[550]&~m[551]&m[552])|(~m[409]&~m[548]&~m[550]&m[551]&m[552])|(m[409]&~m[548]&~m[550]&m[551]&m[552])|(~m[409]&m[548]&~m[550]&m[551]&m[552])|(m[409]&m[548]&~m[550]&m[551]&m[552])|(~m[409]&~m[548]&m[550]&m[551]&m[552])|(m[409]&~m[548]&m[550]&m[551]&m[552])|(m[409]&m[548]&m[550]&m[551]&m[552]))):InitCond[783];
    m[554] = run?((((m[420]&~m[553]&~m[555]&~m[556]&~m[557])|(~m[420]&~m[553]&~m[555]&m[556]&~m[557])|(m[420]&m[553]&~m[555]&m[556]&~m[557])|(m[420]&~m[553]&m[555]&m[556]&~m[557])|(~m[420]&m[553]&~m[555]&~m[556]&m[557])|(~m[420]&~m[553]&m[555]&~m[556]&m[557])|(m[420]&m[553]&m[555]&~m[556]&m[557])|(~m[420]&m[553]&m[555]&m[556]&m[557]))&UnbiasedRNG[257])|((m[420]&~m[553]&~m[555]&m[556]&~m[557])|(~m[420]&~m[553]&~m[555]&~m[556]&m[557])|(m[420]&~m[553]&~m[555]&~m[556]&m[557])|(m[420]&m[553]&~m[555]&~m[556]&m[557])|(m[420]&~m[553]&m[555]&~m[556]&m[557])|(~m[420]&~m[553]&~m[555]&m[556]&m[557])|(m[420]&~m[553]&~m[555]&m[556]&m[557])|(~m[420]&m[553]&~m[555]&m[556]&m[557])|(m[420]&m[553]&~m[555]&m[556]&m[557])|(~m[420]&~m[553]&m[555]&m[556]&m[557])|(m[420]&~m[553]&m[555]&m[556]&m[557])|(m[420]&m[553]&m[555]&m[556]&m[557]))):InitCond[784];
    m[559] = run?((((m[399]&~m[558]&~m[560]&~m[561]&~m[562])|(~m[399]&~m[558]&~m[560]&m[561]&~m[562])|(m[399]&m[558]&~m[560]&m[561]&~m[562])|(m[399]&~m[558]&m[560]&m[561]&~m[562])|(~m[399]&m[558]&~m[560]&~m[561]&m[562])|(~m[399]&~m[558]&m[560]&~m[561]&m[562])|(m[399]&m[558]&m[560]&~m[561]&m[562])|(~m[399]&m[558]&m[560]&m[561]&m[562]))&UnbiasedRNG[258])|((m[399]&~m[558]&~m[560]&m[561]&~m[562])|(~m[399]&~m[558]&~m[560]&~m[561]&m[562])|(m[399]&~m[558]&~m[560]&~m[561]&m[562])|(m[399]&m[558]&~m[560]&~m[561]&m[562])|(m[399]&~m[558]&m[560]&~m[561]&m[562])|(~m[399]&~m[558]&~m[560]&m[561]&m[562])|(m[399]&~m[558]&~m[560]&m[561]&m[562])|(~m[399]&m[558]&~m[560]&m[561]&m[562])|(m[399]&m[558]&~m[560]&m[561]&m[562])|(~m[399]&~m[558]&m[560]&m[561]&m[562])|(m[399]&~m[558]&m[560]&m[561]&m[562])|(m[399]&m[558]&m[560]&m[561]&m[562]))):InitCond[785];
    m[564] = run?((((m[410]&~m[563]&~m[565]&~m[566]&~m[567])|(~m[410]&~m[563]&~m[565]&m[566]&~m[567])|(m[410]&m[563]&~m[565]&m[566]&~m[567])|(m[410]&~m[563]&m[565]&m[566]&~m[567])|(~m[410]&m[563]&~m[565]&~m[566]&m[567])|(~m[410]&~m[563]&m[565]&~m[566]&m[567])|(m[410]&m[563]&m[565]&~m[566]&m[567])|(~m[410]&m[563]&m[565]&m[566]&m[567]))&UnbiasedRNG[259])|((m[410]&~m[563]&~m[565]&m[566]&~m[567])|(~m[410]&~m[563]&~m[565]&~m[566]&m[567])|(m[410]&~m[563]&~m[565]&~m[566]&m[567])|(m[410]&m[563]&~m[565]&~m[566]&m[567])|(m[410]&~m[563]&m[565]&~m[566]&m[567])|(~m[410]&~m[563]&~m[565]&m[566]&m[567])|(m[410]&~m[563]&~m[565]&m[566]&m[567])|(~m[410]&m[563]&~m[565]&m[566]&m[567])|(m[410]&m[563]&~m[565]&m[566]&m[567])|(~m[410]&~m[563]&m[565]&m[566]&m[567])|(m[410]&~m[563]&m[565]&m[566]&m[567])|(m[410]&m[563]&m[565]&m[566]&m[567]))):InitCond[786];
    m[569] = run?((((m[421]&~m[568]&~m[570]&~m[571]&~m[572])|(~m[421]&~m[568]&~m[570]&m[571]&~m[572])|(m[421]&m[568]&~m[570]&m[571]&~m[572])|(m[421]&~m[568]&m[570]&m[571]&~m[572])|(~m[421]&m[568]&~m[570]&~m[571]&m[572])|(~m[421]&~m[568]&m[570]&~m[571]&m[572])|(m[421]&m[568]&m[570]&~m[571]&m[572])|(~m[421]&m[568]&m[570]&m[571]&m[572]))&UnbiasedRNG[260])|((m[421]&~m[568]&~m[570]&m[571]&~m[572])|(~m[421]&~m[568]&~m[570]&~m[571]&m[572])|(m[421]&~m[568]&~m[570]&~m[571]&m[572])|(m[421]&m[568]&~m[570]&~m[571]&m[572])|(m[421]&~m[568]&m[570]&~m[571]&m[572])|(~m[421]&~m[568]&~m[570]&m[571]&m[572])|(m[421]&~m[568]&~m[570]&m[571]&m[572])|(~m[421]&m[568]&~m[570]&m[571]&m[572])|(m[421]&m[568]&~m[570]&m[571]&m[572])|(~m[421]&~m[568]&m[570]&m[571]&m[572])|(m[421]&~m[568]&m[570]&m[571]&m[572])|(m[421]&m[568]&m[570]&m[571]&m[572]))):InitCond[787];
    m[574] = run?((((m[432]&~m[573]&~m[575]&~m[576]&~m[577])|(~m[432]&~m[573]&~m[575]&m[576]&~m[577])|(m[432]&m[573]&~m[575]&m[576]&~m[577])|(m[432]&~m[573]&m[575]&m[576]&~m[577])|(~m[432]&m[573]&~m[575]&~m[576]&m[577])|(~m[432]&~m[573]&m[575]&~m[576]&m[577])|(m[432]&m[573]&m[575]&~m[576]&m[577])|(~m[432]&m[573]&m[575]&m[576]&m[577]))&UnbiasedRNG[261])|((m[432]&~m[573]&~m[575]&m[576]&~m[577])|(~m[432]&~m[573]&~m[575]&~m[576]&m[577])|(m[432]&~m[573]&~m[575]&~m[576]&m[577])|(m[432]&m[573]&~m[575]&~m[576]&m[577])|(m[432]&~m[573]&m[575]&~m[576]&m[577])|(~m[432]&~m[573]&~m[575]&m[576]&m[577])|(m[432]&~m[573]&~m[575]&m[576]&m[577])|(~m[432]&m[573]&~m[575]&m[576]&m[577])|(m[432]&m[573]&~m[575]&m[576]&m[577])|(~m[432]&~m[573]&m[575]&m[576]&m[577])|(m[432]&~m[573]&m[575]&m[576]&m[577])|(m[432]&m[573]&m[575]&m[576]&m[577]))):InitCond[788];
    m[579] = run?((((m[400]&~m[578]&~m[580]&~m[581]&~m[582])|(~m[400]&~m[578]&~m[580]&m[581]&~m[582])|(m[400]&m[578]&~m[580]&m[581]&~m[582])|(m[400]&~m[578]&m[580]&m[581]&~m[582])|(~m[400]&m[578]&~m[580]&~m[581]&m[582])|(~m[400]&~m[578]&m[580]&~m[581]&m[582])|(m[400]&m[578]&m[580]&~m[581]&m[582])|(~m[400]&m[578]&m[580]&m[581]&m[582]))&UnbiasedRNG[262])|((m[400]&~m[578]&~m[580]&m[581]&~m[582])|(~m[400]&~m[578]&~m[580]&~m[581]&m[582])|(m[400]&~m[578]&~m[580]&~m[581]&m[582])|(m[400]&m[578]&~m[580]&~m[581]&m[582])|(m[400]&~m[578]&m[580]&~m[581]&m[582])|(~m[400]&~m[578]&~m[580]&m[581]&m[582])|(m[400]&~m[578]&~m[580]&m[581]&m[582])|(~m[400]&m[578]&~m[580]&m[581]&m[582])|(m[400]&m[578]&~m[580]&m[581]&m[582])|(~m[400]&~m[578]&m[580]&m[581]&m[582])|(m[400]&~m[578]&m[580]&m[581]&m[582])|(m[400]&m[578]&m[580]&m[581]&m[582]))):InitCond[789];
    m[584] = run?((((m[411]&~m[583]&~m[585]&~m[586]&~m[587])|(~m[411]&~m[583]&~m[585]&m[586]&~m[587])|(m[411]&m[583]&~m[585]&m[586]&~m[587])|(m[411]&~m[583]&m[585]&m[586]&~m[587])|(~m[411]&m[583]&~m[585]&~m[586]&m[587])|(~m[411]&~m[583]&m[585]&~m[586]&m[587])|(m[411]&m[583]&m[585]&~m[586]&m[587])|(~m[411]&m[583]&m[585]&m[586]&m[587]))&UnbiasedRNG[263])|((m[411]&~m[583]&~m[585]&m[586]&~m[587])|(~m[411]&~m[583]&~m[585]&~m[586]&m[587])|(m[411]&~m[583]&~m[585]&~m[586]&m[587])|(m[411]&m[583]&~m[585]&~m[586]&m[587])|(m[411]&~m[583]&m[585]&~m[586]&m[587])|(~m[411]&~m[583]&~m[585]&m[586]&m[587])|(m[411]&~m[583]&~m[585]&m[586]&m[587])|(~m[411]&m[583]&~m[585]&m[586]&m[587])|(m[411]&m[583]&~m[585]&m[586]&m[587])|(~m[411]&~m[583]&m[585]&m[586]&m[587])|(m[411]&~m[583]&m[585]&m[586]&m[587])|(m[411]&m[583]&m[585]&m[586]&m[587]))):InitCond[790];
    m[589] = run?((((m[422]&~m[588]&~m[590]&~m[591]&~m[592])|(~m[422]&~m[588]&~m[590]&m[591]&~m[592])|(m[422]&m[588]&~m[590]&m[591]&~m[592])|(m[422]&~m[588]&m[590]&m[591]&~m[592])|(~m[422]&m[588]&~m[590]&~m[591]&m[592])|(~m[422]&~m[588]&m[590]&~m[591]&m[592])|(m[422]&m[588]&m[590]&~m[591]&m[592])|(~m[422]&m[588]&m[590]&m[591]&m[592]))&UnbiasedRNG[264])|((m[422]&~m[588]&~m[590]&m[591]&~m[592])|(~m[422]&~m[588]&~m[590]&~m[591]&m[592])|(m[422]&~m[588]&~m[590]&~m[591]&m[592])|(m[422]&m[588]&~m[590]&~m[591]&m[592])|(m[422]&~m[588]&m[590]&~m[591]&m[592])|(~m[422]&~m[588]&~m[590]&m[591]&m[592])|(m[422]&~m[588]&~m[590]&m[591]&m[592])|(~m[422]&m[588]&~m[590]&m[591]&m[592])|(m[422]&m[588]&~m[590]&m[591]&m[592])|(~m[422]&~m[588]&m[590]&m[591]&m[592])|(m[422]&~m[588]&m[590]&m[591]&m[592])|(m[422]&m[588]&m[590]&m[591]&m[592]))):InitCond[791];
    m[594] = run?((((m[433]&~m[593]&~m[595]&~m[596]&~m[597])|(~m[433]&~m[593]&~m[595]&m[596]&~m[597])|(m[433]&m[593]&~m[595]&m[596]&~m[597])|(m[433]&~m[593]&m[595]&m[596]&~m[597])|(~m[433]&m[593]&~m[595]&~m[596]&m[597])|(~m[433]&~m[593]&m[595]&~m[596]&m[597])|(m[433]&m[593]&m[595]&~m[596]&m[597])|(~m[433]&m[593]&m[595]&m[596]&m[597]))&UnbiasedRNG[265])|((m[433]&~m[593]&~m[595]&m[596]&~m[597])|(~m[433]&~m[593]&~m[595]&~m[596]&m[597])|(m[433]&~m[593]&~m[595]&~m[596]&m[597])|(m[433]&m[593]&~m[595]&~m[596]&m[597])|(m[433]&~m[593]&m[595]&~m[596]&m[597])|(~m[433]&~m[593]&~m[595]&m[596]&m[597])|(m[433]&~m[593]&~m[595]&m[596]&m[597])|(~m[433]&m[593]&~m[595]&m[596]&m[597])|(m[433]&m[593]&~m[595]&m[596]&m[597])|(~m[433]&~m[593]&m[595]&m[596]&m[597])|(m[433]&~m[593]&m[595]&m[596]&m[597])|(m[433]&m[593]&m[595]&m[596]&m[597]))):InitCond[792];
    m[599] = run?((((m[444]&~m[598]&~m[600]&~m[601]&~m[602])|(~m[444]&~m[598]&~m[600]&m[601]&~m[602])|(m[444]&m[598]&~m[600]&m[601]&~m[602])|(m[444]&~m[598]&m[600]&m[601]&~m[602])|(~m[444]&m[598]&~m[600]&~m[601]&m[602])|(~m[444]&~m[598]&m[600]&~m[601]&m[602])|(m[444]&m[598]&m[600]&~m[601]&m[602])|(~m[444]&m[598]&m[600]&m[601]&m[602]))&UnbiasedRNG[266])|((m[444]&~m[598]&~m[600]&m[601]&~m[602])|(~m[444]&~m[598]&~m[600]&~m[601]&m[602])|(m[444]&~m[598]&~m[600]&~m[601]&m[602])|(m[444]&m[598]&~m[600]&~m[601]&m[602])|(m[444]&~m[598]&m[600]&~m[601]&m[602])|(~m[444]&~m[598]&~m[600]&m[601]&m[602])|(m[444]&~m[598]&~m[600]&m[601]&m[602])|(~m[444]&m[598]&~m[600]&m[601]&m[602])|(m[444]&m[598]&~m[600]&m[601]&m[602])|(~m[444]&~m[598]&m[600]&m[601]&m[602])|(m[444]&~m[598]&m[600]&m[601]&m[602])|(m[444]&m[598]&m[600]&m[601]&m[602]))):InitCond[793];
    m[604] = run?((((m[401]&~m[603]&~m[605]&~m[606]&~m[607])|(~m[401]&~m[603]&~m[605]&m[606]&~m[607])|(m[401]&m[603]&~m[605]&m[606]&~m[607])|(m[401]&~m[603]&m[605]&m[606]&~m[607])|(~m[401]&m[603]&~m[605]&~m[606]&m[607])|(~m[401]&~m[603]&m[605]&~m[606]&m[607])|(m[401]&m[603]&m[605]&~m[606]&m[607])|(~m[401]&m[603]&m[605]&m[606]&m[607]))&UnbiasedRNG[267])|((m[401]&~m[603]&~m[605]&m[606]&~m[607])|(~m[401]&~m[603]&~m[605]&~m[606]&m[607])|(m[401]&~m[603]&~m[605]&~m[606]&m[607])|(m[401]&m[603]&~m[605]&~m[606]&m[607])|(m[401]&~m[603]&m[605]&~m[606]&m[607])|(~m[401]&~m[603]&~m[605]&m[606]&m[607])|(m[401]&~m[603]&~m[605]&m[606]&m[607])|(~m[401]&m[603]&~m[605]&m[606]&m[607])|(m[401]&m[603]&~m[605]&m[606]&m[607])|(~m[401]&~m[603]&m[605]&m[606]&m[607])|(m[401]&~m[603]&m[605]&m[606]&m[607])|(m[401]&m[603]&m[605]&m[606]&m[607]))):InitCond[794];
    m[609] = run?((((m[412]&~m[608]&~m[610]&~m[611]&~m[612])|(~m[412]&~m[608]&~m[610]&m[611]&~m[612])|(m[412]&m[608]&~m[610]&m[611]&~m[612])|(m[412]&~m[608]&m[610]&m[611]&~m[612])|(~m[412]&m[608]&~m[610]&~m[611]&m[612])|(~m[412]&~m[608]&m[610]&~m[611]&m[612])|(m[412]&m[608]&m[610]&~m[611]&m[612])|(~m[412]&m[608]&m[610]&m[611]&m[612]))&UnbiasedRNG[268])|((m[412]&~m[608]&~m[610]&m[611]&~m[612])|(~m[412]&~m[608]&~m[610]&~m[611]&m[612])|(m[412]&~m[608]&~m[610]&~m[611]&m[612])|(m[412]&m[608]&~m[610]&~m[611]&m[612])|(m[412]&~m[608]&m[610]&~m[611]&m[612])|(~m[412]&~m[608]&~m[610]&m[611]&m[612])|(m[412]&~m[608]&~m[610]&m[611]&m[612])|(~m[412]&m[608]&~m[610]&m[611]&m[612])|(m[412]&m[608]&~m[610]&m[611]&m[612])|(~m[412]&~m[608]&m[610]&m[611]&m[612])|(m[412]&~m[608]&m[610]&m[611]&m[612])|(m[412]&m[608]&m[610]&m[611]&m[612]))):InitCond[795];
    m[614] = run?((((m[423]&~m[613]&~m[615]&~m[616]&~m[617])|(~m[423]&~m[613]&~m[615]&m[616]&~m[617])|(m[423]&m[613]&~m[615]&m[616]&~m[617])|(m[423]&~m[613]&m[615]&m[616]&~m[617])|(~m[423]&m[613]&~m[615]&~m[616]&m[617])|(~m[423]&~m[613]&m[615]&~m[616]&m[617])|(m[423]&m[613]&m[615]&~m[616]&m[617])|(~m[423]&m[613]&m[615]&m[616]&m[617]))&UnbiasedRNG[269])|((m[423]&~m[613]&~m[615]&m[616]&~m[617])|(~m[423]&~m[613]&~m[615]&~m[616]&m[617])|(m[423]&~m[613]&~m[615]&~m[616]&m[617])|(m[423]&m[613]&~m[615]&~m[616]&m[617])|(m[423]&~m[613]&m[615]&~m[616]&m[617])|(~m[423]&~m[613]&~m[615]&m[616]&m[617])|(m[423]&~m[613]&~m[615]&m[616]&m[617])|(~m[423]&m[613]&~m[615]&m[616]&m[617])|(m[423]&m[613]&~m[615]&m[616]&m[617])|(~m[423]&~m[613]&m[615]&m[616]&m[617])|(m[423]&~m[613]&m[615]&m[616]&m[617])|(m[423]&m[613]&m[615]&m[616]&m[617]))):InitCond[796];
    m[619] = run?((((m[434]&~m[618]&~m[620]&~m[621]&~m[622])|(~m[434]&~m[618]&~m[620]&m[621]&~m[622])|(m[434]&m[618]&~m[620]&m[621]&~m[622])|(m[434]&~m[618]&m[620]&m[621]&~m[622])|(~m[434]&m[618]&~m[620]&~m[621]&m[622])|(~m[434]&~m[618]&m[620]&~m[621]&m[622])|(m[434]&m[618]&m[620]&~m[621]&m[622])|(~m[434]&m[618]&m[620]&m[621]&m[622]))&UnbiasedRNG[270])|((m[434]&~m[618]&~m[620]&m[621]&~m[622])|(~m[434]&~m[618]&~m[620]&~m[621]&m[622])|(m[434]&~m[618]&~m[620]&~m[621]&m[622])|(m[434]&m[618]&~m[620]&~m[621]&m[622])|(m[434]&~m[618]&m[620]&~m[621]&m[622])|(~m[434]&~m[618]&~m[620]&m[621]&m[622])|(m[434]&~m[618]&~m[620]&m[621]&m[622])|(~m[434]&m[618]&~m[620]&m[621]&m[622])|(m[434]&m[618]&~m[620]&m[621]&m[622])|(~m[434]&~m[618]&m[620]&m[621]&m[622])|(m[434]&~m[618]&m[620]&m[621]&m[622])|(m[434]&m[618]&m[620]&m[621]&m[622]))):InitCond[797];
    m[624] = run?((((m[445]&~m[623]&~m[625]&~m[626]&~m[627])|(~m[445]&~m[623]&~m[625]&m[626]&~m[627])|(m[445]&m[623]&~m[625]&m[626]&~m[627])|(m[445]&~m[623]&m[625]&m[626]&~m[627])|(~m[445]&m[623]&~m[625]&~m[626]&m[627])|(~m[445]&~m[623]&m[625]&~m[626]&m[627])|(m[445]&m[623]&m[625]&~m[626]&m[627])|(~m[445]&m[623]&m[625]&m[626]&m[627]))&UnbiasedRNG[271])|((m[445]&~m[623]&~m[625]&m[626]&~m[627])|(~m[445]&~m[623]&~m[625]&~m[626]&m[627])|(m[445]&~m[623]&~m[625]&~m[626]&m[627])|(m[445]&m[623]&~m[625]&~m[626]&m[627])|(m[445]&~m[623]&m[625]&~m[626]&m[627])|(~m[445]&~m[623]&~m[625]&m[626]&m[627])|(m[445]&~m[623]&~m[625]&m[626]&m[627])|(~m[445]&m[623]&~m[625]&m[626]&m[627])|(m[445]&m[623]&~m[625]&m[626]&m[627])|(~m[445]&~m[623]&m[625]&m[626]&m[627])|(m[445]&~m[623]&m[625]&m[626]&m[627])|(m[445]&m[623]&m[625]&m[626]&m[627]))):InitCond[798];
    m[629] = run?((((m[456]&~m[628]&~m[630]&~m[631]&~m[632])|(~m[456]&~m[628]&~m[630]&m[631]&~m[632])|(m[456]&m[628]&~m[630]&m[631]&~m[632])|(m[456]&~m[628]&m[630]&m[631]&~m[632])|(~m[456]&m[628]&~m[630]&~m[631]&m[632])|(~m[456]&~m[628]&m[630]&~m[631]&m[632])|(m[456]&m[628]&m[630]&~m[631]&m[632])|(~m[456]&m[628]&m[630]&m[631]&m[632]))&UnbiasedRNG[272])|((m[456]&~m[628]&~m[630]&m[631]&~m[632])|(~m[456]&~m[628]&~m[630]&~m[631]&m[632])|(m[456]&~m[628]&~m[630]&~m[631]&m[632])|(m[456]&m[628]&~m[630]&~m[631]&m[632])|(m[456]&~m[628]&m[630]&~m[631]&m[632])|(~m[456]&~m[628]&~m[630]&m[631]&m[632])|(m[456]&~m[628]&~m[630]&m[631]&m[632])|(~m[456]&m[628]&~m[630]&m[631]&m[632])|(m[456]&m[628]&~m[630]&m[631]&m[632])|(~m[456]&~m[628]&m[630]&m[631]&m[632])|(m[456]&~m[628]&m[630]&m[631]&m[632])|(m[456]&m[628]&m[630]&m[631]&m[632]))):InitCond[799];
    m[634] = run?((((m[402]&~m[633]&~m[635]&~m[636]&~m[637])|(~m[402]&~m[633]&~m[635]&m[636]&~m[637])|(m[402]&m[633]&~m[635]&m[636]&~m[637])|(m[402]&~m[633]&m[635]&m[636]&~m[637])|(~m[402]&m[633]&~m[635]&~m[636]&m[637])|(~m[402]&~m[633]&m[635]&~m[636]&m[637])|(m[402]&m[633]&m[635]&~m[636]&m[637])|(~m[402]&m[633]&m[635]&m[636]&m[637]))&UnbiasedRNG[273])|((m[402]&~m[633]&~m[635]&m[636]&~m[637])|(~m[402]&~m[633]&~m[635]&~m[636]&m[637])|(m[402]&~m[633]&~m[635]&~m[636]&m[637])|(m[402]&m[633]&~m[635]&~m[636]&m[637])|(m[402]&~m[633]&m[635]&~m[636]&m[637])|(~m[402]&~m[633]&~m[635]&m[636]&m[637])|(m[402]&~m[633]&~m[635]&m[636]&m[637])|(~m[402]&m[633]&~m[635]&m[636]&m[637])|(m[402]&m[633]&~m[635]&m[636]&m[637])|(~m[402]&~m[633]&m[635]&m[636]&m[637])|(m[402]&~m[633]&m[635]&m[636]&m[637])|(m[402]&m[633]&m[635]&m[636]&m[637]))):InitCond[800];
    m[639] = run?((((m[413]&~m[638]&~m[640]&~m[641]&~m[642])|(~m[413]&~m[638]&~m[640]&m[641]&~m[642])|(m[413]&m[638]&~m[640]&m[641]&~m[642])|(m[413]&~m[638]&m[640]&m[641]&~m[642])|(~m[413]&m[638]&~m[640]&~m[641]&m[642])|(~m[413]&~m[638]&m[640]&~m[641]&m[642])|(m[413]&m[638]&m[640]&~m[641]&m[642])|(~m[413]&m[638]&m[640]&m[641]&m[642]))&UnbiasedRNG[274])|((m[413]&~m[638]&~m[640]&m[641]&~m[642])|(~m[413]&~m[638]&~m[640]&~m[641]&m[642])|(m[413]&~m[638]&~m[640]&~m[641]&m[642])|(m[413]&m[638]&~m[640]&~m[641]&m[642])|(m[413]&~m[638]&m[640]&~m[641]&m[642])|(~m[413]&~m[638]&~m[640]&m[641]&m[642])|(m[413]&~m[638]&~m[640]&m[641]&m[642])|(~m[413]&m[638]&~m[640]&m[641]&m[642])|(m[413]&m[638]&~m[640]&m[641]&m[642])|(~m[413]&~m[638]&m[640]&m[641]&m[642])|(m[413]&~m[638]&m[640]&m[641]&m[642])|(m[413]&m[638]&m[640]&m[641]&m[642]))):InitCond[801];
    m[644] = run?((((m[424]&~m[643]&~m[645]&~m[646]&~m[647])|(~m[424]&~m[643]&~m[645]&m[646]&~m[647])|(m[424]&m[643]&~m[645]&m[646]&~m[647])|(m[424]&~m[643]&m[645]&m[646]&~m[647])|(~m[424]&m[643]&~m[645]&~m[646]&m[647])|(~m[424]&~m[643]&m[645]&~m[646]&m[647])|(m[424]&m[643]&m[645]&~m[646]&m[647])|(~m[424]&m[643]&m[645]&m[646]&m[647]))&UnbiasedRNG[275])|((m[424]&~m[643]&~m[645]&m[646]&~m[647])|(~m[424]&~m[643]&~m[645]&~m[646]&m[647])|(m[424]&~m[643]&~m[645]&~m[646]&m[647])|(m[424]&m[643]&~m[645]&~m[646]&m[647])|(m[424]&~m[643]&m[645]&~m[646]&m[647])|(~m[424]&~m[643]&~m[645]&m[646]&m[647])|(m[424]&~m[643]&~m[645]&m[646]&m[647])|(~m[424]&m[643]&~m[645]&m[646]&m[647])|(m[424]&m[643]&~m[645]&m[646]&m[647])|(~m[424]&~m[643]&m[645]&m[646]&m[647])|(m[424]&~m[643]&m[645]&m[646]&m[647])|(m[424]&m[643]&m[645]&m[646]&m[647]))):InitCond[802];
    m[649] = run?((((m[435]&~m[648]&~m[650]&~m[651]&~m[652])|(~m[435]&~m[648]&~m[650]&m[651]&~m[652])|(m[435]&m[648]&~m[650]&m[651]&~m[652])|(m[435]&~m[648]&m[650]&m[651]&~m[652])|(~m[435]&m[648]&~m[650]&~m[651]&m[652])|(~m[435]&~m[648]&m[650]&~m[651]&m[652])|(m[435]&m[648]&m[650]&~m[651]&m[652])|(~m[435]&m[648]&m[650]&m[651]&m[652]))&UnbiasedRNG[276])|((m[435]&~m[648]&~m[650]&m[651]&~m[652])|(~m[435]&~m[648]&~m[650]&~m[651]&m[652])|(m[435]&~m[648]&~m[650]&~m[651]&m[652])|(m[435]&m[648]&~m[650]&~m[651]&m[652])|(m[435]&~m[648]&m[650]&~m[651]&m[652])|(~m[435]&~m[648]&~m[650]&m[651]&m[652])|(m[435]&~m[648]&~m[650]&m[651]&m[652])|(~m[435]&m[648]&~m[650]&m[651]&m[652])|(m[435]&m[648]&~m[650]&m[651]&m[652])|(~m[435]&~m[648]&m[650]&m[651]&m[652])|(m[435]&~m[648]&m[650]&m[651]&m[652])|(m[435]&m[648]&m[650]&m[651]&m[652]))):InitCond[803];
    m[654] = run?((((m[446]&~m[653]&~m[655]&~m[656]&~m[657])|(~m[446]&~m[653]&~m[655]&m[656]&~m[657])|(m[446]&m[653]&~m[655]&m[656]&~m[657])|(m[446]&~m[653]&m[655]&m[656]&~m[657])|(~m[446]&m[653]&~m[655]&~m[656]&m[657])|(~m[446]&~m[653]&m[655]&~m[656]&m[657])|(m[446]&m[653]&m[655]&~m[656]&m[657])|(~m[446]&m[653]&m[655]&m[656]&m[657]))&UnbiasedRNG[277])|((m[446]&~m[653]&~m[655]&m[656]&~m[657])|(~m[446]&~m[653]&~m[655]&~m[656]&m[657])|(m[446]&~m[653]&~m[655]&~m[656]&m[657])|(m[446]&m[653]&~m[655]&~m[656]&m[657])|(m[446]&~m[653]&m[655]&~m[656]&m[657])|(~m[446]&~m[653]&~m[655]&m[656]&m[657])|(m[446]&~m[653]&~m[655]&m[656]&m[657])|(~m[446]&m[653]&~m[655]&m[656]&m[657])|(m[446]&m[653]&~m[655]&m[656]&m[657])|(~m[446]&~m[653]&m[655]&m[656]&m[657])|(m[446]&~m[653]&m[655]&m[656]&m[657])|(m[446]&m[653]&m[655]&m[656]&m[657]))):InitCond[804];
    m[659] = run?((((m[457]&~m[658]&~m[660]&~m[661]&~m[662])|(~m[457]&~m[658]&~m[660]&m[661]&~m[662])|(m[457]&m[658]&~m[660]&m[661]&~m[662])|(m[457]&~m[658]&m[660]&m[661]&~m[662])|(~m[457]&m[658]&~m[660]&~m[661]&m[662])|(~m[457]&~m[658]&m[660]&~m[661]&m[662])|(m[457]&m[658]&m[660]&~m[661]&m[662])|(~m[457]&m[658]&m[660]&m[661]&m[662]))&UnbiasedRNG[278])|((m[457]&~m[658]&~m[660]&m[661]&~m[662])|(~m[457]&~m[658]&~m[660]&~m[661]&m[662])|(m[457]&~m[658]&~m[660]&~m[661]&m[662])|(m[457]&m[658]&~m[660]&~m[661]&m[662])|(m[457]&~m[658]&m[660]&~m[661]&m[662])|(~m[457]&~m[658]&~m[660]&m[661]&m[662])|(m[457]&~m[658]&~m[660]&m[661]&m[662])|(~m[457]&m[658]&~m[660]&m[661]&m[662])|(m[457]&m[658]&~m[660]&m[661]&m[662])|(~m[457]&~m[658]&m[660]&m[661]&m[662])|(m[457]&~m[658]&m[660]&m[661]&m[662])|(m[457]&m[658]&m[660]&m[661]&m[662]))):InitCond[805];
    m[664] = run?((((m[468]&~m[663]&~m[665]&~m[666]&~m[667])|(~m[468]&~m[663]&~m[665]&m[666]&~m[667])|(m[468]&m[663]&~m[665]&m[666]&~m[667])|(m[468]&~m[663]&m[665]&m[666]&~m[667])|(~m[468]&m[663]&~m[665]&~m[666]&m[667])|(~m[468]&~m[663]&m[665]&~m[666]&m[667])|(m[468]&m[663]&m[665]&~m[666]&m[667])|(~m[468]&m[663]&m[665]&m[666]&m[667]))&UnbiasedRNG[279])|((m[468]&~m[663]&~m[665]&m[666]&~m[667])|(~m[468]&~m[663]&~m[665]&~m[666]&m[667])|(m[468]&~m[663]&~m[665]&~m[666]&m[667])|(m[468]&m[663]&~m[665]&~m[666]&m[667])|(m[468]&~m[663]&m[665]&~m[666]&m[667])|(~m[468]&~m[663]&~m[665]&m[666]&m[667])|(m[468]&~m[663]&~m[665]&m[666]&m[667])|(~m[468]&m[663]&~m[665]&m[666]&m[667])|(m[468]&m[663]&~m[665]&m[666]&m[667])|(~m[468]&~m[663]&m[665]&m[666]&m[667])|(m[468]&~m[663]&m[665]&m[666]&m[667])|(m[468]&m[663]&m[665]&m[666]&m[667]))):InitCond[806];
    m[669] = run?((((m[403]&~m[668]&~m[670]&~m[671]&~m[672])|(~m[403]&~m[668]&~m[670]&m[671]&~m[672])|(m[403]&m[668]&~m[670]&m[671]&~m[672])|(m[403]&~m[668]&m[670]&m[671]&~m[672])|(~m[403]&m[668]&~m[670]&~m[671]&m[672])|(~m[403]&~m[668]&m[670]&~m[671]&m[672])|(m[403]&m[668]&m[670]&~m[671]&m[672])|(~m[403]&m[668]&m[670]&m[671]&m[672]))&UnbiasedRNG[280])|((m[403]&~m[668]&~m[670]&m[671]&~m[672])|(~m[403]&~m[668]&~m[670]&~m[671]&m[672])|(m[403]&~m[668]&~m[670]&~m[671]&m[672])|(m[403]&m[668]&~m[670]&~m[671]&m[672])|(m[403]&~m[668]&m[670]&~m[671]&m[672])|(~m[403]&~m[668]&~m[670]&m[671]&m[672])|(m[403]&~m[668]&~m[670]&m[671]&m[672])|(~m[403]&m[668]&~m[670]&m[671]&m[672])|(m[403]&m[668]&~m[670]&m[671]&m[672])|(~m[403]&~m[668]&m[670]&m[671]&m[672])|(m[403]&~m[668]&m[670]&m[671]&m[672])|(m[403]&m[668]&m[670]&m[671]&m[672]))):InitCond[807];
    m[674] = run?((((m[414]&~m[673]&~m[675]&~m[676]&~m[677])|(~m[414]&~m[673]&~m[675]&m[676]&~m[677])|(m[414]&m[673]&~m[675]&m[676]&~m[677])|(m[414]&~m[673]&m[675]&m[676]&~m[677])|(~m[414]&m[673]&~m[675]&~m[676]&m[677])|(~m[414]&~m[673]&m[675]&~m[676]&m[677])|(m[414]&m[673]&m[675]&~m[676]&m[677])|(~m[414]&m[673]&m[675]&m[676]&m[677]))&UnbiasedRNG[281])|((m[414]&~m[673]&~m[675]&m[676]&~m[677])|(~m[414]&~m[673]&~m[675]&~m[676]&m[677])|(m[414]&~m[673]&~m[675]&~m[676]&m[677])|(m[414]&m[673]&~m[675]&~m[676]&m[677])|(m[414]&~m[673]&m[675]&~m[676]&m[677])|(~m[414]&~m[673]&~m[675]&m[676]&m[677])|(m[414]&~m[673]&~m[675]&m[676]&m[677])|(~m[414]&m[673]&~m[675]&m[676]&m[677])|(m[414]&m[673]&~m[675]&m[676]&m[677])|(~m[414]&~m[673]&m[675]&m[676]&m[677])|(m[414]&~m[673]&m[675]&m[676]&m[677])|(m[414]&m[673]&m[675]&m[676]&m[677]))):InitCond[808];
    m[679] = run?((((m[425]&~m[678]&~m[680]&~m[681]&~m[682])|(~m[425]&~m[678]&~m[680]&m[681]&~m[682])|(m[425]&m[678]&~m[680]&m[681]&~m[682])|(m[425]&~m[678]&m[680]&m[681]&~m[682])|(~m[425]&m[678]&~m[680]&~m[681]&m[682])|(~m[425]&~m[678]&m[680]&~m[681]&m[682])|(m[425]&m[678]&m[680]&~m[681]&m[682])|(~m[425]&m[678]&m[680]&m[681]&m[682]))&UnbiasedRNG[282])|((m[425]&~m[678]&~m[680]&m[681]&~m[682])|(~m[425]&~m[678]&~m[680]&~m[681]&m[682])|(m[425]&~m[678]&~m[680]&~m[681]&m[682])|(m[425]&m[678]&~m[680]&~m[681]&m[682])|(m[425]&~m[678]&m[680]&~m[681]&m[682])|(~m[425]&~m[678]&~m[680]&m[681]&m[682])|(m[425]&~m[678]&~m[680]&m[681]&m[682])|(~m[425]&m[678]&~m[680]&m[681]&m[682])|(m[425]&m[678]&~m[680]&m[681]&m[682])|(~m[425]&~m[678]&m[680]&m[681]&m[682])|(m[425]&~m[678]&m[680]&m[681]&m[682])|(m[425]&m[678]&m[680]&m[681]&m[682]))):InitCond[809];
    m[684] = run?((((m[436]&~m[683]&~m[685]&~m[686]&~m[687])|(~m[436]&~m[683]&~m[685]&m[686]&~m[687])|(m[436]&m[683]&~m[685]&m[686]&~m[687])|(m[436]&~m[683]&m[685]&m[686]&~m[687])|(~m[436]&m[683]&~m[685]&~m[686]&m[687])|(~m[436]&~m[683]&m[685]&~m[686]&m[687])|(m[436]&m[683]&m[685]&~m[686]&m[687])|(~m[436]&m[683]&m[685]&m[686]&m[687]))&UnbiasedRNG[283])|((m[436]&~m[683]&~m[685]&m[686]&~m[687])|(~m[436]&~m[683]&~m[685]&~m[686]&m[687])|(m[436]&~m[683]&~m[685]&~m[686]&m[687])|(m[436]&m[683]&~m[685]&~m[686]&m[687])|(m[436]&~m[683]&m[685]&~m[686]&m[687])|(~m[436]&~m[683]&~m[685]&m[686]&m[687])|(m[436]&~m[683]&~m[685]&m[686]&m[687])|(~m[436]&m[683]&~m[685]&m[686]&m[687])|(m[436]&m[683]&~m[685]&m[686]&m[687])|(~m[436]&~m[683]&m[685]&m[686]&m[687])|(m[436]&~m[683]&m[685]&m[686]&m[687])|(m[436]&m[683]&m[685]&m[686]&m[687]))):InitCond[810];
    m[689] = run?((((m[447]&~m[688]&~m[690]&~m[691]&~m[692])|(~m[447]&~m[688]&~m[690]&m[691]&~m[692])|(m[447]&m[688]&~m[690]&m[691]&~m[692])|(m[447]&~m[688]&m[690]&m[691]&~m[692])|(~m[447]&m[688]&~m[690]&~m[691]&m[692])|(~m[447]&~m[688]&m[690]&~m[691]&m[692])|(m[447]&m[688]&m[690]&~m[691]&m[692])|(~m[447]&m[688]&m[690]&m[691]&m[692]))&UnbiasedRNG[284])|((m[447]&~m[688]&~m[690]&m[691]&~m[692])|(~m[447]&~m[688]&~m[690]&~m[691]&m[692])|(m[447]&~m[688]&~m[690]&~m[691]&m[692])|(m[447]&m[688]&~m[690]&~m[691]&m[692])|(m[447]&~m[688]&m[690]&~m[691]&m[692])|(~m[447]&~m[688]&~m[690]&m[691]&m[692])|(m[447]&~m[688]&~m[690]&m[691]&m[692])|(~m[447]&m[688]&~m[690]&m[691]&m[692])|(m[447]&m[688]&~m[690]&m[691]&m[692])|(~m[447]&~m[688]&m[690]&m[691]&m[692])|(m[447]&~m[688]&m[690]&m[691]&m[692])|(m[447]&m[688]&m[690]&m[691]&m[692]))):InitCond[811];
    m[694] = run?((((m[458]&~m[693]&~m[695]&~m[696]&~m[697])|(~m[458]&~m[693]&~m[695]&m[696]&~m[697])|(m[458]&m[693]&~m[695]&m[696]&~m[697])|(m[458]&~m[693]&m[695]&m[696]&~m[697])|(~m[458]&m[693]&~m[695]&~m[696]&m[697])|(~m[458]&~m[693]&m[695]&~m[696]&m[697])|(m[458]&m[693]&m[695]&~m[696]&m[697])|(~m[458]&m[693]&m[695]&m[696]&m[697]))&UnbiasedRNG[285])|((m[458]&~m[693]&~m[695]&m[696]&~m[697])|(~m[458]&~m[693]&~m[695]&~m[696]&m[697])|(m[458]&~m[693]&~m[695]&~m[696]&m[697])|(m[458]&m[693]&~m[695]&~m[696]&m[697])|(m[458]&~m[693]&m[695]&~m[696]&m[697])|(~m[458]&~m[693]&~m[695]&m[696]&m[697])|(m[458]&~m[693]&~m[695]&m[696]&m[697])|(~m[458]&m[693]&~m[695]&m[696]&m[697])|(m[458]&m[693]&~m[695]&m[696]&m[697])|(~m[458]&~m[693]&m[695]&m[696]&m[697])|(m[458]&~m[693]&m[695]&m[696]&m[697])|(m[458]&m[693]&m[695]&m[696]&m[697]))):InitCond[812];
    m[699] = run?((((m[469]&~m[698]&~m[700]&~m[701]&~m[702])|(~m[469]&~m[698]&~m[700]&m[701]&~m[702])|(m[469]&m[698]&~m[700]&m[701]&~m[702])|(m[469]&~m[698]&m[700]&m[701]&~m[702])|(~m[469]&m[698]&~m[700]&~m[701]&m[702])|(~m[469]&~m[698]&m[700]&~m[701]&m[702])|(m[469]&m[698]&m[700]&~m[701]&m[702])|(~m[469]&m[698]&m[700]&m[701]&m[702]))&UnbiasedRNG[286])|((m[469]&~m[698]&~m[700]&m[701]&~m[702])|(~m[469]&~m[698]&~m[700]&~m[701]&m[702])|(m[469]&~m[698]&~m[700]&~m[701]&m[702])|(m[469]&m[698]&~m[700]&~m[701]&m[702])|(m[469]&~m[698]&m[700]&~m[701]&m[702])|(~m[469]&~m[698]&~m[700]&m[701]&m[702])|(m[469]&~m[698]&~m[700]&m[701]&m[702])|(~m[469]&m[698]&~m[700]&m[701]&m[702])|(m[469]&m[698]&~m[700]&m[701]&m[702])|(~m[469]&~m[698]&m[700]&m[701]&m[702])|(m[469]&~m[698]&m[700]&m[701]&m[702])|(m[469]&m[698]&m[700]&m[701]&m[702]))):InitCond[813];
    m[704] = run?((((m[480]&~m[703]&~m[705]&~m[706]&~m[707])|(~m[480]&~m[703]&~m[705]&m[706]&~m[707])|(m[480]&m[703]&~m[705]&m[706]&~m[707])|(m[480]&~m[703]&m[705]&m[706]&~m[707])|(~m[480]&m[703]&~m[705]&~m[706]&m[707])|(~m[480]&~m[703]&m[705]&~m[706]&m[707])|(m[480]&m[703]&m[705]&~m[706]&m[707])|(~m[480]&m[703]&m[705]&m[706]&m[707]))&UnbiasedRNG[287])|((m[480]&~m[703]&~m[705]&m[706]&~m[707])|(~m[480]&~m[703]&~m[705]&~m[706]&m[707])|(m[480]&~m[703]&~m[705]&~m[706]&m[707])|(m[480]&m[703]&~m[705]&~m[706]&m[707])|(m[480]&~m[703]&m[705]&~m[706]&m[707])|(~m[480]&~m[703]&~m[705]&m[706]&m[707])|(m[480]&~m[703]&~m[705]&m[706]&m[707])|(~m[480]&m[703]&~m[705]&m[706]&m[707])|(m[480]&m[703]&~m[705]&m[706]&m[707])|(~m[480]&~m[703]&m[705]&m[706]&m[707])|(m[480]&~m[703]&m[705]&m[706]&m[707])|(m[480]&m[703]&m[705]&m[706]&m[707]))):InitCond[814];
    m[709] = run?((((m[404]&~m[708]&~m[710]&~m[711]&~m[712])|(~m[404]&~m[708]&~m[710]&m[711]&~m[712])|(m[404]&m[708]&~m[710]&m[711]&~m[712])|(m[404]&~m[708]&m[710]&m[711]&~m[712])|(~m[404]&m[708]&~m[710]&~m[711]&m[712])|(~m[404]&~m[708]&m[710]&~m[711]&m[712])|(m[404]&m[708]&m[710]&~m[711]&m[712])|(~m[404]&m[708]&m[710]&m[711]&m[712]))&UnbiasedRNG[288])|((m[404]&~m[708]&~m[710]&m[711]&~m[712])|(~m[404]&~m[708]&~m[710]&~m[711]&m[712])|(m[404]&~m[708]&~m[710]&~m[711]&m[712])|(m[404]&m[708]&~m[710]&~m[711]&m[712])|(m[404]&~m[708]&m[710]&~m[711]&m[712])|(~m[404]&~m[708]&~m[710]&m[711]&m[712])|(m[404]&~m[708]&~m[710]&m[711]&m[712])|(~m[404]&m[708]&~m[710]&m[711]&m[712])|(m[404]&m[708]&~m[710]&m[711]&m[712])|(~m[404]&~m[708]&m[710]&m[711]&m[712])|(m[404]&~m[708]&m[710]&m[711]&m[712])|(m[404]&m[708]&m[710]&m[711]&m[712]))):InitCond[815];
    m[714] = run?((((m[415]&~m[713]&~m[715]&~m[716]&~m[717])|(~m[415]&~m[713]&~m[715]&m[716]&~m[717])|(m[415]&m[713]&~m[715]&m[716]&~m[717])|(m[415]&~m[713]&m[715]&m[716]&~m[717])|(~m[415]&m[713]&~m[715]&~m[716]&m[717])|(~m[415]&~m[713]&m[715]&~m[716]&m[717])|(m[415]&m[713]&m[715]&~m[716]&m[717])|(~m[415]&m[713]&m[715]&m[716]&m[717]))&UnbiasedRNG[289])|((m[415]&~m[713]&~m[715]&m[716]&~m[717])|(~m[415]&~m[713]&~m[715]&~m[716]&m[717])|(m[415]&~m[713]&~m[715]&~m[716]&m[717])|(m[415]&m[713]&~m[715]&~m[716]&m[717])|(m[415]&~m[713]&m[715]&~m[716]&m[717])|(~m[415]&~m[713]&~m[715]&m[716]&m[717])|(m[415]&~m[713]&~m[715]&m[716]&m[717])|(~m[415]&m[713]&~m[715]&m[716]&m[717])|(m[415]&m[713]&~m[715]&m[716]&m[717])|(~m[415]&~m[713]&m[715]&m[716]&m[717])|(m[415]&~m[713]&m[715]&m[716]&m[717])|(m[415]&m[713]&m[715]&m[716]&m[717]))):InitCond[816];
    m[719] = run?((((m[426]&~m[718]&~m[720]&~m[721]&~m[722])|(~m[426]&~m[718]&~m[720]&m[721]&~m[722])|(m[426]&m[718]&~m[720]&m[721]&~m[722])|(m[426]&~m[718]&m[720]&m[721]&~m[722])|(~m[426]&m[718]&~m[720]&~m[721]&m[722])|(~m[426]&~m[718]&m[720]&~m[721]&m[722])|(m[426]&m[718]&m[720]&~m[721]&m[722])|(~m[426]&m[718]&m[720]&m[721]&m[722]))&UnbiasedRNG[290])|((m[426]&~m[718]&~m[720]&m[721]&~m[722])|(~m[426]&~m[718]&~m[720]&~m[721]&m[722])|(m[426]&~m[718]&~m[720]&~m[721]&m[722])|(m[426]&m[718]&~m[720]&~m[721]&m[722])|(m[426]&~m[718]&m[720]&~m[721]&m[722])|(~m[426]&~m[718]&~m[720]&m[721]&m[722])|(m[426]&~m[718]&~m[720]&m[721]&m[722])|(~m[426]&m[718]&~m[720]&m[721]&m[722])|(m[426]&m[718]&~m[720]&m[721]&m[722])|(~m[426]&~m[718]&m[720]&m[721]&m[722])|(m[426]&~m[718]&m[720]&m[721]&m[722])|(m[426]&m[718]&m[720]&m[721]&m[722]))):InitCond[817];
    m[724] = run?((((m[437]&~m[723]&~m[725]&~m[726]&~m[727])|(~m[437]&~m[723]&~m[725]&m[726]&~m[727])|(m[437]&m[723]&~m[725]&m[726]&~m[727])|(m[437]&~m[723]&m[725]&m[726]&~m[727])|(~m[437]&m[723]&~m[725]&~m[726]&m[727])|(~m[437]&~m[723]&m[725]&~m[726]&m[727])|(m[437]&m[723]&m[725]&~m[726]&m[727])|(~m[437]&m[723]&m[725]&m[726]&m[727]))&UnbiasedRNG[291])|((m[437]&~m[723]&~m[725]&m[726]&~m[727])|(~m[437]&~m[723]&~m[725]&~m[726]&m[727])|(m[437]&~m[723]&~m[725]&~m[726]&m[727])|(m[437]&m[723]&~m[725]&~m[726]&m[727])|(m[437]&~m[723]&m[725]&~m[726]&m[727])|(~m[437]&~m[723]&~m[725]&m[726]&m[727])|(m[437]&~m[723]&~m[725]&m[726]&m[727])|(~m[437]&m[723]&~m[725]&m[726]&m[727])|(m[437]&m[723]&~m[725]&m[726]&m[727])|(~m[437]&~m[723]&m[725]&m[726]&m[727])|(m[437]&~m[723]&m[725]&m[726]&m[727])|(m[437]&m[723]&m[725]&m[726]&m[727]))):InitCond[818];
    m[729] = run?((((m[448]&~m[728]&~m[730]&~m[731]&~m[732])|(~m[448]&~m[728]&~m[730]&m[731]&~m[732])|(m[448]&m[728]&~m[730]&m[731]&~m[732])|(m[448]&~m[728]&m[730]&m[731]&~m[732])|(~m[448]&m[728]&~m[730]&~m[731]&m[732])|(~m[448]&~m[728]&m[730]&~m[731]&m[732])|(m[448]&m[728]&m[730]&~m[731]&m[732])|(~m[448]&m[728]&m[730]&m[731]&m[732]))&UnbiasedRNG[292])|((m[448]&~m[728]&~m[730]&m[731]&~m[732])|(~m[448]&~m[728]&~m[730]&~m[731]&m[732])|(m[448]&~m[728]&~m[730]&~m[731]&m[732])|(m[448]&m[728]&~m[730]&~m[731]&m[732])|(m[448]&~m[728]&m[730]&~m[731]&m[732])|(~m[448]&~m[728]&~m[730]&m[731]&m[732])|(m[448]&~m[728]&~m[730]&m[731]&m[732])|(~m[448]&m[728]&~m[730]&m[731]&m[732])|(m[448]&m[728]&~m[730]&m[731]&m[732])|(~m[448]&~m[728]&m[730]&m[731]&m[732])|(m[448]&~m[728]&m[730]&m[731]&m[732])|(m[448]&m[728]&m[730]&m[731]&m[732]))):InitCond[819];
    m[734] = run?((((m[459]&~m[733]&~m[735]&~m[736]&~m[737])|(~m[459]&~m[733]&~m[735]&m[736]&~m[737])|(m[459]&m[733]&~m[735]&m[736]&~m[737])|(m[459]&~m[733]&m[735]&m[736]&~m[737])|(~m[459]&m[733]&~m[735]&~m[736]&m[737])|(~m[459]&~m[733]&m[735]&~m[736]&m[737])|(m[459]&m[733]&m[735]&~m[736]&m[737])|(~m[459]&m[733]&m[735]&m[736]&m[737]))&UnbiasedRNG[293])|((m[459]&~m[733]&~m[735]&m[736]&~m[737])|(~m[459]&~m[733]&~m[735]&~m[736]&m[737])|(m[459]&~m[733]&~m[735]&~m[736]&m[737])|(m[459]&m[733]&~m[735]&~m[736]&m[737])|(m[459]&~m[733]&m[735]&~m[736]&m[737])|(~m[459]&~m[733]&~m[735]&m[736]&m[737])|(m[459]&~m[733]&~m[735]&m[736]&m[737])|(~m[459]&m[733]&~m[735]&m[736]&m[737])|(m[459]&m[733]&~m[735]&m[736]&m[737])|(~m[459]&~m[733]&m[735]&m[736]&m[737])|(m[459]&~m[733]&m[735]&m[736]&m[737])|(m[459]&m[733]&m[735]&m[736]&m[737]))):InitCond[820];
    m[739] = run?((((m[470]&~m[738]&~m[740]&~m[741]&~m[742])|(~m[470]&~m[738]&~m[740]&m[741]&~m[742])|(m[470]&m[738]&~m[740]&m[741]&~m[742])|(m[470]&~m[738]&m[740]&m[741]&~m[742])|(~m[470]&m[738]&~m[740]&~m[741]&m[742])|(~m[470]&~m[738]&m[740]&~m[741]&m[742])|(m[470]&m[738]&m[740]&~m[741]&m[742])|(~m[470]&m[738]&m[740]&m[741]&m[742]))&UnbiasedRNG[294])|((m[470]&~m[738]&~m[740]&m[741]&~m[742])|(~m[470]&~m[738]&~m[740]&~m[741]&m[742])|(m[470]&~m[738]&~m[740]&~m[741]&m[742])|(m[470]&m[738]&~m[740]&~m[741]&m[742])|(m[470]&~m[738]&m[740]&~m[741]&m[742])|(~m[470]&~m[738]&~m[740]&m[741]&m[742])|(m[470]&~m[738]&~m[740]&m[741]&m[742])|(~m[470]&m[738]&~m[740]&m[741]&m[742])|(m[470]&m[738]&~m[740]&m[741]&m[742])|(~m[470]&~m[738]&m[740]&m[741]&m[742])|(m[470]&~m[738]&m[740]&m[741]&m[742])|(m[470]&m[738]&m[740]&m[741]&m[742]))):InitCond[821];
    m[744] = run?((((m[481]&~m[743]&~m[745]&~m[746]&~m[747])|(~m[481]&~m[743]&~m[745]&m[746]&~m[747])|(m[481]&m[743]&~m[745]&m[746]&~m[747])|(m[481]&~m[743]&m[745]&m[746]&~m[747])|(~m[481]&m[743]&~m[745]&~m[746]&m[747])|(~m[481]&~m[743]&m[745]&~m[746]&m[747])|(m[481]&m[743]&m[745]&~m[746]&m[747])|(~m[481]&m[743]&m[745]&m[746]&m[747]))&UnbiasedRNG[295])|((m[481]&~m[743]&~m[745]&m[746]&~m[747])|(~m[481]&~m[743]&~m[745]&~m[746]&m[747])|(m[481]&~m[743]&~m[745]&~m[746]&m[747])|(m[481]&m[743]&~m[745]&~m[746]&m[747])|(m[481]&~m[743]&m[745]&~m[746]&m[747])|(~m[481]&~m[743]&~m[745]&m[746]&m[747])|(m[481]&~m[743]&~m[745]&m[746]&m[747])|(~m[481]&m[743]&~m[745]&m[746]&m[747])|(m[481]&m[743]&~m[745]&m[746]&m[747])|(~m[481]&~m[743]&m[745]&m[746]&m[747])|(m[481]&~m[743]&m[745]&m[746]&m[747])|(m[481]&m[743]&m[745]&m[746]&m[747]))):InitCond[822];
    m[749] = run?((((m[492]&~m[748]&~m[750]&~m[751]&~m[752])|(~m[492]&~m[748]&~m[750]&m[751]&~m[752])|(m[492]&m[748]&~m[750]&m[751]&~m[752])|(m[492]&~m[748]&m[750]&m[751]&~m[752])|(~m[492]&m[748]&~m[750]&~m[751]&m[752])|(~m[492]&~m[748]&m[750]&~m[751]&m[752])|(m[492]&m[748]&m[750]&~m[751]&m[752])|(~m[492]&m[748]&m[750]&m[751]&m[752]))&UnbiasedRNG[296])|((m[492]&~m[748]&~m[750]&m[751]&~m[752])|(~m[492]&~m[748]&~m[750]&~m[751]&m[752])|(m[492]&~m[748]&~m[750]&~m[751]&m[752])|(m[492]&m[748]&~m[750]&~m[751]&m[752])|(m[492]&~m[748]&m[750]&~m[751]&m[752])|(~m[492]&~m[748]&~m[750]&m[751]&m[752])|(m[492]&~m[748]&~m[750]&m[751]&m[752])|(~m[492]&m[748]&~m[750]&m[751]&m[752])|(m[492]&m[748]&~m[750]&m[751]&m[752])|(~m[492]&~m[748]&m[750]&m[751]&m[752])|(m[492]&~m[748]&m[750]&m[751]&m[752])|(m[492]&m[748]&m[750]&m[751]&m[752]))):InitCond[823];
    m[754] = run?((((m[405]&~m[753]&~m[755]&~m[756]&~m[757])|(~m[405]&~m[753]&~m[755]&m[756]&~m[757])|(m[405]&m[753]&~m[755]&m[756]&~m[757])|(m[405]&~m[753]&m[755]&m[756]&~m[757])|(~m[405]&m[753]&~m[755]&~m[756]&m[757])|(~m[405]&~m[753]&m[755]&~m[756]&m[757])|(m[405]&m[753]&m[755]&~m[756]&m[757])|(~m[405]&m[753]&m[755]&m[756]&m[757]))&UnbiasedRNG[297])|((m[405]&~m[753]&~m[755]&m[756]&~m[757])|(~m[405]&~m[753]&~m[755]&~m[756]&m[757])|(m[405]&~m[753]&~m[755]&~m[756]&m[757])|(m[405]&m[753]&~m[755]&~m[756]&m[757])|(m[405]&~m[753]&m[755]&~m[756]&m[757])|(~m[405]&~m[753]&~m[755]&m[756]&m[757])|(m[405]&~m[753]&~m[755]&m[756]&m[757])|(~m[405]&m[753]&~m[755]&m[756]&m[757])|(m[405]&m[753]&~m[755]&m[756]&m[757])|(~m[405]&~m[753]&m[755]&m[756]&m[757])|(m[405]&~m[753]&m[755]&m[756]&m[757])|(m[405]&m[753]&m[755]&m[756]&m[757]))):InitCond[824];
    m[759] = run?((((m[416]&~m[758]&~m[760]&~m[761]&~m[762])|(~m[416]&~m[758]&~m[760]&m[761]&~m[762])|(m[416]&m[758]&~m[760]&m[761]&~m[762])|(m[416]&~m[758]&m[760]&m[761]&~m[762])|(~m[416]&m[758]&~m[760]&~m[761]&m[762])|(~m[416]&~m[758]&m[760]&~m[761]&m[762])|(m[416]&m[758]&m[760]&~m[761]&m[762])|(~m[416]&m[758]&m[760]&m[761]&m[762]))&UnbiasedRNG[298])|((m[416]&~m[758]&~m[760]&m[761]&~m[762])|(~m[416]&~m[758]&~m[760]&~m[761]&m[762])|(m[416]&~m[758]&~m[760]&~m[761]&m[762])|(m[416]&m[758]&~m[760]&~m[761]&m[762])|(m[416]&~m[758]&m[760]&~m[761]&m[762])|(~m[416]&~m[758]&~m[760]&m[761]&m[762])|(m[416]&~m[758]&~m[760]&m[761]&m[762])|(~m[416]&m[758]&~m[760]&m[761]&m[762])|(m[416]&m[758]&~m[760]&m[761]&m[762])|(~m[416]&~m[758]&m[760]&m[761]&m[762])|(m[416]&~m[758]&m[760]&m[761]&m[762])|(m[416]&m[758]&m[760]&m[761]&m[762]))):InitCond[825];
    m[764] = run?((((m[427]&~m[763]&~m[765]&~m[766]&~m[767])|(~m[427]&~m[763]&~m[765]&m[766]&~m[767])|(m[427]&m[763]&~m[765]&m[766]&~m[767])|(m[427]&~m[763]&m[765]&m[766]&~m[767])|(~m[427]&m[763]&~m[765]&~m[766]&m[767])|(~m[427]&~m[763]&m[765]&~m[766]&m[767])|(m[427]&m[763]&m[765]&~m[766]&m[767])|(~m[427]&m[763]&m[765]&m[766]&m[767]))&UnbiasedRNG[299])|((m[427]&~m[763]&~m[765]&m[766]&~m[767])|(~m[427]&~m[763]&~m[765]&~m[766]&m[767])|(m[427]&~m[763]&~m[765]&~m[766]&m[767])|(m[427]&m[763]&~m[765]&~m[766]&m[767])|(m[427]&~m[763]&m[765]&~m[766]&m[767])|(~m[427]&~m[763]&~m[765]&m[766]&m[767])|(m[427]&~m[763]&~m[765]&m[766]&m[767])|(~m[427]&m[763]&~m[765]&m[766]&m[767])|(m[427]&m[763]&~m[765]&m[766]&m[767])|(~m[427]&~m[763]&m[765]&m[766]&m[767])|(m[427]&~m[763]&m[765]&m[766]&m[767])|(m[427]&m[763]&m[765]&m[766]&m[767]))):InitCond[826];
    m[769] = run?((((m[438]&~m[768]&~m[770]&~m[771]&~m[772])|(~m[438]&~m[768]&~m[770]&m[771]&~m[772])|(m[438]&m[768]&~m[770]&m[771]&~m[772])|(m[438]&~m[768]&m[770]&m[771]&~m[772])|(~m[438]&m[768]&~m[770]&~m[771]&m[772])|(~m[438]&~m[768]&m[770]&~m[771]&m[772])|(m[438]&m[768]&m[770]&~m[771]&m[772])|(~m[438]&m[768]&m[770]&m[771]&m[772]))&UnbiasedRNG[300])|((m[438]&~m[768]&~m[770]&m[771]&~m[772])|(~m[438]&~m[768]&~m[770]&~m[771]&m[772])|(m[438]&~m[768]&~m[770]&~m[771]&m[772])|(m[438]&m[768]&~m[770]&~m[771]&m[772])|(m[438]&~m[768]&m[770]&~m[771]&m[772])|(~m[438]&~m[768]&~m[770]&m[771]&m[772])|(m[438]&~m[768]&~m[770]&m[771]&m[772])|(~m[438]&m[768]&~m[770]&m[771]&m[772])|(m[438]&m[768]&~m[770]&m[771]&m[772])|(~m[438]&~m[768]&m[770]&m[771]&m[772])|(m[438]&~m[768]&m[770]&m[771]&m[772])|(m[438]&m[768]&m[770]&m[771]&m[772]))):InitCond[827];
    m[774] = run?((((m[449]&~m[773]&~m[775]&~m[776]&~m[777])|(~m[449]&~m[773]&~m[775]&m[776]&~m[777])|(m[449]&m[773]&~m[775]&m[776]&~m[777])|(m[449]&~m[773]&m[775]&m[776]&~m[777])|(~m[449]&m[773]&~m[775]&~m[776]&m[777])|(~m[449]&~m[773]&m[775]&~m[776]&m[777])|(m[449]&m[773]&m[775]&~m[776]&m[777])|(~m[449]&m[773]&m[775]&m[776]&m[777]))&UnbiasedRNG[301])|((m[449]&~m[773]&~m[775]&m[776]&~m[777])|(~m[449]&~m[773]&~m[775]&~m[776]&m[777])|(m[449]&~m[773]&~m[775]&~m[776]&m[777])|(m[449]&m[773]&~m[775]&~m[776]&m[777])|(m[449]&~m[773]&m[775]&~m[776]&m[777])|(~m[449]&~m[773]&~m[775]&m[776]&m[777])|(m[449]&~m[773]&~m[775]&m[776]&m[777])|(~m[449]&m[773]&~m[775]&m[776]&m[777])|(m[449]&m[773]&~m[775]&m[776]&m[777])|(~m[449]&~m[773]&m[775]&m[776]&m[777])|(m[449]&~m[773]&m[775]&m[776]&m[777])|(m[449]&m[773]&m[775]&m[776]&m[777]))):InitCond[828];
    m[779] = run?((((m[460]&~m[778]&~m[780]&~m[781]&~m[782])|(~m[460]&~m[778]&~m[780]&m[781]&~m[782])|(m[460]&m[778]&~m[780]&m[781]&~m[782])|(m[460]&~m[778]&m[780]&m[781]&~m[782])|(~m[460]&m[778]&~m[780]&~m[781]&m[782])|(~m[460]&~m[778]&m[780]&~m[781]&m[782])|(m[460]&m[778]&m[780]&~m[781]&m[782])|(~m[460]&m[778]&m[780]&m[781]&m[782]))&UnbiasedRNG[302])|((m[460]&~m[778]&~m[780]&m[781]&~m[782])|(~m[460]&~m[778]&~m[780]&~m[781]&m[782])|(m[460]&~m[778]&~m[780]&~m[781]&m[782])|(m[460]&m[778]&~m[780]&~m[781]&m[782])|(m[460]&~m[778]&m[780]&~m[781]&m[782])|(~m[460]&~m[778]&~m[780]&m[781]&m[782])|(m[460]&~m[778]&~m[780]&m[781]&m[782])|(~m[460]&m[778]&~m[780]&m[781]&m[782])|(m[460]&m[778]&~m[780]&m[781]&m[782])|(~m[460]&~m[778]&m[780]&m[781]&m[782])|(m[460]&~m[778]&m[780]&m[781]&m[782])|(m[460]&m[778]&m[780]&m[781]&m[782]))):InitCond[829];
    m[784] = run?((((m[471]&~m[783]&~m[785]&~m[786]&~m[787])|(~m[471]&~m[783]&~m[785]&m[786]&~m[787])|(m[471]&m[783]&~m[785]&m[786]&~m[787])|(m[471]&~m[783]&m[785]&m[786]&~m[787])|(~m[471]&m[783]&~m[785]&~m[786]&m[787])|(~m[471]&~m[783]&m[785]&~m[786]&m[787])|(m[471]&m[783]&m[785]&~m[786]&m[787])|(~m[471]&m[783]&m[785]&m[786]&m[787]))&UnbiasedRNG[303])|((m[471]&~m[783]&~m[785]&m[786]&~m[787])|(~m[471]&~m[783]&~m[785]&~m[786]&m[787])|(m[471]&~m[783]&~m[785]&~m[786]&m[787])|(m[471]&m[783]&~m[785]&~m[786]&m[787])|(m[471]&~m[783]&m[785]&~m[786]&m[787])|(~m[471]&~m[783]&~m[785]&m[786]&m[787])|(m[471]&~m[783]&~m[785]&m[786]&m[787])|(~m[471]&m[783]&~m[785]&m[786]&m[787])|(m[471]&m[783]&~m[785]&m[786]&m[787])|(~m[471]&~m[783]&m[785]&m[786]&m[787])|(m[471]&~m[783]&m[785]&m[786]&m[787])|(m[471]&m[783]&m[785]&m[786]&m[787]))):InitCond[830];
    m[789] = run?((((m[482]&~m[788]&~m[790]&~m[791]&~m[792])|(~m[482]&~m[788]&~m[790]&m[791]&~m[792])|(m[482]&m[788]&~m[790]&m[791]&~m[792])|(m[482]&~m[788]&m[790]&m[791]&~m[792])|(~m[482]&m[788]&~m[790]&~m[791]&m[792])|(~m[482]&~m[788]&m[790]&~m[791]&m[792])|(m[482]&m[788]&m[790]&~m[791]&m[792])|(~m[482]&m[788]&m[790]&m[791]&m[792]))&UnbiasedRNG[304])|((m[482]&~m[788]&~m[790]&m[791]&~m[792])|(~m[482]&~m[788]&~m[790]&~m[791]&m[792])|(m[482]&~m[788]&~m[790]&~m[791]&m[792])|(m[482]&m[788]&~m[790]&~m[791]&m[792])|(m[482]&~m[788]&m[790]&~m[791]&m[792])|(~m[482]&~m[788]&~m[790]&m[791]&m[792])|(m[482]&~m[788]&~m[790]&m[791]&m[792])|(~m[482]&m[788]&~m[790]&m[791]&m[792])|(m[482]&m[788]&~m[790]&m[791]&m[792])|(~m[482]&~m[788]&m[790]&m[791]&m[792])|(m[482]&~m[788]&m[790]&m[791]&m[792])|(m[482]&m[788]&m[790]&m[791]&m[792]))):InitCond[831];
    m[794] = run?((((m[493]&~m[793]&~m[795]&~m[796]&~m[797])|(~m[493]&~m[793]&~m[795]&m[796]&~m[797])|(m[493]&m[793]&~m[795]&m[796]&~m[797])|(m[493]&~m[793]&m[795]&m[796]&~m[797])|(~m[493]&m[793]&~m[795]&~m[796]&m[797])|(~m[493]&~m[793]&m[795]&~m[796]&m[797])|(m[493]&m[793]&m[795]&~m[796]&m[797])|(~m[493]&m[793]&m[795]&m[796]&m[797]))&UnbiasedRNG[305])|((m[493]&~m[793]&~m[795]&m[796]&~m[797])|(~m[493]&~m[793]&~m[795]&~m[796]&m[797])|(m[493]&~m[793]&~m[795]&~m[796]&m[797])|(m[493]&m[793]&~m[795]&~m[796]&m[797])|(m[493]&~m[793]&m[795]&~m[796]&m[797])|(~m[493]&~m[793]&~m[795]&m[796]&m[797])|(m[493]&~m[793]&~m[795]&m[796]&m[797])|(~m[493]&m[793]&~m[795]&m[796]&m[797])|(m[493]&m[793]&~m[795]&m[796]&m[797])|(~m[493]&~m[793]&m[795]&m[796]&m[797])|(m[493]&~m[793]&m[795]&m[796]&m[797])|(m[493]&m[793]&m[795]&m[796]&m[797]))):InitCond[832];
    m[799] = run?((((m[504]&~m[798]&~m[800]&~m[801]&~m[802])|(~m[504]&~m[798]&~m[800]&m[801]&~m[802])|(m[504]&m[798]&~m[800]&m[801]&~m[802])|(m[504]&~m[798]&m[800]&m[801]&~m[802])|(~m[504]&m[798]&~m[800]&~m[801]&m[802])|(~m[504]&~m[798]&m[800]&~m[801]&m[802])|(m[504]&m[798]&m[800]&~m[801]&m[802])|(~m[504]&m[798]&m[800]&m[801]&m[802]))&UnbiasedRNG[306])|((m[504]&~m[798]&~m[800]&m[801]&~m[802])|(~m[504]&~m[798]&~m[800]&~m[801]&m[802])|(m[504]&~m[798]&~m[800]&~m[801]&m[802])|(m[504]&m[798]&~m[800]&~m[801]&m[802])|(m[504]&~m[798]&m[800]&~m[801]&m[802])|(~m[504]&~m[798]&~m[800]&m[801]&m[802])|(m[504]&~m[798]&~m[800]&m[801]&m[802])|(~m[504]&m[798]&~m[800]&m[801]&m[802])|(m[504]&m[798]&~m[800]&m[801]&m[802])|(~m[504]&~m[798]&m[800]&m[801]&m[802])|(m[504]&~m[798]&m[800]&m[801]&m[802])|(m[504]&m[798]&m[800]&m[801]&m[802]))):InitCond[833];
    m[804] = run?((((m[406]&~m[803]&~m[805]&~m[806]&~m[807])|(~m[406]&~m[803]&~m[805]&m[806]&~m[807])|(m[406]&m[803]&~m[805]&m[806]&~m[807])|(m[406]&~m[803]&m[805]&m[806]&~m[807])|(~m[406]&m[803]&~m[805]&~m[806]&m[807])|(~m[406]&~m[803]&m[805]&~m[806]&m[807])|(m[406]&m[803]&m[805]&~m[806]&m[807])|(~m[406]&m[803]&m[805]&m[806]&m[807]))&UnbiasedRNG[307])|((m[406]&~m[803]&~m[805]&m[806]&~m[807])|(~m[406]&~m[803]&~m[805]&~m[806]&m[807])|(m[406]&~m[803]&~m[805]&~m[806]&m[807])|(m[406]&m[803]&~m[805]&~m[806]&m[807])|(m[406]&~m[803]&m[805]&~m[806]&m[807])|(~m[406]&~m[803]&~m[805]&m[806]&m[807])|(m[406]&~m[803]&~m[805]&m[806]&m[807])|(~m[406]&m[803]&~m[805]&m[806]&m[807])|(m[406]&m[803]&~m[805]&m[806]&m[807])|(~m[406]&~m[803]&m[805]&m[806]&m[807])|(m[406]&~m[803]&m[805]&m[806]&m[807])|(m[406]&m[803]&m[805]&m[806]&m[807]))):InitCond[834];
    m[809] = run?((((m[417]&~m[808]&~m[810]&~m[811]&~m[812])|(~m[417]&~m[808]&~m[810]&m[811]&~m[812])|(m[417]&m[808]&~m[810]&m[811]&~m[812])|(m[417]&~m[808]&m[810]&m[811]&~m[812])|(~m[417]&m[808]&~m[810]&~m[811]&m[812])|(~m[417]&~m[808]&m[810]&~m[811]&m[812])|(m[417]&m[808]&m[810]&~m[811]&m[812])|(~m[417]&m[808]&m[810]&m[811]&m[812]))&UnbiasedRNG[308])|((m[417]&~m[808]&~m[810]&m[811]&~m[812])|(~m[417]&~m[808]&~m[810]&~m[811]&m[812])|(m[417]&~m[808]&~m[810]&~m[811]&m[812])|(m[417]&m[808]&~m[810]&~m[811]&m[812])|(m[417]&~m[808]&m[810]&~m[811]&m[812])|(~m[417]&~m[808]&~m[810]&m[811]&m[812])|(m[417]&~m[808]&~m[810]&m[811]&m[812])|(~m[417]&m[808]&~m[810]&m[811]&m[812])|(m[417]&m[808]&~m[810]&m[811]&m[812])|(~m[417]&~m[808]&m[810]&m[811]&m[812])|(m[417]&~m[808]&m[810]&m[811]&m[812])|(m[417]&m[808]&m[810]&m[811]&m[812]))):InitCond[835];
    m[814] = run?((((m[428]&~m[813]&~m[815]&~m[816]&~m[817])|(~m[428]&~m[813]&~m[815]&m[816]&~m[817])|(m[428]&m[813]&~m[815]&m[816]&~m[817])|(m[428]&~m[813]&m[815]&m[816]&~m[817])|(~m[428]&m[813]&~m[815]&~m[816]&m[817])|(~m[428]&~m[813]&m[815]&~m[816]&m[817])|(m[428]&m[813]&m[815]&~m[816]&m[817])|(~m[428]&m[813]&m[815]&m[816]&m[817]))&UnbiasedRNG[309])|((m[428]&~m[813]&~m[815]&m[816]&~m[817])|(~m[428]&~m[813]&~m[815]&~m[816]&m[817])|(m[428]&~m[813]&~m[815]&~m[816]&m[817])|(m[428]&m[813]&~m[815]&~m[816]&m[817])|(m[428]&~m[813]&m[815]&~m[816]&m[817])|(~m[428]&~m[813]&~m[815]&m[816]&m[817])|(m[428]&~m[813]&~m[815]&m[816]&m[817])|(~m[428]&m[813]&~m[815]&m[816]&m[817])|(m[428]&m[813]&~m[815]&m[816]&m[817])|(~m[428]&~m[813]&m[815]&m[816]&m[817])|(m[428]&~m[813]&m[815]&m[816]&m[817])|(m[428]&m[813]&m[815]&m[816]&m[817]))):InitCond[836];
    m[819] = run?((((m[439]&~m[818]&~m[820]&~m[821]&~m[822])|(~m[439]&~m[818]&~m[820]&m[821]&~m[822])|(m[439]&m[818]&~m[820]&m[821]&~m[822])|(m[439]&~m[818]&m[820]&m[821]&~m[822])|(~m[439]&m[818]&~m[820]&~m[821]&m[822])|(~m[439]&~m[818]&m[820]&~m[821]&m[822])|(m[439]&m[818]&m[820]&~m[821]&m[822])|(~m[439]&m[818]&m[820]&m[821]&m[822]))&UnbiasedRNG[310])|((m[439]&~m[818]&~m[820]&m[821]&~m[822])|(~m[439]&~m[818]&~m[820]&~m[821]&m[822])|(m[439]&~m[818]&~m[820]&~m[821]&m[822])|(m[439]&m[818]&~m[820]&~m[821]&m[822])|(m[439]&~m[818]&m[820]&~m[821]&m[822])|(~m[439]&~m[818]&~m[820]&m[821]&m[822])|(m[439]&~m[818]&~m[820]&m[821]&m[822])|(~m[439]&m[818]&~m[820]&m[821]&m[822])|(m[439]&m[818]&~m[820]&m[821]&m[822])|(~m[439]&~m[818]&m[820]&m[821]&m[822])|(m[439]&~m[818]&m[820]&m[821]&m[822])|(m[439]&m[818]&m[820]&m[821]&m[822]))):InitCond[837];
    m[824] = run?((((m[450]&~m[823]&~m[825]&~m[826]&~m[827])|(~m[450]&~m[823]&~m[825]&m[826]&~m[827])|(m[450]&m[823]&~m[825]&m[826]&~m[827])|(m[450]&~m[823]&m[825]&m[826]&~m[827])|(~m[450]&m[823]&~m[825]&~m[826]&m[827])|(~m[450]&~m[823]&m[825]&~m[826]&m[827])|(m[450]&m[823]&m[825]&~m[826]&m[827])|(~m[450]&m[823]&m[825]&m[826]&m[827]))&UnbiasedRNG[311])|((m[450]&~m[823]&~m[825]&m[826]&~m[827])|(~m[450]&~m[823]&~m[825]&~m[826]&m[827])|(m[450]&~m[823]&~m[825]&~m[826]&m[827])|(m[450]&m[823]&~m[825]&~m[826]&m[827])|(m[450]&~m[823]&m[825]&~m[826]&m[827])|(~m[450]&~m[823]&~m[825]&m[826]&m[827])|(m[450]&~m[823]&~m[825]&m[826]&m[827])|(~m[450]&m[823]&~m[825]&m[826]&m[827])|(m[450]&m[823]&~m[825]&m[826]&m[827])|(~m[450]&~m[823]&m[825]&m[826]&m[827])|(m[450]&~m[823]&m[825]&m[826]&m[827])|(m[450]&m[823]&m[825]&m[826]&m[827]))):InitCond[838];
    m[829] = run?((((m[461]&~m[828]&~m[830]&~m[831]&~m[832])|(~m[461]&~m[828]&~m[830]&m[831]&~m[832])|(m[461]&m[828]&~m[830]&m[831]&~m[832])|(m[461]&~m[828]&m[830]&m[831]&~m[832])|(~m[461]&m[828]&~m[830]&~m[831]&m[832])|(~m[461]&~m[828]&m[830]&~m[831]&m[832])|(m[461]&m[828]&m[830]&~m[831]&m[832])|(~m[461]&m[828]&m[830]&m[831]&m[832]))&UnbiasedRNG[312])|((m[461]&~m[828]&~m[830]&m[831]&~m[832])|(~m[461]&~m[828]&~m[830]&~m[831]&m[832])|(m[461]&~m[828]&~m[830]&~m[831]&m[832])|(m[461]&m[828]&~m[830]&~m[831]&m[832])|(m[461]&~m[828]&m[830]&~m[831]&m[832])|(~m[461]&~m[828]&~m[830]&m[831]&m[832])|(m[461]&~m[828]&~m[830]&m[831]&m[832])|(~m[461]&m[828]&~m[830]&m[831]&m[832])|(m[461]&m[828]&~m[830]&m[831]&m[832])|(~m[461]&~m[828]&m[830]&m[831]&m[832])|(m[461]&~m[828]&m[830]&m[831]&m[832])|(m[461]&m[828]&m[830]&m[831]&m[832]))):InitCond[839];
    m[834] = run?((((m[472]&~m[833]&~m[835]&~m[836]&~m[837])|(~m[472]&~m[833]&~m[835]&m[836]&~m[837])|(m[472]&m[833]&~m[835]&m[836]&~m[837])|(m[472]&~m[833]&m[835]&m[836]&~m[837])|(~m[472]&m[833]&~m[835]&~m[836]&m[837])|(~m[472]&~m[833]&m[835]&~m[836]&m[837])|(m[472]&m[833]&m[835]&~m[836]&m[837])|(~m[472]&m[833]&m[835]&m[836]&m[837]))&UnbiasedRNG[313])|((m[472]&~m[833]&~m[835]&m[836]&~m[837])|(~m[472]&~m[833]&~m[835]&~m[836]&m[837])|(m[472]&~m[833]&~m[835]&~m[836]&m[837])|(m[472]&m[833]&~m[835]&~m[836]&m[837])|(m[472]&~m[833]&m[835]&~m[836]&m[837])|(~m[472]&~m[833]&~m[835]&m[836]&m[837])|(m[472]&~m[833]&~m[835]&m[836]&m[837])|(~m[472]&m[833]&~m[835]&m[836]&m[837])|(m[472]&m[833]&~m[835]&m[836]&m[837])|(~m[472]&~m[833]&m[835]&m[836]&m[837])|(m[472]&~m[833]&m[835]&m[836]&m[837])|(m[472]&m[833]&m[835]&m[836]&m[837]))):InitCond[840];
    m[839] = run?((((m[483]&~m[838]&~m[840]&~m[841]&~m[842])|(~m[483]&~m[838]&~m[840]&m[841]&~m[842])|(m[483]&m[838]&~m[840]&m[841]&~m[842])|(m[483]&~m[838]&m[840]&m[841]&~m[842])|(~m[483]&m[838]&~m[840]&~m[841]&m[842])|(~m[483]&~m[838]&m[840]&~m[841]&m[842])|(m[483]&m[838]&m[840]&~m[841]&m[842])|(~m[483]&m[838]&m[840]&m[841]&m[842]))&UnbiasedRNG[314])|((m[483]&~m[838]&~m[840]&m[841]&~m[842])|(~m[483]&~m[838]&~m[840]&~m[841]&m[842])|(m[483]&~m[838]&~m[840]&~m[841]&m[842])|(m[483]&m[838]&~m[840]&~m[841]&m[842])|(m[483]&~m[838]&m[840]&~m[841]&m[842])|(~m[483]&~m[838]&~m[840]&m[841]&m[842])|(m[483]&~m[838]&~m[840]&m[841]&m[842])|(~m[483]&m[838]&~m[840]&m[841]&m[842])|(m[483]&m[838]&~m[840]&m[841]&m[842])|(~m[483]&~m[838]&m[840]&m[841]&m[842])|(m[483]&~m[838]&m[840]&m[841]&m[842])|(m[483]&m[838]&m[840]&m[841]&m[842]))):InitCond[841];
    m[844] = run?((((m[494]&~m[843]&~m[845]&~m[846]&~m[847])|(~m[494]&~m[843]&~m[845]&m[846]&~m[847])|(m[494]&m[843]&~m[845]&m[846]&~m[847])|(m[494]&~m[843]&m[845]&m[846]&~m[847])|(~m[494]&m[843]&~m[845]&~m[846]&m[847])|(~m[494]&~m[843]&m[845]&~m[846]&m[847])|(m[494]&m[843]&m[845]&~m[846]&m[847])|(~m[494]&m[843]&m[845]&m[846]&m[847]))&UnbiasedRNG[315])|((m[494]&~m[843]&~m[845]&m[846]&~m[847])|(~m[494]&~m[843]&~m[845]&~m[846]&m[847])|(m[494]&~m[843]&~m[845]&~m[846]&m[847])|(m[494]&m[843]&~m[845]&~m[846]&m[847])|(m[494]&~m[843]&m[845]&~m[846]&m[847])|(~m[494]&~m[843]&~m[845]&m[846]&m[847])|(m[494]&~m[843]&~m[845]&m[846]&m[847])|(~m[494]&m[843]&~m[845]&m[846]&m[847])|(m[494]&m[843]&~m[845]&m[846]&m[847])|(~m[494]&~m[843]&m[845]&m[846]&m[847])|(m[494]&~m[843]&m[845]&m[846]&m[847])|(m[494]&m[843]&m[845]&m[846]&m[847]))):InitCond[842];
    m[849] = run?((((m[505]&~m[848]&~m[850]&~m[851]&~m[852])|(~m[505]&~m[848]&~m[850]&m[851]&~m[852])|(m[505]&m[848]&~m[850]&m[851]&~m[852])|(m[505]&~m[848]&m[850]&m[851]&~m[852])|(~m[505]&m[848]&~m[850]&~m[851]&m[852])|(~m[505]&~m[848]&m[850]&~m[851]&m[852])|(m[505]&m[848]&m[850]&~m[851]&m[852])|(~m[505]&m[848]&m[850]&m[851]&m[852]))&UnbiasedRNG[316])|((m[505]&~m[848]&~m[850]&m[851]&~m[852])|(~m[505]&~m[848]&~m[850]&~m[851]&m[852])|(m[505]&~m[848]&~m[850]&~m[851]&m[852])|(m[505]&m[848]&~m[850]&~m[851]&m[852])|(m[505]&~m[848]&m[850]&~m[851]&m[852])|(~m[505]&~m[848]&~m[850]&m[851]&m[852])|(m[505]&~m[848]&~m[850]&m[851]&m[852])|(~m[505]&m[848]&~m[850]&m[851]&m[852])|(m[505]&m[848]&~m[850]&m[851]&m[852])|(~m[505]&~m[848]&m[850]&m[851]&m[852])|(m[505]&~m[848]&m[850]&m[851]&m[852])|(m[505]&m[848]&m[850]&m[851]&m[852]))):InitCond[843];
    m[854] = run?((((m[516]&~m[853]&~m[855]&~m[856]&~m[857])|(~m[516]&~m[853]&~m[855]&m[856]&~m[857])|(m[516]&m[853]&~m[855]&m[856]&~m[857])|(m[516]&~m[853]&m[855]&m[856]&~m[857])|(~m[516]&m[853]&~m[855]&~m[856]&m[857])|(~m[516]&~m[853]&m[855]&~m[856]&m[857])|(m[516]&m[853]&m[855]&~m[856]&m[857])|(~m[516]&m[853]&m[855]&m[856]&m[857]))&UnbiasedRNG[317])|((m[516]&~m[853]&~m[855]&m[856]&~m[857])|(~m[516]&~m[853]&~m[855]&~m[856]&m[857])|(m[516]&~m[853]&~m[855]&~m[856]&m[857])|(m[516]&m[853]&~m[855]&~m[856]&m[857])|(m[516]&~m[853]&m[855]&~m[856]&m[857])|(~m[516]&~m[853]&~m[855]&m[856]&m[857])|(m[516]&~m[853]&~m[855]&m[856]&m[857])|(~m[516]&m[853]&~m[855]&m[856]&m[857])|(m[516]&m[853]&~m[855]&m[856]&m[857])|(~m[516]&~m[853]&m[855]&m[856]&m[857])|(m[516]&~m[853]&m[855]&m[856]&m[857])|(m[516]&m[853]&m[855]&m[856]&m[857]))):InitCond[844];
    m[859] = run?((((m[407]&~m[858]&~m[860]&~m[861]&~m[862])|(~m[407]&~m[858]&~m[860]&m[861]&~m[862])|(m[407]&m[858]&~m[860]&m[861]&~m[862])|(m[407]&~m[858]&m[860]&m[861]&~m[862])|(~m[407]&m[858]&~m[860]&~m[861]&m[862])|(~m[407]&~m[858]&m[860]&~m[861]&m[862])|(m[407]&m[858]&m[860]&~m[861]&m[862])|(~m[407]&m[858]&m[860]&m[861]&m[862]))&UnbiasedRNG[318])|((m[407]&~m[858]&~m[860]&m[861]&~m[862])|(~m[407]&~m[858]&~m[860]&~m[861]&m[862])|(m[407]&~m[858]&~m[860]&~m[861]&m[862])|(m[407]&m[858]&~m[860]&~m[861]&m[862])|(m[407]&~m[858]&m[860]&~m[861]&m[862])|(~m[407]&~m[858]&~m[860]&m[861]&m[862])|(m[407]&~m[858]&~m[860]&m[861]&m[862])|(~m[407]&m[858]&~m[860]&m[861]&m[862])|(m[407]&m[858]&~m[860]&m[861]&m[862])|(~m[407]&~m[858]&m[860]&m[861]&m[862])|(m[407]&~m[858]&m[860]&m[861]&m[862])|(m[407]&m[858]&m[860]&m[861]&m[862]))):InitCond[845];
    m[864] = run?((((m[418]&~m[863]&~m[865]&~m[866]&~m[867])|(~m[418]&~m[863]&~m[865]&m[866]&~m[867])|(m[418]&m[863]&~m[865]&m[866]&~m[867])|(m[418]&~m[863]&m[865]&m[866]&~m[867])|(~m[418]&m[863]&~m[865]&~m[866]&m[867])|(~m[418]&~m[863]&m[865]&~m[866]&m[867])|(m[418]&m[863]&m[865]&~m[866]&m[867])|(~m[418]&m[863]&m[865]&m[866]&m[867]))&UnbiasedRNG[319])|((m[418]&~m[863]&~m[865]&m[866]&~m[867])|(~m[418]&~m[863]&~m[865]&~m[866]&m[867])|(m[418]&~m[863]&~m[865]&~m[866]&m[867])|(m[418]&m[863]&~m[865]&~m[866]&m[867])|(m[418]&~m[863]&m[865]&~m[866]&m[867])|(~m[418]&~m[863]&~m[865]&m[866]&m[867])|(m[418]&~m[863]&~m[865]&m[866]&m[867])|(~m[418]&m[863]&~m[865]&m[866]&m[867])|(m[418]&m[863]&~m[865]&m[866]&m[867])|(~m[418]&~m[863]&m[865]&m[866]&m[867])|(m[418]&~m[863]&m[865]&m[866]&m[867])|(m[418]&m[863]&m[865]&m[866]&m[867]))):InitCond[846];
    m[869] = run?((((m[429]&~m[868]&~m[870]&~m[871]&~m[872])|(~m[429]&~m[868]&~m[870]&m[871]&~m[872])|(m[429]&m[868]&~m[870]&m[871]&~m[872])|(m[429]&~m[868]&m[870]&m[871]&~m[872])|(~m[429]&m[868]&~m[870]&~m[871]&m[872])|(~m[429]&~m[868]&m[870]&~m[871]&m[872])|(m[429]&m[868]&m[870]&~m[871]&m[872])|(~m[429]&m[868]&m[870]&m[871]&m[872]))&UnbiasedRNG[320])|((m[429]&~m[868]&~m[870]&m[871]&~m[872])|(~m[429]&~m[868]&~m[870]&~m[871]&m[872])|(m[429]&~m[868]&~m[870]&~m[871]&m[872])|(m[429]&m[868]&~m[870]&~m[871]&m[872])|(m[429]&~m[868]&m[870]&~m[871]&m[872])|(~m[429]&~m[868]&~m[870]&m[871]&m[872])|(m[429]&~m[868]&~m[870]&m[871]&m[872])|(~m[429]&m[868]&~m[870]&m[871]&m[872])|(m[429]&m[868]&~m[870]&m[871]&m[872])|(~m[429]&~m[868]&m[870]&m[871]&m[872])|(m[429]&~m[868]&m[870]&m[871]&m[872])|(m[429]&m[868]&m[870]&m[871]&m[872]))):InitCond[847];
    m[874] = run?((((m[440]&~m[873]&~m[875]&~m[876]&~m[877])|(~m[440]&~m[873]&~m[875]&m[876]&~m[877])|(m[440]&m[873]&~m[875]&m[876]&~m[877])|(m[440]&~m[873]&m[875]&m[876]&~m[877])|(~m[440]&m[873]&~m[875]&~m[876]&m[877])|(~m[440]&~m[873]&m[875]&~m[876]&m[877])|(m[440]&m[873]&m[875]&~m[876]&m[877])|(~m[440]&m[873]&m[875]&m[876]&m[877]))&UnbiasedRNG[321])|((m[440]&~m[873]&~m[875]&m[876]&~m[877])|(~m[440]&~m[873]&~m[875]&~m[876]&m[877])|(m[440]&~m[873]&~m[875]&~m[876]&m[877])|(m[440]&m[873]&~m[875]&~m[876]&m[877])|(m[440]&~m[873]&m[875]&~m[876]&m[877])|(~m[440]&~m[873]&~m[875]&m[876]&m[877])|(m[440]&~m[873]&~m[875]&m[876]&m[877])|(~m[440]&m[873]&~m[875]&m[876]&m[877])|(m[440]&m[873]&~m[875]&m[876]&m[877])|(~m[440]&~m[873]&m[875]&m[876]&m[877])|(m[440]&~m[873]&m[875]&m[876]&m[877])|(m[440]&m[873]&m[875]&m[876]&m[877]))):InitCond[848];
    m[879] = run?((((m[451]&~m[878]&~m[880]&~m[881]&~m[882])|(~m[451]&~m[878]&~m[880]&m[881]&~m[882])|(m[451]&m[878]&~m[880]&m[881]&~m[882])|(m[451]&~m[878]&m[880]&m[881]&~m[882])|(~m[451]&m[878]&~m[880]&~m[881]&m[882])|(~m[451]&~m[878]&m[880]&~m[881]&m[882])|(m[451]&m[878]&m[880]&~m[881]&m[882])|(~m[451]&m[878]&m[880]&m[881]&m[882]))&UnbiasedRNG[322])|((m[451]&~m[878]&~m[880]&m[881]&~m[882])|(~m[451]&~m[878]&~m[880]&~m[881]&m[882])|(m[451]&~m[878]&~m[880]&~m[881]&m[882])|(m[451]&m[878]&~m[880]&~m[881]&m[882])|(m[451]&~m[878]&m[880]&~m[881]&m[882])|(~m[451]&~m[878]&~m[880]&m[881]&m[882])|(m[451]&~m[878]&~m[880]&m[881]&m[882])|(~m[451]&m[878]&~m[880]&m[881]&m[882])|(m[451]&m[878]&~m[880]&m[881]&m[882])|(~m[451]&~m[878]&m[880]&m[881]&m[882])|(m[451]&~m[878]&m[880]&m[881]&m[882])|(m[451]&m[878]&m[880]&m[881]&m[882]))):InitCond[849];
    m[884] = run?((((m[462]&~m[883]&~m[885]&~m[886]&~m[887])|(~m[462]&~m[883]&~m[885]&m[886]&~m[887])|(m[462]&m[883]&~m[885]&m[886]&~m[887])|(m[462]&~m[883]&m[885]&m[886]&~m[887])|(~m[462]&m[883]&~m[885]&~m[886]&m[887])|(~m[462]&~m[883]&m[885]&~m[886]&m[887])|(m[462]&m[883]&m[885]&~m[886]&m[887])|(~m[462]&m[883]&m[885]&m[886]&m[887]))&UnbiasedRNG[323])|((m[462]&~m[883]&~m[885]&m[886]&~m[887])|(~m[462]&~m[883]&~m[885]&~m[886]&m[887])|(m[462]&~m[883]&~m[885]&~m[886]&m[887])|(m[462]&m[883]&~m[885]&~m[886]&m[887])|(m[462]&~m[883]&m[885]&~m[886]&m[887])|(~m[462]&~m[883]&~m[885]&m[886]&m[887])|(m[462]&~m[883]&~m[885]&m[886]&m[887])|(~m[462]&m[883]&~m[885]&m[886]&m[887])|(m[462]&m[883]&~m[885]&m[886]&m[887])|(~m[462]&~m[883]&m[885]&m[886]&m[887])|(m[462]&~m[883]&m[885]&m[886]&m[887])|(m[462]&m[883]&m[885]&m[886]&m[887]))):InitCond[850];
    m[889] = run?((((m[473]&~m[888]&~m[890]&~m[891]&~m[892])|(~m[473]&~m[888]&~m[890]&m[891]&~m[892])|(m[473]&m[888]&~m[890]&m[891]&~m[892])|(m[473]&~m[888]&m[890]&m[891]&~m[892])|(~m[473]&m[888]&~m[890]&~m[891]&m[892])|(~m[473]&~m[888]&m[890]&~m[891]&m[892])|(m[473]&m[888]&m[890]&~m[891]&m[892])|(~m[473]&m[888]&m[890]&m[891]&m[892]))&UnbiasedRNG[324])|((m[473]&~m[888]&~m[890]&m[891]&~m[892])|(~m[473]&~m[888]&~m[890]&~m[891]&m[892])|(m[473]&~m[888]&~m[890]&~m[891]&m[892])|(m[473]&m[888]&~m[890]&~m[891]&m[892])|(m[473]&~m[888]&m[890]&~m[891]&m[892])|(~m[473]&~m[888]&~m[890]&m[891]&m[892])|(m[473]&~m[888]&~m[890]&m[891]&m[892])|(~m[473]&m[888]&~m[890]&m[891]&m[892])|(m[473]&m[888]&~m[890]&m[891]&m[892])|(~m[473]&~m[888]&m[890]&m[891]&m[892])|(m[473]&~m[888]&m[890]&m[891]&m[892])|(m[473]&m[888]&m[890]&m[891]&m[892]))):InitCond[851];
    m[894] = run?((((m[484]&~m[893]&~m[895]&~m[896]&~m[897])|(~m[484]&~m[893]&~m[895]&m[896]&~m[897])|(m[484]&m[893]&~m[895]&m[896]&~m[897])|(m[484]&~m[893]&m[895]&m[896]&~m[897])|(~m[484]&m[893]&~m[895]&~m[896]&m[897])|(~m[484]&~m[893]&m[895]&~m[896]&m[897])|(m[484]&m[893]&m[895]&~m[896]&m[897])|(~m[484]&m[893]&m[895]&m[896]&m[897]))&UnbiasedRNG[325])|((m[484]&~m[893]&~m[895]&m[896]&~m[897])|(~m[484]&~m[893]&~m[895]&~m[896]&m[897])|(m[484]&~m[893]&~m[895]&~m[896]&m[897])|(m[484]&m[893]&~m[895]&~m[896]&m[897])|(m[484]&~m[893]&m[895]&~m[896]&m[897])|(~m[484]&~m[893]&~m[895]&m[896]&m[897])|(m[484]&~m[893]&~m[895]&m[896]&m[897])|(~m[484]&m[893]&~m[895]&m[896]&m[897])|(m[484]&m[893]&~m[895]&m[896]&m[897])|(~m[484]&~m[893]&m[895]&m[896]&m[897])|(m[484]&~m[893]&m[895]&m[896]&m[897])|(m[484]&m[893]&m[895]&m[896]&m[897]))):InitCond[852];
    m[899] = run?((((m[495]&~m[898]&~m[900]&~m[901]&~m[902])|(~m[495]&~m[898]&~m[900]&m[901]&~m[902])|(m[495]&m[898]&~m[900]&m[901]&~m[902])|(m[495]&~m[898]&m[900]&m[901]&~m[902])|(~m[495]&m[898]&~m[900]&~m[901]&m[902])|(~m[495]&~m[898]&m[900]&~m[901]&m[902])|(m[495]&m[898]&m[900]&~m[901]&m[902])|(~m[495]&m[898]&m[900]&m[901]&m[902]))&UnbiasedRNG[326])|((m[495]&~m[898]&~m[900]&m[901]&~m[902])|(~m[495]&~m[898]&~m[900]&~m[901]&m[902])|(m[495]&~m[898]&~m[900]&~m[901]&m[902])|(m[495]&m[898]&~m[900]&~m[901]&m[902])|(m[495]&~m[898]&m[900]&~m[901]&m[902])|(~m[495]&~m[898]&~m[900]&m[901]&m[902])|(m[495]&~m[898]&~m[900]&m[901]&m[902])|(~m[495]&m[898]&~m[900]&m[901]&m[902])|(m[495]&m[898]&~m[900]&m[901]&m[902])|(~m[495]&~m[898]&m[900]&m[901]&m[902])|(m[495]&~m[898]&m[900]&m[901]&m[902])|(m[495]&m[898]&m[900]&m[901]&m[902]))):InitCond[853];
    m[904] = run?((((m[506]&~m[903]&~m[905]&~m[906]&~m[907])|(~m[506]&~m[903]&~m[905]&m[906]&~m[907])|(m[506]&m[903]&~m[905]&m[906]&~m[907])|(m[506]&~m[903]&m[905]&m[906]&~m[907])|(~m[506]&m[903]&~m[905]&~m[906]&m[907])|(~m[506]&~m[903]&m[905]&~m[906]&m[907])|(m[506]&m[903]&m[905]&~m[906]&m[907])|(~m[506]&m[903]&m[905]&m[906]&m[907]))&UnbiasedRNG[327])|((m[506]&~m[903]&~m[905]&m[906]&~m[907])|(~m[506]&~m[903]&~m[905]&~m[906]&m[907])|(m[506]&~m[903]&~m[905]&~m[906]&m[907])|(m[506]&m[903]&~m[905]&~m[906]&m[907])|(m[506]&~m[903]&m[905]&~m[906]&m[907])|(~m[506]&~m[903]&~m[905]&m[906]&m[907])|(m[506]&~m[903]&~m[905]&m[906]&m[907])|(~m[506]&m[903]&~m[905]&m[906]&m[907])|(m[506]&m[903]&~m[905]&m[906]&m[907])|(~m[506]&~m[903]&m[905]&m[906]&m[907])|(m[506]&~m[903]&m[905]&m[906]&m[907])|(m[506]&m[903]&m[905]&m[906]&m[907]))):InitCond[854];
    m[909] = run?((((m[517]&~m[908]&~m[910]&~m[911]&~m[912])|(~m[517]&~m[908]&~m[910]&m[911]&~m[912])|(m[517]&m[908]&~m[910]&m[911]&~m[912])|(m[517]&~m[908]&m[910]&m[911]&~m[912])|(~m[517]&m[908]&~m[910]&~m[911]&m[912])|(~m[517]&~m[908]&m[910]&~m[911]&m[912])|(m[517]&m[908]&m[910]&~m[911]&m[912])|(~m[517]&m[908]&m[910]&m[911]&m[912]))&UnbiasedRNG[328])|((m[517]&~m[908]&~m[910]&m[911]&~m[912])|(~m[517]&~m[908]&~m[910]&~m[911]&m[912])|(m[517]&~m[908]&~m[910]&~m[911]&m[912])|(m[517]&m[908]&~m[910]&~m[911]&m[912])|(m[517]&~m[908]&m[910]&~m[911]&m[912])|(~m[517]&~m[908]&~m[910]&m[911]&m[912])|(m[517]&~m[908]&~m[910]&m[911]&m[912])|(~m[517]&m[908]&~m[910]&m[911]&m[912])|(m[517]&m[908]&~m[910]&m[911]&m[912])|(~m[517]&~m[908]&m[910]&m[911]&m[912])|(m[517]&~m[908]&m[910]&m[911]&m[912])|(m[517]&m[908]&m[910]&m[911]&m[912]))):InitCond[855];
    m[914] = run?((((m[419]&~m[913]&~m[915]&~m[916]&~m[917])|(~m[419]&~m[913]&~m[915]&m[916]&~m[917])|(m[419]&m[913]&~m[915]&m[916]&~m[917])|(m[419]&~m[913]&m[915]&m[916]&~m[917])|(~m[419]&m[913]&~m[915]&~m[916]&m[917])|(~m[419]&~m[913]&m[915]&~m[916]&m[917])|(m[419]&m[913]&m[915]&~m[916]&m[917])|(~m[419]&m[913]&m[915]&m[916]&m[917]))&UnbiasedRNG[329])|((m[419]&~m[913]&~m[915]&m[916]&~m[917])|(~m[419]&~m[913]&~m[915]&~m[916]&m[917])|(m[419]&~m[913]&~m[915]&~m[916]&m[917])|(m[419]&m[913]&~m[915]&~m[916]&m[917])|(m[419]&~m[913]&m[915]&~m[916]&m[917])|(~m[419]&~m[913]&~m[915]&m[916]&m[917])|(m[419]&~m[913]&~m[915]&m[916]&m[917])|(~m[419]&m[913]&~m[915]&m[916]&m[917])|(m[419]&m[913]&~m[915]&m[916]&m[917])|(~m[419]&~m[913]&m[915]&m[916]&m[917])|(m[419]&~m[913]&m[915]&m[916]&m[917])|(m[419]&m[913]&m[915]&m[916]&m[917]))):InitCond[856];
    m[919] = run?((((m[430]&~m[918]&~m[920]&~m[921]&~m[922])|(~m[430]&~m[918]&~m[920]&m[921]&~m[922])|(m[430]&m[918]&~m[920]&m[921]&~m[922])|(m[430]&~m[918]&m[920]&m[921]&~m[922])|(~m[430]&m[918]&~m[920]&~m[921]&m[922])|(~m[430]&~m[918]&m[920]&~m[921]&m[922])|(m[430]&m[918]&m[920]&~m[921]&m[922])|(~m[430]&m[918]&m[920]&m[921]&m[922]))&UnbiasedRNG[330])|((m[430]&~m[918]&~m[920]&m[921]&~m[922])|(~m[430]&~m[918]&~m[920]&~m[921]&m[922])|(m[430]&~m[918]&~m[920]&~m[921]&m[922])|(m[430]&m[918]&~m[920]&~m[921]&m[922])|(m[430]&~m[918]&m[920]&~m[921]&m[922])|(~m[430]&~m[918]&~m[920]&m[921]&m[922])|(m[430]&~m[918]&~m[920]&m[921]&m[922])|(~m[430]&m[918]&~m[920]&m[921]&m[922])|(m[430]&m[918]&~m[920]&m[921]&m[922])|(~m[430]&~m[918]&m[920]&m[921]&m[922])|(m[430]&~m[918]&m[920]&m[921]&m[922])|(m[430]&m[918]&m[920]&m[921]&m[922]))):InitCond[857];
    m[924] = run?((((m[441]&~m[923]&~m[925]&~m[926]&~m[927])|(~m[441]&~m[923]&~m[925]&m[926]&~m[927])|(m[441]&m[923]&~m[925]&m[926]&~m[927])|(m[441]&~m[923]&m[925]&m[926]&~m[927])|(~m[441]&m[923]&~m[925]&~m[926]&m[927])|(~m[441]&~m[923]&m[925]&~m[926]&m[927])|(m[441]&m[923]&m[925]&~m[926]&m[927])|(~m[441]&m[923]&m[925]&m[926]&m[927]))&UnbiasedRNG[331])|((m[441]&~m[923]&~m[925]&m[926]&~m[927])|(~m[441]&~m[923]&~m[925]&~m[926]&m[927])|(m[441]&~m[923]&~m[925]&~m[926]&m[927])|(m[441]&m[923]&~m[925]&~m[926]&m[927])|(m[441]&~m[923]&m[925]&~m[926]&m[927])|(~m[441]&~m[923]&~m[925]&m[926]&m[927])|(m[441]&~m[923]&~m[925]&m[926]&m[927])|(~m[441]&m[923]&~m[925]&m[926]&m[927])|(m[441]&m[923]&~m[925]&m[926]&m[927])|(~m[441]&~m[923]&m[925]&m[926]&m[927])|(m[441]&~m[923]&m[925]&m[926]&m[927])|(m[441]&m[923]&m[925]&m[926]&m[927]))):InitCond[858];
    m[929] = run?((((m[452]&~m[928]&~m[930]&~m[931]&~m[932])|(~m[452]&~m[928]&~m[930]&m[931]&~m[932])|(m[452]&m[928]&~m[930]&m[931]&~m[932])|(m[452]&~m[928]&m[930]&m[931]&~m[932])|(~m[452]&m[928]&~m[930]&~m[931]&m[932])|(~m[452]&~m[928]&m[930]&~m[931]&m[932])|(m[452]&m[928]&m[930]&~m[931]&m[932])|(~m[452]&m[928]&m[930]&m[931]&m[932]))&UnbiasedRNG[332])|((m[452]&~m[928]&~m[930]&m[931]&~m[932])|(~m[452]&~m[928]&~m[930]&~m[931]&m[932])|(m[452]&~m[928]&~m[930]&~m[931]&m[932])|(m[452]&m[928]&~m[930]&~m[931]&m[932])|(m[452]&~m[928]&m[930]&~m[931]&m[932])|(~m[452]&~m[928]&~m[930]&m[931]&m[932])|(m[452]&~m[928]&~m[930]&m[931]&m[932])|(~m[452]&m[928]&~m[930]&m[931]&m[932])|(m[452]&m[928]&~m[930]&m[931]&m[932])|(~m[452]&~m[928]&m[930]&m[931]&m[932])|(m[452]&~m[928]&m[930]&m[931]&m[932])|(m[452]&m[928]&m[930]&m[931]&m[932]))):InitCond[859];
    m[934] = run?((((m[463]&~m[933]&~m[935]&~m[936]&~m[937])|(~m[463]&~m[933]&~m[935]&m[936]&~m[937])|(m[463]&m[933]&~m[935]&m[936]&~m[937])|(m[463]&~m[933]&m[935]&m[936]&~m[937])|(~m[463]&m[933]&~m[935]&~m[936]&m[937])|(~m[463]&~m[933]&m[935]&~m[936]&m[937])|(m[463]&m[933]&m[935]&~m[936]&m[937])|(~m[463]&m[933]&m[935]&m[936]&m[937]))&UnbiasedRNG[333])|((m[463]&~m[933]&~m[935]&m[936]&~m[937])|(~m[463]&~m[933]&~m[935]&~m[936]&m[937])|(m[463]&~m[933]&~m[935]&~m[936]&m[937])|(m[463]&m[933]&~m[935]&~m[936]&m[937])|(m[463]&~m[933]&m[935]&~m[936]&m[937])|(~m[463]&~m[933]&~m[935]&m[936]&m[937])|(m[463]&~m[933]&~m[935]&m[936]&m[937])|(~m[463]&m[933]&~m[935]&m[936]&m[937])|(m[463]&m[933]&~m[935]&m[936]&m[937])|(~m[463]&~m[933]&m[935]&m[936]&m[937])|(m[463]&~m[933]&m[935]&m[936]&m[937])|(m[463]&m[933]&m[935]&m[936]&m[937]))):InitCond[860];
    m[939] = run?((((m[474]&~m[938]&~m[940]&~m[941]&~m[942])|(~m[474]&~m[938]&~m[940]&m[941]&~m[942])|(m[474]&m[938]&~m[940]&m[941]&~m[942])|(m[474]&~m[938]&m[940]&m[941]&~m[942])|(~m[474]&m[938]&~m[940]&~m[941]&m[942])|(~m[474]&~m[938]&m[940]&~m[941]&m[942])|(m[474]&m[938]&m[940]&~m[941]&m[942])|(~m[474]&m[938]&m[940]&m[941]&m[942]))&UnbiasedRNG[334])|((m[474]&~m[938]&~m[940]&m[941]&~m[942])|(~m[474]&~m[938]&~m[940]&~m[941]&m[942])|(m[474]&~m[938]&~m[940]&~m[941]&m[942])|(m[474]&m[938]&~m[940]&~m[941]&m[942])|(m[474]&~m[938]&m[940]&~m[941]&m[942])|(~m[474]&~m[938]&~m[940]&m[941]&m[942])|(m[474]&~m[938]&~m[940]&m[941]&m[942])|(~m[474]&m[938]&~m[940]&m[941]&m[942])|(m[474]&m[938]&~m[940]&m[941]&m[942])|(~m[474]&~m[938]&m[940]&m[941]&m[942])|(m[474]&~m[938]&m[940]&m[941]&m[942])|(m[474]&m[938]&m[940]&m[941]&m[942]))):InitCond[861];
    m[944] = run?((((m[485]&~m[943]&~m[945]&~m[946]&~m[947])|(~m[485]&~m[943]&~m[945]&m[946]&~m[947])|(m[485]&m[943]&~m[945]&m[946]&~m[947])|(m[485]&~m[943]&m[945]&m[946]&~m[947])|(~m[485]&m[943]&~m[945]&~m[946]&m[947])|(~m[485]&~m[943]&m[945]&~m[946]&m[947])|(m[485]&m[943]&m[945]&~m[946]&m[947])|(~m[485]&m[943]&m[945]&m[946]&m[947]))&UnbiasedRNG[335])|((m[485]&~m[943]&~m[945]&m[946]&~m[947])|(~m[485]&~m[943]&~m[945]&~m[946]&m[947])|(m[485]&~m[943]&~m[945]&~m[946]&m[947])|(m[485]&m[943]&~m[945]&~m[946]&m[947])|(m[485]&~m[943]&m[945]&~m[946]&m[947])|(~m[485]&~m[943]&~m[945]&m[946]&m[947])|(m[485]&~m[943]&~m[945]&m[946]&m[947])|(~m[485]&m[943]&~m[945]&m[946]&m[947])|(m[485]&m[943]&~m[945]&m[946]&m[947])|(~m[485]&~m[943]&m[945]&m[946]&m[947])|(m[485]&~m[943]&m[945]&m[946]&m[947])|(m[485]&m[943]&m[945]&m[946]&m[947]))):InitCond[862];
    m[949] = run?((((m[496]&~m[948]&~m[950]&~m[951]&~m[952])|(~m[496]&~m[948]&~m[950]&m[951]&~m[952])|(m[496]&m[948]&~m[950]&m[951]&~m[952])|(m[496]&~m[948]&m[950]&m[951]&~m[952])|(~m[496]&m[948]&~m[950]&~m[951]&m[952])|(~m[496]&~m[948]&m[950]&~m[951]&m[952])|(m[496]&m[948]&m[950]&~m[951]&m[952])|(~m[496]&m[948]&m[950]&m[951]&m[952]))&UnbiasedRNG[336])|((m[496]&~m[948]&~m[950]&m[951]&~m[952])|(~m[496]&~m[948]&~m[950]&~m[951]&m[952])|(m[496]&~m[948]&~m[950]&~m[951]&m[952])|(m[496]&m[948]&~m[950]&~m[951]&m[952])|(m[496]&~m[948]&m[950]&~m[951]&m[952])|(~m[496]&~m[948]&~m[950]&m[951]&m[952])|(m[496]&~m[948]&~m[950]&m[951]&m[952])|(~m[496]&m[948]&~m[950]&m[951]&m[952])|(m[496]&m[948]&~m[950]&m[951]&m[952])|(~m[496]&~m[948]&m[950]&m[951]&m[952])|(m[496]&~m[948]&m[950]&m[951]&m[952])|(m[496]&m[948]&m[950]&m[951]&m[952]))):InitCond[863];
    m[954] = run?((((m[507]&~m[953]&~m[955]&~m[956]&~m[957])|(~m[507]&~m[953]&~m[955]&m[956]&~m[957])|(m[507]&m[953]&~m[955]&m[956]&~m[957])|(m[507]&~m[953]&m[955]&m[956]&~m[957])|(~m[507]&m[953]&~m[955]&~m[956]&m[957])|(~m[507]&~m[953]&m[955]&~m[956]&m[957])|(m[507]&m[953]&m[955]&~m[956]&m[957])|(~m[507]&m[953]&m[955]&m[956]&m[957]))&UnbiasedRNG[337])|((m[507]&~m[953]&~m[955]&m[956]&~m[957])|(~m[507]&~m[953]&~m[955]&~m[956]&m[957])|(m[507]&~m[953]&~m[955]&~m[956]&m[957])|(m[507]&m[953]&~m[955]&~m[956]&m[957])|(m[507]&~m[953]&m[955]&~m[956]&m[957])|(~m[507]&~m[953]&~m[955]&m[956]&m[957])|(m[507]&~m[953]&~m[955]&m[956]&m[957])|(~m[507]&m[953]&~m[955]&m[956]&m[957])|(m[507]&m[953]&~m[955]&m[956]&m[957])|(~m[507]&~m[953]&m[955]&m[956]&m[957])|(m[507]&~m[953]&m[955]&m[956]&m[957])|(m[507]&m[953]&m[955]&m[956]&m[957]))):InitCond[864];
    m[959] = run?((((m[518]&~m[958]&~m[960]&~m[961]&~m[962])|(~m[518]&~m[958]&~m[960]&m[961]&~m[962])|(m[518]&m[958]&~m[960]&m[961]&~m[962])|(m[518]&~m[958]&m[960]&m[961]&~m[962])|(~m[518]&m[958]&~m[960]&~m[961]&m[962])|(~m[518]&~m[958]&m[960]&~m[961]&m[962])|(m[518]&m[958]&m[960]&~m[961]&m[962])|(~m[518]&m[958]&m[960]&m[961]&m[962]))&UnbiasedRNG[338])|((m[518]&~m[958]&~m[960]&m[961]&~m[962])|(~m[518]&~m[958]&~m[960]&~m[961]&m[962])|(m[518]&~m[958]&~m[960]&~m[961]&m[962])|(m[518]&m[958]&~m[960]&~m[961]&m[962])|(m[518]&~m[958]&m[960]&~m[961]&m[962])|(~m[518]&~m[958]&~m[960]&m[961]&m[962])|(m[518]&~m[958]&~m[960]&m[961]&m[962])|(~m[518]&m[958]&~m[960]&m[961]&m[962])|(m[518]&m[958]&~m[960]&m[961]&m[962])|(~m[518]&~m[958]&m[960]&m[961]&m[962])|(m[518]&~m[958]&m[960]&m[961]&m[962])|(m[518]&m[958]&m[960]&m[961]&m[962]))):InitCond[865];
    m[964] = run?((((m[431]&~m[963]&~m[965]&~m[966]&~m[967])|(~m[431]&~m[963]&~m[965]&m[966]&~m[967])|(m[431]&m[963]&~m[965]&m[966]&~m[967])|(m[431]&~m[963]&m[965]&m[966]&~m[967])|(~m[431]&m[963]&~m[965]&~m[966]&m[967])|(~m[431]&~m[963]&m[965]&~m[966]&m[967])|(m[431]&m[963]&m[965]&~m[966]&m[967])|(~m[431]&m[963]&m[965]&m[966]&m[967]))&UnbiasedRNG[339])|((m[431]&~m[963]&~m[965]&m[966]&~m[967])|(~m[431]&~m[963]&~m[965]&~m[966]&m[967])|(m[431]&~m[963]&~m[965]&~m[966]&m[967])|(m[431]&m[963]&~m[965]&~m[966]&m[967])|(m[431]&~m[963]&m[965]&~m[966]&m[967])|(~m[431]&~m[963]&~m[965]&m[966]&m[967])|(m[431]&~m[963]&~m[965]&m[966]&m[967])|(~m[431]&m[963]&~m[965]&m[966]&m[967])|(m[431]&m[963]&~m[965]&m[966]&m[967])|(~m[431]&~m[963]&m[965]&m[966]&m[967])|(m[431]&~m[963]&m[965]&m[966]&m[967])|(m[431]&m[963]&m[965]&m[966]&m[967]))):InitCond[866];
    m[969] = run?((((m[442]&~m[968]&~m[970]&~m[971]&~m[972])|(~m[442]&~m[968]&~m[970]&m[971]&~m[972])|(m[442]&m[968]&~m[970]&m[971]&~m[972])|(m[442]&~m[968]&m[970]&m[971]&~m[972])|(~m[442]&m[968]&~m[970]&~m[971]&m[972])|(~m[442]&~m[968]&m[970]&~m[971]&m[972])|(m[442]&m[968]&m[970]&~m[971]&m[972])|(~m[442]&m[968]&m[970]&m[971]&m[972]))&UnbiasedRNG[340])|((m[442]&~m[968]&~m[970]&m[971]&~m[972])|(~m[442]&~m[968]&~m[970]&~m[971]&m[972])|(m[442]&~m[968]&~m[970]&~m[971]&m[972])|(m[442]&m[968]&~m[970]&~m[971]&m[972])|(m[442]&~m[968]&m[970]&~m[971]&m[972])|(~m[442]&~m[968]&~m[970]&m[971]&m[972])|(m[442]&~m[968]&~m[970]&m[971]&m[972])|(~m[442]&m[968]&~m[970]&m[971]&m[972])|(m[442]&m[968]&~m[970]&m[971]&m[972])|(~m[442]&~m[968]&m[970]&m[971]&m[972])|(m[442]&~m[968]&m[970]&m[971]&m[972])|(m[442]&m[968]&m[970]&m[971]&m[972]))):InitCond[867];
    m[974] = run?((((m[453]&~m[973]&~m[975]&~m[976]&~m[977])|(~m[453]&~m[973]&~m[975]&m[976]&~m[977])|(m[453]&m[973]&~m[975]&m[976]&~m[977])|(m[453]&~m[973]&m[975]&m[976]&~m[977])|(~m[453]&m[973]&~m[975]&~m[976]&m[977])|(~m[453]&~m[973]&m[975]&~m[976]&m[977])|(m[453]&m[973]&m[975]&~m[976]&m[977])|(~m[453]&m[973]&m[975]&m[976]&m[977]))&UnbiasedRNG[341])|((m[453]&~m[973]&~m[975]&m[976]&~m[977])|(~m[453]&~m[973]&~m[975]&~m[976]&m[977])|(m[453]&~m[973]&~m[975]&~m[976]&m[977])|(m[453]&m[973]&~m[975]&~m[976]&m[977])|(m[453]&~m[973]&m[975]&~m[976]&m[977])|(~m[453]&~m[973]&~m[975]&m[976]&m[977])|(m[453]&~m[973]&~m[975]&m[976]&m[977])|(~m[453]&m[973]&~m[975]&m[976]&m[977])|(m[453]&m[973]&~m[975]&m[976]&m[977])|(~m[453]&~m[973]&m[975]&m[976]&m[977])|(m[453]&~m[973]&m[975]&m[976]&m[977])|(m[453]&m[973]&m[975]&m[976]&m[977]))):InitCond[868];
    m[979] = run?((((m[464]&~m[978]&~m[980]&~m[981]&~m[982])|(~m[464]&~m[978]&~m[980]&m[981]&~m[982])|(m[464]&m[978]&~m[980]&m[981]&~m[982])|(m[464]&~m[978]&m[980]&m[981]&~m[982])|(~m[464]&m[978]&~m[980]&~m[981]&m[982])|(~m[464]&~m[978]&m[980]&~m[981]&m[982])|(m[464]&m[978]&m[980]&~m[981]&m[982])|(~m[464]&m[978]&m[980]&m[981]&m[982]))&UnbiasedRNG[342])|((m[464]&~m[978]&~m[980]&m[981]&~m[982])|(~m[464]&~m[978]&~m[980]&~m[981]&m[982])|(m[464]&~m[978]&~m[980]&~m[981]&m[982])|(m[464]&m[978]&~m[980]&~m[981]&m[982])|(m[464]&~m[978]&m[980]&~m[981]&m[982])|(~m[464]&~m[978]&~m[980]&m[981]&m[982])|(m[464]&~m[978]&~m[980]&m[981]&m[982])|(~m[464]&m[978]&~m[980]&m[981]&m[982])|(m[464]&m[978]&~m[980]&m[981]&m[982])|(~m[464]&~m[978]&m[980]&m[981]&m[982])|(m[464]&~m[978]&m[980]&m[981]&m[982])|(m[464]&m[978]&m[980]&m[981]&m[982]))):InitCond[869];
    m[984] = run?((((m[475]&~m[983]&~m[985]&~m[986]&~m[987])|(~m[475]&~m[983]&~m[985]&m[986]&~m[987])|(m[475]&m[983]&~m[985]&m[986]&~m[987])|(m[475]&~m[983]&m[985]&m[986]&~m[987])|(~m[475]&m[983]&~m[985]&~m[986]&m[987])|(~m[475]&~m[983]&m[985]&~m[986]&m[987])|(m[475]&m[983]&m[985]&~m[986]&m[987])|(~m[475]&m[983]&m[985]&m[986]&m[987]))&UnbiasedRNG[343])|((m[475]&~m[983]&~m[985]&m[986]&~m[987])|(~m[475]&~m[983]&~m[985]&~m[986]&m[987])|(m[475]&~m[983]&~m[985]&~m[986]&m[987])|(m[475]&m[983]&~m[985]&~m[986]&m[987])|(m[475]&~m[983]&m[985]&~m[986]&m[987])|(~m[475]&~m[983]&~m[985]&m[986]&m[987])|(m[475]&~m[983]&~m[985]&m[986]&m[987])|(~m[475]&m[983]&~m[985]&m[986]&m[987])|(m[475]&m[983]&~m[985]&m[986]&m[987])|(~m[475]&~m[983]&m[985]&m[986]&m[987])|(m[475]&~m[983]&m[985]&m[986]&m[987])|(m[475]&m[983]&m[985]&m[986]&m[987]))):InitCond[870];
    m[989] = run?((((m[486]&~m[988]&~m[990]&~m[991]&~m[992])|(~m[486]&~m[988]&~m[990]&m[991]&~m[992])|(m[486]&m[988]&~m[990]&m[991]&~m[992])|(m[486]&~m[988]&m[990]&m[991]&~m[992])|(~m[486]&m[988]&~m[990]&~m[991]&m[992])|(~m[486]&~m[988]&m[990]&~m[991]&m[992])|(m[486]&m[988]&m[990]&~m[991]&m[992])|(~m[486]&m[988]&m[990]&m[991]&m[992]))&UnbiasedRNG[344])|((m[486]&~m[988]&~m[990]&m[991]&~m[992])|(~m[486]&~m[988]&~m[990]&~m[991]&m[992])|(m[486]&~m[988]&~m[990]&~m[991]&m[992])|(m[486]&m[988]&~m[990]&~m[991]&m[992])|(m[486]&~m[988]&m[990]&~m[991]&m[992])|(~m[486]&~m[988]&~m[990]&m[991]&m[992])|(m[486]&~m[988]&~m[990]&m[991]&m[992])|(~m[486]&m[988]&~m[990]&m[991]&m[992])|(m[486]&m[988]&~m[990]&m[991]&m[992])|(~m[486]&~m[988]&m[990]&m[991]&m[992])|(m[486]&~m[988]&m[990]&m[991]&m[992])|(m[486]&m[988]&m[990]&m[991]&m[992]))):InitCond[871];
    m[994] = run?((((m[497]&~m[993]&~m[995]&~m[996]&~m[997])|(~m[497]&~m[993]&~m[995]&m[996]&~m[997])|(m[497]&m[993]&~m[995]&m[996]&~m[997])|(m[497]&~m[993]&m[995]&m[996]&~m[997])|(~m[497]&m[993]&~m[995]&~m[996]&m[997])|(~m[497]&~m[993]&m[995]&~m[996]&m[997])|(m[497]&m[993]&m[995]&~m[996]&m[997])|(~m[497]&m[993]&m[995]&m[996]&m[997]))&UnbiasedRNG[345])|((m[497]&~m[993]&~m[995]&m[996]&~m[997])|(~m[497]&~m[993]&~m[995]&~m[996]&m[997])|(m[497]&~m[993]&~m[995]&~m[996]&m[997])|(m[497]&m[993]&~m[995]&~m[996]&m[997])|(m[497]&~m[993]&m[995]&~m[996]&m[997])|(~m[497]&~m[993]&~m[995]&m[996]&m[997])|(m[497]&~m[993]&~m[995]&m[996]&m[997])|(~m[497]&m[993]&~m[995]&m[996]&m[997])|(m[497]&m[993]&~m[995]&m[996]&m[997])|(~m[497]&~m[993]&m[995]&m[996]&m[997])|(m[497]&~m[993]&m[995]&m[996]&m[997])|(m[497]&m[993]&m[995]&m[996]&m[997]))):InitCond[872];
    m[999] = run?((((m[508]&~m[998]&~m[1000]&~m[1001]&~m[1002])|(~m[508]&~m[998]&~m[1000]&m[1001]&~m[1002])|(m[508]&m[998]&~m[1000]&m[1001]&~m[1002])|(m[508]&~m[998]&m[1000]&m[1001]&~m[1002])|(~m[508]&m[998]&~m[1000]&~m[1001]&m[1002])|(~m[508]&~m[998]&m[1000]&~m[1001]&m[1002])|(m[508]&m[998]&m[1000]&~m[1001]&m[1002])|(~m[508]&m[998]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[346])|((m[508]&~m[998]&~m[1000]&m[1001]&~m[1002])|(~m[508]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[508]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[508]&m[998]&~m[1000]&~m[1001]&m[1002])|(m[508]&~m[998]&m[1000]&~m[1001]&m[1002])|(~m[508]&~m[998]&~m[1000]&m[1001]&m[1002])|(m[508]&~m[998]&~m[1000]&m[1001]&m[1002])|(~m[508]&m[998]&~m[1000]&m[1001]&m[1002])|(m[508]&m[998]&~m[1000]&m[1001]&m[1002])|(~m[508]&~m[998]&m[1000]&m[1001]&m[1002])|(m[508]&~m[998]&m[1000]&m[1001]&m[1002])|(m[508]&m[998]&m[1000]&m[1001]&m[1002]))):InitCond[873];
    m[1004] = run?((((m[519]&~m[1003]&~m[1005]&~m[1006]&~m[1007])|(~m[519]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(m[519]&m[1003]&~m[1005]&m[1006]&~m[1007])|(m[519]&~m[1003]&m[1005]&m[1006]&~m[1007])|(~m[519]&m[1003]&~m[1005]&~m[1006]&m[1007])|(~m[519]&~m[1003]&m[1005]&~m[1006]&m[1007])|(m[519]&m[1003]&m[1005]&~m[1006]&m[1007])|(~m[519]&m[1003]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[347])|((m[519]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(~m[519]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[519]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[519]&m[1003]&~m[1005]&~m[1006]&m[1007])|(m[519]&~m[1003]&m[1005]&~m[1006]&m[1007])|(~m[519]&~m[1003]&~m[1005]&m[1006]&m[1007])|(m[519]&~m[1003]&~m[1005]&m[1006]&m[1007])|(~m[519]&m[1003]&~m[1005]&m[1006]&m[1007])|(m[519]&m[1003]&~m[1005]&m[1006]&m[1007])|(~m[519]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[519]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[519]&m[1003]&m[1005]&m[1006]&m[1007]))):InitCond[874];
    m[1009] = run?((((m[443]&~m[1008]&~m[1010]&~m[1011]&~m[1012])|(~m[443]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(m[443]&m[1008]&~m[1010]&m[1011]&~m[1012])|(m[443]&~m[1008]&m[1010]&m[1011]&~m[1012])|(~m[443]&m[1008]&~m[1010]&~m[1011]&m[1012])|(~m[443]&~m[1008]&m[1010]&~m[1011]&m[1012])|(m[443]&m[1008]&m[1010]&~m[1011]&m[1012])|(~m[443]&m[1008]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[348])|((m[443]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(~m[443]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[443]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[443]&m[1008]&~m[1010]&~m[1011]&m[1012])|(m[443]&~m[1008]&m[1010]&~m[1011]&m[1012])|(~m[443]&~m[1008]&~m[1010]&m[1011]&m[1012])|(m[443]&~m[1008]&~m[1010]&m[1011]&m[1012])|(~m[443]&m[1008]&~m[1010]&m[1011]&m[1012])|(m[443]&m[1008]&~m[1010]&m[1011]&m[1012])|(~m[443]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[443]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[443]&m[1008]&m[1010]&m[1011]&m[1012]))):InitCond[875];
    m[1014] = run?((((m[454]&~m[1013]&~m[1015]&~m[1016]&~m[1017])|(~m[454]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(m[454]&m[1013]&~m[1015]&m[1016]&~m[1017])|(m[454]&~m[1013]&m[1015]&m[1016]&~m[1017])|(~m[454]&m[1013]&~m[1015]&~m[1016]&m[1017])|(~m[454]&~m[1013]&m[1015]&~m[1016]&m[1017])|(m[454]&m[1013]&m[1015]&~m[1016]&m[1017])|(~m[454]&m[1013]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[349])|((m[454]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(~m[454]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[454]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[454]&m[1013]&~m[1015]&~m[1016]&m[1017])|(m[454]&~m[1013]&m[1015]&~m[1016]&m[1017])|(~m[454]&~m[1013]&~m[1015]&m[1016]&m[1017])|(m[454]&~m[1013]&~m[1015]&m[1016]&m[1017])|(~m[454]&m[1013]&~m[1015]&m[1016]&m[1017])|(m[454]&m[1013]&~m[1015]&m[1016]&m[1017])|(~m[454]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[454]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[454]&m[1013]&m[1015]&m[1016]&m[1017]))):InitCond[876];
    m[1019] = run?((((m[465]&~m[1018]&~m[1020]&~m[1021]&~m[1022])|(~m[465]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(m[465]&m[1018]&~m[1020]&m[1021]&~m[1022])|(m[465]&~m[1018]&m[1020]&m[1021]&~m[1022])|(~m[465]&m[1018]&~m[1020]&~m[1021]&m[1022])|(~m[465]&~m[1018]&m[1020]&~m[1021]&m[1022])|(m[465]&m[1018]&m[1020]&~m[1021]&m[1022])|(~m[465]&m[1018]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[350])|((m[465]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(~m[465]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[465]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[465]&m[1018]&~m[1020]&~m[1021]&m[1022])|(m[465]&~m[1018]&m[1020]&~m[1021]&m[1022])|(~m[465]&~m[1018]&~m[1020]&m[1021]&m[1022])|(m[465]&~m[1018]&~m[1020]&m[1021]&m[1022])|(~m[465]&m[1018]&~m[1020]&m[1021]&m[1022])|(m[465]&m[1018]&~m[1020]&m[1021]&m[1022])|(~m[465]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[465]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[465]&m[1018]&m[1020]&m[1021]&m[1022]))):InitCond[877];
    m[1024] = run?((((m[476]&~m[1023]&~m[1025]&~m[1026]&~m[1027])|(~m[476]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(m[476]&m[1023]&~m[1025]&m[1026]&~m[1027])|(m[476]&~m[1023]&m[1025]&m[1026]&~m[1027])|(~m[476]&m[1023]&~m[1025]&~m[1026]&m[1027])|(~m[476]&~m[1023]&m[1025]&~m[1026]&m[1027])|(m[476]&m[1023]&m[1025]&~m[1026]&m[1027])|(~m[476]&m[1023]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[351])|((m[476]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(~m[476]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[476]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[476]&m[1023]&~m[1025]&~m[1026]&m[1027])|(m[476]&~m[1023]&m[1025]&~m[1026]&m[1027])|(~m[476]&~m[1023]&~m[1025]&m[1026]&m[1027])|(m[476]&~m[1023]&~m[1025]&m[1026]&m[1027])|(~m[476]&m[1023]&~m[1025]&m[1026]&m[1027])|(m[476]&m[1023]&~m[1025]&m[1026]&m[1027])|(~m[476]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[476]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[476]&m[1023]&m[1025]&m[1026]&m[1027]))):InitCond[878];
    m[1029] = run?((((m[487]&~m[1028]&~m[1030]&~m[1031]&~m[1032])|(~m[487]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(m[487]&m[1028]&~m[1030]&m[1031]&~m[1032])|(m[487]&~m[1028]&m[1030]&m[1031]&~m[1032])|(~m[487]&m[1028]&~m[1030]&~m[1031]&m[1032])|(~m[487]&~m[1028]&m[1030]&~m[1031]&m[1032])|(m[487]&m[1028]&m[1030]&~m[1031]&m[1032])|(~m[487]&m[1028]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[352])|((m[487]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(~m[487]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[487]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[487]&m[1028]&~m[1030]&~m[1031]&m[1032])|(m[487]&~m[1028]&m[1030]&~m[1031]&m[1032])|(~m[487]&~m[1028]&~m[1030]&m[1031]&m[1032])|(m[487]&~m[1028]&~m[1030]&m[1031]&m[1032])|(~m[487]&m[1028]&~m[1030]&m[1031]&m[1032])|(m[487]&m[1028]&~m[1030]&m[1031]&m[1032])|(~m[487]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[487]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[487]&m[1028]&m[1030]&m[1031]&m[1032]))):InitCond[879];
    m[1034] = run?((((m[498]&~m[1033]&~m[1035]&~m[1036]&~m[1037])|(~m[498]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(m[498]&m[1033]&~m[1035]&m[1036]&~m[1037])|(m[498]&~m[1033]&m[1035]&m[1036]&~m[1037])|(~m[498]&m[1033]&~m[1035]&~m[1036]&m[1037])|(~m[498]&~m[1033]&m[1035]&~m[1036]&m[1037])|(m[498]&m[1033]&m[1035]&~m[1036]&m[1037])|(~m[498]&m[1033]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[353])|((m[498]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(~m[498]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[498]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[498]&m[1033]&~m[1035]&~m[1036]&m[1037])|(m[498]&~m[1033]&m[1035]&~m[1036]&m[1037])|(~m[498]&~m[1033]&~m[1035]&m[1036]&m[1037])|(m[498]&~m[1033]&~m[1035]&m[1036]&m[1037])|(~m[498]&m[1033]&~m[1035]&m[1036]&m[1037])|(m[498]&m[1033]&~m[1035]&m[1036]&m[1037])|(~m[498]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[498]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[498]&m[1033]&m[1035]&m[1036]&m[1037]))):InitCond[880];
    m[1039] = run?((((m[509]&~m[1038]&~m[1040]&~m[1041]&~m[1042])|(~m[509]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(m[509]&m[1038]&~m[1040]&m[1041]&~m[1042])|(m[509]&~m[1038]&m[1040]&m[1041]&~m[1042])|(~m[509]&m[1038]&~m[1040]&~m[1041]&m[1042])|(~m[509]&~m[1038]&m[1040]&~m[1041]&m[1042])|(m[509]&m[1038]&m[1040]&~m[1041]&m[1042])|(~m[509]&m[1038]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[354])|((m[509]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(~m[509]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[509]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[509]&m[1038]&~m[1040]&~m[1041]&m[1042])|(m[509]&~m[1038]&m[1040]&~m[1041]&m[1042])|(~m[509]&~m[1038]&~m[1040]&m[1041]&m[1042])|(m[509]&~m[1038]&~m[1040]&m[1041]&m[1042])|(~m[509]&m[1038]&~m[1040]&m[1041]&m[1042])|(m[509]&m[1038]&~m[1040]&m[1041]&m[1042])|(~m[509]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[509]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[509]&m[1038]&m[1040]&m[1041]&m[1042]))):InitCond[881];
    m[1044] = run?((((m[520]&~m[1043]&~m[1045]&~m[1046]&~m[1047])|(~m[520]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(m[520]&m[1043]&~m[1045]&m[1046]&~m[1047])|(m[520]&~m[1043]&m[1045]&m[1046]&~m[1047])|(~m[520]&m[1043]&~m[1045]&~m[1046]&m[1047])|(~m[520]&~m[1043]&m[1045]&~m[1046]&m[1047])|(m[520]&m[1043]&m[1045]&~m[1046]&m[1047])|(~m[520]&m[1043]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[355])|((m[520]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(~m[520]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[520]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[520]&m[1043]&~m[1045]&~m[1046]&m[1047])|(m[520]&~m[1043]&m[1045]&~m[1046]&m[1047])|(~m[520]&~m[1043]&~m[1045]&m[1046]&m[1047])|(m[520]&~m[1043]&~m[1045]&m[1046]&m[1047])|(~m[520]&m[1043]&~m[1045]&m[1046]&m[1047])|(m[520]&m[1043]&~m[1045]&m[1046]&m[1047])|(~m[520]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[520]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[520]&m[1043]&m[1045]&m[1046]&m[1047]))):InitCond[882];
    m[1049] = run?((((m[455]&~m[1048]&~m[1050]&~m[1051]&~m[1052])|(~m[455]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(m[455]&m[1048]&~m[1050]&m[1051]&~m[1052])|(m[455]&~m[1048]&m[1050]&m[1051]&~m[1052])|(~m[455]&m[1048]&~m[1050]&~m[1051]&m[1052])|(~m[455]&~m[1048]&m[1050]&~m[1051]&m[1052])|(m[455]&m[1048]&m[1050]&~m[1051]&m[1052])|(~m[455]&m[1048]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[356])|((m[455]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(~m[455]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[455]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[455]&m[1048]&~m[1050]&~m[1051]&m[1052])|(m[455]&~m[1048]&m[1050]&~m[1051]&m[1052])|(~m[455]&~m[1048]&~m[1050]&m[1051]&m[1052])|(m[455]&~m[1048]&~m[1050]&m[1051]&m[1052])|(~m[455]&m[1048]&~m[1050]&m[1051]&m[1052])|(m[455]&m[1048]&~m[1050]&m[1051]&m[1052])|(~m[455]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[455]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[455]&m[1048]&m[1050]&m[1051]&m[1052]))):InitCond[883];
    m[1054] = run?((((m[466]&~m[1053]&~m[1055]&~m[1056]&~m[1057])|(~m[466]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(m[466]&m[1053]&~m[1055]&m[1056]&~m[1057])|(m[466]&~m[1053]&m[1055]&m[1056]&~m[1057])|(~m[466]&m[1053]&~m[1055]&~m[1056]&m[1057])|(~m[466]&~m[1053]&m[1055]&~m[1056]&m[1057])|(m[466]&m[1053]&m[1055]&~m[1056]&m[1057])|(~m[466]&m[1053]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[357])|((m[466]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(~m[466]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[466]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[466]&m[1053]&~m[1055]&~m[1056]&m[1057])|(m[466]&~m[1053]&m[1055]&~m[1056]&m[1057])|(~m[466]&~m[1053]&~m[1055]&m[1056]&m[1057])|(m[466]&~m[1053]&~m[1055]&m[1056]&m[1057])|(~m[466]&m[1053]&~m[1055]&m[1056]&m[1057])|(m[466]&m[1053]&~m[1055]&m[1056]&m[1057])|(~m[466]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[466]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[466]&m[1053]&m[1055]&m[1056]&m[1057]))):InitCond[884];
    m[1059] = run?((((m[477]&~m[1058]&~m[1060]&~m[1061]&~m[1062])|(~m[477]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(m[477]&m[1058]&~m[1060]&m[1061]&~m[1062])|(m[477]&~m[1058]&m[1060]&m[1061]&~m[1062])|(~m[477]&m[1058]&~m[1060]&~m[1061]&m[1062])|(~m[477]&~m[1058]&m[1060]&~m[1061]&m[1062])|(m[477]&m[1058]&m[1060]&~m[1061]&m[1062])|(~m[477]&m[1058]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[358])|((m[477]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(~m[477]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[477]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[477]&m[1058]&~m[1060]&~m[1061]&m[1062])|(m[477]&~m[1058]&m[1060]&~m[1061]&m[1062])|(~m[477]&~m[1058]&~m[1060]&m[1061]&m[1062])|(m[477]&~m[1058]&~m[1060]&m[1061]&m[1062])|(~m[477]&m[1058]&~m[1060]&m[1061]&m[1062])|(m[477]&m[1058]&~m[1060]&m[1061]&m[1062])|(~m[477]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[477]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[477]&m[1058]&m[1060]&m[1061]&m[1062]))):InitCond[885];
    m[1064] = run?((((m[488]&~m[1063]&~m[1065]&~m[1066]&~m[1067])|(~m[488]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(m[488]&m[1063]&~m[1065]&m[1066]&~m[1067])|(m[488]&~m[1063]&m[1065]&m[1066]&~m[1067])|(~m[488]&m[1063]&~m[1065]&~m[1066]&m[1067])|(~m[488]&~m[1063]&m[1065]&~m[1066]&m[1067])|(m[488]&m[1063]&m[1065]&~m[1066]&m[1067])|(~m[488]&m[1063]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[359])|((m[488]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(~m[488]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[488]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[488]&m[1063]&~m[1065]&~m[1066]&m[1067])|(m[488]&~m[1063]&m[1065]&~m[1066]&m[1067])|(~m[488]&~m[1063]&~m[1065]&m[1066]&m[1067])|(m[488]&~m[1063]&~m[1065]&m[1066]&m[1067])|(~m[488]&m[1063]&~m[1065]&m[1066]&m[1067])|(m[488]&m[1063]&~m[1065]&m[1066]&m[1067])|(~m[488]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[488]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[488]&m[1063]&m[1065]&m[1066]&m[1067]))):InitCond[886];
    m[1069] = run?((((m[499]&~m[1068]&~m[1070]&~m[1071]&~m[1072])|(~m[499]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(m[499]&m[1068]&~m[1070]&m[1071]&~m[1072])|(m[499]&~m[1068]&m[1070]&m[1071]&~m[1072])|(~m[499]&m[1068]&~m[1070]&~m[1071]&m[1072])|(~m[499]&~m[1068]&m[1070]&~m[1071]&m[1072])|(m[499]&m[1068]&m[1070]&~m[1071]&m[1072])|(~m[499]&m[1068]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[360])|((m[499]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(~m[499]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[499]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[499]&m[1068]&~m[1070]&~m[1071]&m[1072])|(m[499]&~m[1068]&m[1070]&~m[1071]&m[1072])|(~m[499]&~m[1068]&~m[1070]&m[1071]&m[1072])|(m[499]&~m[1068]&~m[1070]&m[1071]&m[1072])|(~m[499]&m[1068]&~m[1070]&m[1071]&m[1072])|(m[499]&m[1068]&~m[1070]&m[1071]&m[1072])|(~m[499]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[499]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[499]&m[1068]&m[1070]&m[1071]&m[1072]))):InitCond[887];
    m[1074] = run?((((m[510]&~m[1073]&~m[1075]&~m[1076]&~m[1077])|(~m[510]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(m[510]&m[1073]&~m[1075]&m[1076]&~m[1077])|(m[510]&~m[1073]&m[1075]&m[1076]&~m[1077])|(~m[510]&m[1073]&~m[1075]&~m[1076]&m[1077])|(~m[510]&~m[1073]&m[1075]&~m[1076]&m[1077])|(m[510]&m[1073]&m[1075]&~m[1076]&m[1077])|(~m[510]&m[1073]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[361])|((m[510]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(~m[510]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[510]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[510]&m[1073]&~m[1075]&~m[1076]&m[1077])|(m[510]&~m[1073]&m[1075]&~m[1076]&m[1077])|(~m[510]&~m[1073]&~m[1075]&m[1076]&m[1077])|(m[510]&~m[1073]&~m[1075]&m[1076]&m[1077])|(~m[510]&m[1073]&~m[1075]&m[1076]&m[1077])|(m[510]&m[1073]&~m[1075]&m[1076]&m[1077])|(~m[510]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[510]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[510]&m[1073]&m[1075]&m[1076]&m[1077]))):InitCond[888];
    m[1079] = run?((((m[521]&~m[1078]&~m[1080]&~m[1081]&~m[1082])|(~m[521]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(m[521]&m[1078]&~m[1080]&m[1081]&~m[1082])|(m[521]&~m[1078]&m[1080]&m[1081]&~m[1082])|(~m[521]&m[1078]&~m[1080]&~m[1081]&m[1082])|(~m[521]&~m[1078]&m[1080]&~m[1081]&m[1082])|(m[521]&m[1078]&m[1080]&~m[1081]&m[1082])|(~m[521]&m[1078]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[362])|((m[521]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(~m[521]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[521]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[521]&m[1078]&~m[1080]&~m[1081]&m[1082])|(m[521]&~m[1078]&m[1080]&~m[1081]&m[1082])|(~m[521]&~m[1078]&~m[1080]&m[1081]&m[1082])|(m[521]&~m[1078]&~m[1080]&m[1081]&m[1082])|(~m[521]&m[1078]&~m[1080]&m[1081]&m[1082])|(m[521]&m[1078]&~m[1080]&m[1081]&m[1082])|(~m[521]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[521]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[521]&m[1078]&m[1080]&m[1081]&m[1082]))):InitCond[889];
    m[1084] = run?((((m[467]&~m[1083]&~m[1085]&~m[1086]&~m[1087])|(~m[467]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(m[467]&m[1083]&~m[1085]&m[1086]&~m[1087])|(m[467]&~m[1083]&m[1085]&m[1086]&~m[1087])|(~m[467]&m[1083]&~m[1085]&~m[1086]&m[1087])|(~m[467]&~m[1083]&m[1085]&~m[1086]&m[1087])|(m[467]&m[1083]&m[1085]&~m[1086]&m[1087])|(~m[467]&m[1083]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[363])|((m[467]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(~m[467]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[467]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[467]&m[1083]&~m[1085]&~m[1086]&m[1087])|(m[467]&~m[1083]&m[1085]&~m[1086]&m[1087])|(~m[467]&~m[1083]&~m[1085]&m[1086]&m[1087])|(m[467]&~m[1083]&~m[1085]&m[1086]&m[1087])|(~m[467]&m[1083]&~m[1085]&m[1086]&m[1087])|(m[467]&m[1083]&~m[1085]&m[1086]&m[1087])|(~m[467]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[467]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[467]&m[1083]&m[1085]&m[1086]&m[1087]))):InitCond[890];
    m[1089] = run?((((m[478]&~m[1088]&~m[1090]&~m[1091]&~m[1092])|(~m[478]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(m[478]&m[1088]&~m[1090]&m[1091]&~m[1092])|(m[478]&~m[1088]&m[1090]&m[1091]&~m[1092])|(~m[478]&m[1088]&~m[1090]&~m[1091]&m[1092])|(~m[478]&~m[1088]&m[1090]&~m[1091]&m[1092])|(m[478]&m[1088]&m[1090]&~m[1091]&m[1092])|(~m[478]&m[1088]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[364])|((m[478]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(~m[478]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[478]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[478]&m[1088]&~m[1090]&~m[1091]&m[1092])|(m[478]&~m[1088]&m[1090]&~m[1091]&m[1092])|(~m[478]&~m[1088]&~m[1090]&m[1091]&m[1092])|(m[478]&~m[1088]&~m[1090]&m[1091]&m[1092])|(~m[478]&m[1088]&~m[1090]&m[1091]&m[1092])|(m[478]&m[1088]&~m[1090]&m[1091]&m[1092])|(~m[478]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[478]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[478]&m[1088]&m[1090]&m[1091]&m[1092]))):InitCond[891];
    m[1094] = run?((((m[489]&~m[1093]&~m[1095]&~m[1096]&~m[1097])|(~m[489]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(m[489]&m[1093]&~m[1095]&m[1096]&~m[1097])|(m[489]&~m[1093]&m[1095]&m[1096]&~m[1097])|(~m[489]&m[1093]&~m[1095]&~m[1096]&m[1097])|(~m[489]&~m[1093]&m[1095]&~m[1096]&m[1097])|(m[489]&m[1093]&m[1095]&~m[1096]&m[1097])|(~m[489]&m[1093]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[365])|((m[489]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(~m[489]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[489]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[489]&m[1093]&~m[1095]&~m[1096]&m[1097])|(m[489]&~m[1093]&m[1095]&~m[1096]&m[1097])|(~m[489]&~m[1093]&~m[1095]&m[1096]&m[1097])|(m[489]&~m[1093]&~m[1095]&m[1096]&m[1097])|(~m[489]&m[1093]&~m[1095]&m[1096]&m[1097])|(m[489]&m[1093]&~m[1095]&m[1096]&m[1097])|(~m[489]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[489]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[489]&m[1093]&m[1095]&m[1096]&m[1097]))):InitCond[892];
    m[1099] = run?((((m[500]&~m[1098]&~m[1100]&~m[1101]&~m[1102])|(~m[500]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(m[500]&m[1098]&~m[1100]&m[1101]&~m[1102])|(m[500]&~m[1098]&m[1100]&m[1101]&~m[1102])|(~m[500]&m[1098]&~m[1100]&~m[1101]&m[1102])|(~m[500]&~m[1098]&m[1100]&~m[1101]&m[1102])|(m[500]&m[1098]&m[1100]&~m[1101]&m[1102])|(~m[500]&m[1098]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[366])|((m[500]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(~m[500]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[500]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[500]&m[1098]&~m[1100]&~m[1101]&m[1102])|(m[500]&~m[1098]&m[1100]&~m[1101]&m[1102])|(~m[500]&~m[1098]&~m[1100]&m[1101]&m[1102])|(m[500]&~m[1098]&~m[1100]&m[1101]&m[1102])|(~m[500]&m[1098]&~m[1100]&m[1101]&m[1102])|(m[500]&m[1098]&~m[1100]&m[1101]&m[1102])|(~m[500]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[500]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[500]&m[1098]&m[1100]&m[1101]&m[1102]))):InitCond[893];
    m[1104] = run?((((m[511]&~m[1103]&~m[1105]&~m[1106]&~m[1107])|(~m[511]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(m[511]&m[1103]&~m[1105]&m[1106]&~m[1107])|(m[511]&~m[1103]&m[1105]&m[1106]&~m[1107])|(~m[511]&m[1103]&~m[1105]&~m[1106]&m[1107])|(~m[511]&~m[1103]&m[1105]&~m[1106]&m[1107])|(m[511]&m[1103]&m[1105]&~m[1106]&m[1107])|(~m[511]&m[1103]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[367])|((m[511]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(~m[511]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[511]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[511]&m[1103]&~m[1105]&~m[1106]&m[1107])|(m[511]&~m[1103]&m[1105]&~m[1106]&m[1107])|(~m[511]&~m[1103]&~m[1105]&m[1106]&m[1107])|(m[511]&~m[1103]&~m[1105]&m[1106]&m[1107])|(~m[511]&m[1103]&~m[1105]&m[1106]&m[1107])|(m[511]&m[1103]&~m[1105]&m[1106]&m[1107])|(~m[511]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[511]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[511]&m[1103]&m[1105]&m[1106]&m[1107]))):InitCond[894];
    m[1109] = run?((((m[522]&~m[1108]&~m[1110]&~m[1111]&~m[1112])|(~m[522]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(m[522]&m[1108]&~m[1110]&m[1111]&~m[1112])|(m[522]&~m[1108]&m[1110]&m[1111]&~m[1112])|(~m[522]&m[1108]&~m[1110]&~m[1111]&m[1112])|(~m[522]&~m[1108]&m[1110]&~m[1111]&m[1112])|(m[522]&m[1108]&m[1110]&~m[1111]&m[1112])|(~m[522]&m[1108]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[368])|((m[522]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(~m[522]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[522]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[522]&m[1108]&~m[1110]&~m[1111]&m[1112])|(m[522]&~m[1108]&m[1110]&~m[1111]&m[1112])|(~m[522]&~m[1108]&~m[1110]&m[1111]&m[1112])|(m[522]&~m[1108]&~m[1110]&m[1111]&m[1112])|(~m[522]&m[1108]&~m[1110]&m[1111]&m[1112])|(m[522]&m[1108]&~m[1110]&m[1111]&m[1112])|(~m[522]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[522]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[522]&m[1108]&m[1110]&m[1111]&m[1112]))):InitCond[895];
    m[1114] = run?((((m[479]&~m[1113]&~m[1115]&~m[1116]&~m[1117])|(~m[479]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(m[479]&m[1113]&~m[1115]&m[1116]&~m[1117])|(m[479]&~m[1113]&m[1115]&m[1116]&~m[1117])|(~m[479]&m[1113]&~m[1115]&~m[1116]&m[1117])|(~m[479]&~m[1113]&m[1115]&~m[1116]&m[1117])|(m[479]&m[1113]&m[1115]&~m[1116]&m[1117])|(~m[479]&m[1113]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[369])|((m[479]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(~m[479]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[479]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[479]&m[1113]&~m[1115]&~m[1116]&m[1117])|(m[479]&~m[1113]&m[1115]&~m[1116]&m[1117])|(~m[479]&~m[1113]&~m[1115]&m[1116]&m[1117])|(m[479]&~m[1113]&~m[1115]&m[1116]&m[1117])|(~m[479]&m[1113]&~m[1115]&m[1116]&m[1117])|(m[479]&m[1113]&~m[1115]&m[1116]&m[1117])|(~m[479]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[479]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[479]&m[1113]&m[1115]&m[1116]&m[1117]))):InitCond[896];
    m[1119] = run?((((m[490]&~m[1118]&~m[1120]&~m[1121]&~m[1122])|(~m[490]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(m[490]&m[1118]&~m[1120]&m[1121]&~m[1122])|(m[490]&~m[1118]&m[1120]&m[1121]&~m[1122])|(~m[490]&m[1118]&~m[1120]&~m[1121]&m[1122])|(~m[490]&~m[1118]&m[1120]&~m[1121]&m[1122])|(m[490]&m[1118]&m[1120]&~m[1121]&m[1122])|(~m[490]&m[1118]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[370])|((m[490]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(~m[490]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[490]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[490]&m[1118]&~m[1120]&~m[1121]&m[1122])|(m[490]&~m[1118]&m[1120]&~m[1121]&m[1122])|(~m[490]&~m[1118]&~m[1120]&m[1121]&m[1122])|(m[490]&~m[1118]&~m[1120]&m[1121]&m[1122])|(~m[490]&m[1118]&~m[1120]&m[1121]&m[1122])|(m[490]&m[1118]&~m[1120]&m[1121]&m[1122])|(~m[490]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[490]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[490]&m[1118]&m[1120]&m[1121]&m[1122]))):InitCond[897];
    m[1124] = run?((((m[501]&~m[1123]&~m[1125]&~m[1126]&~m[1127])|(~m[501]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(m[501]&m[1123]&~m[1125]&m[1126]&~m[1127])|(m[501]&~m[1123]&m[1125]&m[1126]&~m[1127])|(~m[501]&m[1123]&~m[1125]&~m[1126]&m[1127])|(~m[501]&~m[1123]&m[1125]&~m[1126]&m[1127])|(m[501]&m[1123]&m[1125]&~m[1126]&m[1127])|(~m[501]&m[1123]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[371])|((m[501]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(~m[501]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[501]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[501]&m[1123]&~m[1125]&~m[1126]&m[1127])|(m[501]&~m[1123]&m[1125]&~m[1126]&m[1127])|(~m[501]&~m[1123]&~m[1125]&m[1126]&m[1127])|(m[501]&~m[1123]&~m[1125]&m[1126]&m[1127])|(~m[501]&m[1123]&~m[1125]&m[1126]&m[1127])|(m[501]&m[1123]&~m[1125]&m[1126]&m[1127])|(~m[501]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[501]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[501]&m[1123]&m[1125]&m[1126]&m[1127]))):InitCond[898];
    m[1129] = run?((((m[512]&~m[1128]&~m[1130]&~m[1131]&~m[1132])|(~m[512]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(m[512]&m[1128]&~m[1130]&m[1131]&~m[1132])|(m[512]&~m[1128]&m[1130]&m[1131]&~m[1132])|(~m[512]&m[1128]&~m[1130]&~m[1131]&m[1132])|(~m[512]&~m[1128]&m[1130]&~m[1131]&m[1132])|(m[512]&m[1128]&m[1130]&~m[1131]&m[1132])|(~m[512]&m[1128]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[372])|((m[512]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(~m[512]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[512]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[512]&m[1128]&~m[1130]&~m[1131]&m[1132])|(m[512]&~m[1128]&m[1130]&~m[1131]&m[1132])|(~m[512]&~m[1128]&~m[1130]&m[1131]&m[1132])|(m[512]&~m[1128]&~m[1130]&m[1131]&m[1132])|(~m[512]&m[1128]&~m[1130]&m[1131]&m[1132])|(m[512]&m[1128]&~m[1130]&m[1131]&m[1132])|(~m[512]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[512]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[512]&m[1128]&m[1130]&m[1131]&m[1132]))):InitCond[899];
    m[1134] = run?((((m[523]&~m[1133]&~m[1135]&~m[1136]&~m[1137])|(~m[523]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(m[523]&m[1133]&~m[1135]&m[1136]&~m[1137])|(m[523]&~m[1133]&m[1135]&m[1136]&~m[1137])|(~m[523]&m[1133]&~m[1135]&~m[1136]&m[1137])|(~m[523]&~m[1133]&m[1135]&~m[1136]&m[1137])|(m[523]&m[1133]&m[1135]&~m[1136]&m[1137])|(~m[523]&m[1133]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[373])|((m[523]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(~m[523]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[523]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[523]&m[1133]&~m[1135]&~m[1136]&m[1137])|(m[523]&~m[1133]&m[1135]&~m[1136]&m[1137])|(~m[523]&~m[1133]&~m[1135]&m[1136]&m[1137])|(m[523]&~m[1133]&~m[1135]&m[1136]&m[1137])|(~m[523]&m[1133]&~m[1135]&m[1136]&m[1137])|(m[523]&m[1133]&~m[1135]&m[1136]&m[1137])|(~m[523]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[523]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[523]&m[1133]&m[1135]&m[1136]&m[1137]))):InitCond[900];
    m[1139] = run?((((m[491]&~m[1138]&~m[1140]&~m[1141]&~m[1142])|(~m[491]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(m[491]&m[1138]&~m[1140]&m[1141]&~m[1142])|(m[491]&~m[1138]&m[1140]&m[1141]&~m[1142])|(~m[491]&m[1138]&~m[1140]&~m[1141]&m[1142])|(~m[491]&~m[1138]&m[1140]&~m[1141]&m[1142])|(m[491]&m[1138]&m[1140]&~m[1141]&m[1142])|(~m[491]&m[1138]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[374])|((m[491]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(~m[491]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[491]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[491]&m[1138]&~m[1140]&~m[1141]&m[1142])|(m[491]&~m[1138]&m[1140]&~m[1141]&m[1142])|(~m[491]&~m[1138]&~m[1140]&m[1141]&m[1142])|(m[491]&~m[1138]&~m[1140]&m[1141]&m[1142])|(~m[491]&m[1138]&~m[1140]&m[1141]&m[1142])|(m[491]&m[1138]&~m[1140]&m[1141]&m[1142])|(~m[491]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[491]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[491]&m[1138]&m[1140]&m[1141]&m[1142]))):InitCond[901];
    m[1144] = run?((((m[502]&~m[1143]&~m[1145]&~m[1146]&~m[1147])|(~m[502]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(m[502]&m[1143]&~m[1145]&m[1146]&~m[1147])|(m[502]&~m[1143]&m[1145]&m[1146]&~m[1147])|(~m[502]&m[1143]&~m[1145]&~m[1146]&m[1147])|(~m[502]&~m[1143]&m[1145]&~m[1146]&m[1147])|(m[502]&m[1143]&m[1145]&~m[1146]&m[1147])|(~m[502]&m[1143]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[375])|((m[502]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(~m[502]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[502]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[502]&m[1143]&~m[1145]&~m[1146]&m[1147])|(m[502]&~m[1143]&m[1145]&~m[1146]&m[1147])|(~m[502]&~m[1143]&~m[1145]&m[1146]&m[1147])|(m[502]&~m[1143]&~m[1145]&m[1146]&m[1147])|(~m[502]&m[1143]&~m[1145]&m[1146]&m[1147])|(m[502]&m[1143]&~m[1145]&m[1146]&m[1147])|(~m[502]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[502]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[502]&m[1143]&m[1145]&m[1146]&m[1147]))):InitCond[902];
    m[1149] = run?((((m[513]&~m[1148]&~m[1150]&~m[1151]&~m[1152])|(~m[513]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(m[513]&m[1148]&~m[1150]&m[1151]&~m[1152])|(m[513]&~m[1148]&m[1150]&m[1151]&~m[1152])|(~m[513]&m[1148]&~m[1150]&~m[1151]&m[1152])|(~m[513]&~m[1148]&m[1150]&~m[1151]&m[1152])|(m[513]&m[1148]&m[1150]&~m[1151]&m[1152])|(~m[513]&m[1148]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[376])|((m[513]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(~m[513]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[513]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[513]&m[1148]&~m[1150]&~m[1151]&m[1152])|(m[513]&~m[1148]&m[1150]&~m[1151]&m[1152])|(~m[513]&~m[1148]&~m[1150]&m[1151]&m[1152])|(m[513]&~m[1148]&~m[1150]&m[1151]&m[1152])|(~m[513]&m[1148]&~m[1150]&m[1151]&m[1152])|(m[513]&m[1148]&~m[1150]&m[1151]&m[1152])|(~m[513]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[513]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[513]&m[1148]&m[1150]&m[1151]&m[1152]))):InitCond[903];
    m[1154] = run?((((m[524]&~m[1153]&~m[1155]&~m[1156]&~m[1157])|(~m[524]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(m[524]&m[1153]&~m[1155]&m[1156]&~m[1157])|(m[524]&~m[1153]&m[1155]&m[1156]&~m[1157])|(~m[524]&m[1153]&~m[1155]&~m[1156]&m[1157])|(~m[524]&~m[1153]&m[1155]&~m[1156]&m[1157])|(m[524]&m[1153]&m[1155]&~m[1156]&m[1157])|(~m[524]&m[1153]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[377])|((m[524]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(~m[524]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[524]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[524]&m[1153]&~m[1155]&~m[1156]&m[1157])|(m[524]&~m[1153]&m[1155]&~m[1156]&m[1157])|(~m[524]&~m[1153]&~m[1155]&m[1156]&m[1157])|(m[524]&~m[1153]&~m[1155]&m[1156]&m[1157])|(~m[524]&m[1153]&~m[1155]&m[1156]&m[1157])|(m[524]&m[1153]&~m[1155]&m[1156]&m[1157])|(~m[524]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[524]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[524]&m[1153]&m[1155]&m[1156]&m[1157]))):InitCond[904];
    m[1159] = run?((((m[503]&~m[1158]&~m[1160]&~m[1161]&~m[1162])|(~m[503]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(m[503]&m[1158]&~m[1160]&m[1161]&~m[1162])|(m[503]&~m[1158]&m[1160]&m[1161]&~m[1162])|(~m[503]&m[1158]&~m[1160]&~m[1161]&m[1162])|(~m[503]&~m[1158]&m[1160]&~m[1161]&m[1162])|(m[503]&m[1158]&m[1160]&~m[1161]&m[1162])|(~m[503]&m[1158]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[378])|((m[503]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(~m[503]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[503]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[503]&m[1158]&~m[1160]&~m[1161]&m[1162])|(m[503]&~m[1158]&m[1160]&~m[1161]&m[1162])|(~m[503]&~m[1158]&~m[1160]&m[1161]&m[1162])|(m[503]&~m[1158]&~m[1160]&m[1161]&m[1162])|(~m[503]&m[1158]&~m[1160]&m[1161]&m[1162])|(m[503]&m[1158]&~m[1160]&m[1161]&m[1162])|(~m[503]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[503]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[503]&m[1158]&m[1160]&m[1161]&m[1162]))):InitCond[905];
    m[1164] = run?((((m[514]&~m[1163]&~m[1165]&~m[1166]&~m[1167])|(~m[514]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(m[514]&m[1163]&~m[1165]&m[1166]&~m[1167])|(m[514]&~m[1163]&m[1165]&m[1166]&~m[1167])|(~m[514]&m[1163]&~m[1165]&~m[1166]&m[1167])|(~m[514]&~m[1163]&m[1165]&~m[1166]&m[1167])|(m[514]&m[1163]&m[1165]&~m[1166]&m[1167])|(~m[514]&m[1163]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[379])|((m[514]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(~m[514]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[514]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[514]&m[1163]&~m[1165]&~m[1166]&m[1167])|(m[514]&~m[1163]&m[1165]&~m[1166]&m[1167])|(~m[514]&~m[1163]&~m[1165]&m[1166]&m[1167])|(m[514]&~m[1163]&~m[1165]&m[1166]&m[1167])|(~m[514]&m[1163]&~m[1165]&m[1166]&m[1167])|(m[514]&m[1163]&~m[1165]&m[1166]&m[1167])|(~m[514]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[514]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[514]&m[1163]&m[1165]&m[1166]&m[1167]))):InitCond[906];
    m[1169] = run?((((m[525]&~m[1168]&~m[1170]&~m[1171]&~m[1172])|(~m[525]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(m[525]&m[1168]&~m[1170]&m[1171]&~m[1172])|(m[525]&~m[1168]&m[1170]&m[1171]&~m[1172])|(~m[525]&m[1168]&~m[1170]&~m[1171]&m[1172])|(~m[525]&~m[1168]&m[1170]&~m[1171]&m[1172])|(m[525]&m[1168]&m[1170]&~m[1171]&m[1172])|(~m[525]&m[1168]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[380])|((m[525]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(~m[525]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[525]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[525]&m[1168]&~m[1170]&~m[1171]&m[1172])|(m[525]&~m[1168]&m[1170]&~m[1171]&m[1172])|(~m[525]&~m[1168]&~m[1170]&m[1171]&m[1172])|(m[525]&~m[1168]&~m[1170]&m[1171]&m[1172])|(~m[525]&m[1168]&~m[1170]&m[1171]&m[1172])|(m[525]&m[1168]&~m[1170]&m[1171]&m[1172])|(~m[525]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[525]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[525]&m[1168]&m[1170]&m[1171]&m[1172]))):InitCond[907];
    m[1174] = run?((((m[515]&~m[1173]&~m[1175]&~m[1176]&~m[1177])|(~m[515]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(m[515]&m[1173]&~m[1175]&m[1176]&~m[1177])|(m[515]&~m[1173]&m[1175]&m[1176]&~m[1177])|(~m[515]&m[1173]&~m[1175]&~m[1176]&m[1177])|(~m[515]&~m[1173]&m[1175]&~m[1176]&m[1177])|(m[515]&m[1173]&m[1175]&~m[1176]&m[1177])|(~m[515]&m[1173]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[381])|((m[515]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(~m[515]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[515]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[515]&m[1173]&~m[1175]&~m[1176]&m[1177])|(m[515]&~m[1173]&m[1175]&~m[1176]&m[1177])|(~m[515]&~m[1173]&~m[1175]&m[1176]&m[1177])|(m[515]&~m[1173]&~m[1175]&m[1176]&m[1177])|(~m[515]&m[1173]&~m[1175]&m[1176]&m[1177])|(m[515]&m[1173]&~m[1175]&m[1176]&m[1177])|(~m[515]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[515]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[515]&m[1173]&m[1175]&m[1176]&m[1177]))):InitCond[908];
    m[1179] = run?((((m[526]&~m[1178]&~m[1180]&~m[1181]&~m[1182])|(~m[526]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(m[526]&m[1178]&~m[1180]&m[1181]&~m[1182])|(m[526]&~m[1178]&m[1180]&m[1181]&~m[1182])|(~m[526]&m[1178]&~m[1180]&~m[1181]&m[1182])|(~m[526]&~m[1178]&m[1180]&~m[1181]&m[1182])|(m[526]&m[1178]&m[1180]&~m[1181]&m[1182])|(~m[526]&m[1178]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[382])|((m[526]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(~m[526]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[526]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[526]&m[1178]&~m[1180]&~m[1181]&m[1182])|(m[526]&~m[1178]&m[1180]&~m[1181]&m[1182])|(~m[526]&~m[1178]&~m[1180]&m[1181]&m[1182])|(m[526]&~m[1178]&~m[1180]&m[1181]&m[1182])|(~m[526]&m[1178]&~m[1180]&m[1181]&m[1182])|(m[526]&m[1178]&~m[1180]&m[1181]&m[1182])|(~m[526]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[526]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[526]&m[1178]&m[1180]&m[1181]&m[1182]))):InitCond[909];
    m[1184] = run?((((m[527]&~m[1183]&~m[1185]&~m[1186]&~m[1187])|(~m[527]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(m[527]&m[1183]&~m[1185]&m[1186]&~m[1187])|(m[527]&~m[1183]&m[1185]&m[1186]&~m[1187])|(~m[527]&m[1183]&~m[1185]&~m[1186]&m[1187])|(~m[527]&~m[1183]&m[1185]&~m[1186]&m[1187])|(m[527]&m[1183]&m[1185]&~m[1186]&m[1187])|(~m[527]&m[1183]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[383])|((m[527]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(~m[527]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[527]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[527]&m[1183]&~m[1185]&~m[1186]&m[1187])|(m[527]&~m[1183]&m[1185]&~m[1186]&m[1187])|(~m[527]&~m[1183]&~m[1185]&m[1186]&m[1187])|(m[527]&~m[1183]&~m[1185]&m[1186]&m[1187])|(~m[527]&m[1183]&~m[1185]&m[1186]&m[1187])|(m[527]&m[1183]&~m[1185]&m[1186]&m[1187])|(~m[527]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[527]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[527]&m[1183]&m[1185]&m[1186]&m[1187]))):InitCond[910];
end

always @(posedge color3_clk) begin
    m[536] = run?((((m[533]&~m[534]&~m[535]&~m[537]&~m[538])|(~m[533]&m[534]&~m[535]&~m[537]&~m[538])|(~m[533]&~m[534]&m[535]&~m[537]&~m[538])|(m[533]&m[534]&m[535]&m[537]&~m[538])|(~m[533]&~m[534]&~m[535]&~m[537]&m[538])|(m[533]&m[534]&~m[535]&m[537]&m[538])|(m[533]&~m[534]&m[535]&m[537]&m[538])|(~m[533]&m[534]&m[535]&m[537]&m[538]))&UnbiasedRNG[384])|((m[533]&m[534]&~m[535]&~m[537]&~m[538])|(m[533]&~m[534]&m[535]&~m[537]&~m[538])|(~m[533]&m[534]&m[535]&~m[537]&~m[538])|(m[533]&m[534]&m[535]&~m[537]&~m[538])|(m[533]&~m[534]&~m[535]&~m[537]&m[538])|(~m[533]&m[534]&~m[535]&~m[537]&m[538])|(m[533]&m[534]&~m[535]&~m[537]&m[538])|(~m[533]&~m[534]&m[535]&~m[537]&m[538])|(m[533]&~m[534]&m[535]&~m[537]&m[538])|(~m[533]&m[534]&m[535]&~m[537]&m[538])|(m[533]&m[534]&m[535]&~m[537]&m[538])|(m[533]&m[534]&m[535]&m[537]&m[538]))):InitCond[911];
    m[546] = run?((((m[543]&~m[544]&~m[545]&~m[547]&~m[548])|(~m[543]&m[544]&~m[545]&~m[547]&~m[548])|(~m[543]&~m[544]&m[545]&~m[547]&~m[548])|(m[543]&m[544]&m[545]&m[547]&~m[548])|(~m[543]&~m[544]&~m[545]&~m[547]&m[548])|(m[543]&m[544]&~m[545]&m[547]&m[548])|(m[543]&~m[544]&m[545]&m[547]&m[548])|(~m[543]&m[544]&m[545]&m[547]&m[548]))&UnbiasedRNG[385])|((m[543]&m[544]&~m[545]&~m[547]&~m[548])|(m[543]&~m[544]&m[545]&~m[547]&~m[548])|(~m[543]&m[544]&m[545]&~m[547]&~m[548])|(m[543]&m[544]&m[545]&~m[547]&~m[548])|(m[543]&~m[544]&~m[545]&~m[547]&m[548])|(~m[543]&m[544]&~m[545]&~m[547]&m[548])|(m[543]&m[544]&~m[545]&~m[547]&m[548])|(~m[543]&~m[544]&m[545]&~m[547]&m[548])|(m[543]&~m[544]&m[545]&~m[547]&m[548])|(~m[543]&m[544]&m[545]&~m[547]&m[548])|(m[543]&m[544]&m[545]&~m[547]&m[548])|(m[543]&m[544]&m[545]&m[547]&m[548]))):InitCond[912];
    m[551] = run?((((m[548]&~m[549]&~m[550]&~m[552]&~m[553])|(~m[548]&m[549]&~m[550]&~m[552]&~m[553])|(~m[548]&~m[549]&m[550]&~m[552]&~m[553])|(m[548]&m[549]&m[550]&m[552]&~m[553])|(~m[548]&~m[549]&~m[550]&~m[552]&m[553])|(m[548]&m[549]&~m[550]&m[552]&m[553])|(m[548]&~m[549]&m[550]&m[552]&m[553])|(~m[548]&m[549]&m[550]&m[552]&m[553]))&UnbiasedRNG[386])|((m[548]&m[549]&~m[550]&~m[552]&~m[553])|(m[548]&~m[549]&m[550]&~m[552]&~m[553])|(~m[548]&m[549]&m[550]&~m[552]&~m[553])|(m[548]&m[549]&m[550]&~m[552]&~m[553])|(m[548]&~m[549]&~m[550]&~m[552]&m[553])|(~m[548]&m[549]&~m[550]&~m[552]&m[553])|(m[548]&m[549]&~m[550]&~m[552]&m[553])|(~m[548]&~m[549]&m[550]&~m[552]&m[553])|(m[548]&~m[549]&m[550]&~m[552]&m[553])|(~m[548]&m[549]&m[550]&~m[552]&m[553])|(m[548]&m[549]&m[550]&~m[552]&m[553])|(m[548]&m[549]&m[550]&m[552]&m[553]))):InitCond[913];
    m[561] = run?((((m[558]&~m[559]&~m[560]&~m[562]&~m[563])|(~m[558]&m[559]&~m[560]&~m[562]&~m[563])|(~m[558]&~m[559]&m[560]&~m[562]&~m[563])|(m[558]&m[559]&m[560]&m[562]&~m[563])|(~m[558]&~m[559]&~m[560]&~m[562]&m[563])|(m[558]&m[559]&~m[560]&m[562]&m[563])|(m[558]&~m[559]&m[560]&m[562]&m[563])|(~m[558]&m[559]&m[560]&m[562]&m[563]))&UnbiasedRNG[387])|((m[558]&m[559]&~m[560]&~m[562]&~m[563])|(m[558]&~m[559]&m[560]&~m[562]&~m[563])|(~m[558]&m[559]&m[560]&~m[562]&~m[563])|(m[558]&m[559]&m[560]&~m[562]&~m[563])|(m[558]&~m[559]&~m[560]&~m[562]&m[563])|(~m[558]&m[559]&~m[560]&~m[562]&m[563])|(m[558]&m[559]&~m[560]&~m[562]&m[563])|(~m[558]&~m[559]&m[560]&~m[562]&m[563])|(m[558]&~m[559]&m[560]&~m[562]&m[563])|(~m[558]&m[559]&m[560]&~m[562]&m[563])|(m[558]&m[559]&m[560]&~m[562]&m[563])|(m[558]&m[559]&m[560]&m[562]&m[563]))):InitCond[914];
    m[566] = run?((((m[563]&~m[564]&~m[565]&~m[567]&~m[568])|(~m[563]&m[564]&~m[565]&~m[567]&~m[568])|(~m[563]&~m[564]&m[565]&~m[567]&~m[568])|(m[563]&m[564]&m[565]&m[567]&~m[568])|(~m[563]&~m[564]&~m[565]&~m[567]&m[568])|(m[563]&m[564]&~m[565]&m[567]&m[568])|(m[563]&~m[564]&m[565]&m[567]&m[568])|(~m[563]&m[564]&m[565]&m[567]&m[568]))&UnbiasedRNG[388])|((m[563]&m[564]&~m[565]&~m[567]&~m[568])|(m[563]&~m[564]&m[565]&~m[567]&~m[568])|(~m[563]&m[564]&m[565]&~m[567]&~m[568])|(m[563]&m[564]&m[565]&~m[567]&~m[568])|(m[563]&~m[564]&~m[565]&~m[567]&m[568])|(~m[563]&m[564]&~m[565]&~m[567]&m[568])|(m[563]&m[564]&~m[565]&~m[567]&m[568])|(~m[563]&~m[564]&m[565]&~m[567]&m[568])|(m[563]&~m[564]&m[565]&~m[567]&m[568])|(~m[563]&m[564]&m[565]&~m[567]&m[568])|(m[563]&m[564]&m[565]&~m[567]&m[568])|(m[563]&m[564]&m[565]&m[567]&m[568]))):InitCond[915];
    m[571] = run?((((m[568]&~m[569]&~m[570]&~m[572]&~m[573])|(~m[568]&m[569]&~m[570]&~m[572]&~m[573])|(~m[568]&~m[569]&m[570]&~m[572]&~m[573])|(m[568]&m[569]&m[570]&m[572]&~m[573])|(~m[568]&~m[569]&~m[570]&~m[572]&m[573])|(m[568]&m[569]&~m[570]&m[572]&m[573])|(m[568]&~m[569]&m[570]&m[572]&m[573])|(~m[568]&m[569]&m[570]&m[572]&m[573]))&UnbiasedRNG[389])|((m[568]&m[569]&~m[570]&~m[572]&~m[573])|(m[568]&~m[569]&m[570]&~m[572]&~m[573])|(~m[568]&m[569]&m[570]&~m[572]&~m[573])|(m[568]&m[569]&m[570]&~m[572]&~m[573])|(m[568]&~m[569]&~m[570]&~m[572]&m[573])|(~m[568]&m[569]&~m[570]&~m[572]&m[573])|(m[568]&m[569]&~m[570]&~m[572]&m[573])|(~m[568]&~m[569]&m[570]&~m[572]&m[573])|(m[568]&~m[569]&m[570]&~m[572]&m[573])|(~m[568]&m[569]&m[570]&~m[572]&m[573])|(m[568]&m[569]&m[570]&~m[572]&m[573])|(m[568]&m[569]&m[570]&m[572]&m[573]))):InitCond[916];
    m[581] = run?((((m[578]&~m[579]&~m[580]&~m[582]&~m[583])|(~m[578]&m[579]&~m[580]&~m[582]&~m[583])|(~m[578]&~m[579]&m[580]&~m[582]&~m[583])|(m[578]&m[579]&m[580]&m[582]&~m[583])|(~m[578]&~m[579]&~m[580]&~m[582]&m[583])|(m[578]&m[579]&~m[580]&m[582]&m[583])|(m[578]&~m[579]&m[580]&m[582]&m[583])|(~m[578]&m[579]&m[580]&m[582]&m[583]))&UnbiasedRNG[390])|((m[578]&m[579]&~m[580]&~m[582]&~m[583])|(m[578]&~m[579]&m[580]&~m[582]&~m[583])|(~m[578]&m[579]&m[580]&~m[582]&~m[583])|(m[578]&m[579]&m[580]&~m[582]&~m[583])|(m[578]&~m[579]&~m[580]&~m[582]&m[583])|(~m[578]&m[579]&~m[580]&~m[582]&m[583])|(m[578]&m[579]&~m[580]&~m[582]&m[583])|(~m[578]&~m[579]&m[580]&~m[582]&m[583])|(m[578]&~m[579]&m[580]&~m[582]&m[583])|(~m[578]&m[579]&m[580]&~m[582]&m[583])|(m[578]&m[579]&m[580]&~m[582]&m[583])|(m[578]&m[579]&m[580]&m[582]&m[583]))):InitCond[917];
    m[586] = run?((((m[583]&~m[584]&~m[585]&~m[587]&~m[588])|(~m[583]&m[584]&~m[585]&~m[587]&~m[588])|(~m[583]&~m[584]&m[585]&~m[587]&~m[588])|(m[583]&m[584]&m[585]&m[587]&~m[588])|(~m[583]&~m[584]&~m[585]&~m[587]&m[588])|(m[583]&m[584]&~m[585]&m[587]&m[588])|(m[583]&~m[584]&m[585]&m[587]&m[588])|(~m[583]&m[584]&m[585]&m[587]&m[588]))&UnbiasedRNG[391])|((m[583]&m[584]&~m[585]&~m[587]&~m[588])|(m[583]&~m[584]&m[585]&~m[587]&~m[588])|(~m[583]&m[584]&m[585]&~m[587]&~m[588])|(m[583]&m[584]&m[585]&~m[587]&~m[588])|(m[583]&~m[584]&~m[585]&~m[587]&m[588])|(~m[583]&m[584]&~m[585]&~m[587]&m[588])|(m[583]&m[584]&~m[585]&~m[587]&m[588])|(~m[583]&~m[584]&m[585]&~m[587]&m[588])|(m[583]&~m[584]&m[585]&~m[587]&m[588])|(~m[583]&m[584]&m[585]&~m[587]&m[588])|(m[583]&m[584]&m[585]&~m[587]&m[588])|(m[583]&m[584]&m[585]&m[587]&m[588]))):InitCond[918];
    m[591] = run?((((m[588]&~m[589]&~m[590]&~m[592]&~m[593])|(~m[588]&m[589]&~m[590]&~m[592]&~m[593])|(~m[588]&~m[589]&m[590]&~m[592]&~m[593])|(m[588]&m[589]&m[590]&m[592]&~m[593])|(~m[588]&~m[589]&~m[590]&~m[592]&m[593])|(m[588]&m[589]&~m[590]&m[592]&m[593])|(m[588]&~m[589]&m[590]&m[592]&m[593])|(~m[588]&m[589]&m[590]&m[592]&m[593]))&UnbiasedRNG[392])|((m[588]&m[589]&~m[590]&~m[592]&~m[593])|(m[588]&~m[589]&m[590]&~m[592]&~m[593])|(~m[588]&m[589]&m[590]&~m[592]&~m[593])|(m[588]&m[589]&m[590]&~m[592]&~m[593])|(m[588]&~m[589]&~m[590]&~m[592]&m[593])|(~m[588]&m[589]&~m[590]&~m[592]&m[593])|(m[588]&m[589]&~m[590]&~m[592]&m[593])|(~m[588]&~m[589]&m[590]&~m[592]&m[593])|(m[588]&~m[589]&m[590]&~m[592]&m[593])|(~m[588]&m[589]&m[590]&~m[592]&m[593])|(m[588]&m[589]&m[590]&~m[592]&m[593])|(m[588]&m[589]&m[590]&m[592]&m[593]))):InitCond[919];
    m[596] = run?((((m[593]&~m[594]&~m[595]&~m[597]&~m[598])|(~m[593]&m[594]&~m[595]&~m[597]&~m[598])|(~m[593]&~m[594]&m[595]&~m[597]&~m[598])|(m[593]&m[594]&m[595]&m[597]&~m[598])|(~m[593]&~m[594]&~m[595]&~m[597]&m[598])|(m[593]&m[594]&~m[595]&m[597]&m[598])|(m[593]&~m[594]&m[595]&m[597]&m[598])|(~m[593]&m[594]&m[595]&m[597]&m[598]))&UnbiasedRNG[393])|((m[593]&m[594]&~m[595]&~m[597]&~m[598])|(m[593]&~m[594]&m[595]&~m[597]&~m[598])|(~m[593]&m[594]&m[595]&~m[597]&~m[598])|(m[593]&m[594]&m[595]&~m[597]&~m[598])|(m[593]&~m[594]&~m[595]&~m[597]&m[598])|(~m[593]&m[594]&~m[595]&~m[597]&m[598])|(m[593]&m[594]&~m[595]&~m[597]&m[598])|(~m[593]&~m[594]&m[595]&~m[597]&m[598])|(m[593]&~m[594]&m[595]&~m[597]&m[598])|(~m[593]&m[594]&m[595]&~m[597]&m[598])|(m[593]&m[594]&m[595]&~m[597]&m[598])|(m[593]&m[594]&m[595]&m[597]&m[598]))):InitCond[920];
    m[606] = run?((((m[603]&~m[604]&~m[605]&~m[607]&~m[608])|(~m[603]&m[604]&~m[605]&~m[607]&~m[608])|(~m[603]&~m[604]&m[605]&~m[607]&~m[608])|(m[603]&m[604]&m[605]&m[607]&~m[608])|(~m[603]&~m[604]&~m[605]&~m[607]&m[608])|(m[603]&m[604]&~m[605]&m[607]&m[608])|(m[603]&~m[604]&m[605]&m[607]&m[608])|(~m[603]&m[604]&m[605]&m[607]&m[608]))&UnbiasedRNG[394])|((m[603]&m[604]&~m[605]&~m[607]&~m[608])|(m[603]&~m[604]&m[605]&~m[607]&~m[608])|(~m[603]&m[604]&m[605]&~m[607]&~m[608])|(m[603]&m[604]&m[605]&~m[607]&~m[608])|(m[603]&~m[604]&~m[605]&~m[607]&m[608])|(~m[603]&m[604]&~m[605]&~m[607]&m[608])|(m[603]&m[604]&~m[605]&~m[607]&m[608])|(~m[603]&~m[604]&m[605]&~m[607]&m[608])|(m[603]&~m[604]&m[605]&~m[607]&m[608])|(~m[603]&m[604]&m[605]&~m[607]&m[608])|(m[603]&m[604]&m[605]&~m[607]&m[608])|(m[603]&m[604]&m[605]&m[607]&m[608]))):InitCond[921];
    m[611] = run?((((m[608]&~m[609]&~m[610]&~m[612]&~m[613])|(~m[608]&m[609]&~m[610]&~m[612]&~m[613])|(~m[608]&~m[609]&m[610]&~m[612]&~m[613])|(m[608]&m[609]&m[610]&m[612]&~m[613])|(~m[608]&~m[609]&~m[610]&~m[612]&m[613])|(m[608]&m[609]&~m[610]&m[612]&m[613])|(m[608]&~m[609]&m[610]&m[612]&m[613])|(~m[608]&m[609]&m[610]&m[612]&m[613]))&UnbiasedRNG[395])|((m[608]&m[609]&~m[610]&~m[612]&~m[613])|(m[608]&~m[609]&m[610]&~m[612]&~m[613])|(~m[608]&m[609]&m[610]&~m[612]&~m[613])|(m[608]&m[609]&m[610]&~m[612]&~m[613])|(m[608]&~m[609]&~m[610]&~m[612]&m[613])|(~m[608]&m[609]&~m[610]&~m[612]&m[613])|(m[608]&m[609]&~m[610]&~m[612]&m[613])|(~m[608]&~m[609]&m[610]&~m[612]&m[613])|(m[608]&~m[609]&m[610]&~m[612]&m[613])|(~m[608]&m[609]&m[610]&~m[612]&m[613])|(m[608]&m[609]&m[610]&~m[612]&m[613])|(m[608]&m[609]&m[610]&m[612]&m[613]))):InitCond[922];
    m[616] = run?((((m[613]&~m[614]&~m[615]&~m[617]&~m[618])|(~m[613]&m[614]&~m[615]&~m[617]&~m[618])|(~m[613]&~m[614]&m[615]&~m[617]&~m[618])|(m[613]&m[614]&m[615]&m[617]&~m[618])|(~m[613]&~m[614]&~m[615]&~m[617]&m[618])|(m[613]&m[614]&~m[615]&m[617]&m[618])|(m[613]&~m[614]&m[615]&m[617]&m[618])|(~m[613]&m[614]&m[615]&m[617]&m[618]))&UnbiasedRNG[396])|((m[613]&m[614]&~m[615]&~m[617]&~m[618])|(m[613]&~m[614]&m[615]&~m[617]&~m[618])|(~m[613]&m[614]&m[615]&~m[617]&~m[618])|(m[613]&m[614]&m[615]&~m[617]&~m[618])|(m[613]&~m[614]&~m[615]&~m[617]&m[618])|(~m[613]&m[614]&~m[615]&~m[617]&m[618])|(m[613]&m[614]&~m[615]&~m[617]&m[618])|(~m[613]&~m[614]&m[615]&~m[617]&m[618])|(m[613]&~m[614]&m[615]&~m[617]&m[618])|(~m[613]&m[614]&m[615]&~m[617]&m[618])|(m[613]&m[614]&m[615]&~m[617]&m[618])|(m[613]&m[614]&m[615]&m[617]&m[618]))):InitCond[923];
    m[621] = run?((((m[618]&~m[619]&~m[620]&~m[622]&~m[623])|(~m[618]&m[619]&~m[620]&~m[622]&~m[623])|(~m[618]&~m[619]&m[620]&~m[622]&~m[623])|(m[618]&m[619]&m[620]&m[622]&~m[623])|(~m[618]&~m[619]&~m[620]&~m[622]&m[623])|(m[618]&m[619]&~m[620]&m[622]&m[623])|(m[618]&~m[619]&m[620]&m[622]&m[623])|(~m[618]&m[619]&m[620]&m[622]&m[623]))&UnbiasedRNG[397])|((m[618]&m[619]&~m[620]&~m[622]&~m[623])|(m[618]&~m[619]&m[620]&~m[622]&~m[623])|(~m[618]&m[619]&m[620]&~m[622]&~m[623])|(m[618]&m[619]&m[620]&~m[622]&~m[623])|(m[618]&~m[619]&~m[620]&~m[622]&m[623])|(~m[618]&m[619]&~m[620]&~m[622]&m[623])|(m[618]&m[619]&~m[620]&~m[622]&m[623])|(~m[618]&~m[619]&m[620]&~m[622]&m[623])|(m[618]&~m[619]&m[620]&~m[622]&m[623])|(~m[618]&m[619]&m[620]&~m[622]&m[623])|(m[618]&m[619]&m[620]&~m[622]&m[623])|(m[618]&m[619]&m[620]&m[622]&m[623]))):InitCond[924];
    m[626] = run?((((m[623]&~m[624]&~m[625]&~m[627]&~m[628])|(~m[623]&m[624]&~m[625]&~m[627]&~m[628])|(~m[623]&~m[624]&m[625]&~m[627]&~m[628])|(m[623]&m[624]&m[625]&m[627]&~m[628])|(~m[623]&~m[624]&~m[625]&~m[627]&m[628])|(m[623]&m[624]&~m[625]&m[627]&m[628])|(m[623]&~m[624]&m[625]&m[627]&m[628])|(~m[623]&m[624]&m[625]&m[627]&m[628]))&UnbiasedRNG[398])|((m[623]&m[624]&~m[625]&~m[627]&~m[628])|(m[623]&~m[624]&m[625]&~m[627]&~m[628])|(~m[623]&m[624]&m[625]&~m[627]&~m[628])|(m[623]&m[624]&m[625]&~m[627]&~m[628])|(m[623]&~m[624]&~m[625]&~m[627]&m[628])|(~m[623]&m[624]&~m[625]&~m[627]&m[628])|(m[623]&m[624]&~m[625]&~m[627]&m[628])|(~m[623]&~m[624]&m[625]&~m[627]&m[628])|(m[623]&~m[624]&m[625]&~m[627]&m[628])|(~m[623]&m[624]&m[625]&~m[627]&m[628])|(m[623]&m[624]&m[625]&~m[627]&m[628])|(m[623]&m[624]&m[625]&m[627]&m[628]))):InitCond[925];
    m[636] = run?((((m[633]&~m[634]&~m[635]&~m[637]&~m[638])|(~m[633]&m[634]&~m[635]&~m[637]&~m[638])|(~m[633]&~m[634]&m[635]&~m[637]&~m[638])|(m[633]&m[634]&m[635]&m[637]&~m[638])|(~m[633]&~m[634]&~m[635]&~m[637]&m[638])|(m[633]&m[634]&~m[635]&m[637]&m[638])|(m[633]&~m[634]&m[635]&m[637]&m[638])|(~m[633]&m[634]&m[635]&m[637]&m[638]))&UnbiasedRNG[399])|((m[633]&m[634]&~m[635]&~m[637]&~m[638])|(m[633]&~m[634]&m[635]&~m[637]&~m[638])|(~m[633]&m[634]&m[635]&~m[637]&~m[638])|(m[633]&m[634]&m[635]&~m[637]&~m[638])|(m[633]&~m[634]&~m[635]&~m[637]&m[638])|(~m[633]&m[634]&~m[635]&~m[637]&m[638])|(m[633]&m[634]&~m[635]&~m[637]&m[638])|(~m[633]&~m[634]&m[635]&~m[637]&m[638])|(m[633]&~m[634]&m[635]&~m[637]&m[638])|(~m[633]&m[634]&m[635]&~m[637]&m[638])|(m[633]&m[634]&m[635]&~m[637]&m[638])|(m[633]&m[634]&m[635]&m[637]&m[638]))):InitCond[926];
    m[641] = run?((((m[638]&~m[639]&~m[640]&~m[642]&~m[643])|(~m[638]&m[639]&~m[640]&~m[642]&~m[643])|(~m[638]&~m[639]&m[640]&~m[642]&~m[643])|(m[638]&m[639]&m[640]&m[642]&~m[643])|(~m[638]&~m[639]&~m[640]&~m[642]&m[643])|(m[638]&m[639]&~m[640]&m[642]&m[643])|(m[638]&~m[639]&m[640]&m[642]&m[643])|(~m[638]&m[639]&m[640]&m[642]&m[643]))&UnbiasedRNG[400])|((m[638]&m[639]&~m[640]&~m[642]&~m[643])|(m[638]&~m[639]&m[640]&~m[642]&~m[643])|(~m[638]&m[639]&m[640]&~m[642]&~m[643])|(m[638]&m[639]&m[640]&~m[642]&~m[643])|(m[638]&~m[639]&~m[640]&~m[642]&m[643])|(~m[638]&m[639]&~m[640]&~m[642]&m[643])|(m[638]&m[639]&~m[640]&~m[642]&m[643])|(~m[638]&~m[639]&m[640]&~m[642]&m[643])|(m[638]&~m[639]&m[640]&~m[642]&m[643])|(~m[638]&m[639]&m[640]&~m[642]&m[643])|(m[638]&m[639]&m[640]&~m[642]&m[643])|(m[638]&m[639]&m[640]&m[642]&m[643]))):InitCond[927];
    m[646] = run?((((m[643]&~m[644]&~m[645]&~m[647]&~m[648])|(~m[643]&m[644]&~m[645]&~m[647]&~m[648])|(~m[643]&~m[644]&m[645]&~m[647]&~m[648])|(m[643]&m[644]&m[645]&m[647]&~m[648])|(~m[643]&~m[644]&~m[645]&~m[647]&m[648])|(m[643]&m[644]&~m[645]&m[647]&m[648])|(m[643]&~m[644]&m[645]&m[647]&m[648])|(~m[643]&m[644]&m[645]&m[647]&m[648]))&UnbiasedRNG[401])|((m[643]&m[644]&~m[645]&~m[647]&~m[648])|(m[643]&~m[644]&m[645]&~m[647]&~m[648])|(~m[643]&m[644]&m[645]&~m[647]&~m[648])|(m[643]&m[644]&m[645]&~m[647]&~m[648])|(m[643]&~m[644]&~m[645]&~m[647]&m[648])|(~m[643]&m[644]&~m[645]&~m[647]&m[648])|(m[643]&m[644]&~m[645]&~m[647]&m[648])|(~m[643]&~m[644]&m[645]&~m[647]&m[648])|(m[643]&~m[644]&m[645]&~m[647]&m[648])|(~m[643]&m[644]&m[645]&~m[647]&m[648])|(m[643]&m[644]&m[645]&~m[647]&m[648])|(m[643]&m[644]&m[645]&m[647]&m[648]))):InitCond[928];
    m[651] = run?((((m[648]&~m[649]&~m[650]&~m[652]&~m[653])|(~m[648]&m[649]&~m[650]&~m[652]&~m[653])|(~m[648]&~m[649]&m[650]&~m[652]&~m[653])|(m[648]&m[649]&m[650]&m[652]&~m[653])|(~m[648]&~m[649]&~m[650]&~m[652]&m[653])|(m[648]&m[649]&~m[650]&m[652]&m[653])|(m[648]&~m[649]&m[650]&m[652]&m[653])|(~m[648]&m[649]&m[650]&m[652]&m[653]))&UnbiasedRNG[402])|((m[648]&m[649]&~m[650]&~m[652]&~m[653])|(m[648]&~m[649]&m[650]&~m[652]&~m[653])|(~m[648]&m[649]&m[650]&~m[652]&~m[653])|(m[648]&m[649]&m[650]&~m[652]&~m[653])|(m[648]&~m[649]&~m[650]&~m[652]&m[653])|(~m[648]&m[649]&~m[650]&~m[652]&m[653])|(m[648]&m[649]&~m[650]&~m[652]&m[653])|(~m[648]&~m[649]&m[650]&~m[652]&m[653])|(m[648]&~m[649]&m[650]&~m[652]&m[653])|(~m[648]&m[649]&m[650]&~m[652]&m[653])|(m[648]&m[649]&m[650]&~m[652]&m[653])|(m[648]&m[649]&m[650]&m[652]&m[653]))):InitCond[929];
    m[656] = run?((((m[653]&~m[654]&~m[655]&~m[657]&~m[658])|(~m[653]&m[654]&~m[655]&~m[657]&~m[658])|(~m[653]&~m[654]&m[655]&~m[657]&~m[658])|(m[653]&m[654]&m[655]&m[657]&~m[658])|(~m[653]&~m[654]&~m[655]&~m[657]&m[658])|(m[653]&m[654]&~m[655]&m[657]&m[658])|(m[653]&~m[654]&m[655]&m[657]&m[658])|(~m[653]&m[654]&m[655]&m[657]&m[658]))&UnbiasedRNG[403])|((m[653]&m[654]&~m[655]&~m[657]&~m[658])|(m[653]&~m[654]&m[655]&~m[657]&~m[658])|(~m[653]&m[654]&m[655]&~m[657]&~m[658])|(m[653]&m[654]&m[655]&~m[657]&~m[658])|(m[653]&~m[654]&~m[655]&~m[657]&m[658])|(~m[653]&m[654]&~m[655]&~m[657]&m[658])|(m[653]&m[654]&~m[655]&~m[657]&m[658])|(~m[653]&~m[654]&m[655]&~m[657]&m[658])|(m[653]&~m[654]&m[655]&~m[657]&m[658])|(~m[653]&m[654]&m[655]&~m[657]&m[658])|(m[653]&m[654]&m[655]&~m[657]&m[658])|(m[653]&m[654]&m[655]&m[657]&m[658]))):InitCond[930];
    m[661] = run?((((m[658]&~m[659]&~m[660]&~m[662]&~m[663])|(~m[658]&m[659]&~m[660]&~m[662]&~m[663])|(~m[658]&~m[659]&m[660]&~m[662]&~m[663])|(m[658]&m[659]&m[660]&m[662]&~m[663])|(~m[658]&~m[659]&~m[660]&~m[662]&m[663])|(m[658]&m[659]&~m[660]&m[662]&m[663])|(m[658]&~m[659]&m[660]&m[662]&m[663])|(~m[658]&m[659]&m[660]&m[662]&m[663]))&UnbiasedRNG[404])|((m[658]&m[659]&~m[660]&~m[662]&~m[663])|(m[658]&~m[659]&m[660]&~m[662]&~m[663])|(~m[658]&m[659]&m[660]&~m[662]&~m[663])|(m[658]&m[659]&m[660]&~m[662]&~m[663])|(m[658]&~m[659]&~m[660]&~m[662]&m[663])|(~m[658]&m[659]&~m[660]&~m[662]&m[663])|(m[658]&m[659]&~m[660]&~m[662]&m[663])|(~m[658]&~m[659]&m[660]&~m[662]&m[663])|(m[658]&~m[659]&m[660]&~m[662]&m[663])|(~m[658]&m[659]&m[660]&~m[662]&m[663])|(m[658]&m[659]&m[660]&~m[662]&m[663])|(m[658]&m[659]&m[660]&m[662]&m[663]))):InitCond[931];
    m[671] = run?((((m[668]&~m[669]&~m[670]&~m[672]&~m[673])|(~m[668]&m[669]&~m[670]&~m[672]&~m[673])|(~m[668]&~m[669]&m[670]&~m[672]&~m[673])|(m[668]&m[669]&m[670]&m[672]&~m[673])|(~m[668]&~m[669]&~m[670]&~m[672]&m[673])|(m[668]&m[669]&~m[670]&m[672]&m[673])|(m[668]&~m[669]&m[670]&m[672]&m[673])|(~m[668]&m[669]&m[670]&m[672]&m[673]))&UnbiasedRNG[405])|((m[668]&m[669]&~m[670]&~m[672]&~m[673])|(m[668]&~m[669]&m[670]&~m[672]&~m[673])|(~m[668]&m[669]&m[670]&~m[672]&~m[673])|(m[668]&m[669]&m[670]&~m[672]&~m[673])|(m[668]&~m[669]&~m[670]&~m[672]&m[673])|(~m[668]&m[669]&~m[670]&~m[672]&m[673])|(m[668]&m[669]&~m[670]&~m[672]&m[673])|(~m[668]&~m[669]&m[670]&~m[672]&m[673])|(m[668]&~m[669]&m[670]&~m[672]&m[673])|(~m[668]&m[669]&m[670]&~m[672]&m[673])|(m[668]&m[669]&m[670]&~m[672]&m[673])|(m[668]&m[669]&m[670]&m[672]&m[673]))):InitCond[932];
    m[676] = run?((((m[673]&~m[674]&~m[675]&~m[677]&~m[678])|(~m[673]&m[674]&~m[675]&~m[677]&~m[678])|(~m[673]&~m[674]&m[675]&~m[677]&~m[678])|(m[673]&m[674]&m[675]&m[677]&~m[678])|(~m[673]&~m[674]&~m[675]&~m[677]&m[678])|(m[673]&m[674]&~m[675]&m[677]&m[678])|(m[673]&~m[674]&m[675]&m[677]&m[678])|(~m[673]&m[674]&m[675]&m[677]&m[678]))&UnbiasedRNG[406])|((m[673]&m[674]&~m[675]&~m[677]&~m[678])|(m[673]&~m[674]&m[675]&~m[677]&~m[678])|(~m[673]&m[674]&m[675]&~m[677]&~m[678])|(m[673]&m[674]&m[675]&~m[677]&~m[678])|(m[673]&~m[674]&~m[675]&~m[677]&m[678])|(~m[673]&m[674]&~m[675]&~m[677]&m[678])|(m[673]&m[674]&~m[675]&~m[677]&m[678])|(~m[673]&~m[674]&m[675]&~m[677]&m[678])|(m[673]&~m[674]&m[675]&~m[677]&m[678])|(~m[673]&m[674]&m[675]&~m[677]&m[678])|(m[673]&m[674]&m[675]&~m[677]&m[678])|(m[673]&m[674]&m[675]&m[677]&m[678]))):InitCond[933];
    m[681] = run?((((m[678]&~m[679]&~m[680]&~m[682]&~m[683])|(~m[678]&m[679]&~m[680]&~m[682]&~m[683])|(~m[678]&~m[679]&m[680]&~m[682]&~m[683])|(m[678]&m[679]&m[680]&m[682]&~m[683])|(~m[678]&~m[679]&~m[680]&~m[682]&m[683])|(m[678]&m[679]&~m[680]&m[682]&m[683])|(m[678]&~m[679]&m[680]&m[682]&m[683])|(~m[678]&m[679]&m[680]&m[682]&m[683]))&UnbiasedRNG[407])|((m[678]&m[679]&~m[680]&~m[682]&~m[683])|(m[678]&~m[679]&m[680]&~m[682]&~m[683])|(~m[678]&m[679]&m[680]&~m[682]&~m[683])|(m[678]&m[679]&m[680]&~m[682]&~m[683])|(m[678]&~m[679]&~m[680]&~m[682]&m[683])|(~m[678]&m[679]&~m[680]&~m[682]&m[683])|(m[678]&m[679]&~m[680]&~m[682]&m[683])|(~m[678]&~m[679]&m[680]&~m[682]&m[683])|(m[678]&~m[679]&m[680]&~m[682]&m[683])|(~m[678]&m[679]&m[680]&~m[682]&m[683])|(m[678]&m[679]&m[680]&~m[682]&m[683])|(m[678]&m[679]&m[680]&m[682]&m[683]))):InitCond[934];
    m[686] = run?((((m[683]&~m[684]&~m[685]&~m[687]&~m[688])|(~m[683]&m[684]&~m[685]&~m[687]&~m[688])|(~m[683]&~m[684]&m[685]&~m[687]&~m[688])|(m[683]&m[684]&m[685]&m[687]&~m[688])|(~m[683]&~m[684]&~m[685]&~m[687]&m[688])|(m[683]&m[684]&~m[685]&m[687]&m[688])|(m[683]&~m[684]&m[685]&m[687]&m[688])|(~m[683]&m[684]&m[685]&m[687]&m[688]))&UnbiasedRNG[408])|((m[683]&m[684]&~m[685]&~m[687]&~m[688])|(m[683]&~m[684]&m[685]&~m[687]&~m[688])|(~m[683]&m[684]&m[685]&~m[687]&~m[688])|(m[683]&m[684]&m[685]&~m[687]&~m[688])|(m[683]&~m[684]&~m[685]&~m[687]&m[688])|(~m[683]&m[684]&~m[685]&~m[687]&m[688])|(m[683]&m[684]&~m[685]&~m[687]&m[688])|(~m[683]&~m[684]&m[685]&~m[687]&m[688])|(m[683]&~m[684]&m[685]&~m[687]&m[688])|(~m[683]&m[684]&m[685]&~m[687]&m[688])|(m[683]&m[684]&m[685]&~m[687]&m[688])|(m[683]&m[684]&m[685]&m[687]&m[688]))):InitCond[935];
    m[691] = run?((((m[688]&~m[689]&~m[690]&~m[692]&~m[693])|(~m[688]&m[689]&~m[690]&~m[692]&~m[693])|(~m[688]&~m[689]&m[690]&~m[692]&~m[693])|(m[688]&m[689]&m[690]&m[692]&~m[693])|(~m[688]&~m[689]&~m[690]&~m[692]&m[693])|(m[688]&m[689]&~m[690]&m[692]&m[693])|(m[688]&~m[689]&m[690]&m[692]&m[693])|(~m[688]&m[689]&m[690]&m[692]&m[693]))&UnbiasedRNG[409])|((m[688]&m[689]&~m[690]&~m[692]&~m[693])|(m[688]&~m[689]&m[690]&~m[692]&~m[693])|(~m[688]&m[689]&m[690]&~m[692]&~m[693])|(m[688]&m[689]&m[690]&~m[692]&~m[693])|(m[688]&~m[689]&~m[690]&~m[692]&m[693])|(~m[688]&m[689]&~m[690]&~m[692]&m[693])|(m[688]&m[689]&~m[690]&~m[692]&m[693])|(~m[688]&~m[689]&m[690]&~m[692]&m[693])|(m[688]&~m[689]&m[690]&~m[692]&m[693])|(~m[688]&m[689]&m[690]&~m[692]&m[693])|(m[688]&m[689]&m[690]&~m[692]&m[693])|(m[688]&m[689]&m[690]&m[692]&m[693]))):InitCond[936];
    m[696] = run?((((m[693]&~m[694]&~m[695]&~m[697]&~m[698])|(~m[693]&m[694]&~m[695]&~m[697]&~m[698])|(~m[693]&~m[694]&m[695]&~m[697]&~m[698])|(m[693]&m[694]&m[695]&m[697]&~m[698])|(~m[693]&~m[694]&~m[695]&~m[697]&m[698])|(m[693]&m[694]&~m[695]&m[697]&m[698])|(m[693]&~m[694]&m[695]&m[697]&m[698])|(~m[693]&m[694]&m[695]&m[697]&m[698]))&UnbiasedRNG[410])|((m[693]&m[694]&~m[695]&~m[697]&~m[698])|(m[693]&~m[694]&m[695]&~m[697]&~m[698])|(~m[693]&m[694]&m[695]&~m[697]&~m[698])|(m[693]&m[694]&m[695]&~m[697]&~m[698])|(m[693]&~m[694]&~m[695]&~m[697]&m[698])|(~m[693]&m[694]&~m[695]&~m[697]&m[698])|(m[693]&m[694]&~m[695]&~m[697]&m[698])|(~m[693]&~m[694]&m[695]&~m[697]&m[698])|(m[693]&~m[694]&m[695]&~m[697]&m[698])|(~m[693]&m[694]&m[695]&~m[697]&m[698])|(m[693]&m[694]&m[695]&~m[697]&m[698])|(m[693]&m[694]&m[695]&m[697]&m[698]))):InitCond[937];
    m[701] = run?((((m[698]&~m[699]&~m[700]&~m[702]&~m[703])|(~m[698]&m[699]&~m[700]&~m[702]&~m[703])|(~m[698]&~m[699]&m[700]&~m[702]&~m[703])|(m[698]&m[699]&m[700]&m[702]&~m[703])|(~m[698]&~m[699]&~m[700]&~m[702]&m[703])|(m[698]&m[699]&~m[700]&m[702]&m[703])|(m[698]&~m[699]&m[700]&m[702]&m[703])|(~m[698]&m[699]&m[700]&m[702]&m[703]))&UnbiasedRNG[411])|((m[698]&m[699]&~m[700]&~m[702]&~m[703])|(m[698]&~m[699]&m[700]&~m[702]&~m[703])|(~m[698]&m[699]&m[700]&~m[702]&~m[703])|(m[698]&m[699]&m[700]&~m[702]&~m[703])|(m[698]&~m[699]&~m[700]&~m[702]&m[703])|(~m[698]&m[699]&~m[700]&~m[702]&m[703])|(m[698]&m[699]&~m[700]&~m[702]&m[703])|(~m[698]&~m[699]&m[700]&~m[702]&m[703])|(m[698]&~m[699]&m[700]&~m[702]&m[703])|(~m[698]&m[699]&m[700]&~m[702]&m[703])|(m[698]&m[699]&m[700]&~m[702]&m[703])|(m[698]&m[699]&m[700]&m[702]&m[703]))):InitCond[938];
    m[711] = run?((((m[708]&~m[709]&~m[710]&~m[712]&~m[713])|(~m[708]&m[709]&~m[710]&~m[712]&~m[713])|(~m[708]&~m[709]&m[710]&~m[712]&~m[713])|(m[708]&m[709]&m[710]&m[712]&~m[713])|(~m[708]&~m[709]&~m[710]&~m[712]&m[713])|(m[708]&m[709]&~m[710]&m[712]&m[713])|(m[708]&~m[709]&m[710]&m[712]&m[713])|(~m[708]&m[709]&m[710]&m[712]&m[713]))&UnbiasedRNG[412])|((m[708]&m[709]&~m[710]&~m[712]&~m[713])|(m[708]&~m[709]&m[710]&~m[712]&~m[713])|(~m[708]&m[709]&m[710]&~m[712]&~m[713])|(m[708]&m[709]&m[710]&~m[712]&~m[713])|(m[708]&~m[709]&~m[710]&~m[712]&m[713])|(~m[708]&m[709]&~m[710]&~m[712]&m[713])|(m[708]&m[709]&~m[710]&~m[712]&m[713])|(~m[708]&~m[709]&m[710]&~m[712]&m[713])|(m[708]&~m[709]&m[710]&~m[712]&m[713])|(~m[708]&m[709]&m[710]&~m[712]&m[713])|(m[708]&m[709]&m[710]&~m[712]&m[713])|(m[708]&m[709]&m[710]&m[712]&m[713]))):InitCond[939];
    m[716] = run?((((m[713]&~m[714]&~m[715]&~m[717]&~m[718])|(~m[713]&m[714]&~m[715]&~m[717]&~m[718])|(~m[713]&~m[714]&m[715]&~m[717]&~m[718])|(m[713]&m[714]&m[715]&m[717]&~m[718])|(~m[713]&~m[714]&~m[715]&~m[717]&m[718])|(m[713]&m[714]&~m[715]&m[717]&m[718])|(m[713]&~m[714]&m[715]&m[717]&m[718])|(~m[713]&m[714]&m[715]&m[717]&m[718]))&UnbiasedRNG[413])|((m[713]&m[714]&~m[715]&~m[717]&~m[718])|(m[713]&~m[714]&m[715]&~m[717]&~m[718])|(~m[713]&m[714]&m[715]&~m[717]&~m[718])|(m[713]&m[714]&m[715]&~m[717]&~m[718])|(m[713]&~m[714]&~m[715]&~m[717]&m[718])|(~m[713]&m[714]&~m[715]&~m[717]&m[718])|(m[713]&m[714]&~m[715]&~m[717]&m[718])|(~m[713]&~m[714]&m[715]&~m[717]&m[718])|(m[713]&~m[714]&m[715]&~m[717]&m[718])|(~m[713]&m[714]&m[715]&~m[717]&m[718])|(m[713]&m[714]&m[715]&~m[717]&m[718])|(m[713]&m[714]&m[715]&m[717]&m[718]))):InitCond[940];
    m[721] = run?((((m[718]&~m[719]&~m[720]&~m[722]&~m[723])|(~m[718]&m[719]&~m[720]&~m[722]&~m[723])|(~m[718]&~m[719]&m[720]&~m[722]&~m[723])|(m[718]&m[719]&m[720]&m[722]&~m[723])|(~m[718]&~m[719]&~m[720]&~m[722]&m[723])|(m[718]&m[719]&~m[720]&m[722]&m[723])|(m[718]&~m[719]&m[720]&m[722]&m[723])|(~m[718]&m[719]&m[720]&m[722]&m[723]))&UnbiasedRNG[414])|((m[718]&m[719]&~m[720]&~m[722]&~m[723])|(m[718]&~m[719]&m[720]&~m[722]&~m[723])|(~m[718]&m[719]&m[720]&~m[722]&~m[723])|(m[718]&m[719]&m[720]&~m[722]&~m[723])|(m[718]&~m[719]&~m[720]&~m[722]&m[723])|(~m[718]&m[719]&~m[720]&~m[722]&m[723])|(m[718]&m[719]&~m[720]&~m[722]&m[723])|(~m[718]&~m[719]&m[720]&~m[722]&m[723])|(m[718]&~m[719]&m[720]&~m[722]&m[723])|(~m[718]&m[719]&m[720]&~m[722]&m[723])|(m[718]&m[719]&m[720]&~m[722]&m[723])|(m[718]&m[719]&m[720]&m[722]&m[723]))):InitCond[941];
    m[726] = run?((((m[723]&~m[724]&~m[725]&~m[727]&~m[728])|(~m[723]&m[724]&~m[725]&~m[727]&~m[728])|(~m[723]&~m[724]&m[725]&~m[727]&~m[728])|(m[723]&m[724]&m[725]&m[727]&~m[728])|(~m[723]&~m[724]&~m[725]&~m[727]&m[728])|(m[723]&m[724]&~m[725]&m[727]&m[728])|(m[723]&~m[724]&m[725]&m[727]&m[728])|(~m[723]&m[724]&m[725]&m[727]&m[728]))&UnbiasedRNG[415])|((m[723]&m[724]&~m[725]&~m[727]&~m[728])|(m[723]&~m[724]&m[725]&~m[727]&~m[728])|(~m[723]&m[724]&m[725]&~m[727]&~m[728])|(m[723]&m[724]&m[725]&~m[727]&~m[728])|(m[723]&~m[724]&~m[725]&~m[727]&m[728])|(~m[723]&m[724]&~m[725]&~m[727]&m[728])|(m[723]&m[724]&~m[725]&~m[727]&m[728])|(~m[723]&~m[724]&m[725]&~m[727]&m[728])|(m[723]&~m[724]&m[725]&~m[727]&m[728])|(~m[723]&m[724]&m[725]&~m[727]&m[728])|(m[723]&m[724]&m[725]&~m[727]&m[728])|(m[723]&m[724]&m[725]&m[727]&m[728]))):InitCond[942];
    m[731] = run?((((m[728]&~m[729]&~m[730]&~m[732]&~m[733])|(~m[728]&m[729]&~m[730]&~m[732]&~m[733])|(~m[728]&~m[729]&m[730]&~m[732]&~m[733])|(m[728]&m[729]&m[730]&m[732]&~m[733])|(~m[728]&~m[729]&~m[730]&~m[732]&m[733])|(m[728]&m[729]&~m[730]&m[732]&m[733])|(m[728]&~m[729]&m[730]&m[732]&m[733])|(~m[728]&m[729]&m[730]&m[732]&m[733]))&UnbiasedRNG[416])|((m[728]&m[729]&~m[730]&~m[732]&~m[733])|(m[728]&~m[729]&m[730]&~m[732]&~m[733])|(~m[728]&m[729]&m[730]&~m[732]&~m[733])|(m[728]&m[729]&m[730]&~m[732]&~m[733])|(m[728]&~m[729]&~m[730]&~m[732]&m[733])|(~m[728]&m[729]&~m[730]&~m[732]&m[733])|(m[728]&m[729]&~m[730]&~m[732]&m[733])|(~m[728]&~m[729]&m[730]&~m[732]&m[733])|(m[728]&~m[729]&m[730]&~m[732]&m[733])|(~m[728]&m[729]&m[730]&~m[732]&m[733])|(m[728]&m[729]&m[730]&~m[732]&m[733])|(m[728]&m[729]&m[730]&m[732]&m[733]))):InitCond[943];
    m[736] = run?((((m[733]&~m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&~m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&m[737]&~m[738])|(~m[733]&~m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&m[737]&m[738])|(m[733]&~m[734]&m[735]&m[737]&m[738])|(~m[733]&m[734]&m[735]&m[737]&m[738]))&UnbiasedRNG[417])|((m[733]&m[734]&~m[735]&~m[737]&~m[738])|(m[733]&~m[734]&m[735]&~m[737]&~m[738])|(~m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&~m[734]&~m[735]&~m[737]&m[738])|(~m[733]&m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&~m[737]&m[738])|(~m[733]&~m[734]&m[735]&~m[737]&m[738])|(m[733]&~m[734]&m[735]&~m[737]&m[738])|(~m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&m[737]&m[738]))):InitCond[944];
    m[741] = run?((((m[738]&~m[739]&~m[740]&~m[742]&~m[743])|(~m[738]&m[739]&~m[740]&~m[742]&~m[743])|(~m[738]&~m[739]&m[740]&~m[742]&~m[743])|(m[738]&m[739]&m[740]&m[742]&~m[743])|(~m[738]&~m[739]&~m[740]&~m[742]&m[743])|(m[738]&m[739]&~m[740]&m[742]&m[743])|(m[738]&~m[739]&m[740]&m[742]&m[743])|(~m[738]&m[739]&m[740]&m[742]&m[743]))&UnbiasedRNG[418])|((m[738]&m[739]&~m[740]&~m[742]&~m[743])|(m[738]&~m[739]&m[740]&~m[742]&~m[743])|(~m[738]&m[739]&m[740]&~m[742]&~m[743])|(m[738]&m[739]&m[740]&~m[742]&~m[743])|(m[738]&~m[739]&~m[740]&~m[742]&m[743])|(~m[738]&m[739]&~m[740]&~m[742]&m[743])|(m[738]&m[739]&~m[740]&~m[742]&m[743])|(~m[738]&~m[739]&m[740]&~m[742]&m[743])|(m[738]&~m[739]&m[740]&~m[742]&m[743])|(~m[738]&m[739]&m[740]&~m[742]&m[743])|(m[738]&m[739]&m[740]&~m[742]&m[743])|(m[738]&m[739]&m[740]&m[742]&m[743]))):InitCond[945];
    m[746] = run?((((m[743]&~m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&~m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&m[747]&~m[748])|(~m[743]&~m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&m[747]&m[748])|(m[743]&~m[744]&m[745]&m[747]&m[748])|(~m[743]&m[744]&m[745]&m[747]&m[748]))&UnbiasedRNG[419])|((m[743]&m[744]&~m[745]&~m[747]&~m[748])|(m[743]&~m[744]&m[745]&~m[747]&~m[748])|(~m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&~m[744]&~m[745]&~m[747]&m[748])|(~m[743]&m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&~m[747]&m[748])|(~m[743]&~m[744]&m[745]&~m[747]&m[748])|(m[743]&~m[744]&m[745]&~m[747]&m[748])|(~m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&m[747]&m[748]))):InitCond[946];
    m[756] = run?((((m[753]&~m[754]&~m[755]&~m[757]&~m[758])|(~m[753]&m[754]&~m[755]&~m[757]&~m[758])|(~m[753]&~m[754]&m[755]&~m[757]&~m[758])|(m[753]&m[754]&m[755]&m[757]&~m[758])|(~m[753]&~m[754]&~m[755]&~m[757]&m[758])|(m[753]&m[754]&~m[755]&m[757]&m[758])|(m[753]&~m[754]&m[755]&m[757]&m[758])|(~m[753]&m[754]&m[755]&m[757]&m[758]))&UnbiasedRNG[420])|((m[753]&m[754]&~m[755]&~m[757]&~m[758])|(m[753]&~m[754]&m[755]&~m[757]&~m[758])|(~m[753]&m[754]&m[755]&~m[757]&~m[758])|(m[753]&m[754]&m[755]&~m[757]&~m[758])|(m[753]&~m[754]&~m[755]&~m[757]&m[758])|(~m[753]&m[754]&~m[755]&~m[757]&m[758])|(m[753]&m[754]&~m[755]&~m[757]&m[758])|(~m[753]&~m[754]&m[755]&~m[757]&m[758])|(m[753]&~m[754]&m[755]&~m[757]&m[758])|(~m[753]&m[754]&m[755]&~m[757]&m[758])|(m[753]&m[754]&m[755]&~m[757]&m[758])|(m[753]&m[754]&m[755]&m[757]&m[758]))):InitCond[947];
    m[761] = run?((((m[758]&~m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&~m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&m[762]&~m[763])|(~m[758]&~m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&m[762]&m[763])|(m[758]&~m[759]&m[760]&m[762]&m[763])|(~m[758]&m[759]&m[760]&m[762]&m[763]))&UnbiasedRNG[421])|((m[758]&m[759]&~m[760]&~m[762]&~m[763])|(m[758]&~m[759]&m[760]&~m[762]&~m[763])|(~m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&~m[759]&~m[760]&~m[762]&m[763])|(~m[758]&m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&~m[762]&m[763])|(~m[758]&~m[759]&m[760]&~m[762]&m[763])|(m[758]&~m[759]&m[760]&~m[762]&m[763])|(~m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&m[762]&m[763]))):InitCond[948];
    m[766] = run?((((m[763]&~m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&~m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&m[767]&~m[768])|(~m[763]&~m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&m[767]&m[768])|(m[763]&~m[764]&m[765]&m[767]&m[768])|(~m[763]&m[764]&m[765]&m[767]&m[768]))&UnbiasedRNG[422])|((m[763]&m[764]&~m[765]&~m[767]&~m[768])|(m[763]&~m[764]&m[765]&~m[767]&~m[768])|(~m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&~m[764]&~m[765]&~m[767]&m[768])|(~m[763]&m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&~m[767]&m[768])|(~m[763]&~m[764]&m[765]&~m[767]&m[768])|(m[763]&~m[764]&m[765]&~m[767]&m[768])|(~m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&m[767]&m[768]))):InitCond[949];
    m[771] = run?((((m[768]&~m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&~m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&m[772]&~m[773])|(~m[768]&~m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&m[772]&m[773])|(m[768]&~m[769]&m[770]&m[772]&m[773])|(~m[768]&m[769]&m[770]&m[772]&m[773]))&UnbiasedRNG[423])|((m[768]&m[769]&~m[770]&~m[772]&~m[773])|(m[768]&~m[769]&m[770]&~m[772]&~m[773])|(~m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&~m[769]&~m[770]&~m[772]&m[773])|(~m[768]&m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&~m[772]&m[773])|(~m[768]&~m[769]&m[770]&~m[772]&m[773])|(m[768]&~m[769]&m[770]&~m[772]&m[773])|(~m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&m[772]&m[773]))):InitCond[950];
    m[776] = run?((((m[773]&~m[774]&~m[775]&~m[777]&~m[778])|(~m[773]&m[774]&~m[775]&~m[777]&~m[778])|(~m[773]&~m[774]&m[775]&~m[777]&~m[778])|(m[773]&m[774]&m[775]&m[777]&~m[778])|(~m[773]&~m[774]&~m[775]&~m[777]&m[778])|(m[773]&m[774]&~m[775]&m[777]&m[778])|(m[773]&~m[774]&m[775]&m[777]&m[778])|(~m[773]&m[774]&m[775]&m[777]&m[778]))&UnbiasedRNG[424])|((m[773]&m[774]&~m[775]&~m[777]&~m[778])|(m[773]&~m[774]&m[775]&~m[777]&~m[778])|(~m[773]&m[774]&m[775]&~m[777]&~m[778])|(m[773]&m[774]&m[775]&~m[777]&~m[778])|(m[773]&~m[774]&~m[775]&~m[777]&m[778])|(~m[773]&m[774]&~m[775]&~m[777]&m[778])|(m[773]&m[774]&~m[775]&~m[777]&m[778])|(~m[773]&~m[774]&m[775]&~m[777]&m[778])|(m[773]&~m[774]&m[775]&~m[777]&m[778])|(~m[773]&m[774]&m[775]&~m[777]&m[778])|(m[773]&m[774]&m[775]&~m[777]&m[778])|(m[773]&m[774]&m[775]&m[777]&m[778]))):InitCond[951];
    m[781] = run?((((m[778]&~m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&~m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&m[782]&~m[783])|(~m[778]&~m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&m[782]&m[783])|(m[778]&~m[779]&m[780]&m[782]&m[783])|(~m[778]&m[779]&m[780]&m[782]&m[783]))&UnbiasedRNG[425])|((m[778]&m[779]&~m[780]&~m[782]&~m[783])|(m[778]&~m[779]&m[780]&~m[782]&~m[783])|(~m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&~m[779]&~m[780]&~m[782]&m[783])|(~m[778]&m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&~m[782]&m[783])|(~m[778]&~m[779]&m[780]&~m[782]&m[783])|(m[778]&~m[779]&m[780]&~m[782]&m[783])|(~m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&m[782]&m[783]))):InitCond[952];
    m[786] = run?((((m[783]&~m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&~m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&m[787]&~m[788])|(~m[783]&~m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&m[787]&m[788])|(m[783]&~m[784]&m[785]&m[787]&m[788])|(~m[783]&m[784]&m[785]&m[787]&m[788]))&UnbiasedRNG[426])|((m[783]&m[784]&~m[785]&~m[787]&~m[788])|(m[783]&~m[784]&m[785]&~m[787]&~m[788])|(~m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&~m[784]&~m[785]&~m[787]&m[788])|(~m[783]&m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&~m[787]&m[788])|(~m[783]&~m[784]&m[785]&~m[787]&m[788])|(m[783]&~m[784]&m[785]&~m[787]&m[788])|(~m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&m[787]&m[788]))):InitCond[953];
    m[791] = run?((((m[788]&~m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&~m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&m[792]&~m[793])|(~m[788]&~m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&m[792]&m[793])|(m[788]&~m[789]&m[790]&m[792]&m[793])|(~m[788]&m[789]&m[790]&m[792]&m[793]))&UnbiasedRNG[427])|((m[788]&m[789]&~m[790]&~m[792]&~m[793])|(m[788]&~m[789]&m[790]&~m[792]&~m[793])|(~m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&~m[789]&~m[790]&~m[792]&m[793])|(~m[788]&m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&~m[792]&m[793])|(~m[788]&~m[789]&m[790]&~m[792]&m[793])|(m[788]&~m[789]&m[790]&~m[792]&m[793])|(~m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&m[792]&m[793]))):InitCond[954];
    m[796] = run?((((m[793]&~m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&~m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&m[797]&~m[798])|(~m[793]&~m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&m[797]&m[798])|(m[793]&~m[794]&m[795]&m[797]&m[798])|(~m[793]&m[794]&m[795]&m[797]&m[798]))&UnbiasedRNG[428])|((m[793]&m[794]&~m[795]&~m[797]&~m[798])|(m[793]&~m[794]&m[795]&~m[797]&~m[798])|(~m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&~m[794]&~m[795]&~m[797]&m[798])|(~m[793]&m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&~m[797]&m[798])|(~m[793]&~m[794]&m[795]&~m[797]&m[798])|(m[793]&~m[794]&m[795]&~m[797]&m[798])|(~m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&m[797]&m[798]))):InitCond[955];
    m[806] = run?((((m[803]&~m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&~m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&m[807]&~m[808])|(~m[803]&~m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&m[807]&m[808])|(m[803]&~m[804]&m[805]&m[807]&m[808])|(~m[803]&m[804]&m[805]&m[807]&m[808]))&UnbiasedRNG[429])|((m[803]&m[804]&~m[805]&~m[807]&~m[808])|(m[803]&~m[804]&m[805]&~m[807]&~m[808])|(~m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&~m[804]&~m[805]&~m[807]&m[808])|(~m[803]&m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&~m[807]&m[808])|(~m[803]&~m[804]&m[805]&~m[807]&m[808])|(m[803]&~m[804]&m[805]&~m[807]&m[808])|(~m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&m[807]&m[808]))):InitCond[956];
    m[811] = run?((((m[808]&~m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&~m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&m[812]&~m[813])|(~m[808]&~m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&m[812]&m[813])|(m[808]&~m[809]&m[810]&m[812]&m[813])|(~m[808]&m[809]&m[810]&m[812]&m[813]))&UnbiasedRNG[430])|((m[808]&m[809]&~m[810]&~m[812]&~m[813])|(m[808]&~m[809]&m[810]&~m[812]&~m[813])|(~m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&~m[809]&~m[810]&~m[812]&m[813])|(~m[808]&m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&~m[812]&m[813])|(~m[808]&~m[809]&m[810]&~m[812]&m[813])|(m[808]&~m[809]&m[810]&~m[812]&m[813])|(~m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&m[812]&m[813]))):InitCond[957];
    m[816] = run?((((m[813]&~m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&~m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&m[817]&~m[818])|(~m[813]&~m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&m[817]&m[818])|(m[813]&~m[814]&m[815]&m[817]&m[818])|(~m[813]&m[814]&m[815]&m[817]&m[818]))&UnbiasedRNG[431])|((m[813]&m[814]&~m[815]&~m[817]&~m[818])|(m[813]&~m[814]&m[815]&~m[817]&~m[818])|(~m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&~m[814]&~m[815]&~m[817]&m[818])|(~m[813]&m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&~m[817]&m[818])|(~m[813]&~m[814]&m[815]&~m[817]&m[818])|(m[813]&~m[814]&m[815]&~m[817]&m[818])|(~m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&m[817]&m[818]))):InitCond[958];
    m[821] = run?((((m[818]&~m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&~m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&m[822]&~m[823])|(~m[818]&~m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&m[822]&m[823])|(m[818]&~m[819]&m[820]&m[822]&m[823])|(~m[818]&m[819]&m[820]&m[822]&m[823]))&UnbiasedRNG[432])|((m[818]&m[819]&~m[820]&~m[822]&~m[823])|(m[818]&~m[819]&m[820]&~m[822]&~m[823])|(~m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&~m[819]&~m[820]&~m[822]&m[823])|(~m[818]&m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&~m[822]&m[823])|(~m[818]&~m[819]&m[820]&~m[822]&m[823])|(m[818]&~m[819]&m[820]&~m[822]&m[823])|(~m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&m[822]&m[823]))):InitCond[959];
    m[826] = run?((((m[823]&~m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&~m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&m[827]&~m[828])|(~m[823]&~m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&m[827]&m[828])|(m[823]&~m[824]&m[825]&m[827]&m[828])|(~m[823]&m[824]&m[825]&m[827]&m[828]))&UnbiasedRNG[433])|((m[823]&m[824]&~m[825]&~m[827]&~m[828])|(m[823]&~m[824]&m[825]&~m[827]&~m[828])|(~m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&~m[824]&~m[825]&~m[827]&m[828])|(~m[823]&m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&~m[827]&m[828])|(~m[823]&~m[824]&m[825]&~m[827]&m[828])|(m[823]&~m[824]&m[825]&~m[827]&m[828])|(~m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&m[827]&m[828]))):InitCond[960];
    m[831] = run?((((m[828]&~m[829]&~m[830]&~m[832]&~m[833])|(~m[828]&m[829]&~m[830]&~m[832]&~m[833])|(~m[828]&~m[829]&m[830]&~m[832]&~m[833])|(m[828]&m[829]&m[830]&m[832]&~m[833])|(~m[828]&~m[829]&~m[830]&~m[832]&m[833])|(m[828]&m[829]&~m[830]&m[832]&m[833])|(m[828]&~m[829]&m[830]&m[832]&m[833])|(~m[828]&m[829]&m[830]&m[832]&m[833]))&UnbiasedRNG[434])|((m[828]&m[829]&~m[830]&~m[832]&~m[833])|(m[828]&~m[829]&m[830]&~m[832]&~m[833])|(~m[828]&m[829]&m[830]&~m[832]&~m[833])|(m[828]&m[829]&m[830]&~m[832]&~m[833])|(m[828]&~m[829]&~m[830]&~m[832]&m[833])|(~m[828]&m[829]&~m[830]&~m[832]&m[833])|(m[828]&m[829]&~m[830]&~m[832]&m[833])|(~m[828]&~m[829]&m[830]&~m[832]&m[833])|(m[828]&~m[829]&m[830]&~m[832]&m[833])|(~m[828]&m[829]&m[830]&~m[832]&m[833])|(m[828]&m[829]&m[830]&~m[832]&m[833])|(m[828]&m[829]&m[830]&m[832]&m[833]))):InitCond[961];
    m[836] = run?((((m[833]&~m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&~m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&m[837]&~m[838])|(~m[833]&~m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&m[837]&m[838])|(m[833]&~m[834]&m[835]&m[837]&m[838])|(~m[833]&m[834]&m[835]&m[837]&m[838]))&UnbiasedRNG[435])|((m[833]&m[834]&~m[835]&~m[837]&~m[838])|(m[833]&~m[834]&m[835]&~m[837]&~m[838])|(~m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&~m[834]&~m[835]&~m[837]&m[838])|(~m[833]&m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&~m[837]&m[838])|(~m[833]&~m[834]&m[835]&~m[837]&m[838])|(m[833]&~m[834]&m[835]&~m[837]&m[838])|(~m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&m[837]&m[838]))):InitCond[962];
    m[841] = run?((((m[838]&~m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&~m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&m[842]&~m[843])|(~m[838]&~m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&m[842]&m[843])|(m[838]&~m[839]&m[840]&m[842]&m[843])|(~m[838]&m[839]&m[840]&m[842]&m[843]))&UnbiasedRNG[436])|((m[838]&m[839]&~m[840]&~m[842]&~m[843])|(m[838]&~m[839]&m[840]&~m[842]&~m[843])|(~m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&~m[839]&~m[840]&~m[842]&m[843])|(~m[838]&m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&~m[842]&m[843])|(~m[838]&~m[839]&m[840]&~m[842]&m[843])|(m[838]&~m[839]&m[840]&~m[842]&m[843])|(~m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&m[842]&m[843]))):InitCond[963];
    m[846] = run?((((m[843]&~m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&~m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&m[847]&~m[848])|(~m[843]&~m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&m[847]&m[848])|(m[843]&~m[844]&m[845]&m[847]&m[848])|(~m[843]&m[844]&m[845]&m[847]&m[848]))&UnbiasedRNG[437])|((m[843]&m[844]&~m[845]&~m[847]&~m[848])|(m[843]&~m[844]&m[845]&~m[847]&~m[848])|(~m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&~m[844]&~m[845]&~m[847]&m[848])|(~m[843]&m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&~m[847]&m[848])|(~m[843]&~m[844]&m[845]&~m[847]&m[848])|(m[843]&~m[844]&m[845]&~m[847]&m[848])|(~m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&m[847]&m[848]))):InitCond[964];
    m[851] = run?((((m[848]&~m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&~m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&m[852]&~m[853])|(~m[848]&~m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&m[852]&m[853])|(m[848]&~m[849]&m[850]&m[852]&m[853])|(~m[848]&m[849]&m[850]&m[852]&m[853]))&UnbiasedRNG[438])|((m[848]&m[849]&~m[850]&~m[852]&~m[853])|(m[848]&~m[849]&m[850]&~m[852]&~m[853])|(~m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&~m[849]&~m[850]&~m[852]&m[853])|(~m[848]&m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&~m[852]&m[853])|(~m[848]&~m[849]&m[850]&~m[852]&m[853])|(m[848]&~m[849]&m[850]&~m[852]&m[853])|(~m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&m[852]&m[853]))):InitCond[965];
    m[861] = run?((((m[858]&~m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&~m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&m[862]&~m[863])|(~m[858]&~m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&m[862]&m[863])|(m[858]&~m[859]&m[860]&m[862]&m[863])|(~m[858]&m[859]&m[860]&m[862]&m[863]))&UnbiasedRNG[439])|((m[858]&m[859]&~m[860]&~m[862]&~m[863])|(m[858]&~m[859]&m[860]&~m[862]&~m[863])|(~m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&~m[859]&~m[860]&~m[862]&m[863])|(~m[858]&m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&~m[862]&m[863])|(~m[858]&~m[859]&m[860]&~m[862]&m[863])|(m[858]&~m[859]&m[860]&~m[862]&m[863])|(~m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&m[862]&m[863]))):InitCond[966];
    m[866] = run?((((m[863]&~m[864]&~m[865]&~m[867]&~m[868])|(~m[863]&m[864]&~m[865]&~m[867]&~m[868])|(~m[863]&~m[864]&m[865]&~m[867]&~m[868])|(m[863]&m[864]&m[865]&m[867]&~m[868])|(~m[863]&~m[864]&~m[865]&~m[867]&m[868])|(m[863]&m[864]&~m[865]&m[867]&m[868])|(m[863]&~m[864]&m[865]&m[867]&m[868])|(~m[863]&m[864]&m[865]&m[867]&m[868]))&UnbiasedRNG[440])|((m[863]&m[864]&~m[865]&~m[867]&~m[868])|(m[863]&~m[864]&m[865]&~m[867]&~m[868])|(~m[863]&m[864]&m[865]&~m[867]&~m[868])|(m[863]&m[864]&m[865]&~m[867]&~m[868])|(m[863]&~m[864]&~m[865]&~m[867]&m[868])|(~m[863]&m[864]&~m[865]&~m[867]&m[868])|(m[863]&m[864]&~m[865]&~m[867]&m[868])|(~m[863]&~m[864]&m[865]&~m[867]&m[868])|(m[863]&~m[864]&m[865]&~m[867]&m[868])|(~m[863]&m[864]&m[865]&~m[867]&m[868])|(m[863]&m[864]&m[865]&~m[867]&m[868])|(m[863]&m[864]&m[865]&m[867]&m[868]))):InitCond[967];
    m[871] = run?((((m[868]&~m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&~m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&m[872]&~m[873])|(~m[868]&~m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&m[872]&m[873])|(m[868]&~m[869]&m[870]&m[872]&m[873])|(~m[868]&m[869]&m[870]&m[872]&m[873]))&UnbiasedRNG[441])|((m[868]&m[869]&~m[870]&~m[872]&~m[873])|(m[868]&~m[869]&m[870]&~m[872]&~m[873])|(~m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&~m[869]&~m[870]&~m[872]&m[873])|(~m[868]&m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&~m[872]&m[873])|(~m[868]&~m[869]&m[870]&~m[872]&m[873])|(m[868]&~m[869]&m[870]&~m[872]&m[873])|(~m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&m[872]&m[873]))):InitCond[968];
    m[876] = run?((((m[873]&~m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&~m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&m[877]&~m[878])|(~m[873]&~m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&m[877]&m[878])|(m[873]&~m[874]&m[875]&m[877]&m[878])|(~m[873]&m[874]&m[875]&m[877]&m[878]))&UnbiasedRNG[442])|((m[873]&m[874]&~m[875]&~m[877]&~m[878])|(m[873]&~m[874]&m[875]&~m[877]&~m[878])|(~m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&~m[874]&~m[875]&~m[877]&m[878])|(~m[873]&m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&~m[877]&m[878])|(~m[873]&~m[874]&m[875]&~m[877]&m[878])|(m[873]&~m[874]&m[875]&~m[877]&m[878])|(~m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&m[877]&m[878]))):InitCond[969];
    m[881] = run?((((m[878]&~m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&~m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&m[882]&~m[883])|(~m[878]&~m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&m[882]&m[883])|(m[878]&~m[879]&m[880]&m[882]&m[883])|(~m[878]&m[879]&m[880]&m[882]&m[883]))&UnbiasedRNG[443])|((m[878]&m[879]&~m[880]&~m[882]&~m[883])|(m[878]&~m[879]&m[880]&~m[882]&~m[883])|(~m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&~m[879]&~m[880]&~m[882]&m[883])|(~m[878]&m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&~m[882]&m[883])|(~m[878]&~m[879]&m[880]&~m[882]&m[883])|(m[878]&~m[879]&m[880]&~m[882]&m[883])|(~m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&m[882]&m[883]))):InitCond[970];
    m[886] = run?((((m[883]&~m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&~m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&m[887]&~m[888])|(~m[883]&~m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&m[887]&m[888])|(m[883]&~m[884]&m[885]&m[887]&m[888])|(~m[883]&m[884]&m[885]&m[887]&m[888]))&UnbiasedRNG[444])|((m[883]&m[884]&~m[885]&~m[887]&~m[888])|(m[883]&~m[884]&m[885]&~m[887]&~m[888])|(~m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&~m[884]&~m[885]&~m[887]&m[888])|(~m[883]&m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&~m[887]&m[888])|(~m[883]&~m[884]&m[885]&~m[887]&m[888])|(m[883]&~m[884]&m[885]&~m[887]&m[888])|(~m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&m[887]&m[888]))):InitCond[971];
    m[891] = run?((((m[888]&~m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&~m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&m[892]&~m[893])|(~m[888]&~m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&m[892]&m[893])|(m[888]&~m[889]&m[890]&m[892]&m[893])|(~m[888]&m[889]&m[890]&m[892]&m[893]))&UnbiasedRNG[445])|((m[888]&m[889]&~m[890]&~m[892]&~m[893])|(m[888]&~m[889]&m[890]&~m[892]&~m[893])|(~m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&~m[889]&~m[890]&~m[892]&m[893])|(~m[888]&m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&~m[892]&m[893])|(~m[888]&~m[889]&m[890]&~m[892]&m[893])|(m[888]&~m[889]&m[890]&~m[892]&m[893])|(~m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&m[892]&m[893]))):InitCond[972];
    m[896] = run?((((m[893]&~m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&~m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&m[897]&~m[898])|(~m[893]&~m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&m[897]&m[898])|(m[893]&~m[894]&m[895]&m[897]&m[898])|(~m[893]&m[894]&m[895]&m[897]&m[898]))&UnbiasedRNG[446])|((m[893]&m[894]&~m[895]&~m[897]&~m[898])|(m[893]&~m[894]&m[895]&~m[897]&~m[898])|(~m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&~m[894]&~m[895]&~m[897]&m[898])|(~m[893]&m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&~m[897]&m[898])|(~m[893]&~m[894]&m[895]&~m[897]&m[898])|(m[893]&~m[894]&m[895]&~m[897]&m[898])|(~m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&m[897]&m[898]))):InitCond[973];
    m[901] = run?((((m[898]&~m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&~m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&m[902]&~m[903])|(~m[898]&~m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&m[902]&m[903])|(m[898]&~m[899]&m[900]&m[902]&m[903])|(~m[898]&m[899]&m[900]&m[902]&m[903]))&UnbiasedRNG[447])|((m[898]&m[899]&~m[900]&~m[902]&~m[903])|(m[898]&~m[899]&m[900]&~m[902]&~m[903])|(~m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&~m[899]&~m[900]&~m[902]&m[903])|(~m[898]&m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&~m[902]&m[903])|(~m[898]&~m[899]&m[900]&~m[902]&m[903])|(m[898]&~m[899]&m[900]&~m[902]&m[903])|(~m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&m[902]&m[903]))):InitCond[974];
    m[906] = run?((((m[903]&~m[904]&~m[905]&~m[907]&~m[908])|(~m[903]&m[904]&~m[905]&~m[907]&~m[908])|(~m[903]&~m[904]&m[905]&~m[907]&~m[908])|(m[903]&m[904]&m[905]&m[907]&~m[908])|(~m[903]&~m[904]&~m[905]&~m[907]&m[908])|(m[903]&m[904]&~m[905]&m[907]&m[908])|(m[903]&~m[904]&m[905]&m[907]&m[908])|(~m[903]&m[904]&m[905]&m[907]&m[908]))&UnbiasedRNG[448])|((m[903]&m[904]&~m[905]&~m[907]&~m[908])|(m[903]&~m[904]&m[905]&~m[907]&~m[908])|(~m[903]&m[904]&m[905]&~m[907]&~m[908])|(m[903]&m[904]&m[905]&~m[907]&~m[908])|(m[903]&~m[904]&~m[905]&~m[907]&m[908])|(~m[903]&m[904]&~m[905]&~m[907]&m[908])|(m[903]&m[904]&~m[905]&~m[907]&m[908])|(~m[903]&~m[904]&m[905]&~m[907]&m[908])|(m[903]&~m[904]&m[905]&~m[907]&m[908])|(~m[903]&m[904]&m[905]&~m[907]&m[908])|(m[903]&m[904]&m[905]&~m[907]&m[908])|(m[903]&m[904]&m[905]&m[907]&m[908]))):InitCond[975];
    m[916] = run?((((m[913]&~m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&~m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&m[917]&~m[918])|(~m[913]&~m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&m[917]&m[918])|(m[913]&~m[914]&m[915]&m[917]&m[918])|(~m[913]&m[914]&m[915]&m[917]&m[918]))&UnbiasedRNG[449])|((m[913]&m[914]&~m[915]&~m[917]&~m[918])|(m[913]&~m[914]&m[915]&~m[917]&~m[918])|(~m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&~m[914]&~m[915]&~m[917]&m[918])|(~m[913]&m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&~m[917]&m[918])|(~m[913]&~m[914]&m[915]&~m[917]&m[918])|(m[913]&~m[914]&m[915]&~m[917]&m[918])|(~m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&m[917]&m[918]))):InitCond[976];
    m[921] = run?((((m[918]&~m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&~m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&m[922]&~m[923])|(~m[918]&~m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&m[922]&m[923])|(m[918]&~m[919]&m[920]&m[922]&m[923])|(~m[918]&m[919]&m[920]&m[922]&m[923]))&UnbiasedRNG[450])|((m[918]&m[919]&~m[920]&~m[922]&~m[923])|(m[918]&~m[919]&m[920]&~m[922]&~m[923])|(~m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&~m[919]&~m[920]&~m[922]&m[923])|(~m[918]&m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&~m[922]&m[923])|(~m[918]&~m[919]&m[920]&~m[922]&m[923])|(m[918]&~m[919]&m[920]&~m[922]&m[923])|(~m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&m[922]&m[923]))):InitCond[977];
    m[926] = run?((((m[923]&~m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&~m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&m[927]&~m[928])|(~m[923]&~m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&m[927]&m[928])|(m[923]&~m[924]&m[925]&m[927]&m[928])|(~m[923]&m[924]&m[925]&m[927]&m[928]))&UnbiasedRNG[451])|((m[923]&m[924]&~m[925]&~m[927]&~m[928])|(m[923]&~m[924]&m[925]&~m[927]&~m[928])|(~m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&~m[924]&~m[925]&~m[927]&m[928])|(~m[923]&m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&~m[927]&m[928])|(~m[923]&~m[924]&m[925]&~m[927]&m[928])|(m[923]&~m[924]&m[925]&~m[927]&m[928])|(~m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&m[927]&m[928]))):InitCond[978];
    m[931] = run?((((m[928]&~m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&~m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&m[932]&~m[933])|(~m[928]&~m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&m[932]&m[933])|(m[928]&~m[929]&m[930]&m[932]&m[933])|(~m[928]&m[929]&m[930]&m[932]&m[933]))&UnbiasedRNG[452])|((m[928]&m[929]&~m[930]&~m[932]&~m[933])|(m[928]&~m[929]&m[930]&~m[932]&~m[933])|(~m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&~m[929]&~m[930]&~m[932]&m[933])|(~m[928]&m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&~m[932]&m[933])|(~m[928]&~m[929]&m[930]&~m[932]&m[933])|(m[928]&~m[929]&m[930]&~m[932]&m[933])|(~m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&m[932]&m[933]))):InitCond[979];
    m[936] = run?((((m[933]&~m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&~m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&m[937]&~m[938])|(~m[933]&~m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&m[937]&m[938])|(m[933]&~m[934]&m[935]&m[937]&m[938])|(~m[933]&m[934]&m[935]&m[937]&m[938]))&UnbiasedRNG[453])|((m[933]&m[934]&~m[935]&~m[937]&~m[938])|(m[933]&~m[934]&m[935]&~m[937]&~m[938])|(~m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&~m[934]&~m[935]&~m[937]&m[938])|(~m[933]&m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&~m[937]&m[938])|(~m[933]&~m[934]&m[935]&~m[937]&m[938])|(m[933]&~m[934]&m[935]&~m[937]&m[938])|(~m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&m[937]&m[938]))):InitCond[980];
    m[941] = run?((((m[938]&~m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&~m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&m[942]&~m[943])|(~m[938]&~m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&m[942]&m[943])|(m[938]&~m[939]&m[940]&m[942]&m[943])|(~m[938]&m[939]&m[940]&m[942]&m[943]))&UnbiasedRNG[454])|((m[938]&m[939]&~m[940]&~m[942]&~m[943])|(m[938]&~m[939]&m[940]&~m[942]&~m[943])|(~m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&~m[939]&~m[940]&~m[942]&m[943])|(~m[938]&m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&~m[942]&m[943])|(~m[938]&~m[939]&m[940]&~m[942]&m[943])|(m[938]&~m[939]&m[940]&~m[942]&m[943])|(~m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&m[942]&m[943]))):InitCond[981];
    m[946] = run?((((m[943]&~m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&~m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&m[947]&~m[948])|(~m[943]&~m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&m[947]&m[948])|(m[943]&~m[944]&m[945]&m[947]&m[948])|(~m[943]&m[944]&m[945]&m[947]&m[948]))&UnbiasedRNG[455])|((m[943]&m[944]&~m[945]&~m[947]&~m[948])|(m[943]&~m[944]&m[945]&~m[947]&~m[948])|(~m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&~m[944]&~m[945]&~m[947]&m[948])|(~m[943]&m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&~m[947]&m[948])|(~m[943]&~m[944]&m[945]&~m[947]&m[948])|(m[943]&~m[944]&m[945]&~m[947]&m[948])|(~m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&m[947]&m[948]))):InitCond[982];
    m[951] = run?((((m[948]&~m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&~m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&m[952]&~m[953])|(~m[948]&~m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&m[952]&m[953])|(m[948]&~m[949]&m[950]&m[952]&m[953])|(~m[948]&m[949]&m[950]&m[952]&m[953]))&UnbiasedRNG[456])|((m[948]&m[949]&~m[950]&~m[952]&~m[953])|(m[948]&~m[949]&m[950]&~m[952]&~m[953])|(~m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&~m[949]&~m[950]&~m[952]&m[953])|(~m[948]&m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&~m[952]&m[953])|(~m[948]&~m[949]&m[950]&~m[952]&m[953])|(m[948]&~m[949]&m[950]&~m[952]&m[953])|(~m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&m[952]&m[953]))):InitCond[983];
    m[956] = run?((((m[953]&~m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&~m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&m[957]&~m[958])|(~m[953]&~m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&m[957]&m[958])|(m[953]&~m[954]&m[955]&m[957]&m[958])|(~m[953]&m[954]&m[955]&m[957]&m[958]))&UnbiasedRNG[457])|((m[953]&m[954]&~m[955]&~m[957]&~m[958])|(m[953]&~m[954]&m[955]&~m[957]&~m[958])|(~m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&~m[954]&~m[955]&~m[957]&m[958])|(~m[953]&m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&~m[957]&m[958])|(~m[953]&~m[954]&m[955]&~m[957]&m[958])|(m[953]&~m[954]&m[955]&~m[957]&m[958])|(~m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&m[957]&m[958]))):InitCond[984];
    m[966] = run?((((m[963]&~m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&~m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&m[967]&~m[968])|(~m[963]&~m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&m[967]&m[968])|(m[963]&~m[964]&m[965]&m[967]&m[968])|(~m[963]&m[964]&m[965]&m[967]&m[968]))&UnbiasedRNG[458])|((m[963]&m[964]&~m[965]&~m[967]&~m[968])|(m[963]&~m[964]&m[965]&~m[967]&~m[968])|(~m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&~m[964]&~m[965]&~m[967]&m[968])|(~m[963]&m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&~m[967]&m[968])|(~m[963]&~m[964]&m[965]&~m[967]&m[968])|(m[963]&~m[964]&m[965]&~m[967]&m[968])|(~m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&m[967]&m[968]))):InitCond[985];
    m[971] = run?((((m[968]&~m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&~m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&m[972]&~m[973])|(~m[968]&~m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&m[972]&m[973])|(m[968]&~m[969]&m[970]&m[972]&m[973])|(~m[968]&m[969]&m[970]&m[972]&m[973]))&UnbiasedRNG[459])|((m[968]&m[969]&~m[970]&~m[972]&~m[973])|(m[968]&~m[969]&m[970]&~m[972]&~m[973])|(~m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&~m[969]&~m[970]&~m[972]&m[973])|(~m[968]&m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&~m[972]&m[973])|(~m[968]&~m[969]&m[970]&~m[972]&m[973])|(m[968]&~m[969]&m[970]&~m[972]&m[973])|(~m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&m[972]&m[973]))):InitCond[986];
    m[976] = run?((((m[973]&~m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&~m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&m[977]&~m[978])|(~m[973]&~m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&m[977]&m[978])|(m[973]&~m[974]&m[975]&m[977]&m[978])|(~m[973]&m[974]&m[975]&m[977]&m[978]))&UnbiasedRNG[460])|((m[973]&m[974]&~m[975]&~m[977]&~m[978])|(m[973]&~m[974]&m[975]&~m[977]&~m[978])|(~m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&~m[974]&~m[975]&~m[977]&m[978])|(~m[973]&m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&~m[977]&m[978])|(~m[973]&~m[974]&m[975]&~m[977]&m[978])|(m[973]&~m[974]&m[975]&~m[977]&m[978])|(~m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&m[977]&m[978]))):InitCond[987];
    m[981] = run?((((m[978]&~m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&~m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&m[982]&~m[983])|(~m[978]&~m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&m[982]&m[983])|(m[978]&~m[979]&m[980]&m[982]&m[983])|(~m[978]&m[979]&m[980]&m[982]&m[983]))&UnbiasedRNG[461])|((m[978]&m[979]&~m[980]&~m[982]&~m[983])|(m[978]&~m[979]&m[980]&~m[982]&~m[983])|(~m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&~m[979]&~m[980]&~m[982]&m[983])|(~m[978]&m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&~m[982]&m[983])|(~m[978]&~m[979]&m[980]&~m[982]&m[983])|(m[978]&~m[979]&m[980]&~m[982]&m[983])|(~m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&m[982]&m[983]))):InitCond[988];
    m[986] = run?((((m[983]&~m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&~m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&m[987]&~m[988])|(~m[983]&~m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&m[987]&m[988])|(m[983]&~m[984]&m[985]&m[987]&m[988])|(~m[983]&m[984]&m[985]&m[987]&m[988]))&UnbiasedRNG[462])|((m[983]&m[984]&~m[985]&~m[987]&~m[988])|(m[983]&~m[984]&m[985]&~m[987]&~m[988])|(~m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&~m[984]&~m[985]&~m[987]&m[988])|(~m[983]&m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&~m[987]&m[988])|(~m[983]&~m[984]&m[985]&~m[987]&m[988])|(m[983]&~m[984]&m[985]&~m[987]&m[988])|(~m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&m[987]&m[988]))):InitCond[989];
    m[991] = run?((((m[988]&~m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&~m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&m[992]&~m[993])|(~m[988]&~m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&m[992]&m[993])|(m[988]&~m[989]&m[990]&m[992]&m[993])|(~m[988]&m[989]&m[990]&m[992]&m[993]))&UnbiasedRNG[463])|((m[988]&m[989]&~m[990]&~m[992]&~m[993])|(m[988]&~m[989]&m[990]&~m[992]&~m[993])|(~m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&~m[989]&~m[990]&~m[992]&m[993])|(~m[988]&m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&~m[992]&m[993])|(~m[988]&~m[989]&m[990]&~m[992]&m[993])|(m[988]&~m[989]&m[990]&~m[992]&m[993])|(~m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&m[992]&m[993]))):InitCond[990];
    m[996] = run?((((m[993]&~m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&~m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&m[997]&~m[998])|(~m[993]&~m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&m[997]&m[998])|(m[993]&~m[994]&m[995]&m[997]&m[998])|(~m[993]&m[994]&m[995]&m[997]&m[998]))&UnbiasedRNG[464])|((m[993]&m[994]&~m[995]&~m[997]&~m[998])|(m[993]&~m[994]&m[995]&~m[997]&~m[998])|(~m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&~m[994]&~m[995]&~m[997]&m[998])|(~m[993]&m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&~m[997]&m[998])|(~m[993]&~m[994]&m[995]&~m[997]&m[998])|(m[993]&~m[994]&m[995]&~m[997]&m[998])|(~m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&m[997]&m[998]))):InitCond[991];
    m[1001] = run?((((m[998]&~m[999]&~m[1000]&~m[1002]&~m[1003])|(~m[998]&m[999]&~m[1000]&~m[1002]&~m[1003])|(~m[998]&~m[999]&m[1000]&~m[1002]&~m[1003])|(m[998]&m[999]&m[1000]&m[1002]&~m[1003])|(~m[998]&~m[999]&~m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&~m[1000]&m[1002]&m[1003])|(m[998]&~m[999]&m[1000]&m[1002]&m[1003])|(~m[998]&m[999]&m[1000]&m[1002]&m[1003]))&UnbiasedRNG[465])|((m[998]&m[999]&~m[1000]&~m[1002]&~m[1003])|(m[998]&~m[999]&m[1000]&~m[1002]&~m[1003])|(~m[998]&m[999]&m[1000]&~m[1002]&~m[1003])|(m[998]&m[999]&m[1000]&~m[1002]&~m[1003])|(m[998]&~m[999]&~m[1000]&~m[1002]&m[1003])|(~m[998]&m[999]&~m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&~m[1000]&~m[1002]&m[1003])|(~m[998]&~m[999]&m[1000]&~m[1002]&m[1003])|(m[998]&~m[999]&m[1000]&~m[1002]&m[1003])|(~m[998]&m[999]&m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&m[1000]&m[1002]&m[1003]))):InitCond[992];
    m[1011] = run?((((m[1008]&~m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&~m[1013])|(~m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))&UnbiasedRNG[466])|((m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))):InitCond[993];
    m[1016] = run?((((m[1013]&~m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&~m[1018])|(~m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))&UnbiasedRNG[467])|((m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))):InitCond[994];
    m[1021] = run?((((m[1018]&~m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&~m[1023])|(~m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))&UnbiasedRNG[468])|((m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))):InitCond[995];
    m[1026] = run?((((m[1023]&~m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&~m[1028])|(~m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))&UnbiasedRNG[469])|((m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))):InitCond[996];
    m[1031] = run?((((m[1028]&~m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&~m[1033])|(~m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&m[1032]&m[1033]))&UnbiasedRNG[470])|((m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&m[1033]))):InitCond[997];
    m[1036] = run?((((m[1033]&~m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&~m[1038])|(~m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))&UnbiasedRNG[471])|((m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))):InitCond[998];
    m[1041] = run?((((m[1038]&~m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&~m[1043])|(~m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))&UnbiasedRNG[472])|((m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))):InitCond[999];
    m[1051] = run?((((m[1048]&~m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&~m[1053])|(~m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))&UnbiasedRNG[473])|((m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))):InitCond[1000];
    m[1056] = run?((((m[1053]&~m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&~m[1058])|(~m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&m[1057]&m[1058]))&UnbiasedRNG[474])|((m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&m[1058]))):InitCond[1001];
    m[1061] = run?((((m[1058]&~m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&~m[1063])|(~m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))&UnbiasedRNG[475])|((m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))):InitCond[1002];
    m[1066] = run?((((m[1063]&~m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&~m[1068])|(~m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&m[1067]&m[1068]))&UnbiasedRNG[476])|((m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&m[1068]))):InitCond[1003];
    m[1071] = run?((((m[1068]&~m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&~m[1073])|(~m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))&UnbiasedRNG[477])|((m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))):InitCond[1004];
    m[1076] = run?((((m[1073]&~m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&~m[1078])|(~m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))&UnbiasedRNG[478])|((m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))):InitCond[1005];
    m[1086] = run?((((m[1083]&~m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&~m[1088])|(~m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))&UnbiasedRNG[479])|((m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))):InitCond[1006];
    m[1091] = run?((((m[1088]&~m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&~m[1093])|(~m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))&UnbiasedRNG[480])|((m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))):InitCond[1007];
    m[1096] = run?((((m[1093]&~m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&~m[1098])|(~m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))&UnbiasedRNG[481])|((m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))):InitCond[1008];
    m[1101] = run?((((m[1098]&~m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&~m[1103])|(~m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))&UnbiasedRNG[482])|((m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))):InitCond[1009];
    m[1106] = run?((((m[1103]&~m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&~m[1108])|(~m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&m[1107]&m[1108]))&UnbiasedRNG[483])|((m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&m[1108]))):InitCond[1010];
    m[1116] = run?((((m[1113]&~m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&~m[1118])|(~m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&m[1117]&m[1118]))&UnbiasedRNG[484])|((m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&m[1118]))):InitCond[1011];
    m[1121] = run?((((m[1118]&~m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&~m[1123])|(~m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))&UnbiasedRNG[485])|((m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))):InitCond[1012];
    m[1126] = run?((((m[1123]&~m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&~m[1128])|(~m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))&UnbiasedRNG[486])|((m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))):InitCond[1013];
    m[1131] = run?((((m[1128]&~m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&~m[1133])|(~m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))&UnbiasedRNG[487])|((m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))):InitCond[1014];
    m[1141] = run?((((m[1138]&~m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&~m[1143])|(~m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))&UnbiasedRNG[488])|((m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))):InitCond[1015];
    m[1146] = run?((((m[1143]&~m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&~m[1148])|(~m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))&UnbiasedRNG[489])|((m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))):InitCond[1016];
    m[1151] = run?((((m[1148]&~m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&~m[1153])|(~m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&m[1152]&m[1153]))&UnbiasedRNG[490])|((m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&m[1153]))):InitCond[1017];
    m[1161] = run?((((m[1158]&~m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&~m[1163])|(~m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))&UnbiasedRNG[491])|((m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))):InitCond[1018];
    m[1166] = run?((((m[1163]&~m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&~m[1168])|(~m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))&UnbiasedRNG[492])|((m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))):InitCond[1019];
    m[1176] = run?((((m[1173]&~m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&~m[1178])|(~m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))&UnbiasedRNG[493])|((m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))):InitCond[1020];
end

always @(posedge color4_clk) begin
    m[532] = run?((((m[528]&~m[529]&~m[530]&~m[531]&~m[535])|(~m[528]&m[529]&~m[530]&~m[531]&~m[535])|(~m[528]&~m[529]&m[530]&~m[531]&~m[535])|(m[528]&m[529]&~m[530]&m[531]&~m[535])|(m[528]&~m[529]&m[530]&m[531]&~m[535])|(~m[528]&m[529]&m[530]&m[531]&~m[535]))&BiasedRNG[527])|(((m[528]&~m[529]&~m[530]&~m[531]&m[535])|(~m[528]&m[529]&~m[530]&~m[531]&m[535])|(~m[528]&~m[529]&m[530]&~m[531]&m[535])|(m[528]&m[529]&~m[530]&m[531]&m[535])|(m[528]&~m[529]&m[530]&m[531]&m[535])|(~m[528]&m[529]&m[530]&m[531]&m[535]))&~BiasedRNG[527])|((m[528]&m[529]&~m[530]&~m[531]&~m[535])|(m[528]&~m[529]&m[530]&~m[531]&~m[535])|(~m[528]&m[529]&m[530]&~m[531]&~m[535])|(m[528]&m[529]&m[530]&~m[531]&~m[535])|(m[528]&m[529]&m[530]&m[531]&~m[535])|(m[528]&m[529]&~m[530]&~m[531]&m[535])|(m[528]&~m[529]&m[530]&~m[531]&m[535])|(~m[528]&m[529]&m[530]&~m[531]&m[535])|(m[528]&m[529]&m[530]&~m[531]&m[535])|(m[528]&m[529]&m[530]&m[531]&m[535]))):InitCond[1021];
    m[537] = run?((((m[533]&~m[534]&~m[535]&~m[536]&~m[545])|(~m[533]&m[534]&~m[535]&~m[536]&~m[545])|(~m[533]&~m[534]&m[535]&~m[536]&~m[545])|(m[533]&m[534]&~m[535]&m[536]&~m[545])|(m[533]&~m[534]&m[535]&m[536]&~m[545])|(~m[533]&m[534]&m[535]&m[536]&~m[545]))&BiasedRNG[528])|(((m[533]&~m[534]&~m[535]&~m[536]&m[545])|(~m[533]&m[534]&~m[535]&~m[536]&m[545])|(~m[533]&~m[534]&m[535]&~m[536]&m[545])|(m[533]&m[534]&~m[535]&m[536]&m[545])|(m[533]&~m[534]&m[535]&m[536]&m[545])|(~m[533]&m[534]&m[535]&m[536]&m[545]))&~BiasedRNG[528])|((m[533]&m[534]&~m[535]&~m[536]&~m[545])|(m[533]&~m[534]&m[535]&~m[536]&~m[545])|(~m[533]&m[534]&m[535]&~m[536]&~m[545])|(m[533]&m[534]&m[535]&~m[536]&~m[545])|(m[533]&m[534]&m[535]&m[536]&~m[545])|(m[533]&m[534]&~m[535]&~m[536]&m[545])|(m[533]&~m[534]&m[535]&~m[536]&m[545])|(~m[533]&m[534]&m[535]&~m[536]&m[545])|(m[533]&m[534]&m[535]&~m[536]&m[545])|(m[533]&m[534]&m[535]&m[536]&m[545]))):InitCond[1022];
    m[542] = run?((((m[538]&~m[539]&~m[540]&~m[541]&~m[550])|(~m[538]&m[539]&~m[540]&~m[541]&~m[550])|(~m[538]&~m[539]&m[540]&~m[541]&~m[550])|(m[538]&m[539]&~m[540]&m[541]&~m[550])|(m[538]&~m[539]&m[540]&m[541]&~m[550])|(~m[538]&m[539]&m[540]&m[541]&~m[550]))&BiasedRNG[529])|(((m[538]&~m[539]&~m[540]&~m[541]&m[550])|(~m[538]&m[539]&~m[540]&~m[541]&m[550])|(~m[538]&~m[539]&m[540]&~m[541]&m[550])|(m[538]&m[539]&~m[540]&m[541]&m[550])|(m[538]&~m[539]&m[540]&m[541]&m[550])|(~m[538]&m[539]&m[540]&m[541]&m[550]))&~BiasedRNG[529])|((m[538]&m[539]&~m[540]&~m[541]&~m[550])|(m[538]&~m[539]&m[540]&~m[541]&~m[550])|(~m[538]&m[539]&m[540]&~m[541]&~m[550])|(m[538]&m[539]&m[540]&~m[541]&~m[550])|(m[538]&m[539]&m[540]&m[541]&~m[550])|(m[538]&m[539]&~m[540]&~m[541]&m[550])|(m[538]&~m[539]&m[540]&~m[541]&m[550])|(~m[538]&m[539]&m[540]&~m[541]&m[550])|(m[538]&m[539]&m[540]&~m[541]&m[550])|(m[538]&m[539]&m[540]&m[541]&m[550]))):InitCond[1023];
    m[547] = run?((((m[543]&~m[544]&~m[545]&~m[546]&~m[560])|(~m[543]&m[544]&~m[545]&~m[546]&~m[560])|(~m[543]&~m[544]&m[545]&~m[546]&~m[560])|(m[543]&m[544]&~m[545]&m[546]&~m[560])|(m[543]&~m[544]&m[545]&m[546]&~m[560])|(~m[543]&m[544]&m[545]&m[546]&~m[560]))&BiasedRNG[530])|(((m[543]&~m[544]&~m[545]&~m[546]&m[560])|(~m[543]&m[544]&~m[545]&~m[546]&m[560])|(~m[543]&~m[544]&m[545]&~m[546]&m[560])|(m[543]&m[544]&~m[545]&m[546]&m[560])|(m[543]&~m[544]&m[545]&m[546]&m[560])|(~m[543]&m[544]&m[545]&m[546]&m[560]))&~BiasedRNG[530])|((m[543]&m[544]&~m[545]&~m[546]&~m[560])|(m[543]&~m[544]&m[545]&~m[546]&~m[560])|(~m[543]&m[544]&m[545]&~m[546]&~m[560])|(m[543]&m[544]&m[545]&~m[546]&~m[560])|(m[543]&m[544]&m[545]&m[546]&~m[560])|(m[543]&m[544]&~m[545]&~m[546]&m[560])|(m[543]&~m[544]&m[545]&~m[546]&m[560])|(~m[543]&m[544]&m[545]&~m[546]&m[560])|(m[543]&m[544]&m[545]&~m[546]&m[560])|(m[543]&m[544]&m[545]&m[546]&m[560]))):InitCond[1024];
    m[552] = run?((((m[548]&~m[549]&~m[550]&~m[551]&~m[565])|(~m[548]&m[549]&~m[550]&~m[551]&~m[565])|(~m[548]&~m[549]&m[550]&~m[551]&~m[565])|(m[548]&m[549]&~m[550]&m[551]&~m[565])|(m[548]&~m[549]&m[550]&m[551]&~m[565])|(~m[548]&m[549]&m[550]&m[551]&~m[565]))&BiasedRNG[531])|(((m[548]&~m[549]&~m[550]&~m[551]&m[565])|(~m[548]&m[549]&~m[550]&~m[551]&m[565])|(~m[548]&~m[549]&m[550]&~m[551]&m[565])|(m[548]&m[549]&~m[550]&m[551]&m[565])|(m[548]&~m[549]&m[550]&m[551]&m[565])|(~m[548]&m[549]&m[550]&m[551]&m[565]))&~BiasedRNG[531])|((m[548]&m[549]&~m[550]&~m[551]&~m[565])|(m[548]&~m[549]&m[550]&~m[551]&~m[565])|(~m[548]&m[549]&m[550]&~m[551]&~m[565])|(m[548]&m[549]&m[550]&~m[551]&~m[565])|(m[548]&m[549]&m[550]&m[551]&~m[565])|(m[548]&m[549]&~m[550]&~m[551]&m[565])|(m[548]&~m[549]&m[550]&~m[551]&m[565])|(~m[548]&m[549]&m[550]&~m[551]&m[565])|(m[548]&m[549]&m[550]&~m[551]&m[565])|(m[548]&m[549]&m[550]&m[551]&m[565]))):InitCond[1025];
    m[557] = run?((((m[553]&~m[554]&~m[555]&~m[556]&~m[570])|(~m[553]&m[554]&~m[555]&~m[556]&~m[570])|(~m[553]&~m[554]&m[555]&~m[556]&~m[570])|(m[553]&m[554]&~m[555]&m[556]&~m[570])|(m[553]&~m[554]&m[555]&m[556]&~m[570])|(~m[553]&m[554]&m[555]&m[556]&~m[570]))&BiasedRNG[532])|(((m[553]&~m[554]&~m[555]&~m[556]&m[570])|(~m[553]&m[554]&~m[555]&~m[556]&m[570])|(~m[553]&~m[554]&m[555]&~m[556]&m[570])|(m[553]&m[554]&~m[555]&m[556]&m[570])|(m[553]&~m[554]&m[555]&m[556]&m[570])|(~m[553]&m[554]&m[555]&m[556]&m[570]))&~BiasedRNG[532])|((m[553]&m[554]&~m[555]&~m[556]&~m[570])|(m[553]&~m[554]&m[555]&~m[556]&~m[570])|(~m[553]&m[554]&m[555]&~m[556]&~m[570])|(m[553]&m[554]&m[555]&~m[556]&~m[570])|(m[553]&m[554]&m[555]&m[556]&~m[570])|(m[553]&m[554]&~m[555]&~m[556]&m[570])|(m[553]&~m[554]&m[555]&~m[556]&m[570])|(~m[553]&m[554]&m[555]&~m[556]&m[570])|(m[553]&m[554]&m[555]&~m[556]&m[570])|(m[553]&m[554]&m[555]&m[556]&m[570]))):InitCond[1026];
    m[562] = run?((((m[558]&~m[559]&~m[560]&~m[561]&~m[580])|(~m[558]&m[559]&~m[560]&~m[561]&~m[580])|(~m[558]&~m[559]&m[560]&~m[561]&~m[580])|(m[558]&m[559]&~m[560]&m[561]&~m[580])|(m[558]&~m[559]&m[560]&m[561]&~m[580])|(~m[558]&m[559]&m[560]&m[561]&~m[580]))&BiasedRNG[533])|(((m[558]&~m[559]&~m[560]&~m[561]&m[580])|(~m[558]&m[559]&~m[560]&~m[561]&m[580])|(~m[558]&~m[559]&m[560]&~m[561]&m[580])|(m[558]&m[559]&~m[560]&m[561]&m[580])|(m[558]&~m[559]&m[560]&m[561]&m[580])|(~m[558]&m[559]&m[560]&m[561]&m[580]))&~BiasedRNG[533])|((m[558]&m[559]&~m[560]&~m[561]&~m[580])|(m[558]&~m[559]&m[560]&~m[561]&~m[580])|(~m[558]&m[559]&m[560]&~m[561]&~m[580])|(m[558]&m[559]&m[560]&~m[561]&~m[580])|(m[558]&m[559]&m[560]&m[561]&~m[580])|(m[558]&m[559]&~m[560]&~m[561]&m[580])|(m[558]&~m[559]&m[560]&~m[561]&m[580])|(~m[558]&m[559]&m[560]&~m[561]&m[580])|(m[558]&m[559]&m[560]&~m[561]&m[580])|(m[558]&m[559]&m[560]&m[561]&m[580]))):InitCond[1027];
    m[567] = run?((((m[563]&~m[564]&~m[565]&~m[566]&~m[585])|(~m[563]&m[564]&~m[565]&~m[566]&~m[585])|(~m[563]&~m[564]&m[565]&~m[566]&~m[585])|(m[563]&m[564]&~m[565]&m[566]&~m[585])|(m[563]&~m[564]&m[565]&m[566]&~m[585])|(~m[563]&m[564]&m[565]&m[566]&~m[585]))&BiasedRNG[534])|(((m[563]&~m[564]&~m[565]&~m[566]&m[585])|(~m[563]&m[564]&~m[565]&~m[566]&m[585])|(~m[563]&~m[564]&m[565]&~m[566]&m[585])|(m[563]&m[564]&~m[565]&m[566]&m[585])|(m[563]&~m[564]&m[565]&m[566]&m[585])|(~m[563]&m[564]&m[565]&m[566]&m[585]))&~BiasedRNG[534])|((m[563]&m[564]&~m[565]&~m[566]&~m[585])|(m[563]&~m[564]&m[565]&~m[566]&~m[585])|(~m[563]&m[564]&m[565]&~m[566]&~m[585])|(m[563]&m[564]&m[565]&~m[566]&~m[585])|(m[563]&m[564]&m[565]&m[566]&~m[585])|(m[563]&m[564]&~m[565]&~m[566]&m[585])|(m[563]&~m[564]&m[565]&~m[566]&m[585])|(~m[563]&m[564]&m[565]&~m[566]&m[585])|(m[563]&m[564]&m[565]&~m[566]&m[585])|(m[563]&m[564]&m[565]&m[566]&m[585]))):InitCond[1028];
    m[572] = run?((((m[568]&~m[569]&~m[570]&~m[571]&~m[590])|(~m[568]&m[569]&~m[570]&~m[571]&~m[590])|(~m[568]&~m[569]&m[570]&~m[571]&~m[590])|(m[568]&m[569]&~m[570]&m[571]&~m[590])|(m[568]&~m[569]&m[570]&m[571]&~m[590])|(~m[568]&m[569]&m[570]&m[571]&~m[590]))&BiasedRNG[535])|(((m[568]&~m[569]&~m[570]&~m[571]&m[590])|(~m[568]&m[569]&~m[570]&~m[571]&m[590])|(~m[568]&~m[569]&m[570]&~m[571]&m[590])|(m[568]&m[569]&~m[570]&m[571]&m[590])|(m[568]&~m[569]&m[570]&m[571]&m[590])|(~m[568]&m[569]&m[570]&m[571]&m[590]))&~BiasedRNG[535])|((m[568]&m[569]&~m[570]&~m[571]&~m[590])|(m[568]&~m[569]&m[570]&~m[571]&~m[590])|(~m[568]&m[569]&m[570]&~m[571]&~m[590])|(m[568]&m[569]&m[570]&~m[571]&~m[590])|(m[568]&m[569]&m[570]&m[571]&~m[590])|(m[568]&m[569]&~m[570]&~m[571]&m[590])|(m[568]&~m[569]&m[570]&~m[571]&m[590])|(~m[568]&m[569]&m[570]&~m[571]&m[590])|(m[568]&m[569]&m[570]&~m[571]&m[590])|(m[568]&m[569]&m[570]&m[571]&m[590]))):InitCond[1029];
    m[577] = run?((((m[573]&~m[574]&~m[575]&~m[576]&~m[595])|(~m[573]&m[574]&~m[575]&~m[576]&~m[595])|(~m[573]&~m[574]&m[575]&~m[576]&~m[595])|(m[573]&m[574]&~m[575]&m[576]&~m[595])|(m[573]&~m[574]&m[575]&m[576]&~m[595])|(~m[573]&m[574]&m[575]&m[576]&~m[595]))&BiasedRNG[536])|(((m[573]&~m[574]&~m[575]&~m[576]&m[595])|(~m[573]&m[574]&~m[575]&~m[576]&m[595])|(~m[573]&~m[574]&m[575]&~m[576]&m[595])|(m[573]&m[574]&~m[575]&m[576]&m[595])|(m[573]&~m[574]&m[575]&m[576]&m[595])|(~m[573]&m[574]&m[575]&m[576]&m[595]))&~BiasedRNG[536])|((m[573]&m[574]&~m[575]&~m[576]&~m[595])|(m[573]&~m[574]&m[575]&~m[576]&~m[595])|(~m[573]&m[574]&m[575]&~m[576]&~m[595])|(m[573]&m[574]&m[575]&~m[576]&~m[595])|(m[573]&m[574]&m[575]&m[576]&~m[595])|(m[573]&m[574]&~m[575]&~m[576]&m[595])|(m[573]&~m[574]&m[575]&~m[576]&m[595])|(~m[573]&m[574]&m[575]&~m[576]&m[595])|(m[573]&m[574]&m[575]&~m[576]&m[595])|(m[573]&m[574]&m[575]&m[576]&m[595]))):InitCond[1030];
    m[582] = run?((((m[578]&~m[579]&~m[580]&~m[581]&~m[605])|(~m[578]&m[579]&~m[580]&~m[581]&~m[605])|(~m[578]&~m[579]&m[580]&~m[581]&~m[605])|(m[578]&m[579]&~m[580]&m[581]&~m[605])|(m[578]&~m[579]&m[580]&m[581]&~m[605])|(~m[578]&m[579]&m[580]&m[581]&~m[605]))&BiasedRNG[537])|(((m[578]&~m[579]&~m[580]&~m[581]&m[605])|(~m[578]&m[579]&~m[580]&~m[581]&m[605])|(~m[578]&~m[579]&m[580]&~m[581]&m[605])|(m[578]&m[579]&~m[580]&m[581]&m[605])|(m[578]&~m[579]&m[580]&m[581]&m[605])|(~m[578]&m[579]&m[580]&m[581]&m[605]))&~BiasedRNG[537])|((m[578]&m[579]&~m[580]&~m[581]&~m[605])|(m[578]&~m[579]&m[580]&~m[581]&~m[605])|(~m[578]&m[579]&m[580]&~m[581]&~m[605])|(m[578]&m[579]&m[580]&~m[581]&~m[605])|(m[578]&m[579]&m[580]&m[581]&~m[605])|(m[578]&m[579]&~m[580]&~m[581]&m[605])|(m[578]&~m[579]&m[580]&~m[581]&m[605])|(~m[578]&m[579]&m[580]&~m[581]&m[605])|(m[578]&m[579]&m[580]&~m[581]&m[605])|(m[578]&m[579]&m[580]&m[581]&m[605]))):InitCond[1031];
    m[587] = run?((((m[583]&~m[584]&~m[585]&~m[586]&~m[610])|(~m[583]&m[584]&~m[585]&~m[586]&~m[610])|(~m[583]&~m[584]&m[585]&~m[586]&~m[610])|(m[583]&m[584]&~m[585]&m[586]&~m[610])|(m[583]&~m[584]&m[585]&m[586]&~m[610])|(~m[583]&m[584]&m[585]&m[586]&~m[610]))&BiasedRNG[538])|(((m[583]&~m[584]&~m[585]&~m[586]&m[610])|(~m[583]&m[584]&~m[585]&~m[586]&m[610])|(~m[583]&~m[584]&m[585]&~m[586]&m[610])|(m[583]&m[584]&~m[585]&m[586]&m[610])|(m[583]&~m[584]&m[585]&m[586]&m[610])|(~m[583]&m[584]&m[585]&m[586]&m[610]))&~BiasedRNG[538])|((m[583]&m[584]&~m[585]&~m[586]&~m[610])|(m[583]&~m[584]&m[585]&~m[586]&~m[610])|(~m[583]&m[584]&m[585]&~m[586]&~m[610])|(m[583]&m[584]&m[585]&~m[586]&~m[610])|(m[583]&m[584]&m[585]&m[586]&~m[610])|(m[583]&m[584]&~m[585]&~m[586]&m[610])|(m[583]&~m[584]&m[585]&~m[586]&m[610])|(~m[583]&m[584]&m[585]&~m[586]&m[610])|(m[583]&m[584]&m[585]&~m[586]&m[610])|(m[583]&m[584]&m[585]&m[586]&m[610]))):InitCond[1032];
    m[592] = run?((((m[588]&~m[589]&~m[590]&~m[591]&~m[615])|(~m[588]&m[589]&~m[590]&~m[591]&~m[615])|(~m[588]&~m[589]&m[590]&~m[591]&~m[615])|(m[588]&m[589]&~m[590]&m[591]&~m[615])|(m[588]&~m[589]&m[590]&m[591]&~m[615])|(~m[588]&m[589]&m[590]&m[591]&~m[615]))&BiasedRNG[539])|(((m[588]&~m[589]&~m[590]&~m[591]&m[615])|(~m[588]&m[589]&~m[590]&~m[591]&m[615])|(~m[588]&~m[589]&m[590]&~m[591]&m[615])|(m[588]&m[589]&~m[590]&m[591]&m[615])|(m[588]&~m[589]&m[590]&m[591]&m[615])|(~m[588]&m[589]&m[590]&m[591]&m[615]))&~BiasedRNG[539])|((m[588]&m[589]&~m[590]&~m[591]&~m[615])|(m[588]&~m[589]&m[590]&~m[591]&~m[615])|(~m[588]&m[589]&m[590]&~m[591]&~m[615])|(m[588]&m[589]&m[590]&~m[591]&~m[615])|(m[588]&m[589]&m[590]&m[591]&~m[615])|(m[588]&m[589]&~m[590]&~m[591]&m[615])|(m[588]&~m[589]&m[590]&~m[591]&m[615])|(~m[588]&m[589]&m[590]&~m[591]&m[615])|(m[588]&m[589]&m[590]&~m[591]&m[615])|(m[588]&m[589]&m[590]&m[591]&m[615]))):InitCond[1033];
    m[597] = run?((((m[593]&~m[594]&~m[595]&~m[596]&~m[620])|(~m[593]&m[594]&~m[595]&~m[596]&~m[620])|(~m[593]&~m[594]&m[595]&~m[596]&~m[620])|(m[593]&m[594]&~m[595]&m[596]&~m[620])|(m[593]&~m[594]&m[595]&m[596]&~m[620])|(~m[593]&m[594]&m[595]&m[596]&~m[620]))&BiasedRNG[540])|(((m[593]&~m[594]&~m[595]&~m[596]&m[620])|(~m[593]&m[594]&~m[595]&~m[596]&m[620])|(~m[593]&~m[594]&m[595]&~m[596]&m[620])|(m[593]&m[594]&~m[595]&m[596]&m[620])|(m[593]&~m[594]&m[595]&m[596]&m[620])|(~m[593]&m[594]&m[595]&m[596]&m[620]))&~BiasedRNG[540])|((m[593]&m[594]&~m[595]&~m[596]&~m[620])|(m[593]&~m[594]&m[595]&~m[596]&~m[620])|(~m[593]&m[594]&m[595]&~m[596]&~m[620])|(m[593]&m[594]&m[595]&~m[596]&~m[620])|(m[593]&m[594]&m[595]&m[596]&~m[620])|(m[593]&m[594]&~m[595]&~m[596]&m[620])|(m[593]&~m[594]&m[595]&~m[596]&m[620])|(~m[593]&m[594]&m[595]&~m[596]&m[620])|(m[593]&m[594]&m[595]&~m[596]&m[620])|(m[593]&m[594]&m[595]&m[596]&m[620]))):InitCond[1034];
    m[602] = run?((((m[598]&~m[599]&~m[600]&~m[601]&~m[625])|(~m[598]&m[599]&~m[600]&~m[601]&~m[625])|(~m[598]&~m[599]&m[600]&~m[601]&~m[625])|(m[598]&m[599]&~m[600]&m[601]&~m[625])|(m[598]&~m[599]&m[600]&m[601]&~m[625])|(~m[598]&m[599]&m[600]&m[601]&~m[625]))&BiasedRNG[541])|(((m[598]&~m[599]&~m[600]&~m[601]&m[625])|(~m[598]&m[599]&~m[600]&~m[601]&m[625])|(~m[598]&~m[599]&m[600]&~m[601]&m[625])|(m[598]&m[599]&~m[600]&m[601]&m[625])|(m[598]&~m[599]&m[600]&m[601]&m[625])|(~m[598]&m[599]&m[600]&m[601]&m[625]))&~BiasedRNG[541])|((m[598]&m[599]&~m[600]&~m[601]&~m[625])|(m[598]&~m[599]&m[600]&~m[601]&~m[625])|(~m[598]&m[599]&m[600]&~m[601]&~m[625])|(m[598]&m[599]&m[600]&~m[601]&~m[625])|(m[598]&m[599]&m[600]&m[601]&~m[625])|(m[598]&m[599]&~m[600]&~m[601]&m[625])|(m[598]&~m[599]&m[600]&~m[601]&m[625])|(~m[598]&m[599]&m[600]&~m[601]&m[625])|(m[598]&m[599]&m[600]&~m[601]&m[625])|(m[598]&m[599]&m[600]&m[601]&m[625]))):InitCond[1035];
    m[607] = run?((((m[603]&~m[604]&~m[605]&~m[606]&~m[635])|(~m[603]&m[604]&~m[605]&~m[606]&~m[635])|(~m[603]&~m[604]&m[605]&~m[606]&~m[635])|(m[603]&m[604]&~m[605]&m[606]&~m[635])|(m[603]&~m[604]&m[605]&m[606]&~m[635])|(~m[603]&m[604]&m[605]&m[606]&~m[635]))&BiasedRNG[542])|(((m[603]&~m[604]&~m[605]&~m[606]&m[635])|(~m[603]&m[604]&~m[605]&~m[606]&m[635])|(~m[603]&~m[604]&m[605]&~m[606]&m[635])|(m[603]&m[604]&~m[605]&m[606]&m[635])|(m[603]&~m[604]&m[605]&m[606]&m[635])|(~m[603]&m[604]&m[605]&m[606]&m[635]))&~BiasedRNG[542])|((m[603]&m[604]&~m[605]&~m[606]&~m[635])|(m[603]&~m[604]&m[605]&~m[606]&~m[635])|(~m[603]&m[604]&m[605]&~m[606]&~m[635])|(m[603]&m[604]&m[605]&~m[606]&~m[635])|(m[603]&m[604]&m[605]&m[606]&~m[635])|(m[603]&m[604]&~m[605]&~m[606]&m[635])|(m[603]&~m[604]&m[605]&~m[606]&m[635])|(~m[603]&m[604]&m[605]&~m[606]&m[635])|(m[603]&m[604]&m[605]&~m[606]&m[635])|(m[603]&m[604]&m[605]&m[606]&m[635]))):InitCond[1036];
    m[612] = run?((((m[608]&~m[609]&~m[610]&~m[611]&~m[640])|(~m[608]&m[609]&~m[610]&~m[611]&~m[640])|(~m[608]&~m[609]&m[610]&~m[611]&~m[640])|(m[608]&m[609]&~m[610]&m[611]&~m[640])|(m[608]&~m[609]&m[610]&m[611]&~m[640])|(~m[608]&m[609]&m[610]&m[611]&~m[640]))&BiasedRNG[543])|(((m[608]&~m[609]&~m[610]&~m[611]&m[640])|(~m[608]&m[609]&~m[610]&~m[611]&m[640])|(~m[608]&~m[609]&m[610]&~m[611]&m[640])|(m[608]&m[609]&~m[610]&m[611]&m[640])|(m[608]&~m[609]&m[610]&m[611]&m[640])|(~m[608]&m[609]&m[610]&m[611]&m[640]))&~BiasedRNG[543])|((m[608]&m[609]&~m[610]&~m[611]&~m[640])|(m[608]&~m[609]&m[610]&~m[611]&~m[640])|(~m[608]&m[609]&m[610]&~m[611]&~m[640])|(m[608]&m[609]&m[610]&~m[611]&~m[640])|(m[608]&m[609]&m[610]&m[611]&~m[640])|(m[608]&m[609]&~m[610]&~m[611]&m[640])|(m[608]&~m[609]&m[610]&~m[611]&m[640])|(~m[608]&m[609]&m[610]&~m[611]&m[640])|(m[608]&m[609]&m[610]&~m[611]&m[640])|(m[608]&m[609]&m[610]&m[611]&m[640]))):InitCond[1037];
    m[617] = run?((((m[613]&~m[614]&~m[615]&~m[616]&~m[645])|(~m[613]&m[614]&~m[615]&~m[616]&~m[645])|(~m[613]&~m[614]&m[615]&~m[616]&~m[645])|(m[613]&m[614]&~m[615]&m[616]&~m[645])|(m[613]&~m[614]&m[615]&m[616]&~m[645])|(~m[613]&m[614]&m[615]&m[616]&~m[645]))&BiasedRNG[544])|(((m[613]&~m[614]&~m[615]&~m[616]&m[645])|(~m[613]&m[614]&~m[615]&~m[616]&m[645])|(~m[613]&~m[614]&m[615]&~m[616]&m[645])|(m[613]&m[614]&~m[615]&m[616]&m[645])|(m[613]&~m[614]&m[615]&m[616]&m[645])|(~m[613]&m[614]&m[615]&m[616]&m[645]))&~BiasedRNG[544])|((m[613]&m[614]&~m[615]&~m[616]&~m[645])|(m[613]&~m[614]&m[615]&~m[616]&~m[645])|(~m[613]&m[614]&m[615]&~m[616]&~m[645])|(m[613]&m[614]&m[615]&~m[616]&~m[645])|(m[613]&m[614]&m[615]&m[616]&~m[645])|(m[613]&m[614]&~m[615]&~m[616]&m[645])|(m[613]&~m[614]&m[615]&~m[616]&m[645])|(~m[613]&m[614]&m[615]&~m[616]&m[645])|(m[613]&m[614]&m[615]&~m[616]&m[645])|(m[613]&m[614]&m[615]&m[616]&m[645]))):InitCond[1038];
    m[622] = run?((((m[618]&~m[619]&~m[620]&~m[621]&~m[650])|(~m[618]&m[619]&~m[620]&~m[621]&~m[650])|(~m[618]&~m[619]&m[620]&~m[621]&~m[650])|(m[618]&m[619]&~m[620]&m[621]&~m[650])|(m[618]&~m[619]&m[620]&m[621]&~m[650])|(~m[618]&m[619]&m[620]&m[621]&~m[650]))&BiasedRNG[545])|(((m[618]&~m[619]&~m[620]&~m[621]&m[650])|(~m[618]&m[619]&~m[620]&~m[621]&m[650])|(~m[618]&~m[619]&m[620]&~m[621]&m[650])|(m[618]&m[619]&~m[620]&m[621]&m[650])|(m[618]&~m[619]&m[620]&m[621]&m[650])|(~m[618]&m[619]&m[620]&m[621]&m[650]))&~BiasedRNG[545])|((m[618]&m[619]&~m[620]&~m[621]&~m[650])|(m[618]&~m[619]&m[620]&~m[621]&~m[650])|(~m[618]&m[619]&m[620]&~m[621]&~m[650])|(m[618]&m[619]&m[620]&~m[621]&~m[650])|(m[618]&m[619]&m[620]&m[621]&~m[650])|(m[618]&m[619]&~m[620]&~m[621]&m[650])|(m[618]&~m[619]&m[620]&~m[621]&m[650])|(~m[618]&m[619]&m[620]&~m[621]&m[650])|(m[618]&m[619]&m[620]&~m[621]&m[650])|(m[618]&m[619]&m[620]&m[621]&m[650]))):InitCond[1039];
    m[627] = run?((((m[623]&~m[624]&~m[625]&~m[626]&~m[655])|(~m[623]&m[624]&~m[625]&~m[626]&~m[655])|(~m[623]&~m[624]&m[625]&~m[626]&~m[655])|(m[623]&m[624]&~m[625]&m[626]&~m[655])|(m[623]&~m[624]&m[625]&m[626]&~m[655])|(~m[623]&m[624]&m[625]&m[626]&~m[655]))&BiasedRNG[546])|(((m[623]&~m[624]&~m[625]&~m[626]&m[655])|(~m[623]&m[624]&~m[625]&~m[626]&m[655])|(~m[623]&~m[624]&m[625]&~m[626]&m[655])|(m[623]&m[624]&~m[625]&m[626]&m[655])|(m[623]&~m[624]&m[625]&m[626]&m[655])|(~m[623]&m[624]&m[625]&m[626]&m[655]))&~BiasedRNG[546])|((m[623]&m[624]&~m[625]&~m[626]&~m[655])|(m[623]&~m[624]&m[625]&~m[626]&~m[655])|(~m[623]&m[624]&m[625]&~m[626]&~m[655])|(m[623]&m[624]&m[625]&~m[626]&~m[655])|(m[623]&m[624]&m[625]&m[626]&~m[655])|(m[623]&m[624]&~m[625]&~m[626]&m[655])|(m[623]&~m[624]&m[625]&~m[626]&m[655])|(~m[623]&m[624]&m[625]&~m[626]&m[655])|(m[623]&m[624]&m[625]&~m[626]&m[655])|(m[623]&m[624]&m[625]&m[626]&m[655]))):InitCond[1040];
    m[632] = run?((((m[628]&~m[629]&~m[630]&~m[631]&~m[660])|(~m[628]&m[629]&~m[630]&~m[631]&~m[660])|(~m[628]&~m[629]&m[630]&~m[631]&~m[660])|(m[628]&m[629]&~m[630]&m[631]&~m[660])|(m[628]&~m[629]&m[630]&m[631]&~m[660])|(~m[628]&m[629]&m[630]&m[631]&~m[660]))&BiasedRNG[547])|(((m[628]&~m[629]&~m[630]&~m[631]&m[660])|(~m[628]&m[629]&~m[630]&~m[631]&m[660])|(~m[628]&~m[629]&m[630]&~m[631]&m[660])|(m[628]&m[629]&~m[630]&m[631]&m[660])|(m[628]&~m[629]&m[630]&m[631]&m[660])|(~m[628]&m[629]&m[630]&m[631]&m[660]))&~BiasedRNG[547])|((m[628]&m[629]&~m[630]&~m[631]&~m[660])|(m[628]&~m[629]&m[630]&~m[631]&~m[660])|(~m[628]&m[629]&m[630]&~m[631]&~m[660])|(m[628]&m[629]&m[630]&~m[631]&~m[660])|(m[628]&m[629]&m[630]&m[631]&~m[660])|(m[628]&m[629]&~m[630]&~m[631]&m[660])|(m[628]&~m[629]&m[630]&~m[631]&m[660])|(~m[628]&m[629]&m[630]&~m[631]&m[660])|(m[628]&m[629]&m[630]&~m[631]&m[660])|(m[628]&m[629]&m[630]&m[631]&m[660]))):InitCond[1041];
    m[637] = run?((((m[633]&~m[634]&~m[635]&~m[636]&~m[670])|(~m[633]&m[634]&~m[635]&~m[636]&~m[670])|(~m[633]&~m[634]&m[635]&~m[636]&~m[670])|(m[633]&m[634]&~m[635]&m[636]&~m[670])|(m[633]&~m[634]&m[635]&m[636]&~m[670])|(~m[633]&m[634]&m[635]&m[636]&~m[670]))&BiasedRNG[548])|(((m[633]&~m[634]&~m[635]&~m[636]&m[670])|(~m[633]&m[634]&~m[635]&~m[636]&m[670])|(~m[633]&~m[634]&m[635]&~m[636]&m[670])|(m[633]&m[634]&~m[635]&m[636]&m[670])|(m[633]&~m[634]&m[635]&m[636]&m[670])|(~m[633]&m[634]&m[635]&m[636]&m[670]))&~BiasedRNG[548])|((m[633]&m[634]&~m[635]&~m[636]&~m[670])|(m[633]&~m[634]&m[635]&~m[636]&~m[670])|(~m[633]&m[634]&m[635]&~m[636]&~m[670])|(m[633]&m[634]&m[635]&~m[636]&~m[670])|(m[633]&m[634]&m[635]&m[636]&~m[670])|(m[633]&m[634]&~m[635]&~m[636]&m[670])|(m[633]&~m[634]&m[635]&~m[636]&m[670])|(~m[633]&m[634]&m[635]&~m[636]&m[670])|(m[633]&m[634]&m[635]&~m[636]&m[670])|(m[633]&m[634]&m[635]&m[636]&m[670]))):InitCond[1042];
    m[642] = run?((((m[638]&~m[639]&~m[640]&~m[641]&~m[675])|(~m[638]&m[639]&~m[640]&~m[641]&~m[675])|(~m[638]&~m[639]&m[640]&~m[641]&~m[675])|(m[638]&m[639]&~m[640]&m[641]&~m[675])|(m[638]&~m[639]&m[640]&m[641]&~m[675])|(~m[638]&m[639]&m[640]&m[641]&~m[675]))&BiasedRNG[549])|(((m[638]&~m[639]&~m[640]&~m[641]&m[675])|(~m[638]&m[639]&~m[640]&~m[641]&m[675])|(~m[638]&~m[639]&m[640]&~m[641]&m[675])|(m[638]&m[639]&~m[640]&m[641]&m[675])|(m[638]&~m[639]&m[640]&m[641]&m[675])|(~m[638]&m[639]&m[640]&m[641]&m[675]))&~BiasedRNG[549])|((m[638]&m[639]&~m[640]&~m[641]&~m[675])|(m[638]&~m[639]&m[640]&~m[641]&~m[675])|(~m[638]&m[639]&m[640]&~m[641]&~m[675])|(m[638]&m[639]&m[640]&~m[641]&~m[675])|(m[638]&m[639]&m[640]&m[641]&~m[675])|(m[638]&m[639]&~m[640]&~m[641]&m[675])|(m[638]&~m[639]&m[640]&~m[641]&m[675])|(~m[638]&m[639]&m[640]&~m[641]&m[675])|(m[638]&m[639]&m[640]&~m[641]&m[675])|(m[638]&m[639]&m[640]&m[641]&m[675]))):InitCond[1043];
    m[647] = run?((((m[643]&~m[644]&~m[645]&~m[646]&~m[680])|(~m[643]&m[644]&~m[645]&~m[646]&~m[680])|(~m[643]&~m[644]&m[645]&~m[646]&~m[680])|(m[643]&m[644]&~m[645]&m[646]&~m[680])|(m[643]&~m[644]&m[645]&m[646]&~m[680])|(~m[643]&m[644]&m[645]&m[646]&~m[680]))&BiasedRNG[550])|(((m[643]&~m[644]&~m[645]&~m[646]&m[680])|(~m[643]&m[644]&~m[645]&~m[646]&m[680])|(~m[643]&~m[644]&m[645]&~m[646]&m[680])|(m[643]&m[644]&~m[645]&m[646]&m[680])|(m[643]&~m[644]&m[645]&m[646]&m[680])|(~m[643]&m[644]&m[645]&m[646]&m[680]))&~BiasedRNG[550])|((m[643]&m[644]&~m[645]&~m[646]&~m[680])|(m[643]&~m[644]&m[645]&~m[646]&~m[680])|(~m[643]&m[644]&m[645]&~m[646]&~m[680])|(m[643]&m[644]&m[645]&~m[646]&~m[680])|(m[643]&m[644]&m[645]&m[646]&~m[680])|(m[643]&m[644]&~m[645]&~m[646]&m[680])|(m[643]&~m[644]&m[645]&~m[646]&m[680])|(~m[643]&m[644]&m[645]&~m[646]&m[680])|(m[643]&m[644]&m[645]&~m[646]&m[680])|(m[643]&m[644]&m[645]&m[646]&m[680]))):InitCond[1044];
    m[652] = run?((((m[648]&~m[649]&~m[650]&~m[651]&~m[685])|(~m[648]&m[649]&~m[650]&~m[651]&~m[685])|(~m[648]&~m[649]&m[650]&~m[651]&~m[685])|(m[648]&m[649]&~m[650]&m[651]&~m[685])|(m[648]&~m[649]&m[650]&m[651]&~m[685])|(~m[648]&m[649]&m[650]&m[651]&~m[685]))&BiasedRNG[551])|(((m[648]&~m[649]&~m[650]&~m[651]&m[685])|(~m[648]&m[649]&~m[650]&~m[651]&m[685])|(~m[648]&~m[649]&m[650]&~m[651]&m[685])|(m[648]&m[649]&~m[650]&m[651]&m[685])|(m[648]&~m[649]&m[650]&m[651]&m[685])|(~m[648]&m[649]&m[650]&m[651]&m[685]))&~BiasedRNG[551])|((m[648]&m[649]&~m[650]&~m[651]&~m[685])|(m[648]&~m[649]&m[650]&~m[651]&~m[685])|(~m[648]&m[649]&m[650]&~m[651]&~m[685])|(m[648]&m[649]&m[650]&~m[651]&~m[685])|(m[648]&m[649]&m[650]&m[651]&~m[685])|(m[648]&m[649]&~m[650]&~m[651]&m[685])|(m[648]&~m[649]&m[650]&~m[651]&m[685])|(~m[648]&m[649]&m[650]&~m[651]&m[685])|(m[648]&m[649]&m[650]&~m[651]&m[685])|(m[648]&m[649]&m[650]&m[651]&m[685]))):InitCond[1045];
    m[657] = run?((((m[653]&~m[654]&~m[655]&~m[656]&~m[690])|(~m[653]&m[654]&~m[655]&~m[656]&~m[690])|(~m[653]&~m[654]&m[655]&~m[656]&~m[690])|(m[653]&m[654]&~m[655]&m[656]&~m[690])|(m[653]&~m[654]&m[655]&m[656]&~m[690])|(~m[653]&m[654]&m[655]&m[656]&~m[690]))&BiasedRNG[552])|(((m[653]&~m[654]&~m[655]&~m[656]&m[690])|(~m[653]&m[654]&~m[655]&~m[656]&m[690])|(~m[653]&~m[654]&m[655]&~m[656]&m[690])|(m[653]&m[654]&~m[655]&m[656]&m[690])|(m[653]&~m[654]&m[655]&m[656]&m[690])|(~m[653]&m[654]&m[655]&m[656]&m[690]))&~BiasedRNG[552])|((m[653]&m[654]&~m[655]&~m[656]&~m[690])|(m[653]&~m[654]&m[655]&~m[656]&~m[690])|(~m[653]&m[654]&m[655]&~m[656]&~m[690])|(m[653]&m[654]&m[655]&~m[656]&~m[690])|(m[653]&m[654]&m[655]&m[656]&~m[690])|(m[653]&m[654]&~m[655]&~m[656]&m[690])|(m[653]&~m[654]&m[655]&~m[656]&m[690])|(~m[653]&m[654]&m[655]&~m[656]&m[690])|(m[653]&m[654]&m[655]&~m[656]&m[690])|(m[653]&m[654]&m[655]&m[656]&m[690]))):InitCond[1046];
    m[662] = run?((((m[658]&~m[659]&~m[660]&~m[661]&~m[695])|(~m[658]&m[659]&~m[660]&~m[661]&~m[695])|(~m[658]&~m[659]&m[660]&~m[661]&~m[695])|(m[658]&m[659]&~m[660]&m[661]&~m[695])|(m[658]&~m[659]&m[660]&m[661]&~m[695])|(~m[658]&m[659]&m[660]&m[661]&~m[695]))&BiasedRNG[553])|(((m[658]&~m[659]&~m[660]&~m[661]&m[695])|(~m[658]&m[659]&~m[660]&~m[661]&m[695])|(~m[658]&~m[659]&m[660]&~m[661]&m[695])|(m[658]&m[659]&~m[660]&m[661]&m[695])|(m[658]&~m[659]&m[660]&m[661]&m[695])|(~m[658]&m[659]&m[660]&m[661]&m[695]))&~BiasedRNG[553])|((m[658]&m[659]&~m[660]&~m[661]&~m[695])|(m[658]&~m[659]&m[660]&~m[661]&~m[695])|(~m[658]&m[659]&m[660]&~m[661]&~m[695])|(m[658]&m[659]&m[660]&~m[661]&~m[695])|(m[658]&m[659]&m[660]&m[661]&~m[695])|(m[658]&m[659]&~m[660]&~m[661]&m[695])|(m[658]&~m[659]&m[660]&~m[661]&m[695])|(~m[658]&m[659]&m[660]&~m[661]&m[695])|(m[658]&m[659]&m[660]&~m[661]&m[695])|(m[658]&m[659]&m[660]&m[661]&m[695]))):InitCond[1047];
    m[667] = run?((((m[663]&~m[664]&~m[665]&~m[666]&~m[700])|(~m[663]&m[664]&~m[665]&~m[666]&~m[700])|(~m[663]&~m[664]&m[665]&~m[666]&~m[700])|(m[663]&m[664]&~m[665]&m[666]&~m[700])|(m[663]&~m[664]&m[665]&m[666]&~m[700])|(~m[663]&m[664]&m[665]&m[666]&~m[700]))&BiasedRNG[554])|(((m[663]&~m[664]&~m[665]&~m[666]&m[700])|(~m[663]&m[664]&~m[665]&~m[666]&m[700])|(~m[663]&~m[664]&m[665]&~m[666]&m[700])|(m[663]&m[664]&~m[665]&m[666]&m[700])|(m[663]&~m[664]&m[665]&m[666]&m[700])|(~m[663]&m[664]&m[665]&m[666]&m[700]))&~BiasedRNG[554])|((m[663]&m[664]&~m[665]&~m[666]&~m[700])|(m[663]&~m[664]&m[665]&~m[666]&~m[700])|(~m[663]&m[664]&m[665]&~m[666]&~m[700])|(m[663]&m[664]&m[665]&~m[666]&~m[700])|(m[663]&m[664]&m[665]&m[666]&~m[700])|(m[663]&m[664]&~m[665]&~m[666]&m[700])|(m[663]&~m[664]&m[665]&~m[666]&m[700])|(~m[663]&m[664]&m[665]&~m[666]&m[700])|(m[663]&m[664]&m[665]&~m[666]&m[700])|(m[663]&m[664]&m[665]&m[666]&m[700]))):InitCond[1048];
    m[672] = run?((((m[668]&~m[669]&~m[670]&~m[671]&~m[710])|(~m[668]&m[669]&~m[670]&~m[671]&~m[710])|(~m[668]&~m[669]&m[670]&~m[671]&~m[710])|(m[668]&m[669]&~m[670]&m[671]&~m[710])|(m[668]&~m[669]&m[670]&m[671]&~m[710])|(~m[668]&m[669]&m[670]&m[671]&~m[710]))&BiasedRNG[555])|(((m[668]&~m[669]&~m[670]&~m[671]&m[710])|(~m[668]&m[669]&~m[670]&~m[671]&m[710])|(~m[668]&~m[669]&m[670]&~m[671]&m[710])|(m[668]&m[669]&~m[670]&m[671]&m[710])|(m[668]&~m[669]&m[670]&m[671]&m[710])|(~m[668]&m[669]&m[670]&m[671]&m[710]))&~BiasedRNG[555])|((m[668]&m[669]&~m[670]&~m[671]&~m[710])|(m[668]&~m[669]&m[670]&~m[671]&~m[710])|(~m[668]&m[669]&m[670]&~m[671]&~m[710])|(m[668]&m[669]&m[670]&~m[671]&~m[710])|(m[668]&m[669]&m[670]&m[671]&~m[710])|(m[668]&m[669]&~m[670]&~m[671]&m[710])|(m[668]&~m[669]&m[670]&~m[671]&m[710])|(~m[668]&m[669]&m[670]&~m[671]&m[710])|(m[668]&m[669]&m[670]&~m[671]&m[710])|(m[668]&m[669]&m[670]&m[671]&m[710]))):InitCond[1049];
    m[677] = run?((((m[673]&~m[674]&~m[675]&~m[676]&~m[715])|(~m[673]&m[674]&~m[675]&~m[676]&~m[715])|(~m[673]&~m[674]&m[675]&~m[676]&~m[715])|(m[673]&m[674]&~m[675]&m[676]&~m[715])|(m[673]&~m[674]&m[675]&m[676]&~m[715])|(~m[673]&m[674]&m[675]&m[676]&~m[715]))&BiasedRNG[556])|(((m[673]&~m[674]&~m[675]&~m[676]&m[715])|(~m[673]&m[674]&~m[675]&~m[676]&m[715])|(~m[673]&~m[674]&m[675]&~m[676]&m[715])|(m[673]&m[674]&~m[675]&m[676]&m[715])|(m[673]&~m[674]&m[675]&m[676]&m[715])|(~m[673]&m[674]&m[675]&m[676]&m[715]))&~BiasedRNG[556])|((m[673]&m[674]&~m[675]&~m[676]&~m[715])|(m[673]&~m[674]&m[675]&~m[676]&~m[715])|(~m[673]&m[674]&m[675]&~m[676]&~m[715])|(m[673]&m[674]&m[675]&~m[676]&~m[715])|(m[673]&m[674]&m[675]&m[676]&~m[715])|(m[673]&m[674]&~m[675]&~m[676]&m[715])|(m[673]&~m[674]&m[675]&~m[676]&m[715])|(~m[673]&m[674]&m[675]&~m[676]&m[715])|(m[673]&m[674]&m[675]&~m[676]&m[715])|(m[673]&m[674]&m[675]&m[676]&m[715]))):InitCond[1050];
    m[682] = run?((((m[678]&~m[679]&~m[680]&~m[681]&~m[720])|(~m[678]&m[679]&~m[680]&~m[681]&~m[720])|(~m[678]&~m[679]&m[680]&~m[681]&~m[720])|(m[678]&m[679]&~m[680]&m[681]&~m[720])|(m[678]&~m[679]&m[680]&m[681]&~m[720])|(~m[678]&m[679]&m[680]&m[681]&~m[720]))&BiasedRNG[557])|(((m[678]&~m[679]&~m[680]&~m[681]&m[720])|(~m[678]&m[679]&~m[680]&~m[681]&m[720])|(~m[678]&~m[679]&m[680]&~m[681]&m[720])|(m[678]&m[679]&~m[680]&m[681]&m[720])|(m[678]&~m[679]&m[680]&m[681]&m[720])|(~m[678]&m[679]&m[680]&m[681]&m[720]))&~BiasedRNG[557])|((m[678]&m[679]&~m[680]&~m[681]&~m[720])|(m[678]&~m[679]&m[680]&~m[681]&~m[720])|(~m[678]&m[679]&m[680]&~m[681]&~m[720])|(m[678]&m[679]&m[680]&~m[681]&~m[720])|(m[678]&m[679]&m[680]&m[681]&~m[720])|(m[678]&m[679]&~m[680]&~m[681]&m[720])|(m[678]&~m[679]&m[680]&~m[681]&m[720])|(~m[678]&m[679]&m[680]&~m[681]&m[720])|(m[678]&m[679]&m[680]&~m[681]&m[720])|(m[678]&m[679]&m[680]&m[681]&m[720]))):InitCond[1051];
    m[687] = run?((((m[683]&~m[684]&~m[685]&~m[686]&~m[725])|(~m[683]&m[684]&~m[685]&~m[686]&~m[725])|(~m[683]&~m[684]&m[685]&~m[686]&~m[725])|(m[683]&m[684]&~m[685]&m[686]&~m[725])|(m[683]&~m[684]&m[685]&m[686]&~m[725])|(~m[683]&m[684]&m[685]&m[686]&~m[725]))&BiasedRNG[558])|(((m[683]&~m[684]&~m[685]&~m[686]&m[725])|(~m[683]&m[684]&~m[685]&~m[686]&m[725])|(~m[683]&~m[684]&m[685]&~m[686]&m[725])|(m[683]&m[684]&~m[685]&m[686]&m[725])|(m[683]&~m[684]&m[685]&m[686]&m[725])|(~m[683]&m[684]&m[685]&m[686]&m[725]))&~BiasedRNG[558])|((m[683]&m[684]&~m[685]&~m[686]&~m[725])|(m[683]&~m[684]&m[685]&~m[686]&~m[725])|(~m[683]&m[684]&m[685]&~m[686]&~m[725])|(m[683]&m[684]&m[685]&~m[686]&~m[725])|(m[683]&m[684]&m[685]&m[686]&~m[725])|(m[683]&m[684]&~m[685]&~m[686]&m[725])|(m[683]&~m[684]&m[685]&~m[686]&m[725])|(~m[683]&m[684]&m[685]&~m[686]&m[725])|(m[683]&m[684]&m[685]&~m[686]&m[725])|(m[683]&m[684]&m[685]&m[686]&m[725]))):InitCond[1052];
    m[692] = run?((((m[688]&~m[689]&~m[690]&~m[691]&~m[730])|(~m[688]&m[689]&~m[690]&~m[691]&~m[730])|(~m[688]&~m[689]&m[690]&~m[691]&~m[730])|(m[688]&m[689]&~m[690]&m[691]&~m[730])|(m[688]&~m[689]&m[690]&m[691]&~m[730])|(~m[688]&m[689]&m[690]&m[691]&~m[730]))&BiasedRNG[559])|(((m[688]&~m[689]&~m[690]&~m[691]&m[730])|(~m[688]&m[689]&~m[690]&~m[691]&m[730])|(~m[688]&~m[689]&m[690]&~m[691]&m[730])|(m[688]&m[689]&~m[690]&m[691]&m[730])|(m[688]&~m[689]&m[690]&m[691]&m[730])|(~m[688]&m[689]&m[690]&m[691]&m[730]))&~BiasedRNG[559])|((m[688]&m[689]&~m[690]&~m[691]&~m[730])|(m[688]&~m[689]&m[690]&~m[691]&~m[730])|(~m[688]&m[689]&m[690]&~m[691]&~m[730])|(m[688]&m[689]&m[690]&~m[691]&~m[730])|(m[688]&m[689]&m[690]&m[691]&~m[730])|(m[688]&m[689]&~m[690]&~m[691]&m[730])|(m[688]&~m[689]&m[690]&~m[691]&m[730])|(~m[688]&m[689]&m[690]&~m[691]&m[730])|(m[688]&m[689]&m[690]&~m[691]&m[730])|(m[688]&m[689]&m[690]&m[691]&m[730]))):InitCond[1053];
    m[697] = run?((((m[693]&~m[694]&~m[695]&~m[696]&~m[735])|(~m[693]&m[694]&~m[695]&~m[696]&~m[735])|(~m[693]&~m[694]&m[695]&~m[696]&~m[735])|(m[693]&m[694]&~m[695]&m[696]&~m[735])|(m[693]&~m[694]&m[695]&m[696]&~m[735])|(~m[693]&m[694]&m[695]&m[696]&~m[735]))&BiasedRNG[560])|(((m[693]&~m[694]&~m[695]&~m[696]&m[735])|(~m[693]&m[694]&~m[695]&~m[696]&m[735])|(~m[693]&~m[694]&m[695]&~m[696]&m[735])|(m[693]&m[694]&~m[695]&m[696]&m[735])|(m[693]&~m[694]&m[695]&m[696]&m[735])|(~m[693]&m[694]&m[695]&m[696]&m[735]))&~BiasedRNG[560])|((m[693]&m[694]&~m[695]&~m[696]&~m[735])|(m[693]&~m[694]&m[695]&~m[696]&~m[735])|(~m[693]&m[694]&m[695]&~m[696]&~m[735])|(m[693]&m[694]&m[695]&~m[696]&~m[735])|(m[693]&m[694]&m[695]&m[696]&~m[735])|(m[693]&m[694]&~m[695]&~m[696]&m[735])|(m[693]&~m[694]&m[695]&~m[696]&m[735])|(~m[693]&m[694]&m[695]&~m[696]&m[735])|(m[693]&m[694]&m[695]&~m[696]&m[735])|(m[693]&m[694]&m[695]&m[696]&m[735]))):InitCond[1054];
    m[702] = run?((((m[698]&~m[699]&~m[700]&~m[701]&~m[740])|(~m[698]&m[699]&~m[700]&~m[701]&~m[740])|(~m[698]&~m[699]&m[700]&~m[701]&~m[740])|(m[698]&m[699]&~m[700]&m[701]&~m[740])|(m[698]&~m[699]&m[700]&m[701]&~m[740])|(~m[698]&m[699]&m[700]&m[701]&~m[740]))&BiasedRNG[561])|(((m[698]&~m[699]&~m[700]&~m[701]&m[740])|(~m[698]&m[699]&~m[700]&~m[701]&m[740])|(~m[698]&~m[699]&m[700]&~m[701]&m[740])|(m[698]&m[699]&~m[700]&m[701]&m[740])|(m[698]&~m[699]&m[700]&m[701]&m[740])|(~m[698]&m[699]&m[700]&m[701]&m[740]))&~BiasedRNG[561])|((m[698]&m[699]&~m[700]&~m[701]&~m[740])|(m[698]&~m[699]&m[700]&~m[701]&~m[740])|(~m[698]&m[699]&m[700]&~m[701]&~m[740])|(m[698]&m[699]&m[700]&~m[701]&~m[740])|(m[698]&m[699]&m[700]&m[701]&~m[740])|(m[698]&m[699]&~m[700]&~m[701]&m[740])|(m[698]&~m[699]&m[700]&~m[701]&m[740])|(~m[698]&m[699]&m[700]&~m[701]&m[740])|(m[698]&m[699]&m[700]&~m[701]&m[740])|(m[698]&m[699]&m[700]&m[701]&m[740]))):InitCond[1055];
    m[707] = run?((((m[703]&~m[704]&~m[705]&~m[706]&~m[745])|(~m[703]&m[704]&~m[705]&~m[706]&~m[745])|(~m[703]&~m[704]&m[705]&~m[706]&~m[745])|(m[703]&m[704]&~m[705]&m[706]&~m[745])|(m[703]&~m[704]&m[705]&m[706]&~m[745])|(~m[703]&m[704]&m[705]&m[706]&~m[745]))&BiasedRNG[562])|(((m[703]&~m[704]&~m[705]&~m[706]&m[745])|(~m[703]&m[704]&~m[705]&~m[706]&m[745])|(~m[703]&~m[704]&m[705]&~m[706]&m[745])|(m[703]&m[704]&~m[705]&m[706]&m[745])|(m[703]&~m[704]&m[705]&m[706]&m[745])|(~m[703]&m[704]&m[705]&m[706]&m[745]))&~BiasedRNG[562])|((m[703]&m[704]&~m[705]&~m[706]&~m[745])|(m[703]&~m[704]&m[705]&~m[706]&~m[745])|(~m[703]&m[704]&m[705]&~m[706]&~m[745])|(m[703]&m[704]&m[705]&~m[706]&~m[745])|(m[703]&m[704]&m[705]&m[706]&~m[745])|(m[703]&m[704]&~m[705]&~m[706]&m[745])|(m[703]&~m[704]&m[705]&~m[706]&m[745])|(~m[703]&m[704]&m[705]&~m[706]&m[745])|(m[703]&m[704]&m[705]&~m[706]&m[745])|(m[703]&m[704]&m[705]&m[706]&m[745]))):InitCond[1056];
    m[712] = run?((((m[708]&~m[709]&~m[710]&~m[711]&~m[755])|(~m[708]&m[709]&~m[710]&~m[711]&~m[755])|(~m[708]&~m[709]&m[710]&~m[711]&~m[755])|(m[708]&m[709]&~m[710]&m[711]&~m[755])|(m[708]&~m[709]&m[710]&m[711]&~m[755])|(~m[708]&m[709]&m[710]&m[711]&~m[755]))&BiasedRNG[563])|(((m[708]&~m[709]&~m[710]&~m[711]&m[755])|(~m[708]&m[709]&~m[710]&~m[711]&m[755])|(~m[708]&~m[709]&m[710]&~m[711]&m[755])|(m[708]&m[709]&~m[710]&m[711]&m[755])|(m[708]&~m[709]&m[710]&m[711]&m[755])|(~m[708]&m[709]&m[710]&m[711]&m[755]))&~BiasedRNG[563])|((m[708]&m[709]&~m[710]&~m[711]&~m[755])|(m[708]&~m[709]&m[710]&~m[711]&~m[755])|(~m[708]&m[709]&m[710]&~m[711]&~m[755])|(m[708]&m[709]&m[710]&~m[711]&~m[755])|(m[708]&m[709]&m[710]&m[711]&~m[755])|(m[708]&m[709]&~m[710]&~m[711]&m[755])|(m[708]&~m[709]&m[710]&~m[711]&m[755])|(~m[708]&m[709]&m[710]&~m[711]&m[755])|(m[708]&m[709]&m[710]&~m[711]&m[755])|(m[708]&m[709]&m[710]&m[711]&m[755]))):InitCond[1057];
    m[717] = run?((((m[713]&~m[714]&~m[715]&~m[716]&~m[760])|(~m[713]&m[714]&~m[715]&~m[716]&~m[760])|(~m[713]&~m[714]&m[715]&~m[716]&~m[760])|(m[713]&m[714]&~m[715]&m[716]&~m[760])|(m[713]&~m[714]&m[715]&m[716]&~m[760])|(~m[713]&m[714]&m[715]&m[716]&~m[760]))&BiasedRNG[564])|(((m[713]&~m[714]&~m[715]&~m[716]&m[760])|(~m[713]&m[714]&~m[715]&~m[716]&m[760])|(~m[713]&~m[714]&m[715]&~m[716]&m[760])|(m[713]&m[714]&~m[715]&m[716]&m[760])|(m[713]&~m[714]&m[715]&m[716]&m[760])|(~m[713]&m[714]&m[715]&m[716]&m[760]))&~BiasedRNG[564])|((m[713]&m[714]&~m[715]&~m[716]&~m[760])|(m[713]&~m[714]&m[715]&~m[716]&~m[760])|(~m[713]&m[714]&m[715]&~m[716]&~m[760])|(m[713]&m[714]&m[715]&~m[716]&~m[760])|(m[713]&m[714]&m[715]&m[716]&~m[760])|(m[713]&m[714]&~m[715]&~m[716]&m[760])|(m[713]&~m[714]&m[715]&~m[716]&m[760])|(~m[713]&m[714]&m[715]&~m[716]&m[760])|(m[713]&m[714]&m[715]&~m[716]&m[760])|(m[713]&m[714]&m[715]&m[716]&m[760]))):InitCond[1058];
    m[722] = run?((((m[718]&~m[719]&~m[720]&~m[721]&~m[765])|(~m[718]&m[719]&~m[720]&~m[721]&~m[765])|(~m[718]&~m[719]&m[720]&~m[721]&~m[765])|(m[718]&m[719]&~m[720]&m[721]&~m[765])|(m[718]&~m[719]&m[720]&m[721]&~m[765])|(~m[718]&m[719]&m[720]&m[721]&~m[765]))&BiasedRNG[565])|(((m[718]&~m[719]&~m[720]&~m[721]&m[765])|(~m[718]&m[719]&~m[720]&~m[721]&m[765])|(~m[718]&~m[719]&m[720]&~m[721]&m[765])|(m[718]&m[719]&~m[720]&m[721]&m[765])|(m[718]&~m[719]&m[720]&m[721]&m[765])|(~m[718]&m[719]&m[720]&m[721]&m[765]))&~BiasedRNG[565])|((m[718]&m[719]&~m[720]&~m[721]&~m[765])|(m[718]&~m[719]&m[720]&~m[721]&~m[765])|(~m[718]&m[719]&m[720]&~m[721]&~m[765])|(m[718]&m[719]&m[720]&~m[721]&~m[765])|(m[718]&m[719]&m[720]&m[721]&~m[765])|(m[718]&m[719]&~m[720]&~m[721]&m[765])|(m[718]&~m[719]&m[720]&~m[721]&m[765])|(~m[718]&m[719]&m[720]&~m[721]&m[765])|(m[718]&m[719]&m[720]&~m[721]&m[765])|(m[718]&m[719]&m[720]&m[721]&m[765]))):InitCond[1059];
    m[727] = run?((((m[723]&~m[724]&~m[725]&~m[726]&~m[770])|(~m[723]&m[724]&~m[725]&~m[726]&~m[770])|(~m[723]&~m[724]&m[725]&~m[726]&~m[770])|(m[723]&m[724]&~m[725]&m[726]&~m[770])|(m[723]&~m[724]&m[725]&m[726]&~m[770])|(~m[723]&m[724]&m[725]&m[726]&~m[770]))&BiasedRNG[566])|(((m[723]&~m[724]&~m[725]&~m[726]&m[770])|(~m[723]&m[724]&~m[725]&~m[726]&m[770])|(~m[723]&~m[724]&m[725]&~m[726]&m[770])|(m[723]&m[724]&~m[725]&m[726]&m[770])|(m[723]&~m[724]&m[725]&m[726]&m[770])|(~m[723]&m[724]&m[725]&m[726]&m[770]))&~BiasedRNG[566])|((m[723]&m[724]&~m[725]&~m[726]&~m[770])|(m[723]&~m[724]&m[725]&~m[726]&~m[770])|(~m[723]&m[724]&m[725]&~m[726]&~m[770])|(m[723]&m[724]&m[725]&~m[726]&~m[770])|(m[723]&m[724]&m[725]&m[726]&~m[770])|(m[723]&m[724]&~m[725]&~m[726]&m[770])|(m[723]&~m[724]&m[725]&~m[726]&m[770])|(~m[723]&m[724]&m[725]&~m[726]&m[770])|(m[723]&m[724]&m[725]&~m[726]&m[770])|(m[723]&m[724]&m[725]&m[726]&m[770]))):InitCond[1060];
    m[732] = run?((((m[728]&~m[729]&~m[730]&~m[731]&~m[775])|(~m[728]&m[729]&~m[730]&~m[731]&~m[775])|(~m[728]&~m[729]&m[730]&~m[731]&~m[775])|(m[728]&m[729]&~m[730]&m[731]&~m[775])|(m[728]&~m[729]&m[730]&m[731]&~m[775])|(~m[728]&m[729]&m[730]&m[731]&~m[775]))&BiasedRNG[567])|(((m[728]&~m[729]&~m[730]&~m[731]&m[775])|(~m[728]&m[729]&~m[730]&~m[731]&m[775])|(~m[728]&~m[729]&m[730]&~m[731]&m[775])|(m[728]&m[729]&~m[730]&m[731]&m[775])|(m[728]&~m[729]&m[730]&m[731]&m[775])|(~m[728]&m[729]&m[730]&m[731]&m[775]))&~BiasedRNG[567])|((m[728]&m[729]&~m[730]&~m[731]&~m[775])|(m[728]&~m[729]&m[730]&~m[731]&~m[775])|(~m[728]&m[729]&m[730]&~m[731]&~m[775])|(m[728]&m[729]&m[730]&~m[731]&~m[775])|(m[728]&m[729]&m[730]&m[731]&~m[775])|(m[728]&m[729]&~m[730]&~m[731]&m[775])|(m[728]&~m[729]&m[730]&~m[731]&m[775])|(~m[728]&m[729]&m[730]&~m[731]&m[775])|(m[728]&m[729]&m[730]&~m[731]&m[775])|(m[728]&m[729]&m[730]&m[731]&m[775]))):InitCond[1061];
    m[737] = run?((((m[733]&~m[734]&~m[735]&~m[736]&~m[780])|(~m[733]&m[734]&~m[735]&~m[736]&~m[780])|(~m[733]&~m[734]&m[735]&~m[736]&~m[780])|(m[733]&m[734]&~m[735]&m[736]&~m[780])|(m[733]&~m[734]&m[735]&m[736]&~m[780])|(~m[733]&m[734]&m[735]&m[736]&~m[780]))&BiasedRNG[568])|(((m[733]&~m[734]&~m[735]&~m[736]&m[780])|(~m[733]&m[734]&~m[735]&~m[736]&m[780])|(~m[733]&~m[734]&m[735]&~m[736]&m[780])|(m[733]&m[734]&~m[735]&m[736]&m[780])|(m[733]&~m[734]&m[735]&m[736]&m[780])|(~m[733]&m[734]&m[735]&m[736]&m[780]))&~BiasedRNG[568])|((m[733]&m[734]&~m[735]&~m[736]&~m[780])|(m[733]&~m[734]&m[735]&~m[736]&~m[780])|(~m[733]&m[734]&m[735]&~m[736]&~m[780])|(m[733]&m[734]&m[735]&~m[736]&~m[780])|(m[733]&m[734]&m[735]&m[736]&~m[780])|(m[733]&m[734]&~m[735]&~m[736]&m[780])|(m[733]&~m[734]&m[735]&~m[736]&m[780])|(~m[733]&m[734]&m[735]&~m[736]&m[780])|(m[733]&m[734]&m[735]&~m[736]&m[780])|(m[733]&m[734]&m[735]&m[736]&m[780]))):InitCond[1062];
    m[742] = run?((((m[738]&~m[739]&~m[740]&~m[741]&~m[785])|(~m[738]&m[739]&~m[740]&~m[741]&~m[785])|(~m[738]&~m[739]&m[740]&~m[741]&~m[785])|(m[738]&m[739]&~m[740]&m[741]&~m[785])|(m[738]&~m[739]&m[740]&m[741]&~m[785])|(~m[738]&m[739]&m[740]&m[741]&~m[785]))&BiasedRNG[569])|(((m[738]&~m[739]&~m[740]&~m[741]&m[785])|(~m[738]&m[739]&~m[740]&~m[741]&m[785])|(~m[738]&~m[739]&m[740]&~m[741]&m[785])|(m[738]&m[739]&~m[740]&m[741]&m[785])|(m[738]&~m[739]&m[740]&m[741]&m[785])|(~m[738]&m[739]&m[740]&m[741]&m[785]))&~BiasedRNG[569])|((m[738]&m[739]&~m[740]&~m[741]&~m[785])|(m[738]&~m[739]&m[740]&~m[741]&~m[785])|(~m[738]&m[739]&m[740]&~m[741]&~m[785])|(m[738]&m[739]&m[740]&~m[741]&~m[785])|(m[738]&m[739]&m[740]&m[741]&~m[785])|(m[738]&m[739]&~m[740]&~m[741]&m[785])|(m[738]&~m[739]&m[740]&~m[741]&m[785])|(~m[738]&m[739]&m[740]&~m[741]&m[785])|(m[738]&m[739]&m[740]&~m[741]&m[785])|(m[738]&m[739]&m[740]&m[741]&m[785]))):InitCond[1063];
    m[747] = run?((((m[743]&~m[744]&~m[745]&~m[746]&~m[790])|(~m[743]&m[744]&~m[745]&~m[746]&~m[790])|(~m[743]&~m[744]&m[745]&~m[746]&~m[790])|(m[743]&m[744]&~m[745]&m[746]&~m[790])|(m[743]&~m[744]&m[745]&m[746]&~m[790])|(~m[743]&m[744]&m[745]&m[746]&~m[790]))&BiasedRNG[570])|(((m[743]&~m[744]&~m[745]&~m[746]&m[790])|(~m[743]&m[744]&~m[745]&~m[746]&m[790])|(~m[743]&~m[744]&m[745]&~m[746]&m[790])|(m[743]&m[744]&~m[745]&m[746]&m[790])|(m[743]&~m[744]&m[745]&m[746]&m[790])|(~m[743]&m[744]&m[745]&m[746]&m[790]))&~BiasedRNG[570])|((m[743]&m[744]&~m[745]&~m[746]&~m[790])|(m[743]&~m[744]&m[745]&~m[746]&~m[790])|(~m[743]&m[744]&m[745]&~m[746]&~m[790])|(m[743]&m[744]&m[745]&~m[746]&~m[790])|(m[743]&m[744]&m[745]&m[746]&~m[790])|(m[743]&m[744]&~m[745]&~m[746]&m[790])|(m[743]&~m[744]&m[745]&~m[746]&m[790])|(~m[743]&m[744]&m[745]&~m[746]&m[790])|(m[743]&m[744]&m[745]&~m[746]&m[790])|(m[743]&m[744]&m[745]&m[746]&m[790]))):InitCond[1064];
    m[752] = run?((((m[748]&~m[749]&~m[750]&~m[751]&~m[795])|(~m[748]&m[749]&~m[750]&~m[751]&~m[795])|(~m[748]&~m[749]&m[750]&~m[751]&~m[795])|(m[748]&m[749]&~m[750]&m[751]&~m[795])|(m[748]&~m[749]&m[750]&m[751]&~m[795])|(~m[748]&m[749]&m[750]&m[751]&~m[795]))&BiasedRNG[571])|(((m[748]&~m[749]&~m[750]&~m[751]&m[795])|(~m[748]&m[749]&~m[750]&~m[751]&m[795])|(~m[748]&~m[749]&m[750]&~m[751]&m[795])|(m[748]&m[749]&~m[750]&m[751]&m[795])|(m[748]&~m[749]&m[750]&m[751]&m[795])|(~m[748]&m[749]&m[750]&m[751]&m[795]))&~BiasedRNG[571])|((m[748]&m[749]&~m[750]&~m[751]&~m[795])|(m[748]&~m[749]&m[750]&~m[751]&~m[795])|(~m[748]&m[749]&m[750]&~m[751]&~m[795])|(m[748]&m[749]&m[750]&~m[751]&~m[795])|(m[748]&m[749]&m[750]&m[751]&~m[795])|(m[748]&m[749]&~m[750]&~m[751]&m[795])|(m[748]&~m[749]&m[750]&~m[751]&m[795])|(~m[748]&m[749]&m[750]&~m[751]&m[795])|(m[748]&m[749]&m[750]&~m[751]&m[795])|(m[748]&m[749]&m[750]&m[751]&m[795]))):InitCond[1065];
    m[757] = run?((((m[753]&~m[754]&~m[755]&~m[756]&~m[805])|(~m[753]&m[754]&~m[755]&~m[756]&~m[805])|(~m[753]&~m[754]&m[755]&~m[756]&~m[805])|(m[753]&m[754]&~m[755]&m[756]&~m[805])|(m[753]&~m[754]&m[755]&m[756]&~m[805])|(~m[753]&m[754]&m[755]&m[756]&~m[805]))&BiasedRNG[572])|(((m[753]&~m[754]&~m[755]&~m[756]&m[805])|(~m[753]&m[754]&~m[755]&~m[756]&m[805])|(~m[753]&~m[754]&m[755]&~m[756]&m[805])|(m[753]&m[754]&~m[755]&m[756]&m[805])|(m[753]&~m[754]&m[755]&m[756]&m[805])|(~m[753]&m[754]&m[755]&m[756]&m[805]))&~BiasedRNG[572])|((m[753]&m[754]&~m[755]&~m[756]&~m[805])|(m[753]&~m[754]&m[755]&~m[756]&~m[805])|(~m[753]&m[754]&m[755]&~m[756]&~m[805])|(m[753]&m[754]&m[755]&~m[756]&~m[805])|(m[753]&m[754]&m[755]&m[756]&~m[805])|(m[753]&m[754]&~m[755]&~m[756]&m[805])|(m[753]&~m[754]&m[755]&~m[756]&m[805])|(~m[753]&m[754]&m[755]&~m[756]&m[805])|(m[753]&m[754]&m[755]&~m[756]&m[805])|(m[753]&m[754]&m[755]&m[756]&m[805]))):InitCond[1066];
    m[762] = run?((((m[758]&~m[759]&~m[760]&~m[761]&~m[810])|(~m[758]&m[759]&~m[760]&~m[761]&~m[810])|(~m[758]&~m[759]&m[760]&~m[761]&~m[810])|(m[758]&m[759]&~m[760]&m[761]&~m[810])|(m[758]&~m[759]&m[760]&m[761]&~m[810])|(~m[758]&m[759]&m[760]&m[761]&~m[810]))&BiasedRNG[573])|(((m[758]&~m[759]&~m[760]&~m[761]&m[810])|(~m[758]&m[759]&~m[760]&~m[761]&m[810])|(~m[758]&~m[759]&m[760]&~m[761]&m[810])|(m[758]&m[759]&~m[760]&m[761]&m[810])|(m[758]&~m[759]&m[760]&m[761]&m[810])|(~m[758]&m[759]&m[760]&m[761]&m[810]))&~BiasedRNG[573])|((m[758]&m[759]&~m[760]&~m[761]&~m[810])|(m[758]&~m[759]&m[760]&~m[761]&~m[810])|(~m[758]&m[759]&m[760]&~m[761]&~m[810])|(m[758]&m[759]&m[760]&~m[761]&~m[810])|(m[758]&m[759]&m[760]&m[761]&~m[810])|(m[758]&m[759]&~m[760]&~m[761]&m[810])|(m[758]&~m[759]&m[760]&~m[761]&m[810])|(~m[758]&m[759]&m[760]&~m[761]&m[810])|(m[758]&m[759]&m[760]&~m[761]&m[810])|(m[758]&m[759]&m[760]&m[761]&m[810]))):InitCond[1067];
    m[767] = run?((((m[763]&~m[764]&~m[765]&~m[766]&~m[815])|(~m[763]&m[764]&~m[765]&~m[766]&~m[815])|(~m[763]&~m[764]&m[765]&~m[766]&~m[815])|(m[763]&m[764]&~m[765]&m[766]&~m[815])|(m[763]&~m[764]&m[765]&m[766]&~m[815])|(~m[763]&m[764]&m[765]&m[766]&~m[815]))&BiasedRNG[574])|(((m[763]&~m[764]&~m[765]&~m[766]&m[815])|(~m[763]&m[764]&~m[765]&~m[766]&m[815])|(~m[763]&~m[764]&m[765]&~m[766]&m[815])|(m[763]&m[764]&~m[765]&m[766]&m[815])|(m[763]&~m[764]&m[765]&m[766]&m[815])|(~m[763]&m[764]&m[765]&m[766]&m[815]))&~BiasedRNG[574])|((m[763]&m[764]&~m[765]&~m[766]&~m[815])|(m[763]&~m[764]&m[765]&~m[766]&~m[815])|(~m[763]&m[764]&m[765]&~m[766]&~m[815])|(m[763]&m[764]&m[765]&~m[766]&~m[815])|(m[763]&m[764]&m[765]&m[766]&~m[815])|(m[763]&m[764]&~m[765]&~m[766]&m[815])|(m[763]&~m[764]&m[765]&~m[766]&m[815])|(~m[763]&m[764]&m[765]&~m[766]&m[815])|(m[763]&m[764]&m[765]&~m[766]&m[815])|(m[763]&m[764]&m[765]&m[766]&m[815]))):InitCond[1068];
    m[772] = run?((((m[768]&~m[769]&~m[770]&~m[771]&~m[820])|(~m[768]&m[769]&~m[770]&~m[771]&~m[820])|(~m[768]&~m[769]&m[770]&~m[771]&~m[820])|(m[768]&m[769]&~m[770]&m[771]&~m[820])|(m[768]&~m[769]&m[770]&m[771]&~m[820])|(~m[768]&m[769]&m[770]&m[771]&~m[820]))&BiasedRNG[575])|(((m[768]&~m[769]&~m[770]&~m[771]&m[820])|(~m[768]&m[769]&~m[770]&~m[771]&m[820])|(~m[768]&~m[769]&m[770]&~m[771]&m[820])|(m[768]&m[769]&~m[770]&m[771]&m[820])|(m[768]&~m[769]&m[770]&m[771]&m[820])|(~m[768]&m[769]&m[770]&m[771]&m[820]))&~BiasedRNG[575])|((m[768]&m[769]&~m[770]&~m[771]&~m[820])|(m[768]&~m[769]&m[770]&~m[771]&~m[820])|(~m[768]&m[769]&m[770]&~m[771]&~m[820])|(m[768]&m[769]&m[770]&~m[771]&~m[820])|(m[768]&m[769]&m[770]&m[771]&~m[820])|(m[768]&m[769]&~m[770]&~m[771]&m[820])|(m[768]&~m[769]&m[770]&~m[771]&m[820])|(~m[768]&m[769]&m[770]&~m[771]&m[820])|(m[768]&m[769]&m[770]&~m[771]&m[820])|(m[768]&m[769]&m[770]&m[771]&m[820]))):InitCond[1069];
    m[777] = run?((((m[773]&~m[774]&~m[775]&~m[776]&~m[825])|(~m[773]&m[774]&~m[775]&~m[776]&~m[825])|(~m[773]&~m[774]&m[775]&~m[776]&~m[825])|(m[773]&m[774]&~m[775]&m[776]&~m[825])|(m[773]&~m[774]&m[775]&m[776]&~m[825])|(~m[773]&m[774]&m[775]&m[776]&~m[825]))&BiasedRNG[576])|(((m[773]&~m[774]&~m[775]&~m[776]&m[825])|(~m[773]&m[774]&~m[775]&~m[776]&m[825])|(~m[773]&~m[774]&m[775]&~m[776]&m[825])|(m[773]&m[774]&~m[775]&m[776]&m[825])|(m[773]&~m[774]&m[775]&m[776]&m[825])|(~m[773]&m[774]&m[775]&m[776]&m[825]))&~BiasedRNG[576])|((m[773]&m[774]&~m[775]&~m[776]&~m[825])|(m[773]&~m[774]&m[775]&~m[776]&~m[825])|(~m[773]&m[774]&m[775]&~m[776]&~m[825])|(m[773]&m[774]&m[775]&~m[776]&~m[825])|(m[773]&m[774]&m[775]&m[776]&~m[825])|(m[773]&m[774]&~m[775]&~m[776]&m[825])|(m[773]&~m[774]&m[775]&~m[776]&m[825])|(~m[773]&m[774]&m[775]&~m[776]&m[825])|(m[773]&m[774]&m[775]&~m[776]&m[825])|(m[773]&m[774]&m[775]&m[776]&m[825]))):InitCond[1070];
    m[782] = run?((((m[778]&~m[779]&~m[780]&~m[781]&~m[830])|(~m[778]&m[779]&~m[780]&~m[781]&~m[830])|(~m[778]&~m[779]&m[780]&~m[781]&~m[830])|(m[778]&m[779]&~m[780]&m[781]&~m[830])|(m[778]&~m[779]&m[780]&m[781]&~m[830])|(~m[778]&m[779]&m[780]&m[781]&~m[830]))&BiasedRNG[577])|(((m[778]&~m[779]&~m[780]&~m[781]&m[830])|(~m[778]&m[779]&~m[780]&~m[781]&m[830])|(~m[778]&~m[779]&m[780]&~m[781]&m[830])|(m[778]&m[779]&~m[780]&m[781]&m[830])|(m[778]&~m[779]&m[780]&m[781]&m[830])|(~m[778]&m[779]&m[780]&m[781]&m[830]))&~BiasedRNG[577])|((m[778]&m[779]&~m[780]&~m[781]&~m[830])|(m[778]&~m[779]&m[780]&~m[781]&~m[830])|(~m[778]&m[779]&m[780]&~m[781]&~m[830])|(m[778]&m[779]&m[780]&~m[781]&~m[830])|(m[778]&m[779]&m[780]&m[781]&~m[830])|(m[778]&m[779]&~m[780]&~m[781]&m[830])|(m[778]&~m[779]&m[780]&~m[781]&m[830])|(~m[778]&m[779]&m[780]&~m[781]&m[830])|(m[778]&m[779]&m[780]&~m[781]&m[830])|(m[778]&m[779]&m[780]&m[781]&m[830]))):InitCond[1071];
    m[787] = run?((((m[783]&~m[784]&~m[785]&~m[786]&~m[835])|(~m[783]&m[784]&~m[785]&~m[786]&~m[835])|(~m[783]&~m[784]&m[785]&~m[786]&~m[835])|(m[783]&m[784]&~m[785]&m[786]&~m[835])|(m[783]&~m[784]&m[785]&m[786]&~m[835])|(~m[783]&m[784]&m[785]&m[786]&~m[835]))&BiasedRNG[578])|(((m[783]&~m[784]&~m[785]&~m[786]&m[835])|(~m[783]&m[784]&~m[785]&~m[786]&m[835])|(~m[783]&~m[784]&m[785]&~m[786]&m[835])|(m[783]&m[784]&~m[785]&m[786]&m[835])|(m[783]&~m[784]&m[785]&m[786]&m[835])|(~m[783]&m[784]&m[785]&m[786]&m[835]))&~BiasedRNG[578])|((m[783]&m[784]&~m[785]&~m[786]&~m[835])|(m[783]&~m[784]&m[785]&~m[786]&~m[835])|(~m[783]&m[784]&m[785]&~m[786]&~m[835])|(m[783]&m[784]&m[785]&~m[786]&~m[835])|(m[783]&m[784]&m[785]&m[786]&~m[835])|(m[783]&m[784]&~m[785]&~m[786]&m[835])|(m[783]&~m[784]&m[785]&~m[786]&m[835])|(~m[783]&m[784]&m[785]&~m[786]&m[835])|(m[783]&m[784]&m[785]&~m[786]&m[835])|(m[783]&m[784]&m[785]&m[786]&m[835]))):InitCond[1072];
    m[792] = run?((((m[788]&~m[789]&~m[790]&~m[791]&~m[840])|(~m[788]&m[789]&~m[790]&~m[791]&~m[840])|(~m[788]&~m[789]&m[790]&~m[791]&~m[840])|(m[788]&m[789]&~m[790]&m[791]&~m[840])|(m[788]&~m[789]&m[790]&m[791]&~m[840])|(~m[788]&m[789]&m[790]&m[791]&~m[840]))&BiasedRNG[579])|(((m[788]&~m[789]&~m[790]&~m[791]&m[840])|(~m[788]&m[789]&~m[790]&~m[791]&m[840])|(~m[788]&~m[789]&m[790]&~m[791]&m[840])|(m[788]&m[789]&~m[790]&m[791]&m[840])|(m[788]&~m[789]&m[790]&m[791]&m[840])|(~m[788]&m[789]&m[790]&m[791]&m[840]))&~BiasedRNG[579])|((m[788]&m[789]&~m[790]&~m[791]&~m[840])|(m[788]&~m[789]&m[790]&~m[791]&~m[840])|(~m[788]&m[789]&m[790]&~m[791]&~m[840])|(m[788]&m[789]&m[790]&~m[791]&~m[840])|(m[788]&m[789]&m[790]&m[791]&~m[840])|(m[788]&m[789]&~m[790]&~m[791]&m[840])|(m[788]&~m[789]&m[790]&~m[791]&m[840])|(~m[788]&m[789]&m[790]&~m[791]&m[840])|(m[788]&m[789]&m[790]&~m[791]&m[840])|(m[788]&m[789]&m[790]&m[791]&m[840]))):InitCond[1073];
    m[797] = run?((((m[793]&~m[794]&~m[795]&~m[796]&~m[845])|(~m[793]&m[794]&~m[795]&~m[796]&~m[845])|(~m[793]&~m[794]&m[795]&~m[796]&~m[845])|(m[793]&m[794]&~m[795]&m[796]&~m[845])|(m[793]&~m[794]&m[795]&m[796]&~m[845])|(~m[793]&m[794]&m[795]&m[796]&~m[845]))&BiasedRNG[580])|(((m[793]&~m[794]&~m[795]&~m[796]&m[845])|(~m[793]&m[794]&~m[795]&~m[796]&m[845])|(~m[793]&~m[794]&m[795]&~m[796]&m[845])|(m[793]&m[794]&~m[795]&m[796]&m[845])|(m[793]&~m[794]&m[795]&m[796]&m[845])|(~m[793]&m[794]&m[795]&m[796]&m[845]))&~BiasedRNG[580])|((m[793]&m[794]&~m[795]&~m[796]&~m[845])|(m[793]&~m[794]&m[795]&~m[796]&~m[845])|(~m[793]&m[794]&m[795]&~m[796]&~m[845])|(m[793]&m[794]&m[795]&~m[796]&~m[845])|(m[793]&m[794]&m[795]&m[796]&~m[845])|(m[793]&m[794]&~m[795]&~m[796]&m[845])|(m[793]&~m[794]&m[795]&~m[796]&m[845])|(~m[793]&m[794]&m[795]&~m[796]&m[845])|(m[793]&m[794]&m[795]&~m[796]&m[845])|(m[793]&m[794]&m[795]&m[796]&m[845]))):InitCond[1074];
    m[802] = run?((((m[798]&~m[799]&~m[800]&~m[801]&~m[850])|(~m[798]&m[799]&~m[800]&~m[801]&~m[850])|(~m[798]&~m[799]&m[800]&~m[801]&~m[850])|(m[798]&m[799]&~m[800]&m[801]&~m[850])|(m[798]&~m[799]&m[800]&m[801]&~m[850])|(~m[798]&m[799]&m[800]&m[801]&~m[850]))&BiasedRNG[581])|(((m[798]&~m[799]&~m[800]&~m[801]&m[850])|(~m[798]&m[799]&~m[800]&~m[801]&m[850])|(~m[798]&~m[799]&m[800]&~m[801]&m[850])|(m[798]&m[799]&~m[800]&m[801]&m[850])|(m[798]&~m[799]&m[800]&m[801]&m[850])|(~m[798]&m[799]&m[800]&m[801]&m[850]))&~BiasedRNG[581])|((m[798]&m[799]&~m[800]&~m[801]&~m[850])|(m[798]&~m[799]&m[800]&~m[801]&~m[850])|(~m[798]&m[799]&m[800]&~m[801]&~m[850])|(m[798]&m[799]&m[800]&~m[801]&~m[850])|(m[798]&m[799]&m[800]&m[801]&~m[850])|(m[798]&m[799]&~m[800]&~m[801]&m[850])|(m[798]&~m[799]&m[800]&~m[801]&m[850])|(~m[798]&m[799]&m[800]&~m[801]&m[850])|(m[798]&m[799]&m[800]&~m[801]&m[850])|(m[798]&m[799]&m[800]&m[801]&m[850]))):InitCond[1075];
    m[807] = run?((((m[803]&~m[804]&~m[805]&~m[806]&~m[860])|(~m[803]&m[804]&~m[805]&~m[806]&~m[860])|(~m[803]&~m[804]&m[805]&~m[806]&~m[860])|(m[803]&m[804]&~m[805]&m[806]&~m[860])|(m[803]&~m[804]&m[805]&m[806]&~m[860])|(~m[803]&m[804]&m[805]&m[806]&~m[860]))&BiasedRNG[582])|(((m[803]&~m[804]&~m[805]&~m[806]&m[860])|(~m[803]&m[804]&~m[805]&~m[806]&m[860])|(~m[803]&~m[804]&m[805]&~m[806]&m[860])|(m[803]&m[804]&~m[805]&m[806]&m[860])|(m[803]&~m[804]&m[805]&m[806]&m[860])|(~m[803]&m[804]&m[805]&m[806]&m[860]))&~BiasedRNG[582])|((m[803]&m[804]&~m[805]&~m[806]&~m[860])|(m[803]&~m[804]&m[805]&~m[806]&~m[860])|(~m[803]&m[804]&m[805]&~m[806]&~m[860])|(m[803]&m[804]&m[805]&~m[806]&~m[860])|(m[803]&m[804]&m[805]&m[806]&~m[860])|(m[803]&m[804]&~m[805]&~m[806]&m[860])|(m[803]&~m[804]&m[805]&~m[806]&m[860])|(~m[803]&m[804]&m[805]&~m[806]&m[860])|(m[803]&m[804]&m[805]&~m[806]&m[860])|(m[803]&m[804]&m[805]&m[806]&m[860]))):InitCond[1076];
    m[812] = run?((((m[808]&~m[809]&~m[810]&~m[811]&~m[865])|(~m[808]&m[809]&~m[810]&~m[811]&~m[865])|(~m[808]&~m[809]&m[810]&~m[811]&~m[865])|(m[808]&m[809]&~m[810]&m[811]&~m[865])|(m[808]&~m[809]&m[810]&m[811]&~m[865])|(~m[808]&m[809]&m[810]&m[811]&~m[865]))&BiasedRNG[583])|(((m[808]&~m[809]&~m[810]&~m[811]&m[865])|(~m[808]&m[809]&~m[810]&~m[811]&m[865])|(~m[808]&~m[809]&m[810]&~m[811]&m[865])|(m[808]&m[809]&~m[810]&m[811]&m[865])|(m[808]&~m[809]&m[810]&m[811]&m[865])|(~m[808]&m[809]&m[810]&m[811]&m[865]))&~BiasedRNG[583])|((m[808]&m[809]&~m[810]&~m[811]&~m[865])|(m[808]&~m[809]&m[810]&~m[811]&~m[865])|(~m[808]&m[809]&m[810]&~m[811]&~m[865])|(m[808]&m[809]&m[810]&~m[811]&~m[865])|(m[808]&m[809]&m[810]&m[811]&~m[865])|(m[808]&m[809]&~m[810]&~m[811]&m[865])|(m[808]&~m[809]&m[810]&~m[811]&m[865])|(~m[808]&m[809]&m[810]&~m[811]&m[865])|(m[808]&m[809]&m[810]&~m[811]&m[865])|(m[808]&m[809]&m[810]&m[811]&m[865]))):InitCond[1077];
    m[817] = run?((((m[813]&~m[814]&~m[815]&~m[816]&~m[870])|(~m[813]&m[814]&~m[815]&~m[816]&~m[870])|(~m[813]&~m[814]&m[815]&~m[816]&~m[870])|(m[813]&m[814]&~m[815]&m[816]&~m[870])|(m[813]&~m[814]&m[815]&m[816]&~m[870])|(~m[813]&m[814]&m[815]&m[816]&~m[870]))&BiasedRNG[584])|(((m[813]&~m[814]&~m[815]&~m[816]&m[870])|(~m[813]&m[814]&~m[815]&~m[816]&m[870])|(~m[813]&~m[814]&m[815]&~m[816]&m[870])|(m[813]&m[814]&~m[815]&m[816]&m[870])|(m[813]&~m[814]&m[815]&m[816]&m[870])|(~m[813]&m[814]&m[815]&m[816]&m[870]))&~BiasedRNG[584])|((m[813]&m[814]&~m[815]&~m[816]&~m[870])|(m[813]&~m[814]&m[815]&~m[816]&~m[870])|(~m[813]&m[814]&m[815]&~m[816]&~m[870])|(m[813]&m[814]&m[815]&~m[816]&~m[870])|(m[813]&m[814]&m[815]&m[816]&~m[870])|(m[813]&m[814]&~m[815]&~m[816]&m[870])|(m[813]&~m[814]&m[815]&~m[816]&m[870])|(~m[813]&m[814]&m[815]&~m[816]&m[870])|(m[813]&m[814]&m[815]&~m[816]&m[870])|(m[813]&m[814]&m[815]&m[816]&m[870]))):InitCond[1078];
    m[822] = run?((((m[818]&~m[819]&~m[820]&~m[821]&~m[875])|(~m[818]&m[819]&~m[820]&~m[821]&~m[875])|(~m[818]&~m[819]&m[820]&~m[821]&~m[875])|(m[818]&m[819]&~m[820]&m[821]&~m[875])|(m[818]&~m[819]&m[820]&m[821]&~m[875])|(~m[818]&m[819]&m[820]&m[821]&~m[875]))&BiasedRNG[585])|(((m[818]&~m[819]&~m[820]&~m[821]&m[875])|(~m[818]&m[819]&~m[820]&~m[821]&m[875])|(~m[818]&~m[819]&m[820]&~m[821]&m[875])|(m[818]&m[819]&~m[820]&m[821]&m[875])|(m[818]&~m[819]&m[820]&m[821]&m[875])|(~m[818]&m[819]&m[820]&m[821]&m[875]))&~BiasedRNG[585])|((m[818]&m[819]&~m[820]&~m[821]&~m[875])|(m[818]&~m[819]&m[820]&~m[821]&~m[875])|(~m[818]&m[819]&m[820]&~m[821]&~m[875])|(m[818]&m[819]&m[820]&~m[821]&~m[875])|(m[818]&m[819]&m[820]&m[821]&~m[875])|(m[818]&m[819]&~m[820]&~m[821]&m[875])|(m[818]&~m[819]&m[820]&~m[821]&m[875])|(~m[818]&m[819]&m[820]&~m[821]&m[875])|(m[818]&m[819]&m[820]&~m[821]&m[875])|(m[818]&m[819]&m[820]&m[821]&m[875]))):InitCond[1079];
    m[827] = run?((((m[823]&~m[824]&~m[825]&~m[826]&~m[880])|(~m[823]&m[824]&~m[825]&~m[826]&~m[880])|(~m[823]&~m[824]&m[825]&~m[826]&~m[880])|(m[823]&m[824]&~m[825]&m[826]&~m[880])|(m[823]&~m[824]&m[825]&m[826]&~m[880])|(~m[823]&m[824]&m[825]&m[826]&~m[880]))&BiasedRNG[586])|(((m[823]&~m[824]&~m[825]&~m[826]&m[880])|(~m[823]&m[824]&~m[825]&~m[826]&m[880])|(~m[823]&~m[824]&m[825]&~m[826]&m[880])|(m[823]&m[824]&~m[825]&m[826]&m[880])|(m[823]&~m[824]&m[825]&m[826]&m[880])|(~m[823]&m[824]&m[825]&m[826]&m[880]))&~BiasedRNG[586])|((m[823]&m[824]&~m[825]&~m[826]&~m[880])|(m[823]&~m[824]&m[825]&~m[826]&~m[880])|(~m[823]&m[824]&m[825]&~m[826]&~m[880])|(m[823]&m[824]&m[825]&~m[826]&~m[880])|(m[823]&m[824]&m[825]&m[826]&~m[880])|(m[823]&m[824]&~m[825]&~m[826]&m[880])|(m[823]&~m[824]&m[825]&~m[826]&m[880])|(~m[823]&m[824]&m[825]&~m[826]&m[880])|(m[823]&m[824]&m[825]&~m[826]&m[880])|(m[823]&m[824]&m[825]&m[826]&m[880]))):InitCond[1080];
    m[832] = run?((((m[828]&~m[829]&~m[830]&~m[831]&~m[885])|(~m[828]&m[829]&~m[830]&~m[831]&~m[885])|(~m[828]&~m[829]&m[830]&~m[831]&~m[885])|(m[828]&m[829]&~m[830]&m[831]&~m[885])|(m[828]&~m[829]&m[830]&m[831]&~m[885])|(~m[828]&m[829]&m[830]&m[831]&~m[885]))&BiasedRNG[587])|(((m[828]&~m[829]&~m[830]&~m[831]&m[885])|(~m[828]&m[829]&~m[830]&~m[831]&m[885])|(~m[828]&~m[829]&m[830]&~m[831]&m[885])|(m[828]&m[829]&~m[830]&m[831]&m[885])|(m[828]&~m[829]&m[830]&m[831]&m[885])|(~m[828]&m[829]&m[830]&m[831]&m[885]))&~BiasedRNG[587])|((m[828]&m[829]&~m[830]&~m[831]&~m[885])|(m[828]&~m[829]&m[830]&~m[831]&~m[885])|(~m[828]&m[829]&m[830]&~m[831]&~m[885])|(m[828]&m[829]&m[830]&~m[831]&~m[885])|(m[828]&m[829]&m[830]&m[831]&~m[885])|(m[828]&m[829]&~m[830]&~m[831]&m[885])|(m[828]&~m[829]&m[830]&~m[831]&m[885])|(~m[828]&m[829]&m[830]&~m[831]&m[885])|(m[828]&m[829]&m[830]&~m[831]&m[885])|(m[828]&m[829]&m[830]&m[831]&m[885]))):InitCond[1081];
    m[837] = run?((((m[833]&~m[834]&~m[835]&~m[836]&~m[890])|(~m[833]&m[834]&~m[835]&~m[836]&~m[890])|(~m[833]&~m[834]&m[835]&~m[836]&~m[890])|(m[833]&m[834]&~m[835]&m[836]&~m[890])|(m[833]&~m[834]&m[835]&m[836]&~m[890])|(~m[833]&m[834]&m[835]&m[836]&~m[890]))&BiasedRNG[588])|(((m[833]&~m[834]&~m[835]&~m[836]&m[890])|(~m[833]&m[834]&~m[835]&~m[836]&m[890])|(~m[833]&~m[834]&m[835]&~m[836]&m[890])|(m[833]&m[834]&~m[835]&m[836]&m[890])|(m[833]&~m[834]&m[835]&m[836]&m[890])|(~m[833]&m[834]&m[835]&m[836]&m[890]))&~BiasedRNG[588])|((m[833]&m[834]&~m[835]&~m[836]&~m[890])|(m[833]&~m[834]&m[835]&~m[836]&~m[890])|(~m[833]&m[834]&m[835]&~m[836]&~m[890])|(m[833]&m[834]&m[835]&~m[836]&~m[890])|(m[833]&m[834]&m[835]&m[836]&~m[890])|(m[833]&m[834]&~m[835]&~m[836]&m[890])|(m[833]&~m[834]&m[835]&~m[836]&m[890])|(~m[833]&m[834]&m[835]&~m[836]&m[890])|(m[833]&m[834]&m[835]&~m[836]&m[890])|(m[833]&m[834]&m[835]&m[836]&m[890]))):InitCond[1082];
    m[842] = run?((((m[838]&~m[839]&~m[840]&~m[841]&~m[895])|(~m[838]&m[839]&~m[840]&~m[841]&~m[895])|(~m[838]&~m[839]&m[840]&~m[841]&~m[895])|(m[838]&m[839]&~m[840]&m[841]&~m[895])|(m[838]&~m[839]&m[840]&m[841]&~m[895])|(~m[838]&m[839]&m[840]&m[841]&~m[895]))&BiasedRNG[589])|(((m[838]&~m[839]&~m[840]&~m[841]&m[895])|(~m[838]&m[839]&~m[840]&~m[841]&m[895])|(~m[838]&~m[839]&m[840]&~m[841]&m[895])|(m[838]&m[839]&~m[840]&m[841]&m[895])|(m[838]&~m[839]&m[840]&m[841]&m[895])|(~m[838]&m[839]&m[840]&m[841]&m[895]))&~BiasedRNG[589])|((m[838]&m[839]&~m[840]&~m[841]&~m[895])|(m[838]&~m[839]&m[840]&~m[841]&~m[895])|(~m[838]&m[839]&m[840]&~m[841]&~m[895])|(m[838]&m[839]&m[840]&~m[841]&~m[895])|(m[838]&m[839]&m[840]&m[841]&~m[895])|(m[838]&m[839]&~m[840]&~m[841]&m[895])|(m[838]&~m[839]&m[840]&~m[841]&m[895])|(~m[838]&m[839]&m[840]&~m[841]&m[895])|(m[838]&m[839]&m[840]&~m[841]&m[895])|(m[838]&m[839]&m[840]&m[841]&m[895]))):InitCond[1083];
    m[847] = run?((((m[843]&~m[844]&~m[845]&~m[846]&~m[900])|(~m[843]&m[844]&~m[845]&~m[846]&~m[900])|(~m[843]&~m[844]&m[845]&~m[846]&~m[900])|(m[843]&m[844]&~m[845]&m[846]&~m[900])|(m[843]&~m[844]&m[845]&m[846]&~m[900])|(~m[843]&m[844]&m[845]&m[846]&~m[900]))&BiasedRNG[590])|(((m[843]&~m[844]&~m[845]&~m[846]&m[900])|(~m[843]&m[844]&~m[845]&~m[846]&m[900])|(~m[843]&~m[844]&m[845]&~m[846]&m[900])|(m[843]&m[844]&~m[845]&m[846]&m[900])|(m[843]&~m[844]&m[845]&m[846]&m[900])|(~m[843]&m[844]&m[845]&m[846]&m[900]))&~BiasedRNG[590])|((m[843]&m[844]&~m[845]&~m[846]&~m[900])|(m[843]&~m[844]&m[845]&~m[846]&~m[900])|(~m[843]&m[844]&m[845]&~m[846]&~m[900])|(m[843]&m[844]&m[845]&~m[846]&~m[900])|(m[843]&m[844]&m[845]&m[846]&~m[900])|(m[843]&m[844]&~m[845]&~m[846]&m[900])|(m[843]&~m[844]&m[845]&~m[846]&m[900])|(~m[843]&m[844]&m[845]&~m[846]&m[900])|(m[843]&m[844]&m[845]&~m[846]&m[900])|(m[843]&m[844]&m[845]&m[846]&m[900]))):InitCond[1084];
    m[852] = run?((((m[848]&~m[849]&~m[850]&~m[851]&~m[905])|(~m[848]&m[849]&~m[850]&~m[851]&~m[905])|(~m[848]&~m[849]&m[850]&~m[851]&~m[905])|(m[848]&m[849]&~m[850]&m[851]&~m[905])|(m[848]&~m[849]&m[850]&m[851]&~m[905])|(~m[848]&m[849]&m[850]&m[851]&~m[905]))&BiasedRNG[591])|(((m[848]&~m[849]&~m[850]&~m[851]&m[905])|(~m[848]&m[849]&~m[850]&~m[851]&m[905])|(~m[848]&~m[849]&m[850]&~m[851]&m[905])|(m[848]&m[849]&~m[850]&m[851]&m[905])|(m[848]&~m[849]&m[850]&m[851]&m[905])|(~m[848]&m[849]&m[850]&m[851]&m[905]))&~BiasedRNG[591])|((m[848]&m[849]&~m[850]&~m[851]&~m[905])|(m[848]&~m[849]&m[850]&~m[851]&~m[905])|(~m[848]&m[849]&m[850]&~m[851]&~m[905])|(m[848]&m[849]&m[850]&~m[851]&~m[905])|(m[848]&m[849]&m[850]&m[851]&~m[905])|(m[848]&m[849]&~m[850]&~m[851]&m[905])|(m[848]&~m[849]&m[850]&~m[851]&m[905])|(~m[848]&m[849]&m[850]&~m[851]&m[905])|(m[848]&m[849]&m[850]&~m[851]&m[905])|(m[848]&m[849]&m[850]&m[851]&m[905]))):InitCond[1085];
    m[857] = run?((((m[853]&~m[854]&~m[855]&~m[856]&~m[910])|(~m[853]&m[854]&~m[855]&~m[856]&~m[910])|(~m[853]&~m[854]&m[855]&~m[856]&~m[910])|(m[853]&m[854]&~m[855]&m[856]&~m[910])|(m[853]&~m[854]&m[855]&m[856]&~m[910])|(~m[853]&m[854]&m[855]&m[856]&~m[910]))&BiasedRNG[592])|(((m[853]&~m[854]&~m[855]&~m[856]&m[910])|(~m[853]&m[854]&~m[855]&~m[856]&m[910])|(~m[853]&~m[854]&m[855]&~m[856]&m[910])|(m[853]&m[854]&~m[855]&m[856]&m[910])|(m[853]&~m[854]&m[855]&m[856]&m[910])|(~m[853]&m[854]&m[855]&m[856]&m[910]))&~BiasedRNG[592])|((m[853]&m[854]&~m[855]&~m[856]&~m[910])|(m[853]&~m[854]&m[855]&~m[856]&~m[910])|(~m[853]&m[854]&m[855]&~m[856]&~m[910])|(m[853]&m[854]&m[855]&~m[856]&~m[910])|(m[853]&m[854]&m[855]&m[856]&~m[910])|(m[853]&m[854]&~m[855]&~m[856]&m[910])|(m[853]&~m[854]&m[855]&~m[856]&m[910])|(~m[853]&m[854]&m[855]&~m[856]&m[910])|(m[853]&m[854]&m[855]&~m[856]&m[910])|(m[853]&m[854]&m[855]&m[856]&m[910]))):InitCond[1086];
    m[862] = run?((((m[858]&~m[859]&~m[860]&~m[861]&~m[913])|(~m[858]&m[859]&~m[860]&~m[861]&~m[913])|(~m[858]&~m[859]&m[860]&~m[861]&~m[913])|(m[858]&m[859]&~m[860]&m[861]&~m[913])|(m[858]&~m[859]&m[860]&m[861]&~m[913])|(~m[858]&m[859]&m[860]&m[861]&~m[913]))&BiasedRNG[593])|(((m[858]&~m[859]&~m[860]&~m[861]&m[913])|(~m[858]&m[859]&~m[860]&~m[861]&m[913])|(~m[858]&~m[859]&m[860]&~m[861]&m[913])|(m[858]&m[859]&~m[860]&m[861]&m[913])|(m[858]&~m[859]&m[860]&m[861]&m[913])|(~m[858]&m[859]&m[860]&m[861]&m[913]))&~BiasedRNG[593])|((m[858]&m[859]&~m[860]&~m[861]&~m[913])|(m[858]&~m[859]&m[860]&~m[861]&~m[913])|(~m[858]&m[859]&m[860]&~m[861]&~m[913])|(m[858]&m[859]&m[860]&~m[861]&~m[913])|(m[858]&m[859]&m[860]&m[861]&~m[913])|(m[858]&m[859]&~m[860]&~m[861]&m[913])|(m[858]&~m[859]&m[860]&~m[861]&m[913])|(~m[858]&m[859]&m[860]&~m[861]&m[913])|(m[858]&m[859]&m[860]&~m[861]&m[913])|(m[858]&m[859]&m[860]&m[861]&m[913]))):InitCond[1087];
    m[867] = run?((((m[863]&~m[864]&~m[865]&~m[866]&~m[915])|(~m[863]&m[864]&~m[865]&~m[866]&~m[915])|(~m[863]&~m[864]&m[865]&~m[866]&~m[915])|(m[863]&m[864]&~m[865]&m[866]&~m[915])|(m[863]&~m[864]&m[865]&m[866]&~m[915])|(~m[863]&m[864]&m[865]&m[866]&~m[915]))&BiasedRNG[594])|(((m[863]&~m[864]&~m[865]&~m[866]&m[915])|(~m[863]&m[864]&~m[865]&~m[866]&m[915])|(~m[863]&~m[864]&m[865]&~m[866]&m[915])|(m[863]&m[864]&~m[865]&m[866]&m[915])|(m[863]&~m[864]&m[865]&m[866]&m[915])|(~m[863]&m[864]&m[865]&m[866]&m[915]))&~BiasedRNG[594])|((m[863]&m[864]&~m[865]&~m[866]&~m[915])|(m[863]&~m[864]&m[865]&~m[866]&~m[915])|(~m[863]&m[864]&m[865]&~m[866]&~m[915])|(m[863]&m[864]&m[865]&~m[866]&~m[915])|(m[863]&m[864]&m[865]&m[866]&~m[915])|(m[863]&m[864]&~m[865]&~m[866]&m[915])|(m[863]&~m[864]&m[865]&~m[866]&m[915])|(~m[863]&m[864]&m[865]&~m[866]&m[915])|(m[863]&m[864]&m[865]&~m[866]&m[915])|(m[863]&m[864]&m[865]&m[866]&m[915]))):InitCond[1088];
    m[872] = run?((((m[868]&~m[869]&~m[870]&~m[871]&~m[920])|(~m[868]&m[869]&~m[870]&~m[871]&~m[920])|(~m[868]&~m[869]&m[870]&~m[871]&~m[920])|(m[868]&m[869]&~m[870]&m[871]&~m[920])|(m[868]&~m[869]&m[870]&m[871]&~m[920])|(~m[868]&m[869]&m[870]&m[871]&~m[920]))&BiasedRNG[595])|(((m[868]&~m[869]&~m[870]&~m[871]&m[920])|(~m[868]&m[869]&~m[870]&~m[871]&m[920])|(~m[868]&~m[869]&m[870]&~m[871]&m[920])|(m[868]&m[869]&~m[870]&m[871]&m[920])|(m[868]&~m[869]&m[870]&m[871]&m[920])|(~m[868]&m[869]&m[870]&m[871]&m[920]))&~BiasedRNG[595])|((m[868]&m[869]&~m[870]&~m[871]&~m[920])|(m[868]&~m[869]&m[870]&~m[871]&~m[920])|(~m[868]&m[869]&m[870]&~m[871]&~m[920])|(m[868]&m[869]&m[870]&~m[871]&~m[920])|(m[868]&m[869]&m[870]&m[871]&~m[920])|(m[868]&m[869]&~m[870]&~m[871]&m[920])|(m[868]&~m[869]&m[870]&~m[871]&m[920])|(~m[868]&m[869]&m[870]&~m[871]&m[920])|(m[868]&m[869]&m[870]&~m[871]&m[920])|(m[868]&m[869]&m[870]&m[871]&m[920]))):InitCond[1089];
    m[877] = run?((((m[873]&~m[874]&~m[875]&~m[876]&~m[925])|(~m[873]&m[874]&~m[875]&~m[876]&~m[925])|(~m[873]&~m[874]&m[875]&~m[876]&~m[925])|(m[873]&m[874]&~m[875]&m[876]&~m[925])|(m[873]&~m[874]&m[875]&m[876]&~m[925])|(~m[873]&m[874]&m[875]&m[876]&~m[925]))&BiasedRNG[596])|(((m[873]&~m[874]&~m[875]&~m[876]&m[925])|(~m[873]&m[874]&~m[875]&~m[876]&m[925])|(~m[873]&~m[874]&m[875]&~m[876]&m[925])|(m[873]&m[874]&~m[875]&m[876]&m[925])|(m[873]&~m[874]&m[875]&m[876]&m[925])|(~m[873]&m[874]&m[875]&m[876]&m[925]))&~BiasedRNG[596])|((m[873]&m[874]&~m[875]&~m[876]&~m[925])|(m[873]&~m[874]&m[875]&~m[876]&~m[925])|(~m[873]&m[874]&m[875]&~m[876]&~m[925])|(m[873]&m[874]&m[875]&~m[876]&~m[925])|(m[873]&m[874]&m[875]&m[876]&~m[925])|(m[873]&m[874]&~m[875]&~m[876]&m[925])|(m[873]&~m[874]&m[875]&~m[876]&m[925])|(~m[873]&m[874]&m[875]&~m[876]&m[925])|(m[873]&m[874]&m[875]&~m[876]&m[925])|(m[873]&m[874]&m[875]&m[876]&m[925]))):InitCond[1090];
    m[882] = run?((((m[878]&~m[879]&~m[880]&~m[881]&~m[930])|(~m[878]&m[879]&~m[880]&~m[881]&~m[930])|(~m[878]&~m[879]&m[880]&~m[881]&~m[930])|(m[878]&m[879]&~m[880]&m[881]&~m[930])|(m[878]&~m[879]&m[880]&m[881]&~m[930])|(~m[878]&m[879]&m[880]&m[881]&~m[930]))&BiasedRNG[597])|(((m[878]&~m[879]&~m[880]&~m[881]&m[930])|(~m[878]&m[879]&~m[880]&~m[881]&m[930])|(~m[878]&~m[879]&m[880]&~m[881]&m[930])|(m[878]&m[879]&~m[880]&m[881]&m[930])|(m[878]&~m[879]&m[880]&m[881]&m[930])|(~m[878]&m[879]&m[880]&m[881]&m[930]))&~BiasedRNG[597])|((m[878]&m[879]&~m[880]&~m[881]&~m[930])|(m[878]&~m[879]&m[880]&~m[881]&~m[930])|(~m[878]&m[879]&m[880]&~m[881]&~m[930])|(m[878]&m[879]&m[880]&~m[881]&~m[930])|(m[878]&m[879]&m[880]&m[881]&~m[930])|(m[878]&m[879]&~m[880]&~m[881]&m[930])|(m[878]&~m[879]&m[880]&~m[881]&m[930])|(~m[878]&m[879]&m[880]&~m[881]&m[930])|(m[878]&m[879]&m[880]&~m[881]&m[930])|(m[878]&m[879]&m[880]&m[881]&m[930]))):InitCond[1091];
    m[887] = run?((((m[883]&~m[884]&~m[885]&~m[886]&~m[935])|(~m[883]&m[884]&~m[885]&~m[886]&~m[935])|(~m[883]&~m[884]&m[885]&~m[886]&~m[935])|(m[883]&m[884]&~m[885]&m[886]&~m[935])|(m[883]&~m[884]&m[885]&m[886]&~m[935])|(~m[883]&m[884]&m[885]&m[886]&~m[935]))&BiasedRNG[598])|(((m[883]&~m[884]&~m[885]&~m[886]&m[935])|(~m[883]&m[884]&~m[885]&~m[886]&m[935])|(~m[883]&~m[884]&m[885]&~m[886]&m[935])|(m[883]&m[884]&~m[885]&m[886]&m[935])|(m[883]&~m[884]&m[885]&m[886]&m[935])|(~m[883]&m[884]&m[885]&m[886]&m[935]))&~BiasedRNG[598])|((m[883]&m[884]&~m[885]&~m[886]&~m[935])|(m[883]&~m[884]&m[885]&~m[886]&~m[935])|(~m[883]&m[884]&m[885]&~m[886]&~m[935])|(m[883]&m[884]&m[885]&~m[886]&~m[935])|(m[883]&m[884]&m[885]&m[886]&~m[935])|(m[883]&m[884]&~m[885]&~m[886]&m[935])|(m[883]&~m[884]&m[885]&~m[886]&m[935])|(~m[883]&m[884]&m[885]&~m[886]&m[935])|(m[883]&m[884]&m[885]&~m[886]&m[935])|(m[883]&m[884]&m[885]&m[886]&m[935]))):InitCond[1092];
    m[892] = run?((((m[888]&~m[889]&~m[890]&~m[891]&~m[940])|(~m[888]&m[889]&~m[890]&~m[891]&~m[940])|(~m[888]&~m[889]&m[890]&~m[891]&~m[940])|(m[888]&m[889]&~m[890]&m[891]&~m[940])|(m[888]&~m[889]&m[890]&m[891]&~m[940])|(~m[888]&m[889]&m[890]&m[891]&~m[940]))&BiasedRNG[599])|(((m[888]&~m[889]&~m[890]&~m[891]&m[940])|(~m[888]&m[889]&~m[890]&~m[891]&m[940])|(~m[888]&~m[889]&m[890]&~m[891]&m[940])|(m[888]&m[889]&~m[890]&m[891]&m[940])|(m[888]&~m[889]&m[890]&m[891]&m[940])|(~m[888]&m[889]&m[890]&m[891]&m[940]))&~BiasedRNG[599])|((m[888]&m[889]&~m[890]&~m[891]&~m[940])|(m[888]&~m[889]&m[890]&~m[891]&~m[940])|(~m[888]&m[889]&m[890]&~m[891]&~m[940])|(m[888]&m[889]&m[890]&~m[891]&~m[940])|(m[888]&m[889]&m[890]&m[891]&~m[940])|(m[888]&m[889]&~m[890]&~m[891]&m[940])|(m[888]&~m[889]&m[890]&~m[891]&m[940])|(~m[888]&m[889]&m[890]&~m[891]&m[940])|(m[888]&m[889]&m[890]&~m[891]&m[940])|(m[888]&m[889]&m[890]&m[891]&m[940]))):InitCond[1093];
    m[897] = run?((((m[893]&~m[894]&~m[895]&~m[896]&~m[945])|(~m[893]&m[894]&~m[895]&~m[896]&~m[945])|(~m[893]&~m[894]&m[895]&~m[896]&~m[945])|(m[893]&m[894]&~m[895]&m[896]&~m[945])|(m[893]&~m[894]&m[895]&m[896]&~m[945])|(~m[893]&m[894]&m[895]&m[896]&~m[945]))&BiasedRNG[600])|(((m[893]&~m[894]&~m[895]&~m[896]&m[945])|(~m[893]&m[894]&~m[895]&~m[896]&m[945])|(~m[893]&~m[894]&m[895]&~m[896]&m[945])|(m[893]&m[894]&~m[895]&m[896]&m[945])|(m[893]&~m[894]&m[895]&m[896]&m[945])|(~m[893]&m[894]&m[895]&m[896]&m[945]))&~BiasedRNG[600])|((m[893]&m[894]&~m[895]&~m[896]&~m[945])|(m[893]&~m[894]&m[895]&~m[896]&~m[945])|(~m[893]&m[894]&m[895]&~m[896]&~m[945])|(m[893]&m[894]&m[895]&~m[896]&~m[945])|(m[893]&m[894]&m[895]&m[896]&~m[945])|(m[893]&m[894]&~m[895]&~m[896]&m[945])|(m[893]&~m[894]&m[895]&~m[896]&m[945])|(~m[893]&m[894]&m[895]&~m[896]&m[945])|(m[893]&m[894]&m[895]&~m[896]&m[945])|(m[893]&m[894]&m[895]&m[896]&m[945]))):InitCond[1094];
    m[902] = run?((((m[898]&~m[899]&~m[900]&~m[901]&~m[950])|(~m[898]&m[899]&~m[900]&~m[901]&~m[950])|(~m[898]&~m[899]&m[900]&~m[901]&~m[950])|(m[898]&m[899]&~m[900]&m[901]&~m[950])|(m[898]&~m[899]&m[900]&m[901]&~m[950])|(~m[898]&m[899]&m[900]&m[901]&~m[950]))&BiasedRNG[601])|(((m[898]&~m[899]&~m[900]&~m[901]&m[950])|(~m[898]&m[899]&~m[900]&~m[901]&m[950])|(~m[898]&~m[899]&m[900]&~m[901]&m[950])|(m[898]&m[899]&~m[900]&m[901]&m[950])|(m[898]&~m[899]&m[900]&m[901]&m[950])|(~m[898]&m[899]&m[900]&m[901]&m[950]))&~BiasedRNG[601])|((m[898]&m[899]&~m[900]&~m[901]&~m[950])|(m[898]&~m[899]&m[900]&~m[901]&~m[950])|(~m[898]&m[899]&m[900]&~m[901]&~m[950])|(m[898]&m[899]&m[900]&~m[901]&~m[950])|(m[898]&m[899]&m[900]&m[901]&~m[950])|(m[898]&m[899]&~m[900]&~m[901]&m[950])|(m[898]&~m[899]&m[900]&~m[901]&m[950])|(~m[898]&m[899]&m[900]&~m[901]&m[950])|(m[898]&m[899]&m[900]&~m[901]&m[950])|(m[898]&m[899]&m[900]&m[901]&m[950]))):InitCond[1095];
    m[907] = run?((((m[903]&~m[904]&~m[905]&~m[906]&~m[955])|(~m[903]&m[904]&~m[905]&~m[906]&~m[955])|(~m[903]&~m[904]&m[905]&~m[906]&~m[955])|(m[903]&m[904]&~m[905]&m[906]&~m[955])|(m[903]&~m[904]&m[905]&m[906]&~m[955])|(~m[903]&m[904]&m[905]&m[906]&~m[955]))&BiasedRNG[602])|(((m[903]&~m[904]&~m[905]&~m[906]&m[955])|(~m[903]&m[904]&~m[905]&~m[906]&m[955])|(~m[903]&~m[904]&m[905]&~m[906]&m[955])|(m[903]&m[904]&~m[905]&m[906]&m[955])|(m[903]&~m[904]&m[905]&m[906]&m[955])|(~m[903]&m[904]&m[905]&m[906]&m[955]))&~BiasedRNG[602])|((m[903]&m[904]&~m[905]&~m[906]&~m[955])|(m[903]&~m[904]&m[905]&~m[906]&~m[955])|(~m[903]&m[904]&m[905]&~m[906]&~m[955])|(m[903]&m[904]&m[905]&~m[906]&~m[955])|(m[903]&m[904]&m[905]&m[906]&~m[955])|(m[903]&m[904]&~m[905]&~m[906]&m[955])|(m[903]&~m[904]&m[905]&~m[906]&m[955])|(~m[903]&m[904]&m[905]&~m[906]&m[955])|(m[903]&m[904]&m[905]&~m[906]&m[955])|(m[903]&m[904]&m[905]&m[906]&m[955]))):InitCond[1096];
    m[912] = run?((((m[908]&~m[909]&~m[910]&~m[911]&~m[960])|(~m[908]&m[909]&~m[910]&~m[911]&~m[960])|(~m[908]&~m[909]&m[910]&~m[911]&~m[960])|(m[908]&m[909]&~m[910]&m[911]&~m[960])|(m[908]&~m[909]&m[910]&m[911]&~m[960])|(~m[908]&m[909]&m[910]&m[911]&~m[960]))&BiasedRNG[603])|(((m[908]&~m[909]&~m[910]&~m[911]&m[960])|(~m[908]&m[909]&~m[910]&~m[911]&m[960])|(~m[908]&~m[909]&m[910]&~m[911]&m[960])|(m[908]&m[909]&~m[910]&m[911]&m[960])|(m[908]&~m[909]&m[910]&m[911]&m[960])|(~m[908]&m[909]&m[910]&m[911]&m[960]))&~BiasedRNG[603])|((m[908]&m[909]&~m[910]&~m[911]&~m[960])|(m[908]&~m[909]&m[910]&~m[911]&~m[960])|(~m[908]&m[909]&m[910]&~m[911]&~m[960])|(m[908]&m[909]&m[910]&~m[911]&~m[960])|(m[908]&m[909]&m[910]&m[911]&~m[960])|(m[908]&m[909]&~m[910]&~m[911]&m[960])|(m[908]&~m[909]&m[910]&~m[911]&m[960])|(~m[908]&m[909]&m[910]&~m[911]&m[960])|(m[908]&m[909]&m[910]&~m[911]&m[960])|(m[908]&m[909]&m[910]&m[911]&m[960]))):InitCond[1097];
    m[917] = run?((((m[913]&~m[914]&~m[915]&~m[916]&~m[963])|(~m[913]&m[914]&~m[915]&~m[916]&~m[963])|(~m[913]&~m[914]&m[915]&~m[916]&~m[963])|(m[913]&m[914]&~m[915]&m[916]&~m[963])|(m[913]&~m[914]&m[915]&m[916]&~m[963])|(~m[913]&m[914]&m[915]&m[916]&~m[963]))&BiasedRNG[604])|(((m[913]&~m[914]&~m[915]&~m[916]&m[963])|(~m[913]&m[914]&~m[915]&~m[916]&m[963])|(~m[913]&~m[914]&m[915]&~m[916]&m[963])|(m[913]&m[914]&~m[915]&m[916]&m[963])|(m[913]&~m[914]&m[915]&m[916]&m[963])|(~m[913]&m[914]&m[915]&m[916]&m[963]))&~BiasedRNG[604])|((m[913]&m[914]&~m[915]&~m[916]&~m[963])|(m[913]&~m[914]&m[915]&~m[916]&~m[963])|(~m[913]&m[914]&m[915]&~m[916]&~m[963])|(m[913]&m[914]&m[915]&~m[916]&~m[963])|(m[913]&m[914]&m[915]&m[916]&~m[963])|(m[913]&m[914]&~m[915]&~m[916]&m[963])|(m[913]&~m[914]&m[915]&~m[916]&m[963])|(~m[913]&m[914]&m[915]&~m[916]&m[963])|(m[913]&m[914]&m[915]&~m[916]&m[963])|(m[913]&m[914]&m[915]&m[916]&m[963]))):InitCond[1098];
    m[922] = run?((((m[918]&~m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&~m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&~m[920]&m[921]&~m[965])|(m[918]&~m[919]&m[920]&m[921]&~m[965])|(~m[918]&m[919]&m[920]&m[921]&~m[965]))&BiasedRNG[605])|(((m[918]&~m[919]&~m[920]&~m[921]&m[965])|(~m[918]&m[919]&~m[920]&~m[921]&m[965])|(~m[918]&~m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&~m[920]&m[921]&m[965])|(m[918]&~m[919]&m[920]&m[921]&m[965])|(~m[918]&m[919]&m[920]&m[921]&m[965]))&~BiasedRNG[605])|((m[918]&m[919]&~m[920]&~m[921]&~m[965])|(m[918]&~m[919]&m[920]&~m[921]&~m[965])|(~m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&m[921]&~m[965])|(m[918]&m[919]&~m[920]&~m[921]&m[965])|(m[918]&~m[919]&m[920]&~m[921]&m[965])|(~m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&m[921]&m[965]))):InitCond[1099];
    m[927] = run?((((m[923]&~m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&~m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&~m[925]&m[926]&~m[970])|(m[923]&~m[924]&m[925]&m[926]&~m[970])|(~m[923]&m[924]&m[925]&m[926]&~m[970]))&BiasedRNG[606])|(((m[923]&~m[924]&~m[925]&~m[926]&m[970])|(~m[923]&m[924]&~m[925]&~m[926]&m[970])|(~m[923]&~m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&~m[925]&m[926]&m[970])|(m[923]&~m[924]&m[925]&m[926]&m[970])|(~m[923]&m[924]&m[925]&m[926]&m[970]))&~BiasedRNG[606])|((m[923]&m[924]&~m[925]&~m[926]&~m[970])|(m[923]&~m[924]&m[925]&~m[926]&~m[970])|(~m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&m[926]&~m[970])|(m[923]&m[924]&~m[925]&~m[926]&m[970])|(m[923]&~m[924]&m[925]&~m[926]&m[970])|(~m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&m[926]&m[970]))):InitCond[1100];
    m[932] = run?((((m[928]&~m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&~m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&~m[930]&m[931]&~m[975])|(m[928]&~m[929]&m[930]&m[931]&~m[975])|(~m[928]&m[929]&m[930]&m[931]&~m[975]))&BiasedRNG[607])|(((m[928]&~m[929]&~m[930]&~m[931]&m[975])|(~m[928]&m[929]&~m[930]&~m[931]&m[975])|(~m[928]&~m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&~m[930]&m[931]&m[975])|(m[928]&~m[929]&m[930]&m[931]&m[975])|(~m[928]&m[929]&m[930]&m[931]&m[975]))&~BiasedRNG[607])|((m[928]&m[929]&~m[930]&~m[931]&~m[975])|(m[928]&~m[929]&m[930]&~m[931]&~m[975])|(~m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&m[931]&~m[975])|(m[928]&m[929]&~m[930]&~m[931]&m[975])|(m[928]&~m[929]&m[930]&~m[931]&m[975])|(~m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&m[931]&m[975]))):InitCond[1101];
    m[937] = run?((((m[933]&~m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&~m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&~m[935]&m[936]&~m[980])|(m[933]&~m[934]&m[935]&m[936]&~m[980])|(~m[933]&m[934]&m[935]&m[936]&~m[980]))&BiasedRNG[608])|(((m[933]&~m[934]&~m[935]&~m[936]&m[980])|(~m[933]&m[934]&~m[935]&~m[936]&m[980])|(~m[933]&~m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&~m[935]&m[936]&m[980])|(m[933]&~m[934]&m[935]&m[936]&m[980])|(~m[933]&m[934]&m[935]&m[936]&m[980]))&~BiasedRNG[608])|((m[933]&m[934]&~m[935]&~m[936]&~m[980])|(m[933]&~m[934]&m[935]&~m[936]&~m[980])|(~m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&m[936]&~m[980])|(m[933]&m[934]&~m[935]&~m[936]&m[980])|(m[933]&~m[934]&m[935]&~m[936]&m[980])|(~m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&m[936]&m[980]))):InitCond[1102];
    m[942] = run?((((m[938]&~m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&~m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&~m[940]&m[941]&~m[985])|(m[938]&~m[939]&m[940]&m[941]&~m[985])|(~m[938]&m[939]&m[940]&m[941]&~m[985]))&BiasedRNG[609])|(((m[938]&~m[939]&~m[940]&~m[941]&m[985])|(~m[938]&m[939]&~m[940]&~m[941]&m[985])|(~m[938]&~m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&~m[940]&m[941]&m[985])|(m[938]&~m[939]&m[940]&m[941]&m[985])|(~m[938]&m[939]&m[940]&m[941]&m[985]))&~BiasedRNG[609])|((m[938]&m[939]&~m[940]&~m[941]&~m[985])|(m[938]&~m[939]&m[940]&~m[941]&~m[985])|(~m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&m[941]&~m[985])|(m[938]&m[939]&~m[940]&~m[941]&m[985])|(m[938]&~m[939]&m[940]&~m[941]&m[985])|(~m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&m[941]&m[985]))):InitCond[1103];
    m[947] = run?((((m[943]&~m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&~m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&~m[945]&m[946]&~m[990])|(m[943]&~m[944]&m[945]&m[946]&~m[990])|(~m[943]&m[944]&m[945]&m[946]&~m[990]))&BiasedRNG[610])|(((m[943]&~m[944]&~m[945]&~m[946]&m[990])|(~m[943]&m[944]&~m[945]&~m[946]&m[990])|(~m[943]&~m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&~m[945]&m[946]&m[990])|(m[943]&~m[944]&m[945]&m[946]&m[990])|(~m[943]&m[944]&m[945]&m[946]&m[990]))&~BiasedRNG[610])|((m[943]&m[944]&~m[945]&~m[946]&~m[990])|(m[943]&~m[944]&m[945]&~m[946]&~m[990])|(~m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&m[946]&~m[990])|(m[943]&m[944]&~m[945]&~m[946]&m[990])|(m[943]&~m[944]&m[945]&~m[946]&m[990])|(~m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&m[946]&m[990]))):InitCond[1104];
    m[952] = run?((((m[948]&~m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&~m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&~m[950]&m[951]&~m[995])|(m[948]&~m[949]&m[950]&m[951]&~m[995])|(~m[948]&m[949]&m[950]&m[951]&~m[995]))&BiasedRNG[611])|(((m[948]&~m[949]&~m[950]&~m[951]&m[995])|(~m[948]&m[949]&~m[950]&~m[951]&m[995])|(~m[948]&~m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&~m[950]&m[951]&m[995])|(m[948]&~m[949]&m[950]&m[951]&m[995])|(~m[948]&m[949]&m[950]&m[951]&m[995]))&~BiasedRNG[611])|((m[948]&m[949]&~m[950]&~m[951]&~m[995])|(m[948]&~m[949]&m[950]&~m[951]&~m[995])|(~m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&m[951]&~m[995])|(m[948]&m[949]&~m[950]&~m[951]&m[995])|(m[948]&~m[949]&m[950]&~m[951]&m[995])|(~m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&m[951]&m[995]))):InitCond[1105];
    m[957] = run?((((m[953]&~m[954]&~m[955]&~m[956]&~m[1000])|(~m[953]&m[954]&~m[955]&~m[956]&~m[1000])|(~m[953]&~m[954]&m[955]&~m[956]&~m[1000])|(m[953]&m[954]&~m[955]&m[956]&~m[1000])|(m[953]&~m[954]&m[955]&m[956]&~m[1000])|(~m[953]&m[954]&m[955]&m[956]&~m[1000]))&BiasedRNG[612])|(((m[953]&~m[954]&~m[955]&~m[956]&m[1000])|(~m[953]&m[954]&~m[955]&~m[956]&m[1000])|(~m[953]&~m[954]&m[955]&~m[956]&m[1000])|(m[953]&m[954]&~m[955]&m[956]&m[1000])|(m[953]&~m[954]&m[955]&m[956]&m[1000])|(~m[953]&m[954]&m[955]&m[956]&m[1000]))&~BiasedRNG[612])|((m[953]&m[954]&~m[955]&~m[956]&~m[1000])|(m[953]&~m[954]&m[955]&~m[956]&~m[1000])|(~m[953]&m[954]&m[955]&~m[956]&~m[1000])|(m[953]&m[954]&m[955]&~m[956]&~m[1000])|(m[953]&m[954]&m[955]&m[956]&~m[1000])|(m[953]&m[954]&~m[955]&~m[956]&m[1000])|(m[953]&~m[954]&m[955]&~m[956]&m[1000])|(~m[953]&m[954]&m[955]&~m[956]&m[1000])|(m[953]&m[954]&m[955]&~m[956]&m[1000])|(m[953]&m[954]&m[955]&m[956]&m[1000]))):InitCond[1106];
    m[962] = run?((((m[958]&~m[959]&~m[960]&~m[961]&~m[1005])|(~m[958]&m[959]&~m[960]&~m[961]&~m[1005])|(~m[958]&~m[959]&m[960]&~m[961]&~m[1005])|(m[958]&m[959]&~m[960]&m[961]&~m[1005])|(m[958]&~m[959]&m[960]&m[961]&~m[1005])|(~m[958]&m[959]&m[960]&m[961]&~m[1005]))&BiasedRNG[613])|(((m[958]&~m[959]&~m[960]&~m[961]&m[1005])|(~m[958]&m[959]&~m[960]&~m[961]&m[1005])|(~m[958]&~m[959]&m[960]&~m[961]&m[1005])|(m[958]&m[959]&~m[960]&m[961]&m[1005])|(m[958]&~m[959]&m[960]&m[961]&m[1005])|(~m[958]&m[959]&m[960]&m[961]&m[1005]))&~BiasedRNG[613])|((m[958]&m[959]&~m[960]&~m[961]&~m[1005])|(m[958]&~m[959]&m[960]&~m[961]&~m[1005])|(~m[958]&m[959]&m[960]&~m[961]&~m[1005])|(m[958]&m[959]&m[960]&~m[961]&~m[1005])|(m[958]&m[959]&m[960]&m[961]&~m[1005])|(m[958]&m[959]&~m[960]&~m[961]&m[1005])|(m[958]&~m[959]&m[960]&~m[961]&m[1005])|(~m[958]&m[959]&m[960]&~m[961]&m[1005])|(m[958]&m[959]&m[960]&~m[961]&m[1005])|(m[958]&m[959]&m[960]&m[961]&m[1005]))):InitCond[1107];
    m[967] = run?((((m[963]&~m[964]&~m[965]&~m[966]&~m[1008])|(~m[963]&m[964]&~m[965]&~m[966]&~m[1008])|(~m[963]&~m[964]&m[965]&~m[966]&~m[1008])|(m[963]&m[964]&~m[965]&m[966]&~m[1008])|(m[963]&~m[964]&m[965]&m[966]&~m[1008])|(~m[963]&m[964]&m[965]&m[966]&~m[1008]))&BiasedRNG[614])|(((m[963]&~m[964]&~m[965]&~m[966]&m[1008])|(~m[963]&m[964]&~m[965]&~m[966]&m[1008])|(~m[963]&~m[964]&m[965]&~m[966]&m[1008])|(m[963]&m[964]&~m[965]&m[966]&m[1008])|(m[963]&~m[964]&m[965]&m[966]&m[1008])|(~m[963]&m[964]&m[965]&m[966]&m[1008]))&~BiasedRNG[614])|((m[963]&m[964]&~m[965]&~m[966]&~m[1008])|(m[963]&~m[964]&m[965]&~m[966]&~m[1008])|(~m[963]&m[964]&m[965]&~m[966]&~m[1008])|(m[963]&m[964]&m[965]&~m[966]&~m[1008])|(m[963]&m[964]&m[965]&m[966]&~m[1008])|(m[963]&m[964]&~m[965]&~m[966]&m[1008])|(m[963]&~m[964]&m[965]&~m[966]&m[1008])|(~m[963]&m[964]&m[965]&~m[966]&m[1008])|(m[963]&m[964]&m[965]&~m[966]&m[1008])|(m[963]&m[964]&m[965]&m[966]&m[1008]))):InitCond[1108];
    m[972] = run?((((m[968]&~m[969]&~m[970]&~m[971]&~m[1010])|(~m[968]&m[969]&~m[970]&~m[971]&~m[1010])|(~m[968]&~m[969]&m[970]&~m[971]&~m[1010])|(m[968]&m[969]&~m[970]&m[971]&~m[1010])|(m[968]&~m[969]&m[970]&m[971]&~m[1010])|(~m[968]&m[969]&m[970]&m[971]&~m[1010]))&BiasedRNG[615])|(((m[968]&~m[969]&~m[970]&~m[971]&m[1010])|(~m[968]&m[969]&~m[970]&~m[971]&m[1010])|(~m[968]&~m[969]&m[970]&~m[971]&m[1010])|(m[968]&m[969]&~m[970]&m[971]&m[1010])|(m[968]&~m[969]&m[970]&m[971]&m[1010])|(~m[968]&m[969]&m[970]&m[971]&m[1010]))&~BiasedRNG[615])|((m[968]&m[969]&~m[970]&~m[971]&~m[1010])|(m[968]&~m[969]&m[970]&~m[971]&~m[1010])|(~m[968]&m[969]&m[970]&~m[971]&~m[1010])|(m[968]&m[969]&m[970]&~m[971]&~m[1010])|(m[968]&m[969]&m[970]&m[971]&~m[1010])|(m[968]&m[969]&~m[970]&~m[971]&m[1010])|(m[968]&~m[969]&m[970]&~m[971]&m[1010])|(~m[968]&m[969]&m[970]&~m[971]&m[1010])|(m[968]&m[969]&m[970]&~m[971]&m[1010])|(m[968]&m[969]&m[970]&m[971]&m[1010]))):InitCond[1109];
    m[977] = run?((((m[973]&~m[974]&~m[975]&~m[976]&~m[1015])|(~m[973]&m[974]&~m[975]&~m[976]&~m[1015])|(~m[973]&~m[974]&m[975]&~m[976]&~m[1015])|(m[973]&m[974]&~m[975]&m[976]&~m[1015])|(m[973]&~m[974]&m[975]&m[976]&~m[1015])|(~m[973]&m[974]&m[975]&m[976]&~m[1015]))&BiasedRNG[616])|(((m[973]&~m[974]&~m[975]&~m[976]&m[1015])|(~m[973]&m[974]&~m[975]&~m[976]&m[1015])|(~m[973]&~m[974]&m[975]&~m[976]&m[1015])|(m[973]&m[974]&~m[975]&m[976]&m[1015])|(m[973]&~m[974]&m[975]&m[976]&m[1015])|(~m[973]&m[974]&m[975]&m[976]&m[1015]))&~BiasedRNG[616])|((m[973]&m[974]&~m[975]&~m[976]&~m[1015])|(m[973]&~m[974]&m[975]&~m[976]&~m[1015])|(~m[973]&m[974]&m[975]&~m[976]&~m[1015])|(m[973]&m[974]&m[975]&~m[976]&~m[1015])|(m[973]&m[974]&m[975]&m[976]&~m[1015])|(m[973]&m[974]&~m[975]&~m[976]&m[1015])|(m[973]&~m[974]&m[975]&~m[976]&m[1015])|(~m[973]&m[974]&m[975]&~m[976]&m[1015])|(m[973]&m[974]&m[975]&~m[976]&m[1015])|(m[973]&m[974]&m[975]&m[976]&m[1015]))):InitCond[1110];
    m[982] = run?((((m[978]&~m[979]&~m[980]&~m[981]&~m[1020])|(~m[978]&m[979]&~m[980]&~m[981]&~m[1020])|(~m[978]&~m[979]&m[980]&~m[981]&~m[1020])|(m[978]&m[979]&~m[980]&m[981]&~m[1020])|(m[978]&~m[979]&m[980]&m[981]&~m[1020])|(~m[978]&m[979]&m[980]&m[981]&~m[1020]))&BiasedRNG[617])|(((m[978]&~m[979]&~m[980]&~m[981]&m[1020])|(~m[978]&m[979]&~m[980]&~m[981]&m[1020])|(~m[978]&~m[979]&m[980]&~m[981]&m[1020])|(m[978]&m[979]&~m[980]&m[981]&m[1020])|(m[978]&~m[979]&m[980]&m[981]&m[1020])|(~m[978]&m[979]&m[980]&m[981]&m[1020]))&~BiasedRNG[617])|((m[978]&m[979]&~m[980]&~m[981]&~m[1020])|(m[978]&~m[979]&m[980]&~m[981]&~m[1020])|(~m[978]&m[979]&m[980]&~m[981]&~m[1020])|(m[978]&m[979]&m[980]&~m[981]&~m[1020])|(m[978]&m[979]&m[980]&m[981]&~m[1020])|(m[978]&m[979]&~m[980]&~m[981]&m[1020])|(m[978]&~m[979]&m[980]&~m[981]&m[1020])|(~m[978]&m[979]&m[980]&~m[981]&m[1020])|(m[978]&m[979]&m[980]&~m[981]&m[1020])|(m[978]&m[979]&m[980]&m[981]&m[1020]))):InitCond[1111];
    m[987] = run?((((m[983]&~m[984]&~m[985]&~m[986]&~m[1025])|(~m[983]&m[984]&~m[985]&~m[986]&~m[1025])|(~m[983]&~m[984]&m[985]&~m[986]&~m[1025])|(m[983]&m[984]&~m[985]&m[986]&~m[1025])|(m[983]&~m[984]&m[985]&m[986]&~m[1025])|(~m[983]&m[984]&m[985]&m[986]&~m[1025]))&BiasedRNG[618])|(((m[983]&~m[984]&~m[985]&~m[986]&m[1025])|(~m[983]&m[984]&~m[985]&~m[986]&m[1025])|(~m[983]&~m[984]&m[985]&~m[986]&m[1025])|(m[983]&m[984]&~m[985]&m[986]&m[1025])|(m[983]&~m[984]&m[985]&m[986]&m[1025])|(~m[983]&m[984]&m[985]&m[986]&m[1025]))&~BiasedRNG[618])|((m[983]&m[984]&~m[985]&~m[986]&~m[1025])|(m[983]&~m[984]&m[985]&~m[986]&~m[1025])|(~m[983]&m[984]&m[985]&~m[986]&~m[1025])|(m[983]&m[984]&m[985]&~m[986]&~m[1025])|(m[983]&m[984]&m[985]&m[986]&~m[1025])|(m[983]&m[984]&~m[985]&~m[986]&m[1025])|(m[983]&~m[984]&m[985]&~m[986]&m[1025])|(~m[983]&m[984]&m[985]&~m[986]&m[1025])|(m[983]&m[984]&m[985]&~m[986]&m[1025])|(m[983]&m[984]&m[985]&m[986]&m[1025]))):InitCond[1112];
    m[992] = run?((((m[988]&~m[989]&~m[990]&~m[991]&~m[1030])|(~m[988]&m[989]&~m[990]&~m[991]&~m[1030])|(~m[988]&~m[989]&m[990]&~m[991]&~m[1030])|(m[988]&m[989]&~m[990]&m[991]&~m[1030])|(m[988]&~m[989]&m[990]&m[991]&~m[1030])|(~m[988]&m[989]&m[990]&m[991]&~m[1030]))&BiasedRNG[619])|(((m[988]&~m[989]&~m[990]&~m[991]&m[1030])|(~m[988]&m[989]&~m[990]&~m[991]&m[1030])|(~m[988]&~m[989]&m[990]&~m[991]&m[1030])|(m[988]&m[989]&~m[990]&m[991]&m[1030])|(m[988]&~m[989]&m[990]&m[991]&m[1030])|(~m[988]&m[989]&m[990]&m[991]&m[1030]))&~BiasedRNG[619])|((m[988]&m[989]&~m[990]&~m[991]&~m[1030])|(m[988]&~m[989]&m[990]&~m[991]&~m[1030])|(~m[988]&m[989]&m[990]&~m[991]&~m[1030])|(m[988]&m[989]&m[990]&~m[991]&~m[1030])|(m[988]&m[989]&m[990]&m[991]&~m[1030])|(m[988]&m[989]&~m[990]&~m[991]&m[1030])|(m[988]&~m[989]&m[990]&~m[991]&m[1030])|(~m[988]&m[989]&m[990]&~m[991]&m[1030])|(m[988]&m[989]&m[990]&~m[991]&m[1030])|(m[988]&m[989]&m[990]&m[991]&m[1030]))):InitCond[1113];
    m[997] = run?((((m[993]&~m[994]&~m[995]&~m[996]&~m[1035])|(~m[993]&m[994]&~m[995]&~m[996]&~m[1035])|(~m[993]&~m[994]&m[995]&~m[996]&~m[1035])|(m[993]&m[994]&~m[995]&m[996]&~m[1035])|(m[993]&~m[994]&m[995]&m[996]&~m[1035])|(~m[993]&m[994]&m[995]&m[996]&~m[1035]))&BiasedRNG[620])|(((m[993]&~m[994]&~m[995]&~m[996]&m[1035])|(~m[993]&m[994]&~m[995]&~m[996]&m[1035])|(~m[993]&~m[994]&m[995]&~m[996]&m[1035])|(m[993]&m[994]&~m[995]&m[996]&m[1035])|(m[993]&~m[994]&m[995]&m[996]&m[1035])|(~m[993]&m[994]&m[995]&m[996]&m[1035]))&~BiasedRNG[620])|((m[993]&m[994]&~m[995]&~m[996]&~m[1035])|(m[993]&~m[994]&m[995]&~m[996]&~m[1035])|(~m[993]&m[994]&m[995]&~m[996]&~m[1035])|(m[993]&m[994]&m[995]&~m[996]&~m[1035])|(m[993]&m[994]&m[995]&m[996]&~m[1035])|(m[993]&m[994]&~m[995]&~m[996]&m[1035])|(m[993]&~m[994]&m[995]&~m[996]&m[1035])|(~m[993]&m[994]&m[995]&~m[996]&m[1035])|(m[993]&m[994]&m[995]&~m[996]&m[1035])|(m[993]&m[994]&m[995]&m[996]&m[1035]))):InitCond[1114];
    m[1002] = run?((((m[998]&~m[999]&~m[1000]&~m[1001]&~m[1040])|(~m[998]&m[999]&~m[1000]&~m[1001]&~m[1040])|(~m[998]&~m[999]&m[1000]&~m[1001]&~m[1040])|(m[998]&m[999]&~m[1000]&m[1001]&~m[1040])|(m[998]&~m[999]&m[1000]&m[1001]&~m[1040])|(~m[998]&m[999]&m[1000]&m[1001]&~m[1040]))&BiasedRNG[621])|(((m[998]&~m[999]&~m[1000]&~m[1001]&m[1040])|(~m[998]&m[999]&~m[1000]&~m[1001]&m[1040])|(~m[998]&~m[999]&m[1000]&~m[1001]&m[1040])|(m[998]&m[999]&~m[1000]&m[1001]&m[1040])|(m[998]&~m[999]&m[1000]&m[1001]&m[1040])|(~m[998]&m[999]&m[1000]&m[1001]&m[1040]))&~BiasedRNG[621])|((m[998]&m[999]&~m[1000]&~m[1001]&~m[1040])|(m[998]&~m[999]&m[1000]&~m[1001]&~m[1040])|(~m[998]&m[999]&m[1000]&~m[1001]&~m[1040])|(m[998]&m[999]&m[1000]&~m[1001]&~m[1040])|(m[998]&m[999]&m[1000]&m[1001]&~m[1040])|(m[998]&m[999]&~m[1000]&~m[1001]&m[1040])|(m[998]&~m[999]&m[1000]&~m[1001]&m[1040])|(~m[998]&m[999]&m[1000]&~m[1001]&m[1040])|(m[998]&m[999]&m[1000]&~m[1001]&m[1040])|(m[998]&m[999]&m[1000]&m[1001]&m[1040]))):InitCond[1115];
    m[1007] = run?((((m[1003]&~m[1004]&~m[1005]&~m[1006]&~m[1045])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1045])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1045])|(m[1003]&m[1004]&~m[1005]&m[1006]&~m[1045])|(m[1003]&~m[1004]&m[1005]&m[1006]&~m[1045])|(~m[1003]&m[1004]&m[1005]&m[1006]&~m[1045]))&BiasedRNG[622])|(((m[1003]&~m[1004]&~m[1005]&~m[1006]&m[1045])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&m[1045])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&m[1045])|(m[1003]&m[1004]&~m[1005]&m[1006]&m[1045])|(m[1003]&~m[1004]&m[1005]&m[1006]&m[1045])|(~m[1003]&m[1004]&m[1005]&m[1006]&m[1045]))&~BiasedRNG[622])|((m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1045])|(m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1045])|(~m[1003]&m[1004]&m[1005]&~m[1006]&~m[1045])|(m[1003]&m[1004]&m[1005]&~m[1006]&~m[1045])|(m[1003]&m[1004]&m[1005]&m[1006]&~m[1045])|(m[1003]&m[1004]&~m[1005]&~m[1006]&m[1045])|(m[1003]&~m[1004]&m[1005]&~m[1006]&m[1045])|(~m[1003]&m[1004]&m[1005]&~m[1006]&m[1045])|(m[1003]&m[1004]&m[1005]&~m[1006]&m[1045])|(m[1003]&m[1004]&m[1005]&m[1006]&m[1045]))):InitCond[1116];
    m[1012] = run?((((m[1008]&~m[1009]&~m[1010]&~m[1011]&~m[1048])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1048])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1048])|(m[1008]&m[1009]&~m[1010]&m[1011]&~m[1048])|(m[1008]&~m[1009]&m[1010]&m[1011]&~m[1048])|(~m[1008]&m[1009]&m[1010]&m[1011]&~m[1048]))&BiasedRNG[623])|(((m[1008]&~m[1009]&~m[1010]&~m[1011]&m[1048])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&m[1048])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&m[1048])|(m[1008]&m[1009]&~m[1010]&m[1011]&m[1048])|(m[1008]&~m[1009]&m[1010]&m[1011]&m[1048])|(~m[1008]&m[1009]&m[1010]&m[1011]&m[1048]))&~BiasedRNG[623])|((m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1048])|(m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1048])|(~m[1008]&m[1009]&m[1010]&~m[1011]&~m[1048])|(m[1008]&m[1009]&m[1010]&~m[1011]&~m[1048])|(m[1008]&m[1009]&m[1010]&m[1011]&~m[1048])|(m[1008]&m[1009]&~m[1010]&~m[1011]&m[1048])|(m[1008]&~m[1009]&m[1010]&~m[1011]&m[1048])|(~m[1008]&m[1009]&m[1010]&~m[1011]&m[1048])|(m[1008]&m[1009]&m[1010]&~m[1011]&m[1048])|(m[1008]&m[1009]&m[1010]&m[1011]&m[1048]))):InitCond[1117];
    m[1017] = run?((((m[1013]&~m[1014]&~m[1015]&~m[1016]&~m[1050])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1050])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1050])|(m[1013]&m[1014]&~m[1015]&m[1016]&~m[1050])|(m[1013]&~m[1014]&m[1015]&m[1016]&~m[1050])|(~m[1013]&m[1014]&m[1015]&m[1016]&~m[1050]))&BiasedRNG[624])|(((m[1013]&~m[1014]&~m[1015]&~m[1016]&m[1050])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&m[1050])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&m[1050])|(m[1013]&m[1014]&~m[1015]&m[1016]&m[1050])|(m[1013]&~m[1014]&m[1015]&m[1016]&m[1050])|(~m[1013]&m[1014]&m[1015]&m[1016]&m[1050]))&~BiasedRNG[624])|((m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1050])|(m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1050])|(~m[1013]&m[1014]&m[1015]&~m[1016]&~m[1050])|(m[1013]&m[1014]&m[1015]&~m[1016]&~m[1050])|(m[1013]&m[1014]&m[1015]&m[1016]&~m[1050])|(m[1013]&m[1014]&~m[1015]&~m[1016]&m[1050])|(m[1013]&~m[1014]&m[1015]&~m[1016]&m[1050])|(~m[1013]&m[1014]&m[1015]&~m[1016]&m[1050])|(m[1013]&m[1014]&m[1015]&~m[1016]&m[1050])|(m[1013]&m[1014]&m[1015]&m[1016]&m[1050]))):InitCond[1118];
    m[1022] = run?((((m[1018]&~m[1019]&~m[1020]&~m[1021]&~m[1055])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1055])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1055])|(m[1018]&m[1019]&~m[1020]&m[1021]&~m[1055])|(m[1018]&~m[1019]&m[1020]&m[1021]&~m[1055])|(~m[1018]&m[1019]&m[1020]&m[1021]&~m[1055]))&BiasedRNG[625])|(((m[1018]&~m[1019]&~m[1020]&~m[1021]&m[1055])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&m[1055])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&m[1055])|(m[1018]&m[1019]&~m[1020]&m[1021]&m[1055])|(m[1018]&~m[1019]&m[1020]&m[1021]&m[1055])|(~m[1018]&m[1019]&m[1020]&m[1021]&m[1055]))&~BiasedRNG[625])|((m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1055])|(m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1055])|(~m[1018]&m[1019]&m[1020]&~m[1021]&~m[1055])|(m[1018]&m[1019]&m[1020]&~m[1021]&~m[1055])|(m[1018]&m[1019]&m[1020]&m[1021]&~m[1055])|(m[1018]&m[1019]&~m[1020]&~m[1021]&m[1055])|(m[1018]&~m[1019]&m[1020]&~m[1021]&m[1055])|(~m[1018]&m[1019]&m[1020]&~m[1021]&m[1055])|(m[1018]&m[1019]&m[1020]&~m[1021]&m[1055])|(m[1018]&m[1019]&m[1020]&m[1021]&m[1055]))):InitCond[1119];
    m[1027] = run?((((m[1023]&~m[1024]&~m[1025]&~m[1026]&~m[1060])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1060])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1060])|(m[1023]&m[1024]&~m[1025]&m[1026]&~m[1060])|(m[1023]&~m[1024]&m[1025]&m[1026]&~m[1060])|(~m[1023]&m[1024]&m[1025]&m[1026]&~m[1060]))&BiasedRNG[626])|(((m[1023]&~m[1024]&~m[1025]&~m[1026]&m[1060])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&m[1060])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&m[1060])|(m[1023]&m[1024]&~m[1025]&m[1026]&m[1060])|(m[1023]&~m[1024]&m[1025]&m[1026]&m[1060])|(~m[1023]&m[1024]&m[1025]&m[1026]&m[1060]))&~BiasedRNG[626])|((m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1060])|(m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1060])|(~m[1023]&m[1024]&m[1025]&~m[1026]&~m[1060])|(m[1023]&m[1024]&m[1025]&~m[1026]&~m[1060])|(m[1023]&m[1024]&m[1025]&m[1026]&~m[1060])|(m[1023]&m[1024]&~m[1025]&~m[1026]&m[1060])|(m[1023]&~m[1024]&m[1025]&~m[1026]&m[1060])|(~m[1023]&m[1024]&m[1025]&~m[1026]&m[1060])|(m[1023]&m[1024]&m[1025]&~m[1026]&m[1060])|(m[1023]&m[1024]&m[1025]&m[1026]&m[1060]))):InitCond[1120];
    m[1032] = run?((((m[1028]&~m[1029]&~m[1030]&~m[1031]&~m[1065])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1065])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1065])|(m[1028]&m[1029]&~m[1030]&m[1031]&~m[1065])|(m[1028]&~m[1029]&m[1030]&m[1031]&~m[1065])|(~m[1028]&m[1029]&m[1030]&m[1031]&~m[1065]))&BiasedRNG[627])|(((m[1028]&~m[1029]&~m[1030]&~m[1031]&m[1065])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&m[1065])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&m[1065])|(m[1028]&m[1029]&~m[1030]&m[1031]&m[1065])|(m[1028]&~m[1029]&m[1030]&m[1031]&m[1065])|(~m[1028]&m[1029]&m[1030]&m[1031]&m[1065]))&~BiasedRNG[627])|((m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1065])|(m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1065])|(~m[1028]&m[1029]&m[1030]&~m[1031]&~m[1065])|(m[1028]&m[1029]&m[1030]&~m[1031]&~m[1065])|(m[1028]&m[1029]&m[1030]&m[1031]&~m[1065])|(m[1028]&m[1029]&~m[1030]&~m[1031]&m[1065])|(m[1028]&~m[1029]&m[1030]&~m[1031]&m[1065])|(~m[1028]&m[1029]&m[1030]&~m[1031]&m[1065])|(m[1028]&m[1029]&m[1030]&~m[1031]&m[1065])|(m[1028]&m[1029]&m[1030]&m[1031]&m[1065]))):InitCond[1121];
    m[1037] = run?((((m[1033]&~m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&~m[1070]))&BiasedRNG[628])|(((m[1033]&~m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&m[1070]))&~BiasedRNG[628])|((m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&m[1070]))):InitCond[1122];
    m[1042] = run?((((m[1038]&~m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&~m[1075]))&BiasedRNG[629])|(((m[1038]&~m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&m[1075]))&~BiasedRNG[629])|((m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&m[1075]))):InitCond[1123];
    m[1047] = run?((((m[1043]&~m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&~m[1080]))&BiasedRNG[630])|(((m[1043]&~m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&m[1080]))&~BiasedRNG[630])|((m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&m[1080]))):InitCond[1124];
    m[1052] = run?((((m[1048]&~m[1049]&~m[1050]&~m[1051]&~m[1083])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1083])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1083])|(m[1048]&m[1049]&~m[1050]&m[1051]&~m[1083])|(m[1048]&~m[1049]&m[1050]&m[1051]&~m[1083])|(~m[1048]&m[1049]&m[1050]&m[1051]&~m[1083]))&BiasedRNG[631])|(((m[1048]&~m[1049]&~m[1050]&~m[1051]&m[1083])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&m[1083])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&m[1083])|(m[1048]&m[1049]&~m[1050]&m[1051]&m[1083])|(m[1048]&~m[1049]&m[1050]&m[1051]&m[1083])|(~m[1048]&m[1049]&m[1050]&m[1051]&m[1083]))&~BiasedRNG[631])|((m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1083])|(m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1083])|(~m[1048]&m[1049]&m[1050]&~m[1051]&~m[1083])|(m[1048]&m[1049]&m[1050]&~m[1051]&~m[1083])|(m[1048]&m[1049]&m[1050]&m[1051]&~m[1083])|(m[1048]&m[1049]&~m[1050]&~m[1051]&m[1083])|(m[1048]&~m[1049]&m[1050]&~m[1051]&m[1083])|(~m[1048]&m[1049]&m[1050]&~m[1051]&m[1083])|(m[1048]&m[1049]&m[1050]&~m[1051]&m[1083])|(m[1048]&m[1049]&m[1050]&m[1051]&m[1083]))):InitCond[1125];
    m[1057] = run?((((m[1053]&~m[1054]&~m[1055]&~m[1056]&~m[1085])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1085])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1085])|(m[1053]&m[1054]&~m[1055]&m[1056]&~m[1085])|(m[1053]&~m[1054]&m[1055]&m[1056]&~m[1085])|(~m[1053]&m[1054]&m[1055]&m[1056]&~m[1085]))&BiasedRNG[632])|(((m[1053]&~m[1054]&~m[1055]&~m[1056]&m[1085])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&m[1085])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&m[1085])|(m[1053]&m[1054]&~m[1055]&m[1056]&m[1085])|(m[1053]&~m[1054]&m[1055]&m[1056]&m[1085])|(~m[1053]&m[1054]&m[1055]&m[1056]&m[1085]))&~BiasedRNG[632])|((m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1085])|(m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1085])|(~m[1053]&m[1054]&m[1055]&~m[1056]&~m[1085])|(m[1053]&m[1054]&m[1055]&~m[1056]&~m[1085])|(m[1053]&m[1054]&m[1055]&m[1056]&~m[1085])|(m[1053]&m[1054]&~m[1055]&~m[1056]&m[1085])|(m[1053]&~m[1054]&m[1055]&~m[1056]&m[1085])|(~m[1053]&m[1054]&m[1055]&~m[1056]&m[1085])|(m[1053]&m[1054]&m[1055]&~m[1056]&m[1085])|(m[1053]&m[1054]&m[1055]&m[1056]&m[1085]))):InitCond[1126];
    m[1062] = run?((((m[1058]&~m[1059]&~m[1060]&~m[1061]&~m[1090])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1090])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1090])|(m[1058]&m[1059]&~m[1060]&m[1061]&~m[1090])|(m[1058]&~m[1059]&m[1060]&m[1061]&~m[1090])|(~m[1058]&m[1059]&m[1060]&m[1061]&~m[1090]))&BiasedRNG[633])|(((m[1058]&~m[1059]&~m[1060]&~m[1061]&m[1090])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&m[1090])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&m[1090])|(m[1058]&m[1059]&~m[1060]&m[1061]&m[1090])|(m[1058]&~m[1059]&m[1060]&m[1061]&m[1090])|(~m[1058]&m[1059]&m[1060]&m[1061]&m[1090]))&~BiasedRNG[633])|((m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1090])|(m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1090])|(~m[1058]&m[1059]&m[1060]&~m[1061]&~m[1090])|(m[1058]&m[1059]&m[1060]&~m[1061]&~m[1090])|(m[1058]&m[1059]&m[1060]&m[1061]&~m[1090])|(m[1058]&m[1059]&~m[1060]&~m[1061]&m[1090])|(m[1058]&~m[1059]&m[1060]&~m[1061]&m[1090])|(~m[1058]&m[1059]&m[1060]&~m[1061]&m[1090])|(m[1058]&m[1059]&m[1060]&~m[1061]&m[1090])|(m[1058]&m[1059]&m[1060]&m[1061]&m[1090]))):InitCond[1127];
    m[1067] = run?((((m[1063]&~m[1064]&~m[1065]&~m[1066]&~m[1095])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1095])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1095])|(m[1063]&m[1064]&~m[1065]&m[1066]&~m[1095])|(m[1063]&~m[1064]&m[1065]&m[1066]&~m[1095])|(~m[1063]&m[1064]&m[1065]&m[1066]&~m[1095]))&BiasedRNG[634])|(((m[1063]&~m[1064]&~m[1065]&~m[1066]&m[1095])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&m[1095])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&m[1095])|(m[1063]&m[1064]&~m[1065]&m[1066]&m[1095])|(m[1063]&~m[1064]&m[1065]&m[1066]&m[1095])|(~m[1063]&m[1064]&m[1065]&m[1066]&m[1095]))&~BiasedRNG[634])|((m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1095])|(m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1095])|(~m[1063]&m[1064]&m[1065]&~m[1066]&~m[1095])|(m[1063]&m[1064]&m[1065]&~m[1066]&~m[1095])|(m[1063]&m[1064]&m[1065]&m[1066]&~m[1095])|(m[1063]&m[1064]&~m[1065]&~m[1066]&m[1095])|(m[1063]&~m[1064]&m[1065]&~m[1066]&m[1095])|(~m[1063]&m[1064]&m[1065]&~m[1066]&m[1095])|(m[1063]&m[1064]&m[1065]&~m[1066]&m[1095])|(m[1063]&m[1064]&m[1065]&m[1066]&m[1095]))):InitCond[1128];
    m[1072] = run?((((m[1068]&~m[1069]&~m[1070]&~m[1071]&~m[1100])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1100])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1100])|(m[1068]&m[1069]&~m[1070]&m[1071]&~m[1100])|(m[1068]&~m[1069]&m[1070]&m[1071]&~m[1100])|(~m[1068]&m[1069]&m[1070]&m[1071]&~m[1100]))&BiasedRNG[635])|(((m[1068]&~m[1069]&~m[1070]&~m[1071]&m[1100])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&m[1100])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&m[1100])|(m[1068]&m[1069]&~m[1070]&m[1071]&m[1100])|(m[1068]&~m[1069]&m[1070]&m[1071]&m[1100])|(~m[1068]&m[1069]&m[1070]&m[1071]&m[1100]))&~BiasedRNG[635])|((m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1100])|(m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1100])|(~m[1068]&m[1069]&m[1070]&~m[1071]&~m[1100])|(m[1068]&m[1069]&m[1070]&~m[1071]&~m[1100])|(m[1068]&m[1069]&m[1070]&m[1071]&~m[1100])|(m[1068]&m[1069]&~m[1070]&~m[1071]&m[1100])|(m[1068]&~m[1069]&m[1070]&~m[1071]&m[1100])|(~m[1068]&m[1069]&m[1070]&~m[1071]&m[1100])|(m[1068]&m[1069]&m[1070]&~m[1071]&m[1100])|(m[1068]&m[1069]&m[1070]&m[1071]&m[1100]))):InitCond[1129];
    m[1077] = run?((((m[1073]&~m[1074]&~m[1075]&~m[1076]&~m[1105])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1105])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1105])|(m[1073]&m[1074]&~m[1075]&m[1076]&~m[1105])|(m[1073]&~m[1074]&m[1075]&m[1076]&~m[1105])|(~m[1073]&m[1074]&m[1075]&m[1076]&~m[1105]))&BiasedRNG[636])|(((m[1073]&~m[1074]&~m[1075]&~m[1076]&m[1105])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&m[1105])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&m[1105])|(m[1073]&m[1074]&~m[1075]&m[1076]&m[1105])|(m[1073]&~m[1074]&m[1075]&m[1076]&m[1105])|(~m[1073]&m[1074]&m[1075]&m[1076]&m[1105]))&~BiasedRNG[636])|((m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1105])|(m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1105])|(~m[1073]&m[1074]&m[1075]&~m[1076]&~m[1105])|(m[1073]&m[1074]&m[1075]&~m[1076]&~m[1105])|(m[1073]&m[1074]&m[1075]&m[1076]&~m[1105])|(m[1073]&m[1074]&~m[1075]&~m[1076]&m[1105])|(m[1073]&~m[1074]&m[1075]&~m[1076]&m[1105])|(~m[1073]&m[1074]&m[1075]&~m[1076]&m[1105])|(m[1073]&m[1074]&m[1075]&~m[1076]&m[1105])|(m[1073]&m[1074]&m[1075]&m[1076]&m[1105]))):InitCond[1130];
    m[1082] = run?((((m[1078]&~m[1079]&~m[1080]&~m[1081]&~m[1110])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1110])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1110])|(m[1078]&m[1079]&~m[1080]&m[1081]&~m[1110])|(m[1078]&~m[1079]&m[1080]&m[1081]&~m[1110])|(~m[1078]&m[1079]&m[1080]&m[1081]&~m[1110]))&BiasedRNG[637])|(((m[1078]&~m[1079]&~m[1080]&~m[1081]&m[1110])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&m[1110])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&m[1110])|(m[1078]&m[1079]&~m[1080]&m[1081]&m[1110])|(m[1078]&~m[1079]&m[1080]&m[1081]&m[1110])|(~m[1078]&m[1079]&m[1080]&m[1081]&m[1110]))&~BiasedRNG[637])|((m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1110])|(m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1110])|(~m[1078]&m[1079]&m[1080]&~m[1081]&~m[1110])|(m[1078]&m[1079]&m[1080]&~m[1081]&~m[1110])|(m[1078]&m[1079]&m[1080]&m[1081]&~m[1110])|(m[1078]&m[1079]&~m[1080]&~m[1081]&m[1110])|(m[1078]&~m[1079]&m[1080]&~m[1081]&m[1110])|(~m[1078]&m[1079]&m[1080]&~m[1081]&m[1110])|(m[1078]&m[1079]&m[1080]&~m[1081]&m[1110])|(m[1078]&m[1079]&m[1080]&m[1081]&m[1110]))):InitCond[1131];
    m[1087] = run?((((m[1083]&~m[1084]&~m[1085]&~m[1086]&~m[1113])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1113])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1113])|(m[1083]&m[1084]&~m[1085]&m[1086]&~m[1113])|(m[1083]&~m[1084]&m[1085]&m[1086]&~m[1113])|(~m[1083]&m[1084]&m[1085]&m[1086]&~m[1113]))&BiasedRNG[638])|(((m[1083]&~m[1084]&~m[1085]&~m[1086]&m[1113])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&m[1113])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&m[1113])|(m[1083]&m[1084]&~m[1085]&m[1086]&m[1113])|(m[1083]&~m[1084]&m[1085]&m[1086]&m[1113])|(~m[1083]&m[1084]&m[1085]&m[1086]&m[1113]))&~BiasedRNG[638])|((m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1113])|(m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1113])|(~m[1083]&m[1084]&m[1085]&~m[1086]&~m[1113])|(m[1083]&m[1084]&m[1085]&~m[1086]&~m[1113])|(m[1083]&m[1084]&m[1085]&m[1086]&~m[1113])|(m[1083]&m[1084]&~m[1085]&~m[1086]&m[1113])|(m[1083]&~m[1084]&m[1085]&~m[1086]&m[1113])|(~m[1083]&m[1084]&m[1085]&~m[1086]&m[1113])|(m[1083]&m[1084]&m[1085]&~m[1086]&m[1113])|(m[1083]&m[1084]&m[1085]&m[1086]&m[1113]))):InitCond[1132];
    m[1092] = run?((((m[1088]&~m[1089]&~m[1090]&~m[1091]&~m[1115])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1115])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1115])|(m[1088]&m[1089]&~m[1090]&m[1091]&~m[1115])|(m[1088]&~m[1089]&m[1090]&m[1091]&~m[1115])|(~m[1088]&m[1089]&m[1090]&m[1091]&~m[1115]))&BiasedRNG[639])|(((m[1088]&~m[1089]&~m[1090]&~m[1091]&m[1115])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&m[1115])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&m[1115])|(m[1088]&m[1089]&~m[1090]&m[1091]&m[1115])|(m[1088]&~m[1089]&m[1090]&m[1091]&m[1115])|(~m[1088]&m[1089]&m[1090]&m[1091]&m[1115]))&~BiasedRNG[639])|((m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1115])|(m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1115])|(~m[1088]&m[1089]&m[1090]&~m[1091]&~m[1115])|(m[1088]&m[1089]&m[1090]&~m[1091]&~m[1115])|(m[1088]&m[1089]&m[1090]&m[1091]&~m[1115])|(m[1088]&m[1089]&~m[1090]&~m[1091]&m[1115])|(m[1088]&~m[1089]&m[1090]&~m[1091]&m[1115])|(~m[1088]&m[1089]&m[1090]&~m[1091]&m[1115])|(m[1088]&m[1089]&m[1090]&~m[1091]&m[1115])|(m[1088]&m[1089]&m[1090]&m[1091]&m[1115]))):InitCond[1133];
    m[1097] = run?((((m[1093]&~m[1094]&~m[1095]&~m[1096]&~m[1120])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1120])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1120])|(m[1093]&m[1094]&~m[1095]&m[1096]&~m[1120])|(m[1093]&~m[1094]&m[1095]&m[1096]&~m[1120])|(~m[1093]&m[1094]&m[1095]&m[1096]&~m[1120]))&BiasedRNG[640])|(((m[1093]&~m[1094]&~m[1095]&~m[1096]&m[1120])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&m[1120])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&m[1120])|(m[1093]&m[1094]&~m[1095]&m[1096]&m[1120])|(m[1093]&~m[1094]&m[1095]&m[1096]&m[1120])|(~m[1093]&m[1094]&m[1095]&m[1096]&m[1120]))&~BiasedRNG[640])|((m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1120])|(m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1120])|(~m[1093]&m[1094]&m[1095]&~m[1096]&~m[1120])|(m[1093]&m[1094]&m[1095]&~m[1096]&~m[1120])|(m[1093]&m[1094]&m[1095]&m[1096]&~m[1120])|(m[1093]&m[1094]&~m[1095]&~m[1096]&m[1120])|(m[1093]&~m[1094]&m[1095]&~m[1096]&m[1120])|(~m[1093]&m[1094]&m[1095]&~m[1096]&m[1120])|(m[1093]&m[1094]&m[1095]&~m[1096]&m[1120])|(m[1093]&m[1094]&m[1095]&m[1096]&m[1120]))):InitCond[1134];
    m[1102] = run?((((m[1098]&~m[1099]&~m[1100]&~m[1101]&~m[1125])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1125])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1125])|(m[1098]&m[1099]&~m[1100]&m[1101]&~m[1125])|(m[1098]&~m[1099]&m[1100]&m[1101]&~m[1125])|(~m[1098]&m[1099]&m[1100]&m[1101]&~m[1125]))&BiasedRNG[641])|(((m[1098]&~m[1099]&~m[1100]&~m[1101]&m[1125])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&m[1125])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&m[1125])|(m[1098]&m[1099]&~m[1100]&m[1101]&m[1125])|(m[1098]&~m[1099]&m[1100]&m[1101]&m[1125])|(~m[1098]&m[1099]&m[1100]&m[1101]&m[1125]))&~BiasedRNG[641])|((m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1125])|(m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1125])|(~m[1098]&m[1099]&m[1100]&~m[1101]&~m[1125])|(m[1098]&m[1099]&m[1100]&~m[1101]&~m[1125])|(m[1098]&m[1099]&m[1100]&m[1101]&~m[1125])|(m[1098]&m[1099]&~m[1100]&~m[1101]&m[1125])|(m[1098]&~m[1099]&m[1100]&~m[1101]&m[1125])|(~m[1098]&m[1099]&m[1100]&~m[1101]&m[1125])|(m[1098]&m[1099]&m[1100]&~m[1101]&m[1125])|(m[1098]&m[1099]&m[1100]&m[1101]&m[1125]))):InitCond[1135];
    m[1107] = run?((((m[1103]&~m[1104]&~m[1105]&~m[1106]&~m[1130])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1130])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1130])|(m[1103]&m[1104]&~m[1105]&m[1106]&~m[1130])|(m[1103]&~m[1104]&m[1105]&m[1106]&~m[1130])|(~m[1103]&m[1104]&m[1105]&m[1106]&~m[1130]))&BiasedRNG[642])|(((m[1103]&~m[1104]&~m[1105]&~m[1106]&m[1130])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&m[1130])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&m[1130])|(m[1103]&m[1104]&~m[1105]&m[1106]&m[1130])|(m[1103]&~m[1104]&m[1105]&m[1106]&m[1130])|(~m[1103]&m[1104]&m[1105]&m[1106]&m[1130]))&~BiasedRNG[642])|((m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1130])|(m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1130])|(~m[1103]&m[1104]&m[1105]&~m[1106]&~m[1130])|(m[1103]&m[1104]&m[1105]&~m[1106]&~m[1130])|(m[1103]&m[1104]&m[1105]&m[1106]&~m[1130])|(m[1103]&m[1104]&~m[1105]&~m[1106]&m[1130])|(m[1103]&~m[1104]&m[1105]&~m[1106]&m[1130])|(~m[1103]&m[1104]&m[1105]&~m[1106]&m[1130])|(m[1103]&m[1104]&m[1105]&~m[1106]&m[1130])|(m[1103]&m[1104]&m[1105]&m[1106]&m[1130]))):InitCond[1136];
    m[1112] = run?((((m[1108]&~m[1109]&~m[1110]&~m[1111]&~m[1135])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1135])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1135])|(m[1108]&m[1109]&~m[1110]&m[1111]&~m[1135])|(m[1108]&~m[1109]&m[1110]&m[1111]&~m[1135])|(~m[1108]&m[1109]&m[1110]&m[1111]&~m[1135]))&BiasedRNG[643])|(((m[1108]&~m[1109]&~m[1110]&~m[1111]&m[1135])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&m[1135])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&m[1135])|(m[1108]&m[1109]&~m[1110]&m[1111]&m[1135])|(m[1108]&~m[1109]&m[1110]&m[1111]&m[1135])|(~m[1108]&m[1109]&m[1110]&m[1111]&m[1135]))&~BiasedRNG[643])|((m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1135])|(m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1135])|(~m[1108]&m[1109]&m[1110]&~m[1111]&~m[1135])|(m[1108]&m[1109]&m[1110]&~m[1111]&~m[1135])|(m[1108]&m[1109]&m[1110]&m[1111]&~m[1135])|(m[1108]&m[1109]&~m[1110]&~m[1111]&m[1135])|(m[1108]&~m[1109]&m[1110]&~m[1111]&m[1135])|(~m[1108]&m[1109]&m[1110]&~m[1111]&m[1135])|(m[1108]&m[1109]&m[1110]&~m[1111]&m[1135])|(m[1108]&m[1109]&m[1110]&m[1111]&m[1135]))):InitCond[1137];
    m[1117] = run?((((m[1113]&~m[1114]&~m[1115]&~m[1116]&~m[1138])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1138])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1138])|(m[1113]&m[1114]&~m[1115]&m[1116]&~m[1138])|(m[1113]&~m[1114]&m[1115]&m[1116]&~m[1138])|(~m[1113]&m[1114]&m[1115]&m[1116]&~m[1138]))&BiasedRNG[644])|(((m[1113]&~m[1114]&~m[1115]&~m[1116]&m[1138])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&m[1138])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&m[1138])|(m[1113]&m[1114]&~m[1115]&m[1116]&m[1138])|(m[1113]&~m[1114]&m[1115]&m[1116]&m[1138])|(~m[1113]&m[1114]&m[1115]&m[1116]&m[1138]))&~BiasedRNG[644])|((m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1138])|(m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1138])|(~m[1113]&m[1114]&m[1115]&~m[1116]&~m[1138])|(m[1113]&m[1114]&m[1115]&~m[1116]&~m[1138])|(m[1113]&m[1114]&m[1115]&m[1116]&~m[1138])|(m[1113]&m[1114]&~m[1115]&~m[1116]&m[1138])|(m[1113]&~m[1114]&m[1115]&~m[1116]&m[1138])|(~m[1113]&m[1114]&m[1115]&~m[1116]&m[1138])|(m[1113]&m[1114]&m[1115]&~m[1116]&m[1138])|(m[1113]&m[1114]&m[1115]&m[1116]&m[1138]))):InitCond[1138];
    m[1122] = run?((((m[1118]&~m[1119]&~m[1120]&~m[1121]&~m[1140])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1140])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1140])|(m[1118]&m[1119]&~m[1120]&m[1121]&~m[1140])|(m[1118]&~m[1119]&m[1120]&m[1121]&~m[1140])|(~m[1118]&m[1119]&m[1120]&m[1121]&~m[1140]))&BiasedRNG[645])|(((m[1118]&~m[1119]&~m[1120]&~m[1121]&m[1140])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&m[1140])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&m[1140])|(m[1118]&m[1119]&~m[1120]&m[1121]&m[1140])|(m[1118]&~m[1119]&m[1120]&m[1121]&m[1140])|(~m[1118]&m[1119]&m[1120]&m[1121]&m[1140]))&~BiasedRNG[645])|((m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1140])|(m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1140])|(~m[1118]&m[1119]&m[1120]&~m[1121]&~m[1140])|(m[1118]&m[1119]&m[1120]&~m[1121]&~m[1140])|(m[1118]&m[1119]&m[1120]&m[1121]&~m[1140])|(m[1118]&m[1119]&~m[1120]&~m[1121]&m[1140])|(m[1118]&~m[1119]&m[1120]&~m[1121]&m[1140])|(~m[1118]&m[1119]&m[1120]&~m[1121]&m[1140])|(m[1118]&m[1119]&m[1120]&~m[1121]&m[1140])|(m[1118]&m[1119]&m[1120]&m[1121]&m[1140]))):InitCond[1139];
    m[1127] = run?((((m[1123]&~m[1124]&~m[1125]&~m[1126]&~m[1145])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1145])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1145])|(m[1123]&m[1124]&~m[1125]&m[1126]&~m[1145])|(m[1123]&~m[1124]&m[1125]&m[1126]&~m[1145])|(~m[1123]&m[1124]&m[1125]&m[1126]&~m[1145]))&BiasedRNG[646])|(((m[1123]&~m[1124]&~m[1125]&~m[1126]&m[1145])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&m[1145])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&m[1145])|(m[1123]&m[1124]&~m[1125]&m[1126]&m[1145])|(m[1123]&~m[1124]&m[1125]&m[1126]&m[1145])|(~m[1123]&m[1124]&m[1125]&m[1126]&m[1145]))&~BiasedRNG[646])|((m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1145])|(m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1145])|(~m[1123]&m[1124]&m[1125]&~m[1126]&~m[1145])|(m[1123]&m[1124]&m[1125]&~m[1126]&~m[1145])|(m[1123]&m[1124]&m[1125]&m[1126]&~m[1145])|(m[1123]&m[1124]&~m[1125]&~m[1126]&m[1145])|(m[1123]&~m[1124]&m[1125]&~m[1126]&m[1145])|(~m[1123]&m[1124]&m[1125]&~m[1126]&m[1145])|(m[1123]&m[1124]&m[1125]&~m[1126]&m[1145])|(m[1123]&m[1124]&m[1125]&m[1126]&m[1145]))):InitCond[1140];
    m[1132] = run?((((m[1128]&~m[1129]&~m[1130]&~m[1131]&~m[1150])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1150])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1150])|(m[1128]&m[1129]&~m[1130]&m[1131]&~m[1150])|(m[1128]&~m[1129]&m[1130]&m[1131]&~m[1150])|(~m[1128]&m[1129]&m[1130]&m[1131]&~m[1150]))&BiasedRNG[647])|(((m[1128]&~m[1129]&~m[1130]&~m[1131]&m[1150])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&m[1150])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&m[1150])|(m[1128]&m[1129]&~m[1130]&m[1131]&m[1150])|(m[1128]&~m[1129]&m[1130]&m[1131]&m[1150])|(~m[1128]&m[1129]&m[1130]&m[1131]&m[1150]))&~BiasedRNG[647])|((m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1150])|(m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1150])|(~m[1128]&m[1129]&m[1130]&~m[1131]&~m[1150])|(m[1128]&m[1129]&m[1130]&~m[1131]&~m[1150])|(m[1128]&m[1129]&m[1130]&m[1131]&~m[1150])|(m[1128]&m[1129]&~m[1130]&~m[1131]&m[1150])|(m[1128]&~m[1129]&m[1130]&~m[1131]&m[1150])|(~m[1128]&m[1129]&m[1130]&~m[1131]&m[1150])|(m[1128]&m[1129]&m[1130]&~m[1131]&m[1150])|(m[1128]&m[1129]&m[1130]&m[1131]&m[1150]))):InitCond[1141];
    m[1137] = run?((((m[1133]&~m[1134]&~m[1135]&~m[1136]&~m[1155])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1155])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1155])|(m[1133]&m[1134]&~m[1135]&m[1136]&~m[1155])|(m[1133]&~m[1134]&m[1135]&m[1136]&~m[1155])|(~m[1133]&m[1134]&m[1135]&m[1136]&~m[1155]))&BiasedRNG[648])|(((m[1133]&~m[1134]&~m[1135]&~m[1136]&m[1155])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&m[1155])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&m[1155])|(m[1133]&m[1134]&~m[1135]&m[1136]&m[1155])|(m[1133]&~m[1134]&m[1135]&m[1136]&m[1155])|(~m[1133]&m[1134]&m[1135]&m[1136]&m[1155]))&~BiasedRNG[648])|((m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1155])|(m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1155])|(~m[1133]&m[1134]&m[1135]&~m[1136]&~m[1155])|(m[1133]&m[1134]&m[1135]&~m[1136]&~m[1155])|(m[1133]&m[1134]&m[1135]&m[1136]&~m[1155])|(m[1133]&m[1134]&~m[1135]&~m[1136]&m[1155])|(m[1133]&~m[1134]&m[1135]&~m[1136]&m[1155])|(~m[1133]&m[1134]&m[1135]&~m[1136]&m[1155])|(m[1133]&m[1134]&m[1135]&~m[1136]&m[1155])|(m[1133]&m[1134]&m[1135]&m[1136]&m[1155]))):InitCond[1142];
    m[1142] = run?((((m[1138]&~m[1139]&~m[1140]&~m[1141]&~m[1158])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1158])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1158])|(m[1138]&m[1139]&~m[1140]&m[1141]&~m[1158])|(m[1138]&~m[1139]&m[1140]&m[1141]&~m[1158])|(~m[1138]&m[1139]&m[1140]&m[1141]&~m[1158]))&BiasedRNG[649])|(((m[1138]&~m[1139]&~m[1140]&~m[1141]&m[1158])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&m[1158])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&m[1158])|(m[1138]&m[1139]&~m[1140]&m[1141]&m[1158])|(m[1138]&~m[1139]&m[1140]&m[1141]&m[1158])|(~m[1138]&m[1139]&m[1140]&m[1141]&m[1158]))&~BiasedRNG[649])|((m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1158])|(m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1158])|(~m[1138]&m[1139]&m[1140]&~m[1141]&~m[1158])|(m[1138]&m[1139]&m[1140]&~m[1141]&~m[1158])|(m[1138]&m[1139]&m[1140]&m[1141]&~m[1158])|(m[1138]&m[1139]&~m[1140]&~m[1141]&m[1158])|(m[1138]&~m[1139]&m[1140]&~m[1141]&m[1158])|(~m[1138]&m[1139]&m[1140]&~m[1141]&m[1158])|(m[1138]&m[1139]&m[1140]&~m[1141]&m[1158])|(m[1138]&m[1139]&m[1140]&m[1141]&m[1158]))):InitCond[1143];
    m[1147] = run?((((m[1143]&~m[1144]&~m[1145]&~m[1146]&~m[1160])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1160])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1160])|(m[1143]&m[1144]&~m[1145]&m[1146]&~m[1160])|(m[1143]&~m[1144]&m[1145]&m[1146]&~m[1160])|(~m[1143]&m[1144]&m[1145]&m[1146]&~m[1160]))&BiasedRNG[650])|(((m[1143]&~m[1144]&~m[1145]&~m[1146]&m[1160])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&m[1160])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&m[1160])|(m[1143]&m[1144]&~m[1145]&m[1146]&m[1160])|(m[1143]&~m[1144]&m[1145]&m[1146]&m[1160])|(~m[1143]&m[1144]&m[1145]&m[1146]&m[1160]))&~BiasedRNG[650])|((m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1160])|(m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1160])|(~m[1143]&m[1144]&m[1145]&~m[1146]&~m[1160])|(m[1143]&m[1144]&m[1145]&~m[1146]&~m[1160])|(m[1143]&m[1144]&m[1145]&m[1146]&~m[1160])|(m[1143]&m[1144]&~m[1145]&~m[1146]&m[1160])|(m[1143]&~m[1144]&m[1145]&~m[1146]&m[1160])|(~m[1143]&m[1144]&m[1145]&~m[1146]&m[1160])|(m[1143]&m[1144]&m[1145]&~m[1146]&m[1160])|(m[1143]&m[1144]&m[1145]&m[1146]&m[1160]))):InitCond[1144];
    m[1152] = run?((((m[1148]&~m[1149]&~m[1150]&~m[1151]&~m[1165])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1165])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1165])|(m[1148]&m[1149]&~m[1150]&m[1151]&~m[1165])|(m[1148]&~m[1149]&m[1150]&m[1151]&~m[1165])|(~m[1148]&m[1149]&m[1150]&m[1151]&~m[1165]))&BiasedRNG[651])|(((m[1148]&~m[1149]&~m[1150]&~m[1151]&m[1165])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&m[1165])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&m[1165])|(m[1148]&m[1149]&~m[1150]&m[1151]&m[1165])|(m[1148]&~m[1149]&m[1150]&m[1151]&m[1165])|(~m[1148]&m[1149]&m[1150]&m[1151]&m[1165]))&~BiasedRNG[651])|((m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1165])|(m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1165])|(~m[1148]&m[1149]&m[1150]&~m[1151]&~m[1165])|(m[1148]&m[1149]&m[1150]&~m[1151]&~m[1165])|(m[1148]&m[1149]&m[1150]&m[1151]&~m[1165])|(m[1148]&m[1149]&~m[1150]&~m[1151]&m[1165])|(m[1148]&~m[1149]&m[1150]&~m[1151]&m[1165])|(~m[1148]&m[1149]&m[1150]&~m[1151]&m[1165])|(m[1148]&m[1149]&m[1150]&~m[1151]&m[1165])|(m[1148]&m[1149]&m[1150]&m[1151]&m[1165]))):InitCond[1145];
    m[1157] = run?((((m[1153]&~m[1154]&~m[1155]&~m[1156]&~m[1170])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1170])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1170])|(m[1153]&m[1154]&~m[1155]&m[1156]&~m[1170])|(m[1153]&~m[1154]&m[1155]&m[1156]&~m[1170])|(~m[1153]&m[1154]&m[1155]&m[1156]&~m[1170]))&BiasedRNG[652])|(((m[1153]&~m[1154]&~m[1155]&~m[1156]&m[1170])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&m[1170])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&m[1170])|(m[1153]&m[1154]&~m[1155]&m[1156]&m[1170])|(m[1153]&~m[1154]&m[1155]&m[1156]&m[1170])|(~m[1153]&m[1154]&m[1155]&m[1156]&m[1170]))&~BiasedRNG[652])|((m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1170])|(m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1170])|(~m[1153]&m[1154]&m[1155]&~m[1156]&~m[1170])|(m[1153]&m[1154]&m[1155]&~m[1156]&~m[1170])|(m[1153]&m[1154]&m[1155]&m[1156]&~m[1170])|(m[1153]&m[1154]&~m[1155]&~m[1156]&m[1170])|(m[1153]&~m[1154]&m[1155]&~m[1156]&m[1170])|(~m[1153]&m[1154]&m[1155]&~m[1156]&m[1170])|(m[1153]&m[1154]&m[1155]&~m[1156]&m[1170])|(m[1153]&m[1154]&m[1155]&m[1156]&m[1170]))):InitCond[1146];
    m[1162] = run?((((m[1158]&~m[1159]&~m[1160]&~m[1161]&~m[1173])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1173])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1173])|(m[1158]&m[1159]&~m[1160]&m[1161]&~m[1173])|(m[1158]&~m[1159]&m[1160]&m[1161]&~m[1173])|(~m[1158]&m[1159]&m[1160]&m[1161]&~m[1173]))&BiasedRNG[653])|(((m[1158]&~m[1159]&~m[1160]&~m[1161]&m[1173])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&m[1173])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&m[1173])|(m[1158]&m[1159]&~m[1160]&m[1161]&m[1173])|(m[1158]&~m[1159]&m[1160]&m[1161]&m[1173])|(~m[1158]&m[1159]&m[1160]&m[1161]&m[1173]))&~BiasedRNG[653])|((m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1173])|(m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1173])|(~m[1158]&m[1159]&m[1160]&~m[1161]&~m[1173])|(m[1158]&m[1159]&m[1160]&~m[1161]&~m[1173])|(m[1158]&m[1159]&m[1160]&m[1161]&~m[1173])|(m[1158]&m[1159]&~m[1160]&~m[1161]&m[1173])|(m[1158]&~m[1159]&m[1160]&~m[1161]&m[1173])|(~m[1158]&m[1159]&m[1160]&~m[1161]&m[1173])|(m[1158]&m[1159]&m[1160]&~m[1161]&m[1173])|(m[1158]&m[1159]&m[1160]&m[1161]&m[1173]))):InitCond[1147];
    m[1167] = run?((((m[1163]&~m[1164]&~m[1165]&~m[1166]&~m[1175])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1175])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1175])|(m[1163]&m[1164]&~m[1165]&m[1166]&~m[1175])|(m[1163]&~m[1164]&m[1165]&m[1166]&~m[1175])|(~m[1163]&m[1164]&m[1165]&m[1166]&~m[1175]))&BiasedRNG[654])|(((m[1163]&~m[1164]&~m[1165]&~m[1166]&m[1175])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&m[1175])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&m[1175])|(m[1163]&m[1164]&~m[1165]&m[1166]&m[1175])|(m[1163]&~m[1164]&m[1165]&m[1166]&m[1175])|(~m[1163]&m[1164]&m[1165]&m[1166]&m[1175]))&~BiasedRNG[654])|((m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1175])|(m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1175])|(~m[1163]&m[1164]&m[1165]&~m[1166]&~m[1175])|(m[1163]&m[1164]&m[1165]&~m[1166]&~m[1175])|(m[1163]&m[1164]&m[1165]&m[1166]&~m[1175])|(m[1163]&m[1164]&~m[1165]&~m[1166]&m[1175])|(m[1163]&~m[1164]&m[1165]&~m[1166]&m[1175])|(~m[1163]&m[1164]&m[1165]&~m[1166]&m[1175])|(m[1163]&m[1164]&m[1165]&~m[1166]&m[1175])|(m[1163]&m[1164]&m[1165]&m[1166]&m[1175]))):InitCond[1148];
    m[1172] = run?((((m[1168]&~m[1169]&~m[1170]&~m[1171]&~m[1180])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1180])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1180])|(m[1168]&m[1169]&~m[1170]&m[1171]&~m[1180])|(m[1168]&~m[1169]&m[1170]&m[1171]&~m[1180])|(~m[1168]&m[1169]&m[1170]&m[1171]&~m[1180]))&BiasedRNG[655])|(((m[1168]&~m[1169]&~m[1170]&~m[1171]&m[1180])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&m[1180])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&m[1180])|(m[1168]&m[1169]&~m[1170]&m[1171]&m[1180])|(m[1168]&~m[1169]&m[1170]&m[1171]&m[1180])|(~m[1168]&m[1169]&m[1170]&m[1171]&m[1180]))&~BiasedRNG[655])|((m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1180])|(m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1180])|(~m[1168]&m[1169]&m[1170]&~m[1171]&~m[1180])|(m[1168]&m[1169]&m[1170]&~m[1171]&~m[1180])|(m[1168]&m[1169]&m[1170]&m[1171]&~m[1180])|(m[1168]&m[1169]&~m[1170]&~m[1171]&m[1180])|(m[1168]&~m[1169]&m[1170]&~m[1171]&m[1180])|(~m[1168]&m[1169]&m[1170]&~m[1171]&m[1180])|(m[1168]&m[1169]&m[1170]&~m[1171]&m[1180])|(m[1168]&m[1169]&m[1170]&m[1171]&m[1180]))):InitCond[1149];
    m[1177] = run?((((m[1173]&~m[1174]&~m[1175]&~m[1176]&~m[1183])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1183])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1183])|(m[1173]&m[1174]&~m[1175]&m[1176]&~m[1183])|(m[1173]&~m[1174]&m[1175]&m[1176]&~m[1183])|(~m[1173]&m[1174]&m[1175]&m[1176]&~m[1183]))&BiasedRNG[656])|(((m[1173]&~m[1174]&~m[1175]&~m[1176]&m[1183])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&m[1183])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&m[1183])|(m[1173]&m[1174]&~m[1175]&m[1176]&m[1183])|(m[1173]&~m[1174]&m[1175]&m[1176]&m[1183])|(~m[1173]&m[1174]&m[1175]&m[1176]&m[1183]))&~BiasedRNG[656])|((m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1183])|(m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1183])|(~m[1173]&m[1174]&m[1175]&~m[1176]&~m[1183])|(m[1173]&m[1174]&m[1175]&~m[1176]&~m[1183])|(m[1173]&m[1174]&m[1175]&m[1176]&~m[1183])|(m[1173]&m[1174]&~m[1175]&~m[1176]&m[1183])|(m[1173]&~m[1174]&m[1175]&~m[1176]&m[1183])|(~m[1173]&m[1174]&m[1175]&~m[1176]&m[1183])|(m[1173]&m[1174]&m[1175]&~m[1176]&m[1183])|(m[1173]&m[1174]&m[1175]&m[1176]&m[1183]))):InitCond[1150];
    m[1182] = run?((((m[1178]&~m[1179]&~m[1180]&~m[1181]&~m[1185])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1185])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1185])|(m[1178]&m[1179]&~m[1180]&m[1181]&~m[1185])|(m[1178]&~m[1179]&m[1180]&m[1181]&~m[1185])|(~m[1178]&m[1179]&m[1180]&m[1181]&~m[1185]))&BiasedRNG[657])|(((m[1178]&~m[1179]&~m[1180]&~m[1181]&m[1185])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&m[1185])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&m[1185])|(m[1178]&m[1179]&~m[1180]&m[1181]&m[1185])|(m[1178]&~m[1179]&m[1180]&m[1181]&m[1185])|(~m[1178]&m[1179]&m[1180]&m[1181]&m[1185]))&~BiasedRNG[657])|((m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1185])|(m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1185])|(~m[1178]&m[1179]&m[1180]&~m[1181]&~m[1185])|(m[1178]&m[1179]&m[1180]&~m[1181]&~m[1185])|(m[1178]&m[1179]&m[1180]&m[1181]&~m[1185])|(m[1178]&m[1179]&~m[1180]&~m[1181]&m[1185])|(m[1178]&~m[1179]&m[1180]&~m[1181]&m[1185])|(~m[1178]&m[1179]&m[1180]&~m[1181]&m[1185])|(m[1178]&m[1179]&m[1180]&~m[1181]&m[1185])|(m[1178]&m[1179]&m[1180]&m[1181]&m[1185]))):InitCond[1151];
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[109]&LFSRcolor0[274]&LFSRcolor0[582]);
    BiasedRNG[1] = (LFSRcolor0[124]&LFSRcolor0[211]&LFSRcolor0[443]);
    BiasedRNG[2] = (LFSRcolor0[473]&LFSRcolor0[110]&LFSRcolor0[400]);
    BiasedRNG[3] = (LFSRcolor0[526]&LFSRcolor0[578]&LFSRcolor0[604]);
    BiasedRNG[4] = (LFSRcolor0[261]&LFSRcolor0[481]&LFSRcolor0[310]);
    BiasedRNG[5] = (LFSRcolor0[525]&LFSRcolor0[237]&LFSRcolor0[123]);
    BiasedRNG[6] = (LFSRcolor0[133]&LFSRcolor0[98]&LFSRcolor0[6]);
    BiasedRNG[7] = (LFSRcolor0[329]&LFSRcolor0[411]&LFSRcolor0[511]);
    BiasedRNG[8] = (LFSRcolor0[149]&LFSRcolor0[77]&LFSRcolor0[167]);
    BiasedRNG[9] = (LFSRcolor0[279]&LFSRcolor0[560]&LFSRcolor0[20]);
    BiasedRNG[10] = (LFSRcolor0[242]&LFSRcolor0[491]&LFSRcolor0[386]);
    BiasedRNG[11] = (LFSRcolor0[224]&LFSRcolor0[436]&LFSRcolor0[565]);
    BiasedRNG[12] = (LFSRcolor0[137]&LFSRcolor0[379]&LFSRcolor0[212]);
    BiasedRNG[13] = (LFSRcolor0[332]&LFSRcolor0[451]&LFSRcolor0[99]);
    BiasedRNG[14] = (LFSRcolor0[394]&LFSRcolor0[160]&LFSRcolor0[81]);
    BiasedRNG[15] = (LFSRcolor0[267]&LFSRcolor0[170]&LFSRcolor0[221]);
    BiasedRNG[16] = (LFSRcolor0[157]&LFSRcolor0[186]&LFSRcolor0[402]);
    BiasedRNG[17] = (LFSRcolor0[58]&LFSRcolor0[487]&LFSRcolor0[255]);
    BiasedRNG[18] = (LFSRcolor0[201]&LFSRcolor0[388]&LFSRcolor0[333]);
    BiasedRNG[19] = (LFSRcolor0[0]&LFSRcolor0[638]&LFSRcolor0[609]);
    BiasedRNG[20] = (LFSRcolor0[340]&LFSRcolor0[338]&LFSRcolor0[571]);
    BiasedRNG[21] = (LFSRcolor0[629]&LFSRcolor0[618]&LFSRcolor0[189]);
    BiasedRNG[22] = (LFSRcolor0[492]&LFSRcolor0[430]&LFSRcolor0[431]);
    BiasedRNG[23] = (LFSRcolor0[320]&LFSRcolor0[464]&LFSRcolor0[193]);
    BiasedRNG[24] = (LFSRcolor0[302]&LFSRcolor0[74]&LFSRcolor0[566]);
    BiasedRNG[25] = (LFSRcolor0[512]&LFSRcolor0[420]&LFSRcolor0[327]);
    BiasedRNG[26] = (LFSRcolor0[115]&LFSRcolor0[184]&LFSRcolor0[369]);
    BiasedRNG[27] = (LFSRcolor0[544]&LFSRcolor0[312]&LFSRcolor0[469]);
    BiasedRNG[28] = (LFSRcolor0[631]&LFSRcolor0[396]&LFSRcolor0[60]);
    BiasedRNG[29] = (LFSRcolor0[276]&LFSRcolor0[513]&LFSRcolor0[19]);
    BiasedRNG[30] = (LFSRcolor0[514]&LFSRcolor0[527]&LFSRcolor0[387]);
    BiasedRNG[31] = (LFSRcolor0[277]&LFSRcolor0[105]&LFSRcolor0[561]);
    BiasedRNG[32] = (LFSRcolor0[307]&LFSRcolor0[182]&LFSRcolor0[410]);
    BiasedRNG[33] = (LFSRcolor0[367]&LFSRcolor0[57]&LFSRcolor0[465]);
    BiasedRNG[34] = (LFSRcolor0[100]&LFSRcolor0[96]&LFSRcolor0[381]);
    BiasedRNG[35] = (LFSRcolor0[401]&LFSRcolor0[339]&LFSRcolor0[342]);
    BiasedRNG[36] = (LFSRcolor0[48]&LFSRcolor0[59]&LFSRcolor0[501]);
    BiasedRNG[37] = (LFSRcolor0[523]&LFSRcolor0[608]&LFSRcolor0[572]);
    BiasedRNG[38] = (LFSRcolor0[304]&LFSRcolor0[321]&LFSRcolor0[116]);
    BiasedRNG[39] = (LFSRcolor0[169]&LFSRcolor0[43]&LFSRcolor0[318]);
    BiasedRNG[40] = (LFSRcolor0[426]&LFSRcolor0[2]&LFSRcolor0[223]);
    BiasedRNG[41] = (LFSRcolor0[29]&LFSRcolor0[150]&LFSRcolor0[245]);
    BiasedRNG[42] = (LFSRcolor0[493]&LFSRcolor0[90]&LFSRcolor0[603]);
    BiasedRNG[43] = (LFSRcolor0[591]&LFSRcolor0[536]&LFSRcolor0[219]);
    BiasedRNG[44] = (LFSRcolor0[635]&LFSRcolor0[268]&LFSRcolor0[1]);
    BiasedRNG[45] = (LFSRcolor0[642]&LFSRcolor0[534]&LFSRcolor0[637]);
    BiasedRNG[46] = (LFSRcolor0[370]&LFSRcolor0[611]&LFSRcolor0[50]);
    BiasedRNG[47] = (LFSRcolor0[437]&LFSRcolor0[295]&LFSRcolor0[73]);
    BiasedRNG[48] = (LFSRcolor0[587]&LFSRcolor0[78]&LFSRcolor0[432]);
    BiasedRNG[49] = (LFSRcolor0[89]&LFSRcolor0[383]&LFSRcolor0[68]);
    BiasedRNG[50] = (LFSRcolor0[517]&LFSRcolor0[316]&LFSRcolor0[232]);
    BiasedRNG[51] = (LFSRcolor0[380]&LFSRcolor0[417]&LFSRcolor0[577]);
    BiasedRNG[52] = (LFSRcolor0[282]&LFSRcolor0[489]&LFSRcolor0[500]);
    BiasedRNG[53] = (LFSRcolor0[305]&LFSRcolor0[583]&LFSRcolor0[357]);
    BiasedRNG[54] = (LFSRcolor0[217]&LFSRcolor0[484]&LFSRcolor0[197]);
    BiasedRNG[55] = (LFSRcolor0[288]&LFSRcolor0[529]&LFSRcolor0[117]);
    BiasedRNG[56] = (LFSRcolor0[7]&LFSRcolor0[438]&LFSRcolor0[272]);
    BiasedRNG[57] = (LFSRcolor0[128]&LFSRcolor0[238]&LFSRcolor0[522]);
    BiasedRNG[58] = (LFSRcolor0[331]&LFSRcolor0[102]&LFSRcolor0[630]);
    BiasedRNG[59] = (LFSRcolor0[207]&LFSRcolor0[356]&LFSRcolor0[176]);
    BiasedRNG[60] = (LFSRcolor0[270]&LFSRcolor0[414]&LFSRcolor0[28]);
    BiasedRNG[61] = (LFSRcolor0[328]&LFSRcolor0[247]&LFSRcolor0[472]);
    BiasedRNG[62] = (LFSRcolor0[343]&LFSRcolor0[4]&LFSRcolor0[138]);
    BiasedRNG[63] = (LFSRcolor0[289]&LFSRcolor0[290]&LFSRcolor0[434]);
    BiasedRNG[64] = (LFSRcolor0[549]&LFSRcolor0[161]&LFSRcolor0[163]);
    BiasedRNG[65] = (LFSRcolor0[15]&LFSRcolor0[38]&LFSRcolor0[459]);
    BiasedRNG[66] = (LFSRcolor0[558]&LFSRcolor0[252]&LFSRcolor0[65]);
    BiasedRNG[67] = (LFSRcolor0[446]&LFSRcolor0[415]&LFSRcolor0[580]);
    BiasedRNG[68] = (LFSRcolor0[361]&LFSRcolor0[480]&LFSRcolor0[21]);
    BiasedRNG[69] = (LFSRcolor0[111]&LFSRcolor0[405]&LFSRcolor0[376]);
    BiasedRNG[70] = (LFSRcolor0[323]&LFSRcolor0[130]&LFSRcolor0[398]);
    BiasedRNG[71] = (LFSRcolor0[563]&LFSRcolor0[249]&LFSRcolor0[265]);
    BiasedRNG[72] = (LFSRcolor0[449]&LFSRcolor0[168]&LFSRcolor0[260]);
    BiasedRNG[73] = (LFSRcolor0[222]&LFSRcolor0[435]&LFSRcolor0[300]);
    BiasedRNG[74] = (LFSRcolor0[142]&LFSRcolor0[395]&LFSRcolor0[588]);
    BiasedRNG[75] = (LFSRcolor0[240]&LFSRcolor0[225]&LFSRcolor0[208]);
    BiasedRNG[76] = (LFSRcolor0[542]&LFSRcolor0[205]&LFSRcolor0[546]);
    BiasedRNG[77] = (LFSRcolor0[94]&LFSRcolor0[551]&LFSRcolor0[362]);
    BiasedRNG[78] = (LFSRcolor0[605]&LFSRcolor0[334]&LFSRcolor0[27]);
    BiasedRNG[79] = (LFSRcolor0[524]&LFSRcolor0[594]&LFSRcolor0[421]);
    BiasedRNG[80] = (LFSRcolor0[363]&LFSRcolor0[423]&LFSRcolor0[155]);
    BiasedRNG[81] = (LFSRcolor0[34]&LFSRcolor0[624]&LFSRcolor0[241]);
    BiasedRNG[82] = (LFSRcolor0[204]&LFSRcolor0[151]&LFSRcolor0[425]);
    BiasedRNG[83] = (LFSRcolor0[453]&LFSRcolor0[385]&LFSRcolor0[203]);
    BiasedRNG[84] = (LFSRcolor0[570]&LFSRcolor0[519]&LFSRcolor0[234]);
    BiasedRNG[85] = (LFSRcolor0[424]&LFSRcolor0[298]&LFSRcolor0[456]);
    BiasedRNG[86] = (LFSRcolor0[403]&LFSRcolor0[462]&LFSRcolor0[346]);
    BiasedRNG[87] = (LFSRcolor0[56]&LFSRcolor0[541]&LFSRcolor0[538]);
    BiasedRNG[88] = (LFSRcolor0[602]&LFSRcolor0[141]&LFSRcolor0[72]);
    BiasedRNG[89] = (LFSRcolor0[273]&LFSRcolor0[470]&LFSRcolor0[474]);
    BiasedRNG[90] = (LFSRcolor0[627]&LFSRcolor0[303]&LFSRcolor0[353]);
    BiasedRNG[91] = (LFSRcolor0[291]&LFSRcolor0[496]&LFSRcolor0[589]);
    BiasedRNG[92] = (LFSRcolor0[409]&LFSRcolor0[40]&LFSRcolor0[412]);
    BiasedRNG[93] = (LFSRcolor0[145]&LFSRcolor0[122]&LFSRcolor0[358]);
    BiasedRNG[94] = (LFSRcolor0[45]&LFSRcolor0[520]&LFSRcolor0[528]);
    BiasedRNG[95] = (LFSRcolor0[69]&LFSRcolor0[550]&LFSRcolor0[159]);
    BiasedRNG[96] = (LFSRcolor0[485]&LFSRcolor0[299]&LFSRcolor0[278]);
    BiasedRNG[97] = (LFSRcolor0[239]&LFSRcolor0[294]&LFSRcolor0[475]);
    BiasedRNG[98] = (LFSRcolor0[359]&LFSRcolor0[350]&LFSRcolor0[18]);
    BiasedRNG[99] = (LFSRcolor0[505]&LFSRcolor0[601]&LFSRcolor0[621]);
    BiasedRNG[100] = (LFSRcolor0[336]&LFSRcolor0[119]&LFSRcolor0[557]);
    BiasedRNG[101] = (LFSRcolor0[576]&LFSRcolor0[344]&LFSRcolor0[131]);
    BiasedRNG[102] = (LFSRcolor0[132]&LFSRcolor0[498]&LFSRcolor0[226]);
    BiasedRNG[103] = (LFSRcolor0[548]&LFSRcolor0[372]&LFSRcolor0[44]);
    BiasedRNG[104] = (LFSRcolor0[552]&LFSRcolor0[171]&LFSRcolor0[228]);
    BiasedRNG[105] = (LFSRcolor0[619]&LFSRcolor0[190]&LFSRcolor0[553]);
    BiasedRNG[106] = (LFSRcolor0[17]&LFSRcolor0[82]&LFSRcolor0[134]);
    BiasedRNG[107] = (LFSRcolor0[482]&LFSRcolor0[172]&LFSRcolor0[384]);
    BiasedRNG[108] = (LFSRcolor0[354]&LFSRcolor0[508]&LFSRcolor0[97]);
    BiasedRNG[109] = (LFSRcolor0[216]&LFSRcolor0[313]&LFSRcolor0[61]);
    BiasedRNG[110] = (LFSRcolor0[194]&LFSRcolor0[214]&LFSRcolor0[486]);
    BiasedRNG[111] = (LFSRcolor0[626]&LFSRcolor0[259]&LFSRcolor0[269]);
    BiasedRNG[112] = (LFSRcolor0[399]&LFSRcolor0[140]&LFSRcolor0[191]);
    BiasedRNG[113] = (LFSRcolor0[337]&LFSRcolor0[539]&LFSRcolor0[573]);
    BiasedRNG[114] = (LFSRcolor0[515]&LFSRcolor0[63]&LFSRcolor0[562]);
    BiasedRNG[115] = (LFSRcolor0[187]&LFSRcolor0[66]&LFSRcolor0[64]);
    BiasedRNG[116] = (LFSRcolor0[46]&LFSRcolor0[506]&LFSRcolor0[364]);
    BiasedRNG[117] = (LFSRcolor0[227]&LFSRcolor0[585]&LFSRcolor0[596]);
    BiasedRNG[118] = (LFSRcolor0[5]&LFSRcolor0[617]&LFSRcolor0[545]);
    BiasedRNG[119] = (LFSRcolor0[389]&LFSRcolor0[590]&LFSRcolor0[91]);
    BiasedRNG[120] = (LFSRcolor0[174]&LFSRcolor0[341]&LFSRcolor0[628]);
    BiasedRNG[121] = (LFSRcolor0[112]&LFSRcolor0[88]&LFSRcolor0[445]);
    BiasedRNG[122] = (LFSRcolor0[251]&LFSRcolor0[62]&LFSRcolor0[407]);
    BiasedRNG[123] = (LFSRcolor0[375]&LFSRcolor0[166]&LFSRcolor0[218]);
    BiasedRNG[124] = (LFSRcolor0[153]&LFSRcolor0[236]&LFSRcolor0[429]);
    BiasedRNG[125] = (LFSRcolor0[139]&LFSRcolor0[80]&LFSRcolor0[510]);
    BiasedRNG[126] = (LFSRcolor0[8]&LFSRcolor0[3]&LFSRcolor0[324]);
    BiasedRNG[127] = (LFSRcolor0[285]&LFSRcolor0[450]&LFSRcolor0[365]);
    BiasedRNG[128] = (LFSRcolor0[579]&LFSRcolor0[360]&LFSRcolor0[185]);
    BiasedRNG[129] = (LFSRcolor0[250]&LFSRcolor0[556]&LFSRcolor0[607]);
    BiasedRNG[130] = (LFSRcolor0[537]&LFSRcolor0[235]&LFSRcolor0[49]);
    BiasedRNG[131] = (LFSRcolor0[559]&LFSRcolor0[547]&LFSRcolor0[516]);
    BiasedRNG[132] = (LFSRcolor0[416]&LFSRcolor0[92]&LFSRcolor0[317]);
    BiasedRNG[133] = (LFSRcolor0[366]&LFSRcolor0[467]&LFSRcolor0[455]);
    BiasedRNG[134] = (LFSRcolor0[30]&LFSRcolor0[67]&LFSRcolor0[292]);
    BiasedRNG[135] = (LFSRcolor0[85]&LFSRcolor0[36]&LFSRcolor0[616]);
    BiasedRNG[136] = (LFSRcolor0[136]&LFSRcolor0[23]&LFSRcolor0[502]);
    BiasedRNG[137] = (LFSRcolor0[640]&LFSRcolor0[35]&LFSRcolor0[54]);
    BiasedRNG[138] = (LFSRcolor0[256]&LFSRcolor0[597]&LFSRcolor0[419]);
    BiasedRNG[139] = (LFSRcolor0[495]&LFSRcolor0[271]&LFSRcolor0[206]);
    BiasedRNG[140] = (LFSRcolor0[293]&LFSRcolor0[404]&LFSRcolor0[262]);
    BiasedRNG[141] = (LFSRcolor0[377]&LFSRcolor0[352]&LFSRcolor0[483]);
    BiasedRNG[142] = (LFSRcolor0[322]&LFSRcolor0[413]&LFSRcolor0[518]);
    BiasedRNG[143] = (LFSRcolor0[543]&LFSRcolor0[574]&LFSRcolor0[118]);
    BiasedRNG[144] = (LFSRcolor0[24]&LFSRcolor0[22]&LFSRcolor0[106]);
    BiasedRNG[145] = (LFSRcolor0[25]&LFSRcolor0[230]&LFSRcolor0[266]);
    BiasedRNG[146] = (LFSRcolor0[32]&LFSRcolor0[220]&LFSRcolor0[593]);
    BiasedRNG[147] = (LFSRcolor0[215]&LFSRcolor0[397]&LFSRcolor0[144]);
    BiasedRNG[148] = (LFSRcolor0[427]&LFSRcolor0[636]&LFSRcolor0[355]);
    BiasedRNG[149] = (LFSRcolor0[504]&LFSRcolor0[507]&LFSRcolor0[532]);
    BiasedRNG[150] = (LFSRcolor0[433]&LFSRcolor0[554]&LFSRcolor0[535]);
    BiasedRNG[151] = (LFSRcolor0[633]&LFSRcolor0[326]&LFSRcolor0[39]);
    BiasedRNG[152] = (LFSRcolor0[599]&LFSRcolor0[392]&LFSRcolor0[615]);
    BiasedRNG[153] = (LFSRcolor0[463]&LFSRcolor0[308]&LFSRcolor0[127]);
    BiasedRNG[154] = (LFSRcolor0[441]&LFSRcolor0[101]&LFSRcolor0[188]);
    BiasedRNG[155] = (LFSRcolor0[108]&LFSRcolor0[373]&LFSRcolor0[374]);
    BiasedRNG[156] = (LFSRcolor0[143]&LFSRcolor0[70]&LFSRcolor0[9]);
    BiasedRNG[157] = (LFSRcolor0[233]&LFSRcolor0[564]&LFSRcolor0[202]);
    BiasedRNG[158] = (LFSRcolor0[477]&LFSRcolor0[76]&LFSRcolor0[620]);
    BiasedRNG[159] = (LFSRcolor0[448]&LFSRcolor0[598]&LFSRcolor0[595]);
    BiasedRNG[160] = (LFSRcolor0[154]&LFSRcolor0[52]&LFSRcolor0[531]);
    BiasedRNG[161] = (LFSRcolor0[643]&LFSRcolor0[192]&LFSRcolor0[349]);
    BiasedRNG[162] = (LFSRcolor0[13]&LFSRcolor0[345]&LFSRcolor0[584]);
    BiasedRNG[163] = (LFSRcolor0[229]&LFSRcolor0[263]&LFSRcolor0[14]);
    BiasedRNG[164] = (LFSRcolor0[209]&LFSRcolor0[103]&LFSRcolor0[568]);
    BiasedRNG[165] = (LFSRcolor0[31]&LFSRcolor0[47]&LFSRcolor0[391]);
    BiasedRNG[166] = (LFSRcolor0[503]&LFSRcolor0[129]&LFSRcolor0[95]);
    BiasedRNG[167] = (LFSRcolor0[33]&LFSRcolor0[569]&LFSRcolor0[210]);
    UnbiasedRNG[0] = LFSRcolor0[113];
    UnbiasedRNG[1] = LFSRcolor0[125];
    UnbiasedRNG[2] = LFSRcolor0[55];
    UnbiasedRNG[3] = LFSRcolor0[213];
    UnbiasedRNG[4] = LFSRcolor0[264];
    UnbiasedRNG[5] = LFSRcolor0[490];
    UnbiasedRNG[6] = LFSRcolor0[86];
    UnbiasedRNG[7] = LFSRcolor0[378];
    UnbiasedRNG[8] = LFSRcolor0[280];
    UnbiasedRNG[9] = LFSRcolor0[444];
    UnbiasedRNG[10] = LFSRcolor0[382];
    UnbiasedRNG[11] = LFSRcolor0[606];
    UnbiasedRNG[12] = LFSRcolor0[439];
    UnbiasedRNG[13] = LFSRcolor0[120];
    UnbiasedRNG[14] = LFSRcolor0[93];
    UnbiasedRNG[15] = LFSRcolor0[126];
    UnbiasedRNG[16] = LFSRcolor0[87];
    UnbiasedRNG[17] = LFSRcolor0[471];
    UnbiasedRNG[18] = LFSRcolor0[296];
    UnbiasedRNG[19] = LFSRcolor0[180];
    UnbiasedRNG[20] = LFSRcolor0[319];
    UnbiasedRNG[21] = LFSRcolor0[555];
    UnbiasedRNG[22] = LFSRcolor0[297];
    UnbiasedRNG[23] = LFSRcolor0[499];
    UnbiasedRNG[24] = LFSRcolor0[315];
    UnbiasedRNG[25] = LFSRcolor0[393];
    UnbiasedRNG[26] = LFSRcolor0[83];
    UnbiasedRNG[27] = LFSRcolor0[179];
    UnbiasedRNG[28] = LFSRcolor0[521];
    UnbiasedRNG[29] = LFSRcolor0[200];
    UnbiasedRNG[30] = LFSRcolor0[610];
    UnbiasedRNG[31] = LFSRcolor0[175];
    UnbiasedRNG[32] = LFSRcolor0[16];
    UnbiasedRNG[33] = LFSRcolor0[283];
    UnbiasedRNG[34] = LFSRcolor0[600];
    UnbiasedRNG[35] = LFSRcolor0[11];
    UnbiasedRNG[36] = LFSRcolor0[581];
    UnbiasedRNG[37] = LFSRcolor0[478];
    UnbiasedRNG[38] = LFSRcolor0[177];
    UnbiasedRNG[39] = LFSRcolor0[351];
    UnbiasedRNG[40] = LFSRcolor0[479];
    UnbiasedRNG[41] = LFSRcolor0[287];
    UnbiasedRNG[42] = LFSRcolor0[79];
    UnbiasedRNG[43] = LFSRcolor0[164];
    UnbiasedRNG[44] = LFSRcolor0[612];
    UnbiasedRNG[45] = LFSRcolor0[248];
    UnbiasedRNG[46] = LFSRcolor0[135];
    UnbiasedRNG[47] = LFSRcolor0[488];
    UnbiasedRNG[48] = LFSRcolor0[53];
    UnbiasedRNG[49] = LFSRcolor0[497];
    UnbiasedRNG[50] = LFSRcolor0[641];
    UnbiasedRNG[51] = LFSRcolor0[461];
    UnbiasedRNG[52] = LFSRcolor0[422];
    UnbiasedRNG[53] = LFSRcolor0[309];
    UnbiasedRNG[54] = LFSRcolor0[457];
    UnbiasedRNG[55] = LFSRcolor0[623];
    UnbiasedRNG[56] = LFSRcolor0[466];
    UnbiasedRNG[57] = LFSRcolor0[148];
    UnbiasedRNG[58] = LFSRcolor0[284];
    UnbiasedRNG[59] = LFSRcolor0[254];
    UnbiasedRNG[60] = LFSRcolor0[314];
    UnbiasedRNG[61] = LFSRcolor0[301];
    UnbiasedRNG[62] = LFSRcolor0[281];
    UnbiasedRNG[63] = LFSRcolor0[51];
    UnbiasedRNG[64] = LFSRcolor0[146];
    UnbiasedRNG[65] = LFSRcolor0[198];
    UnbiasedRNG[66] = LFSRcolor0[390];
    UnbiasedRNG[67] = LFSRcolor0[509];
    UnbiasedRNG[68] = LFSRcolor0[165];
    UnbiasedRNG[69] = LFSRcolor0[71];
    UnbiasedRNG[70] = LFSRcolor0[75];
    UnbiasedRNG[71] = LFSRcolor0[632];
    UnbiasedRNG[72] = LFSRcolor0[196];
    UnbiasedRNG[73] = LFSRcolor0[440];
    UnbiasedRNG[74] = LFSRcolor0[447];
    UnbiasedRNG[75] = LFSRcolor0[347];
    UnbiasedRNG[76] = LFSRcolor0[26];
    UnbiasedRNG[77] = LFSRcolor0[458];
    UnbiasedRNG[78] = LFSRcolor0[41];
    UnbiasedRNG[79] = LFSRcolor0[592];
    UnbiasedRNG[80] = LFSRcolor0[199];
    UnbiasedRNG[81] = LFSRcolor0[540];
    UnbiasedRNG[82] = LFSRcolor0[152];
    UnbiasedRNG[83] = LFSRcolor0[614];
    UnbiasedRNG[84] = LFSRcolor0[253];
    UnbiasedRNG[85] = LFSRcolor0[10];
    UnbiasedRNG[86] = LFSRcolor0[442];
    UnbiasedRNG[87] = LFSRcolor0[348];
    UnbiasedRNG[88] = LFSRcolor0[371];
    UnbiasedRNG[89] = LFSRcolor0[575];
    UnbiasedRNG[90] = LFSRcolor0[625];
    UnbiasedRNG[91] = LFSRcolor0[418];
    UnbiasedRNG[92] = LFSRcolor0[533];
    UnbiasedRNG[93] = LFSRcolor0[325];
    UnbiasedRNG[94] = LFSRcolor0[408];
    UnbiasedRNG[95] = LFSRcolor0[12];
    UnbiasedRNG[96] = LFSRcolor0[406];
    UnbiasedRNG[97] = LFSRcolor0[181];
    UnbiasedRNG[98] = LFSRcolor0[121];
    UnbiasedRNG[99] = LFSRcolor0[286];
    UnbiasedRNG[100] = LFSRcolor0[634];
    UnbiasedRNG[101] = LFSRcolor0[530];
    UnbiasedRNG[102] = LFSRcolor0[428];
    UnbiasedRNG[103] = LFSRcolor0[84];
    UnbiasedRNG[104] = LFSRcolor0[368];
    UnbiasedRNG[105] = LFSRcolor0[178];
    UnbiasedRNG[106] = LFSRcolor0[639];
    UnbiasedRNG[107] = LFSRcolor0[147];
    UnbiasedRNG[108] = LFSRcolor0[306];
    UnbiasedRNG[109] = LFSRcolor0[258];
    UnbiasedRNG[110] = LFSRcolor0[622];
    UnbiasedRNG[111] = LFSRcolor0[476];
    UnbiasedRNG[112] = LFSRcolor0[162];
    UnbiasedRNG[113] = LFSRcolor0[243];
    UnbiasedRNG[114] = LFSRcolor0[183];
    UnbiasedRNG[115] = LFSRcolor0[246];
    UnbiasedRNG[116] = LFSRcolor0[158];
    UnbiasedRNG[117] = LFSRcolor0[454];
    UnbiasedRNG[118] = LFSRcolor0[37];
    UnbiasedRNG[119] = LFSRcolor0[173];
    UnbiasedRNG[120] = LFSRcolor0[330];
    UnbiasedRNG[121] = LFSRcolor0[494];
    UnbiasedRNG[122] = LFSRcolor0[244];
    UnbiasedRNG[123] = LFSRcolor0[311];
    UnbiasedRNG[124] = LFSRcolor0[114];
    UnbiasedRNG[125] = LFSRcolor0[104];
    UnbiasedRNG[126] = LFSRcolor0[452];
    UnbiasedRNG[127] = LFSRcolor0[156];
    UnbiasedRNG[128] = LFSRcolor0[586];
    UnbiasedRNG[129] = LFSRcolor0[107];
    UnbiasedRNG[130] = LFSRcolor0[335];
end

always @(posedge color0_clk) begin
    BiasedRNG[168] = (LFSRcolor1[503]&LFSRcolor1[545]&LFSRcolor1[762]);
    BiasedRNG[169] = (LFSRcolor1[675]&LFSRcolor1[103]&LFSRcolor1[42]);
    BiasedRNG[170] = (LFSRcolor1[370]&LFSRcolor1[36]&LFSRcolor1[653]);
    BiasedRNG[171] = (LFSRcolor1[289]&LFSRcolor1[62]&LFSRcolor1[747]);
    BiasedRNG[172] = (LFSRcolor1[296]&LFSRcolor1[603]&LFSRcolor1[219]);
    BiasedRNG[173] = (LFSRcolor1[70]&LFSRcolor1[418]&LFSRcolor1[487]);
    BiasedRNG[174] = (LFSRcolor1[215]&LFSRcolor1[224]&LFSRcolor1[507]);
    BiasedRNG[175] = (LFSRcolor1[148]&LFSRcolor1[302]&LFSRcolor1[321]);
    BiasedRNG[176] = (LFSRcolor1[447]&LFSRcolor1[22]&LFSRcolor1[65]);
    BiasedRNG[177] = (LFSRcolor1[526]&LFSRcolor1[268]&LFSRcolor1[43]);
    BiasedRNG[178] = (LFSRcolor1[244]&LFSRcolor1[615]&LFSRcolor1[543]);
    BiasedRNG[179] = (LFSRcolor1[27]&LFSRcolor1[635]&LFSRcolor1[195]);
    BiasedRNG[180] = (LFSRcolor1[368]&LFSRcolor1[79]&LFSRcolor1[452]);
    BiasedRNG[181] = (LFSRcolor1[456]&LFSRcolor1[40]&LFSRcolor1[620]);
    BiasedRNG[182] = (LFSRcolor1[254]&LFSRcolor1[176]&LFSRcolor1[274]);
    BiasedRNG[183] = (LFSRcolor1[598]&LFSRcolor1[749]&LFSRcolor1[280]);
    BiasedRNG[184] = (LFSRcolor1[484]&LFSRcolor1[674]&LFSRcolor1[396]);
    BiasedRNG[185] = (LFSRcolor1[333]&LFSRcolor1[765]&LFSRcolor1[137]);
    BiasedRNG[186] = (LFSRcolor1[4]&LFSRcolor1[21]&LFSRcolor1[400]);
    BiasedRNG[187] = (LFSRcolor1[681]&LFSRcolor1[694]&LFSRcolor1[56]);
    BiasedRNG[188] = (LFSRcolor1[455]&LFSRcolor1[386]&LFSRcolor1[23]);
    BiasedRNG[189] = (LFSRcolor1[351]&LFSRcolor1[668]&LFSRcolor1[637]);
    BiasedRNG[190] = (LFSRcolor1[573]&LFSRcolor1[322]&LFSRcolor1[652]);
    BiasedRNG[191] = (LFSRcolor1[555]&LFSRcolor1[240]&LFSRcolor1[531]);
    BiasedRNG[192] = (LFSRcolor1[290]&LFSRcolor1[771]&LFSRcolor1[593]);
    BiasedRNG[193] = (LFSRcolor1[232]&LFSRcolor1[724]&LFSRcolor1[63]);
    BiasedRNG[194] = (LFSRcolor1[489]&LFSRcolor1[314]&LFSRcolor1[661]);
    BiasedRNG[195] = (LFSRcolor1[374]&LFSRcolor1[752]&LFSRcolor1[291]);
    BiasedRNG[196] = (LFSRcolor1[435]&LFSRcolor1[6]&LFSRcolor1[679]);
    BiasedRNG[197] = (LFSRcolor1[494]&LFSRcolor1[278]&LFSRcolor1[380]);
    BiasedRNG[198] = (LFSRcolor1[379]&LFSRcolor1[376]&LFSRcolor1[569]);
    BiasedRNG[199] = (LFSRcolor1[336]&LFSRcolor1[721]&LFSRcolor1[537]);
    BiasedRNG[200] = (LFSRcolor1[535]&LFSRcolor1[756]&LFSRcolor1[209]);
    BiasedRNG[201] = (LFSRcolor1[742]&LFSRcolor1[504]&LFSRcolor1[389]);
    BiasedRNG[202] = (LFSRcolor1[92]&LFSRcolor1[115]&LFSRcolor1[57]);
    BiasedRNG[203] = (LFSRcolor1[364]&LFSRcolor1[478]&LFSRcolor1[217]);
    BiasedRNG[204] = (LFSRcolor1[483]&LFSRcolor1[331]&LFSRcolor1[301]);
    BiasedRNG[205] = (LFSRcolor1[18]&LFSRcolor1[127]&LFSRcolor1[411]);
    BiasedRNG[206] = (LFSRcolor1[399]&LFSRcolor1[517]&LFSRcolor1[521]);
    BiasedRNG[207] = (LFSRcolor1[665]&LFSRcolor1[764]&LFSRcolor1[621]);
    BiasedRNG[208] = (LFSRcolor1[99]&LFSRcolor1[260]&LFSRcolor1[464]);
    BiasedRNG[209] = (LFSRcolor1[446]&LFSRcolor1[574]&LFSRcolor1[472]);
    BiasedRNG[210] = (LFSRcolor1[473]&LFSRcolor1[168]&LFSRcolor1[48]);
    BiasedRNG[211] = (LFSRcolor1[760]&LFSRcolor1[619]&LFSRcolor1[408]);
    BiasedRNG[212] = (LFSRcolor1[305]&LFSRcolor1[711]&LFSRcolor1[470]);
    BiasedRNG[213] = (LFSRcolor1[710]&LFSRcolor1[167]&LFSRcolor1[343]);
    BiasedRNG[214] = (LFSRcolor1[757]&LFSRcolor1[94]&LFSRcolor1[709]);
    BiasedRNG[215] = (LFSRcolor1[107]&LFSRcolor1[361]&LFSRcolor1[753]);
    BiasedRNG[216] = (LFSRcolor1[394]&LFSRcolor1[235]&LFSRcolor1[706]);
    BiasedRNG[217] = (LFSRcolor1[726]&LFSRcolor1[363]&LFSRcolor1[193]);
    BiasedRNG[218] = (LFSRcolor1[310]&LFSRcolor1[371]&LFSRcolor1[3]);
    BiasedRNG[219] = (LFSRcolor1[85]&LFSRcolor1[142]&LFSRcolor1[689]);
    BiasedRNG[220] = (LFSRcolor1[247]&LFSRcolor1[281]&LFSRcolor1[414]);
    BiasedRNG[221] = (LFSRcolor1[469]&LFSRcolor1[166]&LFSRcolor1[84]);
    BiasedRNG[222] = (LFSRcolor1[300]&LFSRcolor1[73]&LFSRcolor1[471]);
    BiasedRNG[223] = (LFSRcolor1[236]&LFSRcolor1[673]&LFSRcolor1[69]);
    BiasedRNG[224] = (LFSRcolor1[434]&LFSRcolor1[377]&LFSRcolor1[781]);
    BiasedRNG[225] = (LFSRcolor1[499]&LFSRcolor1[248]&LFSRcolor1[382]);
    BiasedRNG[226] = (LFSRcolor1[658]&LFSRcolor1[387]&LFSRcolor1[493]);
    BiasedRNG[227] = (LFSRcolor1[568]&LFSRcolor1[67]&LFSRcolor1[185]);
    BiasedRNG[228] = (LFSRcolor1[39]&LFSRcolor1[746]&LFSRcolor1[457]);
    BiasedRNG[229] = (LFSRcolor1[147]&LFSRcolor1[202]&LFSRcolor1[32]);
    BiasedRNG[230] = (LFSRcolor1[221]&LFSRcolor1[163]&LFSRcolor1[252]);
    BiasedRNG[231] = (LFSRcolor1[258]&LFSRcolor1[425]&LFSRcolor1[663]);
    BiasedRNG[232] = (LFSRcolor1[579]&LFSRcolor1[479]&LFSRcolor1[566]);
    BiasedRNG[233] = (LFSRcolor1[359]&LFSRcolor1[450]&LFSRcolor1[727]);
    BiasedRNG[234] = (LFSRcolor1[256]&LFSRcolor1[66]&LFSRcolor1[656]);
    BiasedRNG[235] = (LFSRcolor1[372]&LFSRcolor1[459]&LFSRcolor1[397]);
    BiasedRNG[236] = (LFSRcolor1[439]&LFSRcolor1[309]&LFSRcolor1[345]);
    BiasedRNG[237] = (LFSRcolor1[218]&LFSRcolor1[667]&LFSRcolor1[522]);
    BiasedRNG[238] = (LFSRcolor1[24]&LFSRcolor1[182]&LFSRcolor1[592]);
    BiasedRNG[239] = (LFSRcolor1[304]&LFSRcolor1[261]&LFSRcolor1[743]);
    BiasedRNG[240] = (LFSRcolor1[45]&LFSRcolor1[768]&LFSRcolor1[208]);
    BiasedRNG[241] = (LFSRcolor1[740]&LFSRcolor1[773]&LFSRcolor1[154]);
    BiasedRNG[242] = (LFSRcolor1[31]&LFSRcolor1[750]&LFSRcolor1[64]);
    BiasedRNG[243] = (LFSRcolor1[775]&LFSRcolor1[170]&LFSRcolor1[365]);
    BiasedRNG[244] = (LFSRcolor1[245]&LFSRcolor1[482]&LFSRcolor1[583]);
    BiasedRNG[245] = (LFSRcolor1[687]&LFSRcolor1[87]&LFSRcolor1[181]);
    BiasedRNG[246] = (LFSRcolor1[676]&LFSRcolor1[572]&LFSRcolor1[72]);
    BiasedRNG[247] = (LFSRcolor1[431]&LFSRcolor1[755]&LFSRcolor1[356]);
    BiasedRNG[248] = (LFSRcolor1[428]&LFSRcolor1[284]&LFSRcolor1[91]);
    BiasedRNG[249] = (LFSRcolor1[201]&LFSRcolor1[59]&LFSRcolor1[12]);
    BiasedRNG[250] = (LFSRcolor1[46]&LFSRcolor1[50]&LFSRcolor1[13]);
    BiasedRNG[251] = (LFSRcolor1[509]&LFSRcolor1[714]&LFSRcolor1[298]);
    BiasedRNG[252] = (LFSRcolor1[184]&LFSRcolor1[602]&LFSRcolor1[442]);
    BiasedRNG[253] = (LFSRcolor1[15]&LFSRcolor1[308]&LFSRcolor1[594]);
    BiasedRNG[254] = (LFSRcolor1[530]&LFSRcolor1[536]&LFSRcolor1[349]);
    BiasedRNG[255] = (LFSRcolor1[651]&LFSRcolor1[596]&LFSRcolor1[454]);
    BiasedRNG[256] = (LFSRcolor1[383]&LFSRcolor1[180]&LFSRcolor1[644]);
    BiasedRNG[257] = (LFSRcolor1[662]&LFSRcolor1[229]&LFSRcolor1[0]);
    BiasedRNG[258] = (LFSRcolor1[645]&LFSRcolor1[608]&LFSRcolor1[725]);
    BiasedRNG[259] = (LFSRcolor1[553]&LFSRcolor1[360]&LFSRcolor1[265]);
    BiasedRNG[260] = (LFSRcolor1[285]&LFSRcolor1[134]&LFSRcolor1[119]);
    BiasedRNG[261] = (LFSRcolor1[41]&LFSRcolor1[563]&LFSRcolor1[664]);
    BiasedRNG[262] = (LFSRcolor1[337]&LFSRcolor1[82]&LFSRcolor1[582]);
    BiasedRNG[263] = (LFSRcolor1[388]&LFSRcolor1[696]&LFSRcolor1[506]);
    BiasedRNG[264] = (LFSRcolor1[95]&LFSRcolor1[691]&LFSRcolor1[423]);
    BiasedRNG[265] = (LFSRcolor1[160]&LFSRcolor1[595]&LFSRcolor1[677]);
    BiasedRNG[266] = (LFSRcolor1[540]&LFSRcolor1[173]&LFSRcolor1[684]);
    BiasedRNG[267] = (LFSRcolor1[720]&LFSRcolor1[548]&LFSRcolor1[267]);
    BiasedRNG[268] = (LFSRcolor1[477]&LFSRcolor1[632]&LFSRcolor1[420]);
    BiasedRNG[269] = (LFSRcolor1[636]&LFSRcolor1[307]&LFSRcolor1[678]);
    BiasedRNG[270] = (LFSRcolor1[451]&LFSRcolor1[323]&LFSRcolor1[212]);
    BiasedRNG[271] = (LFSRcolor1[395]&LFSRcolor1[144]&LFSRcolor1[549]);
    BiasedRNG[272] = (LFSRcolor1[682]&LFSRcolor1[524]&LFSRcolor1[106]);
    BiasedRNG[273] = (LFSRcolor1[161]&LFSRcolor1[200]&LFSRcolor1[419]);
    BiasedRNG[274] = (LFSRcolor1[199]&LFSRcolor1[624]&LFSRcolor1[225]);
    BiasedRNG[275] = (LFSRcolor1[10]&LFSRcolor1[463]&LFSRcolor1[384]);
    BiasedRNG[276] = (LFSRcolor1[444]&LFSRcolor1[700]&LFSRcolor1[528]);
    BiasedRNG[277] = (LFSRcolor1[179]&LFSRcolor1[55]&LFSRcolor1[295]);
    BiasedRNG[278] = (LFSRcolor1[178]&LFSRcolor1[288]&LFSRcolor1[342]);
    BiasedRNG[279] = (LFSRcolor1[138]&LFSRcolor1[97]&LFSRcolor1[74]);
    BiasedRNG[280] = (LFSRcolor1[120]&LFSRcolor1[312]&LFSRcolor1[37]);
    BiasedRNG[281] = (LFSRcolor1[354]&LFSRcolor1[17]&LFSRcolor1[601]);
    BiasedRNG[282] = (LFSRcolor1[758]&LFSRcolor1[695]&LFSRcolor1[557]);
    BiasedRNG[283] = (LFSRcolor1[575]&LFSRcolor1[177]&LFSRcolor1[640]);
    BiasedRNG[284] = (LFSRcolor1[410]&LFSRcolor1[516]&LFSRcolor1[567]);
    BiasedRNG[285] = (LFSRcolor1[329]&LFSRcolor1[81]&LFSRcolor1[242]);
    BiasedRNG[286] = (LFSRcolor1[352]&LFSRcolor1[745]&LFSRcolor1[718]);
    BiasedRNG[287] = (LFSRcolor1[259]&LFSRcolor1[722]&LFSRcolor1[649]);
    BiasedRNG[288] = (LFSRcolor1[117]&LFSRcolor1[172]&LFSRcolor1[80]);
    BiasedRNG[289] = (LFSRcolor1[654]&LFSRcolor1[49]&LFSRcolor1[7]);
    BiasedRNG[290] = (LFSRcolor1[779]&LFSRcolor1[707]&LFSRcolor1[311]);
    BiasedRNG[291] = (LFSRcolor1[449]&LFSRcolor1[693]&LFSRcolor1[600]);
    BiasedRNG[292] = (LFSRcolor1[585]&LFSRcolor1[544]&LFSRcolor1[239]);
    BiasedRNG[293] = (LFSRcolor1[9]&LFSRcolor1[381]&LFSRcolor1[589]);
    BiasedRNG[294] = (LFSRcolor1[96]&LFSRcolor1[194]&LFSRcolor1[58]);
    BiasedRNG[295] = (LFSRcolor1[539]&LFSRcolor1[191]&LFSRcolor1[560]);
    BiasedRNG[296] = (LFSRcolor1[581]&LFSRcolor1[458]&LFSRcolor1[401]);
    BiasedRNG[297] = (LFSRcolor1[273]&LFSRcolor1[53]&LFSRcolor1[228]);
    BiasedRNG[298] = (LFSRcolor1[44]&LFSRcolor1[576]&LFSRcolor1[324]);
    BiasedRNG[299] = (LFSRcolor1[216]&LFSRcolor1[634]&LFSRcolor1[130]);
    BiasedRNG[300] = (LFSRcolor1[210]&LFSRcolor1[139]&LFSRcolor1[437]);
    BiasedRNG[301] = (LFSRcolor1[362]&LFSRcolor1[606]&LFSRcolor1[222]);
    BiasedRNG[302] = (LFSRcolor1[61]&LFSRcolor1[378]&LFSRcolor1[475]);
    BiasedRNG[303] = (LFSRcolor1[488]&LFSRcolor1[466]&LFSRcolor1[169]);
    BiasedRNG[304] = (LFSRcolor1[223]&LFSRcolor1[297]&LFSRcolor1[703]);
    BiasedRNG[305] = (LFSRcolor1[481]&LFSRcolor1[164]&LFSRcolor1[93]);
    BiasedRNG[306] = (LFSRcolor1[629]&LFSRcolor1[373]&LFSRcolor1[186]);
    BiasedRNG[307] = (LFSRcolor1[86]&LFSRcolor1[625]&LFSRcolor1[460]);
    BiasedRNG[308] = (LFSRcolor1[554]&LFSRcolor1[511]&LFSRcolor1[33]);
    BiasedRNG[309] = (LFSRcolor1[510]&LFSRcolor1[730]&LFSRcolor1[776]);
    BiasedRNG[310] = (LFSRcolor1[319]&LFSRcolor1[605]&LFSRcolor1[146]);
    BiasedRNG[311] = (LFSRcolor1[88]&LFSRcolor1[465]&LFSRcolor1[697]);
    BiasedRNG[312] = (LFSRcolor1[716]&LFSRcolor1[112]&LFSRcolor1[541]);
    BiasedRNG[313] = (LFSRcolor1[417]&LFSRcolor1[647]&LFSRcolor1[20]);
    BiasedRNG[314] = (LFSRcolor1[198]&LFSRcolor1[123]&LFSRcolor1[686]);
    BiasedRNG[315] = (LFSRcolor1[630]&LFSRcolor1[264]&LFSRcolor1[767]);
    BiasedRNG[316] = (LFSRcolor1[231]&LFSRcolor1[28]&LFSRcolor1[570]);
    BiasedRNG[317] = (LFSRcolor1[512]&LFSRcolor1[559]&LFSRcolor1[590]);
    BiasedRNG[318] = (LFSRcolor1[206]&LFSRcolor1[344]&LFSRcolor1[175]);
    BiasedRNG[319] = (LFSRcolor1[338]&LFSRcolor1[214]&LFSRcolor1[739]);
    BiasedRNG[320] = (LFSRcolor1[213]&LFSRcolor1[398]&LFSRcolor1[149]);
    BiasedRNG[321] = (LFSRcolor1[83]&LFSRcolor1[628]&LFSRcolor1[550]);
    BiasedRNG[322] = (LFSRcolor1[76]&LFSRcolor1[108]&LFSRcolor1[405]);
    BiasedRNG[323] = (LFSRcolor1[627]&LFSRcolor1[436]&LFSRcolor1[111]);
    BiasedRNG[324] = (LFSRcolor1[2]&LFSRcolor1[403]&LFSRcolor1[617]);
    BiasedRNG[325] = (LFSRcolor1[586]&LFSRcolor1[287]&LFSRcolor1[286]);
    BiasedRNG[326] = (LFSRcolor1[205]&LFSRcolor1[580]&LFSRcolor1[604]);
    BiasedRNG[327] = (LFSRcolor1[547]&LFSRcolor1[326]&LFSRcolor1[705]);
    BiasedRNG[328] = (LFSRcolor1[375]&LFSRcolor1[334]&LFSRcolor1[292]);
    BiasedRNG[329] = (LFSRcolor1[132]&LFSRcolor1[335]&LFSRcolor1[688]);
    BiasedRNG[330] = (LFSRcolor1[421]&LFSRcolor1[279]&LFSRcolor1[52]);
    BiasedRNG[331] = (LFSRcolor1[116]&LFSRcolor1[114]&LFSRcolor1[751]);
    BiasedRNG[332] = (LFSRcolor1[129]&LFSRcolor1[690]&LFSRcolor1[683]);
    BiasedRNG[333] = (LFSRcolor1[234]&LFSRcolor1[29]&LFSRcolor1[250]);
    BiasedRNG[334] = (LFSRcolor1[272]&LFSRcolor1[54]&LFSRcolor1[719]);
    BiasedRNG[335] = (LFSRcolor1[538]&LFSRcolor1[599]&LFSRcolor1[584]);
    BiasedRNG[336] = (LFSRcolor1[480]&LFSRcolor1[341]&LFSRcolor1[348]);
    BiasedRNG[337] = (LFSRcolor1[51]&LFSRcolor1[171]&LFSRcolor1[270]);
    BiasedRNG[338] = (LFSRcolor1[155]&LFSRcolor1[492]&LFSRcolor1[699]);
    BiasedRNG[339] = (LFSRcolor1[476]&LFSRcolor1[672]&LFSRcolor1[769]);
    BiasedRNG[340] = (LFSRcolor1[277]&LFSRcolor1[571]&LFSRcolor1[197]);
    BiasedRNG[341] = (LFSRcolor1[622]&LFSRcolor1[692]&LFSRcolor1[441]);
    BiasedRNG[342] = (LFSRcolor1[728]&LFSRcolor1[358]&LFSRcolor1[497]);
    BiasedRNG[343] = (LFSRcolor1[233]&LFSRcolor1[597]&LFSRcolor1[612]);
    BiasedRNG[344] = (LFSRcolor1[8]&LFSRcolor1[520]&LFSRcolor1[502]);
    BiasedRNG[345] = (LFSRcolor1[350]&LFSRcolor1[430]&LFSRcolor1[429]);
    BiasedRNG[346] = (LFSRcolor1[68]&LFSRcolor1[204]&LFSRcolor1[515]);
    BiasedRNG[347] = (LFSRcolor1[614]&LFSRcolor1[35]&LFSRcolor1[735]);
    BiasedRNG[348] = (LFSRcolor1[152]&LFSRcolor1[122]&LFSRcolor1[102]);
    BiasedRNG[349] = (LFSRcolor1[145]&LFSRcolor1[761]&LFSRcolor1[527]);
    BiasedRNG[350] = (LFSRcolor1[157]&LFSRcolor1[607]&LFSRcolor1[263]);
    BiasedRNG[351] = (LFSRcolor1[158]&LFSRcolor1[670]&LFSRcolor1[525]);
    BiasedRNG[352] = (LFSRcolor1[467]&LFSRcolor1[211]&LFSRcolor1[468]);
    BiasedRNG[353] = (LFSRcolor1[412]&LFSRcolor1[445]&LFSRcolor1[490]);
    BiasedRNG[354] = (LFSRcolor1[110]&LFSRcolor1[650]&LFSRcolor1[415]);
    BiasedRNG[355] = (LFSRcolor1[558]&LFSRcolor1[657]&LFSRcolor1[514]);
    BiasedRNG[356] = (LFSRcolor1[347]&LFSRcolor1[98]&LFSRcolor1[203]);
    BiasedRNG[357] = (LFSRcolor1[534]&LFSRcolor1[262]&LFSRcolor1[546]);
    BiasedRNG[358] = (LFSRcolor1[407]&LFSRcolor1[648]&LFSRcolor1[513]);
    BiasedRNG[359] = (LFSRcolor1[402]&LFSRcolor1[780]&LFSRcolor1[519]);
    BiasedRNG[360] = (LFSRcolor1[729]&LFSRcolor1[143]&LFSRcolor1[159]);
    BiasedRNG[361] = (LFSRcolor1[255]&LFSRcolor1[60]&LFSRcolor1[551]);
    BiasedRNG[362] = (LFSRcolor1[47]&LFSRcolor1[357]&LFSRcolor1[237]);
    BiasedRNG[363] = (LFSRcolor1[611]&LFSRcolor1[121]&LFSRcolor1[778]);
    BiasedRNG[364] = (LFSRcolor1[643]&LFSRcolor1[744]&LFSRcolor1[701]);
    BiasedRNG[365] = (LFSRcolor1[128]&LFSRcolor1[30]&LFSRcolor1[646]);
    BiasedRNG[366] = (LFSRcolor1[669]&LFSRcolor1[723]&LFSRcolor1[11]);
    BiasedRNG[367] = (LFSRcolor1[704]&LFSRcolor1[409]&LFSRcolor1[390]);
    BiasedRNG[368] = (LFSRcolor1[562]&LFSRcolor1[104]&LFSRcolor1[306]);
    BiasedRNG[369] = (LFSRcolor1[238]&LFSRcolor1[257]&LFSRcolor1[89]);
    BiasedRNG[370] = (LFSRcolor1[578]&LFSRcolor1[564]&LFSRcolor1[294]);
    BiasedRNG[371] = (LFSRcolor1[367]&LFSRcolor1[426]&LFSRcolor1[346]);
    BiasedRNG[372] = (LFSRcolor1[276]&LFSRcolor1[443]&LFSRcolor1[71]);
    BiasedRNG[373] = (LFSRcolor1[282]&LFSRcolor1[325]&LFSRcolor1[698]);
    BiasedRNG[374] = (LFSRcolor1[474]&LFSRcolor1[518]&LFSRcolor1[275]);
    BiasedRNG[375] = (LFSRcolor1[486]&LFSRcolor1[253]&LFSRcolor1[220]);
    BiasedRNG[376] = (LFSRcolor1[588]&LFSRcolor1[556]&LFSRcolor1[318]);
    BiasedRNG[377] = (LFSRcolor1[135]&LFSRcolor1[741]&LFSRcolor1[101]);
    BiasedRNG[378] = (LFSRcolor1[416]&LFSRcolor1[422]&LFSRcolor1[165]);
    BiasedRNG[379] = (LFSRcolor1[623]&LFSRcolor1[616]&LFSRcolor1[183]);
    BiasedRNG[380] = (LFSRcolor1[156]&LFSRcolor1[491]&LFSRcolor1[126]);
    BiasedRNG[381] = (LFSRcolor1[702]&LFSRcolor1[495]&LFSRcolor1[385]);
    BiasedRNG[382] = (LFSRcolor1[162]&LFSRcolor1[641]&LFSRcolor1[770]);
    UnbiasedRNG[131] = LFSRcolor1[299];
    UnbiasedRNG[132] = LFSRcolor1[748];
    UnbiasedRNG[133] = LFSRcolor1[207];
    UnbiasedRNG[134] = LFSRcolor1[317];
    UnbiasedRNG[135] = LFSRcolor1[587];
    UnbiasedRNG[136] = LFSRcolor1[715];
    UnbiasedRNG[137] = LFSRcolor1[671];
    UnbiasedRNG[138] = LFSRcolor1[271];
    UnbiasedRNG[139] = LFSRcolor1[153];
    UnbiasedRNG[140] = LFSRcolor1[266];
    UnbiasedRNG[141] = LFSRcolor1[124];
    UnbiasedRNG[142] = LFSRcolor1[618];
    UnbiasedRNG[143] = LFSRcolor1[100];
    UnbiasedRNG[144] = LFSRcolor1[424];
    UnbiasedRNG[145] = LFSRcolor1[251];
    UnbiasedRNG[146] = LFSRcolor1[561];
    UnbiasedRNG[147] = LFSRcolor1[712];
    UnbiasedRNG[148] = LFSRcolor1[631];
    UnbiasedRNG[149] = LFSRcolor1[188];
    UnbiasedRNG[150] = LFSRcolor1[141];
    UnbiasedRNG[151] = LFSRcolor1[433];
    UnbiasedRNG[152] = LFSRcolor1[777];
    UnbiasedRNG[153] = LFSRcolor1[226];
    UnbiasedRNG[154] = LFSRcolor1[369];
    UnbiasedRNG[155] = LFSRcolor1[105];
    UnbiasedRNG[156] = LFSRcolor1[432];
    UnbiasedRNG[157] = LFSRcolor1[26];
    UnbiasedRNG[158] = LFSRcolor1[391];
    UnbiasedRNG[159] = LFSRcolor1[25];
    UnbiasedRNG[160] = LFSRcolor1[759];
    UnbiasedRNG[161] = LFSRcolor1[14];
    UnbiasedRNG[162] = LFSRcolor1[140];
    UnbiasedRNG[163] = LFSRcolor1[734];
    UnbiasedRNG[164] = LFSRcolor1[189];
    UnbiasedRNG[165] = LFSRcolor1[609];
    UnbiasedRNG[166] = LFSRcolor1[552];
    UnbiasedRNG[167] = LFSRcolor1[113];
    UnbiasedRNG[168] = LFSRcolor1[187];
    UnbiasedRNG[169] = LFSRcolor1[249];
    UnbiasedRNG[170] = LFSRcolor1[330];
    UnbiasedRNG[171] = LFSRcolor1[174];
    UnbiasedRNG[172] = LFSRcolor1[732];
    UnbiasedRNG[173] = LFSRcolor1[150];
    UnbiasedRNG[174] = LFSRcolor1[90];
    UnbiasedRNG[175] = LFSRcolor1[542];
    UnbiasedRNG[176] = LFSRcolor1[639];
    UnbiasedRNG[177] = LFSRcolor1[438];
    UnbiasedRNG[178] = LFSRcolor1[633];
    UnbiasedRNG[179] = LFSRcolor1[328];
    UnbiasedRNG[180] = LFSRcolor1[626];
    UnbiasedRNG[181] = LFSRcolor1[448];
    UnbiasedRNG[182] = LFSRcolor1[772];
    UnbiasedRNG[183] = LFSRcolor1[565];
    UnbiasedRNG[184] = LFSRcolor1[642];
    UnbiasedRNG[185] = LFSRcolor1[332];
    UnbiasedRNG[186] = LFSRcolor1[427];
    UnbiasedRNG[187] = LFSRcolor1[680];
    UnbiasedRNG[188] = LFSRcolor1[532];
    UnbiasedRNG[189] = LFSRcolor1[774];
    UnbiasedRNG[190] = LFSRcolor1[339];
    UnbiasedRNG[191] = LFSRcolor1[131];
    UnbiasedRNG[192] = LFSRcolor1[577];
    UnbiasedRNG[193] = LFSRcolor1[685];
    UnbiasedRNG[194] = LFSRcolor1[733];
    UnbiasedRNG[195] = LFSRcolor1[713];
    UnbiasedRNG[196] = LFSRcolor1[34];
    UnbiasedRNG[197] = LFSRcolor1[392];
    UnbiasedRNG[198] = LFSRcolor1[610];
    UnbiasedRNG[199] = LFSRcolor1[227];
    UnbiasedRNG[200] = LFSRcolor1[505];
    UnbiasedRNG[201] = LFSRcolor1[613];
    UnbiasedRNG[202] = LFSRcolor1[453];
    UnbiasedRNG[203] = LFSRcolor1[246];
    UnbiasedRNG[204] = LFSRcolor1[508];
    UnbiasedRNG[205] = LFSRcolor1[523];
    UnbiasedRNG[206] = LFSRcolor1[500];
    UnbiasedRNG[207] = LFSRcolor1[591];
    UnbiasedRNG[208] = LFSRcolor1[763];
    UnbiasedRNG[209] = LFSRcolor1[731];
    UnbiasedRNG[210] = LFSRcolor1[241];
    UnbiasedRNG[211] = LFSRcolor1[190];
    UnbiasedRNG[212] = LFSRcolor1[496];
    UnbiasedRNG[213] = LFSRcolor1[736];
    UnbiasedRNG[214] = LFSRcolor1[355];
    UnbiasedRNG[215] = LFSRcolor1[708];
    UnbiasedRNG[216] = LFSRcolor1[440];
    UnbiasedRNG[217] = LFSRcolor1[393];
    UnbiasedRNG[218] = LFSRcolor1[75];
    UnbiasedRNG[219] = LFSRcolor1[109];
    UnbiasedRNG[220] = LFSRcolor1[313];
    UnbiasedRNG[221] = LFSRcolor1[659];
    UnbiasedRNG[222] = LFSRcolor1[125];
    UnbiasedRNG[223] = LFSRcolor1[230];
    UnbiasedRNG[224] = LFSRcolor1[754];
    UnbiasedRNG[225] = LFSRcolor1[461];
    UnbiasedRNG[226] = LFSRcolor1[462];
    UnbiasedRNG[227] = LFSRcolor1[533];
    UnbiasedRNG[228] = LFSRcolor1[485];
    UnbiasedRNG[229] = LFSRcolor1[136];
    UnbiasedRNG[230] = LFSRcolor1[737];
    UnbiasedRNG[231] = LFSRcolor1[293];
    UnbiasedRNG[232] = LFSRcolor1[529];
    UnbiasedRNG[233] = LFSRcolor1[283];
    UnbiasedRNG[234] = LFSRcolor1[655];
    UnbiasedRNG[235] = LFSRcolor1[151];
    UnbiasedRNG[236] = LFSRcolor1[406];
    UnbiasedRNG[237] = LFSRcolor1[413];
    UnbiasedRNG[238] = LFSRcolor1[738];
    UnbiasedRNG[239] = LFSRcolor1[766];
    UnbiasedRNG[240] = LFSRcolor1[19];
    UnbiasedRNG[241] = LFSRcolor1[243];
    UnbiasedRNG[242] = LFSRcolor1[320];
    UnbiasedRNG[243] = LFSRcolor1[666];
    UnbiasedRNG[244] = LFSRcolor1[16];
    UnbiasedRNG[245] = LFSRcolor1[404];
    UnbiasedRNG[246] = LFSRcolor1[638];
    UnbiasedRNG[247] = LFSRcolor1[660];
    UnbiasedRNG[248] = LFSRcolor1[118];
    UnbiasedRNG[249] = LFSRcolor1[192];
    UnbiasedRNG[250] = LFSRcolor1[315];
    UnbiasedRNG[251] = LFSRcolor1[340];
end

always @(posedge color1_clk) begin
    BiasedRNG[383] = (LFSRcolor2[178]&LFSRcolor2[307]&LFSRcolor2[31]);
    BiasedRNG[384] = (LFSRcolor2[597]&LFSRcolor2[354]&LFSRcolor2[170]);
    BiasedRNG[385] = (LFSRcolor2[585]&LFSRcolor2[75]&LFSRcolor2[186]);
    BiasedRNG[386] = (LFSRcolor2[224]&LFSRcolor2[44]&LFSRcolor2[42]);
    BiasedRNG[387] = (LFSRcolor2[378]&LFSRcolor2[470]&LFSRcolor2[221]);
    BiasedRNG[388] = (LFSRcolor2[548]&LFSRcolor2[522]&LFSRcolor2[351]);
    BiasedRNG[389] = (LFSRcolor2[7]&LFSRcolor2[549]&LFSRcolor2[265]);
    BiasedRNG[390] = (LFSRcolor2[385]&LFSRcolor2[171]&LFSRcolor2[505]);
    BiasedRNG[391] = (LFSRcolor2[500]&LFSRcolor2[564]&LFSRcolor2[240]);
    BiasedRNG[392] = (LFSRcolor2[432]&LFSRcolor2[108]&LFSRcolor2[94]);
    BiasedRNG[393] = (LFSRcolor2[302]&LFSRcolor2[409]&LFSRcolor2[47]);
    BiasedRNG[394] = (LFSRcolor2[519]&LFSRcolor2[273]&LFSRcolor2[64]);
    BiasedRNG[395] = (LFSRcolor2[227]&LFSRcolor2[413]&LFSRcolor2[421]);
    BiasedRNG[396] = (LFSRcolor2[592]&LFSRcolor2[242]&LFSRcolor2[164]);
    BiasedRNG[397] = (LFSRcolor2[112]&LFSRcolor2[429]&LFSRcolor2[148]);
    BiasedRNG[398] = (LFSRcolor2[575]&LFSRcolor2[109]&LFSRcolor2[418]);
    BiasedRNG[399] = (LFSRcolor2[325]&LFSRcolor2[347]&LFSRcolor2[527]);
    BiasedRNG[400] = (LFSRcolor2[536]&LFSRcolor2[591]&LFSRcolor2[211]);
    BiasedRNG[401] = (LFSRcolor2[292]&LFSRcolor2[147]&LFSRcolor2[63]);
    BiasedRNG[402] = (LFSRcolor2[136]&LFSRcolor2[533]&LFSRcolor2[453]);
    BiasedRNG[403] = (LFSRcolor2[45]&LFSRcolor2[263]&LFSRcolor2[162]);
    BiasedRNG[404] = (LFSRcolor2[29]&LFSRcolor2[234]&LFSRcolor2[83]);
    BiasedRNG[405] = (LFSRcolor2[367]&LFSRcolor2[285]&LFSRcolor2[249]);
    BiasedRNG[406] = (LFSRcolor2[67]&LFSRcolor2[475]&LFSRcolor2[417]);
    BiasedRNG[407] = (LFSRcolor2[580]&LFSRcolor2[431]&LFSRcolor2[191]);
    BiasedRNG[408] = (LFSRcolor2[458]&LFSRcolor2[41]&LFSRcolor2[311]);
    BiasedRNG[409] = (LFSRcolor2[471]&LFSRcolor2[398]&LFSRcolor2[356]);
    BiasedRNG[410] = (LFSRcolor2[43]&LFSRcolor2[144]&LFSRcolor2[559]);
    BiasedRNG[411] = (LFSRcolor2[81]&LFSRcolor2[433]&LFSRcolor2[54]);
    BiasedRNG[412] = (LFSRcolor2[328]&LFSRcolor2[389]&LFSRcolor2[380]);
    BiasedRNG[413] = (LFSRcolor2[18]&LFSRcolor2[179]&LFSRcolor2[248]);
    BiasedRNG[414] = (LFSRcolor2[133]&LFSRcolor2[74]&LFSRcolor2[80]);
    BiasedRNG[415] = (LFSRcolor2[76]&LFSRcolor2[344]&LFSRcolor2[135]);
    BiasedRNG[416] = (LFSRcolor2[161]&LFSRcolor2[317]&LFSRcolor2[262]);
    BiasedRNG[417] = (LFSRcolor2[309]&LFSRcolor2[23]&LFSRcolor2[126]);
    BiasedRNG[418] = (LFSRcolor2[93]&LFSRcolor2[270]&LFSRcolor2[165]);
    BiasedRNG[419] = (LFSRcolor2[456]&LFSRcolor2[287]&LFSRcolor2[231]);
    BiasedRNG[420] = (LFSRcolor2[58]&LFSRcolor2[379]&LFSRcolor2[449]);
    BiasedRNG[421] = (LFSRcolor2[232]&LFSRcolor2[100]&LFSRcolor2[0]);
    BiasedRNG[422] = (LFSRcolor2[40]&LFSRcolor2[127]&LFSRcolor2[114]);
    BiasedRNG[423] = (LFSRcolor2[541]&LFSRcolor2[176]&LFSRcolor2[391]);
    BiasedRNG[424] = (LFSRcolor2[352]&LFSRcolor2[312]&LFSRcolor2[525]);
    BiasedRNG[425] = (LFSRcolor2[111]&LFSRcolor2[172]&LFSRcolor2[382]);
    BiasedRNG[426] = (LFSRcolor2[92]&LFSRcolor2[370]&LFSRcolor2[571]);
    BiasedRNG[427] = (LFSRcolor2[174]&LFSRcolor2[466]&LFSRcolor2[528]);
    BiasedRNG[428] = (LFSRcolor2[57]&LFSRcolor2[65]&LFSRcolor2[343]);
    BiasedRNG[429] = (LFSRcolor2[365]&LFSRcolor2[233]&LFSRcolor2[331]);
    BiasedRNG[430] = (LFSRcolor2[142]&LFSRcolor2[520]&LFSRcolor2[188]);
    BiasedRNG[431] = (LFSRcolor2[346]&LFSRcolor2[141]&LFSRcolor2[338]);
    BiasedRNG[432] = (LFSRcolor2[574]&LFSRcolor2[425]&LFSRcolor2[422]);
    BiasedRNG[433] = (LFSRcolor2[284]&LFSRcolor2[194]&LFSRcolor2[465]);
    BiasedRNG[434] = (LFSRcolor2[567]&LFSRcolor2[219]&LFSRcolor2[116]);
    BiasedRNG[435] = (LFSRcolor2[371]&LFSRcolor2[545]&LFSRcolor2[215]);
    BiasedRNG[436] = (LFSRcolor2[539]&LFSRcolor2[275]&LFSRcolor2[488]);
    BiasedRNG[437] = (LFSRcolor2[372]&LFSRcolor2[340]&LFSRcolor2[308]);
    BiasedRNG[438] = (LFSRcolor2[572]&LFSRcolor2[281]&LFSRcolor2[9]);
    BiasedRNG[439] = (LFSRcolor2[524]&LFSRcolor2[440]&LFSRcolor2[288]);
    BiasedRNG[440] = (LFSRcolor2[52]&LFSRcolor2[274]&LFSRcolor2[30]);
    BiasedRNG[441] = (LFSRcolor2[426]&LFSRcolor2[91]&LFSRcolor2[167]);
    BiasedRNG[442] = (LFSRcolor2[269]&LFSRcolor2[137]&LFSRcolor2[483]);
    BiasedRNG[443] = (LFSRcolor2[241]&LFSRcolor2[105]&LFSRcolor2[320]);
    BiasedRNG[444] = (LFSRcolor2[146]&LFSRcolor2[132]&LFSRcolor2[214]);
    BiasedRNG[445] = (LFSRcolor2[438]&LFSRcolor2[218]&LFSRcolor2[402]);
    BiasedRNG[446] = (LFSRcolor2[280]&LFSRcolor2[563]&LFSRcolor2[490]);
    BiasedRNG[447] = (LFSRcolor2[386]&LFSRcolor2[236]&LFSRcolor2[551]);
    BiasedRNG[448] = (LFSRcolor2[305]&LFSRcolor2[204]&LFSRcolor2[318]);
    BiasedRNG[449] = (LFSRcolor2[430]&LFSRcolor2[381]&LFSRcolor2[55]);
    BiasedRNG[450] = (LFSRcolor2[565]&LFSRcolor2[376]&LFSRcolor2[264]);
    BiasedRNG[451] = (LFSRcolor2[117]&LFSRcolor2[145]&LFSRcolor2[424]);
    BiasedRNG[452] = (LFSRcolor2[330]&LFSRcolor2[46]&LFSRcolor2[532]);
    BiasedRNG[453] = (LFSRcolor2[360]&LFSRcolor2[399]&LFSRcolor2[300]);
    BiasedRNG[454] = (LFSRcolor2[21]&LFSRcolor2[303]&LFSRcolor2[295]);
    BiasedRNG[455] = (LFSRcolor2[492]&LFSRcolor2[129]&LFSRcolor2[408]);
    BiasedRNG[456] = (LFSRcolor2[387]&LFSRcolor2[448]&LFSRcolor2[79]);
    BiasedRNG[457] = (LFSRcolor2[27]&LFSRcolor2[357]&LFSRcolor2[553]);
    BiasedRNG[458] = (LFSRcolor2[350]&LFSRcolor2[258]&LFSRcolor2[78]);
    BiasedRNG[459] = (LFSRcolor2[552]&LFSRcolor2[230]&LFSRcolor2[415]);
    BiasedRNG[460] = (LFSRcolor2[531]&LFSRcolor2[200]&LFSRcolor2[250]);
    BiasedRNG[461] = (LFSRcolor2[359]&LFSRcolor2[12]&LFSRcolor2[450]);
    BiasedRNG[462] = (LFSRcolor2[485]&LFSRcolor2[276]&LFSRcolor2[119]);
    BiasedRNG[463] = (LFSRcolor2[315]&LFSRcolor2[70]&LFSRcolor2[20]);
    BiasedRNG[464] = (LFSRcolor2[156]&LFSRcolor2[183]&LFSRcolor2[196]);
    BiasedRNG[465] = (LFSRcolor2[260]&LFSRcolor2[319]&LFSRcolor2[293]);
    BiasedRNG[466] = (LFSRcolor2[169]&LFSRcolor2[467]&LFSRcolor2[277]);
    BiasedRNG[467] = (LFSRcolor2[554]&LFSRcolor2[237]&LFSRcolor2[36]);
    BiasedRNG[468] = (LFSRcolor2[557]&LFSRcolor2[122]&LFSRcolor2[62]);
    BiasedRNG[469] = (LFSRcolor2[77]&LFSRcolor2[301]&LFSRcolor2[411]);
    BiasedRNG[470] = (LFSRcolor2[337]&LFSRcolor2[477]&LFSRcolor2[410]);
    BiasedRNG[471] = (LFSRcolor2[181]&LFSRcolor2[212]&LFSRcolor2[474]);
    BiasedRNG[472] = (LFSRcolor2[154]&LFSRcolor2[345]&LFSRcolor2[461]);
    BiasedRNG[473] = (LFSRcolor2[239]&LFSRcolor2[469]&LFSRcolor2[68]);
    BiasedRNG[474] = (LFSRcolor2[404]&LFSRcolor2[168]&LFSRcolor2[420]);
    BiasedRNG[475] = (LFSRcolor2[513]&LFSRcolor2[510]&LFSRcolor2[37]);
    BiasedRNG[476] = (LFSRcolor2[401]&LFSRcolor2[491]&LFSRcolor2[251]);
    BiasedRNG[477] = (LFSRcolor2[498]&LFSRcolor2[254]&LFSRcolor2[578]);
    BiasedRNG[478] = (LFSRcolor2[569]&LFSRcolor2[534]&LFSRcolor2[502]);
    BiasedRNG[479] = (LFSRcolor2[223]&LFSRcolor2[50]&LFSRcolor2[297]);
    BiasedRNG[480] = (LFSRcolor2[427]&LFSRcolor2[481]&LFSRcolor2[266]);
    BiasedRNG[481] = (LFSRcolor2[95]&LFSRcolor2[348]&LFSRcolor2[447]);
    BiasedRNG[482] = (LFSRcolor2[523]&LFSRcolor2[358]&LFSRcolor2[368]);
    BiasedRNG[483] = (LFSRcolor2[326]&LFSRcolor2[89]&LFSRcolor2[103]);
    BiasedRNG[484] = (LFSRcolor2[60]&LFSRcolor2[558]&LFSRcolor2[457]);
    BiasedRNG[485] = (LFSRcolor2[538]&LFSRcolor2[153]&LFSRcolor2[587]);
    BiasedRNG[486] = (LFSRcolor2[4]&LFSRcolor2[479]&LFSRcolor2[462]);
    BiasedRNG[487] = (LFSRcolor2[59]&LFSRcolor2[546]&LFSRcolor2[82]);
    BiasedRNG[488] = (LFSRcolor2[198]&LFSRcolor2[349]&LFSRcolor2[362]);
    BiasedRNG[489] = (LFSRcolor2[195]&LFSRcolor2[374]&LFSRcolor2[208]);
    BiasedRNG[490] = (LFSRcolor2[497]&LFSRcolor2[66]&LFSRcolor2[106]);
    BiasedRNG[491] = (LFSRcolor2[253]&LFSRcolor2[203]&LFSRcolor2[487]);
    BiasedRNG[492] = (LFSRcolor2[48]&LFSRcolor2[143]&LFSRcolor2[90]);
    BiasedRNG[493] = (LFSRcolor2[120]&LFSRcolor2[570]&LFSRcolor2[26]);
    BiasedRNG[494] = (LFSRcolor2[193]&LFSRcolor2[182]&LFSRcolor2[416]);
    BiasedRNG[495] = (LFSRcolor2[375]&LFSRcolor2[526]&LFSRcolor2[99]);
    BiasedRNG[496] = (LFSRcolor2[403]&LFSRcolor2[123]&LFSRcolor2[149]);
    BiasedRNG[497] = (LFSRcolor2[501]&LFSRcolor2[19]&LFSRcolor2[530]);
    BiasedRNG[498] = (LFSRcolor2[56]&LFSRcolor2[220]&LFSRcolor2[291]);
    BiasedRNG[499] = (LFSRcolor2[3]&LFSRcolor2[464]&LFSRcolor2[88]);
    BiasedRNG[500] = (LFSRcolor2[529]&LFSRcolor2[256]&LFSRcolor2[296]);
    BiasedRNG[501] = (LFSRcolor2[128]&LFSRcolor2[562]&LFSRcolor2[339]);
    BiasedRNG[502] = (LFSRcolor2[394]&LFSRcolor2[332]&LFSRcolor2[259]);
    BiasedRNG[503] = (LFSRcolor2[102]&LFSRcolor2[366]&LFSRcolor2[210]);
    BiasedRNG[504] = (LFSRcolor2[323]&LFSRcolor2[428]&LFSRcolor2[434]);
    BiasedRNG[505] = (LFSRcolor2[217]&LFSRcolor2[468]&LFSRcolor2[229]);
    BiasedRNG[506] = (LFSRcolor2[134]&LFSRcolor2[355]&LFSRcolor2[113]);
    BiasedRNG[507] = (LFSRcolor2[118]&LFSRcolor2[441]&LFSRcolor2[290]);
    BiasedRNG[508] = (LFSRcolor2[24]&LFSRcolor2[85]&LFSRcolor2[140]);
    BiasedRNG[509] = (LFSRcolor2[187]&LFSRcolor2[540]&LFSRcolor2[435]);
    BiasedRNG[510] = (LFSRcolor2[86]&LFSRcolor2[363]&LFSRcolor2[560]);
    BiasedRNG[511] = (LFSRcolor2[255]&LFSRcolor2[489]&LFSRcolor2[173]);
    BiasedRNG[512] = (LFSRcolor2[573]&LFSRcolor2[566]&LFSRcolor2[206]);
    BiasedRNG[513] = (LFSRcolor2[207]&LFSRcolor2[98]&LFSRcolor2[473]);
    BiasedRNG[514] = (LFSRcolor2[157]&LFSRcolor2[190]&LFSRcolor2[14]);
    BiasedRNG[515] = (LFSRcolor2[96]&LFSRcolor2[353]&LFSRcolor2[247]);
    BiasedRNG[516] = (LFSRcolor2[228]&LFSRcolor2[322]&LFSRcolor2[412]);
    BiasedRNG[517] = (LFSRcolor2[299]&LFSRcolor2[521]&LFSRcolor2[327]);
    BiasedRNG[518] = (LFSRcolor2[484]&LFSRcolor2[499]&LFSRcolor2[316]);
    BiasedRNG[519] = (LFSRcolor2[139]&LFSRcolor2[494]&LFSRcolor2[452]);
    BiasedRNG[520] = (LFSRcolor2[15]&LFSRcolor2[201]&LFSRcolor2[279]);
    BiasedRNG[521] = (LFSRcolor2[496]&LFSRcolor2[364]&LFSRcolor2[463]);
    BiasedRNG[522] = (LFSRcolor2[324]&LFSRcolor2[406]&LFSRcolor2[584]);
    BiasedRNG[523] = (LFSRcolor2[10]&LFSRcolor2[590]&LFSRcolor2[121]);
    BiasedRNG[524] = (LFSRcolor2[25]&LFSRcolor2[28]&LFSRcolor2[369]);
    BiasedRNG[525] = (LFSRcolor2[423]&LFSRcolor2[568]&LFSRcolor2[596]);
    BiasedRNG[526] = (LFSRcolor2[537]&LFSRcolor2[516]&LFSRcolor2[33]);
    UnbiasedRNG[252] = LFSRcolor2[373];
    UnbiasedRNG[253] = LFSRcolor2[582];
    UnbiasedRNG[254] = LFSRcolor2[53];
    UnbiasedRNG[255] = LFSRcolor2[268];
    UnbiasedRNG[256] = LFSRcolor2[226];
    UnbiasedRNG[257] = LFSRcolor2[294];
    UnbiasedRNG[258] = LFSRcolor2[511];
    UnbiasedRNG[259] = LFSRcolor2[185];
    UnbiasedRNG[260] = LFSRcolor2[125];
    UnbiasedRNG[261] = LFSRcolor2[550];
    UnbiasedRNG[262] = LFSRcolor2[444];
    UnbiasedRNG[263] = LFSRcolor2[152];
    UnbiasedRNG[264] = LFSRcolor2[437];
    UnbiasedRNG[265] = LFSRcolor2[202];
    UnbiasedRNG[266] = LFSRcolor2[71];
    UnbiasedRNG[267] = LFSRcolor2[384];
    UnbiasedRNG[268] = LFSRcolor2[333];
    UnbiasedRNG[269] = LFSRcolor2[395];
    UnbiasedRNG[270] = LFSRcolor2[514];
    UnbiasedRNG[271] = LFSRcolor2[13];
    UnbiasedRNG[272] = LFSRcolor2[51];
    UnbiasedRNG[273] = LFSRcolor2[115];
    UnbiasedRNG[274] = LFSRcolor2[138];
    UnbiasedRNG[275] = LFSRcolor2[267];
    UnbiasedRNG[276] = LFSRcolor2[11];
    UnbiasedRNG[277] = LFSRcolor2[388];
    UnbiasedRNG[278] = LFSRcolor2[298];
    UnbiasedRNG[279] = LFSRcolor2[397];
    UnbiasedRNG[280] = LFSRcolor2[446];
    UnbiasedRNG[281] = LFSRcolor2[22];
    UnbiasedRNG[282] = LFSRcolor2[213];
    UnbiasedRNG[283] = LFSRcolor2[304];
    UnbiasedRNG[284] = LFSRcolor2[205];
    UnbiasedRNG[285] = LFSRcolor2[493];
    UnbiasedRNG[286] = LFSRcolor2[595];
    UnbiasedRNG[287] = LFSRcolor2[225];
    UnbiasedRNG[288] = LFSRcolor2[306];
    UnbiasedRNG[289] = LFSRcolor2[310];
    UnbiasedRNG[290] = LFSRcolor2[506];
    UnbiasedRNG[291] = LFSRcolor2[478];
    UnbiasedRNG[292] = LFSRcolor2[289];
    UnbiasedRNG[293] = LFSRcolor2[589];
    UnbiasedRNG[294] = LFSRcolor2[110];
    UnbiasedRNG[295] = LFSRcolor2[393];
    UnbiasedRNG[296] = LFSRcolor2[577];
    UnbiasedRNG[297] = LFSRcolor2[335];
    UnbiasedRNG[298] = LFSRcolor2[257];
    UnbiasedRNG[299] = LFSRcolor2[445];
    UnbiasedRNG[300] = LFSRcolor2[158];
    UnbiasedRNG[301] = LFSRcolor2[192];
    UnbiasedRNG[302] = LFSRcolor2[2];
    UnbiasedRNG[303] = LFSRcolor2[547];
    UnbiasedRNG[304] = LFSRcolor2[377];
    UnbiasedRNG[305] = LFSRcolor2[107];
    UnbiasedRNG[306] = LFSRcolor2[459];
    UnbiasedRNG[307] = LFSRcolor2[407];
    UnbiasedRNG[308] = LFSRcolor2[49];
    UnbiasedRNG[309] = LFSRcolor2[87];
    UnbiasedRNG[310] = LFSRcolor2[283];
    UnbiasedRNG[311] = LFSRcolor2[507];
    UnbiasedRNG[312] = LFSRcolor2[454];
    UnbiasedRNG[313] = LFSRcolor2[518];
    UnbiasedRNG[314] = LFSRcolor2[517];
    UnbiasedRNG[315] = LFSRcolor2[495];
    UnbiasedRNG[316] = LFSRcolor2[189];
    UnbiasedRNG[317] = LFSRcolor2[282];
    UnbiasedRNG[318] = LFSRcolor2[512];
    UnbiasedRNG[319] = LFSRcolor2[16];
    UnbiasedRNG[320] = LFSRcolor2[34];
    UnbiasedRNG[321] = LFSRcolor2[244];
    UnbiasedRNG[322] = LFSRcolor2[396];
    UnbiasedRNG[323] = LFSRcolor2[515];
    UnbiasedRNG[324] = LFSRcolor2[361];
    UnbiasedRNG[325] = LFSRcolor2[17];
    UnbiasedRNG[326] = LFSRcolor2[439];
    UnbiasedRNG[327] = LFSRcolor2[336];
    UnbiasedRNG[328] = LFSRcolor2[150];
    UnbiasedRNG[329] = LFSRcolor2[593];
    UnbiasedRNG[330] = LFSRcolor2[101];
    UnbiasedRNG[331] = LFSRcolor2[32];
    UnbiasedRNG[332] = LFSRcolor2[97];
    UnbiasedRNG[333] = LFSRcolor2[392];
    UnbiasedRNG[334] = LFSRcolor2[443];
    UnbiasedRNG[335] = LFSRcolor2[535];
    UnbiasedRNG[336] = LFSRcolor2[73];
    UnbiasedRNG[337] = LFSRcolor2[271];
    UnbiasedRNG[338] = LFSRcolor2[480];
    UnbiasedRNG[339] = LFSRcolor2[543];
    UnbiasedRNG[340] = LFSRcolor2[199];
    UnbiasedRNG[341] = LFSRcolor2[278];
    UnbiasedRNG[342] = LFSRcolor2[180];
    UnbiasedRNG[343] = LFSRcolor2[246];
    UnbiasedRNG[344] = LFSRcolor2[476];
    UnbiasedRNG[345] = LFSRcolor2[6];
    UnbiasedRNG[346] = LFSRcolor2[166];
    UnbiasedRNG[347] = LFSRcolor2[272];
    UnbiasedRNG[348] = LFSRcolor2[130];
    UnbiasedRNG[349] = LFSRcolor2[8];
    UnbiasedRNG[350] = LFSRcolor2[261];
    UnbiasedRNG[351] = LFSRcolor2[390];
    UnbiasedRNG[352] = LFSRcolor2[104];
    UnbiasedRNG[353] = LFSRcolor2[243];
    UnbiasedRNG[354] = LFSRcolor2[151];
    UnbiasedRNG[355] = LFSRcolor2[556];
    UnbiasedRNG[356] = LFSRcolor2[160];
    UnbiasedRNG[357] = LFSRcolor2[216];
    UnbiasedRNG[358] = LFSRcolor2[245];
    UnbiasedRNG[359] = LFSRcolor2[314];
    UnbiasedRNG[360] = LFSRcolor2[252];
    UnbiasedRNG[361] = LFSRcolor2[544];
    UnbiasedRNG[362] = LFSRcolor2[588];
    UnbiasedRNG[363] = LFSRcolor2[460];
    UnbiasedRNG[364] = LFSRcolor2[159];
    UnbiasedRNG[365] = LFSRcolor2[238];
    UnbiasedRNG[366] = LFSRcolor2[414];
    UnbiasedRNG[367] = LFSRcolor2[581];
    UnbiasedRNG[368] = LFSRcolor2[286];
    UnbiasedRNG[369] = LFSRcolor2[455];
    UnbiasedRNG[370] = LFSRcolor2[39];
    UnbiasedRNG[371] = LFSRcolor2[329];
    UnbiasedRNG[372] = LFSRcolor2[451];
    UnbiasedRNG[373] = LFSRcolor2[442];
    UnbiasedRNG[374] = LFSRcolor2[321];
    UnbiasedRNG[375] = LFSRcolor2[482];
    UnbiasedRNG[376] = LFSRcolor2[313];
    UnbiasedRNG[377] = LFSRcolor2[235];
    UnbiasedRNG[378] = LFSRcolor2[124];
    UnbiasedRNG[379] = LFSRcolor2[61];
    UnbiasedRNG[380] = LFSRcolor2[504];
    UnbiasedRNG[381] = LFSRcolor2[486];
    UnbiasedRNG[382] = LFSRcolor2[184];
    UnbiasedRNG[383] = LFSRcolor2[436];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[384] = LFSRcolor3[47];
    UnbiasedRNG[385] = LFSRcolor3[19];
    UnbiasedRNG[386] = LFSRcolor3[64];
    UnbiasedRNG[387] = LFSRcolor3[21];
    UnbiasedRNG[388] = LFSRcolor3[62];
    UnbiasedRNG[389] = LFSRcolor3[27];
    UnbiasedRNG[390] = LFSRcolor3[94];
    UnbiasedRNG[391] = LFSRcolor3[131];
    UnbiasedRNG[392] = LFSRcolor3[50];
    UnbiasedRNG[393] = LFSRcolor3[53];
    UnbiasedRNG[394] = LFSRcolor3[128];
    UnbiasedRNG[395] = LFSRcolor3[130];
    UnbiasedRNG[396] = LFSRcolor3[18];
    UnbiasedRNG[397] = LFSRcolor3[98];
    UnbiasedRNG[398] = LFSRcolor3[104];
    UnbiasedRNG[399] = LFSRcolor3[81];
    UnbiasedRNG[400] = LFSRcolor3[120];
    UnbiasedRNG[401] = LFSRcolor3[113];
    UnbiasedRNG[402] = LFSRcolor3[66];
    UnbiasedRNG[403] = LFSRcolor3[110];
    UnbiasedRNG[404] = LFSRcolor3[79];
    UnbiasedRNG[405] = LFSRcolor3[2];
    UnbiasedRNG[406] = LFSRcolor3[75];
    UnbiasedRNG[407] = LFSRcolor3[89];
    UnbiasedRNG[408] = LFSRcolor3[26];
    UnbiasedRNG[409] = LFSRcolor3[91];
    UnbiasedRNG[410] = LFSRcolor3[126];
    UnbiasedRNG[411] = LFSRcolor3[67];
    UnbiasedRNG[412] = LFSRcolor3[83];
    UnbiasedRNG[413] = LFSRcolor3[86];
    UnbiasedRNG[414] = LFSRcolor3[60];
    UnbiasedRNG[415] = LFSRcolor3[84];
    UnbiasedRNG[416] = LFSRcolor3[107];
    UnbiasedRNG[417] = LFSRcolor3[16];
    UnbiasedRNG[418] = LFSRcolor3[121];
    UnbiasedRNG[419] = LFSRcolor3[108];
    UnbiasedRNG[420] = LFSRcolor3[43];
    UnbiasedRNG[421] = LFSRcolor3[6];
    UnbiasedRNG[422] = LFSRcolor3[102];
    UnbiasedRNG[423] = LFSRcolor3[97];
    UnbiasedRNG[424] = LFSRcolor3[36];
    UnbiasedRNG[425] = LFSRcolor3[88];
    UnbiasedRNG[426] = LFSRcolor3[134];
    UnbiasedRNG[427] = LFSRcolor3[127];
    UnbiasedRNG[428] = LFSRcolor3[17];
    UnbiasedRNG[429] = LFSRcolor3[8];
    UnbiasedRNG[430] = LFSRcolor3[3];
    UnbiasedRNG[431] = LFSRcolor3[45];
    UnbiasedRNG[432] = LFSRcolor3[115];
    UnbiasedRNG[433] = LFSRcolor3[137];
    UnbiasedRNG[434] = LFSRcolor3[38];
    UnbiasedRNG[435] = LFSRcolor3[70];
    UnbiasedRNG[436] = LFSRcolor3[20];
    UnbiasedRNG[437] = LFSRcolor3[12];
    UnbiasedRNG[438] = LFSRcolor3[135];
    UnbiasedRNG[439] = LFSRcolor3[122];
    UnbiasedRNG[440] = LFSRcolor3[39];
    UnbiasedRNG[441] = LFSRcolor3[28];
    UnbiasedRNG[442] = LFSRcolor3[24];
    UnbiasedRNG[443] = LFSRcolor3[74];
    UnbiasedRNG[444] = LFSRcolor3[9];
    UnbiasedRNG[445] = LFSRcolor3[54];
    UnbiasedRNG[446] = LFSRcolor3[34];
    UnbiasedRNG[447] = LFSRcolor3[32];
    UnbiasedRNG[448] = LFSRcolor3[95];
    UnbiasedRNG[449] = LFSRcolor3[40];
    UnbiasedRNG[450] = LFSRcolor3[124];
    UnbiasedRNG[451] = LFSRcolor3[10];
    UnbiasedRNG[452] = LFSRcolor3[41];
    UnbiasedRNG[453] = LFSRcolor3[116];
    UnbiasedRNG[454] = LFSRcolor3[56];
    UnbiasedRNG[455] = LFSRcolor3[80];
    UnbiasedRNG[456] = LFSRcolor3[42];
    UnbiasedRNG[457] = LFSRcolor3[109];
    UnbiasedRNG[458] = LFSRcolor3[15];
    UnbiasedRNG[459] = LFSRcolor3[117];
    UnbiasedRNG[460] = LFSRcolor3[100];
    UnbiasedRNG[461] = LFSRcolor3[92];
    UnbiasedRNG[462] = LFSRcolor3[99];
    UnbiasedRNG[463] = LFSRcolor3[125];
    UnbiasedRNG[464] = LFSRcolor3[5];
    UnbiasedRNG[465] = LFSRcolor3[63];
    UnbiasedRNG[466] = LFSRcolor3[31];
    UnbiasedRNG[467] = LFSRcolor3[133];
    UnbiasedRNG[468] = LFSRcolor3[78];
    UnbiasedRNG[469] = LFSRcolor3[96];
    UnbiasedRNG[470] = LFSRcolor3[68];
    UnbiasedRNG[471] = LFSRcolor3[132];
    UnbiasedRNG[472] = LFSRcolor3[51];
    UnbiasedRNG[473] = LFSRcolor3[114];
    UnbiasedRNG[474] = LFSRcolor3[46];
    UnbiasedRNG[475] = LFSRcolor3[76];
    UnbiasedRNG[476] = LFSRcolor3[59];
    UnbiasedRNG[477] = LFSRcolor3[48];
    UnbiasedRNG[478] = LFSRcolor3[119];
    UnbiasedRNG[479] = LFSRcolor3[22];
    UnbiasedRNG[480] = LFSRcolor3[103];
    UnbiasedRNG[481] = LFSRcolor3[1];
    UnbiasedRNG[482] = LFSRcolor3[101];
    UnbiasedRNG[483] = LFSRcolor3[69];
    UnbiasedRNG[484] = LFSRcolor3[123];
    UnbiasedRNG[485] = LFSRcolor3[52];
    UnbiasedRNG[486] = LFSRcolor3[65];
    UnbiasedRNG[487] = LFSRcolor3[57];
    UnbiasedRNG[488] = LFSRcolor3[33];
    UnbiasedRNG[489] = LFSRcolor3[71];
    UnbiasedRNG[490] = LFSRcolor3[7];
    UnbiasedRNG[491] = LFSRcolor3[58];
    UnbiasedRNG[492] = LFSRcolor3[106];
    UnbiasedRNG[493] = LFSRcolor3[37];
end

always @(posedge color3_clk) begin
    BiasedRNG[527] = (LFSRcolor4[386]&LFSRcolor4[261]&LFSRcolor4[45]);
    BiasedRNG[528] = (LFSRcolor4[400]&LFSRcolor4[384]&LFSRcolor4[327]);
    BiasedRNG[529] = (LFSRcolor4[217]&LFSRcolor4[186]&LFSRcolor4[15]);
    BiasedRNG[530] = (LFSRcolor4[212]&LFSRcolor4[226]&LFSRcolor4[388]);
    BiasedRNG[531] = (LFSRcolor4[32]&LFSRcolor4[239]&LFSRcolor4[246]);
    BiasedRNG[532] = (LFSRcolor4[373]&LFSRcolor4[266]&LFSRcolor4[284]);
    BiasedRNG[533] = (LFSRcolor4[248]&LFSRcolor4[335]&LFSRcolor4[289]);
    BiasedRNG[534] = (LFSRcolor4[259]&LFSRcolor4[91]&LFSRcolor4[110]);
    BiasedRNG[535] = (LFSRcolor4[68]&LFSRcolor4[75]&LFSRcolor4[378]);
    BiasedRNG[536] = (LFSRcolor4[182]&LFSRcolor4[256]&LFSRcolor4[340]);
    BiasedRNG[537] = (LFSRcolor4[1]&LFSRcolor4[58]&LFSRcolor4[407]);
    BiasedRNG[538] = (LFSRcolor4[316]&LFSRcolor4[9]&LFSRcolor4[319]);
    BiasedRNG[539] = (LFSRcolor4[69]&LFSRcolor4[62]&LFSRcolor4[325]);
    BiasedRNG[540] = (LFSRcolor4[338]&LFSRcolor4[118]&LFSRcolor4[161]);
    BiasedRNG[541] = (LFSRcolor4[123]&LFSRcolor4[374]&LFSRcolor4[257]);
    BiasedRNG[542] = (LFSRcolor4[241]&LFSRcolor4[0]&LFSRcolor4[55]);
    BiasedRNG[543] = (LFSRcolor4[23]&LFSRcolor4[119]&LFSRcolor4[385]);
    BiasedRNG[544] = (LFSRcolor4[64]&LFSRcolor4[357]&LFSRcolor4[323]);
    BiasedRNG[545] = (LFSRcolor4[121]&LFSRcolor4[376]&LFSRcolor4[331]);
    BiasedRNG[546] = (LFSRcolor4[162]&LFSRcolor4[200]&LFSRcolor4[41]);
    BiasedRNG[547] = (LFSRcolor4[28]&LFSRcolor4[107]&LFSRcolor4[356]);
    BiasedRNG[548] = (LFSRcolor4[272]&LFSRcolor4[330]&LFSRcolor4[105]);
    BiasedRNG[549] = (LFSRcolor4[132]&LFSRcolor4[146]&LFSRcolor4[5]);
    BiasedRNG[550] = (LFSRcolor4[125]&LFSRcolor4[19]&LFSRcolor4[133]);
    BiasedRNG[551] = (LFSRcolor4[329]&LFSRcolor4[22]&LFSRcolor4[265]);
    BiasedRNG[552] = (LFSRcolor4[2]&LFSRcolor4[315]&LFSRcolor4[179]);
    BiasedRNG[553] = (LFSRcolor4[215]&LFSRcolor4[298]&LFSRcolor4[366]);
    BiasedRNG[554] = (LFSRcolor4[78]&LFSRcolor4[303]&LFSRcolor4[109]);
    BiasedRNG[555] = (LFSRcolor4[170]&LFSRcolor4[258]&LFSRcolor4[282]);
    BiasedRNG[556] = (LFSRcolor4[43]&LFSRcolor4[11]&LFSRcolor4[52]);
    BiasedRNG[557] = (LFSRcolor4[67]&LFSRcolor4[326]&LFSRcolor4[302]);
    BiasedRNG[558] = (LFSRcolor4[364]&LFSRcolor4[42]&LFSRcolor4[101]);
    BiasedRNG[559] = (LFSRcolor4[347]&LFSRcolor4[237]&LFSRcolor4[233]);
    BiasedRNG[560] = (LFSRcolor4[250]&LFSRcolor4[145]&LFSRcolor4[273]);
    BiasedRNG[561] = (LFSRcolor4[232]&LFSRcolor4[409]&LFSRcolor4[71]);
    BiasedRNG[562] = (LFSRcolor4[194]&LFSRcolor4[20]&LFSRcolor4[6]);
    BiasedRNG[563] = (LFSRcolor4[252]&LFSRcolor4[404]&LFSRcolor4[314]);
    BiasedRNG[564] = (LFSRcolor4[142]&LFSRcolor4[86]&LFSRcolor4[143]);
    BiasedRNG[565] = (LFSRcolor4[39]&LFSRcolor4[251]&LFSRcolor4[137]);
    BiasedRNG[566] = (LFSRcolor4[150]&LFSRcolor4[304]&LFSRcolor4[283]);
    BiasedRNG[567] = (LFSRcolor4[108]&LFSRcolor4[130]&LFSRcolor4[216]);
    BiasedRNG[568] = (LFSRcolor4[346]&LFSRcolor4[93]&LFSRcolor4[46]);
    BiasedRNG[569] = (LFSRcolor4[344]&LFSRcolor4[117]&LFSRcolor4[353]);
    BiasedRNG[570] = (LFSRcolor4[249]&LFSRcolor4[180]&LFSRcolor4[106]);
    BiasedRNG[571] = (LFSRcolor4[191]&LFSRcolor4[222]&LFSRcolor4[379]);
    BiasedRNG[572] = (LFSRcolor4[207]&LFSRcolor4[70]&LFSRcolor4[134]);
    BiasedRNG[573] = (LFSRcolor4[230]&LFSRcolor4[192]&LFSRcolor4[141]);
    BiasedRNG[574] = (LFSRcolor4[63]&LFSRcolor4[190]&LFSRcolor4[131]);
    BiasedRNG[575] = (LFSRcolor4[354]&LFSRcolor4[213]&LFSRcolor4[4]);
    BiasedRNG[576] = (LFSRcolor4[29]&LFSRcolor4[263]&LFSRcolor4[157]);
    BiasedRNG[577] = (LFSRcolor4[13]&LFSRcolor4[18]&LFSRcolor4[56]);
    BiasedRNG[578] = (LFSRcolor4[99]&LFSRcolor4[290]&LFSRcolor4[287]);
    BiasedRNG[579] = (LFSRcolor4[260]&LFSRcolor4[318]&LFSRcolor4[111]);
    BiasedRNG[580] = (LFSRcolor4[115]&LFSRcolor4[411]&LFSRcolor4[299]);
    BiasedRNG[581] = (LFSRcolor4[274]&LFSRcolor4[95]&LFSRcolor4[380]);
    BiasedRNG[582] = (LFSRcolor4[209]&LFSRcolor4[163]&LFSRcolor4[59]);
    BiasedRNG[583] = (LFSRcolor4[148]&LFSRcolor4[34]&LFSRcolor4[204]);
    BiasedRNG[584] = (LFSRcolor4[113]&LFSRcolor4[8]&LFSRcolor4[269]);
    BiasedRNG[585] = (LFSRcolor4[35]&LFSRcolor4[372]&LFSRcolor4[268]);
    BiasedRNG[586] = (LFSRcolor4[66]&LFSRcolor4[51]&LFSRcolor4[206]);
    BiasedRNG[587] = (LFSRcolor4[149]&LFSRcolor4[324]&LFSRcolor4[309]);
    BiasedRNG[588] = (LFSRcolor4[81]&LFSRcolor4[202]&LFSRcolor4[223]);
    BiasedRNG[589] = (LFSRcolor4[305]&LFSRcolor4[221]&LFSRcolor4[124]);
    BiasedRNG[590] = (LFSRcolor4[363]&LFSRcolor4[310]&LFSRcolor4[16]);
    BiasedRNG[591] = (LFSRcolor4[355]&LFSRcolor4[79]&LFSRcolor4[360]);
    BiasedRNG[592] = (LFSRcolor4[122]&LFSRcolor4[311]&LFSRcolor4[185]);
    BiasedRNG[593] = (LFSRcolor4[61]&LFSRcolor4[74]&LFSRcolor4[96]);
    BiasedRNG[594] = (LFSRcolor4[285]&LFSRcolor4[349]&LFSRcolor4[49]);
    BiasedRNG[595] = (LFSRcolor4[235]&LFSRcolor4[189]&LFSRcolor4[33]);
    BiasedRNG[596] = (LFSRcolor4[40]&LFSRcolor4[164]&LFSRcolor4[177]);
    BiasedRNG[597] = (LFSRcolor4[328]&LFSRcolor4[155]&LFSRcolor4[389]);
    BiasedRNG[598] = (LFSRcolor4[135]&LFSRcolor4[405]&LFSRcolor4[301]);
    BiasedRNG[599] = (LFSRcolor4[367]&LFSRcolor4[225]&LFSRcolor4[97]);
    BiasedRNG[600] = (LFSRcolor4[308]&LFSRcolor4[178]&LFSRcolor4[156]);
    BiasedRNG[601] = (LFSRcolor4[187]&LFSRcolor4[271]&LFSRcolor4[129]);
    BiasedRNG[602] = (LFSRcolor4[85]&LFSRcolor4[210]&LFSRcolor4[396]);
    BiasedRNG[603] = (LFSRcolor4[402]&LFSRcolor4[50]&LFSRcolor4[390]);
    BiasedRNG[604] = (LFSRcolor4[10]&LFSRcolor4[82]&LFSRcolor4[398]);
    BiasedRNG[605] = (LFSRcolor4[114]&LFSRcolor4[220]&LFSRcolor4[102]);
    BiasedRNG[606] = (LFSRcolor4[88]&LFSRcolor4[76]&LFSRcolor4[26]);
    BiasedRNG[607] = (LFSRcolor4[351]&LFSRcolor4[174]&LFSRcolor4[294]);
    BiasedRNG[608] = (LFSRcolor4[195]&LFSRcolor4[393]&LFSRcolor4[214]);
    BiasedRNG[609] = (LFSRcolor4[57]&LFSRcolor4[291]&LFSRcolor4[307]);
    BiasedRNG[610] = (LFSRcolor4[151]&LFSRcolor4[262]&LFSRcolor4[196]);
    BiasedRNG[611] = (LFSRcolor4[65]&LFSRcolor4[100]&LFSRcolor4[138]);
    BiasedRNG[612] = (LFSRcolor4[236]&LFSRcolor4[30]&LFSRcolor4[47]);
    BiasedRNG[613] = (LFSRcolor4[188]&LFSRcolor4[54]&LFSRcolor4[73]);
    BiasedRNG[614] = (LFSRcolor4[339]&LFSRcolor4[77]&LFSRcolor4[397]);
    BiasedRNG[615] = (LFSRcolor4[345]&LFSRcolor4[403]&LFSRcolor4[406]);
    BiasedRNG[616] = (LFSRcolor4[152]&LFSRcolor4[254]&LFSRcolor4[264]);
    BiasedRNG[617] = (LFSRcolor4[306]&LFSRcolor4[392]&LFSRcolor4[288]);
    BiasedRNG[618] = (LFSRcolor4[343]&LFSRcolor4[38]&LFSRcolor4[321]);
    BiasedRNG[619] = (LFSRcolor4[169]&LFSRcolor4[48]&LFSRcolor4[391]);
    BiasedRNG[620] = (LFSRcolor4[37]&LFSRcolor4[322]&LFSRcolor4[375]);
    BiasedRNG[621] = (LFSRcolor4[172]&LFSRcolor4[90]&LFSRcolor4[348]);
    BiasedRNG[622] = (LFSRcolor4[242]&LFSRcolor4[153]&LFSRcolor4[165]);
    BiasedRNG[623] = (LFSRcolor4[173]&LFSRcolor4[89]&LFSRcolor4[3]);
    BiasedRNG[624] = (LFSRcolor4[381]&LFSRcolor4[92]&LFSRcolor4[317]);
    BiasedRNG[625] = (LFSRcolor4[255]&LFSRcolor4[413]&LFSRcolor4[276]);
    BiasedRNG[626] = (LFSRcolor4[371]&LFSRcolor4[140]&LFSRcolor4[293]);
    BiasedRNG[627] = (LFSRcolor4[154]&LFSRcolor4[126]&LFSRcolor4[229]);
    BiasedRNG[628] = (LFSRcolor4[292]&LFSRcolor4[300]&LFSRcolor4[224]);
    BiasedRNG[629] = (LFSRcolor4[112]&LFSRcolor4[296]&LFSRcolor4[139]);
    BiasedRNG[630] = (LFSRcolor4[84]&LFSRcolor4[231]&LFSRcolor4[228]);
    BiasedRNG[631] = (LFSRcolor4[80]&LFSRcolor4[240]&LFSRcolor4[234]);
    BiasedRNG[632] = (LFSRcolor4[183]&LFSRcolor4[104]&LFSRcolor4[368]);
    BiasedRNG[633] = (LFSRcolor4[144]&LFSRcolor4[401]&LFSRcolor4[275]);
    BiasedRNG[634] = (LFSRcolor4[53]&LFSRcolor4[175]&LFSRcolor4[399]);
    BiasedRNG[635] = (LFSRcolor4[358]&LFSRcolor4[116]&LFSRcolor4[408]);
    BiasedRNG[636] = (LFSRcolor4[218]&LFSRcolor4[267]&LFSRcolor4[336]);
    BiasedRNG[637] = (LFSRcolor4[203]&LFSRcolor4[147]&LFSRcolor4[297]);
    BiasedRNG[638] = (LFSRcolor4[184]&LFSRcolor4[332]&LFSRcolor4[94]);
    BiasedRNG[639] = (LFSRcolor4[36]&LFSRcolor4[160]&LFSRcolor4[387]);
    BiasedRNG[640] = (LFSRcolor4[369]&LFSRcolor4[136]&LFSRcolor4[60]);
    BiasedRNG[641] = (LFSRcolor4[219]&LFSRcolor4[412]&LFSRcolor4[370]);
    BiasedRNG[642] = (LFSRcolor4[127]&LFSRcolor4[365]&LFSRcolor4[197]);
    BiasedRNG[643] = (LFSRcolor4[243]&LFSRcolor4[158]&LFSRcolor4[312]);
    BiasedRNG[644] = (LFSRcolor4[17]&LFSRcolor4[21]&LFSRcolor4[342]);
    BiasedRNG[645] = (LFSRcolor4[334]&LFSRcolor4[253]&LFSRcolor4[278]);
    BiasedRNG[646] = (LFSRcolor4[383]&LFSRcolor4[128]&LFSRcolor4[199]);
    BiasedRNG[647] = (LFSRcolor4[211]&LFSRcolor4[333]&LFSRcolor4[359]);
    BiasedRNG[648] = (LFSRcolor4[281]&LFSRcolor4[24]&LFSRcolor4[352]);
    BiasedRNG[649] = (LFSRcolor4[313]&LFSRcolor4[244]&LFSRcolor4[198]);
    BiasedRNG[650] = (LFSRcolor4[166]&LFSRcolor4[171]&LFSRcolor4[201]);
    BiasedRNG[651] = (LFSRcolor4[27]&LFSRcolor4[247]&LFSRcolor4[394]);
    BiasedRNG[652] = (LFSRcolor4[7]&LFSRcolor4[31]&LFSRcolor4[25]);
    BiasedRNG[653] = (LFSRcolor4[410]&LFSRcolor4[167]&LFSRcolor4[286]);
    BiasedRNG[654] = (LFSRcolor4[362]&LFSRcolor4[337]&LFSRcolor4[377]);
    BiasedRNG[655] = (LFSRcolor4[395]&LFSRcolor4[87]&LFSRcolor4[238]);
    BiasedRNG[656] = (LFSRcolor4[83]&LFSRcolor4[361]&LFSRcolor4[168]);
    BiasedRNG[657] = (LFSRcolor4[280]&LFSRcolor4[205]&LFSRcolor4[12]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

//Generate the ILA for data collection:
ila_0 ILAinst(.clk(sample_clk),.probe0(run),.probe1(solution_flag),.probe2(failure),.probe3(counter[37:0]));

//Instantiate VIO:
vio_0 VIOinst (.clk(sample_clk),.probe_out0(reset),.probe_out1(solution_set[23:0]));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule