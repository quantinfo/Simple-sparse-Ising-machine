//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [37:0] counter;
initial counter = 38'b0;
reg [27:0] solution;
reg [27:0] solution_check;
wire [27:0] solution_set;
initial solution_check = 28'b1111110011100010001001000111;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
reg [0:1595] InitCond;
reg run;
wire [965:0] LFSRcolor0;
wire [965:0] LFSRcolor1;
wire [781:0] LFSRcolor2;
wire [183:0] LFSRcolor3;
wire [551:0] LFSRcolor4;
reg [879:0] BiasedRNG;       //For I=+/-1 cases
reg [715:0] UnbiasedRNG;   //For I=0 cases
reg [0:1637] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[532] = 1'b1;
initial m[731] = 1'b1;
initial m[741] = 1'b1;
initial m[756] = 1'b0;
initial m[776] = 1'b0;
initial m[801] = 1'b0;
initial m[831] = 1'b1;
initial m[866] = 1'b0;
initial m[906] = 1'b0;
initial m[951] = 1'b1;
initial m[1001] = 1'b0;
initial m[1056] = 1'b0;
initial m[1116] = 1'b0;
initial m[1181] = 1'b1;
initial m[1246] = 1'b0;
initial m[1306] = 1'b0;
initial m[1361] = 1'b0;
initial m[1411] = 1'b1;
initial m[1456] = 1'b1;
initial m[1496] = 1'b1;
initial m[1531] = 1'b0;
initial m[1561] = 1'b0;
initial m[1586] = 1'b1;
initial m[1606] = 1'b1;
initial m[1621] = 1'b1;
initial m[1631] = 1'b1;
initial m[1636] = 1'b1;
initial m[1637] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[730] = 1'b0;
initial m[740] = 1'b0;
initial m[755] = 1'b0;
initial m[775] = 1'b0;
initial m[800] = 1'b0;
initial m[830] = 1'b0;
initial m[865] = 1'b0;
initial m[905] = 1'b0;
initial m[950] = 1'b0;
initial m[1000] = 1'b0;
initial m[1055] = 1'b0;
initial m[1115] = 1'b0;
initial m[1180] = 1'b0;
initial m[1183] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR0_11(.LFSRregister(LFSRcolor0[551:506]),.clk(sample_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR0_12(.LFSRregister(LFSRcolor0[597:552]),.clk(sample_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR0_13(.LFSRregister(LFSRcolor0[643:598]),.clk(sample_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR0_14(.LFSRregister(LFSRcolor0[689:644]),.clk(sample_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR0_15(.LFSRregister(LFSRcolor0[735:690]),.clk(sample_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR0_16(.LFSRregister(LFSRcolor0[781:736]),.clk(sample_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR0_17(.LFSRregister(LFSRcolor0[827:782]),.clk(sample_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR0_18(.LFSRregister(LFSRcolor0[873:828]),.clk(sample_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR0_19(.LFSRregister(LFSRcolor0[919:874]),.clk(sample_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR0_20(.LFSRregister(LFSRcolor0[965:920]),.clk(sample_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR1_15(.LFSRregister(LFSRcolor1[735:690]),.clk(color0_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR1_16(.LFSRregister(LFSRcolor1[781:736]),.clk(color0_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR1_17(.LFSRregister(LFSRcolor1[827:782]),.clk(color0_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR1_18(.LFSRregister(LFSRcolor1[873:828]),.clk(color0_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR1_19(.LFSRregister(LFSRcolor1[919:874]),.clk(color0_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR1_20(.LFSRregister(LFSRcolor1[965:920]),.clk(color0_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0011001000010001001111001110101111011111000110)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b0101000110100000010101001000010000101101100110)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b1110011010010011001010111010100101111111100000)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b1001111000010100100001100010110000001111101011)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b0011101001111100110111000000010000101100111110)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b1010111010001100001100010110010011100100101100)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b1101010000110001000001011010110100010000110101)) LFSR2_11(.LFSRregister(LFSRcolor2[551:506]),.clk(color1_clk));
lfsr #(.seed(46'b0111111000001001010001100011001110110101101001)) LFSR2_12(.LFSRregister(LFSRcolor2[597:552]),.clk(color1_clk));
lfsr #(.seed(46'b0111011110101100100001111000001001111001010010)) LFSR2_13(.LFSRregister(LFSRcolor2[643:598]),.clk(color1_clk));
lfsr #(.seed(46'b0110010001011011111100000000110011011110000100)) LFSR2_14(.LFSRregister(LFSRcolor2[689:644]),.clk(color1_clk));
lfsr #(.seed(46'b1100101101001001110010011101110000001110111111)) LFSR2_15(.LFSRregister(LFSRcolor2[735:690]),.clk(color1_clk));
lfsr #(.seed(46'b1110010100000011100111110011000001001000000101)) LFSR2_16(.LFSRregister(LFSRcolor2[781:736]),.clk(color1_clk));
lfsr #(.seed(46'b1100111110111110000101110101010111111010101000)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1101101000110111001110111111011011100011111101)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b1011100111101011110000001101111100001111100011)) LFSR3_2(.LFSRregister(LFSRcolor3[137:92]),.clk(color2_clk));
lfsr #(.seed(46'b1000011101010100110111010000000111000111010111)) LFSR3_3(.LFSRregister(LFSRcolor3[183:138]),.clk(color2_clk));
lfsr #(.seed(46'b0011001001101100101110110001011100100100110000)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b0011110010011101000111111110100110110100101000)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1100000100011100010111001011000000101100110100)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b1001101001101101001001111001110100110001100010)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b1000000000001101011011010100000001101001001111)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b1000011000100000010011100100110100001010000001)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b0101000011110010010110011011111101010101011010)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b0011111001110010110000110100101000000000100010)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));
lfsr #(.seed(46'b0011101001110100101101111100101010101100110000)) LFSR4_8(.LFSRregister(LFSRcolor4[413:368]),.clk(color3_clk));
lfsr #(.seed(46'b1100111100001111010111011100011110001010110011)) LFSR4_9(.LFSRregister(LFSRcolor4[459:414]),.clk(color3_clk));
lfsr #(.seed(46'b0101101111111000101111101010111101100011110011)) LFSR4_10(.LFSRregister(LFSRcolor4[505:460]),.clk(color3_clk));
lfsr #(.seed(46'b1100101101101111100100111011110111010010100100)) LFSR4_11(.LFSRregister(LFSRcolor4[551:506]),.clk(color3_clk));
//To control whether the system runs or resets using VIO and counter:
always @(posedge sample_clk) begin
    if (reset) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 28'b0;
        failure = 1'b0;
        solution_check = solution_set;
        m[532] = solution_set[0];
        m[731] = solution_set[1];
        m[741] = solution_set[2];
        m[756] = solution_set[3];
        m[776] = solution_set[4];
        m[801] = solution_set[5];
        m[831] = solution_set[6];
        m[866] = solution_set[7];
        m[906] = solution_set[8];
        m[951] = solution_set[9];
        m[1001] = solution_set[10];
        m[1056] = solution_set[11];
        m[1116] = solution_set[12];
        m[1181] = solution_set[13];
        m[1246] = solution_set[14];
        m[1306] = solution_set[15];
        m[1361] = solution_set[16];
        m[1411] = solution_set[17];
        m[1456] = solution_set[18];
        m[1496] = solution_set[19];
        m[1531] = solution_set[20];
        m[1561] = solution_set[21];
        m[1586] = solution_set[22];
        m[1606] = solution_set[23];
        m[1621] = solution_set[24];
        m[1631] = solution_set[25];
        m[1636] = solution_set[26];
        m[1637] = solution_set[27];
    end else if (solution_flag) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 28'b0;
        failure = 1'b0;
    end else if (counter < 38'b11111111111111111111111111111111111111) begin
        if (counter == 1) begin
            InitCond[0] = UnbiasedRNG[0];
            InitCond[1] = UnbiasedRNG[1];
            InitCond[2] = UnbiasedRNG[2];
            InitCond[3] = UnbiasedRNG[3];
            InitCond[4] = UnbiasedRNG[4];
            InitCond[5] = UnbiasedRNG[5];
            InitCond[6] = UnbiasedRNG[6];
            InitCond[7] = UnbiasedRNG[7];
            InitCond[8] = UnbiasedRNG[8];
            InitCond[9] = UnbiasedRNG[9];
            InitCond[10] = UnbiasedRNG[10];
            InitCond[11] = UnbiasedRNG[11];
            InitCond[12] = UnbiasedRNG[12];
            InitCond[13] = UnbiasedRNG[13];
            InitCond[14] = UnbiasedRNG[14];
            InitCond[15] = UnbiasedRNG[15];
            InitCond[16] = UnbiasedRNG[16];
            InitCond[17] = UnbiasedRNG[17];
            InitCond[18] = UnbiasedRNG[18];
            InitCond[19] = UnbiasedRNG[19];
            InitCond[20] = UnbiasedRNG[20];
            InitCond[21] = UnbiasedRNG[21];
            InitCond[22] = UnbiasedRNG[22];
            InitCond[23] = UnbiasedRNG[23];
            InitCond[24] = UnbiasedRNG[24];
            InitCond[25] = UnbiasedRNG[25];
            InitCond[26] = UnbiasedRNG[26];
            InitCond[27] = UnbiasedRNG[27];
            InitCond[28] = UnbiasedRNG[28];
            InitCond[29] = UnbiasedRNG[29];
            InitCond[30] = UnbiasedRNG[30];
            InitCond[31] = UnbiasedRNG[31];
            InitCond[32] = UnbiasedRNG[32];
            InitCond[33] = UnbiasedRNG[33];
            InitCond[34] = UnbiasedRNG[34];
            InitCond[35] = UnbiasedRNG[35];
            InitCond[36] = UnbiasedRNG[36];
            InitCond[37] = UnbiasedRNG[37];
            InitCond[38] = UnbiasedRNG[38];
            InitCond[39] = UnbiasedRNG[39];
            InitCond[40] = UnbiasedRNG[40];
            InitCond[41] = UnbiasedRNG[41];
            InitCond[42] = UnbiasedRNG[42];
            InitCond[43] = UnbiasedRNG[43];
            InitCond[44] = UnbiasedRNG[44];
            InitCond[45] = UnbiasedRNG[45];
            InitCond[46] = UnbiasedRNG[46];
            InitCond[47] = UnbiasedRNG[47];
            InitCond[48] = UnbiasedRNG[48];
            InitCond[49] = UnbiasedRNG[49];
            InitCond[50] = UnbiasedRNG[50];
            InitCond[51] = UnbiasedRNG[51];
            InitCond[52] = UnbiasedRNG[52];
            InitCond[53] = UnbiasedRNG[53];
            InitCond[54] = UnbiasedRNG[54];
            InitCond[55] = UnbiasedRNG[55];
            InitCond[56] = UnbiasedRNG[56];
            InitCond[57] = UnbiasedRNG[57];
            InitCond[58] = UnbiasedRNG[58];
            InitCond[59] = UnbiasedRNG[59];
            InitCond[60] = UnbiasedRNG[60];
            InitCond[61] = UnbiasedRNG[61];
            InitCond[62] = UnbiasedRNG[62];
            InitCond[63] = UnbiasedRNG[63];
            InitCond[64] = UnbiasedRNG[64];
            InitCond[65] = UnbiasedRNG[65];
            InitCond[66] = UnbiasedRNG[66];
            InitCond[67] = UnbiasedRNG[67];
            InitCond[68] = UnbiasedRNG[68];
            InitCond[69] = UnbiasedRNG[69];
            InitCond[70] = UnbiasedRNG[70];
            InitCond[71] = UnbiasedRNG[71];
            InitCond[72] = UnbiasedRNG[72];
            InitCond[73] = UnbiasedRNG[73];
            InitCond[74] = UnbiasedRNG[74];
            InitCond[75] = UnbiasedRNG[75];
            InitCond[76] = UnbiasedRNG[76];
            InitCond[77] = UnbiasedRNG[77];
            InitCond[78] = UnbiasedRNG[78];
            InitCond[79] = UnbiasedRNG[79];
            InitCond[80] = UnbiasedRNG[80];
            InitCond[81] = UnbiasedRNG[81];
            InitCond[82] = UnbiasedRNG[82];
            InitCond[83] = UnbiasedRNG[83];
            InitCond[84] = UnbiasedRNG[84];
            InitCond[85] = UnbiasedRNG[85];
            InitCond[86] = UnbiasedRNG[86];
            InitCond[87] = UnbiasedRNG[87];
            InitCond[88] = UnbiasedRNG[88];
            InitCond[89] = UnbiasedRNG[89];
            InitCond[90] = UnbiasedRNG[90];
            InitCond[91] = UnbiasedRNG[91];
            InitCond[92] = UnbiasedRNG[92];
            InitCond[93] = UnbiasedRNG[93];
            InitCond[94] = UnbiasedRNG[94];
            InitCond[95] = UnbiasedRNG[95];
            InitCond[96] = UnbiasedRNG[96];
            InitCond[97] = UnbiasedRNG[97];
            InitCond[98] = UnbiasedRNG[98];
            InitCond[99] = UnbiasedRNG[99];
            InitCond[100] = UnbiasedRNG[100];
            InitCond[101] = UnbiasedRNG[101];
            InitCond[102] = UnbiasedRNG[102];
            InitCond[103] = UnbiasedRNG[103];
            InitCond[104] = UnbiasedRNG[104];
            InitCond[105] = UnbiasedRNG[105];
            InitCond[106] = UnbiasedRNG[106];
            InitCond[107] = UnbiasedRNG[107];
            InitCond[108] = UnbiasedRNG[108];
            InitCond[109] = UnbiasedRNG[109];
            InitCond[110] = UnbiasedRNG[110];
            InitCond[111] = UnbiasedRNG[111];
            InitCond[112] = UnbiasedRNG[112];
            InitCond[113] = UnbiasedRNG[113];
            InitCond[114] = UnbiasedRNG[114];
            InitCond[115] = UnbiasedRNG[115];
            InitCond[116] = UnbiasedRNG[116];
            InitCond[117] = UnbiasedRNG[117];
            InitCond[118] = UnbiasedRNG[118];
            InitCond[119] = UnbiasedRNG[119];
            InitCond[120] = UnbiasedRNG[120];
            InitCond[121] = UnbiasedRNG[121];
            InitCond[122] = UnbiasedRNG[122];
            InitCond[123] = UnbiasedRNG[123];
            InitCond[124] = UnbiasedRNG[124];
            InitCond[125] = UnbiasedRNG[125];
            InitCond[126] = UnbiasedRNG[126];
            InitCond[127] = UnbiasedRNG[127];
            InitCond[128] = UnbiasedRNG[128];
            InitCond[129] = UnbiasedRNG[129];
            InitCond[130] = UnbiasedRNG[130];
            InitCond[131] = UnbiasedRNG[131];
            InitCond[132] = UnbiasedRNG[132];
            InitCond[133] = UnbiasedRNG[133];
            InitCond[134] = UnbiasedRNG[134];
            InitCond[135] = UnbiasedRNG[135];
            InitCond[136] = UnbiasedRNG[136];
            InitCond[137] = UnbiasedRNG[137];
            InitCond[138] = UnbiasedRNG[138];
            InitCond[139] = UnbiasedRNG[139];
            InitCond[140] = UnbiasedRNG[140];
            InitCond[141] = UnbiasedRNG[141];
            InitCond[142] = UnbiasedRNG[142];
            InitCond[143] = UnbiasedRNG[143];
            InitCond[144] = UnbiasedRNG[144];
            InitCond[145] = UnbiasedRNG[145];
            InitCond[146] = UnbiasedRNG[146];
            InitCond[147] = UnbiasedRNG[147];
            InitCond[148] = UnbiasedRNG[148];
            InitCond[149] = UnbiasedRNG[149];
            InitCond[150] = UnbiasedRNG[150];
            InitCond[151] = UnbiasedRNG[151];
            InitCond[152] = UnbiasedRNG[152];
            InitCond[153] = UnbiasedRNG[153];
            InitCond[154] = UnbiasedRNG[154];
            InitCond[155] = UnbiasedRNG[155];
            InitCond[156] = UnbiasedRNG[156];
            InitCond[157] = UnbiasedRNG[157];
            InitCond[158] = UnbiasedRNG[158];
            InitCond[159] = UnbiasedRNG[159];
            InitCond[160] = UnbiasedRNG[160];
            InitCond[161] = UnbiasedRNG[161];
            InitCond[162] = UnbiasedRNG[162];
            InitCond[163] = UnbiasedRNG[163];
            InitCond[164] = UnbiasedRNG[164];
            InitCond[165] = UnbiasedRNG[165];
            InitCond[166] = UnbiasedRNG[166];
            InitCond[167] = UnbiasedRNG[167];
            InitCond[168] = UnbiasedRNG[168];
            InitCond[169] = UnbiasedRNG[169];
            InitCond[170] = UnbiasedRNG[170];
            InitCond[171] = UnbiasedRNG[171];
            InitCond[172] = UnbiasedRNG[172];
            InitCond[173] = UnbiasedRNG[173];
            InitCond[174] = UnbiasedRNG[174];
            InitCond[175] = UnbiasedRNG[175];
            InitCond[176] = UnbiasedRNG[176];
            InitCond[177] = UnbiasedRNG[177];
            InitCond[178] = UnbiasedRNG[178];
            InitCond[179] = UnbiasedRNG[179];
            InitCond[180] = UnbiasedRNG[180];
            InitCond[181] = UnbiasedRNG[181];
            InitCond[182] = UnbiasedRNG[182];
            InitCond[183] = UnbiasedRNG[183];
            InitCond[184] = UnbiasedRNG[184];
            InitCond[185] = UnbiasedRNG[185];
            InitCond[186] = UnbiasedRNG[186];
            InitCond[187] = UnbiasedRNG[187];
            InitCond[188] = UnbiasedRNG[188];
            InitCond[189] = UnbiasedRNG[189];
            InitCond[190] = UnbiasedRNG[190];
            InitCond[191] = UnbiasedRNG[191];
            InitCond[192] = UnbiasedRNG[192];
            InitCond[193] = UnbiasedRNG[193];
            InitCond[194] = UnbiasedRNG[194];
            InitCond[195] = UnbiasedRNG[195];
            InitCond[196] = UnbiasedRNG[196];
            InitCond[197] = UnbiasedRNG[197];
            InitCond[198] = UnbiasedRNG[198];
            InitCond[199] = UnbiasedRNG[199];
            InitCond[200] = UnbiasedRNG[200];
            InitCond[201] = UnbiasedRNG[201];
            InitCond[202] = UnbiasedRNG[202];
            InitCond[203] = UnbiasedRNG[203];
            InitCond[204] = UnbiasedRNG[204];
            InitCond[205] = UnbiasedRNG[205];
            InitCond[206] = UnbiasedRNG[206];
            InitCond[207] = UnbiasedRNG[207];
            InitCond[208] = UnbiasedRNG[208];
            InitCond[209] = UnbiasedRNG[209];
            InitCond[210] = UnbiasedRNG[210];
            InitCond[211] = UnbiasedRNG[211];
            InitCond[212] = UnbiasedRNG[212];
            InitCond[213] = UnbiasedRNG[213];
            InitCond[214] = UnbiasedRNG[214];
            InitCond[215] = UnbiasedRNG[215];
            InitCond[216] = UnbiasedRNG[216];
            InitCond[217] = UnbiasedRNG[217];
            InitCond[218] = UnbiasedRNG[218];
            InitCond[219] = UnbiasedRNG[219];
            InitCond[220] = UnbiasedRNG[220];
            InitCond[221] = UnbiasedRNG[221];
            InitCond[222] = UnbiasedRNG[222];
            InitCond[223] = UnbiasedRNG[223];
            InitCond[224] = UnbiasedRNG[224];
            InitCond[225] = UnbiasedRNG[225];
            InitCond[226] = UnbiasedRNG[226];
            InitCond[227] = UnbiasedRNG[227];
            InitCond[228] = UnbiasedRNG[228];
            InitCond[229] = UnbiasedRNG[229];
            InitCond[230] = UnbiasedRNG[230];
            InitCond[231] = UnbiasedRNG[231];
            InitCond[232] = UnbiasedRNG[232];
            InitCond[233] = UnbiasedRNG[233];
            InitCond[234] = UnbiasedRNG[234];
            InitCond[235] = UnbiasedRNG[235];
            InitCond[236] = UnbiasedRNG[236];
            InitCond[237] = UnbiasedRNG[237];
            InitCond[238] = UnbiasedRNG[238];
            InitCond[239] = UnbiasedRNG[239];
            InitCond[240] = UnbiasedRNG[240];
            InitCond[241] = UnbiasedRNG[241];
            InitCond[242] = UnbiasedRNG[242];
            InitCond[243] = UnbiasedRNG[243];
            InitCond[244] = UnbiasedRNG[244];
            InitCond[245] = UnbiasedRNG[245];
            InitCond[246] = UnbiasedRNG[246];
            InitCond[247] = UnbiasedRNG[247];
            InitCond[248] = UnbiasedRNG[248];
            InitCond[249] = UnbiasedRNG[249];
            InitCond[250] = UnbiasedRNG[250];
            InitCond[251] = UnbiasedRNG[251];
            InitCond[252] = UnbiasedRNG[252];
            InitCond[253] = UnbiasedRNG[253];
            InitCond[254] = UnbiasedRNG[254];
            InitCond[255] = UnbiasedRNG[255];
            InitCond[256] = UnbiasedRNG[256];
            InitCond[257] = UnbiasedRNG[257];
            InitCond[258] = UnbiasedRNG[258];
            InitCond[259] = UnbiasedRNG[259];
            InitCond[260] = UnbiasedRNG[260];
            InitCond[261] = UnbiasedRNG[261];
            InitCond[262] = UnbiasedRNG[262];
            InitCond[263] = UnbiasedRNG[263];
            InitCond[264] = UnbiasedRNG[264];
            InitCond[265] = UnbiasedRNG[265];
            InitCond[266] = UnbiasedRNG[266];
            InitCond[267] = UnbiasedRNG[267];
            InitCond[268] = UnbiasedRNG[268];
            InitCond[269] = UnbiasedRNG[269];
            InitCond[270] = UnbiasedRNG[270];
            InitCond[271] = UnbiasedRNG[271];
            InitCond[272] = UnbiasedRNG[272];
            InitCond[273] = UnbiasedRNG[273];
            InitCond[274] = UnbiasedRNG[274];
            InitCond[275] = UnbiasedRNG[275];
            InitCond[276] = UnbiasedRNG[276];
            InitCond[277] = UnbiasedRNG[277];
            InitCond[278] = UnbiasedRNG[278];
            InitCond[279] = UnbiasedRNG[279];
            InitCond[280] = UnbiasedRNG[280];
            InitCond[281] = UnbiasedRNG[281];
            InitCond[282] = UnbiasedRNG[282];
            InitCond[283] = UnbiasedRNG[283];
            InitCond[284] = UnbiasedRNG[284];
            InitCond[285] = UnbiasedRNG[285];
            InitCond[286] = UnbiasedRNG[286];
            InitCond[287] = UnbiasedRNG[287];
            InitCond[288] = UnbiasedRNG[288];
            InitCond[289] = UnbiasedRNG[289];
            InitCond[290] = UnbiasedRNG[290];
            InitCond[291] = UnbiasedRNG[291];
            InitCond[292] = UnbiasedRNG[292];
            InitCond[293] = UnbiasedRNG[293];
            InitCond[294] = UnbiasedRNG[294];
            InitCond[295] = UnbiasedRNG[295];
            InitCond[296] = UnbiasedRNG[296];
            InitCond[297] = UnbiasedRNG[297];
            InitCond[298] = UnbiasedRNG[298];
            InitCond[299] = UnbiasedRNG[299];
            InitCond[300] = UnbiasedRNG[300];
            InitCond[301] = UnbiasedRNG[301];
            InitCond[302] = UnbiasedRNG[302];
            InitCond[303] = UnbiasedRNG[303];
            InitCond[304] = UnbiasedRNG[304];
            InitCond[305] = UnbiasedRNG[305];
            InitCond[306] = UnbiasedRNG[306];
            InitCond[307] = UnbiasedRNG[307];
            InitCond[308] = UnbiasedRNG[308];
            InitCond[309] = UnbiasedRNG[309];
            InitCond[310] = UnbiasedRNG[310];
            InitCond[311] = UnbiasedRNG[311];
            InitCond[312] = UnbiasedRNG[312];
            InitCond[313] = UnbiasedRNG[313];
            InitCond[314] = UnbiasedRNG[314];
            InitCond[315] = UnbiasedRNG[315];
            InitCond[316] = UnbiasedRNG[316];
            InitCond[317] = UnbiasedRNG[317];
            InitCond[318] = UnbiasedRNG[318];
            InitCond[319] = UnbiasedRNG[319];
            InitCond[320] = UnbiasedRNG[320];
            InitCond[321] = UnbiasedRNG[321];
            InitCond[322] = UnbiasedRNG[322];
            InitCond[323] = UnbiasedRNG[323];
            InitCond[324] = UnbiasedRNG[324];
            InitCond[325] = UnbiasedRNG[325];
            InitCond[326] = UnbiasedRNG[326];
            InitCond[327] = UnbiasedRNG[327];
            InitCond[328] = UnbiasedRNG[328];
            InitCond[329] = UnbiasedRNG[329];
            InitCond[330] = UnbiasedRNG[330];
            InitCond[331] = UnbiasedRNG[331];
            InitCond[332] = UnbiasedRNG[332];
            InitCond[333] = UnbiasedRNG[333];
            InitCond[334] = UnbiasedRNG[334];
            InitCond[335] = UnbiasedRNG[335];
            InitCond[336] = UnbiasedRNG[336];
            InitCond[337] = UnbiasedRNG[337];
            InitCond[338] = UnbiasedRNG[338];
            InitCond[339] = UnbiasedRNG[339];
            InitCond[340] = UnbiasedRNG[340];
            InitCond[341] = UnbiasedRNG[341];
            InitCond[342] = UnbiasedRNG[342];
            InitCond[343] = UnbiasedRNG[343];
            InitCond[344] = UnbiasedRNG[344];
            InitCond[345] = UnbiasedRNG[345];
            InitCond[346] = UnbiasedRNG[346];
            InitCond[347] = UnbiasedRNG[347];
            InitCond[348] = UnbiasedRNG[348];
            InitCond[349] = UnbiasedRNG[349];
            InitCond[350] = UnbiasedRNG[350];
            InitCond[351] = UnbiasedRNG[351];
            InitCond[352] = UnbiasedRNG[352];
            InitCond[353] = UnbiasedRNG[353];
            InitCond[354] = UnbiasedRNG[354];
            InitCond[355] = UnbiasedRNG[355];
            InitCond[356] = UnbiasedRNG[356];
            InitCond[357] = UnbiasedRNG[357];
            InitCond[358] = UnbiasedRNG[358];
            InitCond[359] = UnbiasedRNG[359];
            InitCond[360] = UnbiasedRNG[360];
            InitCond[361] = UnbiasedRNG[361];
            InitCond[362] = UnbiasedRNG[362];
            InitCond[363] = UnbiasedRNG[363];
            InitCond[364] = UnbiasedRNG[364];
            InitCond[365] = UnbiasedRNG[365];
            InitCond[366] = UnbiasedRNG[366];
            InitCond[367] = UnbiasedRNG[367];
            InitCond[368] = UnbiasedRNG[368];
            InitCond[369] = UnbiasedRNG[369];
            InitCond[370] = UnbiasedRNG[370];
            InitCond[371] = UnbiasedRNG[371];
            InitCond[372] = UnbiasedRNG[372];
            InitCond[373] = UnbiasedRNG[373];
            InitCond[374] = UnbiasedRNG[374];
            InitCond[375] = UnbiasedRNG[375];
            InitCond[376] = UnbiasedRNG[376];
            InitCond[377] = UnbiasedRNG[377];
            InitCond[378] = UnbiasedRNG[378];
            InitCond[379] = UnbiasedRNG[379];
            InitCond[380] = UnbiasedRNG[380];
            InitCond[381] = UnbiasedRNG[381];
            InitCond[382] = UnbiasedRNG[382];
            InitCond[383] = UnbiasedRNG[383];
            InitCond[384] = UnbiasedRNG[384];
            InitCond[385] = UnbiasedRNG[385];
            InitCond[386] = UnbiasedRNG[386];
            InitCond[387] = UnbiasedRNG[387];
            InitCond[388] = UnbiasedRNG[388];
            InitCond[389] = UnbiasedRNG[389];
            InitCond[390] = UnbiasedRNG[390];
            InitCond[391] = UnbiasedRNG[391];
            InitCond[392] = UnbiasedRNG[392];
            InitCond[393] = UnbiasedRNG[393];
            InitCond[394] = UnbiasedRNG[394];
            InitCond[395] = UnbiasedRNG[395];
            InitCond[396] = UnbiasedRNG[396];
            InitCond[397] = UnbiasedRNG[397];
            InitCond[398] = UnbiasedRNG[398];
            InitCond[399] = UnbiasedRNG[399];
            InitCond[400] = UnbiasedRNG[400];
            InitCond[401] = UnbiasedRNG[401];
            InitCond[402] = UnbiasedRNG[402];
            InitCond[403] = UnbiasedRNG[403];
            InitCond[404] = UnbiasedRNG[404];
            InitCond[405] = UnbiasedRNG[405];
            InitCond[406] = UnbiasedRNG[406];
            InitCond[407] = UnbiasedRNG[407];
            InitCond[408] = UnbiasedRNG[408];
            InitCond[409] = UnbiasedRNG[409];
            InitCond[410] = UnbiasedRNG[410];
            InitCond[411] = UnbiasedRNG[411];
            InitCond[412] = UnbiasedRNG[412];
            InitCond[413] = UnbiasedRNG[413];
            InitCond[414] = UnbiasedRNG[414];
            InitCond[415] = UnbiasedRNG[415];
            InitCond[416] = UnbiasedRNG[416];
            InitCond[417] = UnbiasedRNG[417];
            InitCond[418] = UnbiasedRNG[418];
            InitCond[419] = UnbiasedRNG[419];
            InitCond[420] = UnbiasedRNG[420];
            InitCond[421] = UnbiasedRNG[421];
            InitCond[422] = UnbiasedRNG[422];
            InitCond[423] = UnbiasedRNG[423];
            InitCond[424] = UnbiasedRNG[424];
            InitCond[425] = UnbiasedRNG[425];
            InitCond[426] = UnbiasedRNG[426];
            InitCond[427] = UnbiasedRNG[427];
            InitCond[428] = UnbiasedRNG[428];
            InitCond[429] = UnbiasedRNG[429];
            InitCond[430] = UnbiasedRNG[430];
            InitCond[431] = UnbiasedRNG[431];
            InitCond[432] = UnbiasedRNG[432];
            InitCond[433] = UnbiasedRNG[433];
            InitCond[434] = UnbiasedRNG[434];
            InitCond[435] = UnbiasedRNG[435];
            InitCond[436] = UnbiasedRNG[436];
            InitCond[437] = UnbiasedRNG[437];
            InitCond[438] = UnbiasedRNG[438];
            InitCond[439] = UnbiasedRNG[439];
            InitCond[440] = UnbiasedRNG[440];
            InitCond[441] = UnbiasedRNG[441];
            InitCond[442] = UnbiasedRNG[442];
            InitCond[443] = UnbiasedRNG[443];
            InitCond[444] = UnbiasedRNG[444];
            InitCond[445] = UnbiasedRNG[445];
            InitCond[446] = UnbiasedRNG[446];
            InitCond[447] = UnbiasedRNG[447];
            InitCond[448] = UnbiasedRNG[448];
            InitCond[449] = UnbiasedRNG[449];
            InitCond[450] = UnbiasedRNG[450];
            InitCond[451] = UnbiasedRNG[451];
            InitCond[452] = UnbiasedRNG[452];
            InitCond[453] = UnbiasedRNG[453];
            InitCond[454] = UnbiasedRNG[454];
            InitCond[455] = UnbiasedRNG[455];
            InitCond[456] = UnbiasedRNG[456];
            InitCond[457] = UnbiasedRNG[457];
            InitCond[458] = UnbiasedRNG[458];
            InitCond[459] = UnbiasedRNG[459];
            InitCond[460] = UnbiasedRNG[460];
            InitCond[461] = UnbiasedRNG[461];
            InitCond[462] = UnbiasedRNG[462];
            InitCond[463] = UnbiasedRNG[463];
            InitCond[464] = UnbiasedRNG[464];
            InitCond[465] = UnbiasedRNG[465];
            InitCond[466] = UnbiasedRNG[466];
            InitCond[467] = UnbiasedRNG[467];
            InitCond[468] = UnbiasedRNG[468];
            InitCond[469] = UnbiasedRNG[469];
            InitCond[470] = UnbiasedRNG[470];
            InitCond[471] = UnbiasedRNG[471];
            InitCond[472] = UnbiasedRNG[472];
            InitCond[473] = UnbiasedRNG[473];
            InitCond[474] = UnbiasedRNG[474];
            InitCond[475] = UnbiasedRNG[475];
            InitCond[476] = UnbiasedRNG[476];
            InitCond[477] = UnbiasedRNG[477];
            InitCond[478] = UnbiasedRNG[478];
            InitCond[479] = UnbiasedRNG[479];
            InitCond[480] = UnbiasedRNG[480];
            InitCond[481] = UnbiasedRNG[481];
            InitCond[482] = UnbiasedRNG[482];
            InitCond[483] = UnbiasedRNG[483];
            InitCond[484] = UnbiasedRNG[484];
            InitCond[485] = UnbiasedRNG[485];
            InitCond[486] = UnbiasedRNG[486];
            InitCond[487] = UnbiasedRNG[487];
            InitCond[488] = UnbiasedRNG[488];
            InitCond[489] = UnbiasedRNG[489];
            InitCond[490] = UnbiasedRNG[490];
            InitCond[491] = UnbiasedRNG[491];
            InitCond[492] = UnbiasedRNG[492];
            InitCond[493] = UnbiasedRNG[493];
            InitCond[494] = UnbiasedRNG[494];
            InitCond[495] = UnbiasedRNG[495];
            InitCond[496] = UnbiasedRNG[496];
            InitCond[497] = UnbiasedRNG[497];
            InitCond[498] = UnbiasedRNG[498];
            InitCond[499] = UnbiasedRNG[499];
            InitCond[500] = UnbiasedRNG[500];
            InitCond[501] = UnbiasedRNG[501];
            InitCond[502] = UnbiasedRNG[502];
            InitCond[503] = UnbiasedRNG[503];
            InitCond[504] = UnbiasedRNG[504];
            InitCond[505] = UnbiasedRNG[505];
            InitCond[506] = UnbiasedRNG[506];
            InitCond[507] = UnbiasedRNG[507];
            InitCond[508] = UnbiasedRNG[508];
            InitCond[509] = UnbiasedRNG[509];
            InitCond[510] = UnbiasedRNG[510];
            InitCond[511] = UnbiasedRNG[511];
            InitCond[512] = UnbiasedRNG[512];
            InitCond[513] = UnbiasedRNG[513];
            InitCond[514] = UnbiasedRNG[514];
            InitCond[515] = UnbiasedRNG[515];
            InitCond[516] = UnbiasedRNG[516];
            InitCond[517] = UnbiasedRNG[517];
            InitCond[518] = UnbiasedRNG[518];
            InitCond[519] = UnbiasedRNG[519];
            InitCond[520] = UnbiasedRNG[520];
            InitCond[521] = UnbiasedRNG[521];
            InitCond[522] = UnbiasedRNG[522];
            InitCond[523] = UnbiasedRNG[523];
            InitCond[524] = UnbiasedRNG[524];
            InitCond[525] = UnbiasedRNG[525];
            InitCond[526] = UnbiasedRNG[526];
            InitCond[527] = UnbiasedRNG[527];
            InitCond[528] = UnbiasedRNG[528];
            InitCond[529] = UnbiasedRNG[529];
            InitCond[530] = UnbiasedRNG[530];
            InitCond[531] = UnbiasedRNG[531];
            InitCond[532] = UnbiasedRNG[532];
            InitCond[533] = UnbiasedRNG[533];
            InitCond[534] = UnbiasedRNG[534];
            InitCond[535] = UnbiasedRNG[535];
            InitCond[536] = UnbiasedRNG[536];
            InitCond[537] = UnbiasedRNG[537];
            InitCond[538] = UnbiasedRNG[538];
            InitCond[539] = UnbiasedRNG[539];
            InitCond[540] = UnbiasedRNG[540];
            InitCond[541] = UnbiasedRNG[541];
            InitCond[542] = UnbiasedRNG[542];
            InitCond[543] = UnbiasedRNG[543];
            InitCond[544] = UnbiasedRNG[544];
            InitCond[545] = UnbiasedRNG[545];
            InitCond[546] = UnbiasedRNG[546];
            InitCond[547] = UnbiasedRNG[547];
            InitCond[548] = UnbiasedRNG[548];
            InitCond[549] = UnbiasedRNG[549];
            InitCond[550] = UnbiasedRNG[550];
            InitCond[551] = UnbiasedRNG[551];
            InitCond[552] = UnbiasedRNG[552];
            InitCond[553] = UnbiasedRNG[553];
            InitCond[554] = UnbiasedRNG[554];
            InitCond[555] = UnbiasedRNG[555];
            InitCond[556] = UnbiasedRNG[556];
            InitCond[557] = UnbiasedRNG[557];
            InitCond[558] = UnbiasedRNG[558];
            InitCond[559] = UnbiasedRNG[559];
            InitCond[560] = UnbiasedRNG[560];
            InitCond[561] = UnbiasedRNG[561];
            InitCond[562] = UnbiasedRNG[562];
            InitCond[563] = UnbiasedRNG[563];
            InitCond[564] = UnbiasedRNG[564];
            InitCond[565] = UnbiasedRNG[565];
            InitCond[566] = UnbiasedRNG[566];
            InitCond[567] = UnbiasedRNG[567];
            InitCond[568] = UnbiasedRNG[568];
            InitCond[569] = UnbiasedRNG[569];
            InitCond[570] = UnbiasedRNG[570];
            InitCond[571] = UnbiasedRNG[571];
            InitCond[572] = UnbiasedRNG[572];
            InitCond[573] = UnbiasedRNG[573];
            InitCond[574] = UnbiasedRNG[574];
            InitCond[575] = UnbiasedRNG[575];
            InitCond[576] = UnbiasedRNG[576];
            InitCond[577] = UnbiasedRNG[577];
            InitCond[578] = UnbiasedRNG[578];
            InitCond[579] = UnbiasedRNG[579];
            InitCond[580] = UnbiasedRNG[580];
            InitCond[581] = UnbiasedRNG[581];
            InitCond[582] = UnbiasedRNG[582];
            InitCond[583] = UnbiasedRNG[583];
            InitCond[584] = UnbiasedRNG[584];
            InitCond[585] = UnbiasedRNG[585];
            InitCond[586] = UnbiasedRNG[586];
            InitCond[587] = UnbiasedRNG[587];
            InitCond[588] = UnbiasedRNG[588];
            InitCond[589] = UnbiasedRNG[589];
            InitCond[590] = UnbiasedRNG[590];
            InitCond[591] = UnbiasedRNG[591];
            InitCond[592] = UnbiasedRNG[592];
            InitCond[593] = UnbiasedRNG[593];
            InitCond[594] = UnbiasedRNG[594];
            InitCond[595] = UnbiasedRNG[595];
            InitCond[596] = UnbiasedRNG[596];
            InitCond[597] = UnbiasedRNG[597];
            InitCond[598] = UnbiasedRNG[598];
            InitCond[599] = UnbiasedRNG[599];
            InitCond[600] = UnbiasedRNG[600];
            InitCond[601] = UnbiasedRNG[601];
            InitCond[602] = UnbiasedRNG[602];
            InitCond[603] = UnbiasedRNG[603];
            InitCond[604] = UnbiasedRNG[604];
            InitCond[605] = UnbiasedRNG[605];
            InitCond[606] = UnbiasedRNG[606];
            InitCond[607] = UnbiasedRNG[607];
            InitCond[608] = UnbiasedRNG[608];
            InitCond[609] = UnbiasedRNG[609];
            InitCond[610] = UnbiasedRNG[610];
            InitCond[611] = UnbiasedRNG[611];
            InitCond[612] = UnbiasedRNG[612];
            InitCond[613] = UnbiasedRNG[613];
            InitCond[614] = UnbiasedRNG[614];
            InitCond[615] = UnbiasedRNG[615];
            InitCond[616] = UnbiasedRNG[616];
            InitCond[617] = UnbiasedRNG[617];
            InitCond[618] = UnbiasedRNG[618];
            InitCond[619] = UnbiasedRNG[619];
            InitCond[620] = UnbiasedRNG[620];
            InitCond[621] = UnbiasedRNG[621];
            InitCond[622] = UnbiasedRNG[622];
            InitCond[623] = UnbiasedRNG[623];
            InitCond[624] = UnbiasedRNG[624];
            InitCond[625] = UnbiasedRNG[625];
            InitCond[626] = UnbiasedRNG[626];
            InitCond[627] = UnbiasedRNG[627];
            InitCond[628] = UnbiasedRNG[628];
            InitCond[629] = UnbiasedRNG[629];
            InitCond[630] = UnbiasedRNG[630];
            InitCond[631] = UnbiasedRNG[631];
            InitCond[632] = UnbiasedRNG[632];
            InitCond[633] = UnbiasedRNG[633];
            InitCond[634] = UnbiasedRNG[634];
            InitCond[635] = UnbiasedRNG[635];
            InitCond[636] = UnbiasedRNG[636];
            InitCond[637] = UnbiasedRNG[637];
            InitCond[638] = UnbiasedRNG[638];
            InitCond[639] = UnbiasedRNG[639];
            InitCond[640] = UnbiasedRNG[640];
            InitCond[641] = UnbiasedRNG[641];
            InitCond[642] = UnbiasedRNG[642];
            InitCond[643] = UnbiasedRNG[643];
            InitCond[644] = UnbiasedRNG[644];
            InitCond[645] = UnbiasedRNG[645];
            InitCond[646] = UnbiasedRNG[646];
            InitCond[647] = UnbiasedRNG[647];
            InitCond[648] = UnbiasedRNG[648];
            InitCond[649] = UnbiasedRNG[649];
            InitCond[650] = UnbiasedRNG[650];
            InitCond[651] = UnbiasedRNG[651];
            InitCond[652] = UnbiasedRNG[652];
            InitCond[653] = UnbiasedRNG[653];
            InitCond[654] = UnbiasedRNG[654];
            InitCond[655] = UnbiasedRNG[655];
            InitCond[656] = UnbiasedRNG[656];
            InitCond[657] = UnbiasedRNG[657];
            InitCond[658] = UnbiasedRNG[658];
            InitCond[659] = UnbiasedRNG[659];
            InitCond[660] = UnbiasedRNG[660];
            InitCond[661] = UnbiasedRNG[661];
            InitCond[662] = UnbiasedRNG[662];
            InitCond[663] = UnbiasedRNG[663];
            InitCond[664] = UnbiasedRNG[664];
            InitCond[665] = UnbiasedRNG[665];
            InitCond[666] = UnbiasedRNG[666];
            InitCond[667] = UnbiasedRNG[667];
            InitCond[668] = UnbiasedRNG[668];
            InitCond[669] = UnbiasedRNG[669];
            InitCond[670] = UnbiasedRNG[670];
            InitCond[671] = UnbiasedRNG[671];
            InitCond[672] = UnbiasedRNG[672];
            InitCond[673] = UnbiasedRNG[673];
            InitCond[674] = UnbiasedRNG[674];
            InitCond[675] = UnbiasedRNG[675];
            InitCond[676] = UnbiasedRNG[676];
            InitCond[677] = UnbiasedRNG[677];
            InitCond[678] = UnbiasedRNG[678];
            InitCond[679] = UnbiasedRNG[679];
            InitCond[680] = UnbiasedRNG[680];
            InitCond[681] = UnbiasedRNG[681];
            InitCond[682] = UnbiasedRNG[682];
            InitCond[683] = UnbiasedRNG[683];
            InitCond[684] = UnbiasedRNG[684];
            InitCond[685] = UnbiasedRNG[685];
            InitCond[686] = UnbiasedRNG[686];
            InitCond[687] = UnbiasedRNG[687];
            InitCond[688] = UnbiasedRNG[688];
            InitCond[689] = UnbiasedRNG[689];
            InitCond[690] = UnbiasedRNG[690];
            InitCond[691] = UnbiasedRNG[691];
            InitCond[692] = UnbiasedRNG[692];
            InitCond[693] = UnbiasedRNG[693];
            InitCond[694] = UnbiasedRNG[694];
            InitCond[695] = UnbiasedRNG[695];
            InitCond[696] = UnbiasedRNG[696];
            InitCond[697] = UnbiasedRNG[697];
            InitCond[698] = UnbiasedRNG[698];
            InitCond[699] = UnbiasedRNG[699];
            InitCond[700] = UnbiasedRNG[700];
            InitCond[701] = UnbiasedRNG[701];
            InitCond[702] = UnbiasedRNG[702];
            InitCond[703] = UnbiasedRNG[703];
            InitCond[704] = UnbiasedRNG[704];
            InitCond[705] = UnbiasedRNG[705];
            InitCond[706] = UnbiasedRNG[706];
            InitCond[707] = UnbiasedRNG[707];
            InitCond[708] = UnbiasedRNG[708];
            InitCond[709] = UnbiasedRNG[709];
            InitCond[710] = UnbiasedRNG[710];
            InitCond[711] = UnbiasedRNG[711];
            InitCond[712] = UnbiasedRNG[712];
            InitCond[713] = UnbiasedRNG[713];
            InitCond[714] = UnbiasedRNG[714];
            InitCond[715] = UnbiasedRNG[715];
        end
        else if (counter == 2) begin
            InitCond[716] = UnbiasedRNG[0];
            InitCond[717] = UnbiasedRNG[1];
            InitCond[718] = UnbiasedRNG[2];
            InitCond[719] = UnbiasedRNG[3];
            InitCond[720] = UnbiasedRNG[4];
            InitCond[721] = UnbiasedRNG[5];
            InitCond[722] = UnbiasedRNG[6];
            InitCond[723] = UnbiasedRNG[7];
            InitCond[724] = UnbiasedRNG[8];
            InitCond[725] = UnbiasedRNG[9];
            InitCond[726] = UnbiasedRNG[10];
            InitCond[727] = UnbiasedRNG[11];
            InitCond[728] = UnbiasedRNG[12];
            InitCond[729] = UnbiasedRNG[13];
            InitCond[730] = UnbiasedRNG[14];
            InitCond[731] = UnbiasedRNG[15];
            InitCond[732] = UnbiasedRNG[16];
            InitCond[733] = UnbiasedRNG[17];
            InitCond[734] = UnbiasedRNG[18];
            InitCond[735] = UnbiasedRNG[19];
            InitCond[736] = UnbiasedRNG[20];
            InitCond[737] = UnbiasedRNG[21];
            InitCond[738] = UnbiasedRNG[22];
            InitCond[739] = UnbiasedRNG[23];
            InitCond[740] = UnbiasedRNG[24];
            InitCond[741] = UnbiasedRNG[25];
            InitCond[742] = UnbiasedRNG[26];
            InitCond[743] = UnbiasedRNG[27];
            InitCond[744] = UnbiasedRNG[28];
            InitCond[745] = UnbiasedRNG[29];
            InitCond[746] = UnbiasedRNG[30];
            InitCond[747] = UnbiasedRNG[31];
            InitCond[748] = UnbiasedRNG[32];
            InitCond[749] = UnbiasedRNG[33];
            InitCond[750] = UnbiasedRNG[34];
            InitCond[751] = UnbiasedRNG[35];
            InitCond[752] = UnbiasedRNG[36];
            InitCond[753] = UnbiasedRNG[37];
            InitCond[754] = UnbiasedRNG[38];
            InitCond[755] = UnbiasedRNG[39];
            InitCond[756] = UnbiasedRNG[40];
            InitCond[757] = UnbiasedRNG[41];
            InitCond[758] = UnbiasedRNG[42];
            InitCond[759] = UnbiasedRNG[43];
            InitCond[760] = UnbiasedRNG[44];
            InitCond[761] = UnbiasedRNG[45];
            InitCond[762] = UnbiasedRNG[46];
            InitCond[763] = UnbiasedRNG[47];
            InitCond[764] = UnbiasedRNG[48];
            InitCond[765] = UnbiasedRNG[49];
            InitCond[766] = UnbiasedRNG[50];
            InitCond[767] = UnbiasedRNG[51];
            InitCond[768] = UnbiasedRNG[52];
            InitCond[769] = UnbiasedRNG[53];
            InitCond[770] = UnbiasedRNG[54];
            InitCond[771] = UnbiasedRNG[55];
            InitCond[772] = UnbiasedRNG[56];
            InitCond[773] = UnbiasedRNG[57];
            InitCond[774] = UnbiasedRNG[58];
            InitCond[775] = UnbiasedRNG[59];
            InitCond[776] = UnbiasedRNG[60];
            InitCond[777] = UnbiasedRNG[61];
            InitCond[778] = UnbiasedRNG[62];
            InitCond[779] = UnbiasedRNG[63];
            InitCond[780] = UnbiasedRNG[64];
            InitCond[781] = UnbiasedRNG[65];
            InitCond[782] = UnbiasedRNG[66];
            InitCond[783] = UnbiasedRNG[67];
            InitCond[784] = UnbiasedRNG[68];
            InitCond[785] = UnbiasedRNG[69];
            InitCond[786] = UnbiasedRNG[70];
            InitCond[787] = UnbiasedRNG[71];
            InitCond[788] = UnbiasedRNG[72];
            InitCond[789] = UnbiasedRNG[73];
            InitCond[790] = UnbiasedRNG[74];
            InitCond[791] = UnbiasedRNG[75];
            InitCond[792] = UnbiasedRNG[76];
            InitCond[793] = UnbiasedRNG[77];
            InitCond[794] = UnbiasedRNG[78];
            InitCond[795] = UnbiasedRNG[79];
            InitCond[796] = UnbiasedRNG[80];
            InitCond[797] = UnbiasedRNG[81];
            InitCond[798] = UnbiasedRNG[82];
            InitCond[799] = UnbiasedRNG[83];
            InitCond[800] = UnbiasedRNG[84];
            InitCond[801] = UnbiasedRNG[85];
            InitCond[802] = UnbiasedRNG[86];
            InitCond[803] = UnbiasedRNG[87];
            InitCond[804] = UnbiasedRNG[88];
            InitCond[805] = UnbiasedRNG[89];
            InitCond[806] = UnbiasedRNG[90];
            InitCond[807] = UnbiasedRNG[91];
            InitCond[808] = UnbiasedRNG[92];
            InitCond[809] = UnbiasedRNG[93];
            InitCond[810] = UnbiasedRNG[94];
            InitCond[811] = UnbiasedRNG[95];
            InitCond[812] = UnbiasedRNG[96];
            InitCond[813] = UnbiasedRNG[97];
            InitCond[814] = UnbiasedRNG[98];
            InitCond[815] = UnbiasedRNG[99];
            InitCond[816] = UnbiasedRNG[100];
            InitCond[817] = UnbiasedRNG[101];
            InitCond[818] = UnbiasedRNG[102];
            InitCond[819] = UnbiasedRNG[103];
            InitCond[820] = UnbiasedRNG[104];
            InitCond[821] = UnbiasedRNG[105];
            InitCond[822] = UnbiasedRNG[106];
            InitCond[823] = UnbiasedRNG[107];
            InitCond[824] = UnbiasedRNG[108];
            InitCond[825] = UnbiasedRNG[109];
            InitCond[826] = UnbiasedRNG[110];
            InitCond[827] = UnbiasedRNG[111];
            InitCond[828] = UnbiasedRNG[112];
            InitCond[829] = UnbiasedRNG[113];
            InitCond[830] = UnbiasedRNG[114];
            InitCond[831] = UnbiasedRNG[115];
            InitCond[832] = UnbiasedRNG[116];
            InitCond[833] = UnbiasedRNG[117];
            InitCond[834] = UnbiasedRNG[118];
            InitCond[835] = UnbiasedRNG[119];
            InitCond[836] = UnbiasedRNG[120];
            InitCond[837] = UnbiasedRNG[121];
            InitCond[838] = UnbiasedRNG[122];
            InitCond[839] = UnbiasedRNG[123];
            InitCond[840] = UnbiasedRNG[124];
            InitCond[841] = UnbiasedRNG[125];
            InitCond[842] = UnbiasedRNG[126];
            InitCond[843] = UnbiasedRNG[127];
            InitCond[844] = UnbiasedRNG[128];
            InitCond[845] = UnbiasedRNG[129];
            InitCond[846] = UnbiasedRNG[130];
            InitCond[847] = UnbiasedRNG[131];
            InitCond[848] = UnbiasedRNG[132];
            InitCond[849] = UnbiasedRNG[133];
            InitCond[850] = UnbiasedRNG[134];
            InitCond[851] = UnbiasedRNG[135];
            InitCond[852] = UnbiasedRNG[136];
            InitCond[853] = UnbiasedRNG[137];
            InitCond[854] = UnbiasedRNG[138];
            InitCond[855] = UnbiasedRNG[139];
            InitCond[856] = UnbiasedRNG[140];
            InitCond[857] = UnbiasedRNG[141];
            InitCond[858] = UnbiasedRNG[142];
            InitCond[859] = UnbiasedRNG[143];
            InitCond[860] = UnbiasedRNG[144];
            InitCond[861] = UnbiasedRNG[145];
            InitCond[862] = UnbiasedRNG[146];
            InitCond[863] = UnbiasedRNG[147];
            InitCond[864] = UnbiasedRNG[148];
            InitCond[865] = UnbiasedRNG[149];
            InitCond[866] = UnbiasedRNG[150];
            InitCond[867] = UnbiasedRNG[151];
            InitCond[868] = UnbiasedRNG[152];
            InitCond[869] = UnbiasedRNG[153];
            InitCond[870] = UnbiasedRNG[154];
            InitCond[871] = UnbiasedRNG[155];
            InitCond[872] = UnbiasedRNG[156];
            InitCond[873] = UnbiasedRNG[157];
            InitCond[874] = UnbiasedRNG[158];
            InitCond[875] = UnbiasedRNG[159];
            InitCond[876] = UnbiasedRNG[160];
            InitCond[877] = UnbiasedRNG[161];
            InitCond[878] = UnbiasedRNG[162];
            InitCond[879] = UnbiasedRNG[163];
            InitCond[880] = UnbiasedRNG[164];
            InitCond[881] = UnbiasedRNG[165];
            InitCond[882] = UnbiasedRNG[166];
            InitCond[883] = UnbiasedRNG[167];
            InitCond[884] = UnbiasedRNG[168];
            InitCond[885] = UnbiasedRNG[169];
            InitCond[886] = UnbiasedRNG[170];
            InitCond[887] = UnbiasedRNG[171];
            InitCond[888] = UnbiasedRNG[172];
            InitCond[889] = UnbiasedRNG[173];
            InitCond[890] = UnbiasedRNG[174];
            InitCond[891] = UnbiasedRNG[175];
            InitCond[892] = UnbiasedRNG[176];
            InitCond[893] = UnbiasedRNG[177];
            InitCond[894] = UnbiasedRNG[178];
            InitCond[895] = UnbiasedRNG[179];
            InitCond[896] = UnbiasedRNG[180];
            InitCond[897] = UnbiasedRNG[181];
            InitCond[898] = UnbiasedRNG[182];
            InitCond[899] = UnbiasedRNG[183];
            InitCond[900] = UnbiasedRNG[184];
            InitCond[901] = UnbiasedRNG[185];
            InitCond[902] = UnbiasedRNG[186];
            InitCond[903] = UnbiasedRNG[187];
            InitCond[904] = UnbiasedRNG[188];
            InitCond[905] = UnbiasedRNG[189];
            InitCond[906] = UnbiasedRNG[190];
            InitCond[907] = UnbiasedRNG[191];
            InitCond[908] = UnbiasedRNG[192];
            InitCond[909] = UnbiasedRNG[193];
            InitCond[910] = UnbiasedRNG[194];
            InitCond[911] = UnbiasedRNG[195];
            InitCond[912] = UnbiasedRNG[196];
            InitCond[913] = UnbiasedRNG[197];
            InitCond[914] = UnbiasedRNG[198];
            InitCond[915] = UnbiasedRNG[199];
            InitCond[916] = UnbiasedRNG[200];
            InitCond[917] = UnbiasedRNG[201];
            InitCond[918] = UnbiasedRNG[202];
            InitCond[919] = UnbiasedRNG[203];
            InitCond[920] = UnbiasedRNG[204];
            InitCond[921] = UnbiasedRNG[205];
            InitCond[922] = UnbiasedRNG[206];
            InitCond[923] = UnbiasedRNG[207];
            InitCond[924] = UnbiasedRNG[208];
            InitCond[925] = UnbiasedRNG[209];
            InitCond[926] = UnbiasedRNG[210];
            InitCond[927] = UnbiasedRNG[211];
            InitCond[928] = UnbiasedRNG[212];
            InitCond[929] = UnbiasedRNG[213];
            InitCond[930] = UnbiasedRNG[214];
            InitCond[931] = UnbiasedRNG[215];
            InitCond[932] = UnbiasedRNG[216];
            InitCond[933] = UnbiasedRNG[217];
            InitCond[934] = UnbiasedRNG[218];
            InitCond[935] = UnbiasedRNG[219];
            InitCond[936] = UnbiasedRNG[220];
            InitCond[937] = UnbiasedRNG[221];
            InitCond[938] = UnbiasedRNG[222];
            InitCond[939] = UnbiasedRNG[223];
            InitCond[940] = UnbiasedRNG[224];
            InitCond[941] = UnbiasedRNG[225];
            InitCond[942] = UnbiasedRNG[226];
            InitCond[943] = UnbiasedRNG[227];
            InitCond[944] = UnbiasedRNG[228];
            InitCond[945] = UnbiasedRNG[229];
            InitCond[946] = UnbiasedRNG[230];
            InitCond[947] = UnbiasedRNG[231];
            InitCond[948] = UnbiasedRNG[232];
            InitCond[949] = UnbiasedRNG[233];
            InitCond[950] = UnbiasedRNG[234];
            InitCond[951] = UnbiasedRNG[235];
            InitCond[952] = UnbiasedRNG[236];
            InitCond[953] = UnbiasedRNG[237];
            InitCond[954] = UnbiasedRNG[238];
            InitCond[955] = UnbiasedRNG[239];
            InitCond[956] = UnbiasedRNG[240];
            InitCond[957] = UnbiasedRNG[241];
            InitCond[958] = UnbiasedRNG[242];
            InitCond[959] = UnbiasedRNG[243];
            InitCond[960] = UnbiasedRNG[244];
            InitCond[961] = UnbiasedRNG[245];
            InitCond[962] = UnbiasedRNG[246];
            InitCond[963] = UnbiasedRNG[247];
            InitCond[964] = UnbiasedRNG[248];
            InitCond[965] = UnbiasedRNG[249];
            InitCond[966] = UnbiasedRNG[250];
            InitCond[967] = UnbiasedRNG[251];
            InitCond[968] = UnbiasedRNG[252];
            InitCond[969] = UnbiasedRNG[253];
            InitCond[970] = UnbiasedRNG[254];
            InitCond[971] = UnbiasedRNG[255];
            InitCond[972] = UnbiasedRNG[256];
            InitCond[973] = UnbiasedRNG[257];
            InitCond[974] = UnbiasedRNG[258];
            InitCond[975] = UnbiasedRNG[259];
            InitCond[976] = UnbiasedRNG[260];
            InitCond[977] = UnbiasedRNG[261];
            InitCond[978] = UnbiasedRNG[262];
            InitCond[979] = UnbiasedRNG[263];
            InitCond[980] = UnbiasedRNG[264];
            InitCond[981] = UnbiasedRNG[265];
            InitCond[982] = UnbiasedRNG[266];
            InitCond[983] = UnbiasedRNG[267];
            InitCond[984] = UnbiasedRNG[268];
            InitCond[985] = UnbiasedRNG[269];
            InitCond[986] = UnbiasedRNG[270];
            InitCond[987] = UnbiasedRNG[271];
            InitCond[988] = UnbiasedRNG[272];
            InitCond[989] = UnbiasedRNG[273];
            InitCond[990] = UnbiasedRNG[274];
            InitCond[991] = UnbiasedRNG[275];
            InitCond[992] = UnbiasedRNG[276];
            InitCond[993] = UnbiasedRNG[277];
            InitCond[994] = UnbiasedRNG[278];
            InitCond[995] = UnbiasedRNG[279];
            InitCond[996] = UnbiasedRNG[280];
            InitCond[997] = UnbiasedRNG[281];
            InitCond[998] = UnbiasedRNG[282];
            InitCond[999] = UnbiasedRNG[283];
            InitCond[1000] = UnbiasedRNG[284];
            InitCond[1001] = UnbiasedRNG[285];
            InitCond[1002] = UnbiasedRNG[286];
            InitCond[1003] = UnbiasedRNG[287];
            InitCond[1004] = UnbiasedRNG[288];
            InitCond[1005] = UnbiasedRNG[289];
            InitCond[1006] = UnbiasedRNG[290];
            InitCond[1007] = UnbiasedRNG[291];
            InitCond[1008] = UnbiasedRNG[292];
            InitCond[1009] = UnbiasedRNG[293];
            InitCond[1010] = UnbiasedRNG[294];
            InitCond[1011] = UnbiasedRNG[295];
            InitCond[1012] = UnbiasedRNG[296];
            InitCond[1013] = UnbiasedRNG[297];
            InitCond[1014] = UnbiasedRNG[298];
            InitCond[1015] = UnbiasedRNG[299];
            InitCond[1016] = UnbiasedRNG[300];
            InitCond[1017] = UnbiasedRNG[301];
            InitCond[1018] = UnbiasedRNG[302];
            InitCond[1019] = UnbiasedRNG[303];
            InitCond[1020] = UnbiasedRNG[304];
            InitCond[1021] = UnbiasedRNG[305];
            InitCond[1022] = UnbiasedRNG[306];
            InitCond[1023] = UnbiasedRNG[307];
            InitCond[1024] = UnbiasedRNG[308];
            InitCond[1025] = UnbiasedRNG[309];
            InitCond[1026] = UnbiasedRNG[310];
            InitCond[1027] = UnbiasedRNG[311];
            InitCond[1028] = UnbiasedRNG[312];
            InitCond[1029] = UnbiasedRNG[313];
            InitCond[1030] = UnbiasedRNG[314];
            InitCond[1031] = UnbiasedRNG[315];
            InitCond[1032] = UnbiasedRNG[316];
            InitCond[1033] = UnbiasedRNG[317];
            InitCond[1034] = UnbiasedRNG[318];
            InitCond[1035] = UnbiasedRNG[319];
            InitCond[1036] = UnbiasedRNG[320];
            InitCond[1037] = UnbiasedRNG[321];
            InitCond[1038] = UnbiasedRNG[322];
            InitCond[1039] = UnbiasedRNG[323];
            InitCond[1040] = UnbiasedRNG[324];
            InitCond[1041] = UnbiasedRNG[325];
            InitCond[1042] = UnbiasedRNG[326];
            InitCond[1043] = UnbiasedRNG[327];
            InitCond[1044] = UnbiasedRNG[328];
            InitCond[1045] = UnbiasedRNG[329];
            InitCond[1046] = UnbiasedRNG[330];
            InitCond[1047] = UnbiasedRNG[331];
            InitCond[1048] = UnbiasedRNG[332];
            InitCond[1049] = UnbiasedRNG[333];
            InitCond[1050] = UnbiasedRNG[334];
            InitCond[1051] = UnbiasedRNG[335];
            InitCond[1052] = UnbiasedRNG[336];
            InitCond[1053] = UnbiasedRNG[337];
            InitCond[1054] = UnbiasedRNG[338];
            InitCond[1055] = UnbiasedRNG[339];
            InitCond[1056] = UnbiasedRNG[340];
            InitCond[1057] = UnbiasedRNG[341];
            InitCond[1058] = UnbiasedRNG[342];
            InitCond[1059] = UnbiasedRNG[343];
            InitCond[1060] = UnbiasedRNG[344];
            InitCond[1061] = UnbiasedRNG[345];
            InitCond[1062] = UnbiasedRNG[346];
            InitCond[1063] = UnbiasedRNG[347];
            InitCond[1064] = UnbiasedRNG[348];
            InitCond[1065] = UnbiasedRNG[349];
            InitCond[1066] = UnbiasedRNG[350];
            InitCond[1067] = UnbiasedRNG[351];
            InitCond[1068] = UnbiasedRNG[352];
            InitCond[1069] = UnbiasedRNG[353];
            InitCond[1070] = UnbiasedRNG[354];
            InitCond[1071] = UnbiasedRNG[355];
            InitCond[1072] = UnbiasedRNG[356];
            InitCond[1073] = UnbiasedRNG[357];
            InitCond[1074] = UnbiasedRNG[358];
            InitCond[1075] = UnbiasedRNG[359];
            InitCond[1076] = UnbiasedRNG[360];
            InitCond[1077] = UnbiasedRNG[361];
            InitCond[1078] = UnbiasedRNG[362];
            InitCond[1079] = UnbiasedRNG[363];
            InitCond[1080] = UnbiasedRNG[364];
            InitCond[1081] = UnbiasedRNG[365];
            InitCond[1082] = UnbiasedRNG[366];
            InitCond[1083] = UnbiasedRNG[367];
            InitCond[1084] = UnbiasedRNG[368];
            InitCond[1085] = UnbiasedRNG[369];
            InitCond[1086] = UnbiasedRNG[370];
            InitCond[1087] = UnbiasedRNG[371];
            InitCond[1088] = UnbiasedRNG[372];
            InitCond[1089] = UnbiasedRNG[373];
            InitCond[1090] = UnbiasedRNG[374];
            InitCond[1091] = UnbiasedRNG[375];
            InitCond[1092] = UnbiasedRNG[376];
            InitCond[1093] = UnbiasedRNG[377];
            InitCond[1094] = UnbiasedRNG[378];
            InitCond[1095] = UnbiasedRNG[379];
            InitCond[1096] = UnbiasedRNG[380];
            InitCond[1097] = UnbiasedRNG[381];
            InitCond[1098] = UnbiasedRNG[382];
            InitCond[1099] = UnbiasedRNG[383];
            InitCond[1100] = UnbiasedRNG[384];
            InitCond[1101] = UnbiasedRNG[385];
            InitCond[1102] = UnbiasedRNG[386];
            InitCond[1103] = UnbiasedRNG[387];
            InitCond[1104] = UnbiasedRNG[388];
            InitCond[1105] = UnbiasedRNG[389];
            InitCond[1106] = UnbiasedRNG[390];
            InitCond[1107] = UnbiasedRNG[391];
            InitCond[1108] = UnbiasedRNG[392];
            InitCond[1109] = UnbiasedRNG[393];
            InitCond[1110] = UnbiasedRNG[394];
            InitCond[1111] = UnbiasedRNG[395];
            InitCond[1112] = UnbiasedRNG[396];
            InitCond[1113] = UnbiasedRNG[397];
            InitCond[1114] = UnbiasedRNG[398];
            InitCond[1115] = UnbiasedRNG[399];
            InitCond[1116] = UnbiasedRNG[400];
            InitCond[1117] = UnbiasedRNG[401];
            InitCond[1118] = UnbiasedRNG[402];
            InitCond[1119] = UnbiasedRNG[403];
            InitCond[1120] = UnbiasedRNG[404];
            InitCond[1121] = UnbiasedRNG[405];
            InitCond[1122] = UnbiasedRNG[406];
            InitCond[1123] = UnbiasedRNG[407];
            InitCond[1124] = UnbiasedRNG[408];
            InitCond[1125] = UnbiasedRNG[409];
            InitCond[1126] = UnbiasedRNG[410];
            InitCond[1127] = UnbiasedRNG[411];
            InitCond[1128] = UnbiasedRNG[412];
            InitCond[1129] = UnbiasedRNG[413];
            InitCond[1130] = UnbiasedRNG[414];
            InitCond[1131] = UnbiasedRNG[415];
            InitCond[1132] = UnbiasedRNG[416];
            InitCond[1133] = UnbiasedRNG[417];
            InitCond[1134] = UnbiasedRNG[418];
            InitCond[1135] = UnbiasedRNG[419];
            InitCond[1136] = UnbiasedRNG[420];
            InitCond[1137] = UnbiasedRNG[421];
            InitCond[1138] = UnbiasedRNG[422];
            InitCond[1139] = UnbiasedRNG[423];
            InitCond[1140] = UnbiasedRNG[424];
            InitCond[1141] = UnbiasedRNG[425];
            InitCond[1142] = UnbiasedRNG[426];
            InitCond[1143] = UnbiasedRNG[427];
            InitCond[1144] = UnbiasedRNG[428];
            InitCond[1145] = UnbiasedRNG[429];
            InitCond[1146] = UnbiasedRNG[430];
            InitCond[1147] = UnbiasedRNG[431];
            InitCond[1148] = UnbiasedRNG[432];
            InitCond[1149] = UnbiasedRNG[433];
            InitCond[1150] = UnbiasedRNG[434];
            InitCond[1151] = UnbiasedRNG[435];
            InitCond[1152] = UnbiasedRNG[436];
            InitCond[1153] = UnbiasedRNG[437];
            InitCond[1154] = UnbiasedRNG[438];
            InitCond[1155] = UnbiasedRNG[439];
            InitCond[1156] = UnbiasedRNG[440];
            InitCond[1157] = UnbiasedRNG[441];
            InitCond[1158] = UnbiasedRNG[442];
            InitCond[1159] = UnbiasedRNG[443];
            InitCond[1160] = UnbiasedRNG[444];
            InitCond[1161] = UnbiasedRNG[445];
            InitCond[1162] = UnbiasedRNG[446];
            InitCond[1163] = UnbiasedRNG[447];
            InitCond[1164] = UnbiasedRNG[448];
            InitCond[1165] = UnbiasedRNG[449];
            InitCond[1166] = UnbiasedRNG[450];
            InitCond[1167] = UnbiasedRNG[451];
            InitCond[1168] = UnbiasedRNG[452];
            InitCond[1169] = UnbiasedRNG[453];
            InitCond[1170] = UnbiasedRNG[454];
            InitCond[1171] = UnbiasedRNG[455];
            InitCond[1172] = UnbiasedRNG[456];
            InitCond[1173] = UnbiasedRNG[457];
            InitCond[1174] = UnbiasedRNG[458];
            InitCond[1175] = UnbiasedRNG[459];
            InitCond[1176] = UnbiasedRNG[460];
            InitCond[1177] = UnbiasedRNG[461];
            InitCond[1178] = UnbiasedRNG[462];
            InitCond[1179] = UnbiasedRNG[463];
            InitCond[1180] = UnbiasedRNG[464];
            InitCond[1181] = UnbiasedRNG[465];
            InitCond[1182] = UnbiasedRNG[466];
            InitCond[1183] = UnbiasedRNG[467];
            InitCond[1184] = UnbiasedRNG[468];
            InitCond[1185] = UnbiasedRNG[469];
            InitCond[1186] = UnbiasedRNG[470];
            InitCond[1187] = UnbiasedRNG[471];
            InitCond[1188] = UnbiasedRNG[472];
            InitCond[1189] = UnbiasedRNG[473];
            InitCond[1190] = UnbiasedRNG[474];
            InitCond[1191] = UnbiasedRNG[475];
            InitCond[1192] = UnbiasedRNG[476];
            InitCond[1193] = UnbiasedRNG[477];
            InitCond[1194] = UnbiasedRNG[478];
            InitCond[1195] = UnbiasedRNG[479];
            InitCond[1196] = UnbiasedRNG[480];
            InitCond[1197] = UnbiasedRNG[481];
            InitCond[1198] = UnbiasedRNG[482];
            InitCond[1199] = UnbiasedRNG[483];
            InitCond[1200] = UnbiasedRNG[484];
            InitCond[1201] = UnbiasedRNG[485];
            InitCond[1202] = UnbiasedRNG[486];
            InitCond[1203] = UnbiasedRNG[487];
            InitCond[1204] = UnbiasedRNG[488];
            InitCond[1205] = UnbiasedRNG[489];
            InitCond[1206] = UnbiasedRNG[490];
            InitCond[1207] = UnbiasedRNG[491];
            InitCond[1208] = UnbiasedRNG[492];
            InitCond[1209] = UnbiasedRNG[493];
            InitCond[1210] = UnbiasedRNG[494];
            InitCond[1211] = UnbiasedRNG[495];
            InitCond[1212] = UnbiasedRNG[496];
            InitCond[1213] = UnbiasedRNG[497];
            InitCond[1214] = UnbiasedRNG[498];
            InitCond[1215] = UnbiasedRNG[499];
            InitCond[1216] = UnbiasedRNG[500];
            InitCond[1217] = UnbiasedRNG[501];
            InitCond[1218] = UnbiasedRNG[502];
            InitCond[1219] = UnbiasedRNG[503];
            InitCond[1220] = UnbiasedRNG[504];
            InitCond[1221] = UnbiasedRNG[505];
            InitCond[1222] = UnbiasedRNG[506];
            InitCond[1223] = UnbiasedRNG[507];
            InitCond[1224] = UnbiasedRNG[508];
            InitCond[1225] = UnbiasedRNG[509];
            InitCond[1226] = UnbiasedRNG[510];
            InitCond[1227] = UnbiasedRNG[511];
            InitCond[1228] = UnbiasedRNG[512];
            InitCond[1229] = UnbiasedRNG[513];
            InitCond[1230] = UnbiasedRNG[514];
            InitCond[1231] = UnbiasedRNG[515];
            InitCond[1232] = UnbiasedRNG[516];
            InitCond[1233] = UnbiasedRNG[517];
            InitCond[1234] = UnbiasedRNG[518];
            InitCond[1235] = UnbiasedRNG[519];
            InitCond[1236] = UnbiasedRNG[520];
            InitCond[1237] = UnbiasedRNG[521];
            InitCond[1238] = UnbiasedRNG[522];
            InitCond[1239] = UnbiasedRNG[523];
            InitCond[1240] = UnbiasedRNG[524];
            InitCond[1241] = UnbiasedRNG[525];
            InitCond[1242] = UnbiasedRNG[526];
            InitCond[1243] = UnbiasedRNG[527];
            InitCond[1244] = UnbiasedRNG[528];
            InitCond[1245] = UnbiasedRNG[529];
            InitCond[1246] = UnbiasedRNG[530];
            InitCond[1247] = UnbiasedRNG[531];
            InitCond[1248] = UnbiasedRNG[532];
            InitCond[1249] = UnbiasedRNG[533];
            InitCond[1250] = UnbiasedRNG[534];
            InitCond[1251] = UnbiasedRNG[535];
            InitCond[1252] = UnbiasedRNG[536];
            InitCond[1253] = UnbiasedRNG[537];
            InitCond[1254] = UnbiasedRNG[538];
            InitCond[1255] = UnbiasedRNG[539];
            InitCond[1256] = UnbiasedRNG[540];
            InitCond[1257] = UnbiasedRNG[541];
            InitCond[1258] = UnbiasedRNG[542];
            InitCond[1259] = UnbiasedRNG[543];
            InitCond[1260] = UnbiasedRNG[544];
            InitCond[1261] = UnbiasedRNG[545];
            InitCond[1262] = UnbiasedRNG[546];
            InitCond[1263] = UnbiasedRNG[547];
            InitCond[1264] = UnbiasedRNG[548];
            InitCond[1265] = UnbiasedRNG[549];
            InitCond[1266] = UnbiasedRNG[550];
            InitCond[1267] = UnbiasedRNG[551];
            InitCond[1268] = UnbiasedRNG[552];
            InitCond[1269] = UnbiasedRNG[553];
            InitCond[1270] = UnbiasedRNG[554];
            InitCond[1271] = UnbiasedRNG[555];
            InitCond[1272] = UnbiasedRNG[556];
            InitCond[1273] = UnbiasedRNG[557];
            InitCond[1274] = UnbiasedRNG[558];
            InitCond[1275] = UnbiasedRNG[559];
            InitCond[1276] = UnbiasedRNG[560];
            InitCond[1277] = UnbiasedRNG[561];
            InitCond[1278] = UnbiasedRNG[562];
            InitCond[1279] = UnbiasedRNG[563];
            InitCond[1280] = UnbiasedRNG[564];
            InitCond[1281] = UnbiasedRNG[565];
            InitCond[1282] = UnbiasedRNG[566];
            InitCond[1283] = UnbiasedRNG[567];
            InitCond[1284] = UnbiasedRNG[568];
            InitCond[1285] = UnbiasedRNG[569];
            InitCond[1286] = UnbiasedRNG[570];
            InitCond[1287] = UnbiasedRNG[571];
            InitCond[1288] = UnbiasedRNG[572];
            InitCond[1289] = UnbiasedRNG[573];
            InitCond[1290] = UnbiasedRNG[574];
            InitCond[1291] = UnbiasedRNG[575];
            InitCond[1292] = UnbiasedRNG[576];
            InitCond[1293] = UnbiasedRNG[577];
            InitCond[1294] = UnbiasedRNG[578];
            InitCond[1295] = UnbiasedRNG[579];
            InitCond[1296] = UnbiasedRNG[580];
            InitCond[1297] = UnbiasedRNG[581];
            InitCond[1298] = UnbiasedRNG[582];
            InitCond[1299] = UnbiasedRNG[583];
            InitCond[1300] = UnbiasedRNG[584];
            InitCond[1301] = UnbiasedRNG[585];
            InitCond[1302] = UnbiasedRNG[586];
            InitCond[1303] = UnbiasedRNG[587];
            InitCond[1304] = UnbiasedRNG[588];
            InitCond[1305] = UnbiasedRNG[589];
            InitCond[1306] = UnbiasedRNG[590];
            InitCond[1307] = UnbiasedRNG[591];
            InitCond[1308] = UnbiasedRNG[592];
            InitCond[1309] = UnbiasedRNG[593];
            InitCond[1310] = UnbiasedRNG[594];
            InitCond[1311] = UnbiasedRNG[595];
            InitCond[1312] = UnbiasedRNG[596];
            InitCond[1313] = UnbiasedRNG[597];
            InitCond[1314] = UnbiasedRNG[598];
            InitCond[1315] = UnbiasedRNG[599];
            InitCond[1316] = UnbiasedRNG[600];
            InitCond[1317] = UnbiasedRNG[601];
            InitCond[1318] = UnbiasedRNG[602];
            InitCond[1319] = UnbiasedRNG[603];
            InitCond[1320] = UnbiasedRNG[604];
            InitCond[1321] = UnbiasedRNG[605];
            InitCond[1322] = UnbiasedRNG[606];
            InitCond[1323] = UnbiasedRNG[607];
            InitCond[1324] = UnbiasedRNG[608];
            InitCond[1325] = UnbiasedRNG[609];
            InitCond[1326] = UnbiasedRNG[610];
            InitCond[1327] = UnbiasedRNG[611];
            InitCond[1328] = UnbiasedRNG[612];
            InitCond[1329] = UnbiasedRNG[613];
            InitCond[1330] = UnbiasedRNG[614];
            InitCond[1331] = UnbiasedRNG[615];
            InitCond[1332] = UnbiasedRNG[616];
            InitCond[1333] = UnbiasedRNG[617];
            InitCond[1334] = UnbiasedRNG[618];
            InitCond[1335] = UnbiasedRNG[619];
            InitCond[1336] = UnbiasedRNG[620];
            InitCond[1337] = UnbiasedRNG[621];
            InitCond[1338] = UnbiasedRNG[622];
            InitCond[1339] = UnbiasedRNG[623];
            InitCond[1340] = UnbiasedRNG[624];
            InitCond[1341] = UnbiasedRNG[625];
            InitCond[1342] = UnbiasedRNG[626];
            InitCond[1343] = UnbiasedRNG[627];
            InitCond[1344] = UnbiasedRNG[628];
            InitCond[1345] = UnbiasedRNG[629];
            InitCond[1346] = UnbiasedRNG[630];
            InitCond[1347] = UnbiasedRNG[631];
            InitCond[1348] = UnbiasedRNG[632];
            InitCond[1349] = UnbiasedRNG[633];
            InitCond[1350] = UnbiasedRNG[634];
            InitCond[1351] = UnbiasedRNG[635];
            InitCond[1352] = UnbiasedRNG[636];
            InitCond[1353] = UnbiasedRNG[637];
            InitCond[1354] = UnbiasedRNG[638];
            InitCond[1355] = UnbiasedRNG[639];
            InitCond[1356] = UnbiasedRNG[640];
            InitCond[1357] = UnbiasedRNG[641];
            InitCond[1358] = UnbiasedRNG[642];
            InitCond[1359] = UnbiasedRNG[643];
            InitCond[1360] = UnbiasedRNG[644];
            InitCond[1361] = UnbiasedRNG[645];
            InitCond[1362] = UnbiasedRNG[646];
            InitCond[1363] = UnbiasedRNG[647];
            InitCond[1364] = UnbiasedRNG[648];
            InitCond[1365] = UnbiasedRNG[649];
            InitCond[1366] = UnbiasedRNG[650];
            InitCond[1367] = UnbiasedRNG[651];
            InitCond[1368] = UnbiasedRNG[652];
            InitCond[1369] = UnbiasedRNG[653];
            InitCond[1370] = UnbiasedRNG[654];
            InitCond[1371] = UnbiasedRNG[655];
            InitCond[1372] = UnbiasedRNG[656];
            InitCond[1373] = UnbiasedRNG[657];
            InitCond[1374] = UnbiasedRNG[658];
            InitCond[1375] = UnbiasedRNG[659];
            InitCond[1376] = UnbiasedRNG[660];
            InitCond[1377] = UnbiasedRNG[661];
            InitCond[1378] = UnbiasedRNG[662];
            InitCond[1379] = UnbiasedRNG[663];
            InitCond[1380] = UnbiasedRNG[664];
            InitCond[1381] = UnbiasedRNG[665];
            InitCond[1382] = UnbiasedRNG[666];
            InitCond[1383] = UnbiasedRNG[667];
            InitCond[1384] = UnbiasedRNG[668];
            InitCond[1385] = UnbiasedRNG[669];
            InitCond[1386] = UnbiasedRNG[670];
            InitCond[1387] = UnbiasedRNG[671];
            InitCond[1388] = UnbiasedRNG[672];
            InitCond[1389] = UnbiasedRNG[673];
            InitCond[1390] = UnbiasedRNG[674];
            InitCond[1391] = UnbiasedRNG[675];
            InitCond[1392] = UnbiasedRNG[676];
            InitCond[1393] = UnbiasedRNG[677];
            InitCond[1394] = UnbiasedRNG[678];
            InitCond[1395] = UnbiasedRNG[679];
            InitCond[1396] = UnbiasedRNG[680];
            InitCond[1397] = UnbiasedRNG[681];
            InitCond[1398] = UnbiasedRNG[682];
            InitCond[1399] = UnbiasedRNG[683];
            InitCond[1400] = UnbiasedRNG[684];
            InitCond[1401] = UnbiasedRNG[685];
            InitCond[1402] = UnbiasedRNG[686];
            InitCond[1403] = UnbiasedRNG[687];
            InitCond[1404] = UnbiasedRNG[688];
            InitCond[1405] = UnbiasedRNG[689];
            InitCond[1406] = UnbiasedRNG[690];
            InitCond[1407] = UnbiasedRNG[691];
            InitCond[1408] = UnbiasedRNG[692];
            InitCond[1409] = UnbiasedRNG[693];
            InitCond[1410] = UnbiasedRNG[694];
            InitCond[1411] = UnbiasedRNG[695];
            InitCond[1412] = UnbiasedRNG[696];
            InitCond[1413] = UnbiasedRNG[697];
            InitCond[1414] = UnbiasedRNG[698];
            InitCond[1415] = UnbiasedRNG[699];
            InitCond[1416] = UnbiasedRNG[700];
            InitCond[1417] = UnbiasedRNG[701];
            InitCond[1418] = UnbiasedRNG[702];
            InitCond[1419] = UnbiasedRNG[703];
            InitCond[1420] = UnbiasedRNG[704];
            InitCond[1421] = UnbiasedRNG[705];
            InitCond[1422] = UnbiasedRNG[706];
            InitCond[1423] = UnbiasedRNG[707];
            InitCond[1424] = UnbiasedRNG[708];
            InitCond[1425] = UnbiasedRNG[709];
            InitCond[1426] = UnbiasedRNG[710];
            InitCond[1427] = UnbiasedRNG[711];
            InitCond[1428] = UnbiasedRNG[712];
            InitCond[1429] = UnbiasedRNG[713];
            InitCond[1430] = UnbiasedRNG[714];
            InitCond[1431] = UnbiasedRNG[715];
        end
        else if (counter == 3) begin
            InitCond[1432] = UnbiasedRNG[0];
            InitCond[1433] = UnbiasedRNG[1];
            InitCond[1434] = UnbiasedRNG[2];
            InitCond[1435] = UnbiasedRNG[3];
            InitCond[1436] = UnbiasedRNG[4];
            InitCond[1437] = UnbiasedRNG[5];
            InitCond[1438] = UnbiasedRNG[6];
            InitCond[1439] = UnbiasedRNG[7];
            InitCond[1440] = UnbiasedRNG[8];
            InitCond[1441] = UnbiasedRNG[9];
            InitCond[1442] = UnbiasedRNG[10];
            InitCond[1443] = UnbiasedRNG[11];
            InitCond[1444] = UnbiasedRNG[12];
            InitCond[1445] = UnbiasedRNG[13];
            InitCond[1446] = UnbiasedRNG[14];
            InitCond[1447] = UnbiasedRNG[15];
            InitCond[1448] = UnbiasedRNG[16];
            InitCond[1449] = UnbiasedRNG[17];
            InitCond[1450] = UnbiasedRNG[18];
            InitCond[1451] = UnbiasedRNG[19];
            InitCond[1452] = UnbiasedRNG[20];
            InitCond[1453] = UnbiasedRNG[21];
            InitCond[1454] = UnbiasedRNG[22];
            InitCond[1455] = UnbiasedRNG[23];
            InitCond[1456] = UnbiasedRNG[24];
            InitCond[1457] = UnbiasedRNG[25];
            InitCond[1458] = UnbiasedRNG[26];
            InitCond[1459] = UnbiasedRNG[27];
            InitCond[1460] = UnbiasedRNG[28];
            InitCond[1461] = UnbiasedRNG[29];
            InitCond[1462] = UnbiasedRNG[30];
            InitCond[1463] = UnbiasedRNG[31];
            InitCond[1464] = UnbiasedRNG[32];
            InitCond[1465] = UnbiasedRNG[33];
            InitCond[1466] = UnbiasedRNG[34];
            InitCond[1467] = UnbiasedRNG[35];
            InitCond[1468] = UnbiasedRNG[36];
            InitCond[1469] = UnbiasedRNG[37];
            InitCond[1470] = UnbiasedRNG[38];
            InitCond[1471] = UnbiasedRNG[39];
            InitCond[1472] = UnbiasedRNG[40];
            InitCond[1473] = UnbiasedRNG[41];
            InitCond[1474] = UnbiasedRNG[42];
            InitCond[1475] = UnbiasedRNG[43];
            InitCond[1476] = UnbiasedRNG[44];
            InitCond[1477] = UnbiasedRNG[45];
            InitCond[1478] = UnbiasedRNG[46];
            InitCond[1479] = UnbiasedRNG[47];
            InitCond[1480] = UnbiasedRNG[48];
            InitCond[1481] = UnbiasedRNG[49];
            InitCond[1482] = UnbiasedRNG[50];
            InitCond[1483] = UnbiasedRNG[51];
            InitCond[1484] = UnbiasedRNG[52];
            InitCond[1485] = UnbiasedRNG[53];
            InitCond[1486] = UnbiasedRNG[54];
            InitCond[1487] = UnbiasedRNG[55];
            InitCond[1488] = UnbiasedRNG[56];
            InitCond[1489] = UnbiasedRNG[57];
            InitCond[1490] = UnbiasedRNG[58];
            InitCond[1491] = UnbiasedRNG[59];
            InitCond[1492] = UnbiasedRNG[60];
            InitCond[1493] = UnbiasedRNG[61];
            InitCond[1494] = UnbiasedRNG[62];
            InitCond[1495] = UnbiasedRNG[63];
            InitCond[1496] = UnbiasedRNG[64];
            InitCond[1497] = UnbiasedRNG[65];
            InitCond[1498] = UnbiasedRNG[66];
            InitCond[1499] = UnbiasedRNG[67];
            InitCond[1500] = UnbiasedRNG[68];
            InitCond[1501] = UnbiasedRNG[69];
            InitCond[1502] = UnbiasedRNG[70];
            InitCond[1503] = UnbiasedRNG[71];
            InitCond[1504] = UnbiasedRNG[72];
            InitCond[1505] = UnbiasedRNG[73];
            InitCond[1506] = UnbiasedRNG[74];
            InitCond[1507] = UnbiasedRNG[75];
            InitCond[1508] = UnbiasedRNG[76];
            InitCond[1509] = UnbiasedRNG[77];
            InitCond[1510] = UnbiasedRNG[78];
            InitCond[1511] = UnbiasedRNG[79];
            InitCond[1512] = UnbiasedRNG[80];
            InitCond[1513] = UnbiasedRNG[81];
            InitCond[1514] = UnbiasedRNG[82];
            InitCond[1515] = UnbiasedRNG[83];
            InitCond[1516] = UnbiasedRNG[84];
            InitCond[1517] = UnbiasedRNG[85];
            InitCond[1518] = UnbiasedRNG[86];
            InitCond[1519] = UnbiasedRNG[87];
            InitCond[1520] = UnbiasedRNG[88];
            InitCond[1521] = UnbiasedRNG[89];
            InitCond[1522] = UnbiasedRNG[90];
            InitCond[1523] = UnbiasedRNG[91];
            InitCond[1524] = UnbiasedRNG[92];
            InitCond[1525] = UnbiasedRNG[93];
            InitCond[1526] = UnbiasedRNG[94];
            InitCond[1527] = UnbiasedRNG[95];
            InitCond[1528] = UnbiasedRNG[96];
            InitCond[1529] = UnbiasedRNG[97];
            InitCond[1530] = UnbiasedRNG[98];
            InitCond[1531] = UnbiasedRNG[99];
            InitCond[1532] = UnbiasedRNG[100];
            InitCond[1533] = UnbiasedRNG[101];
            InitCond[1534] = UnbiasedRNG[102];
            InitCond[1535] = UnbiasedRNG[103];
            InitCond[1536] = UnbiasedRNG[104];
            InitCond[1537] = UnbiasedRNG[105];
            InitCond[1538] = UnbiasedRNG[106];
            InitCond[1539] = UnbiasedRNG[107];
            InitCond[1540] = UnbiasedRNG[108];
            InitCond[1541] = UnbiasedRNG[109];
            InitCond[1542] = UnbiasedRNG[110];
            InitCond[1543] = UnbiasedRNG[111];
            InitCond[1544] = UnbiasedRNG[112];
            InitCond[1545] = UnbiasedRNG[113];
            InitCond[1546] = UnbiasedRNG[114];
            InitCond[1547] = UnbiasedRNG[115];
            InitCond[1548] = UnbiasedRNG[116];
            InitCond[1549] = UnbiasedRNG[117];
            InitCond[1550] = UnbiasedRNG[118];
            InitCond[1551] = UnbiasedRNG[119];
            InitCond[1552] = UnbiasedRNG[120];
            InitCond[1553] = UnbiasedRNG[121];
            InitCond[1554] = UnbiasedRNG[122];
            InitCond[1555] = UnbiasedRNG[123];
            InitCond[1556] = UnbiasedRNG[124];
            InitCond[1557] = UnbiasedRNG[125];
            InitCond[1558] = UnbiasedRNG[126];
            InitCond[1559] = UnbiasedRNG[127];
            InitCond[1560] = UnbiasedRNG[128];
            InitCond[1561] = UnbiasedRNG[129];
            InitCond[1562] = UnbiasedRNG[130];
            InitCond[1563] = UnbiasedRNG[131];
            InitCond[1564] = UnbiasedRNG[132];
            InitCond[1565] = UnbiasedRNG[133];
            InitCond[1566] = UnbiasedRNG[134];
            InitCond[1567] = UnbiasedRNG[135];
            InitCond[1568] = UnbiasedRNG[136];
            InitCond[1569] = UnbiasedRNG[137];
            InitCond[1570] = UnbiasedRNG[138];
            InitCond[1571] = UnbiasedRNG[139];
            InitCond[1572] = UnbiasedRNG[140];
            InitCond[1573] = UnbiasedRNG[141];
            InitCond[1574] = UnbiasedRNG[142];
            InitCond[1575] = UnbiasedRNG[143];
            InitCond[1576] = UnbiasedRNG[144];
            InitCond[1577] = UnbiasedRNG[145];
            InitCond[1578] = UnbiasedRNG[146];
            InitCond[1579] = UnbiasedRNG[147];
            InitCond[1580] = UnbiasedRNG[148];
            InitCond[1581] = UnbiasedRNG[149];
            InitCond[1582] = UnbiasedRNG[150];
            InitCond[1583] = UnbiasedRNG[151];
            InitCond[1584] = UnbiasedRNG[152];
            InitCond[1585] = UnbiasedRNG[153];
            InitCond[1586] = UnbiasedRNG[154];
            InitCond[1587] = UnbiasedRNG[155];
            InitCond[1588] = UnbiasedRNG[156];
            InitCond[1589] = UnbiasedRNG[157];
            InitCond[1590] = UnbiasedRNG[158];
            InitCond[1591] = UnbiasedRNG[159];
            InitCond[1592] = UnbiasedRNG[160];
            InitCond[1593] = UnbiasedRNG[161];
            InitCond[1594] = UnbiasedRNG[162];
            InitCond[1595] = UnbiasedRNG[163];
        end
        else if (counter==5)
            run = 1'b1;
        counter = counter+38'b1;
        solution = {m[13],m[12],m[11],m[10],m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[27],m[26],m[25],m[24],m[23],m[22],m[21],m[20],m[19],m[18],m[17],m[16],m[15],m[14]};
    end else begin 
        counter = 38'b0;
        failure = 1'b1;
        run = 1'b0;
    end
end

//To measure on only the last step using ILA:
always @(negedge sample_clk) begin
    if (solution_flag)
        solution_flag = 1'b0;
    else if ((run & (solution == solution_check)) | failure)
        solution_flag = 1'b1;
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = run?((((m[28]&~m[56])|(~m[28]&m[56]))&UnbiasedRNG[0])|((m[28]&m[56]))):InitCond[0];
    m[1] = run?((((m[29]&~m[59])|(~m[29]&m[59]))&UnbiasedRNG[1])|((m[29]&m[59]))):InitCond[1];
    m[2] = run?((((m[30]&~m[62])|(~m[30]&m[62]))&UnbiasedRNG[2])|((m[30]&m[62]))):InitCond[2];
    m[3] = run?((((m[31]&~m[65])|(~m[31]&m[65]))&UnbiasedRNG[3])|((m[31]&m[65]))):InitCond[3];
    m[4] = run?((((m[32]&~m[68])|(~m[32]&m[68]))&UnbiasedRNG[4])|((m[32]&m[68]))):InitCond[4];
    m[5] = run?((((m[33]&~m[71])|(~m[33]&m[71]))&UnbiasedRNG[5])|((m[33]&m[71]))):InitCond[5];
    m[6] = run?((((m[34]&~m[74])|(~m[34]&m[74]))&UnbiasedRNG[6])|((m[34]&m[74]))):InitCond[6];
    m[7] = run?((((m[35]&~m[77])|(~m[35]&m[77]))&UnbiasedRNG[7])|((m[35]&m[77]))):InitCond[7];
    m[8] = run?((((m[36]&~m[80])|(~m[36]&m[80]))&UnbiasedRNG[8])|((m[36]&m[80]))):InitCond[8];
    m[9] = run?((((m[37]&~m[83])|(~m[37]&m[83]))&UnbiasedRNG[9])|((m[37]&m[83]))):InitCond[9];
    m[10] = run?((((m[38]&~m[86])|(~m[38]&m[86]))&UnbiasedRNG[10])|((m[38]&m[86]))):InitCond[10];
    m[11] = run?((((m[39]&~m[89])|(~m[39]&m[89]))&UnbiasedRNG[11])|((m[39]&m[89]))):InitCond[11];
    m[12] = run?((((m[40]&~m[92])|(~m[40]&m[92]))&UnbiasedRNG[12])|((m[40]&m[92]))):InitCond[12];
    m[13] = run?((((m[41]&~m[95])|(~m[41]&m[95]))&UnbiasedRNG[13])|((m[41]&m[95]))):InitCond[13];
    m[14] = run?((((m[42]&~m[98])|(~m[42]&m[98]))&UnbiasedRNG[14])|((m[42]&m[98]))):InitCond[14];
    m[15] = run?((((m[43]&~m[101])|(~m[43]&m[101]))&UnbiasedRNG[15])|((m[43]&m[101]))):InitCond[15];
    m[16] = run?((((m[44]&~m[104])|(~m[44]&m[104]))&UnbiasedRNG[16])|((m[44]&m[104]))):InitCond[16];
    m[17] = run?((((m[45]&~m[107])|(~m[45]&m[107]))&UnbiasedRNG[17])|((m[45]&m[107]))):InitCond[17];
    m[18] = run?((((m[46]&~m[110])|(~m[46]&m[110]))&UnbiasedRNG[18])|((m[46]&m[110]))):InitCond[18];
    m[19] = run?((((m[47]&~m[113])|(~m[47]&m[113]))&UnbiasedRNG[19])|((m[47]&m[113]))):InitCond[19];
    m[20] = run?((((m[48]&~m[116])|(~m[48]&m[116]))&UnbiasedRNG[20])|((m[48]&m[116]))):InitCond[20];
    m[21] = run?((((m[49]&~m[119])|(~m[49]&m[119]))&UnbiasedRNG[21])|((m[49]&m[119]))):InitCond[21];
    m[22] = run?((((m[50]&~m[122])|(~m[50]&m[122]))&UnbiasedRNG[22])|((m[50]&m[122]))):InitCond[22];
    m[23] = run?((((m[51]&~m[125])|(~m[51]&m[125]))&UnbiasedRNG[23])|((m[51]&m[125]))):InitCond[23];
    m[24] = run?((((m[52]&~m[128])|(~m[52]&m[128]))&UnbiasedRNG[24])|((m[52]&m[128]))):InitCond[24];
    m[25] = run?((((m[53]&~m[131])|(~m[53]&m[131]))&UnbiasedRNG[25])|((m[53]&m[131]))):InitCond[25];
    m[26] = run?((((m[54]&~m[134])|(~m[54]&m[134]))&UnbiasedRNG[26])|((m[54]&m[134]))):InitCond[26];
    m[27] = run?((((m[55]&~m[137])|(~m[55]&m[137]))&UnbiasedRNG[27])|((m[55]&m[137]))):InitCond[27];
    m[57] = run?((((m[28]&m[146]&~m[147]&~m[148]&~m[149])|(m[28]&~m[146]&m[147]&~m[148]&~m[149])|(~m[28]&m[146]&m[147]&~m[148]&~m[149])|(m[28]&~m[146]&~m[147]&m[148]&~m[149])|(~m[28]&m[146]&~m[147]&m[148]&~m[149])|(~m[28]&~m[146]&m[147]&m[148]&~m[149])|(m[28]&~m[146]&~m[147]&~m[148]&m[149])|(~m[28]&m[146]&~m[147]&~m[148]&m[149])|(~m[28]&~m[146]&m[147]&~m[148]&m[149])|(~m[28]&~m[146]&~m[147]&m[148]&m[149]))&BiasedRNG[0])|(((m[28]&m[146]&m[147]&~m[148]&~m[149])|(m[28]&m[146]&~m[147]&m[148]&~m[149])|(m[28]&~m[146]&m[147]&m[148]&~m[149])|(~m[28]&m[146]&m[147]&m[148]&~m[149])|(m[28]&m[146]&~m[147]&~m[148]&m[149])|(m[28]&~m[146]&m[147]&~m[148]&m[149])|(~m[28]&m[146]&m[147]&~m[148]&m[149])|(m[28]&~m[146]&~m[147]&m[148]&m[149])|(~m[28]&m[146]&~m[147]&m[148]&m[149])|(~m[28]&~m[146]&m[147]&m[148]&m[149]))&~BiasedRNG[0])|((m[28]&m[146]&m[147]&m[148]&~m[149])|(m[28]&m[146]&m[147]&~m[148]&m[149])|(m[28]&m[146]&~m[147]&m[148]&m[149])|(m[28]&~m[146]&m[147]&m[148]&m[149])|(~m[28]&m[146]&m[147]&m[148]&m[149])|(m[28]&m[146]&m[147]&m[148]&m[149]))):InitCond[28];
    m[58] = run?((((m[28]&m[150]&~m[151]&~m[152]&~m[153])|(m[28]&~m[150]&m[151]&~m[152]&~m[153])|(~m[28]&m[150]&m[151]&~m[152]&~m[153])|(m[28]&~m[150]&~m[151]&m[152]&~m[153])|(~m[28]&m[150]&~m[151]&m[152]&~m[153])|(~m[28]&~m[150]&m[151]&m[152]&~m[153])|(m[28]&~m[150]&~m[151]&~m[152]&m[153])|(~m[28]&m[150]&~m[151]&~m[152]&m[153])|(~m[28]&~m[150]&m[151]&~m[152]&m[153])|(~m[28]&~m[150]&~m[151]&m[152]&m[153]))&BiasedRNG[1])|(((m[28]&m[150]&m[151]&~m[152]&~m[153])|(m[28]&m[150]&~m[151]&m[152]&~m[153])|(m[28]&~m[150]&m[151]&m[152]&~m[153])|(~m[28]&m[150]&m[151]&m[152]&~m[153])|(m[28]&m[150]&~m[151]&~m[152]&m[153])|(m[28]&~m[150]&m[151]&~m[152]&m[153])|(~m[28]&m[150]&m[151]&~m[152]&m[153])|(m[28]&~m[150]&~m[151]&m[152]&m[153])|(~m[28]&m[150]&~m[151]&m[152]&m[153])|(~m[28]&~m[150]&m[151]&m[152]&m[153]))&~BiasedRNG[1])|((m[28]&m[150]&m[151]&m[152]&~m[153])|(m[28]&m[150]&m[151]&~m[152]&m[153])|(m[28]&m[150]&~m[151]&m[152]&m[153])|(m[28]&~m[150]&m[151]&m[152]&m[153])|(~m[28]&m[150]&m[151]&m[152]&m[153])|(m[28]&m[150]&m[151]&m[152]&m[153]))):InitCond[29];
    m[60] = run?((((m[29]&m[160]&~m[161]&~m[162]&~m[163])|(m[29]&~m[160]&m[161]&~m[162]&~m[163])|(~m[29]&m[160]&m[161]&~m[162]&~m[163])|(m[29]&~m[160]&~m[161]&m[162]&~m[163])|(~m[29]&m[160]&~m[161]&m[162]&~m[163])|(~m[29]&~m[160]&m[161]&m[162]&~m[163])|(m[29]&~m[160]&~m[161]&~m[162]&m[163])|(~m[29]&m[160]&~m[161]&~m[162]&m[163])|(~m[29]&~m[160]&m[161]&~m[162]&m[163])|(~m[29]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[2])|(((m[29]&m[160]&m[161]&~m[162]&~m[163])|(m[29]&m[160]&~m[161]&m[162]&~m[163])|(m[29]&~m[160]&m[161]&m[162]&~m[163])|(~m[29]&m[160]&m[161]&m[162]&~m[163])|(m[29]&m[160]&~m[161]&~m[162]&m[163])|(m[29]&~m[160]&m[161]&~m[162]&m[163])|(~m[29]&m[160]&m[161]&~m[162]&m[163])|(m[29]&~m[160]&~m[161]&m[162]&m[163])|(~m[29]&m[160]&~m[161]&m[162]&m[163])|(~m[29]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[2])|((m[29]&m[160]&m[161]&m[162]&~m[163])|(m[29]&m[160]&m[161]&~m[162]&m[163])|(m[29]&m[160]&~m[161]&m[162]&m[163])|(m[29]&~m[160]&m[161]&m[162]&m[163])|(~m[29]&m[160]&m[161]&m[162]&m[163])|(m[29]&m[160]&m[161]&m[162]&m[163]))):InitCond[30];
    m[61] = run?((((m[29]&m[164]&~m[165]&~m[166]&~m[167])|(m[29]&~m[164]&m[165]&~m[166]&~m[167])|(~m[29]&m[164]&m[165]&~m[166]&~m[167])|(m[29]&~m[164]&~m[165]&m[166]&~m[167])|(~m[29]&m[164]&~m[165]&m[166]&~m[167])|(~m[29]&~m[164]&m[165]&m[166]&~m[167])|(m[29]&~m[164]&~m[165]&~m[166]&m[167])|(~m[29]&m[164]&~m[165]&~m[166]&m[167])|(~m[29]&~m[164]&m[165]&~m[166]&m[167])|(~m[29]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[3])|(((m[29]&m[164]&m[165]&~m[166]&~m[167])|(m[29]&m[164]&~m[165]&m[166]&~m[167])|(m[29]&~m[164]&m[165]&m[166]&~m[167])|(~m[29]&m[164]&m[165]&m[166]&~m[167])|(m[29]&m[164]&~m[165]&~m[166]&m[167])|(m[29]&~m[164]&m[165]&~m[166]&m[167])|(~m[29]&m[164]&m[165]&~m[166]&m[167])|(m[29]&~m[164]&~m[165]&m[166]&m[167])|(~m[29]&m[164]&~m[165]&m[166]&m[167])|(~m[29]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[3])|((m[29]&m[164]&m[165]&m[166]&~m[167])|(m[29]&m[164]&m[165]&~m[166]&m[167])|(m[29]&m[164]&~m[165]&m[166]&m[167])|(m[29]&~m[164]&m[165]&m[166]&m[167])|(~m[29]&m[164]&m[165]&m[166]&m[167])|(m[29]&m[164]&m[165]&m[166]&m[167]))):InitCond[31];
    m[63] = run?((((m[30]&m[174]&~m[175]&~m[176]&~m[177])|(m[30]&~m[174]&m[175]&~m[176]&~m[177])|(~m[30]&m[174]&m[175]&~m[176]&~m[177])|(m[30]&~m[174]&~m[175]&m[176]&~m[177])|(~m[30]&m[174]&~m[175]&m[176]&~m[177])|(~m[30]&~m[174]&m[175]&m[176]&~m[177])|(m[30]&~m[174]&~m[175]&~m[176]&m[177])|(~m[30]&m[174]&~m[175]&~m[176]&m[177])|(~m[30]&~m[174]&m[175]&~m[176]&m[177])|(~m[30]&~m[174]&~m[175]&m[176]&m[177]))&BiasedRNG[4])|(((m[30]&m[174]&m[175]&~m[176]&~m[177])|(m[30]&m[174]&~m[175]&m[176]&~m[177])|(m[30]&~m[174]&m[175]&m[176]&~m[177])|(~m[30]&m[174]&m[175]&m[176]&~m[177])|(m[30]&m[174]&~m[175]&~m[176]&m[177])|(m[30]&~m[174]&m[175]&~m[176]&m[177])|(~m[30]&m[174]&m[175]&~m[176]&m[177])|(m[30]&~m[174]&~m[175]&m[176]&m[177])|(~m[30]&m[174]&~m[175]&m[176]&m[177])|(~m[30]&~m[174]&m[175]&m[176]&m[177]))&~BiasedRNG[4])|((m[30]&m[174]&m[175]&m[176]&~m[177])|(m[30]&m[174]&m[175]&~m[176]&m[177])|(m[30]&m[174]&~m[175]&m[176]&m[177])|(m[30]&~m[174]&m[175]&m[176]&m[177])|(~m[30]&m[174]&m[175]&m[176]&m[177])|(m[30]&m[174]&m[175]&m[176]&m[177]))):InitCond[32];
    m[64] = run?((((m[30]&m[178]&~m[179]&~m[180]&~m[181])|(m[30]&~m[178]&m[179]&~m[180]&~m[181])|(~m[30]&m[178]&m[179]&~m[180]&~m[181])|(m[30]&~m[178]&~m[179]&m[180]&~m[181])|(~m[30]&m[178]&~m[179]&m[180]&~m[181])|(~m[30]&~m[178]&m[179]&m[180]&~m[181])|(m[30]&~m[178]&~m[179]&~m[180]&m[181])|(~m[30]&m[178]&~m[179]&~m[180]&m[181])|(~m[30]&~m[178]&m[179]&~m[180]&m[181])|(~m[30]&~m[178]&~m[179]&m[180]&m[181]))&BiasedRNG[5])|(((m[30]&m[178]&m[179]&~m[180]&~m[181])|(m[30]&m[178]&~m[179]&m[180]&~m[181])|(m[30]&~m[178]&m[179]&m[180]&~m[181])|(~m[30]&m[178]&m[179]&m[180]&~m[181])|(m[30]&m[178]&~m[179]&~m[180]&m[181])|(m[30]&~m[178]&m[179]&~m[180]&m[181])|(~m[30]&m[178]&m[179]&~m[180]&m[181])|(m[30]&~m[178]&~m[179]&m[180]&m[181])|(~m[30]&m[178]&~m[179]&m[180]&m[181])|(~m[30]&~m[178]&m[179]&m[180]&m[181]))&~BiasedRNG[5])|((m[30]&m[178]&m[179]&m[180]&~m[181])|(m[30]&m[178]&m[179]&~m[180]&m[181])|(m[30]&m[178]&~m[179]&m[180]&m[181])|(m[30]&~m[178]&m[179]&m[180]&m[181])|(~m[30]&m[178]&m[179]&m[180]&m[181])|(m[30]&m[178]&m[179]&m[180]&m[181]))):InitCond[33];
    m[66] = run?((((m[31]&m[188]&~m[189]&~m[190]&~m[191])|(m[31]&~m[188]&m[189]&~m[190]&~m[191])|(~m[31]&m[188]&m[189]&~m[190]&~m[191])|(m[31]&~m[188]&~m[189]&m[190]&~m[191])|(~m[31]&m[188]&~m[189]&m[190]&~m[191])|(~m[31]&~m[188]&m[189]&m[190]&~m[191])|(m[31]&~m[188]&~m[189]&~m[190]&m[191])|(~m[31]&m[188]&~m[189]&~m[190]&m[191])|(~m[31]&~m[188]&m[189]&~m[190]&m[191])|(~m[31]&~m[188]&~m[189]&m[190]&m[191]))&BiasedRNG[6])|(((m[31]&m[188]&m[189]&~m[190]&~m[191])|(m[31]&m[188]&~m[189]&m[190]&~m[191])|(m[31]&~m[188]&m[189]&m[190]&~m[191])|(~m[31]&m[188]&m[189]&m[190]&~m[191])|(m[31]&m[188]&~m[189]&~m[190]&m[191])|(m[31]&~m[188]&m[189]&~m[190]&m[191])|(~m[31]&m[188]&m[189]&~m[190]&m[191])|(m[31]&~m[188]&~m[189]&m[190]&m[191])|(~m[31]&m[188]&~m[189]&m[190]&m[191])|(~m[31]&~m[188]&m[189]&m[190]&m[191]))&~BiasedRNG[6])|((m[31]&m[188]&m[189]&m[190]&~m[191])|(m[31]&m[188]&m[189]&~m[190]&m[191])|(m[31]&m[188]&~m[189]&m[190]&m[191])|(m[31]&~m[188]&m[189]&m[190]&m[191])|(~m[31]&m[188]&m[189]&m[190]&m[191])|(m[31]&m[188]&m[189]&m[190]&m[191]))):InitCond[34];
    m[67] = run?((((m[31]&m[192]&~m[193]&~m[194]&~m[195])|(m[31]&~m[192]&m[193]&~m[194]&~m[195])|(~m[31]&m[192]&m[193]&~m[194]&~m[195])|(m[31]&~m[192]&~m[193]&m[194]&~m[195])|(~m[31]&m[192]&~m[193]&m[194]&~m[195])|(~m[31]&~m[192]&m[193]&m[194]&~m[195])|(m[31]&~m[192]&~m[193]&~m[194]&m[195])|(~m[31]&m[192]&~m[193]&~m[194]&m[195])|(~m[31]&~m[192]&m[193]&~m[194]&m[195])|(~m[31]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[7])|(((m[31]&m[192]&m[193]&~m[194]&~m[195])|(m[31]&m[192]&~m[193]&m[194]&~m[195])|(m[31]&~m[192]&m[193]&m[194]&~m[195])|(~m[31]&m[192]&m[193]&m[194]&~m[195])|(m[31]&m[192]&~m[193]&~m[194]&m[195])|(m[31]&~m[192]&m[193]&~m[194]&m[195])|(~m[31]&m[192]&m[193]&~m[194]&m[195])|(m[31]&~m[192]&~m[193]&m[194]&m[195])|(~m[31]&m[192]&~m[193]&m[194]&m[195])|(~m[31]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[7])|((m[31]&m[192]&m[193]&m[194]&~m[195])|(m[31]&m[192]&m[193]&~m[194]&m[195])|(m[31]&m[192]&~m[193]&m[194]&m[195])|(m[31]&~m[192]&m[193]&m[194]&m[195])|(~m[31]&m[192]&m[193]&m[194]&m[195])|(m[31]&m[192]&m[193]&m[194]&m[195]))):InitCond[35];
    m[69] = run?((((m[32]&m[202]&~m[203]&~m[204]&~m[205])|(m[32]&~m[202]&m[203]&~m[204]&~m[205])|(~m[32]&m[202]&m[203]&~m[204]&~m[205])|(m[32]&~m[202]&~m[203]&m[204]&~m[205])|(~m[32]&m[202]&~m[203]&m[204]&~m[205])|(~m[32]&~m[202]&m[203]&m[204]&~m[205])|(m[32]&~m[202]&~m[203]&~m[204]&m[205])|(~m[32]&m[202]&~m[203]&~m[204]&m[205])|(~m[32]&~m[202]&m[203]&~m[204]&m[205])|(~m[32]&~m[202]&~m[203]&m[204]&m[205]))&BiasedRNG[8])|(((m[32]&m[202]&m[203]&~m[204]&~m[205])|(m[32]&m[202]&~m[203]&m[204]&~m[205])|(m[32]&~m[202]&m[203]&m[204]&~m[205])|(~m[32]&m[202]&m[203]&m[204]&~m[205])|(m[32]&m[202]&~m[203]&~m[204]&m[205])|(m[32]&~m[202]&m[203]&~m[204]&m[205])|(~m[32]&m[202]&m[203]&~m[204]&m[205])|(m[32]&~m[202]&~m[203]&m[204]&m[205])|(~m[32]&m[202]&~m[203]&m[204]&m[205])|(~m[32]&~m[202]&m[203]&m[204]&m[205]))&~BiasedRNG[8])|((m[32]&m[202]&m[203]&m[204]&~m[205])|(m[32]&m[202]&m[203]&~m[204]&m[205])|(m[32]&m[202]&~m[203]&m[204]&m[205])|(m[32]&~m[202]&m[203]&m[204]&m[205])|(~m[32]&m[202]&m[203]&m[204]&m[205])|(m[32]&m[202]&m[203]&m[204]&m[205]))):InitCond[36];
    m[70] = run?((((m[32]&m[206]&~m[207]&~m[208]&~m[209])|(m[32]&~m[206]&m[207]&~m[208]&~m[209])|(~m[32]&m[206]&m[207]&~m[208]&~m[209])|(m[32]&~m[206]&~m[207]&m[208]&~m[209])|(~m[32]&m[206]&~m[207]&m[208]&~m[209])|(~m[32]&~m[206]&m[207]&m[208]&~m[209])|(m[32]&~m[206]&~m[207]&~m[208]&m[209])|(~m[32]&m[206]&~m[207]&~m[208]&m[209])|(~m[32]&~m[206]&m[207]&~m[208]&m[209])|(~m[32]&~m[206]&~m[207]&m[208]&m[209]))&BiasedRNG[9])|(((m[32]&m[206]&m[207]&~m[208]&~m[209])|(m[32]&m[206]&~m[207]&m[208]&~m[209])|(m[32]&~m[206]&m[207]&m[208]&~m[209])|(~m[32]&m[206]&m[207]&m[208]&~m[209])|(m[32]&m[206]&~m[207]&~m[208]&m[209])|(m[32]&~m[206]&m[207]&~m[208]&m[209])|(~m[32]&m[206]&m[207]&~m[208]&m[209])|(m[32]&~m[206]&~m[207]&m[208]&m[209])|(~m[32]&m[206]&~m[207]&m[208]&m[209])|(~m[32]&~m[206]&m[207]&m[208]&m[209]))&~BiasedRNG[9])|((m[32]&m[206]&m[207]&m[208]&~m[209])|(m[32]&m[206]&m[207]&~m[208]&m[209])|(m[32]&m[206]&~m[207]&m[208]&m[209])|(m[32]&~m[206]&m[207]&m[208]&m[209])|(~m[32]&m[206]&m[207]&m[208]&m[209])|(m[32]&m[206]&m[207]&m[208]&m[209]))):InitCond[37];
    m[72] = run?((((m[33]&m[216]&~m[217]&~m[218]&~m[219])|(m[33]&~m[216]&m[217]&~m[218]&~m[219])|(~m[33]&m[216]&m[217]&~m[218]&~m[219])|(m[33]&~m[216]&~m[217]&m[218]&~m[219])|(~m[33]&m[216]&~m[217]&m[218]&~m[219])|(~m[33]&~m[216]&m[217]&m[218]&~m[219])|(m[33]&~m[216]&~m[217]&~m[218]&m[219])|(~m[33]&m[216]&~m[217]&~m[218]&m[219])|(~m[33]&~m[216]&m[217]&~m[218]&m[219])|(~m[33]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[10])|(((m[33]&m[216]&m[217]&~m[218]&~m[219])|(m[33]&m[216]&~m[217]&m[218]&~m[219])|(m[33]&~m[216]&m[217]&m[218]&~m[219])|(~m[33]&m[216]&m[217]&m[218]&~m[219])|(m[33]&m[216]&~m[217]&~m[218]&m[219])|(m[33]&~m[216]&m[217]&~m[218]&m[219])|(~m[33]&m[216]&m[217]&~m[218]&m[219])|(m[33]&~m[216]&~m[217]&m[218]&m[219])|(~m[33]&m[216]&~m[217]&m[218]&m[219])|(~m[33]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[10])|((m[33]&m[216]&m[217]&m[218]&~m[219])|(m[33]&m[216]&m[217]&~m[218]&m[219])|(m[33]&m[216]&~m[217]&m[218]&m[219])|(m[33]&~m[216]&m[217]&m[218]&m[219])|(~m[33]&m[216]&m[217]&m[218]&m[219])|(m[33]&m[216]&m[217]&m[218]&m[219]))):InitCond[38];
    m[73] = run?((((m[33]&m[220]&~m[221]&~m[222]&~m[223])|(m[33]&~m[220]&m[221]&~m[222]&~m[223])|(~m[33]&m[220]&m[221]&~m[222]&~m[223])|(m[33]&~m[220]&~m[221]&m[222]&~m[223])|(~m[33]&m[220]&~m[221]&m[222]&~m[223])|(~m[33]&~m[220]&m[221]&m[222]&~m[223])|(m[33]&~m[220]&~m[221]&~m[222]&m[223])|(~m[33]&m[220]&~m[221]&~m[222]&m[223])|(~m[33]&~m[220]&m[221]&~m[222]&m[223])|(~m[33]&~m[220]&~m[221]&m[222]&m[223]))&BiasedRNG[11])|(((m[33]&m[220]&m[221]&~m[222]&~m[223])|(m[33]&m[220]&~m[221]&m[222]&~m[223])|(m[33]&~m[220]&m[221]&m[222]&~m[223])|(~m[33]&m[220]&m[221]&m[222]&~m[223])|(m[33]&m[220]&~m[221]&~m[222]&m[223])|(m[33]&~m[220]&m[221]&~m[222]&m[223])|(~m[33]&m[220]&m[221]&~m[222]&m[223])|(m[33]&~m[220]&~m[221]&m[222]&m[223])|(~m[33]&m[220]&~m[221]&m[222]&m[223])|(~m[33]&~m[220]&m[221]&m[222]&m[223]))&~BiasedRNG[11])|((m[33]&m[220]&m[221]&m[222]&~m[223])|(m[33]&m[220]&m[221]&~m[222]&m[223])|(m[33]&m[220]&~m[221]&m[222]&m[223])|(m[33]&~m[220]&m[221]&m[222]&m[223])|(~m[33]&m[220]&m[221]&m[222]&m[223])|(m[33]&m[220]&m[221]&m[222]&m[223]))):InitCond[39];
    m[75] = run?((((m[34]&m[230]&~m[231]&~m[232]&~m[233])|(m[34]&~m[230]&m[231]&~m[232]&~m[233])|(~m[34]&m[230]&m[231]&~m[232]&~m[233])|(m[34]&~m[230]&~m[231]&m[232]&~m[233])|(~m[34]&m[230]&~m[231]&m[232]&~m[233])|(~m[34]&~m[230]&m[231]&m[232]&~m[233])|(m[34]&~m[230]&~m[231]&~m[232]&m[233])|(~m[34]&m[230]&~m[231]&~m[232]&m[233])|(~m[34]&~m[230]&m[231]&~m[232]&m[233])|(~m[34]&~m[230]&~m[231]&m[232]&m[233]))&BiasedRNG[12])|(((m[34]&m[230]&m[231]&~m[232]&~m[233])|(m[34]&m[230]&~m[231]&m[232]&~m[233])|(m[34]&~m[230]&m[231]&m[232]&~m[233])|(~m[34]&m[230]&m[231]&m[232]&~m[233])|(m[34]&m[230]&~m[231]&~m[232]&m[233])|(m[34]&~m[230]&m[231]&~m[232]&m[233])|(~m[34]&m[230]&m[231]&~m[232]&m[233])|(m[34]&~m[230]&~m[231]&m[232]&m[233])|(~m[34]&m[230]&~m[231]&m[232]&m[233])|(~m[34]&~m[230]&m[231]&m[232]&m[233]))&~BiasedRNG[12])|((m[34]&m[230]&m[231]&m[232]&~m[233])|(m[34]&m[230]&m[231]&~m[232]&m[233])|(m[34]&m[230]&~m[231]&m[232]&m[233])|(m[34]&~m[230]&m[231]&m[232]&m[233])|(~m[34]&m[230]&m[231]&m[232]&m[233])|(m[34]&m[230]&m[231]&m[232]&m[233]))):InitCond[40];
    m[76] = run?((((m[34]&m[234]&~m[235]&~m[236]&~m[237])|(m[34]&~m[234]&m[235]&~m[236]&~m[237])|(~m[34]&m[234]&m[235]&~m[236]&~m[237])|(m[34]&~m[234]&~m[235]&m[236]&~m[237])|(~m[34]&m[234]&~m[235]&m[236]&~m[237])|(~m[34]&~m[234]&m[235]&m[236]&~m[237])|(m[34]&~m[234]&~m[235]&~m[236]&m[237])|(~m[34]&m[234]&~m[235]&~m[236]&m[237])|(~m[34]&~m[234]&m[235]&~m[236]&m[237])|(~m[34]&~m[234]&~m[235]&m[236]&m[237]))&BiasedRNG[13])|(((m[34]&m[234]&m[235]&~m[236]&~m[237])|(m[34]&m[234]&~m[235]&m[236]&~m[237])|(m[34]&~m[234]&m[235]&m[236]&~m[237])|(~m[34]&m[234]&m[235]&m[236]&~m[237])|(m[34]&m[234]&~m[235]&~m[236]&m[237])|(m[34]&~m[234]&m[235]&~m[236]&m[237])|(~m[34]&m[234]&m[235]&~m[236]&m[237])|(m[34]&~m[234]&~m[235]&m[236]&m[237])|(~m[34]&m[234]&~m[235]&m[236]&m[237])|(~m[34]&~m[234]&m[235]&m[236]&m[237]))&~BiasedRNG[13])|((m[34]&m[234]&m[235]&m[236]&~m[237])|(m[34]&m[234]&m[235]&~m[236]&m[237])|(m[34]&m[234]&~m[235]&m[236]&m[237])|(m[34]&~m[234]&m[235]&m[236]&m[237])|(~m[34]&m[234]&m[235]&m[236]&m[237])|(m[34]&m[234]&m[235]&m[236]&m[237]))):InitCond[41];
    m[78] = run?((((m[35]&m[244]&~m[245]&~m[246]&~m[247])|(m[35]&~m[244]&m[245]&~m[246]&~m[247])|(~m[35]&m[244]&m[245]&~m[246]&~m[247])|(m[35]&~m[244]&~m[245]&m[246]&~m[247])|(~m[35]&m[244]&~m[245]&m[246]&~m[247])|(~m[35]&~m[244]&m[245]&m[246]&~m[247])|(m[35]&~m[244]&~m[245]&~m[246]&m[247])|(~m[35]&m[244]&~m[245]&~m[246]&m[247])|(~m[35]&~m[244]&m[245]&~m[246]&m[247])|(~m[35]&~m[244]&~m[245]&m[246]&m[247]))&BiasedRNG[14])|(((m[35]&m[244]&m[245]&~m[246]&~m[247])|(m[35]&m[244]&~m[245]&m[246]&~m[247])|(m[35]&~m[244]&m[245]&m[246]&~m[247])|(~m[35]&m[244]&m[245]&m[246]&~m[247])|(m[35]&m[244]&~m[245]&~m[246]&m[247])|(m[35]&~m[244]&m[245]&~m[246]&m[247])|(~m[35]&m[244]&m[245]&~m[246]&m[247])|(m[35]&~m[244]&~m[245]&m[246]&m[247])|(~m[35]&m[244]&~m[245]&m[246]&m[247])|(~m[35]&~m[244]&m[245]&m[246]&m[247]))&~BiasedRNG[14])|((m[35]&m[244]&m[245]&m[246]&~m[247])|(m[35]&m[244]&m[245]&~m[246]&m[247])|(m[35]&m[244]&~m[245]&m[246]&m[247])|(m[35]&~m[244]&m[245]&m[246]&m[247])|(~m[35]&m[244]&m[245]&m[246]&m[247])|(m[35]&m[244]&m[245]&m[246]&m[247]))):InitCond[42];
    m[79] = run?((((m[35]&m[248]&~m[249]&~m[250]&~m[251])|(m[35]&~m[248]&m[249]&~m[250]&~m[251])|(~m[35]&m[248]&m[249]&~m[250]&~m[251])|(m[35]&~m[248]&~m[249]&m[250]&~m[251])|(~m[35]&m[248]&~m[249]&m[250]&~m[251])|(~m[35]&~m[248]&m[249]&m[250]&~m[251])|(m[35]&~m[248]&~m[249]&~m[250]&m[251])|(~m[35]&m[248]&~m[249]&~m[250]&m[251])|(~m[35]&~m[248]&m[249]&~m[250]&m[251])|(~m[35]&~m[248]&~m[249]&m[250]&m[251]))&BiasedRNG[15])|(((m[35]&m[248]&m[249]&~m[250]&~m[251])|(m[35]&m[248]&~m[249]&m[250]&~m[251])|(m[35]&~m[248]&m[249]&m[250]&~m[251])|(~m[35]&m[248]&m[249]&m[250]&~m[251])|(m[35]&m[248]&~m[249]&~m[250]&m[251])|(m[35]&~m[248]&m[249]&~m[250]&m[251])|(~m[35]&m[248]&m[249]&~m[250]&m[251])|(m[35]&~m[248]&~m[249]&m[250]&m[251])|(~m[35]&m[248]&~m[249]&m[250]&m[251])|(~m[35]&~m[248]&m[249]&m[250]&m[251]))&~BiasedRNG[15])|((m[35]&m[248]&m[249]&m[250]&~m[251])|(m[35]&m[248]&m[249]&~m[250]&m[251])|(m[35]&m[248]&~m[249]&m[250]&m[251])|(m[35]&~m[248]&m[249]&m[250]&m[251])|(~m[35]&m[248]&m[249]&m[250]&m[251])|(m[35]&m[248]&m[249]&m[250]&m[251]))):InitCond[43];
    m[81] = run?((((m[36]&m[258]&~m[259]&~m[260]&~m[261])|(m[36]&~m[258]&m[259]&~m[260]&~m[261])|(~m[36]&m[258]&m[259]&~m[260]&~m[261])|(m[36]&~m[258]&~m[259]&m[260]&~m[261])|(~m[36]&m[258]&~m[259]&m[260]&~m[261])|(~m[36]&~m[258]&m[259]&m[260]&~m[261])|(m[36]&~m[258]&~m[259]&~m[260]&m[261])|(~m[36]&m[258]&~m[259]&~m[260]&m[261])|(~m[36]&~m[258]&m[259]&~m[260]&m[261])|(~m[36]&~m[258]&~m[259]&m[260]&m[261]))&BiasedRNG[16])|(((m[36]&m[258]&m[259]&~m[260]&~m[261])|(m[36]&m[258]&~m[259]&m[260]&~m[261])|(m[36]&~m[258]&m[259]&m[260]&~m[261])|(~m[36]&m[258]&m[259]&m[260]&~m[261])|(m[36]&m[258]&~m[259]&~m[260]&m[261])|(m[36]&~m[258]&m[259]&~m[260]&m[261])|(~m[36]&m[258]&m[259]&~m[260]&m[261])|(m[36]&~m[258]&~m[259]&m[260]&m[261])|(~m[36]&m[258]&~m[259]&m[260]&m[261])|(~m[36]&~m[258]&m[259]&m[260]&m[261]))&~BiasedRNG[16])|((m[36]&m[258]&m[259]&m[260]&~m[261])|(m[36]&m[258]&m[259]&~m[260]&m[261])|(m[36]&m[258]&~m[259]&m[260]&m[261])|(m[36]&~m[258]&m[259]&m[260]&m[261])|(~m[36]&m[258]&m[259]&m[260]&m[261])|(m[36]&m[258]&m[259]&m[260]&m[261]))):InitCond[44];
    m[82] = run?((((m[36]&m[262]&~m[263]&~m[264]&~m[265])|(m[36]&~m[262]&m[263]&~m[264]&~m[265])|(~m[36]&m[262]&m[263]&~m[264]&~m[265])|(m[36]&~m[262]&~m[263]&m[264]&~m[265])|(~m[36]&m[262]&~m[263]&m[264]&~m[265])|(~m[36]&~m[262]&m[263]&m[264]&~m[265])|(m[36]&~m[262]&~m[263]&~m[264]&m[265])|(~m[36]&m[262]&~m[263]&~m[264]&m[265])|(~m[36]&~m[262]&m[263]&~m[264]&m[265])|(~m[36]&~m[262]&~m[263]&m[264]&m[265]))&BiasedRNG[17])|(((m[36]&m[262]&m[263]&~m[264]&~m[265])|(m[36]&m[262]&~m[263]&m[264]&~m[265])|(m[36]&~m[262]&m[263]&m[264]&~m[265])|(~m[36]&m[262]&m[263]&m[264]&~m[265])|(m[36]&m[262]&~m[263]&~m[264]&m[265])|(m[36]&~m[262]&m[263]&~m[264]&m[265])|(~m[36]&m[262]&m[263]&~m[264]&m[265])|(m[36]&~m[262]&~m[263]&m[264]&m[265])|(~m[36]&m[262]&~m[263]&m[264]&m[265])|(~m[36]&~m[262]&m[263]&m[264]&m[265]))&~BiasedRNG[17])|((m[36]&m[262]&m[263]&m[264]&~m[265])|(m[36]&m[262]&m[263]&~m[264]&m[265])|(m[36]&m[262]&~m[263]&m[264]&m[265])|(m[36]&~m[262]&m[263]&m[264]&m[265])|(~m[36]&m[262]&m[263]&m[264]&m[265])|(m[36]&m[262]&m[263]&m[264]&m[265]))):InitCond[45];
    m[84] = run?((((m[37]&m[272]&~m[273]&~m[274]&~m[275])|(m[37]&~m[272]&m[273]&~m[274]&~m[275])|(~m[37]&m[272]&m[273]&~m[274]&~m[275])|(m[37]&~m[272]&~m[273]&m[274]&~m[275])|(~m[37]&m[272]&~m[273]&m[274]&~m[275])|(~m[37]&~m[272]&m[273]&m[274]&~m[275])|(m[37]&~m[272]&~m[273]&~m[274]&m[275])|(~m[37]&m[272]&~m[273]&~m[274]&m[275])|(~m[37]&~m[272]&m[273]&~m[274]&m[275])|(~m[37]&~m[272]&~m[273]&m[274]&m[275]))&BiasedRNG[18])|(((m[37]&m[272]&m[273]&~m[274]&~m[275])|(m[37]&m[272]&~m[273]&m[274]&~m[275])|(m[37]&~m[272]&m[273]&m[274]&~m[275])|(~m[37]&m[272]&m[273]&m[274]&~m[275])|(m[37]&m[272]&~m[273]&~m[274]&m[275])|(m[37]&~m[272]&m[273]&~m[274]&m[275])|(~m[37]&m[272]&m[273]&~m[274]&m[275])|(m[37]&~m[272]&~m[273]&m[274]&m[275])|(~m[37]&m[272]&~m[273]&m[274]&m[275])|(~m[37]&~m[272]&m[273]&m[274]&m[275]))&~BiasedRNG[18])|((m[37]&m[272]&m[273]&m[274]&~m[275])|(m[37]&m[272]&m[273]&~m[274]&m[275])|(m[37]&m[272]&~m[273]&m[274]&m[275])|(m[37]&~m[272]&m[273]&m[274]&m[275])|(~m[37]&m[272]&m[273]&m[274]&m[275])|(m[37]&m[272]&m[273]&m[274]&m[275]))):InitCond[46];
    m[85] = run?((((m[37]&m[276]&~m[277]&~m[278]&~m[279])|(m[37]&~m[276]&m[277]&~m[278]&~m[279])|(~m[37]&m[276]&m[277]&~m[278]&~m[279])|(m[37]&~m[276]&~m[277]&m[278]&~m[279])|(~m[37]&m[276]&~m[277]&m[278]&~m[279])|(~m[37]&~m[276]&m[277]&m[278]&~m[279])|(m[37]&~m[276]&~m[277]&~m[278]&m[279])|(~m[37]&m[276]&~m[277]&~m[278]&m[279])|(~m[37]&~m[276]&m[277]&~m[278]&m[279])|(~m[37]&~m[276]&~m[277]&m[278]&m[279]))&BiasedRNG[19])|(((m[37]&m[276]&m[277]&~m[278]&~m[279])|(m[37]&m[276]&~m[277]&m[278]&~m[279])|(m[37]&~m[276]&m[277]&m[278]&~m[279])|(~m[37]&m[276]&m[277]&m[278]&~m[279])|(m[37]&m[276]&~m[277]&~m[278]&m[279])|(m[37]&~m[276]&m[277]&~m[278]&m[279])|(~m[37]&m[276]&m[277]&~m[278]&m[279])|(m[37]&~m[276]&~m[277]&m[278]&m[279])|(~m[37]&m[276]&~m[277]&m[278]&m[279])|(~m[37]&~m[276]&m[277]&m[278]&m[279]))&~BiasedRNG[19])|((m[37]&m[276]&m[277]&m[278]&~m[279])|(m[37]&m[276]&m[277]&~m[278]&m[279])|(m[37]&m[276]&~m[277]&m[278]&m[279])|(m[37]&~m[276]&m[277]&m[278]&m[279])|(~m[37]&m[276]&m[277]&m[278]&m[279])|(m[37]&m[276]&m[277]&m[278]&m[279]))):InitCond[47];
    m[87] = run?((((m[38]&m[286]&~m[287]&~m[288]&~m[289])|(m[38]&~m[286]&m[287]&~m[288]&~m[289])|(~m[38]&m[286]&m[287]&~m[288]&~m[289])|(m[38]&~m[286]&~m[287]&m[288]&~m[289])|(~m[38]&m[286]&~m[287]&m[288]&~m[289])|(~m[38]&~m[286]&m[287]&m[288]&~m[289])|(m[38]&~m[286]&~m[287]&~m[288]&m[289])|(~m[38]&m[286]&~m[287]&~m[288]&m[289])|(~m[38]&~m[286]&m[287]&~m[288]&m[289])|(~m[38]&~m[286]&~m[287]&m[288]&m[289]))&BiasedRNG[20])|(((m[38]&m[286]&m[287]&~m[288]&~m[289])|(m[38]&m[286]&~m[287]&m[288]&~m[289])|(m[38]&~m[286]&m[287]&m[288]&~m[289])|(~m[38]&m[286]&m[287]&m[288]&~m[289])|(m[38]&m[286]&~m[287]&~m[288]&m[289])|(m[38]&~m[286]&m[287]&~m[288]&m[289])|(~m[38]&m[286]&m[287]&~m[288]&m[289])|(m[38]&~m[286]&~m[287]&m[288]&m[289])|(~m[38]&m[286]&~m[287]&m[288]&m[289])|(~m[38]&~m[286]&m[287]&m[288]&m[289]))&~BiasedRNG[20])|((m[38]&m[286]&m[287]&m[288]&~m[289])|(m[38]&m[286]&m[287]&~m[288]&m[289])|(m[38]&m[286]&~m[287]&m[288]&m[289])|(m[38]&~m[286]&m[287]&m[288]&m[289])|(~m[38]&m[286]&m[287]&m[288]&m[289])|(m[38]&m[286]&m[287]&m[288]&m[289]))):InitCond[48];
    m[88] = run?((((m[38]&m[290]&~m[291]&~m[292]&~m[293])|(m[38]&~m[290]&m[291]&~m[292]&~m[293])|(~m[38]&m[290]&m[291]&~m[292]&~m[293])|(m[38]&~m[290]&~m[291]&m[292]&~m[293])|(~m[38]&m[290]&~m[291]&m[292]&~m[293])|(~m[38]&~m[290]&m[291]&m[292]&~m[293])|(m[38]&~m[290]&~m[291]&~m[292]&m[293])|(~m[38]&m[290]&~m[291]&~m[292]&m[293])|(~m[38]&~m[290]&m[291]&~m[292]&m[293])|(~m[38]&~m[290]&~m[291]&m[292]&m[293]))&BiasedRNG[21])|(((m[38]&m[290]&m[291]&~m[292]&~m[293])|(m[38]&m[290]&~m[291]&m[292]&~m[293])|(m[38]&~m[290]&m[291]&m[292]&~m[293])|(~m[38]&m[290]&m[291]&m[292]&~m[293])|(m[38]&m[290]&~m[291]&~m[292]&m[293])|(m[38]&~m[290]&m[291]&~m[292]&m[293])|(~m[38]&m[290]&m[291]&~m[292]&m[293])|(m[38]&~m[290]&~m[291]&m[292]&m[293])|(~m[38]&m[290]&~m[291]&m[292]&m[293])|(~m[38]&~m[290]&m[291]&m[292]&m[293]))&~BiasedRNG[21])|((m[38]&m[290]&m[291]&m[292]&~m[293])|(m[38]&m[290]&m[291]&~m[292]&m[293])|(m[38]&m[290]&~m[291]&m[292]&m[293])|(m[38]&~m[290]&m[291]&m[292]&m[293])|(~m[38]&m[290]&m[291]&m[292]&m[293])|(m[38]&m[290]&m[291]&m[292]&m[293]))):InitCond[49];
    m[90] = run?((((m[39]&m[300]&~m[301]&~m[302]&~m[303])|(m[39]&~m[300]&m[301]&~m[302]&~m[303])|(~m[39]&m[300]&m[301]&~m[302]&~m[303])|(m[39]&~m[300]&~m[301]&m[302]&~m[303])|(~m[39]&m[300]&~m[301]&m[302]&~m[303])|(~m[39]&~m[300]&m[301]&m[302]&~m[303])|(m[39]&~m[300]&~m[301]&~m[302]&m[303])|(~m[39]&m[300]&~m[301]&~m[302]&m[303])|(~m[39]&~m[300]&m[301]&~m[302]&m[303])|(~m[39]&~m[300]&~m[301]&m[302]&m[303]))&BiasedRNG[22])|(((m[39]&m[300]&m[301]&~m[302]&~m[303])|(m[39]&m[300]&~m[301]&m[302]&~m[303])|(m[39]&~m[300]&m[301]&m[302]&~m[303])|(~m[39]&m[300]&m[301]&m[302]&~m[303])|(m[39]&m[300]&~m[301]&~m[302]&m[303])|(m[39]&~m[300]&m[301]&~m[302]&m[303])|(~m[39]&m[300]&m[301]&~m[302]&m[303])|(m[39]&~m[300]&~m[301]&m[302]&m[303])|(~m[39]&m[300]&~m[301]&m[302]&m[303])|(~m[39]&~m[300]&m[301]&m[302]&m[303]))&~BiasedRNG[22])|((m[39]&m[300]&m[301]&m[302]&~m[303])|(m[39]&m[300]&m[301]&~m[302]&m[303])|(m[39]&m[300]&~m[301]&m[302]&m[303])|(m[39]&~m[300]&m[301]&m[302]&m[303])|(~m[39]&m[300]&m[301]&m[302]&m[303])|(m[39]&m[300]&m[301]&m[302]&m[303]))):InitCond[50];
    m[91] = run?((((m[39]&m[304]&~m[305]&~m[306]&~m[307])|(m[39]&~m[304]&m[305]&~m[306]&~m[307])|(~m[39]&m[304]&m[305]&~m[306]&~m[307])|(m[39]&~m[304]&~m[305]&m[306]&~m[307])|(~m[39]&m[304]&~m[305]&m[306]&~m[307])|(~m[39]&~m[304]&m[305]&m[306]&~m[307])|(m[39]&~m[304]&~m[305]&~m[306]&m[307])|(~m[39]&m[304]&~m[305]&~m[306]&m[307])|(~m[39]&~m[304]&m[305]&~m[306]&m[307])|(~m[39]&~m[304]&~m[305]&m[306]&m[307]))&BiasedRNG[23])|(((m[39]&m[304]&m[305]&~m[306]&~m[307])|(m[39]&m[304]&~m[305]&m[306]&~m[307])|(m[39]&~m[304]&m[305]&m[306]&~m[307])|(~m[39]&m[304]&m[305]&m[306]&~m[307])|(m[39]&m[304]&~m[305]&~m[306]&m[307])|(m[39]&~m[304]&m[305]&~m[306]&m[307])|(~m[39]&m[304]&m[305]&~m[306]&m[307])|(m[39]&~m[304]&~m[305]&m[306]&m[307])|(~m[39]&m[304]&~m[305]&m[306]&m[307])|(~m[39]&~m[304]&m[305]&m[306]&m[307]))&~BiasedRNG[23])|((m[39]&m[304]&m[305]&m[306]&~m[307])|(m[39]&m[304]&m[305]&~m[306]&m[307])|(m[39]&m[304]&~m[305]&m[306]&m[307])|(m[39]&~m[304]&m[305]&m[306]&m[307])|(~m[39]&m[304]&m[305]&m[306]&m[307])|(m[39]&m[304]&m[305]&m[306]&m[307]))):InitCond[51];
    m[93] = run?((((m[40]&m[314]&~m[315]&~m[316]&~m[317])|(m[40]&~m[314]&m[315]&~m[316]&~m[317])|(~m[40]&m[314]&m[315]&~m[316]&~m[317])|(m[40]&~m[314]&~m[315]&m[316]&~m[317])|(~m[40]&m[314]&~m[315]&m[316]&~m[317])|(~m[40]&~m[314]&m[315]&m[316]&~m[317])|(m[40]&~m[314]&~m[315]&~m[316]&m[317])|(~m[40]&m[314]&~m[315]&~m[316]&m[317])|(~m[40]&~m[314]&m[315]&~m[316]&m[317])|(~m[40]&~m[314]&~m[315]&m[316]&m[317]))&BiasedRNG[24])|(((m[40]&m[314]&m[315]&~m[316]&~m[317])|(m[40]&m[314]&~m[315]&m[316]&~m[317])|(m[40]&~m[314]&m[315]&m[316]&~m[317])|(~m[40]&m[314]&m[315]&m[316]&~m[317])|(m[40]&m[314]&~m[315]&~m[316]&m[317])|(m[40]&~m[314]&m[315]&~m[316]&m[317])|(~m[40]&m[314]&m[315]&~m[316]&m[317])|(m[40]&~m[314]&~m[315]&m[316]&m[317])|(~m[40]&m[314]&~m[315]&m[316]&m[317])|(~m[40]&~m[314]&m[315]&m[316]&m[317]))&~BiasedRNG[24])|((m[40]&m[314]&m[315]&m[316]&~m[317])|(m[40]&m[314]&m[315]&~m[316]&m[317])|(m[40]&m[314]&~m[315]&m[316]&m[317])|(m[40]&~m[314]&m[315]&m[316]&m[317])|(~m[40]&m[314]&m[315]&m[316]&m[317])|(m[40]&m[314]&m[315]&m[316]&m[317]))):InitCond[52];
    m[94] = run?((((m[40]&m[318]&~m[319]&~m[320]&~m[321])|(m[40]&~m[318]&m[319]&~m[320]&~m[321])|(~m[40]&m[318]&m[319]&~m[320]&~m[321])|(m[40]&~m[318]&~m[319]&m[320]&~m[321])|(~m[40]&m[318]&~m[319]&m[320]&~m[321])|(~m[40]&~m[318]&m[319]&m[320]&~m[321])|(m[40]&~m[318]&~m[319]&~m[320]&m[321])|(~m[40]&m[318]&~m[319]&~m[320]&m[321])|(~m[40]&~m[318]&m[319]&~m[320]&m[321])|(~m[40]&~m[318]&~m[319]&m[320]&m[321]))&BiasedRNG[25])|(((m[40]&m[318]&m[319]&~m[320]&~m[321])|(m[40]&m[318]&~m[319]&m[320]&~m[321])|(m[40]&~m[318]&m[319]&m[320]&~m[321])|(~m[40]&m[318]&m[319]&m[320]&~m[321])|(m[40]&m[318]&~m[319]&~m[320]&m[321])|(m[40]&~m[318]&m[319]&~m[320]&m[321])|(~m[40]&m[318]&m[319]&~m[320]&m[321])|(m[40]&~m[318]&~m[319]&m[320]&m[321])|(~m[40]&m[318]&~m[319]&m[320]&m[321])|(~m[40]&~m[318]&m[319]&m[320]&m[321]))&~BiasedRNG[25])|((m[40]&m[318]&m[319]&m[320]&~m[321])|(m[40]&m[318]&m[319]&~m[320]&m[321])|(m[40]&m[318]&~m[319]&m[320]&m[321])|(m[40]&~m[318]&m[319]&m[320]&m[321])|(~m[40]&m[318]&m[319]&m[320]&m[321])|(m[40]&m[318]&m[319]&m[320]&m[321]))):InitCond[53];
    m[96] = run?((((m[41]&m[328]&~m[329]&~m[330]&~m[331])|(m[41]&~m[328]&m[329]&~m[330]&~m[331])|(~m[41]&m[328]&m[329]&~m[330]&~m[331])|(m[41]&~m[328]&~m[329]&m[330]&~m[331])|(~m[41]&m[328]&~m[329]&m[330]&~m[331])|(~m[41]&~m[328]&m[329]&m[330]&~m[331])|(m[41]&~m[328]&~m[329]&~m[330]&m[331])|(~m[41]&m[328]&~m[329]&~m[330]&m[331])|(~m[41]&~m[328]&m[329]&~m[330]&m[331])|(~m[41]&~m[328]&~m[329]&m[330]&m[331]))&BiasedRNG[26])|(((m[41]&m[328]&m[329]&~m[330]&~m[331])|(m[41]&m[328]&~m[329]&m[330]&~m[331])|(m[41]&~m[328]&m[329]&m[330]&~m[331])|(~m[41]&m[328]&m[329]&m[330]&~m[331])|(m[41]&m[328]&~m[329]&~m[330]&m[331])|(m[41]&~m[328]&m[329]&~m[330]&m[331])|(~m[41]&m[328]&m[329]&~m[330]&m[331])|(m[41]&~m[328]&~m[329]&m[330]&m[331])|(~m[41]&m[328]&~m[329]&m[330]&m[331])|(~m[41]&~m[328]&m[329]&m[330]&m[331]))&~BiasedRNG[26])|((m[41]&m[328]&m[329]&m[330]&~m[331])|(m[41]&m[328]&m[329]&~m[330]&m[331])|(m[41]&m[328]&~m[329]&m[330]&m[331])|(m[41]&~m[328]&m[329]&m[330]&m[331])|(~m[41]&m[328]&m[329]&m[330]&m[331])|(m[41]&m[328]&m[329]&m[330]&m[331]))):InitCond[54];
    m[97] = run?((((m[41]&m[332]&~m[333]&~m[334]&~m[335])|(m[41]&~m[332]&m[333]&~m[334]&~m[335])|(~m[41]&m[332]&m[333]&~m[334]&~m[335])|(m[41]&~m[332]&~m[333]&m[334]&~m[335])|(~m[41]&m[332]&~m[333]&m[334]&~m[335])|(~m[41]&~m[332]&m[333]&m[334]&~m[335])|(m[41]&~m[332]&~m[333]&~m[334]&m[335])|(~m[41]&m[332]&~m[333]&~m[334]&m[335])|(~m[41]&~m[332]&m[333]&~m[334]&m[335])|(~m[41]&~m[332]&~m[333]&m[334]&m[335]))&BiasedRNG[27])|(((m[41]&m[332]&m[333]&~m[334]&~m[335])|(m[41]&m[332]&~m[333]&m[334]&~m[335])|(m[41]&~m[332]&m[333]&m[334]&~m[335])|(~m[41]&m[332]&m[333]&m[334]&~m[335])|(m[41]&m[332]&~m[333]&~m[334]&m[335])|(m[41]&~m[332]&m[333]&~m[334]&m[335])|(~m[41]&m[332]&m[333]&~m[334]&m[335])|(m[41]&~m[332]&~m[333]&m[334]&m[335])|(~m[41]&m[332]&~m[333]&m[334]&m[335])|(~m[41]&~m[332]&m[333]&m[334]&m[335]))&~BiasedRNG[27])|((m[41]&m[332]&m[333]&m[334]&~m[335])|(m[41]&m[332]&m[333]&~m[334]&m[335])|(m[41]&m[332]&~m[333]&m[334]&m[335])|(m[41]&~m[332]&m[333]&m[334]&m[335])|(~m[41]&m[332]&m[333]&m[334]&m[335])|(m[41]&m[332]&m[333]&m[334]&m[335]))):InitCond[55];
    m[99] = run?((((m[42]&m[342]&~m[343]&~m[344]&~m[345])|(m[42]&~m[342]&m[343]&~m[344]&~m[345])|(~m[42]&m[342]&m[343]&~m[344]&~m[345])|(m[42]&~m[342]&~m[343]&m[344]&~m[345])|(~m[42]&m[342]&~m[343]&m[344]&~m[345])|(~m[42]&~m[342]&m[343]&m[344]&~m[345])|(m[42]&~m[342]&~m[343]&~m[344]&m[345])|(~m[42]&m[342]&~m[343]&~m[344]&m[345])|(~m[42]&~m[342]&m[343]&~m[344]&m[345])|(~m[42]&~m[342]&~m[343]&m[344]&m[345]))&BiasedRNG[28])|(((m[42]&m[342]&m[343]&~m[344]&~m[345])|(m[42]&m[342]&~m[343]&m[344]&~m[345])|(m[42]&~m[342]&m[343]&m[344]&~m[345])|(~m[42]&m[342]&m[343]&m[344]&~m[345])|(m[42]&m[342]&~m[343]&~m[344]&m[345])|(m[42]&~m[342]&m[343]&~m[344]&m[345])|(~m[42]&m[342]&m[343]&~m[344]&m[345])|(m[42]&~m[342]&~m[343]&m[344]&m[345])|(~m[42]&m[342]&~m[343]&m[344]&m[345])|(~m[42]&~m[342]&m[343]&m[344]&m[345]))&~BiasedRNG[28])|((m[42]&m[342]&m[343]&m[344]&~m[345])|(m[42]&m[342]&m[343]&~m[344]&m[345])|(m[42]&m[342]&~m[343]&m[344]&m[345])|(m[42]&~m[342]&m[343]&m[344]&m[345])|(~m[42]&m[342]&m[343]&m[344]&m[345])|(m[42]&m[342]&m[343]&m[344]&m[345]))):InitCond[56];
    m[100] = run?((((m[42]&m[346]&~m[347]&~m[348]&~m[349])|(m[42]&~m[346]&m[347]&~m[348]&~m[349])|(~m[42]&m[346]&m[347]&~m[348]&~m[349])|(m[42]&~m[346]&~m[347]&m[348]&~m[349])|(~m[42]&m[346]&~m[347]&m[348]&~m[349])|(~m[42]&~m[346]&m[347]&m[348]&~m[349])|(m[42]&~m[346]&~m[347]&~m[348]&m[349])|(~m[42]&m[346]&~m[347]&~m[348]&m[349])|(~m[42]&~m[346]&m[347]&~m[348]&m[349])|(~m[42]&~m[346]&~m[347]&m[348]&m[349]))&BiasedRNG[29])|(((m[42]&m[346]&m[347]&~m[348]&~m[349])|(m[42]&m[346]&~m[347]&m[348]&~m[349])|(m[42]&~m[346]&m[347]&m[348]&~m[349])|(~m[42]&m[346]&m[347]&m[348]&~m[349])|(m[42]&m[346]&~m[347]&~m[348]&m[349])|(m[42]&~m[346]&m[347]&~m[348]&m[349])|(~m[42]&m[346]&m[347]&~m[348]&m[349])|(m[42]&~m[346]&~m[347]&m[348]&m[349])|(~m[42]&m[346]&~m[347]&m[348]&m[349])|(~m[42]&~m[346]&m[347]&m[348]&m[349]))&~BiasedRNG[29])|((m[42]&m[346]&m[347]&m[348]&~m[349])|(m[42]&m[346]&m[347]&~m[348]&m[349])|(m[42]&m[346]&~m[347]&m[348]&m[349])|(m[42]&~m[346]&m[347]&m[348]&m[349])|(~m[42]&m[346]&m[347]&m[348]&m[349])|(m[42]&m[346]&m[347]&m[348]&m[349]))):InitCond[57];
    m[102] = run?((((m[43]&m[356]&~m[357]&~m[358]&~m[359])|(m[43]&~m[356]&m[357]&~m[358]&~m[359])|(~m[43]&m[356]&m[357]&~m[358]&~m[359])|(m[43]&~m[356]&~m[357]&m[358]&~m[359])|(~m[43]&m[356]&~m[357]&m[358]&~m[359])|(~m[43]&~m[356]&m[357]&m[358]&~m[359])|(m[43]&~m[356]&~m[357]&~m[358]&m[359])|(~m[43]&m[356]&~m[357]&~m[358]&m[359])|(~m[43]&~m[356]&m[357]&~m[358]&m[359])|(~m[43]&~m[356]&~m[357]&m[358]&m[359]))&BiasedRNG[30])|(((m[43]&m[356]&m[357]&~m[358]&~m[359])|(m[43]&m[356]&~m[357]&m[358]&~m[359])|(m[43]&~m[356]&m[357]&m[358]&~m[359])|(~m[43]&m[356]&m[357]&m[358]&~m[359])|(m[43]&m[356]&~m[357]&~m[358]&m[359])|(m[43]&~m[356]&m[357]&~m[358]&m[359])|(~m[43]&m[356]&m[357]&~m[358]&m[359])|(m[43]&~m[356]&~m[357]&m[358]&m[359])|(~m[43]&m[356]&~m[357]&m[358]&m[359])|(~m[43]&~m[356]&m[357]&m[358]&m[359]))&~BiasedRNG[30])|((m[43]&m[356]&m[357]&m[358]&~m[359])|(m[43]&m[356]&m[357]&~m[358]&m[359])|(m[43]&m[356]&~m[357]&m[358]&m[359])|(m[43]&~m[356]&m[357]&m[358]&m[359])|(~m[43]&m[356]&m[357]&m[358]&m[359])|(m[43]&m[356]&m[357]&m[358]&m[359]))):InitCond[58];
    m[103] = run?((((m[43]&m[360]&~m[361]&~m[362]&~m[363])|(m[43]&~m[360]&m[361]&~m[362]&~m[363])|(~m[43]&m[360]&m[361]&~m[362]&~m[363])|(m[43]&~m[360]&~m[361]&m[362]&~m[363])|(~m[43]&m[360]&~m[361]&m[362]&~m[363])|(~m[43]&~m[360]&m[361]&m[362]&~m[363])|(m[43]&~m[360]&~m[361]&~m[362]&m[363])|(~m[43]&m[360]&~m[361]&~m[362]&m[363])|(~m[43]&~m[360]&m[361]&~m[362]&m[363])|(~m[43]&~m[360]&~m[361]&m[362]&m[363]))&BiasedRNG[31])|(((m[43]&m[360]&m[361]&~m[362]&~m[363])|(m[43]&m[360]&~m[361]&m[362]&~m[363])|(m[43]&~m[360]&m[361]&m[362]&~m[363])|(~m[43]&m[360]&m[361]&m[362]&~m[363])|(m[43]&m[360]&~m[361]&~m[362]&m[363])|(m[43]&~m[360]&m[361]&~m[362]&m[363])|(~m[43]&m[360]&m[361]&~m[362]&m[363])|(m[43]&~m[360]&~m[361]&m[362]&m[363])|(~m[43]&m[360]&~m[361]&m[362]&m[363])|(~m[43]&~m[360]&m[361]&m[362]&m[363]))&~BiasedRNG[31])|((m[43]&m[360]&m[361]&m[362]&~m[363])|(m[43]&m[360]&m[361]&~m[362]&m[363])|(m[43]&m[360]&~m[361]&m[362]&m[363])|(m[43]&~m[360]&m[361]&m[362]&m[363])|(~m[43]&m[360]&m[361]&m[362]&m[363])|(m[43]&m[360]&m[361]&m[362]&m[363]))):InitCond[59];
    m[105] = run?((((m[44]&m[370]&~m[371]&~m[372]&~m[373])|(m[44]&~m[370]&m[371]&~m[372]&~m[373])|(~m[44]&m[370]&m[371]&~m[372]&~m[373])|(m[44]&~m[370]&~m[371]&m[372]&~m[373])|(~m[44]&m[370]&~m[371]&m[372]&~m[373])|(~m[44]&~m[370]&m[371]&m[372]&~m[373])|(m[44]&~m[370]&~m[371]&~m[372]&m[373])|(~m[44]&m[370]&~m[371]&~m[372]&m[373])|(~m[44]&~m[370]&m[371]&~m[372]&m[373])|(~m[44]&~m[370]&~m[371]&m[372]&m[373]))&BiasedRNG[32])|(((m[44]&m[370]&m[371]&~m[372]&~m[373])|(m[44]&m[370]&~m[371]&m[372]&~m[373])|(m[44]&~m[370]&m[371]&m[372]&~m[373])|(~m[44]&m[370]&m[371]&m[372]&~m[373])|(m[44]&m[370]&~m[371]&~m[372]&m[373])|(m[44]&~m[370]&m[371]&~m[372]&m[373])|(~m[44]&m[370]&m[371]&~m[372]&m[373])|(m[44]&~m[370]&~m[371]&m[372]&m[373])|(~m[44]&m[370]&~m[371]&m[372]&m[373])|(~m[44]&~m[370]&m[371]&m[372]&m[373]))&~BiasedRNG[32])|((m[44]&m[370]&m[371]&m[372]&~m[373])|(m[44]&m[370]&m[371]&~m[372]&m[373])|(m[44]&m[370]&~m[371]&m[372]&m[373])|(m[44]&~m[370]&m[371]&m[372]&m[373])|(~m[44]&m[370]&m[371]&m[372]&m[373])|(m[44]&m[370]&m[371]&m[372]&m[373]))):InitCond[60];
    m[106] = run?((((m[44]&m[374]&~m[375]&~m[376]&~m[377])|(m[44]&~m[374]&m[375]&~m[376]&~m[377])|(~m[44]&m[374]&m[375]&~m[376]&~m[377])|(m[44]&~m[374]&~m[375]&m[376]&~m[377])|(~m[44]&m[374]&~m[375]&m[376]&~m[377])|(~m[44]&~m[374]&m[375]&m[376]&~m[377])|(m[44]&~m[374]&~m[375]&~m[376]&m[377])|(~m[44]&m[374]&~m[375]&~m[376]&m[377])|(~m[44]&~m[374]&m[375]&~m[376]&m[377])|(~m[44]&~m[374]&~m[375]&m[376]&m[377]))&BiasedRNG[33])|(((m[44]&m[374]&m[375]&~m[376]&~m[377])|(m[44]&m[374]&~m[375]&m[376]&~m[377])|(m[44]&~m[374]&m[375]&m[376]&~m[377])|(~m[44]&m[374]&m[375]&m[376]&~m[377])|(m[44]&m[374]&~m[375]&~m[376]&m[377])|(m[44]&~m[374]&m[375]&~m[376]&m[377])|(~m[44]&m[374]&m[375]&~m[376]&m[377])|(m[44]&~m[374]&~m[375]&m[376]&m[377])|(~m[44]&m[374]&~m[375]&m[376]&m[377])|(~m[44]&~m[374]&m[375]&m[376]&m[377]))&~BiasedRNG[33])|((m[44]&m[374]&m[375]&m[376]&~m[377])|(m[44]&m[374]&m[375]&~m[376]&m[377])|(m[44]&m[374]&~m[375]&m[376]&m[377])|(m[44]&~m[374]&m[375]&m[376]&m[377])|(~m[44]&m[374]&m[375]&m[376]&m[377])|(m[44]&m[374]&m[375]&m[376]&m[377]))):InitCond[61];
    m[108] = run?((((m[45]&m[384]&~m[385]&~m[386]&~m[387])|(m[45]&~m[384]&m[385]&~m[386]&~m[387])|(~m[45]&m[384]&m[385]&~m[386]&~m[387])|(m[45]&~m[384]&~m[385]&m[386]&~m[387])|(~m[45]&m[384]&~m[385]&m[386]&~m[387])|(~m[45]&~m[384]&m[385]&m[386]&~m[387])|(m[45]&~m[384]&~m[385]&~m[386]&m[387])|(~m[45]&m[384]&~m[385]&~m[386]&m[387])|(~m[45]&~m[384]&m[385]&~m[386]&m[387])|(~m[45]&~m[384]&~m[385]&m[386]&m[387]))&BiasedRNG[34])|(((m[45]&m[384]&m[385]&~m[386]&~m[387])|(m[45]&m[384]&~m[385]&m[386]&~m[387])|(m[45]&~m[384]&m[385]&m[386]&~m[387])|(~m[45]&m[384]&m[385]&m[386]&~m[387])|(m[45]&m[384]&~m[385]&~m[386]&m[387])|(m[45]&~m[384]&m[385]&~m[386]&m[387])|(~m[45]&m[384]&m[385]&~m[386]&m[387])|(m[45]&~m[384]&~m[385]&m[386]&m[387])|(~m[45]&m[384]&~m[385]&m[386]&m[387])|(~m[45]&~m[384]&m[385]&m[386]&m[387]))&~BiasedRNG[34])|((m[45]&m[384]&m[385]&m[386]&~m[387])|(m[45]&m[384]&m[385]&~m[386]&m[387])|(m[45]&m[384]&~m[385]&m[386]&m[387])|(m[45]&~m[384]&m[385]&m[386]&m[387])|(~m[45]&m[384]&m[385]&m[386]&m[387])|(m[45]&m[384]&m[385]&m[386]&m[387]))):InitCond[62];
    m[109] = run?((((m[45]&m[388]&~m[389]&~m[390]&~m[391])|(m[45]&~m[388]&m[389]&~m[390]&~m[391])|(~m[45]&m[388]&m[389]&~m[390]&~m[391])|(m[45]&~m[388]&~m[389]&m[390]&~m[391])|(~m[45]&m[388]&~m[389]&m[390]&~m[391])|(~m[45]&~m[388]&m[389]&m[390]&~m[391])|(m[45]&~m[388]&~m[389]&~m[390]&m[391])|(~m[45]&m[388]&~m[389]&~m[390]&m[391])|(~m[45]&~m[388]&m[389]&~m[390]&m[391])|(~m[45]&~m[388]&~m[389]&m[390]&m[391]))&BiasedRNG[35])|(((m[45]&m[388]&m[389]&~m[390]&~m[391])|(m[45]&m[388]&~m[389]&m[390]&~m[391])|(m[45]&~m[388]&m[389]&m[390]&~m[391])|(~m[45]&m[388]&m[389]&m[390]&~m[391])|(m[45]&m[388]&~m[389]&~m[390]&m[391])|(m[45]&~m[388]&m[389]&~m[390]&m[391])|(~m[45]&m[388]&m[389]&~m[390]&m[391])|(m[45]&~m[388]&~m[389]&m[390]&m[391])|(~m[45]&m[388]&~m[389]&m[390]&m[391])|(~m[45]&~m[388]&m[389]&m[390]&m[391]))&~BiasedRNG[35])|((m[45]&m[388]&m[389]&m[390]&~m[391])|(m[45]&m[388]&m[389]&~m[390]&m[391])|(m[45]&m[388]&~m[389]&m[390]&m[391])|(m[45]&~m[388]&m[389]&m[390]&m[391])|(~m[45]&m[388]&m[389]&m[390]&m[391])|(m[45]&m[388]&m[389]&m[390]&m[391]))):InitCond[63];
    m[111] = run?((((m[46]&m[398]&~m[399]&~m[400]&~m[401])|(m[46]&~m[398]&m[399]&~m[400]&~m[401])|(~m[46]&m[398]&m[399]&~m[400]&~m[401])|(m[46]&~m[398]&~m[399]&m[400]&~m[401])|(~m[46]&m[398]&~m[399]&m[400]&~m[401])|(~m[46]&~m[398]&m[399]&m[400]&~m[401])|(m[46]&~m[398]&~m[399]&~m[400]&m[401])|(~m[46]&m[398]&~m[399]&~m[400]&m[401])|(~m[46]&~m[398]&m[399]&~m[400]&m[401])|(~m[46]&~m[398]&~m[399]&m[400]&m[401]))&BiasedRNG[36])|(((m[46]&m[398]&m[399]&~m[400]&~m[401])|(m[46]&m[398]&~m[399]&m[400]&~m[401])|(m[46]&~m[398]&m[399]&m[400]&~m[401])|(~m[46]&m[398]&m[399]&m[400]&~m[401])|(m[46]&m[398]&~m[399]&~m[400]&m[401])|(m[46]&~m[398]&m[399]&~m[400]&m[401])|(~m[46]&m[398]&m[399]&~m[400]&m[401])|(m[46]&~m[398]&~m[399]&m[400]&m[401])|(~m[46]&m[398]&~m[399]&m[400]&m[401])|(~m[46]&~m[398]&m[399]&m[400]&m[401]))&~BiasedRNG[36])|((m[46]&m[398]&m[399]&m[400]&~m[401])|(m[46]&m[398]&m[399]&~m[400]&m[401])|(m[46]&m[398]&~m[399]&m[400]&m[401])|(m[46]&~m[398]&m[399]&m[400]&m[401])|(~m[46]&m[398]&m[399]&m[400]&m[401])|(m[46]&m[398]&m[399]&m[400]&m[401]))):InitCond[64];
    m[112] = run?((((m[46]&m[402]&~m[403]&~m[404]&~m[405])|(m[46]&~m[402]&m[403]&~m[404]&~m[405])|(~m[46]&m[402]&m[403]&~m[404]&~m[405])|(m[46]&~m[402]&~m[403]&m[404]&~m[405])|(~m[46]&m[402]&~m[403]&m[404]&~m[405])|(~m[46]&~m[402]&m[403]&m[404]&~m[405])|(m[46]&~m[402]&~m[403]&~m[404]&m[405])|(~m[46]&m[402]&~m[403]&~m[404]&m[405])|(~m[46]&~m[402]&m[403]&~m[404]&m[405])|(~m[46]&~m[402]&~m[403]&m[404]&m[405]))&BiasedRNG[37])|(((m[46]&m[402]&m[403]&~m[404]&~m[405])|(m[46]&m[402]&~m[403]&m[404]&~m[405])|(m[46]&~m[402]&m[403]&m[404]&~m[405])|(~m[46]&m[402]&m[403]&m[404]&~m[405])|(m[46]&m[402]&~m[403]&~m[404]&m[405])|(m[46]&~m[402]&m[403]&~m[404]&m[405])|(~m[46]&m[402]&m[403]&~m[404]&m[405])|(m[46]&~m[402]&~m[403]&m[404]&m[405])|(~m[46]&m[402]&~m[403]&m[404]&m[405])|(~m[46]&~m[402]&m[403]&m[404]&m[405]))&~BiasedRNG[37])|((m[46]&m[402]&m[403]&m[404]&~m[405])|(m[46]&m[402]&m[403]&~m[404]&m[405])|(m[46]&m[402]&~m[403]&m[404]&m[405])|(m[46]&~m[402]&m[403]&m[404]&m[405])|(~m[46]&m[402]&m[403]&m[404]&m[405])|(m[46]&m[402]&m[403]&m[404]&m[405]))):InitCond[65];
    m[114] = run?((((m[47]&m[412]&~m[413]&~m[414]&~m[415])|(m[47]&~m[412]&m[413]&~m[414]&~m[415])|(~m[47]&m[412]&m[413]&~m[414]&~m[415])|(m[47]&~m[412]&~m[413]&m[414]&~m[415])|(~m[47]&m[412]&~m[413]&m[414]&~m[415])|(~m[47]&~m[412]&m[413]&m[414]&~m[415])|(m[47]&~m[412]&~m[413]&~m[414]&m[415])|(~m[47]&m[412]&~m[413]&~m[414]&m[415])|(~m[47]&~m[412]&m[413]&~m[414]&m[415])|(~m[47]&~m[412]&~m[413]&m[414]&m[415]))&BiasedRNG[38])|(((m[47]&m[412]&m[413]&~m[414]&~m[415])|(m[47]&m[412]&~m[413]&m[414]&~m[415])|(m[47]&~m[412]&m[413]&m[414]&~m[415])|(~m[47]&m[412]&m[413]&m[414]&~m[415])|(m[47]&m[412]&~m[413]&~m[414]&m[415])|(m[47]&~m[412]&m[413]&~m[414]&m[415])|(~m[47]&m[412]&m[413]&~m[414]&m[415])|(m[47]&~m[412]&~m[413]&m[414]&m[415])|(~m[47]&m[412]&~m[413]&m[414]&m[415])|(~m[47]&~m[412]&m[413]&m[414]&m[415]))&~BiasedRNG[38])|((m[47]&m[412]&m[413]&m[414]&~m[415])|(m[47]&m[412]&m[413]&~m[414]&m[415])|(m[47]&m[412]&~m[413]&m[414]&m[415])|(m[47]&~m[412]&m[413]&m[414]&m[415])|(~m[47]&m[412]&m[413]&m[414]&m[415])|(m[47]&m[412]&m[413]&m[414]&m[415]))):InitCond[66];
    m[115] = run?((((m[47]&m[416]&~m[417]&~m[418]&~m[419])|(m[47]&~m[416]&m[417]&~m[418]&~m[419])|(~m[47]&m[416]&m[417]&~m[418]&~m[419])|(m[47]&~m[416]&~m[417]&m[418]&~m[419])|(~m[47]&m[416]&~m[417]&m[418]&~m[419])|(~m[47]&~m[416]&m[417]&m[418]&~m[419])|(m[47]&~m[416]&~m[417]&~m[418]&m[419])|(~m[47]&m[416]&~m[417]&~m[418]&m[419])|(~m[47]&~m[416]&m[417]&~m[418]&m[419])|(~m[47]&~m[416]&~m[417]&m[418]&m[419]))&BiasedRNG[39])|(((m[47]&m[416]&m[417]&~m[418]&~m[419])|(m[47]&m[416]&~m[417]&m[418]&~m[419])|(m[47]&~m[416]&m[417]&m[418]&~m[419])|(~m[47]&m[416]&m[417]&m[418]&~m[419])|(m[47]&m[416]&~m[417]&~m[418]&m[419])|(m[47]&~m[416]&m[417]&~m[418]&m[419])|(~m[47]&m[416]&m[417]&~m[418]&m[419])|(m[47]&~m[416]&~m[417]&m[418]&m[419])|(~m[47]&m[416]&~m[417]&m[418]&m[419])|(~m[47]&~m[416]&m[417]&m[418]&m[419]))&~BiasedRNG[39])|((m[47]&m[416]&m[417]&m[418]&~m[419])|(m[47]&m[416]&m[417]&~m[418]&m[419])|(m[47]&m[416]&~m[417]&m[418]&m[419])|(m[47]&~m[416]&m[417]&m[418]&m[419])|(~m[47]&m[416]&m[417]&m[418]&m[419])|(m[47]&m[416]&m[417]&m[418]&m[419]))):InitCond[67];
    m[117] = run?((((m[48]&m[426]&~m[427]&~m[428]&~m[429])|(m[48]&~m[426]&m[427]&~m[428]&~m[429])|(~m[48]&m[426]&m[427]&~m[428]&~m[429])|(m[48]&~m[426]&~m[427]&m[428]&~m[429])|(~m[48]&m[426]&~m[427]&m[428]&~m[429])|(~m[48]&~m[426]&m[427]&m[428]&~m[429])|(m[48]&~m[426]&~m[427]&~m[428]&m[429])|(~m[48]&m[426]&~m[427]&~m[428]&m[429])|(~m[48]&~m[426]&m[427]&~m[428]&m[429])|(~m[48]&~m[426]&~m[427]&m[428]&m[429]))&BiasedRNG[40])|(((m[48]&m[426]&m[427]&~m[428]&~m[429])|(m[48]&m[426]&~m[427]&m[428]&~m[429])|(m[48]&~m[426]&m[427]&m[428]&~m[429])|(~m[48]&m[426]&m[427]&m[428]&~m[429])|(m[48]&m[426]&~m[427]&~m[428]&m[429])|(m[48]&~m[426]&m[427]&~m[428]&m[429])|(~m[48]&m[426]&m[427]&~m[428]&m[429])|(m[48]&~m[426]&~m[427]&m[428]&m[429])|(~m[48]&m[426]&~m[427]&m[428]&m[429])|(~m[48]&~m[426]&m[427]&m[428]&m[429]))&~BiasedRNG[40])|((m[48]&m[426]&m[427]&m[428]&~m[429])|(m[48]&m[426]&m[427]&~m[428]&m[429])|(m[48]&m[426]&~m[427]&m[428]&m[429])|(m[48]&~m[426]&m[427]&m[428]&m[429])|(~m[48]&m[426]&m[427]&m[428]&m[429])|(m[48]&m[426]&m[427]&m[428]&m[429]))):InitCond[68];
    m[118] = run?((((m[48]&m[430]&~m[431]&~m[432]&~m[433])|(m[48]&~m[430]&m[431]&~m[432]&~m[433])|(~m[48]&m[430]&m[431]&~m[432]&~m[433])|(m[48]&~m[430]&~m[431]&m[432]&~m[433])|(~m[48]&m[430]&~m[431]&m[432]&~m[433])|(~m[48]&~m[430]&m[431]&m[432]&~m[433])|(m[48]&~m[430]&~m[431]&~m[432]&m[433])|(~m[48]&m[430]&~m[431]&~m[432]&m[433])|(~m[48]&~m[430]&m[431]&~m[432]&m[433])|(~m[48]&~m[430]&~m[431]&m[432]&m[433]))&BiasedRNG[41])|(((m[48]&m[430]&m[431]&~m[432]&~m[433])|(m[48]&m[430]&~m[431]&m[432]&~m[433])|(m[48]&~m[430]&m[431]&m[432]&~m[433])|(~m[48]&m[430]&m[431]&m[432]&~m[433])|(m[48]&m[430]&~m[431]&~m[432]&m[433])|(m[48]&~m[430]&m[431]&~m[432]&m[433])|(~m[48]&m[430]&m[431]&~m[432]&m[433])|(m[48]&~m[430]&~m[431]&m[432]&m[433])|(~m[48]&m[430]&~m[431]&m[432]&m[433])|(~m[48]&~m[430]&m[431]&m[432]&m[433]))&~BiasedRNG[41])|((m[48]&m[430]&m[431]&m[432]&~m[433])|(m[48]&m[430]&m[431]&~m[432]&m[433])|(m[48]&m[430]&~m[431]&m[432]&m[433])|(m[48]&~m[430]&m[431]&m[432]&m[433])|(~m[48]&m[430]&m[431]&m[432]&m[433])|(m[48]&m[430]&m[431]&m[432]&m[433]))):InitCond[69];
    m[120] = run?((((m[49]&m[440]&~m[441]&~m[442]&~m[443])|(m[49]&~m[440]&m[441]&~m[442]&~m[443])|(~m[49]&m[440]&m[441]&~m[442]&~m[443])|(m[49]&~m[440]&~m[441]&m[442]&~m[443])|(~m[49]&m[440]&~m[441]&m[442]&~m[443])|(~m[49]&~m[440]&m[441]&m[442]&~m[443])|(m[49]&~m[440]&~m[441]&~m[442]&m[443])|(~m[49]&m[440]&~m[441]&~m[442]&m[443])|(~m[49]&~m[440]&m[441]&~m[442]&m[443])|(~m[49]&~m[440]&~m[441]&m[442]&m[443]))&BiasedRNG[42])|(((m[49]&m[440]&m[441]&~m[442]&~m[443])|(m[49]&m[440]&~m[441]&m[442]&~m[443])|(m[49]&~m[440]&m[441]&m[442]&~m[443])|(~m[49]&m[440]&m[441]&m[442]&~m[443])|(m[49]&m[440]&~m[441]&~m[442]&m[443])|(m[49]&~m[440]&m[441]&~m[442]&m[443])|(~m[49]&m[440]&m[441]&~m[442]&m[443])|(m[49]&~m[440]&~m[441]&m[442]&m[443])|(~m[49]&m[440]&~m[441]&m[442]&m[443])|(~m[49]&~m[440]&m[441]&m[442]&m[443]))&~BiasedRNG[42])|((m[49]&m[440]&m[441]&m[442]&~m[443])|(m[49]&m[440]&m[441]&~m[442]&m[443])|(m[49]&m[440]&~m[441]&m[442]&m[443])|(m[49]&~m[440]&m[441]&m[442]&m[443])|(~m[49]&m[440]&m[441]&m[442]&m[443])|(m[49]&m[440]&m[441]&m[442]&m[443]))):InitCond[70];
    m[121] = run?((((m[49]&m[444]&~m[445]&~m[446]&~m[447])|(m[49]&~m[444]&m[445]&~m[446]&~m[447])|(~m[49]&m[444]&m[445]&~m[446]&~m[447])|(m[49]&~m[444]&~m[445]&m[446]&~m[447])|(~m[49]&m[444]&~m[445]&m[446]&~m[447])|(~m[49]&~m[444]&m[445]&m[446]&~m[447])|(m[49]&~m[444]&~m[445]&~m[446]&m[447])|(~m[49]&m[444]&~m[445]&~m[446]&m[447])|(~m[49]&~m[444]&m[445]&~m[446]&m[447])|(~m[49]&~m[444]&~m[445]&m[446]&m[447]))&BiasedRNG[43])|(((m[49]&m[444]&m[445]&~m[446]&~m[447])|(m[49]&m[444]&~m[445]&m[446]&~m[447])|(m[49]&~m[444]&m[445]&m[446]&~m[447])|(~m[49]&m[444]&m[445]&m[446]&~m[447])|(m[49]&m[444]&~m[445]&~m[446]&m[447])|(m[49]&~m[444]&m[445]&~m[446]&m[447])|(~m[49]&m[444]&m[445]&~m[446]&m[447])|(m[49]&~m[444]&~m[445]&m[446]&m[447])|(~m[49]&m[444]&~m[445]&m[446]&m[447])|(~m[49]&~m[444]&m[445]&m[446]&m[447]))&~BiasedRNG[43])|((m[49]&m[444]&m[445]&m[446]&~m[447])|(m[49]&m[444]&m[445]&~m[446]&m[447])|(m[49]&m[444]&~m[445]&m[446]&m[447])|(m[49]&~m[444]&m[445]&m[446]&m[447])|(~m[49]&m[444]&m[445]&m[446]&m[447])|(m[49]&m[444]&m[445]&m[446]&m[447]))):InitCond[71];
    m[123] = run?((((m[50]&m[454]&~m[455]&~m[456]&~m[457])|(m[50]&~m[454]&m[455]&~m[456]&~m[457])|(~m[50]&m[454]&m[455]&~m[456]&~m[457])|(m[50]&~m[454]&~m[455]&m[456]&~m[457])|(~m[50]&m[454]&~m[455]&m[456]&~m[457])|(~m[50]&~m[454]&m[455]&m[456]&~m[457])|(m[50]&~m[454]&~m[455]&~m[456]&m[457])|(~m[50]&m[454]&~m[455]&~m[456]&m[457])|(~m[50]&~m[454]&m[455]&~m[456]&m[457])|(~m[50]&~m[454]&~m[455]&m[456]&m[457]))&BiasedRNG[44])|(((m[50]&m[454]&m[455]&~m[456]&~m[457])|(m[50]&m[454]&~m[455]&m[456]&~m[457])|(m[50]&~m[454]&m[455]&m[456]&~m[457])|(~m[50]&m[454]&m[455]&m[456]&~m[457])|(m[50]&m[454]&~m[455]&~m[456]&m[457])|(m[50]&~m[454]&m[455]&~m[456]&m[457])|(~m[50]&m[454]&m[455]&~m[456]&m[457])|(m[50]&~m[454]&~m[455]&m[456]&m[457])|(~m[50]&m[454]&~m[455]&m[456]&m[457])|(~m[50]&~m[454]&m[455]&m[456]&m[457]))&~BiasedRNG[44])|((m[50]&m[454]&m[455]&m[456]&~m[457])|(m[50]&m[454]&m[455]&~m[456]&m[457])|(m[50]&m[454]&~m[455]&m[456]&m[457])|(m[50]&~m[454]&m[455]&m[456]&m[457])|(~m[50]&m[454]&m[455]&m[456]&m[457])|(m[50]&m[454]&m[455]&m[456]&m[457]))):InitCond[72];
    m[124] = run?((((m[50]&m[458]&~m[459]&~m[460]&~m[461])|(m[50]&~m[458]&m[459]&~m[460]&~m[461])|(~m[50]&m[458]&m[459]&~m[460]&~m[461])|(m[50]&~m[458]&~m[459]&m[460]&~m[461])|(~m[50]&m[458]&~m[459]&m[460]&~m[461])|(~m[50]&~m[458]&m[459]&m[460]&~m[461])|(m[50]&~m[458]&~m[459]&~m[460]&m[461])|(~m[50]&m[458]&~m[459]&~m[460]&m[461])|(~m[50]&~m[458]&m[459]&~m[460]&m[461])|(~m[50]&~m[458]&~m[459]&m[460]&m[461]))&BiasedRNG[45])|(((m[50]&m[458]&m[459]&~m[460]&~m[461])|(m[50]&m[458]&~m[459]&m[460]&~m[461])|(m[50]&~m[458]&m[459]&m[460]&~m[461])|(~m[50]&m[458]&m[459]&m[460]&~m[461])|(m[50]&m[458]&~m[459]&~m[460]&m[461])|(m[50]&~m[458]&m[459]&~m[460]&m[461])|(~m[50]&m[458]&m[459]&~m[460]&m[461])|(m[50]&~m[458]&~m[459]&m[460]&m[461])|(~m[50]&m[458]&~m[459]&m[460]&m[461])|(~m[50]&~m[458]&m[459]&m[460]&m[461]))&~BiasedRNG[45])|((m[50]&m[458]&m[459]&m[460]&~m[461])|(m[50]&m[458]&m[459]&~m[460]&m[461])|(m[50]&m[458]&~m[459]&m[460]&m[461])|(m[50]&~m[458]&m[459]&m[460]&m[461])|(~m[50]&m[458]&m[459]&m[460]&m[461])|(m[50]&m[458]&m[459]&m[460]&m[461]))):InitCond[73];
    m[126] = run?((((m[51]&m[468]&~m[469]&~m[470]&~m[471])|(m[51]&~m[468]&m[469]&~m[470]&~m[471])|(~m[51]&m[468]&m[469]&~m[470]&~m[471])|(m[51]&~m[468]&~m[469]&m[470]&~m[471])|(~m[51]&m[468]&~m[469]&m[470]&~m[471])|(~m[51]&~m[468]&m[469]&m[470]&~m[471])|(m[51]&~m[468]&~m[469]&~m[470]&m[471])|(~m[51]&m[468]&~m[469]&~m[470]&m[471])|(~m[51]&~m[468]&m[469]&~m[470]&m[471])|(~m[51]&~m[468]&~m[469]&m[470]&m[471]))&BiasedRNG[46])|(((m[51]&m[468]&m[469]&~m[470]&~m[471])|(m[51]&m[468]&~m[469]&m[470]&~m[471])|(m[51]&~m[468]&m[469]&m[470]&~m[471])|(~m[51]&m[468]&m[469]&m[470]&~m[471])|(m[51]&m[468]&~m[469]&~m[470]&m[471])|(m[51]&~m[468]&m[469]&~m[470]&m[471])|(~m[51]&m[468]&m[469]&~m[470]&m[471])|(m[51]&~m[468]&~m[469]&m[470]&m[471])|(~m[51]&m[468]&~m[469]&m[470]&m[471])|(~m[51]&~m[468]&m[469]&m[470]&m[471]))&~BiasedRNG[46])|((m[51]&m[468]&m[469]&m[470]&~m[471])|(m[51]&m[468]&m[469]&~m[470]&m[471])|(m[51]&m[468]&~m[469]&m[470]&m[471])|(m[51]&~m[468]&m[469]&m[470]&m[471])|(~m[51]&m[468]&m[469]&m[470]&m[471])|(m[51]&m[468]&m[469]&m[470]&m[471]))):InitCond[74];
    m[127] = run?((((m[51]&m[472]&~m[473]&~m[474]&~m[475])|(m[51]&~m[472]&m[473]&~m[474]&~m[475])|(~m[51]&m[472]&m[473]&~m[474]&~m[475])|(m[51]&~m[472]&~m[473]&m[474]&~m[475])|(~m[51]&m[472]&~m[473]&m[474]&~m[475])|(~m[51]&~m[472]&m[473]&m[474]&~m[475])|(m[51]&~m[472]&~m[473]&~m[474]&m[475])|(~m[51]&m[472]&~m[473]&~m[474]&m[475])|(~m[51]&~m[472]&m[473]&~m[474]&m[475])|(~m[51]&~m[472]&~m[473]&m[474]&m[475]))&BiasedRNG[47])|(((m[51]&m[472]&m[473]&~m[474]&~m[475])|(m[51]&m[472]&~m[473]&m[474]&~m[475])|(m[51]&~m[472]&m[473]&m[474]&~m[475])|(~m[51]&m[472]&m[473]&m[474]&~m[475])|(m[51]&m[472]&~m[473]&~m[474]&m[475])|(m[51]&~m[472]&m[473]&~m[474]&m[475])|(~m[51]&m[472]&m[473]&~m[474]&m[475])|(m[51]&~m[472]&~m[473]&m[474]&m[475])|(~m[51]&m[472]&~m[473]&m[474]&m[475])|(~m[51]&~m[472]&m[473]&m[474]&m[475]))&~BiasedRNG[47])|((m[51]&m[472]&m[473]&m[474]&~m[475])|(m[51]&m[472]&m[473]&~m[474]&m[475])|(m[51]&m[472]&~m[473]&m[474]&m[475])|(m[51]&~m[472]&m[473]&m[474]&m[475])|(~m[51]&m[472]&m[473]&m[474]&m[475])|(m[51]&m[472]&m[473]&m[474]&m[475]))):InitCond[75];
    m[129] = run?((((m[52]&m[482]&~m[483]&~m[484]&~m[485])|(m[52]&~m[482]&m[483]&~m[484]&~m[485])|(~m[52]&m[482]&m[483]&~m[484]&~m[485])|(m[52]&~m[482]&~m[483]&m[484]&~m[485])|(~m[52]&m[482]&~m[483]&m[484]&~m[485])|(~m[52]&~m[482]&m[483]&m[484]&~m[485])|(m[52]&~m[482]&~m[483]&~m[484]&m[485])|(~m[52]&m[482]&~m[483]&~m[484]&m[485])|(~m[52]&~m[482]&m[483]&~m[484]&m[485])|(~m[52]&~m[482]&~m[483]&m[484]&m[485]))&BiasedRNG[48])|(((m[52]&m[482]&m[483]&~m[484]&~m[485])|(m[52]&m[482]&~m[483]&m[484]&~m[485])|(m[52]&~m[482]&m[483]&m[484]&~m[485])|(~m[52]&m[482]&m[483]&m[484]&~m[485])|(m[52]&m[482]&~m[483]&~m[484]&m[485])|(m[52]&~m[482]&m[483]&~m[484]&m[485])|(~m[52]&m[482]&m[483]&~m[484]&m[485])|(m[52]&~m[482]&~m[483]&m[484]&m[485])|(~m[52]&m[482]&~m[483]&m[484]&m[485])|(~m[52]&~m[482]&m[483]&m[484]&m[485]))&~BiasedRNG[48])|((m[52]&m[482]&m[483]&m[484]&~m[485])|(m[52]&m[482]&m[483]&~m[484]&m[485])|(m[52]&m[482]&~m[483]&m[484]&m[485])|(m[52]&~m[482]&m[483]&m[484]&m[485])|(~m[52]&m[482]&m[483]&m[484]&m[485])|(m[52]&m[482]&m[483]&m[484]&m[485]))):InitCond[76];
    m[130] = run?((((m[52]&m[486]&~m[487]&~m[488]&~m[489])|(m[52]&~m[486]&m[487]&~m[488]&~m[489])|(~m[52]&m[486]&m[487]&~m[488]&~m[489])|(m[52]&~m[486]&~m[487]&m[488]&~m[489])|(~m[52]&m[486]&~m[487]&m[488]&~m[489])|(~m[52]&~m[486]&m[487]&m[488]&~m[489])|(m[52]&~m[486]&~m[487]&~m[488]&m[489])|(~m[52]&m[486]&~m[487]&~m[488]&m[489])|(~m[52]&~m[486]&m[487]&~m[488]&m[489])|(~m[52]&~m[486]&~m[487]&m[488]&m[489]))&BiasedRNG[49])|(((m[52]&m[486]&m[487]&~m[488]&~m[489])|(m[52]&m[486]&~m[487]&m[488]&~m[489])|(m[52]&~m[486]&m[487]&m[488]&~m[489])|(~m[52]&m[486]&m[487]&m[488]&~m[489])|(m[52]&m[486]&~m[487]&~m[488]&m[489])|(m[52]&~m[486]&m[487]&~m[488]&m[489])|(~m[52]&m[486]&m[487]&~m[488]&m[489])|(m[52]&~m[486]&~m[487]&m[488]&m[489])|(~m[52]&m[486]&~m[487]&m[488]&m[489])|(~m[52]&~m[486]&m[487]&m[488]&m[489]))&~BiasedRNG[49])|((m[52]&m[486]&m[487]&m[488]&~m[489])|(m[52]&m[486]&m[487]&~m[488]&m[489])|(m[52]&m[486]&~m[487]&m[488]&m[489])|(m[52]&~m[486]&m[487]&m[488]&m[489])|(~m[52]&m[486]&m[487]&m[488]&m[489])|(m[52]&m[486]&m[487]&m[488]&m[489]))):InitCond[77];
    m[132] = run?((((m[53]&m[496]&~m[497]&~m[498]&~m[499])|(m[53]&~m[496]&m[497]&~m[498]&~m[499])|(~m[53]&m[496]&m[497]&~m[498]&~m[499])|(m[53]&~m[496]&~m[497]&m[498]&~m[499])|(~m[53]&m[496]&~m[497]&m[498]&~m[499])|(~m[53]&~m[496]&m[497]&m[498]&~m[499])|(m[53]&~m[496]&~m[497]&~m[498]&m[499])|(~m[53]&m[496]&~m[497]&~m[498]&m[499])|(~m[53]&~m[496]&m[497]&~m[498]&m[499])|(~m[53]&~m[496]&~m[497]&m[498]&m[499]))&BiasedRNG[50])|(((m[53]&m[496]&m[497]&~m[498]&~m[499])|(m[53]&m[496]&~m[497]&m[498]&~m[499])|(m[53]&~m[496]&m[497]&m[498]&~m[499])|(~m[53]&m[496]&m[497]&m[498]&~m[499])|(m[53]&m[496]&~m[497]&~m[498]&m[499])|(m[53]&~m[496]&m[497]&~m[498]&m[499])|(~m[53]&m[496]&m[497]&~m[498]&m[499])|(m[53]&~m[496]&~m[497]&m[498]&m[499])|(~m[53]&m[496]&~m[497]&m[498]&m[499])|(~m[53]&~m[496]&m[497]&m[498]&m[499]))&~BiasedRNG[50])|((m[53]&m[496]&m[497]&m[498]&~m[499])|(m[53]&m[496]&m[497]&~m[498]&m[499])|(m[53]&m[496]&~m[497]&m[498]&m[499])|(m[53]&~m[496]&m[497]&m[498]&m[499])|(~m[53]&m[496]&m[497]&m[498]&m[499])|(m[53]&m[496]&m[497]&m[498]&m[499]))):InitCond[78];
    m[133] = run?((((m[53]&m[500]&~m[501]&~m[502]&~m[503])|(m[53]&~m[500]&m[501]&~m[502]&~m[503])|(~m[53]&m[500]&m[501]&~m[502]&~m[503])|(m[53]&~m[500]&~m[501]&m[502]&~m[503])|(~m[53]&m[500]&~m[501]&m[502]&~m[503])|(~m[53]&~m[500]&m[501]&m[502]&~m[503])|(m[53]&~m[500]&~m[501]&~m[502]&m[503])|(~m[53]&m[500]&~m[501]&~m[502]&m[503])|(~m[53]&~m[500]&m[501]&~m[502]&m[503])|(~m[53]&~m[500]&~m[501]&m[502]&m[503]))&BiasedRNG[51])|(((m[53]&m[500]&m[501]&~m[502]&~m[503])|(m[53]&m[500]&~m[501]&m[502]&~m[503])|(m[53]&~m[500]&m[501]&m[502]&~m[503])|(~m[53]&m[500]&m[501]&m[502]&~m[503])|(m[53]&m[500]&~m[501]&~m[502]&m[503])|(m[53]&~m[500]&m[501]&~m[502]&m[503])|(~m[53]&m[500]&m[501]&~m[502]&m[503])|(m[53]&~m[500]&~m[501]&m[502]&m[503])|(~m[53]&m[500]&~m[501]&m[502]&m[503])|(~m[53]&~m[500]&m[501]&m[502]&m[503]))&~BiasedRNG[51])|((m[53]&m[500]&m[501]&m[502]&~m[503])|(m[53]&m[500]&m[501]&~m[502]&m[503])|(m[53]&m[500]&~m[501]&m[502]&m[503])|(m[53]&~m[500]&m[501]&m[502]&m[503])|(~m[53]&m[500]&m[501]&m[502]&m[503])|(m[53]&m[500]&m[501]&m[502]&m[503]))):InitCond[79];
    m[135] = run?((((m[54]&m[510]&~m[511]&~m[512]&~m[513])|(m[54]&~m[510]&m[511]&~m[512]&~m[513])|(~m[54]&m[510]&m[511]&~m[512]&~m[513])|(m[54]&~m[510]&~m[511]&m[512]&~m[513])|(~m[54]&m[510]&~m[511]&m[512]&~m[513])|(~m[54]&~m[510]&m[511]&m[512]&~m[513])|(m[54]&~m[510]&~m[511]&~m[512]&m[513])|(~m[54]&m[510]&~m[511]&~m[512]&m[513])|(~m[54]&~m[510]&m[511]&~m[512]&m[513])|(~m[54]&~m[510]&~m[511]&m[512]&m[513]))&BiasedRNG[52])|(((m[54]&m[510]&m[511]&~m[512]&~m[513])|(m[54]&m[510]&~m[511]&m[512]&~m[513])|(m[54]&~m[510]&m[511]&m[512]&~m[513])|(~m[54]&m[510]&m[511]&m[512]&~m[513])|(m[54]&m[510]&~m[511]&~m[512]&m[513])|(m[54]&~m[510]&m[511]&~m[512]&m[513])|(~m[54]&m[510]&m[511]&~m[512]&m[513])|(m[54]&~m[510]&~m[511]&m[512]&m[513])|(~m[54]&m[510]&~m[511]&m[512]&m[513])|(~m[54]&~m[510]&m[511]&m[512]&m[513]))&~BiasedRNG[52])|((m[54]&m[510]&m[511]&m[512]&~m[513])|(m[54]&m[510]&m[511]&~m[512]&m[513])|(m[54]&m[510]&~m[511]&m[512]&m[513])|(m[54]&~m[510]&m[511]&m[512]&m[513])|(~m[54]&m[510]&m[511]&m[512]&m[513])|(m[54]&m[510]&m[511]&m[512]&m[513]))):InitCond[80];
    m[136] = run?((((m[54]&m[514]&~m[515]&~m[516]&~m[517])|(m[54]&~m[514]&m[515]&~m[516]&~m[517])|(~m[54]&m[514]&m[515]&~m[516]&~m[517])|(m[54]&~m[514]&~m[515]&m[516]&~m[517])|(~m[54]&m[514]&~m[515]&m[516]&~m[517])|(~m[54]&~m[514]&m[515]&m[516]&~m[517])|(m[54]&~m[514]&~m[515]&~m[516]&m[517])|(~m[54]&m[514]&~m[515]&~m[516]&m[517])|(~m[54]&~m[514]&m[515]&~m[516]&m[517])|(~m[54]&~m[514]&~m[515]&m[516]&m[517]))&BiasedRNG[53])|(((m[54]&m[514]&m[515]&~m[516]&~m[517])|(m[54]&m[514]&~m[515]&m[516]&~m[517])|(m[54]&~m[514]&m[515]&m[516]&~m[517])|(~m[54]&m[514]&m[515]&m[516]&~m[517])|(m[54]&m[514]&~m[515]&~m[516]&m[517])|(m[54]&~m[514]&m[515]&~m[516]&m[517])|(~m[54]&m[514]&m[515]&~m[516]&m[517])|(m[54]&~m[514]&~m[515]&m[516]&m[517])|(~m[54]&m[514]&~m[515]&m[516]&m[517])|(~m[54]&~m[514]&m[515]&m[516]&m[517]))&~BiasedRNG[53])|((m[54]&m[514]&m[515]&m[516]&~m[517])|(m[54]&m[514]&m[515]&~m[516]&m[517])|(m[54]&m[514]&~m[515]&m[516]&m[517])|(m[54]&~m[514]&m[515]&m[516]&m[517])|(~m[54]&m[514]&m[515]&m[516]&m[517])|(m[54]&m[514]&m[515]&m[516]&m[517]))):InitCond[81];
    m[138] = run?((((m[55]&m[524]&~m[525]&~m[526]&~m[527])|(m[55]&~m[524]&m[525]&~m[526]&~m[527])|(~m[55]&m[524]&m[525]&~m[526]&~m[527])|(m[55]&~m[524]&~m[525]&m[526]&~m[527])|(~m[55]&m[524]&~m[525]&m[526]&~m[527])|(~m[55]&~m[524]&m[525]&m[526]&~m[527])|(m[55]&~m[524]&~m[525]&~m[526]&m[527])|(~m[55]&m[524]&~m[525]&~m[526]&m[527])|(~m[55]&~m[524]&m[525]&~m[526]&m[527])|(~m[55]&~m[524]&~m[525]&m[526]&m[527]))&BiasedRNG[54])|(((m[55]&m[524]&m[525]&~m[526]&~m[527])|(m[55]&m[524]&~m[525]&m[526]&~m[527])|(m[55]&~m[524]&m[525]&m[526]&~m[527])|(~m[55]&m[524]&m[525]&m[526]&~m[527])|(m[55]&m[524]&~m[525]&~m[526]&m[527])|(m[55]&~m[524]&m[525]&~m[526]&m[527])|(~m[55]&m[524]&m[525]&~m[526]&m[527])|(m[55]&~m[524]&~m[525]&m[526]&m[527])|(~m[55]&m[524]&~m[525]&m[526]&m[527])|(~m[55]&~m[524]&m[525]&m[526]&m[527]))&~BiasedRNG[54])|((m[55]&m[524]&m[525]&m[526]&~m[527])|(m[55]&m[524]&m[525]&~m[526]&m[527])|(m[55]&m[524]&~m[525]&m[526]&m[527])|(m[55]&~m[524]&m[525]&m[526]&m[527])|(~m[55]&m[524]&m[525]&m[526]&m[527])|(m[55]&m[524]&m[525]&m[526]&m[527]))):InitCond[82];
    m[139] = run?((((m[55]&m[528]&~m[529]&~m[530]&~m[531])|(m[55]&~m[528]&m[529]&~m[530]&~m[531])|(~m[55]&m[528]&m[529]&~m[530]&~m[531])|(m[55]&~m[528]&~m[529]&m[530]&~m[531])|(~m[55]&m[528]&~m[529]&m[530]&~m[531])|(~m[55]&~m[528]&m[529]&m[530]&~m[531])|(m[55]&~m[528]&~m[529]&~m[530]&m[531])|(~m[55]&m[528]&~m[529]&~m[530]&m[531])|(~m[55]&~m[528]&m[529]&~m[530]&m[531])|(~m[55]&~m[528]&~m[529]&m[530]&m[531]))&BiasedRNG[55])|(((m[55]&m[528]&m[529]&~m[530]&~m[531])|(m[55]&m[528]&~m[529]&m[530]&~m[531])|(m[55]&~m[528]&m[529]&m[530]&~m[531])|(~m[55]&m[528]&m[529]&m[530]&~m[531])|(m[55]&m[528]&~m[529]&~m[530]&m[531])|(m[55]&~m[528]&m[529]&~m[530]&m[531])|(~m[55]&m[528]&m[529]&~m[530]&m[531])|(m[55]&~m[528]&~m[529]&m[530]&m[531])|(~m[55]&m[528]&~m[529]&m[530]&m[531])|(~m[55]&~m[528]&m[529]&m[530]&m[531]))&~BiasedRNG[55])|((m[55]&m[528]&m[529]&m[530]&~m[531])|(m[55]&m[528]&m[529]&~m[530]&m[531])|(m[55]&m[528]&~m[529]&m[530]&m[531])|(m[55]&~m[528]&m[529]&m[530]&m[531])|(~m[55]&m[528]&m[529]&m[530]&m[531])|(m[55]&m[528]&m[529]&m[530]&m[531]))):InitCond[83];
    m[140] = run?((((~m[28]&~m[336]&~m[532])|(m[28]&m[336]&~m[532]))&BiasedRNG[56])|(((m[28]&~m[336]&~m[532])|(~m[28]&m[336]&m[532]))&~BiasedRNG[56])|((~m[28]&~m[336]&m[532])|(m[28]&~m[336]&m[532])|(m[28]&m[336]&m[532]))):InitCond[84];
    m[141] = run?((((~m[28]&~m[350]&~m[546])|(m[28]&m[350]&~m[546]))&BiasedRNG[57])|(((m[28]&~m[350]&~m[546])|(~m[28]&m[350]&m[546]))&~BiasedRNG[57])|((~m[28]&~m[350]&m[546])|(m[28]&~m[350]&m[546])|(m[28]&m[350]&m[546]))):InitCond[85];
    m[142] = run?((((~m[56]&~m[364]&~m[560])|(m[56]&m[364]&~m[560]))&BiasedRNG[58])|(((m[56]&~m[364]&~m[560])|(~m[56]&m[364]&m[560]))&~BiasedRNG[58])|((~m[56]&~m[364]&m[560])|(m[56]&~m[364]&m[560])|(m[56]&m[364]&m[560]))):InitCond[86];
    m[143] = run?((((~m[56]&~m[378]&~m[574])|(m[56]&m[378]&~m[574]))&BiasedRNG[59])|(((m[56]&~m[378]&~m[574])|(~m[56]&m[378]&m[574]))&~BiasedRNG[59])|((~m[56]&~m[378]&m[574])|(m[56]&~m[378]&m[574])|(m[56]&m[378]&m[574]))):InitCond[87];
    m[144] = run?((((~m[56]&~m[392]&~m[588])|(m[56]&m[392]&~m[588]))&BiasedRNG[60])|(((m[56]&~m[392]&~m[588])|(~m[56]&m[392]&m[588]))&~BiasedRNG[60])|((~m[56]&~m[392]&m[588])|(m[56]&~m[392]&m[588])|(m[56]&m[392]&m[588]))):InitCond[88];
    m[145] = run?((((~m[56]&~m[406]&~m[602])|(m[56]&m[406]&~m[602]))&BiasedRNG[61])|(((m[56]&~m[406]&~m[602])|(~m[56]&m[406]&m[602]))&~BiasedRNG[61])|((~m[56]&~m[406]&m[602])|(m[56]&~m[406]&m[602])|(m[56]&m[406]&m[602]))):InitCond[89];
    m[154] = run?((((~m[29]&~m[337]&~m[533])|(m[29]&m[337]&~m[533]))&BiasedRNG[62])|(((m[29]&~m[337]&~m[533])|(~m[29]&m[337]&m[533]))&~BiasedRNG[62])|((~m[29]&~m[337]&m[533])|(m[29]&~m[337]&m[533])|(m[29]&m[337]&m[533]))):InitCond[90];
    m[155] = run?((((~m[29]&~m[351]&~m[547])|(m[29]&m[351]&~m[547]))&BiasedRNG[63])|(((m[29]&~m[351]&~m[547])|(~m[29]&m[351]&m[547]))&~BiasedRNG[63])|((~m[29]&~m[351]&m[547])|(m[29]&~m[351]&m[547])|(m[29]&m[351]&m[547]))):InitCond[91];
    m[156] = run?((((~m[59]&~m[365]&~m[561])|(m[59]&m[365]&~m[561]))&BiasedRNG[64])|(((m[59]&~m[365]&~m[561])|(~m[59]&m[365]&m[561]))&~BiasedRNG[64])|((~m[59]&~m[365]&m[561])|(m[59]&~m[365]&m[561])|(m[59]&m[365]&m[561]))):InitCond[92];
    m[157] = run?((((~m[59]&~m[379]&~m[575])|(m[59]&m[379]&~m[575]))&BiasedRNG[65])|(((m[59]&~m[379]&~m[575])|(~m[59]&m[379]&m[575]))&~BiasedRNG[65])|((~m[59]&~m[379]&m[575])|(m[59]&~m[379]&m[575])|(m[59]&m[379]&m[575]))):InitCond[93];
    m[158] = run?((((~m[59]&~m[393]&~m[589])|(m[59]&m[393]&~m[589]))&BiasedRNG[66])|(((m[59]&~m[393]&~m[589])|(~m[59]&m[393]&m[589]))&~BiasedRNG[66])|((~m[59]&~m[393]&m[589])|(m[59]&~m[393]&m[589])|(m[59]&m[393]&m[589]))):InitCond[94];
    m[159] = run?((((~m[59]&~m[407]&~m[603])|(m[59]&m[407]&~m[603]))&BiasedRNG[67])|(((m[59]&~m[407]&~m[603])|(~m[59]&m[407]&m[603]))&~BiasedRNG[67])|((~m[59]&~m[407]&m[603])|(m[59]&~m[407]&m[603])|(m[59]&m[407]&m[603]))):InitCond[95];
    m[168] = run?((((~m[30]&~m[338]&~m[534])|(m[30]&m[338]&~m[534]))&BiasedRNG[68])|(((m[30]&~m[338]&~m[534])|(~m[30]&m[338]&m[534]))&~BiasedRNG[68])|((~m[30]&~m[338]&m[534])|(m[30]&~m[338]&m[534])|(m[30]&m[338]&m[534]))):InitCond[96];
    m[169] = run?((((~m[30]&~m[352]&~m[548])|(m[30]&m[352]&~m[548]))&BiasedRNG[69])|(((m[30]&~m[352]&~m[548])|(~m[30]&m[352]&m[548]))&~BiasedRNG[69])|((~m[30]&~m[352]&m[548])|(m[30]&~m[352]&m[548])|(m[30]&m[352]&m[548]))):InitCond[97];
    m[170] = run?((((~m[62]&~m[366]&~m[562])|(m[62]&m[366]&~m[562]))&BiasedRNG[70])|(((m[62]&~m[366]&~m[562])|(~m[62]&m[366]&m[562]))&~BiasedRNG[70])|((~m[62]&~m[366]&m[562])|(m[62]&~m[366]&m[562])|(m[62]&m[366]&m[562]))):InitCond[98];
    m[171] = run?((((~m[62]&~m[380]&~m[576])|(m[62]&m[380]&~m[576]))&BiasedRNG[71])|(((m[62]&~m[380]&~m[576])|(~m[62]&m[380]&m[576]))&~BiasedRNG[71])|((~m[62]&~m[380]&m[576])|(m[62]&~m[380]&m[576])|(m[62]&m[380]&m[576]))):InitCond[99];
    m[172] = run?((((~m[62]&~m[394]&~m[590])|(m[62]&m[394]&~m[590]))&BiasedRNG[72])|(((m[62]&~m[394]&~m[590])|(~m[62]&m[394]&m[590]))&~BiasedRNG[72])|((~m[62]&~m[394]&m[590])|(m[62]&~m[394]&m[590])|(m[62]&m[394]&m[590]))):InitCond[100];
    m[173] = run?((((~m[62]&~m[408]&~m[604])|(m[62]&m[408]&~m[604]))&BiasedRNG[73])|(((m[62]&~m[408]&~m[604])|(~m[62]&m[408]&m[604]))&~BiasedRNG[73])|((~m[62]&~m[408]&m[604])|(m[62]&~m[408]&m[604])|(m[62]&m[408]&m[604]))):InitCond[101];
    m[182] = run?((((~m[31]&~m[339]&~m[535])|(m[31]&m[339]&~m[535]))&BiasedRNG[74])|(((m[31]&~m[339]&~m[535])|(~m[31]&m[339]&m[535]))&~BiasedRNG[74])|((~m[31]&~m[339]&m[535])|(m[31]&~m[339]&m[535])|(m[31]&m[339]&m[535]))):InitCond[102];
    m[183] = run?((((~m[31]&~m[353]&~m[549])|(m[31]&m[353]&~m[549]))&BiasedRNG[75])|(((m[31]&~m[353]&~m[549])|(~m[31]&m[353]&m[549]))&~BiasedRNG[75])|((~m[31]&~m[353]&m[549])|(m[31]&~m[353]&m[549])|(m[31]&m[353]&m[549]))):InitCond[103];
    m[184] = run?((((~m[65]&~m[367]&~m[563])|(m[65]&m[367]&~m[563]))&BiasedRNG[76])|(((m[65]&~m[367]&~m[563])|(~m[65]&m[367]&m[563]))&~BiasedRNG[76])|((~m[65]&~m[367]&m[563])|(m[65]&~m[367]&m[563])|(m[65]&m[367]&m[563]))):InitCond[104];
    m[185] = run?((((~m[65]&~m[381]&~m[577])|(m[65]&m[381]&~m[577]))&BiasedRNG[77])|(((m[65]&~m[381]&~m[577])|(~m[65]&m[381]&m[577]))&~BiasedRNG[77])|((~m[65]&~m[381]&m[577])|(m[65]&~m[381]&m[577])|(m[65]&m[381]&m[577]))):InitCond[105];
    m[186] = run?((((~m[65]&~m[395]&~m[591])|(m[65]&m[395]&~m[591]))&BiasedRNG[78])|(((m[65]&~m[395]&~m[591])|(~m[65]&m[395]&m[591]))&~BiasedRNG[78])|((~m[65]&~m[395]&m[591])|(m[65]&~m[395]&m[591])|(m[65]&m[395]&m[591]))):InitCond[106];
    m[187] = run?((((~m[65]&~m[409]&~m[605])|(m[65]&m[409]&~m[605]))&BiasedRNG[79])|(((m[65]&~m[409]&~m[605])|(~m[65]&m[409]&m[605]))&~BiasedRNG[79])|((~m[65]&~m[409]&m[605])|(m[65]&~m[409]&m[605])|(m[65]&m[409]&m[605]))):InitCond[107];
    m[196] = run?((((~m[32]&~m[340]&~m[536])|(m[32]&m[340]&~m[536]))&BiasedRNG[80])|(((m[32]&~m[340]&~m[536])|(~m[32]&m[340]&m[536]))&~BiasedRNG[80])|((~m[32]&~m[340]&m[536])|(m[32]&~m[340]&m[536])|(m[32]&m[340]&m[536]))):InitCond[108];
    m[197] = run?((((~m[32]&~m[354]&~m[550])|(m[32]&m[354]&~m[550]))&BiasedRNG[81])|(((m[32]&~m[354]&~m[550])|(~m[32]&m[354]&m[550]))&~BiasedRNG[81])|((~m[32]&~m[354]&m[550])|(m[32]&~m[354]&m[550])|(m[32]&m[354]&m[550]))):InitCond[109];
    m[198] = run?((((~m[68]&~m[368]&~m[564])|(m[68]&m[368]&~m[564]))&BiasedRNG[82])|(((m[68]&~m[368]&~m[564])|(~m[68]&m[368]&m[564]))&~BiasedRNG[82])|((~m[68]&~m[368]&m[564])|(m[68]&~m[368]&m[564])|(m[68]&m[368]&m[564]))):InitCond[110];
    m[199] = run?((((~m[68]&~m[382]&~m[578])|(m[68]&m[382]&~m[578]))&BiasedRNG[83])|(((m[68]&~m[382]&~m[578])|(~m[68]&m[382]&m[578]))&~BiasedRNG[83])|((~m[68]&~m[382]&m[578])|(m[68]&~m[382]&m[578])|(m[68]&m[382]&m[578]))):InitCond[111];
    m[200] = run?((((~m[68]&~m[396]&~m[592])|(m[68]&m[396]&~m[592]))&BiasedRNG[84])|(((m[68]&~m[396]&~m[592])|(~m[68]&m[396]&m[592]))&~BiasedRNG[84])|((~m[68]&~m[396]&m[592])|(m[68]&~m[396]&m[592])|(m[68]&m[396]&m[592]))):InitCond[112];
    m[201] = run?((((~m[68]&~m[410]&~m[606])|(m[68]&m[410]&~m[606]))&BiasedRNG[85])|(((m[68]&~m[410]&~m[606])|(~m[68]&m[410]&m[606]))&~BiasedRNG[85])|((~m[68]&~m[410]&m[606])|(m[68]&~m[410]&m[606])|(m[68]&m[410]&m[606]))):InitCond[113];
    m[210] = run?((((~m[33]&~m[341]&~m[537])|(m[33]&m[341]&~m[537]))&BiasedRNG[86])|(((m[33]&~m[341]&~m[537])|(~m[33]&m[341]&m[537]))&~BiasedRNG[86])|((~m[33]&~m[341]&m[537])|(m[33]&~m[341]&m[537])|(m[33]&m[341]&m[537]))):InitCond[114];
    m[211] = run?((((~m[33]&~m[355]&~m[551])|(m[33]&m[355]&~m[551]))&BiasedRNG[87])|(((m[33]&~m[355]&~m[551])|(~m[33]&m[355]&m[551]))&~BiasedRNG[87])|((~m[33]&~m[355]&m[551])|(m[33]&~m[355]&m[551])|(m[33]&m[355]&m[551]))):InitCond[115];
    m[212] = run?((((~m[71]&~m[369]&~m[565])|(m[71]&m[369]&~m[565]))&BiasedRNG[88])|(((m[71]&~m[369]&~m[565])|(~m[71]&m[369]&m[565]))&~BiasedRNG[88])|((~m[71]&~m[369]&m[565])|(m[71]&~m[369]&m[565])|(m[71]&m[369]&m[565]))):InitCond[116];
    m[213] = run?((((~m[71]&~m[383]&~m[579])|(m[71]&m[383]&~m[579]))&BiasedRNG[89])|(((m[71]&~m[383]&~m[579])|(~m[71]&m[383]&m[579]))&~BiasedRNG[89])|((~m[71]&~m[383]&m[579])|(m[71]&~m[383]&m[579])|(m[71]&m[383]&m[579]))):InitCond[117];
    m[214] = run?((((~m[71]&~m[397]&~m[593])|(m[71]&m[397]&~m[593]))&BiasedRNG[90])|(((m[71]&~m[397]&~m[593])|(~m[71]&m[397]&m[593]))&~BiasedRNG[90])|((~m[71]&~m[397]&m[593])|(m[71]&~m[397]&m[593])|(m[71]&m[397]&m[593]))):InitCond[118];
    m[215] = run?((((~m[71]&~m[411]&~m[607])|(m[71]&m[411]&~m[607]))&BiasedRNG[91])|(((m[71]&~m[411]&~m[607])|(~m[71]&m[411]&m[607]))&~BiasedRNG[91])|((~m[71]&~m[411]&m[607])|(m[71]&~m[411]&m[607])|(m[71]&m[411]&m[607]))):InitCond[119];
    m[224] = run?((((~m[34]&~m[342]&~m[538])|(m[34]&m[342]&~m[538]))&BiasedRNG[92])|(((m[34]&~m[342]&~m[538])|(~m[34]&m[342]&m[538]))&~BiasedRNG[92])|((~m[34]&~m[342]&m[538])|(m[34]&~m[342]&m[538])|(m[34]&m[342]&m[538]))):InitCond[120];
    m[225] = run?((((~m[34]&~m[356]&~m[552])|(m[34]&m[356]&~m[552]))&BiasedRNG[93])|(((m[34]&~m[356]&~m[552])|(~m[34]&m[356]&m[552]))&~BiasedRNG[93])|((~m[34]&~m[356]&m[552])|(m[34]&~m[356]&m[552])|(m[34]&m[356]&m[552]))):InitCond[121];
    m[226] = run?((((~m[74]&~m[370]&~m[566])|(m[74]&m[370]&~m[566]))&BiasedRNG[94])|(((m[74]&~m[370]&~m[566])|(~m[74]&m[370]&m[566]))&~BiasedRNG[94])|((~m[74]&~m[370]&m[566])|(m[74]&~m[370]&m[566])|(m[74]&m[370]&m[566]))):InitCond[122];
    m[227] = run?((((~m[74]&~m[384]&~m[580])|(m[74]&m[384]&~m[580]))&BiasedRNG[95])|(((m[74]&~m[384]&~m[580])|(~m[74]&m[384]&m[580]))&~BiasedRNG[95])|((~m[74]&~m[384]&m[580])|(m[74]&~m[384]&m[580])|(m[74]&m[384]&m[580]))):InitCond[123];
    m[228] = run?((((~m[74]&~m[398]&~m[594])|(m[74]&m[398]&~m[594]))&BiasedRNG[96])|(((m[74]&~m[398]&~m[594])|(~m[74]&m[398]&m[594]))&~BiasedRNG[96])|((~m[74]&~m[398]&m[594])|(m[74]&~m[398]&m[594])|(m[74]&m[398]&m[594]))):InitCond[124];
    m[229] = run?((((~m[74]&~m[412]&~m[608])|(m[74]&m[412]&~m[608]))&BiasedRNG[97])|(((m[74]&~m[412]&~m[608])|(~m[74]&m[412]&m[608]))&~BiasedRNG[97])|((~m[74]&~m[412]&m[608])|(m[74]&~m[412]&m[608])|(m[74]&m[412]&m[608]))):InitCond[125];
    m[238] = run?((((~m[35]&~m[343]&~m[539])|(m[35]&m[343]&~m[539]))&BiasedRNG[98])|(((m[35]&~m[343]&~m[539])|(~m[35]&m[343]&m[539]))&~BiasedRNG[98])|((~m[35]&~m[343]&m[539])|(m[35]&~m[343]&m[539])|(m[35]&m[343]&m[539]))):InitCond[126];
    m[239] = run?((((~m[35]&~m[357]&~m[553])|(m[35]&m[357]&~m[553]))&BiasedRNG[99])|(((m[35]&~m[357]&~m[553])|(~m[35]&m[357]&m[553]))&~BiasedRNG[99])|((~m[35]&~m[357]&m[553])|(m[35]&~m[357]&m[553])|(m[35]&m[357]&m[553]))):InitCond[127];
    m[240] = run?((((~m[77]&~m[371]&~m[567])|(m[77]&m[371]&~m[567]))&BiasedRNG[100])|(((m[77]&~m[371]&~m[567])|(~m[77]&m[371]&m[567]))&~BiasedRNG[100])|((~m[77]&~m[371]&m[567])|(m[77]&~m[371]&m[567])|(m[77]&m[371]&m[567]))):InitCond[128];
    m[241] = run?((((~m[77]&~m[385]&~m[581])|(m[77]&m[385]&~m[581]))&BiasedRNG[101])|(((m[77]&~m[385]&~m[581])|(~m[77]&m[385]&m[581]))&~BiasedRNG[101])|((~m[77]&~m[385]&m[581])|(m[77]&~m[385]&m[581])|(m[77]&m[385]&m[581]))):InitCond[129];
    m[242] = run?((((~m[77]&~m[399]&~m[595])|(m[77]&m[399]&~m[595]))&BiasedRNG[102])|(((m[77]&~m[399]&~m[595])|(~m[77]&m[399]&m[595]))&~BiasedRNG[102])|((~m[77]&~m[399]&m[595])|(m[77]&~m[399]&m[595])|(m[77]&m[399]&m[595]))):InitCond[130];
    m[243] = run?((((~m[77]&~m[413]&~m[609])|(m[77]&m[413]&~m[609]))&BiasedRNG[103])|(((m[77]&~m[413]&~m[609])|(~m[77]&m[413]&m[609]))&~BiasedRNG[103])|((~m[77]&~m[413]&m[609])|(m[77]&~m[413]&m[609])|(m[77]&m[413]&m[609]))):InitCond[131];
    m[252] = run?((((~m[36]&~m[344]&~m[540])|(m[36]&m[344]&~m[540]))&BiasedRNG[104])|(((m[36]&~m[344]&~m[540])|(~m[36]&m[344]&m[540]))&~BiasedRNG[104])|((~m[36]&~m[344]&m[540])|(m[36]&~m[344]&m[540])|(m[36]&m[344]&m[540]))):InitCond[132];
    m[253] = run?((((~m[36]&~m[358]&~m[554])|(m[36]&m[358]&~m[554]))&BiasedRNG[105])|(((m[36]&~m[358]&~m[554])|(~m[36]&m[358]&m[554]))&~BiasedRNG[105])|((~m[36]&~m[358]&m[554])|(m[36]&~m[358]&m[554])|(m[36]&m[358]&m[554]))):InitCond[133];
    m[254] = run?((((~m[80]&~m[372]&~m[568])|(m[80]&m[372]&~m[568]))&BiasedRNG[106])|(((m[80]&~m[372]&~m[568])|(~m[80]&m[372]&m[568]))&~BiasedRNG[106])|((~m[80]&~m[372]&m[568])|(m[80]&~m[372]&m[568])|(m[80]&m[372]&m[568]))):InitCond[134];
    m[255] = run?((((~m[80]&~m[386]&~m[582])|(m[80]&m[386]&~m[582]))&BiasedRNG[107])|(((m[80]&~m[386]&~m[582])|(~m[80]&m[386]&m[582]))&~BiasedRNG[107])|((~m[80]&~m[386]&m[582])|(m[80]&~m[386]&m[582])|(m[80]&m[386]&m[582]))):InitCond[135];
    m[256] = run?((((~m[80]&~m[400]&~m[596])|(m[80]&m[400]&~m[596]))&BiasedRNG[108])|(((m[80]&~m[400]&~m[596])|(~m[80]&m[400]&m[596]))&~BiasedRNG[108])|((~m[80]&~m[400]&m[596])|(m[80]&~m[400]&m[596])|(m[80]&m[400]&m[596]))):InitCond[136];
    m[257] = run?((((~m[80]&~m[414]&~m[610])|(m[80]&m[414]&~m[610]))&BiasedRNG[109])|(((m[80]&~m[414]&~m[610])|(~m[80]&m[414]&m[610]))&~BiasedRNG[109])|((~m[80]&~m[414]&m[610])|(m[80]&~m[414]&m[610])|(m[80]&m[414]&m[610]))):InitCond[137];
    m[266] = run?((((~m[37]&~m[345]&~m[541])|(m[37]&m[345]&~m[541]))&BiasedRNG[110])|(((m[37]&~m[345]&~m[541])|(~m[37]&m[345]&m[541]))&~BiasedRNG[110])|((~m[37]&~m[345]&m[541])|(m[37]&~m[345]&m[541])|(m[37]&m[345]&m[541]))):InitCond[138];
    m[267] = run?((((~m[37]&~m[359]&~m[555])|(m[37]&m[359]&~m[555]))&BiasedRNG[111])|(((m[37]&~m[359]&~m[555])|(~m[37]&m[359]&m[555]))&~BiasedRNG[111])|((~m[37]&~m[359]&m[555])|(m[37]&~m[359]&m[555])|(m[37]&m[359]&m[555]))):InitCond[139];
    m[268] = run?((((~m[83]&~m[373]&~m[569])|(m[83]&m[373]&~m[569]))&BiasedRNG[112])|(((m[83]&~m[373]&~m[569])|(~m[83]&m[373]&m[569]))&~BiasedRNG[112])|((~m[83]&~m[373]&m[569])|(m[83]&~m[373]&m[569])|(m[83]&m[373]&m[569]))):InitCond[140];
    m[269] = run?((((~m[83]&~m[387]&~m[583])|(m[83]&m[387]&~m[583]))&BiasedRNG[113])|(((m[83]&~m[387]&~m[583])|(~m[83]&m[387]&m[583]))&~BiasedRNG[113])|((~m[83]&~m[387]&m[583])|(m[83]&~m[387]&m[583])|(m[83]&m[387]&m[583]))):InitCond[141];
    m[270] = run?((((~m[83]&~m[401]&~m[597])|(m[83]&m[401]&~m[597]))&BiasedRNG[114])|(((m[83]&~m[401]&~m[597])|(~m[83]&m[401]&m[597]))&~BiasedRNG[114])|((~m[83]&~m[401]&m[597])|(m[83]&~m[401]&m[597])|(m[83]&m[401]&m[597]))):InitCond[142];
    m[271] = run?((((~m[83]&~m[415]&~m[611])|(m[83]&m[415]&~m[611]))&BiasedRNG[115])|(((m[83]&~m[415]&~m[611])|(~m[83]&m[415]&m[611]))&~BiasedRNG[115])|((~m[83]&~m[415]&m[611])|(m[83]&~m[415]&m[611])|(m[83]&m[415]&m[611]))):InitCond[143];
    m[280] = run?((((~m[38]&~m[346]&~m[542])|(m[38]&m[346]&~m[542]))&BiasedRNG[116])|(((m[38]&~m[346]&~m[542])|(~m[38]&m[346]&m[542]))&~BiasedRNG[116])|((~m[38]&~m[346]&m[542])|(m[38]&~m[346]&m[542])|(m[38]&m[346]&m[542]))):InitCond[144];
    m[281] = run?((((~m[38]&~m[360]&~m[556])|(m[38]&m[360]&~m[556]))&BiasedRNG[117])|(((m[38]&~m[360]&~m[556])|(~m[38]&m[360]&m[556]))&~BiasedRNG[117])|((~m[38]&~m[360]&m[556])|(m[38]&~m[360]&m[556])|(m[38]&m[360]&m[556]))):InitCond[145];
    m[282] = run?((((~m[86]&~m[374]&~m[570])|(m[86]&m[374]&~m[570]))&BiasedRNG[118])|(((m[86]&~m[374]&~m[570])|(~m[86]&m[374]&m[570]))&~BiasedRNG[118])|((~m[86]&~m[374]&m[570])|(m[86]&~m[374]&m[570])|(m[86]&m[374]&m[570]))):InitCond[146];
    m[283] = run?((((~m[86]&~m[388]&~m[584])|(m[86]&m[388]&~m[584]))&BiasedRNG[119])|(((m[86]&~m[388]&~m[584])|(~m[86]&m[388]&m[584]))&~BiasedRNG[119])|((~m[86]&~m[388]&m[584])|(m[86]&~m[388]&m[584])|(m[86]&m[388]&m[584]))):InitCond[147];
    m[284] = run?((((~m[86]&~m[402]&~m[598])|(m[86]&m[402]&~m[598]))&BiasedRNG[120])|(((m[86]&~m[402]&~m[598])|(~m[86]&m[402]&m[598]))&~BiasedRNG[120])|((~m[86]&~m[402]&m[598])|(m[86]&~m[402]&m[598])|(m[86]&m[402]&m[598]))):InitCond[148];
    m[285] = run?((((~m[86]&~m[416]&~m[612])|(m[86]&m[416]&~m[612]))&BiasedRNG[121])|(((m[86]&~m[416]&~m[612])|(~m[86]&m[416]&m[612]))&~BiasedRNG[121])|((~m[86]&~m[416]&m[612])|(m[86]&~m[416]&m[612])|(m[86]&m[416]&m[612]))):InitCond[149];
    m[294] = run?((((~m[39]&~m[347]&~m[543])|(m[39]&m[347]&~m[543]))&BiasedRNG[122])|(((m[39]&~m[347]&~m[543])|(~m[39]&m[347]&m[543]))&~BiasedRNG[122])|((~m[39]&~m[347]&m[543])|(m[39]&~m[347]&m[543])|(m[39]&m[347]&m[543]))):InitCond[150];
    m[295] = run?((((~m[39]&~m[361]&~m[557])|(m[39]&m[361]&~m[557]))&BiasedRNG[123])|(((m[39]&~m[361]&~m[557])|(~m[39]&m[361]&m[557]))&~BiasedRNG[123])|((~m[39]&~m[361]&m[557])|(m[39]&~m[361]&m[557])|(m[39]&m[361]&m[557]))):InitCond[151];
    m[296] = run?((((~m[89]&~m[375]&~m[571])|(m[89]&m[375]&~m[571]))&BiasedRNG[124])|(((m[89]&~m[375]&~m[571])|(~m[89]&m[375]&m[571]))&~BiasedRNG[124])|((~m[89]&~m[375]&m[571])|(m[89]&~m[375]&m[571])|(m[89]&m[375]&m[571]))):InitCond[152];
    m[297] = run?((((~m[89]&~m[389]&~m[585])|(m[89]&m[389]&~m[585]))&BiasedRNG[125])|(((m[89]&~m[389]&~m[585])|(~m[89]&m[389]&m[585]))&~BiasedRNG[125])|((~m[89]&~m[389]&m[585])|(m[89]&~m[389]&m[585])|(m[89]&m[389]&m[585]))):InitCond[153];
    m[298] = run?((((~m[89]&~m[403]&~m[599])|(m[89]&m[403]&~m[599]))&BiasedRNG[126])|(((m[89]&~m[403]&~m[599])|(~m[89]&m[403]&m[599]))&~BiasedRNG[126])|((~m[89]&~m[403]&m[599])|(m[89]&~m[403]&m[599])|(m[89]&m[403]&m[599]))):InitCond[154];
    m[299] = run?((((~m[89]&~m[417]&~m[613])|(m[89]&m[417]&~m[613]))&BiasedRNG[127])|(((m[89]&~m[417]&~m[613])|(~m[89]&m[417]&m[613]))&~BiasedRNG[127])|((~m[89]&~m[417]&m[613])|(m[89]&~m[417]&m[613])|(m[89]&m[417]&m[613]))):InitCond[155];
    m[308] = run?((((~m[40]&~m[348]&~m[544])|(m[40]&m[348]&~m[544]))&BiasedRNG[128])|(((m[40]&~m[348]&~m[544])|(~m[40]&m[348]&m[544]))&~BiasedRNG[128])|((~m[40]&~m[348]&m[544])|(m[40]&~m[348]&m[544])|(m[40]&m[348]&m[544]))):InitCond[156];
    m[309] = run?((((~m[40]&~m[362]&~m[558])|(m[40]&m[362]&~m[558]))&BiasedRNG[129])|(((m[40]&~m[362]&~m[558])|(~m[40]&m[362]&m[558]))&~BiasedRNG[129])|((~m[40]&~m[362]&m[558])|(m[40]&~m[362]&m[558])|(m[40]&m[362]&m[558]))):InitCond[157];
    m[310] = run?((((~m[92]&~m[376]&~m[572])|(m[92]&m[376]&~m[572]))&BiasedRNG[130])|(((m[92]&~m[376]&~m[572])|(~m[92]&m[376]&m[572]))&~BiasedRNG[130])|((~m[92]&~m[376]&m[572])|(m[92]&~m[376]&m[572])|(m[92]&m[376]&m[572]))):InitCond[158];
    m[311] = run?((((~m[92]&~m[390]&~m[586])|(m[92]&m[390]&~m[586]))&BiasedRNG[131])|(((m[92]&~m[390]&~m[586])|(~m[92]&m[390]&m[586]))&~BiasedRNG[131])|((~m[92]&~m[390]&m[586])|(m[92]&~m[390]&m[586])|(m[92]&m[390]&m[586]))):InitCond[159];
    m[312] = run?((((~m[92]&~m[404]&~m[600])|(m[92]&m[404]&~m[600]))&BiasedRNG[132])|(((m[92]&~m[404]&~m[600])|(~m[92]&m[404]&m[600]))&~BiasedRNG[132])|((~m[92]&~m[404]&m[600])|(m[92]&~m[404]&m[600])|(m[92]&m[404]&m[600]))):InitCond[160];
    m[313] = run?((((~m[92]&~m[418]&~m[614])|(m[92]&m[418]&~m[614]))&BiasedRNG[133])|(((m[92]&~m[418]&~m[614])|(~m[92]&m[418]&m[614]))&~BiasedRNG[133])|((~m[92]&~m[418]&m[614])|(m[92]&~m[418]&m[614])|(m[92]&m[418]&m[614]))):InitCond[161];
    m[322] = run?((((~m[41]&~m[349]&~m[545])|(m[41]&m[349]&~m[545]))&BiasedRNG[134])|(((m[41]&~m[349]&~m[545])|(~m[41]&m[349]&m[545]))&~BiasedRNG[134])|((~m[41]&~m[349]&m[545])|(m[41]&~m[349]&m[545])|(m[41]&m[349]&m[545]))):InitCond[162];
    m[323] = run?((((~m[41]&~m[363]&~m[559])|(m[41]&m[363]&~m[559]))&BiasedRNG[135])|(((m[41]&~m[363]&~m[559])|(~m[41]&m[363]&m[559]))&~BiasedRNG[135])|((~m[41]&~m[363]&m[559])|(m[41]&~m[363]&m[559])|(m[41]&m[363]&m[559]))):InitCond[163];
    m[324] = run?((((~m[95]&~m[377]&~m[573])|(m[95]&m[377]&~m[573]))&BiasedRNG[136])|(((m[95]&~m[377]&~m[573])|(~m[95]&m[377]&m[573]))&~BiasedRNG[136])|((~m[95]&~m[377]&m[573])|(m[95]&~m[377]&m[573])|(m[95]&m[377]&m[573]))):InitCond[164];
    m[325] = run?((((~m[95]&~m[391]&~m[587])|(m[95]&m[391]&~m[587]))&BiasedRNG[137])|(((m[95]&~m[391]&~m[587])|(~m[95]&m[391]&m[587]))&~BiasedRNG[137])|((~m[95]&~m[391]&m[587])|(m[95]&~m[391]&m[587])|(m[95]&m[391]&m[587]))):InitCond[165];
    m[326] = run?((((~m[95]&~m[405]&~m[601])|(m[95]&m[405]&~m[601]))&BiasedRNG[138])|(((m[95]&~m[405]&~m[601])|(~m[95]&m[405]&m[601]))&~BiasedRNG[138])|((~m[95]&~m[405]&m[601])|(m[95]&~m[405]&m[601])|(m[95]&m[405]&m[601]))):InitCond[166];
    m[327] = run?((((~m[95]&~m[419]&~m[615])|(m[95]&m[419]&~m[615]))&BiasedRNG[139])|(((m[95]&~m[419]&~m[615])|(~m[95]&m[419]&m[615]))&~BiasedRNG[139])|((~m[95]&~m[419]&m[615])|(m[95]&~m[419]&m[615])|(m[95]&m[419]&m[615]))):InitCond[167];
    m[420] = run?((((~m[48]&~m[146]&~m[616])|(m[48]&m[146]&~m[616]))&BiasedRNG[140])|(((m[48]&~m[146]&~m[616])|(~m[48]&m[146]&m[616]))&~BiasedRNG[140])|((~m[48]&~m[146]&m[616])|(m[48]&~m[146]&m[616])|(m[48]&m[146]&m[616]))):InitCond[168];
    m[421] = run?((((~m[48]&~m[160]&~m[617])|(m[48]&m[160]&~m[617]))&BiasedRNG[141])|(((m[48]&~m[160]&~m[617])|(~m[48]&m[160]&m[617]))&~BiasedRNG[141])|((~m[48]&~m[160]&m[617])|(m[48]&~m[160]&m[617])|(m[48]&m[160]&m[617]))):InitCond[169];
    m[422] = run?((((~m[116]&~m[174]&~m[618])|(m[116]&m[174]&~m[618]))&BiasedRNG[142])|(((m[116]&~m[174]&~m[618])|(~m[116]&m[174]&m[618]))&~BiasedRNG[142])|((~m[116]&~m[174]&m[618])|(m[116]&~m[174]&m[618])|(m[116]&m[174]&m[618]))):InitCond[170];
    m[423] = run?((((~m[116]&~m[188]&~m[619])|(m[116]&m[188]&~m[619]))&BiasedRNG[143])|(((m[116]&~m[188]&~m[619])|(~m[116]&m[188]&m[619]))&~BiasedRNG[143])|((~m[116]&~m[188]&m[619])|(m[116]&~m[188]&m[619])|(m[116]&m[188]&m[619]))):InitCond[171];
    m[424] = run?((((~m[116]&~m[202]&~m[620])|(m[116]&m[202]&~m[620]))&BiasedRNG[144])|(((m[116]&~m[202]&~m[620])|(~m[116]&m[202]&m[620]))&~BiasedRNG[144])|((~m[116]&~m[202]&m[620])|(m[116]&~m[202]&m[620])|(m[116]&m[202]&m[620]))):InitCond[172];
    m[425] = run?((((~m[116]&~m[216]&~m[621])|(m[116]&m[216]&~m[621]))&BiasedRNG[145])|(((m[116]&~m[216]&~m[621])|(~m[116]&m[216]&m[621]))&~BiasedRNG[145])|((~m[116]&~m[216]&m[621])|(m[116]&~m[216]&m[621])|(m[116]&m[216]&m[621]))):InitCond[173];
    m[434] = run?((((~m[49]&~m[147]&~m[630])|(m[49]&m[147]&~m[630]))&BiasedRNG[146])|(((m[49]&~m[147]&~m[630])|(~m[49]&m[147]&m[630]))&~BiasedRNG[146])|((~m[49]&~m[147]&m[630])|(m[49]&~m[147]&m[630])|(m[49]&m[147]&m[630]))):InitCond[174];
    m[435] = run?((((~m[49]&~m[161]&~m[631])|(m[49]&m[161]&~m[631]))&BiasedRNG[147])|(((m[49]&~m[161]&~m[631])|(~m[49]&m[161]&m[631]))&~BiasedRNG[147])|((~m[49]&~m[161]&m[631])|(m[49]&~m[161]&m[631])|(m[49]&m[161]&m[631]))):InitCond[175];
    m[436] = run?((((~m[119]&~m[175]&~m[632])|(m[119]&m[175]&~m[632]))&BiasedRNG[148])|(((m[119]&~m[175]&~m[632])|(~m[119]&m[175]&m[632]))&~BiasedRNG[148])|((~m[119]&~m[175]&m[632])|(m[119]&~m[175]&m[632])|(m[119]&m[175]&m[632]))):InitCond[176];
    m[437] = run?((((~m[119]&~m[189]&~m[633])|(m[119]&m[189]&~m[633]))&BiasedRNG[149])|(((m[119]&~m[189]&~m[633])|(~m[119]&m[189]&m[633]))&~BiasedRNG[149])|((~m[119]&~m[189]&m[633])|(m[119]&~m[189]&m[633])|(m[119]&m[189]&m[633]))):InitCond[177];
    m[438] = run?((((~m[119]&~m[203]&~m[634])|(m[119]&m[203]&~m[634]))&BiasedRNG[150])|(((m[119]&~m[203]&~m[634])|(~m[119]&m[203]&m[634]))&~BiasedRNG[150])|((~m[119]&~m[203]&m[634])|(m[119]&~m[203]&m[634])|(m[119]&m[203]&m[634]))):InitCond[178];
    m[439] = run?((((~m[119]&~m[217]&~m[635])|(m[119]&m[217]&~m[635]))&BiasedRNG[151])|(((m[119]&~m[217]&~m[635])|(~m[119]&m[217]&m[635]))&~BiasedRNG[151])|((~m[119]&~m[217]&m[635])|(m[119]&~m[217]&m[635])|(m[119]&m[217]&m[635]))):InitCond[179];
    m[448] = run?((((~m[50]&~m[148]&~m[644])|(m[50]&m[148]&~m[644]))&BiasedRNG[152])|(((m[50]&~m[148]&~m[644])|(~m[50]&m[148]&m[644]))&~BiasedRNG[152])|((~m[50]&~m[148]&m[644])|(m[50]&~m[148]&m[644])|(m[50]&m[148]&m[644]))):InitCond[180];
    m[449] = run?((((~m[50]&~m[162]&~m[645])|(m[50]&m[162]&~m[645]))&BiasedRNG[153])|(((m[50]&~m[162]&~m[645])|(~m[50]&m[162]&m[645]))&~BiasedRNG[153])|((~m[50]&~m[162]&m[645])|(m[50]&~m[162]&m[645])|(m[50]&m[162]&m[645]))):InitCond[181];
    m[450] = run?((((~m[122]&~m[176]&~m[646])|(m[122]&m[176]&~m[646]))&BiasedRNG[154])|(((m[122]&~m[176]&~m[646])|(~m[122]&m[176]&m[646]))&~BiasedRNG[154])|((~m[122]&~m[176]&m[646])|(m[122]&~m[176]&m[646])|(m[122]&m[176]&m[646]))):InitCond[182];
    m[451] = run?((((~m[122]&~m[190]&~m[647])|(m[122]&m[190]&~m[647]))&BiasedRNG[155])|(((m[122]&~m[190]&~m[647])|(~m[122]&m[190]&m[647]))&~BiasedRNG[155])|((~m[122]&~m[190]&m[647])|(m[122]&~m[190]&m[647])|(m[122]&m[190]&m[647]))):InitCond[183];
    m[452] = run?((((~m[122]&~m[204]&~m[648])|(m[122]&m[204]&~m[648]))&BiasedRNG[156])|(((m[122]&~m[204]&~m[648])|(~m[122]&m[204]&m[648]))&~BiasedRNG[156])|((~m[122]&~m[204]&m[648])|(m[122]&~m[204]&m[648])|(m[122]&m[204]&m[648]))):InitCond[184];
    m[453] = run?((((~m[122]&~m[218]&~m[649])|(m[122]&m[218]&~m[649]))&BiasedRNG[157])|(((m[122]&~m[218]&~m[649])|(~m[122]&m[218]&m[649]))&~BiasedRNG[157])|((~m[122]&~m[218]&m[649])|(m[122]&~m[218]&m[649])|(m[122]&m[218]&m[649]))):InitCond[185];
    m[462] = run?((((~m[51]&~m[149]&~m[658])|(m[51]&m[149]&~m[658]))&BiasedRNG[158])|(((m[51]&~m[149]&~m[658])|(~m[51]&m[149]&m[658]))&~BiasedRNG[158])|((~m[51]&~m[149]&m[658])|(m[51]&~m[149]&m[658])|(m[51]&m[149]&m[658]))):InitCond[186];
    m[463] = run?((((~m[51]&~m[163]&~m[659])|(m[51]&m[163]&~m[659]))&BiasedRNG[159])|(((m[51]&~m[163]&~m[659])|(~m[51]&m[163]&m[659]))&~BiasedRNG[159])|((~m[51]&~m[163]&m[659])|(m[51]&~m[163]&m[659])|(m[51]&m[163]&m[659]))):InitCond[187];
    m[464] = run?((((~m[125]&~m[177]&~m[660])|(m[125]&m[177]&~m[660]))&BiasedRNG[160])|(((m[125]&~m[177]&~m[660])|(~m[125]&m[177]&m[660]))&~BiasedRNG[160])|((~m[125]&~m[177]&m[660])|(m[125]&~m[177]&m[660])|(m[125]&m[177]&m[660]))):InitCond[188];
    m[465] = run?((((~m[125]&~m[191]&~m[661])|(m[125]&m[191]&~m[661]))&BiasedRNG[161])|(((m[125]&~m[191]&~m[661])|(~m[125]&m[191]&m[661]))&~BiasedRNG[161])|((~m[125]&~m[191]&m[661])|(m[125]&~m[191]&m[661])|(m[125]&m[191]&m[661]))):InitCond[189];
    m[466] = run?((((~m[125]&~m[205]&~m[662])|(m[125]&m[205]&~m[662]))&BiasedRNG[162])|(((m[125]&~m[205]&~m[662])|(~m[125]&m[205]&m[662]))&~BiasedRNG[162])|((~m[125]&~m[205]&m[662])|(m[125]&~m[205]&m[662])|(m[125]&m[205]&m[662]))):InitCond[190];
    m[467] = run?((((~m[125]&~m[219]&~m[663])|(m[125]&m[219]&~m[663]))&BiasedRNG[163])|(((m[125]&~m[219]&~m[663])|(~m[125]&m[219]&m[663]))&~BiasedRNG[163])|((~m[125]&~m[219]&m[663])|(m[125]&~m[219]&m[663])|(m[125]&m[219]&m[663]))):InitCond[191];
    m[476] = run?((((~m[52]&~m[150]&~m[672])|(m[52]&m[150]&~m[672]))&BiasedRNG[164])|(((m[52]&~m[150]&~m[672])|(~m[52]&m[150]&m[672]))&~BiasedRNG[164])|((~m[52]&~m[150]&m[672])|(m[52]&~m[150]&m[672])|(m[52]&m[150]&m[672]))):InitCond[192];
    m[477] = run?((((~m[52]&~m[164]&~m[673])|(m[52]&m[164]&~m[673]))&BiasedRNG[165])|(((m[52]&~m[164]&~m[673])|(~m[52]&m[164]&m[673]))&~BiasedRNG[165])|((~m[52]&~m[164]&m[673])|(m[52]&~m[164]&m[673])|(m[52]&m[164]&m[673]))):InitCond[193];
    m[478] = run?((((~m[128]&~m[178]&~m[674])|(m[128]&m[178]&~m[674]))&BiasedRNG[166])|(((m[128]&~m[178]&~m[674])|(~m[128]&m[178]&m[674]))&~BiasedRNG[166])|((~m[128]&~m[178]&m[674])|(m[128]&~m[178]&m[674])|(m[128]&m[178]&m[674]))):InitCond[194];
    m[479] = run?((((~m[128]&~m[192]&~m[675])|(m[128]&m[192]&~m[675]))&BiasedRNG[167])|(((m[128]&~m[192]&~m[675])|(~m[128]&m[192]&m[675]))&~BiasedRNG[167])|((~m[128]&~m[192]&m[675])|(m[128]&~m[192]&m[675])|(m[128]&m[192]&m[675]))):InitCond[195];
    m[480] = run?((((~m[128]&~m[206]&~m[676])|(m[128]&m[206]&~m[676]))&BiasedRNG[168])|(((m[128]&~m[206]&~m[676])|(~m[128]&m[206]&m[676]))&~BiasedRNG[168])|((~m[128]&~m[206]&m[676])|(m[128]&~m[206]&m[676])|(m[128]&m[206]&m[676]))):InitCond[196];
    m[481] = run?((((~m[128]&~m[220]&~m[677])|(m[128]&m[220]&~m[677]))&BiasedRNG[169])|(((m[128]&~m[220]&~m[677])|(~m[128]&m[220]&m[677]))&~BiasedRNG[169])|((~m[128]&~m[220]&m[677])|(m[128]&~m[220]&m[677])|(m[128]&m[220]&m[677]))):InitCond[197];
    m[490] = run?((((~m[53]&~m[151]&~m[686])|(m[53]&m[151]&~m[686]))&BiasedRNG[170])|(((m[53]&~m[151]&~m[686])|(~m[53]&m[151]&m[686]))&~BiasedRNG[170])|((~m[53]&~m[151]&m[686])|(m[53]&~m[151]&m[686])|(m[53]&m[151]&m[686]))):InitCond[198];
    m[491] = run?((((~m[53]&~m[165]&~m[687])|(m[53]&m[165]&~m[687]))&BiasedRNG[171])|(((m[53]&~m[165]&~m[687])|(~m[53]&m[165]&m[687]))&~BiasedRNG[171])|((~m[53]&~m[165]&m[687])|(m[53]&~m[165]&m[687])|(m[53]&m[165]&m[687]))):InitCond[199];
    m[492] = run?((((~m[131]&~m[179]&~m[688])|(m[131]&m[179]&~m[688]))&BiasedRNG[172])|(((m[131]&~m[179]&~m[688])|(~m[131]&m[179]&m[688]))&~BiasedRNG[172])|((~m[131]&~m[179]&m[688])|(m[131]&~m[179]&m[688])|(m[131]&m[179]&m[688]))):InitCond[200];
    m[493] = run?((((~m[131]&~m[193]&~m[689])|(m[131]&m[193]&~m[689]))&BiasedRNG[173])|(((m[131]&~m[193]&~m[689])|(~m[131]&m[193]&m[689]))&~BiasedRNG[173])|((~m[131]&~m[193]&m[689])|(m[131]&~m[193]&m[689])|(m[131]&m[193]&m[689]))):InitCond[201];
    m[494] = run?((((~m[131]&~m[207]&~m[690])|(m[131]&m[207]&~m[690]))&BiasedRNG[174])|(((m[131]&~m[207]&~m[690])|(~m[131]&m[207]&m[690]))&~BiasedRNG[174])|((~m[131]&~m[207]&m[690])|(m[131]&~m[207]&m[690])|(m[131]&m[207]&m[690]))):InitCond[202];
    m[495] = run?((((~m[131]&~m[221]&~m[691])|(m[131]&m[221]&~m[691]))&BiasedRNG[175])|(((m[131]&~m[221]&~m[691])|(~m[131]&m[221]&m[691]))&~BiasedRNG[175])|((~m[131]&~m[221]&m[691])|(m[131]&~m[221]&m[691])|(m[131]&m[221]&m[691]))):InitCond[203];
    m[504] = run?((((~m[54]&~m[152]&~m[700])|(m[54]&m[152]&~m[700]))&BiasedRNG[176])|(((m[54]&~m[152]&~m[700])|(~m[54]&m[152]&m[700]))&~BiasedRNG[176])|((~m[54]&~m[152]&m[700])|(m[54]&~m[152]&m[700])|(m[54]&m[152]&m[700]))):InitCond[204];
    m[505] = run?((((~m[54]&~m[166]&~m[701])|(m[54]&m[166]&~m[701]))&BiasedRNG[177])|(((m[54]&~m[166]&~m[701])|(~m[54]&m[166]&m[701]))&~BiasedRNG[177])|((~m[54]&~m[166]&m[701])|(m[54]&~m[166]&m[701])|(m[54]&m[166]&m[701]))):InitCond[205];
    m[506] = run?((((~m[134]&~m[180]&~m[702])|(m[134]&m[180]&~m[702]))&BiasedRNG[178])|(((m[134]&~m[180]&~m[702])|(~m[134]&m[180]&m[702]))&~BiasedRNG[178])|((~m[134]&~m[180]&m[702])|(m[134]&~m[180]&m[702])|(m[134]&m[180]&m[702]))):InitCond[206];
    m[507] = run?((((~m[134]&~m[194]&~m[703])|(m[134]&m[194]&~m[703]))&BiasedRNG[179])|(((m[134]&~m[194]&~m[703])|(~m[134]&m[194]&m[703]))&~BiasedRNG[179])|((~m[134]&~m[194]&m[703])|(m[134]&~m[194]&m[703])|(m[134]&m[194]&m[703]))):InitCond[207];
    m[508] = run?((((~m[134]&~m[208]&~m[704])|(m[134]&m[208]&~m[704]))&BiasedRNG[180])|(((m[134]&~m[208]&~m[704])|(~m[134]&m[208]&m[704]))&~BiasedRNG[180])|((~m[134]&~m[208]&m[704])|(m[134]&~m[208]&m[704])|(m[134]&m[208]&m[704]))):InitCond[208];
    m[509] = run?((((~m[134]&~m[222]&~m[705])|(m[134]&m[222]&~m[705]))&BiasedRNG[181])|(((m[134]&~m[222]&~m[705])|(~m[134]&m[222]&m[705]))&~BiasedRNG[181])|((~m[134]&~m[222]&m[705])|(m[134]&~m[222]&m[705])|(m[134]&m[222]&m[705]))):InitCond[209];
    m[518] = run?((((~m[55]&~m[153]&~m[714])|(m[55]&m[153]&~m[714]))&BiasedRNG[182])|(((m[55]&~m[153]&~m[714])|(~m[55]&m[153]&m[714]))&~BiasedRNG[182])|((~m[55]&~m[153]&m[714])|(m[55]&~m[153]&m[714])|(m[55]&m[153]&m[714]))):InitCond[210];
    m[519] = run?((((~m[55]&~m[167]&~m[715])|(m[55]&m[167]&~m[715]))&BiasedRNG[183])|(((m[55]&~m[167]&~m[715])|(~m[55]&m[167]&m[715]))&~BiasedRNG[183])|((~m[55]&~m[167]&m[715])|(m[55]&~m[167]&m[715])|(m[55]&m[167]&m[715]))):InitCond[211];
    m[520] = run?((((~m[137]&~m[181]&~m[716])|(m[137]&m[181]&~m[716]))&BiasedRNG[184])|(((m[137]&~m[181]&~m[716])|(~m[137]&m[181]&m[716]))&~BiasedRNG[184])|((~m[137]&~m[181]&m[716])|(m[137]&~m[181]&m[716])|(m[137]&m[181]&m[716]))):InitCond[212];
    m[521] = run?((((~m[137]&~m[195]&~m[717])|(m[137]&m[195]&~m[717]))&BiasedRNG[185])|(((m[137]&~m[195]&~m[717])|(~m[137]&m[195]&m[717]))&~BiasedRNG[185])|((~m[137]&~m[195]&m[717])|(m[137]&~m[195]&m[717])|(m[137]&m[195]&m[717]))):InitCond[213];
    m[522] = run?((((~m[137]&~m[209]&~m[718])|(m[137]&m[209]&~m[718]))&BiasedRNG[186])|(((m[137]&~m[209]&~m[718])|(~m[137]&m[209]&m[718]))&~BiasedRNG[186])|((~m[137]&~m[209]&m[718])|(m[137]&~m[209]&m[718])|(m[137]&m[209]&m[718]))):InitCond[214];
    m[523] = run?((((~m[137]&~m[223]&~m[719])|(m[137]&m[223]&~m[719]))&BiasedRNG[187])|(((m[137]&~m[223]&~m[719])|(~m[137]&m[223]&m[719]))&~BiasedRNG[187])|((~m[137]&~m[223]&m[719])|(m[137]&~m[223]&m[719])|(m[137]&m[223]&m[719]))):InitCond[215];
    m[622] = run?((((m[230]&~m[426]&m[1084])|(~m[230]&m[426]&m[1084]))&BiasedRNG[188])|(((m[230]&m[426]&~m[1084]))&~BiasedRNG[188])|((m[230]&m[426]&m[1084]))):InitCond[216];
    m[623] = run?((((m[244]&~m[427]&m[1144])|(~m[244]&m[427]&m[1144]))&BiasedRNG[189])|(((m[244]&m[427]&~m[1144]))&~BiasedRNG[189])|((m[244]&m[427]&m[1144]))):InitCond[217];
    m[624] = run?((((m[258]&~m[428]&m[1209])|(~m[258]&m[428]&m[1209]))&BiasedRNG[190])|(((m[258]&m[428]&~m[1209]))&~BiasedRNG[190])|((m[258]&m[428]&m[1209]))):InitCond[218];
    m[625] = run?((((m[272]&~m[429]&m[1269])|(~m[272]&m[429]&m[1269]))&BiasedRNG[191])|(((m[272]&m[429]&~m[1269]))&~BiasedRNG[191])|((m[272]&m[429]&m[1269]))):InitCond[219];
    m[626] = run?((((m[286]&~m[430]&m[1324])|(~m[286]&m[430]&m[1324]))&BiasedRNG[192])|(((m[286]&m[430]&~m[1324]))&~BiasedRNG[192])|((m[286]&m[430]&m[1324]))):InitCond[220];
    m[627] = run?((((m[300]&~m[431]&m[1374])|(~m[300]&m[431]&m[1374]))&BiasedRNG[193])|(((m[300]&m[431]&~m[1374]))&~BiasedRNG[193])|((m[300]&m[431]&m[1374]))):InitCond[221];
    m[628] = run?((((m[314]&~m[432]&m[1419])|(~m[314]&m[432]&m[1419]))&BiasedRNG[194])|(((m[314]&m[432]&~m[1419]))&~BiasedRNG[194])|((m[314]&m[432]&m[1419]))):InitCond[222];
    m[629] = run?((((m[328]&~m[433]&m[1459])|(~m[328]&m[433]&m[1459]))&BiasedRNG[195])|(((m[328]&m[433]&~m[1459]))&~BiasedRNG[195])|((m[328]&m[433]&m[1459]))):InitCond[223];
    m[636] = run?((((m[231]&~m[440]&m[1149])|(~m[231]&m[440]&m[1149]))&BiasedRNG[196])|(((m[231]&m[440]&~m[1149]))&~BiasedRNG[196])|((m[231]&m[440]&m[1149]))):InitCond[224];
    m[637] = run?((((m[245]&~m[441]&m[1214])|(~m[245]&m[441]&m[1214]))&BiasedRNG[197])|(((m[245]&m[441]&~m[1214]))&~BiasedRNG[197])|((m[245]&m[441]&m[1214]))):InitCond[225];
    m[638] = run?((((m[259]&~m[442]&m[1274])|(~m[259]&m[442]&m[1274]))&BiasedRNG[198])|(((m[259]&m[442]&~m[1274]))&~BiasedRNG[198])|((m[259]&m[442]&m[1274]))):InitCond[226];
    m[639] = run?((((m[273]&~m[443]&m[1329])|(~m[273]&m[443]&m[1329]))&BiasedRNG[199])|(((m[273]&m[443]&~m[1329]))&~BiasedRNG[199])|((m[273]&m[443]&m[1329]))):InitCond[227];
    m[640] = run?((((m[287]&~m[444]&m[1379])|(~m[287]&m[444]&m[1379]))&BiasedRNG[200])|(((m[287]&m[444]&~m[1379]))&~BiasedRNG[200])|((m[287]&m[444]&m[1379]))):InitCond[228];
    m[641] = run?((((m[301]&~m[445]&m[1424])|(~m[301]&m[445]&m[1424]))&BiasedRNG[201])|(((m[301]&m[445]&~m[1424]))&~BiasedRNG[201])|((m[301]&m[445]&m[1424]))):InitCond[229];
    m[642] = run?((((m[315]&~m[446]&m[1464])|(~m[315]&m[446]&m[1464]))&BiasedRNG[202])|(((m[315]&m[446]&~m[1464]))&~BiasedRNG[202])|((m[315]&m[446]&m[1464]))):InitCond[230];
    m[643] = run?((((m[329]&~m[447]&m[1499])|(~m[329]&m[447]&m[1499]))&BiasedRNG[203])|(((m[329]&m[447]&~m[1499]))&~BiasedRNG[203])|((m[329]&m[447]&m[1499]))):InitCond[231];
    m[650] = run?((((m[232]&~m[454]&m[1219])|(~m[232]&m[454]&m[1219]))&BiasedRNG[204])|(((m[232]&m[454]&~m[1219]))&~BiasedRNG[204])|((m[232]&m[454]&m[1219]))):InitCond[232];
    m[651] = run?((((m[246]&~m[455]&m[1279])|(~m[246]&m[455]&m[1279]))&BiasedRNG[205])|(((m[246]&m[455]&~m[1279]))&~BiasedRNG[205])|((m[246]&m[455]&m[1279]))):InitCond[233];
    m[652] = run?((((m[260]&~m[456]&m[1334])|(~m[260]&m[456]&m[1334]))&BiasedRNG[206])|(((m[260]&m[456]&~m[1334]))&~BiasedRNG[206])|((m[260]&m[456]&m[1334]))):InitCond[234];
    m[653] = run?((((m[274]&~m[457]&m[1384])|(~m[274]&m[457]&m[1384]))&BiasedRNG[207])|(((m[274]&m[457]&~m[1384]))&~BiasedRNG[207])|((m[274]&m[457]&m[1384]))):InitCond[235];
    m[654] = run?((((m[288]&~m[458]&m[1429])|(~m[288]&m[458]&m[1429]))&BiasedRNG[208])|(((m[288]&m[458]&~m[1429]))&~BiasedRNG[208])|((m[288]&m[458]&m[1429]))):InitCond[236];
    m[655] = run?((((m[302]&~m[459]&m[1469])|(~m[302]&m[459]&m[1469]))&BiasedRNG[209])|(((m[302]&m[459]&~m[1469]))&~BiasedRNG[209])|((m[302]&m[459]&m[1469]))):InitCond[237];
    m[656] = run?((((m[316]&~m[460]&m[1504])|(~m[316]&m[460]&m[1504]))&BiasedRNG[210])|(((m[316]&m[460]&~m[1504]))&~BiasedRNG[210])|((m[316]&m[460]&m[1504]))):InitCond[238];
    m[657] = run?((((m[330]&~m[461]&m[1534])|(~m[330]&m[461]&m[1534]))&BiasedRNG[211])|(((m[330]&m[461]&~m[1534]))&~BiasedRNG[211])|((m[330]&m[461]&m[1534]))):InitCond[239];
    m[664] = run?((((m[233]&~m[468]&m[1284])|(~m[233]&m[468]&m[1284]))&BiasedRNG[212])|(((m[233]&m[468]&~m[1284]))&~BiasedRNG[212])|((m[233]&m[468]&m[1284]))):InitCond[240];
    m[665] = run?((((m[247]&~m[469]&m[1339])|(~m[247]&m[469]&m[1339]))&BiasedRNG[213])|(((m[247]&m[469]&~m[1339]))&~BiasedRNG[213])|((m[247]&m[469]&m[1339]))):InitCond[241];
    m[666] = run?((((m[261]&~m[470]&m[1389])|(~m[261]&m[470]&m[1389]))&BiasedRNG[214])|(((m[261]&m[470]&~m[1389]))&~BiasedRNG[214])|((m[261]&m[470]&m[1389]))):InitCond[242];
    m[667] = run?((((m[275]&~m[471]&m[1434])|(~m[275]&m[471]&m[1434]))&BiasedRNG[215])|(((m[275]&m[471]&~m[1434]))&~BiasedRNG[215])|((m[275]&m[471]&m[1434]))):InitCond[243];
    m[668] = run?((((m[289]&~m[472]&m[1474])|(~m[289]&m[472]&m[1474]))&BiasedRNG[216])|(((m[289]&m[472]&~m[1474]))&~BiasedRNG[216])|((m[289]&m[472]&m[1474]))):InitCond[244];
    m[669] = run?((((m[303]&~m[473]&m[1509])|(~m[303]&m[473]&m[1509]))&BiasedRNG[217])|(((m[303]&m[473]&~m[1509]))&~BiasedRNG[217])|((m[303]&m[473]&m[1509]))):InitCond[245];
    m[670] = run?((((m[317]&~m[474]&m[1539])|(~m[317]&m[474]&m[1539]))&BiasedRNG[218])|(((m[317]&m[474]&~m[1539]))&~BiasedRNG[218])|((m[317]&m[474]&m[1539]))):InitCond[246];
    m[671] = run?((((m[331]&~m[475]&m[1564])|(~m[331]&m[475]&m[1564]))&BiasedRNG[219])|(((m[331]&m[475]&~m[1564]))&~BiasedRNG[219])|((m[331]&m[475]&m[1564]))):InitCond[247];
    m[678] = run?((((m[234]&~m[482]&m[1344])|(~m[234]&m[482]&m[1344]))&BiasedRNG[220])|(((m[234]&m[482]&~m[1344]))&~BiasedRNG[220])|((m[234]&m[482]&m[1344]))):InitCond[248];
    m[679] = run?((((m[248]&~m[483]&m[1394])|(~m[248]&m[483]&m[1394]))&BiasedRNG[221])|(((m[248]&m[483]&~m[1394]))&~BiasedRNG[221])|((m[248]&m[483]&m[1394]))):InitCond[249];
    m[680] = run?((((m[262]&~m[484]&m[1439])|(~m[262]&m[484]&m[1439]))&BiasedRNG[222])|(((m[262]&m[484]&~m[1439]))&~BiasedRNG[222])|((m[262]&m[484]&m[1439]))):InitCond[250];
    m[681] = run?((((m[276]&~m[485]&m[1479])|(~m[276]&m[485]&m[1479]))&BiasedRNG[223])|(((m[276]&m[485]&~m[1479]))&~BiasedRNG[223])|((m[276]&m[485]&m[1479]))):InitCond[251];
    m[682] = run?((((m[290]&~m[486]&m[1514])|(~m[290]&m[486]&m[1514]))&BiasedRNG[224])|(((m[290]&m[486]&~m[1514]))&~BiasedRNG[224])|((m[290]&m[486]&m[1514]))):InitCond[252];
    m[683] = run?((((m[304]&~m[487]&m[1544])|(~m[304]&m[487]&m[1544]))&BiasedRNG[225])|(((m[304]&m[487]&~m[1544]))&~BiasedRNG[225])|((m[304]&m[487]&m[1544]))):InitCond[253];
    m[684] = run?((((m[318]&~m[488]&m[1569])|(~m[318]&m[488]&m[1569]))&BiasedRNG[226])|(((m[318]&m[488]&~m[1569]))&~BiasedRNG[226])|((m[318]&m[488]&m[1569]))):InitCond[254];
    m[685] = run?((((m[332]&~m[489]&m[1589])|(~m[332]&m[489]&m[1589]))&BiasedRNG[227])|(((m[332]&m[489]&~m[1589]))&~BiasedRNG[227])|((m[332]&m[489]&m[1589]))):InitCond[255];
    m[692] = run?((((m[235]&~m[496]&m[1399])|(~m[235]&m[496]&m[1399]))&BiasedRNG[228])|(((m[235]&m[496]&~m[1399]))&~BiasedRNG[228])|((m[235]&m[496]&m[1399]))):InitCond[256];
    m[693] = run?((((m[249]&~m[497]&m[1444])|(~m[249]&m[497]&m[1444]))&BiasedRNG[229])|(((m[249]&m[497]&~m[1444]))&~BiasedRNG[229])|((m[249]&m[497]&m[1444]))):InitCond[257];
    m[694] = run?((((m[263]&~m[498]&m[1484])|(~m[263]&m[498]&m[1484]))&BiasedRNG[230])|(((m[263]&m[498]&~m[1484]))&~BiasedRNG[230])|((m[263]&m[498]&m[1484]))):InitCond[258];
    m[695] = run?((((m[277]&~m[499]&m[1519])|(~m[277]&m[499]&m[1519]))&BiasedRNG[231])|(((m[277]&m[499]&~m[1519]))&~BiasedRNG[231])|((m[277]&m[499]&m[1519]))):InitCond[259];
    m[696] = run?((((m[291]&~m[500]&m[1549])|(~m[291]&m[500]&m[1549]))&BiasedRNG[232])|(((m[291]&m[500]&~m[1549]))&~BiasedRNG[232])|((m[291]&m[500]&m[1549]))):InitCond[260];
    m[697] = run?((((m[305]&~m[501]&m[1574])|(~m[305]&m[501]&m[1574]))&BiasedRNG[233])|(((m[305]&m[501]&~m[1574]))&~BiasedRNG[233])|((m[305]&m[501]&m[1574]))):InitCond[261];
    m[698] = run?((((m[319]&~m[502]&m[1594])|(~m[319]&m[502]&m[1594]))&BiasedRNG[234])|(((m[319]&m[502]&~m[1594]))&~BiasedRNG[234])|((m[319]&m[502]&m[1594]))):InitCond[262];
    m[699] = run?((((m[333]&~m[503]&m[1609])|(~m[333]&m[503]&m[1609]))&BiasedRNG[235])|(((m[333]&m[503]&~m[1609]))&~BiasedRNG[235])|((m[333]&m[503]&m[1609]))):InitCond[263];
    m[706] = run?((((m[236]&~m[510]&m[1449])|(~m[236]&m[510]&m[1449]))&BiasedRNG[236])|(((m[236]&m[510]&~m[1449]))&~BiasedRNG[236])|((m[236]&m[510]&m[1449]))):InitCond[264];
    m[707] = run?((((m[250]&~m[511]&m[1489])|(~m[250]&m[511]&m[1489]))&BiasedRNG[237])|(((m[250]&m[511]&~m[1489]))&~BiasedRNG[237])|((m[250]&m[511]&m[1489]))):InitCond[265];
    m[708] = run?((((m[264]&~m[512]&m[1524])|(~m[264]&m[512]&m[1524]))&BiasedRNG[238])|(((m[264]&m[512]&~m[1524]))&~BiasedRNG[238])|((m[264]&m[512]&m[1524]))):InitCond[266];
    m[709] = run?((((m[278]&~m[513]&m[1554])|(~m[278]&m[513]&m[1554]))&BiasedRNG[239])|(((m[278]&m[513]&~m[1554]))&~BiasedRNG[239])|((m[278]&m[513]&m[1554]))):InitCond[267];
    m[710] = run?((((m[292]&~m[514]&m[1579])|(~m[292]&m[514]&m[1579]))&BiasedRNG[240])|(((m[292]&m[514]&~m[1579]))&~BiasedRNG[240])|((m[292]&m[514]&m[1579]))):InitCond[268];
    m[711] = run?((((m[306]&~m[515]&m[1599])|(~m[306]&m[515]&m[1599]))&BiasedRNG[241])|(((m[306]&m[515]&~m[1599]))&~BiasedRNG[241])|((m[306]&m[515]&m[1599]))):InitCond[269];
    m[712] = run?((((m[320]&~m[516]&m[1614])|(~m[320]&m[516]&m[1614]))&BiasedRNG[242])|(((m[320]&m[516]&~m[1614]))&~BiasedRNG[242])|((m[320]&m[516]&m[1614]))):InitCond[270];
    m[713] = run?((((m[334]&~m[517]&m[1624])|(~m[334]&m[517]&m[1624]))&BiasedRNG[243])|(((m[334]&m[517]&~m[1624]))&~BiasedRNG[243])|((m[334]&m[517]&m[1624]))):InitCond[271];
    m[720] = run?((((m[237]&~m[524]&m[1494])|(~m[237]&m[524]&m[1494]))&BiasedRNG[244])|(((m[237]&m[524]&~m[1494]))&~BiasedRNG[244])|((m[237]&m[524]&m[1494]))):InitCond[272];
    m[721] = run?((((m[251]&~m[525]&m[1529])|(~m[251]&m[525]&m[1529]))&BiasedRNG[245])|(((m[251]&m[525]&~m[1529]))&~BiasedRNG[245])|((m[251]&m[525]&m[1529]))):InitCond[273];
    m[722] = run?((((m[265]&~m[526]&m[1559])|(~m[265]&m[526]&m[1559]))&BiasedRNG[246])|(((m[265]&m[526]&~m[1559]))&~BiasedRNG[246])|((m[265]&m[526]&m[1559]))):InitCond[274];
    m[723] = run?((((m[279]&~m[527]&m[1584])|(~m[279]&m[527]&m[1584]))&BiasedRNG[247])|(((m[279]&m[527]&~m[1584]))&~BiasedRNG[247])|((m[279]&m[527]&m[1584]))):InitCond[275];
    m[724] = run?((((m[293]&~m[528]&m[1604])|(~m[293]&m[528]&m[1604]))&BiasedRNG[248])|(((m[293]&m[528]&~m[1604]))&~BiasedRNG[248])|((m[293]&m[528]&m[1604]))):InitCond[276];
    m[725] = run?((((m[307]&~m[529]&m[1619])|(~m[307]&m[529]&m[1619]))&BiasedRNG[249])|(((m[307]&m[529]&~m[1619]))&~BiasedRNG[249])|((m[307]&m[529]&m[1619]))):InitCond[277];
    m[726] = run?((((m[321]&~m[530]&m[1629])|(~m[321]&m[530]&m[1629]))&BiasedRNG[250])|(((m[321]&m[530]&~m[1629]))&~BiasedRNG[250])|((m[321]&m[530]&m[1629]))):InitCond[278];
    m[727] = run?((((m[335]&~m[531]&m[1634])|(~m[335]&m[531]&m[1634]))&BiasedRNG[251])|(((m[335]&m[531]&~m[1634]))&~BiasedRNG[251])|((m[335]&m[531]&m[1634]))):InitCond[279];
    m[728] = run?((((m[533]&~m[729]&~m[730]&~m[731]&~m[732])|(~m[533]&~m[729]&~m[730]&m[731]&~m[732])|(m[533]&m[729]&~m[730]&m[731]&~m[732])|(m[533]&~m[729]&m[730]&m[731]&~m[732])|(~m[533]&m[729]&~m[730]&~m[731]&m[732])|(~m[533]&~m[729]&m[730]&~m[731]&m[732])|(m[533]&m[729]&m[730]&~m[731]&m[732])|(~m[533]&m[729]&m[730]&m[731]&m[732]))&UnbiasedRNG[28])|((m[533]&~m[729]&~m[730]&m[731]&~m[732])|(~m[533]&~m[729]&~m[730]&~m[731]&m[732])|(m[533]&~m[729]&~m[730]&~m[731]&m[732])|(m[533]&m[729]&~m[730]&~m[731]&m[732])|(m[533]&~m[729]&m[730]&~m[731]&m[732])|(~m[533]&~m[729]&~m[730]&m[731]&m[732])|(m[533]&~m[729]&~m[730]&m[731]&m[732])|(~m[533]&m[729]&~m[730]&m[731]&m[732])|(m[533]&m[729]&~m[730]&m[731]&m[732])|(~m[533]&~m[729]&m[730]&m[731]&m[732])|(m[533]&~m[729]&m[730]&m[731]&m[732])|(m[533]&m[729]&m[730]&m[731]&m[732]))):InitCond[280];
    m[733] = run?((((m[534]&~m[734]&~m[735]&~m[736]&~m[737])|(~m[534]&~m[734]&~m[735]&m[736]&~m[737])|(m[534]&m[734]&~m[735]&m[736]&~m[737])|(m[534]&~m[734]&m[735]&m[736]&~m[737])|(~m[534]&m[734]&~m[735]&~m[736]&m[737])|(~m[534]&~m[734]&m[735]&~m[736]&m[737])|(m[534]&m[734]&m[735]&~m[736]&m[737])|(~m[534]&m[734]&m[735]&m[736]&m[737]))&UnbiasedRNG[29])|((m[534]&~m[734]&~m[735]&m[736]&~m[737])|(~m[534]&~m[734]&~m[735]&~m[736]&m[737])|(m[534]&~m[734]&~m[735]&~m[736]&m[737])|(m[534]&m[734]&~m[735]&~m[736]&m[737])|(m[534]&~m[734]&m[735]&~m[736]&m[737])|(~m[534]&~m[734]&~m[735]&m[736]&m[737])|(m[534]&~m[734]&~m[735]&m[736]&m[737])|(~m[534]&m[734]&~m[735]&m[736]&m[737])|(m[534]&m[734]&~m[735]&m[736]&m[737])|(~m[534]&~m[734]&m[735]&m[736]&m[737])|(m[534]&~m[734]&m[735]&m[736]&m[737])|(m[534]&m[734]&m[735]&m[736]&m[737]))):InitCond[281];
    m[738] = run?((((m[736]&~m[739]&~m[740]&~m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&m[741]&~m[742])|(m[736]&m[739]&~m[740]&m[741]&~m[742])|(m[736]&~m[739]&m[740]&m[741]&~m[742])|(~m[736]&m[739]&~m[740]&~m[741]&m[742])|(~m[736]&~m[739]&m[740]&~m[741]&m[742])|(m[736]&m[739]&m[740]&~m[741]&m[742])|(~m[736]&m[739]&m[740]&m[741]&m[742]))&UnbiasedRNG[30])|((m[736]&~m[739]&~m[740]&m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&m[740]&~m[741]&m[742])|(~m[736]&~m[739]&~m[740]&m[741]&m[742])|(m[736]&~m[739]&~m[740]&m[741]&m[742])|(~m[736]&m[739]&~m[740]&m[741]&m[742])|(m[736]&m[739]&~m[740]&m[741]&m[742])|(~m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&m[739]&m[740]&m[741]&m[742]))):InitCond[282];
    m[743] = run?((((m[535]&~m[744]&~m[745]&~m[746]&~m[747])|(~m[535]&~m[744]&~m[745]&m[746]&~m[747])|(m[535]&m[744]&~m[745]&m[746]&~m[747])|(m[535]&~m[744]&m[745]&m[746]&~m[747])|(~m[535]&m[744]&~m[745]&~m[746]&m[747])|(~m[535]&~m[744]&m[745]&~m[746]&m[747])|(m[535]&m[744]&m[745]&~m[746]&m[747])|(~m[535]&m[744]&m[745]&m[746]&m[747]))&UnbiasedRNG[31])|((m[535]&~m[744]&~m[745]&m[746]&~m[747])|(~m[535]&~m[744]&~m[745]&~m[746]&m[747])|(m[535]&~m[744]&~m[745]&~m[746]&m[747])|(m[535]&m[744]&~m[745]&~m[746]&m[747])|(m[535]&~m[744]&m[745]&~m[746]&m[747])|(~m[535]&~m[744]&~m[745]&m[746]&m[747])|(m[535]&~m[744]&~m[745]&m[746]&m[747])|(~m[535]&m[744]&~m[745]&m[746]&m[747])|(m[535]&m[744]&~m[745]&m[746]&m[747])|(~m[535]&~m[744]&m[745]&m[746]&m[747])|(m[535]&~m[744]&m[745]&m[746]&m[747])|(m[535]&m[744]&m[745]&m[746]&m[747]))):InitCond[283];
    m[748] = run?((((m[746]&~m[749]&~m[750]&~m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&m[751]&~m[752])|(m[746]&m[749]&~m[750]&m[751]&~m[752])|(m[746]&~m[749]&m[750]&m[751]&~m[752])|(~m[746]&m[749]&~m[750]&~m[751]&m[752])|(~m[746]&~m[749]&m[750]&~m[751]&m[752])|(m[746]&m[749]&m[750]&~m[751]&m[752])|(~m[746]&m[749]&m[750]&m[751]&m[752]))&UnbiasedRNG[32])|((m[746]&~m[749]&~m[750]&m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&m[750]&~m[751]&m[752])|(~m[746]&~m[749]&~m[750]&m[751]&m[752])|(m[746]&~m[749]&~m[750]&m[751]&m[752])|(~m[746]&m[749]&~m[750]&m[751]&m[752])|(m[746]&m[749]&~m[750]&m[751]&m[752])|(~m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&m[749]&m[750]&m[751]&m[752]))):InitCond[284];
    m[753] = run?((((m[751]&~m[754]&~m[755]&~m[756]&~m[757])|(~m[751]&~m[754]&~m[755]&m[756]&~m[757])|(m[751]&m[754]&~m[755]&m[756]&~m[757])|(m[751]&~m[754]&m[755]&m[756]&~m[757])|(~m[751]&m[754]&~m[755]&~m[756]&m[757])|(~m[751]&~m[754]&m[755]&~m[756]&m[757])|(m[751]&m[754]&m[755]&~m[756]&m[757])|(~m[751]&m[754]&m[755]&m[756]&m[757]))&UnbiasedRNG[33])|((m[751]&~m[754]&~m[755]&m[756]&~m[757])|(~m[751]&~m[754]&~m[755]&~m[756]&m[757])|(m[751]&~m[754]&~m[755]&~m[756]&m[757])|(m[751]&m[754]&~m[755]&~m[756]&m[757])|(m[751]&~m[754]&m[755]&~m[756]&m[757])|(~m[751]&~m[754]&~m[755]&m[756]&m[757])|(m[751]&~m[754]&~m[755]&m[756]&m[757])|(~m[751]&m[754]&~m[755]&m[756]&m[757])|(m[751]&m[754]&~m[755]&m[756]&m[757])|(~m[751]&~m[754]&m[755]&m[756]&m[757])|(m[751]&~m[754]&m[755]&m[756]&m[757])|(m[751]&m[754]&m[755]&m[756]&m[757]))):InitCond[285];
    m[758] = run?((((m[536]&~m[759]&~m[760]&~m[761]&~m[762])|(~m[536]&~m[759]&~m[760]&m[761]&~m[762])|(m[536]&m[759]&~m[760]&m[761]&~m[762])|(m[536]&~m[759]&m[760]&m[761]&~m[762])|(~m[536]&m[759]&~m[760]&~m[761]&m[762])|(~m[536]&~m[759]&m[760]&~m[761]&m[762])|(m[536]&m[759]&m[760]&~m[761]&m[762])|(~m[536]&m[759]&m[760]&m[761]&m[762]))&UnbiasedRNG[34])|((m[536]&~m[759]&~m[760]&m[761]&~m[762])|(~m[536]&~m[759]&~m[760]&~m[761]&m[762])|(m[536]&~m[759]&~m[760]&~m[761]&m[762])|(m[536]&m[759]&~m[760]&~m[761]&m[762])|(m[536]&~m[759]&m[760]&~m[761]&m[762])|(~m[536]&~m[759]&~m[760]&m[761]&m[762])|(m[536]&~m[759]&~m[760]&m[761]&m[762])|(~m[536]&m[759]&~m[760]&m[761]&m[762])|(m[536]&m[759]&~m[760]&m[761]&m[762])|(~m[536]&~m[759]&m[760]&m[761]&m[762])|(m[536]&~m[759]&m[760]&m[761]&m[762])|(m[536]&m[759]&m[760]&m[761]&m[762]))):InitCond[286];
    m[763] = run?((((m[761]&~m[764]&~m[765]&~m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&m[766]&~m[767])|(m[761]&m[764]&~m[765]&m[766]&~m[767])|(m[761]&~m[764]&m[765]&m[766]&~m[767])|(~m[761]&m[764]&~m[765]&~m[766]&m[767])|(~m[761]&~m[764]&m[765]&~m[766]&m[767])|(m[761]&m[764]&m[765]&~m[766]&m[767])|(~m[761]&m[764]&m[765]&m[766]&m[767]))&UnbiasedRNG[35])|((m[761]&~m[764]&~m[765]&m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&m[765]&~m[766]&m[767])|(~m[761]&~m[764]&~m[765]&m[766]&m[767])|(m[761]&~m[764]&~m[765]&m[766]&m[767])|(~m[761]&m[764]&~m[765]&m[766]&m[767])|(m[761]&m[764]&~m[765]&m[766]&m[767])|(~m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&m[764]&m[765]&m[766]&m[767]))):InitCond[287];
    m[768] = run?((((m[766]&~m[769]&~m[770]&~m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&m[771]&~m[772])|(m[766]&m[769]&~m[770]&m[771]&~m[772])|(m[766]&~m[769]&m[770]&m[771]&~m[772])|(~m[766]&m[769]&~m[770]&~m[771]&m[772])|(~m[766]&~m[769]&m[770]&~m[771]&m[772])|(m[766]&m[769]&m[770]&~m[771]&m[772])|(~m[766]&m[769]&m[770]&m[771]&m[772]))&UnbiasedRNG[36])|((m[766]&~m[769]&~m[770]&m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&m[770]&~m[771]&m[772])|(~m[766]&~m[769]&~m[770]&m[771]&m[772])|(m[766]&~m[769]&~m[770]&m[771]&m[772])|(~m[766]&m[769]&~m[770]&m[771]&m[772])|(m[766]&m[769]&~m[770]&m[771]&m[772])|(~m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&m[769]&m[770]&m[771]&m[772]))):InitCond[288];
    m[773] = run?((((m[771]&~m[774]&~m[775]&~m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&m[776]&~m[777])|(m[771]&m[774]&~m[775]&m[776]&~m[777])|(m[771]&~m[774]&m[775]&m[776]&~m[777])|(~m[771]&m[774]&~m[775]&~m[776]&m[777])|(~m[771]&~m[774]&m[775]&~m[776]&m[777])|(m[771]&m[774]&m[775]&~m[776]&m[777])|(~m[771]&m[774]&m[775]&m[776]&m[777]))&UnbiasedRNG[37])|((m[771]&~m[774]&~m[775]&m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&m[775]&~m[776]&m[777])|(~m[771]&~m[774]&~m[775]&m[776]&m[777])|(m[771]&~m[774]&~m[775]&m[776]&m[777])|(~m[771]&m[774]&~m[775]&m[776]&m[777])|(m[771]&m[774]&~m[775]&m[776]&m[777])|(~m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&m[774]&m[775]&m[776]&m[777]))):InitCond[289];
    m[778] = run?((((m[537]&~m[779]&~m[780]&~m[781]&~m[782])|(~m[537]&~m[779]&~m[780]&m[781]&~m[782])|(m[537]&m[779]&~m[780]&m[781]&~m[782])|(m[537]&~m[779]&m[780]&m[781]&~m[782])|(~m[537]&m[779]&~m[780]&~m[781]&m[782])|(~m[537]&~m[779]&m[780]&~m[781]&m[782])|(m[537]&m[779]&m[780]&~m[781]&m[782])|(~m[537]&m[779]&m[780]&m[781]&m[782]))&UnbiasedRNG[38])|((m[537]&~m[779]&~m[780]&m[781]&~m[782])|(~m[537]&~m[779]&~m[780]&~m[781]&m[782])|(m[537]&~m[779]&~m[780]&~m[781]&m[782])|(m[537]&m[779]&~m[780]&~m[781]&m[782])|(m[537]&~m[779]&m[780]&~m[781]&m[782])|(~m[537]&~m[779]&~m[780]&m[781]&m[782])|(m[537]&~m[779]&~m[780]&m[781]&m[782])|(~m[537]&m[779]&~m[780]&m[781]&m[782])|(m[537]&m[779]&~m[780]&m[781]&m[782])|(~m[537]&~m[779]&m[780]&m[781]&m[782])|(m[537]&~m[779]&m[780]&m[781]&m[782])|(m[537]&m[779]&m[780]&m[781]&m[782]))):InitCond[290];
    m[783] = run?((((m[781]&~m[784]&~m[785]&~m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&m[786]&~m[787])|(m[781]&m[784]&~m[785]&m[786]&~m[787])|(m[781]&~m[784]&m[785]&m[786]&~m[787])|(~m[781]&m[784]&~m[785]&~m[786]&m[787])|(~m[781]&~m[784]&m[785]&~m[786]&m[787])|(m[781]&m[784]&m[785]&~m[786]&m[787])|(~m[781]&m[784]&m[785]&m[786]&m[787]))&UnbiasedRNG[39])|((m[781]&~m[784]&~m[785]&m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&m[785]&~m[786]&m[787])|(~m[781]&~m[784]&~m[785]&m[786]&m[787])|(m[781]&~m[784]&~m[785]&m[786]&m[787])|(~m[781]&m[784]&~m[785]&m[786]&m[787])|(m[781]&m[784]&~m[785]&m[786]&m[787])|(~m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&m[784]&m[785]&m[786]&m[787]))):InitCond[291];
    m[788] = run?((((m[786]&~m[789]&~m[790]&~m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&m[791]&~m[792])|(m[786]&m[789]&~m[790]&m[791]&~m[792])|(m[786]&~m[789]&m[790]&m[791]&~m[792])|(~m[786]&m[789]&~m[790]&~m[791]&m[792])|(~m[786]&~m[789]&m[790]&~m[791]&m[792])|(m[786]&m[789]&m[790]&~m[791]&m[792])|(~m[786]&m[789]&m[790]&m[791]&m[792]))&UnbiasedRNG[40])|((m[786]&~m[789]&~m[790]&m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&m[790]&~m[791]&m[792])|(~m[786]&~m[789]&~m[790]&m[791]&m[792])|(m[786]&~m[789]&~m[790]&m[791]&m[792])|(~m[786]&m[789]&~m[790]&m[791]&m[792])|(m[786]&m[789]&~m[790]&m[791]&m[792])|(~m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&m[789]&m[790]&m[791]&m[792]))):InitCond[292];
    m[793] = run?((((m[791]&~m[794]&~m[795]&~m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&m[796]&~m[797])|(m[791]&m[794]&~m[795]&m[796]&~m[797])|(m[791]&~m[794]&m[795]&m[796]&~m[797])|(~m[791]&m[794]&~m[795]&~m[796]&m[797])|(~m[791]&~m[794]&m[795]&~m[796]&m[797])|(m[791]&m[794]&m[795]&~m[796]&m[797])|(~m[791]&m[794]&m[795]&m[796]&m[797]))&UnbiasedRNG[41])|((m[791]&~m[794]&~m[795]&m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&m[795]&~m[796]&m[797])|(~m[791]&~m[794]&~m[795]&m[796]&m[797])|(m[791]&~m[794]&~m[795]&m[796]&m[797])|(~m[791]&m[794]&~m[795]&m[796]&m[797])|(m[791]&m[794]&~m[795]&m[796]&m[797])|(~m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&m[794]&m[795]&m[796]&m[797]))):InitCond[293];
    m[798] = run?((((m[796]&~m[799]&~m[800]&~m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&m[801]&~m[802])|(m[796]&m[799]&~m[800]&m[801]&~m[802])|(m[796]&~m[799]&m[800]&m[801]&~m[802])|(~m[796]&m[799]&~m[800]&~m[801]&m[802])|(~m[796]&~m[799]&m[800]&~m[801]&m[802])|(m[796]&m[799]&m[800]&~m[801]&m[802])|(~m[796]&m[799]&m[800]&m[801]&m[802]))&UnbiasedRNG[42])|((m[796]&~m[799]&~m[800]&m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&m[800]&~m[801]&m[802])|(~m[796]&~m[799]&~m[800]&m[801]&m[802])|(m[796]&~m[799]&~m[800]&m[801]&m[802])|(~m[796]&m[799]&~m[800]&m[801]&m[802])|(m[796]&m[799]&~m[800]&m[801]&m[802])|(~m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&m[799]&m[800]&m[801]&m[802]))):InitCond[294];
    m[803] = run?((((m[538]&~m[804]&~m[805]&~m[806]&~m[807])|(~m[538]&~m[804]&~m[805]&m[806]&~m[807])|(m[538]&m[804]&~m[805]&m[806]&~m[807])|(m[538]&~m[804]&m[805]&m[806]&~m[807])|(~m[538]&m[804]&~m[805]&~m[806]&m[807])|(~m[538]&~m[804]&m[805]&~m[806]&m[807])|(m[538]&m[804]&m[805]&~m[806]&m[807])|(~m[538]&m[804]&m[805]&m[806]&m[807]))&UnbiasedRNG[43])|((m[538]&~m[804]&~m[805]&m[806]&~m[807])|(~m[538]&~m[804]&~m[805]&~m[806]&m[807])|(m[538]&~m[804]&~m[805]&~m[806]&m[807])|(m[538]&m[804]&~m[805]&~m[806]&m[807])|(m[538]&~m[804]&m[805]&~m[806]&m[807])|(~m[538]&~m[804]&~m[805]&m[806]&m[807])|(m[538]&~m[804]&~m[805]&m[806]&m[807])|(~m[538]&m[804]&~m[805]&m[806]&m[807])|(m[538]&m[804]&~m[805]&m[806]&m[807])|(~m[538]&~m[804]&m[805]&m[806]&m[807])|(m[538]&~m[804]&m[805]&m[806]&m[807])|(m[538]&m[804]&m[805]&m[806]&m[807]))):InitCond[295];
    m[808] = run?((((m[806]&~m[809]&~m[810]&~m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&m[811]&~m[812])|(m[806]&m[809]&~m[810]&m[811]&~m[812])|(m[806]&~m[809]&m[810]&m[811]&~m[812])|(~m[806]&m[809]&~m[810]&~m[811]&m[812])|(~m[806]&~m[809]&m[810]&~m[811]&m[812])|(m[806]&m[809]&m[810]&~m[811]&m[812])|(~m[806]&m[809]&m[810]&m[811]&m[812]))&UnbiasedRNG[44])|((m[806]&~m[809]&~m[810]&m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&m[810]&~m[811]&m[812])|(~m[806]&~m[809]&~m[810]&m[811]&m[812])|(m[806]&~m[809]&~m[810]&m[811]&m[812])|(~m[806]&m[809]&~m[810]&m[811]&m[812])|(m[806]&m[809]&~m[810]&m[811]&m[812])|(~m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&m[809]&m[810]&m[811]&m[812]))):InitCond[296];
    m[813] = run?((((m[811]&~m[814]&~m[815]&~m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&m[816]&~m[817])|(m[811]&m[814]&~m[815]&m[816]&~m[817])|(m[811]&~m[814]&m[815]&m[816]&~m[817])|(~m[811]&m[814]&~m[815]&~m[816]&m[817])|(~m[811]&~m[814]&m[815]&~m[816]&m[817])|(m[811]&m[814]&m[815]&~m[816]&m[817])|(~m[811]&m[814]&m[815]&m[816]&m[817]))&UnbiasedRNG[45])|((m[811]&~m[814]&~m[815]&m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&m[815]&~m[816]&m[817])|(~m[811]&~m[814]&~m[815]&m[816]&m[817])|(m[811]&~m[814]&~m[815]&m[816]&m[817])|(~m[811]&m[814]&~m[815]&m[816]&m[817])|(m[811]&m[814]&~m[815]&m[816]&m[817])|(~m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&m[814]&m[815]&m[816]&m[817]))):InitCond[297];
    m[818] = run?((((m[816]&~m[819]&~m[820]&~m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&m[821]&~m[822])|(m[816]&m[819]&~m[820]&m[821]&~m[822])|(m[816]&~m[819]&m[820]&m[821]&~m[822])|(~m[816]&m[819]&~m[820]&~m[821]&m[822])|(~m[816]&~m[819]&m[820]&~m[821]&m[822])|(m[816]&m[819]&m[820]&~m[821]&m[822])|(~m[816]&m[819]&m[820]&m[821]&m[822]))&UnbiasedRNG[46])|((m[816]&~m[819]&~m[820]&m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&m[820]&~m[821]&m[822])|(~m[816]&~m[819]&~m[820]&m[821]&m[822])|(m[816]&~m[819]&~m[820]&m[821]&m[822])|(~m[816]&m[819]&~m[820]&m[821]&m[822])|(m[816]&m[819]&~m[820]&m[821]&m[822])|(~m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&m[819]&m[820]&m[821]&m[822]))):InitCond[298];
    m[823] = run?((((m[821]&~m[824]&~m[825]&~m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&m[826]&~m[827])|(m[821]&m[824]&~m[825]&m[826]&~m[827])|(m[821]&~m[824]&m[825]&m[826]&~m[827])|(~m[821]&m[824]&~m[825]&~m[826]&m[827])|(~m[821]&~m[824]&m[825]&~m[826]&m[827])|(m[821]&m[824]&m[825]&~m[826]&m[827])|(~m[821]&m[824]&m[825]&m[826]&m[827]))&UnbiasedRNG[47])|((m[821]&~m[824]&~m[825]&m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&m[825]&~m[826]&m[827])|(~m[821]&~m[824]&~m[825]&m[826]&m[827])|(m[821]&~m[824]&~m[825]&m[826]&m[827])|(~m[821]&m[824]&~m[825]&m[826]&m[827])|(m[821]&m[824]&~m[825]&m[826]&m[827])|(~m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&m[824]&m[825]&m[826]&m[827]))):InitCond[299];
    m[828] = run?((((m[826]&~m[829]&~m[830]&~m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&m[831]&~m[832])|(m[826]&m[829]&~m[830]&m[831]&~m[832])|(m[826]&~m[829]&m[830]&m[831]&~m[832])|(~m[826]&m[829]&~m[830]&~m[831]&m[832])|(~m[826]&~m[829]&m[830]&~m[831]&m[832])|(m[826]&m[829]&m[830]&~m[831]&m[832])|(~m[826]&m[829]&m[830]&m[831]&m[832]))&UnbiasedRNG[48])|((m[826]&~m[829]&~m[830]&m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&m[830]&~m[831]&m[832])|(~m[826]&~m[829]&~m[830]&m[831]&m[832])|(m[826]&~m[829]&~m[830]&m[831]&m[832])|(~m[826]&m[829]&~m[830]&m[831]&m[832])|(m[826]&m[829]&~m[830]&m[831]&m[832])|(~m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&m[829]&m[830]&m[831]&m[832]))):InitCond[300];
    m[833] = run?((((m[539]&~m[834]&~m[835]&~m[836]&~m[837])|(~m[539]&~m[834]&~m[835]&m[836]&~m[837])|(m[539]&m[834]&~m[835]&m[836]&~m[837])|(m[539]&~m[834]&m[835]&m[836]&~m[837])|(~m[539]&m[834]&~m[835]&~m[836]&m[837])|(~m[539]&~m[834]&m[835]&~m[836]&m[837])|(m[539]&m[834]&m[835]&~m[836]&m[837])|(~m[539]&m[834]&m[835]&m[836]&m[837]))&UnbiasedRNG[49])|((m[539]&~m[834]&~m[835]&m[836]&~m[837])|(~m[539]&~m[834]&~m[835]&~m[836]&m[837])|(m[539]&~m[834]&~m[835]&~m[836]&m[837])|(m[539]&m[834]&~m[835]&~m[836]&m[837])|(m[539]&~m[834]&m[835]&~m[836]&m[837])|(~m[539]&~m[834]&~m[835]&m[836]&m[837])|(m[539]&~m[834]&~m[835]&m[836]&m[837])|(~m[539]&m[834]&~m[835]&m[836]&m[837])|(m[539]&m[834]&~m[835]&m[836]&m[837])|(~m[539]&~m[834]&m[835]&m[836]&m[837])|(m[539]&~m[834]&m[835]&m[836]&m[837])|(m[539]&m[834]&m[835]&m[836]&m[837]))):InitCond[301];
    m[838] = run?((((m[836]&~m[839]&~m[840]&~m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&m[841]&~m[842])|(m[836]&m[839]&~m[840]&m[841]&~m[842])|(m[836]&~m[839]&m[840]&m[841]&~m[842])|(~m[836]&m[839]&~m[840]&~m[841]&m[842])|(~m[836]&~m[839]&m[840]&~m[841]&m[842])|(m[836]&m[839]&m[840]&~m[841]&m[842])|(~m[836]&m[839]&m[840]&m[841]&m[842]))&UnbiasedRNG[50])|((m[836]&~m[839]&~m[840]&m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&m[840]&~m[841]&m[842])|(~m[836]&~m[839]&~m[840]&m[841]&m[842])|(m[836]&~m[839]&~m[840]&m[841]&m[842])|(~m[836]&m[839]&~m[840]&m[841]&m[842])|(m[836]&m[839]&~m[840]&m[841]&m[842])|(~m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&m[839]&m[840]&m[841]&m[842]))):InitCond[302];
    m[843] = run?((((m[841]&~m[844]&~m[845]&~m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&m[846]&~m[847])|(m[841]&m[844]&~m[845]&m[846]&~m[847])|(m[841]&~m[844]&m[845]&m[846]&~m[847])|(~m[841]&m[844]&~m[845]&~m[846]&m[847])|(~m[841]&~m[844]&m[845]&~m[846]&m[847])|(m[841]&m[844]&m[845]&~m[846]&m[847])|(~m[841]&m[844]&m[845]&m[846]&m[847]))&UnbiasedRNG[51])|((m[841]&~m[844]&~m[845]&m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&m[845]&~m[846]&m[847])|(~m[841]&~m[844]&~m[845]&m[846]&m[847])|(m[841]&~m[844]&~m[845]&m[846]&m[847])|(~m[841]&m[844]&~m[845]&m[846]&m[847])|(m[841]&m[844]&~m[845]&m[846]&m[847])|(~m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&m[844]&m[845]&m[846]&m[847]))):InitCond[303];
    m[848] = run?((((m[846]&~m[849]&~m[850]&~m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&m[851]&~m[852])|(m[846]&m[849]&~m[850]&m[851]&~m[852])|(m[846]&~m[849]&m[850]&m[851]&~m[852])|(~m[846]&m[849]&~m[850]&~m[851]&m[852])|(~m[846]&~m[849]&m[850]&~m[851]&m[852])|(m[846]&m[849]&m[850]&~m[851]&m[852])|(~m[846]&m[849]&m[850]&m[851]&m[852]))&UnbiasedRNG[52])|((m[846]&~m[849]&~m[850]&m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&m[850]&~m[851]&m[852])|(~m[846]&~m[849]&~m[850]&m[851]&m[852])|(m[846]&~m[849]&~m[850]&m[851]&m[852])|(~m[846]&m[849]&~m[850]&m[851]&m[852])|(m[846]&m[849]&~m[850]&m[851]&m[852])|(~m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&m[849]&m[850]&m[851]&m[852]))):InitCond[304];
    m[853] = run?((((m[851]&~m[854]&~m[855]&~m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&m[856]&~m[857])|(m[851]&m[854]&~m[855]&m[856]&~m[857])|(m[851]&~m[854]&m[855]&m[856]&~m[857])|(~m[851]&m[854]&~m[855]&~m[856]&m[857])|(~m[851]&~m[854]&m[855]&~m[856]&m[857])|(m[851]&m[854]&m[855]&~m[856]&m[857])|(~m[851]&m[854]&m[855]&m[856]&m[857]))&UnbiasedRNG[53])|((m[851]&~m[854]&~m[855]&m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&m[855]&~m[856]&m[857])|(~m[851]&~m[854]&~m[855]&m[856]&m[857])|(m[851]&~m[854]&~m[855]&m[856]&m[857])|(~m[851]&m[854]&~m[855]&m[856]&m[857])|(m[851]&m[854]&~m[855]&m[856]&m[857])|(~m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&m[854]&m[855]&m[856]&m[857]))):InitCond[305];
    m[858] = run?((((m[856]&~m[859]&~m[860]&~m[861]&~m[862])|(~m[856]&~m[859]&~m[860]&m[861]&~m[862])|(m[856]&m[859]&~m[860]&m[861]&~m[862])|(m[856]&~m[859]&m[860]&m[861]&~m[862])|(~m[856]&m[859]&~m[860]&~m[861]&m[862])|(~m[856]&~m[859]&m[860]&~m[861]&m[862])|(m[856]&m[859]&m[860]&~m[861]&m[862])|(~m[856]&m[859]&m[860]&m[861]&m[862]))&UnbiasedRNG[54])|((m[856]&~m[859]&~m[860]&m[861]&~m[862])|(~m[856]&~m[859]&~m[860]&~m[861]&m[862])|(m[856]&~m[859]&~m[860]&~m[861]&m[862])|(m[856]&m[859]&~m[860]&~m[861]&m[862])|(m[856]&~m[859]&m[860]&~m[861]&m[862])|(~m[856]&~m[859]&~m[860]&m[861]&m[862])|(m[856]&~m[859]&~m[860]&m[861]&m[862])|(~m[856]&m[859]&~m[860]&m[861]&m[862])|(m[856]&m[859]&~m[860]&m[861]&m[862])|(~m[856]&~m[859]&m[860]&m[861]&m[862])|(m[856]&~m[859]&m[860]&m[861]&m[862])|(m[856]&m[859]&m[860]&m[861]&m[862]))):InitCond[306];
    m[863] = run?((((m[861]&~m[864]&~m[865]&~m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&m[866]&~m[867])|(m[861]&m[864]&~m[865]&m[866]&~m[867])|(m[861]&~m[864]&m[865]&m[866]&~m[867])|(~m[861]&m[864]&~m[865]&~m[866]&m[867])|(~m[861]&~m[864]&m[865]&~m[866]&m[867])|(m[861]&m[864]&m[865]&~m[866]&m[867])|(~m[861]&m[864]&m[865]&m[866]&m[867]))&UnbiasedRNG[55])|((m[861]&~m[864]&~m[865]&m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&m[865]&~m[866]&m[867])|(~m[861]&~m[864]&~m[865]&m[866]&m[867])|(m[861]&~m[864]&~m[865]&m[866]&m[867])|(~m[861]&m[864]&~m[865]&m[866]&m[867])|(m[861]&m[864]&~m[865]&m[866]&m[867])|(~m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&m[864]&m[865]&m[866]&m[867]))):InitCond[307];
    m[868] = run?((((m[540]&~m[869]&~m[870]&~m[871]&~m[872])|(~m[540]&~m[869]&~m[870]&m[871]&~m[872])|(m[540]&m[869]&~m[870]&m[871]&~m[872])|(m[540]&~m[869]&m[870]&m[871]&~m[872])|(~m[540]&m[869]&~m[870]&~m[871]&m[872])|(~m[540]&~m[869]&m[870]&~m[871]&m[872])|(m[540]&m[869]&m[870]&~m[871]&m[872])|(~m[540]&m[869]&m[870]&m[871]&m[872]))&UnbiasedRNG[56])|((m[540]&~m[869]&~m[870]&m[871]&~m[872])|(~m[540]&~m[869]&~m[870]&~m[871]&m[872])|(m[540]&~m[869]&~m[870]&~m[871]&m[872])|(m[540]&m[869]&~m[870]&~m[871]&m[872])|(m[540]&~m[869]&m[870]&~m[871]&m[872])|(~m[540]&~m[869]&~m[870]&m[871]&m[872])|(m[540]&~m[869]&~m[870]&m[871]&m[872])|(~m[540]&m[869]&~m[870]&m[871]&m[872])|(m[540]&m[869]&~m[870]&m[871]&m[872])|(~m[540]&~m[869]&m[870]&m[871]&m[872])|(m[540]&~m[869]&m[870]&m[871]&m[872])|(m[540]&m[869]&m[870]&m[871]&m[872]))):InitCond[308];
    m[873] = run?((((m[871]&~m[874]&~m[875]&~m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&m[876]&~m[877])|(m[871]&m[874]&~m[875]&m[876]&~m[877])|(m[871]&~m[874]&m[875]&m[876]&~m[877])|(~m[871]&m[874]&~m[875]&~m[876]&m[877])|(~m[871]&~m[874]&m[875]&~m[876]&m[877])|(m[871]&m[874]&m[875]&~m[876]&m[877])|(~m[871]&m[874]&m[875]&m[876]&m[877]))&UnbiasedRNG[57])|((m[871]&~m[874]&~m[875]&m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&m[875]&~m[876]&m[877])|(~m[871]&~m[874]&~m[875]&m[876]&m[877])|(m[871]&~m[874]&~m[875]&m[876]&m[877])|(~m[871]&m[874]&~m[875]&m[876]&m[877])|(m[871]&m[874]&~m[875]&m[876]&m[877])|(~m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&m[874]&m[875]&m[876]&m[877]))):InitCond[309];
    m[878] = run?((((m[876]&~m[879]&~m[880]&~m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&m[881]&~m[882])|(m[876]&m[879]&~m[880]&m[881]&~m[882])|(m[876]&~m[879]&m[880]&m[881]&~m[882])|(~m[876]&m[879]&~m[880]&~m[881]&m[882])|(~m[876]&~m[879]&m[880]&~m[881]&m[882])|(m[876]&m[879]&m[880]&~m[881]&m[882])|(~m[876]&m[879]&m[880]&m[881]&m[882]))&UnbiasedRNG[58])|((m[876]&~m[879]&~m[880]&m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&m[880]&~m[881]&m[882])|(~m[876]&~m[879]&~m[880]&m[881]&m[882])|(m[876]&~m[879]&~m[880]&m[881]&m[882])|(~m[876]&m[879]&~m[880]&m[881]&m[882])|(m[876]&m[879]&~m[880]&m[881]&m[882])|(~m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&m[879]&m[880]&m[881]&m[882]))):InitCond[310];
    m[883] = run?((((m[881]&~m[884]&~m[885]&~m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&m[886]&~m[887])|(m[881]&m[884]&~m[885]&m[886]&~m[887])|(m[881]&~m[884]&m[885]&m[886]&~m[887])|(~m[881]&m[884]&~m[885]&~m[886]&m[887])|(~m[881]&~m[884]&m[885]&~m[886]&m[887])|(m[881]&m[884]&m[885]&~m[886]&m[887])|(~m[881]&m[884]&m[885]&m[886]&m[887]))&UnbiasedRNG[59])|((m[881]&~m[884]&~m[885]&m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&m[885]&~m[886]&m[887])|(~m[881]&~m[884]&~m[885]&m[886]&m[887])|(m[881]&~m[884]&~m[885]&m[886]&m[887])|(~m[881]&m[884]&~m[885]&m[886]&m[887])|(m[881]&m[884]&~m[885]&m[886]&m[887])|(~m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&m[884]&m[885]&m[886]&m[887]))):InitCond[311];
    m[888] = run?((((m[886]&~m[889]&~m[890]&~m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&m[891]&~m[892])|(m[886]&m[889]&~m[890]&m[891]&~m[892])|(m[886]&~m[889]&m[890]&m[891]&~m[892])|(~m[886]&m[889]&~m[890]&~m[891]&m[892])|(~m[886]&~m[889]&m[890]&~m[891]&m[892])|(m[886]&m[889]&m[890]&~m[891]&m[892])|(~m[886]&m[889]&m[890]&m[891]&m[892]))&UnbiasedRNG[60])|((m[886]&~m[889]&~m[890]&m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&m[890]&~m[891]&m[892])|(~m[886]&~m[889]&~m[890]&m[891]&m[892])|(m[886]&~m[889]&~m[890]&m[891]&m[892])|(~m[886]&m[889]&~m[890]&m[891]&m[892])|(m[886]&m[889]&~m[890]&m[891]&m[892])|(~m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&m[889]&m[890]&m[891]&m[892]))):InitCond[312];
    m[893] = run?((((m[891]&~m[894]&~m[895]&~m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&m[896]&~m[897])|(m[891]&m[894]&~m[895]&m[896]&~m[897])|(m[891]&~m[894]&m[895]&m[896]&~m[897])|(~m[891]&m[894]&~m[895]&~m[896]&m[897])|(~m[891]&~m[894]&m[895]&~m[896]&m[897])|(m[891]&m[894]&m[895]&~m[896]&m[897])|(~m[891]&m[894]&m[895]&m[896]&m[897]))&UnbiasedRNG[61])|((m[891]&~m[894]&~m[895]&m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&m[895]&~m[896]&m[897])|(~m[891]&~m[894]&~m[895]&m[896]&m[897])|(m[891]&~m[894]&~m[895]&m[896]&m[897])|(~m[891]&m[894]&~m[895]&m[896]&m[897])|(m[891]&m[894]&~m[895]&m[896]&m[897])|(~m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&m[894]&m[895]&m[896]&m[897]))):InitCond[313];
    m[898] = run?((((m[896]&~m[899]&~m[900]&~m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&m[901]&~m[902])|(m[896]&m[899]&~m[900]&m[901]&~m[902])|(m[896]&~m[899]&m[900]&m[901]&~m[902])|(~m[896]&m[899]&~m[900]&~m[901]&m[902])|(~m[896]&~m[899]&m[900]&~m[901]&m[902])|(m[896]&m[899]&m[900]&~m[901]&m[902])|(~m[896]&m[899]&m[900]&m[901]&m[902]))&UnbiasedRNG[62])|((m[896]&~m[899]&~m[900]&m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&m[900]&~m[901]&m[902])|(~m[896]&~m[899]&~m[900]&m[901]&m[902])|(m[896]&~m[899]&~m[900]&m[901]&m[902])|(~m[896]&m[899]&~m[900]&m[901]&m[902])|(m[896]&m[899]&~m[900]&m[901]&m[902])|(~m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&m[899]&m[900]&m[901]&m[902]))):InitCond[314];
    m[903] = run?((((m[901]&~m[904]&~m[905]&~m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&m[906]&~m[907])|(m[901]&m[904]&~m[905]&m[906]&~m[907])|(m[901]&~m[904]&m[905]&m[906]&~m[907])|(~m[901]&m[904]&~m[905]&~m[906]&m[907])|(~m[901]&~m[904]&m[905]&~m[906]&m[907])|(m[901]&m[904]&m[905]&~m[906]&m[907])|(~m[901]&m[904]&m[905]&m[906]&m[907]))&UnbiasedRNG[63])|((m[901]&~m[904]&~m[905]&m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&m[905]&~m[906]&m[907])|(~m[901]&~m[904]&~m[905]&m[906]&m[907])|(m[901]&~m[904]&~m[905]&m[906]&m[907])|(~m[901]&m[904]&~m[905]&m[906]&m[907])|(m[901]&m[904]&~m[905]&m[906]&m[907])|(~m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&m[904]&m[905]&m[906]&m[907]))):InitCond[315];
    m[908] = run?((((m[541]&~m[909]&~m[910]&~m[911]&~m[912])|(~m[541]&~m[909]&~m[910]&m[911]&~m[912])|(m[541]&m[909]&~m[910]&m[911]&~m[912])|(m[541]&~m[909]&m[910]&m[911]&~m[912])|(~m[541]&m[909]&~m[910]&~m[911]&m[912])|(~m[541]&~m[909]&m[910]&~m[911]&m[912])|(m[541]&m[909]&m[910]&~m[911]&m[912])|(~m[541]&m[909]&m[910]&m[911]&m[912]))&UnbiasedRNG[64])|((m[541]&~m[909]&~m[910]&m[911]&~m[912])|(~m[541]&~m[909]&~m[910]&~m[911]&m[912])|(m[541]&~m[909]&~m[910]&~m[911]&m[912])|(m[541]&m[909]&~m[910]&~m[911]&m[912])|(m[541]&~m[909]&m[910]&~m[911]&m[912])|(~m[541]&~m[909]&~m[910]&m[911]&m[912])|(m[541]&~m[909]&~m[910]&m[911]&m[912])|(~m[541]&m[909]&~m[910]&m[911]&m[912])|(m[541]&m[909]&~m[910]&m[911]&m[912])|(~m[541]&~m[909]&m[910]&m[911]&m[912])|(m[541]&~m[909]&m[910]&m[911]&m[912])|(m[541]&m[909]&m[910]&m[911]&m[912]))):InitCond[316];
    m[913] = run?((((m[911]&~m[914]&~m[915]&~m[916]&~m[917])|(~m[911]&~m[914]&~m[915]&m[916]&~m[917])|(m[911]&m[914]&~m[915]&m[916]&~m[917])|(m[911]&~m[914]&m[915]&m[916]&~m[917])|(~m[911]&m[914]&~m[915]&~m[916]&m[917])|(~m[911]&~m[914]&m[915]&~m[916]&m[917])|(m[911]&m[914]&m[915]&~m[916]&m[917])|(~m[911]&m[914]&m[915]&m[916]&m[917]))&UnbiasedRNG[65])|((m[911]&~m[914]&~m[915]&m[916]&~m[917])|(~m[911]&~m[914]&~m[915]&~m[916]&m[917])|(m[911]&~m[914]&~m[915]&~m[916]&m[917])|(m[911]&m[914]&~m[915]&~m[916]&m[917])|(m[911]&~m[914]&m[915]&~m[916]&m[917])|(~m[911]&~m[914]&~m[915]&m[916]&m[917])|(m[911]&~m[914]&~m[915]&m[916]&m[917])|(~m[911]&m[914]&~m[915]&m[916]&m[917])|(m[911]&m[914]&~m[915]&m[916]&m[917])|(~m[911]&~m[914]&m[915]&m[916]&m[917])|(m[911]&~m[914]&m[915]&m[916]&m[917])|(m[911]&m[914]&m[915]&m[916]&m[917]))):InitCond[317];
    m[918] = run?((((m[916]&~m[919]&~m[920]&~m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&m[921]&~m[922])|(m[916]&m[919]&~m[920]&m[921]&~m[922])|(m[916]&~m[919]&m[920]&m[921]&~m[922])|(~m[916]&m[919]&~m[920]&~m[921]&m[922])|(~m[916]&~m[919]&m[920]&~m[921]&m[922])|(m[916]&m[919]&m[920]&~m[921]&m[922])|(~m[916]&m[919]&m[920]&m[921]&m[922]))&UnbiasedRNG[66])|((m[916]&~m[919]&~m[920]&m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&m[920]&~m[921]&m[922])|(~m[916]&~m[919]&~m[920]&m[921]&m[922])|(m[916]&~m[919]&~m[920]&m[921]&m[922])|(~m[916]&m[919]&~m[920]&m[921]&m[922])|(m[916]&m[919]&~m[920]&m[921]&m[922])|(~m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&m[919]&m[920]&m[921]&m[922]))):InitCond[318];
    m[923] = run?((((m[921]&~m[924]&~m[925]&~m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&m[926]&~m[927])|(m[921]&m[924]&~m[925]&m[926]&~m[927])|(m[921]&~m[924]&m[925]&m[926]&~m[927])|(~m[921]&m[924]&~m[925]&~m[926]&m[927])|(~m[921]&~m[924]&m[925]&~m[926]&m[927])|(m[921]&m[924]&m[925]&~m[926]&m[927])|(~m[921]&m[924]&m[925]&m[926]&m[927]))&UnbiasedRNG[67])|((m[921]&~m[924]&~m[925]&m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&m[925]&~m[926]&m[927])|(~m[921]&~m[924]&~m[925]&m[926]&m[927])|(m[921]&~m[924]&~m[925]&m[926]&m[927])|(~m[921]&m[924]&~m[925]&m[926]&m[927])|(m[921]&m[924]&~m[925]&m[926]&m[927])|(~m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&m[924]&m[925]&m[926]&m[927]))):InitCond[319];
    m[928] = run?((((m[926]&~m[929]&~m[930]&~m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&m[931]&~m[932])|(m[926]&m[929]&~m[930]&m[931]&~m[932])|(m[926]&~m[929]&m[930]&m[931]&~m[932])|(~m[926]&m[929]&~m[930]&~m[931]&m[932])|(~m[926]&~m[929]&m[930]&~m[931]&m[932])|(m[926]&m[929]&m[930]&~m[931]&m[932])|(~m[926]&m[929]&m[930]&m[931]&m[932]))&UnbiasedRNG[68])|((m[926]&~m[929]&~m[930]&m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&m[930]&~m[931]&m[932])|(~m[926]&~m[929]&~m[930]&m[931]&m[932])|(m[926]&~m[929]&~m[930]&m[931]&m[932])|(~m[926]&m[929]&~m[930]&m[931]&m[932])|(m[926]&m[929]&~m[930]&m[931]&m[932])|(~m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&m[929]&m[930]&m[931]&m[932]))):InitCond[320];
    m[933] = run?((((m[931]&~m[934]&~m[935]&~m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&m[936]&~m[937])|(m[931]&m[934]&~m[935]&m[936]&~m[937])|(m[931]&~m[934]&m[935]&m[936]&~m[937])|(~m[931]&m[934]&~m[935]&~m[936]&m[937])|(~m[931]&~m[934]&m[935]&~m[936]&m[937])|(m[931]&m[934]&m[935]&~m[936]&m[937])|(~m[931]&m[934]&m[935]&m[936]&m[937]))&UnbiasedRNG[69])|((m[931]&~m[934]&~m[935]&m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&m[935]&~m[936]&m[937])|(~m[931]&~m[934]&~m[935]&m[936]&m[937])|(m[931]&~m[934]&~m[935]&m[936]&m[937])|(~m[931]&m[934]&~m[935]&m[936]&m[937])|(m[931]&m[934]&~m[935]&m[936]&m[937])|(~m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&m[934]&m[935]&m[936]&m[937]))):InitCond[321];
    m[938] = run?((((m[936]&~m[939]&~m[940]&~m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&m[941]&~m[942])|(m[936]&m[939]&~m[940]&m[941]&~m[942])|(m[936]&~m[939]&m[940]&m[941]&~m[942])|(~m[936]&m[939]&~m[940]&~m[941]&m[942])|(~m[936]&~m[939]&m[940]&~m[941]&m[942])|(m[936]&m[939]&m[940]&~m[941]&m[942])|(~m[936]&m[939]&m[940]&m[941]&m[942]))&UnbiasedRNG[70])|((m[936]&~m[939]&~m[940]&m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&m[940]&~m[941]&m[942])|(~m[936]&~m[939]&~m[940]&m[941]&m[942])|(m[936]&~m[939]&~m[940]&m[941]&m[942])|(~m[936]&m[939]&~m[940]&m[941]&m[942])|(m[936]&m[939]&~m[940]&m[941]&m[942])|(~m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&m[939]&m[940]&m[941]&m[942]))):InitCond[322];
    m[943] = run?((((m[941]&~m[944]&~m[945]&~m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&m[946]&~m[947])|(m[941]&m[944]&~m[945]&m[946]&~m[947])|(m[941]&~m[944]&m[945]&m[946]&~m[947])|(~m[941]&m[944]&~m[945]&~m[946]&m[947])|(~m[941]&~m[944]&m[945]&~m[946]&m[947])|(m[941]&m[944]&m[945]&~m[946]&m[947])|(~m[941]&m[944]&m[945]&m[946]&m[947]))&UnbiasedRNG[71])|((m[941]&~m[944]&~m[945]&m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&m[945]&~m[946]&m[947])|(~m[941]&~m[944]&~m[945]&m[946]&m[947])|(m[941]&~m[944]&~m[945]&m[946]&m[947])|(~m[941]&m[944]&~m[945]&m[946]&m[947])|(m[941]&m[944]&~m[945]&m[946]&m[947])|(~m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&m[944]&m[945]&m[946]&m[947]))):InitCond[323];
    m[948] = run?((((m[946]&~m[949]&~m[950]&~m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&m[951]&~m[952])|(m[946]&m[949]&~m[950]&m[951]&~m[952])|(m[946]&~m[949]&m[950]&m[951]&~m[952])|(~m[946]&m[949]&~m[950]&~m[951]&m[952])|(~m[946]&~m[949]&m[950]&~m[951]&m[952])|(m[946]&m[949]&m[950]&~m[951]&m[952])|(~m[946]&m[949]&m[950]&m[951]&m[952]))&UnbiasedRNG[72])|((m[946]&~m[949]&~m[950]&m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&m[950]&~m[951]&m[952])|(~m[946]&~m[949]&~m[950]&m[951]&m[952])|(m[946]&~m[949]&~m[950]&m[951]&m[952])|(~m[946]&m[949]&~m[950]&m[951]&m[952])|(m[946]&m[949]&~m[950]&m[951]&m[952])|(~m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&m[949]&m[950]&m[951]&m[952]))):InitCond[324];
    m[953] = run?((((m[542]&~m[954]&~m[955]&~m[956]&~m[957])|(~m[542]&~m[954]&~m[955]&m[956]&~m[957])|(m[542]&m[954]&~m[955]&m[956]&~m[957])|(m[542]&~m[954]&m[955]&m[956]&~m[957])|(~m[542]&m[954]&~m[955]&~m[956]&m[957])|(~m[542]&~m[954]&m[955]&~m[956]&m[957])|(m[542]&m[954]&m[955]&~m[956]&m[957])|(~m[542]&m[954]&m[955]&m[956]&m[957]))&UnbiasedRNG[73])|((m[542]&~m[954]&~m[955]&m[956]&~m[957])|(~m[542]&~m[954]&~m[955]&~m[956]&m[957])|(m[542]&~m[954]&~m[955]&~m[956]&m[957])|(m[542]&m[954]&~m[955]&~m[956]&m[957])|(m[542]&~m[954]&m[955]&~m[956]&m[957])|(~m[542]&~m[954]&~m[955]&m[956]&m[957])|(m[542]&~m[954]&~m[955]&m[956]&m[957])|(~m[542]&m[954]&~m[955]&m[956]&m[957])|(m[542]&m[954]&~m[955]&m[956]&m[957])|(~m[542]&~m[954]&m[955]&m[956]&m[957])|(m[542]&~m[954]&m[955]&m[956]&m[957])|(m[542]&m[954]&m[955]&m[956]&m[957]))):InitCond[325];
    m[958] = run?((((m[956]&~m[959]&~m[960]&~m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&m[961]&~m[962])|(m[956]&m[959]&~m[960]&m[961]&~m[962])|(m[956]&~m[959]&m[960]&m[961]&~m[962])|(~m[956]&m[959]&~m[960]&~m[961]&m[962])|(~m[956]&~m[959]&m[960]&~m[961]&m[962])|(m[956]&m[959]&m[960]&~m[961]&m[962])|(~m[956]&m[959]&m[960]&m[961]&m[962]))&UnbiasedRNG[74])|((m[956]&~m[959]&~m[960]&m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&m[960]&~m[961]&m[962])|(~m[956]&~m[959]&~m[960]&m[961]&m[962])|(m[956]&~m[959]&~m[960]&m[961]&m[962])|(~m[956]&m[959]&~m[960]&m[961]&m[962])|(m[956]&m[959]&~m[960]&m[961]&m[962])|(~m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&m[959]&m[960]&m[961]&m[962]))):InitCond[326];
    m[963] = run?((((m[961]&~m[964]&~m[965]&~m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&m[966]&~m[967])|(m[961]&m[964]&~m[965]&m[966]&~m[967])|(m[961]&~m[964]&m[965]&m[966]&~m[967])|(~m[961]&m[964]&~m[965]&~m[966]&m[967])|(~m[961]&~m[964]&m[965]&~m[966]&m[967])|(m[961]&m[964]&m[965]&~m[966]&m[967])|(~m[961]&m[964]&m[965]&m[966]&m[967]))&UnbiasedRNG[75])|((m[961]&~m[964]&~m[965]&m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&m[965]&~m[966]&m[967])|(~m[961]&~m[964]&~m[965]&m[966]&m[967])|(m[961]&~m[964]&~m[965]&m[966]&m[967])|(~m[961]&m[964]&~m[965]&m[966]&m[967])|(m[961]&m[964]&~m[965]&m[966]&m[967])|(~m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&m[964]&m[965]&m[966]&m[967]))):InitCond[327];
    m[968] = run?((((m[966]&~m[969]&~m[970]&~m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&m[971]&~m[972])|(m[966]&m[969]&~m[970]&m[971]&~m[972])|(m[966]&~m[969]&m[970]&m[971]&~m[972])|(~m[966]&m[969]&~m[970]&~m[971]&m[972])|(~m[966]&~m[969]&m[970]&~m[971]&m[972])|(m[966]&m[969]&m[970]&~m[971]&m[972])|(~m[966]&m[969]&m[970]&m[971]&m[972]))&UnbiasedRNG[76])|((m[966]&~m[969]&~m[970]&m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&m[970]&~m[971]&m[972])|(~m[966]&~m[969]&~m[970]&m[971]&m[972])|(m[966]&~m[969]&~m[970]&m[971]&m[972])|(~m[966]&m[969]&~m[970]&m[971]&m[972])|(m[966]&m[969]&~m[970]&m[971]&m[972])|(~m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&m[969]&m[970]&m[971]&m[972]))):InitCond[328];
    m[973] = run?((((m[971]&~m[974]&~m[975]&~m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&m[976]&~m[977])|(m[971]&m[974]&~m[975]&m[976]&~m[977])|(m[971]&~m[974]&m[975]&m[976]&~m[977])|(~m[971]&m[974]&~m[975]&~m[976]&m[977])|(~m[971]&~m[974]&m[975]&~m[976]&m[977])|(m[971]&m[974]&m[975]&~m[976]&m[977])|(~m[971]&m[974]&m[975]&m[976]&m[977]))&UnbiasedRNG[77])|((m[971]&~m[974]&~m[975]&m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&m[975]&~m[976]&m[977])|(~m[971]&~m[974]&~m[975]&m[976]&m[977])|(m[971]&~m[974]&~m[975]&m[976]&m[977])|(~m[971]&m[974]&~m[975]&m[976]&m[977])|(m[971]&m[974]&~m[975]&m[976]&m[977])|(~m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&m[974]&m[975]&m[976]&m[977]))):InitCond[329];
    m[978] = run?((((m[976]&~m[979]&~m[980]&~m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&m[981]&~m[982])|(m[976]&m[979]&~m[980]&m[981]&~m[982])|(m[976]&~m[979]&m[980]&m[981]&~m[982])|(~m[976]&m[979]&~m[980]&~m[981]&m[982])|(~m[976]&~m[979]&m[980]&~m[981]&m[982])|(m[976]&m[979]&m[980]&~m[981]&m[982])|(~m[976]&m[979]&m[980]&m[981]&m[982]))&UnbiasedRNG[78])|((m[976]&~m[979]&~m[980]&m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&m[980]&~m[981]&m[982])|(~m[976]&~m[979]&~m[980]&m[981]&m[982])|(m[976]&~m[979]&~m[980]&m[981]&m[982])|(~m[976]&m[979]&~m[980]&m[981]&m[982])|(m[976]&m[979]&~m[980]&m[981]&m[982])|(~m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&m[979]&m[980]&m[981]&m[982]))):InitCond[330];
    m[983] = run?((((m[981]&~m[984]&~m[985]&~m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&m[986]&~m[987])|(m[981]&m[984]&~m[985]&m[986]&~m[987])|(m[981]&~m[984]&m[985]&m[986]&~m[987])|(~m[981]&m[984]&~m[985]&~m[986]&m[987])|(~m[981]&~m[984]&m[985]&~m[986]&m[987])|(m[981]&m[984]&m[985]&~m[986]&m[987])|(~m[981]&m[984]&m[985]&m[986]&m[987]))&UnbiasedRNG[79])|((m[981]&~m[984]&~m[985]&m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&m[985]&~m[986]&m[987])|(~m[981]&~m[984]&~m[985]&m[986]&m[987])|(m[981]&~m[984]&~m[985]&m[986]&m[987])|(~m[981]&m[984]&~m[985]&m[986]&m[987])|(m[981]&m[984]&~m[985]&m[986]&m[987])|(~m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&m[984]&m[985]&m[986]&m[987]))):InitCond[331];
    m[988] = run?((((m[986]&~m[989]&~m[990]&~m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&m[991]&~m[992])|(m[986]&m[989]&~m[990]&m[991]&~m[992])|(m[986]&~m[989]&m[990]&m[991]&~m[992])|(~m[986]&m[989]&~m[990]&~m[991]&m[992])|(~m[986]&~m[989]&m[990]&~m[991]&m[992])|(m[986]&m[989]&m[990]&~m[991]&m[992])|(~m[986]&m[989]&m[990]&m[991]&m[992]))&UnbiasedRNG[80])|((m[986]&~m[989]&~m[990]&m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&m[990]&~m[991]&m[992])|(~m[986]&~m[989]&~m[990]&m[991]&m[992])|(m[986]&~m[989]&~m[990]&m[991]&m[992])|(~m[986]&m[989]&~m[990]&m[991]&m[992])|(m[986]&m[989]&~m[990]&m[991]&m[992])|(~m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&m[989]&m[990]&m[991]&m[992]))):InitCond[332];
    m[993] = run?((((m[991]&~m[994]&~m[995]&~m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&m[996]&~m[997])|(m[991]&m[994]&~m[995]&m[996]&~m[997])|(m[991]&~m[994]&m[995]&m[996]&~m[997])|(~m[991]&m[994]&~m[995]&~m[996]&m[997])|(~m[991]&~m[994]&m[995]&~m[996]&m[997])|(m[991]&m[994]&m[995]&~m[996]&m[997])|(~m[991]&m[994]&m[995]&m[996]&m[997]))&UnbiasedRNG[81])|((m[991]&~m[994]&~m[995]&m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&m[995]&~m[996]&m[997])|(~m[991]&~m[994]&~m[995]&m[996]&m[997])|(m[991]&~m[994]&~m[995]&m[996]&m[997])|(~m[991]&m[994]&~m[995]&m[996]&m[997])|(m[991]&m[994]&~m[995]&m[996]&m[997])|(~m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&m[994]&m[995]&m[996]&m[997]))):InitCond[333];
    m[998] = run?((((m[996]&~m[999]&~m[1000]&~m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&~m[1002])|(~m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&m[999]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[82])|((m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&m[999]&m[1000]&m[1001]&m[1002]))):InitCond[334];
    m[1003] = run?((((m[543]&~m[1004]&~m[1005]&~m[1006]&~m[1007])|(~m[543]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(m[543]&m[1004]&~m[1005]&m[1006]&~m[1007])|(m[543]&~m[1004]&m[1005]&m[1006]&~m[1007])|(~m[543]&m[1004]&~m[1005]&~m[1006]&m[1007])|(~m[543]&~m[1004]&m[1005]&~m[1006]&m[1007])|(m[543]&m[1004]&m[1005]&~m[1006]&m[1007])|(~m[543]&m[1004]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[83])|((m[543]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(~m[543]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[543]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[543]&m[1004]&~m[1005]&~m[1006]&m[1007])|(m[543]&~m[1004]&m[1005]&~m[1006]&m[1007])|(~m[543]&~m[1004]&~m[1005]&m[1006]&m[1007])|(m[543]&~m[1004]&~m[1005]&m[1006]&m[1007])|(~m[543]&m[1004]&~m[1005]&m[1006]&m[1007])|(m[543]&m[1004]&~m[1005]&m[1006]&m[1007])|(~m[543]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[543]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[543]&m[1004]&m[1005]&m[1006]&m[1007]))):InitCond[335];
    m[1008] = run?((((m[1006]&~m[1009]&~m[1010]&~m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&~m[1012])|(~m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&m[1009]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[84])|((m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&m[1011]&m[1012]))):InitCond[336];
    m[1013] = run?((((m[1011]&~m[1014]&~m[1015]&~m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&~m[1017])|(~m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[85])|((m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))):InitCond[337];
    m[1018] = run?((((m[1016]&~m[1019]&~m[1020]&~m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&~m[1022])|(~m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[86])|((m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))):InitCond[338];
    m[1023] = run?((((m[1021]&~m[1024]&~m[1025]&~m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&~m[1027])|(~m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[87])|((m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))):InitCond[339];
    m[1028] = run?((((m[1026]&~m[1029]&~m[1030]&~m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&~m[1032])|(~m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[88])|((m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))):InitCond[340];
    m[1033] = run?((((m[1031]&~m[1034]&~m[1035]&~m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&~m[1037])|(~m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&m[1034]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[89])|((m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&m[1036]&m[1037]))):InitCond[341];
    m[1038] = run?((((m[1036]&~m[1039]&~m[1040]&~m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&~m[1042])|(~m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[90])|((m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))):InitCond[342];
    m[1043] = run?((((m[1041]&~m[1044]&~m[1045]&~m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&~m[1047])|(~m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[91])|((m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))):InitCond[343];
    m[1048] = run?((((m[1046]&~m[1049]&~m[1050]&~m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&~m[1052])|(~m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&m[1049]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[92])|((m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&m[1051]&m[1052]))):InitCond[344];
    m[1053] = run?((((m[1051]&~m[1054]&~m[1055]&~m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&~m[1057])|(~m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[93])|((m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))):InitCond[345];
    m[1058] = run?((((m[544]&~m[1059]&~m[1060]&~m[1061]&~m[1062])|(~m[544]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(m[544]&m[1059]&~m[1060]&m[1061]&~m[1062])|(m[544]&~m[1059]&m[1060]&m[1061]&~m[1062])|(~m[544]&m[1059]&~m[1060]&~m[1061]&m[1062])|(~m[544]&~m[1059]&m[1060]&~m[1061]&m[1062])|(m[544]&m[1059]&m[1060]&~m[1061]&m[1062])|(~m[544]&m[1059]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[94])|((m[544]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(~m[544]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[544]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[544]&m[1059]&~m[1060]&~m[1061]&m[1062])|(m[544]&~m[1059]&m[1060]&~m[1061]&m[1062])|(~m[544]&~m[1059]&~m[1060]&m[1061]&m[1062])|(m[544]&~m[1059]&~m[1060]&m[1061]&m[1062])|(~m[544]&m[1059]&~m[1060]&m[1061]&m[1062])|(m[544]&m[1059]&~m[1060]&m[1061]&m[1062])|(~m[544]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[544]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[544]&m[1059]&m[1060]&m[1061]&m[1062]))):InitCond[346];
    m[1063] = run?((((m[1061]&~m[1064]&~m[1065]&~m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&~m[1067])|(~m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[95])|((m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))):InitCond[347];
    m[1068] = run?((((m[1066]&~m[1069]&~m[1070]&~m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&~m[1072])|(~m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&m[1069]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[96])|((m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&m[1071]&m[1072]))):InitCond[348];
    m[1073] = run?((((m[1071]&~m[1074]&~m[1075]&~m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&~m[1077])|(~m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[97])|((m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))):InitCond[349];
    m[1078] = run?((((m[1076]&~m[1079]&~m[1080]&~m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&~m[1082])|(~m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[98])|((m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))):InitCond[350];
    m[1083] = run?((((m[1081]&~m[1084]&~m[1085]&~m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&~m[1087])|(~m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&m[1084]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[99])|((m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&m[1086]&m[1087]))):InitCond[351];
    m[1088] = run?((((m[1086]&~m[1089]&~m[1090]&~m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&~m[1092])|(~m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[100])|((m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))):InitCond[352];
    m[1093] = run?((((m[1091]&~m[1094]&~m[1095]&~m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&~m[1097])|(~m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[101])|((m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))):InitCond[353];
    m[1098] = run?((((m[1096]&~m[1099]&~m[1100]&~m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&~m[1102])|(~m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[102])|((m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))):InitCond[354];
    m[1103] = run?((((m[1101]&~m[1104]&~m[1105]&~m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&~m[1107])|(~m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[103])|((m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))):InitCond[355];
    m[1108] = run?((((m[1106]&~m[1109]&~m[1110]&~m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&~m[1112])|(~m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&m[1109]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[104])|((m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&m[1111]&m[1112]))):InitCond[356];
    m[1113] = run?((((m[1111]&~m[1114]&~m[1115]&~m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&~m[1117])|(~m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&m[1114]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[105])|((m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&m[1116]&m[1117]))):InitCond[357];
    m[1118] = run?((((m[545]&~m[1119]&~m[1120]&~m[1121]&~m[1122])|(~m[545]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(m[545]&m[1119]&~m[1120]&m[1121]&~m[1122])|(m[545]&~m[1119]&m[1120]&m[1121]&~m[1122])|(~m[545]&m[1119]&~m[1120]&~m[1121]&m[1122])|(~m[545]&~m[1119]&m[1120]&~m[1121]&m[1122])|(m[545]&m[1119]&m[1120]&~m[1121]&m[1122])|(~m[545]&m[1119]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[106])|((m[545]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(~m[545]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[545]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[545]&m[1119]&~m[1120]&~m[1121]&m[1122])|(m[545]&~m[1119]&m[1120]&~m[1121]&m[1122])|(~m[545]&~m[1119]&~m[1120]&m[1121]&m[1122])|(m[545]&~m[1119]&~m[1120]&m[1121]&m[1122])|(~m[545]&m[1119]&~m[1120]&m[1121]&m[1122])|(m[545]&m[1119]&~m[1120]&m[1121]&m[1122])|(~m[545]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[545]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[545]&m[1119]&m[1120]&m[1121]&m[1122]))):InitCond[358];
    m[1123] = run?((((m[1121]&~m[1124]&~m[1125]&~m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&~m[1127])|(~m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[107])|((m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))):InitCond[359];
    m[1128] = run?((((m[1126]&~m[1129]&~m[1130]&~m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&~m[1132])|(~m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[108])|((m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))):InitCond[360];
    m[1133] = run?((((m[1131]&~m[1134]&~m[1135]&~m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&~m[1137])|(~m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[109])|((m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))):InitCond[361];
    m[1138] = run?((((m[1136]&~m[1139]&~m[1140]&~m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&~m[1142])|(~m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&m[1139]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[110])|((m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&m[1141]&m[1142]))):InitCond[362];
    m[1143] = run?((((m[1141]&~m[1144]&~m[1145]&~m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&~m[1147])|(~m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[111])|((m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))):InitCond[363];
    m[1148] = run?((((m[1146]&~m[1149]&~m[1150]&~m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&~m[1152])|(~m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[112])|((m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))):InitCond[364];
    m[1153] = run?((((m[1151]&~m[1154]&~m[1155]&~m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&~m[1157])|(~m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&m[1154]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[113])|((m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&m[1156]&m[1157]))):InitCond[365];
    m[1158] = run?((((m[1156]&~m[1159]&~m[1160]&~m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&~m[1162])|(~m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&m[1159]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[114])|((m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&m[1161]&m[1162]))):InitCond[366];
    m[1163] = run?((((m[1161]&~m[1164]&~m[1165]&~m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&~m[1167])|(~m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[115])|((m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))):InitCond[367];
    m[1168] = run?((((m[1166]&~m[1169]&~m[1170]&~m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&~m[1172])|(~m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[116])|((m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))):InitCond[368];
    m[1173] = run?((((m[1171]&~m[1174]&~m[1175]&~m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&~m[1177])|(~m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&m[1174]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[117])|((m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&m[1176]&m[1177]))):InitCond[369];
    m[1178] = run?((((m[1176]&~m[1179]&~m[1180]&~m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&~m[1182])|(~m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[118])|((m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))):InitCond[370];
    m[1188] = run?((((m[1186]&~m[1189]&~m[1190]&~m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&~m[1192])|(~m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&m[1189]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[119])|((m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&m[1191]&m[1192]))):InitCond[371];
    m[1193] = run?((((m[1191]&~m[1194]&~m[1195]&~m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&~m[1197])|(~m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&m[1194]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[120])|((m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&m[1196]&m[1197]))):InitCond[372];
    m[1198] = run?((((m[1196]&~m[1199]&~m[1200]&~m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&~m[1202])|(~m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&m[1199]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[121])|((m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&m[1201]&m[1202]))):InitCond[373];
    m[1203] = run?((((m[1201]&~m[1204]&~m[1205]&~m[1206]&~m[1207])|(~m[1201]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(m[1201]&m[1204]&~m[1205]&m[1206]&~m[1207])|(m[1201]&~m[1204]&m[1205]&m[1206]&~m[1207])|(~m[1201]&m[1204]&~m[1205]&~m[1206]&m[1207])|(~m[1201]&~m[1204]&m[1205]&~m[1206]&m[1207])|(m[1201]&m[1204]&m[1205]&~m[1206]&m[1207])|(~m[1201]&m[1204]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[122])|((m[1201]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(~m[1201]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[1201]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[1201]&m[1204]&~m[1205]&~m[1206]&m[1207])|(m[1201]&~m[1204]&m[1205]&~m[1206]&m[1207])|(~m[1201]&~m[1204]&~m[1205]&m[1206]&m[1207])|(m[1201]&~m[1204]&~m[1205]&m[1206]&m[1207])|(~m[1201]&m[1204]&~m[1205]&m[1206]&m[1207])|(m[1201]&m[1204]&~m[1205]&m[1206]&m[1207])|(~m[1201]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[1201]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[1201]&m[1204]&m[1205]&m[1206]&m[1207]))):InitCond[374];
    m[1208] = run?((((m[1206]&~m[1209]&~m[1210]&~m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&~m[1212])|(~m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&m[1209]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[123])|((m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&m[1211]&m[1212]))):InitCond[375];
    m[1213] = run?((((m[1211]&~m[1214]&~m[1215]&~m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&~m[1217])|(~m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&m[1214]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[124])|((m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&m[1216]&m[1217]))):InitCond[376];
    m[1218] = run?((((m[1216]&~m[1219]&~m[1220]&~m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&~m[1222])|(~m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&m[1219]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[125])|((m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&m[1221]&m[1222]))):InitCond[377];
    m[1223] = run?((((m[1221]&~m[1224]&~m[1225]&~m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&~m[1227])|(~m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&m[1224]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[126])|((m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&m[1226]&m[1227]))):InitCond[378];
    m[1228] = run?((((m[1226]&~m[1229]&~m[1230]&~m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&~m[1232])|(~m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&m[1229]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[127])|((m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&m[1231]&m[1232]))):InitCond[379];
    m[1233] = run?((((m[1231]&~m[1234]&~m[1235]&~m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&~m[1237])|(~m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&m[1234]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[128])|((m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&m[1236]&m[1237]))):InitCond[380];
    m[1238] = run?((((m[1236]&~m[1239]&~m[1240]&~m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&~m[1242])|(~m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&m[1239]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[129])|((m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&m[1241]&m[1242]))):InitCond[381];
    m[1243] = run?((((m[1241]&~m[1244]&~m[1245]&~m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&~m[1247])|(~m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&m[1244]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[130])|((m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&m[1246]&m[1247]))):InitCond[382];
    m[1248] = run?((((m[1187]&~m[1249]&~m[1250]&~m[1251]&~m[1252])|(~m[1187]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1187]&m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1187]&~m[1249]&m[1250]&m[1251]&~m[1252])|(~m[1187]&m[1249]&~m[1250]&~m[1251]&m[1252])|(~m[1187]&~m[1249]&m[1250]&~m[1251]&m[1252])|(m[1187]&m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1187]&m[1249]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[131])|((m[1187]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(~m[1187]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1187]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1187]&m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1187]&~m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1187]&~m[1249]&~m[1250]&m[1251]&m[1252])|(m[1187]&~m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1187]&m[1249]&~m[1250]&m[1251]&m[1252])|(m[1187]&m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1187]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1187]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1187]&m[1249]&m[1250]&m[1251]&m[1252]))):InitCond[383];
    m[1253] = run?((((m[1251]&~m[1254]&~m[1255]&~m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&~m[1257])|(~m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&m[1254]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[132])|((m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&m[1256]&m[1257]))):InitCond[384];
    m[1258] = run?((((m[1256]&~m[1259]&~m[1260]&~m[1261]&~m[1262])|(~m[1256]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(m[1256]&m[1259]&~m[1260]&m[1261]&~m[1262])|(m[1256]&~m[1259]&m[1260]&m[1261]&~m[1262])|(~m[1256]&m[1259]&~m[1260]&~m[1261]&m[1262])|(~m[1256]&~m[1259]&m[1260]&~m[1261]&m[1262])|(m[1256]&m[1259]&m[1260]&~m[1261]&m[1262])|(~m[1256]&m[1259]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[133])|((m[1256]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(~m[1256]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[1256]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[1256]&m[1259]&~m[1260]&~m[1261]&m[1262])|(m[1256]&~m[1259]&m[1260]&~m[1261]&m[1262])|(~m[1256]&~m[1259]&~m[1260]&m[1261]&m[1262])|(m[1256]&~m[1259]&~m[1260]&m[1261]&m[1262])|(~m[1256]&m[1259]&~m[1260]&m[1261]&m[1262])|(m[1256]&m[1259]&~m[1260]&m[1261]&m[1262])|(~m[1256]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[1256]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[1256]&m[1259]&m[1260]&m[1261]&m[1262]))):InitCond[385];
    m[1263] = run?((((m[1261]&~m[1264]&~m[1265]&~m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&~m[1267])|(~m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&m[1264]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[134])|((m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&m[1266]&m[1267]))):InitCond[386];
    m[1268] = run?((((m[1266]&~m[1269]&~m[1270]&~m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&~m[1272])|(~m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&m[1269]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[135])|((m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&m[1271]&m[1272]))):InitCond[387];
    m[1273] = run?((((m[1271]&~m[1274]&~m[1275]&~m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&~m[1277])|(~m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&m[1274]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[136])|((m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&m[1276]&m[1277]))):InitCond[388];
    m[1278] = run?((((m[1276]&~m[1279]&~m[1280]&~m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&~m[1282])|(~m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&m[1279]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[137])|((m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&m[1281]&m[1282]))):InitCond[389];
    m[1283] = run?((((m[1281]&~m[1284]&~m[1285]&~m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&~m[1287])|(~m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&m[1284]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[138])|((m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&m[1286]&m[1287]))):InitCond[390];
    m[1288] = run?((((m[1286]&~m[1289]&~m[1290]&~m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&~m[1292])|(~m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&m[1289]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[139])|((m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&m[1291]&m[1292]))):InitCond[391];
    m[1293] = run?((((m[1291]&~m[1294]&~m[1295]&~m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&~m[1297])|(~m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&m[1294]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[140])|((m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&m[1296]&m[1297]))):InitCond[392];
    m[1298] = run?((((m[1296]&~m[1299]&~m[1300]&~m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&~m[1302])|(~m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&m[1299]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[141])|((m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&m[1301]&m[1302]))):InitCond[393];
    m[1303] = run?((((m[1301]&~m[1304]&~m[1305]&~m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&~m[1307])|(~m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&m[1304]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[142])|((m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&m[1306]&m[1307]))):InitCond[394];
    m[1308] = run?((((m[1252]&~m[1309]&~m[1310]&~m[1311]&~m[1312])|(~m[1252]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1252]&m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1252]&~m[1309]&m[1310]&m[1311]&~m[1312])|(~m[1252]&m[1309]&~m[1310]&~m[1311]&m[1312])|(~m[1252]&~m[1309]&m[1310]&~m[1311]&m[1312])|(m[1252]&m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1252]&m[1309]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[143])|((m[1252]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(~m[1252]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1252]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1252]&m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1252]&~m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1252]&~m[1309]&~m[1310]&m[1311]&m[1312])|(m[1252]&~m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1252]&m[1309]&~m[1310]&m[1311]&m[1312])|(m[1252]&m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1252]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1252]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1252]&m[1309]&m[1310]&m[1311]&m[1312]))):InitCond[395];
    m[1313] = run?((((m[1311]&~m[1314]&~m[1315]&~m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&~m[1317])|(~m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&m[1314]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[144])|((m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&m[1316]&m[1317]))):InitCond[396];
    m[1318] = run?((((m[1316]&~m[1319]&~m[1320]&~m[1321]&~m[1322])|(~m[1316]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(m[1316]&m[1319]&~m[1320]&m[1321]&~m[1322])|(m[1316]&~m[1319]&m[1320]&m[1321]&~m[1322])|(~m[1316]&m[1319]&~m[1320]&~m[1321]&m[1322])|(~m[1316]&~m[1319]&m[1320]&~m[1321]&m[1322])|(m[1316]&m[1319]&m[1320]&~m[1321]&m[1322])|(~m[1316]&m[1319]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[145])|((m[1316]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(~m[1316]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[1316]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[1316]&m[1319]&~m[1320]&~m[1321]&m[1322])|(m[1316]&~m[1319]&m[1320]&~m[1321]&m[1322])|(~m[1316]&~m[1319]&~m[1320]&m[1321]&m[1322])|(m[1316]&~m[1319]&~m[1320]&m[1321]&m[1322])|(~m[1316]&m[1319]&~m[1320]&m[1321]&m[1322])|(m[1316]&m[1319]&~m[1320]&m[1321]&m[1322])|(~m[1316]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[1316]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[1316]&m[1319]&m[1320]&m[1321]&m[1322]))):InitCond[397];
    m[1323] = run?((((m[1321]&~m[1324]&~m[1325]&~m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&~m[1327])|(~m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&m[1324]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[146])|((m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&m[1326]&m[1327]))):InitCond[398];
    m[1328] = run?((((m[1326]&~m[1329]&~m[1330]&~m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&~m[1332])|(~m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&m[1329]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[147])|((m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&m[1331]&m[1332]))):InitCond[399];
    m[1333] = run?((((m[1331]&~m[1334]&~m[1335]&~m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&~m[1337])|(~m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&m[1334]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[148])|((m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&m[1336]&m[1337]))):InitCond[400];
    m[1338] = run?((((m[1336]&~m[1339]&~m[1340]&~m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&~m[1342])|(~m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&m[1339]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[149])|((m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&m[1341]&m[1342]))):InitCond[401];
    m[1343] = run?((((m[1341]&~m[1344]&~m[1345]&~m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&~m[1347])|(~m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&m[1344]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[150])|((m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&m[1346]&m[1347]))):InitCond[402];
    m[1348] = run?((((m[1346]&~m[1349]&~m[1350]&~m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&~m[1352])|(~m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&m[1349]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[151])|((m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&m[1351]&m[1352]))):InitCond[403];
    m[1353] = run?((((m[1351]&~m[1354]&~m[1355]&~m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&~m[1357])|(~m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&m[1354]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[152])|((m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&m[1356]&m[1357]))):InitCond[404];
    m[1358] = run?((((m[1356]&~m[1359]&~m[1360]&~m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&~m[1362])|(~m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&m[1359]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[153])|((m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&m[1361]&m[1362]))):InitCond[405];
    m[1363] = run?((((m[1312]&~m[1364]&~m[1365]&~m[1366]&~m[1367])|(~m[1312]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1312]&m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1312]&~m[1364]&m[1365]&m[1366]&~m[1367])|(~m[1312]&m[1364]&~m[1365]&~m[1366]&m[1367])|(~m[1312]&~m[1364]&m[1365]&~m[1366]&m[1367])|(m[1312]&m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1312]&m[1364]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[154])|((m[1312]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(~m[1312]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1312]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1312]&m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1312]&~m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1312]&~m[1364]&~m[1365]&m[1366]&m[1367])|(m[1312]&~m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1312]&m[1364]&~m[1365]&m[1366]&m[1367])|(m[1312]&m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1312]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1312]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1312]&m[1364]&m[1365]&m[1366]&m[1367]))):InitCond[406];
    m[1368] = run?((((m[1366]&~m[1369]&~m[1370]&~m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&~m[1372])|(~m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&m[1369]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[155])|((m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&m[1371]&m[1372]))):InitCond[407];
    m[1373] = run?((((m[1371]&~m[1374]&~m[1375]&~m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&~m[1377])|(~m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&m[1374]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[156])|((m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&m[1376]&m[1377]))):InitCond[408];
    m[1378] = run?((((m[1376]&~m[1379]&~m[1380]&~m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&~m[1382])|(~m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&m[1379]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[157])|((m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&m[1381]&m[1382]))):InitCond[409];
    m[1383] = run?((((m[1381]&~m[1384]&~m[1385]&~m[1386]&~m[1387])|(~m[1381]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(m[1381]&m[1384]&~m[1385]&m[1386]&~m[1387])|(m[1381]&~m[1384]&m[1385]&m[1386]&~m[1387])|(~m[1381]&m[1384]&~m[1385]&~m[1386]&m[1387])|(~m[1381]&~m[1384]&m[1385]&~m[1386]&m[1387])|(m[1381]&m[1384]&m[1385]&~m[1386]&m[1387])|(~m[1381]&m[1384]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[158])|((m[1381]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(~m[1381]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[1381]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[1381]&m[1384]&~m[1385]&~m[1386]&m[1387])|(m[1381]&~m[1384]&m[1385]&~m[1386]&m[1387])|(~m[1381]&~m[1384]&~m[1385]&m[1386]&m[1387])|(m[1381]&~m[1384]&~m[1385]&m[1386]&m[1387])|(~m[1381]&m[1384]&~m[1385]&m[1386]&m[1387])|(m[1381]&m[1384]&~m[1385]&m[1386]&m[1387])|(~m[1381]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[1381]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[1381]&m[1384]&m[1385]&m[1386]&m[1387]))):InitCond[410];
    m[1388] = run?((((m[1386]&~m[1389]&~m[1390]&~m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&~m[1392])|(~m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&m[1389]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[159])|((m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&m[1391]&m[1392]))):InitCond[411];
    m[1393] = run?((((m[1391]&~m[1394]&~m[1395]&~m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&~m[1397])|(~m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&m[1394]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[160])|((m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&m[1396]&m[1397]))):InitCond[412];
    m[1398] = run?((((m[1396]&~m[1399]&~m[1400]&~m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&~m[1402])|(~m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&m[1399]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[161])|((m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&m[1401]&m[1402]))):InitCond[413];
    m[1403] = run?((((m[1401]&~m[1404]&~m[1405]&~m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&~m[1407])|(~m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&m[1404]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[162])|((m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&m[1406]&m[1407]))):InitCond[414];
    m[1408] = run?((((m[1406]&~m[1409]&~m[1410]&~m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&~m[1412])|(~m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&m[1409]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[163])|((m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&m[1411]&m[1412]))):InitCond[415];
    m[1413] = run?((((m[1367]&~m[1414]&~m[1415]&~m[1416]&~m[1417])|(~m[1367]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1367]&m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1367]&~m[1414]&m[1415]&m[1416]&~m[1417])|(~m[1367]&m[1414]&~m[1415]&~m[1416]&m[1417])|(~m[1367]&~m[1414]&m[1415]&~m[1416]&m[1417])|(m[1367]&m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1367]&m[1414]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[164])|((m[1367]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(~m[1367]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1367]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1367]&m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1367]&~m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1367]&~m[1414]&~m[1415]&m[1416]&m[1417])|(m[1367]&~m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1367]&m[1414]&~m[1415]&m[1416]&m[1417])|(m[1367]&m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1367]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1367]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1367]&m[1414]&m[1415]&m[1416]&m[1417]))):InitCond[416];
    m[1418] = run?((((m[1416]&~m[1419]&~m[1420]&~m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&~m[1422])|(~m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&m[1419]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[165])|((m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&m[1421]&m[1422]))):InitCond[417];
    m[1423] = run?((((m[1421]&~m[1424]&~m[1425]&~m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&~m[1427])|(~m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&m[1424]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[166])|((m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&m[1426]&m[1427]))):InitCond[418];
    m[1428] = run?((((m[1426]&~m[1429]&~m[1430]&~m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&~m[1432])|(~m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&m[1429]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[167])|((m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&m[1431]&m[1432]))):InitCond[419];
    m[1433] = run?((((m[1431]&~m[1434]&~m[1435]&~m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&~m[1437])|(~m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&m[1434]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[168])|((m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&m[1436]&m[1437]))):InitCond[420];
    m[1438] = run?((((m[1436]&~m[1439]&~m[1440]&~m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&~m[1442])|(~m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&m[1439]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[169])|((m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&m[1441]&m[1442]))):InitCond[421];
    m[1443] = run?((((m[1441]&~m[1444]&~m[1445]&~m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&~m[1447])|(~m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&m[1444]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[170])|((m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&m[1446]&m[1447]))):InitCond[422];
    m[1448] = run?((((m[1446]&~m[1449]&~m[1450]&~m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&~m[1452])|(~m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&m[1449]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[171])|((m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&m[1451]&m[1452]))):InitCond[423];
    m[1453] = run?((((m[1451]&~m[1454]&~m[1455]&~m[1456]&~m[1457])|(~m[1451]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(m[1451]&m[1454]&~m[1455]&m[1456]&~m[1457])|(m[1451]&~m[1454]&m[1455]&m[1456]&~m[1457])|(~m[1451]&m[1454]&~m[1455]&~m[1456]&m[1457])|(~m[1451]&~m[1454]&m[1455]&~m[1456]&m[1457])|(m[1451]&m[1454]&m[1455]&~m[1456]&m[1457])|(~m[1451]&m[1454]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[172])|((m[1451]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(~m[1451]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[1451]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[1451]&m[1454]&~m[1455]&~m[1456]&m[1457])|(m[1451]&~m[1454]&m[1455]&~m[1456]&m[1457])|(~m[1451]&~m[1454]&~m[1455]&m[1456]&m[1457])|(m[1451]&~m[1454]&~m[1455]&m[1456]&m[1457])|(~m[1451]&m[1454]&~m[1455]&m[1456]&m[1457])|(m[1451]&m[1454]&~m[1455]&m[1456]&m[1457])|(~m[1451]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[1451]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[1451]&m[1454]&m[1455]&m[1456]&m[1457]))):InitCond[424];
    m[1458] = run?((((m[1417]&~m[1459]&~m[1460]&~m[1461]&~m[1462])|(~m[1417]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1417]&m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1417]&~m[1459]&m[1460]&m[1461]&~m[1462])|(~m[1417]&m[1459]&~m[1460]&~m[1461]&m[1462])|(~m[1417]&~m[1459]&m[1460]&~m[1461]&m[1462])|(m[1417]&m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1417]&m[1459]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[173])|((m[1417]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(~m[1417]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1417]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1417]&m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1417]&~m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1417]&~m[1459]&~m[1460]&m[1461]&m[1462])|(m[1417]&~m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1417]&m[1459]&~m[1460]&m[1461]&m[1462])|(m[1417]&m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1417]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1417]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1417]&m[1459]&m[1460]&m[1461]&m[1462]))):InitCond[425];
    m[1463] = run?((((m[1461]&~m[1464]&~m[1465]&~m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&~m[1467])|(~m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&m[1464]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[174])|((m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&m[1466]&m[1467]))):InitCond[426];
    m[1468] = run?((((m[1466]&~m[1469]&~m[1470]&~m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&~m[1472])|(~m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&m[1469]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[175])|((m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&m[1471]&m[1472]))):InitCond[427];
    m[1473] = run?((((m[1471]&~m[1474]&~m[1475]&~m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&~m[1477])|(~m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&m[1474]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[176])|((m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&m[1476]&m[1477]))):InitCond[428];
    m[1478] = run?((((m[1476]&~m[1479]&~m[1480]&~m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&~m[1482])|(~m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&m[1479]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[177])|((m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&m[1481]&m[1482]))):InitCond[429];
    m[1483] = run?((((m[1481]&~m[1484]&~m[1485]&~m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&~m[1487])|(~m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&m[1484]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[178])|((m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&m[1486]&m[1487]))):InitCond[430];
    m[1488] = run?((((m[1486]&~m[1489]&~m[1490]&~m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&~m[1492])|(~m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&m[1489]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[179])|((m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&m[1491]&m[1492]))):InitCond[431];
    m[1493] = run?((((m[1491]&~m[1494]&~m[1495]&~m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&~m[1497])|(~m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&m[1494]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[180])|((m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&m[1496]&m[1497]))):InitCond[432];
    m[1498] = run?((((m[1462]&~m[1499]&~m[1500]&~m[1501]&~m[1502])|(~m[1462]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1462]&m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1462]&~m[1499]&m[1500]&m[1501]&~m[1502])|(~m[1462]&m[1499]&~m[1500]&~m[1501]&m[1502])|(~m[1462]&~m[1499]&m[1500]&~m[1501]&m[1502])|(m[1462]&m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1462]&m[1499]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[181])|((m[1462]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(~m[1462]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1462]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1462]&m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1462]&~m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1462]&~m[1499]&~m[1500]&m[1501]&m[1502])|(m[1462]&~m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1462]&m[1499]&~m[1500]&m[1501]&m[1502])|(m[1462]&m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1462]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1462]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1462]&m[1499]&m[1500]&m[1501]&m[1502]))):InitCond[433];
    m[1503] = run?((((m[1501]&~m[1504]&~m[1505]&~m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&~m[1507])|(~m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&m[1504]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[182])|((m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&m[1506]&m[1507]))):InitCond[434];
    m[1508] = run?((((m[1506]&~m[1509]&~m[1510]&~m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&~m[1512])|(~m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&m[1509]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[183])|((m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&m[1511]&m[1512]))):InitCond[435];
    m[1513] = run?((((m[1511]&~m[1514]&~m[1515]&~m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&~m[1517])|(~m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&m[1514]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[184])|((m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&m[1516]&m[1517]))):InitCond[436];
    m[1518] = run?((((m[1516]&~m[1519]&~m[1520]&~m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&~m[1522])|(~m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&m[1519]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[185])|((m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&m[1521]&m[1522]))):InitCond[437];
    m[1523] = run?((((m[1521]&~m[1524]&~m[1525]&~m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&~m[1527])|(~m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&m[1524]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[186])|((m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&m[1526]&m[1527]))):InitCond[438];
    m[1528] = run?((((m[1526]&~m[1529]&~m[1530]&~m[1531]&~m[1532])|(~m[1526]&~m[1529]&~m[1530]&m[1531]&~m[1532])|(m[1526]&m[1529]&~m[1530]&m[1531]&~m[1532])|(m[1526]&~m[1529]&m[1530]&m[1531]&~m[1532])|(~m[1526]&m[1529]&~m[1530]&~m[1531]&m[1532])|(~m[1526]&~m[1529]&m[1530]&~m[1531]&m[1532])|(m[1526]&m[1529]&m[1530]&~m[1531]&m[1532])|(~m[1526]&m[1529]&m[1530]&m[1531]&m[1532]))&UnbiasedRNG[187])|((m[1526]&~m[1529]&~m[1530]&m[1531]&~m[1532])|(~m[1526]&~m[1529]&~m[1530]&~m[1531]&m[1532])|(m[1526]&~m[1529]&~m[1530]&~m[1531]&m[1532])|(m[1526]&m[1529]&~m[1530]&~m[1531]&m[1532])|(m[1526]&~m[1529]&m[1530]&~m[1531]&m[1532])|(~m[1526]&~m[1529]&~m[1530]&m[1531]&m[1532])|(m[1526]&~m[1529]&~m[1530]&m[1531]&m[1532])|(~m[1526]&m[1529]&~m[1530]&m[1531]&m[1532])|(m[1526]&m[1529]&~m[1530]&m[1531]&m[1532])|(~m[1526]&~m[1529]&m[1530]&m[1531]&m[1532])|(m[1526]&~m[1529]&m[1530]&m[1531]&m[1532])|(m[1526]&m[1529]&m[1530]&m[1531]&m[1532]))):InitCond[439];
    m[1533] = run?((((m[1502]&~m[1534]&~m[1535]&~m[1536]&~m[1537])|(~m[1502]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1502]&m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1502]&~m[1534]&m[1535]&m[1536]&~m[1537])|(~m[1502]&m[1534]&~m[1535]&~m[1536]&m[1537])|(~m[1502]&~m[1534]&m[1535]&~m[1536]&m[1537])|(m[1502]&m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1502]&m[1534]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[188])|((m[1502]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(~m[1502]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1502]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1502]&m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1502]&~m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1502]&~m[1534]&~m[1535]&m[1536]&m[1537])|(m[1502]&~m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1502]&m[1534]&~m[1535]&m[1536]&m[1537])|(m[1502]&m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1502]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1502]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1502]&m[1534]&m[1535]&m[1536]&m[1537]))):InitCond[440];
    m[1538] = run?((((m[1536]&~m[1539]&~m[1540]&~m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&~m[1542])|(~m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&m[1539]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[189])|((m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&m[1541]&m[1542]))):InitCond[441];
    m[1543] = run?((((m[1541]&~m[1544]&~m[1545]&~m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&~m[1547])|(~m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&m[1544]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[190])|((m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&m[1546]&m[1547]))):InitCond[442];
    m[1548] = run?((((m[1546]&~m[1549]&~m[1550]&~m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&~m[1552])|(~m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&m[1549]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[191])|((m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&m[1551]&m[1552]))):InitCond[443];
    m[1553] = run?((((m[1551]&~m[1554]&~m[1555]&~m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&~m[1557])|(~m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&m[1554]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[192])|((m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&m[1556]&m[1557]))):InitCond[444];
    m[1558] = run?((((m[1556]&~m[1559]&~m[1560]&~m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&~m[1562])|(~m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&m[1559]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[193])|((m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&m[1561]&m[1562]))):InitCond[445];
    m[1563] = run?((((m[1537]&~m[1564]&~m[1565]&~m[1566]&~m[1567])|(~m[1537]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1537]&m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1537]&~m[1564]&m[1565]&m[1566]&~m[1567])|(~m[1537]&m[1564]&~m[1565]&~m[1566]&m[1567])|(~m[1537]&~m[1564]&m[1565]&~m[1566]&m[1567])|(m[1537]&m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1537]&m[1564]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[194])|((m[1537]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(~m[1537]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1537]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1537]&m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1537]&~m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1537]&~m[1564]&~m[1565]&m[1566]&m[1567])|(m[1537]&~m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1537]&m[1564]&~m[1565]&m[1566]&m[1567])|(m[1537]&m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1537]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1537]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1537]&m[1564]&m[1565]&m[1566]&m[1567]))):InitCond[446];
    m[1568] = run?((((m[1566]&~m[1569]&~m[1570]&~m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&~m[1572])|(~m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&m[1569]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[195])|((m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&m[1571]&m[1572]))):InitCond[447];
    m[1573] = run?((((m[1571]&~m[1574]&~m[1575]&~m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&~m[1577])|(~m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&m[1574]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[196])|((m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&m[1576]&m[1577]))):InitCond[448];
    m[1578] = run?((((m[1576]&~m[1579]&~m[1580]&~m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&~m[1582])|(~m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&m[1579]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[197])|((m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&m[1581]&m[1582]))):InitCond[449];
    m[1583] = run?((((m[1581]&~m[1584]&~m[1585]&~m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&~m[1587])|(~m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&m[1584]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[198])|((m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&m[1586]&m[1587]))):InitCond[450];
    m[1588] = run?((((m[1567]&~m[1589]&~m[1590]&~m[1591]&~m[1592])|(~m[1567]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1567]&m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1567]&~m[1589]&m[1590]&m[1591]&~m[1592])|(~m[1567]&m[1589]&~m[1590]&~m[1591]&m[1592])|(~m[1567]&~m[1589]&m[1590]&~m[1591]&m[1592])|(m[1567]&m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1567]&m[1589]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[199])|((m[1567]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(~m[1567]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1567]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1567]&m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1567]&~m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1567]&~m[1589]&~m[1590]&m[1591]&m[1592])|(m[1567]&~m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1567]&m[1589]&~m[1590]&m[1591]&m[1592])|(m[1567]&m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1567]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1567]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1567]&m[1589]&m[1590]&m[1591]&m[1592]))):InitCond[451];
    m[1593] = run?((((m[1591]&~m[1594]&~m[1595]&~m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&~m[1597])|(~m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&m[1594]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[200])|((m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&m[1596]&m[1597]))):InitCond[452];
    m[1598] = run?((((m[1596]&~m[1599]&~m[1600]&~m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&~m[1602])|(~m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&m[1599]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[201])|((m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&m[1601]&m[1602]))):InitCond[453];
    m[1603] = run?((((m[1601]&~m[1604]&~m[1605]&~m[1606]&~m[1607])|(~m[1601]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1601]&m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1601]&~m[1604]&m[1605]&m[1606]&~m[1607])|(~m[1601]&m[1604]&~m[1605]&~m[1606]&m[1607])|(~m[1601]&~m[1604]&m[1605]&~m[1606]&m[1607])|(m[1601]&m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1601]&m[1604]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[202])|((m[1601]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(~m[1601]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1601]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1601]&m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1601]&~m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1601]&~m[1604]&~m[1605]&m[1606]&m[1607])|(m[1601]&~m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1601]&m[1604]&~m[1605]&m[1606]&m[1607])|(m[1601]&m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1601]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1601]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1601]&m[1604]&m[1605]&m[1606]&m[1607]))):InitCond[454];
    m[1608] = run?((((m[1592]&~m[1609]&~m[1610]&~m[1611]&~m[1612])|(~m[1592]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1592]&m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1592]&~m[1609]&m[1610]&m[1611]&~m[1612])|(~m[1592]&m[1609]&~m[1610]&~m[1611]&m[1612])|(~m[1592]&~m[1609]&m[1610]&~m[1611]&m[1612])|(m[1592]&m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1592]&m[1609]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[203])|((m[1592]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(~m[1592]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1592]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1592]&m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1592]&~m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1592]&~m[1609]&~m[1610]&m[1611]&m[1612])|(m[1592]&~m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1592]&m[1609]&~m[1610]&m[1611]&m[1612])|(m[1592]&m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1592]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1592]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1592]&m[1609]&m[1610]&m[1611]&m[1612]))):InitCond[455];
    m[1613] = run?((((m[1611]&~m[1614]&~m[1615]&~m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&~m[1617])|(~m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&m[1614]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[204])|((m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&m[1616]&m[1617]))):InitCond[456];
    m[1618] = run?((((m[1616]&~m[1619]&~m[1620]&~m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&~m[1622])|(~m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&m[1619]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[205])|((m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&m[1621]&m[1622]))):InitCond[457];
    m[1623] = run?((((m[1612]&~m[1624]&~m[1625]&~m[1626]&~m[1627])|(~m[1612]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1612]&m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1612]&~m[1624]&m[1625]&m[1626]&~m[1627])|(~m[1612]&m[1624]&~m[1625]&~m[1626]&m[1627])|(~m[1612]&~m[1624]&m[1625]&~m[1626]&m[1627])|(m[1612]&m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1612]&m[1624]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[206])|((m[1612]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(~m[1612]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1612]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1612]&m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1612]&~m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1612]&~m[1624]&~m[1625]&m[1626]&m[1627])|(m[1612]&~m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1612]&m[1624]&~m[1625]&m[1626]&m[1627])|(m[1612]&m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1612]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1612]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1612]&m[1624]&m[1625]&m[1626]&m[1627]))):InitCond[458];
    m[1628] = run?((((m[1626]&~m[1629]&~m[1630]&~m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&~m[1632])|(~m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&m[1629]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[207])|((m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&m[1631]&m[1632]))):InitCond[459];
    m[1633] = run?((((m[1627]&~m[1634]&~m[1635]&~m[1636]&~m[1637])|(~m[1627]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1627]&m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1627]&~m[1634]&m[1635]&m[1636]&~m[1637])|(~m[1627]&m[1634]&~m[1635]&~m[1636]&m[1637])|(~m[1627]&~m[1634]&m[1635]&~m[1636]&m[1637])|(m[1627]&m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1627]&m[1634]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[208])|((m[1627]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(~m[1627]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1627]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1627]&m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1627]&~m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1627]&~m[1634]&~m[1635]&m[1636]&m[1637])|(m[1627]&~m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1627]&m[1634]&~m[1635]&m[1636]&m[1637])|(m[1627]&m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1627]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1627]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1627]&m[1634]&m[1635]&m[1636]&m[1637]))):InitCond[460];
end

always @(posedge color1_clk) begin
    m[28] = run?((((m[0]&m[57]&~m[58]&~m[140]&~m[141])|(m[0]&~m[57]&m[58]&~m[140]&~m[141])|(~m[0]&m[57]&m[58]&~m[140]&~m[141])|(m[0]&~m[57]&~m[58]&m[140]&~m[141])|(~m[0]&m[57]&~m[58]&m[140]&~m[141])|(~m[0]&~m[57]&m[58]&m[140]&~m[141])|(m[0]&~m[57]&~m[58]&~m[140]&m[141])|(~m[0]&m[57]&~m[58]&~m[140]&m[141])|(~m[0]&~m[57]&m[58]&~m[140]&m[141])|(~m[0]&~m[57]&~m[58]&m[140]&m[141]))&BiasedRNG[252])|(((m[0]&m[57]&m[58]&~m[140]&~m[141])|(m[0]&m[57]&~m[58]&m[140]&~m[141])|(m[0]&~m[57]&m[58]&m[140]&~m[141])|(~m[0]&m[57]&m[58]&m[140]&~m[141])|(m[0]&m[57]&~m[58]&~m[140]&m[141])|(m[0]&~m[57]&m[58]&~m[140]&m[141])|(~m[0]&m[57]&m[58]&~m[140]&m[141])|(m[0]&~m[57]&~m[58]&m[140]&m[141])|(~m[0]&m[57]&~m[58]&m[140]&m[141])|(~m[0]&~m[57]&m[58]&m[140]&m[141]))&~BiasedRNG[252])|((m[0]&m[57]&m[58]&m[140]&~m[141])|(m[0]&m[57]&m[58]&~m[140]&m[141])|(m[0]&m[57]&~m[58]&m[140]&m[141])|(m[0]&~m[57]&m[58]&m[140]&m[141])|(~m[0]&m[57]&m[58]&m[140]&m[141])|(m[0]&m[57]&m[58]&m[140]&m[141]))):InitCond[461];
    m[29] = run?((((m[1]&m[60]&~m[61]&~m[154]&~m[155])|(m[1]&~m[60]&m[61]&~m[154]&~m[155])|(~m[1]&m[60]&m[61]&~m[154]&~m[155])|(m[1]&~m[60]&~m[61]&m[154]&~m[155])|(~m[1]&m[60]&~m[61]&m[154]&~m[155])|(~m[1]&~m[60]&m[61]&m[154]&~m[155])|(m[1]&~m[60]&~m[61]&~m[154]&m[155])|(~m[1]&m[60]&~m[61]&~m[154]&m[155])|(~m[1]&~m[60]&m[61]&~m[154]&m[155])|(~m[1]&~m[60]&~m[61]&m[154]&m[155]))&BiasedRNG[253])|(((m[1]&m[60]&m[61]&~m[154]&~m[155])|(m[1]&m[60]&~m[61]&m[154]&~m[155])|(m[1]&~m[60]&m[61]&m[154]&~m[155])|(~m[1]&m[60]&m[61]&m[154]&~m[155])|(m[1]&m[60]&~m[61]&~m[154]&m[155])|(m[1]&~m[60]&m[61]&~m[154]&m[155])|(~m[1]&m[60]&m[61]&~m[154]&m[155])|(m[1]&~m[60]&~m[61]&m[154]&m[155])|(~m[1]&m[60]&~m[61]&m[154]&m[155])|(~m[1]&~m[60]&m[61]&m[154]&m[155]))&~BiasedRNG[253])|((m[1]&m[60]&m[61]&m[154]&~m[155])|(m[1]&m[60]&m[61]&~m[154]&m[155])|(m[1]&m[60]&~m[61]&m[154]&m[155])|(m[1]&~m[60]&m[61]&m[154]&m[155])|(~m[1]&m[60]&m[61]&m[154]&m[155])|(m[1]&m[60]&m[61]&m[154]&m[155]))):InitCond[462];
    m[30] = run?((((m[2]&m[63]&~m[64]&~m[168]&~m[169])|(m[2]&~m[63]&m[64]&~m[168]&~m[169])|(~m[2]&m[63]&m[64]&~m[168]&~m[169])|(m[2]&~m[63]&~m[64]&m[168]&~m[169])|(~m[2]&m[63]&~m[64]&m[168]&~m[169])|(~m[2]&~m[63]&m[64]&m[168]&~m[169])|(m[2]&~m[63]&~m[64]&~m[168]&m[169])|(~m[2]&m[63]&~m[64]&~m[168]&m[169])|(~m[2]&~m[63]&m[64]&~m[168]&m[169])|(~m[2]&~m[63]&~m[64]&m[168]&m[169]))&BiasedRNG[254])|(((m[2]&m[63]&m[64]&~m[168]&~m[169])|(m[2]&m[63]&~m[64]&m[168]&~m[169])|(m[2]&~m[63]&m[64]&m[168]&~m[169])|(~m[2]&m[63]&m[64]&m[168]&~m[169])|(m[2]&m[63]&~m[64]&~m[168]&m[169])|(m[2]&~m[63]&m[64]&~m[168]&m[169])|(~m[2]&m[63]&m[64]&~m[168]&m[169])|(m[2]&~m[63]&~m[64]&m[168]&m[169])|(~m[2]&m[63]&~m[64]&m[168]&m[169])|(~m[2]&~m[63]&m[64]&m[168]&m[169]))&~BiasedRNG[254])|((m[2]&m[63]&m[64]&m[168]&~m[169])|(m[2]&m[63]&m[64]&~m[168]&m[169])|(m[2]&m[63]&~m[64]&m[168]&m[169])|(m[2]&~m[63]&m[64]&m[168]&m[169])|(~m[2]&m[63]&m[64]&m[168]&m[169])|(m[2]&m[63]&m[64]&m[168]&m[169]))):InitCond[463];
    m[31] = run?((((m[3]&m[66]&~m[67]&~m[182]&~m[183])|(m[3]&~m[66]&m[67]&~m[182]&~m[183])|(~m[3]&m[66]&m[67]&~m[182]&~m[183])|(m[3]&~m[66]&~m[67]&m[182]&~m[183])|(~m[3]&m[66]&~m[67]&m[182]&~m[183])|(~m[3]&~m[66]&m[67]&m[182]&~m[183])|(m[3]&~m[66]&~m[67]&~m[182]&m[183])|(~m[3]&m[66]&~m[67]&~m[182]&m[183])|(~m[3]&~m[66]&m[67]&~m[182]&m[183])|(~m[3]&~m[66]&~m[67]&m[182]&m[183]))&BiasedRNG[255])|(((m[3]&m[66]&m[67]&~m[182]&~m[183])|(m[3]&m[66]&~m[67]&m[182]&~m[183])|(m[3]&~m[66]&m[67]&m[182]&~m[183])|(~m[3]&m[66]&m[67]&m[182]&~m[183])|(m[3]&m[66]&~m[67]&~m[182]&m[183])|(m[3]&~m[66]&m[67]&~m[182]&m[183])|(~m[3]&m[66]&m[67]&~m[182]&m[183])|(m[3]&~m[66]&~m[67]&m[182]&m[183])|(~m[3]&m[66]&~m[67]&m[182]&m[183])|(~m[3]&~m[66]&m[67]&m[182]&m[183]))&~BiasedRNG[255])|((m[3]&m[66]&m[67]&m[182]&~m[183])|(m[3]&m[66]&m[67]&~m[182]&m[183])|(m[3]&m[66]&~m[67]&m[182]&m[183])|(m[3]&~m[66]&m[67]&m[182]&m[183])|(~m[3]&m[66]&m[67]&m[182]&m[183])|(m[3]&m[66]&m[67]&m[182]&m[183]))):InitCond[464];
    m[32] = run?((((m[4]&m[69]&~m[70]&~m[196]&~m[197])|(m[4]&~m[69]&m[70]&~m[196]&~m[197])|(~m[4]&m[69]&m[70]&~m[196]&~m[197])|(m[4]&~m[69]&~m[70]&m[196]&~m[197])|(~m[4]&m[69]&~m[70]&m[196]&~m[197])|(~m[4]&~m[69]&m[70]&m[196]&~m[197])|(m[4]&~m[69]&~m[70]&~m[196]&m[197])|(~m[4]&m[69]&~m[70]&~m[196]&m[197])|(~m[4]&~m[69]&m[70]&~m[196]&m[197])|(~m[4]&~m[69]&~m[70]&m[196]&m[197]))&BiasedRNG[256])|(((m[4]&m[69]&m[70]&~m[196]&~m[197])|(m[4]&m[69]&~m[70]&m[196]&~m[197])|(m[4]&~m[69]&m[70]&m[196]&~m[197])|(~m[4]&m[69]&m[70]&m[196]&~m[197])|(m[4]&m[69]&~m[70]&~m[196]&m[197])|(m[4]&~m[69]&m[70]&~m[196]&m[197])|(~m[4]&m[69]&m[70]&~m[196]&m[197])|(m[4]&~m[69]&~m[70]&m[196]&m[197])|(~m[4]&m[69]&~m[70]&m[196]&m[197])|(~m[4]&~m[69]&m[70]&m[196]&m[197]))&~BiasedRNG[256])|((m[4]&m[69]&m[70]&m[196]&~m[197])|(m[4]&m[69]&m[70]&~m[196]&m[197])|(m[4]&m[69]&~m[70]&m[196]&m[197])|(m[4]&~m[69]&m[70]&m[196]&m[197])|(~m[4]&m[69]&m[70]&m[196]&m[197])|(m[4]&m[69]&m[70]&m[196]&m[197]))):InitCond[465];
    m[33] = run?((((m[5]&m[72]&~m[73]&~m[210]&~m[211])|(m[5]&~m[72]&m[73]&~m[210]&~m[211])|(~m[5]&m[72]&m[73]&~m[210]&~m[211])|(m[5]&~m[72]&~m[73]&m[210]&~m[211])|(~m[5]&m[72]&~m[73]&m[210]&~m[211])|(~m[5]&~m[72]&m[73]&m[210]&~m[211])|(m[5]&~m[72]&~m[73]&~m[210]&m[211])|(~m[5]&m[72]&~m[73]&~m[210]&m[211])|(~m[5]&~m[72]&m[73]&~m[210]&m[211])|(~m[5]&~m[72]&~m[73]&m[210]&m[211]))&BiasedRNG[257])|(((m[5]&m[72]&m[73]&~m[210]&~m[211])|(m[5]&m[72]&~m[73]&m[210]&~m[211])|(m[5]&~m[72]&m[73]&m[210]&~m[211])|(~m[5]&m[72]&m[73]&m[210]&~m[211])|(m[5]&m[72]&~m[73]&~m[210]&m[211])|(m[5]&~m[72]&m[73]&~m[210]&m[211])|(~m[5]&m[72]&m[73]&~m[210]&m[211])|(m[5]&~m[72]&~m[73]&m[210]&m[211])|(~m[5]&m[72]&~m[73]&m[210]&m[211])|(~m[5]&~m[72]&m[73]&m[210]&m[211]))&~BiasedRNG[257])|((m[5]&m[72]&m[73]&m[210]&~m[211])|(m[5]&m[72]&m[73]&~m[210]&m[211])|(m[5]&m[72]&~m[73]&m[210]&m[211])|(m[5]&~m[72]&m[73]&m[210]&m[211])|(~m[5]&m[72]&m[73]&m[210]&m[211])|(m[5]&m[72]&m[73]&m[210]&m[211]))):InitCond[466];
    m[34] = run?((((m[6]&m[75]&~m[76]&~m[224]&~m[225])|(m[6]&~m[75]&m[76]&~m[224]&~m[225])|(~m[6]&m[75]&m[76]&~m[224]&~m[225])|(m[6]&~m[75]&~m[76]&m[224]&~m[225])|(~m[6]&m[75]&~m[76]&m[224]&~m[225])|(~m[6]&~m[75]&m[76]&m[224]&~m[225])|(m[6]&~m[75]&~m[76]&~m[224]&m[225])|(~m[6]&m[75]&~m[76]&~m[224]&m[225])|(~m[6]&~m[75]&m[76]&~m[224]&m[225])|(~m[6]&~m[75]&~m[76]&m[224]&m[225]))&BiasedRNG[258])|(((m[6]&m[75]&m[76]&~m[224]&~m[225])|(m[6]&m[75]&~m[76]&m[224]&~m[225])|(m[6]&~m[75]&m[76]&m[224]&~m[225])|(~m[6]&m[75]&m[76]&m[224]&~m[225])|(m[6]&m[75]&~m[76]&~m[224]&m[225])|(m[6]&~m[75]&m[76]&~m[224]&m[225])|(~m[6]&m[75]&m[76]&~m[224]&m[225])|(m[6]&~m[75]&~m[76]&m[224]&m[225])|(~m[6]&m[75]&~m[76]&m[224]&m[225])|(~m[6]&~m[75]&m[76]&m[224]&m[225]))&~BiasedRNG[258])|((m[6]&m[75]&m[76]&m[224]&~m[225])|(m[6]&m[75]&m[76]&~m[224]&m[225])|(m[6]&m[75]&~m[76]&m[224]&m[225])|(m[6]&~m[75]&m[76]&m[224]&m[225])|(~m[6]&m[75]&m[76]&m[224]&m[225])|(m[6]&m[75]&m[76]&m[224]&m[225]))):InitCond[467];
    m[35] = run?((((m[7]&m[78]&~m[79]&~m[238]&~m[239])|(m[7]&~m[78]&m[79]&~m[238]&~m[239])|(~m[7]&m[78]&m[79]&~m[238]&~m[239])|(m[7]&~m[78]&~m[79]&m[238]&~m[239])|(~m[7]&m[78]&~m[79]&m[238]&~m[239])|(~m[7]&~m[78]&m[79]&m[238]&~m[239])|(m[7]&~m[78]&~m[79]&~m[238]&m[239])|(~m[7]&m[78]&~m[79]&~m[238]&m[239])|(~m[7]&~m[78]&m[79]&~m[238]&m[239])|(~m[7]&~m[78]&~m[79]&m[238]&m[239]))&BiasedRNG[259])|(((m[7]&m[78]&m[79]&~m[238]&~m[239])|(m[7]&m[78]&~m[79]&m[238]&~m[239])|(m[7]&~m[78]&m[79]&m[238]&~m[239])|(~m[7]&m[78]&m[79]&m[238]&~m[239])|(m[7]&m[78]&~m[79]&~m[238]&m[239])|(m[7]&~m[78]&m[79]&~m[238]&m[239])|(~m[7]&m[78]&m[79]&~m[238]&m[239])|(m[7]&~m[78]&~m[79]&m[238]&m[239])|(~m[7]&m[78]&~m[79]&m[238]&m[239])|(~m[7]&~m[78]&m[79]&m[238]&m[239]))&~BiasedRNG[259])|((m[7]&m[78]&m[79]&m[238]&~m[239])|(m[7]&m[78]&m[79]&~m[238]&m[239])|(m[7]&m[78]&~m[79]&m[238]&m[239])|(m[7]&~m[78]&m[79]&m[238]&m[239])|(~m[7]&m[78]&m[79]&m[238]&m[239])|(m[7]&m[78]&m[79]&m[238]&m[239]))):InitCond[468];
    m[36] = run?((((m[8]&m[81]&~m[82]&~m[252]&~m[253])|(m[8]&~m[81]&m[82]&~m[252]&~m[253])|(~m[8]&m[81]&m[82]&~m[252]&~m[253])|(m[8]&~m[81]&~m[82]&m[252]&~m[253])|(~m[8]&m[81]&~m[82]&m[252]&~m[253])|(~m[8]&~m[81]&m[82]&m[252]&~m[253])|(m[8]&~m[81]&~m[82]&~m[252]&m[253])|(~m[8]&m[81]&~m[82]&~m[252]&m[253])|(~m[8]&~m[81]&m[82]&~m[252]&m[253])|(~m[8]&~m[81]&~m[82]&m[252]&m[253]))&BiasedRNG[260])|(((m[8]&m[81]&m[82]&~m[252]&~m[253])|(m[8]&m[81]&~m[82]&m[252]&~m[253])|(m[8]&~m[81]&m[82]&m[252]&~m[253])|(~m[8]&m[81]&m[82]&m[252]&~m[253])|(m[8]&m[81]&~m[82]&~m[252]&m[253])|(m[8]&~m[81]&m[82]&~m[252]&m[253])|(~m[8]&m[81]&m[82]&~m[252]&m[253])|(m[8]&~m[81]&~m[82]&m[252]&m[253])|(~m[8]&m[81]&~m[82]&m[252]&m[253])|(~m[8]&~m[81]&m[82]&m[252]&m[253]))&~BiasedRNG[260])|((m[8]&m[81]&m[82]&m[252]&~m[253])|(m[8]&m[81]&m[82]&~m[252]&m[253])|(m[8]&m[81]&~m[82]&m[252]&m[253])|(m[8]&~m[81]&m[82]&m[252]&m[253])|(~m[8]&m[81]&m[82]&m[252]&m[253])|(m[8]&m[81]&m[82]&m[252]&m[253]))):InitCond[469];
    m[37] = run?((((m[9]&m[84]&~m[85]&~m[266]&~m[267])|(m[9]&~m[84]&m[85]&~m[266]&~m[267])|(~m[9]&m[84]&m[85]&~m[266]&~m[267])|(m[9]&~m[84]&~m[85]&m[266]&~m[267])|(~m[9]&m[84]&~m[85]&m[266]&~m[267])|(~m[9]&~m[84]&m[85]&m[266]&~m[267])|(m[9]&~m[84]&~m[85]&~m[266]&m[267])|(~m[9]&m[84]&~m[85]&~m[266]&m[267])|(~m[9]&~m[84]&m[85]&~m[266]&m[267])|(~m[9]&~m[84]&~m[85]&m[266]&m[267]))&BiasedRNG[261])|(((m[9]&m[84]&m[85]&~m[266]&~m[267])|(m[9]&m[84]&~m[85]&m[266]&~m[267])|(m[9]&~m[84]&m[85]&m[266]&~m[267])|(~m[9]&m[84]&m[85]&m[266]&~m[267])|(m[9]&m[84]&~m[85]&~m[266]&m[267])|(m[9]&~m[84]&m[85]&~m[266]&m[267])|(~m[9]&m[84]&m[85]&~m[266]&m[267])|(m[9]&~m[84]&~m[85]&m[266]&m[267])|(~m[9]&m[84]&~m[85]&m[266]&m[267])|(~m[9]&~m[84]&m[85]&m[266]&m[267]))&~BiasedRNG[261])|((m[9]&m[84]&m[85]&m[266]&~m[267])|(m[9]&m[84]&m[85]&~m[266]&m[267])|(m[9]&m[84]&~m[85]&m[266]&m[267])|(m[9]&~m[84]&m[85]&m[266]&m[267])|(~m[9]&m[84]&m[85]&m[266]&m[267])|(m[9]&m[84]&m[85]&m[266]&m[267]))):InitCond[470];
    m[38] = run?((((m[10]&m[87]&~m[88]&~m[280]&~m[281])|(m[10]&~m[87]&m[88]&~m[280]&~m[281])|(~m[10]&m[87]&m[88]&~m[280]&~m[281])|(m[10]&~m[87]&~m[88]&m[280]&~m[281])|(~m[10]&m[87]&~m[88]&m[280]&~m[281])|(~m[10]&~m[87]&m[88]&m[280]&~m[281])|(m[10]&~m[87]&~m[88]&~m[280]&m[281])|(~m[10]&m[87]&~m[88]&~m[280]&m[281])|(~m[10]&~m[87]&m[88]&~m[280]&m[281])|(~m[10]&~m[87]&~m[88]&m[280]&m[281]))&BiasedRNG[262])|(((m[10]&m[87]&m[88]&~m[280]&~m[281])|(m[10]&m[87]&~m[88]&m[280]&~m[281])|(m[10]&~m[87]&m[88]&m[280]&~m[281])|(~m[10]&m[87]&m[88]&m[280]&~m[281])|(m[10]&m[87]&~m[88]&~m[280]&m[281])|(m[10]&~m[87]&m[88]&~m[280]&m[281])|(~m[10]&m[87]&m[88]&~m[280]&m[281])|(m[10]&~m[87]&~m[88]&m[280]&m[281])|(~m[10]&m[87]&~m[88]&m[280]&m[281])|(~m[10]&~m[87]&m[88]&m[280]&m[281]))&~BiasedRNG[262])|((m[10]&m[87]&m[88]&m[280]&~m[281])|(m[10]&m[87]&m[88]&~m[280]&m[281])|(m[10]&m[87]&~m[88]&m[280]&m[281])|(m[10]&~m[87]&m[88]&m[280]&m[281])|(~m[10]&m[87]&m[88]&m[280]&m[281])|(m[10]&m[87]&m[88]&m[280]&m[281]))):InitCond[471];
    m[39] = run?((((m[11]&m[90]&~m[91]&~m[294]&~m[295])|(m[11]&~m[90]&m[91]&~m[294]&~m[295])|(~m[11]&m[90]&m[91]&~m[294]&~m[295])|(m[11]&~m[90]&~m[91]&m[294]&~m[295])|(~m[11]&m[90]&~m[91]&m[294]&~m[295])|(~m[11]&~m[90]&m[91]&m[294]&~m[295])|(m[11]&~m[90]&~m[91]&~m[294]&m[295])|(~m[11]&m[90]&~m[91]&~m[294]&m[295])|(~m[11]&~m[90]&m[91]&~m[294]&m[295])|(~m[11]&~m[90]&~m[91]&m[294]&m[295]))&BiasedRNG[263])|(((m[11]&m[90]&m[91]&~m[294]&~m[295])|(m[11]&m[90]&~m[91]&m[294]&~m[295])|(m[11]&~m[90]&m[91]&m[294]&~m[295])|(~m[11]&m[90]&m[91]&m[294]&~m[295])|(m[11]&m[90]&~m[91]&~m[294]&m[295])|(m[11]&~m[90]&m[91]&~m[294]&m[295])|(~m[11]&m[90]&m[91]&~m[294]&m[295])|(m[11]&~m[90]&~m[91]&m[294]&m[295])|(~m[11]&m[90]&~m[91]&m[294]&m[295])|(~m[11]&~m[90]&m[91]&m[294]&m[295]))&~BiasedRNG[263])|((m[11]&m[90]&m[91]&m[294]&~m[295])|(m[11]&m[90]&m[91]&~m[294]&m[295])|(m[11]&m[90]&~m[91]&m[294]&m[295])|(m[11]&~m[90]&m[91]&m[294]&m[295])|(~m[11]&m[90]&m[91]&m[294]&m[295])|(m[11]&m[90]&m[91]&m[294]&m[295]))):InitCond[472];
    m[40] = run?((((m[12]&m[93]&~m[94]&~m[308]&~m[309])|(m[12]&~m[93]&m[94]&~m[308]&~m[309])|(~m[12]&m[93]&m[94]&~m[308]&~m[309])|(m[12]&~m[93]&~m[94]&m[308]&~m[309])|(~m[12]&m[93]&~m[94]&m[308]&~m[309])|(~m[12]&~m[93]&m[94]&m[308]&~m[309])|(m[12]&~m[93]&~m[94]&~m[308]&m[309])|(~m[12]&m[93]&~m[94]&~m[308]&m[309])|(~m[12]&~m[93]&m[94]&~m[308]&m[309])|(~m[12]&~m[93]&~m[94]&m[308]&m[309]))&BiasedRNG[264])|(((m[12]&m[93]&m[94]&~m[308]&~m[309])|(m[12]&m[93]&~m[94]&m[308]&~m[309])|(m[12]&~m[93]&m[94]&m[308]&~m[309])|(~m[12]&m[93]&m[94]&m[308]&~m[309])|(m[12]&m[93]&~m[94]&~m[308]&m[309])|(m[12]&~m[93]&m[94]&~m[308]&m[309])|(~m[12]&m[93]&m[94]&~m[308]&m[309])|(m[12]&~m[93]&~m[94]&m[308]&m[309])|(~m[12]&m[93]&~m[94]&m[308]&m[309])|(~m[12]&~m[93]&m[94]&m[308]&m[309]))&~BiasedRNG[264])|((m[12]&m[93]&m[94]&m[308]&~m[309])|(m[12]&m[93]&m[94]&~m[308]&m[309])|(m[12]&m[93]&~m[94]&m[308]&m[309])|(m[12]&~m[93]&m[94]&m[308]&m[309])|(~m[12]&m[93]&m[94]&m[308]&m[309])|(m[12]&m[93]&m[94]&m[308]&m[309]))):InitCond[473];
    m[41] = run?((((m[13]&m[96]&~m[97]&~m[322]&~m[323])|(m[13]&~m[96]&m[97]&~m[322]&~m[323])|(~m[13]&m[96]&m[97]&~m[322]&~m[323])|(m[13]&~m[96]&~m[97]&m[322]&~m[323])|(~m[13]&m[96]&~m[97]&m[322]&~m[323])|(~m[13]&~m[96]&m[97]&m[322]&~m[323])|(m[13]&~m[96]&~m[97]&~m[322]&m[323])|(~m[13]&m[96]&~m[97]&~m[322]&m[323])|(~m[13]&~m[96]&m[97]&~m[322]&m[323])|(~m[13]&~m[96]&~m[97]&m[322]&m[323]))&BiasedRNG[265])|(((m[13]&m[96]&m[97]&~m[322]&~m[323])|(m[13]&m[96]&~m[97]&m[322]&~m[323])|(m[13]&~m[96]&m[97]&m[322]&~m[323])|(~m[13]&m[96]&m[97]&m[322]&~m[323])|(m[13]&m[96]&~m[97]&~m[322]&m[323])|(m[13]&~m[96]&m[97]&~m[322]&m[323])|(~m[13]&m[96]&m[97]&~m[322]&m[323])|(m[13]&~m[96]&~m[97]&m[322]&m[323])|(~m[13]&m[96]&~m[97]&m[322]&m[323])|(~m[13]&~m[96]&m[97]&m[322]&m[323]))&~BiasedRNG[265])|((m[13]&m[96]&m[97]&m[322]&~m[323])|(m[13]&m[96]&m[97]&~m[322]&m[323])|(m[13]&m[96]&~m[97]&m[322]&m[323])|(m[13]&~m[96]&m[97]&m[322]&m[323])|(~m[13]&m[96]&m[97]&m[322]&m[323])|(m[13]&m[96]&m[97]&m[322]&m[323]))):InitCond[474];
    m[42] = run?((((m[14]&m[99]&~m[100]&~m[336]&~m[337])|(m[14]&~m[99]&m[100]&~m[336]&~m[337])|(~m[14]&m[99]&m[100]&~m[336]&~m[337])|(m[14]&~m[99]&~m[100]&m[336]&~m[337])|(~m[14]&m[99]&~m[100]&m[336]&~m[337])|(~m[14]&~m[99]&m[100]&m[336]&~m[337])|(m[14]&~m[99]&~m[100]&~m[336]&m[337])|(~m[14]&m[99]&~m[100]&~m[336]&m[337])|(~m[14]&~m[99]&m[100]&~m[336]&m[337])|(~m[14]&~m[99]&~m[100]&m[336]&m[337]))&BiasedRNG[266])|(((m[14]&m[99]&m[100]&~m[336]&~m[337])|(m[14]&m[99]&~m[100]&m[336]&~m[337])|(m[14]&~m[99]&m[100]&m[336]&~m[337])|(~m[14]&m[99]&m[100]&m[336]&~m[337])|(m[14]&m[99]&~m[100]&~m[336]&m[337])|(m[14]&~m[99]&m[100]&~m[336]&m[337])|(~m[14]&m[99]&m[100]&~m[336]&m[337])|(m[14]&~m[99]&~m[100]&m[336]&m[337])|(~m[14]&m[99]&~m[100]&m[336]&m[337])|(~m[14]&~m[99]&m[100]&m[336]&m[337]))&~BiasedRNG[266])|((m[14]&m[99]&m[100]&m[336]&~m[337])|(m[14]&m[99]&m[100]&~m[336]&m[337])|(m[14]&m[99]&~m[100]&m[336]&m[337])|(m[14]&~m[99]&m[100]&m[336]&m[337])|(~m[14]&m[99]&m[100]&m[336]&m[337])|(m[14]&m[99]&m[100]&m[336]&m[337]))):InitCond[475];
    m[43] = run?((((m[15]&m[102]&~m[103]&~m[350]&~m[351])|(m[15]&~m[102]&m[103]&~m[350]&~m[351])|(~m[15]&m[102]&m[103]&~m[350]&~m[351])|(m[15]&~m[102]&~m[103]&m[350]&~m[351])|(~m[15]&m[102]&~m[103]&m[350]&~m[351])|(~m[15]&~m[102]&m[103]&m[350]&~m[351])|(m[15]&~m[102]&~m[103]&~m[350]&m[351])|(~m[15]&m[102]&~m[103]&~m[350]&m[351])|(~m[15]&~m[102]&m[103]&~m[350]&m[351])|(~m[15]&~m[102]&~m[103]&m[350]&m[351]))&BiasedRNG[267])|(((m[15]&m[102]&m[103]&~m[350]&~m[351])|(m[15]&m[102]&~m[103]&m[350]&~m[351])|(m[15]&~m[102]&m[103]&m[350]&~m[351])|(~m[15]&m[102]&m[103]&m[350]&~m[351])|(m[15]&m[102]&~m[103]&~m[350]&m[351])|(m[15]&~m[102]&m[103]&~m[350]&m[351])|(~m[15]&m[102]&m[103]&~m[350]&m[351])|(m[15]&~m[102]&~m[103]&m[350]&m[351])|(~m[15]&m[102]&~m[103]&m[350]&m[351])|(~m[15]&~m[102]&m[103]&m[350]&m[351]))&~BiasedRNG[267])|((m[15]&m[102]&m[103]&m[350]&~m[351])|(m[15]&m[102]&m[103]&~m[350]&m[351])|(m[15]&m[102]&~m[103]&m[350]&m[351])|(m[15]&~m[102]&m[103]&m[350]&m[351])|(~m[15]&m[102]&m[103]&m[350]&m[351])|(m[15]&m[102]&m[103]&m[350]&m[351]))):InitCond[476];
    m[44] = run?((((m[16]&m[105]&~m[106]&~m[364]&~m[365])|(m[16]&~m[105]&m[106]&~m[364]&~m[365])|(~m[16]&m[105]&m[106]&~m[364]&~m[365])|(m[16]&~m[105]&~m[106]&m[364]&~m[365])|(~m[16]&m[105]&~m[106]&m[364]&~m[365])|(~m[16]&~m[105]&m[106]&m[364]&~m[365])|(m[16]&~m[105]&~m[106]&~m[364]&m[365])|(~m[16]&m[105]&~m[106]&~m[364]&m[365])|(~m[16]&~m[105]&m[106]&~m[364]&m[365])|(~m[16]&~m[105]&~m[106]&m[364]&m[365]))&BiasedRNG[268])|(((m[16]&m[105]&m[106]&~m[364]&~m[365])|(m[16]&m[105]&~m[106]&m[364]&~m[365])|(m[16]&~m[105]&m[106]&m[364]&~m[365])|(~m[16]&m[105]&m[106]&m[364]&~m[365])|(m[16]&m[105]&~m[106]&~m[364]&m[365])|(m[16]&~m[105]&m[106]&~m[364]&m[365])|(~m[16]&m[105]&m[106]&~m[364]&m[365])|(m[16]&~m[105]&~m[106]&m[364]&m[365])|(~m[16]&m[105]&~m[106]&m[364]&m[365])|(~m[16]&~m[105]&m[106]&m[364]&m[365]))&~BiasedRNG[268])|((m[16]&m[105]&m[106]&m[364]&~m[365])|(m[16]&m[105]&m[106]&~m[364]&m[365])|(m[16]&m[105]&~m[106]&m[364]&m[365])|(m[16]&~m[105]&m[106]&m[364]&m[365])|(~m[16]&m[105]&m[106]&m[364]&m[365])|(m[16]&m[105]&m[106]&m[364]&m[365]))):InitCond[477];
    m[45] = run?((((m[17]&m[108]&~m[109]&~m[378]&~m[379])|(m[17]&~m[108]&m[109]&~m[378]&~m[379])|(~m[17]&m[108]&m[109]&~m[378]&~m[379])|(m[17]&~m[108]&~m[109]&m[378]&~m[379])|(~m[17]&m[108]&~m[109]&m[378]&~m[379])|(~m[17]&~m[108]&m[109]&m[378]&~m[379])|(m[17]&~m[108]&~m[109]&~m[378]&m[379])|(~m[17]&m[108]&~m[109]&~m[378]&m[379])|(~m[17]&~m[108]&m[109]&~m[378]&m[379])|(~m[17]&~m[108]&~m[109]&m[378]&m[379]))&BiasedRNG[269])|(((m[17]&m[108]&m[109]&~m[378]&~m[379])|(m[17]&m[108]&~m[109]&m[378]&~m[379])|(m[17]&~m[108]&m[109]&m[378]&~m[379])|(~m[17]&m[108]&m[109]&m[378]&~m[379])|(m[17]&m[108]&~m[109]&~m[378]&m[379])|(m[17]&~m[108]&m[109]&~m[378]&m[379])|(~m[17]&m[108]&m[109]&~m[378]&m[379])|(m[17]&~m[108]&~m[109]&m[378]&m[379])|(~m[17]&m[108]&~m[109]&m[378]&m[379])|(~m[17]&~m[108]&m[109]&m[378]&m[379]))&~BiasedRNG[269])|((m[17]&m[108]&m[109]&m[378]&~m[379])|(m[17]&m[108]&m[109]&~m[378]&m[379])|(m[17]&m[108]&~m[109]&m[378]&m[379])|(m[17]&~m[108]&m[109]&m[378]&m[379])|(~m[17]&m[108]&m[109]&m[378]&m[379])|(m[17]&m[108]&m[109]&m[378]&m[379]))):InitCond[478];
    m[46] = run?((((m[18]&m[111]&~m[112]&~m[392]&~m[393])|(m[18]&~m[111]&m[112]&~m[392]&~m[393])|(~m[18]&m[111]&m[112]&~m[392]&~m[393])|(m[18]&~m[111]&~m[112]&m[392]&~m[393])|(~m[18]&m[111]&~m[112]&m[392]&~m[393])|(~m[18]&~m[111]&m[112]&m[392]&~m[393])|(m[18]&~m[111]&~m[112]&~m[392]&m[393])|(~m[18]&m[111]&~m[112]&~m[392]&m[393])|(~m[18]&~m[111]&m[112]&~m[392]&m[393])|(~m[18]&~m[111]&~m[112]&m[392]&m[393]))&BiasedRNG[270])|(((m[18]&m[111]&m[112]&~m[392]&~m[393])|(m[18]&m[111]&~m[112]&m[392]&~m[393])|(m[18]&~m[111]&m[112]&m[392]&~m[393])|(~m[18]&m[111]&m[112]&m[392]&~m[393])|(m[18]&m[111]&~m[112]&~m[392]&m[393])|(m[18]&~m[111]&m[112]&~m[392]&m[393])|(~m[18]&m[111]&m[112]&~m[392]&m[393])|(m[18]&~m[111]&~m[112]&m[392]&m[393])|(~m[18]&m[111]&~m[112]&m[392]&m[393])|(~m[18]&~m[111]&m[112]&m[392]&m[393]))&~BiasedRNG[270])|((m[18]&m[111]&m[112]&m[392]&~m[393])|(m[18]&m[111]&m[112]&~m[392]&m[393])|(m[18]&m[111]&~m[112]&m[392]&m[393])|(m[18]&~m[111]&m[112]&m[392]&m[393])|(~m[18]&m[111]&m[112]&m[392]&m[393])|(m[18]&m[111]&m[112]&m[392]&m[393]))):InitCond[479];
    m[47] = run?((((m[19]&m[114]&~m[115]&~m[406]&~m[407])|(m[19]&~m[114]&m[115]&~m[406]&~m[407])|(~m[19]&m[114]&m[115]&~m[406]&~m[407])|(m[19]&~m[114]&~m[115]&m[406]&~m[407])|(~m[19]&m[114]&~m[115]&m[406]&~m[407])|(~m[19]&~m[114]&m[115]&m[406]&~m[407])|(m[19]&~m[114]&~m[115]&~m[406]&m[407])|(~m[19]&m[114]&~m[115]&~m[406]&m[407])|(~m[19]&~m[114]&m[115]&~m[406]&m[407])|(~m[19]&~m[114]&~m[115]&m[406]&m[407]))&BiasedRNG[271])|(((m[19]&m[114]&m[115]&~m[406]&~m[407])|(m[19]&m[114]&~m[115]&m[406]&~m[407])|(m[19]&~m[114]&m[115]&m[406]&~m[407])|(~m[19]&m[114]&m[115]&m[406]&~m[407])|(m[19]&m[114]&~m[115]&~m[406]&m[407])|(m[19]&~m[114]&m[115]&~m[406]&m[407])|(~m[19]&m[114]&m[115]&~m[406]&m[407])|(m[19]&~m[114]&~m[115]&m[406]&m[407])|(~m[19]&m[114]&~m[115]&m[406]&m[407])|(~m[19]&~m[114]&m[115]&m[406]&m[407]))&~BiasedRNG[271])|((m[19]&m[114]&m[115]&m[406]&~m[407])|(m[19]&m[114]&m[115]&~m[406]&m[407])|(m[19]&m[114]&~m[115]&m[406]&m[407])|(m[19]&~m[114]&m[115]&m[406]&m[407])|(~m[19]&m[114]&m[115]&m[406]&m[407])|(m[19]&m[114]&m[115]&m[406]&m[407]))):InitCond[480];
    m[48] = run?((((m[20]&m[117]&~m[118]&~m[420]&~m[421])|(m[20]&~m[117]&m[118]&~m[420]&~m[421])|(~m[20]&m[117]&m[118]&~m[420]&~m[421])|(m[20]&~m[117]&~m[118]&m[420]&~m[421])|(~m[20]&m[117]&~m[118]&m[420]&~m[421])|(~m[20]&~m[117]&m[118]&m[420]&~m[421])|(m[20]&~m[117]&~m[118]&~m[420]&m[421])|(~m[20]&m[117]&~m[118]&~m[420]&m[421])|(~m[20]&~m[117]&m[118]&~m[420]&m[421])|(~m[20]&~m[117]&~m[118]&m[420]&m[421]))&BiasedRNG[272])|(((m[20]&m[117]&m[118]&~m[420]&~m[421])|(m[20]&m[117]&~m[118]&m[420]&~m[421])|(m[20]&~m[117]&m[118]&m[420]&~m[421])|(~m[20]&m[117]&m[118]&m[420]&~m[421])|(m[20]&m[117]&~m[118]&~m[420]&m[421])|(m[20]&~m[117]&m[118]&~m[420]&m[421])|(~m[20]&m[117]&m[118]&~m[420]&m[421])|(m[20]&~m[117]&~m[118]&m[420]&m[421])|(~m[20]&m[117]&~m[118]&m[420]&m[421])|(~m[20]&~m[117]&m[118]&m[420]&m[421]))&~BiasedRNG[272])|((m[20]&m[117]&m[118]&m[420]&~m[421])|(m[20]&m[117]&m[118]&~m[420]&m[421])|(m[20]&m[117]&~m[118]&m[420]&m[421])|(m[20]&~m[117]&m[118]&m[420]&m[421])|(~m[20]&m[117]&m[118]&m[420]&m[421])|(m[20]&m[117]&m[118]&m[420]&m[421]))):InitCond[481];
    m[49] = run?((((m[21]&m[120]&~m[121]&~m[434]&~m[435])|(m[21]&~m[120]&m[121]&~m[434]&~m[435])|(~m[21]&m[120]&m[121]&~m[434]&~m[435])|(m[21]&~m[120]&~m[121]&m[434]&~m[435])|(~m[21]&m[120]&~m[121]&m[434]&~m[435])|(~m[21]&~m[120]&m[121]&m[434]&~m[435])|(m[21]&~m[120]&~m[121]&~m[434]&m[435])|(~m[21]&m[120]&~m[121]&~m[434]&m[435])|(~m[21]&~m[120]&m[121]&~m[434]&m[435])|(~m[21]&~m[120]&~m[121]&m[434]&m[435]))&BiasedRNG[273])|(((m[21]&m[120]&m[121]&~m[434]&~m[435])|(m[21]&m[120]&~m[121]&m[434]&~m[435])|(m[21]&~m[120]&m[121]&m[434]&~m[435])|(~m[21]&m[120]&m[121]&m[434]&~m[435])|(m[21]&m[120]&~m[121]&~m[434]&m[435])|(m[21]&~m[120]&m[121]&~m[434]&m[435])|(~m[21]&m[120]&m[121]&~m[434]&m[435])|(m[21]&~m[120]&~m[121]&m[434]&m[435])|(~m[21]&m[120]&~m[121]&m[434]&m[435])|(~m[21]&~m[120]&m[121]&m[434]&m[435]))&~BiasedRNG[273])|((m[21]&m[120]&m[121]&m[434]&~m[435])|(m[21]&m[120]&m[121]&~m[434]&m[435])|(m[21]&m[120]&~m[121]&m[434]&m[435])|(m[21]&~m[120]&m[121]&m[434]&m[435])|(~m[21]&m[120]&m[121]&m[434]&m[435])|(m[21]&m[120]&m[121]&m[434]&m[435]))):InitCond[482];
    m[50] = run?((((m[22]&m[123]&~m[124]&~m[448]&~m[449])|(m[22]&~m[123]&m[124]&~m[448]&~m[449])|(~m[22]&m[123]&m[124]&~m[448]&~m[449])|(m[22]&~m[123]&~m[124]&m[448]&~m[449])|(~m[22]&m[123]&~m[124]&m[448]&~m[449])|(~m[22]&~m[123]&m[124]&m[448]&~m[449])|(m[22]&~m[123]&~m[124]&~m[448]&m[449])|(~m[22]&m[123]&~m[124]&~m[448]&m[449])|(~m[22]&~m[123]&m[124]&~m[448]&m[449])|(~m[22]&~m[123]&~m[124]&m[448]&m[449]))&BiasedRNG[274])|(((m[22]&m[123]&m[124]&~m[448]&~m[449])|(m[22]&m[123]&~m[124]&m[448]&~m[449])|(m[22]&~m[123]&m[124]&m[448]&~m[449])|(~m[22]&m[123]&m[124]&m[448]&~m[449])|(m[22]&m[123]&~m[124]&~m[448]&m[449])|(m[22]&~m[123]&m[124]&~m[448]&m[449])|(~m[22]&m[123]&m[124]&~m[448]&m[449])|(m[22]&~m[123]&~m[124]&m[448]&m[449])|(~m[22]&m[123]&~m[124]&m[448]&m[449])|(~m[22]&~m[123]&m[124]&m[448]&m[449]))&~BiasedRNG[274])|((m[22]&m[123]&m[124]&m[448]&~m[449])|(m[22]&m[123]&m[124]&~m[448]&m[449])|(m[22]&m[123]&~m[124]&m[448]&m[449])|(m[22]&~m[123]&m[124]&m[448]&m[449])|(~m[22]&m[123]&m[124]&m[448]&m[449])|(m[22]&m[123]&m[124]&m[448]&m[449]))):InitCond[483];
    m[51] = run?((((m[23]&m[126]&~m[127]&~m[462]&~m[463])|(m[23]&~m[126]&m[127]&~m[462]&~m[463])|(~m[23]&m[126]&m[127]&~m[462]&~m[463])|(m[23]&~m[126]&~m[127]&m[462]&~m[463])|(~m[23]&m[126]&~m[127]&m[462]&~m[463])|(~m[23]&~m[126]&m[127]&m[462]&~m[463])|(m[23]&~m[126]&~m[127]&~m[462]&m[463])|(~m[23]&m[126]&~m[127]&~m[462]&m[463])|(~m[23]&~m[126]&m[127]&~m[462]&m[463])|(~m[23]&~m[126]&~m[127]&m[462]&m[463]))&BiasedRNG[275])|(((m[23]&m[126]&m[127]&~m[462]&~m[463])|(m[23]&m[126]&~m[127]&m[462]&~m[463])|(m[23]&~m[126]&m[127]&m[462]&~m[463])|(~m[23]&m[126]&m[127]&m[462]&~m[463])|(m[23]&m[126]&~m[127]&~m[462]&m[463])|(m[23]&~m[126]&m[127]&~m[462]&m[463])|(~m[23]&m[126]&m[127]&~m[462]&m[463])|(m[23]&~m[126]&~m[127]&m[462]&m[463])|(~m[23]&m[126]&~m[127]&m[462]&m[463])|(~m[23]&~m[126]&m[127]&m[462]&m[463]))&~BiasedRNG[275])|((m[23]&m[126]&m[127]&m[462]&~m[463])|(m[23]&m[126]&m[127]&~m[462]&m[463])|(m[23]&m[126]&~m[127]&m[462]&m[463])|(m[23]&~m[126]&m[127]&m[462]&m[463])|(~m[23]&m[126]&m[127]&m[462]&m[463])|(m[23]&m[126]&m[127]&m[462]&m[463]))):InitCond[484];
    m[52] = run?((((m[24]&m[129]&~m[130]&~m[476]&~m[477])|(m[24]&~m[129]&m[130]&~m[476]&~m[477])|(~m[24]&m[129]&m[130]&~m[476]&~m[477])|(m[24]&~m[129]&~m[130]&m[476]&~m[477])|(~m[24]&m[129]&~m[130]&m[476]&~m[477])|(~m[24]&~m[129]&m[130]&m[476]&~m[477])|(m[24]&~m[129]&~m[130]&~m[476]&m[477])|(~m[24]&m[129]&~m[130]&~m[476]&m[477])|(~m[24]&~m[129]&m[130]&~m[476]&m[477])|(~m[24]&~m[129]&~m[130]&m[476]&m[477]))&BiasedRNG[276])|(((m[24]&m[129]&m[130]&~m[476]&~m[477])|(m[24]&m[129]&~m[130]&m[476]&~m[477])|(m[24]&~m[129]&m[130]&m[476]&~m[477])|(~m[24]&m[129]&m[130]&m[476]&~m[477])|(m[24]&m[129]&~m[130]&~m[476]&m[477])|(m[24]&~m[129]&m[130]&~m[476]&m[477])|(~m[24]&m[129]&m[130]&~m[476]&m[477])|(m[24]&~m[129]&~m[130]&m[476]&m[477])|(~m[24]&m[129]&~m[130]&m[476]&m[477])|(~m[24]&~m[129]&m[130]&m[476]&m[477]))&~BiasedRNG[276])|((m[24]&m[129]&m[130]&m[476]&~m[477])|(m[24]&m[129]&m[130]&~m[476]&m[477])|(m[24]&m[129]&~m[130]&m[476]&m[477])|(m[24]&~m[129]&m[130]&m[476]&m[477])|(~m[24]&m[129]&m[130]&m[476]&m[477])|(m[24]&m[129]&m[130]&m[476]&m[477]))):InitCond[485];
    m[53] = run?((((m[25]&m[132]&~m[133]&~m[490]&~m[491])|(m[25]&~m[132]&m[133]&~m[490]&~m[491])|(~m[25]&m[132]&m[133]&~m[490]&~m[491])|(m[25]&~m[132]&~m[133]&m[490]&~m[491])|(~m[25]&m[132]&~m[133]&m[490]&~m[491])|(~m[25]&~m[132]&m[133]&m[490]&~m[491])|(m[25]&~m[132]&~m[133]&~m[490]&m[491])|(~m[25]&m[132]&~m[133]&~m[490]&m[491])|(~m[25]&~m[132]&m[133]&~m[490]&m[491])|(~m[25]&~m[132]&~m[133]&m[490]&m[491]))&BiasedRNG[277])|(((m[25]&m[132]&m[133]&~m[490]&~m[491])|(m[25]&m[132]&~m[133]&m[490]&~m[491])|(m[25]&~m[132]&m[133]&m[490]&~m[491])|(~m[25]&m[132]&m[133]&m[490]&~m[491])|(m[25]&m[132]&~m[133]&~m[490]&m[491])|(m[25]&~m[132]&m[133]&~m[490]&m[491])|(~m[25]&m[132]&m[133]&~m[490]&m[491])|(m[25]&~m[132]&~m[133]&m[490]&m[491])|(~m[25]&m[132]&~m[133]&m[490]&m[491])|(~m[25]&~m[132]&m[133]&m[490]&m[491]))&~BiasedRNG[277])|((m[25]&m[132]&m[133]&m[490]&~m[491])|(m[25]&m[132]&m[133]&~m[490]&m[491])|(m[25]&m[132]&~m[133]&m[490]&m[491])|(m[25]&~m[132]&m[133]&m[490]&m[491])|(~m[25]&m[132]&m[133]&m[490]&m[491])|(m[25]&m[132]&m[133]&m[490]&m[491]))):InitCond[486];
    m[54] = run?((((m[26]&m[135]&~m[136]&~m[504]&~m[505])|(m[26]&~m[135]&m[136]&~m[504]&~m[505])|(~m[26]&m[135]&m[136]&~m[504]&~m[505])|(m[26]&~m[135]&~m[136]&m[504]&~m[505])|(~m[26]&m[135]&~m[136]&m[504]&~m[505])|(~m[26]&~m[135]&m[136]&m[504]&~m[505])|(m[26]&~m[135]&~m[136]&~m[504]&m[505])|(~m[26]&m[135]&~m[136]&~m[504]&m[505])|(~m[26]&~m[135]&m[136]&~m[504]&m[505])|(~m[26]&~m[135]&~m[136]&m[504]&m[505]))&BiasedRNG[278])|(((m[26]&m[135]&m[136]&~m[504]&~m[505])|(m[26]&m[135]&~m[136]&m[504]&~m[505])|(m[26]&~m[135]&m[136]&m[504]&~m[505])|(~m[26]&m[135]&m[136]&m[504]&~m[505])|(m[26]&m[135]&~m[136]&~m[504]&m[505])|(m[26]&~m[135]&m[136]&~m[504]&m[505])|(~m[26]&m[135]&m[136]&~m[504]&m[505])|(m[26]&~m[135]&~m[136]&m[504]&m[505])|(~m[26]&m[135]&~m[136]&m[504]&m[505])|(~m[26]&~m[135]&m[136]&m[504]&m[505]))&~BiasedRNG[278])|((m[26]&m[135]&m[136]&m[504]&~m[505])|(m[26]&m[135]&m[136]&~m[504]&m[505])|(m[26]&m[135]&~m[136]&m[504]&m[505])|(m[26]&~m[135]&m[136]&m[504]&m[505])|(~m[26]&m[135]&m[136]&m[504]&m[505])|(m[26]&m[135]&m[136]&m[504]&m[505]))):InitCond[487];
    m[55] = run?((((m[27]&m[138]&~m[139]&~m[518]&~m[519])|(m[27]&~m[138]&m[139]&~m[518]&~m[519])|(~m[27]&m[138]&m[139]&~m[518]&~m[519])|(m[27]&~m[138]&~m[139]&m[518]&~m[519])|(~m[27]&m[138]&~m[139]&m[518]&~m[519])|(~m[27]&~m[138]&m[139]&m[518]&~m[519])|(m[27]&~m[138]&~m[139]&~m[518]&m[519])|(~m[27]&m[138]&~m[139]&~m[518]&m[519])|(~m[27]&~m[138]&m[139]&~m[518]&m[519])|(~m[27]&~m[138]&~m[139]&m[518]&m[519]))&BiasedRNG[279])|(((m[27]&m[138]&m[139]&~m[518]&~m[519])|(m[27]&m[138]&~m[139]&m[518]&~m[519])|(m[27]&~m[138]&m[139]&m[518]&~m[519])|(~m[27]&m[138]&m[139]&m[518]&~m[519])|(m[27]&m[138]&~m[139]&~m[518]&m[519])|(m[27]&~m[138]&m[139]&~m[518]&m[519])|(~m[27]&m[138]&m[139]&~m[518]&m[519])|(m[27]&~m[138]&~m[139]&m[518]&m[519])|(~m[27]&m[138]&~m[139]&m[518]&m[519])|(~m[27]&~m[138]&m[139]&m[518]&m[519]))&~BiasedRNG[279])|((m[27]&m[138]&m[139]&m[518]&~m[519])|(m[27]&m[138]&m[139]&~m[518]&m[519])|(m[27]&m[138]&~m[139]&m[518]&m[519])|(m[27]&~m[138]&m[139]&m[518]&m[519])|(~m[27]&m[138]&m[139]&m[518]&m[519])|(m[27]&m[138]&m[139]&m[518]&m[519]))):InitCond[488];
    m[56] = run?((((m[0]&m[142]&~m[143]&~m[144]&~m[145])|(m[0]&~m[142]&m[143]&~m[144]&~m[145])|(~m[0]&m[142]&m[143]&~m[144]&~m[145])|(m[0]&~m[142]&~m[143]&m[144]&~m[145])|(~m[0]&m[142]&~m[143]&m[144]&~m[145])|(~m[0]&~m[142]&m[143]&m[144]&~m[145])|(m[0]&~m[142]&~m[143]&~m[144]&m[145])|(~m[0]&m[142]&~m[143]&~m[144]&m[145])|(~m[0]&~m[142]&m[143]&~m[144]&m[145])|(~m[0]&~m[142]&~m[143]&m[144]&m[145]))&BiasedRNG[280])|(((m[0]&m[142]&m[143]&~m[144]&~m[145])|(m[0]&m[142]&~m[143]&m[144]&~m[145])|(m[0]&~m[142]&m[143]&m[144]&~m[145])|(~m[0]&m[142]&m[143]&m[144]&~m[145])|(m[0]&m[142]&~m[143]&~m[144]&m[145])|(m[0]&~m[142]&m[143]&~m[144]&m[145])|(~m[0]&m[142]&m[143]&~m[144]&m[145])|(m[0]&~m[142]&~m[143]&m[144]&m[145])|(~m[0]&m[142]&~m[143]&m[144]&m[145])|(~m[0]&~m[142]&m[143]&m[144]&m[145]))&~BiasedRNG[280])|((m[0]&m[142]&m[143]&m[144]&~m[145])|(m[0]&m[142]&m[143]&~m[144]&m[145])|(m[0]&m[142]&~m[143]&m[144]&m[145])|(m[0]&~m[142]&m[143]&m[144]&m[145])|(~m[0]&m[142]&m[143]&m[144]&m[145])|(m[0]&m[142]&m[143]&m[144]&m[145]))):InitCond[489];
    m[59] = run?((((m[1]&m[156]&~m[157]&~m[158]&~m[159])|(m[1]&~m[156]&m[157]&~m[158]&~m[159])|(~m[1]&m[156]&m[157]&~m[158]&~m[159])|(m[1]&~m[156]&~m[157]&m[158]&~m[159])|(~m[1]&m[156]&~m[157]&m[158]&~m[159])|(~m[1]&~m[156]&m[157]&m[158]&~m[159])|(m[1]&~m[156]&~m[157]&~m[158]&m[159])|(~m[1]&m[156]&~m[157]&~m[158]&m[159])|(~m[1]&~m[156]&m[157]&~m[158]&m[159])|(~m[1]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[281])|(((m[1]&m[156]&m[157]&~m[158]&~m[159])|(m[1]&m[156]&~m[157]&m[158]&~m[159])|(m[1]&~m[156]&m[157]&m[158]&~m[159])|(~m[1]&m[156]&m[157]&m[158]&~m[159])|(m[1]&m[156]&~m[157]&~m[158]&m[159])|(m[1]&~m[156]&m[157]&~m[158]&m[159])|(~m[1]&m[156]&m[157]&~m[158]&m[159])|(m[1]&~m[156]&~m[157]&m[158]&m[159])|(~m[1]&m[156]&~m[157]&m[158]&m[159])|(~m[1]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[281])|((m[1]&m[156]&m[157]&m[158]&~m[159])|(m[1]&m[156]&m[157]&~m[158]&m[159])|(m[1]&m[156]&~m[157]&m[158]&m[159])|(m[1]&~m[156]&m[157]&m[158]&m[159])|(~m[1]&m[156]&m[157]&m[158]&m[159])|(m[1]&m[156]&m[157]&m[158]&m[159]))):InitCond[490];
    m[62] = run?((((m[2]&m[170]&~m[171]&~m[172]&~m[173])|(m[2]&~m[170]&m[171]&~m[172]&~m[173])|(~m[2]&m[170]&m[171]&~m[172]&~m[173])|(m[2]&~m[170]&~m[171]&m[172]&~m[173])|(~m[2]&m[170]&~m[171]&m[172]&~m[173])|(~m[2]&~m[170]&m[171]&m[172]&~m[173])|(m[2]&~m[170]&~m[171]&~m[172]&m[173])|(~m[2]&m[170]&~m[171]&~m[172]&m[173])|(~m[2]&~m[170]&m[171]&~m[172]&m[173])|(~m[2]&~m[170]&~m[171]&m[172]&m[173]))&BiasedRNG[282])|(((m[2]&m[170]&m[171]&~m[172]&~m[173])|(m[2]&m[170]&~m[171]&m[172]&~m[173])|(m[2]&~m[170]&m[171]&m[172]&~m[173])|(~m[2]&m[170]&m[171]&m[172]&~m[173])|(m[2]&m[170]&~m[171]&~m[172]&m[173])|(m[2]&~m[170]&m[171]&~m[172]&m[173])|(~m[2]&m[170]&m[171]&~m[172]&m[173])|(m[2]&~m[170]&~m[171]&m[172]&m[173])|(~m[2]&m[170]&~m[171]&m[172]&m[173])|(~m[2]&~m[170]&m[171]&m[172]&m[173]))&~BiasedRNG[282])|((m[2]&m[170]&m[171]&m[172]&~m[173])|(m[2]&m[170]&m[171]&~m[172]&m[173])|(m[2]&m[170]&~m[171]&m[172]&m[173])|(m[2]&~m[170]&m[171]&m[172]&m[173])|(~m[2]&m[170]&m[171]&m[172]&m[173])|(m[2]&m[170]&m[171]&m[172]&m[173]))):InitCond[491];
    m[65] = run?((((m[3]&m[184]&~m[185]&~m[186]&~m[187])|(m[3]&~m[184]&m[185]&~m[186]&~m[187])|(~m[3]&m[184]&m[185]&~m[186]&~m[187])|(m[3]&~m[184]&~m[185]&m[186]&~m[187])|(~m[3]&m[184]&~m[185]&m[186]&~m[187])|(~m[3]&~m[184]&m[185]&m[186]&~m[187])|(m[3]&~m[184]&~m[185]&~m[186]&m[187])|(~m[3]&m[184]&~m[185]&~m[186]&m[187])|(~m[3]&~m[184]&m[185]&~m[186]&m[187])|(~m[3]&~m[184]&~m[185]&m[186]&m[187]))&BiasedRNG[283])|(((m[3]&m[184]&m[185]&~m[186]&~m[187])|(m[3]&m[184]&~m[185]&m[186]&~m[187])|(m[3]&~m[184]&m[185]&m[186]&~m[187])|(~m[3]&m[184]&m[185]&m[186]&~m[187])|(m[3]&m[184]&~m[185]&~m[186]&m[187])|(m[3]&~m[184]&m[185]&~m[186]&m[187])|(~m[3]&m[184]&m[185]&~m[186]&m[187])|(m[3]&~m[184]&~m[185]&m[186]&m[187])|(~m[3]&m[184]&~m[185]&m[186]&m[187])|(~m[3]&~m[184]&m[185]&m[186]&m[187]))&~BiasedRNG[283])|((m[3]&m[184]&m[185]&m[186]&~m[187])|(m[3]&m[184]&m[185]&~m[186]&m[187])|(m[3]&m[184]&~m[185]&m[186]&m[187])|(m[3]&~m[184]&m[185]&m[186]&m[187])|(~m[3]&m[184]&m[185]&m[186]&m[187])|(m[3]&m[184]&m[185]&m[186]&m[187]))):InitCond[492];
    m[68] = run?((((m[4]&m[198]&~m[199]&~m[200]&~m[201])|(m[4]&~m[198]&m[199]&~m[200]&~m[201])|(~m[4]&m[198]&m[199]&~m[200]&~m[201])|(m[4]&~m[198]&~m[199]&m[200]&~m[201])|(~m[4]&m[198]&~m[199]&m[200]&~m[201])|(~m[4]&~m[198]&m[199]&m[200]&~m[201])|(m[4]&~m[198]&~m[199]&~m[200]&m[201])|(~m[4]&m[198]&~m[199]&~m[200]&m[201])|(~m[4]&~m[198]&m[199]&~m[200]&m[201])|(~m[4]&~m[198]&~m[199]&m[200]&m[201]))&BiasedRNG[284])|(((m[4]&m[198]&m[199]&~m[200]&~m[201])|(m[4]&m[198]&~m[199]&m[200]&~m[201])|(m[4]&~m[198]&m[199]&m[200]&~m[201])|(~m[4]&m[198]&m[199]&m[200]&~m[201])|(m[4]&m[198]&~m[199]&~m[200]&m[201])|(m[4]&~m[198]&m[199]&~m[200]&m[201])|(~m[4]&m[198]&m[199]&~m[200]&m[201])|(m[4]&~m[198]&~m[199]&m[200]&m[201])|(~m[4]&m[198]&~m[199]&m[200]&m[201])|(~m[4]&~m[198]&m[199]&m[200]&m[201]))&~BiasedRNG[284])|((m[4]&m[198]&m[199]&m[200]&~m[201])|(m[4]&m[198]&m[199]&~m[200]&m[201])|(m[4]&m[198]&~m[199]&m[200]&m[201])|(m[4]&~m[198]&m[199]&m[200]&m[201])|(~m[4]&m[198]&m[199]&m[200]&m[201])|(m[4]&m[198]&m[199]&m[200]&m[201]))):InitCond[493];
    m[71] = run?((((m[5]&m[212]&~m[213]&~m[214]&~m[215])|(m[5]&~m[212]&m[213]&~m[214]&~m[215])|(~m[5]&m[212]&m[213]&~m[214]&~m[215])|(m[5]&~m[212]&~m[213]&m[214]&~m[215])|(~m[5]&m[212]&~m[213]&m[214]&~m[215])|(~m[5]&~m[212]&m[213]&m[214]&~m[215])|(m[5]&~m[212]&~m[213]&~m[214]&m[215])|(~m[5]&m[212]&~m[213]&~m[214]&m[215])|(~m[5]&~m[212]&m[213]&~m[214]&m[215])|(~m[5]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[285])|(((m[5]&m[212]&m[213]&~m[214]&~m[215])|(m[5]&m[212]&~m[213]&m[214]&~m[215])|(m[5]&~m[212]&m[213]&m[214]&~m[215])|(~m[5]&m[212]&m[213]&m[214]&~m[215])|(m[5]&m[212]&~m[213]&~m[214]&m[215])|(m[5]&~m[212]&m[213]&~m[214]&m[215])|(~m[5]&m[212]&m[213]&~m[214]&m[215])|(m[5]&~m[212]&~m[213]&m[214]&m[215])|(~m[5]&m[212]&~m[213]&m[214]&m[215])|(~m[5]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[285])|((m[5]&m[212]&m[213]&m[214]&~m[215])|(m[5]&m[212]&m[213]&~m[214]&m[215])|(m[5]&m[212]&~m[213]&m[214]&m[215])|(m[5]&~m[212]&m[213]&m[214]&m[215])|(~m[5]&m[212]&m[213]&m[214]&m[215])|(m[5]&m[212]&m[213]&m[214]&m[215]))):InitCond[494];
    m[74] = run?((((m[6]&m[226]&~m[227]&~m[228]&~m[229])|(m[6]&~m[226]&m[227]&~m[228]&~m[229])|(~m[6]&m[226]&m[227]&~m[228]&~m[229])|(m[6]&~m[226]&~m[227]&m[228]&~m[229])|(~m[6]&m[226]&~m[227]&m[228]&~m[229])|(~m[6]&~m[226]&m[227]&m[228]&~m[229])|(m[6]&~m[226]&~m[227]&~m[228]&m[229])|(~m[6]&m[226]&~m[227]&~m[228]&m[229])|(~m[6]&~m[226]&m[227]&~m[228]&m[229])|(~m[6]&~m[226]&~m[227]&m[228]&m[229]))&BiasedRNG[286])|(((m[6]&m[226]&m[227]&~m[228]&~m[229])|(m[6]&m[226]&~m[227]&m[228]&~m[229])|(m[6]&~m[226]&m[227]&m[228]&~m[229])|(~m[6]&m[226]&m[227]&m[228]&~m[229])|(m[6]&m[226]&~m[227]&~m[228]&m[229])|(m[6]&~m[226]&m[227]&~m[228]&m[229])|(~m[6]&m[226]&m[227]&~m[228]&m[229])|(m[6]&~m[226]&~m[227]&m[228]&m[229])|(~m[6]&m[226]&~m[227]&m[228]&m[229])|(~m[6]&~m[226]&m[227]&m[228]&m[229]))&~BiasedRNG[286])|((m[6]&m[226]&m[227]&m[228]&~m[229])|(m[6]&m[226]&m[227]&~m[228]&m[229])|(m[6]&m[226]&~m[227]&m[228]&m[229])|(m[6]&~m[226]&m[227]&m[228]&m[229])|(~m[6]&m[226]&m[227]&m[228]&m[229])|(m[6]&m[226]&m[227]&m[228]&m[229]))):InitCond[495];
    m[77] = run?((((m[7]&m[240]&~m[241]&~m[242]&~m[243])|(m[7]&~m[240]&m[241]&~m[242]&~m[243])|(~m[7]&m[240]&m[241]&~m[242]&~m[243])|(m[7]&~m[240]&~m[241]&m[242]&~m[243])|(~m[7]&m[240]&~m[241]&m[242]&~m[243])|(~m[7]&~m[240]&m[241]&m[242]&~m[243])|(m[7]&~m[240]&~m[241]&~m[242]&m[243])|(~m[7]&m[240]&~m[241]&~m[242]&m[243])|(~m[7]&~m[240]&m[241]&~m[242]&m[243])|(~m[7]&~m[240]&~m[241]&m[242]&m[243]))&BiasedRNG[287])|(((m[7]&m[240]&m[241]&~m[242]&~m[243])|(m[7]&m[240]&~m[241]&m[242]&~m[243])|(m[7]&~m[240]&m[241]&m[242]&~m[243])|(~m[7]&m[240]&m[241]&m[242]&~m[243])|(m[7]&m[240]&~m[241]&~m[242]&m[243])|(m[7]&~m[240]&m[241]&~m[242]&m[243])|(~m[7]&m[240]&m[241]&~m[242]&m[243])|(m[7]&~m[240]&~m[241]&m[242]&m[243])|(~m[7]&m[240]&~m[241]&m[242]&m[243])|(~m[7]&~m[240]&m[241]&m[242]&m[243]))&~BiasedRNG[287])|((m[7]&m[240]&m[241]&m[242]&~m[243])|(m[7]&m[240]&m[241]&~m[242]&m[243])|(m[7]&m[240]&~m[241]&m[242]&m[243])|(m[7]&~m[240]&m[241]&m[242]&m[243])|(~m[7]&m[240]&m[241]&m[242]&m[243])|(m[7]&m[240]&m[241]&m[242]&m[243]))):InitCond[496];
    m[80] = run?((((m[8]&m[254]&~m[255]&~m[256]&~m[257])|(m[8]&~m[254]&m[255]&~m[256]&~m[257])|(~m[8]&m[254]&m[255]&~m[256]&~m[257])|(m[8]&~m[254]&~m[255]&m[256]&~m[257])|(~m[8]&m[254]&~m[255]&m[256]&~m[257])|(~m[8]&~m[254]&m[255]&m[256]&~m[257])|(m[8]&~m[254]&~m[255]&~m[256]&m[257])|(~m[8]&m[254]&~m[255]&~m[256]&m[257])|(~m[8]&~m[254]&m[255]&~m[256]&m[257])|(~m[8]&~m[254]&~m[255]&m[256]&m[257]))&BiasedRNG[288])|(((m[8]&m[254]&m[255]&~m[256]&~m[257])|(m[8]&m[254]&~m[255]&m[256]&~m[257])|(m[8]&~m[254]&m[255]&m[256]&~m[257])|(~m[8]&m[254]&m[255]&m[256]&~m[257])|(m[8]&m[254]&~m[255]&~m[256]&m[257])|(m[8]&~m[254]&m[255]&~m[256]&m[257])|(~m[8]&m[254]&m[255]&~m[256]&m[257])|(m[8]&~m[254]&~m[255]&m[256]&m[257])|(~m[8]&m[254]&~m[255]&m[256]&m[257])|(~m[8]&~m[254]&m[255]&m[256]&m[257]))&~BiasedRNG[288])|((m[8]&m[254]&m[255]&m[256]&~m[257])|(m[8]&m[254]&m[255]&~m[256]&m[257])|(m[8]&m[254]&~m[255]&m[256]&m[257])|(m[8]&~m[254]&m[255]&m[256]&m[257])|(~m[8]&m[254]&m[255]&m[256]&m[257])|(m[8]&m[254]&m[255]&m[256]&m[257]))):InitCond[497];
    m[83] = run?((((m[9]&m[268]&~m[269]&~m[270]&~m[271])|(m[9]&~m[268]&m[269]&~m[270]&~m[271])|(~m[9]&m[268]&m[269]&~m[270]&~m[271])|(m[9]&~m[268]&~m[269]&m[270]&~m[271])|(~m[9]&m[268]&~m[269]&m[270]&~m[271])|(~m[9]&~m[268]&m[269]&m[270]&~m[271])|(m[9]&~m[268]&~m[269]&~m[270]&m[271])|(~m[9]&m[268]&~m[269]&~m[270]&m[271])|(~m[9]&~m[268]&m[269]&~m[270]&m[271])|(~m[9]&~m[268]&~m[269]&m[270]&m[271]))&BiasedRNG[289])|(((m[9]&m[268]&m[269]&~m[270]&~m[271])|(m[9]&m[268]&~m[269]&m[270]&~m[271])|(m[9]&~m[268]&m[269]&m[270]&~m[271])|(~m[9]&m[268]&m[269]&m[270]&~m[271])|(m[9]&m[268]&~m[269]&~m[270]&m[271])|(m[9]&~m[268]&m[269]&~m[270]&m[271])|(~m[9]&m[268]&m[269]&~m[270]&m[271])|(m[9]&~m[268]&~m[269]&m[270]&m[271])|(~m[9]&m[268]&~m[269]&m[270]&m[271])|(~m[9]&~m[268]&m[269]&m[270]&m[271]))&~BiasedRNG[289])|((m[9]&m[268]&m[269]&m[270]&~m[271])|(m[9]&m[268]&m[269]&~m[270]&m[271])|(m[9]&m[268]&~m[269]&m[270]&m[271])|(m[9]&~m[268]&m[269]&m[270]&m[271])|(~m[9]&m[268]&m[269]&m[270]&m[271])|(m[9]&m[268]&m[269]&m[270]&m[271]))):InitCond[498];
    m[86] = run?((((m[10]&m[282]&~m[283]&~m[284]&~m[285])|(m[10]&~m[282]&m[283]&~m[284]&~m[285])|(~m[10]&m[282]&m[283]&~m[284]&~m[285])|(m[10]&~m[282]&~m[283]&m[284]&~m[285])|(~m[10]&m[282]&~m[283]&m[284]&~m[285])|(~m[10]&~m[282]&m[283]&m[284]&~m[285])|(m[10]&~m[282]&~m[283]&~m[284]&m[285])|(~m[10]&m[282]&~m[283]&~m[284]&m[285])|(~m[10]&~m[282]&m[283]&~m[284]&m[285])|(~m[10]&~m[282]&~m[283]&m[284]&m[285]))&BiasedRNG[290])|(((m[10]&m[282]&m[283]&~m[284]&~m[285])|(m[10]&m[282]&~m[283]&m[284]&~m[285])|(m[10]&~m[282]&m[283]&m[284]&~m[285])|(~m[10]&m[282]&m[283]&m[284]&~m[285])|(m[10]&m[282]&~m[283]&~m[284]&m[285])|(m[10]&~m[282]&m[283]&~m[284]&m[285])|(~m[10]&m[282]&m[283]&~m[284]&m[285])|(m[10]&~m[282]&~m[283]&m[284]&m[285])|(~m[10]&m[282]&~m[283]&m[284]&m[285])|(~m[10]&~m[282]&m[283]&m[284]&m[285]))&~BiasedRNG[290])|((m[10]&m[282]&m[283]&m[284]&~m[285])|(m[10]&m[282]&m[283]&~m[284]&m[285])|(m[10]&m[282]&~m[283]&m[284]&m[285])|(m[10]&~m[282]&m[283]&m[284]&m[285])|(~m[10]&m[282]&m[283]&m[284]&m[285])|(m[10]&m[282]&m[283]&m[284]&m[285]))):InitCond[499];
    m[89] = run?((((m[11]&m[296]&~m[297]&~m[298]&~m[299])|(m[11]&~m[296]&m[297]&~m[298]&~m[299])|(~m[11]&m[296]&m[297]&~m[298]&~m[299])|(m[11]&~m[296]&~m[297]&m[298]&~m[299])|(~m[11]&m[296]&~m[297]&m[298]&~m[299])|(~m[11]&~m[296]&m[297]&m[298]&~m[299])|(m[11]&~m[296]&~m[297]&~m[298]&m[299])|(~m[11]&m[296]&~m[297]&~m[298]&m[299])|(~m[11]&~m[296]&m[297]&~m[298]&m[299])|(~m[11]&~m[296]&~m[297]&m[298]&m[299]))&BiasedRNG[291])|(((m[11]&m[296]&m[297]&~m[298]&~m[299])|(m[11]&m[296]&~m[297]&m[298]&~m[299])|(m[11]&~m[296]&m[297]&m[298]&~m[299])|(~m[11]&m[296]&m[297]&m[298]&~m[299])|(m[11]&m[296]&~m[297]&~m[298]&m[299])|(m[11]&~m[296]&m[297]&~m[298]&m[299])|(~m[11]&m[296]&m[297]&~m[298]&m[299])|(m[11]&~m[296]&~m[297]&m[298]&m[299])|(~m[11]&m[296]&~m[297]&m[298]&m[299])|(~m[11]&~m[296]&m[297]&m[298]&m[299]))&~BiasedRNG[291])|((m[11]&m[296]&m[297]&m[298]&~m[299])|(m[11]&m[296]&m[297]&~m[298]&m[299])|(m[11]&m[296]&~m[297]&m[298]&m[299])|(m[11]&~m[296]&m[297]&m[298]&m[299])|(~m[11]&m[296]&m[297]&m[298]&m[299])|(m[11]&m[296]&m[297]&m[298]&m[299]))):InitCond[500];
    m[92] = run?((((m[12]&m[310]&~m[311]&~m[312]&~m[313])|(m[12]&~m[310]&m[311]&~m[312]&~m[313])|(~m[12]&m[310]&m[311]&~m[312]&~m[313])|(m[12]&~m[310]&~m[311]&m[312]&~m[313])|(~m[12]&m[310]&~m[311]&m[312]&~m[313])|(~m[12]&~m[310]&m[311]&m[312]&~m[313])|(m[12]&~m[310]&~m[311]&~m[312]&m[313])|(~m[12]&m[310]&~m[311]&~m[312]&m[313])|(~m[12]&~m[310]&m[311]&~m[312]&m[313])|(~m[12]&~m[310]&~m[311]&m[312]&m[313]))&BiasedRNG[292])|(((m[12]&m[310]&m[311]&~m[312]&~m[313])|(m[12]&m[310]&~m[311]&m[312]&~m[313])|(m[12]&~m[310]&m[311]&m[312]&~m[313])|(~m[12]&m[310]&m[311]&m[312]&~m[313])|(m[12]&m[310]&~m[311]&~m[312]&m[313])|(m[12]&~m[310]&m[311]&~m[312]&m[313])|(~m[12]&m[310]&m[311]&~m[312]&m[313])|(m[12]&~m[310]&~m[311]&m[312]&m[313])|(~m[12]&m[310]&~m[311]&m[312]&m[313])|(~m[12]&~m[310]&m[311]&m[312]&m[313]))&~BiasedRNG[292])|((m[12]&m[310]&m[311]&m[312]&~m[313])|(m[12]&m[310]&m[311]&~m[312]&m[313])|(m[12]&m[310]&~m[311]&m[312]&m[313])|(m[12]&~m[310]&m[311]&m[312]&m[313])|(~m[12]&m[310]&m[311]&m[312]&m[313])|(m[12]&m[310]&m[311]&m[312]&m[313]))):InitCond[501];
    m[95] = run?((((m[13]&m[324]&~m[325]&~m[326]&~m[327])|(m[13]&~m[324]&m[325]&~m[326]&~m[327])|(~m[13]&m[324]&m[325]&~m[326]&~m[327])|(m[13]&~m[324]&~m[325]&m[326]&~m[327])|(~m[13]&m[324]&~m[325]&m[326]&~m[327])|(~m[13]&~m[324]&m[325]&m[326]&~m[327])|(m[13]&~m[324]&~m[325]&~m[326]&m[327])|(~m[13]&m[324]&~m[325]&~m[326]&m[327])|(~m[13]&~m[324]&m[325]&~m[326]&m[327])|(~m[13]&~m[324]&~m[325]&m[326]&m[327]))&BiasedRNG[293])|(((m[13]&m[324]&m[325]&~m[326]&~m[327])|(m[13]&m[324]&~m[325]&m[326]&~m[327])|(m[13]&~m[324]&m[325]&m[326]&~m[327])|(~m[13]&m[324]&m[325]&m[326]&~m[327])|(m[13]&m[324]&~m[325]&~m[326]&m[327])|(m[13]&~m[324]&m[325]&~m[326]&m[327])|(~m[13]&m[324]&m[325]&~m[326]&m[327])|(m[13]&~m[324]&~m[325]&m[326]&m[327])|(~m[13]&m[324]&~m[325]&m[326]&m[327])|(~m[13]&~m[324]&m[325]&m[326]&m[327]))&~BiasedRNG[293])|((m[13]&m[324]&m[325]&m[326]&~m[327])|(m[13]&m[324]&m[325]&~m[326]&m[327])|(m[13]&m[324]&~m[325]&m[326]&m[327])|(m[13]&~m[324]&m[325]&m[326]&m[327])|(~m[13]&m[324]&m[325]&m[326]&m[327])|(m[13]&m[324]&m[325]&m[326]&m[327]))):InitCond[502];
    m[98] = run?((((m[14]&m[338]&~m[339]&~m[340]&~m[341])|(m[14]&~m[338]&m[339]&~m[340]&~m[341])|(~m[14]&m[338]&m[339]&~m[340]&~m[341])|(m[14]&~m[338]&~m[339]&m[340]&~m[341])|(~m[14]&m[338]&~m[339]&m[340]&~m[341])|(~m[14]&~m[338]&m[339]&m[340]&~m[341])|(m[14]&~m[338]&~m[339]&~m[340]&m[341])|(~m[14]&m[338]&~m[339]&~m[340]&m[341])|(~m[14]&~m[338]&m[339]&~m[340]&m[341])|(~m[14]&~m[338]&~m[339]&m[340]&m[341]))&BiasedRNG[294])|(((m[14]&m[338]&m[339]&~m[340]&~m[341])|(m[14]&m[338]&~m[339]&m[340]&~m[341])|(m[14]&~m[338]&m[339]&m[340]&~m[341])|(~m[14]&m[338]&m[339]&m[340]&~m[341])|(m[14]&m[338]&~m[339]&~m[340]&m[341])|(m[14]&~m[338]&m[339]&~m[340]&m[341])|(~m[14]&m[338]&m[339]&~m[340]&m[341])|(m[14]&~m[338]&~m[339]&m[340]&m[341])|(~m[14]&m[338]&~m[339]&m[340]&m[341])|(~m[14]&~m[338]&m[339]&m[340]&m[341]))&~BiasedRNG[294])|((m[14]&m[338]&m[339]&m[340]&~m[341])|(m[14]&m[338]&m[339]&~m[340]&m[341])|(m[14]&m[338]&~m[339]&m[340]&m[341])|(m[14]&~m[338]&m[339]&m[340]&m[341])|(~m[14]&m[338]&m[339]&m[340]&m[341])|(m[14]&m[338]&m[339]&m[340]&m[341]))):InitCond[503];
    m[101] = run?((((m[15]&m[352]&~m[353]&~m[354]&~m[355])|(m[15]&~m[352]&m[353]&~m[354]&~m[355])|(~m[15]&m[352]&m[353]&~m[354]&~m[355])|(m[15]&~m[352]&~m[353]&m[354]&~m[355])|(~m[15]&m[352]&~m[353]&m[354]&~m[355])|(~m[15]&~m[352]&m[353]&m[354]&~m[355])|(m[15]&~m[352]&~m[353]&~m[354]&m[355])|(~m[15]&m[352]&~m[353]&~m[354]&m[355])|(~m[15]&~m[352]&m[353]&~m[354]&m[355])|(~m[15]&~m[352]&~m[353]&m[354]&m[355]))&BiasedRNG[295])|(((m[15]&m[352]&m[353]&~m[354]&~m[355])|(m[15]&m[352]&~m[353]&m[354]&~m[355])|(m[15]&~m[352]&m[353]&m[354]&~m[355])|(~m[15]&m[352]&m[353]&m[354]&~m[355])|(m[15]&m[352]&~m[353]&~m[354]&m[355])|(m[15]&~m[352]&m[353]&~m[354]&m[355])|(~m[15]&m[352]&m[353]&~m[354]&m[355])|(m[15]&~m[352]&~m[353]&m[354]&m[355])|(~m[15]&m[352]&~m[353]&m[354]&m[355])|(~m[15]&~m[352]&m[353]&m[354]&m[355]))&~BiasedRNG[295])|((m[15]&m[352]&m[353]&m[354]&~m[355])|(m[15]&m[352]&m[353]&~m[354]&m[355])|(m[15]&m[352]&~m[353]&m[354]&m[355])|(m[15]&~m[352]&m[353]&m[354]&m[355])|(~m[15]&m[352]&m[353]&m[354]&m[355])|(m[15]&m[352]&m[353]&m[354]&m[355]))):InitCond[504];
    m[104] = run?((((m[16]&m[366]&~m[367]&~m[368]&~m[369])|(m[16]&~m[366]&m[367]&~m[368]&~m[369])|(~m[16]&m[366]&m[367]&~m[368]&~m[369])|(m[16]&~m[366]&~m[367]&m[368]&~m[369])|(~m[16]&m[366]&~m[367]&m[368]&~m[369])|(~m[16]&~m[366]&m[367]&m[368]&~m[369])|(m[16]&~m[366]&~m[367]&~m[368]&m[369])|(~m[16]&m[366]&~m[367]&~m[368]&m[369])|(~m[16]&~m[366]&m[367]&~m[368]&m[369])|(~m[16]&~m[366]&~m[367]&m[368]&m[369]))&BiasedRNG[296])|(((m[16]&m[366]&m[367]&~m[368]&~m[369])|(m[16]&m[366]&~m[367]&m[368]&~m[369])|(m[16]&~m[366]&m[367]&m[368]&~m[369])|(~m[16]&m[366]&m[367]&m[368]&~m[369])|(m[16]&m[366]&~m[367]&~m[368]&m[369])|(m[16]&~m[366]&m[367]&~m[368]&m[369])|(~m[16]&m[366]&m[367]&~m[368]&m[369])|(m[16]&~m[366]&~m[367]&m[368]&m[369])|(~m[16]&m[366]&~m[367]&m[368]&m[369])|(~m[16]&~m[366]&m[367]&m[368]&m[369]))&~BiasedRNG[296])|((m[16]&m[366]&m[367]&m[368]&~m[369])|(m[16]&m[366]&m[367]&~m[368]&m[369])|(m[16]&m[366]&~m[367]&m[368]&m[369])|(m[16]&~m[366]&m[367]&m[368]&m[369])|(~m[16]&m[366]&m[367]&m[368]&m[369])|(m[16]&m[366]&m[367]&m[368]&m[369]))):InitCond[505];
    m[107] = run?((((m[17]&m[380]&~m[381]&~m[382]&~m[383])|(m[17]&~m[380]&m[381]&~m[382]&~m[383])|(~m[17]&m[380]&m[381]&~m[382]&~m[383])|(m[17]&~m[380]&~m[381]&m[382]&~m[383])|(~m[17]&m[380]&~m[381]&m[382]&~m[383])|(~m[17]&~m[380]&m[381]&m[382]&~m[383])|(m[17]&~m[380]&~m[381]&~m[382]&m[383])|(~m[17]&m[380]&~m[381]&~m[382]&m[383])|(~m[17]&~m[380]&m[381]&~m[382]&m[383])|(~m[17]&~m[380]&~m[381]&m[382]&m[383]))&BiasedRNG[297])|(((m[17]&m[380]&m[381]&~m[382]&~m[383])|(m[17]&m[380]&~m[381]&m[382]&~m[383])|(m[17]&~m[380]&m[381]&m[382]&~m[383])|(~m[17]&m[380]&m[381]&m[382]&~m[383])|(m[17]&m[380]&~m[381]&~m[382]&m[383])|(m[17]&~m[380]&m[381]&~m[382]&m[383])|(~m[17]&m[380]&m[381]&~m[382]&m[383])|(m[17]&~m[380]&~m[381]&m[382]&m[383])|(~m[17]&m[380]&~m[381]&m[382]&m[383])|(~m[17]&~m[380]&m[381]&m[382]&m[383]))&~BiasedRNG[297])|((m[17]&m[380]&m[381]&m[382]&~m[383])|(m[17]&m[380]&m[381]&~m[382]&m[383])|(m[17]&m[380]&~m[381]&m[382]&m[383])|(m[17]&~m[380]&m[381]&m[382]&m[383])|(~m[17]&m[380]&m[381]&m[382]&m[383])|(m[17]&m[380]&m[381]&m[382]&m[383]))):InitCond[506];
    m[110] = run?((((m[18]&m[394]&~m[395]&~m[396]&~m[397])|(m[18]&~m[394]&m[395]&~m[396]&~m[397])|(~m[18]&m[394]&m[395]&~m[396]&~m[397])|(m[18]&~m[394]&~m[395]&m[396]&~m[397])|(~m[18]&m[394]&~m[395]&m[396]&~m[397])|(~m[18]&~m[394]&m[395]&m[396]&~m[397])|(m[18]&~m[394]&~m[395]&~m[396]&m[397])|(~m[18]&m[394]&~m[395]&~m[396]&m[397])|(~m[18]&~m[394]&m[395]&~m[396]&m[397])|(~m[18]&~m[394]&~m[395]&m[396]&m[397]))&BiasedRNG[298])|(((m[18]&m[394]&m[395]&~m[396]&~m[397])|(m[18]&m[394]&~m[395]&m[396]&~m[397])|(m[18]&~m[394]&m[395]&m[396]&~m[397])|(~m[18]&m[394]&m[395]&m[396]&~m[397])|(m[18]&m[394]&~m[395]&~m[396]&m[397])|(m[18]&~m[394]&m[395]&~m[396]&m[397])|(~m[18]&m[394]&m[395]&~m[396]&m[397])|(m[18]&~m[394]&~m[395]&m[396]&m[397])|(~m[18]&m[394]&~m[395]&m[396]&m[397])|(~m[18]&~m[394]&m[395]&m[396]&m[397]))&~BiasedRNG[298])|((m[18]&m[394]&m[395]&m[396]&~m[397])|(m[18]&m[394]&m[395]&~m[396]&m[397])|(m[18]&m[394]&~m[395]&m[396]&m[397])|(m[18]&~m[394]&m[395]&m[396]&m[397])|(~m[18]&m[394]&m[395]&m[396]&m[397])|(m[18]&m[394]&m[395]&m[396]&m[397]))):InitCond[507];
    m[113] = run?((((m[19]&m[408]&~m[409]&~m[410]&~m[411])|(m[19]&~m[408]&m[409]&~m[410]&~m[411])|(~m[19]&m[408]&m[409]&~m[410]&~m[411])|(m[19]&~m[408]&~m[409]&m[410]&~m[411])|(~m[19]&m[408]&~m[409]&m[410]&~m[411])|(~m[19]&~m[408]&m[409]&m[410]&~m[411])|(m[19]&~m[408]&~m[409]&~m[410]&m[411])|(~m[19]&m[408]&~m[409]&~m[410]&m[411])|(~m[19]&~m[408]&m[409]&~m[410]&m[411])|(~m[19]&~m[408]&~m[409]&m[410]&m[411]))&BiasedRNG[299])|(((m[19]&m[408]&m[409]&~m[410]&~m[411])|(m[19]&m[408]&~m[409]&m[410]&~m[411])|(m[19]&~m[408]&m[409]&m[410]&~m[411])|(~m[19]&m[408]&m[409]&m[410]&~m[411])|(m[19]&m[408]&~m[409]&~m[410]&m[411])|(m[19]&~m[408]&m[409]&~m[410]&m[411])|(~m[19]&m[408]&m[409]&~m[410]&m[411])|(m[19]&~m[408]&~m[409]&m[410]&m[411])|(~m[19]&m[408]&~m[409]&m[410]&m[411])|(~m[19]&~m[408]&m[409]&m[410]&m[411]))&~BiasedRNG[299])|((m[19]&m[408]&m[409]&m[410]&~m[411])|(m[19]&m[408]&m[409]&~m[410]&m[411])|(m[19]&m[408]&~m[409]&m[410]&m[411])|(m[19]&~m[408]&m[409]&m[410]&m[411])|(~m[19]&m[408]&m[409]&m[410]&m[411])|(m[19]&m[408]&m[409]&m[410]&m[411]))):InitCond[508];
    m[116] = run?((((m[20]&m[422]&~m[423]&~m[424]&~m[425])|(m[20]&~m[422]&m[423]&~m[424]&~m[425])|(~m[20]&m[422]&m[423]&~m[424]&~m[425])|(m[20]&~m[422]&~m[423]&m[424]&~m[425])|(~m[20]&m[422]&~m[423]&m[424]&~m[425])|(~m[20]&~m[422]&m[423]&m[424]&~m[425])|(m[20]&~m[422]&~m[423]&~m[424]&m[425])|(~m[20]&m[422]&~m[423]&~m[424]&m[425])|(~m[20]&~m[422]&m[423]&~m[424]&m[425])|(~m[20]&~m[422]&~m[423]&m[424]&m[425]))&BiasedRNG[300])|(((m[20]&m[422]&m[423]&~m[424]&~m[425])|(m[20]&m[422]&~m[423]&m[424]&~m[425])|(m[20]&~m[422]&m[423]&m[424]&~m[425])|(~m[20]&m[422]&m[423]&m[424]&~m[425])|(m[20]&m[422]&~m[423]&~m[424]&m[425])|(m[20]&~m[422]&m[423]&~m[424]&m[425])|(~m[20]&m[422]&m[423]&~m[424]&m[425])|(m[20]&~m[422]&~m[423]&m[424]&m[425])|(~m[20]&m[422]&~m[423]&m[424]&m[425])|(~m[20]&~m[422]&m[423]&m[424]&m[425]))&~BiasedRNG[300])|((m[20]&m[422]&m[423]&m[424]&~m[425])|(m[20]&m[422]&m[423]&~m[424]&m[425])|(m[20]&m[422]&~m[423]&m[424]&m[425])|(m[20]&~m[422]&m[423]&m[424]&m[425])|(~m[20]&m[422]&m[423]&m[424]&m[425])|(m[20]&m[422]&m[423]&m[424]&m[425]))):InitCond[509];
    m[119] = run?((((m[21]&m[436]&~m[437]&~m[438]&~m[439])|(m[21]&~m[436]&m[437]&~m[438]&~m[439])|(~m[21]&m[436]&m[437]&~m[438]&~m[439])|(m[21]&~m[436]&~m[437]&m[438]&~m[439])|(~m[21]&m[436]&~m[437]&m[438]&~m[439])|(~m[21]&~m[436]&m[437]&m[438]&~m[439])|(m[21]&~m[436]&~m[437]&~m[438]&m[439])|(~m[21]&m[436]&~m[437]&~m[438]&m[439])|(~m[21]&~m[436]&m[437]&~m[438]&m[439])|(~m[21]&~m[436]&~m[437]&m[438]&m[439]))&BiasedRNG[301])|(((m[21]&m[436]&m[437]&~m[438]&~m[439])|(m[21]&m[436]&~m[437]&m[438]&~m[439])|(m[21]&~m[436]&m[437]&m[438]&~m[439])|(~m[21]&m[436]&m[437]&m[438]&~m[439])|(m[21]&m[436]&~m[437]&~m[438]&m[439])|(m[21]&~m[436]&m[437]&~m[438]&m[439])|(~m[21]&m[436]&m[437]&~m[438]&m[439])|(m[21]&~m[436]&~m[437]&m[438]&m[439])|(~m[21]&m[436]&~m[437]&m[438]&m[439])|(~m[21]&~m[436]&m[437]&m[438]&m[439]))&~BiasedRNG[301])|((m[21]&m[436]&m[437]&m[438]&~m[439])|(m[21]&m[436]&m[437]&~m[438]&m[439])|(m[21]&m[436]&~m[437]&m[438]&m[439])|(m[21]&~m[436]&m[437]&m[438]&m[439])|(~m[21]&m[436]&m[437]&m[438]&m[439])|(m[21]&m[436]&m[437]&m[438]&m[439]))):InitCond[510];
    m[122] = run?((((m[22]&m[450]&~m[451]&~m[452]&~m[453])|(m[22]&~m[450]&m[451]&~m[452]&~m[453])|(~m[22]&m[450]&m[451]&~m[452]&~m[453])|(m[22]&~m[450]&~m[451]&m[452]&~m[453])|(~m[22]&m[450]&~m[451]&m[452]&~m[453])|(~m[22]&~m[450]&m[451]&m[452]&~m[453])|(m[22]&~m[450]&~m[451]&~m[452]&m[453])|(~m[22]&m[450]&~m[451]&~m[452]&m[453])|(~m[22]&~m[450]&m[451]&~m[452]&m[453])|(~m[22]&~m[450]&~m[451]&m[452]&m[453]))&BiasedRNG[302])|(((m[22]&m[450]&m[451]&~m[452]&~m[453])|(m[22]&m[450]&~m[451]&m[452]&~m[453])|(m[22]&~m[450]&m[451]&m[452]&~m[453])|(~m[22]&m[450]&m[451]&m[452]&~m[453])|(m[22]&m[450]&~m[451]&~m[452]&m[453])|(m[22]&~m[450]&m[451]&~m[452]&m[453])|(~m[22]&m[450]&m[451]&~m[452]&m[453])|(m[22]&~m[450]&~m[451]&m[452]&m[453])|(~m[22]&m[450]&~m[451]&m[452]&m[453])|(~m[22]&~m[450]&m[451]&m[452]&m[453]))&~BiasedRNG[302])|((m[22]&m[450]&m[451]&m[452]&~m[453])|(m[22]&m[450]&m[451]&~m[452]&m[453])|(m[22]&m[450]&~m[451]&m[452]&m[453])|(m[22]&~m[450]&m[451]&m[452]&m[453])|(~m[22]&m[450]&m[451]&m[452]&m[453])|(m[22]&m[450]&m[451]&m[452]&m[453]))):InitCond[511];
    m[125] = run?((((m[23]&m[464]&~m[465]&~m[466]&~m[467])|(m[23]&~m[464]&m[465]&~m[466]&~m[467])|(~m[23]&m[464]&m[465]&~m[466]&~m[467])|(m[23]&~m[464]&~m[465]&m[466]&~m[467])|(~m[23]&m[464]&~m[465]&m[466]&~m[467])|(~m[23]&~m[464]&m[465]&m[466]&~m[467])|(m[23]&~m[464]&~m[465]&~m[466]&m[467])|(~m[23]&m[464]&~m[465]&~m[466]&m[467])|(~m[23]&~m[464]&m[465]&~m[466]&m[467])|(~m[23]&~m[464]&~m[465]&m[466]&m[467]))&BiasedRNG[303])|(((m[23]&m[464]&m[465]&~m[466]&~m[467])|(m[23]&m[464]&~m[465]&m[466]&~m[467])|(m[23]&~m[464]&m[465]&m[466]&~m[467])|(~m[23]&m[464]&m[465]&m[466]&~m[467])|(m[23]&m[464]&~m[465]&~m[466]&m[467])|(m[23]&~m[464]&m[465]&~m[466]&m[467])|(~m[23]&m[464]&m[465]&~m[466]&m[467])|(m[23]&~m[464]&~m[465]&m[466]&m[467])|(~m[23]&m[464]&~m[465]&m[466]&m[467])|(~m[23]&~m[464]&m[465]&m[466]&m[467]))&~BiasedRNG[303])|((m[23]&m[464]&m[465]&m[466]&~m[467])|(m[23]&m[464]&m[465]&~m[466]&m[467])|(m[23]&m[464]&~m[465]&m[466]&m[467])|(m[23]&~m[464]&m[465]&m[466]&m[467])|(~m[23]&m[464]&m[465]&m[466]&m[467])|(m[23]&m[464]&m[465]&m[466]&m[467]))):InitCond[512];
    m[128] = run?((((m[24]&m[478]&~m[479]&~m[480]&~m[481])|(m[24]&~m[478]&m[479]&~m[480]&~m[481])|(~m[24]&m[478]&m[479]&~m[480]&~m[481])|(m[24]&~m[478]&~m[479]&m[480]&~m[481])|(~m[24]&m[478]&~m[479]&m[480]&~m[481])|(~m[24]&~m[478]&m[479]&m[480]&~m[481])|(m[24]&~m[478]&~m[479]&~m[480]&m[481])|(~m[24]&m[478]&~m[479]&~m[480]&m[481])|(~m[24]&~m[478]&m[479]&~m[480]&m[481])|(~m[24]&~m[478]&~m[479]&m[480]&m[481]))&BiasedRNG[304])|(((m[24]&m[478]&m[479]&~m[480]&~m[481])|(m[24]&m[478]&~m[479]&m[480]&~m[481])|(m[24]&~m[478]&m[479]&m[480]&~m[481])|(~m[24]&m[478]&m[479]&m[480]&~m[481])|(m[24]&m[478]&~m[479]&~m[480]&m[481])|(m[24]&~m[478]&m[479]&~m[480]&m[481])|(~m[24]&m[478]&m[479]&~m[480]&m[481])|(m[24]&~m[478]&~m[479]&m[480]&m[481])|(~m[24]&m[478]&~m[479]&m[480]&m[481])|(~m[24]&~m[478]&m[479]&m[480]&m[481]))&~BiasedRNG[304])|((m[24]&m[478]&m[479]&m[480]&~m[481])|(m[24]&m[478]&m[479]&~m[480]&m[481])|(m[24]&m[478]&~m[479]&m[480]&m[481])|(m[24]&~m[478]&m[479]&m[480]&m[481])|(~m[24]&m[478]&m[479]&m[480]&m[481])|(m[24]&m[478]&m[479]&m[480]&m[481]))):InitCond[513];
    m[131] = run?((((m[25]&m[492]&~m[493]&~m[494]&~m[495])|(m[25]&~m[492]&m[493]&~m[494]&~m[495])|(~m[25]&m[492]&m[493]&~m[494]&~m[495])|(m[25]&~m[492]&~m[493]&m[494]&~m[495])|(~m[25]&m[492]&~m[493]&m[494]&~m[495])|(~m[25]&~m[492]&m[493]&m[494]&~m[495])|(m[25]&~m[492]&~m[493]&~m[494]&m[495])|(~m[25]&m[492]&~m[493]&~m[494]&m[495])|(~m[25]&~m[492]&m[493]&~m[494]&m[495])|(~m[25]&~m[492]&~m[493]&m[494]&m[495]))&BiasedRNG[305])|(((m[25]&m[492]&m[493]&~m[494]&~m[495])|(m[25]&m[492]&~m[493]&m[494]&~m[495])|(m[25]&~m[492]&m[493]&m[494]&~m[495])|(~m[25]&m[492]&m[493]&m[494]&~m[495])|(m[25]&m[492]&~m[493]&~m[494]&m[495])|(m[25]&~m[492]&m[493]&~m[494]&m[495])|(~m[25]&m[492]&m[493]&~m[494]&m[495])|(m[25]&~m[492]&~m[493]&m[494]&m[495])|(~m[25]&m[492]&~m[493]&m[494]&m[495])|(~m[25]&~m[492]&m[493]&m[494]&m[495]))&~BiasedRNG[305])|((m[25]&m[492]&m[493]&m[494]&~m[495])|(m[25]&m[492]&m[493]&~m[494]&m[495])|(m[25]&m[492]&~m[493]&m[494]&m[495])|(m[25]&~m[492]&m[493]&m[494]&m[495])|(~m[25]&m[492]&m[493]&m[494]&m[495])|(m[25]&m[492]&m[493]&m[494]&m[495]))):InitCond[514];
    m[134] = run?((((m[26]&m[506]&~m[507]&~m[508]&~m[509])|(m[26]&~m[506]&m[507]&~m[508]&~m[509])|(~m[26]&m[506]&m[507]&~m[508]&~m[509])|(m[26]&~m[506]&~m[507]&m[508]&~m[509])|(~m[26]&m[506]&~m[507]&m[508]&~m[509])|(~m[26]&~m[506]&m[507]&m[508]&~m[509])|(m[26]&~m[506]&~m[507]&~m[508]&m[509])|(~m[26]&m[506]&~m[507]&~m[508]&m[509])|(~m[26]&~m[506]&m[507]&~m[508]&m[509])|(~m[26]&~m[506]&~m[507]&m[508]&m[509]))&BiasedRNG[306])|(((m[26]&m[506]&m[507]&~m[508]&~m[509])|(m[26]&m[506]&~m[507]&m[508]&~m[509])|(m[26]&~m[506]&m[507]&m[508]&~m[509])|(~m[26]&m[506]&m[507]&m[508]&~m[509])|(m[26]&m[506]&~m[507]&~m[508]&m[509])|(m[26]&~m[506]&m[507]&~m[508]&m[509])|(~m[26]&m[506]&m[507]&~m[508]&m[509])|(m[26]&~m[506]&~m[507]&m[508]&m[509])|(~m[26]&m[506]&~m[507]&m[508]&m[509])|(~m[26]&~m[506]&m[507]&m[508]&m[509]))&~BiasedRNG[306])|((m[26]&m[506]&m[507]&m[508]&~m[509])|(m[26]&m[506]&m[507]&~m[508]&m[509])|(m[26]&m[506]&~m[507]&m[508]&m[509])|(m[26]&~m[506]&m[507]&m[508]&m[509])|(~m[26]&m[506]&m[507]&m[508]&m[509])|(m[26]&m[506]&m[507]&m[508]&m[509]))):InitCond[515];
    m[137] = run?((((m[27]&m[520]&~m[521]&~m[522]&~m[523])|(m[27]&~m[520]&m[521]&~m[522]&~m[523])|(~m[27]&m[520]&m[521]&~m[522]&~m[523])|(m[27]&~m[520]&~m[521]&m[522]&~m[523])|(~m[27]&m[520]&~m[521]&m[522]&~m[523])|(~m[27]&~m[520]&m[521]&m[522]&~m[523])|(m[27]&~m[520]&~m[521]&~m[522]&m[523])|(~m[27]&m[520]&~m[521]&~m[522]&m[523])|(~m[27]&~m[520]&m[521]&~m[522]&m[523])|(~m[27]&~m[520]&~m[521]&m[522]&m[523]))&BiasedRNG[307])|(((m[27]&m[520]&m[521]&~m[522]&~m[523])|(m[27]&m[520]&~m[521]&m[522]&~m[523])|(m[27]&~m[520]&m[521]&m[522]&~m[523])|(~m[27]&m[520]&m[521]&m[522]&~m[523])|(m[27]&m[520]&~m[521]&~m[522]&m[523])|(m[27]&~m[520]&m[521]&~m[522]&m[523])|(~m[27]&m[520]&m[521]&~m[522]&m[523])|(m[27]&~m[520]&~m[521]&m[522]&m[523])|(~m[27]&m[520]&~m[521]&m[522]&m[523])|(~m[27]&~m[520]&m[521]&m[522]&m[523]))&~BiasedRNG[307])|((m[27]&m[520]&m[521]&m[522]&~m[523])|(m[27]&m[520]&m[521]&~m[522]&m[523])|(m[27]&m[520]&~m[521]&m[522]&m[523])|(m[27]&~m[520]&m[521]&m[522]&m[523])|(~m[27]&m[520]&m[521]&m[522]&m[523])|(m[27]&m[520]&m[521]&m[522]&m[523]))):InitCond[516];
    m[146] = run?((((~m[57]&~m[420]&~m[616])|(m[57]&m[420]&~m[616]))&BiasedRNG[308])|(((m[57]&~m[420]&~m[616])|(~m[57]&m[420]&m[616]))&~BiasedRNG[308])|((~m[57]&~m[420]&m[616])|(m[57]&~m[420]&m[616])|(m[57]&m[420]&m[616]))):InitCond[517];
    m[147] = run?((((~m[57]&~m[434]&~m[630])|(m[57]&m[434]&~m[630]))&BiasedRNG[309])|(((m[57]&~m[434]&~m[630])|(~m[57]&m[434]&m[630]))&~BiasedRNG[309])|((~m[57]&~m[434]&m[630])|(m[57]&~m[434]&m[630])|(m[57]&m[434]&m[630]))):InitCond[518];
    m[148] = run?((((~m[57]&~m[448]&~m[644])|(m[57]&m[448]&~m[644]))&BiasedRNG[310])|(((m[57]&~m[448]&~m[644])|(~m[57]&m[448]&m[644]))&~BiasedRNG[310])|((~m[57]&~m[448]&m[644])|(m[57]&~m[448]&m[644])|(m[57]&m[448]&m[644]))):InitCond[519];
    m[149] = run?((((~m[57]&~m[462]&~m[658])|(m[57]&m[462]&~m[658]))&BiasedRNG[311])|(((m[57]&~m[462]&~m[658])|(~m[57]&m[462]&m[658]))&~BiasedRNG[311])|((~m[57]&~m[462]&m[658])|(m[57]&~m[462]&m[658])|(m[57]&m[462]&m[658]))):InitCond[520];
    m[150] = run?((((~m[58]&~m[476]&~m[672])|(m[58]&m[476]&~m[672]))&BiasedRNG[312])|(((m[58]&~m[476]&~m[672])|(~m[58]&m[476]&m[672]))&~BiasedRNG[312])|((~m[58]&~m[476]&m[672])|(m[58]&~m[476]&m[672])|(m[58]&m[476]&m[672]))):InitCond[521];
    m[151] = run?((((~m[58]&~m[490]&~m[686])|(m[58]&m[490]&~m[686]))&BiasedRNG[313])|(((m[58]&~m[490]&~m[686])|(~m[58]&m[490]&m[686]))&~BiasedRNG[313])|((~m[58]&~m[490]&m[686])|(m[58]&~m[490]&m[686])|(m[58]&m[490]&m[686]))):InitCond[522];
    m[152] = run?((((~m[58]&~m[504]&~m[700])|(m[58]&m[504]&~m[700]))&BiasedRNG[314])|(((m[58]&~m[504]&~m[700])|(~m[58]&m[504]&m[700]))&~BiasedRNG[314])|((~m[58]&~m[504]&m[700])|(m[58]&~m[504]&m[700])|(m[58]&m[504]&m[700]))):InitCond[523];
    m[153] = run?((((~m[58]&~m[518]&~m[714])|(m[58]&m[518]&~m[714]))&BiasedRNG[315])|(((m[58]&~m[518]&~m[714])|(~m[58]&m[518]&m[714]))&~BiasedRNG[315])|((~m[58]&~m[518]&m[714])|(m[58]&~m[518]&m[714])|(m[58]&m[518]&m[714]))):InitCond[524];
    m[160] = run?((((~m[60]&~m[421]&~m[617])|(m[60]&m[421]&~m[617]))&BiasedRNG[316])|(((m[60]&~m[421]&~m[617])|(~m[60]&m[421]&m[617]))&~BiasedRNG[316])|((~m[60]&~m[421]&m[617])|(m[60]&~m[421]&m[617])|(m[60]&m[421]&m[617]))):InitCond[525];
    m[161] = run?((((~m[60]&~m[435]&~m[631])|(m[60]&m[435]&~m[631]))&BiasedRNG[317])|(((m[60]&~m[435]&~m[631])|(~m[60]&m[435]&m[631]))&~BiasedRNG[317])|((~m[60]&~m[435]&m[631])|(m[60]&~m[435]&m[631])|(m[60]&m[435]&m[631]))):InitCond[526];
    m[162] = run?((((~m[60]&~m[449]&~m[645])|(m[60]&m[449]&~m[645]))&BiasedRNG[318])|(((m[60]&~m[449]&~m[645])|(~m[60]&m[449]&m[645]))&~BiasedRNG[318])|((~m[60]&~m[449]&m[645])|(m[60]&~m[449]&m[645])|(m[60]&m[449]&m[645]))):InitCond[527];
    m[163] = run?((((~m[60]&~m[463]&~m[659])|(m[60]&m[463]&~m[659]))&BiasedRNG[319])|(((m[60]&~m[463]&~m[659])|(~m[60]&m[463]&m[659]))&~BiasedRNG[319])|((~m[60]&~m[463]&m[659])|(m[60]&~m[463]&m[659])|(m[60]&m[463]&m[659]))):InitCond[528];
    m[164] = run?((((~m[61]&~m[477]&~m[673])|(m[61]&m[477]&~m[673]))&BiasedRNG[320])|(((m[61]&~m[477]&~m[673])|(~m[61]&m[477]&m[673]))&~BiasedRNG[320])|((~m[61]&~m[477]&m[673])|(m[61]&~m[477]&m[673])|(m[61]&m[477]&m[673]))):InitCond[529];
    m[165] = run?((((~m[61]&~m[491]&~m[687])|(m[61]&m[491]&~m[687]))&BiasedRNG[321])|(((m[61]&~m[491]&~m[687])|(~m[61]&m[491]&m[687]))&~BiasedRNG[321])|((~m[61]&~m[491]&m[687])|(m[61]&~m[491]&m[687])|(m[61]&m[491]&m[687]))):InitCond[530];
    m[166] = run?((((~m[61]&~m[505]&~m[701])|(m[61]&m[505]&~m[701]))&BiasedRNG[322])|(((m[61]&~m[505]&~m[701])|(~m[61]&m[505]&m[701]))&~BiasedRNG[322])|((~m[61]&~m[505]&m[701])|(m[61]&~m[505]&m[701])|(m[61]&m[505]&m[701]))):InitCond[531];
    m[167] = run?((((~m[61]&~m[519]&~m[715])|(m[61]&m[519]&~m[715]))&BiasedRNG[323])|(((m[61]&~m[519]&~m[715])|(~m[61]&m[519]&m[715]))&~BiasedRNG[323])|((~m[61]&~m[519]&m[715])|(m[61]&~m[519]&m[715])|(m[61]&m[519]&m[715]))):InitCond[532];
    m[174] = run?((((~m[63]&~m[422]&~m[618])|(m[63]&m[422]&~m[618]))&BiasedRNG[324])|(((m[63]&~m[422]&~m[618])|(~m[63]&m[422]&m[618]))&~BiasedRNG[324])|((~m[63]&~m[422]&m[618])|(m[63]&~m[422]&m[618])|(m[63]&m[422]&m[618]))):InitCond[533];
    m[175] = run?((((~m[63]&~m[436]&~m[632])|(m[63]&m[436]&~m[632]))&BiasedRNG[325])|(((m[63]&~m[436]&~m[632])|(~m[63]&m[436]&m[632]))&~BiasedRNG[325])|((~m[63]&~m[436]&m[632])|(m[63]&~m[436]&m[632])|(m[63]&m[436]&m[632]))):InitCond[534];
    m[176] = run?((((~m[63]&~m[450]&~m[646])|(m[63]&m[450]&~m[646]))&BiasedRNG[326])|(((m[63]&~m[450]&~m[646])|(~m[63]&m[450]&m[646]))&~BiasedRNG[326])|((~m[63]&~m[450]&m[646])|(m[63]&~m[450]&m[646])|(m[63]&m[450]&m[646]))):InitCond[535];
    m[177] = run?((((~m[63]&~m[464]&~m[660])|(m[63]&m[464]&~m[660]))&BiasedRNG[327])|(((m[63]&~m[464]&~m[660])|(~m[63]&m[464]&m[660]))&~BiasedRNG[327])|((~m[63]&~m[464]&m[660])|(m[63]&~m[464]&m[660])|(m[63]&m[464]&m[660]))):InitCond[536];
    m[178] = run?((((~m[64]&~m[478]&~m[674])|(m[64]&m[478]&~m[674]))&BiasedRNG[328])|(((m[64]&~m[478]&~m[674])|(~m[64]&m[478]&m[674]))&~BiasedRNG[328])|((~m[64]&~m[478]&m[674])|(m[64]&~m[478]&m[674])|(m[64]&m[478]&m[674]))):InitCond[537];
    m[179] = run?((((~m[64]&~m[492]&~m[688])|(m[64]&m[492]&~m[688]))&BiasedRNG[329])|(((m[64]&~m[492]&~m[688])|(~m[64]&m[492]&m[688]))&~BiasedRNG[329])|((~m[64]&~m[492]&m[688])|(m[64]&~m[492]&m[688])|(m[64]&m[492]&m[688]))):InitCond[538];
    m[180] = run?((((~m[64]&~m[506]&~m[702])|(m[64]&m[506]&~m[702]))&BiasedRNG[330])|(((m[64]&~m[506]&~m[702])|(~m[64]&m[506]&m[702]))&~BiasedRNG[330])|((~m[64]&~m[506]&m[702])|(m[64]&~m[506]&m[702])|(m[64]&m[506]&m[702]))):InitCond[539];
    m[181] = run?((((~m[64]&~m[520]&~m[716])|(m[64]&m[520]&~m[716]))&BiasedRNG[331])|(((m[64]&~m[520]&~m[716])|(~m[64]&m[520]&m[716]))&~BiasedRNG[331])|((~m[64]&~m[520]&m[716])|(m[64]&~m[520]&m[716])|(m[64]&m[520]&m[716]))):InitCond[540];
    m[188] = run?((((~m[66]&~m[423]&~m[619])|(m[66]&m[423]&~m[619]))&BiasedRNG[332])|(((m[66]&~m[423]&~m[619])|(~m[66]&m[423]&m[619]))&~BiasedRNG[332])|((~m[66]&~m[423]&m[619])|(m[66]&~m[423]&m[619])|(m[66]&m[423]&m[619]))):InitCond[541];
    m[189] = run?((((~m[66]&~m[437]&~m[633])|(m[66]&m[437]&~m[633]))&BiasedRNG[333])|(((m[66]&~m[437]&~m[633])|(~m[66]&m[437]&m[633]))&~BiasedRNG[333])|((~m[66]&~m[437]&m[633])|(m[66]&~m[437]&m[633])|(m[66]&m[437]&m[633]))):InitCond[542];
    m[190] = run?((((~m[66]&~m[451]&~m[647])|(m[66]&m[451]&~m[647]))&BiasedRNG[334])|(((m[66]&~m[451]&~m[647])|(~m[66]&m[451]&m[647]))&~BiasedRNG[334])|((~m[66]&~m[451]&m[647])|(m[66]&~m[451]&m[647])|(m[66]&m[451]&m[647]))):InitCond[543];
    m[191] = run?((((~m[66]&~m[465]&~m[661])|(m[66]&m[465]&~m[661]))&BiasedRNG[335])|(((m[66]&~m[465]&~m[661])|(~m[66]&m[465]&m[661]))&~BiasedRNG[335])|((~m[66]&~m[465]&m[661])|(m[66]&~m[465]&m[661])|(m[66]&m[465]&m[661]))):InitCond[544];
    m[192] = run?((((~m[67]&~m[479]&~m[675])|(m[67]&m[479]&~m[675]))&BiasedRNG[336])|(((m[67]&~m[479]&~m[675])|(~m[67]&m[479]&m[675]))&~BiasedRNG[336])|((~m[67]&~m[479]&m[675])|(m[67]&~m[479]&m[675])|(m[67]&m[479]&m[675]))):InitCond[545];
    m[193] = run?((((~m[67]&~m[493]&~m[689])|(m[67]&m[493]&~m[689]))&BiasedRNG[337])|(((m[67]&~m[493]&~m[689])|(~m[67]&m[493]&m[689]))&~BiasedRNG[337])|((~m[67]&~m[493]&m[689])|(m[67]&~m[493]&m[689])|(m[67]&m[493]&m[689]))):InitCond[546];
    m[194] = run?((((~m[67]&~m[507]&~m[703])|(m[67]&m[507]&~m[703]))&BiasedRNG[338])|(((m[67]&~m[507]&~m[703])|(~m[67]&m[507]&m[703]))&~BiasedRNG[338])|((~m[67]&~m[507]&m[703])|(m[67]&~m[507]&m[703])|(m[67]&m[507]&m[703]))):InitCond[547];
    m[195] = run?((((~m[67]&~m[521]&~m[717])|(m[67]&m[521]&~m[717]))&BiasedRNG[339])|(((m[67]&~m[521]&~m[717])|(~m[67]&m[521]&m[717]))&~BiasedRNG[339])|((~m[67]&~m[521]&m[717])|(m[67]&~m[521]&m[717])|(m[67]&m[521]&m[717]))):InitCond[548];
    m[202] = run?((((~m[69]&~m[424]&~m[620])|(m[69]&m[424]&~m[620]))&BiasedRNG[340])|(((m[69]&~m[424]&~m[620])|(~m[69]&m[424]&m[620]))&~BiasedRNG[340])|((~m[69]&~m[424]&m[620])|(m[69]&~m[424]&m[620])|(m[69]&m[424]&m[620]))):InitCond[549];
    m[203] = run?((((~m[69]&~m[438]&~m[634])|(m[69]&m[438]&~m[634]))&BiasedRNG[341])|(((m[69]&~m[438]&~m[634])|(~m[69]&m[438]&m[634]))&~BiasedRNG[341])|((~m[69]&~m[438]&m[634])|(m[69]&~m[438]&m[634])|(m[69]&m[438]&m[634]))):InitCond[550];
    m[204] = run?((((~m[69]&~m[452]&~m[648])|(m[69]&m[452]&~m[648]))&BiasedRNG[342])|(((m[69]&~m[452]&~m[648])|(~m[69]&m[452]&m[648]))&~BiasedRNG[342])|((~m[69]&~m[452]&m[648])|(m[69]&~m[452]&m[648])|(m[69]&m[452]&m[648]))):InitCond[551];
    m[205] = run?((((~m[69]&~m[466]&~m[662])|(m[69]&m[466]&~m[662]))&BiasedRNG[343])|(((m[69]&~m[466]&~m[662])|(~m[69]&m[466]&m[662]))&~BiasedRNG[343])|((~m[69]&~m[466]&m[662])|(m[69]&~m[466]&m[662])|(m[69]&m[466]&m[662]))):InitCond[552];
    m[206] = run?((((~m[70]&~m[480]&~m[676])|(m[70]&m[480]&~m[676]))&BiasedRNG[344])|(((m[70]&~m[480]&~m[676])|(~m[70]&m[480]&m[676]))&~BiasedRNG[344])|((~m[70]&~m[480]&m[676])|(m[70]&~m[480]&m[676])|(m[70]&m[480]&m[676]))):InitCond[553];
    m[207] = run?((((~m[70]&~m[494]&~m[690])|(m[70]&m[494]&~m[690]))&BiasedRNG[345])|(((m[70]&~m[494]&~m[690])|(~m[70]&m[494]&m[690]))&~BiasedRNG[345])|((~m[70]&~m[494]&m[690])|(m[70]&~m[494]&m[690])|(m[70]&m[494]&m[690]))):InitCond[554];
    m[208] = run?((((~m[70]&~m[508]&~m[704])|(m[70]&m[508]&~m[704]))&BiasedRNG[346])|(((m[70]&~m[508]&~m[704])|(~m[70]&m[508]&m[704]))&~BiasedRNG[346])|((~m[70]&~m[508]&m[704])|(m[70]&~m[508]&m[704])|(m[70]&m[508]&m[704]))):InitCond[555];
    m[209] = run?((((~m[70]&~m[522]&~m[718])|(m[70]&m[522]&~m[718]))&BiasedRNG[347])|(((m[70]&~m[522]&~m[718])|(~m[70]&m[522]&m[718]))&~BiasedRNG[347])|((~m[70]&~m[522]&m[718])|(m[70]&~m[522]&m[718])|(m[70]&m[522]&m[718]))):InitCond[556];
    m[216] = run?((((~m[72]&~m[425]&~m[621])|(m[72]&m[425]&~m[621]))&BiasedRNG[348])|(((m[72]&~m[425]&~m[621])|(~m[72]&m[425]&m[621]))&~BiasedRNG[348])|((~m[72]&~m[425]&m[621])|(m[72]&~m[425]&m[621])|(m[72]&m[425]&m[621]))):InitCond[557];
    m[217] = run?((((~m[72]&~m[439]&~m[635])|(m[72]&m[439]&~m[635]))&BiasedRNG[349])|(((m[72]&~m[439]&~m[635])|(~m[72]&m[439]&m[635]))&~BiasedRNG[349])|((~m[72]&~m[439]&m[635])|(m[72]&~m[439]&m[635])|(m[72]&m[439]&m[635]))):InitCond[558];
    m[218] = run?((((~m[72]&~m[453]&~m[649])|(m[72]&m[453]&~m[649]))&BiasedRNG[350])|(((m[72]&~m[453]&~m[649])|(~m[72]&m[453]&m[649]))&~BiasedRNG[350])|((~m[72]&~m[453]&m[649])|(m[72]&~m[453]&m[649])|(m[72]&m[453]&m[649]))):InitCond[559];
    m[219] = run?((((~m[72]&~m[467]&~m[663])|(m[72]&m[467]&~m[663]))&BiasedRNG[351])|(((m[72]&~m[467]&~m[663])|(~m[72]&m[467]&m[663]))&~BiasedRNG[351])|((~m[72]&~m[467]&m[663])|(m[72]&~m[467]&m[663])|(m[72]&m[467]&m[663]))):InitCond[560];
    m[220] = run?((((~m[73]&~m[481]&~m[677])|(m[73]&m[481]&~m[677]))&BiasedRNG[352])|(((m[73]&~m[481]&~m[677])|(~m[73]&m[481]&m[677]))&~BiasedRNG[352])|((~m[73]&~m[481]&m[677])|(m[73]&~m[481]&m[677])|(m[73]&m[481]&m[677]))):InitCond[561];
    m[221] = run?((((~m[73]&~m[495]&~m[691])|(m[73]&m[495]&~m[691]))&BiasedRNG[353])|(((m[73]&~m[495]&~m[691])|(~m[73]&m[495]&m[691]))&~BiasedRNG[353])|((~m[73]&~m[495]&m[691])|(m[73]&~m[495]&m[691])|(m[73]&m[495]&m[691]))):InitCond[562];
    m[222] = run?((((~m[73]&~m[509]&~m[705])|(m[73]&m[509]&~m[705]))&BiasedRNG[354])|(((m[73]&~m[509]&~m[705])|(~m[73]&m[509]&m[705]))&~BiasedRNG[354])|((~m[73]&~m[509]&m[705])|(m[73]&~m[509]&m[705])|(m[73]&m[509]&m[705]))):InitCond[563];
    m[223] = run?((((~m[73]&~m[523]&~m[719])|(m[73]&m[523]&~m[719]))&BiasedRNG[355])|(((m[73]&~m[523]&~m[719])|(~m[73]&m[523]&m[719]))&~BiasedRNG[355])|((~m[73]&~m[523]&m[719])|(m[73]&~m[523]&m[719])|(m[73]&m[523]&m[719]))):InitCond[564];
    m[230] = run?((((~m[75]&~m[426]&~m[622])|(m[75]&m[426]&~m[622]))&BiasedRNG[356])|(((m[75]&~m[426]&~m[622])|(~m[75]&m[426]&m[622]))&~BiasedRNG[356])|((~m[75]&~m[426]&m[622])|(m[75]&~m[426]&m[622])|(m[75]&m[426]&m[622]))):InitCond[565];
    m[231] = run?((((~m[75]&~m[440]&~m[636])|(m[75]&m[440]&~m[636]))&BiasedRNG[357])|(((m[75]&~m[440]&~m[636])|(~m[75]&m[440]&m[636]))&~BiasedRNG[357])|((~m[75]&~m[440]&m[636])|(m[75]&~m[440]&m[636])|(m[75]&m[440]&m[636]))):InitCond[566];
    m[232] = run?((((~m[75]&~m[454]&~m[650])|(m[75]&m[454]&~m[650]))&BiasedRNG[358])|(((m[75]&~m[454]&~m[650])|(~m[75]&m[454]&m[650]))&~BiasedRNG[358])|((~m[75]&~m[454]&m[650])|(m[75]&~m[454]&m[650])|(m[75]&m[454]&m[650]))):InitCond[567];
    m[233] = run?((((~m[75]&~m[468]&~m[664])|(m[75]&m[468]&~m[664]))&BiasedRNG[359])|(((m[75]&~m[468]&~m[664])|(~m[75]&m[468]&m[664]))&~BiasedRNG[359])|((~m[75]&~m[468]&m[664])|(m[75]&~m[468]&m[664])|(m[75]&m[468]&m[664]))):InitCond[568];
    m[234] = run?((((~m[76]&~m[482]&~m[678])|(m[76]&m[482]&~m[678]))&BiasedRNG[360])|(((m[76]&~m[482]&~m[678])|(~m[76]&m[482]&m[678]))&~BiasedRNG[360])|((~m[76]&~m[482]&m[678])|(m[76]&~m[482]&m[678])|(m[76]&m[482]&m[678]))):InitCond[569];
    m[235] = run?((((~m[76]&~m[496]&~m[692])|(m[76]&m[496]&~m[692]))&BiasedRNG[361])|(((m[76]&~m[496]&~m[692])|(~m[76]&m[496]&m[692]))&~BiasedRNG[361])|((~m[76]&~m[496]&m[692])|(m[76]&~m[496]&m[692])|(m[76]&m[496]&m[692]))):InitCond[570];
    m[236] = run?((((~m[76]&~m[510]&~m[706])|(m[76]&m[510]&~m[706]))&BiasedRNG[362])|(((m[76]&~m[510]&~m[706])|(~m[76]&m[510]&m[706]))&~BiasedRNG[362])|((~m[76]&~m[510]&m[706])|(m[76]&~m[510]&m[706])|(m[76]&m[510]&m[706]))):InitCond[571];
    m[237] = run?((((~m[76]&~m[524]&~m[720])|(m[76]&m[524]&~m[720]))&BiasedRNG[363])|(((m[76]&~m[524]&~m[720])|(~m[76]&m[524]&m[720]))&~BiasedRNG[363])|((~m[76]&~m[524]&m[720])|(m[76]&~m[524]&m[720])|(m[76]&m[524]&m[720]))):InitCond[572];
    m[244] = run?((((~m[78]&~m[427]&~m[623])|(m[78]&m[427]&~m[623]))&BiasedRNG[364])|(((m[78]&~m[427]&~m[623])|(~m[78]&m[427]&m[623]))&~BiasedRNG[364])|((~m[78]&~m[427]&m[623])|(m[78]&~m[427]&m[623])|(m[78]&m[427]&m[623]))):InitCond[573];
    m[245] = run?((((~m[78]&~m[441]&~m[637])|(m[78]&m[441]&~m[637]))&BiasedRNG[365])|(((m[78]&~m[441]&~m[637])|(~m[78]&m[441]&m[637]))&~BiasedRNG[365])|((~m[78]&~m[441]&m[637])|(m[78]&~m[441]&m[637])|(m[78]&m[441]&m[637]))):InitCond[574];
    m[246] = run?((((~m[78]&~m[455]&~m[651])|(m[78]&m[455]&~m[651]))&BiasedRNG[366])|(((m[78]&~m[455]&~m[651])|(~m[78]&m[455]&m[651]))&~BiasedRNG[366])|((~m[78]&~m[455]&m[651])|(m[78]&~m[455]&m[651])|(m[78]&m[455]&m[651]))):InitCond[575];
    m[247] = run?((((~m[78]&~m[469]&~m[665])|(m[78]&m[469]&~m[665]))&BiasedRNG[367])|(((m[78]&~m[469]&~m[665])|(~m[78]&m[469]&m[665]))&~BiasedRNG[367])|((~m[78]&~m[469]&m[665])|(m[78]&~m[469]&m[665])|(m[78]&m[469]&m[665]))):InitCond[576];
    m[248] = run?((((~m[79]&~m[483]&~m[679])|(m[79]&m[483]&~m[679]))&BiasedRNG[368])|(((m[79]&~m[483]&~m[679])|(~m[79]&m[483]&m[679]))&~BiasedRNG[368])|((~m[79]&~m[483]&m[679])|(m[79]&~m[483]&m[679])|(m[79]&m[483]&m[679]))):InitCond[577];
    m[249] = run?((((~m[79]&~m[497]&~m[693])|(m[79]&m[497]&~m[693]))&BiasedRNG[369])|(((m[79]&~m[497]&~m[693])|(~m[79]&m[497]&m[693]))&~BiasedRNG[369])|((~m[79]&~m[497]&m[693])|(m[79]&~m[497]&m[693])|(m[79]&m[497]&m[693]))):InitCond[578];
    m[250] = run?((((~m[79]&~m[511]&~m[707])|(m[79]&m[511]&~m[707]))&BiasedRNG[370])|(((m[79]&~m[511]&~m[707])|(~m[79]&m[511]&m[707]))&~BiasedRNG[370])|((~m[79]&~m[511]&m[707])|(m[79]&~m[511]&m[707])|(m[79]&m[511]&m[707]))):InitCond[579];
    m[251] = run?((((~m[79]&~m[525]&~m[721])|(m[79]&m[525]&~m[721]))&BiasedRNG[371])|(((m[79]&~m[525]&~m[721])|(~m[79]&m[525]&m[721]))&~BiasedRNG[371])|((~m[79]&~m[525]&m[721])|(m[79]&~m[525]&m[721])|(m[79]&m[525]&m[721]))):InitCond[580];
    m[258] = run?((((~m[81]&~m[428]&~m[624])|(m[81]&m[428]&~m[624]))&BiasedRNG[372])|(((m[81]&~m[428]&~m[624])|(~m[81]&m[428]&m[624]))&~BiasedRNG[372])|((~m[81]&~m[428]&m[624])|(m[81]&~m[428]&m[624])|(m[81]&m[428]&m[624]))):InitCond[581];
    m[259] = run?((((~m[81]&~m[442]&~m[638])|(m[81]&m[442]&~m[638]))&BiasedRNG[373])|(((m[81]&~m[442]&~m[638])|(~m[81]&m[442]&m[638]))&~BiasedRNG[373])|((~m[81]&~m[442]&m[638])|(m[81]&~m[442]&m[638])|(m[81]&m[442]&m[638]))):InitCond[582];
    m[260] = run?((((~m[81]&~m[456]&~m[652])|(m[81]&m[456]&~m[652]))&BiasedRNG[374])|(((m[81]&~m[456]&~m[652])|(~m[81]&m[456]&m[652]))&~BiasedRNG[374])|((~m[81]&~m[456]&m[652])|(m[81]&~m[456]&m[652])|(m[81]&m[456]&m[652]))):InitCond[583];
    m[261] = run?((((~m[81]&~m[470]&~m[666])|(m[81]&m[470]&~m[666]))&BiasedRNG[375])|(((m[81]&~m[470]&~m[666])|(~m[81]&m[470]&m[666]))&~BiasedRNG[375])|((~m[81]&~m[470]&m[666])|(m[81]&~m[470]&m[666])|(m[81]&m[470]&m[666]))):InitCond[584];
    m[262] = run?((((~m[82]&~m[484]&~m[680])|(m[82]&m[484]&~m[680]))&BiasedRNG[376])|(((m[82]&~m[484]&~m[680])|(~m[82]&m[484]&m[680]))&~BiasedRNG[376])|((~m[82]&~m[484]&m[680])|(m[82]&~m[484]&m[680])|(m[82]&m[484]&m[680]))):InitCond[585];
    m[263] = run?((((~m[82]&~m[498]&~m[694])|(m[82]&m[498]&~m[694]))&BiasedRNG[377])|(((m[82]&~m[498]&~m[694])|(~m[82]&m[498]&m[694]))&~BiasedRNG[377])|((~m[82]&~m[498]&m[694])|(m[82]&~m[498]&m[694])|(m[82]&m[498]&m[694]))):InitCond[586];
    m[264] = run?((((~m[82]&~m[512]&~m[708])|(m[82]&m[512]&~m[708]))&BiasedRNG[378])|(((m[82]&~m[512]&~m[708])|(~m[82]&m[512]&m[708]))&~BiasedRNG[378])|((~m[82]&~m[512]&m[708])|(m[82]&~m[512]&m[708])|(m[82]&m[512]&m[708]))):InitCond[587];
    m[265] = run?((((~m[82]&~m[526]&~m[722])|(m[82]&m[526]&~m[722]))&BiasedRNG[379])|(((m[82]&~m[526]&~m[722])|(~m[82]&m[526]&m[722]))&~BiasedRNG[379])|((~m[82]&~m[526]&m[722])|(m[82]&~m[526]&m[722])|(m[82]&m[526]&m[722]))):InitCond[588];
    m[272] = run?((((~m[84]&~m[429]&~m[625])|(m[84]&m[429]&~m[625]))&BiasedRNG[380])|(((m[84]&~m[429]&~m[625])|(~m[84]&m[429]&m[625]))&~BiasedRNG[380])|((~m[84]&~m[429]&m[625])|(m[84]&~m[429]&m[625])|(m[84]&m[429]&m[625]))):InitCond[589];
    m[273] = run?((((~m[84]&~m[443]&~m[639])|(m[84]&m[443]&~m[639]))&BiasedRNG[381])|(((m[84]&~m[443]&~m[639])|(~m[84]&m[443]&m[639]))&~BiasedRNG[381])|((~m[84]&~m[443]&m[639])|(m[84]&~m[443]&m[639])|(m[84]&m[443]&m[639]))):InitCond[590];
    m[274] = run?((((~m[84]&~m[457]&~m[653])|(m[84]&m[457]&~m[653]))&BiasedRNG[382])|(((m[84]&~m[457]&~m[653])|(~m[84]&m[457]&m[653]))&~BiasedRNG[382])|((~m[84]&~m[457]&m[653])|(m[84]&~m[457]&m[653])|(m[84]&m[457]&m[653]))):InitCond[591];
    m[275] = run?((((~m[84]&~m[471]&~m[667])|(m[84]&m[471]&~m[667]))&BiasedRNG[383])|(((m[84]&~m[471]&~m[667])|(~m[84]&m[471]&m[667]))&~BiasedRNG[383])|((~m[84]&~m[471]&m[667])|(m[84]&~m[471]&m[667])|(m[84]&m[471]&m[667]))):InitCond[592];
    m[276] = run?((((~m[85]&~m[485]&~m[681])|(m[85]&m[485]&~m[681]))&BiasedRNG[384])|(((m[85]&~m[485]&~m[681])|(~m[85]&m[485]&m[681]))&~BiasedRNG[384])|((~m[85]&~m[485]&m[681])|(m[85]&~m[485]&m[681])|(m[85]&m[485]&m[681]))):InitCond[593];
    m[277] = run?((((~m[85]&~m[499]&~m[695])|(m[85]&m[499]&~m[695]))&BiasedRNG[385])|(((m[85]&~m[499]&~m[695])|(~m[85]&m[499]&m[695]))&~BiasedRNG[385])|((~m[85]&~m[499]&m[695])|(m[85]&~m[499]&m[695])|(m[85]&m[499]&m[695]))):InitCond[594];
    m[278] = run?((((~m[85]&~m[513]&~m[709])|(m[85]&m[513]&~m[709]))&BiasedRNG[386])|(((m[85]&~m[513]&~m[709])|(~m[85]&m[513]&m[709]))&~BiasedRNG[386])|((~m[85]&~m[513]&m[709])|(m[85]&~m[513]&m[709])|(m[85]&m[513]&m[709]))):InitCond[595];
    m[279] = run?((((~m[85]&~m[527]&~m[723])|(m[85]&m[527]&~m[723]))&BiasedRNG[387])|(((m[85]&~m[527]&~m[723])|(~m[85]&m[527]&m[723]))&~BiasedRNG[387])|((~m[85]&~m[527]&m[723])|(m[85]&~m[527]&m[723])|(m[85]&m[527]&m[723]))):InitCond[596];
    m[286] = run?((((~m[87]&~m[430]&~m[626])|(m[87]&m[430]&~m[626]))&BiasedRNG[388])|(((m[87]&~m[430]&~m[626])|(~m[87]&m[430]&m[626]))&~BiasedRNG[388])|((~m[87]&~m[430]&m[626])|(m[87]&~m[430]&m[626])|(m[87]&m[430]&m[626]))):InitCond[597];
    m[287] = run?((((~m[87]&~m[444]&~m[640])|(m[87]&m[444]&~m[640]))&BiasedRNG[389])|(((m[87]&~m[444]&~m[640])|(~m[87]&m[444]&m[640]))&~BiasedRNG[389])|((~m[87]&~m[444]&m[640])|(m[87]&~m[444]&m[640])|(m[87]&m[444]&m[640]))):InitCond[598];
    m[288] = run?((((~m[87]&~m[458]&~m[654])|(m[87]&m[458]&~m[654]))&BiasedRNG[390])|(((m[87]&~m[458]&~m[654])|(~m[87]&m[458]&m[654]))&~BiasedRNG[390])|((~m[87]&~m[458]&m[654])|(m[87]&~m[458]&m[654])|(m[87]&m[458]&m[654]))):InitCond[599];
    m[289] = run?((((~m[87]&~m[472]&~m[668])|(m[87]&m[472]&~m[668]))&BiasedRNG[391])|(((m[87]&~m[472]&~m[668])|(~m[87]&m[472]&m[668]))&~BiasedRNG[391])|((~m[87]&~m[472]&m[668])|(m[87]&~m[472]&m[668])|(m[87]&m[472]&m[668]))):InitCond[600];
    m[290] = run?((((~m[88]&~m[486]&~m[682])|(m[88]&m[486]&~m[682]))&BiasedRNG[392])|(((m[88]&~m[486]&~m[682])|(~m[88]&m[486]&m[682]))&~BiasedRNG[392])|((~m[88]&~m[486]&m[682])|(m[88]&~m[486]&m[682])|(m[88]&m[486]&m[682]))):InitCond[601];
    m[291] = run?((((~m[88]&~m[500]&~m[696])|(m[88]&m[500]&~m[696]))&BiasedRNG[393])|(((m[88]&~m[500]&~m[696])|(~m[88]&m[500]&m[696]))&~BiasedRNG[393])|((~m[88]&~m[500]&m[696])|(m[88]&~m[500]&m[696])|(m[88]&m[500]&m[696]))):InitCond[602];
    m[292] = run?((((~m[88]&~m[514]&~m[710])|(m[88]&m[514]&~m[710]))&BiasedRNG[394])|(((m[88]&~m[514]&~m[710])|(~m[88]&m[514]&m[710]))&~BiasedRNG[394])|((~m[88]&~m[514]&m[710])|(m[88]&~m[514]&m[710])|(m[88]&m[514]&m[710]))):InitCond[603];
    m[293] = run?((((~m[88]&~m[528]&~m[724])|(m[88]&m[528]&~m[724]))&BiasedRNG[395])|(((m[88]&~m[528]&~m[724])|(~m[88]&m[528]&m[724]))&~BiasedRNG[395])|((~m[88]&~m[528]&m[724])|(m[88]&~m[528]&m[724])|(m[88]&m[528]&m[724]))):InitCond[604];
    m[300] = run?((((~m[90]&~m[431]&~m[627])|(m[90]&m[431]&~m[627]))&BiasedRNG[396])|(((m[90]&~m[431]&~m[627])|(~m[90]&m[431]&m[627]))&~BiasedRNG[396])|((~m[90]&~m[431]&m[627])|(m[90]&~m[431]&m[627])|(m[90]&m[431]&m[627]))):InitCond[605];
    m[301] = run?((((~m[90]&~m[445]&~m[641])|(m[90]&m[445]&~m[641]))&BiasedRNG[397])|(((m[90]&~m[445]&~m[641])|(~m[90]&m[445]&m[641]))&~BiasedRNG[397])|((~m[90]&~m[445]&m[641])|(m[90]&~m[445]&m[641])|(m[90]&m[445]&m[641]))):InitCond[606];
    m[302] = run?((((~m[90]&~m[459]&~m[655])|(m[90]&m[459]&~m[655]))&BiasedRNG[398])|(((m[90]&~m[459]&~m[655])|(~m[90]&m[459]&m[655]))&~BiasedRNG[398])|((~m[90]&~m[459]&m[655])|(m[90]&~m[459]&m[655])|(m[90]&m[459]&m[655]))):InitCond[607];
    m[303] = run?((((~m[90]&~m[473]&~m[669])|(m[90]&m[473]&~m[669]))&BiasedRNG[399])|(((m[90]&~m[473]&~m[669])|(~m[90]&m[473]&m[669]))&~BiasedRNG[399])|((~m[90]&~m[473]&m[669])|(m[90]&~m[473]&m[669])|(m[90]&m[473]&m[669]))):InitCond[608];
    m[304] = run?((((~m[91]&~m[487]&~m[683])|(m[91]&m[487]&~m[683]))&BiasedRNG[400])|(((m[91]&~m[487]&~m[683])|(~m[91]&m[487]&m[683]))&~BiasedRNG[400])|((~m[91]&~m[487]&m[683])|(m[91]&~m[487]&m[683])|(m[91]&m[487]&m[683]))):InitCond[609];
    m[305] = run?((((~m[91]&~m[501]&~m[697])|(m[91]&m[501]&~m[697]))&BiasedRNG[401])|(((m[91]&~m[501]&~m[697])|(~m[91]&m[501]&m[697]))&~BiasedRNG[401])|((~m[91]&~m[501]&m[697])|(m[91]&~m[501]&m[697])|(m[91]&m[501]&m[697]))):InitCond[610];
    m[306] = run?((((~m[91]&~m[515]&~m[711])|(m[91]&m[515]&~m[711]))&BiasedRNG[402])|(((m[91]&~m[515]&~m[711])|(~m[91]&m[515]&m[711]))&~BiasedRNG[402])|((~m[91]&~m[515]&m[711])|(m[91]&~m[515]&m[711])|(m[91]&m[515]&m[711]))):InitCond[611];
    m[307] = run?((((~m[91]&~m[529]&~m[725])|(m[91]&m[529]&~m[725]))&BiasedRNG[403])|(((m[91]&~m[529]&~m[725])|(~m[91]&m[529]&m[725]))&~BiasedRNG[403])|((~m[91]&~m[529]&m[725])|(m[91]&~m[529]&m[725])|(m[91]&m[529]&m[725]))):InitCond[612];
    m[314] = run?((((~m[93]&~m[432]&~m[628])|(m[93]&m[432]&~m[628]))&BiasedRNG[404])|(((m[93]&~m[432]&~m[628])|(~m[93]&m[432]&m[628]))&~BiasedRNG[404])|((~m[93]&~m[432]&m[628])|(m[93]&~m[432]&m[628])|(m[93]&m[432]&m[628]))):InitCond[613];
    m[315] = run?((((~m[93]&~m[446]&~m[642])|(m[93]&m[446]&~m[642]))&BiasedRNG[405])|(((m[93]&~m[446]&~m[642])|(~m[93]&m[446]&m[642]))&~BiasedRNG[405])|((~m[93]&~m[446]&m[642])|(m[93]&~m[446]&m[642])|(m[93]&m[446]&m[642]))):InitCond[614];
    m[316] = run?((((~m[93]&~m[460]&~m[656])|(m[93]&m[460]&~m[656]))&BiasedRNG[406])|(((m[93]&~m[460]&~m[656])|(~m[93]&m[460]&m[656]))&~BiasedRNG[406])|((~m[93]&~m[460]&m[656])|(m[93]&~m[460]&m[656])|(m[93]&m[460]&m[656]))):InitCond[615];
    m[317] = run?((((~m[93]&~m[474]&~m[670])|(m[93]&m[474]&~m[670]))&BiasedRNG[407])|(((m[93]&~m[474]&~m[670])|(~m[93]&m[474]&m[670]))&~BiasedRNG[407])|((~m[93]&~m[474]&m[670])|(m[93]&~m[474]&m[670])|(m[93]&m[474]&m[670]))):InitCond[616];
    m[318] = run?((((~m[94]&~m[488]&~m[684])|(m[94]&m[488]&~m[684]))&BiasedRNG[408])|(((m[94]&~m[488]&~m[684])|(~m[94]&m[488]&m[684]))&~BiasedRNG[408])|((~m[94]&~m[488]&m[684])|(m[94]&~m[488]&m[684])|(m[94]&m[488]&m[684]))):InitCond[617];
    m[319] = run?((((~m[94]&~m[502]&~m[698])|(m[94]&m[502]&~m[698]))&BiasedRNG[409])|(((m[94]&~m[502]&~m[698])|(~m[94]&m[502]&m[698]))&~BiasedRNG[409])|((~m[94]&~m[502]&m[698])|(m[94]&~m[502]&m[698])|(m[94]&m[502]&m[698]))):InitCond[618];
    m[320] = run?((((~m[94]&~m[516]&~m[712])|(m[94]&m[516]&~m[712]))&BiasedRNG[410])|(((m[94]&~m[516]&~m[712])|(~m[94]&m[516]&m[712]))&~BiasedRNG[410])|((~m[94]&~m[516]&m[712])|(m[94]&~m[516]&m[712])|(m[94]&m[516]&m[712]))):InitCond[619];
    m[321] = run?((((~m[94]&~m[530]&~m[726])|(m[94]&m[530]&~m[726]))&BiasedRNG[411])|(((m[94]&~m[530]&~m[726])|(~m[94]&m[530]&m[726]))&~BiasedRNG[411])|((~m[94]&~m[530]&m[726])|(m[94]&~m[530]&m[726])|(m[94]&m[530]&m[726]))):InitCond[620];
    m[328] = run?((((~m[96]&~m[433]&~m[629])|(m[96]&m[433]&~m[629]))&BiasedRNG[412])|(((m[96]&~m[433]&~m[629])|(~m[96]&m[433]&m[629]))&~BiasedRNG[412])|((~m[96]&~m[433]&m[629])|(m[96]&~m[433]&m[629])|(m[96]&m[433]&m[629]))):InitCond[621];
    m[329] = run?((((~m[96]&~m[447]&~m[643])|(m[96]&m[447]&~m[643]))&BiasedRNG[413])|(((m[96]&~m[447]&~m[643])|(~m[96]&m[447]&m[643]))&~BiasedRNG[413])|((~m[96]&~m[447]&m[643])|(m[96]&~m[447]&m[643])|(m[96]&m[447]&m[643]))):InitCond[622];
    m[330] = run?((((~m[96]&~m[461]&~m[657])|(m[96]&m[461]&~m[657]))&BiasedRNG[414])|(((m[96]&~m[461]&~m[657])|(~m[96]&m[461]&m[657]))&~BiasedRNG[414])|((~m[96]&~m[461]&m[657])|(m[96]&~m[461]&m[657])|(m[96]&m[461]&m[657]))):InitCond[623];
    m[331] = run?((((~m[96]&~m[475]&~m[671])|(m[96]&m[475]&~m[671]))&BiasedRNG[415])|(((m[96]&~m[475]&~m[671])|(~m[96]&m[475]&m[671]))&~BiasedRNG[415])|((~m[96]&~m[475]&m[671])|(m[96]&~m[475]&m[671])|(m[96]&m[475]&m[671]))):InitCond[624];
    m[332] = run?((((~m[97]&~m[489]&~m[685])|(m[97]&m[489]&~m[685]))&BiasedRNG[416])|(((m[97]&~m[489]&~m[685])|(~m[97]&m[489]&m[685]))&~BiasedRNG[416])|((~m[97]&~m[489]&m[685])|(m[97]&~m[489]&m[685])|(m[97]&m[489]&m[685]))):InitCond[625];
    m[333] = run?((((~m[97]&~m[503]&~m[699])|(m[97]&m[503]&~m[699]))&BiasedRNG[417])|(((m[97]&~m[503]&~m[699])|(~m[97]&m[503]&m[699]))&~BiasedRNG[417])|((~m[97]&~m[503]&m[699])|(m[97]&~m[503]&m[699])|(m[97]&m[503]&m[699]))):InitCond[626];
    m[334] = run?((((~m[97]&~m[517]&~m[713])|(m[97]&m[517]&~m[713]))&BiasedRNG[418])|(((m[97]&~m[517]&~m[713])|(~m[97]&m[517]&m[713]))&~BiasedRNG[418])|((~m[97]&~m[517]&m[713])|(m[97]&~m[517]&m[713])|(m[97]&m[517]&m[713]))):InitCond[627];
    m[335] = run?((((~m[97]&~m[531]&~m[727])|(m[97]&m[531]&~m[727]))&BiasedRNG[419])|(((m[97]&~m[531]&~m[727])|(~m[97]&m[531]&m[727]))&~BiasedRNG[419])|((~m[97]&~m[531]&m[727])|(m[97]&~m[531]&m[727])|(m[97]&m[531]&m[727]))):InitCond[628];
    m[342] = run?((((~m[99]&~m[224]&~m[538])|(m[99]&m[224]&~m[538]))&BiasedRNG[420])|(((m[99]&~m[224]&~m[538])|(~m[99]&m[224]&m[538]))&~BiasedRNG[420])|((~m[99]&~m[224]&m[538])|(m[99]&~m[224]&m[538])|(m[99]&m[224]&m[538]))):InitCond[629];
    m[343] = run?((((~m[99]&~m[238]&~m[539])|(m[99]&m[238]&~m[539]))&BiasedRNG[421])|(((m[99]&~m[238]&~m[539])|(~m[99]&m[238]&m[539]))&~BiasedRNG[421])|((~m[99]&~m[238]&m[539])|(m[99]&~m[238]&m[539])|(m[99]&m[238]&m[539]))):InitCond[630];
    m[344] = run?((((~m[99]&~m[252]&~m[540])|(m[99]&m[252]&~m[540]))&BiasedRNG[422])|(((m[99]&~m[252]&~m[540])|(~m[99]&m[252]&m[540]))&~BiasedRNG[422])|((~m[99]&~m[252]&m[540])|(m[99]&~m[252]&m[540])|(m[99]&m[252]&m[540]))):InitCond[631];
    m[345] = run?((((~m[99]&~m[266]&~m[541])|(m[99]&m[266]&~m[541]))&BiasedRNG[423])|(((m[99]&~m[266]&~m[541])|(~m[99]&m[266]&m[541]))&~BiasedRNG[423])|((~m[99]&~m[266]&m[541])|(m[99]&~m[266]&m[541])|(m[99]&m[266]&m[541]))):InitCond[632];
    m[346] = run?((((~m[100]&~m[280]&~m[542])|(m[100]&m[280]&~m[542]))&BiasedRNG[424])|(((m[100]&~m[280]&~m[542])|(~m[100]&m[280]&m[542]))&~BiasedRNG[424])|((~m[100]&~m[280]&m[542])|(m[100]&~m[280]&m[542])|(m[100]&m[280]&m[542]))):InitCond[633];
    m[347] = run?((((~m[100]&~m[294]&~m[543])|(m[100]&m[294]&~m[543]))&BiasedRNG[425])|(((m[100]&~m[294]&~m[543])|(~m[100]&m[294]&m[543]))&~BiasedRNG[425])|((~m[100]&~m[294]&m[543])|(m[100]&~m[294]&m[543])|(m[100]&m[294]&m[543]))):InitCond[634];
    m[348] = run?((((~m[100]&~m[308]&~m[544])|(m[100]&m[308]&~m[544]))&BiasedRNG[426])|(((m[100]&~m[308]&~m[544])|(~m[100]&m[308]&m[544]))&~BiasedRNG[426])|((~m[100]&~m[308]&m[544])|(m[100]&~m[308]&m[544])|(m[100]&m[308]&m[544]))):InitCond[635];
    m[349] = run?((((~m[100]&~m[322]&~m[545])|(m[100]&m[322]&~m[545]))&BiasedRNG[427])|(((m[100]&~m[322]&~m[545])|(~m[100]&m[322]&m[545]))&~BiasedRNG[427])|((~m[100]&~m[322]&m[545])|(m[100]&~m[322]&m[545])|(m[100]&m[322]&m[545]))):InitCond[636];
    m[356] = run?((((~m[102]&~m[225]&~m[552])|(m[102]&m[225]&~m[552]))&BiasedRNG[428])|(((m[102]&~m[225]&~m[552])|(~m[102]&m[225]&m[552]))&~BiasedRNG[428])|((~m[102]&~m[225]&m[552])|(m[102]&~m[225]&m[552])|(m[102]&m[225]&m[552]))):InitCond[637];
    m[357] = run?((((~m[102]&~m[239]&~m[553])|(m[102]&m[239]&~m[553]))&BiasedRNG[429])|(((m[102]&~m[239]&~m[553])|(~m[102]&m[239]&m[553]))&~BiasedRNG[429])|((~m[102]&~m[239]&m[553])|(m[102]&~m[239]&m[553])|(m[102]&m[239]&m[553]))):InitCond[638];
    m[358] = run?((((~m[102]&~m[253]&~m[554])|(m[102]&m[253]&~m[554]))&BiasedRNG[430])|(((m[102]&~m[253]&~m[554])|(~m[102]&m[253]&m[554]))&~BiasedRNG[430])|((~m[102]&~m[253]&m[554])|(m[102]&~m[253]&m[554])|(m[102]&m[253]&m[554]))):InitCond[639];
    m[359] = run?((((~m[102]&~m[267]&~m[555])|(m[102]&m[267]&~m[555]))&BiasedRNG[431])|(((m[102]&~m[267]&~m[555])|(~m[102]&m[267]&m[555]))&~BiasedRNG[431])|((~m[102]&~m[267]&m[555])|(m[102]&~m[267]&m[555])|(m[102]&m[267]&m[555]))):InitCond[640];
    m[360] = run?((((~m[103]&~m[281]&~m[556])|(m[103]&m[281]&~m[556]))&BiasedRNG[432])|(((m[103]&~m[281]&~m[556])|(~m[103]&m[281]&m[556]))&~BiasedRNG[432])|((~m[103]&~m[281]&m[556])|(m[103]&~m[281]&m[556])|(m[103]&m[281]&m[556]))):InitCond[641];
    m[361] = run?((((~m[103]&~m[295]&~m[557])|(m[103]&m[295]&~m[557]))&BiasedRNG[433])|(((m[103]&~m[295]&~m[557])|(~m[103]&m[295]&m[557]))&~BiasedRNG[433])|((~m[103]&~m[295]&m[557])|(m[103]&~m[295]&m[557])|(m[103]&m[295]&m[557]))):InitCond[642];
    m[362] = run?((((~m[103]&~m[309]&~m[558])|(m[103]&m[309]&~m[558]))&BiasedRNG[434])|(((m[103]&~m[309]&~m[558])|(~m[103]&m[309]&m[558]))&~BiasedRNG[434])|((~m[103]&~m[309]&m[558])|(m[103]&~m[309]&m[558])|(m[103]&m[309]&m[558]))):InitCond[643];
    m[363] = run?((((~m[103]&~m[323]&~m[559])|(m[103]&m[323]&~m[559]))&BiasedRNG[435])|(((m[103]&~m[323]&~m[559])|(~m[103]&m[323]&m[559]))&~BiasedRNG[435])|((~m[103]&~m[323]&m[559])|(m[103]&~m[323]&m[559])|(m[103]&m[323]&m[559]))):InitCond[644];
    m[370] = run?((((~m[105]&~m[226]&~m[566])|(m[105]&m[226]&~m[566]))&BiasedRNG[436])|(((m[105]&~m[226]&~m[566])|(~m[105]&m[226]&m[566]))&~BiasedRNG[436])|((~m[105]&~m[226]&m[566])|(m[105]&~m[226]&m[566])|(m[105]&m[226]&m[566]))):InitCond[645];
    m[371] = run?((((~m[105]&~m[240]&~m[567])|(m[105]&m[240]&~m[567]))&BiasedRNG[437])|(((m[105]&~m[240]&~m[567])|(~m[105]&m[240]&m[567]))&~BiasedRNG[437])|((~m[105]&~m[240]&m[567])|(m[105]&~m[240]&m[567])|(m[105]&m[240]&m[567]))):InitCond[646];
    m[372] = run?((((~m[105]&~m[254]&~m[568])|(m[105]&m[254]&~m[568]))&BiasedRNG[438])|(((m[105]&~m[254]&~m[568])|(~m[105]&m[254]&m[568]))&~BiasedRNG[438])|((~m[105]&~m[254]&m[568])|(m[105]&~m[254]&m[568])|(m[105]&m[254]&m[568]))):InitCond[647];
    m[373] = run?((((~m[105]&~m[268]&~m[569])|(m[105]&m[268]&~m[569]))&BiasedRNG[439])|(((m[105]&~m[268]&~m[569])|(~m[105]&m[268]&m[569]))&~BiasedRNG[439])|((~m[105]&~m[268]&m[569])|(m[105]&~m[268]&m[569])|(m[105]&m[268]&m[569]))):InitCond[648];
    m[374] = run?((((~m[106]&~m[282]&~m[570])|(m[106]&m[282]&~m[570]))&BiasedRNG[440])|(((m[106]&~m[282]&~m[570])|(~m[106]&m[282]&m[570]))&~BiasedRNG[440])|((~m[106]&~m[282]&m[570])|(m[106]&~m[282]&m[570])|(m[106]&m[282]&m[570]))):InitCond[649];
    m[375] = run?((((~m[106]&~m[296]&~m[571])|(m[106]&m[296]&~m[571]))&BiasedRNG[441])|(((m[106]&~m[296]&~m[571])|(~m[106]&m[296]&m[571]))&~BiasedRNG[441])|((~m[106]&~m[296]&m[571])|(m[106]&~m[296]&m[571])|(m[106]&m[296]&m[571]))):InitCond[650];
    m[376] = run?((((~m[106]&~m[310]&~m[572])|(m[106]&m[310]&~m[572]))&BiasedRNG[442])|(((m[106]&~m[310]&~m[572])|(~m[106]&m[310]&m[572]))&~BiasedRNG[442])|((~m[106]&~m[310]&m[572])|(m[106]&~m[310]&m[572])|(m[106]&m[310]&m[572]))):InitCond[651];
    m[377] = run?((((~m[106]&~m[324]&~m[573])|(m[106]&m[324]&~m[573]))&BiasedRNG[443])|(((m[106]&~m[324]&~m[573])|(~m[106]&m[324]&m[573]))&~BiasedRNG[443])|((~m[106]&~m[324]&m[573])|(m[106]&~m[324]&m[573])|(m[106]&m[324]&m[573]))):InitCond[652];
    m[384] = run?((((~m[108]&~m[227]&~m[580])|(m[108]&m[227]&~m[580]))&BiasedRNG[444])|(((m[108]&~m[227]&~m[580])|(~m[108]&m[227]&m[580]))&~BiasedRNG[444])|((~m[108]&~m[227]&m[580])|(m[108]&~m[227]&m[580])|(m[108]&m[227]&m[580]))):InitCond[653];
    m[385] = run?((((~m[108]&~m[241]&~m[581])|(m[108]&m[241]&~m[581]))&BiasedRNG[445])|(((m[108]&~m[241]&~m[581])|(~m[108]&m[241]&m[581]))&~BiasedRNG[445])|((~m[108]&~m[241]&m[581])|(m[108]&~m[241]&m[581])|(m[108]&m[241]&m[581]))):InitCond[654];
    m[386] = run?((((~m[108]&~m[255]&~m[582])|(m[108]&m[255]&~m[582]))&BiasedRNG[446])|(((m[108]&~m[255]&~m[582])|(~m[108]&m[255]&m[582]))&~BiasedRNG[446])|((~m[108]&~m[255]&m[582])|(m[108]&~m[255]&m[582])|(m[108]&m[255]&m[582]))):InitCond[655];
    m[387] = run?((((~m[108]&~m[269]&~m[583])|(m[108]&m[269]&~m[583]))&BiasedRNG[447])|(((m[108]&~m[269]&~m[583])|(~m[108]&m[269]&m[583]))&~BiasedRNG[447])|((~m[108]&~m[269]&m[583])|(m[108]&~m[269]&m[583])|(m[108]&m[269]&m[583]))):InitCond[656];
    m[388] = run?((((~m[109]&~m[283]&~m[584])|(m[109]&m[283]&~m[584]))&BiasedRNG[448])|(((m[109]&~m[283]&~m[584])|(~m[109]&m[283]&m[584]))&~BiasedRNG[448])|((~m[109]&~m[283]&m[584])|(m[109]&~m[283]&m[584])|(m[109]&m[283]&m[584]))):InitCond[657];
    m[389] = run?((((~m[109]&~m[297]&~m[585])|(m[109]&m[297]&~m[585]))&BiasedRNG[449])|(((m[109]&~m[297]&~m[585])|(~m[109]&m[297]&m[585]))&~BiasedRNG[449])|((~m[109]&~m[297]&m[585])|(m[109]&~m[297]&m[585])|(m[109]&m[297]&m[585]))):InitCond[658];
    m[390] = run?((((~m[109]&~m[311]&~m[586])|(m[109]&m[311]&~m[586]))&BiasedRNG[450])|(((m[109]&~m[311]&~m[586])|(~m[109]&m[311]&m[586]))&~BiasedRNG[450])|((~m[109]&~m[311]&m[586])|(m[109]&~m[311]&m[586])|(m[109]&m[311]&m[586]))):InitCond[659];
    m[391] = run?((((~m[109]&~m[325]&~m[587])|(m[109]&m[325]&~m[587]))&BiasedRNG[451])|(((m[109]&~m[325]&~m[587])|(~m[109]&m[325]&m[587]))&~BiasedRNG[451])|((~m[109]&~m[325]&m[587])|(m[109]&~m[325]&m[587])|(m[109]&m[325]&m[587]))):InitCond[660];
    m[398] = run?((((~m[111]&~m[228]&~m[594])|(m[111]&m[228]&~m[594]))&BiasedRNG[452])|(((m[111]&~m[228]&~m[594])|(~m[111]&m[228]&m[594]))&~BiasedRNG[452])|((~m[111]&~m[228]&m[594])|(m[111]&~m[228]&m[594])|(m[111]&m[228]&m[594]))):InitCond[661];
    m[399] = run?((((~m[111]&~m[242]&~m[595])|(m[111]&m[242]&~m[595]))&BiasedRNG[453])|(((m[111]&~m[242]&~m[595])|(~m[111]&m[242]&m[595]))&~BiasedRNG[453])|((~m[111]&~m[242]&m[595])|(m[111]&~m[242]&m[595])|(m[111]&m[242]&m[595]))):InitCond[662];
    m[400] = run?((((~m[111]&~m[256]&~m[596])|(m[111]&m[256]&~m[596]))&BiasedRNG[454])|(((m[111]&~m[256]&~m[596])|(~m[111]&m[256]&m[596]))&~BiasedRNG[454])|((~m[111]&~m[256]&m[596])|(m[111]&~m[256]&m[596])|(m[111]&m[256]&m[596]))):InitCond[663];
    m[401] = run?((((~m[111]&~m[270]&~m[597])|(m[111]&m[270]&~m[597]))&BiasedRNG[455])|(((m[111]&~m[270]&~m[597])|(~m[111]&m[270]&m[597]))&~BiasedRNG[455])|((~m[111]&~m[270]&m[597])|(m[111]&~m[270]&m[597])|(m[111]&m[270]&m[597]))):InitCond[664];
    m[402] = run?((((~m[112]&~m[284]&~m[598])|(m[112]&m[284]&~m[598]))&BiasedRNG[456])|(((m[112]&~m[284]&~m[598])|(~m[112]&m[284]&m[598]))&~BiasedRNG[456])|((~m[112]&~m[284]&m[598])|(m[112]&~m[284]&m[598])|(m[112]&m[284]&m[598]))):InitCond[665];
    m[403] = run?((((~m[112]&~m[298]&~m[599])|(m[112]&m[298]&~m[599]))&BiasedRNG[457])|(((m[112]&~m[298]&~m[599])|(~m[112]&m[298]&m[599]))&~BiasedRNG[457])|((~m[112]&~m[298]&m[599])|(m[112]&~m[298]&m[599])|(m[112]&m[298]&m[599]))):InitCond[666];
    m[404] = run?((((~m[112]&~m[312]&~m[600])|(m[112]&m[312]&~m[600]))&BiasedRNG[458])|(((m[112]&~m[312]&~m[600])|(~m[112]&m[312]&m[600]))&~BiasedRNG[458])|((~m[112]&~m[312]&m[600])|(m[112]&~m[312]&m[600])|(m[112]&m[312]&m[600]))):InitCond[667];
    m[405] = run?((((~m[112]&~m[326]&~m[601])|(m[112]&m[326]&~m[601]))&BiasedRNG[459])|(((m[112]&~m[326]&~m[601])|(~m[112]&m[326]&m[601]))&~BiasedRNG[459])|((~m[112]&~m[326]&m[601])|(m[112]&~m[326]&m[601])|(m[112]&m[326]&m[601]))):InitCond[668];
    m[412] = run?((((~m[114]&~m[229]&~m[608])|(m[114]&m[229]&~m[608]))&BiasedRNG[460])|(((m[114]&~m[229]&~m[608])|(~m[114]&m[229]&m[608]))&~BiasedRNG[460])|((~m[114]&~m[229]&m[608])|(m[114]&~m[229]&m[608])|(m[114]&m[229]&m[608]))):InitCond[669];
    m[413] = run?((((~m[114]&~m[243]&~m[609])|(m[114]&m[243]&~m[609]))&BiasedRNG[461])|(((m[114]&~m[243]&~m[609])|(~m[114]&m[243]&m[609]))&~BiasedRNG[461])|((~m[114]&~m[243]&m[609])|(m[114]&~m[243]&m[609])|(m[114]&m[243]&m[609]))):InitCond[670];
    m[414] = run?((((~m[114]&~m[257]&~m[610])|(m[114]&m[257]&~m[610]))&BiasedRNG[462])|(((m[114]&~m[257]&~m[610])|(~m[114]&m[257]&m[610]))&~BiasedRNG[462])|((~m[114]&~m[257]&m[610])|(m[114]&~m[257]&m[610])|(m[114]&m[257]&m[610]))):InitCond[671];
    m[415] = run?((((~m[114]&~m[271]&~m[611])|(m[114]&m[271]&~m[611]))&BiasedRNG[463])|(((m[114]&~m[271]&~m[611])|(~m[114]&m[271]&m[611]))&~BiasedRNG[463])|((~m[114]&~m[271]&m[611])|(m[114]&~m[271]&m[611])|(m[114]&m[271]&m[611]))):InitCond[672];
    m[416] = run?((((~m[115]&~m[285]&~m[612])|(m[115]&m[285]&~m[612]))&BiasedRNG[464])|(((m[115]&~m[285]&~m[612])|(~m[115]&m[285]&m[612]))&~BiasedRNG[464])|((~m[115]&~m[285]&m[612])|(m[115]&~m[285]&m[612])|(m[115]&m[285]&m[612]))):InitCond[673];
    m[417] = run?((((~m[115]&~m[299]&~m[613])|(m[115]&m[299]&~m[613]))&BiasedRNG[465])|(((m[115]&~m[299]&~m[613])|(~m[115]&m[299]&m[613]))&~BiasedRNG[465])|((~m[115]&~m[299]&m[613])|(m[115]&~m[299]&m[613])|(m[115]&m[299]&m[613]))):InitCond[674];
    m[418] = run?((((~m[115]&~m[313]&~m[614])|(m[115]&m[313]&~m[614]))&BiasedRNG[466])|(((m[115]&~m[313]&~m[614])|(~m[115]&m[313]&m[614]))&~BiasedRNG[466])|((~m[115]&~m[313]&m[614])|(m[115]&~m[313]&m[614])|(m[115]&m[313]&m[614]))):InitCond[675];
    m[419] = run?((((~m[115]&~m[327]&~m[615])|(m[115]&m[327]&~m[615]))&BiasedRNG[467])|(((m[115]&~m[327]&~m[615])|(~m[115]&m[327]&m[615]))&~BiasedRNG[467])|((~m[115]&~m[327]&m[615])|(m[115]&~m[327]&m[615])|(m[115]&m[327]&m[615]))):InitCond[676];
    m[533] = run?((((m[154]&~m[337]&m[728])|(~m[154]&m[337]&m[728]))&BiasedRNG[468])|(((m[154]&m[337]&~m[728]))&~BiasedRNG[468])|((m[154]&m[337]&m[728]))):InitCond[677];
    m[534] = run?((((m[168]&~m[338]&m[733])|(~m[168]&m[338]&m[733]))&BiasedRNG[469])|(((m[168]&m[338]&~m[733]))&~BiasedRNG[469])|((m[168]&m[338]&m[733]))):InitCond[678];
    m[535] = run?((((m[182]&~m[339]&m[743])|(~m[182]&m[339]&m[743]))&BiasedRNG[470])|(((m[182]&m[339]&~m[743]))&~BiasedRNG[470])|((m[182]&m[339]&m[743]))):InitCond[679];
    m[536] = run?((((m[196]&~m[340]&m[758])|(~m[196]&m[340]&m[758]))&BiasedRNG[471])|(((m[196]&m[340]&~m[758]))&~BiasedRNG[471])|((m[196]&m[340]&m[758]))):InitCond[680];
    m[537] = run?((((m[210]&~m[341]&m[778])|(~m[210]&m[341]&m[778]))&BiasedRNG[472])|(((m[210]&m[341]&~m[778]))&~BiasedRNG[472])|((m[210]&m[341]&m[778]))):InitCond[681];
    m[546] = run?((((m[141]&~m[350]&m[729])|(~m[141]&m[350]&m[729]))&BiasedRNG[473])|(((m[141]&m[350]&~m[729]))&~BiasedRNG[473])|((m[141]&m[350]&m[729]))):InitCond[682];
    m[547] = run?((((m[155]&~m[351]&m[734])|(~m[155]&m[351]&m[734]))&BiasedRNG[474])|(((m[155]&m[351]&~m[734]))&~BiasedRNG[474])|((m[155]&m[351]&m[734]))):InitCond[683];
    m[548] = run?((((m[169]&~m[352]&m[744])|(~m[169]&m[352]&m[744]))&BiasedRNG[475])|(((m[169]&m[352]&~m[744]))&~BiasedRNG[475])|((m[169]&m[352]&m[744]))):InitCond[684];
    m[549] = run?((((m[183]&~m[353]&m[759])|(~m[183]&m[353]&m[759]))&BiasedRNG[476])|(((m[183]&m[353]&~m[759]))&~BiasedRNG[476])|((m[183]&m[353]&m[759]))):InitCond[685];
    m[550] = run?((((m[197]&~m[354]&m[779])|(~m[197]&m[354]&m[779]))&BiasedRNG[477])|(((m[197]&m[354]&~m[779]))&~BiasedRNG[477])|((m[197]&m[354]&m[779]))):InitCond[686];
    m[551] = run?((((m[211]&~m[355]&m[804])|(~m[211]&m[355]&m[804]))&BiasedRNG[478])|(((m[211]&m[355]&~m[804]))&~BiasedRNG[478])|((m[211]&m[355]&m[804]))):InitCond[687];
    m[560] = run?((((m[142]&~m[364]&m[739])|(~m[142]&m[364]&m[739]))&BiasedRNG[479])|(((m[142]&m[364]&~m[739]))&~BiasedRNG[479])|((m[142]&m[364]&m[739]))):InitCond[688];
    m[561] = run?((((m[156]&~m[365]&m[749])|(~m[156]&m[365]&m[749]))&BiasedRNG[480])|(((m[156]&m[365]&~m[749]))&~BiasedRNG[480])|((m[156]&m[365]&m[749]))):InitCond[689];
    m[562] = run?((((m[170]&~m[366]&m[764])|(~m[170]&m[366]&m[764]))&BiasedRNG[481])|(((m[170]&m[366]&~m[764]))&~BiasedRNG[481])|((m[170]&m[366]&m[764]))):InitCond[690];
    m[563] = run?((((m[184]&~m[367]&m[784])|(~m[184]&m[367]&m[784]))&BiasedRNG[482])|(((m[184]&m[367]&~m[784]))&~BiasedRNG[482])|((m[184]&m[367]&m[784]))):InitCond[691];
    m[564] = run?((((m[198]&~m[368]&m[809])|(~m[198]&m[368]&m[809]))&BiasedRNG[483])|(((m[198]&m[368]&~m[809]))&~BiasedRNG[483])|((m[198]&m[368]&m[809]))):InitCond[692];
    m[565] = run?((((m[212]&~m[369]&m[839])|(~m[212]&m[369]&m[839]))&BiasedRNG[484])|(((m[212]&m[369]&~m[839]))&~BiasedRNG[484])|((m[212]&m[369]&m[839]))):InitCond[693];
    m[574] = run?((((m[143]&~m[378]&m[754])|(~m[143]&m[378]&m[754]))&BiasedRNG[485])|(((m[143]&m[378]&~m[754]))&~BiasedRNG[485])|((m[143]&m[378]&m[754]))):InitCond[694];
    m[575] = run?((((m[157]&~m[379]&m[769])|(~m[157]&m[379]&m[769]))&BiasedRNG[486])|(((m[157]&m[379]&~m[769]))&~BiasedRNG[486])|((m[157]&m[379]&m[769]))):InitCond[695];
    m[576] = run?((((m[171]&~m[380]&m[789])|(~m[171]&m[380]&m[789]))&BiasedRNG[487])|(((m[171]&m[380]&~m[789]))&~BiasedRNG[487])|((m[171]&m[380]&m[789]))):InitCond[696];
    m[577] = run?((((m[185]&~m[381]&m[814])|(~m[185]&m[381]&m[814]))&BiasedRNG[488])|(((m[185]&m[381]&~m[814]))&~BiasedRNG[488])|((m[185]&m[381]&m[814]))):InitCond[697];
    m[578] = run?((((m[199]&~m[382]&m[844])|(~m[199]&m[382]&m[844]))&BiasedRNG[489])|(((m[199]&m[382]&~m[844]))&~BiasedRNG[489])|((m[199]&m[382]&m[844]))):InitCond[698];
    m[579] = run?((((m[213]&~m[383]&m[879])|(~m[213]&m[383]&m[879]))&BiasedRNG[490])|(((m[213]&m[383]&~m[879]))&~BiasedRNG[490])|((m[213]&m[383]&m[879]))):InitCond[699];
    m[588] = run?((((m[144]&~m[392]&m[774])|(~m[144]&m[392]&m[774]))&BiasedRNG[491])|(((m[144]&m[392]&~m[774]))&~BiasedRNG[491])|((m[144]&m[392]&m[774]))):InitCond[700];
    m[589] = run?((((m[158]&~m[393]&m[794])|(~m[158]&m[393]&m[794]))&BiasedRNG[492])|(((m[158]&m[393]&~m[794]))&~BiasedRNG[492])|((m[158]&m[393]&m[794]))):InitCond[701];
    m[590] = run?((((m[172]&~m[394]&m[819])|(~m[172]&m[394]&m[819]))&BiasedRNG[493])|(((m[172]&m[394]&~m[819]))&~BiasedRNG[493])|((m[172]&m[394]&m[819]))):InitCond[702];
    m[591] = run?((((m[186]&~m[395]&m[849])|(~m[186]&m[395]&m[849]))&BiasedRNG[494])|(((m[186]&m[395]&~m[849]))&~BiasedRNG[494])|((m[186]&m[395]&m[849]))):InitCond[703];
    m[592] = run?((((m[200]&~m[396]&m[884])|(~m[200]&m[396]&m[884]))&BiasedRNG[495])|(((m[200]&m[396]&~m[884]))&~BiasedRNG[495])|((m[200]&m[396]&m[884]))):InitCond[704];
    m[593] = run?((((m[214]&~m[397]&m[924])|(~m[214]&m[397]&m[924]))&BiasedRNG[496])|(((m[214]&m[397]&~m[924]))&~BiasedRNG[496])|((m[214]&m[397]&m[924]))):InitCond[705];
    m[602] = run?((((m[145]&~m[406]&m[799])|(~m[145]&m[406]&m[799]))&BiasedRNG[497])|(((m[145]&m[406]&~m[799]))&~BiasedRNG[497])|((m[145]&m[406]&m[799]))):InitCond[706];
    m[603] = run?((((m[159]&~m[407]&m[824])|(~m[159]&m[407]&m[824]))&BiasedRNG[498])|(((m[159]&m[407]&~m[824]))&~BiasedRNG[498])|((m[159]&m[407]&m[824]))):InitCond[707];
    m[604] = run?((((m[173]&~m[408]&m[854])|(~m[173]&m[408]&m[854]))&BiasedRNG[499])|(((m[173]&m[408]&~m[854]))&~BiasedRNG[499])|((m[173]&m[408]&m[854]))):InitCond[708];
    m[605] = run?((((m[187]&~m[409]&m[889])|(~m[187]&m[409]&m[889]))&BiasedRNG[500])|(((m[187]&m[409]&~m[889]))&~BiasedRNG[500])|((m[187]&m[409]&m[889]))):InitCond[709];
    m[606] = run?((((m[201]&~m[410]&m[929])|(~m[201]&m[410]&m[929]))&BiasedRNG[501])|(((m[201]&m[410]&~m[929]))&~BiasedRNG[501])|((m[201]&m[410]&m[929]))):InitCond[710];
    m[607] = run?((((m[215]&~m[411]&m[974])|(~m[215]&m[411]&m[974]))&BiasedRNG[502])|(((m[215]&m[411]&~m[974]))&~BiasedRNG[502])|((m[215]&m[411]&m[974]))):InitCond[711];
    m[735] = run?((((m[732]&~m[733]&~m[734]&~m[736]&~m[737])|(~m[732]&~m[733]&~m[734]&m[736]&~m[737])|(m[732]&m[733]&~m[734]&m[736]&~m[737])|(m[732]&~m[733]&m[734]&m[736]&~m[737])|(~m[732]&m[733]&~m[734]&~m[736]&m[737])|(~m[732]&~m[733]&m[734]&~m[736]&m[737])|(m[732]&m[733]&m[734]&~m[736]&m[737])|(~m[732]&m[733]&m[734]&m[736]&m[737]))&UnbiasedRNG[209])|((m[732]&~m[733]&~m[734]&m[736]&~m[737])|(~m[732]&~m[733]&~m[734]&~m[736]&m[737])|(m[732]&~m[733]&~m[734]&~m[736]&m[737])|(m[732]&m[733]&~m[734]&~m[736]&m[737])|(m[732]&~m[733]&m[734]&~m[736]&m[737])|(~m[732]&~m[733]&~m[734]&m[736]&m[737])|(m[732]&~m[733]&~m[734]&m[736]&m[737])|(~m[732]&m[733]&~m[734]&m[736]&m[737])|(m[732]&m[733]&~m[734]&m[736]&m[737])|(~m[732]&~m[733]&m[734]&m[736]&m[737])|(m[732]&~m[733]&m[734]&m[736]&m[737])|(m[732]&m[733]&m[734]&m[736]&m[737]))):InitCond[712];
    m[745] = run?((((m[737]&~m[743]&~m[744]&~m[746]&~m[747])|(~m[737]&~m[743]&~m[744]&m[746]&~m[747])|(m[737]&m[743]&~m[744]&m[746]&~m[747])|(m[737]&~m[743]&m[744]&m[746]&~m[747])|(~m[737]&m[743]&~m[744]&~m[746]&m[747])|(~m[737]&~m[743]&m[744]&~m[746]&m[747])|(m[737]&m[743]&m[744]&~m[746]&m[747])|(~m[737]&m[743]&m[744]&m[746]&m[747]))&UnbiasedRNG[210])|((m[737]&~m[743]&~m[744]&m[746]&~m[747])|(~m[737]&~m[743]&~m[744]&~m[746]&m[747])|(m[737]&~m[743]&~m[744]&~m[746]&m[747])|(m[737]&m[743]&~m[744]&~m[746]&m[747])|(m[737]&~m[743]&m[744]&~m[746]&m[747])|(~m[737]&~m[743]&~m[744]&m[746]&m[747])|(m[737]&~m[743]&~m[744]&m[746]&m[747])|(~m[737]&m[743]&~m[744]&m[746]&m[747])|(m[737]&m[743]&~m[744]&m[746]&m[747])|(~m[737]&~m[743]&m[744]&m[746]&m[747])|(m[737]&~m[743]&m[744]&m[746]&m[747])|(m[737]&m[743]&m[744]&m[746]&m[747]))):InitCond[713];
    m[750] = run?((((m[742]&~m[748]&~m[749]&~m[751]&~m[752])|(~m[742]&~m[748]&~m[749]&m[751]&~m[752])|(m[742]&m[748]&~m[749]&m[751]&~m[752])|(m[742]&~m[748]&m[749]&m[751]&~m[752])|(~m[742]&m[748]&~m[749]&~m[751]&m[752])|(~m[742]&~m[748]&m[749]&~m[751]&m[752])|(m[742]&m[748]&m[749]&~m[751]&m[752])|(~m[742]&m[748]&m[749]&m[751]&m[752]))&UnbiasedRNG[211])|((m[742]&~m[748]&~m[749]&m[751]&~m[752])|(~m[742]&~m[748]&~m[749]&~m[751]&m[752])|(m[742]&~m[748]&~m[749]&~m[751]&m[752])|(m[742]&m[748]&~m[749]&~m[751]&m[752])|(m[742]&~m[748]&m[749]&~m[751]&m[752])|(~m[742]&~m[748]&~m[749]&m[751]&m[752])|(m[742]&~m[748]&~m[749]&m[751]&m[752])|(~m[742]&m[748]&~m[749]&m[751]&m[752])|(m[742]&m[748]&~m[749]&m[751]&m[752])|(~m[742]&~m[748]&m[749]&m[751]&m[752])|(m[742]&~m[748]&m[749]&m[751]&m[752])|(m[742]&m[748]&m[749]&m[751]&m[752]))):InitCond[714];
    m[760] = run?((((m[747]&~m[758]&~m[759]&~m[761]&~m[762])|(~m[747]&~m[758]&~m[759]&m[761]&~m[762])|(m[747]&m[758]&~m[759]&m[761]&~m[762])|(m[747]&~m[758]&m[759]&m[761]&~m[762])|(~m[747]&m[758]&~m[759]&~m[761]&m[762])|(~m[747]&~m[758]&m[759]&~m[761]&m[762])|(m[747]&m[758]&m[759]&~m[761]&m[762])|(~m[747]&m[758]&m[759]&m[761]&m[762]))&UnbiasedRNG[212])|((m[747]&~m[758]&~m[759]&m[761]&~m[762])|(~m[747]&~m[758]&~m[759]&~m[761]&m[762])|(m[747]&~m[758]&~m[759]&~m[761]&m[762])|(m[747]&m[758]&~m[759]&~m[761]&m[762])|(m[747]&~m[758]&m[759]&~m[761]&m[762])|(~m[747]&~m[758]&~m[759]&m[761]&m[762])|(m[747]&~m[758]&~m[759]&m[761]&m[762])|(~m[747]&m[758]&~m[759]&m[761]&m[762])|(m[747]&m[758]&~m[759]&m[761]&m[762])|(~m[747]&~m[758]&m[759]&m[761]&m[762])|(m[747]&~m[758]&m[759]&m[761]&m[762])|(m[747]&m[758]&m[759]&m[761]&m[762]))):InitCond[715];
    m[765] = run?((((m[752]&~m[763]&~m[764]&~m[766]&~m[767])|(~m[752]&~m[763]&~m[764]&m[766]&~m[767])|(m[752]&m[763]&~m[764]&m[766]&~m[767])|(m[752]&~m[763]&m[764]&m[766]&~m[767])|(~m[752]&m[763]&~m[764]&~m[766]&m[767])|(~m[752]&~m[763]&m[764]&~m[766]&m[767])|(m[752]&m[763]&m[764]&~m[766]&m[767])|(~m[752]&m[763]&m[764]&m[766]&m[767]))&UnbiasedRNG[213])|((m[752]&~m[763]&~m[764]&m[766]&~m[767])|(~m[752]&~m[763]&~m[764]&~m[766]&m[767])|(m[752]&~m[763]&~m[764]&~m[766]&m[767])|(m[752]&m[763]&~m[764]&~m[766]&m[767])|(m[752]&~m[763]&m[764]&~m[766]&m[767])|(~m[752]&~m[763]&~m[764]&m[766]&m[767])|(m[752]&~m[763]&~m[764]&m[766]&m[767])|(~m[752]&m[763]&~m[764]&m[766]&m[767])|(m[752]&m[763]&~m[764]&m[766]&m[767])|(~m[752]&~m[763]&m[764]&m[766]&m[767])|(m[752]&~m[763]&m[764]&m[766]&m[767])|(m[752]&m[763]&m[764]&m[766]&m[767]))):InitCond[716];
    m[770] = run?((((m[757]&~m[768]&~m[769]&~m[771]&~m[772])|(~m[757]&~m[768]&~m[769]&m[771]&~m[772])|(m[757]&m[768]&~m[769]&m[771]&~m[772])|(m[757]&~m[768]&m[769]&m[771]&~m[772])|(~m[757]&m[768]&~m[769]&~m[771]&m[772])|(~m[757]&~m[768]&m[769]&~m[771]&m[772])|(m[757]&m[768]&m[769]&~m[771]&m[772])|(~m[757]&m[768]&m[769]&m[771]&m[772]))&UnbiasedRNG[214])|((m[757]&~m[768]&~m[769]&m[771]&~m[772])|(~m[757]&~m[768]&~m[769]&~m[771]&m[772])|(m[757]&~m[768]&~m[769]&~m[771]&m[772])|(m[757]&m[768]&~m[769]&~m[771]&m[772])|(m[757]&~m[768]&m[769]&~m[771]&m[772])|(~m[757]&~m[768]&~m[769]&m[771]&m[772])|(m[757]&~m[768]&~m[769]&m[771]&m[772])|(~m[757]&m[768]&~m[769]&m[771]&m[772])|(m[757]&m[768]&~m[769]&m[771]&m[772])|(~m[757]&~m[768]&m[769]&m[771]&m[772])|(m[757]&~m[768]&m[769]&m[771]&m[772])|(m[757]&m[768]&m[769]&m[771]&m[772]))):InitCond[717];
    m[780] = run?((((m[762]&~m[778]&~m[779]&~m[781]&~m[782])|(~m[762]&~m[778]&~m[779]&m[781]&~m[782])|(m[762]&m[778]&~m[779]&m[781]&~m[782])|(m[762]&~m[778]&m[779]&m[781]&~m[782])|(~m[762]&m[778]&~m[779]&~m[781]&m[782])|(~m[762]&~m[778]&m[779]&~m[781]&m[782])|(m[762]&m[778]&m[779]&~m[781]&m[782])|(~m[762]&m[778]&m[779]&m[781]&m[782]))&UnbiasedRNG[215])|((m[762]&~m[778]&~m[779]&m[781]&~m[782])|(~m[762]&~m[778]&~m[779]&~m[781]&m[782])|(m[762]&~m[778]&~m[779]&~m[781]&m[782])|(m[762]&m[778]&~m[779]&~m[781]&m[782])|(m[762]&~m[778]&m[779]&~m[781]&m[782])|(~m[762]&~m[778]&~m[779]&m[781]&m[782])|(m[762]&~m[778]&~m[779]&m[781]&m[782])|(~m[762]&m[778]&~m[779]&m[781]&m[782])|(m[762]&m[778]&~m[779]&m[781]&m[782])|(~m[762]&~m[778]&m[779]&m[781]&m[782])|(m[762]&~m[778]&m[779]&m[781]&m[782])|(m[762]&m[778]&m[779]&m[781]&m[782]))):InitCond[718];
    m[785] = run?((((m[767]&~m[783]&~m[784]&~m[786]&~m[787])|(~m[767]&~m[783]&~m[784]&m[786]&~m[787])|(m[767]&m[783]&~m[784]&m[786]&~m[787])|(m[767]&~m[783]&m[784]&m[786]&~m[787])|(~m[767]&m[783]&~m[784]&~m[786]&m[787])|(~m[767]&~m[783]&m[784]&~m[786]&m[787])|(m[767]&m[783]&m[784]&~m[786]&m[787])|(~m[767]&m[783]&m[784]&m[786]&m[787]))&UnbiasedRNG[216])|((m[767]&~m[783]&~m[784]&m[786]&~m[787])|(~m[767]&~m[783]&~m[784]&~m[786]&m[787])|(m[767]&~m[783]&~m[784]&~m[786]&m[787])|(m[767]&m[783]&~m[784]&~m[786]&m[787])|(m[767]&~m[783]&m[784]&~m[786]&m[787])|(~m[767]&~m[783]&~m[784]&m[786]&m[787])|(m[767]&~m[783]&~m[784]&m[786]&m[787])|(~m[767]&m[783]&~m[784]&m[786]&m[787])|(m[767]&m[783]&~m[784]&m[786]&m[787])|(~m[767]&~m[783]&m[784]&m[786]&m[787])|(m[767]&~m[783]&m[784]&m[786]&m[787])|(m[767]&m[783]&m[784]&m[786]&m[787]))):InitCond[719];
    m[790] = run?((((m[772]&~m[788]&~m[789]&~m[791]&~m[792])|(~m[772]&~m[788]&~m[789]&m[791]&~m[792])|(m[772]&m[788]&~m[789]&m[791]&~m[792])|(m[772]&~m[788]&m[789]&m[791]&~m[792])|(~m[772]&m[788]&~m[789]&~m[791]&m[792])|(~m[772]&~m[788]&m[789]&~m[791]&m[792])|(m[772]&m[788]&m[789]&~m[791]&m[792])|(~m[772]&m[788]&m[789]&m[791]&m[792]))&UnbiasedRNG[217])|((m[772]&~m[788]&~m[789]&m[791]&~m[792])|(~m[772]&~m[788]&~m[789]&~m[791]&m[792])|(m[772]&~m[788]&~m[789]&~m[791]&m[792])|(m[772]&m[788]&~m[789]&~m[791]&m[792])|(m[772]&~m[788]&m[789]&~m[791]&m[792])|(~m[772]&~m[788]&~m[789]&m[791]&m[792])|(m[772]&~m[788]&~m[789]&m[791]&m[792])|(~m[772]&m[788]&~m[789]&m[791]&m[792])|(m[772]&m[788]&~m[789]&m[791]&m[792])|(~m[772]&~m[788]&m[789]&m[791]&m[792])|(m[772]&~m[788]&m[789]&m[791]&m[792])|(m[772]&m[788]&m[789]&m[791]&m[792]))):InitCond[720];
    m[795] = run?((((m[777]&~m[793]&~m[794]&~m[796]&~m[797])|(~m[777]&~m[793]&~m[794]&m[796]&~m[797])|(m[777]&m[793]&~m[794]&m[796]&~m[797])|(m[777]&~m[793]&m[794]&m[796]&~m[797])|(~m[777]&m[793]&~m[794]&~m[796]&m[797])|(~m[777]&~m[793]&m[794]&~m[796]&m[797])|(m[777]&m[793]&m[794]&~m[796]&m[797])|(~m[777]&m[793]&m[794]&m[796]&m[797]))&UnbiasedRNG[218])|((m[777]&~m[793]&~m[794]&m[796]&~m[797])|(~m[777]&~m[793]&~m[794]&~m[796]&m[797])|(m[777]&~m[793]&~m[794]&~m[796]&m[797])|(m[777]&m[793]&~m[794]&~m[796]&m[797])|(m[777]&~m[793]&m[794]&~m[796]&m[797])|(~m[777]&~m[793]&~m[794]&m[796]&m[797])|(m[777]&~m[793]&~m[794]&m[796]&m[797])|(~m[777]&m[793]&~m[794]&m[796]&m[797])|(m[777]&m[793]&~m[794]&m[796]&m[797])|(~m[777]&~m[793]&m[794]&m[796]&m[797])|(m[777]&~m[793]&m[794]&m[796]&m[797])|(m[777]&m[793]&m[794]&m[796]&m[797]))):InitCond[721];
    m[805] = run?((((m[782]&~m[803]&~m[804]&~m[806]&~m[807])|(~m[782]&~m[803]&~m[804]&m[806]&~m[807])|(m[782]&m[803]&~m[804]&m[806]&~m[807])|(m[782]&~m[803]&m[804]&m[806]&~m[807])|(~m[782]&m[803]&~m[804]&~m[806]&m[807])|(~m[782]&~m[803]&m[804]&~m[806]&m[807])|(m[782]&m[803]&m[804]&~m[806]&m[807])|(~m[782]&m[803]&m[804]&m[806]&m[807]))&UnbiasedRNG[219])|((m[782]&~m[803]&~m[804]&m[806]&~m[807])|(~m[782]&~m[803]&~m[804]&~m[806]&m[807])|(m[782]&~m[803]&~m[804]&~m[806]&m[807])|(m[782]&m[803]&~m[804]&~m[806]&m[807])|(m[782]&~m[803]&m[804]&~m[806]&m[807])|(~m[782]&~m[803]&~m[804]&m[806]&m[807])|(m[782]&~m[803]&~m[804]&m[806]&m[807])|(~m[782]&m[803]&~m[804]&m[806]&m[807])|(m[782]&m[803]&~m[804]&m[806]&m[807])|(~m[782]&~m[803]&m[804]&m[806]&m[807])|(m[782]&~m[803]&m[804]&m[806]&m[807])|(m[782]&m[803]&m[804]&m[806]&m[807]))):InitCond[722];
    m[810] = run?((((m[787]&~m[808]&~m[809]&~m[811]&~m[812])|(~m[787]&~m[808]&~m[809]&m[811]&~m[812])|(m[787]&m[808]&~m[809]&m[811]&~m[812])|(m[787]&~m[808]&m[809]&m[811]&~m[812])|(~m[787]&m[808]&~m[809]&~m[811]&m[812])|(~m[787]&~m[808]&m[809]&~m[811]&m[812])|(m[787]&m[808]&m[809]&~m[811]&m[812])|(~m[787]&m[808]&m[809]&m[811]&m[812]))&UnbiasedRNG[220])|((m[787]&~m[808]&~m[809]&m[811]&~m[812])|(~m[787]&~m[808]&~m[809]&~m[811]&m[812])|(m[787]&~m[808]&~m[809]&~m[811]&m[812])|(m[787]&m[808]&~m[809]&~m[811]&m[812])|(m[787]&~m[808]&m[809]&~m[811]&m[812])|(~m[787]&~m[808]&~m[809]&m[811]&m[812])|(m[787]&~m[808]&~m[809]&m[811]&m[812])|(~m[787]&m[808]&~m[809]&m[811]&m[812])|(m[787]&m[808]&~m[809]&m[811]&m[812])|(~m[787]&~m[808]&m[809]&m[811]&m[812])|(m[787]&~m[808]&m[809]&m[811]&m[812])|(m[787]&m[808]&m[809]&m[811]&m[812]))):InitCond[723];
    m[815] = run?((((m[792]&~m[813]&~m[814]&~m[816]&~m[817])|(~m[792]&~m[813]&~m[814]&m[816]&~m[817])|(m[792]&m[813]&~m[814]&m[816]&~m[817])|(m[792]&~m[813]&m[814]&m[816]&~m[817])|(~m[792]&m[813]&~m[814]&~m[816]&m[817])|(~m[792]&~m[813]&m[814]&~m[816]&m[817])|(m[792]&m[813]&m[814]&~m[816]&m[817])|(~m[792]&m[813]&m[814]&m[816]&m[817]))&UnbiasedRNG[221])|((m[792]&~m[813]&~m[814]&m[816]&~m[817])|(~m[792]&~m[813]&~m[814]&~m[816]&m[817])|(m[792]&~m[813]&~m[814]&~m[816]&m[817])|(m[792]&m[813]&~m[814]&~m[816]&m[817])|(m[792]&~m[813]&m[814]&~m[816]&m[817])|(~m[792]&~m[813]&~m[814]&m[816]&m[817])|(m[792]&~m[813]&~m[814]&m[816]&m[817])|(~m[792]&m[813]&~m[814]&m[816]&m[817])|(m[792]&m[813]&~m[814]&m[816]&m[817])|(~m[792]&~m[813]&m[814]&m[816]&m[817])|(m[792]&~m[813]&m[814]&m[816]&m[817])|(m[792]&m[813]&m[814]&m[816]&m[817]))):InitCond[724];
    m[820] = run?((((m[797]&~m[818]&~m[819]&~m[821]&~m[822])|(~m[797]&~m[818]&~m[819]&m[821]&~m[822])|(m[797]&m[818]&~m[819]&m[821]&~m[822])|(m[797]&~m[818]&m[819]&m[821]&~m[822])|(~m[797]&m[818]&~m[819]&~m[821]&m[822])|(~m[797]&~m[818]&m[819]&~m[821]&m[822])|(m[797]&m[818]&m[819]&~m[821]&m[822])|(~m[797]&m[818]&m[819]&m[821]&m[822]))&UnbiasedRNG[222])|((m[797]&~m[818]&~m[819]&m[821]&~m[822])|(~m[797]&~m[818]&~m[819]&~m[821]&m[822])|(m[797]&~m[818]&~m[819]&~m[821]&m[822])|(m[797]&m[818]&~m[819]&~m[821]&m[822])|(m[797]&~m[818]&m[819]&~m[821]&m[822])|(~m[797]&~m[818]&~m[819]&m[821]&m[822])|(m[797]&~m[818]&~m[819]&m[821]&m[822])|(~m[797]&m[818]&~m[819]&m[821]&m[822])|(m[797]&m[818]&~m[819]&m[821]&m[822])|(~m[797]&~m[818]&m[819]&m[821]&m[822])|(m[797]&~m[818]&m[819]&m[821]&m[822])|(m[797]&m[818]&m[819]&m[821]&m[822]))):InitCond[725];
    m[825] = run?((((m[802]&~m[823]&~m[824]&~m[826]&~m[827])|(~m[802]&~m[823]&~m[824]&m[826]&~m[827])|(m[802]&m[823]&~m[824]&m[826]&~m[827])|(m[802]&~m[823]&m[824]&m[826]&~m[827])|(~m[802]&m[823]&~m[824]&~m[826]&m[827])|(~m[802]&~m[823]&m[824]&~m[826]&m[827])|(m[802]&m[823]&m[824]&~m[826]&m[827])|(~m[802]&m[823]&m[824]&m[826]&m[827]))&UnbiasedRNG[223])|((m[802]&~m[823]&~m[824]&m[826]&~m[827])|(~m[802]&~m[823]&~m[824]&~m[826]&m[827])|(m[802]&~m[823]&~m[824]&~m[826]&m[827])|(m[802]&m[823]&~m[824]&~m[826]&m[827])|(m[802]&~m[823]&m[824]&~m[826]&m[827])|(~m[802]&~m[823]&~m[824]&m[826]&m[827])|(m[802]&~m[823]&~m[824]&m[826]&m[827])|(~m[802]&m[823]&~m[824]&m[826]&m[827])|(m[802]&m[823]&~m[824]&m[826]&m[827])|(~m[802]&~m[823]&m[824]&m[826]&m[827])|(m[802]&~m[823]&m[824]&m[826]&m[827])|(m[802]&m[823]&m[824]&m[826]&m[827]))):InitCond[726];
    m[829] = run?((((m[616]&~m[828]&~m[830]&~m[831]&~m[832])|(~m[616]&~m[828]&~m[830]&m[831]&~m[832])|(m[616]&m[828]&~m[830]&m[831]&~m[832])|(m[616]&~m[828]&m[830]&m[831]&~m[832])|(~m[616]&m[828]&~m[830]&~m[831]&m[832])|(~m[616]&~m[828]&m[830]&~m[831]&m[832])|(m[616]&m[828]&m[830]&~m[831]&m[832])|(~m[616]&m[828]&m[830]&m[831]&m[832]))&UnbiasedRNG[224])|((m[616]&~m[828]&~m[830]&m[831]&~m[832])|(~m[616]&~m[828]&~m[830]&~m[831]&m[832])|(m[616]&~m[828]&~m[830]&~m[831]&m[832])|(m[616]&m[828]&~m[830]&~m[831]&m[832])|(m[616]&~m[828]&m[830]&~m[831]&m[832])|(~m[616]&~m[828]&~m[830]&m[831]&m[832])|(m[616]&~m[828]&~m[830]&m[831]&m[832])|(~m[616]&m[828]&~m[830]&m[831]&m[832])|(m[616]&m[828]&~m[830]&m[831]&m[832])|(~m[616]&~m[828]&m[830]&m[831]&m[832])|(m[616]&~m[828]&m[830]&m[831]&m[832])|(m[616]&m[828]&m[830]&m[831]&m[832]))):InitCond[727];
    m[834] = run?((((m[552]&~m[833]&~m[835]&~m[836]&~m[837])|(~m[552]&~m[833]&~m[835]&m[836]&~m[837])|(m[552]&m[833]&~m[835]&m[836]&~m[837])|(m[552]&~m[833]&m[835]&m[836]&~m[837])|(~m[552]&m[833]&~m[835]&~m[836]&m[837])|(~m[552]&~m[833]&m[835]&~m[836]&m[837])|(m[552]&m[833]&m[835]&~m[836]&m[837])|(~m[552]&m[833]&m[835]&m[836]&m[837]))&UnbiasedRNG[225])|((m[552]&~m[833]&~m[835]&m[836]&~m[837])|(~m[552]&~m[833]&~m[835]&~m[836]&m[837])|(m[552]&~m[833]&~m[835]&~m[836]&m[837])|(m[552]&m[833]&~m[835]&~m[836]&m[837])|(m[552]&~m[833]&m[835]&~m[836]&m[837])|(~m[552]&~m[833]&~m[835]&m[836]&m[837])|(m[552]&~m[833]&~m[835]&m[836]&m[837])|(~m[552]&m[833]&~m[835]&m[836]&m[837])|(m[552]&m[833]&~m[835]&m[836]&m[837])|(~m[552]&~m[833]&m[835]&m[836]&m[837])|(m[552]&~m[833]&m[835]&m[836]&m[837])|(m[552]&m[833]&m[835]&m[836]&m[837]))):InitCond[728];
    m[840] = run?((((m[812]&~m[838]&~m[839]&~m[841]&~m[842])|(~m[812]&~m[838]&~m[839]&m[841]&~m[842])|(m[812]&m[838]&~m[839]&m[841]&~m[842])|(m[812]&~m[838]&m[839]&m[841]&~m[842])|(~m[812]&m[838]&~m[839]&~m[841]&m[842])|(~m[812]&~m[838]&m[839]&~m[841]&m[842])|(m[812]&m[838]&m[839]&~m[841]&m[842])|(~m[812]&m[838]&m[839]&m[841]&m[842]))&UnbiasedRNG[226])|((m[812]&~m[838]&~m[839]&m[841]&~m[842])|(~m[812]&~m[838]&~m[839]&~m[841]&m[842])|(m[812]&~m[838]&~m[839]&~m[841]&m[842])|(m[812]&m[838]&~m[839]&~m[841]&m[842])|(m[812]&~m[838]&m[839]&~m[841]&m[842])|(~m[812]&~m[838]&~m[839]&m[841]&m[842])|(m[812]&~m[838]&~m[839]&m[841]&m[842])|(~m[812]&m[838]&~m[839]&m[841]&m[842])|(m[812]&m[838]&~m[839]&m[841]&m[842])|(~m[812]&~m[838]&m[839]&m[841]&m[842])|(m[812]&~m[838]&m[839]&m[841]&m[842])|(m[812]&m[838]&m[839]&m[841]&m[842]))):InitCond[729];
    m[845] = run?((((m[817]&~m[843]&~m[844]&~m[846]&~m[847])|(~m[817]&~m[843]&~m[844]&m[846]&~m[847])|(m[817]&m[843]&~m[844]&m[846]&~m[847])|(m[817]&~m[843]&m[844]&m[846]&~m[847])|(~m[817]&m[843]&~m[844]&~m[846]&m[847])|(~m[817]&~m[843]&m[844]&~m[846]&m[847])|(m[817]&m[843]&m[844]&~m[846]&m[847])|(~m[817]&m[843]&m[844]&m[846]&m[847]))&UnbiasedRNG[227])|((m[817]&~m[843]&~m[844]&m[846]&~m[847])|(~m[817]&~m[843]&~m[844]&~m[846]&m[847])|(m[817]&~m[843]&~m[844]&~m[846]&m[847])|(m[817]&m[843]&~m[844]&~m[846]&m[847])|(m[817]&~m[843]&m[844]&~m[846]&m[847])|(~m[817]&~m[843]&~m[844]&m[846]&m[847])|(m[817]&~m[843]&~m[844]&m[846]&m[847])|(~m[817]&m[843]&~m[844]&m[846]&m[847])|(m[817]&m[843]&~m[844]&m[846]&m[847])|(~m[817]&~m[843]&m[844]&m[846]&m[847])|(m[817]&~m[843]&m[844]&m[846]&m[847])|(m[817]&m[843]&m[844]&m[846]&m[847]))):InitCond[730];
    m[850] = run?((((m[822]&~m[848]&~m[849]&~m[851]&~m[852])|(~m[822]&~m[848]&~m[849]&m[851]&~m[852])|(m[822]&m[848]&~m[849]&m[851]&~m[852])|(m[822]&~m[848]&m[849]&m[851]&~m[852])|(~m[822]&m[848]&~m[849]&~m[851]&m[852])|(~m[822]&~m[848]&m[849]&~m[851]&m[852])|(m[822]&m[848]&m[849]&~m[851]&m[852])|(~m[822]&m[848]&m[849]&m[851]&m[852]))&UnbiasedRNG[228])|((m[822]&~m[848]&~m[849]&m[851]&~m[852])|(~m[822]&~m[848]&~m[849]&~m[851]&m[852])|(m[822]&~m[848]&~m[849]&~m[851]&m[852])|(m[822]&m[848]&~m[849]&~m[851]&m[852])|(m[822]&~m[848]&m[849]&~m[851]&m[852])|(~m[822]&~m[848]&~m[849]&m[851]&m[852])|(m[822]&~m[848]&~m[849]&m[851]&m[852])|(~m[822]&m[848]&~m[849]&m[851]&m[852])|(m[822]&m[848]&~m[849]&m[851]&m[852])|(~m[822]&~m[848]&m[849]&m[851]&m[852])|(m[822]&~m[848]&m[849]&m[851]&m[852])|(m[822]&m[848]&m[849]&m[851]&m[852]))):InitCond[731];
    m[855] = run?((((m[827]&~m[853]&~m[854]&~m[856]&~m[857])|(~m[827]&~m[853]&~m[854]&m[856]&~m[857])|(m[827]&m[853]&~m[854]&m[856]&~m[857])|(m[827]&~m[853]&m[854]&m[856]&~m[857])|(~m[827]&m[853]&~m[854]&~m[856]&m[857])|(~m[827]&~m[853]&m[854]&~m[856]&m[857])|(m[827]&m[853]&m[854]&~m[856]&m[857])|(~m[827]&m[853]&m[854]&m[856]&m[857]))&UnbiasedRNG[229])|((m[827]&~m[853]&~m[854]&m[856]&~m[857])|(~m[827]&~m[853]&~m[854]&~m[856]&m[857])|(m[827]&~m[853]&~m[854]&~m[856]&m[857])|(m[827]&m[853]&~m[854]&~m[856]&m[857])|(m[827]&~m[853]&m[854]&~m[856]&m[857])|(~m[827]&~m[853]&~m[854]&m[856]&m[857])|(m[827]&~m[853]&~m[854]&m[856]&m[857])|(~m[827]&m[853]&~m[854]&m[856]&m[857])|(m[827]&m[853]&~m[854]&m[856]&m[857])|(~m[827]&~m[853]&m[854]&m[856]&m[857])|(m[827]&~m[853]&m[854]&m[856]&m[857])|(m[827]&m[853]&m[854]&m[856]&m[857]))):InitCond[732];
    m[859] = run?((((m[617]&~m[858]&~m[860]&~m[861]&~m[862])|(~m[617]&~m[858]&~m[860]&m[861]&~m[862])|(m[617]&m[858]&~m[860]&m[861]&~m[862])|(m[617]&~m[858]&m[860]&m[861]&~m[862])|(~m[617]&m[858]&~m[860]&~m[861]&m[862])|(~m[617]&~m[858]&m[860]&~m[861]&m[862])|(m[617]&m[858]&m[860]&~m[861]&m[862])|(~m[617]&m[858]&m[860]&m[861]&m[862]))&UnbiasedRNG[230])|((m[617]&~m[858]&~m[860]&m[861]&~m[862])|(~m[617]&~m[858]&~m[860]&~m[861]&m[862])|(m[617]&~m[858]&~m[860]&~m[861]&m[862])|(m[617]&m[858]&~m[860]&~m[861]&m[862])|(m[617]&~m[858]&m[860]&~m[861]&m[862])|(~m[617]&~m[858]&~m[860]&m[861]&m[862])|(m[617]&~m[858]&~m[860]&m[861]&m[862])|(~m[617]&m[858]&~m[860]&m[861]&m[862])|(m[617]&m[858]&~m[860]&m[861]&m[862])|(~m[617]&~m[858]&m[860]&m[861]&m[862])|(m[617]&~m[858]&m[860]&m[861]&m[862])|(m[617]&m[858]&m[860]&m[861]&m[862]))):InitCond[733];
    m[864] = run?((((m[630]&~m[863]&~m[865]&~m[866]&~m[867])|(~m[630]&~m[863]&~m[865]&m[866]&~m[867])|(m[630]&m[863]&~m[865]&m[866]&~m[867])|(m[630]&~m[863]&m[865]&m[866]&~m[867])|(~m[630]&m[863]&~m[865]&~m[866]&m[867])|(~m[630]&~m[863]&m[865]&~m[866]&m[867])|(m[630]&m[863]&m[865]&~m[866]&m[867])|(~m[630]&m[863]&m[865]&m[866]&m[867]))&UnbiasedRNG[231])|((m[630]&~m[863]&~m[865]&m[866]&~m[867])|(~m[630]&~m[863]&~m[865]&~m[866]&m[867])|(m[630]&~m[863]&~m[865]&~m[866]&m[867])|(m[630]&m[863]&~m[865]&~m[866]&m[867])|(m[630]&~m[863]&m[865]&~m[866]&m[867])|(~m[630]&~m[863]&~m[865]&m[866]&m[867])|(m[630]&~m[863]&~m[865]&m[866]&m[867])|(~m[630]&m[863]&~m[865]&m[866]&m[867])|(m[630]&m[863]&~m[865]&m[866]&m[867])|(~m[630]&~m[863]&m[865]&m[866]&m[867])|(m[630]&~m[863]&m[865]&m[866]&m[867])|(m[630]&m[863]&m[865]&m[866]&m[867]))):InitCond[734];
    m[869] = run?((((m[553]&~m[868]&~m[870]&~m[871]&~m[872])|(~m[553]&~m[868]&~m[870]&m[871]&~m[872])|(m[553]&m[868]&~m[870]&m[871]&~m[872])|(m[553]&~m[868]&m[870]&m[871]&~m[872])|(~m[553]&m[868]&~m[870]&~m[871]&m[872])|(~m[553]&~m[868]&m[870]&~m[871]&m[872])|(m[553]&m[868]&m[870]&~m[871]&m[872])|(~m[553]&m[868]&m[870]&m[871]&m[872]))&UnbiasedRNG[232])|((m[553]&~m[868]&~m[870]&m[871]&~m[872])|(~m[553]&~m[868]&~m[870]&~m[871]&m[872])|(m[553]&~m[868]&~m[870]&~m[871]&m[872])|(m[553]&m[868]&~m[870]&~m[871]&m[872])|(m[553]&~m[868]&m[870]&~m[871]&m[872])|(~m[553]&~m[868]&~m[870]&m[871]&m[872])|(m[553]&~m[868]&~m[870]&m[871]&m[872])|(~m[553]&m[868]&~m[870]&m[871]&m[872])|(m[553]&m[868]&~m[870]&m[871]&m[872])|(~m[553]&~m[868]&m[870]&m[871]&m[872])|(m[553]&~m[868]&m[870]&m[871]&m[872])|(m[553]&m[868]&m[870]&m[871]&m[872]))):InitCond[735];
    m[874] = run?((((m[566]&~m[873]&~m[875]&~m[876]&~m[877])|(~m[566]&~m[873]&~m[875]&m[876]&~m[877])|(m[566]&m[873]&~m[875]&m[876]&~m[877])|(m[566]&~m[873]&m[875]&m[876]&~m[877])|(~m[566]&m[873]&~m[875]&~m[876]&m[877])|(~m[566]&~m[873]&m[875]&~m[876]&m[877])|(m[566]&m[873]&m[875]&~m[876]&m[877])|(~m[566]&m[873]&m[875]&m[876]&m[877]))&UnbiasedRNG[233])|((m[566]&~m[873]&~m[875]&m[876]&~m[877])|(~m[566]&~m[873]&~m[875]&~m[876]&m[877])|(m[566]&~m[873]&~m[875]&~m[876]&m[877])|(m[566]&m[873]&~m[875]&~m[876]&m[877])|(m[566]&~m[873]&m[875]&~m[876]&m[877])|(~m[566]&~m[873]&~m[875]&m[876]&m[877])|(m[566]&~m[873]&~m[875]&m[876]&m[877])|(~m[566]&m[873]&~m[875]&m[876]&m[877])|(m[566]&m[873]&~m[875]&m[876]&m[877])|(~m[566]&~m[873]&m[875]&m[876]&m[877])|(m[566]&~m[873]&m[875]&m[876]&m[877])|(m[566]&m[873]&m[875]&m[876]&m[877]))):InitCond[736];
    m[880] = run?((((m[847]&~m[878]&~m[879]&~m[881]&~m[882])|(~m[847]&~m[878]&~m[879]&m[881]&~m[882])|(m[847]&m[878]&~m[879]&m[881]&~m[882])|(m[847]&~m[878]&m[879]&m[881]&~m[882])|(~m[847]&m[878]&~m[879]&~m[881]&m[882])|(~m[847]&~m[878]&m[879]&~m[881]&m[882])|(m[847]&m[878]&m[879]&~m[881]&m[882])|(~m[847]&m[878]&m[879]&m[881]&m[882]))&UnbiasedRNG[234])|((m[847]&~m[878]&~m[879]&m[881]&~m[882])|(~m[847]&~m[878]&~m[879]&~m[881]&m[882])|(m[847]&~m[878]&~m[879]&~m[881]&m[882])|(m[847]&m[878]&~m[879]&~m[881]&m[882])|(m[847]&~m[878]&m[879]&~m[881]&m[882])|(~m[847]&~m[878]&~m[879]&m[881]&m[882])|(m[847]&~m[878]&~m[879]&m[881]&m[882])|(~m[847]&m[878]&~m[879]&m[881]&m[882])|(m[847]&m[878]&~m[879]&m[881]&m[882])|(~m[847]&~m[878]&m[879]&m[881]&m[882])|(m[847]&~m[878]&m[879]&m[881]&m[882])|(m[847]&m[878]&m[879]&m[881]&m[882]))):InitCond[737];
    m[885] = run?((((m[852]&~m[883]&~m[884]&~m[886]&~m[887])|(~m[852]&~m[883]&~m[884]&m[886]&~m[887])|(m[852]&m[883]&~m[884]&m[886]&~m[887])|(m[852]&~m[883]&m[884]&m[886]&~m[887])|(~m[852]&m[883]&~m[884]&~m[886]&m[887])|(~m[852]&~m[883]&m[884]&~m[886]&m[887])|(m[852]&m[883]&m[884]&~m[886]&m[887])|(~m[852]&m[883]&m[884]&m[886]&m[887]))&UnbiasedRNG[235])|((m[852]&~m[883]&~m[884]&m[886]&~m[887])|(~m[852]&~m[883]&~m[884]&~m[886]&m[887])|(m[852]&~m[883]&~m[884]&~m[886]&m[887])|(m[852]&m[883]&~m[884]&~m[886]&m[887])|(m[852]&~m[883]&m[884]&~m[886]&m[887])|(~m[852]&~m[883]&~m[884]&m[886]&m[887])|(m[852]&~m[883]&~m[884]&m[886]&m[887])|(~m[852]&m[883]&~m[884]&m[886]&m[887])|(m[852]&m[883]&~m[884]&m[886]&m[887])|(~m[852]&~m[883]&m[884]&m[886]&m[887])|(m[852]&~m[883]&m[884]&m[886]&m[887])|(m[852]&m[883]&m[884]&m[886]&m[887]))):InitCond[738];
    m[890] = run?((((m[857]&~m[888]&~m[889]&~m[891]&~m[892])|(~m[857]&~m[888]&~m[889]&m[891]&~m[892])|(m[857]&m[888]&~m[889]&m[891]&~m[892])|(m[857]&~m[888]&m[889]&m[891]&~m[892])|(~m[857]&m[888]&~m[889]&~m[891]&m[892])|(~m[857]&~m[888]&m[889]&~m[891]&m[892])|(m[857]&m[888]&m[889]&~m[891]&m[892])|(~m[857]&m[888]&m[889]&m[891]&m[892]))&UnbiasedRNG[236])|((m[857]&~m[888]&~m[889]&m[891]&~m[892])|(~m[857]&~m[888]&~m[889]&~m[891]&m[892])|(m[857]&~m[888]&~m[889]&~m[891]&m[892])|(m[857]&m[888]&~m[889]&~m[891]&m[892])|(m[857]&~m[888]&m[889]&~m[891]&m[892])|(~m[857]&~m[888]&~m[889]&m[891]&m[892])|(m[857]&~m[888]&~m[889]&m[891]&m[892])|(~m[857]&m[888]&~m[889]&m[891]&m[892])|(m[857]&m[888]&~m[889]&m[891]&m[892])|(~m[857]&~m[888]&m[889]&m[891]&m[892])|(m[857]&~m[888]&m[889]&m[891]&m[892])|(m[857]&m[888]&m[889]&m[891]&m[892]))):InitCond[739];
    m[894] = run?((((m[618]&~m[893]&~m[895]&~m[896]&~m[897])|(~m[618]&~m[893]&~m[895]&m[896]&~m[897])|(m[618]&m[893]&~m[895]&m[896]&~m[897])|(m[618]&~m[893]&m[895]&m[896]&~m[897])|(~m[618]&m[893]&~m[895]&~m[896]&m[897])|(~m[618]&~m[893]&m[895]&~m[896]&m[897])|(m[618]&m[893]&m[895]&~m[896]&m[897])|(~m[618]&m[893]&m[895]&m[896]&m[897]))&UnbiasedRNG[237])|((m[618]&~m[893]&~m[895]&m[896]&~m[897])|(~m[618]&~m[893]&~m[895]&~m[896]&m[897])|(m[618]&~m[893]&~m[895]&~m[896]&m[897])|(m[618]&m[893]&~m[895]&~m[896]&m[897])|(m[618]&~m[893]&m[895]&~m[896]&m[897])|(~m[618]&~m[893]&~m[895]&m[896]&m[897])|(m[618]&~m[893]&~m[895]&m[896]&m[897])|(~m[618]&m[893]&~m[895]&m[896]&m[897])|(m[618]&m[893]&~m[895]&m[896]&m[897])|(~m[618]&~m[893]&m[895]&m[896]&m[897])|(m[618]&~m[893]&m[895]&m[896]&m[897])|(m[618]&m[893]&m[895]&m[896]&m[897]))):InitCond[740];
    m[899] = run?((((m[631]&~m[898]&~m[900]&~m[901]&~m[902])|(~m[631]&~m[898]&~m[900]&m[901]&~m[902])|(m[631]&m[898]&~m[900]&m[901]&~m[902])|(m[631]&~m[898]&m[900]&m[901]&~m[902])|(~m[631]&m[898]&~m[900]&~m[901]&m[902])|(~m[631]&~m[898]&m[900]&~m[901]&m[902])|(m[631]&m[898]&m[900]&~m[901]&m[902])|(~m[631]&m[898]&m[900]&m[901]&m[902]))&UnbiasedRNG[238])|((m[631]&~m[898]&~m[900]&m[901]&~m[902])|(~m[631]&~m[898]&~m[900]&~m[901]&m[902])|(m[631]&~m[898]&~m[900]&~m[901]&m[902])|(m[631]&m[898]&~m[900]&~m[901]&m[902])|(m[631]&~m[898]&m[900]&~m[901]&m[902])|(~m[631]&~m[898]&~m[900]&m[901]&m[902])|(m[631]&~m[898]&~m[900]&m[901]&m[902])|(~m[631]&m[898]&~m[900]&m[901]&m[902])|(m[631]&m[898]&~m[900]&m[901]&m[902])|(~m[631]&~m[898]&m[900]&m[901]&m[902])|(m[631]&~m[898]&m[900]&m[901]&m[902])|(m[631]&m[898]&m[900]&m[901]&m[902]))):InitCond[741];
    m[904] = run?((((m[644]&~m[903]&~m[905]&~m[906]&~m[907])|(~m[644]&~m[903]&~m[905]&m[906]&~m[907])|(m[644]&m[903]&~m[905]&m[906]&~m[907])|(m[644]&~m[903]&m[905]&m[906]&~m[907])|(~m[644]&m[903]&~m[905]&~m[906]&m[907])|(~m[644]&~m[903]&m[905]&~m[906]&m[907])|(m[644]&m[903]&m[905]&~m[906]&m[907])|(~m[644]&m[903]&m[905]&m[906]&m[907]))&UnbiasedRNG[239])|((m[644]&~m[903]&~m[905]&m[906]&~m[907])|(~m[644]&~m[903]&~m[905]&~m[906]&m[907])|(m[644]&~m[903]&~m[905]&~m[906]&m[907])|(m[644]&m[903]&~m[905]&~m[906]&m[907])|(m[644]&~m[903]&m[905]&~m[906]&m[907])|(~m[644]&~m[903]&~m[905]&m[906]&m[907])|(m[644]&~m[903]&~m[905]&m[906]&m[907])|(~m[644]&m[903]&~m[905]&m[906]&m[907])|(m[644]&m[903]&~m[905]&m[906]&m[907])|(~m[644]&~m[903]&m[905]&m[906]&m[907])|(m[644]&~m[903]&m[905]&m[906]&m[907])|(m[644]&m[903]&m[905]&m[906]&m[907]))):InitCond[742];
    m[909] = run?((((m[554]&~m[908]&~m[910]&~m[911]&~m[912])|(~m[554]&~m[908]&~m[910]&m[911]&~m[912])|(m[554]&m[908]&~m[910]&m[911]&~m[912])|(m[554]&~m[908]&m[910]&m[911]&~m[912])|(~m[554]&m[908]&~m[910]&~m[911]&m[912])|(~m[554]&~m[908]&m[910]&~m[911]&m[912])|(m[554]&m[908]&m[910]&~m[911]&m[912])|(~m[554]&m[908]&m[910]&m[911]&m[912]))&UnbiasedRNG[240])|((m[554]&~m[908]&~m[910]&m[911]&~m[912])|(~m[554]&~m[908]&~m[910]&~m[911]&m[912])|(m[554]&~m[908]&~m[910]&~m[911]&m[912])|(m[554]&m[908]&~m[910]&~m[911]&m[912])|(m[554]&~m[908]&m[910]&~m[911]&m[912])|(~m[554]&~m[908]&~m[910]&m[911]&m[912])|(m[554]&~m[908]&~m[910]&m[911]&m[912])|(~m[554]&m[908]&~m[910]&m[911]&m[912])|(m[554]&m[908]&~m[910]&m[911]&m[912])|(~m[554]&~m[908]&m[910]&m[911]&m[912])|(m[554]&~m[908]&m[910]&m[911]&m[912])|(m[554]&m[908]&m[910]&m[911]&m[912]))):InitCond[743];
    m[914] = run?((((m[567]&~m[913]&~m[915]&~m[916]&~m[917])|(~m[567]&~m[913]&~m[915]&m[916]&~m[917])|(m[567]&m[913]&~m[915]&m[916]&~m[917])|(m[567]&~m[913]&m[915]&m[916]&~m[917])|(~m[567]&m[913]&~m[915]&~m[916]&m[917])|(~m[567]&~m[913]&m[915]&~m[916]&m[917])|(m[567]&m[913]&m[915]&~m[916]&m[917])|(~m[567]&m[913]&m[915]&m[916]&m[917]))&UnbiasedRNG[241])|((m[567]&~m[913]&~m[915]&m[916]&~m[917])|(~m[567]&~m[913]&~m[915]&~m[916]&m[917])|(m[567]&~m[913]&~m[915]&~m[916]&m[917])|(m[567]&m[913]&~m[915]&~m[916]&m[917])|(m[567]&~m[913]&m[915]&~m[916]&m[917])|(~m[567]&~m[913]&~m[915]&m[916]&m[917])|(m[567]&~m[913]&~m[915]&m[916]&m[917])|(~m[567]&m[913]&~m[915]&m[916]&m[917])|(m[567]&m[913]&~m[915]&m[916]&m[917])|(~m[567]&~m[913]&m[915]&m[916]&m[917])|(m[567]&~m[913]&m[915]&m[916]&m[917])|(m[567]&m[913]&m[915]&m[916]&m[917]))):InitCond[744];
    m[919] = run?((((m[580]&~m[918]&~m[920]&~m[921]&~m[922])|(~m[580]&~m[918]&~m[920]&m[921]&~m[922])|(m[580]&m[918]&~m[920]&m[921]&~m[922])|(m[580]&~m[918]&m[920]&m[921]&~m[922])|(~m[580]&m[918]&~m[920]&~m[921]&m[922])|(~m[580]&~m[918]&m[920]&~m[921]&m[922])|(m[580]&m[918]&m[920]&~m[921]&m[922])|(~m[580]&m[918]&m[920]&m[921]&m[922]))&UnbiasedRNG[242])|((m[580]&~m[918]&~m[920]&m[921]&~m[922])|(~m[580]&~m[918]&~m[920]&~m[921]&m[922])|(m[580]&~m[918]&~m[920]&~m[921]&m[922])|(m[580]&m[918]&~m[920]&~m[921]&m[922])|(m[580]&~m[918]&m[920]&~m[921]&m[922])|(~m[580]&~m[918]&~m[920]&m[921]&m[922])|(m[580]&~m[918]&~m[920]&m[921]&m[922])|(~m[580]&m[918]&~m[920]&m[921]&m[922])|(m[580]&m[918]&~m[920]&m[921]&m[922])|(~m[580]&~m[918]&m[920]&m[921]&m[922])|(m[580]&~m[918]&m[920]&m[921]&m[922])|(m[580]&m[918]&m[920]&m[921]&m[922]))):InitCond[745];
    m[925] = run?((((m[887]&~m[923]&~m[924]&~m[926]&~m[927])|(~m[887]&~m[923]&~m[924]&m[926]&~m[927])|(m[887]&m[923]&~m[924]&m[926]&~m[927])|(m[887]&~m[923]&m[924]&m[926]&~m[927])|(~m[887]&m[923]&~m[924]&~m[926]&m[927])|(~m[887]&~m[923]&m[924]&~m[926]&m[927])|(m[887]&m[923]&m[924]&~m[926]&m[927])|(~m[887]&m[923]&m[924]&m[926]&m[927]))&UnbiasedRNG[243])|((m[887]&~m[923]&~m[924]&m[926]&~m[927])|(~m[887]&~m[923]&~m[924]&~m[926]&m[927])|(m[887]&~m[923]&~m[924]&~m[926]&m[927])|(m[887]&m[923]&~m[924]&~m[926]&m[927])|(m[887]&~m[923]&m[924]&~m[926]&m[927])|(~m[887]&~m[923]&~m[924]&m[926]&m[927])|(m[887]&~m[923]&~m[924]&m[926]&m[927])|(~m[887]&m[923]&~m[924]&m[926]&m[927])|(m[887]&m[923]&~m[924]&m[926]&m[927])|(~m[887]&~m[923]&m[924]&m[926]&m[927])|(m[887]&~m[923]&m[924]&m[926]&m[927])|(m[887]&m[923]&m[924]&m[926]&m[927]))):InitCond[746];
    m[930] = run?((((m[892]&~m[928]&~m[929]&~m[931]&~m[932])|(~m[892]&~m[928]&~m[929]&m[931]&~m[932])|(m[892]&m[928]&~m[929]&m[931]&~m[932])|(m[892]&~m[928]&m[929]&m[931]&~m[932])|(~m[892]&m[928]&~m[929]&~m[931]&m[932])|(~m[892]&~m[928]&m[929]&~m[931]&m[932])|(m[892]&m[928]&m[929]&~m[931]&m[932])|(~m[892]&m[928]&m[929]&m[931]&m[932]))&UnbiasedRNG[244])|((m[892]&~m[928]&~m[929]&m[931]&~m[932])|(~m[892]&~m[928]&~m[929]&~m[931]&m[932])|(m[892]&~m[928]&~m[929]&~m[931]&m[932])|(m[892]&m[928]&~m[929]&~m[931]&m[932])|(m[892]&~m[928]&m[929]&~m[931]&m[932])|(~m[892]&~m[928]&~m[929]&m[931]&m[932])|(m[892]&~m[928]&~m[929]&m[931]&m[932])|(~m[892]&m[928]&~m[929]&m[931]&m[932])|(m[892]&m[928]&~m[929]&m[931]&m[932])|(~m[892]&~m[928]&m[929]&m[931]&m[932])|(m[892]&~m[928]&m[929]&m[931]&m[932])|(m[892]&m[928]&m[929]&m[931]&m[932]))):InitCond[747];
    m[934] = run?((((m[619]&~m[933]&~m[935]&~m[936]&~m[937])|(~m[619]&~m[933]&~m[935]&m[936]&~m[937])|(m[619]&m[933]&~m[935]&m[936]&~m[937])|(m[619]&~m[933]&m[935]&m[936]&~m[937])|(~m[619]&m[933]&~m[935]&~m[936]&m[937])|(~m[619]&~m[933]&m[935]&~m[936]&m[937])|(m[619]&m[933]&m[935]&~m[936]&m[937])|(~m[619]&m[933]&m[935]&m[936]&m[937]))&UnbiasedRNG[245])|((m[619]&~m[933]&~m[935]&m[936]&~m[937])|(~m[619]&~m[933]&~m[935]&~m[936]&m[937])|(m[619]&~m[933]&~m[935]&~m[936]&m[937])|(m[619]&m[933]&~m[935]&~m[936]&m[937])|(m[619]&~m[933]&m[935]&~m[936]&m[937])|(~m[619]&~m[933]&~m[935]&m[936]&m[937])|(m[619]&~m[933]&~m[935]&m[936]&m[937])|(~m[619]&m[933]&~m[935]&m[936]&m[937])|(m[619]&m[933]&~m[935]&m[936]&m[937])|(~m[619]&~m[933]&m[935]&m[936]&m[937])|(m[619]&~m[933]&m[935]&m[936]&m[937])|(m[619]&m[933]&m[935]&m[936]&m[937]))):InitCond[748];
    m[939] = run?((((m[632]&~m[938]&~m[940]&~m[941]&~m[942])|(~m[632]&~m[938]&~m[940]&m[941]&~m[942])|(m[632]&m[938]&~m[940]&m[941]&~m[942])|(m[632]&~m[938]&m[940]&m[941]&~m[942])|(~m[632]&m[938]&~m[940]&~m[941]&m[942])|(~m[632]&~m[938]&m[940]&~m[941]&m[942])|(m[632]&m[938]&m[940]&~m[941]&m[942])|(~m[632]&m[938]&m[940]&m[941]&m[942]))&UnbiasedRNG[246])|((m[632]&~m[938]&~m[940]&m[941]&~m[942])|(~m[632]&~m[938]&~m[940]&~m[941]&m[942])|(m[632]&~m[938]&~m[940]&~m[941]&m[942])|(m[632]&m[938]&~m[940]&~m[941]&m[942])|(m[632]&~m[938]&m[940]&~m[941]&m[942])|(~m[632]&~m[938]&~m[940]&m[941]&m[942])|(m[632]&~m[938]&~m[940]&m[941]&m[942])|(~m[632]&m[938]&~m[940]&m[941]&m[942])|(m[632]&m[938]&~m[940]&m[941]&m[942])|(~m[632]&~m[938]&m[940]&m[941]&m[942])|(m[632]&~m[938]&m[940]&m[941]&m[942])|(m[632]&m[938]&m[940]&m[941]&m[942]))):InitCond[749];
    m[944] = run?((((m[645]&~m[943]&~m[945]&~m[946]&~m[947])|(~m[645]&~m[943]&~m[945]&m[946]&~m[947])|(m[645]&m[943]&~m[945]&m[946]&~m[947])|(m[645]&~m[943]&m[945]&m[946]&~m[947])|(~m[645]&m[943]&~m[945]&~m[946]&m[947])|(~m[645]&~m[943]&m[945]&~m[946]&m[947])|(m[645]&m[943]&m[945]&~m[946]&m[947])|(~m[645]&m[943]&m[945]&m[946]&m[947]))&UnbiasedRNG[247])|((m[645]&~m[943]&~m[945]&m[946]&~m[947])|(~m[645]&~m[943]&~m[945]&~m[946]&m[947])|(m[645]&~m[943]&~m[945]&~m[946]&m[947])|(m[645]&m[943]&~m[945]&~m[946]&m[947])|(m[645]&~m[943]&m[945]&~m[946]&m[947])|(~m[645]&~m[943]&~m[945]&m[946]&m[947])|(m[645]&~m[943]&~m[945]&m[946]&m[947])|(~m[645]&m[943]&~m[945]&m[946]&m[947])|(m[645]&m[943]&~m[945]&m[946]&m[947])|(~m[645]&~m[943]&m[945]&m[946]&m[947])|(m[645]&~m[943]&m[945]&m[946]&m[947])|(m[645]&m[943]&m[945]&m[946]&m[947]))):InitCond[750];
    m[949] = run?((((m[658]&~m[948]&~m[950]&~m[951]&~m[952])|(~m[658]&~m[948]&~m[950]&m[951]&~m[952])|(m[658]&m[948]&~m[950]&m[951]&~m[952])|(m[658]&~m[948]&m[950]&m[951]&~m[952])|(~m[658]&m[948]&~m[950]&~m[951]&m[952])|(~m[658]&~m[948]&m[950]&~m[951]&m[952])|(m[658]&m[948]&m[950]&~m[951]&m[952])|(~m[658]&m[948]&m[950]&m[951]&m[952]))&UnbiasedRNG[248])|((m[658]&~m[948]&~m[950]&m[951]&~m[952])|(~m[658]&~m[948]&~m[950]&~m[951]&m[952])|(m[658]&~m[948]&~m[950]&~m[951]&m[952])|(m[658]&m[948]&~m[950]&~m[951]&m[952])|(m[658]&~m[948]&m[950]&~m[951]&m[952])|(~m[658]&~m[948]&~m[950]&m[951]&m[952])|(m[658]&~m[948]&~m[950]&m[951]&m[952])|(~m[658]&m[948]&~m[950]&m[951]&m[952])|(m[658]&m[948]&~m[950]&m[951]&m[952])|(~m[658]&~m[948]&m[950]&m[951]&m[952])|(m[658]&~m[948]&m[950]&m[951]&m[952])|(m[658]&m[948]&m[950]&m[951]&m[952]))):InitCond[751];
    m[954] = run?((((m[555]&~m[953]&~m[955]&~m[956]&~m[957])|(~m[555]&~m[953]&~m[955]&m[956]&~m[957])|(m[555]&m[953]&~m[955]&m[956]&~m[957])|(m[555]&~m[953]&m[955]&m[956]&~m[957])|(~m[555]&m[953]&~m[955]&~m[956]&m[957])|(~m[555]&~m[953]&m[955]&~m[956]&m[957])|(m[555]&m[953]&m[955]&~m[956]&m[957])|(~m[555]&m[953]&m[955]&m[956]&m[957]))&UnbiasedRNG[249])|((m[555]&~m[953]&~m[955]&m[956]&~m[957])|(~m[555]&~m[953]&~m[955]&~m[956]&m[957])|(m[555]&~m[953]&~m[955]&~m[956]&m[957])|(m[555]&m[953]&~m[955]&~m[956]&m[957])|(m[555]&~m[953]&m[955]&~m[956]&m[957])|(~m[555]&~m[953]&~m[955]&m[956]&m[957])|(m[555]&~m[953]&~m[955]&m[956]&m[957])|(~m[555]&m[953]&~m[955]&m[956]&m[957])|(m[555]&m[953]&~m[955]&m[956]&m[957])|(~m[555]&~m[953]&m[955]&m[956]&m[957])|(m[555]&~m[953]&m[955]&m[956]&m[957])|(m[555]&m[953]&m[955]&m[956]&m[957]))):InitCond[752];
    m[959] = run?((((m[568]&~m[958]&~m[960]&~m[961]&~m[962])|(~m[568]&~m[958]&~m[960]&m[961]&~m[962])|(m[568]&m[958]&~m[960]&m[961]&~m[962])|(m[568]&~m[958]&m[960]&m[961]&~m[962])|(~m[568]&m[958]&~m[960]&~m[961]&m[962])|(~m[568]&~m[958]&m[960]&~m[961]&m[962])|(m[568]&m[958]&m[960]&~m[961]&m[962])|(~m[568]&m[958]&m[960]&m[961]&m[962]))&UnbiasedRNG[250])|((m[568]&~m[958]&~m[960]&m[961]&~m[962])|(~m[568]&~m[958]&~m[960]&~m[961]&m[962])|(m[568]&~m[958]&~m[960]&~m[961]&m[962])|(m[568]&m[958]&~m[960]&~m[961]&m[962])|(m[568]&~m[958]&m[960]&~m[961]&m[962])|(~m[568]&~m[958]&~m[960]&m[961]&m[962])|(m[568]&~m[958]&~m[960]&m[961]&m[962])|(~m[568]&m[958]&~m[960]&m[961]&m[962])|(m[568]&m[958]&~m[960]&m[961]&m[962])|(~m[568]&~m[958]&m[960]&m[961]&m[962])|(m[568]&~m[958]&m[960]&m[961]&m[962])|(m[568]&m[958]&m[960]&m[961]&m[962]))):InitCond[753];
    m[964] = run?((((m[581]&~m[963]&~m[965]&~m[966]&~m[967])|(~m[581]&~m[963]&~m[965]&m[966]&~m[967])|(m[581]&m[963]&~m[965]&m[966]&~m[967])|(m[581]&~m[963]&m[965]&m[966]&~m[967])|(~m[581]&m[963]&~m[965]&~m[966]&m[967])|(~m[581]&~m[963]&m[965]&~m[966]&m[967])|(m[581]&m[963]&m[965]&~m[966]&m[967])|(~m[581]&m[963]&m[965]&m[966]&m[967]))&UnbiasedRNG[251])|((m[581]&~m[963]&~m[965]&m[966]&~m[967])|(~m[581]&~m[963]&~m[965]&~m[966]&m[967])|(m[581]&~m[963]&~m[965]&~m[966]&m[967])|(m[581]&m[963]&~m[965]&~m[966]&m[967])|(m[581]&~m[963]&m[965]&~m[966]&m[967])|(~m[581]&~m[963]&~m[965]&m[966]&m[967])|(m[581]&~m[963]&~m[965]&m[966]&m[967])|(~m[581]&m[963]&~m[965]&m[966]&m[967])|(m[581]&m[963]&~m[965]&m[966]&m[967])|(~m[581]&~m[963]&m[965]&m[966]&m[967])|(m[581]&~m[963]&m[965]&m[966]&m[967])|(m[581]&m[963]&m[965]&m[966]&m[967]))):InitCond[754];
    m[969] = run?((((m[594]&~m[968]&~m[970]&~m[971]&~m[972])|(~m[594]&~m[968]&~m[970]&m[971]&~m[972])|(m[594]&m[968]&~m[970]&m[971]&~m[972])|(m[594]&~m[968]&m[970]&m[971]&~m[972])|(~m[594]&m[968]&~m[970]&~m[971]&m[972])|(~m[594]&~m[968]&m[970]&~m[971]&m[972])|(m[594]&m[968]&m[970]&~m[971]&m[972])|(~m[594]&m[968]&m[970]&m[971]&m[972]))&UnbiasedRNG[252])|((m[594]&~m[968]&~m[970]&m[971]&~m[972])|(~m[594]&~m[968]&~m[970]&~m[971]&m[972])|(m[594]&~m[968]&~m[970]&~m[971]&m[972])|(m[594]&m[968]&~m[970]&~m[971]&m[972])|(m[594]&~m[968]&m[970]&~m[971]&m[972])|(~m[594]&~m[968]&~m[970]&m[971]&m[972])|(m[594]&~m[968]&~m[970]&m[971]&m[972])|(~m[594]&m[968]&~m[970]&m[971]&m[972])|(m[594]&m[968]&~m[970]&m[971]&m[972])|(~m[594]&~m[968]&m[970]&m[971]&m[972])|(m[594]&~m[968]&m[970]&m[971]&m[972])|(m[594]&m[968]&m[970]&m[971]&m[972]))):InitCond[755];
    m[975] = run?((((m[932]&~m[973]&~m[974]&~m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&m[976]&~m[977])|(m[932]&m[973]&~m[974]&m[976]&~m[977])|(m[932]&~m[973]&m[974]&m[976]&~m[977])|(~m[932]&m[973]&~m[974]&~m[976]&m[977])|(~m[932]&~m[973]&m[974]&~m[976]&m[977])|(m[932]&m[973]&m[974]&~m[976]&m[977])|(~m[932]&m[973]&m[974]&m[976]&m[977]))&UnbiasedRNG[253])|((m[932]&~m[973]&~m[974]&m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&m[974]&~m[976]&m[977])|(~m[932]&~m[973]&~m[974]&m[976]&m[977])|(m[932]&~m[973]&~m[974]&m[976]&m[977])|(~m[932]&m[973]&~m[974]&m[976]&m[977])|(m[932]&m[973]&~m[974]&m[976]&m[977])|(~m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&m[973]&m[974]&m[976]&m[977]))):InitCond[756];
    m[979] = run?((((m[620]&~m[978]&~m[980]&~m[981]&~m[982])|(~m[620]&~m[978]&~m[980]&m[981]&~m[982])|(m[620]&m[978]&~m[980]&m[981]&~m[982])|(m[620]&~m[978]&m[980]&m[981]&~m[982])|(~m[620]&m[978]&~m[980]&~m[981]&m[982])|(~m[620]&~m[978]&m[980]&~m[981]&m[982])|(m[620]&m[978]&m[980]&~m[981]&m[982])|(~m[620]&m[978]&m[980]&m[981]&m[982]))&UnbiasedRNG[254])|((m[620]&~m[978]&~m[980]&m[981]&~m[982])|(~m[620]&~m[978]&~m[980]&~m[981]&m[982])|(m[620]&~m[978]&~m[980]&~m[981]&m[982])|(m[620]&m[978]&~m[980]&~m[981]&m[982])|(m[620]&~m[978]&m[980]&~m[981]&m[982])|(~m[620]&~m[978]&~m[980]&m[981]&m[982])|(m[620]&~m[978]&~m[980]&m[981]&m[982])|(~m[620]&m[978]&~m[980]&m[981]&m[982])|(m[620]&m[978]&~m[980]&m[981]&m[982])|(~m[620]&~m[978]&m[980]&m[981]&m[982])|(m[620]&~m[978]&m[980]&m[981]&m[982])|(m[620]&m[978]&m[980]&m[981]&m[982]))):InitCond[757];
    m[984] = run?((((m[633]&~m[983]&~m[985]&~m[986]&~m[987])|(~m[633]&~m[983]&~m[985]&m[986]&~m[987])|(m[633]&m[983]&~m[985]&m[986]&~m[987])|(m[633]&~m[983]&m[985]&m[986]&~m[987])|(~m[633]&m[983]&~m[985]&~m[986]&m[987])|(~m[633]&~m[983]&m[985]&~m[986]&m[987])|(m[633]&m[983]&m[985]&~m[986]&m[987])|(~m[633]&m[983]&m[985]&m[986]&m[987]))&UnbiasedRNG[255])|((m[633]&~m[983]&~m[985]&m[986]&~m[987])|(~m[633]&~m[983]&~m[985]&~m[986]&m[987])|(m[633]&~m[983]&~m[985]&~m[986]&m[987])|(m[633]&m[983]&~m[985]&~m[986]&m[987])|(m[633]&~m[983]&m[985]&~m[986]&m[987])|(~m[633]&~m[983]&~m[985]&m[986]&m[987])|(m[633]&~m[983]&~m[985]&m[986]&m[987])|(~m[633]&m[983]&~m[985]&m[986]&m[987])|(m[633]&m[983]&~m[985]&m[986]&m[987])|(~m[633]&~m[983]&m[985]&m[986]&m[987])|(m[633]&~m[983]&m[985]&m[986]&m[987])|(m[633]&m[983]&m[985]&m[986]&m[987]))):InitCond[758];
    m[989] = run?((((m[646]&~m[988]&~m[990]&~m[991]&~m[992])|(~m[646]&~m[988]&~m[990]&m[991]&~m[992])|(m[646]&m[988]&~m[990]&m[991]&~m[992])|(m[646]&~m[988]&m[990]&m[991]&~m[992])|(~m[646]&m[988]&~m[990]&~m[991]&m[992])|(~m[646]&~m[988]&m[990]&~m[991]&m[992])|(m[646]&m[988]&m[990]&~m[991]&m[992])|(~m[646]&m[988]&m[990]&m[991]&m[992]))&UnbiasedRNG[256])|((m[646]&~m[988]&~m[990]&m[991]&~m[992])|(~m[646]&~m[988]&~m[990]&~m[991]&m[992])|(m[646]&~m[988]&~m[990]&~m[991]&m[992])|(m[646]&m[988]&~m[990]&~m[991]&m[992])|(m[646]&~m[988]&m[990]&~m[991]&m[992])|(~m[646]&~m[988]&~m[990]&m[991]&m[992])|(m[646]&~m[988]&~m[990]&m[991]&m[992])|(~m[646]&m[988]&~m[990]&m[991]&m[992])|(m[646]&m[988]&~m[990]&m[991]&m[992])|(~m[646]&~m[988]&m[990]&m[991]&m[992])|(m[646]&~m[988]&m[990]&m[991]&m[992])|(m[646]&m[988]&m[990]&m[991]&m[992]))):InitCond[759];
    m[994] = run?((((m[659]&~m[993]&~m[995]&~m[996]&~m[997])|(~m[659]&~m[993]&~m[995]&m[996]&~m[997])|(m[659]&m[993]&~m[995]&m[996]&~m[997])|(m[659]&~m[993]&m[995]&m[996]&~m[997])|(~m[659]&m[993]&~m[995]&~m[996]&m[997])|(~m[659]&~m[993]&m[995]&~m[996]&m[997])|(m[659]&m[993]&m[995]&~m[996]&m[997])|(~m[659]&m[993]&m[995]&m[996]&m[997]))&UnbiasedRNG[257])|((m[659]&~m[993]&~m[995]&m[996]&~m[997])|(~m[659]&~m[993]&~m[995]&~m[996]&m[997])|(m[659]&~m[993]&~m[995]&~m[996]&m[997])|(m[659]&m[993]&~m[995]&~m[996]&m[997])|(m[659]&~m[993]&m[995]&~m[996]&m[997])|(~m[659]&~m[993]&~m[995]&m[996]&m[997])|(m[659]&~m[993]&~m[995]&m[996]&m[997])|(~m[659]&m[993]&~m[995]&m[996]&m[997])|(m[659]&m[993]&~m[995]&m[996]&m[997])|(~m[659]&~m[993]&m[995]&m[996]&m[997])|(m[659]&~m[993]&m[995]&m[996]&m[997])|(m[659]&m[993]&m[995]&m[996]&m[997]))):InitCond[760];
    m[999] = run?((((m[672]&~m[998]&~m[1000]&~m[1001]&~m[1002])|(~m[672]&~m[998]&~m[1000]&m[1001]&~m[1002])|(m[672]&m[998]&~m[1000]&m[1001]&~m[1002])|(m[672]&~m[998]&m[1000]&m[1001]&~m[1002])|(~m[672]&m[998]&~m[1000]&~m[1001]&m[1002])|(~m[672]&~m[998]&m[1000]&~m[1001]&m[1002])|(m[672]&m[998]&m[1000]&~m[1001]&m[1002])|(~m[672]&m[998]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[258])|((m[672]&~m[998]&~m[1000]&m[1001]&~m[1002])|(~m[672]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[672]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[672]&m[998]&~m[1000]&~m[1001]&m[1002])|(m[672]&~m[998]&m[1000]&~m[1001]&m[1002])|(~m[672]&~m[998]&~m[1000]&m[1001]&m[1002])|(m[672]&~m[998]&~m[1000]&m[1001]&m[1002])|(~m[672]&m[998]&~m[1000]&m[1001]&m[1002])|(m[672]&m[998]&~m[1000]&m[1001]&m[1002])|(~m[672]&~m[998]&m[1000]&m[1001]&m[1002])|(m[672]&~m[998]&m[1000]&m[1001]&m[1002])|(m[672]&m[998]&m[1000]&m[1001]&m[1002]))):InitCond[761];
    m[1004] = run?((((m[556]&~m[1003]&~m[1005]&~m[1006]&~m[1007])|(~m[556]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(m[556]&m[1003]&~m[1005]&m[1006]&~m[1007])|(m[556]&~m[1003]&m[1005]&m[1006]&~m[1007])|(~m[556]&m[1003]&~m[1005]&~m[1006]&m[1007])|(~m[556]&~m[1003]&m[1005]&~m[1006]&m[1007])|(m[556]&m[1003]&m[1005]&~m[1006]&m[1007])|(~m[556]&m[1003]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[259])|((m[556]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(~m[556]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[556]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[556]&m[1003]&~m[1005]&~m[1006]&m[1007])|(m[556]&~m[1003]&m[1005]&~m[1006]&m[1007])|(~m[556]&~m[1003]&~m[1005]&m[1006]&m[1007])|(m[556]&~m[1003]&~m[1005]&m[1006]&m[1007])|(~m[556]&m[1003]&~m[1005]&m[1006]&m[1007])|(m[556]&m[1003]&~m[1005]&m[1006]&m[1007])|(~m[556]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[556]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[556]&m[1003]&m[1005]&m[1006]&m[1007]))):InitCond[762];
    m[1009] = run?((((m[569]&~m[1008]&~m[1010]&~m[1011]&~m[1012])|(~m[569]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(m[569]&m[1008]&~m[1010]&m[1011]&~m[1012])|(m[569]&~m[1008]&m[1010]&m[1011]&~m[1012])|(~m[569]&m[1008]&~m[1010]&~m[1011]&m[1012])|(~m[569]&~m[1008]&m[1010]&~m[1011]&m[1012])|(m[569]&m[1008]&m[1010]&~m[1011]&m[1012])|(~m[569]&m[1008]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[260])|((m[569]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(~m[569]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[569]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[569]&m[1008]&~m[1010]&~m[1011]&m[1012])|(m[569]&~m[1008]&m[1010]&~m[1011]&m[1012])|(~m[569]&~m[1008]&~m[1010]&m[1011]&m[1012])|(m[569]&~m[1008]&~m[1010]&m[1011]&m[1012])|(~m[569]&m[1008]&~m[1010]&m[1011]&m[1012])|(m[569]&m[1008]&~m[1010]&m[1011]&m[1012])|(~m[569]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[569]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[569]&m[1008]&m[1010]&m[1011]&m[1012]))):InitCond[763];
    m[1014] = run?((((m[582]&~m[1013]&~m[1015]&~m[1016]&~m[1017])|(~m[582]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(m[582]&m[1013]&~m[1015]&m[1016]&~m[1017])|(m[582]&~m[1013]&m[1015]&m[1016]&~m[1017])|(~m[582]&m[1013]&~m[1015]&~m[1016]&m[1017])|(~m[582]&~m[1013]&m[1015]&~m[1016]&m[1017])|(m[582]&m[1013]&m[1015]&~m[1016]&m[1017])|(~m[582]&m[1013]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[261])|((m[582]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(~m[582]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[582]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[582]&m[1013]&~m[1015]&~m[1016]&m[1017])|(m[582]&~m[1013]&m[1015]&~m[1016]&m[1017])|(~m[582]&~m[1013]&~m[1015]&m[1016]&m[1017])|(m[582]&~m[1013]&~m[1015]&m[1016]&m[1017])|(~m[582]&m[1013]&~m[1015]&m[1016]&m[1017])|(m[582]&m[1013]&~m[1015]&m[1016]&m[1017])|(~m[582]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[582]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[582]&m[1013]&m[1015]&m[1016]&m[1017]))):InitCond[764];
    m[1019] = run?((((m[595]&~m[1018]&~m[1020]&~m[1021]&~m[1022])|(~m[595]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(m[595]&m[1018]&~m[1020]&m[1021]&~m[1022])|(m[595]&~m[1018]&m[1020]&m[1021]&~m[1022])|(~m[595]&m[1018]&~m[1020]&~m[1021]&m[1022])|(~m[595]&~m[1018]&m[1020]&~m[1021]&m[1022])|(m[595]&m[1018]&m[1020]&~m[1021]&m[1022])|(~m[595]&m[1018]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[262])|((m[595]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(~m[595]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[595]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[595]&m[1018]&~m[1020]&~m[1021]&m[1022])|(m[595]&~m[1018]&m[1020]&~m[1021]&m[1022])|(~m[595]&~m[1018]&~m[1020]&m[1021]&m[1022])|(m[595]&~m[1018]&~m[1020]&m[1021]&m[1022])|(~m[595]&m[1018]&~m[1020]&m[1021]&m[1022])|(m[595]&m[1018]&~m[1020]&m[1021]&m[1022])|(~m[595]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[595]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[595]&m[1018]&m[1020]&m[1021]&m[1022]))):InitCond[765];
    m[1024] = run?((((m[608]&~m[1023]&~m[1025]&~m[1026]&~m[1027])|(~m[608]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(m[608]&m[1023]&~m[1025]&m[1026]&~m[1027])|(m[608]&~m[1023]&m[1025]&m[1026]&~m[1027])|(~m[608]&m[1023]&~m[1025]&~m[1026]&m[1027])|(~m[608]&~m[1023]&m[1025]&~m[1026]&m[1027])|(m[608]&m[1023]&m[1025]&~m[1026]&m[1027])|(~m[608]&m[1023]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[263])|((m[608]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(~m[608]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[608]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[608]&m[1023]&~m[1025]&~m[1026]&m[1027])|(m[608]&~m[1023]&m[1025]&~m[1026]&m[1027])|(~m[608]&~m[1023]&~m[1025]&m[1026]&m[1027])|(m[608]&~m[1023]&~m[1025]&m[1026]&m[1027])|(~m[608]&m[1023]&~m[1025]&m[1026]&m[1027])|(m[608]&m[1023]&~m[1025]&m[1026]&m[1027])|(~m[608]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[608]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[608]&m[1023]&m[1025]&m[1026]&m[1027]))):InitCond[766];
    m[1029] = run?((((m[621]&~m[1028]&~m[1030]&~m[1031]&~m[1032])|(~m[621]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(m[621]&m[1028]&~m[1030]&m[1031]&~m[1032])|(m[621]&~m[1028]&m[1030]&m[1031]&~m[1032])|(~m[621]&m[1028]&~m[1030]&~m[1031]&m[1032])|(~m[621]&~m[1028]&m[1030]&~m[1031]&m[1032])|(m[621]&m[1028]&m[1030]&~m[1031]&m[1032])|(~m[621]&m[1028]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[264])|((m[621]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(~m[621]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[621]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[621]&m[1028]&~m[1030]&~m[1031]&m[1032])|(m[621]&~m[1028]&m[1030]&~m[1031]&m[1032])|(~m[621]&~m[1028]&~m[1030]&m[1031]&m[1032])|(m[621]&~m[1028]&~m[1030]&m[1031]&m[1032])|(~m[621]&m[1028]&~m[1030]&m[1031]&m[1032])|(m[621]&m[1028]&~m[1030]&m[1031]&m[1032])|(~m[621]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[621]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[621]&m[1028]&m[1030]&m[1031]&m[1032]))):InitCond[767];
    m[1034] = run?((((m[634]&~m[1033]&~m[1035]&~m[1036]&~m[1037])|(~m[634]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(m[634]&m[1033]&~m[1035]&m[1036]&~m[1037])|(m[634]&~m[1033]&m[1035]&m[1036]&~m[1037])|(~m[634]&m[1033]&~m[1035]&~m[1036]&m[1037])|(~m[634]&~m[1033]&m[1035]&~m[1036]&m[1037])|(m[634]&m[1033]&m[1035]&~m[1036]&m[1037])|(~m[634]&m[1033]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[265])|((m[634]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(~m[634]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[634]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[634]&m[1033]&~m[1035]&~m[1036]&m[1037])|(m[634]&~m[1033]&m[1035]&~m[1036]&m[1037])|(~m[634]&~m[1033]&~m[1035]&m[1036]&m[1037])|(m[634]&~m[1033]&~m[1035]&m[1036]&m[1037])|(~m[634]&m[1033]&~m[1035]&m[1036]&m[1037])|(m[634]&m[1033]&~m[1035]&m[1036]&m[1037])|(~m[634]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[634]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[634]&m[1033]&m[1035]&m[1036]&m[1037]))):InitCond[768];
    m[1039] = run?((((m[647]&~m[1038]&~m[1040]&~m[1041]&~m[1042])|(~m[647]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(m[647]&m[1038]&~m[1040]&m[1041]&~m[1042])|(m[647]&~m[1038]&m[1040]&m[1041]&~m[1042])|(~m[647]&m[1038]&~m[1040]&~m[1041]&m[1042])|(~m[647]&~m[1038]&m[1040]&~m[1041]&m[1042])|(m[647]&m[1038]&m[1040]&~m[1041]&m[1042])|(~m[647]&m[1038]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[266])|((m[647]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(~m[647]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[647]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[647]&m[1038]&~m[1040]&~m[1041]&m[1042])|(m[647]&~m[1038]&m[1040]&~m[1041]&m[1042])|(~m[647]&~m[1038]&~m[1040]&m[1041]&m[1042])|(m[647]&~m[1038]&~m[1040]&m[1041]&m[1042])|(~m[647]&m[1038]&~m[1040]&m[1041]&m[1042])|(m[647]&m[1038]&~m[1040]&m[1041]&m[1042])|(~m[647]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[647]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[647]&m[1038]&m[1040]&m[1041]&m[1042]))):InitCond[769];
    m[1044] = run?((((m[660]&~m[1043]&~m[1045]&~m[1046]&~m[1047])|(~m[660]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(m[660]&m[1043]&~m[1045]&m[1046]&~m[1047])|(m[660]&~m[1043]&m[1045]&m[1046]&~m[1047])|(~m[660]&m[1043]&~m[1045]&~m[1046]&m[1047])|(~m[660]&~m[1043]&m[1045]&~m[1046]&m[1047])|(m[660]&m[1043]&m[1045]&~m[1046]&m[1047])|(~m[660]&m[1043]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[267])|((m[660]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(~m[660]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[660]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[660]&m[1043]&~m[1045]&~m[1046]&m[1047])|(m[660]&~m[1043]&m[1045]&~m[1046]&m[1047])|(~m[660]&~m[1043]&~m[1045]&m[1046]&m[1047])|(m[660]&~m[1043]&~m[1045]&m[1046]&m[1047])|(~m[660]&m[1043]&~m[1045]&m[1046]&m[1047])|(m[660]&m[1043]&~m[1045]&m[1046]&m[1047])|(~m[660]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[660]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[660]&m[1043]&m[1045]&m[1046]&m[1047]))):InitCond[770];
    m[1049] = run?((((m[673]&~m[1048]&~m[1050]&~m[1051]&~m[1052])|(~m[673]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(m[673]&m[1048]&~m[1050]&m[1051]&~m[1052])|(m[673]&~m[1048]&m[1050]&m[1051]&~m[1052])|(~m[673]&m[1048]&~m[1050]&~m[1051]&m[1052])|(~m[673]&~m[1048]&m[1050]&~m[1051]&m[1052])|(m[673]&m[1048]&m[1050]&~m[1051]&m[1052])|(~m[673]&m[1048]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[268])|((m[673]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(~m[673]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[673]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[673]&m[1048]&~m[1050]&~m[1051]&m[1052])|(m[673]&~m[1048]&m[1050]&~m[1051]&m[1052])|(~m[673]&~m[1048]&~m[1050]&m[1051]&m[1052])|(m[673]&~m[1048]&~m[1050]&m[1051]&m[1052])|(~m[673]&m[1048]&~m[1050]&m[1051]&m[1052])|(m[673]&m[1048]&~m[1050]&m[1051]&m[1052])|(~m[673]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[673]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[673]&m[1048]&m[1050]&m[1051]&m[1052]))):InitCond[771];
    m[1054] = run?((((m[686]&~m[1053]&~m[1055]&~m[1056]&~m[1057])|(~m[686]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(m[686]&m[1053]&~m[1055]&m[1056]&~m[1057])|(m[686]&~m[1053]&m[1055]&m[1056]&~m[1057])|(~m[686]&m[1053]&~m[1055]&~m[1056]&m[1057])|(~m[686]&~m[1053]&m[1055]&~m[1056]&m[1057])|(m[686]&m[1053]&m[1055]&~m[1056]&m[1057])|(~m[686]&m[1053]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[269])|((m[686]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(~m[686]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[686]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[686]&m[1053]&~m[1055]&~m[1056]&m[1057])|(m[686]&~m[1053]&m[1055]&~m[1056]&m[1057])|(~m[686]&~m[1053]&~m[1055]&m[1056]&m[1057])|(m[686]&~m[1053]&~m[1055]&m[1056]&m[1057])|(~m[686]&m[1053]&~m[1055]&m[1056]&m[1057])|(m[686]&m[1053]&~m[1055]&m[1056]&m[1057])|(~m[686]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[686]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[686]&m[1053]&m[1055]&m[1056]&m[1057]))):InitCond[772];
    m[1059] = run?((((m[557]&~m[1058]&~m[1060]&~m[1061]&~m[1062])|(~m[557]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(m[557]&m[1058]&~m[1060]&m[1061]&~m[1062])|(m[557]&~m[1058]&m[1060]&m[1061]&~m[1062])|(~m[557]&m[1058]&~m[1060]&~m[1061]&m[1062])|(~m[557]&~m[1058]&m[1060]&~m[1061]&m[1062])|(m[557]&m[1058]&m[1060]&~m[1061]&m[1062])|(~m[557]&m[1058]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[270])|((m[557]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(~m[557]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[557]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[557]&m[1058]&~m[1060]&~m[1061]&m[1062])|(m[557]&~m[1058]&m[1060]&~m[1061]&m[1062])|(~m[557]&~m[1058]&~m[1060]&m[1061]&m[1062])|(m[557]&~m[1058]&~m[1060]&m[1061]&m[1062])|(~m[557]&m[1058]&~m[1060]&m[1061]&m[1062])|(m[557]&m[1058]&~m[1060]&m[1061]&m[1062])|(~m[557]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[557]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[557]&m[1058]&m[1060]&m[1061]&m[1062]))):InitCond[773];
    m[1064] = run?((((m[570]&~m[1063]&~m[1065]&~m[1066]&~m[1067])|(~m[570]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(m[570]&m[1063]&~m[1065]&m[1066]&~m[1067])|(m[570]&~m[1063]&m[1065]&m[1066]&~m[1067])|(~m[570]&m[1063]&~m[1065]&~m[1066]&m[1067])|(~m[570]&~m[1063]&m[1065]&~m[1066]&m[1067])|(m[570]&m[1063]&m[1065]&~m[1066]&m[1067])|(~m[570]&m[1063]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[271])|((m[570]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(~m[570]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[570]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[570]&m[1063]&~m[1065]&~m[1066]&m[1067])|(m[570]&~m[1063]&m[1065]&~m[1066]&m[1067])|(~m[570]&~m[1063]&~m[1065]&m[1066]&m[1067])|(m[570]&~m[1063]&~m[1065]&m[1066]&m[1067])|(~m[570]&m[1063]&~m[1065]&m[1066]&m[1067])|(m[570]&m[1063]&~m[1065]&m[1066]&m[1067])|(~m[570]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[570]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[570]&m[1063]&m[1065]&m[1066]&m[1067]))):InitCond[774];
    m[1069] = run?((((m[583]&~m[1068]&~m[1070]&~m[1071]&~m[1072])|(~m[583]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(m[583]&m[1068]&~m[1070]&m[1071]&~m[1072])|(m[583]&~m[1068]&m[1070]&m[1071]&~m[1072])|(~m[583]&m[1068]&~m[1070]&~m[1071]&m[1072])|(~m[583]&~m[1068]&m[1070]&~m[1071]&m[1072])|(m[583]&m[1068]&m[1070]&~m[1071]&m[1072])|(~m[583]&m[1068]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[272])|((m[583]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(~m[583]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[583]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[583]&m[1068]&~m[1070]&~m[1071]&m[1072])|(m[583]&~m[1068]&m[1070]&~m[1071]&m[1072])|(~m[583]&~m[1068]&~m[1070]&m[1071]&m[1072])|(m[583]&~m[1068]&~m[1070]&m[1071]&m[1072])|(~m[583]&m[1068]&~m[1070]&m[1071]&m[1072])|(m[583]&m[1068]&~m[1070]&m[1071]&m[1072])|(~m[583]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[583]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[583]&m[1068]&m[1070]&m[1071]&m[1072]))):InitCond[775];
    m[1074] = run?((((m[596]&~m[1073]&~m[1075]&~m[1076]&~m[1077])|(~m[596]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(m[596]&m[1073]&~m[1075]&m[1076]&~m[1077])|(m[596]&~m[1073]&m[1075]&m[1076]&~m[1077])|(~m[596]&m[1073]&~m[1075]&~m[1076]&m[1077])|(~m[596]&~m[1073]&m[1075]&~m[1076]&m[1077])|(m[596]&m[1073]&m[1075]&~m[1076]&m[1077])|(~m[596]&m[1073]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[273])|((m[596]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(~m[596]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[596]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[596]&m[1073]&~m[1075]&~m[1076]&m[1077])|(m[596]&~m[1073]&m[1075]&~m[1076]&m[1077])|(~m[596]&~m[1073]&~m[1075]&m[1076]&m[1077])|(m[596]&~m[1073]&~m[1075]&m[1076]&m[1077])|(~m[596]&m[1073]&~m[1075]&m[1076]&m[1077])|(m[596]&m[1073]&~m[1075]&m[1076]&m[1077])|(~m[596]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[596]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[596]&m[1073]&m[1075]&m[1076]&m[1077]))):InitCond[776];
    m[1079] = run?((((m[609]&~m[1078]&~m[1080]&~m[1081]&~m[1082])|(~m[609]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(m[609]&m[1078]&~m[1080]&m[1081]&~m[1082])|(m[609]&~m[1078]&m[1080]&m[1081]&~m[1082])|(~m[609]&m[1078]&~m[1080]&~m[1081]&m[1082])|(~m[609]&~m[1078]&m[1080]&~m[1081]&m[1082])|(m[609]&m[1078]&m[1080]&~m[1081]&m[1082])|(~m[609]&m[1078]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[274])|((m[609]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(~m[609]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[609]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[609]&m[1078]&~m[1080]&~m[1081]&m[1082])|(m[609]&~m[1078]&m[1080]&~m[1081]&m[1082])|(~m[609]&~m[1078]&~m[1080]&m[1081]&m[1082])|(m[609]&~m[1078]&~m[1080]&m[1081]&m[1082])|(~m[609]&m[1078]&~m[1080]&m[1081]&m[1082])|(m[609]&m[1078]&~m[1080]&m[1081]&m[1082])|(~m[609]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[609]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[609]&m[1078]&m[1080]&m[1081]&m[1082]))):InitCond[777];
    m[1084] = run?((((m[622]&~m[1083]&~m[1085]&~m[1086]&~m[1087])|(~m[622]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(m[622]&m[1083]&~m[1085]&m[1086]&~m[1087])|(m[622]&~m[1083]&m[1085]&m[1086]&~m[1087])|(~m[622]&m[1083]&~m[1085]&~m[1086]&m[1087])|(~m[622]&~m[1083]&m[1085]&~m[1086]&m[1087])|(m[622]&m[1083]&m[1085]&~m[1086]&m[1087])|(~m[622]&m[1083]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[275])|((m[622]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(~m[622]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[622]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[622]&m[1083]&~m[1085]&~m[1086]&m[1087])|(m[622]&~m[1083]&m[1085]&~m[1086]&m[1087])|(~m[622]&~m[1083]&~m[1085]&m[1086]&m[1087])|(m[622]&~m[1083]&~m[1085]&m[1086]&m[1087])|(~m[622]&m[1083]&~m[1085]&m[1086]&m[1087])|(m[622]&m[1083]&~m[1085]&m[1086]&m[1087])|(~m[622]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[622]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[622]&m[1083]&m[1085]&m[1086]&m[1087]))):InitCond[778];
    m[1089] = run?((((m[635]&~m[1088]&~m[1090]&~m[1091]&~m[1092])|(~m[635]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(m[635]&m[1088]&~m[1090]&m[1091]&~m[1092])|(m[635]&~m[1088]&m[1090]&m[1091]&~m[1092])|(~m[635]&m[1088]&~m[1090]&~m[1091]&m[1092])|(~m[635]&~m[1088]&m[1090]&~m[1091]&m[1092])|(m[635]&m[1088]&m[1090]&~m[1091]&m[1092])|(~m[635]&m[1088]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[276])|((m[635]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(~m[635]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[635]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[635]&m[1088]&~m[1090]&~m[1091]&m[1092])|(m[635]&~m[1088]&m[1090]&~m[1091]&m[1092])|(~m[635]&~m[1088]&~m[1090]&m[1091]&m[1092])|(m[635]&~m[1088]&~m[1090]&m[1091]&m[1092])|(~m[635]&m[1088]&~m[1090]&m[1091]&m[1092])|(m[635]&m[1088]&~m[1090]&m[1091]&m[1092])|(~m[635]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[635]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[635]&m[1088]&m[1090]&m[1091]&m[1092]))):InitCond[779];
    m[1094] = run?((((m[648]&~m[1093]&~m[1095]&~m[1096]&~m[1097])|(~m[648]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(m[648]&m[1093]&~m[1095]&m[1096]&~m[1097])|(m[648]&~m[1093]&m[1095]&m[1096]&~m[1097])|(~m[648]&m[1093]&~m[1095]&~m[1096]&m[1097])|(~m[648]&~m[1093]&m[1095]&~m[1096]&m[1097])|(m[648]&m[1093]&m[1095]&~m[1096]&m[1097])|(~m[648]&m[1093]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[277])|((m[648]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(~m[648]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[648]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[648]&m[1093]&~m[1095]&~m[1096]&m[1097])|(m[648]&~m[1093]&m[1095]&~m[1096]&m[1097])|(~m[648]&~m[1093]&~m[1095]&m[1096]&m[1097])|(m[648]&~m[1093]&~m[1095]&m[1096]&m[1097])|(~m[648]&m[1093]&~m[1095]&m[1096]&m[1097])|(m[648]&m[1093]&~m[1095]&m[1096]&m[1097])|(~m[648]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[648]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[648]&m[1093]&m[1095]&m[1096]&m[1097]))):InitCond[780];
    m[1099] = run?((((m[661]&~m[1098]&~m[1100]&~m[1101]&~m[1102])|(~m[661]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(m[661]&m[1098]&~m[1100]&m[1101]&~m[1102])|(m[661]&~m[1098]&m[1100]&m[1101]&~m[1102])|(~m[661]&m[1098]&~m[1100]&~m[1101]&m[1102])|(~m[661]&~m[1098]&m[1100]&~m[1101]&m[1102])|(m[661]&m[1098]&m[1100]&~m[1101]&m[1102])|(~m[661]&m[1098]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[278])|((m[661]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(~m[661]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[661]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[661]&m[1098]&~m[1100]&~m[1101]&m[1102])|(m[661]&~m[1098]&m[1100]&~m[1101]&m[1102])|(~m[661]&~m[1098]&~m[1100]&m[1101]&m[1102])|(m[661]&~m[1098]&~m[1100]&m[1101]&m[1102])|(~m[661]&m[1098]&~m[1100]&m[1101]&m[1102])|(m[661]&m[1098]&~m[1100]&m[1101]&m[1102])|(~m[661]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[661]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[661]&m[1098]&m[1100]&m[1101]&m[1102]))):InitCond[781];
    m[1104] = run?((((m[674]&~m[1103]&~m[1105]&~m[1106]&~m[1107])|(~m[674]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(m[674]&m[1103]&~m[1105]&m[1106]&~m[1107])|(m[674]&~m[1103]&m[1105]&m[1106]&~m[1107])|(~m[674]&m[1103]&~m[1105]&~m[1106]&m[1107])|(~m[674]&~m[1103]&m[1105]&~m[1106]&m[1107])|(m[674]&m[1103]&m[1105]&~m[1106]&m[1107])|(~m[674]&m[1103]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[279])|((m[674]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(~m[674]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[674]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[674]&m[1103]&~m[1105]&~m[1106]&m[1107])|(m[674]&~m[1103]&m[1105]&~m[1106]&m[1107])|(~m[674]&~m[1103]&~m[1105]&m[1106]&m[1107])|(m[674]&~m[1103]&~m[1105]&m[1106]&m[1107])|(~m[674]&m[1103]&~m[1105]&m[1106]&m[1107])|(m[674]&m[1103]&~m[1105]&m[1106]&m[1107])|(~m[674]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[674]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[674]&m[1103]&m[1105]&m[1106]&m[1107]))):InitCond[782];
    m[1109] = run?((((m[687]&~m[1108]&~m[1110]&~m[1111]&~m[1112])|(~m[687]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(m[687]&m[1108]&~m[1110]&m[1111]&~m[1112])|(m[687]&~m[1108]&m[1110]&m[1111]&~m[1112])|(~m[687]&m[1108]&~m[1110]&~m[1111]&m[1112])|(~m[687]&~m[1108]&m[1110]&~m[1111]&m[1112])|(m[687]&m[1108]&m[1110]&~m[1111]&m[1112])|(~m[687]&m[1108]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[280])|((m[687]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(~m[687]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[687]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[687]&m[1108]&~m[1110]&~m[1111]&m[1112])|(m[687]&~m[1108]&m[1110]&~m[1111]&m[1112])|(~m[687]&~m[1108]&~m[1110]&m[1111]&m[1112])|(m[687]&~m[1108]&~m[1110]&m[1111]&m[1112])|(~m[687]&m[1108]&~m[1110]&m[1111]&m[1112])|(m[687]&m[1108]&~m[1110]&m[1111]&m[1112])|(~m[687]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[687]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[687]&m[1108]&m[1110]&m[1111]&m[1112]))):InitCond[783];
    m[1114] = run?((((m[700]&~m[1113]&~m[1115]&~m[1116]&~m[1117])|(~m[700]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(m[700]&m[1113]&~m[1115]&m[1116]&~m[1117])|(m[700]&~m[1113]&m[1115]&m[1116]&~m[1117])|(~m[700]&m[1113]&~m[1115]&~m[1116]&m[1117])|(~m[700]&~m[1113]&m[1115]&~m[1116]&m[1117])|(m[700]&m[1113]&m[1115]&~m[1116]&m[1117])|(~m[700]&m[1113]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[281])|((m[700]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(~m[700]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[700]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[700]&m[1113]&~m[1115]&~m[1116]&m[1117])|(m[700]&~m[1113]&m[1115]&~m[1116]&m[1117])|(~m[700]&~m[1113]&~m[1115]&m[1116]&m[1117])|(m[700]&~m[1113]&~m[1115]&m[1116]&m[1117])|(~m[700]&m[1113]&~m[1115]&m[1116]&m[1117])|(m[700]&m[1113]&~m[1115]&m[1116]&m[1117])|(~m[700]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[700]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[700]&m[1113]&m[1115]&m[1116]&m[1117]))):InitCond[784];
    m[1119] = run?((((m[558]&~m[1118]&~m[1120]&~m[1121]&~m[1122])|(~m[558]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(m[558]&m[1118]&~m[1120]&m[1121]&~m[1122])|(m[558]&~m[1118]&m[1120]&m[1121]&~m[1122])|(~m[558]&m[1118]&~m[1120]&~m[1121]&m[1122])|(~m[558]&~m[1118]&m[1120]&~m[1121]&m[1122])|(m[558]&m[1118]&m[1120]&~m[1121]&m[1122])|(~m[558]&m[1118]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[282])|((m[558]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(~m[558]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[558]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[558]&m[1118]&~m[1120]&~m[1121]&m[1122])|(m[558]&~m[1118]&m[1120]&~m[1121]&m[1122])|(~m[558]&~m[1118]&~m[1120]&m[1121]&m[1122])|(m[558]&~m[1118]&~m[1120]&m[1121]&m[1122])|(~m[558]&m[1118]&~m[1120]&m[1121]&m[1122])|(m[558]&m[1118]&~m[1120]&m[1121]&m[1122])|(~m[558]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[558]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[558]&m[1118]&m[1120]&m[1121]&m[1122]))):InitCond[785];
    m[1124] = run?((((m[571]&~m[1123]&~m[1125]&~m[1126]&~m[1127])|(~m[571]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(m[571]&m[1123]&~m[1125]&m[1126]&~m[1127])|(m[571]&~m[1123]&m[1125]&m[1126]&~m[1127])|(~m[571]&m[1123]&~m[1125]&~m[1126]&m[1127])|(~m[571]&~m[1123]&m[1125]&~m[1126]&m[1127])|(m[571]&m[1123]&m[1125]&~m[1126]&m[1127])|(~m[571]&m[1123]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[283])|((m[571]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(~m[571]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[571]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[571]&m[1123]&~m[1125]&~m[1126]&m[1127])|(m[571]&~m[1123]&m[1125]&~m[1126]&m[1127])|(~m[571]&~m[1123]&~m[1125]&m[1126]&m[1127])|(m[571]&~m[1123]&~m[1125]&m[1126]&m[1127])|(~m[571]&m[1123]&~m[1125]&m[1126]&m[1127])|(m[571]&m[1123]&~m[1125]&m[1126]&m[1127])|(~m[571]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[571]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[571]&m[1123]&m[1125]&m[1126]&m[1127]))):InitCond[786];
    m[1129] = run?((((m[584]&~m[1128]&~m[1130]&~m[1131]&~m[1132])|(~m[584]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(m[584]&m[1128]&~m[1130]&m[1131]&~m[1132])|(m[584]&~m[1128]&m[1130]&m[1131]&~m[1132])|(~m[584]&m[1128]&~m[1130]&~m[1131]&m[1132])|(~m[584]&~m[1128]&m[1130]&~m[1131]&m[1132])|(m[584]&m[1128]&m[1130]&~m[1131]&m[1132])|(~m[584]&m[1128]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[284])|((m[584]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(~m[584]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[584]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[584]&m[1128]&~m[1130]&~m[1131]&m[1132])|(m[584]&~m[1128]&m[1130]&~m[1131]&m[1132])|(~m[584]&~m[1128]&~m[1130]&m[1131]&m[1132])|(m[584]&~m[1128]&~m[1130]&m[1131]&m[1132])|(~m[584]&m[1128]&~m[1130]&m[1131]&m[1132])|(m[584]&m[1128]&~m[1130]&m[1131]&m[1132])|(~m[584]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[584]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[584]&m[1128]&m[1130]&m[1131]&m[1132]))):InitCond[787];
    m[1134] = run?((((m[597]&~m[1133]&~m[1135]&~m[1136]&~m[1137])|(~m[597]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(m[597]&m[1133]&~m[1135]&m[1136]&~m[1137])|(m[597]&~m[1133]&m[1135]&m[1136]&~m[1137])|(~m[597]&m[1133]&~m[1135]&~m[1136]&m[1137])|(~m[597]&~m[1133]&m[1135]&~m[1136]&m[1137])|(m[597]&m[1133]&m[1135]&~m[1136]&m[1137])|(~m[597]&m[1133]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[285])|((m[597]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(~m[597]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[597]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[597]&m[1133]&~m[1135]&~m[1136]&m[1137])|(m[597]&~m[1133]&m[1135]&~m[1136]&m[1137])|(~m[597]&~m[1133]&~m[1135]&m[1136]&m[1137])|(m[597]&~m[1133]&~m[1135]&m[1136]&m[1137])|(~m[597]&m[1133]&~m[1135]&m[1136]&m[1137])|(m[597]&m[1133]&~m[1135]&m[1136]&m[1137])|(~m[597]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[597]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[597]&m[1133]&m[1135]&m[1136]&m[1137]))):InitCond[788];
    m[1139] = run?((((m[610]&~m[1138]&~m[1140]&~m[1141]&~m[1142])|(~m[610]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(m[610]&m[1138]&~m[1140]&m[1141]&~m[1142])|(m[610]&~m[1138]&m[1140]&m[1141]&~m[1142])|(~m[610]&m[1138]&~m[1140]&~m[1141]&m[1142])|(~m[610]&~m[1138]&m[1140]&~m[1141]&m[1142])|(m[610]&m[1138]&m[1140]&~m[1141]&m[1142])|(~m[610]&m[1138]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[286])|((m[610]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(~m[610]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[610]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[610]&m[1138]&~m[1140]&~m[1141]&m[1142])|(m[610]&~m[1138]&m[1140]&~m[1141]&m[1142])|(~m[610]&~m[1138]&~m[1140]&m[1141]&m[1142])|(m[610]&~m[1138]&~m[1140]&m[1141]&m[1142])|(~m[610]&m[1138]&~m[1140]&m[1141]&m[1142])|(m[610]&m[1138]&~m[1140]&m[1141]&m[1142])|(~m[610]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[610]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[610]&m[1138]&m[1140]&m[1141]&m[1142]))):InitCond[789];
    m[1144] = run?((((m[623]&~m[1143]&~m[1145]&~m[1146]&~m[1147])|(~m[623]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(m[623]&m[1143]&~m[1145]&m[1146]&~m[1147])|(m[623]&~m[1143]&m[1145]&m[1146]&~m[1147])|(~m[623]&m[1143]&~m[1145]&~m[1146]&m[1147])|(~m[623]&~m[1143]&m[1145]&~m[1146]&m[1147])|(m[623]&m[1143]&m[1145]&~m[1146]&m[1147])|(~m[623]&m[1143]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[287])|((m[623]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(~m[623]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[623]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[623]&m[1143]&~m[1145]&~m[1146]&m[1147])|(m[623]&~m[1143]&m[1145]&~m[1146]&m[1147])|(~m[623]&~m[1143]&~m[1145]&m[1146]&m[1147])|(m[623]&~m[1143]&~m[1145]&m[1146]&m[1147])|(~m[623]&m[1143]&~m[1145]&m[1146]&m[1147])|(m[623]&m[1143]&~m[1145]&m[1146]&m[1147])|(~m[623]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[623]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[623]&m[1143]&m[1145]&m[1146]&m[1147]))):InitCond[790];
    m[1149] = run?((((m[636]&~m[1148]&~m[1150]&~m[1151]&~m[1152])|(~m[636]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(m[636]&m[1148]&~m[1150]&m[1151]&~m[1152])|(m[636]&~m[1148]&m[1150]&m[1151]&~m[1152])|(~m[636]&m[1148]&~m[1150]&~m[1151]&m[1152])|(~m[636]&~m[1148]&m[1150]&~m[1151]&m[1152])|(m[636]&m[1148]&m[1150]&~m[1151]&m[1152])|(~m[636]&m[1148]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[288])|((m[636]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(~m[636]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[636]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[636]&m[1148]&~m[1150]&~m[1151]&m[1152])|(m[636]&~m[1148]&m[1150]&~m[1151]&m[1152])|(~m[636]&~m[1148]&~m[1150]&m[1151]&m[1152])|(m[636]&~m[1148]&~m[1150]&m[1151]&m[1152])|(~m[636]&m[1148]&~m[1150]&m[1151]&m[1152])|(m[636]&m[1148]&~m[1150]&m[1151]&m[1152])|(~m[636]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[636]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[636]&m[1148]&m[1150]&m[1151]&m[1152]))):InitCond[791];
    m[1154] = run?((((m[649]&~m[1153]&~m[1155]&~m[1156]&~m[1157])|(~m[649]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(m[649]&m[1153]&~m[1155]&m[1156]&~m[1157])|(m[649]&~m[1153]&m[1155]&m[1156]&~m[1157])|(~m[649]&m[1153]&~m[1155]&~m[1156]&m[1157])|(~m[649]&~m[1153]&m[1155]&~m[1156]&m[1157])|(m[649]&m[1153]&m[1155]&~m[1156]&m[1157])|(~m[649]&m[1153]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[289])|((m[649]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(~m[649]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[649]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[649]&m[1153]&~m[1155]&~m[1156]&m[1157])|(m[649]&~m[1153]&m[1155]&~m[1156]&m[1157])|(~m[649]&~m[1153]&~m[1155]&m[1156]&m[1157])|(m[649]&~m[1153]&~m[1155]&m[1156]&m[1157])|(~m[649]&m[1153]&~m[1155]&m[1156]&m[1157])|(m[649]&m[1153]&~m[1155]&m[1156]&m[1157])|(~m[649]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[649]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[649]&m[1153]&m[1155]&m[1156]&m[1157]))):InitCond[792];
    m[1159] = run?((((m[662]&~m[1158]&~m[1160]&~m[1161]&~m[1162])|(~m[662]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(m[662]&m[1158]&~m[1160]&m[1161]&~m[1162])|(m[662]&~m[1158]&m[1160]&m[1161]&~m[1162])|(~m[662]&m[1158]&~m[1160]&~m[1161]&m[1162])|(~m[662]&~m[1158]&m[1160]&~m[1161]&m[1162])|(m[662]&m[1158]&m[1160]&~m[1161]&m[1162])|(~m[662]&m[1158]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[290])|((m[662]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(~m[662]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[662]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[662]&m[1158]&~m[1160]&~m[1161]&m[1162])|(m[662]&~m[1158]&m[1160]&~m[1161]&m[1162])|(~m[662]&~m[1158]&~m[1160]&m[1161]&m[1162])|(m[662]&~m[1158]&~m[1160]&m[1161]&m[1162])|(~m[662]&m[1158]&~m[1160]&m[1161]&m[1162])|(m[662]&m[1158]&~m[1160]&m[1161]&m[1162])|(~m[662]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[662]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[662]&m[1158]&m[1160]&m[1161]&m[1162]))):InitCond[793];
    m[1164] = run?((((m[675]&~m[1163]&~m[1165]&~m[1166]&~m[1167])|(~m[675]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(m[675]&m[1163]&~m[1165]&m[1166]&~m[1167])|(m[675]&~m[1163]&m[1165]&m[1166]&~m[1167])|(~m[675]&m[1163]&~m[1165]&~m[1166]&m[1167])|(~m[675]&~m[1163]&m[1165]&~m[1166]&m[1167])|(m[675]&m[1163]&m[1165]&~m[1166]&m[1167])|(~m[675]&m[1163]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[291])|((m[675]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(~m[675]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[675]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[675]&m[1163]&~m[1165]&~m[1166]&m[1167])|(m[675]&~m[1163]&m[1165]&~m[1166]&m[1167])|(~m[675]&~m[1163]&~m[1165]&m[1166]&m[1167])|(m[675]&~m[1163]&~m[1165]&m[1166]&m[1167])|(~m[675]&m[1163]&~m[1165]&m[1166]&m[1167])|(m[675]&m[1163]&~m[1165]&m[1166]&m[1167])|(~m[675]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[675]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[675]&m[1163]&m[1165]&m[1166]&m[1167]))):InitCond[794];
    m[1169] = run?((((m[688]&~m[1168]&~m[1170]&~m[1171]&~m[1172])|(~m[688]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(m[688]&m[1168]&~m[1170]&m[1171]&~m[1172])|(m[688]&~m[1168]&m[1170]&m[1171]&~m[1172])|(~m[688]&m[1168]&~m[1170]&~m[1171]&m[1172])|(~m[688]&~m[1168]&m[1170]&~m[1171]&m[1172])|(m[688]&m[1168]&m[1170]&~m[1171]&m[1172])|(~m[688]&m[1168]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[292])|((m[688]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(~m[688]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[688]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[688]&m[1168]&~m[1170]&~m[1171]&m[1172])|(m[688]&~m[1168]&m[1170]&~m[1171]&m[1172])|(~m[688]&~m[1168]&~m[1170]&m[1171]&m[1172])|(m[688]&~m[1168]&~m[1170]&m[1171]&m[1172])|(~m[688]&m[1168]&~m[1170]&m[1171]&m[1172])|(m[688]&m[1168]&~m[1170]&m[1171]&m[1172])|(~m[688]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[688]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[688]&m[1168]&m[1170]&m[1171]&m[1172]))):InitCond[795];
    m[1174] = run?((((m[701]&~m[1173]&~m[1175]&~m[1176]&~m[1177])|(~m[701]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(m[701]&m[1173]&~m[1175]&m[1176]&~m[1177])|(m[701]&~m[1173]&m[1175]&m[1176]&~m[1177])|(~m[701]&m[1173]&~m[1175]&~m[1176]&m[1177])|(~m[701]&~m[1173]&m[1175]&~m[1176]&m[1177])|(m[701]&m[1173]&m[1175]&~m[1176]&m[1177])|(~m[701]&m[1173]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[293])|((m[701]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(~m[701]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[701]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[701]&m[1173]&~m[1175]&~m[1176]&m[1177])|(m[701]&~m[1173]&m[1175]&~m[1176]&m[1177])|(~m[701]&~m[1173]&~m[1175]&m[1176]&m[1177])|(m[701]&~m[1173]&~m[1175]&m[1176]&m[1177])|(~m[701]&m[1173]&~m[1175]&m[1176]&m[1177])|(m[701]&m[1173]&~m[1175]&m[1176]&m[1177])|(~m[701]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[701]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[701]&m[1173]&m[1175]&m[1176]&m[1177]))):InitCond[796];
    m[1179] = run?((((m[714]&~m[1178]&~m[1180]&~m[1181]&~m[1182])|(~m[714]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(m[714]&m[1178]&~m[1180]&m[1181]&~m[1182])|(m[714]&~m[1178]&m[1180]&m[1181]&~m[1182])|(~m[714]&m[1178]&~m[1180]&~m[1181]&m[1182])|(~m[714]&~m[1178]&m[1180]&~m[1181]&m[1182])|(m[714]&m[1178]&m[1180]&~m[1181]&m[1182])|(~m[714]&m[1178]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[294])|((m[714]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(~m[714]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[714]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[714]&m[1178]&~m[1180]&~m[1181]&m[1182])|(m[714]&~m[1178]&m[1180]&~m[1181]&m[1182])|(~m[714]&~m[1178]&~m[1180]&m[1181]&m[1182])|(m[714]&~m[1178]&~m[1180]&m[1181]&m[1182])|(~m[714]&m[1178]&~m[1180]&m[1181]&m[1182])|(m[714]&m[1178]&~m[1180]&m[1181]&m[1182])|(~m[714]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[714]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[714]&m[1178]&m[1180]&m[1181]&m[1182]))):InitCond[797];
    m[1184] = run?((((m[559]&~m[1183]&~m[1185]&~m[1186]&~m[1187])|(~m[559]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(m[559]&m[1183]&~m[1185]&m[1186]&~m[1187])|(m[559]&~m[1183]&m[1185]&m[1186]&~m[1187])|(~m[559]&m[1183]&~m[1185]&~m[1186]&m[1187])|(~m[559]&~m[1183]&m[1185]&~m[1186]&m[1187])|(m[559]&m[1183]&m[1185]&~m[1186]&m[1187])|(~m[559]&m[1183]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[295])|((m[559]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(~m[559]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[559]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[559]&m[1183]&~m[1185]&~m[1186]&m[1187])|(m[559]&~m[1183]&m[1185]&~m[1186]&m[1187])|(~m[559]&~m[1183]&~m[1185]&m[1186]&m[1187])|(m[559]&~m[1183]&~m[1185]&m[1186]&m[1187])|(~m[559]&m[1183]&~m[1185]&m[1186]&m[1187])|(m[559]&m[1183]&~m[1185]&m[1186]&m[1187])|(~m[559]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[559]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[559]&m[1183]&m[1185]&m[1186]&m[1187]))):InitCond[798];
    m[1189] = run?((((m[572]&~m[1188]&~m[1190]&~m[1191]&~m[1192])|(~m[572]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(m[572]&m[1188]&~m[1190]&m[1191]&~m[1192])|(m[572]&~m[1188]&m[1190]&m[1191]&~m[1192])|(~m[572]&m[1188]&~m[1190]&~m[1191]&m[1192])|(~m[572]&~m[1188]&m[1190]&~m[1191]&m[1192])|(m[572]&m[1188]&m[1190]&~m[1191]&m[1192])|(~m[572]&m[1188]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[296])|((m[572]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(~m[572]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[572]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[572]&m[1188]&~m[1190]&~m[1191]&m[1192])|(m[572]&~m[1188]&m[1190]&~m[1191]&m[1192])|(~m[572]&~m[1188]&~m[1190]&m[1191]&m[1192])|(m[572]&~m[1188]&~m[1190]&m[1191]&m[1192])|(~m[572]&m[1188]&~m[1190]&m[1191]&m[1192])|(m[572]&m[1188]&~m[1190]&m[1191]&m[1192])|(~m[572]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[572]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[572]&m[1188]&m[1190]&m[1191]&m[1192]))):InitCond[799];
    m[1194] = run?((((m[585]&~m[1193]&~m[1195]&~m[1196]&~m[1197])|(~m[585]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(m[585]&m[1193]&~m[1195]&m[1196]&~m[1197])|(m[585]&~m[1193]&m[1195]&m[1196]&~m[1197])|(~m[585]&m[1193]&~m[1195]&~m[1196]&m[1197])|(~m[585]&~m[1193]&m[1195]&~m[1196]&m[1197])|(m[585]&m[1193]&m[1195]&~m[1196]&m[1197])|(~m[585]&m[1193]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[297])|((m[585]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(~m[585]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[585]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[585]&m[1193]&~m[1195]&~m[1196]&m[1197])|(m[585]&~m[1193]&m[1195]&~m[1196]&m[1197])|(~m[585]&~m[1193]&~m[1195]&m[1196]&m[1197])|(m[585]&~m[1193]&~m[1195]&m[1196]&m[1197])|(~m[585]&m[1193]&~m[1195]&m[1196]&m[1197])|(m[585]&m[1193]&~m[1195]&m[1196]&m[1197])|(~m[585]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[585]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[585]&m[1193]&m[1195]&m[1196]&m[1197]))):InitCond[800];
    m[1199] = run?((((m[598]&~m[1198]&~m[1200]&~m[1201]&~m[1202])|(~m[598]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(m[598]&m[1198]&~m[1200]&m[1201]&~m[1202])|(m[598]&~m[1198]&m[1200]&m[1201]&~m[1202])|(~m[598]&m[1198]&~m[1200]&~m[1201]&m[1202])|(~m[598]&~m[1198]&m[1200]&~m[1201]&m[1202])|(m[598]&m[1198]&m[1200]&~m[1201]&m[1202])|(~m[598]&m[1198]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[298])|((m[598]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(~m[598]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[598]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[598]&m[1198]&~m[1200]&~m[1201]&m[1202])|(m[598]&~m[1198]&m[1200]&~m[1201]&m[1202])|(~m[598]&~m[1198]&~m[1200]&m[1201]&m[1202])|(m[598]&~m[1198]&~m[1200]&m[1201]&m[1202])|(~m[598]&m[1198]&~m[1200]&m[1201]&m[1202])|(m[598]&m[1198]&~m[1200]&m[1201]&m[1202])|(~m[598]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[598]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[598]&m[1198]&m[1200]&m[1201]&m[1202]))):InitCond[801];
    m[1204] = run?((((m[611]&~m[1203]&~m[1205]&~m[1206]&~m[1207])|(~m[611]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(m[611]&m[1203]&~m[1205]&m[1206]&~m[1207])|(m[611]&~m[1203]&m[1205]&m[1206]&~m[1207])|(~m[611]&m[1203]&~m[1205]&~m[1206]&m[1207])|(~m[611]&~m[1203]&m[1205]&~m[1206]&m[1207])|(m[611]&m[1203]&m[1205]&~m[1206]&m[1207])|(~m[611]&m[1203]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[299])|((m[611]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(~m[611]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[611]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[611]&m[1203]&~m[1205]&~m[1206]&m[1207])|(m[611]&~m[1203]&m[1205]&~m[1206]&m[1207])|(~m[611]&~m[1203]&~m[1205]&m[1206]&m[1207])|(m[611]&~m[1203]&~m[1205]&m[1206]&m[1207])|(~m[611]&m[1203]&~m[1205]&m[1206]&m[1207])|(m[611]&m[1203]&~m[1205]&m[1206]&m[1207])|(~m[611]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[611]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[611]&m[1203]&m[1205]&m[1206]&m[1207]))):InitCond[802];
    m[1209] = run?((((m[624]&~m[1208]&~m[1210]&~m[1211]&~m[1212])|(~m[624]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(m[624]&m[1208]&~m[1210]&m[1211]&~m[1212])|(m[624]&~m[1208]&m[1210]&m[1211]&~m[1212])|(~m[624]&m[1208]&~m[1210]&~m[1211]&m[1212])|(~m[624]&~m[1208]&m[1210]&~m[1211]&m[1212])|(m[624]&m[1208]&m[1210]&~m[1211]&m[1212])|(~m[624]&m[1208]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[300])|((m[624]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(~m[624]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[624]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[624]&m[1208]&~m[1210]&~m[1211]&m[1212])|(m[624]&~m[1208]&m[1210]&~m[1211]&m[1212])|(~m[624]&~m[1208]&~m[1210]&m[1211]&m[1212])|(m[624]&~m[1208]&~m[1210]&m[1211]&m[1212])|(~m[624]&m[1208]&~m[1210]&m[1211]&m[1212])|(m[624]&m[1208]&~m[1210]&m[1211]&m[1212])|(~m[624]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[624]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[624]&m[1208]&m[1210]&m[1211]&m[1212]))):InitCond[803];
    m[1214] = run?((((m[637]&~m[1213]&~m[1215]&~m[1216]&~m[1217])|(~m[637]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(m[637]&m[1213]&~m[1215]&m[1216]&~m[1217])|(m[637]&~m[1213]&m[1215]&m[1216]&~m[1217])|(~m[637]&m[1213]&~m[1215]&~m[1216]&m[1217])|(~m[637]&~m[1213]&m[1215]&~m[1216]&m[1217])|(m[637]&m[1213]&m[1215]&~m[1216]&m[1217])|(~m[637]&m[1213]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[301])|((m[637]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(~m[637]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[637]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[637]&m[1213]&~m[1215]&~m[1216]&m[1217])|(m[637]&~m[1213]&m[1215]&~m[1216]&m[1217])|(~m[637]&~m[1213]&~m[1215]&m[1216]&m[1217])|(m[637]&~m[1213]&~m[1215]&m[1216]&m[1217])|(~m[637]&m[1213]&~m[1215]&m[1216]&m[1217])|(m[637]&m[1213]&~m[1215]&m[1216]&m[1217])|(~m[637]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[637]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[637]&m[1213]&m[1215]&m[1216]&m[1217]))):InitCond[804];
    m[1219] = run?((((m[650]&~m[1218]&~m[1220]&~m[1221]&~m[1222])|(~m[650]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(m[650]&m[1218]&~m[1220]&m[1221]&~m[1222])|(m[650]&~m[1218]&m[1220]&m[1221]&~m[1222])|(~m[650]&m[1218]&~m[1220]&~m[1221]&m[1222])|(~m[650]&~m[1218]&m[1220]&~m[1221]&m[1222])|(m[650]&m[1218]&m[1220]&~m[1221]&m[1222])|(~m[650]&m[1218]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[302])|((m[650]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(~m[650]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[650]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[650]&m[1218]&~m[1220]&~m[1221]&m[1222])|(m[650]&~m[1218]&m[1220]&~m[1221]&m[1222])|(~m[650]&~m[1218]&~m[1220]&m[1221]&m[1222])|(m[650]&~m[1218]&~m[1220]&m[1221]&m[1222])|(~m[650]&m[1218]&~m[1220]&m[1221]&m[1222])|(m[650]&m[1218]&~m[1220]&m[1221]&m[1222])|(~m[650]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[650]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[650]&m[1218]&m[1220]&m[1221]&m[1222]))):InitCond[805];
    m[1224] = run?((((m[663]&~m[1223]&~m[1225]&~m[1226]&~m[1227])|(~m[663]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(m[663]&m[1223]&~m[1225]&m[1226]&~m[1227])|(m[663]&~m[1223]&m[1225]&m[1226]&~m[1227])|(~m[663]&m[1223]&~m[1225]&~m[1226]&m[1227])|(~m[663]&~m[1223]&m[1225]&~m[1226]&m[1227])|(m[663]&m[1223]&m[1225]&~m[1226]&m[1227])|(~m[663]&m[1223]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[303])|((m[663]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(~m[663]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[663]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[663]&m[1223]&~m[1225]&~m[1226]&m[1227])|(m[663]&~m[1223]&m[1225]&~m[1226]&m[1227])|(~m[663]&~m[1223]&~m[1225]&m[1226]&m[1227])|(m[663]&~m[1223]&~m[1225]&m[1226]&m[1227])|(~m[663]&m[1223]&~m[1225]&m[1226]&m[1227])|(m[663]&m[1223]&~m[1225]&m[1226]&m[1227])|(~m[663]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[663]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[663]&m[1223]&m[1225]&m[1226]&m[1227]))):InitCond[806];
    m[1229] = run?((((m[676]&~m[1228]&~m[1230]&~m[1231]&~m[1232])|(~m[676]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(m[676]&m[1228]&~m[1230]&m[1231]&~m[1232])|(m[676]&~m[1228]&m[1230]&m[1231]&~m[1232])|(~m[676]&m[1228]&~m[1230]&~m[1231]&m[1232])|(~m[676]&~m[1228]&m[1230]&~m[1231]&m[1232])|(m[676]&m[1228]&m[1230]&~m[1231]&m[1232])|(~m[676]&m[1228]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[304])|((m[676]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(~m[676]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[676]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[676]&m[1228]&~m[1230]&~m[1231]&m[1232])|(m[676]&~m[1228]&m[1230]&~m[1231]&m[1232])|(~m[676]&~m[1228]&~m[1230]&m[1231]&m[1232])|(m[676]&~m[1228]&~m[1230]&m[1231]&m[1232])|(~m[676]&m[1228]&~m[1230]&m[1231]&m[1232])|(m[676]&m[1228]&~m[1230]&m[1231]&m[1232])|(~m[676]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[676]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[676]&m[1228]&m[1230]&m[1231]&m[1232]))):InitCond[807];
    m[1234] = run?((((m[689]&~m[1233]&~m[1235]&~m[1236]&~m[1237])|(~m[689]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(m[689]&m[1233]&~m[1235]&m[1236]&~m[1237])|(m[689]&~m[1233]&m[1235]&m[1236]&~m[1237])|(~m[689]&m[1233]&~m[1235]&~m[1236]&m[1237])|(~m[689]&~m[1233]&m[1235]&~m[1236]&m[1237])|(m[689]&m[1233]&m[1235]&~m[1236]&m[1237])|(~m[689]&m[1233]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[305])|((m[689]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(~m[689]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[689]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[689]&m[1233]&~m[1235]&~m[1236]&m[1237])|(m[689]&~m[1233]&m[1235]&~m[1236]&m[1237])|(~m[689]&~m[1233]&~m[1235]&m[1236]&m[1237])|(m[689]&~m[1233]&~m[1235]&m[1236]&m[1237])|(~m[689]&m[1233]&~m[1235]&m[1236]&m[1237])|(m[689]&m[1233]&~m[1235]&m[1236]&m[1237])|(~m[689]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[689]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[689]&m[1233]&m[1235]&m[1236]&m[1237]))):InitCond[808];
    m[1239] = run?((((m[702]&~m[1238]&~m[1240]&~m[1241]&~m[1242])|(~m[702]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(m[702]&m[1238]&~m[1240]&m[1241]&~m[1242])|(m[702]&~m[1238]&m[1240]&m[1241]&~m[1242])|(~m[702]&m[1238]&~m[1240]&~m[1241]&m[1242])|(~m[702]&~m[1238]&m[1240]&~m[1241]&m[1242])|(m[702]&m[1238]&m[1240]&~m[1241]&m[1242])|(~m[702]&m[1238]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[306])|((m[702]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(~m[702]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[702]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[702]&m[1238]&~m[1240]&~m[1241]&m[1242])|(m[702]&~m[1238]&m[1240]&~m[1241]&m[1242])|(~m[702]&~m[1238]&~m[1240]&m[1241]&m[1242])|(m[702]&~m[1238]&~m[1240]&m[1241]&m[1242])|(~m[702]&m[1238]&~m[1240]&m[1241]&m[1242])|(m[702]&m[1238]&~m[1240]&m[1241]&m[1242])|(~m[702]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[702]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[702]&m[1238]&m[1240]&m[1241]&m[1242]))):InitCond[809];
    m[1244] = run?((((m[715]&~m[1243]&~m[1245]&~m[1246]&~m[1247])|(~m[715]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(m[715]&m[1243]&~m[1245]&m[1246]&~m[1247])|(m[715]&~m[1243]&m[1245]&m[1246]&~m[1247])|(~m[715]&m[1243]&~m[1245]&~m[1246]&m[1247])|(~m[715]&~m[1243]&m[1245]&~m[1246]&m[1247])|(m[715]&m[1243]&m[1245]&~m[1246]&m[1247])|(~m[715]&m[1243]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[307])|((m[715]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(~m[715]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[715]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[715]&m[1243]&~m[1245]&~m[1246]&m[1247])|(m[715]&~m[1243]&m[1245]&~m[1246]&m[1247])|(~m[715]&~m[1243]&~m[1245]&m[1246]&m[1247])|(m[715]&~m[1243]&~m[1245]&m[1246]&m[1247])|(~m[715]&m[1243]&~m[1245]&m[1246]&m[1247])|(m[715]&m[1243]&~m[1245]&m[1246]&m[1247])|(~m[715]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[715]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[715]&m[1243]&m[1245]&m[1246]&m[1247]))):InitCond[810];
    m[1249] = run?((((m[573]&~m[1248]&~m[1250]&~m[1251]&~m[1252])|(~m[573]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(m[573]&m[1248]&~m[1250]&m[1251]&~m[1252])|(m[573]&~m[1248]&m[1250]&m[1251]&~m[1252])|(~m[573]&m[1248]&~m[1250]&~m[1251]&m[1252])|(~m[573]&~m[1248]&m[1250]&~m[1251]&m[1252])|(m[573]&m[1248]&m[1250]&~m[1251]&m[1252])|(~m[573]&m[1248]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[308])|((m[573]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(~m[573]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[573]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[573]&m[1248]&~m[1250]&~m[1251]&m[1252])|(m[573]&~m[1248]&m[1250]&~m[1251]&m[1252])|(~m[573]&~m[1248]&~m[1250]&m[1251]&m[1252])|(m[573]&~m[1248]&~m[1250]&m[1251]&m[1252])|(~m[573]&m[1248]&~m[1250]&m[1251]&m[1252])|(m[573]&m[1248]&~m[1250]&m[1251]&m[1252])|(~m[573]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[573]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[573]&m[1248]&m[1250]&m[1251]&m[1252]))):InitCond[811];
    m[1254] = run?((((m[586]&~m[1253]&~m[1255]&~m[1256]&~m[1257])|(~m[586]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(m[586]&m[1253]&~m[1255]&m[1256]&~m[1257])|(m[586]&~m[1253]&m[1255]&m[1256]&~m[1257])|(~m[586]&m[1253]&~m[1255]&~m[1256]&m[1257])|(~m[586]&~m[1253]&m[1255]&~m[1256]&m[1257])|(m[586]&m[1253]&m[1255]&~m[1256]&m[1257])|(~m[586]&m[1253]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[309])|((m[586]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(~m[586]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[586]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[586]&m[1253]&~m[1255]&~m[1256]&m[1257])|(m[586]&~m[1253]&m[1255]&~m[1256]&m[1257])|(~m[586]&~m[1253]&~m[1255]&m[1256]&m[1257])|(m[586]&~m[1253]&~m[1255]&m[1256]&m[1257])|(~m[586]&m[1253]&~m[1255]&m[1256]&m[1257])|(m[586]&m[1253]&~m[1255]&m[1256]&m[1257])|(~m[586]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[586]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[586]&m[1253]&m[1255]&m[1256]&m[1257]))):InitCond[812];
    m[1259] = run?((((m[599]&~m[1258]&~m[1260]&~m[1261]&~m[1262])|(~m[599]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(m[599]&m[1258]&~m[1260]&m[1261]&~m[1262])|(m[599]&~m[1258]&m[1260]&m[1261]&~m[1262])|(~m[599]&m[1258]&~m[1260]&~m[1261]&m[1262])|(~m[599]&~m[1258]&m[1260]&~m[1261]&m[1262])|(m[599]&m[1258]&m[1260]&~m[1261]&m[1262])|(~m[599]&m[1258]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[310])|((m[599]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(~m[599]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[599]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[599]&m[1258]&~m[1260]&~m[1261]&m[1262])|(m[599]&~m[1258]&m[1260]&~m[1261]&m[1262])|(~m[599]&~m[1258]&~m[1260]&m[1261]&m[1262])|(m[599]&~m[1258]&~m[1260]&m[1261]&m[1262])|(~m[599]&m[1258]&~m[1260]&m[1261]&m[1262])|(m[599]&m[1258]&~m[1260]&m[1261]&m[1262])|(~m[599]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[599]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[599]&m[1258]&m[1260]&m[1261]&m[1262]))):InitCond[813];
    m[1264] = run?((((m[612]&~m[1263]&~m[1265]&~m[1266]&~m[1267])|(~m[612]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(m[612]&m[1263]&~m[1265]&m[1266]&~m[1267])|(m[612]&~m[1263]&m[1265]&m[1266]&~m[1267])|(~m[612]&m[1263]&~m[1265]&~m[1266]&m[1267])|(~m[612]&~m[1263]&m[1265]&~m[1266]&m[1267])|(m[612]&m[1263]&m[1265]&~m[1266]&m[1267])|(~m[612]&m[1263]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[311])|((m[612]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(~m[612]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[612]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[612]&m[1263]&~m[1265]&~m[1266]&m[1267])|(m[612]&~m[1263]&m[1265]&~m[1266]&m[1267])|(~m[612]&~m[1263]&~m[1265]&m[1266]&m[1267])|(m[612]&~m[1263]&~m[1265]&m[1266]&m[1267])|(~m[612]&m[1263]&~m[1265]&m[1266]&m[1267])|(m[612]&m[1263]&~m[1265]&m[1266]&m[1267])|(~m[612]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[612]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[612]&m[1263]&m[1265]&m[1266]&m[1267]))):InitCond[814];
    m[1269] = run?((((m[625]&~m[1268]&~m[1270]&~m[1271]&~m[1272])|(~m[625]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(m[625]&m[1268]&~m[1270]&m[1271]&~m[1272])|(m[625]&~m[1268]&m[1270]&m[1271]&~m[1272])|(~m[625]&m[1268]&~m[1270]&~m[1271]&m[1272])|(~m[625]&~m[1268]&m[1270]&~m[1271]&m[1272])|(m[625]&m[1268]&m[1270]&~m[1271]&m[1272])|(~m[625]&m[1268]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[312])|((m[625]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(~m[625]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[625]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[625]&m[1268]&~m[1270]&~m[1271]&m[1272])|(m[625]&~m[1268]&m[1270]&~m[1271]&m[1272])|(~m[625]&~m[1268]&~m[1270]&m[1271]&m[1272])|(m[625]&~m[1268]&~m[1270]&m[1271]&m[1272])|(~m[625]&m[1268]&~m[1270]&m[1271]&m[1272])|(m[625]&m[1268]&~m[1270]&m[1271]&m[1272])|(~m[625]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[625]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[625]&m[1268]&m[1270]&m[1271]&m[1272]))):InitCond[815];
    m[1274] = run?((((m[638]&~m[1273]&~m[1275]&~m[1276]&~m[1277])|(~m[638]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(m[638]&m[1273]&~m[1275]&m[1276]&~m[1277])|(m[638]&~m[1273]&m[1275]&m[1276]&~m[1277])|(~m[638]&m[1273]&~m[1275]&~m[1276]&m[1277])|(~m[638]&~m[1273]&m[1275]&~m[1276]&m[1277])|(m[638]&m[1273]&m[1275]&~m[1276]&m[1277])|(~m[638]&m[1273]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[313])|((m[638]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(~m[638]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[638]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[638]&m[1273]&~m[1275]&~m[1276]&m[1277])|(m[638]&~m[1273]&m[1275]&~m[1276]&m[1277])|(~m[638]&~m[1273]&~m[1275]&m[1276]&m[1277])|(m[638]&~m[1273]&~m[1275]&m[1276]&m[1277])|(~m[638]&m[1273]&~m[1275]&m[1276]&m[1277])|(m[638]&m[1273]&~m[1275]&m[1276]&m[1277])|(~m[638]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[638]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[638]&m[1273]&m[1275]&m[1276]&m[1277]))):InitCond[816];
    m[1279] = run?((((m[651]&~m[1278]&~m[1280]&~m[1281]&~m[1282])|(~m[651]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(m[651]&m[1278]&~m[1280]&m[1281]&~m[1282])|(m[651]&~m[1278]&m[1280]&m[1281]&~m[1282])|(~m[651]&m[1278]&~m[1280]&~m[1281]&m[1282])|(~m[651]&~m[1278]&m[1280]&~m[1281]&m[1282])|(m[651]&m[1278]&m[1280]&~m[1281]&m[1282])|(~m[651]&m[1278]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[314])|((m[651]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(~m[651]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[651]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[651]&m[1278]&~m[1280]&~m[1281]&m[1282])|(m[651]&~m[1278]&m[1280]&~m[1281]&m[1282])|(~m[651]&~m[1278]&~m[1280]&m[1281]&m[1282])|(m[651]&~m[1278]&~m[1280]&m[1281]&m[1282])|(~m[651]&m[1278]&~m[1280]&m[1281]&m[1282])|(m[651]&m[1278]&~m[1280]&m[1281]&m[1282])|(~m[651]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[651]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[651]&m[1278]&m[1280]&m[1281]&m[1282]))):InitCond[817];
    m[1284] = run?((((m[664]&~m[1283]&~m[1285]&~m[1286]&~m[1287])|(~m[664]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(m[664]&m[1283]&~m[1285]&m[1286]&~m[1287])|(m[664]&~m[1283]&m[1285]&m[1286]&~m[1287])|(~m[664]&m[1283]&~m[1285]&~m[1286]&m[1287])|(~m[664]&~m[1283]&m[1285]&~m[1286]&m[1287])|(m[664]&m[1283]&m[1285]&~m[1286]&m[1287])|(~m[664]&m[1283]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[315])|((m[664]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(~m[664]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[664]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[664]&m[1283]&~m[1285]&~m[1286]&m[1287])|(m[664]&~m[1283]&m[1285]&~m[1286]&m[1287])|(~m[664]&~m[1283]&~m[1285]&m[1286]&m[1287])|(m[664]&~m[1283]&~m[1285]&m[1286]&m[1287])|(~m[664]&m[1283]&~m[1285]&m[1286]&m[1287])|(m[664]&m[1283]&~m[1285]&m[1286]&m[1287])|(~m[664]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[664]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[664]&m[1283]&m[1285]&m[1286]&m[1287]))):InitCond[818];
    m[1289] = run?((((m[677]&~m[1288]&~m[1290]&~m[1291]&~m[1292])|(~m[677]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(m[677]&m[1288]&~m[1290]&m[1291]&~m[1292])|(m[677]&~m[1288]&m[1290]&m[1291]&~m[1292])|(~m[677]&m[1288]&~m[1290]&~m[1291]&m[1292])|(~m[677]&~m[1288]&m[1290]&~m[1291]&m[1292])|(m[677]&m[1288]&m[1290]&~m[1291]&m[1292])|(~m[677]&m[1288]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[316])|((m[677]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(~m[677]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[677]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[677]&m[1288]&~m[1290]&~m[1291]&m[1292])|(m[677]&~m[1288]&m[1290]&~m[1291]&m[1292])|(~m[677]&~m[1288]&~m[1290]&m[1291]&m[1292])|(m[677]&~m[1288]&~m[1290]&m[1291]&m[1292])|(~m[677]&m[1288]&~m[1290]&m[1291]&m[1292])|(m[677]&m[1288]&~m[1290]&m[1291]&m[1292])|(~m[677]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[677]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[677]&m[1288]&m[1290]&m[1291]&m[1292]))):InitCond[819];
    m[1294] = run?((((m[690]&~m[1293]&~m[1295]&~m[1296]&~m[1297])|(~m[690]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(m[690]&m[1293]&~m[1295]&m[1296]&~m[1297])|(m[690]&~m[1293]&m[1295]&m[1296]&~m[1297])|(~m[690]&m[1293]&~m[1295]&~m[1296]&m[1297])|(~m[690]&~m[1293]&m[1295]&~m[1296]&m[1297])|(m[690]&m[1293]&m[1295]&~m[1296]&m[1297])|(~m[690]&m[1293]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[317])|((m[690]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(~m[690]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[690]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[690]&m[1293]&~m[1295]&~m[1296]&m[1297])|(m[690]&~m[1293]&m[1295]&~m[1296]&m[1297])|(~m[690]&~m[1293]&~m[1295]&m[1296]&m[1297])|(m[690]&~m[1293]&~m[1295]&m[1296]&m[1297])|(~m[690]&m[1293]&~m[1295]&m[1296]&m[1297])|(m[690]&m[1293]&~m[1295]&m[1296]&m[1297])|(~m[690]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[690]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[690]&m[1293]&m[1295]&m[1296]&m[1297]))):InitCond[820];
    m[1299] = run?((((m[703]&~m[1298]&~m[1300]&~m[1301]&~m[1302])|(~m[703]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(m[703]&m[1298]&~m[1300]&m[1301]&~m[1302])|(m[703]&~m[1298]&m[1300]&m[1301]&~m[1302])|(~m[703]&m[1298]&~m[1300]&~m[1301]&m[1302])|(~m[703]&~m[1298]&m[1300]&~m[1301]&m[1302])|(m[703]&m[1298]&m[1300]&~m[1301]&m[1302])|(~m[703]&m[1298]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[318])|((m[703]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(~m[703]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[703]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[703]&m[1298]&~m[1300]&~m[1301]&m[1302])|(m[703]&~m[1298]&m[1300]&~m[1301]&m[1302])|(~m[703]&~m[1298]&~m[1300]&m[1301]&m[1302])|(m[703]&~m[1298]&~m[1300]&m[1301]&m[1302])|(~m[703]&m[1298]&~m[1300]&m[1301]&m[1302])|(m[703]&m[1298]&~m[1300]&m[1301]&m[1302])|(~m[703]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[703]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[703]&m[1298]&m[1300]&m[1301]&m[1302]))):InitCond[821];
    m[1304] = run?((((m[716]&~m[1303]&~m[1305]&~m[1306]&~m[1307])|(~m[716]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(m[716]&m[1303]&~m[1305]&m[1306]&~m[1307])|(m[716]&~m[1303]&m[1305]&m[1306]&~m[1307])|(~m[716]&m[1303]&~m[1305]&~m[1306]&m[1307])|(~m[716]&~m[1303]&m[1305]&~m[1306]&m[1307])|(m[716]&m[1303]&m[1305]&~m[1306]&m[1307])|(~m[716]&m[1303]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[319])|((m[716]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(~m[716]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[716]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[716]&m[1303]&~m[1305]&~m[1306]&m[1307])|(m[716]&~m[1303]&m[1305]&~m[1306]&m[1307])|(~m[716]&~m[1303]&~m[1305]&m[1306]&m[1307])|(m[716]&~m[1303]&~m[1305]&m[1306]&m[1307])|(~m[716]&m[1303]&~m[1305]&m[1306]&m[1307])|(m[716]&m[1303]&~m[1305]&m[1306]&m[1307])|(~m[716]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[716]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[716]&m[1303]&m[1305]&m[1306]&m[1307]))):InitCond[822];
    m[1309] = run?((((m[587]&~m[1308]&~m[1310]&~m[1311]&~m[1312])|(~m[587]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(m[587]&m[1308]&~m[1310]&m[1311]&~m[1312])|(m[587]&~m[1308]&m[1310]&m[1311]&~m[1312])|(~m[587]&m[1308]&~m[1310]&~m[1311]&m[1312])|(~m[587]&~m[1308]&m[1310]&~m[1311]&m[1312])|(m[587]&m[1308]&m[1310]&~m[1311]&m[1312])|(~m[587]&m[1308]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[320])|((m[587]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(~m[587]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[587]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[587]&m[1308]&~m[1310]&~m[1311]&m[1312])|(m[587]&~m[1308]&m[1310]&~m[1311]&m[1312])|(~m[587]&~m[1308]&~m[1310]&m[1311]&m[1312])|(m[587]&~m[1308]&~m[1310]&m[1311]&m[1312])|(~m[587]&m[1308]&~m[1310]&m[1311]&m[1312])|(m[587]&m[1308]&~m[1310]&m[1311]&m[1312])|(~m[587]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[587]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[587]&m[1308]&m[1310]&m[1311]&m[1312]))):InitCond[823];
    m[1314] = run?((((m[600]&~m[1313]&~m[1315]&~m[1316]&~m[1317])|(~m[600]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(m[600]&m[1313]&~m[1315]&m[1316]&~m[1317])|(m[600]&~m[1313]&m[1315]&m[1316]&~m[1317])|(~m[600]&m[1313]&~m[1315]&~m[1316]&m[1317])|(~m[600]&~m[1313]&m[1315]&~m[1316]&m[1317])|(m[600]&m[1313]&m[1315]&~m[1316]&m[1317])|(~m[600]&m[1313]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[321])|((m[600]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(~m[600]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[600]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[600]&m[1313]&~m[1315]&~m[1316]&m[1317])|(m[600]&~m[1313]&m[1315]&~m[1316]&m[1317])|(~m[600]&~m[1313]&~m[1315]&m[1316]&m[1317])|(m[600]&~m[1313]&~m[1315]&m[1316]&m[1317])|(~m[600]&m[1313]&~m[1315]&m[1316]&m[1317])|(m[600]&m[1313]&~m[1315]&m[1316]&m[1317])|(~m[600]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[600]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[600]&m[1313]&m[1315]&m[1316]&m[1317]))):InitCond[824];
    m[1319] = run?((((m[613]&~m[1318]&~m[1320]&~m[1321]&~m[1322])|(~m[613]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(m[613]&m[1318]&~m[1320]&m[1321]&~m[1322])|(m[613]&~m[1318]&m[1320]&m[1321]&~m[1322])|(~m[613]&m[1318]&~m[1320]&~m[1321]&m[1322])|(~m[613]&~m[1318]&m[1320]&~m[1321]&m[1322])|(m[613]&m[1318]&m[1320]&~m[1321]&m[1322])|(~m[613]&m[1318]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[322])|((m[613]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(~m[613]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[613]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[613]&m[1318]&~m[1320]&~m[1321]&m[1322])|(m[613]&~m[1318]&m[1320]&~m[1321]&m[1322])|(~m[613]&~m[1318]&~m[1320]&m[1321]&m[1322])|(m[613]&~m[1318]&~m[1320]&m[1321]&m[1322])|(~m[613]&m[1318]&~m[1320]&m[1321]&m[1322])|(m[613]&m[1318]&~m[1320]&m[1321]&m[1322])|(~m[613]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[613]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[613]&m[1318]&m[1320]&m[1321]&m[1322]))):InitCond[825];
    m[1324] = run?((((m[626]&~m[1323]&~m[1325]&~m[1326]&~m[1327])|(~m[626]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(m[626]&m[1323]&~m[1325]&m[1326]&~m[1327])|(m[626]&~m[1323]&m[1325]&m[1326]&~m[1327])|(~m[626]&m[1323]&~m[1325]&~m[1326]&m[1327])|(~m[626]&~m[1323]&m[1325]&~m[1326]&m[1327])|(m[626]&m[1323]&m[1325]&~m[1326]&m[1327])|(~m[626]&m[1323]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[323])|((m[626]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(~m[626]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[626]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[626]&m[1323]&~m[1325]&~m[1326]&m[1327])|(m[626]&~m[1323]&m[1325]&~m[1326]&m[1327])|(~m[626]&~m[1323]&~m[1325]&m[1326]&m[1327])|(m[626]&~m[1323]&~m[1325]&m[1326]&m[1327])|(~m[626]&m[1323]&~m[1325]&m[1326]&m[1327])|(m[626]&m[1323]&~m[1325]&m[1326]&m[1327])|(~m[626]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[626]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[626]&m[1323]&m[1325]&m[1326]&m[1327]))):InitCond[826];
    m[1329] = run?((((m[639]&~m[1328]&~m[1330]&~m[1331]&~m[1332])|(~m[639]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(m[639]&m[1328]&~m[1330]&m[1331]&~m[1332])|(m[639]&~m[1328]&m[1330]&m[1331]&~m[1332])|(~m[639]&m[1328]&~m[1330]&~m[1331]&m[1332])|(~m[639]&~m[1328]&m[1330]&~m[1331]&m[1332])|(m[639]&m[1328]&m[1330]&~m[1331]&m[1332])|(~m[639]&m[1328]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[324])|((m[639]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(~m[639]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[639]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[639]&m[1328]&~m[1330]&~m[1331]&m[1332])|(m[639]&~m[1328]&m[1330]&~m[1331]&m[1332])|(~m[639]&~m[1328]&~m[1330]&m[1331]&m[1332])|(m[639]&~m[1328]&~m[1330]&m[1331]&m[1332])|(~m[639]&m[1328]&~m[1330]&m[1331]&m[1332])|(m[639]&m[1328]&~m[1330]&m[1331]&m[1332])|(~m[639]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[639]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[639]&m[1328]&m[1330]&m[1331]&m[1332]))):InitCond[827];
    m[1334] = run?((((m[652]&~m[1333]&~m[1335]&~m[1336]&~m[1337])|(~m[652]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(m[652]&m[1333]&~m[1335]&m[1336]&~m[1337])|(m[652]&~m[1333]&m[1335]&m[1336]&~m[1337])|(~m[652]&m[1333]&~m[1335]&~m[1336]&m[1337])|(~m[652]&~m[1333]&m[1335]&~m[1336]&m[1337])|(m[652]&m[1333]&m[1335]&~m[1336]&m[1337])|(~m[652]&m[1333]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[325])|((m[652]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(~m[652]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[652]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[652]&m[1333]&~m[1335]&~m[1336]&m[1337])|(m[652]&~m[1333]&m[1335]&~m[1336]&m[1337])|(~m[652]&~m[1333]&~m[1335]&m[1336]&m[1337])|(m[652]&~m[1333]&~m[1335]&m[1336]&m[1337])|(~m[652]&m[1333]&~m[1335]&m[1336]&m[1337])|(m[652]&m[1333]&~m[1335]&m[1336]&m[1337])|(~m[652]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[652]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[652]&m[1333]&m[1335]&m[1336]&m[1337]))):InitCond[828];
    m[1339] = run?((((m[665]&~m[1338]&~m[1340]&~m[1341]&~m[1342])|(~m[665]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(m[665]&m[1338]&~m[1340]&m[1341]&~m[1342])|(m[665]&~m[1338]&m[1340]&m[1341]&~m[1342])|(~m[665]&m[1338]&~m[1340]&~m[1341]&m[1342])|(~m[665]&~m[1338]&m[1340]&~m[1341]&m[1342])|(m[665]&m[1338]&m[1340]&~m[1341]&m[1342])|(~m[665]&m[1338]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[326])|((m[665]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(~m[665]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[665]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[665]&m[1338]&~m[1340]&~m[1341]&m[1342])|(m[665]&~m[1338]&m[1340]&~m[1341]&m[1342])|(~m[665]&~m[1338]&~m[1340]&m[1341]&m[1342])|(m[665]&~m[1338]&~m[1340]&m[1341]&m[1342])|(~m[665]&m[1338]&~m[1340]&m[1341]&m[1342])|(m[665]&m[1338]&~m[1340]&m[1341]&m[1342])|(~m[665]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[665]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[665]&m[1338]&m[1340]&m[1341]&m[1342]))):InitCond[829];
    m[1344] = run?((((m[678]&~m[1343]&~m[1345]&~m[1346]&~m[1347])|(~m[678]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(m[678]&m[1343]&~m[1345]&m[1346]&~m[1347])|(m[678]&~m[1343]&m[1345]&m[1346]&~m[1347])|(~m[678]&m[1343]&~m[1345]&~m[1346]&m[1347])|(~m[678]&~m[1343]&m[1345]&~m[1346]&m[1347])|(m[678]&m[1343]&m[1345]&~m[1346]&m[1347])|(~m[678]&m[1343]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[327])|((m[678]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(~m[678]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[678]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[678]&m[1343]&~m[1345]&~m[1346]&m[1347])|(m[678]&~m[1343]&m[1345]&~m[1346]&m[1347])|(~m[678]&~m[1343]&~m[1345]&m[1346]&m[1347])|(m[678]&~m[1343]&~m[1345]&m[1346]&m[1347])|(~m[678]&m[1343]&~m[1345]&m[1346]&m[1347])|(m[678]&m[1343]&~m[1345]&m[1346]&m[1347])|(~m[678]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[678]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[678]&m[1343]&m[1345]&m[1346]&m[1347]))):InitCond[830];
    m[1349] = run?((((m[691]&~m[1348]&~m[1350]&~m[1351]&~m[1352])|(~m[691]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(m[691]&m[1348]&~m[1350]&m[1351]&~m[1352])|(m[691]&~m[1348]&m[1350]&m[1351]&~m[1352])|(~m[691]&m[1348]&~m[1350]&~m[1351]&m[1352])|(~m[691]&~m[1348]&m[1350]&~m[1351]&m[1352])|(m[691]&m[1348]&m[1350]&~m[1351]&m[1352])|(~m[691]&m[1348]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[328])|((m[691]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(~m[691]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[691]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[691]&m[1348]&~m[1350]&~m[1351]&m[1352])|(m[691]&~m[1348]&m[1350]&~m[1351]&m[1352])|(~m[691]&~m[1348]&~m[1350]&m[1351]&m[1352])|(m[691]&~m[1348]&~m[1350]&m[1351]&m[1352])|(~m[691]&m[1348]&~m[1350]&m[1351]&m[1352])|(m[691]&m[1348]&~m[1350]&m[1351]&m[1352])|(~m[691]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[691]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[691]&m[1348]&m[1350]&m[1351]&m[1352]))):InitCond[831];
    m[1354] = run?((((m[704]&~m[1353]&~m[1355]&~m[1356]&~m[1357])|(~m[704]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(m[704]&m[1353]&~m[1355]&m[1356]&~m[1357])|(m[704]&~m[1353]&m[1355]&m[1356]&~m[1357])|(~m[704]&m[1353]&~m[1355]&~m[1356]&m[1357])|(~m[704]&~m[1353]&m[1355]&~m[1356]&m[1357])|(m[704]&m[1353]&m[1355]&~m[1356]&m[1357])|(~m[704]&m[1353]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[329])|((m[704]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(~m[704]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[704]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[704]&m[1353]&~m[1355]&~m[1356]&m[1357])|(m[704]&~m[1353]&m[1355]&~m[1356]&m[1357])|(~m[704]&~m[1353]&~m[1355]&m[1356]&m[1357])|(m[704]&~m[1353]&~m[1355]&m[1356]&m[1357])|(~m[704]&m[1353]&~m[1355]&m[1356]&m[1357])|(m[704]&m[1353]&~m[1355]&m[1356]&m[1357])|(~m[704]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[704]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[704]&m[1353]&m[1355]&m[1356]&m[1357]))):InitCond[832];
    m[1359] = run?((((m[717]&~m[1358]&~m[1360]&~m[1361]&~m[1362])|(~m[717]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(m[717]&m[1358]&~m[1360]&m[1361]&~m[1362])|(m[717]&~m[1358]&m[1360]&m[1361]&~m[1362])|(~m[717]&m[1358]&~m[1360]&~m[1361]&m[1362])|(~m[717]&~m[1358]&m[1360]&~m[1361]&m[1362])|(m[717]&m[1358]&m[1360]&~m[1361]&m[1362])|(~m[717]&m[1358]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[330])|((m[717]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(~m[717]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[717]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[717]&m[1358]&~m[1360]&~m[1361]&m[1362])|(m[717]&~m[1358]&m[1360]&~m[1361]&m[1362])|(~m[717]&~m[1358]&~m[1360]&m[1361]&m[1362])|(m[717]&~m[1358]&~m[1360]&m[1361]&m[1362])|(~m[717]&m[1358]&~m[1360]&m[1361]&m[1362])|(m[717]&m[1358]&~m[1360]&m[1361]&m[1362])|(~m[717]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[717]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[717]&m[1358]&m[1360]&m[1361]&m[1362]))):InitCond[833];
    m[1364] = run?((((m[601]&~m[1363]&~m[1365]&~m[1366]&~m[1367])|(~m[601]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(m[601]&m[1363]&~m[1365]&m[1366]&~m[1367])|(m[601]&~m[1363]&m[1365]&m[1366]&~m[1367])|(~m[601]&m[1363]&~m[1365]&~m[1366]&m[1367])|(~m[601]&~m[1363]&m[1365]&~m[1366]&m[1367])|(m[601]&m[1363]&m[1365]&~m[1366]&m[1367])|(~m[601]&m[1363]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[331])|((m[601]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(~m[601]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[601]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[601]&m[1363]&~m[1365]&~m[1366]&m[1367])|(m[601]&~m[1363]&m[1365]&~m[1366]&m[1367])|(~m[601]&~m[1363]&~m[1365]&m[1366]&m[1367])|(m[601]&~m[1363]&~m[1365]&m[1366]&m[1367])|(~m[601]&m[1363]&~m[1365]&m[1366]&m[1367])|(m[601]&m[1363]&~m[1365]&m[1366]&m[1367])|(~m[601]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[601]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[601]&m[1363]&m[1365]&m[1366]&m[1367]))):InitCond[834];
    m[1369] = run?((((m[614]&~m[1368]&~m[1370]&~m[1371]&~m[1372])|(~m[614]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(m[614]&m[1368]&~m[1370]&m[1371]&~m[1372])|(m[614]&~m[1368]&m[1370]&m[1371]&~m[1372])|(~m[614]&m[1368]&~m[1370]&~m[1371]&m[1372])|(~m[614]&~m[1368]&m[1370]&~m[1371]&m[1372])|(m[614]&m[1368]&m[1370]&~m[1371]&m[1372])|(~m[614]&m[1368]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[332])|((m[614]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(~m[614]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[614]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[614]&m[1368]&~m[1370]&~m[1371]&m[1372])|(m[614]&~m[1368]&m[1370]&~m[1371]&m[1372])|(~m[614]&~m[1368]&~m[1370]&m[1371]&m[1372])|(m[614]&~m[1368]&~m[1370]&m[1371]&m[1372])|(~m[614]&m[1368]&~m[1370]&m[1371]&m[1372])|(m[614]&m[1368]&~m[1370]&m[1371]&m[1372])|(~m[614]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[614]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[614]&m[1368]&m[1370]&m[1371]&m[1372]))):InitCond[835];
    m[1374] = run?((((m[627]&~m[1373]&~m[1375]&~m[1376]&~m[1377])|(~m[627]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(m[627]&m[1373]&~m[1375]&m[1376]&~m[1377])|(m[627]&~m[1373]&m[1375]&m[1376]&~m[1377])|(~m[627]&m[1373]&~m[1375]&~m[1376]&m[1377])|(~m[627]&~m[1373]&m[1375]&~m[1376]&m[1377])|(m[627]&m[1373]&m[1375]&~m[1376]&m[1377])|(~m[627]&m[1373]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[333])|((m[627]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(~m[627]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[627]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[627]&m[1373]&~m[1375]&~m[1376]&m[1377])|(m[627]&~m[1373]&m[1375]&~m[1376]&m[1377])|(~m[627]&~m[1373]&~m[1375]&m[1376]&m[1377])|(m[627]&~m[1373]&~m[1375]&m[1376]&m[1377])|(~m[627]&m[1373]&~m[1375]&m[1376]&m[1377])|(m[627]&m[1373]&~m[1375]&m[1376]&m[1377])|(~m[627]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[627]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[627]&m[1373]&m[1375]&m[1376]&m[1377]))):InitCond[836];
    m[1379] = run?((((m[640]&~m[1378]&~m[1380]&~m[1381]&~m[1382])|(~m[640]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(m[640]&m[1378]&~m[1380]&m[1381]&~m[1382])|(m[640]&~m[1378]&m[1380]&m[1381]&~m[1382])|(~m[640]&m[1378]&~m[1380]&~m[1381]&m[1382])|(~m[640]&~m[1378]&m[1380]&~m[1381]&m[1382])|(m[640]&m[1378]&m[1380]&~m[1381]&m[1382])|(~m[640]&m[1378]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[334])|((m[640]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(~m[640]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[640]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[640]&m[1378]&~m[1380]&~m[1381]&m[1382])|(m[640]&~m[1378]&m[1380]&~m[1381]&m[1382])|(~m[640]&~m[1378]&~m[1380]&m[1381]&m[1382])|(m[640]&~m[1378]&~m[1380]&m[1381]&m[1382])|(~m[640]&m[1378]&~m[1380]&m[1381]&m[1382])|(m[640]&m[1378]&~m[1380]&m[1381]&m[1382])|(~m[640]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[640]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[640]&m[1378]&m[1380]&m[1381]&m[1382]))):InitCond[837];
    m[1384] = run?((((m[653]&~m[1383]&~m[1385]&~m[1386]&~m[1387])|(~m[653]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(m[653]&m[1383]&~m[1385]&m[1386]&~m[1387])|(m[653]&~m[1383]&m[1385]&m[1386]&~m[1387])|(~m[653]&m[1383]&~m[1385]&~m[1386]&m[1387])|(~m[653]&~m[1383]&m[1385]&~m[1386]&m[1387])|(m[653]&m[1383]&m[1385]&~m[1386]&m[1387])|(~m[653]&m[1383]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[335])|((m[653]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(~m[653]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[653]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[653]&m[1383]&~m[1385]&~m[1386]&m[1387])|(m[653]&~m[1383]&m[1385]&~m[1386]&m[1387])|(~m[653]&~m[1383]&~m[1385]&m[1386]&m[1387])|(m[653]&~m[1383]&~m[1385]&m[1386]&m[1387])|(~m[653]&m[1383]&~m[1385]&m[1386]&m[1387])|(m[653]&m[1383]&~m[1385]&m[1386]&m[1387])|(~m[653]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[653]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[653]&m[1383]&m[1385]&m[1386]&m[1387]))):InitCond[838];
    m[1389] = run?((((m[666]&~m[1388]&~m[1390]&~m[1391]&~m[1392])|(~m[666]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(m[666]&m[1388]&~m[1390]&m[1391]&~m[1392])|(m[666]&~m[1388]&m[1390]&m[1391]&~m[1392])|(~m[666]&m[1388]&~m[1390]&~m[1391]&m[1392])|(~m[666]&~m[1388]&m[1390]&~m[1391]&m[1392])|(m[666]&m[1388]&m[1390]&~m[1391]&m[1392])|(~m[666]&m[1388]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[336])|((m[666]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(~m[666]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[666]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[666]&m[1388]&~m[1390]&~m[1391]&m[1392])|(m[666]&~m[1388]&m[1390]&~m[1391]&m[1392])|(~m[666]&~m[1388]&~m[1390]&m[1391]&m[1392])|(m[666]&~m[1388]&~m[1390]&m[1391]&m[1392])|(~m[666]&m[1388]&~m[1390]&m[1391]&m[1392])|(m[666]&m[1388]&~m[1390]&m[1391]&m[1392])|(~m[666]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[666]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[666]&m[1388]&m[1390]&m[1391]&m[1392]))):InitCond[839];
    m[1394] = run?((((m[679]&~m[1393]&~m[1395]&~m[1396]&~m[1397])|(~m[679]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(m[679]&m[1393]&~m[1395]&m[1396]&~m[1397])|(m[679]&~m[1393]&m[1395]&m[1396]&~m[1397])|(~m[679]&m[1393]&~m[1395]&~m[1396]&m[1397])|(~m[679]&~m[1393]&m[1395]&~m[1396]&m[1397])|(m[679]&m[1393]&m[1395]&~m[1396]&m[1397])|(~m[679]&m[1393]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[337])|((m[679]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(~m[679]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[679]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[679]&m[1393]&~m[1395]&~m[1396]&m[1397])|(m[679]&~m[1393]&m[1395]&~m[1396]&m[1397])|(~m[679]&~m[1393]&~m[1395]&m[1396]&m[1397])|(m[679]&~m[1393]&~m[1395]&m[1396]&m[1397])|(~m[679]&m[1393]&~m[1395]&m[1396]&m[1397])|(m[679]&m[1393]&~m[1395]&m[1396]&m[1397])|(~m[679]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[679]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[679]&m[1393]&m[1395]&m[1396]&m[1397]))):InitCond[840];
    m[1399] = run?((((m[692]&~m[1398]&~m[1400]&~m[1401]&~m[1402])|(~m[692]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(m[692]&m[1398]&~m[1400]&m[1401]&~m[1402])|(m[692]&~m[1398]&m[1400]&m[1401]&~m[1402])|(~m[692]&m[1398]&~m[1400]&~m[1401]&m[1402])|(~m[692]&~m[1398]&m[1400]&~m[1401]&m[1402])|(m[692]&m[1398]&m[1400]&~m[1401]&m[1402])|(~m[692]&m[1398]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[338])|((m[692]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(~m[692]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[692]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[692]&m[1398]&~m[1400]&~m[1401]&m[1402])|(m[692]&~m[1398]&m[1400]&~m[1401]&m[1402])|(~m[692]&~m[1398]&~m[1400]&m[1401]&m[1402])|(m[692]&~m[1398]&~m[1400]&m[1401]&m[1402])|(~m[692]&m[1398]&~m[1400]&m[1401]&m[1402])|(m[692]&m[1398]&~m[1400]&m[1401]&m[1402])|(~m[692]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[692]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[692]&m[1398]&m[1400]&m[1401]&m[1402]))):InitCond[841];
    m[1404] = run?((((m[705]&~m[1403]&~m[1405]&~m[1406]&~m[1407])|(~m[705]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(m[705]&m[1403]&~m[1405]&m[1406]&~m[1407])|(m[705]&~m[1403]&m[1405]&m[1406]&~m[1407])|(~m[705]&m[1403]&~m[1405]&~m[1406]&m[1407])|(~m[705]&~m[1403]&m[1405]&~m[1406]&m[1407])|(m[705]&m[1403]&m[1405]&~m[1406]&m[1407])|(~m[705]&m[1403]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[339])|((m[705]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(~m[705]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[705]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[705]&m[1403]&~m[1405]&~m[1406]&m[1407])|(m[705]&~m[1403]&m[1405]&~m[1406]&m[1407])|(~m[705]&~m[1403]&~m[1405]&m[1406]&m[1407])|(m[705]&~m[1403]&~m[1405]&m[1406]&m[1407])|(~m[705]&m[1403]&~m[1405]&m[1406]&m[1407])|(m[705]&m[1403]&~m[1405]&m[1406]&m[1407])|(~m[705]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[705]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[705]&m[1403]&m[1405]&m[1406]&m[1407]))):InitCond[842];
    m[1409] = run?((((m[718]&~m[1408]&~m[1410]&~m[1411]&~m[1412])|(~m[718]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(m[718]&m[1408]&~m[1410]&m[1411]&~m[1412])|(m[718]&~m[1408]&m[1410]&m[1411]&~m[1412])|(~m[718]&m[1408]&~m[1410]&~m[1411]&m[1412])|(~m[718]&~m[1408]&m[1410]&~m[1411]&m[1412])|(m[718]&m[1408]&m[1410]&~m[1411]&m[1412])|(~m[718]&m[1408]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[340])|((m[718]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(~m[718]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[718]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[718]&m[1408]&~m[1410]&~m[1411]&m[1412])|(m[718]&~m[1408]&m[1410]&~m[1411]&m[1412])|(~m[718]&~m[1408]&~m[1410]&m[1411]&m[1412])|(m[718]&~m[1408]&~m[1410]&m[1411]&m[1412])|(~m[718]&m[1408]&~m[1410]&m[1411]&m[1412])|(m[718]&m[1408]&~m[1410]&m[1411]&m[1412])|(~m[718]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[718]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[718]&m[1408]&m[1410]&m[1411]&m[1412]))):InitCond[843];
    m[1414] = run?((((m[615]&~m[1413]&~m[1415]&~m[1416]&~m[1417])|(~m[615]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(m[615]&m[1413]&~m[1415]&m[1416]&~m[1417])|(m[615]&~m[1413]&m[1415]&m[1416]&~m[1417])|(~m[615]&m[1413]&~m[1415]&~m[1416]&m[1417])|(~m[615]&~m[1413]&m[1415]&~m[1416]&m[1417])|(m[615]&m[1413]&m[1415]&~m[1416]&m[1417])|(~m[615]&m[1413]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[341])|((m[615]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(~m[615]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[615]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[615]&m[1413]&~m[1415]&~m[1416]&m[1417])|(m[615]&~m[1413]&m[1415]&~m[1416]&m[1417])|(~m[615]&~m[1413]&~m[1415]&m[1416]&m[1417])|(m[615]&~m[1413]&~m[1415]&m[1416]&m[1417])|(~m[615]&m[1413]&~m[1415]&m[1416]&m[1417])|(m[615]&m[1413]&~m[1415]&m[1416]&m[1417])|(~m[615]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[615]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[615]&m[1413]&m[1415]&m[1416]&m[1417]))):InitCond[844];
    m[1419] = run?((((m[628]&~m[1418]&~m[1420]&~m[1421]&~m[1422])|(~m[628]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(m[628]&m[1418]&~m[1420]&m[1421]&~m[1422])|(m[628]&~m[1418]&m[1420]&m[1421]&~m[1422])|(~m[628]&m[1418]&~m[1420]&~m[1421]&m[1422])|(~m[628]&~m[1418]&m[1420]&~m[1421]&m[1422])|(m[628]&m[1418]&m[1420]&~m[1421]&m[1422])|(~m[628]&m[1418]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[342])|((m[628]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(~m[628]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[628]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[628]&m[1418]&~m[1420]&~m[1421]&m[1422])|(m[628]&~m[1418]&m[1420]&~m[1421]&m[1422])|(~m[628]&~m[1418]&~m[1420]&m[1421]&m[1422])|(m[628]&~m[1418]&~m[1420]&m[1421]&m[1422])|(~m[628]&m[1418]&~m[1420]&m[1421]&m[1422])|(m[628]&m[1418]&~m[1420]&m[1421]&m[1422])|(~m[628]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[628]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[628]&m[1418]&m[1420]&m[1421]&m[1422]))):InitCond[845];
    m[1424] = run?((((m[641]&~m[1423]&~m[1425]&~m[1426]&~m[1427])|(~m[641]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(m[641]&m[1423]&~m[1425]&m[1426]&~m[1427])|(m[641]&~m[1423]&m[1425]&m[1426]&~m[1427])|(~m[641]&m[1423]&~m[1425]&~m[1426]&m[1427])|(~m[641]&~m[1423]&m[1425]&~m[1426]&m[1427])|(m[641]&m[1423]&m[1425]&~m[1426]&m[1427])|(~m[641]&m[1423]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[343])|((m[641]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(~m[641]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[641]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[641]&m[1423]&~m[1425]&~m[1426]&m[1427])|(m[641]&~m[1423]&m[1425]&~m[1426]&m[1427])|(~m[641]&~m[1423]&~m[1425]&m[1426]&m[1427])|(m[641]&~m[1423]&~m[1425]&m[1426]&m[1427])|(~m[641]&m[1423]&~m[1425]&m[1426]&m[1427])|(m[641]&m[1423]&~m[1425]&m[1426]&m[1427])|(~m[641]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[641]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[641]&m[1423]&m[1425]&m[1426]&m[1427]))):InitCond[846];
    m[1429] = run?((((m[654]&~m[1428]&~m[1430]&~m[1431]&~m[1432])|(~m[654]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(m[654]&m[1428]&~m[1430]&m[1431]&~m[1432])|(m[654]&~m[1428]&m[1430]&m[1431]&~m[1432])|(~m[654]&m[1428]&~m[1430]&~m[1431]&m[1432])|(~m[654]&~m[1428]&m[1430]&~m[1431]&m[1432])|(m[654]&m[1428]&m[1430]&~m[1431]&m[1432])|(~m[654]&m[1428]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[344])|((m[654]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(~m[654]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[654]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[654]&m[1428]&~m[1430]&~m[1431]&m[1432])|(m[654]&~m[1428]&m[1430]&~m[1431]&m[1432])|(~m[654]&~m[1428]&~m[1430]&m[1431]&m[1432])|(m[654]&~m[1428]&~m[1430]&m[1431]&m[1432])|(~m[654]&m[1428]&~m[1430]&m[1431]&m[1432])|(m[654]&m[1428]&~m[1430]&m[1431]&m[1432])|(~m[654]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[654]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[654]&m[1428]&m[1430]&m[1431]&m[1432]))):InitCond[847];
    m[1434] = run?((((m[667]&~m[1433]&~m[1435]&~m[1436]&~m[1437])|(~m[667]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(m[667]&m[1433]&~m[1435]&m[1436]&~m[1437])|(m[667]&~m[1433]&m[1435]&m[1436]&~m[1437])|(~m[667]&m[1433]&~m[1435]&~m[1436]&m[1437])|(~m[667]&~m[1433]&m[1435]&~m[1436]&m[1437])|(m[667]&m[1433]&m[1435]&~m[1436]&m[1437])|(~m[667]&m[1433]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[345])|((m[667]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(~m[667]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[667]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[667]&m[1433]&~m[1435]&~m[1436]&m[1437])|(m[667]&~m[1433]&m[1435]&~m[1436]&m[1437])|(~m[667]&~m[1433]&~m[1435]&m[1436]&m[1437])|(m[667]&~m[1433]&~m[1435]&m[1436]&m[1437])|(~m[667]&m[1433]&~m[1435]&m[1436]&m[1437])|(m[667]&m[1433]&~m[1435]&m[1436]&m[1437])|(~m[667]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[667]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[667]&m[1433]&m[1435]&m[1436]&m[1437]))):InitCond[848];
    m[1439] = run?((((m[680]&~m[1438]&~m[1440]&~m[1441]&~m[1442])|(~m[680]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(m[680]&m[1438]&~m[1440]&m[1441]&~m[1442])|(m[680]&~m[1438]&m[1440]&m[1441]&~m[1442])|(~m[680]&m[1438]&~m[1440]&~m[1441]&m[1442])|(~m[680]&~m[1438]&m[1440]&~m[1441]&m[1442])|(m[680]&m[1438]&m[1440]&~m[1441]&m[1442])|(~m[680]&m[1438]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[346])|((m[680]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(~m[680]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[680]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[680]&m[1438]&~m[1440]&~m[1441]&m[1442])|(m[680]&~m[1438]&m[1440]&~m[1441]&m[1442])|(~m[680]&~m[1438]&~m[1440]&m[1441]&m[1442])|(m[680]&~m[1438]&~m[1440]&m[1441]&m[1442])|(~m[680]&m[1438]&~m[1440]&m[1441]&m[1442])|(m[680]&m[1438]&~m[1440]&m[1441]&m[1442])|(~m[680]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[680]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[680]&m[1438]&m[1440]&m[1441]&m[1442]))):InitCond[849];
    m[1444] = run?((((m[693]&~m[1443]&~m[1445]&~m[1446]&~m[1447])|(~m[693]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(m[693]&m[1443]&~m[1445]&m[1446]&~m[1447])|(m[693]&~m[1443]&m[1445]&m[1446]&~m[1447])|(~m[693]&m[1443]&~m[1445]&~m[1446]&m[1447])|(~m[693]&~m[1443]&m[1445]&~m[1446]&m[1447])|(m[693]&m[1443]&m[1445]&~m[1446]&m[1447])|(~m[693]&m[1443]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[347])|((m[693]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(~m[693]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[693]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[693]&m[1443]&~m[1445]&~m[1446]&m[1447])|(m[693]&~m[1443]&m[1445]&~m[1446]&m[1447])|(~m[693]&~m[1443]&~m[1445]&m[1446]&m[1447])|(m[693]&~m[1443]&~m[1445]&m[1446]&m[1447])|(~m[693]&m[1443]&~m[1445]&m[1446]&m[1447])|(m[693]&m[1443]&~m[1445]&m[1446]&m[1447])|(~m[693]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[693]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[693]&m[1443]&m[1445]&m[1446]&m[1447]))):InitCond[850];
    m[1449] = run?((((m[706]&~m[1448]&~m[1450]&~m[1451]&~m[1452])|(~m[706]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(m[706]&m[1448]&~m[1450]&m[1451]&~m[1452])|(m[706]&~m[1448]&m[1450]&m[1451]&~m[1452])|(~m[706]&m[1448]&~m[1450]&~m[1451]&m[1452])|(~m[706]&~m[1448]&m[1450]&~m[1451]&m[1452])|(m[706]&m[1448]&m[1450]&~m[1451]&m[1452])|(~m[706]&m[1448]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[348])|((m[706]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(~m[706]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[706]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[706]&m[1448]&~m[1450]&~m[1451]&m[1452])|(m[706]&~m[1448]&m[1450]&~m[1451]&m[1452])|(~m[706]&~m[1448]&~m[1450]&m[1451]&m[1452])|(m[706]&~m[1448]&~m[1450]&m[1451]&m[1452])|(~m[706]&m[1448]&~m[1450]&m[1451]&m[1452])|(m[706]&m[1448]&~m[1450]&m[1451]&m[1452])|(~m[706]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[706]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[706]&m[1448]&m[1450]&m[1451]&m[1452]))):InitCond[851];
    m[1454] = run?((((m[719]&~m[1453]&~m[1455]&~m[1456]&~m[1457])|(~m[719]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(m[719]&m[1453]&~m[1455]&m[1456]&~m[1457])|(m[719]&~m[1453]&m[1455]&m[1456]&~m[1457])|(~m[719]&m[1453]&~m[1455]&~m[1456]&m[1457])|(~m[719]&~m[1453]&m[1455]&~m[1456]&m[1457])|(m[719]&m[1453]&m[1455]&~m[1456]&m[1457])|(~m[719]&m[1453]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[349])|((m[719]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(~m[719]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[719]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[719]&m[1453]&~m[1455]&~m[1456]&m[1457])|(m[719]&~m[1453]&m[1455]&~m[1456]&m[1457])|(~m[719]&~m[1453]&~m[1455]&m[1456]&m[1457])|(m[719]&~m[1453]&~m[1455]&m[1456]&m[1457])|(~m[719]&m[1453]&~m[1455]&m[1456]&m[1457])|(m[719]&m[1453]&~m[1455]&m[1456]&m[1457])|(~m[719]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[719]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[719]&m[1453]&m[1455]&m[1456]&m[1457]))):InitCond[852];
    m[1459] = run?((((m[629]&~m[1458]&~m[1460]&~m[1461]&~m[1462])|(~m[629]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(m[629]&m[1458]&~m[1460]&m[1461]&~m[1462])|(m[629]&~m[1458]&m[1460]&m[1461]&~m[1462])|(~m[629]&m[1458]&~m[1460]&~m[1461]&m[1462])|(~m[629]&~m[1458]&m[1460]&~m[1461]&m[1462])|(m[629]&m[1458]&m[1460]&~m[1461]&m[1462])|(~m[629]&m[1458]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[350])|((m[629]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(~m[629]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[629]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[629]&m[1458]&~m[1460]&~m[1461]&m[1462])|(m[629]&~m[1458]&m[1460]&~m[1461]&m[1462])|(~m[629]&~m[1458]&~m[1460]&m[1461]&m[1462])|(m[629]&~m[1458]&~m[1460]&m[1461]&m[1462])|(~m[629]&m[1458]&~m[1460]&m[1461]&m[1462])|(m[629]&m[1458]&~m[1460]&m[1461]&m[1462])|(~m[629]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[629]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[629]&m[1458]&m[1460]&m[1461]&m[1462]))):InitCond[853];
    m[1464] = run?((((m[642]&~m[1463]&~m[1465]&~m[1466]&~m[1467])|(~m[642]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(m[642]&m[1463]&~m[1465]&m[1466]&~m[1467])|(m[642]&~m[1463]&m[1465]&m[1466]&~m[1467])|(~m[642]&m[1463]&~m[1465]&~m[1466]&m[1467])|(~m[642]&~m[1463]&m[1465]&~m[1466]&m[1467])|(m[642]&m[1463]&m[1465]&~m[1466]&m[1467])|(~m[642]&m[1463]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[351])|((m[642]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(~m[642]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[642]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[642]&m[1463]&~m[1465]&~m[1466]&m[1467])|(m[642]&~m[1463]&m[1465]&~m[1466]&m[1467])|(~m[642]&~m[1463]&~m[1465]&m[1466]&m[1467])|(m[642]&~m[1463]&~m[1465]&m[1466]&m[1467])|(~m[642]&m[1463]&~m[1465]&m[1466]&m[1467])|(m[642]&m[1463]&~m[1465]&m[1466]&m[1467])|(~m[642]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[642]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[642]&m[1463]&m[1465]&m[1466]&m[1467]))):InitCond[854];
    m[1469] = run?((((m[655]&~m[1468]&~m[1470]&~m[1471]&~m[1472])|(~m[655]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(m[655]&m[1468]&~m[1470]&m[1471]&~m[1472])|(m[655]&~m[1468]&m[1470]&m[1471]&~m[1472])|(~m[655]&m[1468]&~m[1470]&~m[1471]&m[1472])|(~m[655]&~m[1468]&m[1470]&~m[1471]&m[1472])|(m[655]&m[1468]&m[1470]&~m[1471]&m[1472])|(~m[655]&m[1468]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[352])|((m[655]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(~m[655]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[655]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[655]&m[1468]&~m[1470]&~m[1471]&m[1472])|(m[655]&~m[1468]&m[1470]&~m[1471]&m[1472])|(~m[655]&~m[1468]&~m[1470]&m[1471]&m[1472])|(m[655]&~m[1468]&~m[1470]&m[1471]&m[1472])|(~m[655]&m[1468]&~m[1470]&m[1471]&m[1472])|(m[655]&m[1468]&~m[1470]&m[1471]&m[1472])|(~m[655]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[655]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[655]&m[1468]&m[1470]&m[1471]&m[1472]))):InitCond[855];
    m[1474] = run?((((m[668]&~m[1473]&~m[1475]&~m[1476]&~m[1477])|(~m[668]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(m[668]&m[1473]&~m[1475]&m[1476]&~m[1477])|(m[668]&~m[1473]&m[1475]&m[1476]&~m[1477])|(~m[668]&m[1473]&~m[1475]&~m[1476]&m[1477])|(~m[668]&~m[1473]&m[1475]&~m[1476]&m[1477])|(m[668]&m[1473]&m[1475]&~m[1476]&m[1477])|(~m[668]&m[1473]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[353])|((m[668]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(~m[668]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[668]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[668]&m[1473]&~m[1475]&~m[1476]&m[1477])|(m[668]&~m[1473]&m[1475]&~m[1476]&m[1477])|(~m[668]&~m[1473]&~m[1475]&m[1476]&m[1477])|(m[668]&~m[1473]&~m[1475]&m[1476]&m[1477])|(~m[668]&m[1473]&~m[1475]&m[1476]&m[1477])|(m[668]&m[1473]&~m[1475]&m[1476]&m[1477])|(~m[668]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[668]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[668]&m[1473]&m[1475]&m[1476]&m[1477]))):InitCond[856];
    m[1479] = run?((((m[681]&~m[1478]&~m[1480]&~m[1481]&~m[1482])|(~m[681]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(m[681]&m[1478]&~m[1480]&m[1481]&~m[1482])|(m[681]&~m[1478]&m[1480]&m[1481]&~m[1482])|(~m[681]&m[1478]&~m[1480]&~m[1481]&m[1482])|(~m[681]&~m[1478]&m[1480]&~m[1481]&m[1482])|(m[681]&m[1478]&m[1480]&~m[1481]&m[1482])|(~m[681]&m[1478]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[354])|((m[681]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(~m[681]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[681]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[681]&m[1478]&~m[1480]&~m[1481]&m[1482])|(m[681]&~m[1478]&m[1480]&~m[1481]&m[1482])|(~m[681]&~m[1478]&~m[1480]&m[1481]&m[1482])|(m[681]&~m[1478]&~m[1480]&m[1481]&m[1482])|(~m[681]&m[1478]&~m[1480]&m[1481]&m[1482])|(m[681]&m[1478]&~m[1480]&m[1481]&m[1482])|(~m[681]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[681]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[681]&m[1478]&m[1480]&m[1481]&m[1482]))):InitCond[857];
    m[1484] = run?((((m[694]&~m[1483]&~m[1485]&~m[1486]&~m[1487])|(~m[694]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(m[694]&m[1483]&~m[1485]&m[1486]&~m[1487])|(m[694]&~m[1483]&m[1485]&m[1486]&~m[1487])|(~m[694]&m[1483]&~m[1485]&~m[1486]&m[1487])|(~m[694]&~m[1483]&m[1485]&~m[1486]&m[1487])|(m[694]&m[1483]&m[1485]&~m[1486]&m[1487])|(~m[694]&m[1483]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[355])|((m[694]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(~m[694]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[694]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[694]&m[1483]&~m[1485]&~m[1486]&m[1487])|(m[694]&~m[1483]&m[1485]&~m[1486]&m[1487])|(~m[694]&~m[1483]&~m[1485]&m[1486]&m[1487])|(m[694]&~m[1483]&~m[1485]&m[1486]&m[1487])|(~m[694]&m[1483]&~m[1485]&m[1486]&m[1487])|(m[694]&m[1483]&~m[1485]&m[1486]&m[1487])|(~m[694]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[694]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[694]&m[1483]&m[1485]&m[1486]&m[1487]))):InitCond[858];
    m[1489] = run?((((m[707]&~m[1488]&~m[1490]&~m[1491]&~m[1492])|(~m[707]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(m[707]&m[1488]&~m[1490]&m[1491]&~m[1492])|(m[707]&~m[1488]&m[1490]&m[1491]&~m[1492])|(~m[707]&m[1488]&~m[1490]&~m[1491]&m[1492])|(~m[707]&~m[1488]&m[1490]&~m[1491]&m[1492])|(m[707]&m[1488]&m[1490]&~m[1491]&m[1492])|(~m[707]&m[1488]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[356])|((m[707]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(~m[707]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[707]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[707]&m[1488]&~m[1490]&~m[1491]&m[1492])|(m[707]&~m[1488]&m[1490]&~m[1491]&m[1492])|(~m[707]&~m[1488]&~m[1490]&m[1491]&m[1492])|(m[707]&~m[1488]&~m[1490]&m[1491]&m[1492])|(~m[707]&m[1488]&~m[1490]&m[1491]&m[1492])|(m[707]&m[1488]&~m[1490]&m[1491]&m[1492])|(~m[707]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[707]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[707]&m[1488]&m[1490]&m[1491]&m[1492]))):InitCond[859];
    m[1494] = run?((((m[720]&~m[1493]&~m[1495]&~m[1496]&~m[1497])|(~m[720]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(m[720]&m[1493]&~m[1495]&m[1496]&~m[1497])|(m[720]&~m[1493]&m[1495]&m[1496]&~m[1497])|(~m[720]&m[1493]&~m[1495]&~m[1496]&m[1497])|(~m[720]&~m[1493]&m[1495]&~m[1496]&m[1497])|(m[720]&m[1493]&m[1495]&~m[1496]&m[1497])|(~m[720]&m[1493]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[357])|((m[720]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(~m[720]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[720]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[720]&m[1493]&~m[1495]&~m[1496]&m[1497])|(m[720]&~m[1493]&m[1495]&~m[1496]&m[1497])|(~m[720]&~m[1493]&~m[1495]&m[1496]&m[1497])|(m[720]&~m[1493]&~m[1495]&m[1496]&m[1497])|(~m[720]&m[1493]&~m[1495]&m[1496]&m[1497])|(m[720]&m[1493]&~m[1495]&m[1496]&m[1497])|(~m[720]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[720]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[720]&m[1493]&m[1495]&m[1496]&m[1497]))):InitCond[860];
    m[1499] = run?((((m[643]&~m[1498]&~m[1500]&~m[1501]&~m[1502])|(~m[643]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(m[643]&m[1498]&~m[1500]&m[1501]&~m[1502])|(m[643]&~m[1498]&m[1500]&m[1501]&~m[1502])|(~m[643]&m[1498]&~m[1500]&~m[1501]&m[1502])|(~m[643]&~m[1498]&m[1500]&~m[1501]&m[1502])|(m[643]&m[1498]&m[1500]&~m[1501]&m[1502])|(~m[643]&m[1498]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[358])|((m[643]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(~m[643]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[643]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[643]&m[1498]&~m[1500]&~m[1501]&m[1502])|(m[643]&~m[1498]&m[1500]&~m[1501]&m[1502])|(~m[643]&~m[1498]&~m[1500]&m[1501]&m[1502])|(m[643]&~m[1498]&~m[1500]&m[1501]&m[1502])|(~m[643]&m[1498]&~m[1500]&m[1501]&m[1502])|(m[643]&m[1498]&~m[1500]&m[1501]&m[1502])|(~m[643]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[643]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[643]&m[1498]&m[1500]&m[1501]&m[1502]))):InitCond[861];
    m[1504] = run?((((m[656]&~m[1503]&~m[1505]&~m[1506]&~m[1507])|(~m[656]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(m[656]&m[1503]&~m[1505]&m[1506]&~m[1507])|(m[656]&~m[1503]&m[1505]&m[1506]&~m[1507])|(~m[656]&m[1503]&~m[1505]&~m[1506]&m[1507])|(~m[656]&~m[1503]&m[1505]&~m[1506]&m[1507])|(m[656]&m[1503]&m[1505]&~m[1506]&m[1507])|(~m[656]&m[1503]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[359])|((m[656]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(~m[656]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[656]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[656]&m[1503]&~m[1505]&~m[1506]&m[1507])|(m[656]&~m[1503]&m[1505]&~m[1506]&m[1507])|(~m[656]&~m[1503]&~m[1505]&m[1506]&m[1507])|(m[656]&~m[1503]&~m[1505]&m[1506]&m[1507])|(~m[656]&m[1503]&~m[1505]&m[1506]&m[1507])|(m[656]&m[1503]&~m[1505]&m[1506]&m[1507])|(~m[656]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[656]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[656]&m[1503]&m[1505]&m[1506]&m[1507]))):InitCond[862];
    m[1509] = run?((((m[669]&~m[1508]&~m[1510]&~m[1511]&~m[1512])|(~m[669]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(m[669]&m[1508]&~m[1510]&m[1511]&~m[1512])|(m[669]&~m[1508]&m[1510]&m[1511]&~m[1512])|(~m[669]&m[1508]&~m[1510]&~m[1511]&m[1512])|(~m[669]&~m[1508]&m[1510]&~m[1511]&m[1512])|(m[669]&m[1508]&m[1510]&~m[1511]&m[1512])|(~m[669]&m[1508]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[360])|((m[669]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(~m[669]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[669]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[669]&m[1508]&~m[1510]&~m[1511]&m[1512])|(m[669]&~m[1508]&m[1510]&~m[1511]&m[1512])|(~m[669]&~m[1508]&~m[1510]&m[1511]&m[1512])|(m[669]&~m[1508]&~m[1510]&m[1511]&m[1512])|(~m[669]&m[1508]&~m[1510]&m[1511]&m[1512])|(m[669]&m[1508]&~m[1510]&m[1511]&m[1512])|(~m[669]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[669]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[669]&m[1508]&m[1510]&m[1511]&m[1512]))):InitCond[863];
    m[1514] = run?((((m[682]&~m[1513]&~m[1515]&~m[1516]&~m[1517])|(~m[682]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(m[682]&m[1513]&~m[1515]&m[1516]&~m[1517])|(m[682]&~m[1513]&m[1515]&m[1516]&~m[1517])|(~m[682]&m[1513]&~m[1515]&~m[1516]&m[1517])|(~m[682]&~m[1513]&m[1515]&~m[1516]&m[1517])|(m[682]&m[1513]&m[1515]&~m[1516]&m[1517])|(~m[682]&m[1513]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[361])|((m[682]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(~m[682]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[682]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[682]&m[1513]&~m[1515]&~m[1516]&m[1517])|(m[682]&~m[1513]&m[1515]&~m[1516]&m[1517])|(~m[682]&~m[1513]&~m[1515]&m[1516]&m[1517])|(m[682]&~m[1513]&~m[1515]&m[1516]&m[1517])|(~m[682]&m[1513]&~m[1515]&m[1516]&m[1517])|(m[682]&m[1513]&~m[1515]&m[1516]&m[1517])|(~m[682]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[682]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[682]&m[1513]&m[1515]&m[1516]&m[1517]))):InitCond[864];
    m[1519] = run?((((m[695]&~m[1518]&~m[1520]&~m[1521]&~m[1522])|(~m[695]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(m[695]&m[1518]&~m[1520]&m[1521]&~m[1522])|(m[695]&~m[1518]&m[1520]&m[1521]&~m[1522])|(~m[695]&m[1518]&~m[1520]&~m[1521]&m[1522])|(~m[695]&~m[1518]&m[1520]&~m[1521]&m[1522])|(m[695]&m[1518]&m[1520]&~m[1521]&m[1522])|(~m[695]&m[1518]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[362])|((m[695]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(~m[695]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[695]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[695]&m[1518]&~m[1520]&~m[1521]&m[1522])|(m[695]&~m[1518]&m[1520]&~m[1521]&m[1522])|(~m[695]&~m[1518]&~m[1520]&m[1521]&m[1522])|(m[695]&~m[1518]&~m[1520]&m[1521]&m[1522])|(~m[695]&m[1518]&~m[1520]&m[1521]&m[1522])|(m[695]&m[1518]&~m[1520]&m[1521]&m[1522])|(~m[695]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[695]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[695]&m[1518]&m[1520]&m[1521]&m[1522]))):InitCond[865];
    m[1524] = run?((((m[708]&~m[1523]&~m[1525]&~m[1526]&~m[1527])|(~m[708]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(m[708]&m[1523]&~m[1525]&m[1526]&~m[1527])|(m[708]&~m[1523]&m[1525]&m[1526]&~m[1527])|(~m[708]&m[1523]&~m[1525]&~m[1526]&m[1527])|(~m[708]&~m[1523]&m[1525]&~m[1526]&m[1527])|(m[708]&m[1523]&m[1525]&~m[1526]&m[1527])|(~m[708]&m[1523]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[363])|((m[708]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(~m[708]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[708]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[708]&m[1523]&~m[1525]&~m[1526]&m[1527])|(m[708]&~m[1523]&m[1525]&~m[1526]&m[1527])|(~m[708]&~m[1523]&~m[1525]&m[1526]&m[1527])|(m[708]&~m[1523]&~m[1525]&m[1526]&m[1527])|(~m[708]&m[1523]&~m[1525]&m[1526]&m[1527])|(m[708]&m[1523]&~m[1525]&m[1526]&m[1527])|(~m[708]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[708]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[708]&m[1523]&m[1525]&m[1526]&m[1527]))):InitCond[866];
    m[1529] = run?((((m[721]&~m[1528]&~m[1530]&~m[1531]&~m[1532])|(~m[721]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(m[721]&m[1528]&~m[1530]&m[1531]&~m[1532])|(m[721]&~m[1528]&m[1530]&m[1531]&~m[1532])|(~m[721]&m[1528]&~m[1530]&~m[1531]&m[1532])|(~m[721]&~m[1528]&m[1530]&~m[1531]&m[1532])|(m[721]&m[1528]&m[1530]&~m[1531]&m[1532])|(~m[721]&m[1528]&m[1530]&m[1531]&m[1532]))&UnbiasedRNG[364])|((m[721]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(~m[721]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[721]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[721]&m[1528]&~m[1530]&~m[1531]&m[1532])|(m[721]&~m[1528]&m[1530]&~m[1531]&m[1532])|(~m[721]&~m[1528]&~m[1530]&m[1531]&m[1532])|(m[721]&~m[1528]&~m[1530]&m[1531]&m[1532])|(~m[721]&m[1528]&~m[1530]&m[1531]&m[1532])|(m[721]&m[1528]&~m[1530]&m[1531]&m[1532])|(~m[721]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[721]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[721]&m[1528]&m[1530]&m[1531]&m[1532]))):InitCond[867];
    m[1534] = run?((((m[657]&~m[1533]&~m[1535]&~m[1536]&~m[1537])|(~m[657]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(m[657]&m[1533]&~m[1535]&m[1536]&~m[1537])|(m[657]&~m[1533]&m[1535]&m[1536]&~m[1537])|(~m[657]&m[1533]&~m[1535]&~m[1536]&m[1537])|(~m[657]&~m[1533]&m[1535]&~m[1536]&m[1537])|(m[657]&m[1533]&m[1535]&~m[1536]&m[1537])|(~m[657]&m[1533]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[365])|((m[657]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(~m[657]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[657]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[657]&m[1533]&~m[1535]&~m[1536]&m[1537])|(m[657]&~m[1533]&m[1535]&~m[1536]&m[1537])|(~m[657]&~m[1533]&~m[1535]&m[1536]&m[1537])|(m[657]&~m[1533]&~m[1535]&m[1536]&m[1537])|(~m[657]&m[1533]&~m[1535]&m[1536]&m[1537])|(m[657]&m[1533]&~m[1535]&m[1536]&m[1537])|(~m[657]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[657]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[657]&m[1533]&m[1535]&m[1536]&m[1537]))):InitCond[868];
    m[1539] = run?((((m[670]&~m[1538]&~m[1540]&~m[1541]&~m[1542])|(~m[670]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(m[670]&m[1538]&~m[1540]&m[1541]&~m[1542])|(m[670]&~m[1538]&m[1540]&m[1541]&~m[1542])|(~m[670]&m[1538]&~m[1540]&~m[1541]&m[1542])|(~m[670]&~m[1538]&m[1540]&~m[1541]&m[1542])|(m[670]&m[1538]&m[1540]&~m[1541]&m[1542])|(~m[670]&m[1538]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[366])|((m[670]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(~m[670]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[670]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[670]&m[1538]&~m[1540]&~m[1541]&m[1542])|(m[670]&~m[1538]&m[1540]&~m[1541]&m[1542])|(~m[670]&~m[1538]&~m[1540]&m[1541]&m[1542])|(m[670]&~m[1538]&~m[1540]&m[1541]&m[1542])|(~m[670]&m[1538]&~m[1540]&m[1541]&m[1542])|(m[670]&m[1538]&~m[1540]&m[1541]&m[1542])|(~m[670]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[670]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[670]&m[1538]&m[1540]&m[1541]&m[1542]))):InitCond[869];
    m[1544] = run?((((m[683]&~m[1543]&~m[1545]&~m[1546]&~m[1547])|(~m[683]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(m[683]&m[1543]&~m[1545]&m[1546]&~m[1547])|(m[683]&~m[1543]&m[1545]&m[1546]&~m[1547])|(~m[683]&m[1543]&~m[1545]&~m[1546]&m[1547])|(~m[683]&~m[1543]&m[1545]&~m[1546]&m[1547])|(m[683]&m[1543]&m[1545]&~m[1546]&m[1547])|(~m[683]&m[1543]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[367])|((m[683]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(~m[683]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[683]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[683]&m[1543]&~m[1545]&~m[1546]&m[1547])|(m[683]&~m[1543]&m[1545]&~m[1546]&m[1547])|(~m[683]&~m[1543]&~m[1545]&m[1546]&m[1547])|(m[683]&~m[1543]&~m[1545]&m[1546]&m[1547])|(~m[683]&m[1543]&~m[1545]&m[1546]&m[1547])|(m[683]&m[1543]&~m[1545]&m[1546]&m[1547])|(~m[683]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[683]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[683]&m[1543]&m[1545]&m[1546]&m[1547]))):InitCond[870];
    m[1549] = run?((((m[696]&~m[1548]&~m[1550]&~m[1551]&~m[1552])|(~m[696]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(m[696]&m[1548]&~m[1550]&m[1551]&~m[1552])|(m[696]&~m[1548]&m[1550]&m[1551]&~m[1552])|(~m[696]&m[1548]&~m[1550]&~m[1551]&m[1552])|(~m[696]&~m[1548]&m[1550]&~m[1551]&m[1552])|(m[696]&m[1548]&m[1550]&~m[1551]&m[1552])|(~m[696]&m[1548]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[368])|((m[696]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(~m[696]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[696]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[696]&m[1548]&~m[1550]&~m[1551]&m[1552])|(m[696]&~m[1548]&m[1550]&~m[1551]&m[1552])|(~m[696]&~m[1548]&~m[1550]&m[1551]&m[1552])|(m[696]&~m[1548]&~m[1550]&m[1551]&m[1552])|(~m[696]&m[1548]&~m[1550]&m[1551]&m[1552])|(m[696]&m[1548]&~m[1550]&m[1551]&m[1552])|(~m[696]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[696]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[696]&m[1548]&m[1550]&m[1551]&m[1552]))):InitCond[871];
    m[1554] = run?((((m[709]&~m[1553]&~m[1555]&~m[1556]&~m[1557])|(~m[709]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(m[709]&m[1553]&~m[1555]&m[1556]&~m[1557])|(m[709]&~m[1553]&m[1555]&m[1556]&~m[1557])|(~m[709]&m[1553]&~m[1555]&~m[1556]&m[1557])|(~m[709]&~m[1553]&m[1555]&~m[1556]&m[1557])|(m[709]&m[1553]&m[1555]&~m[1556]&m[1557])|(~m[709]&m[1553]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[369])|((m[709]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(~m[709]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[709]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[709]&m[1553]&~m[1555]&~m[1556]&m[1557])|(m[709]&~m[1553]&m[1555]&~m[1556]&m[1557])|(~m[709]&~m[1553]&~m[1555]&m[1556]&m[1557])|(m[709]&~m[1553]&~m[1555]&m[1556]&m[1557])|(~m[709]&m[1553]&~m[1555]&m[1556]&m[1557])|(m[709]&m[1553]&~m[1555]&m[1556]&m[1557])|(~m[709]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[709]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[709]&m[1553]&m[1555]&m[1556]&m[1557]))):InitCond[872];
    m[1559] = run?((((m[722]&~m[1558]&~m[1560]&~m[1561]&~m[1562])|(~m[722]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(m[722]&m[1558]&~m[1560]&m[1561]&~m[1562])|(m[722]&~m[1558]&m[1560]&m[1561]&~m[1562])|(~m[722]&m[1558]&~m[1560]&~m[1561]&m[1562])|(~m[722]&~m[1558]&m[1560]&~m[1561]&m[1562])|(m[722]&m[1558]&m[1560]&~m[1561]&m[1562])|(~m[722]&m[1558]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[370])|((m[722]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(~m[722]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[722]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[722]&m[1558]&~m[1560]&~m[1561]&m[1562])|(m[722]&~m[1558]&m[1560]&~m[1561]&m[1562])|(~m[722]&~m[1558]&~m[1560]&m[1561]&m[1562])|(m[722]&~m[1558]&~m[1560]&m[1561]&m[1562])|(~m[722]&m[1558]&~m[1560]&m[1561]&m[1562])|(m[722]&m[1558]&~m[1560]&m[1561]&m[1562])|(~m[722]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[722]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[722]&m[1558]&m[1560]&m[1561]&m[1562]))):InitCond[873];
    m[1564] = run?((((m[671]&~m[1563]&~m[1565]&~m[1566]&~m[1567])|(~m[671]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(m[671]&m[1563]&~m[1565]&m[1566]&~m[1567])|(m[671]&~m[1563]&m[1565]&m[1566]&~m[1567])|(~m[671]&m[1563]&~m[1565]&~m[1566]&m[1567])|(~m[671]&~m[1563]&m[1565]&~m[1566]&m[1567])|(m[671]&m[1563]&m[1565]&~m[1566]&m[1567])|(~m[671]&m[1563]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[371])|((m[671]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(~m[671]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[671]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[671]&m[1563]&~m[1565]&~m[1566]&m[1567])|(m[671]&~m[1563]&m[1565]&~m[1566]&m[1567])|(~m[671]&~m[1563]&~m[1565]&m[1566]&m[1567])|(m[671]&~m[1563]&~m[1565]&m[1566]&m[1567])|(~m[671]&m[1563]&~m[1565]&m[1566]&m[1567])|(m[671]&m[1563]&~m[1565]&m[1566]&m[1567])|(~m[671]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[671]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[671]&m[1563]&m[1565]&m[1566]&m[1567]))):InitCond[874];
    m[1569] = run?((((m[684]&~m[1568]&~m[1570]&~m[1571]&~m[1572])|(~m[684]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(m[684]&m[1568]&~m[1570]&m[1571]&~m[1572])|(m[684]&~m[1568]&m[1570]&m[1571]&~m[1572])|(~m[684]&m[1568]&~m[1570]&~m[1571]&m[1572])|(~m[684]&~m[1568]&m[1570]&~m[1571]&m[1572])|(m[684]&m[1568]&m[1570]&~m[1571]&m[1572])|(~m[684]&m[1568]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[372])|((m[684]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(~m[684]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[684]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[684]&m[1568]&~m[1570]&~m[1571]&m[1572])|(m[684]&~m[1568]&m[1570]&~m[1571]&m[1572])|(~m[684]&~m[1568]&~m[1570]&m[1571]&m[1572])|(m[684]&~m[1568]&~m[1570]&m[1571]&m[1572])|(~m[684]&m[1568]&~m[1570]&m[1571]&m[1572])|(m[684]&m[1568]&~m[1570]&m[1571]&m[1572])|(~m[684]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[684]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[684]&m[1568]&m[1570]&m[1571]&m[1572]))):InitCond[875];
    m[1574] = run?((((m[697]&~m[1573]&~m[1575]&~m[1576]&~m[1577])|(~m[697]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(m[697]&m[1573]&~m[1575]&m[1576]&~m[1577])|(m[697]&~m[1573]&m[1575]&m[1576]&~m[1577])|(~m[697]&m[1573]&~m[1575]&~m[1576]&m[1577])|(~m[697]&~m[1573]&m[1575]&~m[1576]&m[1577])|(m[697]&m[1573]&m[1575]&~m[1576]&m[1577])|(~m[697]&m[1573]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[373])|((m[697]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(~m[697]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[697]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[697]&m[1573]&~m[1575]&~m[1576]&m[1577])|(m[697]&~m[1573]&m[1575]&~m[1576]&m[1577])|(~m[697]&~m[1573]&~m[1575]&m[1576]&m[1577])|(m[697]&~m[1573]&~m[1575]&m[1576]&m[1577])|(~m[697]&m[1573]&~m[1575]&m[1576]&m[1577])|(m[697]&m[1573]&~m[1575]&m[1576]&m[1577])|(~m[697]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[697]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[697]&m[1573]&m[1575]&m[1576]&m[1577]))):InitCond[876];
    m[1579] = run?((((m[710]&~m[1578]&~m[1580]&~m[1581]&~m[1582])|(~m[710]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(m[710]&m[1578]&~m[1580]&m[1581]&~m[1582])|(m[710]&~m[1578]&m[1580]&m[1581]&~m[1582])|(~m[710]&m[1578]&~m[1580]&~m[1581]&m[1582])|(~m[710]&~m[1578]&m[1580]&~m[1581]&m[1582])|(m[710]&m[1578]&m[1580]&~m[1581]&m[1582])|(~m[710]&m[1578]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[374])|((m[710]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(~m[710]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[710]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[710]&m[1578]&~m[1580]&~m[1581]&m[1582])|(m[710]&~m[1578]&m[1580]&~m[1581]&m[1582])|(~m[710]&~m[1578]&~m[1580]&m[1581]&m[1582])|(m[710]&~m[1578]&~m[1580]&m[1581]&m[1582])|(~m[710]&m[1578]&~m[1580]&m[1581]&m[1582])|(m[710]&m[1578]&~m[1580]&m[1581]&m[1582])|(~m[710]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[710]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[710]&m[1578]&m[1580]&m[1581]&m[1582]))):InitCond[877];
    m[1584] = run?((((m[723]&~m[1583]&~m[1585]&~m[1586]&~m[1587])|(~m[723]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(m[723]&m[1583]&~m[1585]&m[1586]&~m[1587])|(m[723]&~m[1583]&m[1585]&m[1586]&~m[1587])|(~m[723]&m[1583]&~m[1585]&~m[1586]&m[1587])|(~m[723]&~m[1583]&m[1585]&~m[1586]&m[1587])|(m[723]&m[1583]&m[1585]&~m[1586]&m[1587])|(~m[723]&m[1583]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[375])|((m[723]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(~m[723]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[723]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[723]&m[1583]&~m[1585]&~m[1586]&m[1587])|(m[723]&~m[1583]&m[1585]&~m[1586]&m[1587])|(~m[723]&~m[1583]&~m[1585]&m[1586]&m[1587])|(m[723]&~m[1583]&~m[1585]&m[1586]&m[1587])|(~m[723]&m[1583]&~m[1585]&m[1586]&m[1587])|(m[723]&m[1583]&~m[1585]&m[1586]&m[1587])|(~m[723]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[723]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[723]&m[1583]&m[1585]&m[1586]&m[1587]))):InitCond[878];
    m[1589] = run?((((m[685]&~m[1588]&~m[1590]&~m[1591]&~m[1592])|(~m[685]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(m[685]&m[1588]&~m[1590]&m[1591]&~m[1592])|(m[685]&~m[1588]&m[1590]&m[1591]&~m[1592])|(~m[685]&m[1588]&~m[1590]&~m[1591]&m[1592])|(~m[685]&~m[1588]&m[1590]&~m[1591]&m[1592])|(m[685]&m[1588]&m[1590]&~m[1591]&m[1592])|(~m[685]&m[1588]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[376])|((m[685]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(~m[685]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[685]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[685]&m[1588]&~m[1590]&~m[1591]&m[1592])|(m[685]&~m[1588]&m[1590]&~m[1591]&m[1592])|(~m[685]&~m[1588]&~m[1590]&m[1591]&m[1592])|(m[685]&~m[1588]&~m[1590]&m[1591]&m[1592])|(~m[685]&m[1588]&~m[1590]&m[1591]&m[1592])|(m[685]&m[1588]&~m[1590]&m[1591]&m[1592])|(~m[685]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[685]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[685]&m[1588]&m[1590]&m[1591]&m[1592]))):InitCond[879];
    m[1594] = run?((((m[698]&~m[1593]&~m[1595]&~m[1596]&~m[1597])|(~m[698]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(m[698]&m[1593]&~m[1595]&m[1596]&~m[1597])|(m[698]&~m[1593]&m[1595]&m[1596]&~m[1597])|(~m[698]&m[1593]&~m[1595]&~m[1596]&m[1597])|(~m[698]&~m[1593]&m[1595]&~m[1596]&m[1597])|(m[698]&m[1593]&m[1595]&~m[1596]&m[1597])|(~m[698]&m[1593]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[377])|((m[698]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(~m[698]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[698]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[698]&m[1593]&~m[1595]&~m[1596]&m[1597])|(m[698]&~m[1593]&m[1595]&~m[1596]&m[1597])|(~m[698]&~m[1593]&~m[1595]&m[1596]&m[1597])|(m[698]&~m[1593]&~m[1595]&m[1596]&m[1597])|(~m[698]&m[1593]&~m[1595]&m[1596]&m[1597])|(m[698]&m[1593]&~m[1595]&m[1596]&m[1597])|(~m[698]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[698]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[698]&m[1593]&m[1595]&m[1596]&m[1597]))):InitCond[880];
    m[1599] = run?((((m[711]&~m[1598]&~m[1600]&~m[1601]&~m[1602])|(~m[711]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(m[711]&m[1598]&~m[1600]&m[1601]&~m[1602])|(m[711]&~m[1598]&m[1600]&m[1601]&~m[1602])|(~m[711]&m[1598]&~m[1600]&~m[1601]&m[1602])|(~m[711]&~m[1598]&m[1600]&~m[1601]&m[1602])|(m[711]&m[1598]&m[1600]&~m[1601]&m[1602])|(~m[711]&m[1598]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[378])|((m[711]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(~m[711]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[711]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[711]&m[1598]&~m[1600]&~m[1601]&m[1602])|(m[711]&~m[1598]&m[1600]&~m[1601]&m[1602])|(~m[711]&~m[1598]&~m[1600]&m[1601]&m[1602])|(m[711]&~m[1598]&~m[1600]&m[1601]&m[1602])|(~m[711]&m[1598]&~m[1600]&m[1601]&m[1602])|(m[711]&m[1598]&~m[1600]&m[1601]&m[1602])|(~m[711]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[711]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[711]&m[1598]&m[1600]&m[1601]&m[1602]))):InitCond[881];
    m[1604] = run?((((m[724]&~m[1603]&~m[1605]&~m[1606]&~m[1607])|(~m[724]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(m[724]&m[1603]&~m[1605]&m[1606]&~m[1607])|(m[724]&~m[1603]&m[1605]&m[1606]&~m[1607])|(~m[724]&m[1603]&~m[1605]&~m[1606]&m[1607])|(~m[724]&~m[1603]&m[1605]&~m[1606]&m[1607])|(m[724]&m[1603]&m[1605]&~m[1606]&m[1607])|(~m[724]&m[1603]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[379])|((m[724]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(~m[724]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[724]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[724]&m[1603]&~m[1605]&~m[1606]&m[1607])|(m[724]&~m[1603]&m[1605]&~m[1606]&m[1607])|(~m[724]&~m[1603]&~m[1605]&m[1606]&m[1607])|(m[724]&~m[1603]&~m[1605]&m[1606]&m[1607])|(~m[724]&m[1603]&~m[1605]&m[1606]&m[1607])|(m[724]&m[1603]&~m[1605]&m[1606]&m[1607])|(~m[724]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[724]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[724]&m[1603]&m[1605]&m[1606]&m[1607]))):InitCond[882];
    m[1609] = run?((((m[699]&~m[1608]&~m[1610]&~m[1611]&~m[1612])|(~m[699]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(m[699]&m[1608]&~m[1610]&m[1611]&~m[1612])|(m[699]&~m[1608]&m[1610]&m[1611]&~m[1612])|(~m[699]&m[1608]&~m[1610]&~m[1611]&m[1612])|(~m[699]&~m[1608]&m[1610]&~m[1611]&m[1612])|(m[699]&m[1608]&m[1610]&~m[1611]&m[1612])|(~m[699]&m[1608]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[380])|((m[699]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(~m[699]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[699]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[699]&m[1608]&~m[1610]&~m[1611]&m[1612])|(m[699]&~m[1608]&m[1610]&~m[1611]&m[1612])|(~m[699]&~m[1608]&~m[1610]&m[1611]&m[1612])|(m[699]&~m[1608]&~m[1610]&m[1611]&m[1612])|(~m[699]&m[1608]&~m[1610]&m[1611]&m[1612])|(m[699]&m[1608]&~m[1610]&m[1611]&m[1612])|(~m[699]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[699]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[699]&m[1608]&m[1610]&m[1611]&m[1612]))):InitCond[883];
    m[1614] = run?((((m[712]&~m[1613]&~m[1615]&~m[1616]&~m[1617])|(~m[712]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(m[712]&m[1613]&~m[1615]&m[1616]&~m[1617])|(m[712]&~m[1613]&m[1615]&m[1616]&~m[1617])|(~m[712]&m[1613]&~m[1615]&~m[1616]&m[1617])|(~m[712]&~m[1613]&m[1615]&~m[1616]&m[1617])|(m[712]&m[1613]&m[1615]&~m[1616]&m[1617])|(~m[712]&m[1613]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[381])|((m[712]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(~m[712]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[712]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[712]&m[1613]&~m[1615]&~m[1616]&m[1617])|(m[712]&~m[1613]&m[1615]&~m[1616]&m[1617])|(~m[712]&~m[1613]&~m[1615]&m[1616]&m[1617])|(m[712]&~m[1613]&~m[1615]&m[1616]&m[1617])|(~m[712]&m[1613]&~m[1615]&m[1616]&m[1617])|(m[712]&m[1613]&~m[1615]&m[1616]&m[1617])|(~m[712]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[712]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[712]&m[1613]&m[1615]&m[1616]&m[1617]))):InitCond[884];
    m[1619] = run?((((m[725]&~m[1618]&~m[1620]&~m[1621]&~m[1622])|(~m[725]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(m[725]&m[1618]&~m[1620]&m[1621]&~m[1622])|(m[725]&~m[1618]&m[1620]&m[1621]&~m[1622])|(~m[725]&m[1618]&~m[1620]&~m[1621]&m[1622])|(~m[725]&~m[1618]&m[1620]&~m[1621]&m[1622])|(m[725]&m[1618]&m[1620]&~m[1621]&m[1622])|(~m[725]&m[1618]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[382])|((m[725]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(~m[725]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[725]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[725]&m[1618]&~m[1620]&~m[1621]&m[1622])|(m[725]&~m[1618]&m[1620]&~m[1621]&m[1622])|(~m[725]&~m[1618]&~m[1620]&m[1621]&m[1622])|(m[725]&~m[1618]&~m[1620]&m[1621]&m[1622])|(~m[725]&m[1618]&~m[1620]&m[1621]&m[1622])|(m[725]&m[1618]&~m[1620]&m[1621]&m[1622])|(~m[725]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[725]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[725]&m[1618]&m[1620]&m[1621]&m[1622]))):InitCond[885];
    m[1624] = run?((((m[713]&~m[1623]&~m[1625]&~m[1626]&~m[1627])|(~m[713]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(m[713]&m[1623]&~m[1625]&m[1626]&~m[1627])|(m[713]&~m[1623]&m[1625]&m[1626]&~m[1627])|(~m[713]&m[1623]&~m[1625]&~m[1626]&m[1627])|(~m[713]&~m[1623]&m[1625]&~m[1626]&m[1627])|(m[713]&m[1623]&m[1625]&~m[1626]&m[1627])|(~m[713]&m[1623]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[383])|((m[713]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(~m[713]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[713]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[713]&m[1623]&~m[1625]&~m[1626]&m[1627])|(m[713]&~m[1623]&m[1625]&~m[1626]&m[1627])|(~m[713]&~m[1623]&~m[1625]&m[1626]&m[1627])|(m[713]&~m[1623]&~m[1625]&m[1626]&m[1627])|(~m[713]&m[1623]&~m[1625]&m[1626]&m[1627])|(m[713]&m[1623]&~m[1625]&m[1626]&m[1627])|(~m[713]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[713]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[713]&m[1623]&m[1625]&m[1626]&m[1627]))):InitCond[886];
    m[1629] = run?((((m[726]&~m[1628]&~m[1630]&~m[1631]&~m[1632])|(~m[726]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(m[726]&m[1628]&~m[1630]&m[1631]&~m[1632])|(m[726]&~m[1628]&m[1630]&m[1631]&~m[1632])|(~m[726]&m[1628]&~m[1630]&~m[1631]&m[1632])|(~m[726]&~m[1628]&m[1630]&~m[1631]&m[1632])|(m[726]&m[1628]&m[1630]&~m[1631]&m[1632])|(~m[726]&m[1628]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[384])|((m[726]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(~m[726]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[726]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[726]&m[1628]&~m[1630]&~m[1631]&m[1632])|(m[726]&~m[1628]&m[1630]&~m[1631]&m[1632])|(~m[726]&~m[1628]&~m[1630]&m[1631]&m[1632])|(m[726]&~m[1628]&~m[1630]&m[1631]&m[1632])|(~m[726]&m[1628]&~m[1630]&m[1631]&m[1632])|(m[726]&m[1628]&~m[1630]&m[1631]&m[1632])|(~m[726]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[726]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[726]&m[1628]&m[1630]&m[1631]&m[1632]))):InitCond[887];
    m[1634] = run?((((m[727]&~m[1633]&~m[1635]&~m[1636]&~m[1637])|(~m[727]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(m[727]&m[1633]&~m[1635]&m[1636]&~m[1637])|(m[727]&~m[1633]&m[1635]&m[1636]&~m[1637])|(~m[727]&m[1633]&~m[1635]&~m[1636]&m[1637])|(~m[727]&~m[1633]&m[1635]&~m[1636]&m[1637])|(m[727]&m[1633]&m[1635]&~m[1636]&m[1637])|(~m[727]&m[1633]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[385])|((m[727]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(~m[727]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[727]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[727]&m[1633]&~m[1635]&~m[1636]&m[1637])|(m[727]&~m[1633]&m[1635]&~m[1636]&m[1637])|(~m[727]&~m[1633]&~m[1635]&m[1636]&m[1637])|(m[727]&~m[1633]&~m[1635]&m[1636]&m[1637])|(~m[727]&m[1633]&~m[1635]&m[1636]&m[1637])|(m[727]&m[1633]&~m[1635]&m[1636]&m[1637])|(~m[727]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[727]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[727]&m[1633]&m[1635]&m[1636]&m[1637]))):InitCond[888];
end

always @(posedge color2_clk) begin
    m[336] = run?((((~m[42]&~m[140]&~m[532])|(m[42]&m[140]&~m[532]))&BiasedRNG[503])|(((m[42]&~m[140]&~m[532])|(~m[42]&m[140]&m[532]))&~BiasedRNG[503])|((~m[42]&~m[140]&m[532])|(m[42]&~m[140]&m[532])|(m[42]&m[140]&m[532]))):InitCond[889];
    m[337] = run?((((~m[42]&~m[154]&~m[533])|(m[42]&m[154]&~m[533]))&BiasedRNG[504])|(((m[42]&~m[154]&~m[533])|(~m[42]&m[154]&m[533]))&~BiasedRNG[504])|((~m[42]&~m[154]&m[533])|(m[42]&~m[154]&m[533])|(m[42]&m[154]&m[533]))):InitCond[890];
    m[338] = run?((((~m[98]&~m[168]&~m[534])|(m[98]&m[168]&~m[534]))&BiasedRNG[505])|(((m[98]&~m[168]&~m[534])|(~m[98]&m[168]&m[534]))&~BiasedRNG[505])|((~m[98]&~m[168]&m[534])|(m[98]&~m[168]&m[534])|(m[98]&m[168]&m[534]))):InitCond[891];
    m[339] = run?((((~m[98]&~m[182]&~m[535])|(m[98]&m[182]&~m[535]))&BiasedRNG[506])|(((m[98]&~m[182]&~m[535])|(~m[98]&m[182]&m[535]))&~BiasedRNG[506])|((~m[98]&~m[182]&m[535])|(m[98]&~m[182]&m[535])|(m[98]&m[182]&m[535]))):InitCond[892];
    m[340] = run?((((~m[98]&~m[196]&~m[536])|(m[98]&m[196]&~m[536]))&BiasedRNG[507])|(((m[98]&~m[196]&~m[536])|(~m[98]&m[196]&m[536]))&~BiasedRNG[507])|((~m[98]&~m[196]&m[536])|(m[98]&~m[196]&m[536])|(m[98]&m[196]&m[536]))):InitCond[893];
    m[341] = run?((((~m[98]&~m[210]&~m[537])|(m[98]&m[210]&~m[537]))&BiasedRNG[508])|(((m[98]&~m[210]&~m[537])|(~m[98]&m[210]&m[537]))&~BiasedRNG[508])|((~m[98]&~m[210]&m[537])|(m[98]&~m[210]&m[537])|(m[98]&m[210]&m[537]))):InitCond[894];
    m[350] = run?((((~m[43]&~m[141]&~m[546])|(m[43]&m[141]&~m[546]))&BiasedRNG[509])|(((m[43]&~m[141]&~m[546])|(~m[43]&m[141]&m[546]))&~BiasedRNG[509])|((~m[43]&~m[141]&m[546])|(m[43]&~m[141]&m[546])|(m[43]&m[141]&m[546]))):InitCond[895];
    m[351] = run?((((~m[43]&~m[155]&~m[547])|(m[43]&m[155]&~m[547]))&BiasedRNG[510])|(((m[43]&~m[155]&~m[547])|(~m[43]&m[155]&m[547]))&~BiasedRNG[510])|((~m[43]&~m[155]&m[547])|(m[43]&~m[155]&m[547])|(m[43]&m[155]&m[547]))):InitCond[896];
    m[352] = run?((((~m[101]&~m[169]&~m[548])|(m[101]&m[169]&~m[548]))&BiasedRNG[511])|(((m[101]&~m[169]&~m[548])|(~m[101]&m[169]&m[548]))&~BiasedRNG[511])|((~m[101]&~m[169]&m[548])|(m[101]&~m[169]&m[548])|(m[101]&m[169]&m[548]))):InitCond[897];
    m[353] = run?((((~m[101]&~m[183]&~m[549])|(m[101]&m[183]&~m[549]))&BiasedRNG[512])|(((m[101]&~m[183]&~m[549])|(~m[101]&m[183]&m[549]))&~BiasedRNG[512])|((~m[101]&~m[183]&m[549])|(m[101]&~m[183]&m[549])|(m[101]&m[183]&m[549]))):InitCond[898];
    m[354] = run?((((~m[101]&~m[197]&~m[550])|(m[101]&m[197]&~m[550]))&BiasedRNG[513])|(((m[101]&~m[197]&~m[550])|(~m[101]&m[197]&m[550]))&~BiasedRNG[513])|((~m[101]&~m[197]&m[550])|(m[101]&~m[197]&m[550])|(m[101]&m[197]&m[550]))):InitCond[899];
    m[355] = run?((((~m[101]&~m[211]&~m[551])|(m[101]&m[211]&~m[551]))&BiasedRNG[514])|(((m[101]&~m[211]&~m[551])|(~m[101]&m[211]&m[551]))&~BiasedRNG[514])|((~m[101]&~m[211]&m[551])|(m[101]&~m[211]&m[551])|(m[101]&m[211]&m[551]))):InitCond[900];
    m[364] = run?((((~m[44]&~m[142]&~m[560])|(m[44]&m[142]&~m[560]))&BiasedRNG[515])|(((m[44]&~m[142]&~m[560])|(~m[44]&m[142]&m[560]))&~BiasedRNG[515])|((~m[44]&~m[142]&m[560])|(m[44]&~m[142]&m[560])|(m[44]&m[142]&m[560]))):InitCond[901];
    m[365] = run?((((~m[44]&~m[156]&~m[561])|(m[44]&m[156]&~m[561]))&BiasedRNG[516])|(((m[44]&~m[156]&~m[561])|(~m[44]&m[156]&m[561]))&~BiasedRNG[516])|((~m[44]&~m[156]&m[561])|(m[44]&~m[156]&m[561])|(m[44]&m[156]&m[561]))):InitCond[902];
    m[366] = run?((((~m[104]&~m[170]&~m[562])|(m[104]&m[170]&~m[562]))&BiasedRNG[517])|(((m[104]&~m[170]&~m[562])|(~m[104]&m[170]&m[562]))&~BiasedRNG[517])|((~m[104]&~m[170]&m[562])|(m[104]&~m[170]&m[562])|(m[104]&m[170]&m[562]))):InitCond[903];
    m[367] = run?((((~m[104]&~m[184]&~m[563])|(m[104]&m[184]&~m[563]))&BiasedRNG[518])|(((m[104]&~m[184]&~m[563])|(~m[104]&m[184]&m[563]))&~BiasedRNG[518])|((~m[104]&~m[184]&m[563])|(m[104]&~m[184]&m[563])|(m[104]&m[184]&m[563]))):InitCond[904];
    m[368] = run?((((~m[104]&~m[198]&~m[564])|(m[104]&m[198]&~m[564]))&BiasedRNG[519])|(((m[104]&~m[198]&~m[564])|(~m[104]&m[198]&m[564]))&~BiasedRNG[519])|((~m[104]&~m[198]&m[564])|(m[104]&~m[198]&m[564])|(m[104]&m[198]&m[564]))):InitCond[905];
    m[369] = run?((((~m[104]&~m[212]&~m[565])|(m[104]&m[212]&~m[565]))&BiasedRNG[520])|(((m[104]&~m[212]&~m[565])|(~m[104]&m[212]&m[565]))&~BiasedRNG[520])|((~m[104]&~m[212]&m[565])|(m[104]&~m[212]&m[565])|(m[104]&m[212]&m[565]))):InitCond[906];
    m[378] = run?((((~m[45]&~m[143]&~m[574])|(m[45]&m[143]&~m[574]))&BiasedRNG[521])|(((m[45]&~m[143]&~m[574])|(~m[45]&m[143]&m[574]))&~BiasedRNG[521])|((~m[45]&~m[143]&m[574])|(m[45]&~m[143]&m[574])|(m[45]&m[143]&m[574]))):InitCond[907];
    m[379] = run?((((~m[45]&~m[157]&~m[575])|(m[45]&m[157]&~m[575]))&BiasedRNG[522])|(((m[45]&~m[157]&~m[575])|(~m[45]&m[157]&m[575]))&~BiasedRNG[522])|((~m[45]&~m[157]&m[575])|(m[45]&~m[157]&m[575])|(m[45]&m[157]&m[575]))):InitCond[908];
    m[380] = run?((((~m[107]&~m[171]&~m[576])|(m[107]&m[171]&~m[576]))&BiasedRNG[523])|(((m[107]&~m[171]&~m[576])|(~m[107]&m[171]&m[576]))&~BiasedRNG[523])|((~m[107]&~m[171]&m[576])|(m[107]&~m[171]&m[576])|(m[107]&m[171]&m[576]))):InitCond[909];
    m[381] = run?((((~m[107]&~m[185]&~m[577])|(m[107]&m[185]&~m[577]))&BiasedRNG[524])|(((m[107]&~m[185]&~m[577])|(~m[107]&m[185]&m[577]))&~BiasedRNG[524])|((~m[107]&~m[185]&m[577])|(m[107]&~m[185]&m[577])|(m[107]&m[185]&m[577]))):InitCond[910];
    m[382] = run?((((~m[107]&~m[199]&~m[578])|(m[107]&m[199]&~m[578]))&BiasedRNG[525])|(((m[107]&~m[199]&~m[578])|(~m[107]&m[199]&m[578]))&~BiasedRNG[525])|((~m[107]&~m[199]&m[578])|(m[107]&~m[199]&m[578])|(m[107]&m[199]&m[578]))):InitCond[911];
    m[383] = run?((((~m[107]&~m[213]&~m[579])|(m[107]&m[213]&~m[579]))&BiasedRNG[526])|(((m[107]&~m[213]&~m[579])|(~m[107]&m[213]&m[579]))&~BiasedRNG[526])|((~m[107]&~m[213]&m[579])|(m[107]&~m[213]&m[579])|(m[107]&m[213]&m[579]))):InitCond[912];
    m[392] = run?((((~m[46]&~m[144]&~m[588])|(m[46]&m[144]&~m[588]))&BiasedRNG[527])|(((m[46]&~m[144]&~m[588])|(~m[46]&m[144]&m[588]))&~BiasedRNG[527])|((~m[46]&~m[144]&m[588])|(m[46]&~m[144]&m[588])|(m[46]&m[144]&m[588]))):InitCond[913];
    m[393] = run?((((~m[46]&~m[158]&~m[589])|(m[46]&m[158]&~m[589]))&BiasedRNG[528])|(((m[46]&~m[158]&~m[589])|(~m[46]&m[158]&m[589]))&~BiasedRNG[528])|((~m[46]&~m[158]&m[589])|(m[46]&~m[158]&m[589])|(m[46]&m[158]&m[589]))):InitCond[914];
    m[394] = run?((((~m[110]&~m[172]&~m[590])|(m[110]&m[172]&~m[590]))&BiasedRNG[529])|(((m[110]&~m[172]&~m[590])|(~m[110]&m[172]&m[590]))&~BiasedRNG[529])|((~m[110]&~m[172]&m[590])|(m[110]&~m[172]&m[590])|(m[110]&m[172]&m[590]))):InitCond[915];
    m[395] = run?((((~m[110]&~m[186]&~m[591])|(m[110]&m[186]&~m[591]))&BiasedRNG[530])|(((m[110]&~m[186]&~m[591])|(~m[110]&m[186]&m[591]))&~BiasedRNG[530])|((~m[110]&~m[186]&m[591])|(m[110]&~m[186]&m[591])|(m[110]&m[186]&m[591]))):InitCond[916];
    m[396] = run?((((~m[110]&~m[200]&~m[592])|(m[110]&m[200]&~m[592]))&BiasedRNG[531])|(((m[110]&~m[200]&~m[592])|(~m[110]&m[200]&m[592]))&~BiasedRNG[531])|((~m[110]&~m[200]&m[592])|(m[110]&~m[200]&m[592])|(m[110]&m[200]&m[592]))):InitCond[917];
    m[397] = run?((((~m[110]&~m[214]&~m[593])|(m[110]&m[214]&~m[593]))&BiasedRNG[532])|(((m[110]&~m[214]&~m[593])|(~m[110]&m[214]&m[593]))&~BiasedRNG[532])|((~m[110]&~m[214]&m[593])|(m[110]&~m[214]&m[593])|(m[110]&m[214]&m[593]))):InitCond[918];
    m[406] = run?((((~m[47]&~m[145]&~m[602])|(m[47]&m[145]&~m[602]))&BiasedRNG[533])|(((m[47]&~m[145]&~m[602])|(~m[47]&m[145]&m[602]))&~BiasedRNG[533])|((~m[47]&~m[145]&m[602])|(m[47]&~m[145]&m[602])|(m[47]&m[145]&m[602]))):InitCond[919];
    m[407] = run?((((~m[47]&~m[159]&~m[603])|(m[47]&m[159]&~m[603]))&BiasedRNG[534])|(((m[47]&~m[159]&~m[603])|(~m[47]&m[159]&m[603]))&~BiasedRNG[534])|((~m[47]&~m[159]&m[603])|(m[47]&~m[159]&m[603])|(m[47]&m[159]&m[603]))):InitCond[920];
    m[408] = run?((((~m[113]&~m[173]&~m[604])|(m[113]&m[173]&~m[604]))&BiasedRNG[535])|(((m[113]&~m[173]&~m[604])|(~m[113]&m[173]&m[604]))&~BiasedRNG[535])|((~m[113]&~m[173]&m[604])|(m[113]&~m[173]&m[604])|(m[113]&m[173]&m[604]))):InitCond[921];
    m[409] = run?((((~m[113]&~m[187]&~m[605])|(m[113]&m[187]&~m[605]))&BiasedRNG[536])|(((m[113]&~m[187]&~m[605])|(~m[113]&m[187]&m[605]))&~BiasedRNG[536])|((~m[113]&~m[187]&m[605])|(m[113]&~m[187]&m[605])|(m[113]&m[187]&m[605]))):InitCond[922];
    m[410] = run?((((~m[113]&~m[201]&~m[606])|(m[113]&m[201]&~m[606]))&BiasedRNG[537])|(((m[113]&~m[201]&~m[606])|(~m[113]&m[201]&m[606]))&~BiasedRNG[537])|((~m[113]&~m[201]&m[606])|(m[113]&~m[201]&m[606])|(m[113]&m[201]&m[606]))):InitCond[923];
    m[411] = run?((((~m[113]&~m[215]&~m[607])|(m[113]&m[215]&~m[607]))&BiasedRNG[538])|(((m[113]&~m[215]&~m[607])|(~m[113]&m[215]&m[607]))&~BiasedRNG[538])|((~m[113]&~m[215]&m[607])|(m[113]&~m[215]&m[607])|(m[113]&m[215]&m[607]))):InitCond[924];
    m[426] = run?((((~m[117]&~m[230]&~m[622])|(m[117]&m[230]&~m[622]))&BiasedRNG[539])|(((m[117]&~m[230]&~m[622])|(~m[117]&m[230]&m[622]))&~BiasedRNG[539])|((~m[117]&~m[230]&m[622])|(m[117]&~m[230]&m[622])|(m[117]&m[230]&m[622]))):InitCond[925];
    m[427] = run?((((~m[117]&~m[244]&~m[623])|(m[117]&m[244]&~m[623]))&BiasedRNG[540])|(((m[117]&~m[244]&~m[623])|(~m[117]&m[244]&m[623]))&~BiasedRNG[540])|((~m[117]&~m[244]&m[623])|(m[117]&~m[244]&m[623])|(m[117]&m[244]&m[623]))):InitCond[926];
    m[428] = run?((((~m[117]&~m[258]&~m[624])|(m[117]&m[258]&~m[624]))&BiasedRNG[541])|(((m[117]&~m[258]&~m[624])|(~m[117]&m[258]&m[624]))&~BiasedRNG[541])|((~m[117]&~m[258]&m[624])|(m[117]&~m[258]&m[624])|(m[117]&m[258]&m[624]))):InitCond[927];
    m[429] = run?((((~m[117]&~m[272]&~m[625])|(m[117]&m[272]&~m[625]))&BiasedRNG[542])|(((m[117]&~m[272]&~m[625])|(~m[117]&m[272]&m[625]))&~BiasedRNG[542])|((~m[117]&~m[272]&m[625])|(m[117]&~m[272]&m[625])|(m[117]&m[272]&m[625]))):InitCond[928];
    m[430] = run?((((~m[118]&~m[286]&~m[626])|(m[118]&m[286]&~m[626]))&BiasedRNG[543])|(((m[118]&~m[286]&~m[626])|(~m[118]&m[286]&m[626]))&~BiasedRNG[543])|((~m[118]&~m[286]&m[626])|(m[118]&~m[286]&m[626])|(m[118]&m[286]&m[626]))):InitCond[929];
    m[431] = run?((((~m[118]&~m[300]&~m[627])|(m[118]&m[300]&~m[627]))&BiasedRNG[544])|(((m[118]&~m[300]&~m[627])|(~m[118]&m[300]&m[627]))&~BiasedRNG[544])|((~m[118]&~m[300]&m[627])|(m[118]&~m[300]&m[627])|(m[118]&m[300]&m[627]))):InitCond[930];
    m[432] = run?((((~m[118]&~m[314]&~m[628])|(m[118]&m[314]&~m[628]))&BiasedRNG[545])|(((m[118]&~m[314]&~m[628])|(~m[118]&m[314]&m[628]))&~BiasedRNG[545])|((~m[118]&~m[314]&m[628])|(m[118]&~m[314]&m[628])|(m[118]&m[314]&m[628]))):InitCond[931];
    m[433] = run?((((~m[118]&~m[328]&~m[629])|(m[118]&m[328]&~m[629]))&BiasedRNG[546])|(((m[118]&~m[328]&~m[629])|(~m[118]&m[328]&m[629]))&~BiasedRNG[546])|((~m[118]&~m[328]&m[629])|(m[118]&~m[328]&m[629])|(m[118]&m[328]&m[629]))):InitCond[932];
    m[440] = run?((((~m[120]&~m[231]&~m[636])|(m[120]&m[231]&~m[636]))&BiasedRNG[547])|(((m[120]&~m[231]&~m[636])|(~m[120]&m[231]&m[636]))&~BiasedRNG[547])|((~m[120]&~m[231]&m[636])|(m[120]&~m[231]&m[636])|(m[120]&m[231]&m[636]))):InitCond[933];
    m[441] = run?((((~m[120]&~m[245]&~m[637])|(m[120]&m[245]&~m[637]))&BiasedRNG[548])|(((m[120]&~m[245]&~m[637])|(~m[120]&m[245]&m[637]))&~BiasedRNG[548])|((~m[120]&~m[245]&m[637])|(m[120]&~m[245]&m[637])|(m[120]&m[245]&m[637]))):InitCond[934];
    m[442] = run?((((~m[120]&~m[259]&~m[638])|(m[120]&m[259]&~m[638]))&BiasedRNG[549])|(((m[120]&~m[259]&~m[638])|(~m[120]&m[259]&m[638]))&~BiasedRNG[549])|((~m[120]&~m[259]&m[638])|(m[120]&~m[259]&m[638])|(m[120]&m[259]&m[638]))):InitCond[935];
    m[443] = run?((((~m[120]&~m[273]&~m[639])|(m[120]&m[273]&~m[639]))&BiasedRNG[550])|(((m[120]&~m[273]&~m[639])|(~m[120]&m[273]&m[639]))&~BiasedRNG[550])|((~m[120]&~m[273]&m[639])|(m[120]&~m[273]&m[639])|(m[120]&m[273]&m[639]))):InitCond[936];
    m[444] = run?((((~m[121]&~m[287]&~m[640])|(m[121]&m[287]&~m[640]))&BiasedRNG[551])|(((m[121]&~m[287]&~m[640])|(~m[121]&m[287]&m[640]))&~BiasedRNG[551])|((~m[121]&~m[287]&m[640])|(m[121]&~m[287]&m[640])|(m[121]&m[287]&m[640]))):InitCond[937];
    m[445] = run?((((~m[121]&~m[301]&~m[641])|(m[121]&m[301]&~m[641]))&BiasedRNG[552])|(((m[121]&~m[301]&~m[641])|(~m[121]&m[301]&m[641]))&~BiasedRNG[552])|((~m[121]&~m[301]&m[641])|(m[121]&~m[301]&m[641])|(m[121]&m[301]&m[641]))):InitCond[938];
    m[446] = run?((((~m[121]&~m[315]&~m[642])|(m[121]&m[315]&~m[642]))&BiasedRNG[553])|(((m[121]&~m[315]&~m[642])|(~m[121]&m[315]&m[642]))&~BiasedRNG[553])|((~m[121]&~m[315]&m[642])|(m[121]&~m[315]&m[642])|(m[121]&m[315]&m[642]))):InitCond[939];
    m[447] = run?((((~m[121]&~m[329]&~m[643])|(m[121]&m[329]&~m[643]))&BiasedRNG[554])|(((m[121]&~m[329]&~m[643])|(~m[121]&m[329]&m[643]))&~BiasedRNG[554])|((~m[121]&~m[329]&m[643])|(m[121]&~m[329]&m[643])|(m[121]&m[329]&m[643]))):InitCond[940];
    m[454] = run?((((~m[123]&~m[232]&~m[650])|(m[123]&m[232]&~m[650]))&BiasedRNG[555])|(((m[123]&~m[232]&~m[650])|(~m[123]&m[232]&m[650]))&~BiasedRNG[555])|((~m[123]&~m[232]&m[650])|(m[123]&~m[232]&m[650])|(m[123]&m[232]&m[650]))):InitCond[941];
    m[455] = run?((((~m[123]&~m[246]&~m[651])|(m[123]&m[246]&~m[651]))&BiasedRNG[556])|(((m[123]&~m[246]&~m[651])|(~m[123]&m[246]&m[651]))&~BiasedRNG[556])|((~m[123]&~m[246]&m[651])|(m[123]&~m[246]&m[651])|(m[123]&m[246]&m[651]))):InitCond[942];
    m[456] = run?((((~m[123]&~m[260]&~m[652])|(m[123]&m[260]&~m[652]))&BiasedRNG[557])|(((m[123]&~m[260]&~m[652])|(~m[123]&m[260]&m[652]))&~BiasedRNG[557])|((~m[123]&~m[260]&m[652])|(m[123]&~m[260]&m[652])|(m[123]&m[260]&m[652]))):InitCond[943];
    m[457] = run?((((~m[123]&~m[274]&~m[653])|(m[123]&m[274]&~m[653]))&BiasedRNG[558])|(((m[123]&~m[274]&~m[653])|(~m[123]&m[274]&m[653]))&~BiasedRNG[558])|((~m[123]&~m[274]&m[653])|(m[123]&~m[274]&m[653])|(m[123]&m[274]&m[653]))):InitCond[944];
    m[458] = run?((((~m[124]&~m[288]&~m[654])|(m[124]&m[288]&~m[654]))&BiasedRNG[559])|(((m[124]&~m[288]&~m[654])|(~m[124]&m[288]&m[654]))&~BiasedRNG[559])|((~m[124]&~m[288]&m[654])|(m[124]&~m[288]&m[654])|(m[124]&m[288]&m[654]))):InitCond[945];
    m[459] = run?((((~m[124]&~m[302]&~m[655])|(m[124]&m[302]&~m[655]))&BiasedRNG[560])|(((m[124]&~m[302]&~m[655])|(~m[124]&m[302]&m[655]))&~BiasedRNG[560])|((~m[124]&~m[302]&m[655])|(m[124]&~m[302]&m[655])|(m[124]&m[302]&m[655]))):InitCond[946];
    m[460] = run?((((~m[124]&~m[316]&~m[656])|(m[124]&m[316]&~m[656]))&BiasedRNG[561])|(((m[124]&~m[316]&~m[656])|(~m[124]&m[316]&m[656]))&~BiasedRNG[561])|((~m[124]&~m[316]&m[656])|(m[124]&~m[316]&m[656])|(m[124]&m[316]&m[656]))):InitCond[947];
    m[461] = run?((((~m[124]&~m[330]&~m[657])|(m[124]&m[330]&~m[657]))&BiasedRNG[562])|(((m[124]&~m[330]&~m[657])|(~m[124]&m[330]&m[657]))&~BiasedRNG[562])|((~m[124]&~m[330]&m[657])|(m[124]&~m[330]&m[657])|(m[124]&m[330]&m[657]))):InitCond[948];
    m[468] = run?((((~m[126]&~m[233]&~m[664])|(m[126]&m[233]&~m[664]))&BiasedRNG[563])|(((m[126]&~m[233]&~m[664])|(~m[126]&m[233]&m[664]))&~BiasedRNG[563])|((~m[126]&~m[233]&m[664])|(m[126]&~m[233]&m[664])|(m[126]&m[233]&m[664]))):InitCond[949];
    m[469] = run?((((~m[126]&~m[247]&~m[665])|(m[126]&m[247]&~m[665]))&BiasedRNG[564])|(((m[126]&~m[247]&~m[665])|(~m[126]&m[247]&m[665]))&~BiasedRNG[564])|((~m[126]&~m[247]&m[665])|(m[126]&~m[247]&m[665])|(m[126]&m[247]&m[665]))):InitCond[950];
    m[470] = run?((((~m[126]&~m[261]&~m[666])|(m[126]&m[261]&~m[666]))&BiasedRNG[565])|(((m[126]&~m[261]&~m[666])|(~m[126]&m[261]&m[666]))&~BiasedRNG[565])|((~m[126]&~m[261]&m[666])|(m[126]&~m[261]&m[666])|(m[126]&m[261]&m[666]))):InitCond[951];
    m[471] = run?((((~m[126]&~m[275]&~m[667])|(m[126]&m[275]&~m[667]))&BiasedRNG[566])|(((m[126]&~m[275]&~m[667])|(~m[126]&m[275]&m[667]))&~BiasedRNG[566])|((~m[126]&~m[275]&m[667])|(m[126]&~m[275]&m[667])|(m[126]&m[275]&m[667]))):InitCond[952];
    m[472] = run?((((~m[127]&~m[289]&~m[668])|(m[127]&m[289]&~m[668]))&BiasedRNG[567])|(((m[127]&~m[289]&~m[668])|(~m[127]&m[289]&m[668]))&~BiasedRNG[567])|((~m[127]&~m[289]&m[668])|(m[127]&~m[289]&m[668])|(m[127]&m[289]&m[668]))):InitCond[953];
    m[473] = run?((((~m[127]&~m[303]&~m[669])|(m[127]&m[303]&~m[669]))&BiasedRNG[568])|(((m[127]&~m[303]&~m[669])|(~m[127]&m[303]&m[669]))&~BiasedRNG[568])|((~m[127]&~m[303]&m[669])|(m[127]&~m[303]&m[669])|(m[127]&m[303]&m[669]))):InitCond[954];
    m[474] = run?((((~m[127]&~m[317]&~m[670])|(m[127]&m[317]&~m[670]))&BiasedRNG[569])|(((m[127]&~m[317]&~m[670])|(~m[127]&m[317]&m[670]))&~BiasedRNG[569])|((~m[127]&~m[317]&m[670])|(m[127]&~m[317]&m[670])|(m[127]&m[317]&m[670]))):InitCond[955];
    m[475] = run?((((~m[127]&~m[331]&~m[671])|(m[127]&m[331]&~m[671]))&BiasedRNG[570])|(((m[127]&~m[331]&~m[671])|(~m[127]&m[331]&m[671]))&~BiasedRNG[570])|((~m[127]&~m[331]&m[671])|(m[127]&~m[331]&m[671])|(m[127]&m[331]&m[671]))):InitCond[956];
    m[482] = run?((((~m[129]&~m[234]&~m[678])|(m[129]&m[234]&~m[678]))&BiasedRNG[571])|(((m[129]&~m[234]&~m[678])|(~m[129]&m[234]&m[678]))&~BiasedRNG[571])|((~m[129]&~m[234]&m[678])|(m[129]&~m[234]&m[678])|(m[129]&m[234]&m[678]))):InitCond[957];
    m[483] = run?((((~m[129]&~m[248]&~m[679])|(m[129]&m[248]&~m[679]))&BiasedRNG[572])|(((m[129]&~m[248]&~m[679])|(~m[129]&m[248]&m[679]))&~BiasedRNG[572])|((~m[129]&~m[248]&m[679])|(m[129]&~m[248]&m[679])|(m[129]&m[248]&m[679]))):InitCond[958];
    m[484] = run?((((~m[129]&~m[262]&~m[680])|(m[129]&m[262]&~m[680]))&BiasedRNG[573])|(((m[129]&~m[262]&~m[680])|(~m[129]&m[262]&m[680]))&~BiasedRNG[573])|((~m[129]&~m[262]&m[680])|(m[129]&~m[262]&m[680])|(m[129]&m[262]&m[680]))):InitCond[959];
    m[485] = run?((((~m[129]&~m[276]&~m[681])|(m[129]&m[276]&~m[681]))&BiasedRNG[574])|(((m[129]&~m[276]&~m[681])|(~m[129]&m[276]&m[681]))&~BiasedRNG[574])|((~m[129]&~m[276]&m[681])|(m[129]&~m[276]&m[681])|(m[129]&m[276]&m[681]))):InitCond[960];
    m[486] = run?((((~m[130]&~m[290]&~m[682])|(m[130]&m[290]&~m[682]))&BiasedRNG[575])|(((m[130]&~m[290]&~m[682])|(~m[130]&m[290]&m[682]))&~BiasedRNG[575])|((~m[130]&~m[290]&m[682])|(m[130]&~m[290]&m[682])|(m[130]&m[290]&m[682]))):InitCond[961];
    m[487] = run?((((~m[130]&~m[304]&~m[683])|(m[130]&m[304]&~m[683]))&BiasedRNG[576])|(((m[130]&~m[304]&~m[683])|(~m[130]&m[304]&m[683]))&~BiasedRNG[576])|((~m[130]&~m[304]&m[683])|(m[130]&~m[304]&m[683])|(m[130]&m[304]&m[683]))):InitCond[962];
    m[488] = run?((((~m[130]&~m[318]&~m[684])|(m[130]&m[318]&~m[684]))&BiasedRNG[577])|(((m[130]&~m[318]&~m[684])|(~m[130]&m[318]&m[684]))&~BiasedRNG[577])|((~m[130]&~m[318]&m[684])|(m[130]&~m[318]&m[684])|(m[130]&m[318]&m[684]))):InitCond[963];
    m[489] = run?((((~m[130]&~m[332]&~m[685])|(m[130]&m[332]&~m[685]))&BiasedRNG[578])|(((m[130]&~m[332]&~m[685])|(~m[130]&m[332]&m[685]))&~BiasedRNG[578])|((~m[130]&~m[332]&m[685])|(m[130]&~m[332]&m[685])|(m[130]&m[332]&m[685]))):InitCond[964];
    m[496] = run?((((~m[132]&~m[235]&~m[692])|(m[132]&m[235]&~m[692]))&BiasedRNG[579])|(((m[132]&~m[235]&~m[692])|(~m[132]&m[235]&m[692]))&~BiasedRNG[579])|((~m[132]&~m[235]&m[692])|(m[132]&~m[235]&m[692])|(m[132]&m[235]&m[692]))):InitCond[965];
    m[497] = run?((((~m[132]&~m[249]&~m[693])|(m[132]&m[249]&~m[693]))&BiasedRNG[580])|(((m[132]&~m[249]&~m[693])|(~m[132]&m[249]&m[693]))&~BiasedRNG[580])|((~m[132]&~m[249]&m[693])|(m[132]&~m[249]&m[693])|(m[132]&m[249]&m[693]))):InitCond[966];
    m[498] = run?((((~m[132]&~m[263]&~m[694])|(m[132]&m[263]&~m[694]))&BiasedRNG[581])|(((m[132]&~m[263]&~m[694])|(~m[132]&m[263]&m[694]))&~BiasedRNG[581])|((~m[132]&~m[263]&m[694])|(m[132]&~m[263]&m[694])|(m[132]&m[263]&m[694]))):InitCond[967];
    m[499] = run?((((~m[132]&~m[277]&~m[695])|(m[132]&m[277]&~m[695]))&BiasedRNG[582])|(((m[132]&~m[277]&~m[695])|(~m[132]&m[277]&m[695]))&~BiasedRNG[582])|((~m[132]&~m[277]&m[695])|(m[132]&~m[277]&m[695])|(m[132]&m[277]&m[695]))):InitCond[968];
    m[500] = run?((((~m[133]&~m[291]&~m[696])|(m[133]&m[291]&~m[696]))&BiasedRNG[583])|(((m[133]&~m[291]&~m[696])|(~m[133]&m[291]&m[696]))&~BiasedRNG[583])|((~m[133]&~m[291]&m[696])|(m[133]&~m[291]&m[696])|(m[133]&m[291]&m[696]))):InitCond[969];
    m[501] = run?((((~m[133]&~m[305]&~m[697])|(m[133]&m[305]&~m[697]))&BiasedRNG[584])|(((m[133]&~m[305]&~m[697])|(~m[133]&m[305]&m[697]))&~BiasedRNG[584])|((~m[133]&~m[305]&m[697])|(m[133]&~m[305]&m[697])|(m[133]&m[305]&m[697]))):InitCond[970];
    m[502] = run?((((~m[133]&~m[319]&~m[698])|(m[133]&m[319]&~m[698]))&BiasedRNG[585])|(((m[133]&~m[319]&~m[698])|(~m[133]&m[319]&m[698]))&~BiasedRNG[585])|((~m[133]&~m[319]&m[698])|(m[133]&~m[319]&m[698])|(m[133]&m[319]&m[698]))):InitCond[971];
    m[503] = run?((((~m[133]&~m[333]&~m[699])|(m[133]&m[333]&~m[699]))&BiasedRNG[586])|(((m[133]&~m[333]&~m[699])|(~m[133]&m[333]&m[699]))&~BiasedRNG[586])|((~m[133]&~m[333]&m[699])|(m[133]&~m[333]&m[699])|(m[133]&m[333]&m[699]))):InitCond[972];
    m[510] = run?((((~m[135]&~m[236]&~m[706])|(m[135]&m[236]&~m[706]))&BiasedRNG[587])|(((m[135]&~m[236]&~m[706])|(~m[135]&m[236]&m[706]))&~BiasedRNG[587])|((~m[135]&~m[236]&m[706])|(m[135]&~m[236]&m[706])|(m[135]&m[236]&m[706]))):InitCond[973];
    m[511] = run?((((~m[135]&~m[250]&~m[707])|(m[135]&m[250]&~m[707]))&BiasedRNG[588])|(((m[135]&~m[250]&~m[707])|(~m[135]&m[250]&m[707]))&~BiasedRNG[588])|((~m[135]&~m[250]&m[707])|(m[135]&~m[250]&m[707])|(m[135]&m[250]&m[707]))):InitCond[974];
    m[512] = run?((((~m[135]&~m[264]&~m[708])|(m[135]&m[264]&~m[708]))&BiasedRNG[589])|(((m[135]&~m[264]&~m[708])|(~m[135]&m[264]&m[708]))&~BiasedRNG[589])|((~m[135]&~m[264]&m[708])|(m[135]&~m[264]&m[708])|(m[135]&m[264]&m[708]))):InitCond[975];
    m[513] = run?((((~m[135]&~m[278]&~m[709])|(m[135]&m[278]&~m[709]))&BiasedRNG[590])|(((m[135]&~m[278]&~m[709])|(~m[135]&m[278]&m[709]))&~BiasedRNG[590])|((~m[135]&~m[278]&m[709])|(m[135]&~m[278]&m[709])|(m[135]&m[278]&m[709]))):InitCond[976];
    m[514] = run?((((~m[136]&~m[292]&~m[710])|(m[136]&m[292]&~m[710]))&BiasedRNG[591])|(((m[136]&~m[292]&~m[710])|(~m[136]&m[292]&m[710]))&~BiasedRNG[591])|((~m[136]&~m[292]&m[710])|(m[136]&~m[292]&m[710])|(m[136]&m[292]&m[710]))):InitCond[977];
    m[515] = run?((((~m[136]&~m[306]&~m[711])|(m[136]&m[306]&~m[711]))&BiasedRNG[592])|(((m[136]&~m[306]&~m[711])|(~m[136]&m[306]&m[711]))&~BiasedRNG[592])|((~m[136]&~m[306]&m[711])|(m[136]&~m[306]&m[711])|(m[136]&m[306]&m[711]))):InitCond[978];
    m[516] = run?((((~m[136]&~m[320]&~m[712])|(m[136]&m[320]&~m[712]))&BiasedRNG[593])|(((m[136]&~m[320]&~m[712])|(~m[136]&m[320]&m[712]))&~BiasedRNG[593])|((~m[136]&~m[320]&m[712])|(m[136]&~m[320]&m[712])|(m[136]&m[320]&m[712]))):InitCond[979];
    m[517] = run?((((~m[136]&~m[334]&~m[713])|(m[136]&m[334]&~m[713]))&BiasedRNG[594])|(((m[136]&~m[334]&~m[713])|(~m[136]&m[334]&m[713]))&~BiasedRNG[594])|((~m[136]&~m[334]&m[713])|(m[136]&~m[334]&m[713])|(m[136]&m[334]&m[713]))):InitCond[980];
    m[524] = run?((((~m[138]&~m[237]&~m[720])|(m[138]&m[237]&~m[720]))&BiasedRNG[595])|(((m[138]&~m[237]&~m[720])|(~m[138]&m[237]&m[720]))&~BiasedRNG[595])|((~m[138]&~m[237]&m[720])|(m[138]&~m[237]&m[720])|(m[138]&m[237]&m[720]))):InitCond[981];
    m[525] = run?((((~m[138]&~m[251]&~m[721])|(m[138]&m[251]&~m[721]))&BiasedRNG[596])|(((m[138]&~m[251]&~m[721])|(~m[138]&m[251]&m[721]))&~BiasedRNG[596])|((~m[138]&~m[251]&m[721])|(m[138]&~m[251]&m[721])|(m[138]&m[251]&m[721]))):InitCond[982];
    m[526] = run?((((~m[138]&~m[265]&~m[722])|(m[138]&m[265]&~m[722]))&BiasedRNG[597])|(((m[138]&~m[265]&~m[722])|(~m[138]&m[265]&m[722]))&~BiasedRNG[597])|((~m[138]&~m[265]&m[722])|(m[138]&~m[265]&m[722])|(m[138]&m[265]&m[722]))):InitCond[983];
    m[527] = run?((((~m[138]&~m[279]&~m[723])|(m[138]&m[279]&~m[723]))&BiasedRNG[598])|(((m[138]&~m[279]&~m[723])|(~m[138]&m[279]&m[723]))&~BiasedRNG[598])|((~m[138]&~m[279]&m[723])|(m[138]&~m[279]&m[723])|(m[138]&m[279]&m[723]))):InitCond[984];
    m[528] = run?((((~m[139]&~m[293]&~m[724])|(m[139]&m[293]&~m[724]))&BiasedRNG[599])|(((m[139]&~m[293]&~m[724])|(~m[139]&m[293]&m[724]))&~BiasedRNG[599])|((~m[139]&~m[293]&m[724])|(m[139]&~m[293]&m[724])|(m[139]&m[293]&m[724]))):InitCond[985];
    m[529] = run?((((~m[139]&~m[307]&~m[725])|(m[139]&m[307]&~m[725]))&BiasedRNG[600])|(((m[139]&~m[307]&~m[725])|(~m[139]&m[307]&m[725]))&~BiasedRNG[600])|((~m[139]&~m[307]&m[725])|(m[139]&~m[307]&m[725])|(m[139]&m[307]&m[725]))):InitCond[986];
    m[530] = run?((((~m[139]&~m[321]&~m[726])|(m[139]&m[321]&~m[726]))&BiasedRNG[601])|(((m[139]&~m[321]&~m[726])|(~m[139]&m[321]&m[726]))&~BiasedRNG[601])|((~m[139]&~m[321]&m[726])|(m[139]&~m[321]&m[726])|(m[139]&m[321]&m[726]))):InitCond[987];
    m[531] = run?((((~m[139]&~m[335]&~m[727])|(m[139]&m[335]&~m[727]))&BiasedRNG[602])|(((m[139]&~m[335]&~m[727])|(~m[139]&m[335]&m[727]))&~BiasedRNG[602])|((~m[139]&~m[335]&m[727])|(m[139]&~m[335]&m[727])|(m[139]&m[335]&m[727]))):InitCond[988];
    m[538] = run?((((m[224]&~m[342]&m[803])|(~m[224]&m[342]&m[803]))&BiasedRNG[603])|(((m[224]&m[342]&~m[803]))&~BiasedRNG[603])|((m[224]&m[342]&m[803]))):InitCond[989];
    m[539] = run?((((m[238]&~m[343]&m[833])|(~m[238]&m[343]&m[833]))&BiasedRNG[604])|(((m[238]&m[343]&~m[833]))&~BiasedRNG[604])|((m[238]&m[343]&m[833]))):InitCond[990];
    m[540] = run?((((m[252]&~m[344]&m[868])|(~m[252]&m[344]&m[868]))&BiasedRNG[605])|(((m[252]&m[344]&~m[868]))&~BiasedRNG[605])|((m[252]&m[344]&m[868]))):InitCond[991];
    m[541] = run?((((m[266]&~m[345]&m[908])|(~m[266]&m[345]&m[908]))&BiasedRNG[606])|(((m[266]&m[345]&~m[908]))&~BiasedRNG[606])|((m[266]&m[345]&m[908]))):InitCond[992];
    m[542] = run?((((m[280]&~m[346]&m[953])|(~m[280]&m[346]&m[953]))&BiasedRNG[607])|(((m[280]&m[346]&~m[953]))&~BiasedRNG[607])|((m[280]&m[346]&m[953]))):InitCond[993];
    m[543] = run?((((m[294]&~m[347]&m[1003])|(~m[294]&m[347]&m[1003]))&BiasedRNG[608])|(((m[294]&m[347]&~m[1003]))&~BiasedRNG[608])|((m[294]&m[347]&m[1003]))):InitCond[994];
    m[544] = run?((((m[308]&~m[348]&m[1058])|(~m[308]&m[348]&m[1058]))&BiasedRNG[609])|(((m[308]&m[348]&~m[1058]))&~BiasedRNG[609])|((m[308]&m[348]&m[1058]))):InitCond[995];
    m[545] = run?((((m[322]&~m[349]&m[1118])|(~m[322]&m[349]&m[1118]))&BiasedRNG[610])|(((m[322]&m[349]&~m[1118]))&~BiasedRNG[610])|((m[322]&m[349]&m[1118]))):InitCond[996];
    m[552] = run?((((m[225]&~m[356]&m[834])|(~m[225]&m[356]&m[834]))&BiasedRNG[611])|(((m[225]&m[356]&~m[834]))&~BiasedRNG[611])|((m[225]&m[356]&m[834]))):InitCond[997];
    m[553] = run?((((m[239]&~m[357]&m[869])|(~m[239]&m[357]&m[869]))&BiasedRNG[612])|(((m[239]&m[357]&~m[869]))&~BiasedRNG[612])|((m[239]&m[357]&m[869]))):InitCond[998];
    m[554] = run?((((m[253]&~m[358]&m[909])|(~m[253]&m[358]&m[909]))&BiasedRNG[613])|(((m[253]&m[358]&~m[909]))&~BiasedRNG[613])|((m[253]&m[358]&m[909]))):InitCond[999];
    m[555] = run?((((m[267]&~m[359]&m[954])|(~m[267]&m[359]&m[954]))&BiasedRNG[614])|(((m[267]&m[359]&~m[954]))&~BiasedRNG[614])|((m[267]&m[359]&m[954]))):InitCond[1000];
    m[556] = run?((((m[281]&~m[360]&m[1004])|(~m[281]&m[360]&m[1004]))&BiasedRNG[615])|(((m[281]&m[360]&~m[1004]))&~BiasedRNG[615])|((m[281]&m[360]&m[1004]))):InitCond[1001];
    m[557] = run?((((m[295]&~m[361]&m[1059])|(~m[295]&m[361]&m[1059]))&BiasedRNG[616])|(((m[295]&m[361]&~m[1059]))&~BiasedRNG[616])|((m[295]&m[361]&m[1059]))):InitCond[1002];
    m[558] = run?((((m[309]&~m[362]&m[1119])|(~m[309]&m[362]&m[1119]))&BiasedRNG[617])|(((m[309]&m[362]&~m[1119]))&~BiasedRNG[617])|((m[309]&m[362]&m[1119]))):InitCond[1003];
    m[559] = run?((((m[323]&~m[363]&m[1184])|(~m[323]&m[363]&m[1184]))&BiasedRNG[618])|(((m[323]&m[363]&~m[1184]))&~BiasedRNG[618])|((m[323]&m[363]&m[1184]))):InitCond[1004];
    m[566] = run?((((m[226]&~m[370]&m[874])|(~m[226]&m[370]&m[874]))&BiasedRNG[619])|(((m[226]&m[370]&~m[874]))&~BiasedRNG[619])|((m[226]&m[370]&m[874]))):InitCond[1005];
    m[567] = run?((((m[240]&~m[371]&m[914])|(~m[240]&m[371]&m[914]))&BiasedRNG[620])|(((m[240]&m[371]&~m[914]))&~BiasedRNG[620])|((m[240]&m[371]&m[914]))):InitCond[1006];
    m[568] = run?((((m[254]&~m[372]&m[959])|(~m[254]&m[372]&m[959]))&BiasedRNG[621])|(((m[254]&m[372]&~m[959]))&~BiasedRNG[621])|((m[254]&m[372]&m[959]))):InitCond[1007];
    m[569] = run?((((m[268]&~m[373]&m[1009])|(~m[268]&m[373]&m[1009]))&BiasedRNG[622])|(((m[268]&m[373]&~m[1009]))&~BiasedRNG[622])|((m[268]&m[373]&m[1009]))):InitCond[1008];
    m[570] = run?((((m[282]&~m[374]&m[1064])|(~m[282]&m[374]&m[1064]))&BiasedRNG[623])|(((m[282]&m[374]&~m[1064]))&~BiasedRNG[623])|((m[282]&m[374]&m[1064]))):InitCond[1009];
    m[571] = run?((((m[296]&~m[375]&m[1124])|(~m[296]&m[375]&m[1124]))&BiasedRNG[624])|(((m[296]&m[375]&~m[1124]))&~BiasedRNG[624])|((m[296]&m[375]&m[1124]))):InitCond[1010];
    m[572] = run?((((m[310]&~m[376]&m[1189])|(~m[310]&m[376]&m[1189]))&BiasedRNG[625])|(((m[310]&m[376]&~m[1189]))&~BiasedRNG[625])|((m[310]&m[376]&m[1189]))):InitCond[1011];
    m[573] = run?((((m[324]&~m[377]&m[1249])|(~m[324]&m[377]&m[1249]))&BiasedRNG[626])|(((m[324]&m[377]&~m[1249]))&~BiasedRNG[626])|((m[324]&m[377]&m[1249]))):InitCond[1012];
    m[580] = run?((((m[227]&~m[384]&m[919])|(~m[227]&m[384]&m[919]))&BiasedRNG[627])|(((m[227]&m[384]&~m[919]))&~BiasedRNG[627])|((m[227]&m[384]&m[919]))):InitCond[1013];
    m[581] = run?((((m[241]&~m[385]&m[964])|(~m[241]&m[385]&m[964]))&BiasedRNG[628])|(((m[241]&m[385]&~m[964]))&~BiasedRNG[628])|((m[241]&m[385]&m[964]))):InitCond[1014];
    m[582] = run?((((m[255]&~m[386]&m[1014])|(~m[255]&m[386]&m[1014]))&BiasedRNG[629])|(((m[255]&m[386]&~m[1014]))&~BiasedRNG[629])|((m[255]&m[386]&m[1014]))):InitCond[1015];
    m[583] = run?((((m[269]&~m[387]&m[1069])|(~m[269]&m[387]&m[1069]))&BiasedRNG[630])|(((m[269]&m[387]&~m[1069]))&~BiasedRNG[630])|((m[269]&m[387]&m[1069]))):InitCond[1016];
    m[584] = run?((((m[283]&~m[388]&m[1129])|(~m[283]&m[388]&m[1129]))&BiasedRNG[631])|(((m[283]&m[388]&~m[1129]))&~BiasedRNG[631])|((m[283]&m[388]&m[1129]))):InitCond[1017];
    m[585] = run?((((m[297]&~m[389]&m[1194])|(~m[297]&m[389]&m[1194]))&BiasedRNG[632])|(((m[297]&m[389]&~m[1194]))&~BiasedRNG[632])|((m[297]&m[389]&m[1194]))):InitCond[1018];
    m[586] = run?((((m[311]&~m[390]&m[1254])|(~m[311]&m[390]&m[1254]))&BiasedRNG[633])|(((m[311]&m[390]&~m[1254]))&~BiasedRNG[633])|((m[311]&m[390]&m[1254]))):InitCond[1019];
    m[587] = run?((((m[325]&~m[391]&m[1309])|(~m[325]&m[391]&m[1309]))&BiasedRNG[634])|(((m[325]&m[391]&~m[1309]))&~BiasedRNG[634])|((m[325]&m[391]&m[1309]))):InitCond[1020];
    m[594] = run?((((m[228]&~m[398]&m[969])|(~m[228]&m[398]&m[969]))&BiasedRNG[635])|(((m[228]&m[398]&~m[969]))&~BiasedRNG[635])|((m[228]&m[398]&m[969]))):InitCond[1021];
    m[595] = run?((((m[242]&~m[399]&m[1019])|(~m[242]&m[399]&m[1019]))&BiasedRNG[636])|(((m[242]&m[399]&~m[1019]))&~BiasedRNG[636])|((m[242]&m[399]&m[1019]))):InitCond[1022];
    m[596] = run?((((m[256]&~m[400]&m[1074])|(~m[256]&m[400]&m[1074]))&BiasedRNG[637])|(((m[256]&m[400]&~m[1074]))&~BiasedRNG[637])|((m[256]&m[400]&m[1074]))):InitCond[1023];
    m[597] = run?((((m[270]&~m[401]&m[1134])|(~m[270]&m[401]&m[1134]))&BiasedRNG[638])|(((m[270]&m[401]&~m[1134]))&~BiasedRNG[638])|((m[270]&m[401]&m[1134]))):InitCond[1024];
    m[598] = run?((((m[284]&~m[402]&m[1199])|(~m[284]&m[402]&m[1199]))&BiasedRNG[639])|(((m[284]&m[402]&~m[1199]))&~BiasedRNG[639])|((m[284]&m[402]&m[1199]))):InitCond[1025];
    m[599] = run?((((m[298]&~m[403]&m[1259])|(~m[298]&m[403]&m[1259]))&BiasedRNG[640])|(((m[298]&m[403]&~m[1259]))&~BiasedRNG[640])|((m[298]&m[403]&m[1259]))):InitCond[1026];
    m[600] = run?((((m[312]&~m[404]&m[1314])|(~m[312]&m[404]&m[1314]))&BiasedRNG[641])|(((m[312]&m[404]&~m[1314]))&~BiasedRNG[641])|((m[312]&m[404]&m[1314]))):InitCond[1027];
    m[601] = run?((((m[326]&~m[405]&m[1364])|(~m[326]&m[405]&m[1364]))&BiasedRNG[642])|(((m[326]&m[405]&~m[1364]))&~BiasedRNG[642])|((m[326]&m[405]&m[1364]))):InitCond[1028];
    m[608] = run?((((m[229]&~m[412]&m[1024])|(~m[229]&m[412]&m[1024]))&BiasedRNG[643])|(((m[229]&m[412]&~m[1024]))&~BiasedRNG[643])|((m[229]&m[412]&m[1024]))):InitCond[1029];
    m[609] = run?((((m[243]&~m[413]&m[1079])|(~m[243]&m[413]&m[1079]))&BiasedRNG[644])|(((m[243]&m[413]&~m[1079]))&~BiasedRNG[644])|((m[243]&m[413]&m[1079]))):InitCond[1030];
    m[610] = run?((((m[257]&~m[414]&m[1139])|(~m[257]&m[414]&m[1139]))&BiasedRNG[645])|(((m[257]&m[414]&~m[1139]))&~BiasedRNG[645])|((m[257]&m[414]&m[1139]))):InitCond[1031];
    m[611] = run?((((m[271]&~m[415]&m[1204])|(~m[271]&m[415]&m[1204]))&BiasedRNG[646])|(((m[271]&m[415]&~m[1204]))&~BiasedRNG[646])|((m[271]&m[415]&m[1204]))):InitCond[1032];
    m[612] = run?((((m[285]&~m[416]&m[1264])|(~m[285]&m[416]&m[1264]))&BiasedRNG[647])|(((m[285]&m[416]&~m[1264]))&~BiasedRNG[647])|((m[285]&m[416]&m[1264]))):InitCond[1033];
    m[613] = run?((((m[299]&~m[417]&m[1319])|(~m[299]&m[417]&m[1319]))&BiasedRNG[648])|(((m[299]&m[417]&~m[1319]))&~BiasedRNG[648])|((m[299]&m[417]&m[1319]))):InitCond[1034];
    m[614] = run?((((m[313]&~m[418]&m[1369])|(~m[313]&m[418]&m[1369]))&BiasedRNG[649])|(((m[313]&m[418]&~m[1369]))&~BiasedRNG[649])|((m[313]&m[418]&m[1369]))):InitCond[1035];
    m[615] = run?((((m[327]&~m[419]&m[1414])|(~m[327]&m[419]&m[1414]))&BiasedRNG[650])|(((m[327]&m[419]&~m[1414]))&~BiasedRNG[650])|((m[327]&m[419]&m[1414]))):InitCond[1036];
    m[616] = run?((((m[146]&~m[420]&m[829])|(~m[146]&m[420]&m[829]))&BiasedRNG[651])|(((m[146]&m[420]&~m[829]))&~BiasedRNG[651])|((m[146]&m[420]&m[829]))):InitCond[1037];
    m[617] = run?((((m[160]&~m[421]&m[859])|(~m[160]&m[421]&m[859]))&BiasedRNG[652])|(((m[160]&m[421]&~m[859]))&~BiasedRNG[652])|((m[160]&m[421]&m[859]))):InitCond[1038];
    m[618] = run?((((m[174]&~m[422]&m[894])|(~m[174]&m[422]&m[894]))&BiasedRNG[653])|(((m[174]&m[422]&~m[894]))&~BiasedRNG[653])|((m[174]&m[422]&m[894]))):InitCond[1039];
    m[619] = run?((((m[188]&~m[423]&m[934])|(~m[188]&m[423]&m[934]))&BiasedRNG[654])|(((m[188]&m[423]&~m[934]))&~BiasedRNG[654])|((m[188]&m[423]&m[934]))):InitCond[1040];
    m[620] = run?((((m[202]&~m[424]&m[979])|(~m[202]&m[424]&m[979]))&BiasedRNG[655])|(((m[202]&m[424]&~m[979]))&~BiasedRNG[655])|((m[202]&m[424]&m[979]))):InitCond[1041];
    m[621] = run?((((m[216]&~m[425]&m[1029])|(~m[216]&m[425]&m[1029]))&BiasedRNG[656])|(((m[216]&m[425]&~m[1029]))&~BiasedRNG[656])|((m[216]&m[425]&m[1029]))):InitCond[1042];
    m[630] = run?((((m[147]&~m[434]&m[864])|(~m[147]&m[434]&m[864]))&BiasedRNG[657])|(((m[147]&m[434]&~m[864]))&~BiasedRNG[657])|((m[147]&m[434]&m[864]))):InitCond[1043];
    m[631] = run?((((m[161]&~m[435]&m[899])|(~m[161]&m[435]&m[899]))&BiasedRNG[658])|(((m[161]&m[435]&~m[899]))&~BiasedRNG[658])|((m[161]&m[435]&m[899]))):InitCond[1044];
    m[632] = run?((((m[175]&~m[436]&m[939])|(~m[175]&m[436]&m[939]))&BiasedRNG[659])|(((m[175]&m[436]&~m[939]))&~BiasedRNG[659])|((m[175]&m[436]&m[939]))):InitCond[1045];
    m[633] = run?((((m[189]&~m[437]&m[984])|(~m[189]&m[437]&m[984]))&BiasedRNG[660])|(((m[189]&m[437]&~m[984]))&~BiasedRNG[660])|((m[189]&m[437]&m[984]))):InitCond[1046];
    m[634] = run?((((m[203]&~m[438]&m[1034])|(~m[203]&m[438]&m[1034]))&BiasedRNG[661])|(((m[203]&m[438]&~m[1034]))&~BiasedRNG[661])|((m[203]&m[438]&m[1034]))):InitCond[1047];
    m[635] = run?((((m[217]&~m[439]&m[1089])|(~m[217]&m[439]&m[1089]))&BiasedRNG[662])|(((m[217]&m[439]&~m[1089]))&~BiasedRNG[662])|((m[217]&m[439]&m[1089]))):InitCond[1048];
    m[644] = run?((((m[148]&~m[448]&m[904])|(~m[148]&m[448]&m[904]))&BiasedRNG[663])|(((m[148]&m[448]&~m[904]))&~BiasedRNG[663])|((m[148]&m[448]&m[904]))):InitCond[1049];
    m[645] = run?((((m[162]&~m[449]&m[944])|(~m[162]&m[449]&m[944]))&BiasedRNG[664])|(((m[162]&m[449]&~m[944]))&~BiasedRNG[664])|((m[162]&m[449]&m[944]))):InitCond[1050];
    m[646] = run?((((m[176]&~m[450]&m[989])|(~m[176]&m[450]&m[989]))&BiasedRNG[665])|(((m[176]&m[450]&~m[989]))&~BiasedRNG[665])|((m[176]&m[450]&m[989]))):InitCond[1051];
    m[647] = run?((((m[190]&~m[451]&m[1039])|(~m[190]&m[451]&m[1039]))&BiasedRNG[666])|(((m[190]&m[451]&~m[1039]))&~BiasedRNG[666])|((m[190]&m[451]&m[1039]))):InitCond[1052];
    m[648] = run?((((m[204]&~m[452]&m[1094])|(~m[204]&m[452]&m[1094]))&BiasedRNG[667])|(((m[204]&m[452]&~m[1094]))&~BiasedRNG[667])|((m[204]&m[452]&m[1094]))):InitCond[1053];
    m[649] = run?((((m[218]&~m[453]&m[1154])|(~m[218]&m[453]&m[1154]))&BiasedRNG[668])|(((m[218]&m[453]&~m[1154]))&~BiasedRNG[668])|((m[218]&m[453]&m[1154]))):InitCond[1054];
    m[658] = run?((((m[149]&~m[462]&m[949])|(~m[149]&m[462]&m[949]))&BiasedRNG[669])|(((m[149]&m[462]&~m[949]))&~BiasedRNG[669])|((m[149]&m[462]&m[949]))):InitCond[1055];
    m[659] = run?((((m[163]&~m[463]&m[994])|(~m[163]&m[463]&m[994]))&BiasedRNG[670])|(((m[163]&m[463]&~m[994]))&~BiasedRNG[670])|((m[163]&m[463]&m[994]))):InitCond[1056];
    m[660] = run?((((m[177]&~m[464]&m[1044])|(~m[177]&m[464]&m[1044]))&BiasedRNG[671])|(((m[177]&m[464]&~m[1044]))&~BiasedRNG[671])|((m[177]&m[464]&m[1044]))):InitCond[1057];
    m[661] = run?((((m[191]&~m[465]&m[1099])|(~m[191]&m[465]&m[1099]))&BiasedRNG[672])|(((m[191]&m[465]&~m[1099]))&~BiasedRNG[672])|((m[191]&m[465]&m[1099]))):InitCond[1058];
    m[662] = run?((((m[205]&~m[466]&m[1159])|(~m[205]&m[466]&m[1159]))&BiasedRNG[673])|(((m[205]&m[466]&~m[1159]))&~BiasedRNG[673])|((m[205]&m[466]&m[1159]))):InitCond[1059];
    m[663] = run?((((m[219]&~m[467]&m[1224])|(~m[219]&m[467]&m[1224]))&BiasedRNG[674])|(((m[219]&m[467]&~m[1224]))&~BiasedRNG[674])|((m[219]&m[467]&m[1224]))):InitCond[1060];
    m[672] = run?((((m[150]&~m[476]&m[999])|(~m[150]&m[476]&m[999]))&BiasedRNG[675])|(((m[150]&m[476]&~m[999]))&~BiasedRNG[675])|((m[150]&m[476]&m[999]))):InitCond[1061];
    m[673] = run?((((m[164]&~m[477]&m[1049])|(~m[164]&m[477]&m[1049]))&BiasedRNG[676])|(((m[164]&m[477]&~m[1049]))&~BiasedRNG[676])|((m[164]&m[477]&m[1049]))):InitCond[1062];
    m[674] = run?((((m[178]&~m[478]&m[1104])|(~m[178]&m[478]&m[1104]))&BiasedRNG[677])|(((m[178]&m[478]&~m[1104]))&~BiasedRNG[677])|((m[178]&m[478]&m[1104]))):InitCond[1063];
    m[675] = run?((((m[192]&~m[479]&m[1164])|(~m[192]&m[479]&m[1164]))&BiasedRNG[678])|(((m[192]&m[479]&~m[1164]))&~BiasedRNG[678])|((m[192]&m[479]&m[1164]))):InitCond[1064];
    m[676] = run?((((m[206]&~m[480]&m[1229])|(~m[206]&m[480]&m[1229]))&BiasedRNG[679])|(((m[206]&m[480]&~m[1229]))&~BiasedRNG[679])|((m[206]&m[480]&m[1229]))):InitCond[1065];
    m[677] = run?((((m[220]&~m[481]&m[1289])|(~m[220]&m[481]&m[1289]))&BiasedRNG[680])|(((m[220]&m[481]&~m[1289]))&~BiasedRNG[680])|((m[220]&m[481]&m[1289]))):InitCond[1066];
    m[686] = run?((((m[151]&~m[490]&m[1054])|(~m[151]&m[490]&m[1054]))&BiasedRNG[681])|(((m[151]&m[490]&~m[1054]))&~BiasedRNG[681])|((m[151]&m[490]&m[1054]))):InitCond[1067];
    m[687] = run?((((m[165]&~m[491]&m[1109])|(~m[165]&m[491]&m[1109]))&BiasedRNG[682])|(((m[165]&m[491]&~m[1109]))&~BiasedRNG[682])|((m[165]&m[491]&m[1109]))):InitCond[1068];
    m[688] = run?((((m[179]&~m[492]&m[1169])|(~m[179]&m[492]&m[1169]))&BiasedRNG[683])|(((m[179]&m[492]&~m[1169]))&~BiasedRNG[683])|((m[179]&m[492]&m[1169]))):InitCond[1069];
    m[689] = run?((((m[193]&~m[493]&m[1234])|(~m[193]&m[493]&m[1234]))&BiasedRNG[684])|(((m[193]&m[493]&~m[1234]))&~BiasedRNG[684])|((m[193]&m[493]&m[1234]))):InitCond[1070];
    m[690] = run?((((m[207]&~m[494]&m[1294])|(~m[207]&m[494]&m[1294]))&BiasedRNG[685])|(((m[207]&m[494]&~m[1294]))&~BiasedRNG[685])|((m[207]&m[494]&m[1294]))):InitCond[1071];
    m[691] = run?((((m[221]&~m[495]&m[1349])|(~m[221]&m[495]&m[1349]))&BiasedRNG[686])|(((m[221]&m[495]&~m[1349]))&~BiasedRNG[686])|((m[221]&m[495]&m[1349]))):InitCond[1072];
    m[700] = run?((((m[152]&~m[504]&m[1114])|(~m[152]&m[504]&m[1114]))&BiasedRNG[687])|(((m[152]&m[504]&~m[1114]))&~BiasedRNG[687])|((m[152]&m[504]&m[1114]))):InitCond[1073];
    m[701] = run?((((m[166]&~m[505]&m[1174])|(~m[166]&m[505]&m[1174]))&BiasedRNG[688])|(((m[166]&m[505]&~m[1174]))&~BiasedRNG[688])|((m[166]&m[505]&m[1174]))):InitCond[1074];
    m[702] = run?((((m[180]&~m[506]&m[1239])|(~m[180]&m[506]&m[1239]))&BiasedRNG[689])|(((m[180]&m[506]&~m[1239]))&~BiasedRNG[689])|((m[180]&m[506]&m[1239]))):InitCond[1075];
    m[703] = run?((((m[194]&~m[507]&m[1299])|(~m[194]&m[507]&m[1299]))&BiasedRNG[690])|(((m[194]&m[507]&~m[1299]))&~BiasedRNG[690])|((m[194]&m[507]&m[1299]))):InitCond[1076];
    m[704] = run?((((m[208]&~m[508]&m[1354])|(~m[208]&m[508]&m[1354]))&BiasedRNG[691])|(((m[208]&m[508]&~m[1354]))&~BiasedRNG[691])|((m[208]&m[508]&m[1354]))):InitCond[1077];
    m[705] = run?((((m[222]&~m[509]&m[1404])|(~m[222]&m[509]&m[1404]))&BiasedRNG[692])|(((m[222]&m[509]&~m[1404]))&~BiasedRNG[692])|((m[222]&m[509]&m[1404]))):InitCond[1078];
    m[714] = run?((((m[153]&~m[518]&m[1179])|(~m[153]&m[518]&m[1179]))&BiasedRNG[693])|(((m[153]&m[518]&~m[1179]))&~BiasedRNG[693])|((m[153]&m[518]&m[1179]))):InitCond[1079];
    m[715] = run?((((m[167]&~m[519]&m[1244])|(~m[167]&m[519]&m[1244]))&BiasedRNG[694])|(((m[167]&m[519]&~m[1244]))&~BiasedRNG[694])|((m[167]&m[519]&m[1244]))):InitCond[1080];
    m[716] = run?((((m[181]&~m[520]&m[1304])|(~m[181]&m[520]&m[1304]))&BiasedRNG[695])|(((m[181]&m[520]&~m[1304]))&~BiasedRNG[695])|((m[181]&m[520]&m[1304]))):InitCond[1081];
    m[717] = run?((((m[195]&~m[521]&m[1359])|(~m[195]&m[521]&m[1359]))&BiasedRNG[696])|(((m[195]&m[521]&~m[1359]))&~BiasedRNG[696])|((m[195]&m[521]&m[1359]))):InitCond[1082];
    m[718] = run?((((m[209]&~m[522]&m[1409])|(~m[209]&m[522]&m[1409]))&BiasedRNG[697])|(((m[209]&m[522]&~m[1409]))&~BiasedRNG[697])|((m[209]&m[522]&m[1409]))):InitCond[1083];
    m[719] = run?((((m[223]&~m[523]&m[1454])|(~m[223]&m[523]&m[1454]))&BiasedRNG[698])|(((m[223]&m[523]&~m[1454]))&~BiasedRNG[698])|((m[223]&m[523]&m[1454]))):InitCond[1084];
    m[729] = run?((((m[546]&~m[728]&~m[730]&~m[731]&~m[732])|(~m[546]&~m[728]&~m[730]&m[731]&~m[732])|(m[546]&m[728]&~m[730]&m[731]&~m[732])|(m[546]&~m[728]&m[730]&m[731]&~m[732])|(~m[546]&m[728]&~m[730]&~m[731]&m[732])|(~m[546]&~m[728]&m[730]&~m[731]&m[732])|(m[546]&m[728]&m[730]&~m[731]&m[732])|(~m[546]&m[728]&m[730]&m[731]&m[732]))&UnbiasedRNG[386])|((m[546]&~m[728]&~m[730]&m[731]&~m[732])|(~m[546]&~m[728]&~m[730]&~m[731]&m[732])|(m[546]&~m[728]&~m[730]&~m[731]&m[732])|(m[546]&m[728]&~m[730]&~m[731]&m[732])|(m[546]&~m[728]&m[730]&~m[731]&m[732])|(~m[546]&~m[728]&~m[730]&m[731]&m[732])|(m[546]&~m[728]&~m[730]&m[731]&m[732])|(~m[546]&m[728]&~m[730]&m[731]&m[732])|(m[546]&m[728]&~m[730]&m[731]&m[732])|(~m[546]&~m[728]&m[730]&m[731]&m[732])|(m[546]&~m[728]&m[730]&m[731]&m[732])|(m[546]&m[728]&m[730]&m[731]&m[732]))):InitCond[1085];
    m[734] = run?((((m[547]&~m[733]&~m[735]&~m[736]&~m[737])|(~m[547]&~m[733]&~m[735]&m[736]&~m[737])|(m[547]&m[733]&~m[735]&m[736]&~m[737])|(m[547]&~m[733]&m[735]&m[736]&~m[737])|(~m[547]&m[733]&~m[735]&~m[736]&m[737])|(~m[547]&~m[733]&m[735]&~m[736]&m[737])|(m[547]&m[733]&m[735]&~m[736]&m[737])|(~m[547]&m[733]&m[735]&m[736]&m[737]))&UnbiasedRNG[387])|((m[547]&~m[733]&~m[735]&m[736]&~m[737])|(~m[547]&~m[733]&~m[735]&~m[736]&m[737])|(m[547]&~m[733]&~m[735]&~m[736]&m[737])|(m[547]&m[733]&~m[735]&~m[736]&m[737])|(m[547]&~m[733]&m[735]&~m[736]&m[737])|(~m[547]&~m[733]&~m[735]&m[736]&m[737])|(m[547]&~m[733]&~m[735]&m[736]&m[737])|(~m[547]&m[733]&~m[735]&m[736]&m[737])|(m[547]&m[733]&~m[735]&m[736]&m[737])|(~m[547]&~m[733]&m[735]&m[736]&m[737])|(m[547]&~m[733]&m[735]&m[736]&m[737])|(m[547]&m[733]&m[735]&m[736]&m[737]))):InitCond[1086];
    m[739] = run?((((m[560]&~m[738]&~m[740]&~m[741]&~m[742])|(~m[560]&~m[738]&~m[740]&m[741]&~m[742])|(m[560]&m[738]&~m[740]&m[741]&~m[742])|(m[560]&~m[738]&m[740]&m[741]&~m[742])|(~m[560]&m[738]&~m[740]&~m[741]&m[742])|(~m[560]&~m[738]&m[740]&~m[741]&m[742])|(m[560]&m[738]&m[740]&~m[741]&m[742])|(~m[560]&m[738]&m[740]&m[741]&m[742]))&UnbiasedRNG[388])|((m[560]&~m[738]&~m[740]&m[741]&~m[742])|(~m[560]&~m[738]&~m[740]&~m[741]&m[742])|(m[560]&~m[738]&~m[740]&~m[741]&m[742])|(m[560]&m[738]&~m[740]&~m[741]&m[742])|(m[560]&~m[738]&m[740]&~m[741]&m[742])|(~m[560]&~m[738]&~m[740]&m[741]&m[742])|(m[560]&~m[738]&~m[740]&m[741]&m[742])|(~m[560]&m[738]&~m[740]&m[741]&m[742])|(m[560]&m[738]&~m[740]&m[741]&m[742])|(~m[560]&~m[738]&m[740]&m[741]&m[742])|(m[560]&~m[738]&m[740]&m[741]&m[742])|(m[560]&m[738]&m[740]&m[741]&m[742]))):InitCond[1087];
    m[744] = run?((((m[548]&~m[743]&~m[745]&~m[746]&~m[747])|(~m[548]&~m[743]&~m[745]&m[746]&~m[747])|(m[548]&m[743]&~m[745]&m[746]&~m[747])|(m[548]&~m[743]&m[745]&m[746]&~m[747])|(~m[548]&m[743]&~m[745]&~m[746]&m[747])|(~m[548]&~m[743]&m[745]&~m[746]&m[747])|(m[548]&m[743]&m[745]&~m[746]&m[747])|(~m[548]&m[743]&m[745]&m[746]&m[747]))&UnbiasedRNG[389])|((m[548]&~m[743]&~m[745]&m[746]&~m[747])|(~m[548]&~m[743]&~m[745]&~m[746]&m[747])|(m[548]&~m[743]&~m[745]&~m[746]&m[747])|(m[548]&m[743]&~m[745]&~m[746]&m[747])|(m[548]&~m[743]&m[745]&~m[746]&m[747])|(~m[548]&~m[743]&~m[745]&m[746]&m[747])|(m[548]&~m[743]&~m[745]&m[746]&m[747])|(~m[548]&m[743]&~m[745]&m[746]&m[747])|(m[548]&m[743]&~m[745]&m[746]&m[747])|(~m[548]&~m[743]&m[745]&m[746]&m[747])|(m[548]&~m[743]&m[745]&m[746]&m[747])|(m[548]&m[743]&m[745]&m[746]&m[747]))):InitCond[1088];
    m[749] = run?((((m[561]&~m[748]&~m[750]&~m[751]&~m[752])|(~m[561]&~m[748]&~m[750]&m[751]&~m[752])|(m[561]&m[748]&~m[750]&m[751]&~m[752])|(m[561]&~m[748]&m[750]&m[751]&~m[752])|(~m[561]&m[748]&~m[750]&~m[751]&m[752])|(~m[561]&~m[748]&m[750]&~m[751]&m[752])|(m[561]&m[748]&m[750]&~m[751]&m[752])|(~m[561]&m[748]&m[750]&m[751]&m[752]))&UnbiasedRNG[390])|((m[561]&~m[748]&~m[750]&m[751]&~m[752])|(~m[561]&~m[748]&~m[750]&~m[751]&m[752])|(m[561]&~m[748]&~m[750]&~m[751]&m[752])|(m[561]&m[748]&~m[750]&~m[751]&m[752])|(m[561]&~m[748]&m[750]&~m[751]&m[752])|(~m[561]&~m[748]&~m[750]&m[751]&m[752])|(m[561]&~m[748]&~m[750]&m[751]&m[752])|(~m[561]&m[748]&~m[750]&m[751]&m[752])|(m[561]&m[748]&~m[750]&m[751]&m[752])|(~m[561]&~m[748]&m[750]&m[751]&m[752])|(m[561]&~m[748]&m[750]&m[751]&m[752])|(m[561]&m[748]&m[750]&m[751]&m[752]))):InitCond[1089];
    m[754] = run?((((m[574]&~m[753]&~m[755]&~m[756]&~m[757])|(~m[574]&~m[753]&~m[755]&m[756]&~m[757])|(m[574]&m[753]&~m[755]&m[756]&~m[757])|(m[574]&~m[753]&m[755]&m[756]&~m[757])|(~m[574]&m[753]&~m[755]&~m[756]&m[757])|(~m[574]&~m[753]&m[755]&~m[756]&m[757])|(m[574]&m[753]&m[755]&~m[756]&m[757])|(~m[574]&m[753]&m[755]&m[756]&m[757]))&UnbiasedRNG[391])|((m[574]&~m[753]&~m[755]&m[756]&~m[757])|(~m[574]&~m[753]&~m[755]&~m[756]&m[757])|(m[574]&~m[753]&~m[755]&~m[756]&m[757])|(m[574]&m[753]&~m[755]&~m[756]&m[757])|(m[574]&~m[753]&m[755]&~m[756]&m[757])|(~m[574]&~m[753]&~m[755]&m[756]&m[757])|(m[574]&~m[753]&~m[755]&m[756]&m[757])|(~m[574]&m[753]&~m[755]&m[756]&m[757])|(m[574]&m[753]&~m[755]&m[756]&m[757])|(~m[574]&~m[753]&m[755]&m[756]&m[757])|(m[574]&~m[753]&m[755]&m[756]&m[757])|(m[574]&m[753]&m[755]&m[756]&m[757]))):InitCond[1090];
    m[759] = run?((((m[549]&~m[758]&~m[760]&~m[761]&~m[762])|(~m[549]&~m[758]&~m[760]&m[761]&~m[762])|(m[549]&m[758]&~m[760]&m[761]&~m[762])|(m[549]&~m[758]&m[760]&m[761]&~m[762])|(~m[549]&m[758]&~m[760]&~m[761]&m[762])|(~m[549]&~m[758]&m[760]&~m[761]&m[762])|(m[549]&m[758]&m[760]&~m[761]&m[762])|(~m[549]&m[758]&m[760]&m[761]&m[762]))&UnbiasedRNG[392])|((m[549]&~m[758]&~m[760]&m[761]&~m[762])|(~m[549]&~m[758]&~m[760]&~m[761]&m[762])|(m[549]&~m[758]&~m[760]&~m[761]&m[762])|(m[549]&m[758]&~m[760]&~m[761]&m[762])|(m[549]&~m[758]&m[760]&~m[761]&m[762])|(~m[549]&~m[758]&~m[760]&m[761]&m[762])|(m[549]&~m[758]&~m[760]&m[761]&m[762])|(~m[549]&m[758]&~m[760]&m[761]&m[762])|(m[549]&m[758]&~m[760]&m[761]&m[762])|(~m[549]&~m[758]&m[760]&m[761]&m[762])|(m[549]&~m[758]&m[760]&m[761]&m[762])|(m[549]&m[758]&m[760]&m[761]&m[762]))):InitCond[1091];
    m[764] = run?((((m[562]&~m[763]&~m[765]&~m[766]&~m[767])|(~m[562]&~m[763]&~m[765]&m[766]&~m[767])|(m[562]&m[763]&~m[765]&m[766]&~m[767])|(m[562]&~m[763]&m[765]&m[766]&~m[767])|(~m[562]&m[763]&~m[765]&~m[766]&m[767])|(~m[562]&~m[763]&m[765]&~m[766]&m[767])|(m[562]&m[763]&m[765]&~m[766]&m[767])|(~m[562]&m[763]&m[765]&m[766]&m[767]))&UnbiasedRNG[393])|((m[562]&~m[763]&~m[765]&m[766]&~m[767])|(~m[562]&~m[763]&~m[765]&~m[766]&m[767])|(m[562]&~m[763]&~m[765]&~m[766]&m[767])|(m[562]&m[763]&~m[765]&~m[766]&m[767])|(m[562]&~m[763]&m[765]&~m[766]&m[767])|(~m[562]&~m[763]&~m[765]&m[766]&m[767])|(m[562]&~m[763]&~m[765]&m[766]&m[767])|(~m[562]&m[763]&~m[765]&m[766]&m[767])|(m[562]&m[763]&~m[765]&m[766]&m[767])|(~m[562]&~m[763]&m[765]&m[766]&m[767])|(m[562]&~m[763]&m[765]&m[766]&m[767])|(m[562]&m[763]&m[765]&m[766]&m[767]))):InitCond[1092];
    m[769] = run?((((m[575]&~m[768]&~m[770]&~m[771]&~m[772])|(~m[575]&~m[768]&~m[770]&m[771]&~m[772])|(m[575]&m[768]&~m[770]&m[771]&~m[772])|(m[575]&~m[768]&m[770]&m[771]&~m[772])|(~m[575]&m[768]&~m[770]&~m[771]&m[772])|(~m[575]&~m[768]&m[770]&~m[771]&m[772])|(m[575]&m[768]&m[770]&~m[771]&m[772])|(~m[575]&m[768]&m[770]&m[771]&m[772]))&UnbiasedRNG[394])|((m[575]&~m[768]&~m[770]&m[771]&~m[772])|(~m[575]&~m[768]&~m[770]&~m[771]&m[772])|(m[575]&~m[768]&~m[770]&~m[771]&m[772])|(m[575]&m[768]&~m[770]&~m[771]&m[772])|(m[575]&~m[768]&m[770]&~m[771]&m[772])|(~m[575]&~m[768]&~m[770]&m[771]&m[772])|(m[575]&~m[768]&~m[770]&m[771]&m[772])|(~m[575]&m[768]&~m[770]&m[771]&m[772])|(m[575]&m[768]&~m[770]&m[771]&m[772])|(~m[575]&~m[768]&m[770]&m[771]&m[772])|(m[575]&~m[768]&m[770]&m[771]&m[772])|(m[575]&m[768]&m[770]&m[771]&m[772]))):InitCond[1093];
    m[774] = run?((((m[588]&~m[773]&~m[775]&~m[776]&~m[777])|(~m[588]&~m[773]&~m[775]&m[776]&~m[777])|(m[588]&m[773]&~m[775]&m[776]&~m[777])|(m[588]&~m[773]&m[775]&m[776]&~m[777])|(~m[588]&m[773]&~m[775]&~m[776]&m[777])|(~m[588]&~m[773]&m[775]&~m[776]&m[777])|(m[588]&m[773]&m[775]&~m[776]&m[777])|(~m[588]&m[773]&m[775]&m[776]&m[777]))&UnbiasedRNG[395])|((m[588]&~m[773]&~m[775]&m[776]&~m[777])|(~m[588]&~m[773]&~m[775]&~m[776]&m[777])|(m[588]&~m[773]&~m[775]&~m[776]&m[777])|(m[588]&m[773]&~m[775]&~m[776]&m[777])|(m[588]&~m[773]&m[775]&~m[776]&m[777])|(~m[588]&~m[773]&~m[775]&m[776]&m[777])|(m[588]&~m[773]&~m[775]&m[776]&m[777])|(~m[588]&m[773]&~m[775]&m[776]&m[777])|(m[588]&m[773]&~m[775]&m[776]&m[777])|(~m[588]&~m[773]&m[775]&m[776]&m[777])|(m[588]&~m[773]&m[775]&m[776]&m[777])|(m[588]&m[773]&m[775]&m[776]&m[777]))):InitCond[1094];
    m[779] = run?((((m[550]&~m[778]&~m[780]&~m[781]&~m[782])|(~m[550]&~m[778]&~m[780]&m[781]&~m[782])|(m[550]&m[778]&~m[780]&m[781]&~m[782])|(m[550]&~m[778]&m[780]&m[781]&~m[782])|(~m[550]&m[778]&~m[780]&~m[781]&m[782])|(~m[550]&~m[778]&m[780]&~m[781]&m[782])|(m[550]&m[778]&m[780]&~m[781]&m[782])|(~m[550]&m[778]&m[780]&m[781]&m[782]))&UnbiasedRNG[396])|((m[550]&~m[778]&~m[780]&m[781]&~m[782])|(~m[550]&~m[778]&~m[780]&~m[781]&m[782])|(m[550]&~m[778]&~m[780]&~m[781]&m[782])|(m[550]&m[778]&~m[780]&~m[781]&m[782])|(m[550]&~m[778]&m[780]&~m[781]&m[782])|(~m[550]&~m[778]&~m[780]&m[781]&m[782])|(m[550]&~m[778]&~m[780]&m[781]&m[782])|(~m[550]&m[778]&~m[780]&m[781]&m[782])|(m[550]&m[778]&~m[780]&m[781]&m[782])|(~m[550]&~m[778]&m[780]&m[781]&m[782])|(m[550]&~m[778]&m[780]&m[781]&m[782])|(m[550]&m[778]&m[780]&m[781]&m[782]))):InitCond[1095];
    m[784] = run?((((m[563]&~m[783]&~m[785]&~m[786]&~m[787])|(~m[563]&~m[783]&~m[785]&m[786]&~m[787])|(m[563]&m[783]&~m[785]&m[786]&~m[787])|(m[563]&~m[783]&m[785]&m[786]&~m[787])|(~m[563]&m[783]&~m[785]&~m[786]&m[787])|(~m[563]&~m[783]&m[785]&~m[786]&m[787])|(m[563]&m[783]&m[785]&~m[786]&m[787])|(~m[563]&m[783]&m[785]&m[786]&m[787]))&UnbiasedRNG[397])|((m[563]&~m[783]&~m[785]&m[786]&~m[787])|(~m[563]&~m[783]&~m[785]&~m[786]&m[787])|(m[563]&~m[783]&~m[785]&~m[786]&m[787])|(m[563]&m[783]&~m[785]&~m[786]&m[787])|(m[563]&~m[783]&m[785]&~m[786]&m[787])|(~m[563]&~m[783]&~m[785]&m[786]&m[787])|(m[563]&~m[783]&~m[785]&m[786]&m[787])|(~m[563]&m[783]&~m[785]&m[786]&m[787])|(m[563]&m[783]&~m[785]&m[786]&m[787])|(~m[563]&~m[783]&m[785]&m[786]&m[787])|(m[563]&~m[783]&m[785]&m[786]&m[787])|(m[563]&m[783]&m[785]&m[786]&m[787]))):InitCond[1096];
    m[789] = run?((((m[576]&~m[788]&~m[790]&~m[791]&~m[792])|(~m[576]&~m[788]&~m[790]&m[791]&~m[792])|(m[576]&m[788]&~m[790]&m[791]&~m[792])|(m[576]&~m[788]&m[790]&m[791]&~m[792])|(~m[576]&m[788]&~m[790]&~m[791]&m[792])|(~m[576]&~m[788]&m[790]&~m[791]&m[792])|(m[576]&m[788]&m[790]&~m[791]&m[792])|(~m[576]&m[788]&m[790]&m[791]&m[792]))&UnbiasedRNG[398])|((m[576]&~m[788]&~m[790]&m[791]&~m[792])|(~m[576]&~m[788]&~m[790]&~m[791]&m[792])|(m[576]&~m[788]&~m[790]&~m[791]&m[792])|(m[576]&m[788]&~m[790]&~m[791]&m[792])|(m[576]&~m[788]&m[790]&~m[791]&m[792])|(~m[576]&~m[788]&~m[790]&m[791]&m[792])|(m[576]&~m[788]&~m[790]&m[791]&m[792])|(~m[576]&m[788]&~m[790]&m[791]&m[792])|(m[576]&m[788]&~m[790]&m[791]&m[792])|(~m[576]&~m[788]&m[790]&m[791]&m[792])|(m[576]&~m[788]&m[790]&m[791]&m[792])|(m[576]&m[788]&m[790]&m[791]&m[792]))):InitCond[1097];
    m[794] = run?((((m[589]&~m[793]&~m[795]&~m[796]&~m[797])|(~m[589]&~m[793]&~m[795]&m[796]&~m[797])|(m[589]&m[793]&~m[795]&m[796]&~m[797])|(m[589]&~m[793]&m[795]&m[796]&~m[797])|(~m[589]&m[793]&~m[795]&~m[796]&m[797])|(~m[589]&~m[793]&m[795]&~m[796]&m[797])|(m[589]&m[793]&m[795]&~m[796]&m[797])|(~m[589]&m[793]&m[795]&m[796]&m[797]))&UnbiasedRNG[399])|((m[589]&~m[793]&~m[795]&m[796]&~m[797])|(~m[589]&~m[793]&~m[795]&~m[796]&m[797])|(m[589]&~m[793]&~m[795]&~m[796]&m[797])|(m[589]&m[793]&~m[795]&~m[796]&m[797])|(m[589]&~m[793]&m[795]&~m[796]&m[797])|(~m[589]&~m[793]&~m[795]&m[796]&m[797])|(m[589]&~m[793]&~m[795]&m[796]&m[797])|(~m[589]&m[793]&~m[795]&m[796]&m[797])|(m[589]&m[793]&~m[795]&m[796]&m[797])|(~m[589]&~m[793]&m[795]&m[796]&m[797])|(m[589]&~m[793]&m[795]&m[796]&m[797])|(m[589]&m[793]&m[795]&m[796]&m[797]))):InitCond[1098];
    m[799] = run?((((m[602]&~m[798]&~m[800]&~m[801]&~m[802])|(~m[602]&~m[798]&~m[800]&m[801]&~m[802])|(m[602]&m[798]&~m[800]&m[801]&~m[802])|(m[602]&~m[798]&m[800]&m[801]&~m[802])|(~m[602]&m[798]&~m[800]&~m[801]&m[802])|(~m[602]&~m[798]&m[800]&~m[801]&m[802])|(m[602]&m[798]&m[800]&~m[801]&m[802])|(~m[602]&m[798]&m[800]&m[801]&m[802]))&UnbiasedRNG[400])|((m[602]&~m[798]&~m[800]&m[801]&~m[802])|(~m[602]&~m[798]&~m[800]&~m[801]&m[802])|(m[602]&~m[798]&~m[800]&~m[801]&m[802])|(m[602]&m[798]&~m[800]&~m[801]&m[802])|(m[602]&~m[798]&m[800]&~m[801]&m[802])|(~m[602]&~m[798]&~m[800]&m[801]&m[802])|(m[602]&~m[798]&~m[800]&m[801]&m[802])|(~m[602]&m[798]&~m[800]&m[801]&m[802])|(m[602]&m[798]&~m[800]&m[801]&m[802])|(~m[602]&~m[798]&m[800]&m[801]&m[802])|(m[602]&~m[798]&m[800]&m[801]&m[802])|(m[602]&m[798]&m[800]&m[801]&m[802]))):InitCond[1099];
    m[804] = run?((((m[551]&~m[803]&~m[805]&~m[806]&~m[807])|(~m[551]&~m[803]&~m[805]&m[806]&~m[807])|(m[551]&m[803]&~m[805]&m[806]&~m[807])|(m[551]&~m[803]&m[805]&m[806]&~m[807])|(~m[551]&m[803]&~m[805]&~m[806]&m[807])|(~m[551]&~m[803]&m[805]&~m[806]&m[807])|(m[551]&m[803]&m[805]&~m[806]&m[807])|(~m[551]&m[803]&m[805]&m[806]&m[807]))&UnbiasedRNG[401])|((m[551]&~m[803]&~m[805]&m[806]&~m[807])|(~m[551]&~m[803]&~m[805]&~m[806]&m[807])|(m[551]&~m[803]&~m[805]&~m[806]&m[807])|(m[551]&m[803]&~m[805]&~m[806]&m[807])|(m[551]&~m[803]&m[805]&~m[806]&m[807])|(~m[551]&~m[803]&~m[805]&m[806]&m[807])|(m[551]&~m[803]&~m[805]&m[806]&m[807])|(~m[551]&m[803]&~m[805]&m[806]&m[807])|(m[551]&m[803]&~m[805]&m[806]&m[807])|(~m[551]&~m[803]&m[805]&m[806]&m[807])|(m[551]&~m[803]&m[805]&m[806]&m[807])|(m[551]&m[803]&m[805]&m[806]&m[807]))):InitCond[1100];
    m[809] = run?((((m[564]&~m[808]&~m[810]&~m[811]&~m[812])|(~m[564]&~m[808]&~m[810]&m[811]&~m[812])|(m[564]&m[808]&~m[810]&m[811]&~m[812])|(m[564]&~m[808]&m[810]&m[811]&~m[812])|(~m[564]&m[808]&~m[810]&~m[811]&m[812])|(~m[564]&~m[808]&m[810]&~m[811]&m[812])|(m[564]&m[808]&m[810]&~m[811]&m[812])|(~m[564]&m[808]&m[810]&m[811]&m[812]))&UnbiasedRNG[402])|((m[564]&~m[808]&~m[810]&m[811]&~m[812])|(~m[564]&~m[808]&~m[810]&~m[811]&m[812])|(m[564]&~m[808]&~m[810]&~m[811]&m[812])|(m[564]&m[808]&~m[810]&~m[811]&m[812])|(m[564]&~m[808]&m[810]&~m[811]&m[812])|(~m[564]&~m[808]&~m[810]&m[811]&m[812])|(m[564]&~m[808]&~m[810]&m[811]&m[812])|(~m[564]&m[808]&~m[810]&m[811]&m[812])|(m[564]&m[808]&~m[810]&m[811]&m[812])|(~m[564]&~m[808]&m[810]&m[811]&m[812])|(m[564]&~m[808]&m[810]&m[811]&m[812])|(m[564]&m[808]&m[810]&m[811]&m[812]))):InitCond[1101];
    m[814] = run?((((m[577]&~m[813]&~m[815]&~m[816]&~m[817])|(~m[577]&~m[813]&~m[815]&m[816]&~m[817])|(m[577]&m[813]&~m[815]&m[816]&~m[817])|(m[577]&~m[813]&m[815]&m[816]&~m[817])|(~m[577]&m[813]&~m[815]&~m[816]&m[817])|(~m[577]&~m[813]&m[815]&~m[816]&m[817])|(m[577]&m[813]&m[815]&~m[816]&m[817])|(~m[577]&m[813]&m[815]&m[816]&m[817]))&UnbiasedRNG[403])|((m[577]&~m[813]&~m[815]&m[816]&~m[817])|(~m[577]&~m[813]&~m[815]&~m[816]&m[817])|(m[577]&~m[813]&~m[815]&~m[816]&m[817])|(m[577]&m[813]&~m[815]&~m[816]&m[817])|(m[577]&~m[813]&m[815]&~m[816]&m[817])|(~m[577]&~m[813]&~m[815]&m[816]&m[817])|(m[577]&~m[813]&~m[815]&m[816]&m[817])|(~m[577]&m[813]&~m[815]&m[816]&m[817])|(m[577]&m[813]&~m[815]&m[816]&m[817])|(~m[577]&~m[813]&m[815]&m[816]&m[817])|(m[577]&~m[813]&m[815]&m[816]&m[817])|(m[577]&m[813]&m[815]&m[816]&m[817]))):InitCond[1102];
    m[819] = run?((((m[590]&~m[818]&~m[820]&~m[821]&~m[822])|(~m[590]&~m[818]&~m[820]&m[821]&~m[822])|(m[590]&m[818]&~m[820]&m[821]&~m[822])|(m[590]&~m[818]&m[820]&m[821]&~m[822])|(~m[590]&m[818]&~m[820]&~m[821]&m[822])|(~m[590]&~m[818]&m[820]&~m[821]&m[822])|(m[590]&m[818]&m[820]&~m[821]&m[822])|(~m[590]&m[818]&m[820]&m[821]&m[822]))&UnbiasedRNG[404])|((m[590]&~m[818]&~m[820]&m[821]&~m[822])|(~m[590]&~m[818]&~m[820]&~m[821]&m[822])|(m[590]&~m[818]&~m[820]&~m[821]&m[822])|(m[590]&m[818]&~m[820]&~m[821]&m[822])|(m[590]&~m[818]&m[820]&~m[821]&m[822])|(~m[590]&~m[818]&~m[820]&m[821]&m[822])|(m[590]&~m[818]&~m[820]&m[821]&m[822])|(~m[590]&m[818]&~m[820]&m[821]&m[822])|(m[590]&m[818]&~m[820]&m[821]&m[822])|(~m[590]&~m[818]&m[820]&m[821]&m[822])|(m[590]&~m[818]&m[820]&m[821]&m[822])|(m[590]&m[818]&m[820]&m[821]&m[822]))):InitCond[1103];
    m[824] = run?((((m[603]&~m[823]&~m[825]&~m[826]&~m[827])|(~m[603]&~m[823]&~m[825]&m[826]&~m[827])|(m[603]&m[823]&~m[825]&m[826]&~m[827])|(m[603]&~m[823]&m[825]&m[826]&~m[827])|(~m[603]&m[823]&~m[825]&~m[826]&m[827])|(~m[603]&~m[823]&m[825]&~m[826]&m[827])|(m[603]&m[823]&m[825]&~m[826]&m[827])|(~m[603]&m[823]&m[825]&m[826]&m[827]))&UnbiasedRNG[405])|((m[603]&~m[823]&~m[825]&m[826]&~m[827])|(~m[603]&~m[823]&~m[825]&~m[826]&m[827])|(m[603]&~m[823]&~m[825]&~m[826]&m[827])|(m[603]&m[823]&~m[825]&~m[826]&m[827])|(m[603]&~m[823]&m[825]&~m[826]&m[827])|(~m[603]&~m[823]&~m[825]&m[826]&m[827])|(m[603]&~m[823]&~m[825]&m[826]&m[827])|(~m[603]&m[823]&~m[825]&m[826]&m[827])|(m[603]&m[823]&~m[825]&m[826]&m[827])|(~m[603]&~m[823]&m[825]&m[826]&m[827])|(m[603]&~m[823]&m[825]&m[826]&m[827])|(m[603]&m[823]&m[825]&m[826]&m[827]))):InitCond[1104];
    m[835] = run?((((m[807]&~m[833]&~m[834]&~m[836]&~m[837])|(~m[807]&~m[833]&~m[834]&m[836]&~m[837])|(m[807]&m[833]&~m[834]&m[836]&~m[837])|(m[807]&~m[833]&m[834]&m[836]&~m[837])|(~m[807]&m[833]&~m[834]&~m[836]&m[837])|(~m[807]&~m[833]&m[834]&~m[836]&m[837])|(m[807]&m[833]&m[834]&~m[836]&m[837])|(~m[807]&m[833]&m[834]&m[836]&m[837]))&UnbiasedRNG[406])|((m[807]&~m[833]&~m[834]&m[836]&~m[837])|(~m[807]&~m[833]&~m[834]&~m[836]&m[837])|(m[807]&~m[833]&~m[834]&~m[836]&m[837])|(m[807]&m[833]&~m[834]&~m[836]&m[837])|(m[807]&~m[833]&m[834]&~m[836]&m[837])|(~m[807]&~m[833]&~m[834]&m[836]&m[837])|(m[807]&~m[833]&~m[834]&m[836]&m[837])|(~m[807]&m[833]&~m[834]&m[836]&m[837])|(m[807]&m[833]&~m[834]&m[836]&m[837])|(~m[807]&~m[833]&m[834]&m[836]&m[837])|(m[807]&~m[833]&m[834]&m[836]&m[837])|(m[807]&m[833]&m[834]&m[836]&m[837]))):InitCond[1105];
    m[839] = run?((((m[565]&~m[838]&~m[840]&~m[841]&~m[842])|(~m[565]&~m[838]&~m[840]&m[841]&~m[842])|(m[565]&m[838]&~m[840]&m[841]&~m[842])|(m[565]&~m[838]&m[840]&m[841]&~m[842])|(~m[565]&m[838]&~m[840]&~m[841]&m[842])|(~m[565]&~m[838]&m[840]&~m[841]&m[842])|(m[565]&m[838]&m[840]&~m[841]&m[842])|(~m[565]&m[838]&m[840]&m[841]&m[842]))&UnbiasedRNG[407])|((m[565]&~m[838]&~m[840]&m[841]&~m[842])|(~m[565]&~m[838]&~m[840]&~m[841]&m[842])|(m[565]&~m[838]&~m[840]&~m[841]&m[842])|(m[565]&m[838]&~m[840]&~m[841]&m[842])|(m[565]&~m[838]&m[840]&~m[841]&m[842])|(~m[565]&~m[838]&~m[840]&m[841]&m[842])|(m[565]&~m[838]&~m[840]&m[841]&m[842])|(~m[565]&m[838]&~m[840]&m[841]&m[842])|(m[565]&m[838]&~m[840]&m[841]&m[842])|(~m[565]&~m[838]&m[840]&m[841]&m[842])|(m[565]&~m[838]&m[840]&m[841]&m[842])|(m[565]&m[838]&m[840]&m[841]&m[842]))):InitCond[1106];
    m[844] = run?((((m[578]&~m[843]&~m[845]&~m[846]&~m[847])|(~m[578]&~m[843]&~m[845]&m[846]&~m[847])|(m[578]&m[843]&~m[845]&m[846]&~m[847])|(m[578]&~m[843]&m[845]&m[846]&~m[847])|(~m[578]&m[843]&~m[845]&~m[846]&m[847])|(~m[578]&~m[843]&m[845]&~m[846]&m[847])|(m[578]&m[843]&m[845]&~m[846]&m[847])|(~m[578]&m[843]&m[845]&m[846]&m[847]))&UnbiasedRNG[408])|((m[578]&~m[843]&~m[845]&m[846]&~m[847])|(~m[578]&~m[843]&~m[845]&~m[846]&m[847])|(m[578]&~m[843]&~m[845]&~m[846]&m[847])|(m[578]&m[843]&~m[845]&~m[846]&m[847])|(m[578]&~m[843]&m[845]&~m[846]&m[847])|(~m[578]&~m[843]&~m[845]&m[846]&m[847])|(m[578]&~m[843]&~m[845]&m[846]&m[847])|(~m[578]&m[843]&~m[845]&m[846]&m[847])|(m[578]&m[843]&~m[845]&m[846]&m[847])|(~m[578]&~m[843]&m[845]&m[846]&m[847])|(m[578]&~m[843]&m[845]&m[846]&m[847])|(m[578]&m[843]&m[845]&m[846]&m[847]))):InitCond[1107];
    m[849] = run?((((m[591]&~m[848]&~m[850]&~m[851]&~m[852])|(~m[591]&~m[848]&~m[850]&m[851]&~m[852])|(m[591]&m[848]&~m[850]&m[851]&~m[852])|(m[591]&~m[848]&m[850]&m[851]&~m[852])|(~m[591]&m[848]&~m[850]&~m[851]&m[852])|(~m[591]&~m[848]&m[850]&~m[851]&m[852])|(m[591]&m[848]&m[850]&~m[851]&m[852])|(~m[591]&m[848]&m[850]&m[851]&m[852]))&UnbiasedRNG[409])|((m[591]&~m[848]&~m[850]&m[851]&~m[852])|(~m[591]&~m[848]&~m[850]&~m[851]&m[852])|(m[591]&~m[848]&~m[850]&~m[851]&m[852])|(m[591]&m[848]&~m[850]&~m[851]&m[852])|(m[591]&~m[848]&m[850]&~m[851]&m[852])|(~m[591]&~m[848]&~m[850]&m[851]&m[852])|(m[591]&~m[848]&~m[850]&m[851]&m[852])|(~m[591]&m[848]&~m[850]&m[851]&m[852])|(m[591]&m[848]&~m[850]&m[851]&m[852])|(~m[591]&~m[848]&m[850]&m[851]&m[852])|(m[591]&~m[848]&m[850]&m[851]&m[852])|(m[591]&m[848]&m[850]&m[851]&m[852]))):InitCond[1108];
    m[854] = run?((((m[604]&~m[853]&~m[855]&~m[856]&~m[857])|(~m[604]&~m[853]&~m[855]&m[856]&~m[857])|(m[604]&m[853]&~m[855]&m[856]&~m[857])|(m[604]&~m[853]&m[855]&m[856]&~m[857])|(~m[604]&m[853]&~m[855]&~m[856]&m[857])|(~m[604]&~m[853]&m[855]&~m[856]&m[857])|(m[604]&m[853]&m[855]&~m[856]&m[857])|(~m[604]&m[853]&m[855]&m[856]&m[857]))&UnbiasedRNG[410])|((m[604]&~m[853]&~m[855]&m[856]&~m[857])|(~m[604]&~m[853]&~m[855]&~m[856]&m[857])|(m[604]&~m[853]&~m[855]&~m[856]&m[857])|(m[604]&m[853]&~m[855]&~m[856]&m[857])|(m[604]&~m[853]&m[855]&~m[856]&m[857])|(~m[604]&~m[853]&~m[855]&m[856]&m[857])|(m[604]&~m[853]&~m[855]&m[856]&m[857])|(~m[604]&m[853]&~m[855]&m[856]&m[857])|(m[604]&m[853]&~m[855]&m[856]&m[857])|(~m[604]&~m[853]&m[855]&m[856]&m[857])|(m[604]&~m[853]&m[855]&m[856]&m[857])|(m[604]&m[853]&m[855]&m[856]&m[857]))):InitCond[1109];
    m[860] = run?((((m[832]&~m[858]&~m[859]&~m[861]&~m[862])|(~m[832]&~m[858]&~m[859]&m[861]&~m[862])|(m[832]&m[858]&~m[859]&m[861]&~m[862])|(m[832]&~m[858]&m[859]&m[861]&~m[862])|(~m[832]&m[858]&~m[859]&~m[861]&m[862])|(~m[832]&~m[858]&m[859]&~m[861]&m[862])|(m[832]&m[858]&m[859]&~m[861]&m[862])|(~m[832]&m[858]&m[859]&m[861]&m[862]))&UnbiasedRNG[411])|((m[832]&~m[858]&~m[859]&m[861]&~m[862])|(~m[832]&~m[858]&~m[859]&~m[861]&m[862])|(m[832]&~m[858]&~m[859]&~m[861]&m[862])|(m[832]&m[858]&~m[859]&~m[861]&m[862])|(m[832]&~m[858]&m[859]&~m[861]&m[862])|(~m[832]&~m[858]&~m[859]&m[861]&m[862])|(m[832]&~m[858]&~m[859]&m[861]&m[862])|(~m[832]&m[858]&~m[859]&m[861]&m[862])|(m[832]&m[858]&~m[859]&m[861]&m[862])|(~m[832]&~m[858]&m[859]&m[861]&m[862])|(m[832]&~m[858]&m[859]&m[861]&m[862])|(m[832]&m[858]&m[859]&m[861]&m[862]))):InitCond[1110];
    m[870] = run?((((m[837]&~m[868]&~m[869]&~m[871]&~m[872])|(~m[837]&~m[868]&~m[869]&m[871]&~m[872])|(m[837]&m[868]&~m[869]&m[871]&~m[872])|(m[837]&~m[868]&m[869]&m[871]&~m[872])|(~m[837]&m[868]&~m[869]&~m[871]&m[872])|(~m[837]&~m[868]&m[869]&~m[871]&m[872])|(m[837]&m[868]&m[869]&~m[871]&m[872])|(~m[837]&m[868]&m[869]&m[871]&m[872]))&UnbiasedRNG[412])|((m[837]&~m[868]&~m[869]&m[871]&~m[872])|(~m[837]&~m[868]&~m[869]&~m[871]&m[872])|(m[837]&~m[868]&~m[869]&~m[871]&m[872])|(m[837]&m[868]&~m[869]&~m[871]&m[872])|(m[837]&~m[868]&m[869]&~m[871]&m[872])|(~m[837]&~m[868]&~m[869]&m[871]&m[872])|(m[837]&~m[868]&~m[869]&m[871]&m[872])|(~m[837]&m[868]&~m[869]&m[871]&m[872])|(m[837]&m[868]&~m[869]&m[871]&m[872])|(~m[837]&~m[868]&m[869]&m[871]&m[872])|(m[837]&~m[868]&m[869]&m[871]&m[872])|(m[837]&m[868]&m[869]&m[871]&m[872]))):InitCond[1111];
    m[875] = run?((((m[842]&~m[873]&~m[874]&~m[876]&~m[877])|(~m[842]&~m[873]&~m[874]&m[876]&~m[877])|(m[842]&m[873]&~m[874]&m[876]&~m[877])|(m[842]&~m[873]&m[874]&m[876]&~m[877])|(~m[842]&m[873]&~m[874]&~m[876]&m[877])|(~m[842]&~m[873]&m[874]&~m[876]&m[877])|(m[842]&m[873]&m[874]&~m[876]&m[877])|(~m[842]&m[873]&m[874]&m[876]&m[877]))&UnbiasedRNG[413])|((m[842]&~m[873]&~m[874]&m[876]&~m[877])|(~m[842]&~m[873]&~m[874]&~m[876]&m[877])|(m[842]&~m[873]&~m[874]&~m[876]&m[877])|(m[842]&m[873]&~m[874]&~m[876]&m[877])|(m[842]&~m[873]&m[874]&~m[876]&m[877])|(~m[842]&~m[873]&~m[874]&m[876]&m[877])|(m[842]&~m[873]&~m[874]&m[876]&m[877])|(~m[842]&m[873]&~m[874]&m[876]&m[877])|(m[842]&m[873]&~m[874]&m[876]&m[877])|(~m[842]&~m[873]&m[874]&m[876]&m[877])|(m[842]&~m[873]&m[874]&m[876]&m[877])|(m[842]&m[873]&m[874]&m[876]&m[877]))):InitCond[1112];
    m[879] = run?((((m[579]&~m[878]&~m[880]&~m[881]&~m[882])|(~m[579]&~m[878]&~m[880]&m[881]&~m[882])|(m[579]&m[878]&~m[880]&m[881]&~m[882])|(m[579]&~m[878]&m[880]&m[881]&~m[882])|(~m[579]&m[878]&~m[880]&~m[881]&m[882])|(~m[579]&~m[878]&m[880]&~m[881]&m[882])|(m[579]&m[878]&m[880]&~m[881]&m[882])|(~m[579]&m[878]&m[880]&m[881]&m[882]))&UnbiasedRNG[414])|((m[579]&~m[878]&~m[880]&m[881]&~m[882])|(~m[579]&~m[878]&~m[880]&~m[881]&m[882])|(m[579]&~m[878]&~m[880]&~m[881]&m[882])|(m[579]&m[878]&~m[880]&~m[881]&m[882])|(m[579]&~m[878]&m[880]&~m[881]&m[882])|(~m[579]&~m[878]&~m[880]&m[881]&m[882])|(m[579]&~m[878]&~m[880]&m[881]&m[882])|(~m[579]&m[878]&~m[880]&m[881]&m[882])|(m[579]&m[878]&~m[880]&m[881]&m[882])|(~m[579]&~m[878]&m[880]&m[881]&m[882])|(m[579]&~m[878]&m[880]&m[881]&m[882])|(m[579]&m[878]&m[880]&m[881]&m[882]))):InitCond[1113];
    m[884] = run?((((m[592]&~m[883]&~m[885]&~m[886]&~m[887])|(~m[592]&~m[883]&~m[885]&m[886]&~m[887])|(m[592]&m[883]&~m[885]&m[886]&~m[887])|(m[592]&~m[883]&m[885]&m[886]&~m[887])|(~m[592]&m[883]&~m[885]&~m[886]&m[887])|(~m[592]&~m[883]&m[885]&~m[886]&m[887])|(m[592]&m[883]&m[885]&~m[886]&m[887])|(~m[592]&m[883]&m[885]&m[886]&m[887]))&UnbiasedRNG[415])|((m[592]&~m[883]&~m[885]&m[886]&~m[887])|(~m[592]&~m[883]&~m[885]&~m[886]&m[887])|(m[592]&~m[883]&~m[885]&~m[886]&m[887])|(m[592]&m[883]&~m[885]&~m[886]&m[887])|(m[592]&~m[883]&m[885]&~m[886]&m[887])|(~m[592]&~m[883]&~m[885]&m[886]&m[887])|(m[592]&~m[883]&~m[885]&m[886]&m[887])|(~m[592]&m[883]&~m[885]&m[886]&m[887])|(m[592]&m[883]&~m[885]&m[886]&m[887])|(~m[592]&~m[883]&m[885]&m[886]&m[887])|(m[592]&~m[883]&m[885]&m[886]&m[887])|(m[592]&m[883]&m[885]&m[886]&m[887]))):InitCond[1114];
    m[889] = run?((((m[605]&~m[888]&~m[890]&~m[891]&~m[892])|(~m[605]&~m[888]&~m[890]&m[891]&~m[892])|(m[605]&m[888]&~m[890]&m[891]&~m[892])|(m[605]&~m[888]&m[890]&m[891]&~m[892])|(~m[605]&m[888]&~m[890]&~m[891]&m[892])|(~m[605]&~m[888]&m[890]&~m[891]&m[892])|(m[605]&m[888]&m[890]&~m[891]&m[892])|(~m[605]&m[888]&m[890]&m[891]&m[892]))&UnbiasedRNG[416])|((m[605]&~m[888]&~m[890]&m[891]&~m[892])|(~m[605]&~m[888]&~m[890]&~m[891]&m[892])|(m[605]&~m[888]&~m[890]&~m[891]&m[892])|(m[605]&m[888]&~m[890]&~m[891]&m[892])|(m[605]&~m[888]&m[890]&~m[891]&m[892])|(~m[605]&~m[888]&~m[890]&m[891]&m[892])|(m[605]&~m[888]&~m[890]&m[891]&m[892])|(~m[605]&m[888]&~m[890]&m[891]&m[892])|(m[605]&m[888]&~m[890]&m[891]&m[892])|(~m[605]&~m[888]&m[890]&m[891]&m[892])|(m[605]&~m[888]&m[890]&m[891]&m[892])|(m[605]&m[888]&m[890]&m[891]&m[892]))):InitCond[1115];
    m[895] = run?((((m[862]&~m[893]&~m[894]&~m[896]&~m[897])|(~m[862]&~m[893]&~m[894]&m[896]&~m[897])|(m[862]&m[893]&~m[894]&m[896]&~m[897])|(m[862]&~m[893]&m[894]&m[896]&~m[897])|(~m[862]&m[893]&~m[894]&~m[896]&m[897])|(~m[862]&~m[893]&m[894]&~m[896]&m[897])|(m[862]&m[893]&m[894]&~m[896]&m[897])|(~m[862]&m[893]&m[894]&m[896]&m[897]))&UnbiasedRNG[417])|((m[862]&~m[893]&~m[894]&m[896]&~m[897])|(~m[862]&~m[893]&~m[894]&~m[896]&m[897])|(m[862]&~m[893]&~m[894]&~m[896]&m[897])|(m[862]&m[893]&~m[894]&~m[896]&m[897])|(m[862]&~m[893]&m[894]&~m[896]&m[897])|(~m[862]&~m[893]&~m[894]&m[896]&m[897])|(m[862]&~m[893]&~m[894]&m[896]&m[897])|(~m[862]&m[893]&~m[894]&m[896]&m[897])|(m[862]&m[893]&~m[894]&m[896]&m[897])|(~m[862]&~m[893]&m[894]&m[896]&m[897])|(m[862]&~m[893]&m[894]&m[896]&m[897])|(m[862]&m[893]&m[894]&m[896]&m[897]))):InitCond[1116];
    m[900] = run?((((m[867]&~m[898]&~m[899]&~m[901]&~m[902])|(~m[867]&~m[898]&~m[899]&m[901]&~m[902])|(m[867]&m[898]&~m[899]&m[901]&~m[902])|(m[867]&~m[898]&m[899]&m[901]&~m[902])|(~m[867]&m[898]&~m[899]&~m[901]&m[902])|(~m[867]&~m[898]&m[899]&~m[901]&m[902])|(m[867]&m[898]&m[899]&~m[901]&m[902])|(~m[867]&m[898]&m[899]&m[901]&m[902]))&UnbiasedRNG[418])|((m[867]&~m[898]&~m[899]&m[901]&~m[902])|(~m[867]&~m[898]&~m[899]&~m[901]&m[902])|(m[867]&~m[898]&~m[899]&~m[901]&m[902])|(m[867]&m[898]&~m[899]&~m[901]&m[902])|(m[867]&~m[898]&m[899]&~m[901]&m[902])|(~m[867]&~m[898]&~m[899]&m[901]&m[902])|(m[867]&~m[898]&~m[899]&m[901]&m[902])|(~m[867]&m[898]&~m[899]&m[901]&m[902])|(m[867]&m[898]&~m[899]&m[901]&m[902])|(~m[867]&~m[898]&m[899]&m[901]&m[902])|(m[867]&~m[898]&m[899]&m[901]&m[902])|(m[867]&m[898]&m[899]&m[901]&m[902]))):InitCond[1117];
    m[910] = run?((((m[872]&~m[908]&~m[909]&~m[911]&~m[912])|(~m[872]&~m[908]&~m[909]&m[911]&~m[912])|(m[872]&m[908]&~m[909]&m[911]&~m[912])|(m[872]&~m[908]&m[909]&m[911]&~m[912])|(~m[872]&m[908]&~m[909]&~m[911]&m[912])|(~m[872]&~m[908]&m[909]&~m[911]&m[912])|(m[872]&m[908]&m[909]&~m[911]&m[912])|(~m[872]&m[908]&m[909]&m[911]&m[912]))&UnbiasedRNG[419])|((m[872]&~m[908]&~m[909]&m[911]&~m[912])|(~m[872]&~m[908]&~m[909]&~m[911]&m[912])|(m[872]&~m[908]&~m[909]&~m[911]&m[912])|(m[872]&m[908]&~m[909]&~m[911]&m[912])|(m[872]&~m[908]&m[909]&~m[911]&m[912])|(~m[872]&~m[908]&~m[909]&m[911]&m[912])|(m[872]&~m[908]&~m[909]&m[911]&m[912])|(~m[872]&m[908]&~m[909]&m[911]&m[912])|(m[872]&m[908]&~m[909]&m[911]&m[912])|(~m[872]&~m[908]&m[909]&m[911]&m[912])|(m[872]&~m[908]&m[909]&m[911]&m[912])|(m[872]&m[908]&m[909]&m[911]&m[912]))):InitCond[1118];
    m[915] = run?((((m[877]&~m[913]&~m[914]&~m[916]&~m[917])|(~m[877]&~m[913]&~m[914]&m[916]&~m[917])|(m[877]&m[913]&~m[914]&m[916]&~m[917])|(m[877]&~m[913]&m[914]&m[916]&~m[917])|(~m[877]&m[913]&~m[914]&~m[916]&m[917])|(~m[877]&~m[913]&m[914]&~m[916]&m[917])|(m[877]&m[913]&m[914]&~m[916]&m[917])|(~m[877]&m[913]&m[914]&m[916]&m[917]))&UnbiasedRNG[420])|((m[877]&~m[913]&~m[914]&m[916]&~m[917])|(~m[877]&~m[913]&~m[914]&~m[916]&m[917])|(m[877]&~m[913]&~m[914]&~m[916]&m[917])|(m[877]&m[913]&~m[914]&~m[916]&m[917])|(m[877]&~m[913]&m[914]&~m[916]&m[917])|(~m[877]&~m[913]&~m[914]&m[916]&m[917])|(m[877]&~m[913]&~m[914]&m[916]&m[917])|(~m[877]&m[913]&~m[914]&m[916]&m[917])|(m[877]&m[913]&~m[914]&m[916]&m[917])|(~m[877]&~m[913]&m[914]&m[916]&m[917])|(m[877]&~m[913]&m[914]&m[916]&m[917])|(m[877]&m[913]&m[914]&m[916]&m[917]))):InitCond[1119];
    m[920] = run?((((m[882]&~m[918]&~m[919]&~m[921]&~m[922])|(~m[882]&~m[918]&~m[919]&m[921]&~m[922])|(m[882]&m[918]&~m[919]&m[921]&~m[922])|(m[882]&~m[918]&m[919]&m[921]&~m[922])|(~m[882]&m[918]&~m[919]&~m[921]&m[922])|(~m[882]&~m[918]&m[919]&~m[921]&m[922])|(m[882]&m[918]&m[919]&~m[921]&m[922])|(~m[882]&m[918]&m[919]&m[921]&m[922]))&UnbiasedRNG[421])|((m[882]&~m[918]&~m[919]&m[921]&~m[922])|(~m[882]&~m[918]&~m[919]&~m[921]&m[922])|(m[882]&~m[918]&~m[919]&~m[921]&m[922])|(m[882]&m[918]&~m[919]&~m[921]&m[922])|(m[882]&~m[918]&m[919]&~m[921]&m[922])|(~m[882]&~m[918]&~m[919]&m[921]&m[922])|(m[882]&~m[918]&~m[919]&m[921]&m[922])|(~m[882]&m[918]&~m[919]&m[921]&m[922])|(m[882]&m[918]&~m[919]&m[921]&m[922])|(~m[882]&~m[918]&m[919]&m[921]&m[922])|(m[882]&~m[918]&m[919]&m[921]&m[922])|(m[882]&m[918]&m[919]&m[921]&m[922]))):InitCond[1120];
    m[924] = run?((((m[593]&~m[923]&~m[925]&~m[926]&~m[927])|(~m[593]&~m[923]&~m[925]&m[926]&~m[927])|(m[593]&m[923]&~m[925]&m[926]&~m[927])|(m[593]&~m[923]&m[925]&m[926]&~m[927])|(~m[593]&m[923]&~m[925]&~m[926]&m[927])|(~m[593]&~m[923]&m[925]&~m[926]&m[927])|(m[593]&m[923]&m[925]&~m[926]&m[927])|(~m[593]&m[923]&m[925]&m[926]&m[927]))&UnbiasedRNG[422])|((m[593]&~m[923]&~m[925]&m[926]&~m[927])|(~m[593]&~m[923]&~m[925]&~m[926]&m[927])|(m[593]&~m[923]&~m[925]&~m[926]&m[927])|(m[593]&m[923]&~m[925]&~m[926]&m[927])|(m[593]&~m[923]&m[925]&~m[926]&m[927])|(~m[593]&~m[923]&~m[925]&m[926]&m[927])|(m[593]&~m[923]&~m[925]&m[926]&m[927])|(~m[593]&m[923]&~m[925]&m[926]&m[927])|(m[593]&m[923]&~m[925]&m[926]&m[927])|(~m[593]&~m[923]&m[925]&m[926]&m[927])|(m[593]&~m[923]&m[925]&m[926]&m[927])|(m[593]&m[923]&m[925]&m[926]&m[927]))):InitCond[1121];
    m[929] = run?((((m[606]&~m[928]&~m[930]&~m[931]&~m[932])|(~m[606]&~m[928]&~m[930]&m[931]&~m[932])|(m[606]&m[928]&~m[930]&m[931]&~m[932])|(m[606]&~m[928]&m[930]&m[931]&~m[932])|(~m[606]&m[928]&~m[930]&~m[931]&m[932])|(~m[606]&~m[928]&m[930]&~m[931]&m[932])|(m[606]&m[928]&m[930]&~m[931]&m[932])|(~m[606]&m[928]&m[930]&m[931]&m[932]))&UnbiasedRNG[423])|((m[606]&~m[928]&~m[930]&m[931]&~m[932])|(~m[606]&~m[928]&~m[930]&~m[931]&m[932])|(m[606]&~m[928]&~m[930]&~m[931]&m[932])|(m[606]&m[928]&~m[930]&~m[931]&m[932])|(m[606]&~m[928]&m[930]&~m[931]&m[932])|(~m[606]&~m[928]&~m[930]&m[931]&m[932])|(m[606]&~m[928]&~m[930]&m[931]&m[932])|(~m[606]&m[928]&~m[930]&m[931]&m[932])|(m[606]&m[928]&~m[930]&m[931]&m[932])|(~m[606]&~m[928]&m[930]&m[931]&m[932])|(m[606]&~m[928]&m[930]&m[931]&m[932])|(m[606]&m[928]&m[930]&m[931]&m[932]))):InitCond[1122];
    m[935] = run?((((m[897]&~m[933]&~m[934]&~m[936]&~m[937])|(~m[897]&~m[933]&~m[934]&m[936]&~m[937])|(m[897]&m[933]&~m[934]&m[936]&~m[937])|(m[897]&~m[933]&m[934]&m[936]&~m[937])|(~m[897]&m[933]&~m[934]&~m[936]&m[937])|(~m[897]&~m[933]&m[934]&~m[936]&m[937])|(m[897]&m[933]&m[934]&~m[936]&m[937])|(~m[897]&m[933]&m[934]&m[936]&m[937]))&UnbiasedRNG[424])|((m[897]&~m[933]&~m[934]&m[936]&~m[937])|(~m[897]&~m[933]&~m[934]&~m[936]&m[937])|(m[897]&~m[933]&~m[934]&~m[936]&m[937])|(m[897]&m[933]&~m[934]&~m[936]&m[937])|(m[897]&~m[933]&m[934]&~m[936]&m[937])|(~m[897]&~m[933]&~m[934]&m[936]&m[937])|(m[897]&~m[933]&~m[934]&m[936]&m[937])|(~m[897]&m[933]&~m[934]&m[936]&m[937])|(m[897]&m[933]&~m[934]&m[936]&m[937])|(~m[897]&~m[933]&m[934]&m[936]&m[937])|(m[897]&~m[933]&m[934]&m[936]&m[937])|(m[897]&m[933]&m[934]&m[936]&m[937]))):InitCond[1123];
    m[940] = run?((((m[902]&~m[938]&~m[939]&~m[941]&~m[942])|(~m[902]&~m[938]&~m[939]&m[941]&~m[942])|(m[902]&m[938]&~m[939]&m[941]&~m[942])|(m[902]&~m[938]&m[939]&m[941]&~m[942])|(~m[902]&m[938]&~m[939]&~m[941]&m[942])|(~m[902]&~m[938]&m[939]&~m[941]&m[942])|(m[902]&m[938]&m[939]&~m[941]&m[942])|(~m[902]&m[938]&m[939]&m[941]&m[942]))&UnbiasedRNG[425])|((m[902]&~m[938]&~m[939]&m[941]&~m[942])|(~m[902]&~m[938]&~m[939]&~m[941]&m[942])|(m[902]&~m[938]&~m[939]&~m[941]&m[942])|(m[902]&m[938]&~m[939]&~m[941]&m[942])|(m[902]&~m[938]&m[939]&~m[941]&m[942])|(~m[902]&~m[938]&~m[939]&m[941]&m[942])|(m[902]&~m[938]&~m[939]&m[941]&m[942])|(~m[902]&m[938]&~m[939]&m[941]&m[942])|(m[902]&m[938]&~m[939]&m[941]&m[942])|(~m[902]&~m[938]&m[939]&m[941]&m[942])|(m[902]&~m[938]&m[939]&m[941]&m[942])|(m[902]&m[938]&m[939]&m[941]&m[942]))):InitCond[1124];
    m[945] = run?((((m[907]&~m[943]&~m[944]&~m[946]&~m[947])|(~m[907]&~m[943]&~m[944]&m[946]&~m[947])|(m[907]&m[943]&~m[944]&m[946]&~m[947])|(m[907]&~m[943]&m[944]&m[946]&~m[947])|(~m[907]&m[943]&~m[944]&~m[946]&m[947])|(~m[907]&~m[943]&m[944]&~m[946]&m[947])|(m[907]&m[943]&m[944]&~m[946]&m[947])|(~m[907]&m[943]&m[944]&m[946]&m[947]))&UnbiasedRNG[426])|((m[907]&~m[943]&~m[944]&m[946]&~m[947])|(~m[907]&~m[943]&~m[944]&~m[946]&m[947])|(m[907]&~m[943]&~m[944]&~m[946]&m[947])|(m[907]&m[943]&~m[944]&~m[946]&m[947])|(m[907]&~m[943]&m[944]&~m[946]&m[947])|(~m[907]&~m[943]&~m[944]&m[946]&m[947])|(m[907]&~m[943]&~m[944]&m[946]&m[947])|(~m[907]&m[943]&~m[944]&m[946]&m[947])|(m[907]&m[943]&~m[944]&m[946]&m[947])|(~m[907]&~m[943]&m[944]&m[946]&m[947])|(m[907]&~m[943]&m[944]&m[946]&m[947])|(m[907]&m[943]&m[944]&m[946]&m[947]))):InitCond[1125];
    m[955] = run?((((m[912]&~m[953]&~m[954]&~m[956]&~m[957])|(~m[912]&~m[953]&~m[954]&m[956]&~m[957])|(m[912]&m[953]&~m[954]&m[956]&~m[957])|(m[912]&~m[953]&m[954]&m[956]&~m[957])|(~m[912]&m[953]&~m[954]&~m[956]&m[957])|(~m[912]&~m[953]&m[954]&~m[956]&m[957])|(m[912]&m[953]&m[954]&~m[956]&m[957])|(~m[912]&m[953]&m[954]&m[956]&m[957]))&UnbiasedRNG[427])|((m[912]&~m[953]&~m[954]&m[956]&~m[957])|(~m[912]&~m[953]&~m[954]&~m[956]&m[957])|(m[912]&~m[953]&~m[954]&~m[956]&m[957])|(m[912]&m[953]&~m[954]&~m[956]&m[957])|(m[912]&~m[953]&m[954]&~m[956]&m[957])|(~m[912]&~m[953]&~m[954]&m[956]&m[957])|(m[912]&~m[953]&~m[954]&m[956]&m[957])|(~m[912]&m[953]&~m[954]&m[956]&m[957])|(m[912]&m[953]&~m[954]&m[956]&m[957])|(~m[912]&~m[953]&m[954]&m[956]&m[957])|(m[912]&~m[953]&m[954]&m[956]&m[957])|(m[912]&m[953]&m[954]&m[956]&m[957]))):InitCond[1126];
    m[960] = run?((((m[917]&~m[958]&~m[959]&~m[961]&~m[962])|(~m[917]&~m[958]&~m[959]&m[961]&~m[962])|(m[917]&m[958]&~m[959]&m[961]&~m[962])|(m[917]&~m[958]&m[959]&m[961]&~m[962])|(~m[917]&m[958]&~m[959]&~m[961]&m[962])|(~m[917]&~m[958]&m[959]&~m[961]&m[962])|(m[917]&m[958]&m[959]&~m[961]&m[962])|(~m[917]&m[958]&m[959]&m[961]&m[962]))&UnbiasedRNG[428])|((m[917]&~m[958]&~m[959]&m[961]&~m[962])|(~m[917]&~m[958]&~m[959]&~m[961]&m[962])|(m[917]&~m[958]&~m[959]&~m[961]&m[962])|(m[917]&m[958]&~m[959]&~m[961]&m[962])|(m[917]&~m[958]&m[959]&~m[961]&m[962])|(~m[917]&~m[958]&~m[959]&m[961]&m[962])|(m[917]&~m[958]&~m[959]&m[961]&m[962])|(~m[917]&m[958]&~m[959]&m[961]&m[962])|(m[917]&m[958]&~m[959]&m[961]&m[962])|(~m[917]&~m[958]&m[959]&m[961]&m[962])|(m[917]&~m[958]&m[959]&m[961]&m[962])|(m[917]&m[958]&m[959]&m[961]&m[962]))):InitCond[1127];
    m[965] = run?((((m[922]&~m[963]&~m[964]&~m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&m[966]&~m[967])|(m[922]&m[963]&~m[964]&m[966]&~m[967])|(m[922]&~m[963]&m[964]&m[966]&~m[967])|(~m[922]&m[963]&~m[964]&~m[966]&m[967])|(~m[922]&~m[963]&m[964]&~m[966]&m[967])|(m[922]&m[963]&m[964]&~m[966]&m[967])|(~m[922]&m[963]&m[964]&m[966]&m[967]))&UnbiasedRNG[429])|((m[922]&~m[963]&~m[964]&m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&m[964]&~m[966]&m[967])|(~m[922]&~m[963]&~m[964]&m[966]&m[967])|(m[922]&~m[963]&~m[964]&m[966]&m[967])|(~m[922]&m[963]&~m[964]&m[966]&m[967])|(m[922]&m[963]&~m[964]&m[966]&m[967])|(~m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&m[963]&m[964]&m[966]&m[967]))):InitCond[1128];
    m[970] = run?((((m[927]&~m[968]&~m[969]&~m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&m[971]&~m[972])|(m[927]&m[968]&~m[969]&m[971]&~m[972])|(m[927]&~m[968]&m[969]&m[971]&~m[972])|(~m[927]&m[968]&~m[969]&~m[971]&m[972])|(~m[927]&~m[968]&m[969]&~m[971]&m[972])|(m[927]&m[968]&m[969]&~m[971]&m[972])|(~m[927]&m[968]&m[969]&m[971]&m[972]))&UnbiasedRNG[430])|((m[927]&~m[968]&~m[969]&m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&m[969]&~m[971]&m[972])|(~m[927]&~m[968]&~m[969]&m[971]&m[972])|(m[927]&~m[968]&~m[969]&m[971]&m[972])|(~m[927]&m[968]&~m[969]&m[971]&m[972])|(m[927]&m[968]&~m[969]&m[971]&m[972])|(~m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&m[968]&m[969]&m[971]&m[972]))):InitCond[1129];
    m[974] = run?((((m[607]&~m[973]&~m[975]&~m[976]&~m[977])|(~m[607]&~m[973]&~m[975]&m[976]&~m[977])|(m[607]&m[973]&~m[975]&m[976]&~m[977])|(m[607]&~m[973]&m[975]&m[976]&~m[977])|(~m[607]&m[973]&~m[975]&~m[976]&m[977])|(~m[607]&~m[973]&m[975]&~m[976]&m[977])|(m[607]&m[973]&m[975]&~m[976]&m[977])|(~m[607]&m[973]&m[975]&m[976]&m[977]))&UnbiasedRNG[431])|((m[607]&~m[973]&~m[975]&m[976]&~m[977])|(~m[607]&~m[973]&~m[975]&~m[976]&m[977])|(m[607]&~m[973]&~m[975]&~m[976]&m[977])|(m[607]&m[973]&~m[975]&~m[976]&m[977])|(m[607]&~m[973]&m[975]&~m[976]&m[977])|(~m[607]&~m[973]&~m[975]&m[976]&m[977])|(m[607]&~m[973]&~m[975]&m[976]&m[977])|(~m[607]&m[973]&~m[975]&m[976]&m[977])|(m[607]&m[973]&~m[975]&m[976]&m[977])|(~m[607]&~m[973]&m[975]&m[976]&m[977])|(m[607]&~m[973]&m[975]&m[976]&m[977])|(m[607]&m[973]&m[975]&m[976]&m[977]))):InitCond[1130];
    m[980] = run?((((m[937]&~m[978]&~m[979]&~m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&m[981]&~m[982])|(m[937]&m[978]&~m[979]&m[981]&~m[982])|(m[937]&~m[978]&m[979]&m[981]&~m[982])|(~m[937]&m[978]&~m[979]&~m[981]&m[982])|(~m[937]&~m[978]&m[979]&~m[981]&m[982])|(m[937]&m[978]&m[979]&~m[981]&m[982])|(~m[937]&m[978]&m[979]&m[981]&m[982]))&UnbiasedRNG[432])|((m[937]&~m[978]&~m[979]&m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&m[979]&~m[981]&m[982])|(~m[937]&~m[978]&~m[979]&m[981]&m[982])|(m[937]&~m[978]&~m[979]&m[981]&m[982])|(~m[937]&m[978]&~m[979]&m[981]&m[982])|(m[937]&m[978]&~m[979]&m[981]&m[982])|(~m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&m[978]&m[979]&m[981]&m[982]))):InitCond[1131];
    m[985] = run?((((m[942]&~m[983]&~m[984]&~m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&m[986]&~m[987])|(m[942]&m[983]&~m[984]&m[986]&~m[987])|(m[942]&~m[983]&m[984]&m[986]&~m[987])|(~m[942]&m[983]&~m[984]&~m[986]&m[987])|(~m[942]&~m[983]&m[984]&~m[986]&m[987])|(m[942]&m[983]&m[984]&~m[986]&m[987])|(~m[942]&m[983]&m[984]&m[986]&m[987]))&UnbiasedRNG[433])|((m[942]&~m[983]&~m[984]&m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&m[984]&~m[986]&m[987])|(~m[942]&~m[983]&~m[984]&m[986]&m[987])|(m[942]&~m[983]&~m[984]&m[986]&m[987])|(~m[942]&m[983]&~m[984]&m[986]&m[987])|(m[942]&m[983]&~m[984]&m[986]&m[987])|(~m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&m[983]&m[984]&m[986]&m[987]))):InitCond[1132];
    m[990] = run?((((m[947]&~m[988]&~m[989]&~m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&m[991]&~m[992])|(m[947]&m[988]&~m[989]&m[991]&~m[992])|(m[947]&~m[988]&m[989]&m[991]&~m[992])|(~m[947]&m[988]&~m[989]&~m[991]&m[992])|(~m[947]&~m[988]&m[989]&~m[991]&m[992])|(m[947]&m[988]&m[989]&~m[991]&m[992])|(~m[947]&m[988]&m[989]&m[991]&m[992]))&UnbiasedRNG[434])|((m[947]&~m[988]&~m[989]&m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&m[989]&~m[991]&m[992])|(~m[947]&~m[988]&~m[989]&m[991]&m[992])|(m[947]&~m[988]&~m[989]&m[991]&m[992])|(~m[947]&m[988]&~m[989]&m[991]&m[992])|(m[947]&m[988]&~m[989]&m[991]&m[992])|(~m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&m[988]&m[989]&m[991]&m[992]))):InitCond[1133];
    m[995] = run?((((m[952]&~m[993]&~m[994]&~m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&m[996]&~m[997])|(m[952]&m[993]&~m[994]&m[996]&~m[997])|(m[952]&~m[993]&m[994]&m[996]&~m[997])|(~m[952]&m[993]&~m[994]&~m[996]&m[997])|(~m[952]&~m[993]&m[994]&~m[996]&m[997])|(m[952]&m[993]&m[994]&~m[996]&m[997])|(~m[952]&m[993]&m[994]&m[996]&m[997]))&UnbiasedRNG[435])|((m[952]&~m[993]&~m[994]&m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&m[994]&~m[996]&m[997])|(~m[952]&~m[993]&~m[994]&m[996]&m[997])|(m[952]&~m[993]&~m[994]&m[996]&m[997])|(~m[952]&m[993]&~m[994]&m[996]&m[997])|(m[952]&m[993]&~m[994]&m[996]&m[997])|(~m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&m[993]&m[994]&m[996]&m[997]))):InitCond[1134];
    m[1005] = run?((((m[957]&~m[1003]&~m[1004]&~m[1006]&~m[1007])|(~m[957]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(m[957]&m[1003]&~m[1004]&m[1006]&~m[1007])|(m[957]&~m[1003]&m[1004]&m[1006]&~m[1007])|(~m[957]&m[1003]&~m[1004]&~m[1006]&m[1007])|(~m[957]&~m[1003]&m[1004]&~m[1006]&m[1007])|(m[957]&m[1003]&m[1004]&~m[1006]&m[1007])|(~m[957]&m[1003]&m[1004]&m[1006]&m[1007]))&UnbiasedRNG[436])|((m[957]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(~m[957]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[957]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[957]&m[1003]&~m[1004]&~m[1006]&m[1007])|(m[957]&~m[1003]&m[1004]&~m[1006]&m[1007])|(~m[957]&~m[1003]&~m[1004]&m[1006]&m[1007])|(m[957]&~m[1003]&~m[1004]&m[1006]&m[1007])|(~m[957]&m[1003]&~m[1004]&m[1006]&m[1007])|(m[957]&m[1003]&~m[1004]&m[1006]&m[1007])|(~m[957]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[957]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[957]&m[1003]&m[1004]&m[1006]&m[1007]))):InitCond[1135];
    m[1010] = run?((((m[962]&~m[1008]&~m[1009]&~m[1011]&~m[1012])|(~m[962]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(m[962]&m[1008]&~m[1009]&m[1011]&~m[1012])|(m[962]&~m[1008]&m[1009]&m[1011]&~m[1012])|(~m[962]&m[1008]&~m[1009]&~m[1011]&m[1012])|(~m[962]&~m[1008]&m[1009]&~m[1011]&m[1012])|(m[962]&m[1008]&m[1009]&~m[1011]&m[1012])|(~m[962]&m[1008]&m[1009]&m[1011]&m[1012]))&UnbiasedRNG[437])|((m[962]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(~m[962]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[962]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[962]&m[1008]&~m[1009]&~m[1011]&m[1012])|(m[962]&~m[1008]&m[1009]&~m[1011]&m[1012])|(~m[962]&~m[1008]&~m[1009]&m[1011]&m[1012])|(m[962]&~m[1008]&~m[1009]&m[1011]&m[1012])|(~m[962]&m[1008]&~m[1009]&m[1011]&m[1012])|(m[962]&m[1008]&~m[1009]&m[1011]&m[1012])|(~m[962]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[962]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[962]&m[1008]&m[1009]&m[1011]&m[1012]))):InitCond[1136];
    m[1015] = run?((((m[967]&~m[1013]&~m[1014]&~m[1016]&~m[1017])|(~m[967]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(m[967]&m[1013]&~m[1014]&m[1016]&~m[1017])|(m[967]&~m[1013]&m[1014]&m[1016]&~m[1017])|(~m[967]&m[1013]&~m[1014]&~m[1016]&m[1017])|(~m[967]&~m[1013]&m[1014]&~m[1016]&m[1017])|(m[967]&m[1013]&m[1014]&~m[1016]&m[1017])|(~m[967]&m[1013]&m[1014]&m[1016]&m[1017]))&UnbiasedRNG[438])|((m[967]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(~m[967]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[967]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[967]&m[1013]&~m[1014]&~m[1016]&m[1017])|(m[967]&~m[1013]&m[1014]&~m[1016]&m[1017])|(~m[967]&~m[1013]&~m[1014]&m[1016]&m[1017])|(m[967]&~m[1013]&~m[1014]&m[1016]&m[1017])|(~m[967]&m[1013]&~m[1014]&m[1016]&m[1017])|(m[967]&m[1013]&~m[1014]&m[1016]&m[1017])|(~m[967]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[967]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[967]&m[1013]&m[1014]&m[1016]&m[1017]))):InitCond[1137];
    m[1020] = run?((((m[972]&~m[1018]&~m[1019]&~m[1021]&~m[1022])|(~m[972]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(m[972]&m[1018]&~m[1019]&m[1021]&~m[1022])|(m[972]&~m[1018]&m[1019]&m[1021]&~m[1022])|(~m[972]&m[1018]&~m[1019]&~m[1021]&m[1022])|(~m[972]&~m[1018]&m[1019]&~m[1021]&m[1022])|(m[972]&m[1018]&m[1019]&~m[1021]&m[1022])|(~m[972]&m[1018]&m[1019]&m[1021]&m[1022]))&UnbiasedRNG[439])|((m[972]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(~m[972]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[972]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[972]&m[1018]&~m[1019]&~m[1021]&m[1022])|(m[972]&~m[1018]&m[1019]&~m[1021]&m[1022])|(~m[972]&~m[1018]&~m[1019]&m[1021]&m[1022])|(m[972]&~m[1018]&~m[1019]&m[1021]&m[1022])|(~m[972]&m[1018]&~m[1019]&m[1021]&m[1022])|(m[972]&m[1018]&~m[1019]&m[1021]&m[1022])|(~m[972]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[972]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[972]&m[1018]&m[1019]&m[1021]&m[1022]))):InitCond[1138];
    m[1025] = run?((((m[977]&~m[1023]&~m[1024]&~m[1026]&~m[1027])|(~m[977]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(m[977]&m[1023]&~m[1024]&m[1026]&~m[1027])|(m[977]&~m[1023]&m[1024]&m[1026]&~m[1027])|(~m[977]&m[1023]&~m[1024]&~m[1026]&m[1027])|(~m[977]&~m[1023]&m[1024]&~m[1026]&m[1027])|(m[977]&m[1023]&m[1024]&~m[1026]&m[1027])|(~m[977]&m[1023]&m[1024]&m[1026]&m[1027]))&UnbiasedRNG[440])|((m[977]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(~m[977]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[977]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[977]&m[1023]&~m[1024]&~m[1026]&m[1027])|(m[977]&~m[1023]&m[1024]&~m[1026]&m[1027])|(~m[977]&~m[1023]&~m[1024]&m[1026]&m[1027])|(m[977]&~m[1023]&~m[1024]&m[1026]&m[1027])|(~m[977]&m[1023]&~m[1024]&m[1026]&m[1027])|(m[977]&m[1023]&~m[1024]&m[1026]&m[1027])|(~m[977]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[977]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[977]&m[1023]&m[1024]&m[1026]&m[1027]))):InitCond[1139];
    m[1030] = run?((((m[982]&~m[1028]&~m[1029]&~m[1031]&~m[1032])|(~m[982]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(m[982]&m[1028]&~m[1029]&m[1031]&~m[1032])|(m[982]&~m[1028]&m[1029]&m[1031]&~m[1032])|(~m[982]&m[1028]&~m[1029]&~m[1031]&m[1032])|(~m[982]&~m[1028]&m[1029]&~m[1031]&m[1032])|(m[982]&m[1028]&m[1029]&~m[1031]&m[1032])|(~m[982]&m[1028]&m[1029]&m[1031]&m[1032]))&UnbiasedRNG[441])|((m[982]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(~m[982]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[982]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[982]&m[1028]&~m[1029]&~m[1031]&m[1032])|(m[982]&~m[1028]&m[1029]&~m[1031]&m[1032])|(~m[982]&~m[1028]&~m[1029]&m[1031]&m[1032])|(m[982]&~m[1028]&~m[1029]&m[1031]&m[1032])|(~m[982]&m[1028]&~m[1029]&m[1031]&m[1032])|(m[982]&m[1028]&~m[1029]&m[1031]&m[1032])|(~m[982]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[982]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[982]&m[1028]&m[1029]&m[1031]&m[1032]))):InitCond[1140];
    m[1035] = run?((((m[987]&~m[1033]&~m[1034]&~m[1036]&~m[1037])|(~m[987]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(m[987]&m[1033]&~m[1034]&m[1036]&~m[1037])|(m[987]&~m[1033]&m[1034]&m[1036]&~m[1037])|(~m[987]&m[1033]&~m[1034]&~m[1036]&m[1037])|(~m[987]&~m[1033]&m[1034]&~m[1036]&m[1037])|(m[987]&m[1033]&m[1034]&~m[1036]&m[1037])|(~m[987]&m[1033]&m[1034]&m[1036]&m[1037]))&UnbiasedRNG[442])|((m[987]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(~m[987]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[987]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[987]&m[1033]&~m[1034]&~m[1036]&m[1037])|(m[987]&~m[1033]&m[1034]&~m[1036]&m[1037])|(~m[987]&~m[1033]&~m[1034]&m[1036]&m[1037])|(m[987]&~m[1033]&~m[1034]&m[1036]&m[1037])|(~m[987]&m[1033]&~m[1034]&m[1036]&m[1037])|(m[987]&m[1033]&~m[1034]&m[1036]&m[1037])|(~m[987]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[987]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[987]&m[1033]&m[1034]&m[1036]&m[1037]))):InitCond[1141];
    m[1040] = run?((((m[992]&~m[1038]&~m[1039]&~m[1041]&~m[1042])|(~m[992]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(m[992]&m[1038]&~m[1039]&m[1041]&~m[1042])|(m[992]&~m[1038]&m[1039]&m[1041]&~m[1042])|(~m[992]&m[1038]&~m[1039]&~m[1041]&m[1042])|(~m[992]&~m[1038]&m[1039]&~m[1041]&m[1042])|(m[992]&m[1038]&m[1039]&~m[1041]&m[1042])|(~m[992]&m[1038]&m[1039]&m[1041]&m[1042]))&UnbiasedRNG[443])|((m[992]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(~m[992]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[992]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[992]&m[1038]&~m[1039]&~m[1041]&m[1042])|(m[992]&~m[1038]&m[1039]&~m[1041]&m[1042])|(~m[992]&~m[1038]&~m[1039]&m[1041]&m[1042])|(m[992]&~m[1038]&~m[1039]&m[1041]&m[1042])|(~m[992]&m[1038]&~m[1039]&m[1041]&m[1042])|(m[992]&m[1038]&~m[1039]&m[1041]&m[1042])|(~m[992]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[992]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[992]&m[1038]&m[1039]&m[1041]&m[1042]))):InitCond[1142];
    m[1045] = run?((((m[997]&~m[1043]&~m[1044]&~m[1046]&~m[1047])|(~m[997]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(m[997]&m[1043]&~m[1044]&m[1046]&~m[1047])|(m[997]&~m[1043]&m[1044]&m[1046]&~m[1047])|(~m[997]&m[1043]&~m[1044]&~m[1046]&m[1047])|(~m[997]&~m[1043]&m[1044]&~m[1046]&m[1047])|(m[997]&m[1043]&m[1044]&~m[1046]&m[1047])|(~m[997]&m[1043]&m[1044]&m[1046]&m[1047]))&UnbiasedRNG[444])|((m[997]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(~m[997]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[997]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[997]&m[1043]&~m[1044]&~m[1046]&m[1047])|(m[997]&~m[1043]&m[1044]&~m[1046]&m[1047])|(~m[997]&~m[1043]&~m[1044]&m[1046]&m[1047])|(m[997]&~m[1043]&~m[1044]&m[1046]&m[1047])|(~m[997]&m[1043]&~m[1044]&m[1046]&m[1047])|(m[997]&m[1043]&~m[1044]&m[1046]&m[1047])|(~m[997]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[997]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[997]&m[1043]&m[1044]&m[1046]&m[1047]))):InitCond[1143];
    m[1050] = run?((((m[1002]&~m[1048]&~m[1049]&~m[1051]&~m[1052])|(~m[1002]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1002]&m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1002]&~m[1048]&m[1049]&m[1051]&~m[1052])|(~m[1002]&m[1048]&~m[1049]&~m[1051]&m[1052])|(~m[1002]&~m[1048]&m[1049]&~m[1051]&m[1052])|(m[1002]&m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1002]&m[1048]&m[1049]&m[1051]&m[1052]))&UnbiasedRNG[445])|((m[1002]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(~m[1002]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1002]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1002]&m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1002]&~m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1002]&~m[1048]&~m[1049]&m[1051]&m[1052])|(m[1002]&~m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1002]&m[1048]&~m[1049]&m[1051]&m[1052])|(m[1002]&m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1002]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1002]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1002]&m[1048]&m[1049]&m[1051]&m[1052]))):InitCond[1144];
    m[1060] = run?((((m[1007]&~m[1058]&~m[1059]&~m[1061]&~m[1062])|(~m[1007]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1007]&m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1007]&~m[1058]&m[1059]&m[1061]&~m[1062])|(~m[1007]&m[1058]&~m[1059]&~m[1061]&m[1062])|(~m[1007]&~m[1058]&m[1059]&~m[1061]&m[1062])|(m[1007]&m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1007]&m[1058]&m[1059]&m[1061]&m[1062]))&UnbiasedRNG[446])|((m[1007]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(~m[1007]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1007]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1007]&m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1007]&~m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1007]&~m[1058]&~m[1059]&m[1061]&m[1062])|(m[1007]&~m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1007]&m[1058]&~m[1059]&m[1061]&m[1062])|(m[1007]&m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1007]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1007]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1007]&m[1058]&m[1059]&m[1061]&m[1062]))):InitCond[1145];
    m[1065] = run?((((m[1012]&~m[1063]&~m[1064]&~m[1066]&~m[1067])|(~m[1012]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1012]&m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1012]&~m[1063]&m[1064]&m[1066]&~m[1067])|(~m[1012]&m[1063]&~m[1064]&~m[1066]&m[1067])|(~m[1012]&~m[1063]&m[1064]&~m[1066]&m[1067])|(m[1012]&m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1012]&m[1063]&m[1064]&m[1066]&m[1067]))&UnbiasedRNG[447])|((m[1012]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(~m[1012]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1012]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1012]&m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1012]&~m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1012]&~m[1063]&~m[1064]&m[1066]&m[1067])|(m[1012]&~m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1012]&m[1063]&~m[1064]&m[1066]&m[1067])|(m[1012]&m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1012]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1012]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1012]&m[1063]&m[1064]&m[1066]&m[1067]))):InitCond[1146];
    m[1070] = run?((((m[1017]&~m[1068]&~m[1069]&~m[1071]&~m[1072])|(~m[1017]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1017]&m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1017]&~m[1068]&m[1069]&m[1071]&~m[1072])|(~m[1017]&m[1068]&~m[1069]&~m[1071]&m[1072])|(~m[1017]&~m[1068]&m[1069]&~m[1071]&m[1072])|(m[1017]&m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1017]&m[1068]&m[1069]&m[1071]&m[1072]))&UnbiasedRNG[448])|((m[1017]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(~m[1017]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1017]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1017]&m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1017]&~m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1017]&~m[1068]&~m[1069]&m[1071]&m[1072])|(m[1017]&~m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1017]&m[1068]&~m[1069]&m[1071]&m[1072])|(m[1017]&m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1017]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1017]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1017]&m[1068]&m[1069]&m[1071]&m[1072]))):InitCond[1147];
    m[1075] = run?((((m[1022]&~m[1073]&~m[1074]&~m[1076]&~m[1077])|(~m[1022]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1022]&m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1022]&~m[1073]&m[1074]&m[1076]&~m[1077])|(~m[1022]&m[1073]&~m[1074]&~m[1076]&m[1077])|(~m[1022]&~m[1073]&m[1074]&~m[1076]&m[1077])|(m[1022]&m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1022]&m[1073]&m[1074]&m[1076]&m[1077]))&UnbiasedRNG[449])|((m[1022]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(~m[1022]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1022]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1022]&m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1022]&~m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1022]&~m[1073]&~m[1074]&m[1076]&m[1077])|(m[1022]&~m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1022]&m[1073]&~m[1074]&m[1076]&m[1077])|(m[1022]&m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1022]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1022]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1022]&m[1073]&m[1074]&m[1076]&m[1077]))):InitCond[1148];
    m[1080] = run?((((m[1027]&~m[1078]&~m[1079]&~m[1081]&~m[1082])|(~m[1027]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1027]&m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1027]&~m[1078]&m[1079]&m[1081]&~m[1082])|(~m[1027]&m[1078]&~m[1079]&~m[1081]&m[1082])|(~m[1027]&~m[1078]&m[1079]&~m[1081]&m[1082])|(m[1027]&m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1027]&m[1078]&m[1079]&m[1081]&m[1082]))&UnbiasedRNG[450])|((m[1027]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(~m[1027]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1027]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1027]&m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1027]&~m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1027]&~m[1078]&~m[1079]&m[1081]&m[1082])|(m[1027]&~m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1027]&m[1078]&~m[1079]&m[1081]&m[1082])|(m[1027]&m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1027]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1027]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1027]&m[1078]&m[1079]&m[1081]&m[1082]))):InitCond[1149];
    m[1085] = run?((((m[1032]&~m[1083]&~m[1084]&~m[1086]&~m[1087])|(~m[1032]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1032]&m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1032]&~m[1083]&m[1084]&m[1086]&~m[1087])|(~m[1032]&m[1083]&~m[1084]&~m[1086]&m[1087])|(~m[1032]&~m[1083]&m[1084]&~m[1086]&m[1087])|(m[1032]&m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1032]&m[1083]&m[1084]&m[1086]&m[1087]))&UnbiasedRNG[451])|((m[1032]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(~m[1032]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1032]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1032]&m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1032]&~m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1032]&~m[1083]&~m[1084]&m[1086]&m[1087])|(m[1032]&~m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1032]&m[1083]&~m[1084]&m[1086]&m[1087])|(m[1032]&m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1032]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1032]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1032]&m[1083]&m[1084]&m[1086]&m[1087]))):InitCond[1150];
    m[1090] = run?((((m[1037]&~m[1088]&~m[1089]&~m[1091]&~m[1092])|(~m[1037]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1037]&m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1037]&~m[1088]&m[1089]&m[1091]&~m[1092])|(~m[1037]&m[1088]&~m[1089]&~m[1091]&m[1092])|(~m[1037]&~m[1088]&m[1089]&~m[1091]&m[1092])|(m[1037]&m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1037]&m[1088]&m[1089]&m[1091]&m[1092]))&UnbiasedRNG[452])|((m[1037]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(~m[1037]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1037]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1037]&m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1037]&~m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1037]&~m[1088]&~m[1089]&m[1091]&m[1092])|(m[1037]&~m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1037]&m[1088]&~m[1089]&m[1091]&m[1092])|(m[1037]&m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1037]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1037]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1037]&m[1088]&m[1089]&m[1091]&m[1092]))):InitCond[1151];
    m[1095] = run?((((m[1042]&~m[1093]&~m[1094]&~m[1096]&~m[1097])|(~m[1042]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1042]&m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1042]&~m[1093]&m[1094]&m[1096]&~m[1097])|(~m[1042]&m[1093]&~m[1094]&~m[1096]&m[1097])|(~m[1042]&~m[1093]&m[1094]&~m[1096]&m[1097])|(m[1042]&m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1042]&m[1093]&m[1094]&m[1096]&m[1097]))&UnbiasedRNG[453])|((m[1042]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(~m[1042]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1042]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1042]&m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1042]&~m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1042]&~m[1093]&~m[1094]&m[1096]&m[1097])|(m[1042]&~m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1042]&m[1093]&~m[1094]&m[1096]&m[1097])|(m[1042]&m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1042]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1042]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1042]&m[1093]&m[1094]&m[1096]&m[1097]))):InitCond[1152];
    m[1100] = run?((((m[1047]&~m[1098]&~m[1099]&~m[1101]&~m[1102])|(~m[1047]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1047]&m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1047]&~m[1098]&m[1099]&m[1101]&~m[1102])|(~m[1047]&m[1098]&~m[1099]&~m[1101]&m[1102])|(~m[1047]&~m[1098]&m[1099]&~m[1101]&m[1102])|(m[1047]&m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1047]&m[1098]&m[1099]&m[1101]&m[1102]))&UnbiasedRNG[454])|((m[1047]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(~m[1047]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1047]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1047]&m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1047]&~m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1047]&~m[1098]&~m[1099]&m[1101]&m[1102])|(m[1047]&~m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1047]&m[1098]&~m[1099]&m[1101]&m[1102])|(m[1047]&m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1047]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1047]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1047]&m[1098]&m[1099]&m[1101]&m[1102]))):InitCond[1153];
    m[1105] = run?((((m[1052]&~m[1103]&~m[1104]&~m[1106]&~m[1107])|(~m[1052]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1052]&m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1052]&~m[1103]&m[1104]&m[1106]&~m[1107])|(~m[1052]&m[1103]&~m[1104]&~m[1106]&m[1107])|(~m[1052]&~m[1103]&m[1104]&~m[1106]&m[1107])|(m[1052]&m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1052]&m[1103]&m[1104]&m[1106]&m[1107]))&UnbiasedRNG[455])|((m[1052]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(~m[1052]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1052]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1052]&m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1052]&~m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1052]&~m[1103]&~m[1104]&m[1106]&m[1107])|(m[1052]&~m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1052]&m[1103]&~m[1104]&m[1106]&m[1107])|(m[1052]&m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1052]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1052]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1052]&m[1103]&m[1104]&m[1106]&m[1107]))):InitCond[1154];
    m[1110] = run?((((m[1057]&~m[1108]&~m[1109]&~m[1111]&~m[1112])|(~m[1057]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1057]&m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1057]&~m[1108]&m[1109]&m[1111]&~m[1112])|(~m[1057]&m[1108]&~m[1109]&~m[1111]&m[1112])|(~m[1057]&~m[1108]&m[1109]&~m[1111]&m[1112])|(m[1057]&m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1057]&m[1108]&m[1109]&m[1111]&m[1112]))&UnbiasedRNG[456])|((m[1057]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(~m[1057]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1057]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1057]&m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1057]&~m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1057]&~m[1108]&~m[1109]&m[1111]&m[1112])|(m[1057]&~m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1057]&m[1108]&~m[1109]&m[1111]&m[1112])|(m[1057]&m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1057]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1057]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1057]&m[1108]&m[1109]&m[1111]&m[1112]))):InitCond[1155];
    m[1120] = run?((((m[1062]&~m[1118]&~m[1119]&~m[1121]&~m[1122])|(~m[1062]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1062]&m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1062]&~m[1118]&m[1119]&m[1121]&~m[1122])|(~m[1062]&m[1118]&~m[1119]&~m[1121]&m[1122])|(~m[1062]&~m[1118]&m[1119]&~m[1121]&m[1122])|(m[1062]&m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1062]&m[1118]&m[1119]&m[1121]&m[1122]))&UnbiasedRNG[457])|((m[1062]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(~m[1062]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1062]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1062]&m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1062]&~m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1062]&~m[1118]&~m[1119]&m[1121]&m[1122])|(m[1062]&~m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1062]&m[1118]&~m[1119]&m[1121]&m[1122])|(m[1062]&m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1062]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1062]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1062]&m[1118]&m[1119]&m[1121]&m[1122]))):InitCond[1156];
    m[1125] = run?((((m[1067]&~m[1123]&~m[1124]&~m[1126]&~m[1127])|(~m[1067]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1067]&m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1067]&~m[1123]&m[1124]&m[1126]&~m[1127])|(~m[1067]&m[1123]&~m[1124]&~m[1126]&m[1127])|(~m[1067]&~m[1123]&m[1124]&~m[1126]&m[1127])|(m[1067]&m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1067]&m[1123]&m[1124]&m[1126]&m[1127]))&UnbiasedRNG[458])|((m[1067]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(~m[1067]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1067]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1067]&m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1067]&~m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1067]&~m[1123]&~m[1124]&m[1126]&m[1127])|(m[1067]&~m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1067]&m[1123]&~m[1124]&m[1126]&m[1127])|(m[1067]&m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1067]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1067]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1067]&m[1123]&m[1124]&m[1126]&m[1127]))):InitCond[1157];
    m[1130] = run?((((m[1072]&~m[1128]&~m[1129]&~m[1131]&~m[1132])|(~m[1072]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1072]&m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1072]&~m[1128]&m[1129]&m[1131]&~m[1132])|(~m[1072]&m[1128]&~m[1129]&~m[1131]&m[1132])|(~m[1072]&~m[1128]&m[1129]&~m[1131]&m[1132])|(m[1072]&m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1072]&m[1128]&m[1129]&m[1131]&m[1132]))&UnbiasedRNG[459])|((m[1072]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(~m[1072]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1072]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1072]&m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1072]&~m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1072]&~m[1128]&~m[1129]&m[1131]&m[1132])|(m[1072]&~m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1072]&m[1128]&~m[1129]&m[1131]&m[1132])|(m[1072]&m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1072]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1072]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1072]&m[1128]&m[1129]&m[1131]&m[1132]))):InitCond[1158];
    m[1135] = run?((((m[1077]&~m[1133]&~m[1134]&~m[1136]&~m[1137])|(~m[1077]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1077]&m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1077]&~m[1133]&m[1134]&m[1136]&~m[1137])|(~m[1077]&m[1133]&~m[1134]&~m[1136]&m[1137])|(~m[1077]&~m[1133]&m[1134]&~m[1136]&m[1137])|(m[1077]&m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1077]&m[1133]&m[1134]&m[1136]&m[1137]))&UnbiasedRNG[460])|((m[1077]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(~m[1077]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1077]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1077]&m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1077]&~m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1077]&~m[1133]&~m[1134]&m[1136]&m[1137])|(m[1077]&~m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1077]&m[1133]&~m[1134]&m[1136]&m[1137])|(m[1077]&m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1077]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1077]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1077]&m[1133]&m[1134]&m[1136]&m[1137]))):InitCond[1159];
    m[1140] = run?((((m[1082]&~m[1138]&~m[1139]&~m[1141]&~m[1142])|(~m[1082]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1082]&m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1082]&~m[1138]&m[1139]&m[1141]&~m[1142])|(~m[1082]&m[1138]&~m[1139]&~m[1141]&m[1142])|(~m[1082]&~m[1138]&m[1139]&~m[1141]&m[1142])|(m[1082]&m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1082]&m[1138]&m[1139]&m[1141]&m[1142]))&UnbiasedRNG[461])|((m[1082]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(~m[1082]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1082]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1082]&m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1082]&~m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1082]&~m[1138]&~m[1139]&m[1141]&m[1142])|(m[1082]&~m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1082]&m[1138]&~m[1139]&m[1141]&m[1142])|(m[1082]&m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1082]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1082]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1082]&m[1138]&m[1139]&m[1141]&m[1142]))):InitCond[1160];
    m[1145] = run?((((m[1087]&~m[1143]&~m[1144]&~m[1146]&~m[1147])|(~m[1087]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1087]&m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1087]&~m[1143]&m[1144]&m[1146]&~m[1147])|(~m[1087]&m[1143]&~m[1144]&~m[1146]&m[1147])|(~m[1087]&~m[1143]&m[1144]&~m[1146]&m[1147])|(m[1087]&m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1087]&m[1143]&m[1144]&m[1146]&m[1147]))&UnbiasedRNG[462])|((m[1087]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(~m[1087]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1087]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1087]&m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1087]&~m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1087]&~m[1143]&~m[1144]&m[1146]&m[1147])|(m[1087]&~m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1087]&m[1143]&~m[1144]&m[1146]&m[1147])|(m[1087]&m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1087]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1087]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1087]&m[1143]&m[1144]&m[1146]&m[1147]))):InitCond[1161];
    m[1150] = run?((((m[1092]&~m[1148]&~m[1149]&~m[1151]&~m[1152])|(~m[1092]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1092]&m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1092]&~m[1148]&m[1149]&m[1151]&~m[1152])|(~m[1092]&m[1148]&~m[1149]&~m[1151]&m[1152])|(~m[1092]&~m[1148]&m[1149]&~m[1151]&m[1152])|(m[1092]&m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1092]&m[1148]&m[1149]&m[1151]&m[1152]))&UnbiasedRNG[463])|((m[1092]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(~m[1092]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1092]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1092]&m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1092]&~m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1092]&~m[1148]&~m[1149]&m[1151]&m[1152])|(m[1092]&~m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1092]&m[1148]&~m[1149]&m[1151]&m[1152])|(m[1092]&m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1092]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1092]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1092]&m[1148]&m[1149]&m[1151]&m[1152]))):InitCond[1162];
    m[1155] = run?((((m[1097]&~m[1153]&~m[1154]&~m[1156]&~m[1157])|(~m[1097]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1097]&m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1097]&~m[1153]&m[1154]&m[1156]&~m[1157])|(~m[1097]&m[1153]&~m[1154]&~m[1156]&m[1157])|(~m[1097]&~m[1153]&m[1154]&~m[1156]&m[1157])|(m[1097]&m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1097]&m[1153]&m[1154]&m[1156]&m[1157]))&UnbiasedRNG[464])|((m[1097]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(~m[1097]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1097]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1097]&m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1097]&~m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1097]&~m[1153]&~m[1154]&m[1156]&m[1157])|(m[1097]&~m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1097]&m[1153]&~m[1154]&m[1156]&m[1157])|(m[1097]&m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1097]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1097]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1097]&m[1153]&m[1154]&m[1156]&m[1157]))):InitCond[1163];
    m[1160] = run?((((m[1102]&~m[1158]&~m[1159]&~m[1161]&~m[1162])|(~m[1102]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1102]&m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1102]&~m[1158]&m[1159]&m[1161]&~m[1162])|(~m[1102]&m[1158]&~m[1159]&~m[1161]&m[1162])|(~m[1102]&~m[1158]&m[1159]&~m[1161]&m[1162])|(m[1102]&m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1102]&m[1158]&m[1159]&m[1161]&m[1162]))&UnbiasedRNG[465])|((m[1102]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(~m[1102]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1102]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1102]&m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1102]&~m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1102]&~m[1158]&~m[1159]&m[1161]&m[1162])|(m[1102]&~m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1102]&m[1158]&~m[1159]&m[1161]&m[1162])|(m[1102]&m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1102]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1102]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1102]&m[1158]&m[1159]&m[1161]&m[1162]))):InitCond[1164];
    m[1165] = run?((((m[1107]&~m[1163]&~m[1164]&~m[1166]&~m[1167])|(~m[1107]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1107]&m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1107]&~m[1163]&m[1164]&m[1166]&~m[1167])|(~m[1107]&m[1163]&~m[1164]&~m[1166]&m[1167])|(~m[1107]&~m[1163]&m[1164]&~m[1166]&m[1167])|(m[1107]&m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1107]&m[1163]&m[1164]&m[1166]&m[1167]))&UnbiasedRNG[466])|((m[1107]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(~m[1107]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1107]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1107]&m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1107]&~m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1107]&~m[1163]&~m[1164]&m[1166]&m[1167])|(m[1107]&~m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1107]&m[1163]&~m[1164]&m[1166]&m[1167])|(m[1107]&m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1107]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1107]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1107]&m[1163]&m[1164]&m[1166]&m[1167]))):InitCond[1165];
    m[1170] = run?((((m[1112]&~m[1168]&~m[1169]&~m[1171]&~m[1172])|(~m[1112]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1112]&m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1112]&~m[1168]&m[1169]&m[1171]&~m[1172])|(~m[1112]&m[1168]&~m[1169]&~m[1171]&m[1172])|(~m[1112]&~m[1168]&m[1169]&~m[1171]&m[1172])|(m[1112]&m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1112]&m[1168]&m[1169]&m[1171]&m[1172]))&UnbiasedRNG[467])|((m[1112]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(~m[1112]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1112]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1112]&m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1112]&~m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1112]&~m[1168]&~m[1169]&m[1171]&m[1172])|(m[1112]&~m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1112]&m[1168]&~m[1169]&m[1171]&m[1172])|(m[1112]&m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1112]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1112]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1112]&m[1168]&m[1169]&m[1171]&m[1172]))):InitCond[1166];
    m[1175] = run?((((m[1117]&~m[1173]&~m[1174]&~m[1176]&~m[1177])|(~m[1117]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1117]&m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1117]&~m[1173]&m[1174]&m[1176]&~m[1177])|(~m[1117]&m[1173]&~m[1174]&~m[1176]&m[1177])|(~m[1117]&~m[1173]&m[1174]&~m[1176]&m[1177])|(m[1117]&m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1117]&m[1173]&m[1174]&m[1176]&m[1177]))&UnbiasedRNG[468])|((m[1117]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(~m[1117]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1117]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1117]&m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1117]&~m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1117]&~m[1173]&~m[1174]&m[1176]&m[1177])|(m[1117]&~m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1117]&m[1173]&~m[1174]&m[1176]&m[1177])|(m[1117]&m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1117]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1117]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1117]&m[1173]&m[1174]&m[1176]&m[1177]))):InitCond[1167];
    m[1185] = run?((((m[1122]&~m[1183]&~m[1184]&~m[1186]&~m[1187])|(~m[1122]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1122]&m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1122]&~m[1183]&m[1184]&m[1186]&~m[1187])|(~m[1122]&m[1183]&~m[1184]&~m[1186]&m[1187])|(~m[1122]&~m[1183]&m[1184]&~m[1186]&m[1187])|(m[1122]&m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1122]&m[1183]&m[1184]&m[1186]&m[1187]))&UnbiasedRNG[469])|((m[1122]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(~m[1122]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1122]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1122]&m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1122]&~m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1122]&~m[1183]&~m[1184]&m[1186]&m[1187])|(m[1122]&~m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1122]&m[1183]&~m[1184]&m[1186]&m[1187])|(m[1122]&m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1122]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1122]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1122]&m[1183]&m[1184]&m[1186]&m[1187]))):InitCond[1168];
    m[1190] = run?((((m[1127]&~m[1188]&~m[1189]&~m[1191]&~m[1192])|(~m[1127]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1127]&m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1127]&~m[1188]&m[1189]&m[1191]&~m[1192])|(~m[1127]&m[1188]&~m[1189]&~m[1191]&m[1192])|(~m[1127]&~m[1188]&m[1189]&~m[1191]&m[1192])|(m[1127]&m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1127]&m[1188]&m[1189]&m[1191]&m[1192]))&UnbiasedRNG[470])|((m[1127]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(~m[1127]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1127]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1127]&m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1127]&~m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1127]&~m[1188]&~m[1189]&m[1191]&m[1192])|(m[1127]&~m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1127]&m[1188]&~m[1189]&m[1191]&m[1192])|(m[1127]&m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1127]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1127]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1127]&m[1188]&m[1189]&m[1191]&m[1192]))):InitCond[1169];
    m[1195] = run?((((m[1132]&~m[1193]&~m[1194]&~m[1196]&~m[1197])|(~m[1132]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1132]&m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1132]&~m[1193]&m[1194]&m[1196]&~m[1197])|(~m[1132]&m[1193]&~m[1194]&~m[1196]&m[1197])|(~m[1132]&~m[1193]&m[1194]&~m[1196]&m[1197])|(m[1132]&m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1132]&m[1193]&m[1194]&m[1196]&m[1197]))&UnbiasedRNG[471])|((m[1132]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(~m[1132]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1132]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1132]&m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1132]&~m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1132]&~m[1193]&~m[1194]&m[1196]&m[1197])|(m[1132]&~m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1132]&m[1193]&~m[1194]&m[1196]&m[1197])|(m[1132]&m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1132]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1132]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1132]&m[1193]&m[1194]&m[1196]&m[1197]))):InitCond[1170];
    m[1200] = run?((((m[1137]&~m[1198]&~m[1199]&~m[1201]&~m[1202])|(~m[1137]&~m[1198]&~m[1199]&m[1201]&~m[1202])|(m[1137]&m[1198]&~m[1199]&m[1201]&~m[1202])|(m[1137]&~m[1198]&m[1199]&m[1201]&~m[1202])|(~m[1137]&m[1198]&~m[1199]&~m[1201]&m[1202])|(~m[1137]&~m[1198]&m[1199]&~m[1201]&m[1202])|(m[1137]&m[1198]&m[1199]&~m[1201]&m[1202])|(~m[1137]&m[1198]&m[1199]&m[1201]&m[1202]))&UnbiasedRNG[472])|((m[1137]&~m[1198]&~m[1199]&m[1201]&~m[1202])|(~m[1137]&~m[1198]&~m[1199]&~m[1201]&m[1202])|(m[1137]&~m[1198]&~m[1199]&~m[1201]&m[1202])|(m[1137]&m[1198]&~m[1199]&~m[1201]&m[1202])|(m[1137]&~m[1198]&m[1199]&~m[1201]&m[1202])|(~m[1137]&~m[1198]&~m[1199]&m[1201]&m[1202])|(m[1137]&~m[1198]&~m[1199]&m[1201]&m[1202])|(~m[1137]&m[1198]&~m[1199]&m[1201]&m[1202])|(m[1137]&m[1198]&~m[1199]&m[1201]&m[1202])|(~m[1137]&~m[1198]&m[1199]&m[1201]&m[1202])|(m[1137]&~m[1198]&m[1199]&m[1201]&m[1202])|(m[1137]&m[1198]&m[1199]&m[1201]&m[1202]))):InitCond[1171];
    m[1205] = run?((((m[1142]&~m[1203]&~m[1204]&~m[1206]&~m[1207])|(~m[1142]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1142]&m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1142]&~m[1203]&m[1204]&m[1206]&~m[1207])|(~m[1142]&m[1203]&~m[1204]&~m[1206]&m[1207])|(~m[1142]&~m[1203]&m[1204]&~m[1206]&m[1207])|(m[1142]&m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1142]&m[1203]&m[1204]&m[1206]&m[1207]))&UnbiasedRNG[473])|((m[1142]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(~m[1142]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1142]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1142]&m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1142]&~m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1142]&~m[1203]&~m[1204]&m[1206]&m[1207])|(m[1142]&~m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1142]&m[1203]&~m[1204]&m[1206]&m[1207])|(m[1142]&m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1142]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1142]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1142]&m[1203]&m[1204]&m[1206]&m[1207]))):InitCond[1172];
    m[1210] = run?((((m[1147]&~m[1208]&~m[1209]&~m[1211]&~m[1212])|(~m[1147]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1147]&m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1147]&~m[1208]&m[1209]&m[1211]&~m[1212])|(~m[1147]&m[1208]&~m[1209]&~m[1211]&m[1212])|(~m[1147]&~m[1208]&m[1209]&~m[1211]&m[1212])|(m[1147]&m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1147]&m[1208]&m[1209]&m[1211]&m[1212]))&UnbiasedRNG[474])|((m[1147]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(~m[1147]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1147]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1147]&m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1147]&~m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1147]&~m[1208]&~m[1209]&m[1211]&m[1212])|(m[1147]&~m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1147]&m[1208]&~m[1209]&m[1211]&m[1212])|(m[1147]&m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1147]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1147]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1147]&m[1208]&m[1209]&m[1211]&m[1212]))):InitCond[1173];
    m[1215] = run?((((m[1152]&~m[1213]&~m[1214]&~m[1216]&~m[1217])|(~m[1152]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1152]&m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1152]&~m[1213]&m[1214]&m[1216]&~m[1217])|(~m[1152]&m[1213]&~m[1214]&~m[1216]&m[1217])|(~m[1152]&~m[1213]&m[1214]&~m[1216]&m[1217])|(m[1152]&m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1152]&m[1213]&m[1214]&m[1216]&m[1217]))&UnbiasedRNG[475])|((m[1152]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(~m[1152]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1152]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1152]&m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1152]&~m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1152]&~m[1213]&~m[1214]&m[1216]&m[1217])|(m[1152]&~m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1152]&m[1213]&~m[1214]&m[1216]&m[1217])|(m[1152]&m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1152]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1152]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1152]&m[1213]&m[1214]&m[1216]&m[1217]))):InitCond[1174];
    m[1220] = run?((((m[1157]&~m[1218]&~m[1219]&~m[1221]&~m[1222])|(~m[1157]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1157]&m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1157]&~m[1218]&m[1219]&m[1221]&~m[1222])|(~m[1157]&m[1218]&~m[1219]&~m[1221]&m[1222])|(~m[1157]&~m[1218]&m[1219]&~m[1221]&m[1222])|(m[1157]&m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1157]&m[1218]&m[1219]&m[1221]&m[1222]))&UnbiasedRNG[476])|((m[1157]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(~m[1157]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1157]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1157]&m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1157]&~m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1157]&~m[1218]&~m[1219]&m[1221]&m[1222])|(m[1157]&~m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1157]&m[1218]&~m[1219]&m[1221]&m[1222])|(m[1157]&m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1157]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1157]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1157]&m[1218]&m[1219]&m[1221]&m[1222]))):InitCond[1175];
    m[1225] = run?((((m[1162]&~m[1223]&~m[1224]&~m[1226]&~m[1227])|(~m[1162]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1162]&m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1162]&~m[1223]&m[1224]&m[1226]&~m[1227])|(~m[1162]&m[1223]&~m[1224]&~m[1226]&m[1227])|(~m[1162]&~m[1223]&m[1224]&~m[1226]&m[1227])|(m[1162]&m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1162]&m[1223]&m[1224]&m[1226]&m[1227]))&UnbiasedRNG[477])|((m[1162]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(~m[1162]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1162]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1162]&m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1162]&~m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1162]&~m[1223]&~m[1224]&m[1226]&m[1227])|(m[1162]&~m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1162]&m[1223]&~m[1224]&m[1226]&m[1227])|(m[1162]&m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1162]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1162]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1162]&m[1223]&m[1224]&m[1226]&m[1227]))):InitCond[1176];
    m[1230] = run?((((m[1167]&~m[1228]&~m[1229]&~m[1231]&~m[1232])|(~m[1167]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1167]&m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1167]&~m[1228]&m[1229]&m[1231]&~m[1232])|(~m[1167]&m[1228]&~m[1229]&~m[1231]&m[1232])|(~m[1167]&~m[1228]&m[1229]&~m[1231]&m[1232])|(m[1167]&m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1167]&m[1228]&m[1229]&m[1231]&m[1232]))&UnbiasedRNG[478])|((m[1167]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(~m[1167]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1167]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1167]&m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1167]&~m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1167]&~m[1228]&~m[1229]&m[1231]&m[1232])|(m[1167]&~m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1167]&m[1228]&~m[1229]&m[1231]&m[1232])|(m[1167]&m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1167]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1167]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1167]&m[1228]&m[1229]&m[1231]&m[1232]))):InitCond[1177];
    m[1235] = run?((((m[1172]&~m[1233]&~m[1234]&~m[1236]&~m[1237])|(~m[1172]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1172]&m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1172]&~m[1233]&m[1234]&m[1236]&~m[1237])|(~m[1172]&m[1233]&~m[1234]&~m[1236]&m[1237])|(~m[1172]&~m[1233]&m[1234]&~m[1236]&m[1237])|(m[1172]&m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1172]&m[1233]&m[1234]&m[1236]&m[1237]))&UnbiasedRNG[479])|((m[1172]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(~m[1172]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1172]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1172]&m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1172]&~m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1172]&~m[1233]&~m[1234]&m[1236]&m[1237])|(m[1172]&~m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1172]&m[1233]&~m[1234]&m[1236]&m[1237])|(m[1172]&m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1172]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1172]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1172]&m[1233]&m[1234]&m[1236]&m[1237]))):InitCond[1178];
    m[1240] = run?((((m[1177]&~m[1238]&~m[1239]&~m[1241]&~m[1242])|(~m[1177]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1177]&m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1177]&~m[1238]&m[1239]&m[1241]&~m[1242])|(~m[1177]&m[1238]&~m[1239]&~m[1241]&m[1242])|(~m[1177]&~m[1238]&m[1239]&~m[1241]&m[1242])|(m[1177]&m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1177]&m[1238]&m[1239]&m[1241]&m[1242]))&UnbiasedRNG[480])|((m[1177]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(~m[1177]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1177]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1177]&m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1177]&~m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1177]&~m[1238]&~m[1239]&m[1241]&m[1242])|(m[1177]&~m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1177]&m[1238]&~m[1239]&m[1241]&m[1242])|(m[1177]&m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1177]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1177]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1177]&m[1238]&m[1239]&m[1241]&m[1242]))):InitCond[1179];
    m[1245] = run?((((m[1182]&~m[1243]&~m[1244]&~m[1246]&~m[1247])|(~m[1182]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1182]&m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1182]&~m[1243]&m[1244]&m[1246]&~m[1247])|(~m[1182]&m[1243]&~m[1244]&~m[1246]&m[1247])|(~m[1182]&~m[1243]&m[1244]&~m[1246]&m[1247])|(m[1182]&m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1182]&m[1243]&m[1244]&m[1246]&m[1247]))&UnbiasedRNG[481])|((m[1182]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(~m[1182]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1182]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1182]&m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1182]&~m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1182]&~m[1243]&~m[1244]&m[1246]&m[1247])|(m[1182]&~m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1182]&m[1243]&~m[1244]&m[1246]&m[1247])|(m[1182]&m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1182]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1182]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1182]&m[1243]&m[1244]&m[1246]&m[1247]))):InitCond[1180];
    m[1250] = run?((((m[1192]&~m[1248]&~m[1249]&~m[1251]&~m[1252])|(~m[1192]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1192]&m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1192]&~m[1248]&m[1249]&m[1251]&~m[1252])|(~m[1192]&m[1248]&~m[1249]&~m[1251]&m[1252])|(~m[1192]&~m[1248]&m[1249]&~m[1251]&m[1252])|(m[1192]&m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1192]&m[1248]&m[1249]&m[1251]&m[1252]))&UnbiasedRNG[482])|((m[1192]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(~m[1192]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1192]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1192]&m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1192]&~m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1192]&~m[1248]&~m[1249]&m[1251]&m[1252])|(m[1192]&~m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1192]&m[1248]&~m[1249]&m[1251]&m[1252])|(m[1192]&m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1192]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1192]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1192]&m[1248]&m[1249]&m[1251]&m[1252]))):InitCond[1181];
    m[1255] = run?((((m[1197]&~m[1253]&~m[1254]&~m[1256]&~m[1257])|(~m[1197]&~m[1253]&~m[1254]&m[1256]&~m[1257])|(m[1197]&m[1253]&~m[1254]&m[1256]&~m[1257])|(m[1197]&~m[1253]&m[1254]&m[1256]&~m[1257])|(~m[1197]&m[1253]&~m[1254]&~m[1256]&m[1257])|(~m[1197]&~m[1253]&m[1254]&~m[1256]&m[1257])|(m[1197]&m[1253]&m[1254]&~m[1256]&m[1257])|(~m[1197]&m[1253]&m[1254]&m[1256]&m[1257]))&UnbiasedRNG[483])|((m[1197]&~m[1253]&~m[1254]&m[1256]&~m[1257])|(~m[1197]&~m[1253]&~m[1254]&~m[1256]&m[1257])|(m[1197]&~m[1253]&~m[1254]&~m[1256]&m[1257])|(m[1197]&m[1253]&~m[1254]&~m[1256]&m[1257])|(m[1197]&~m[1253]&m[1254]&~m[1256]&m[1257])|(~m[1197]&~m[1253]&~m[1254]&m[1256]&m[1257])|(m[1197]&~m[1253]&~m[1254]&m[1256]&m[1257])|(~m[1197]&m[1253]&~m[1254]&m[1256]&m[1257])|(m[1197]&m[1253]&~m[1254]&m[1256]&m[1257])|(~m[1197]&~m[1253]&m[1254]&m[1256]&m[1257])|(m[1197]&~m[1253]&m[1254]&m[1256]&m[1257])|(m[1197]&m[1253]&m[1254]&m[1256]&m[1257]))):InitCond[1182];
    m[1260] = run?((((m[1202]&~m[1258]&~m[1259]&~m[1261]&~m[1262])|(~m[1202]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1202]&m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1202]&~m[1258]&m[1259]&m[1261]&~m[1262])|(~m[1202]&m[1258]&~m[1259]&~m[1261]&m[1262])|(~m[1202]&~m[1258]&m[1259]&~m[1261]&m[1262])|(m[1202]&m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1202]&m[1258]&m[1259]&m[1261]&m[1262]))&UnbiasedRNG[484])|((m[1202]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(~m[1202]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1202]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1202]&m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1202]&~m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1202]&~m[1258]&~m[1259]&m[1261]&m[1262])|(m[1202]&~m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1202]&m[1258]&~m[1259]&m[1261]&m[1262])|(m[1202]&m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1202]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1202]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1202]&m[1258]&m[1259]&m[1261]&m[1262]))):InitCond[1183];
    m[1265] = run?((((m[1207]&~m[1263]&~m[1264]&~m[1266]&~m[1267])|(~m[1207]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1207]&m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1207]&~m[1263]&m[1264]&m[1266]&~m[1267])|(~m[1207]&m[1263]&~m[1264]&~m[1266]&m[1267])|(~m[1207]&~m[1263]&m[1264]&~m[1266]&m[1267])|(m[1207]&m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1207]&m[1263]&m[1264]&m[1266]&m[1267]))&UnbiasedRNG[485])|((m[1207]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(~m[1207]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1207]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1207]&m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1207]&~m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1207]&~m[1263]&~m[1264]&m[1266]&m[1267])|(m[1207]&~m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1207]&m[1263]&~m[1264]&m[1266]&m[1267])|(m[1207]&m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1207]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1207]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1207]&m[1263]&m[1264]&m[1266]&m[1267]))):InitCond[1184];
    m[1270] = run?((((m[1212]&~m[1268]&~m[1269]&~m[1271]&~m[1272])|(~m[1212]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1212]&m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1212]&~m[1268]&m[1269]&m[1271]&~m[1272])|(~m[1212]&m[1268]&~m[1269]&~m[1271]&m[1272])|(~m[1212]&~m[1268]&m[1269]&~m[1271]&m[1272])|(m[1212]&m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1212]&m[1268]&m[1269]&m[1271]&m[1272]))&UnbiasedRNG[486])|((m[1212]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(~m[1212]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1212]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1212]&m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1212]&~m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1212]&~m[1268]&~m[1269]&m[1271]&m[1272])|(m[1212]&~m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1212]&m[1268]&~m[1269]&m[1271]&m[1272])|(m[1212]&m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1212]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1212]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1212]&m[1268]&m[1269]&m[1271]&m[1272]))):InitCond[1185];
    m[1275] = run?((((m[1217]&~m[1273]&~m[1274]&~m[1276]&~m[1277])|(~m[1217]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1217]&m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1217]&~m[1273]&m[1274]&m[1276]&~m[1277])|(~m[1217]&m[1273]&~m[1274]&~m[1276]&m[1277])|(~m[1217]&~m[1273]&m[1274]&~m[1276]&m[1277])|(m[1217]&m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1217]&m[1273]&m[1274]&m[1276]&m[1277]))&UnbiasedRNG[487])|((m[1217]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(~m[1217]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1217]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1217]&m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1217]&~m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1217]&~m[1273]&~m[1274]&m[1276]&m[1277])|(m[1217]&~m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1217]&m[1273]&~m[1274]&m[1276]&m[1277])|(m[1217]&m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1217]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1217]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1217]&m[1273]&m[1274]&m[1276]&m[1277]))):InitCond[1186];
    m[1280] = run?((((m[1222]&~m[1278]&~m[1279]&~m[1281]&~m[1282])|(~m[1222]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1222]&m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1222]&~m[1278]&m[1279]&m[1281]&~m[1282])|(~m[1222]&m[1278]&~m[1279]&~m[1281]&m[1282])|(~m[1222]&~m[1278]&m[1279]&~m[1281]&m[1282])|(m[1222]&m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1222]&m[1278]&m[1279]&m[1281]&m[1282]))&UnbiasedRNG[488])|((m[1222]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(~m[1222]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1222]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1222]&m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1222]&~m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1222]&~m[1278]&~m[1279]&m[1281]&m[1282])|(m[1222]&~m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1222]&m[1278]&~m[1279]&m[1281]&m[1282])|(m[1222]&m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1222]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1222]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1222]&m[1278]&m[1279]&m[1281]&m[1282]))):InitCond[1187];
    m[1285] = run?((((m[1227]&~m[1283]&~m[1284]&~m[1286]&~m[1287])|(~m[1227]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1227]&m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1227]&~m[1283]&m[1284]&m[1286]&~m[1287])|(~m[1227]&m[1283]&~m[1284]&~m[1286]&m[1287])|(~m[1227]&~m[1283]&m[1284]&~m[1286]&m[1287])|(m[1227]&m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1227]&m[1283]&m[1284]&m[1286]&m[1287]))&UnbiasedRNG[489])|((m[1227]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(~m[1227]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1227]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1227]&m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1227]&~m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1227]&~m[1283]&~m[1284]&m[1286]&m[1287])|(m[1227]&~m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1227]&m[1283]&~m[1284]&m[1286]&m[1287])|(m[1227]&m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1227]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1227]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1227]&m[1283]&m[1284]&m[1286]&m[1287]))):InitCond[1188];
    m[1290] = run?((((m[1232]&~m[1288]&~m[1289]&~m[1291]&~m[1292])|(~m[1232]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1232]&m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1232]&~m[1288]&m[1289]&m[1291]&~m[1292])|(~m[1232]&m[1288]&~m[1289]&~m[1291]&m[1292])|(~m[1232]&~m[1288]&m[1289]&~m[1291]&m[1292])|(m[1232]&m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1232]&m[1288]&m[1289]&m[1291]&m[1292]))&UnbiasedRNG[490])|((m[1232]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(~m[1232]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1232]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1232]&m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1232]&~m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1232]&~m[1288]&~m[1289]&m[1291]&m[1292])|(m[1232]&~m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1232]&m[1288]&~m[1289]&m[1291]&m[1292])|(m[1232]&m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1232]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1232]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1232]&m[1288]&m[1289]&m[1291]&m[1292]))):InitCond[1189];
    m[1295] = run?((((m[1237]&~m[1293]&~m[1294]&~m[1296]&~m[1297])|(~m[1237]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1237]&m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1237]&~m[1293]&m[1294]&m[1296]&~m[1297])|(~m[1237]&m[1293]&~m[1294]&~m[1296]&m[1297])|(~m[1237]&~m[1293]&m[1294]&~m[1296]&m[1297])|(m[1237]&m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1237]&m[1293]&m[1294]&m[1296]&m[1297]))&UnbiasedRNG[491])|((m[1237]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(~m[1237]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1237]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1237]&m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1237]&~m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1237]&~m[1293]&~m[1294]&m[1296]&m[1297])|(m[1237]&~m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1237]&m[1293]&~m[1294]&m[1296]&m[1297])|(m[1237]&m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1237]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1237]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1237]&m[1293]&m[1294]&m[1296]&m[1297]))):InitCond[1190];
    m[1300] = run?((((m[1242]&~m[1298]&~m[1299]&~m[1301]&~m[1302])|(~m[1242]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1242]&m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1242]&~m[1298]&m[1299]&m[1301]&~m[1302])|(~m[1242]&m[1298]&~m[1299]&~m[1301]&m[1302])|(~m[1242]&~m[1298]&m[1299]&~m[1301]&m[1302])|(m[1242]&m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1242]&m[1298]&m[1299]&m[1301]&m[1302]))&UnbiasedRNG[492])|((m[1242]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(~m[1242]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1242]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1242]&m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1242]&~m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1242]&~m[1298]&~m[1299]&m[1301]&m[1302])|(m[1242]&~m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1242]&m[1298]&~m[1299]&m[1301]&m[1302])|(m[1242]&m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1242]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1242]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1242]&m[1298]&m[1299]&m[1301]&m[1302]))):InitCond[1191];
    m[1305] = run?((((m[1247]&~m[1303]&~m[1304]&~m[1306]&~m[1307])|(~m[1247]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1247]&m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1247]&~m[1303]&m[1304]&m[1306]&~m[1307])|(~m[1247]&m[1303]&~m[1304]&~m[1306]&m[1307])|(~m[1247]&~m[1303]&m[1304]&~m[1306]&m[1307])|(m[1247]&m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1247]&m[1303]&m[1304]&m[1306]&m[1307]))&UnbiasedRNG[493])|((m[1247]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(~m[1247]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1247]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1247]&m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1247]&~m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1247]&~m[1303]&~m[1304]&m[1306]&m[1307])|(m[1247]&~m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1247]&m[1303]&~m[1304]&m[1306]&m[1307])|(m[1247]&m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1247]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1247]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1247]&m[1303]&m[1304]&m[1306]&m[1307]))):InitCond[1192];
    m[1310] = run?((((m[1257]&~m[1308]&~m[1309]&~m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&~m[1312])|(~m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&m[1308]&m[1309]&m[1311]&m[1312]))&UnbiasedRNG[494])|((m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&m[1311]&m[1312]))):InitCond[1193];
    m[1315] = run?((((m[1262]&~m[1313]&~m[1314]&~m[1316]&~m[1317])|(~m[1262]&~m[1313]&~m[1314]&m[1316]&~m[1317])|(m[1262]&m[1313]&~m[1314]&m[1316]&~m[1317])|(m[1262]&~m[1313]&m[1314]&m[1316]&~m[1317])|(~m[1262]&m[1313]&~m[1314]&~m[1316]&m[1317])|(~m[1262]&~m[1313]&m[1314]&~m[1316]&m[1317])|(m[1262]&m[1313]&m[1314]&~m[1316]&m[1317])|(~m[1262]&m[1313]&m[1314]&m[1316]&m[1317]))&UnbiasedRNG[495])|((m[1262]&~m[1313]&~m[1314]&m[1316]&~m[1317])|(~m[1262]&~m[1313]&~m[1314]&~m[1316]&m[1317])|(m[1262]&~m[1313]&~m[1314]&~m[1316]&m[1317])|(m[1262]&m[1313]&~m[1314]&~m[1316]&m[1317])|(m[1262]&~m[1313]&m[1314]&~m[1316]&m[1317])|(~m[1262]&~m[1313]&~m[1314]&m[1316]&m[1317])|(m[1262]&~m[1313]&~m[1314]&m[1316]&m[1317])|(~m[1262]&m[1313]&~m[1314]&m[1316]&m[1317])|(m[1262]&m[1313]&~m[1314]&m[1316]&m[1317])|(~m[1262]&~m[1313]&m[1314]&m[1316]&m[1317])|(m[1262]&~m[1313]&m[1314]&m[1316]&m[1317])|(m[1262]&m[1313]&m[1314]&m[1316]&m[1317]))):InitCond[1194];
    m[1320] = run?((((m[1267]&~m[1318]&~m[1319]&~m[1321]&~m[1322])|(~m[1267]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1267]&m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1267]&~m[1318]&m[1319]&m[1321]&~m[1322])|(~m[1267]&m[1318]&~m[1319]&~m[1321]&m[1322])|(~m[1267]&~m[1318]&m[1319]&~m[1321]&m[1322])|(m[1267]&m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1267]&m[1318]&m[1319]&m[1321]&m[1322]))&UnbiasedRNG[496])|((m[1267]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(~m[1267]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1267]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1267]&m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1267]&~m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1267]&~m[1318]&~m[1319]&m[1321]&m[1322])|(m[1267]&~m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1267]&m[1318]&~m[1319]&m[1321]&m[1322])|(m[1267]&m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1267]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1267]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1267]&m[1318]&m[1319]&m[1321]&m[1322]))):InitCond[1195];
    m[1325] = run?((((m[1272]&~m[1323]&~m[1324]&~m[1326]&~m[1327])|(~m[1272]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1272]&m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1272]&~m[1323]&m[1324]&m[1326]&~m[1327])|(~m[1272]&m[1323]&~m[1324]&~m[1326]&m[1327])|(~m[1272]&~m[1323]&m[1324]&~m[1326]&m[1327])|(m[1272]&m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1272]&m[1323]&m[1324]&m[1326]&m[1327]))&UnbiasedRNG[497])|((m[1272]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(~m[1272]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1272]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1272]&m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1272]&~m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1272]&~m[1323]&~m[1324]&m[1326]&m[1327])|(m[1272]&~m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1272]&m[1323]&~m[1324]&m[1326]&m[1327])|(m[1272]&m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1272]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1272]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1272]&m[1323]&m[1324]&m[1326]&m[1327]))):InitCond[1196];
    m[1330] = run?((((m[1277]&~m[1328]&~m[1329]&~m[1331]&~m[1332])|(~m[1277]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1277]&m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1277]&~m[1328]&m[1329]&m[1331]&~m[1332])|(~m[1277]&m[1328]&~m[1329]&~m[1331]&m[1332])|(~m[1277]&~m[1328]&m[1329]&~m[1331]&m[1332])|(m[1277]&m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1277]&m[1328]&m[1329]&m[1331]&m[1332]))&UnbiasedRNG[498])|((m[1277]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(~m[1277]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1277]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1277]&m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1277]&~m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1277]&~m[1328]&~m[1329]&m[1331]&m[1332])|(m[1277]&~m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1277]&m[1328]&~m[1329]&m[1331]&m[1332])|(m[1277]&m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1277]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1277]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1277]&m[1328]&m[1329]&m[1331]&m[1332]))):InitCond[1197];
    m[1335] = run?((((m[1282]&~m[1333]&~m[1334]&~m[1336]&~m[1337])|(~m[1282]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1282]&m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1282]&~m[1333]&m[1334]&m[1336]&~m[1337])|(~m[1282]&m[1333]&~m[1334]&~m[1336]&m[1337])|(~m[1282]&~m[1333]&m[1334]&~m[1336]&m[1337])|(m[1282]&m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1282]&m[1333]&m[1334]&m[1336]&m[1337]))&UnbiasedRNG[499])|((m[1282]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(~m[1282]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1282]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1282]&m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1282]&~m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1282]&~m[1333]&~m[1334]&m[1336]&m[1337])|(m[1282]&~m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1282]&m[1333]&~m[1334]&m[1336]&m[1337])|(m[1282]&m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1282]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1282]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1282]&m[1333]&m[1334]&m[1336]&m[1337]))):InitCond[1198];
    m[1340] = run?((((m[1287]&~m[1338]&~m[1339]&~m[1341]&~m[1342])|(~m[1287]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1287]&m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1287]&~m[1338]&m[1339]&m[1341]&~m[1342])|(~m[1287]&m[1338]&~m[1339]&~m[1341]&m[1342])|(~m[1287]&~m[1338]&m[1339]&~m[1341]&m[1342])|(m[1287]&m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1287]&m[1338]&m[1339]&m[1341]&m[1342]))&UnbiasedRNG[500])|((m[1287]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(~m[1287]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1287]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1287]&m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1287]&~m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1287]&~m[1338]&~m[1339]&m[1341]&m[1342])|(m[1287]&~m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1287]&m[1338]&~m[1339]&m[1341]&m[1342])|(m[1287]&m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1287]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1287]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1287]&m[1338]&m[1339]&m[1341]&m[1342]))):InitCond[1199];
    m[1345] = run?((((m[1292]&~m[1343]&~m[1344]&~m[1346]&~m[1347])|(~m[1292]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1292]&m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1292]&~m[1343]&m[1344]&m[1346]&~m[1347])|(~m[1292]&m[1343]&~m[1344]&~m[1346]&m[1347])|(~m[1292]&~m[1343]&m[1344]&~m[1346]&m[1347])|(m[1292]&m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1292]&m[1343]&m[1344]&m[1346]&m[1347]))&UnbiasedRNG[501])|((m[1292]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(~m[1292]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1292]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1292]&m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1292]&~m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1292]&~m[1343]&~m[1344]&m[1346]&m[1347])|(m[1292]&~m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1292]&m[1343]&~m[1344]&m[1346]&m[1347])|(m[1292]&m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1292]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1292]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1292]&m[1343]&m[1344]&m[1346]&m[1347]))):InitCond[1200];
    m[1350] = run?((((m[1297]&~m[1348]&~m[1349]&~m[1351]&~m[1352])|(~m[1297]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1297]&m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1297]&~m[1348]&m[1349]&m[1351]&~m[1352])|(~m[1297]&m[1348]&~m[1349]&~m[1351]&m[1352])|(~m[1297]&~m[1348]&m[1349]&~m[1351]&m[1352])|(m[1297]&m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1297]&m[1348]&m[1349]&m[1351]&m[1352]))&UnbiasedRNG[502])|((m[1297]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(~m[1297]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1297]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1297]&m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1297]&~m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1297]&~m[1348]&~m[1349]&m[1351]&m[1352])|(m[1297]&~m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1297]&m[1348]&~m[1349]&m[1351]&m[1352])|(m[1297]&m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1297]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1297]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1297]&m[1348]&m[1349]&m[1351]&m[1352]))):InitCond[1201];
    m[1355] = run?((((m[1302]&~m[1353]&~m[1354]&~m[1356]&~m[1357])|(~m[1302]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1302]&m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1302]&~m[1353]&m[1354]&m[1356]&~m[1357])|(~m[1302]&m[1353]&~m[1354]&~m[1356]&m[1357])|(~m[1302]&~m[1353]&m[1354]&~m[1356]&m[1357])|(m[1302]&m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1302]&m[1353]&m[1354]&m[1356]&m[1357]))&UnbiasedRNG[503])|((m[1302]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(~m[1302]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1302]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1302]&m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1302]&~m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1302]&~m[1353]&~m[1354]&m[1356]&m[1357])|(m[1302]&~m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1302]&m[1353]&~m[1354]&m[1356]&m[1357])|(m[1302]&m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1302]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1302]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1302]&m[1353]&m[1354]&m[1356]&m[1357]))):InitCond[1202];
    m[1360] = run?((((m[1307]&~m[1358]&~m[1359]&~m[1361]&~m[1362])|(~m[1307]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1307]&m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1307]&~m[1358]&m[1359]&m[1361]&~m[1362])|(~m[1307]&m[1358]&~m[1359]&~m[1361]&m[1362])|(~m[1307]&~m[1358]&m[1359]&~m[1361]&m[1362])|(m[1307]&m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1307]&m[1358]&m[1359]&m[1361]&m[1362]))&UnbiasedRNG[504])|((m[1307]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(~m[1307]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1307]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1307]&m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1307]&~m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1307]&~m[1358]&~m[1359]&m[1361]&m[1362])|(m[1307]&~m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1307]&m[1358]&~m[1359]&m[1361]&m[1362])|(m[1307]&m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1307]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1307]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1307]&m[1358]&m[1359]&m[1361]&m[1362]))):InitCond[1203];
    m[1365] = run?((((m[1317]&~m[1363]&~m[1364]&~m[1366]&~m[1367])|(~m[1317]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1317]&m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1317]&~m[1363]&m[1364]&m[1366]&~m[1367])|(~m[1317]&m[1363]&~m[1364]&~m[1366]&m[1367])|(~m[1317]&~m[1363]&m[1364]&~m[1366]&m[1367])|(m[1317]&m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1317]&m[1363]&m[1364]&m[1366]&m[1367]))&UnbiasedRNG[505])|((m[1317]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(~m[1317]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1317]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1317]&m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1317]&~m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1317]&~m[1363]&~m[1364]&m[1366]&m[1367])|(m[1317]&~m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1317]&m[1363]&~m[1364]&m[1366]&m[1367])|(m[1317]&m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1317]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1317]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1317]&m[1363]&m[1364]&m[1366]&m[1367]))):InitCond[1204];
    m[1370] = run?((((m[1322]&~m[1368]&~m[1369]&~m[1371]&~m[1372])|(~m[1322]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1322]&m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1322]&~m[1368]&m[1369]&m[1371]&~m[1372])|(~m[1322]&m[1368]&~m[1369]&~m[1371]&m[1372])|(~m[1322]&~m[1368]&m[1369]&~m[1371]&m[1372])|(m[1322]&m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1322]&m[1368]&m[1369]&m[1371]&m[1372]))&UnbiasedRNG[506])|((m[1322]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(~m[1322]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1322]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1322]&m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1322]&~m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1322]&~m[1368]&~m[1369]&m[1371]&m[1372])|(m[1322]&~m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1322]&m[1368]&~m[1369]&m[1371]&m[1372])|(m[1322]&m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1322]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1322]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1322]&m[1368]&m[1369]&m[1371]&m[1372]))):InitCond[1205];
    m[1375] = run?((((m[1327]&~m[1373]&~m[1374]&~m[1376]&~m[1377])|(~m[1327]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1327]&m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1327]&~m[1373]&m[1374]&m[1376]&~m[1377])|(~m[1327]&m[1373]&~m[1374]&~m[1376]&m[1377])|(~m[1327]&~m[1373]&m[1374]&~m[1376]&m[1377])|(m[1327]&m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1327]&m[1373]&m[1374]&m[1376]&m[1377]))&UnbiasedRNG[507])|((m[1327]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(~m[1327]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1327]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1327]&m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1327]&~m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1327]&~m[1373]&~m[1374]&m[1376]&m[1377])|(m[1327]&~m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1327]&m[1373]&~m[1374]&m[1376]&m[1377])|(m[1327]&m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1327]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1327]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1327]&m[1373]&m[1374]&m[1376]&m[1377]))):InitCond[1206];
    m[1380] = run?((((m[1332]&~m[1378]&~m[1379]&~m[1381]&~m[1382])|(~m[1332]&~m[1378]&~m[1379]&m[1381]&~m[1382])|(m[1332]&m[1378]&~m[1379]&m[1381]&~m[1382])|(m[1332]&~m[1378]&m[1379]&m[1381]&~m[1382])|(~m[1332]&m[1378]&~m[1379]&~m[1381]&m[1382])|(~m[1332]&~m[1378]&m[1379]&~m[1381]&m[1382])|(m[1332]&m[1378]&m[1379]&~m[1381]&m[1382])|(~m[1332]&m[1378]&m[1379]&m[1381]&m[1382]))&UnbiasedRNG[508])|((m[1332]&~m[1378]&~m[1379]&m[1381]&~m[1382])|(~m[1332]&~m[1378]&~m[1379]&~m[1381]&m[1382])|(m[1332]&~m[1378]&~m[1379]&~m[1381]&m[1382])|(m[1332]&m[1378]&~m[1379]&~m[1381]&m[1382])|(m[1332]&~m[1378]&m[1379]&~m[1381]&m[1382])|(~m[1332]&~m[1378]&~m[1379]&m[1381]&m[1382])|(m[1332]&~m[1378]&~m[1379]&m[1381]&m[1382])|(~m[1332]&m[1378]&~m[1379]&m[1381]&m[1382])|(m[1332]&m[1378]&~m[1379]&m[1381]&m[1382])|(~m[1332]&~m[1378]&m[1379]&m[1381]&m[1382])|(m[1332]&~m[1378]&m[1379]&m[1381]&m[1382])|(m[1332]&m[1378]&m[1379]&m[1381]&m[1382]))):InitCond[1207];
    m[1385] = run?((((m[1337]&~m[1383]&~m[1384]&~m[1386]&~m[1387])|(~m[1337]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1337]&m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1337]&~m[1383]&m[1384]&m[1386]&~m[1387])|(~m[1337]&m[1383]&~m[1384]&~m[1386]&m[1387])|(~m[1337]&~m[1383]&m[1384]&~m[1386]&m[1387])|(m[1337]&m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1337]&m[1383]&m[1384]&m[1386]&m[1387]))&UnbiasedRNG[509])|((m[1337]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(~m[1337]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1337]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1337]&m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1337]&~m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1337]&~m[1383]&~m[1384]&m[1386]&m[1387])|(m[1337]&~m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1337]&m[1383]&~m[1384]&m[1386]&m[1387])|(m[1337]&m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1337]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1337]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1337]&m[1383]&m[1384]&m[1386]&m[1387]))):InitCond[1208];
    m[1390] = run?((((m[1342]&~m[1388]&~m[1389]&~m[1391]&~m[1392])|(~m[1342]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1342]&m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1342]&~m[1388]&m[1389]&m[1391]&~m[1392])|(~m[1342]&m[1388]&~m[1389]&~m[1391]&m[1392])|(~m[1342]&~m[1388]&m[1389]&~m[1391]&m[1392])|(m[1342]&m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1342]&m[1388]&m[1389]&m[1391]&m[1392]))&UnbiasedRNG[510])|((m[1342]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(~m[1342]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1342]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1342]&m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1342]&~m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1342]&~m[1388]&~m[1389]&m[1391]&m[1392])|(m[1342]&~m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1342]&m[1388]&~m[1389]&m[1391]&m[1392])|(m[1342]&m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1342]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1342]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1342]&m[1388]&m[1389]&m[1391]&m[1392]))):InitCond[1209];
    m[1395] = run?((((m[1347]&~m[1393]&~m[1394]&~m[1396]&~m[1397])|(~m[1347]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1347]&m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1347]&~m[1393]&m[1394]&m[1396]&~m[1397])|(~m[1347]&m[1393]&~m[1394]&~m[1396]&m[1397])|(~m[1347]&~m[1393]&m[1394]&~m[1396]&m[1397])|(m[1347]&m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1347]&m[1393]&m[1394]&m[1396]&m[1397]))&UnbiasedRNG[511])|((m[1347]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(~m[1347]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1347]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1347]&m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1347]&~m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1347]&~m[1393]&~m[1394]&m[1396]&m[1397])|(m[1347]&~m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1347]&m[1393]&~m[1394]&m[1396]&m[1397])|(m[1347]&m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1347]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1347]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1347]&m[1393]&m[1394]&m[1396]&m[1397]))):InitCond[1210];
    m[1400] = run?((((m[1352]&~m[1398]&~m[1399]&~m[1401]&~m[1402])|(~m[1352]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1352]&m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1352]&~m[1398]&m[1399]&m[1401]&~m[1402])|(~m[1352]&m[1398]&~m[1399]&~m[1401]&m[1402])|(~m[1352]&~m[1398]&m[1399]&~m[1401]&m[1402])|(m[1352]&m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1352]&m[1398]&m[1399]&m[1401]&m[1402]))&UnbiasedRNG[512])|((m[1352]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(~m[1352]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1352]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1352]&m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1352]&~m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1352]&~m[1398]&~m[1399]&m[1401]&m[1402])|(m[1352]&~m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1352]&m[1398]&~m[1399]&m[1401]&m[1402])|(m[1352]&m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1352]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1352]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1352]&m[1398]&m[1399]&m[1401]&m[1402]))):InitCond[1211];
    m[1405] = run?((((m[1357]&~m[1403]&~m[1404]&~m[1406]&~m[1407])|(~m[1357]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1357]&m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1357]&~m[1403]&m[1404]&m[1406]&~m[1407])|(~m[1357]&m[1403]&~m[1404]&~m[1406]&m[1407])|(~m[1357]&~m[1403]&m[1404]&~m[1406]&m[1407])|(m[1357]&m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1357]&m[1403]&m[1404]&m[1406]&m[1407]))&UnbiasedRNG[513])|((m[1357]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(~m[1357]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1357]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1357]&m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1357]&~m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1357]&~m[1403]&~m[1404]&m[1406]&m[1407])|(m[1357]&~m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1357]&m[1403]&~m[1404]&m[1406]&m[1407])|(m[1357]&m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1357]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1357]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1357]&m[1403]&m[1404]&m[1406]&m[1407]))):InitCond[1212];
    m[1410] = run?((((m[1362]&~m[1408]&~m[1409]&~m[1411]&~m[1412])|(~m[1362]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1362]&m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1362]&~m[1408]&m[1409]&m[1411]&~m[1412])|(~m[1362]&m[1408]&~m[1409]&~m[1411]&m[1412])|(~m[1362]&~m[1408]&m[1409]&~m[1411]&m[1412])|(m[1362]&m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1362]&m[1408]&m[1409]&m[1411]&m[1412]))&UnbiasedRNG[514])|((m[1362]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(~m[1362]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1362]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1362]&m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1362]&~m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1362]&~m[1408]&~m[1409]&m[1411]&m[1412])|(m[1362]&~m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1362]&m[1408]&~m[1409]&m[1411]&m[1412])|(m[1362]&m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1362]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1362]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1362]&m[1408]&m[1409]&m[1411]&m[1412]))):InitCond[1213];
    m[1415] = run?((((m[1372]&~m[1413]&~m[1414]&~m[1416]&~m[1417])|(~m[1372]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1372]&m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1372]&~m[1413]&m[1414]&m[1416]&~m[1417])|(~m[1372]&m[1413]&~m[1414]&~m[1416]&m[1417])|(~m[1372]&~m[1413]&m[1414]&~m[1416]&m[1417])|(m[1372]&m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1372]&m[1413]&m[1414]&m[1416]&m[1417]))&UnbiasedRNG[515])|((m[1372]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(~m[1372]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1372]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1372]&m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1372]&~m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1372]&~m[1413]&~m[1414]&m[1416]&m[1417])|(m[1372]&~m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1372]&m[1413]&~m[1414]&m[1416]&m[1417])|(m[1372]&m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1372]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1372]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1372]&m[1413]&m[1414]&m[1416]&m[1417]))):InitCond[1214];
    m[1420] = run?((((m[1377]&~m[1418]&~m[1419]&~m[1421]&~m[1422])|(~m[1377]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1377]&m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1377]&~m[1418]&m[1419]&m[1421]&~m[1422])|(~m[1377]&m[1418]&~m[1419]&~m[1421]&m[1422])|(~m[1377]&~m[1418]&m[1419]&~m[1421]&m[1422])|(m[1377]&m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1377]&m[1418]&m[1419]&m[1421]&m[1422]))&UnbiasedRNG[516])|((m[1377]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(~m[1377]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1377]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1377]&m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1377]&~m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1377]&~m[1418]&~m[1419]&m[1421]&m[1422])|(m[1377]&~m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1377]&m[1418]&~m[1419]&m[1421]&m[1422])|(m[1377]&m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1377]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1377]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1377]&m[1418]&m[1419]&m[1421]&m[1422]))):InitCond[1215];
    m[1425] = run?((((m[1382]&~m[1423]&~m[1424]&~m[1426]&~m[1427])|(~m[1382]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1382]&m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1382]&~m[1423]&m[1424]&m[1426]&~m[1427])|(~m[1382]&m[1423]&~m[1424]&~m[1426]&m[1427])|(~m[1382]&~m[1423]&m[1424]&~m[1426]&m[1427])|(m[1382]&m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1382]&m[1423]&m[1424]&m[1426]&m[1427]))&UnbiasedRNG[517])|((m[1382]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(~m[1382]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1382]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1382]&m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1382]&~m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1382]&~m[1423]&~m[1424]&m[1426]&m[1427])|(m[1382]&~m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1382]&m[1423]&~m[1424]&m[1426]&m[1427])|(m[1382]&m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1382]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1382]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1382]&m[1423]&m[1424]&m[1426]&m[1427]))):InitCond[1216];
    m[1430] = run?((((m[1387]&~m[1428]&~m[1429]&~m[1431]&~m[1432])|(~m[1387]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1387]&m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1387]&~m[1428]&m[1429]&m[1431]&~m[1432])|(~m[1387]&m[1428]&~m[1429]&~m[1431]&m[1432])|(~m[1387]&~m[1428]&m[1429]&~m[1431]&m[1432])|(m[1387]&m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1387]&m[1428]&m[1429]&m[1431]&m[1432]))&UnbiasedRNG[518])|((m[1387]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(~m[1387]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1387]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1387]&m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1387]&~m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1387]&~m[1428]&~m[1429]&m[1431]&m[1432])|(m[1387]&~m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1387]&m[1428]&~m[1429]&m[1431]&m[1432])|(m[1387]&m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1387]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1387]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1387]&m[1428]&m[1429]&m[1431]&m[1432]))):InitCond[1217];
    m[1435] = run?((((m[1392]&~m[1433]&~m[1434]&~m[1436]&~m[1437])|(~m[1392]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1392]&m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1392]&~m[1433]&m[1434]&m[1436]&~m[1437])|(~m[1392]&m[1433]&~m[1434]&~m[1436]&m[1437])|(~m[1392]&~m[1433]&m[1434]&~m[1436]&m[1437])|(m[1392]&m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1392]&m[1433]&m[1434]&m[1436]&m[1437]))&UnbiasedRNG[519])|((m[1392]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(~m[1392]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1392]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1392]&m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1392]&~m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1392]&~m[1433]&~m[1434]&m[1436]&m[1437])|(m[1392]&~m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1392]&m[1433]&~m[1434]&m[1436]&m[1437])|(m[1392]&m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1392]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1392]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1392]&m[1433]&m[1434]&m[1436]&m[1437]))):InitCond[1218];
    m[1440] = run?((((m[1397]&~m[1438]&~m[1439]&~m[1441]&~m[1442])|(~m[1397]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1397]&m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1397]&~m[1438]&m[1439]&m[1441]&~m[1442])|(~m[1397]&m[1438]&~m[1439]&~m[1441]&m[1442])|(~m[1397]&~m[1438]&m[1439]&~m[1441]&m[1442])|(m[1397]&m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1397]&m[1438]&m[1439]&m[1441]&m[1442]))&UnbiasedRNG[520])|((m[1397]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(~m[1397]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1397]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1397]&m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1397]&~m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1397]&~m[1438]&~m[1439]&m[1441]&m[1442])|(m[1397]&~m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1397]&m[1438]&~m[1439]&m[1441]&m[1442])|(m[1397]&m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1397]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1397]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1397]&m[1438]&m[1439]&m[1441]&m[1442]))):InitCond[1219];
    m[1445] = run?((((m[1402]&~m[1443]&~m[1444]&~m[1446]&~m[1447])|(~m[1402]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1402]&m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1402]&~m[1443]&m[1444]&m[1446]&~m[1447])|(~m[1402]&m[1443]&~m[1444]&~m[1446]&m[1447])|(~m[1402]&~m[1443]&m[1444]&~m[1446]&m[1447])|(m[1402]&m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1402]&m[1443]&m[1444]&m[1446]&m[1447]))&UnbiasedRNG[521])|((m[1402]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(~m[1402]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1402]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1402]&m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1402]&~m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1402]&~m[1443]&~m[1444]&m[1446]&m[1447])|(m[1402]&~m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1402]&m[1443]&~m[1444]&m[1446]&m[1447])|(m[1402]&m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1402]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1402]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1402]&m[1443]&m[1444]&m[1446]&m[1447]))):InitCond[1220];
    m[1450] = run?((((m[1407]&~m[1448]&~m[1449]&~m[1451]&~m[1452])|(~m[1407]&~m[1448]&~m[1449]&m[1451]&~m[1452])|(m[1407]&m[1448]&~m[1449]&m[1451]&~m[1452])|(m[1407]&~m[1448]&m[1449]&m[1451]&~m[1452])|(~m[1407]&m[1448]&~m[1449]&~m[1451]&m[1452])|(~m[1407]&~m[1448]&m[1449]&~m[1451]&m[1452])|(m[1407]&m[1448]&m[1449]&~m[1451]&m[1452])|(~m[1407]&m[1448]&m[1449]&m[1451]&m[1452]))&UnbiasedRNG[522])|((m[1407]&~m[1448]&~m[1449]&m[1451]&~m[1452])|(~m[1407]&~m[1448]&~m[1449]&~m[1451]&m[1452])|(m[1407]&~m[1448]&~m[1449]&~m[1451]&m[1452])|(m[1407]&m[1448]&~m[1449]&~m[1451]&m[1452])|(m[1407]&~m[1448]&m[1449]&~m[1451]&m[1452])|(~m[1407]&~m[1448]&~m[1449]&m[1451]&m[1452])|(m[1407]&~m[1448]&~m[1449]&m[1451]&m[1452])|(~m[1407]&m[1448]&~m[1449]&m[1451]&m[1452])|(m[1407]&m[1448]&~m[1449]&m[1451]&m[1452])|(~m[1407]&~m[1448]&m[1449]&m[1451]&m[1452])|(m[1407]&~m[1448]&m[1449]&m[1451]&m[1452])|(m[1407]&m[1448]&m[1449]&m[1451]&m[1452]))):InitCond[1221];
    m[1455] = run?((((m[1412]&~m[1453]&~m[1454]&~m[1456]&~m[1457])|(~m[1412]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1412]&m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1412]&~m[1453]&m[1454]&m[1456]&~m[1457])|(~m[1412]&m[1453]&~m[1454]&~m[1456]&m[1457])|(~m[1412]&~m[1453]&m[1454]&~m[1456]&m[1457])|(m[1412]&m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1412]&m[1453]&m[1454]&m[1456]&m[1457]))&UnbiasedRNG[523])|((m[1412]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(~m[1412]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1412]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1412]&m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1412]&~m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1412]&~m[1453]&~m[1454]&m[1456]&m[1457])|(m[1412]&~m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1412]&m[1453]&~m[1454]&m[1456]&m[1457])|(m[1412]&m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1412]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1412]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1412]&m[1453]&m[1454]&m[1456]&m[1457]))):InitCond[1222];
    m[1460] = run?((((m[1422]&~m[1458]&~m[1459]&~m[1461]&~m[1462])|(~m[1422]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1422]&m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1422]&~m[1458]&m[1459]&m[1461]&~m[1462])|(~m[1422]&m[1458]&~m[1459]&~m[1461]&m[1462])|(~m[1422]&~m[1458]&m[1459]&~m[1461]&m[1462])|(m[1422]&m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1422]&m[1458]&m[1459]&m[1461]&m[1462]))&UnbiasedRNG[524])|((m[1422]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(~m[1422]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1422]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1422]&m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1422]&~m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1422]&~m[1458]&~m[1459]&m[1461]&m[1462])|(m[1422]&~m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1422]&m[1458]&~m[1459]&m[1461]&m[1462])|(m[1422]&m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1422]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1422]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1422]&m[1458]&m[1459]&m[1461]&m[1462]))):InitCond[1223];
    m[1465] = run?((((m[1427]&~m[1463]&~m[1464]&~m[1466]&~m[1467])|(~m[1427]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1427]&m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1427]&~m[1463]&m[1464]&m[1466]&~m[1467])|(~m[1427]&m[1463]&~m[1464]&~m[1466]&m[1467])|(~m[1427]&~m[1463]&m[1464]&~m[1466]&m[1467])|(m[1427]&m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1427]&m[1463]&m[1464]&m[1466]&m[1467]))&UnbiasedRNG[525])|((m[1427]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(~m[1427]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1427]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1427]&m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1427]&~m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1427]&~m[1463]&~m[1464]&m[1466]&m[1467])|(m[1427]&~m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1427]&m[1463]&~m[1464]&m[1466]&m[1467])|(m[1427]&m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1427]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1427]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1427]&m[1463]&m[1464]&m[1466]&m[1467]))):InitCond[1224];
    m[1470] = run?((((m[1432]&~m[1468]&~m[1469]&~m[1471]&~m[1472])|(~m[1432]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1432]&m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1432]&~m[1468]&m[1469]&m[1471]&~m[1472])|(~m[1432]&m[1468]&~m[1469]&~m[1471]&m[1472])|(~m[1432]&~m[1468]&m[1469]&~m[1471]&m[1472])|(m[1432]&m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1432]&m[1468]&m[1469]&m[1471]&m[1472]))&UnbiasedRNG[526])|((m[1432]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(~m[1432]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1432]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1432]&m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1432]&~m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1432]&~m[1468]&~m[1469]&m[1471]&m[1472])|(m[1432]&~m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1432]&m[1468]&~m[1469]&m[1471]&m[1472])|(m[1432]&m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1432]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1432]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1432]&m[1468]&m[1469]&m[1471]&m[1472]))):InitCond[1225];
    m[1475] = run?((((m[1437]&~m[1473]&~m[1474]&~m[1476]&~m[1477])|(~m[1437]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1437]&m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1437]&~m[1473]&m[1474]&m[1476]&~m[1477])|(~m[1437]&m[1473]&~m[1474]&~m[1476]&m[1477])|(~m[1437]&~m[1473]&m[1474]&~m[1476]&m[1477])|(m[1437]&m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1437]&m[1473]&m[1474]&m[1476]&m[1477]))&UnbiasedRNG[527])|((m[1437]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(~m[1437]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1437]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1437]&m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1437]&~m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1437]&~m[1473]&~m[1474]&m[1476]&m[1477])|(m[1437]&~m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1437]&m[1473]&~m[1474]&m[1476]&m[1477])|(m[1437]&m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1437]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1437]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1437]&m[1473]&m[1474]&m[1476]&m[1477]))):InitCond[1226];
    m[1480] = run?((((m[1442]&~m[1478]&~m[1479]&~m[1481]&~m[1482])|(~m[1442]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1442]&m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1442]&~m[1478]&m[1479]&m[1481]&~m[1482])|(~m[1442]&m[1478]&~m[1479]&~m[1481]&m[1482])|(~m[1442]&~m[1478]&m[1479]&~m[1481]&m[1482])|(m[1442]&m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1442]&m[1478]&m[1479]&m[1481]&m[1482]))&UnbiasedRNG[528])|((m[1442]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(~m[1442]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1442]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1442]&m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1442]&~m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1442]&~m[1478]&~m[1479]&m[1481]&m[1482])|(m[1442]&~m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1442]&m[1478]&~m[1479]&m[1481]&m[1482])|(m[1442]&m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1442]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1442]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1442]&m[1478]&m[1479]&m[1481]&m[1482]))):InitCond[1227];
    m[1485] = run?((((m[1447]&~m[1483]&~m[1484]&~m[1486]&~m[1487])|(~m[1447]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1447]&m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1447]&~m[1483]&m[1484]&m[1486]&~m[1487])|(~m[1447]&m[1483]&~m[1484]&~m[1486]&m[1487])|(~m[1447]&~m[1483]&m[1484]&~m[1486]&m[1487])|(m[1447]&m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1447]&m[1483]&m[1484]&m[1486]&m[1487]))&UnbiasedRNG[529])|((m[1447]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(~m[1447]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1447]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1447]&m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1447]&~m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1447]&~m[1483]&~m[1484]&m[1486]&m[1487])|(m[1447]&~m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1447]&m[1483]&~m[1484]&m[1486]&m[1487])|(m[1447]&m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1447]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1447]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1447]&m[1483]&m[1484]&m[1486]&m[1487]))):InitCond[1228];
    m[1490] = run?((((m[1452]&~m[1488]&~m[1489]&~m[1491]&~m[1492])|(~m[1452]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1452]&m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1452]&~m[1488]&m[1489]&m[1491]&~m[1492])|(~m[1452]&m[1488]&~m[1489]&~m[1491]&m[1492])|(~m[1452]&~m[1488]&m[1489]&~m[1491]&m[1492])|(m[1452]&m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1452]&m[1488]&m[1489]&m[1491]&m[1492]))&UnbiasedRNG[530])|((m[1452]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(~m[1452]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1452]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1452]&m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1452]&~m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1452]&~m[1488]&~m[1489]&m[1491]&m[1492])|(m[1452]&~m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1452]&m[1488]&~m[1489]&m[1491]&m[1492])|(m[1452]&m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1452]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1452]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1452]&m[1488]&m[1489]&m[1491]&m[1492]))):InitCond[1229];
    m[1495] = run?((((m[1457]&~m[1493]&~m[1494]&~m[1496]&~m[1497])|(~m[1457]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1457]&m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1457]&~m[1493]&m[1494]&m[1496]&~m[1497])|(~m[1457]&m[1493]&~m[1494]&~m[1496]&m[1497])|(~m[1457]&~m[1493]&m[1494]&~m[1496]&m[1497])|(m[1457]&m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1457]&m[1493]&m[1494]&m[1496]&m[1497]))&UnbiasedRNG[531])|((m[1457]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(~m[1457]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1457]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1457]&m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1457]&~m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1457]&~m[1493]&~m[1494]&m[1496]&m[1497])|(m[1457]&~m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1457]&m[1493]&~m[1494]&m[1496]&m[1497])|(m[1457]&m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1457]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1457]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1457]&m[1493]&m[1494]&m[1496]&m[1497]))):InitCond[1230];
    m[1500] = run?((((m[1467]&~m[1498]&~m[1499]&~m[1501]&~m[1502])|(~m[1467]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1467]&m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1467]&~m[1498]&m[1499]&m[1501]&~m[1502])|(~m[1467]&m[1498]&~m[1499]&~m[1501]&m[1502])|(~m[1467]&~m[1498]&m[1499]&~m[1501]&m[1502])|(m[1467]&m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1467]&m[1498]&m[1499]&m[1501]&m[1502]))&UnbiasedRNG[532])|((m[1467]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(~m[1467]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1467]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1467]&m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1467]&~m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1467]&~m[1498]&~m[1499]&m[1501]&m[1502])|(m[1467]&~m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1467]&m[1498]&~m[1499]&m[1501]&m[1502])|(m[1467]&m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1467]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1467]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1467]&m[1498]&m[1499]&m[1501]&m[1502]))):InitCond[1231];
    m[1505] = run?((((m[1472]&~m[1503]&~m[1504]&~m[1506]&~m[1507])|(~m[1472]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1472]&m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1472]&~m[1503]&m[1504]&m[1506]&~m[1507])|(~m[1472]&m[1503]&~m[1504]&~m[1506]&m[1507])|(~m[1472]&~m[1503]&m[1504]&~m[1506]&m[1507])|(m[1472]&m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1472]&m[1503]&m[1504]&m[1506]&m[1507]))&UnbiasedRNG[533])|((m[1472]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(~m[1472]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1472]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1472]&m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1472]&~m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1472]&~m[1503]&~m[1504]&m[1506]&m[1507])|(m[1472]&~m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1472]&m[1503]&~m[1504]&m[1506]&m[1507])|(m[1472]&m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1472]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1472]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1472]&m[1503]&m[1504]&m[1506]&m[1507]))):InitCond[1232];
    m[1510] = run?((((m[1477]&~m[1508]&~m[1509]&~m[1511]&~m[1512])|(~m[1477]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1477]&m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1477]&~m[1508]&m[1509]&m[1511]&~m[1512])|(~m[1477]&m[1508]&~m[1509]&~m[1511]&m[1512])|(~m[1477]&~m[1508]&m[1509]&~m[1511]&m[1512])|(m[1477]&m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1477]&m[1508]&m[1509]&m[1511]&m[1512]))&UnbiasedRNG[534])|((m[1477]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(~m[1477]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1477]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1477]&m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1477]&~m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1477]&~m[1508]&~m[1509]&m[1511]&m[1512])|(m[1477]&~m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1477]&m[1508]&~m[1509]&m[1511]&m[1512])|(m[1477]&m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1477]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1477]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1477]&m[1508]&m[1509]&m[1511]&m[1512]))):InitCond[1233];
    m[1515] = run?((((m[1482]&~m[1513]&~m[1514]&~m[1516]&~m[1517])|(~m[1482]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1482]&m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1482]&~m[1513]&m[1514]&m[1516]&~m[1517])|(~m[1482]&m[1513]&~m[1514]&~m[1516]&m[1517])|(~m[1482]&~m[1513]&m[1514]&~m[1516]&m[1517])|(m[1482]&m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1482]&m[1513]&m[1514]&m[1516]&m[1517]))&UnbiasedRNG[535])|((m[1482]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(~m[1482]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1482]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1482]&m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1482]&~m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1482]&~m[1513]&~m[1514]&m[1516]&m[1517])|(m[1482]&~m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1482]&m[1513]&~m[1514]&m[1516]&m[1517])|(m[1482]&m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1482]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1482]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1482]&m[1513]&m[1514]&m[1516]&m[1517]))):InitCond[1234];
    m[1520] = run?((((m[1487]&~m[1518]&~m[1519]&~m[1521]&~m[1522])|(~m[1487]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1487]&m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1487]&~m[1518]&m[1519]&m[1521]&~m[1522])|(~m[1487]&m[1518]&~m[1519]&~m[1521]&m[1522])|(~m[1487]&~m[1518]&m[1519]&~m[1521]&m[1522])|(m[1487]&m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1487]&m[1518]&m[1519]&m[1521]&m[1522]))&UnbiasedRNG[536])|((m[1487]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(~m[1487]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1487]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1487]&m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1487]&~m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1487]&~m[1518]&~m[1519]&m[1521]&m[1522])|(m[1487]&~m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1487]&m[1518]&~m[1519]&m[1521]&m[1522])|(m[1487]&m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1487]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1487]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1487]&m[1518]&m[1519]&m[1521]&m[1522]))):InitCond[1235];
    m[1525] = run?((((m[1492]&~m[1523]&~m[1524]&~m[1526]&~m[1527])|(~m[1492]&~m[1523]&~m[1524]&m[1526]&~m[1527])|(m[1492]&m[1523]&~m[1524]&m[1526]&~m[1527])|(m[1492]&~m[1523]&m[1524]&m[1526]&~m[1527])|(~m[1492]&m[1523]&~m[1524]&~m[1526]&m[1527])|(~m[1492]&~m[1523]&m[1524]&~m[1526]&m[1527])|(m[1492]&m[1523]&m[1524]&~m[1526]&m[1527])|(~m[1492]&m[1523]&m[1524]&m[1526]&m[1527]))&UnbiasedRNG[537])|((m[1492]&~m[1523]&~m[1524]&m[1526]&~m[1527])|(~m[1492]&~m[1523]&~m[1524]&~m[1526]&m[1527])|(m[1492]&~m[1523]&~m[1524]&~m[1526]&m[1527])|(m[1492]&m[1523]&~m[1524]&~m[1526]&m[1527])|(m[1492]&~m[1523]&m[1524]&~m[1526]&m[1527])|(~m[1492]&~m[1523]&~m[1524]&m[1526]&m[1527])|(m[1492]&~m[1523]&~m[1524]&m[1526]&m[1527])|(~m[1492]&m[1523]&~m[1524]&m[1526]&m[1527])|(m[1492]&m[1523]&~m[1524]&m[1526]&m[1527])|(~m[1492]&~m[1523]&m[1524]&m[1526]&m[1527])|(m[1492]&~m[1523]&m[1524]&m[1526]&m[1527])|(m[1492]&m[1523]&m[1524]&m[1526]&m[1527]))):InitCond[1236];
    m[1530] = run?((((m[1497]&~m[1528]&~m[1529]&~m[1531]&~m[1532])|(~m[1497]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1497]&m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1497]&~m[1528]&m[1529]&m[1531]&~m[1532])|(~m[1497]&m[1528]&~m[1529]&~m[1531]&m[1532])|(~m[1497]&~m[1528]&m[1529]&~m[1531]&m[1532])|(m[1497]&m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1497]&m[1528]&m[1529]&m[1531]&m[1532]))&UnbiasedRNG[538])|((m[1497]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(~m[1497]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1497]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1497]&m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1497]&~m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1497]&~m[1528]&~m[1529]&m[1531]&m[1532])|(m[1497]&~m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1497]&m[1528]&~m[1529]&m[1531]&m[1532])|(m[1497]&m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1497]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1497]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1497]&m[1528]&m[1529]&m[1531]&m[1532]))):InitCond[1237];
    m[1535] = run?((((m[1507]&~m[1533]&~m[1534]&~m[1536]&~m[1537])|(~m[1507]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1507]&m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1507]&~m[1533]&m[1534]&m[1536]&~m[1537])|(~m[1507]&m[1533]&~m[1534]&~m[1536]&m[1537])|(~m[1507]&~m[1533]&m[1534]&~m[1536]&m[1537])|(m[1507]&m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1507]&m[1533]&m[1534]&m[1536]&m[1537]))&UnbiasedRNG[539])|((m[1507]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(~m[1507]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1507]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1507]&m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1507]&~m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1507]&~m[1533]&~m[1534]&m[1536]&m[1537])|(m[1507]&~m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1507]&m[1533]&~m[1534]&m[1536]&m[1537])|(m[1507]&m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1507]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1507]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1507]&m[1533]&m[1534]&m[1536]&m[1537]))):InitCond[1238];
    m[1540] = run?((((m[1512]&~m[1538]&~m[1539]&~m[1541]&~m[1542])|(~m[1512]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1512]&m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1512]&~m[1538]&m[1539]&m[1541]&~m[1542])|(~m[1512]&m[1538]&~m[1539]&~m[1541]&m[1542])|(~m[1512]&~m[1538]&m[1539]&~m[1541]&m[1542])|(m[1512]&m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1512]&m[1538]&m[1539]&m[1541]&m[1542]))&UnbiasedRNG[540])|((m[1512]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(~m[1512]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1512]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1512]&m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1512]&~m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1512]&~m[1538]&~m[1539]&m[1541]&m[1542])|(m[1512]&~m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1512]&m[1538]&~m[1539]&m[1541]&m[1542])|(m[1512]&m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1512]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1512]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1512]&m[1538]&m[1539]&m[1541]&m[1542]))):InitCond[1239];
    m[1545] = run?((((m[1517]&~m[1543]&~m[1544]&~m[1546]&~m[1547])|(~m[1517]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1517]&m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1517]&~m[1543]&m[1544]&m[1546]&~m[1547])|(~m[1517]&m[1543]&~m[1544]&~m[1546]&m[1547])|(~m[1517]&~m[1543]&m[1544]&~m[1546]&m[1547])|(m[1517]&m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1517]&m[1543]&m[1544]&m[1546]&m[1547]))&UnbiasedRNG[541])|((m[1517]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(~m[1517]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1517]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1517]&m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1517]&~m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1517]&~m[1543]&~m[1544]&m[1546]&m[1547])|(m[1517]&~m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1517]&m[1543]&~m[1544]&m[1546]&m[1547])|(m[1517]&m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1517]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1517]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1517]&m[1543]&m[1544]&m[1546]&m[1547]))):InitCond[1240];
    m[1550] = run?((((m[1522]&~m[1548]&~m[1549]&~m[1551]&~m[1552])|(~m[1522]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1522]&m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1522]&~m[1548]&m[1549]&m[1551]&~m[1552])|(~m[1522]&m[1548]&~m[1549]&~m[1551]&m[1552])|(~m[1522]&~m[1548]&m[1549]&~m[1551]&m[1552])|(m[1522]&m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1522]&m[1548]&m[1549]&m[1551]&m[1552]))&UnbiasedRNG[542])|((m[1522]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(~m[1522]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1522]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1522]&m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1522]&~m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1522]&~m[1548]&~m[1549]&m[1551]&m[1552])|(m[1522]&~m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1522]&m[1548]&~m[1549]&m[1551]&m[1552])|(m[1522]&m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1522]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1522]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1522]&m[1548]&m[1549]&m[1551]&m[1552]))):InitCond[1241];
    m[1555] = run?((((m[1527]&~m[1553]&~m[1554]&~m[1556]&~m[1557])|(~m[1527]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1527]&m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1527]&~m[1553]&m[1554]&m[1556]&~m[1557])|(~m[1527]&m[1553]&~m[1554]&~m[1556]&m[1557])|(~m[1527]&~m[1553]&m[1554]&~m[1556]&m[1557])|(m[1527]&m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1527]&m[1553]&m[1554]&m[1556]&m[1557]))&UnbiasedRNG[543])|((m[1527]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(~m[1527]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1527]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1527]&m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1527]&~m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1527]&~m[1553]&~m[1554]&m[1556]&m[1557])|(m[1527]&~m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1527]&m[1553]&~m[1554]&m[1556]&m[1557])|(m[1527]&m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1527]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1527]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1527]&m[1553]&m[1554]&m[1556]&m[1557]))):InitCond[1242];
    m[1560] = run?((((m[1532]&~m[1558]&~m[1559]&~m[1561]&~m[1562])|(~m[1532]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1532]&m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1532]&~m[1558]&m[1559]&m[1561]&~m[1562])|(~m[1532]&m[1558]&~m[1559]&~m[1561]&m[1562])|(~m[1532]&~m[1558]&m[1559]&~m[1561]&m[1562])|(m[1532]&m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1532]&m[1558]&m[1559]&m[1561]&m[1562]))&UnbiasedRNG[544])|((m[1532]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(~m[1532]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1532]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1532]&m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1532]&~m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1532]&~m[1558]&~m[1559]&m[1561]&m[1562])|(m[1532]&~m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1532]&m[1558]&~m[1559]&m[1561]&m[1562])|(m[1532]&m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1532]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1532]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1532]&m[1558]&m[1559]&m[1561]&m[1562]))):InitCond[1243];
    m[1565] = run?((((m[1542]&~m[1563]&~m[1564]&~m[1566]&~m[1567])|(~m[1542]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1542]&m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1542]&~m[1563]&m[1564]&m[1566]&~m[1567])|(~m[1542]&m[1563]&~m[1564]&~m[1566]&m[1567])|(~m[1542]&~m[1563]&m[1564]&~m[1566]&m[1567])|(m[1542]&m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1542]&m[1563]&m[1564]&m[1566]&m[1567]))&UnbiasedRNG[545])|((m[1542]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(~m[1542]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1542]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1542]&m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1542]&~m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1542]&~m[1563]&~m[1564]&m[1566]&m[1567])|(m[1542]&~m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1542]&m[1563]&~m[1564]&m[1566]&m[1567])|(m[1542]&m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1542]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1542]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1542]&m[1563]&m[1564]&m[1566]&m[1567]))):InitCond[1244];
    m[1570] = run?((((m[1547]&~m[1568]&~m[1569]&~m[1571]&~m[1572])|(~m[1547]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1547]&m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1547]&~m[1568]&m[1569]&m[1571]&~m[1572])|(~m[1547]&m[1568]&~m[1569]&~m[1571]&m[1572])|(~m[1547]&~m[1568]&m[1569]&~m[1571]&m[1572])|(m[1547]&m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1547]&m[1568]&m[1569]&m[1571]&m[1572]))&UnbiasedRNG[546])|((m[1547]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(~m[1547]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1547]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1547]&m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1547]&~m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1547]&~m[1568]&~m[1569]&m[1571]&m[1572])|(m[1547]&~m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1547]&m[1568]&~m[1569]&m[1571]&m[1572])|(m[1547]&m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1547]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1547]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1547]&m[1568]&m[1569]&m[1571]&m[1572]))):InitCond[1245];
    m[1575] = run?((((m[1552]&~m[1573]&~m[1574]&~m[1576]&~m[1577])|(~m[1552]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1552]&m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1552]&~m[1573]&m[1574]&m[1576]&~m[1577])|(~m[1552]&m[1573]&~m[1574]&~m[1576]&m[1577])|(~m[1552]&~m[1573]&m[1574]&~m[1576]&m[1577])|(m[1552]&m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1552]&m[1573]&m[1574]&m[1576]&m[1577]))&UnbiasedRNG[547])|((m[1552]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(~m[1552]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1552]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1552]&m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1552]&~m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1552]&~m[1573]&~m[1574]&m[1576]&m[1577])|(m[1552]&~m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1552]&m[1573]&~m[1574]&m[1576]&m[1577])|(m[1552]&m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1552]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1552]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1552]&m[1573]&m[1574]&m[1576]&m[1577]))):InitCond[1246];
    m[1580] = run?((((m[1557]&~m[1578]&~m[1579]&~m[1581]&~m[1582])|(~m[1557]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1557]&m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1557]&~m[1578]&m[1579]&m[1581]&~m[1582])|(~m[1557]&m[1578]&~m[1579]&~m[1581]&m[1582])|(~m[1557]&~m[1578]&m[1579]&~m[1581]&m[1582])|(m[1557]&m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1557]&m[1578]&m[1579]&m[1581]&m[1582]))&UnbiasedRNG[548])|((m[1557]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(~m[1557]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1557]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1557]&m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1557]&~m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1557]&~m[1578]&~m[1579]&m[1581]&m[1582])|(m[1557]&~m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1557]&m[1578]&~m[1579]&m[1581]&m[1582])|(m[1557]&m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1557]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1557]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1557]&m[1578]&m[1579]&m[1581]&m[1582]))):InitCond[1247];
    m[1585] = run?((((m[1562]&~m[1583]&~m[1584]&~m[1586]&~m[1587])|(~m[1562]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1562]&m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1562]&~m[1583]&m[1584]&m[1586]&~m[1587])|(~m[1562]&m[1583]&~m[1584]&~m[1586]&m[1587])|(~m[1562]&~m[1583]&m[1584]&~m[1586]&m[1587])|(m[1562]&m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1562]&m[1583]&m[1584]&m[1586]&m[1587]))&UnbiasedRNG[549])|((m[1562]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(~m[1562]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1562]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1562]&m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1562]&~m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1562]&~m[1583]&~m[1584]&m[1586]&m[1587])|(m[1562]&~m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1562]&m[1583]&~m[1584]&m[1586]&m[1587])|(m[1562]&m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1562]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1562]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1562]&m[1583]&m[1584]&m[1586]&m[1587]))):InitCond[1248];
    m[1590] = run?((((m[1572]&~m[1588]&~m[1589]&~m[1591]&~m[1592])|(~m[1572]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1572]&m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1572]&~m[1588]&m[1589]&m[1591]&~m[1592])|(~m[1572]&m[1588]&~m[1589]&~m[1591]&m[1592])|(~m[1572]&~m[1588]&m[1589]&~m[1591]&m[1592])|(m[1572]&m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1572]&m[1588]&m[1589]&m[1591]&m[1592]))&UnbiasedRNG[550])|((m[1572]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(~m[1572]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1572]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1572]&m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1572]&~m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1572]&~m[1588]&~m[1589]&m[1591]&m[1592])|(m[1572]&~m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1572]&m[1588]&~m[1589]&m[1591]&m[1592])|(m[1572]&m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1572]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1572]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1572]&m[1588]&m[1589]&m[1591]&m[1592]))):InitCond[1249];
    m[1595] = run?((((m[1577]&~m[1593]&~m[1594]&~m[1596]&~m[1597])|(~m[1577]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1577]&m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1577]&~m[1593]&m[1594]&m[1596]&~m[1597])|(~m[1577]&m[1593]&~m[1594]&~m[1596]&m[1597])|(~m[1577]&~m[1593]&m[1594]&~m[1596]&m[1597])|(m[1577]&m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1577]&m[1593]&m[1594]&m[1596]&m[1597]))&UnbiasedRNG[551])|((m[1577]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(~m[1577]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1577]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1577]&m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1577]&~m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1577]&~m[1593]&~m[1594]&m[1596]&m[1597])|(m[1577]&~m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1577]&m[1593]&~m[1594]&m[1596]&m[1597])|(m[1577]&m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1577]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1577]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1577]&m[1593]&m[1594]&m[1596]&m[1597]))):InitCond[1250];
    m[1600] = run?((((m[1582]&~m[1598]&~m[1599]&~m[1601]&~m[1602])|(~m[1582]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1582]&m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1582]&~m[1598]&m[1599]&m[1601]&~m[1602])|(~m[1582]&m[1598]&~m[1599]&~m[1601]&m[1602])|(~m[1582]&~m[1598]&m[1599]&~m[1601]&m[1602])|(m[1582]&m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1582]&m[1598]&m[1599]&m[1601]&m[1602]))&UnbiasedRNG[552])|((m[1582]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(~m[1582]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1582]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1582]&m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1582]&~m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1582]&~m[1598]&~m[1599]&m[1601]&m[1602])|(m[1582]&~m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1582]&m[1598]&~m[1599]&m[1601]&m[1602])|(m[1582]&m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1582]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1582]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1582]&m[1598]&m[1599]&m[1601]&m[1602]))):InitCond[1251];
    m[1605] = run?((((m[1587]&~m[1603]&~m[1604]&~m[1606]&~m[1607])|(~m[1587]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1587]&m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1587]&~m[1603]&m[1604]&m[1606]&~m[1607])|(~m[1587]&m[1603]&~m[1604]&~m[1606]&m[1607])|(~m[1587]&~m[1603]&m[1604]&~m[1606]&m[1607])|(m[1587]&m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1587]&m[1603]&m[1604]&m[1606]&m[1607]))&UnbiasedRNG[553])|((m[1587]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(~m[1587]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1587]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1587]&m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1587]&~m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1587]&~m[1603]&~m[1604]&m[1606]&m[1607])|(m[1587]&~m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1587]&m[1603]&~m[1604]&m[1606]&m[1607])|(m[1587]&m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1587]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1587]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1587]&m[1603]&m[1604]&m[1606]&m[1607]))):InitCond[1252];
    m[1610] = run?((((m[1597]&~m[1608]&~m[1609]&~m[1611]&~m[1612])|(~m[1597]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1597]&m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1597]&~m[1608]&m[1609]&m[1611]&~m[1612])|(~m[1597]&m[1608]&~m[1609]&~m[1611]&m[1612])|(~m[1597]&~m[1608]&m[1609]&~m[1611]&m[1612])|(m[1597]&m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1597]&m[1608]&m[1609]&m[1611]&m[1612]))&UnbiasedRNG[554])|((m[1597]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(~m[1597]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1597]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1597]&m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1597]&~m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1597]&~m[1608]&~m[1609]&m[1611]&m[1612])|(m[1597]&~m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1597]&m[1608]&~m[1609]&m[1611]&m[1612])|(m[1597]&m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1597]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1597]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1597]&m[1608]&m[1609]&m[1611]&m[1612]))):InitCond[1253];
    m[1615] = run?((((m[1602]&~m[1613]&~m[1614]&~m[1616]&~m[1617])|(~m[1602]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1602]&m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1602]&~m[1613]&m[1614]&m[1616]&~m[1617])|(~m[1602]&m[1613]&~m[1614]&~m[1616]&m[1617])|(~m[1602]&~m[1613]&m[1614]&~m[1616]&m[1617])|(m[1602]&m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1602]&m[1613]&m[1614]&m[1616]&m[1617]))&UnbiasedRNG[555])|((m[1602]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(~m[1602]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1602]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1602]&m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1602]&~m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1602]&~m[1613]&~m[1614]&m[1616]&m[1617])|(m[1602]&~m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1602]&m[1613]&~m[1614]&m[1616]&m[1617])|(m[1602]&m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1602]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1602]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1602]&m[1613]&m[1614]&m[1616]&m[1617]))):InitCond[1254];
    m[1620] = run?((((m[1607]&~m[1618]&~m[1619]&~m[1621]&~m[1622])|(~m[1607]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1607]&m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1607]&~m[1618]&m[1619]&m[1621]&~m[1622])|(~m[1607]&m[1618]&~m[1619]&~m[1621]&m[1622])|(~m[1607]&~m[1618]&m[1619]&~m[1621]&m[1622])|(m[1607]&m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1607]&m[1618]&m[1619]&m[1621]&m[1622]))&UnbiasedRNG[556])|((m[1607]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(~m[1607]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1607]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1607]&m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1607]&~m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1607]&~m[1618]&~m[1619]&m[1621]&m[1622])|(m[1607]&~m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1607]&m[1618]&~m[1619]&m[1621]&m[1622])|(m[1607]&m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1607]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1607]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1607]&m[1618]&m[1619]&m[1621]&m[1622]))):InitCond[1255];
    m[1625] = run?((((m[1617]&~m[1623]&~m[1624]&~m[1626]&~m[1627])|(~m[1617]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1617]&m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1617]&~m[1623]&m[1624]&m[1626]&~m[1627])|(~m[1617]&m[1623]&~m[1624]&~m[1626]&m[1627])|(~m[1617]&~m[1623]&m[1624]&~m[1626]&m[1627])|(m[1617]&m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1617]&m[1623]&m[1624]&m[1626]&m[1627]))&UnbiasedRNG[557])|((m[1617]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(~m[1617]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1617]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1617]&m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1617]&~m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1617]&~m[1623]&~m[1624]&m[1626]&m[1627])|(m[1617]&~m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1617]&m[1623]&~m[1624]&m[1626]&m[1627])|(m[1617]&m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1617]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1617]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1617]&m[1623]&m[1624]&m[1626]&m[1627]))):InitCond[1256];
    m[1630] = run?((((m[1622]&~m[1628]&~m[1629]&~m[1631]&~m[1632])|(~m[1622]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1622]&m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1622]&~m[1628]&m[1629]&m[1631]&~m[1632])|(~m[1622]&m[1628]&~m[1629]&~m[1631]&m[1632])|(~m[1622]&~m[1628]&m[1629]&~m[1631]&m[1632])|(m[1622]&m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1622]&m[1628]&m[1629]&m[1631]&m[1632]))&UnbiasedRNG[558])|((m[1622]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(~m[1622]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1622]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1622]&m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1622]&~m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1622]&~m[1628]&~m[1629]&m[1631]&m[1632])|(m[1622]&~m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1622]&m[1628]&~m[1629]&m[1631]&m[1632])|(m[1622]&m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1622]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1622]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1622]&m[1628]&m[1629]&m[1631]&m[1632]))):InitCond[1257];
    m[1635] = run?((((m[1632]&~m[1633]&~m[1634]&~m[1636]&~m[1637])|(~m[1632]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1632]&m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1632]&~m[1633]&m[1634]&m[1636]&~m[1637])|(~m[1632]&m[1633]&~m[1634]&~m[1636]&m[1637])|(~m[1632]&~m[1633]&m[1634]&~m[1636]&m[1637])|(m[1632]&m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1632]&m[1633]&m[1634]&m[1636]&m[1637]))&UnbiasedRNG[559])|((m[1632]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(~m[1632]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1632]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1632]&m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1632]&~m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1632]&~m[1633]&~m[1634]&m[1636]&m[1637])|(m[1632]&~m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1632]&m[1633]&~m[1634]&m[1636]&m[1637])|(m[1632]&m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1632]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1632]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1632]&m[1633]&m[1634]&m[1636]&m[1637]))):InitCond[1258];
end

always @(posedge color3_clk) begin
    m[736] = run?((((m[733]&~m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&~m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&m[737]&~m[738])|(~m[733]&~m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&m[737]&m[738])|(m[733]&~m[734]&m[735]&m[737]&m[738])|(~m[733]&m[734]&m[735]&m[737]&m[738]))&UnbiasedRNG[560])|((m[733]&m[734]&~m[735]&~m[737]&~m[738])|(m[733]&~m[734]&m[735]&~m[737]&~m[738])|(~m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&~m[734]&~m[735]&~m[737]&m[738])|(~m[733]&m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&~m[737]&m[738])|(~m[733]&~m[734]&m[735]&~m[737]&m[738])|(m[733]&~m[734]&m[735]&~m[737]&m[738])|(~m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&m[737]&m[738]))):InitCond[1259];
    m[746] = run?((((m[743]&~m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&~m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&m[747]&~m[748])|(~m[743]&~m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&m[747]&m[748])|(m[743]&~m[744]&m[745]&m[747]&m[748])|(~m[743]&m[744]&m[745]&m[747]&m[748]))&UnbiasedRNG[561])|((m[743]&m[744]&~m[745]&~m[747]&~m[748])|(m[743]&~m[744]&m[745]&~m[747]&~m[748])|(~m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&~m[744]&~m[745]&~m[747]&m[748])|(~m[743]&m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&~m[747]&m[748])|(~m[743]&~m[744]&m[745]&~m[747]&m[748])|(m[743]&~m[744]&m[745]&~m[747]&m[748])|(~m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&m[747]&m[748]))):InitCond[1260];
    m[751] = run?((((m[748]&~m[749]&~m[750]&~m[752]&~m[753])|(~m[748]&m[749]&~m[750]&~m[752]&~m[753])|(~m[748]&~m[749]&m[750]&~m[752]&~m[753])|(m[748]&m[749]&m[750]&m[752]&~m[753])|(~m[748]&~m[749]&~m[750]&~m[752]&m[753])|(m[748]&m[749]&~m[750]&m[752]&m[753])|(m[748]&~m[749]&m[750]&m[752]&m[753])|(~m[748]&m[749]&m[750]&m[752]&m[753]))&UnbiasedRNG[562])|((m[748]&m[749]&~m[750]&~m[752]&~m[753])|(m[748]&~m[749]&m[750]&~m[752]&~m[753])|(~m[748]&m[749]&m[750]&~m[752]&~m[753])|(m[748]&m[749]&m[750]&~m[752]&~m[753])|(m[748]&~m[749]&~m[750]&~m[752]&m[753])|(~m[748]&m[749]&~m[750]&~m[752]&m[753])|(m[748]&m[749]&~m[750]&~m[752]&m[753])|(~m[748]&~m[749]&m[750]&~m[752]&m[753])|(m[748]&~m[749]&m[750]&~m[752]&m[753])|(~m[748]&m[749]&m[750]&~m[752]&m[753])|(m[748]&m[749]&m[750]&~m[752]&m[753])|(m[748]&m[749]&m[750]&m[752]&m[753]))):InitCond[1261];
    m[761] = run?((((m[758]&~m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&~m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&m[762]&~m[763])|(~m[758]&~m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&m[762]&m[763])|(m[758]&~m[759]&m[760]&m[762]&m[763])|(~m[758]&m[759]&m[760]&m[762]&m[763]))&UnbiasedRNG[563])|((m[758]&m[759]&~m[760]&~m[762]&~m[763])|(m[758]&~m[759]&m[760]&~m[762]&~m[763])|(~m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&~m[759]&~m[760]&~m[762]&m[763])|(~m[758]&m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&~m[762]&m[763])|(~m[758]&~m[759]&m[760]&~m[762]&m[763])|(m[758]&~m[759]&m[760]&~m[762]&m[763])|(~m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&m[762]&m[763]))):InitCond[1262];
    m[766] = run?((((m[763]&~m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&~m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&m[767]&~m[768])|(~m[763]&~m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&m[767]&m[768])|(m[763]&~m[764]&m[765]&m[767]&m[768])|(~m[763]&m[764]&m[765]&m[767]&m[768]))&UnbiasedRNG[564])|((m[763]&m[764]&~m[765]&~m[767]&~m[768])|(m[763]&~m[764]&m[765]&~m[767]&~m[768])|(~m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&~m[764]&~m[765]&~m[767]&m[768])|(~m[763]&m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&~m[767]&m[768])|(~m[763]&~m[764]&m[765]&~m[767]&m[768])|(m[763]&~m[764]&m[765]&~m[767]&m[768])|(~m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&m[767]&m[768]))):InitCond[1263];
    m[771] = run?((((m[768]&~m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&~m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&m[772]&~m[773])|(~m[768]&~m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&m[772]&m[773])|(m[768]&~m[769]&m[770]&m[772]&m[773])|(~m[768]&m[769]&m[770]&m[772]&m[773]))&UnbiasedRNG[565])|((m[768]&m[769]&~m[770]&~m[772]&~m[773])|(m[768]&~m[769]&m[770]&~m[772]&~m[773])|(~m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&~m[769]&~m[770]&~m[772]&m[773])|(~m[768]&m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&~m[772]&m[773])|(~m[768]&~m[769]&m[770]&~m[772]&m[773])|(m[768]&~m[769]&m[770]&~m[772]&m[773])|(~m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&m[772]&m[773]))):InitCond[1264];
    m[781] = run?((((m[778]&~m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&~m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&m[782]&~m[783])|(~m[778]&~m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&m[782]&m[783])|(m[778]&~m[779]&m[780]&m[782]&m[783])|(~m[778]&m[779]&m[780]&m[782]&m[783]))&UnbiasedRNG[566])|((m[778]&m[779]&~m[780]&~m[782]&~m[783])|(m[778]&~m[779]&m[780]&~m[782]&~m[783])|(~m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&~m[779]&~m[780]&~m[782]&m[783])|(~m[778]&m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&~m[782]&m[783])|(~m[778]&~m[779]&m[780]&~m[782]&m[783])|(m[778]&~m[779]&m[780]&~m[782]&m[783])|(~m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&m[782]&m[783]))):InitCond[1265];
    m[786] = run?((((m[783]&~m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&~m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&m[787]&~m[788])|(~m[783]&~m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&m[787]&m[788])|(m[783]&~m[784]&m[785]&m[787]&m[788])|(~m[783]&m[784]&m[785]&m[787]&m[788]))&UnbiasedRNG[567])|((m[783]&m[784]&~m[785]&~m[787]&~m[788])|(m[783]&~m[784]&m[785]&~m[787]&~m[788])|(~m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&~m[784]&~m[785]&~m[787]&m[788])|(~m[783]&m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&~m[787]&m[788])|(~m[783]&~m[784]&m[785]&~m[787]&m[788])|(m[783]&~m[784]&m[785]&~m[787]&m[788])|(~m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&m[787]&m[788]))):InitCond[1266];
    m[791] = run?((((m[788]&~m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&~m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&m[792]&~m[793])|(~m[788]&~m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&m[792]&m[793])|(m[788]&~m[789]&m[790]&m[792]&m[793])|(~m[788]&m[789]&m[790]&m[792]&m[793]))&UnbiasedRNG[568])|((m[788]&m[789]&~m[790]&~m[792]&~m[793])|(m[788]&~m[789]&m[790]&~m[792]&~m[793])|(~m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&~m[789]&~m[790]&~m[792]&m[793])|(~m[788]&m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&~m[792]&m[793])|(~m[788]&~m[789]&m[790]&~m[792]&m[793])|(m[788]&~m[789]&m[790]&~m[792]&m[793])|(~m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&m[792]&m[793]))):InitCond[1267];
    m[796] = run?((((m[793]&~m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&~m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&m[797]&~m[798])|(~m[793]&~m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&m[797]&m[798])|(m[793]&~m[794]&m[795]&m[797]&m[798])|(~m[793]&m[794]&m[795]&m[797]&m[798]))&UnbiasedRNG[569])|((m[793]&m[794]&~m[795]&~m[797]&~m[798])|(m[793]&~m[794]&m[795]&~m[797]&~m[798])|(~m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&~m[794]&~m[795]&~m[797]&m[798])|(~m[793]&m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&~m[797]&m[798])|(~m[793]&~m[794]&m[795]&~m[797]&m[798])|(m[793]&~m[794]&m[795]&~m[797]&m[798])|(~m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&m[797]&m[798]))):InitCond[1268];
    m[806] = run?((((m[803]&~m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&~m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&m[807]&~m[808])|(~m[803]&~m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&m[807]&m[808])|(m[803]&~m[804]&m[805]&m[807]&m[808])|(~m[803]&m[804]&m[805]&m[807]&m[808]))&UnbiasedRNG[570])|((m[803]&m[804]&~m[805]&~m[807]&~m[808])|(m[803]&~m[804]&m[805]&~m[807]&~m[808])|(~m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&~m[804]&~m[805]&~m[807]&m[808])|(~m[803]&m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&~m[807]&m[808])|(~m[803]&~m[804]&m[805]&~m[807]&m[808])|(m[803]&~m[804]&m[805]&~m[807]&m[808])|(~m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&m[807]&m[808]))):InitCond[1269];
    m[811] = run?((((m[808]&~m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&~m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&m[812]&~m[813])|(~m[808]&~m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&m[812]&m[813])|(m[808]&~m[809]&m[810]&m[812]&m[813])|(~m[808]&m[809]&m[810]&m[812]&m[813]))&UnbiasedRNG[571])|((m[808]&m[809]&~m[810]&~m[812]&~m[813])|(m[808]&~m[809]&m[810]&~m[812]&~m[813])|(~m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&~m[809]&~m[810]&~m[812]&m[813])|(~m[808]&m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&~m[812]&m[813])|(~m[808]&~m[809]&m[810]&~m[812]&m[813])|(m[808]&~m[809]&m[810]&~m[812]&m[813])|(~m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&m[812]&m[813]))):InitCond[1270];
    m[816] = run?((((m[813]&~m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&~m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&m[817]&~m[818])|(~m[813]&~m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&m[817]&m[818])|(m[813]&~m[814]&m[815]&m[817]&m[818])|(~m[813]&m[814]&m[815]&m[817]&m[818]))&UnbiasedRNG[572])|((m[813]&m[814]&~m[815]&~m[817]&~m[818])|(m[813]&~m[814]&m[815]&~m[817]&~m[818])|(~m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&~m[814]&~m[815]&~m[817]&m[818])|(~m[813]&m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&~m[817]&m[818])|(~m[813]&~m[814]&m[815]&~m[817]&m[818])|(m[813]&~m[814]&m[815]&~m[817]&m[818])|(~m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&m[817]&m[818]))):InitCond[1271];
    m[821] = run?((((m[818]&~m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&~m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&m[822]&~m[823])|(~m[818]&~m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&m[822]&m[823])|(m[818]&~m[819]&m[820]&m[822]&m[823])|(~m[818]&m[819]&m[820]&m[822]&m[823]))&UnbiasedRNG[573])|((m[818]&m[819]&~m[820]&~m[822]&~m[823])|(m[818]&~m[819]&m[820]&~m[822]&~m[823])|(~m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&~m[819]&~m[820]&~m[822]&m[823])|(~m[818]&m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&~m[822]&m[823])|(~m[818]&~m[819]&m[820]&~m[822]&m[823])|(m[818]&~m[819]&m[820]&~m[822]&m[823])|(~m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&m[822]&m[823]))):InitCond[1272];
    m[826] = run?((((m[823]&~m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&~m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&m[827]&~m[828])|(~m[823]&~m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&m[827]&m[828])|(m[823]&~m[824]&m[825]&m[827]&m[828])|(~m[823]&m[824]&m[825]&m[827]&m[828]))&UnbiasedRNG[574])|((m[823]&m[824]&~m[825]&~m[827]&~m[828])|(m[823]&~m[824]&m[825]&~m[827]&~m[828])|(~m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&~m[824]&~m[825]&~m[827]&m[828])|(~m[823]&m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&~m[827]&m[828])|(~m[823]&~m[824]&m[825]&~m[827]&m[828])|(m[823]&~m[824]&m[825]&~m[827]&m[828])|(~m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&m[827]&m[828]))):InitCond[1273];
    m[836] = run?((((m[833]&~m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&~m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&m[837]&~m[838])|(~m[833]&~m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&m[837]&m[838])|(m[833]&~m[834]&m[835]&m[837]&m[838])|(~m[833]&m[834]&m[835]&m[837]&m[838]))&UnbiasedRNG[575])|((m[833]&m[834]&~m[835]&~m[837]&~m[838])|(m[833]&~m[834]&m[835]&~m[837]&~m[838])|(~m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&~m[834]&~m[835]&~m[837]&m[838])|(~m[833]&m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&~m[837]&m[838])|(~m[833]&~m[834]&m[835]&~m[837]&m[838])|(m[833]&~m[834]&m[835]&~m[837]&m[838])|(~m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&m[837]&m[838]))):InitCond[1274];
    m[841] = run?((((m[838]&~m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&~m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&m[842]&~m[843])|(~m[838]&~m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&m[842]&m[843])|(m[838]&~m[839]&m[840]&m[842]&m[843])|(~m[838]&m[839]&m[840]&m[842]&m[843]))&UnbiasedRNG[576])|((m[838]&m[839]&~m[840]&~m[842]&~m[843])|(m[838]&~m[839]&m[840]&~m[842]&~m[843])|(~m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&~m[839]&~m[840]&~m[842]&m[843])|(~m[838]&m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&~m[842]&m[843])|(~m[838]&~m[839]&m[840]&~m[842]&m[843])|(m[838]&~m[839]&m[840]&~m[842]&m[843])|(~m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&m[842]&m[843]))):InitCond[1275];
    m[846] = run?((((m[843]&~m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&~m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&m[847]&~m[848])|(~m[843]&~m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&m[847]&m[848])|(m[843]&~m[844]&m[845]&m[847]&m[848])|(~m[843]&m[844]&m[845]&m[847]&m[848]))&UnbiasedRNG[577])|((m[843]&m[844]&~m[845]&~m[847]&~m[848])|(m[843]&~m[844]&m[845]&~m[847]&~m[848])|(~m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&~m[844]&~m[845]&~m[847]&m[848])|(~m[843]&m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&~m[847]&m[848])|(~m[843]&~m[844]&m[845]&~m[847]&m[848])|(m[843]&~m[844]&m[845]&~m[847]&m[848])|(~m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&m[847]&m[848]))):InitCond[1276];
    m[851] = run?((((m[848]&~m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&~m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&m[852]&~m[853])|(~m[848]&~m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&m[852]&m[853])|(m[848]&~m[849]&m[850]&m[852]&m[853])|(~m[848]&m[849]&m[850]&m[852]&m[853]))&UnbiasedRNG[578])|((m[848]&m[849]&~m[850]&~m[852]&~m[853])|(m[848]&~m[849]&m[850]&~m[852]&~m[853])|(~m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&~m[849]&~m[850]&~m[852]&m[853])|(~m[848]&m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&~m[852]&m[853])|(~m[848]&~m[849]&m[850]&~m[852]&m[853])|(m[848]&~m[849]&m[850]&~m[852]&m[853])|(~m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&m[852]&m[853]))):InitCond[1277];
    m[856] = run?((((m[853]&~m[854]&~m[855]&~m[857]&~m[858])|(~m[853]&m[854]&~m[855]&~m[857]&~m[858])|(~m[853]&~m[854]&m[855]&~m[857]&~m[858])|(m[853]&m[854]&m[855]&m[857]&~m[858])|(~m[853]&~m[854]&~m[855]&~m[857]&m[858])|(m[853]&m[854]&~m[855]&m[857]&m[858])|(m[853]&~m[854]&m[855]&m[857]&m[858])|(~m[853]&m[854]&m[855]&m[857]&m[858]))&UnbiasedRNG[579])|((m[853]&m[854]&~m[855]&~m[857]&~m[858])|(m[853]&~m[854]&m[855]&~m[857]&~m[858])|(~m[853]&m[854]&m[855]&~m[857]&~m[858])|(m[853]&m[854]&m[855]&~m[857]&~m[858])|(m[853]&~m[854]&~m[855]&~m[857]&m[858])|(~m[853]&m[854]&~m[855]&~m[857]&m[858])|(m[853]&m[854]&~m[855]&~m[857]&m[858])|(~m[853]&~m[854]&m[855]&~m[857]&m[858])|(m[853]&~m[854]&m[855]&~m[857]&m[858])|(~m[853]&m[854]&m[855]&~m[857]&m[858])|(m[853]&m[854]&m[855]&~m[857]&m[858])|(m[853]&m[854]&m[855]&m[857]&m[858]))):InitCond[1278];
    m[861] = run?((((m[858]&~m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&~m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&m[862]&~m[863])|(~m[858]&~m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&m[862]&m[863])|(m[858]&~m[859]&m[860]&m[862]&m[863])|(~m[858]&m[859]&m[860]&m[862]&m[863]))&UnbiasedRNG[580])|((m[858]&m[859]&~m[860]&~m[862]&~m[863])|(m[858]&~m[859]&m[860]&~m[862]&~m[863])|(~m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&~m[859]&~m[860]&~m[862]&m[863])|(~m[858]&m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&~m[862]&m[863])|(~m[858]&~m[859]&m[860]&~m[862]&m[863])|(m[858]&~m[859]&m[860]&~m[862]&m[863])|(~m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&m[862]&m[863]))):InitCond[1279];
    m[871] = run?((((m[868]&~m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&~m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&m[872]&~m[873])|(~m[868]&~m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&m[872]&m[873])|(m[868]&~m[869]&m[870]&m[872]&m[873])|(~m[868]&m[869]&m[870]&m[872]&m[873]))&UnbiasedRNG[581])|((m[868]&m[869]&~m[870]&~m[872]&~m[873])|(m[868]&~m[869]&m[870]&~m[872]&~m[873])|(~m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&~m[869]&~m[870]&~m[872]&m[873])|(~m[868]&m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&~m[872]&m[873])|(~m[868]&~m[869]&m[870]&~m[872]&m[873])|(m[868]&~m[869]&m[870]&~m[872]&m[873])|(~m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&m[872]&m[873]))):InitCond[1280];
    m[876] = run?((((m[873]&~m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&~m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&m[877]&~m[878])|(~m[873]&~m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&m[877]&m[878])|(m[873]&~m[874]&m[875]&m[877]&m[878])|(~m[873]&m[874]&m[875]&m[877]&m[878]))&UnbiasedRNG[582])|((m[873]&m[874]&~m[875]&~m[877]&~m[878])|(m[873]&~m[874]&m[875]&~m[877]&~m[878])|(~m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&~m[874]&~m[875]&~m[877]&m[878])|(~m[873]&m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&~m[877]&m[878])|(~m[873]&~m[874]&m[875]&~m[877]&m[878])|(m[873]&~m[874]&m[875]&~m[877]&m[878])|(~m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&m[877]&m[878]))):InitCond[1281];
    m[881] = run?((((m[878]&~m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&~m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&m[882]&~m[883])|(~m[878]&~m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&m[882]&m[883])|(m[878]&~m[879]&m[880]&m[882]&m[883])|(~m[878]&m[879]&m[880]&m[882]&m[883]))&UnbiasedRNG[583])|((m[878]&m[879]&~m[880]&~m[882]&~m[883])|(m[878]&~m[879]&m[880]&~m[882]&~m[883])|(~m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&~m[879]&~m[880]&~m[882]&m[883])|(~m[878]&m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&~m[882]&m[883])|(~m[878]&~m[879]&m[880]&~m[882]&m[883])|(m[878]&~m[879]&m[880]&~m[882]&m[883])|(~m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&m[882]&m[883]))):InitCond[1282];
    m[886] = run?((((m[883]&~m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&~m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&m[887]&~m[888])|(~m[883]&~m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&m[887]&m[888])|(m[883]&~m[884]&m[885]&m[887]&m[888])|(~m[883]&m[884]&m[885]&m[887]&m[888]))&UnbiasedRNG[584])|((m[883]&m[884]&~m[885]&~m[887]&~m[888])|(m[883]&~m[884]&m[885]&~m[887]&~m[888])|(~m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&~m[884]&~m[885]&~m[887]&m[888])|(~m[883]&m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&~m[887]&m[888])|(~m[883]&~m[884]&m[885]&~m[887]&m[888])|(m[883]&~m[884]&m[885]&~m[887]&m[888])|(~m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&m[887]&m[888]))):InitCond[1283];
    m[891] = run?((((m[888]&~m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&~m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&m[892]&~m[893])|(~m[888]&~m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&m[892]&m[893])|(m[888]&~m[889]&m[890]&m[892]&m[893])|(~m[888]&m[889]&m[890]&m[892]&m[893]))&UnbiasedRNG[585])|((m[888]&m[889]&~m[890]&~m[892]&~m[893])|(m[888]&~m[889]&m[890]&~m[892]&~m[893])|(~m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&~m[889]&~m[890]&~m[892]&m[893])|(~m[888]&m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&~m[892]&m[893])|(~m[888]&~m[889]&m[890]&~m[892]&m[893])|(m[888]&~m[889]&m[890]&~m[892]&m[893])|(~m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&m[892]&m[893]))):InitCond[1284];
    m[896] = run?((((m[893]&~m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&~m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&m[897]&~m[898])|(~m[893]&~m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&m[897]&m[898])|(m[893]&~m[894]&m[895]&m[897]&m[898])|(~m[893]&m[894]&m[895]&m[897]&m[898]))&UnbiasedRNG[586])|((m[893]&m[894]&~m[895]&~m[897]&~m[898])|(m[893]&~m[894]&m[895]&~m[897]&~m[898])|(~m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&~m[894]&~m[895]&~m[897]&m[898])|(~m[893]&m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&~m[897]&m[898])|(~m[893]&~m[894]&m[895]&~m[897]&m[898])|(m[893]&~m[894]&m[895]&~m[897]&m[898])|(~m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&m[897]&m[898]))):InitCond[1285];
    m[901] = run?((((m[898]&~m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&~m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&m[902]&~m[903])|(~m[898]&~m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&m[902]&m[903])|(m[898]&~m[899]&m[900]&m[902]&m[903])|(~m[898]&m[899]&m[900]&m[902]&m[903]))&UnbiasedRNG[587])|((m[898]&m[899]&~m[900]&~m[902]&~m[903])|(m[898]&~m[899]&m[900]&~m[902]&~m[903])|(~m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&~m[899]&~m[900]&~m[902]&m[903])|(~m[898]&m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&~m[902]&m[903])|(~m[898]&~m[899]&m[900]&~m[902]&m[903])|(m[898]&~m[899]&m[900]&~m[902]&m[903])|(~m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&m[902]&m[903]))):InitCond[1286];
    m[911] = run?((((m[908]&~m[909]&~m[910]&~m[912]&~m[913])|(~m[908]&m[909]&~m[910]&~m[912]&~m[913])|(~m[908]&~m[909]&m[910]&~m[912]&~m[913])|(m[908]&m[909]&m[910]&m[912]&~m[913])|(~m[908]&~m[909]&~m[910]&~m[912]&m[913])|(m[908]&m[909]&~m[910]&m[912]&m[913])|(m[908]&~m[909]&m[910]&m[912]&m[913])|(~m[908]&m[909]&m[910]&m[912]&m[913]))&UnbiasedRNG[588])|((m[908]&m[909]&~m[910]&~m[912]&~m[913])|(m[908]&~m[909]&m[910]&~m[912]&~m[913])|(~m[908]&m[909]&m[910]&~m[912]&~m[913])|(m[908]&m[909]&m[910]&~m[912]&~m[913])|(m[908]&~m[909]&~m[910]&~m[912]&m[913])|(~m[908]&m[909]&~m[910]&~m[912]&m[913])|(m[908]&m[909]&~m[910]&~m[912]&m[913])|(~m[908]&~m[909]&m[910]&~m[912]&m[913])|(m[908]&~m[909]&m[910]&~m[912]&m[913])|(~m[908]&m[909]&m[910]&~m[912]&m[913])|(m[908]&m[909]&m[910]&~m[912]&m[913])|(m[908]&m[909]&m[910]&m[912]&m[913]))):InitCond[1287];
    m[916] = run?((((m[913]&~m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&~m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&m[917]&~m[918])|(~m[913]&~m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&m[917]&m[918])|(m[913]&~m[914]&m[915]&m[917]&m[918])|(~m[913]&m[914]&m[915]&m[917]&m[918]))&UnbiasedRNG[589])|((m[913]&m[914]&~m[915]&~m[917]&~m[918])|(m[913]&~m[914]&m[915]&~m[917]&~m[918])|(~m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&~m[914]&~m[915]&~m[917]&m[918])|(~m[913]&m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&~m[917]&m[918])|(~m[913]&~m[914]&m[915]&~m[917]&m[918])|(m[913]&~m[914]&m[915]&~m[917]&m[918])|(~m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&m[917]&m[918]))):InitCond[1288];
    m[921] = run?((((m[918]&~m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&~m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&m[922]&~m[923])|(~m[918]&~m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&m[922]&m[923])|(m[918]&~m[919]&m[920]&m[922]&m[923])|(~m[918]&m[919]&m[920]&m[922]&m[923]))&UnbiasedRNG[590])|((m[918]&m[919]&~m[920]&~m[922]&~m[923])|(m[918]&~m[919]&m[920]&~m[922]&~m[923])|(~m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&~m[919]&~m[920]&~m[922]&m[923])|(~m[918]&m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&~m[922]&m[923])|(~m[918]&~m[919]&m[920]&~m[922]&m[923])|(m[918]&~m[919]&m[920]&~m[922]&m[923])|(~m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&m[922]&m[923]))):InitCond[1289];
    m[926] = run?((((m[923]&~m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&~m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&m[927]&~m[928])|(~m[923]&~m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&m[927]&m[928])|(m[923]&~m[924]&m[925]&m[927]&m[928])|(~m[923]&m[924]&m[925]&m[927]&m[928]))&UnbiasedRNG[591])|((m[923]&m[924]&~m[925]&~m[927]&~m[928])|(m[923]&~m[924]&m[925]&~m[927]&~m[928])|(~m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&~m[924]&~m[925]&~m[927]&m[928])|(~m[923]&m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&~m[927]&m[928])|(~m[923]&~m[924]&m[925]&~m[927]&m[928])|(m[923]&~m[924]&m[925]&~m[927]&m[928])|(~m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&m[927]&m[928]))):InitCond[1290];
    m[931] = run?((((m[928]&~m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&~m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&m[932]&~m[933])|(~m[928]&~m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&m[932]&m[933])|(m[928]&~m[929]&m[930]&m[932]&m[933])|(~m[928]&m[929]&m[930]&m[932]&m[933]))&UnbiasedRNG[592])|((m[928]&m[929]&~m[930]&~m[932]&~m[933])|(m[928]&~m[929]&m[930]&~m[932]&~m[933])|(~m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&~m[929]&~m[930]&~m[932]&m[933])|(~m[928]&m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&~m[932]&m[933])|(~m[928]&~m[929]&m[930]&~m[932]&m[933])|(m[928]&~m[929]&m[930]&~m[932]&m[933])|(~m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&m[932]&m[933]))):InitCond[1291];
    m[936] = run?((((m[933]&~m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&~m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&m[937]&~m[938])|(~m[933]&~m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&m[937]&m[938])|(m[933]&~m[934]&m[935]&m[937]&m[938])|(~m[933]&m[934]&m[935]&m[937]&m[938]))&UnbiasedRNG[593])|((m[933]&m[934]&~m[935]&~m[937]&~m[938])|(m[933]&~m[934]&m[935]&~m[937]&~m[938])|(~m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&~m[934]&~m[935]&~m[937]&m[938])|(~m[933]&m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&~m[937]&m[938])|(~m[933]&~m[934]&m[935]&~m[937]&m[938])|(m[933]&~m[934]&m[935]&~m[937]&m[938])|(~m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&m[937]&m[938]))):InitCond[1292];
    m[941] = run?((((m[938]&~m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&~m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&m[942]&~m[943])|(~m[938]&~m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&m[942]&m[943])|(m[938]&~m[939]&m[940]&m[942]&m[943])|(~m[938]&m[939]&m[940]&m[942]&m[943]))&UnbiasedRNG[594])|((m[938]&m[939]&~m[940]&~m[942]&~m[943])|(m[938]&~m[939]&m[940]&~m[942]&~m[943])|(~m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&~m[939]&~m[940]&~m[942]&m[943])|(~m[938]&m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&~m[942]&m[943])|(~m[938]&~m[939]&m[940]&~m[942]&m[943])|(m[938]&~m[939]&m[940]&~m[942]&m[943])|(~m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&m[942]&m[943]))):InitCond[1293];
    m[946] = run?((((m[943]&~m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&~m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&m[947]&~m[948])|(~m[943]&~m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&m[947]&m[948])|(m[943]&~m[944]&m[945]&m[947]&m[948])|(~m[943]&m[944]&m[945]&m[947]&m[948]))&UnbiasedRNG[595])|((m[943]&m[944]&~m[945]&~m[947]&~m[948])|(m[943]&~m[944]&m[945]&~m[947]&~m[948])|(~m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&~m[944]&~m[945]&~m[947]&m[948])|(~m[943]&m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&~m[947]&m[948])|(~m[943]&~m[944]&m[945]&~m[947]&m[948])|(m[943]&~m[944]&m[945]&~m[947]&m[948])|(~m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&m[947]&m[948]))):InitCond[1294];
    m[956] = run?((((m[953]&~m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&~m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&m[957]&~m[958])|(~m[953]&~m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&m[957]&m[958])|(m[953]&~m[954]&m[955]&m[957]&m[958])|(~m[953]&m[954]&m[955]&m[957]&m[958]))&UnbiasedRNG[596])|((m[953]&m[954]&~m[955]&~m[957]&~m[958])|(m[953]&~m[954]&m[955]&~m[957]&~m[958])|(~m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&~m[954]&~m[955]&~m[957]&m[958])|(~m[953]&m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&~m[957]&m[958])|(~m[953]&~m[954]&m[955]&~m[957]&m[958])|(m[953]&~m[954]&m[955]&~m[957]&m[958])|(~m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&m[957]&m[958]))):InitCond[1295];
    m[961] = run?((((m[958]&~m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&~m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&m[962]&~m[963])|(~m[958]&~m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&m[962]&m[963])|(m[958]&~m[959]&m[960]&m[962]&m[963])|(~m[958]&m[959]&m[960]&m[962]&m[963]))&UnbiasedRNG[597])|((m[958]&m[959]&~m[960]&~m[962]&~m[963])|(m[958]&~m[959]&m[960]&~m[962]&~m[963])|(~m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&~m[959]&~m[960]&~m[962]&m[963])|(~m[958]&m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&~m[962]&m[963])|(~m[958]&~m[959]&m[960]&~m[962]&m[963])|(m[958]&~m[959]&m[960]&~m[962]&m[963])|(~m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&m[962]&m[963]))):InitCond[1296];
    m[966] = run?((((m[963]&~m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&~m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&m[967]&~m[968])|(~m[963]&~m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&m[967]&m[968])|(m[963]&~m[964]&m[965]&m[967]&m[968])|(~m[963]&m[964]&m[965]&m[967]&m[968]))&UnbiasedRNG[598])|((m[963]&m[964]&~m[965]&~m[967]&~m[968])|(m[963]&~m[964]&m[965]&~m[967]&~m[968])|(~m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&~m[964]&~m[965]&~m[967]&m[968])|(~m[963]&m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&~m[967]&m[968])|(~m[963]&~m[964]&m[965]&~m[967]&m[968])|(m[963]&~m[964]&m[965]&~m[967]&m[968])|(~m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&m[967]&m[968]))):InitCond[1297];
    m[971] = run?((((m[968]&~m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&~m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&m[972]&~m[973])|(~m[968]&~m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&m[972]&m[973])|(m[968]&~m[969]&m[970]&m[972]&m[973])|(~m[968]&m[969]&m[970]&m[972]&m[973]))&UnbiasedRNG[599])|((m[968]&m[969]&~m[970]&~m[972]&~m[973])|(m[968]&~m[969]&m[970]&~m[972]&~m[973])|(~m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&~m[969]&~m[970]&~m[972]&m[973])|(~m[968]&m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&~m[972]&m[973])|(~m[968]&~m[969]&m[970]&~m[972]&m[973])|(m[968]&~m[969]&m[970]&~m[972]&m[973])|(~m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&m[972]&m[973]))):InitCond[1298];
    m[976] = run?((((m[973]&~m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&~m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&m[977]&~m[978])|(~m[973]&~m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&m[977]&m[978])|(m[973]&~m[974]&m[975]&m[977]&m[978])|(~m[973]&m[974]&m[975]&m[977]&m[978]))&UnbiasedRNG[600])|((m[973]&m[974]&~m[975]&~m[977]&~m[978])|(m[973]&~m[974]&m[975]&~m[977]&~m[978])|(~m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&~m[974]&~m[975]&~m[977]&m[978])|(~m[973]&m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&~m[977]&m[978])|(~m[973]&~m[974]&m[975]&~m[977]&m[978])|(m[973]&~m[974]&m[975]&~m[977]&m[978])|(~m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&m[977]&m[978]))):InitCond[1299];
    m[981] = run?((((m[978]&~m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&~m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&m[982]&~m[983])|(~m[978]&~m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&m[982]&m[983])|(m[978]&~m[979]&m[980]&m[982]&m[983])|(~m[978]&m[979]&m[980]&m[982]&m[983]))&UnbiasedRNG[601])|((m[978]&m[979]&~m[980]&~m[982]&~m[983])|(m[978]&~m[979]&m[980]&~m[982]&~m[983])|(~m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&~m[979]&~m[980]&~m[982]&m[983])|(~m[978]&m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&~m[982]&m[983])|(~m[978]&~m[979]&m[980]&~m[982]&m[983])|(m[978]&~m[979]&m[980]&~m[982]&m[983])|(~m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&m[982]&m[983]))):InitCond[1300];
    m[986] = run?((((m[983]&~m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&~m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&m[987]&~m[988])|(~m[983]&~m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&m[987]&m[988])|(m[983]&~m[984]&m[985]&m[987]&m[988])|(~m[983]&m[984]&m[985]&m[987]&m[988]))&UnbiasedRNG[602])|((m[983]&m[984]&~m[985]&~m[987]&~m[988])|(m[983]&~m[984]&m[985]&~m[987]&~m[988])|(~m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&~m[984]&~m[985]&~m[987]&m[988])|(~m[983]&m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&~m[987]&m[988])|(~m[983]&~m[984]&m[985]&~m[987]&m[988])|(m[983]&~m[984]&m[985]&~m[987]&m[988])|(~m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&m[987]&m[988]))):InitCond[1301];
    m[991] = run?((((m[988]&~m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&~m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&m[992]&~m[993])|(~m[988]&~m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&m[992]&m[993])|(m[988]&~m[989]&m[990]&m[992]&m[993])|(~m[988]&m[989]&m[990]&m[992]&m[993]))&UnbiasedRNG[603])|((m[988]&m[989]&~m[990]&~m[992]&~m[993])|(m[988]&~m[989]&m[990]&~m[992]&~m[993])|(~m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&~m[989]&~m[990]&~m[992]&m[993])|(~m[988]&m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&~m[992]&m[993])|(~m[988]&~m[989]&m[990]&~m[992]&m[993])|(m[988]&~m[989]&m[990]&~m[992]&m[993])|(~m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&m[992]&m[993]))):InitCond[1302];
    m[996] = run?((((m[993]&~m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&~m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&m[997]&~m[998])|(~m[993]&~m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&m[997]&m[998])|(m[993]&~m[994]&m[995]&m[997]&m[998])|(~m[993]&m[994]&m[995]&m[997]&m[998]))&UnbiasedRNG[604])|((m[993]&m[994]&~m[995]&~m[997]&~m[998])|(m[993]&~m[994]&m[995]&~m[997]&~m[998])|(~m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&~m[994]&~m[995]&~m[997]&m[998])|(~m[993]&m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&~m[997]&m[998])|(~m[993]&~m[994]&m[995]&~m[997]&m[998])|(m[993]&~m[994]&m[995]&~m[997]&m[998])|(~m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&m[997]&m[998]))):InitCond[1303];
    m[1006] = run?((((m[1003]&~m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&~m[1008])|(~m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&m[1007]&m[1008]))&UnbiasedRNG[605])|((m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&m[1008]))):InitCond[1304];
    m[1011] = run?((((m[1008]&~m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&~m[1013])|(~m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))&UnbiasedRNG[606])|((m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))):InitCond[1305];
    m[1016] = run?((((m[1013]&~m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&~m[1018])|(~m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))&UnbiasedRNG[607])|((m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))):InitCond[1306];
    m[1021] = run?((((m[1018]&~m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&~m[1023])|(~m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))&UnbiasedRNG[608])|((m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))):InitCond[1307];
    m[1026] = run?((((m[1023]&~m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&~m[1028])|(~m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))&UnbiasedRNG[609])|((m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))):InitCond[1308];
    m[1031] = run?((((m[1028]&~m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&~m[1033])|(~m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&m[1032]&m[1033]))&UnbiasedRNG[610])|((m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&m[1033]))):InitCond[1309];
    m[1036] = run?((((m[1033]&~m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&~m[1038])|(~m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))&UnbiasedRNG[611])|((m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))):InitCond[1310];
    m[1041] = run?((((m[1038]&~m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&~m[1043])|(~m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))&UnbiasedRNG[612])|((m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))):InitCond[1311];
    m[1046] = run?((((m[1043]&~m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&~m[1048])|(~m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&m[1047]&m[1048]))&UnbiasedRNG[613])|((m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&m[1048]))):InitCond[1312];
    m[1051] = run?((((m[1048]&~m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&~m[1053])|(~m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))&UnbiasedRNG[614])|((m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))):InitCond[1313];
    m[1061] = run?((((m[1058]&~m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&~m[1063])|(~m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))&UnbiasedRNG[615])|((m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))):InitCond[1314];
    m[1066] = run?((((m[1063]&~m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&~m[1068])|(~m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&m[1067]&m[1068]))&UnbiasedRNG[616])|((m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&m[1068]))):InitCond[1315];
    m[1071] = run?((((m[1068]&~m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&~m[1073])|(~m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))&UnbiasedRNG[617])|((m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))):InitCond[1316];
    m[1076] = run?((((m[1073]&~m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&~m[1078])|(~m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))&UnbiasedRNG[618])|((m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))):InitCond[1317];
    m[1081] = run?((((m[1078]&~m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&~m[1083])|(~m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&m[1082]&m[1083]))&UnbiasedRNG[619])|((m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&m[1083]))):InitCond[1318];
    m[1086] = run?((((m[1083]&~m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&~m[1088])|(~m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))&UnbiasedRNG[620])|((m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))):InitCond[1319];
    m[1091] = run?((((m[1088]&~m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&~m[1093])|(~m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))&UnbiasedRNG[621])|((m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))):InitCond[1320];
    m[1096] = run?((((m[1093]&~m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&~m[1098])|(~m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))&UnbiasedRNG[622])|((m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))):InitCond[1321];
    m[1101] = run?((((m[1098]&~m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&~m[1103])|(~m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))&UnbiasedRNG[623])|((m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))):InitCond[1322];
    m[1106] = run?((((m[1103]&~m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&~m[1108])|(~m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&m[1107]&m[1108]))&UnbiasedRNG[624])|((m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&m[1108]))):InitCond[1323];
    m[1111] = run?((((m[1108]&~m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&~m[1113])|(~m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&m[1112]&m[1113]))&UnbiasedRNG[625])|((m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&m[1113]))):InitCond[1324];
    m[1121] = run?((((m[1118]&~m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&~m[1123])|(~m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))&UnbiasedRNG[626])|((m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))):InitCond[1325];
    m[1126] = run?((((m[1123]&~m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&~m[1128])|(~m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))&UnbiasedRNG[627])|((m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))):InitCond[1326];
    m[1131] = run?((((m[1128]&~m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&~m[1133])|(~m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))&UnbiasedRNG[628])|((m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))):InitCond[1327];
    m[1136] = run?((((m[1133]&~m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&~m[1138])|(~m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&m[1137]&m[1138]))&UnbiasedRNG[629])|((m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&m[1138]))):InitCond[1328];
    m[1141] = run?((((m[1138]&~m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&~m[1143])|(~m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))&UnbiasedRNG[630])|((m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))):InitCond[1329];
    m[1146] = run?((((m[1143]&~m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&~m[1148])|(~m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))&UnbiasedRNG[631])|((m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))):InitCond[1330];
    m[1151] = run?((((m[1148]&~m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&~m[1153])|(~m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&m[1152]&m[1153]))&UnbiasedRNG[632])|((m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&m[1153]))):InitCond[1331];
    m[1156] = run?((((m[1153]&~m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&~m[1158])|(~m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&m[1157]&m[1158]))&UnbiasedRNG[633])|((m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&m[1158]))):InitCond[1332];
    m[1161] = run?((((m[1158]&~m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&~m[1163])|(~m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))&UnbiasedRNG[634])|((m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))):InitCond[1333];
    m[1166] = run?((((m[1163]&~m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&~m[1168])|(~m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))&UnbiasedRNG[635])|((m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))):InitCond[1334];
    m[1171] = run?((((m[1168]&~m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&~m[1173])|(~m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&m[1172]&m[1173]))&UnbiasedRNG[636])|((m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&m[1173]))):InitCond[1335];
    m[1176] = run?((((m[1173]&~m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&~m[1178])|(~m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))&UnbiasedRNG[637])|((m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))):InitCond[1336];
    m[1186] = run?((((m[1183]&~m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&~m[1188])|(~m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&m[1187]&m[1188]))&UnbiasedRNG[638])|((m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&m[1188]))):InitCond[1337];
    m[1191] = run?((((m[1188]&~m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&~m[1193])|(~m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&m[1192]&m[1193]))&UnbiasedRNG[639])|((m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&m[1193]))):InitCond[1338];
    m[1196] = run?((((m[1193]&~m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&~m[1198])|(~m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&m[1197]&m[1198]))&UnbiasedRNG[640])|((m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&m[1198]))):InitCond[1339];
    m[1201] = run?((((m[1198]&~m[1199]&~m[1200]&~m[1202]&~m[1203])|(~m[1198]&m[1199]&~m[1200]&~m[1202]&~m[1203])|(~m[1198]&~m[1199]&m[1200]&~m[1202]&~m[1203])|(m[1198]&m[1199]&m[1200]&m[1202]&~m[1203])|(~m[1198]&~m[1199]&~m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&~m[1200]&m[1202]&m[1203])|(m[1198]&~m[1199]&m[1200]&m[1202]&m[1203])|(~m[1198]&m[1199]&m[1200]&m[1202]&m[1203]))&UnbiasedRNG[641])|((m[1198]&m[1199]&~m[1200]&~m[1202]&~m[1203])|(m[1198]&~m[1199]&m[1200]&~m[1202]&~m[1203])|(~m[1198]&m[1199]&m[1200]&~m[1202]&~m[1203])|(m[1198]&m[1199]&m[1200]&~m[1202]&~m[1203])|(m[1198]&~m[1199]&~m[1200]&~m[1202]&m[1203])|(~m[1198]&m[1199]&~m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&~m[1200]&~m[1202]&m[1203])|(~m[1198]&~m[1199]&m[1200]&~m[1202]&m[1203])|(m[1198]&~m[1199]&m[1200]&~m[1202]&m[1203])|(~m[1198]&m[1199]&m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&m[1200]&m[1202]&m[1203]))):InitCond[1340];
    m[1206] = run?((((m[1203]&~m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&~m[1208])|(~m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&m[1207]&m[1208]))&UnbiasedRNG[642])|((m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&m[1208]))):InitCond[1341];
    m[1211] = run?((((m[1208]&~m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&~m[1213])|(~m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&m[1212]&m[1213]))&UnbiasedRNG[643])|((m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&m[1213]))):InitCond[1342];
    m[1216] = run?((((m[1213]&~m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&~m[1218])|(~m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&m[1217]&m[1218]))&UnbiasedRNG[644])|((m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&m[1218]))):InitCond[1343];
    m[1221] = run?((((m[1218]&~m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&~m[1223])|(~m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&m[1222]&m[1223]))&UnbiasedRNG[645])|((m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&m[1223]))):InitCond[1344];
    m[1226] = run?((((m[1223]&~m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&~m[1228])|(~m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&m[1227]&m[1228]))&UnbiasedRNG[646])|((m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&m[1228]))):InitCond[1345];
    m[1231] = run?((((m[1228]&~m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&~m[1233])|(~m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&m[1232]&m[1233]))&UnbiasedRNG[647])|((m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&m[1233]))):InitCond[1346];
    m[1236] = run?((((m[1233]&~m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&~m[1238])|(~m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&m[1237]&m[1238]))&UnbiasedRNG[648])|((m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&m[1238]))):InitCond[1347];
    m[1241] = run?((((m[1238]&~m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&~m[1243])|(~m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&m[1242]&m[1243]))&UnbiasedRNG[649])|((m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&m[1243]))):InitCond[1348];
    m[1251] = run?((((m[1248]&~m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&~m[1253])|(~m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&m[1252]&m[1253]))&UnbiasedRNG[650])|((m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&m[1253]))):InitCond[1349];
    m[1256] = run?((((m[1253]&~m[1254]&~m[1255]&~m[1257]&~m[1258])|(~m[1253]&m[1254]&~m[1255]&~m[1257]&~m[1258])|(~m[1253]&~m[1254]&m[1255]&~m[1257]&~m[1258])|(m[1253]&m[1254]&m[1255]&m[1257]&~m[1258])|(~m[1253]&~m[1254]&~m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&~m[1255]&m[1257]&m[1258])|(m[1253]&~m[1254]&m[1255]&m[1257]&m[1258])|(~m[1253]&m[1254]&m[1255]&m[1257]&m[1258]))&UnbiasedRNG[651])|((m[1253]&m[1254]&~m[1255]&~m[1257]&~m[1258])|(m[1253]&~m[1254]&m[1255]&~m[1257]&~m[1258])|(~m[1253]&m[1254]&m[1255]&~m[1257]&~m[1258])|(m[1253]&m[1254]&m[1255]&~m[1257]&~m[1258])|(m[1253]&~m[1254]&~m[1255]&~m[1257]&m[1258])|(~m[1253]&m[1254]&~m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&~m[1255]&~m[1257]&m[1258])|(~m[1253]&~m[1254]&m[1255]&~m[1257]&m[1258])|(m[1253]&~m[1254]&m[1255]&~m[1257]&m[1258])|(~m[1253]&m[1254]&m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&m[1255]&m[1257]&m[1258]))):InitCond[1350];
    m[1261] = run?((((m[1258]&~m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&~m[1263])|(~m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&m[1262]&m[1263]))&UnbiasedRNG[652])|((m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&m[1263]))):InitCond[1351];
    m[1266] = run?((((m[1263]&~m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&~m[1268])|(~m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&m[1267]&m[1268]))&UnbiasedRNG[653])|((m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&m[1268]))):InitCond[1352];
    m[1271] = run?((((m[1268]&~m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&~m[1273])|(~m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&m[1272]&m[1273]))&UnbiasedRNG[654])|((m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&m[1273]))):InitCond[1353];
    m[1276] = run?((((m[1273]&~m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&~m[1278])|(~m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&m[1277]&m[1278]))&UnbiasedRNG[655])|((m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&m[1278]))):InitCond[1354];
    m[1281] = run?((((m[1278]&~m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&~m[1283])|(~m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&m[1282]&m[1283]))&UnbiasedRNG[656])|((m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&m[1283]))):InitCond[1355];
    m[1286] = run?((((m[1283]&~m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&~m[1288])|(~m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&m[1287]&m[1288]))&UnbiasedRNG[657])|((m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&m[1288]))):InitCond[1356];
    m[1291] = run?((((m[1288]&~m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&~m[1293])|(~m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&m[1292]&m[1293]))&UnbiasedRNG[658])|((m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&m[1293]))):InitCond[1357];
    m[1296] = run?((((m[1293]&~m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&~m[1298])|(~m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&m[1297]&m[1298]))&UnbiasedRNG[659])|((m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&m[1298]))):InitCond[1358];
    m[1301] = run?((((m[1298]&~m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&~m[1303])|(~m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&m[1302]&m[1303]))&UnbiasedRNG[660])|((m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&m[1303]))):InitCond[1359];
    m[1311] = run?((((m[1308]&~m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&~m[1313])|(~m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&m[1312]&m[1313]))&UnbiasedRNG[661])|((m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&m[1313]))):InitCond[1360];
    m[1316] = run?((((m[1313]&~m[1314]&~m[1315]&~m[1317]&~m[1318])|(~m[1313]&m[1314]&~m[1315]&~m[1317]&~m[1318])|(~m[1313]&~m[1314]&m[1315]&~m[1317]&~m[1318])|(m[1313]&m[1314]&m[1315]&m[1317]&~m[1318])|(~m[1313]&~m[1314]&~m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&~m[1315]&m[1317]&m[1318])|(m[1313]&~m[1314]&m[1315]&m[1317]&m[1318])|(~m[1313]&m[1314]&m[1315]&m[1317]&m[1318]))&UnbiasedRNG[662])|((m[1313]&m[1314]&~m[1315]&~m[1317]&~m[1318])|(m[1313]&~m[1314]&m[1315]&~m[1317]&~m[1318])|(~m[1313]&m[1314]&m[1315]&~m[1317]&~m[1318])|(m[1313]&m[1314]&m[1315]&~m[1317]&~m[1318])|(m[1313]&~m[1314]&~m[1315]&~m[1317]&m[1318])|(~m[1313]&m[1314]&~m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&~m[1315]&~m[1317]&m[1318])|(~m[1313]&~m[1314]&m[1315]&~m[1317]&m[1318])|(m[1313]&~m[1314]&m[1315]&~m[1317]&m[1318])|(~m[1313]&m[1314]&m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&m[1315]&m[1317]&m[1318]))):InitCond[1361];
    m[1321] = run?((((m[1318]&~m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&~m[1323])|(~m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&m[1322]&m[1323]))&UnbiasedRNG[663])|((m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&m[1323]))):InitCond[1362];
    m[1326] = run?((((m[1323]&~m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&~m[1328])|(~m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&m[1327]&m[1328]))&UnbiasedRNG[664])|((m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&m[1328]))):InitCond[1363];
    m[1331] = run?((((m[1328]&~m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&~m[1333])|(~m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&m[1332]&m[1333]))&UnbiasedRNG[665])|((m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&m[1333]))):InitCond[1364];
    m[1336] = run?((((m[1333]&~m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&~m[1338])|(~m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&m[1337]&m[1338]))&UnbiasedRNG[666])|((m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&m[1338]))):InitCond[1365];
    m[1341] = run?((((m[1338]&~m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&~m[1343])|(~m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&m[1342]&m[1343]))&UnbiasedRNG[667])|((m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&m[1343]))):InitCond[1366];
    m[1346] = run?((((m[1343]&~m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&~m[1348])|(~m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&m[1347]&m[1348]))&UnbiasedRNG[668])|((m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&m[1348]))):InitCond[1367];
    m[1351] = run?((((m[1348]&~m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&~m[1353])|(~m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&m[1352]&m[1353]))&UnbiasedRNG[669])|((m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&m[1353]))):InitCond[1368];
    m[1356] = run?((((m[1353]&~m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&~m[1358])|(~m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&m[1357]&m[1358]))&UnbiasedRNG[670])|((m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&m[1358]))):InitCond[1369];
    m[1366] = run?((((m[1363]&~m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&~m[1368])|(~m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&m[1367]&m[1368]))&UnbiasedRNG[671])|((m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&m[1368]))):InitCond[1370];
    m[1371] = run?((((m[1368]&~m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&~m[1373])|(~m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&m[1372]&m[1373]))&UnbiasedRNG[672])|((m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&m[1373]))):InitCond[1371];
    m[1376] = run?((((m[1373]&~m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&~m[1378])|(~m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&m[1377]&m[1378]))&UnbiasedRNG[673])|((m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&m[1378]))):InitCond[1372];
    m[1381] = run?((((m[1378]&~m[1379]&~m[1380]&~m[1382]&~m[1383])|(~m[1378]&m[1379]&~m[1380]&~m[1382]&~m[1383])|(~m[1378]&~m[1379]&m[1380]&~m[1382]&~m[1383])|(m[1378]&m[1379]&m[1380]&m[1382]&~m[1383])|(~m[1378]&~m[1379]&~m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&~m[1380]&m[1382]&m[1383])|(m[1378]&~m[1379]&m[1380]&m[1382]&m[1383])|(~m[1378]&m[1379]&m[1380]&m[1382]&m[1383]))&UnbiasedRNG[674])|((m[1378]&m[1379]&~m[1380]&~m[1382]&~m[1383])|(m[1378]&~m[1379]&m[1380]&~m[1382]&~m[1383])|(~m[1378]&m[1379]&m[1380]&~m[1382]&~m[1383])|(m[1378]&m[1379]&m[1380]&~m[1382]&~m[1383])|(m[1378]&~m[1379]&~m[1380]&~m[1382]&m[1383])|(~m[1378]&m[1379]&~m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&~m[1380]&~m[1382]&m[1383])|(~m[1378]&~m[1379]&m[1380]&~m[1382]&m[1383])|(m[1378]&~m[1379]&m[1380]&~m[1382]&m[1383])|(~m[1378]&m[1379]&m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&m[1380]&m[1382]&m[1383]))):InitCond[1373];
    m[1386] = run?((((m[1383]&~m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&~m[1388])|(~m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&m[1387]&m[1388]))&UnbiasedRNG[675])|((m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&m[1388]))):InitCond[1374];
    m[1391] = run?((((m[1388]&~m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&~m[1393])|(~m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&m[1392]&m[1393]))&UnbiasedRNG[676])|((m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&m[1393]))):InitCond[1375];
    m[1396] = run?((((m[1393]&~m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&~m[1398])|(~m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&m[1397]&m[1398]))&UnbiasedRNG[677])|((m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&m[1398]))):InitCond[1376];
    m[1401] = run?((((m[1398]&~m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&~m[1403])|(~m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&m[1402]&m[1403]))&UnbiasedRNG[678])|((m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&m[1403]))):InitCond[1377];
    m[1406] = run?((((m[1403]&~m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&~m[1408])|(~m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&m[1407]&m[1408]))&UnbiasedRNG[679])|((m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&m[1408]))):InitCond[1378];
    m[1416] = run?((((m[1413]&~m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&~m[1418])|(~m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&m[1417]&m[1418]))&UnbiasedRNG[680])|((m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&m[1418]))):InitCond[1379];
    m[1421] = run?((((m[1418]&~m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&~m[1423])|(~m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&m[1422]&m[1423]))&UnbiasedRNG[681])|((m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&m[1423]))):InitCond[1380];
    m[1426] = run?((((m[1423]&~m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&~m[1428])|(~m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&m[1427]&m[1428]))&UnbiasedRNG[682])|((m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&m[1428]))):InitCond[1381];
    m[1431] = run?((((m[1428]&~m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&~m[1433])|(~m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&m[1432]&m[1433]))&UnbiasedRNG[683])|((m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&m[1433]))):InitCond[1382];
    m[1436] = run?((((m[1433]&~m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&~m[1438])|(~m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&m[1437]&m[1438]))&UnbiasedRNG[684])|((m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&m[1438]))):InitCond[1383];
    m[1441] = run?((((m[1438]&~m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&~m[1443])|(~m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&m[1442]&m[1443]))&UnbiasedRNG[685])|((m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&m[1443]))):InitCond[1384];
    m[1446] = run?((((m[1443]&~m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&~m[1448])|(~m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&m[1447]&m[1448]))&UnbiasedRNG[686])|((m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&m[1448]))):InitCond[1385];
    m[1451] = run?((((m[1448]&~m[1449]&~m[1450]&~m[1452]&~m[1453])|(~m[1448]&m[1449]&~m[1450]&~m[1452]&~m[1453])|(~m[1448]&~m[1449]&m[1450]&~m[1452]&~m[1453])|(m[1448]&m[1449]&m[1450]&m[1452]&~m[1453])|(~m[1448]&~m[1449]&~m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&~m[1450]&m[1452]&m[1453])|(m[1448]&~m[1449]&m[1450]&m[1452]&m[1453])|(~m[1448]&m[1449]&m[1450]&m[1452]&m[1453]))&UnbiasedRNG[687])|((m[1448]&m[1449]&~m[1450]&~m[1452]&~m[1453])|(m[1448]&~m[1449]&m[1450]&~m[1452]&~m[1453])|(~m[1448]&m[1449]&m[1450]&~m[1452]&~m[1453])|(m[1448]&m[1449]&m[1450]&~m[1452]&~m[1453])|(m[1448]&~m[1449]&~m[1450]&~m[1452]&m[1453])|(~m[1448]&m[1449]&~m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&~m[1450]&~m[1452]&m[1453])|(~m[1448]&~m[1449]&m[1450]&~m[1452]&m[1453])|(m[1448]&~m[1449]&m[1450]&~m[1452]&m[1453])|(~m[1448]&m[1449]&m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&m[1450]&m[1452]&m[1453]))):InitCond[1386];
    m[1461] = run?((((m[1458]&~m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&~m[1463])|(~m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&m[1462]&m[1463]))&UnbiasedRNG[688])|((m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&m[1463]))):InitCond[1387];
    m[1466] = run?((((m[1463]&~m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&~m[1468])|(~m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&m[1467]&m[1468]))&UnbiasedRNG[689])|((m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&m[1468]))):InitCond[1388];
    m[1471] = run?((((m[1468]&~m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&~m[1473])|(~m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&m[1472]&m[1473]))&UnbiasedRNG[690])|((m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&m[1473]))):InitCond[1389];
    m[1476] = run?((((m[1473]&~m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&~m[1478])|(~m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&m[1477]&m[1478]))&UnbiasedRNG[691])|((m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&m[1478]))):InitCond[1390];
    m[1481] = run?((((m[1478]&~m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&~m[1483])|(~m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&m[1482]&m[1483]))&UnbiasedRNG[692])|((m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&m[1483]))):InitCond[1391];
    m[1486] = run?((((m[1483]&~m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&~m[1488])|(~m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&m[1487]&m[1488]))&UnbiasedRNG[693])|((m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&m[1488]))):InitCond[1392];
    m[1491] = run?((((m[1488]&~m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&~m[1493])|(~m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&m[1492]&m[1493]))&UnbiasedRNG[694])|((m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&m[1493]))):InitCond[1393];
    m[1501] = run?((((m[1498]&~m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&~m[1503])|(~m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&m[1502]&m[1503]))&UnbiasedRNG[695])|((m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&m[1503]))):InitCond[1394];
    m[1506] = run?((((m[1503]&~m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&~m[1508])|(~m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&m[1507]&m[1508]))&UnbiasedRNG[696])|((m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&m[1508]))):InitCond[1395];
    m[1511] = run?((((m[1508]&~m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&~m[1513])|(~m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&m[1512]&m[1513]))&UnbiasedRNG[697])|((m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&m[1513]))):InitCond[1396];
    m[1516] = run?((((m[1513]&~m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&~m[1518])|(~m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&m[1517]&m[1518]))&UnbiasedRNG[698])|((m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&m[1518]))):InitCond[1397];
    m[1521] = run?((((m[1518]&~m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&~m[1523])|(~m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&m[1522]&m[1523]))&UnbiasedRNG[699])|((m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&m[1523]))):InitCond[1398];
    m[1526] = run?((((m[1523]&~m[1524]&~m[1525]&~m[1527]&~m[1528])|(~m[1523]&m[1524]&~m[1525]&~m[1527]&~m[1528])|(~m[1523]&~m[1524]&m[1525]&~m[1527]&~m[1528])|(m[1523]&m[1524]&m[1525]&m[1527]&~m[1528])|(~m[1523]&~m[1524]&~m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&~m[1525]&m[1527]&m[1528])|(m[1523]&~m[1524]&m[1525]&m[1527]&m[1528])|(~m[1523]&m[1524]&m[1525]&m[1527]&m[1528]))&UnbiasedRNG[700])|((m[1523]&m[1524]&~m[1525]&~m[1527]&~m[1528])|(m[1523]&~m[1524]&m[1525]&~m[1527]&~m[1528])|(~m[1523]&m[1524]&m[1525]&~m[1527]&~m[1528])|(m[1523]&m[1524]&m[1525]&~m[1527]&~m[1528])|(m[1523]&~m[1524]&~m[1525]&~m[1527]&m[1528])|(~m[1523]&m[1524]&~m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&~m[1525]&~m[1527]&m[1528])|(~m[1523]&~m[1524]&m[1525]&~m[1527]&m[1528])|(m[1523]&~m[1524]&m[1525]&~m[1527]&m[1528])|(~m[1523]&m[1524]&m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&m[1525]&m[1527]&m[1528]))):InitCond[1399];
    m[1536] = run?((((m[1533]&~m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&~m[1538])|(~m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&m[1537]&m[1538]))&UnbiasedRNG[701])|((m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&m[1538]))):InitCond[1400];
    m[1541] = run?((((m[1538]&~m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&~m[1543])|(~m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&m[1542]&m[1543]))&UnbiasedRNG[702])|((m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&m[1543]))):InitCond[1401];
    m[1546] = run?((((m[1543]&~m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&~m[1548])|(~m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&m[1547]&m[1548]))&UnbiasedRNG[703])|((m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&m[1548]))):InitCond[1402];
    m[1551] = run?((((m[1548]&~m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&~m[1553])|(~m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&m[1552]&m[1553]))&UnbiasedRNG[704])|((m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&m[1553]))):InitCond[1403];
    m[1556] = run?((((m[1553]&~m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&~m[1558])|(~m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&m[1557]&m[1558]))&UnbiasedRNG[705])|((m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&m[1558]))):InitCond[1404];
    m[1566] = run?((((m[1563]&~m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&~m[1568])|(~m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&m[1567]&m[1568]))&UnbiasedRNG[706])|((m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&m[1568]))):InitCond[1405];
    m[1571] = run?((((m[1568]&~m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&~m[1573])|(~m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&m[1572]&m[1573]))&UnbiasedRNG[707])|((m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&m[1573]))):InitCond[1406];
    m[1576] = run?((((m[1573]&~m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&~m[1578])|(~m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&m[1577]&m[1578]))&UnbiasedRNG[708])|((m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&m[1578]))):InitCond[1407];
    m[1581] = run?((((m[1578]&~m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&~m[1583])|(~m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&m[1582]&m[1583]))&UnbiasedRNG[709])|((m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&m[1583]))):InitCond[1408];
    m[1591] = run?((((m[1588]&~m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&~m[1593])|(~m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&m[1592]&m[1593]))&UnbiasedRNG[710])|((m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&m[1593]))):InitCond[1409];
    m[1596] = run?((((m[1593]&~m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&~m[1598])|(~m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&m[1597]&m[1598]))&UnbiasedRNG[711])|((m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&m[1598]))):InitCond[1410];
    m[1601] = run?((((m[1598]&~m[1599]&~m[1600]&~m[1602]&~m[1603])|(~m[1598]&m[1599]&~m[1600]&~m[1602]&~m[1603])|(~m[1598]&~m[1599]&m[1600]&~m[1602]&~m[1603])|(m[1598]&m[1599]&m[1600]&m[1602]&~m[1603])|(~m[1598]&~m[1599]&~m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&~m[1600]&m[1602]&m[1603])|(m[1598]&~m[1599]&m[1600]&m[1602]&m[1603])|(~m[1598]&m[1599]&m[1600]&m[1602]&m[1603]))&UnbiasedRNG[712])|((m[1598]&m[1599]&~m[1600]&~m[1602]&~m[1603])|(m[1598]&~m[1599]&m[1600]&~m[1602]&~m[1603])|(~m[1598]&m[1599]&m[1600]&~m[1602]&~m[1603])|(m[1598]&m[1599]&m[1600]&~m[1602]&~m[1603])|(m[1598]&~m[1599]&~m[1600]&~m[1602]&m[1603])|(~m[1598]&m[1599]&~m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&~m[1600]&~m[1602]&m[1603])|(~m[1598]&~m[1599]&m[1600]&~m[1602]&m[1603])|(m[1598]&~m[1599]&m[1600]&~m[1602]&m[1603])|(~m[1598]&m[1599]&m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&m[1600]&m[1602]&m[1603]))):InitCond[1411];
    m[1611] = run?((((m[1608]&~m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&~m[1613])|(~m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&m[1612]&m[1613]))&UnbiasedRNG[713])|((m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&m[1613]))):InitCond[1412];
    m[1616] = run?((((m[1613]&~m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&~m[1618])|(~m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&m[1617]&m[1618]))&UnbiasedRNG[714])|((m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&m[1618]))):InitCond[1413];
    m[1626] = run?((((m[1623]&~m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&~m[1628])|(~m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&m[1627]&m[1628]))&UnbiasedRNG[715])|((m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&m[1628]))):InitCond[1414];
end

always @(posedge color4_clk) begin
    m[732] = run?((((m[728]&~m[729]&~m[730]&~m[731]&~m[735])|(~m[728]&m[729]&~m[730]&~m[731]&~m[735])|(~m[728]&~m[729]&m[730]&~m[731]&~m[735])|(m[728]&m[729]&~m[730]&m[731]&~m[735])|(m[728]&~m[729]&m[730]&m[731]&~m[735])|(~m[728]&m[729]&m[730]&m[731]&~m[735]))&BiasedRNG[699])|(((m[728]&~m[729]&~m[730]&~m[731]&m[735])|(~m[728]&m[729]&~m[730]&~m[731]&m[735])|(~m[728]&~m[729]&m[730]&~m[731]&m[735])|(m[728]&m[729]&~m[730]&m[731]&m[735])|(m[728]&~m[729]&m[730]&m[731]&m[735])|(~m[728]&m[729]&m[730]&m[731]&m[735]))&~BiasedRNG[699])|((m[728]&m[729]&~m[730]&~m[731]&~m[735])|(m[728]&~m[729]&m[730]&~m[731]&~m[735])|(~m[728]&m[729]&m[730]&~m[731]&~m[735])|(m[728]&m[729]&m[730]&~m[731]&~m[735])|(m[728]&m[729]&m[730]&m[731]&~m[735])|(m[728]&m[729]&~m[730]&~m[731]&m[735])|(m[728]&~m[729]&m[730]&~m[731]&m[735])|(~m[728]&m[729]&m[730]&~m[731]&m[735])|(m[728]&m[729]&m[730]&~m[731]&m[735])|(m[728]&m[729]&m[730]&m[731]&m[735]))):InitCond[1415];
    m[737] = run?((((m[733]&~m[734]&~m[735]&~m[736]&~m[745])|(~m[733]&m[734]&~m[735]&~m[736]&~m[745])|(~m[733]&~m[734]&m[735]&~m[736]&~m[745])|(m[733]&m[734]&~m[735]&m[736]&~m[745])|(m[733]&~m[734]&m[735]&m[736]&~m[745])|(~m[733]&m[734]&m[735]&m[736]&~m[745]))&BiasedRNG[700])|(((m[733]&~m[734]&~m[735]&~m[736]&m[745])|(~m[733]&m[734]&~m[735]&~m[736]&m[745])|(~m[733]&~m[734]&m[735]&~m[736]&m[745])|(m[733]&m[734]&~m[735]&m[736]&m[745])|(m[733]&~m[734]&m[735]&m[736]&m[745])|(~m[733]&m[734]&m[735]&m[736]&m[745]))&~BiasedRNG[700])|((m[733]&m[734]&~m[735]&~m[736]&~m[745])|(m[733]&~m[734]&m[735]&~m[736]&~m[745])|(~m[733]&m[734]&m[735]&~m[736]&~m[745])|(m[733]&m[734]&m[735]&~m[736]&~m[745])|(m[733]&m[734]&m[735]&m[736]&~m[745])|(m[733]&m[734]&~m[735]&~m[736]&m[745])|(m[733]&~m[734]&m[735]&~m[736]&m[745])|(~m[733]&m[734]&m[735]&~m[736]&m[745])|(m[733]&m[734]&m[735]&~m[736]&m[745])|(m[733]&m[734]&m[735]&m[736]&m[745]))):InitCond[1416];
    m[742] = run?((((m[738]&~m[739]&~m[740]&~m[741]&~m[750])|(~m[738]&m[739]&~m[740]&~m[741]&~m[750])|(~m[738]&~m[739]&m[740]&~m[741]&~m[750])|(m[738]&m[739]&~m[740]&m[741]&~m[750])|(m[738]&~m[739]&m[740]&m[741]&~m[750])|(~m[738]&m[739]&m[740]&m[741]&~m[750]))&BiasedRNG[701])|(((m[738]&~m[739]&~m[740]&~m[741]&m[750])|(~m[738]&m[739]&~m[740]&~m[741]&m[750])|(~m[738]&~m[739]&m[740]&~m[741]&m[750])|(m[738]&m[739]&~m[740]&m[741]&m[750])|(m[738]&~m[739]&m[740]&m[741]&m[750])|(~m[738]&m[739]&m[740]&m[741]&m[750]))&~BiasedRNG[701])|((m[738]&m[739]&~m[740]&~m[741]&~m[750])|(m[738]&~m[739]&m[740]&~m[741]&~m[750])|(~m[738]&m[739]&m[740]&~m[741]&~m[750])|(m[738]&m[739]&m[740]&~m[741]&~m[750])|(m[738]&m[739]&m[740]&m[741]&~m[750])|(m[738]&m[739]&~m[740]&~m[741]&m[750])|(m[738]&~m[739]&m[740]&~m[741]&m[750])|(~m[738]&m[739]&m[740]&~m[741]&m[750])|(m[738]&m[739]&m[740]&~m[741]&m[750])|(m[738]&m[739]&m[740]&m[741]&m[750]))):InitCond[1417];
    m[747] = run?((((m[743]&~m[744]&~m[745]&~m[746]&~m[760])|(~m[743]&m[744]&~m[745]&~m[746]&~m[760])|(~m[743]&~m[744]&m[745]&~m[746]&~m[760])|(m[743]&m[744]&~m[745]&m[746]&~m[760])|(m[743]&~m[744]&m[745]&m[746]&~m[760])|(~m[743]&m[744]&m[745]&m[746]&~m[760]))&BiasedRNG[702])|(((m[743]&~m[744]&~m[745]&~m[746]&m[760])|(~m[743]&m[744]&~m[745]&~m[746]&m[760])|(~m[743]&~m[744]&m[745]&~m[746]&m[760])|(m[743]&m[744]&~m[745]&m[746]&m[760])|(m[743]&~m[744]&m[745]&m[746]&m[760])|(~m[743]&m[744]&m[745]&m[746]&m[760]))&~BiasedRNG[702])|((m[743]&m[744]&~m[745]&~m[746]&~m[760])|(m[743]&~m[744]&m[745]&~m[746]&~m[760])|(~m[743]&m[744]&m[745]&~m[746]&~m[760])|(m[743]&m[744]&m[745]&~m[746]&~m[760])|(m[743]&m[744]&m[745]&m[746]&~m[760])|(m[743]&m[744]&~m[745]&~m[746]&m[760])|(m[743]&~m[744]&m[745]&~m[746]&m[760])|(~m[743]&m[744]&m[745]&~m[746]&m[760])|(m[743]&m[744]&m[745]&~m[746]&m[760])|(m[743]&m[744]&m[745]&m[746]&m[760]))):InitCond[1418];
    m[752] = run?((((m[748]&~m[749]&~m[750]&~m[751]&~m[765])|(~m[748]&m[749]&~m[750]&~m[751]&~m[765])|(~m[748]&~m[749]&m[750]&~m[751]&~m[765])|(m[748]&m[749]&~m[750]&m[751]&~m[765])|(m[748]&~m[749]&m[750]&m[751]&~m[765])|(~m[748]&m[749]&m[750]&m[751]&~m[765]))&BiasedRNG[703])|(((m[748]&~m[749]&~m[750]&~m[751]&m[765])|(~m[748]&m[749]&~m[750]&~m[751]&m[765])|(~m[748]&~m[749]&m[750]&~m[751]&m[765])|(m[748]&m[749]&~m[750]&m[751]&m[765])|(m[748]&~m[749]&m[750]&m[751]&m[765])|(~m[748]&m[749]&m[750]&m[751]&m[765]))&~BiasedRNG[703])|((m[748]&m[749]&~m[750]&~m[751]&~m[765])|(m[748]&~m[749]&m[750]&~m[751]&~m[765])|(~m[748]&m[749]&m[750]&~m[751]&~m[765])|(m[748]&m[749]&m[750]&~m[751]&~m[765])|(m[748]&m[749]&m[750]&m[751]&~m[765])|(m[748]&m[749]&~m[750]&~m[751]&m[765])|(m[748]&~m[749]&m[750]&~m[751]&m[765])|(~m[748]&m[749]&m[750]&~m[751]&m[765])|(m[748]&m[749]&m[750]&~m[751]&m[765])|(m[748]&m[749]&m[750]&m[751]&m[765]))):InitCond[1419];
    m[757] = run?((((m[753]&~m[754]&~m[755]&~m[756]&~m[770])|(~m[753]&m[754]&~m[755]&~m[756]&~m[770])|(~m[753]&~m[754]&m[755]&~m[756]&~m[770])|(m[753]&m[754]&~m[755]&m[756]&~m[770])|(m[753]&~m[754]&m[755]&m[756]&~m[770])|(~m[753]&m[754]&m[755]&m[756]&~m[770]))&BiasedRNG[704])|(((m[753]&~m[754]&~m[755]&~m[756]&m[770])|(~m[753]&m[754]&~m[755]&~m[756]&m[770])|(~m[753]&~m[754]&m[755]&~m[756]&m[770])|(m[753]&m[754]&~m[755]&m[756]&m[770])|(m[753]&~m[754]&m[755]&m[756]&m[770])|(~m[753]&m[754]&m[755]&m[756]&m[770]))&~BiasedRNG[704])|((m[753]&m[754]&~m[755]&~m[756]&~m[770])|(m[753]&~m[754]&m[755]&~m[756]&~m[770])|(~m[753]&m[754]&m[755]&~m[756]&~m[770])|(m[753]&m[754]&m[755]&~m[756]&~m[770])|(m[753]&m[754]&m[755]&m[756]&~m[770])|(m[753]&m[754]&~m[755]&~m[756]&m[770])|(m[753]&~m[754]&m[755]&~m[756]&m[770])|(~m[753]&m[754]&m[755]&~m[756]&m[770])|(m[753]&m[754]&m[755]&~m[756]&m[770])|(m[753]&m[754]&m[755]&m[756]&m[770]))):InitCond[1420];
    m[762] = run?((((m[758]&~m[759]&~m[760]&~m[761]&~m[780])|(~m[758]&m[759]&~m[760]&~m[761]&~m[780])|(~m[758]&~m[759]&m[760]&~m[761]&~m[780])|(m[758]&m[759]&~m[760]&m[761]&~m[780])|(m[758]&~m[759]&m[760]&m[761]&~m[780])|(~m[758]&m[759]&m[760]&m[761]&~m[780]))&BiasedRNG[705])|(((m[758]&~m[759]&~m[760]&~m[761]&m[780])|(~m[758]&m[759]&~m[760]&~m[761]&m[780])|(~m[758]&~m[759]&m[760]&~m[761]&m[780])|(m[758]&m[759]&~m[760]&m[761]&m[780])|(m[758]&~m[759]&m[760]&m[761]&m[780])|(~m[758]&m[759]&m[760]&m[761]&m[780]))&~BiasedRNG[705])|((m[758]&m[759]&~m[760]&~m[761]&~m[780])|(m[758]&~m[759]&m[760]&~m[761]&~m[780])|(~m[758]&m[759]&m[760]&~m[761]&~m[780])|(m[758]&m[759]&m[760]&~m[761]&~m[780])|(m[758]&m[759]&m[760]&m[761]&~m[780])|(m[758]&m[759]&~m[760]&~m[761]&m[780])|(m[758]&~m[759]&m[760]&~m[761]&m[780])|(~m[758]&m[759]&m[760]&~m[761]&m[780])|(m[758]&m[759]&m[760]&~m[761]&m[780])|(m[758]&m[759]&m[760]&m[761]&m[780]))):InitCond[1421];
    m[767] = run?((((m[763]&~m[764]&~m[765]&~m[766]&~m[785])|(~m[763]&m[764]&~m[765]&~m[766]&~m[785])|(~m[763]&~m[764]&m[765]&~m[766]&~m[785])|(m[763]&m[764]&~m[765]&m[766]&~m[785])|(m[763]&~m[764]&m[765]&m[766]&~m[785])|(~m[763]&m[764]&m[765]&m[766]&~m[785]))&BiasedRNG[706])|(((m[763]&~m[764]&~m[765]&~m[766]&m[785])|(~m[763]&m[764]&~m[765]&~m[766]&m[785])|(~m[763]&~m[764]&m[765]&~m[766]&m[785])|(m[763]&m[764]&~m[765]&m[766]&m[785])|(m[763]&~m[764]&m[765]&m[766]&m[785])|(~m[763]&m[764]&m[765]&m[766]&m[785]))&~BiasedRNG[706])|((m[763]&m[764]&~m[765]&~m[766]&~m[785])|(m[763]&~m[764]&m[765]&~m[766]&~m[785])|(~m[763]&m[764]&m[765]&~m[766]&~m[785])|(m[763]&m[764]&m[765]&~m[766]&~m[785])|(m[763]&m[764]&m[765]&m[766]&~m[785])|(m[763]&m[764]&~m[765]&~m[766]&m[785])|(m[763]&~m[764]&m[765]&~m[766]&m[785])|(~m[763]&m[764]&m[765]&~m[766]&m[785])|(m[763]&m[764]&m[765]&~m[766]&m[785])|(m[763]&m[764]&m[765]&m[766]&m[785]))):InitCond[1422];
    m[772] = run?((((m[768]&~m[769]&~m[770]&~m[771]&~m[790])|(~m[768]&m[769]&~m[770]&~m[771]&~m[790])|(~m[768]&~m[769]&m[770]&~m[771]&~m[790])|(m[768]&m[769]&~m[770]&m[771]&~m[790])|(m[768]&~m[769]&m[770]&m[771]&~m[790])|(~m[768]&m[769]&m[770]&m[771]&~m[790]))&BiasedRNG[707])|(((m[768]&~m[769]&~m[770]&~m[771]&m[790])|(~m[768]&m[769]&~m[770]&~m[771]&m[790])|(~m[768]&~m[769]&m[770]&~m[771]&m[790])|(m[768]&m[769]&~m[770]&m[771]&m[790])|(m[768]&~m[769]&m[770]&m[771]&m[790])|(~m[768]&m[769]&m[770]&m[771]&m[790]))&~BiasedRNG[707])|((m[768]&m[769]&~m[770]&~m[771]&~m[790])|(m[768]&~m[769]&m[770]&~m[771]&~m[790])|(~m[768]&m[769]&m[770]&~m[771]&~m[790])|(m[768]&m[769]&m[770]&~m[771]&~m[790])|(m[768]&m[769]&m[770]&m[771]&~m[790])|(m[768]&m[769]&~m[770]&~m[771]&m[790])|(m[768]&~m[769]&m[770]&~m[771]&m[790])|(~m[768]&m[769]&m[770]&~m[771]&m[790])|(m[768]&m[769]&m[770]&~m[771]&m[790])|(m[768]&m[769]&m[770]&m[771]&m[790]))):InitCond[1423];
    m[777] = run?((((m[773]&~m[774]&~m[775]&~m[776]&~m[795])|(~m[773]&m[774]&~m[775]&~m[776]&~m[795])|(~m[773]&~m[774]&m[775]&~m[776]&~m[795])|(m[773]&m[774]&~m[775]&m[776]&~m[795])|(m[773]&~m[774]&m[775]&m[776]&~m[795])|(~m[773]&m[774]&m[775]&m[776]&~m[795]))&BiasedRNG[708])|(((m[773]&~m[774]&~m[775]&~m[776]&m[795])|(~m[773]&m[774]&~m[775]&~m[776]&m[795])|(~m[773]&~m[774]&m[775]&~m[776]&m[795])|(m[773]&m[774]&~m[775]&m[776]&m[795])|(m[773]&~m[774]&m[775]&m[776]&m[795])|(~m[773]&m[774]&m[775]&m[776]&m[795]))&~BiasedRNG[708])|((m[773]&m[774]&~m[775]&~m[776]&~m[795])|(m[773]&~m[774]&m[775]&~m[776]&~m[795])|(~m[773]&m[774]&m[775]&~m[776]&~m[795])|(m[773]&m[774]&m[775]&~m[776]&~m[795])|(m[773]&m[774]&m[775]&m[776]&~m[795])|(m[773]&m[774]&~m[775]&~m[776]&m[795])|(m[773]&~m[774]&m[775]&~m[776]&m[795])|(~m[773]&m[774]&m[775]&~m[776]&m[795])|(m[773]&m[774]&m[775]&~m[776]&m[795])|(m[773]&m[774]&m[775]&m[776]&m[795]))):InitCond[1424];
    m[782] = run?((((m[778]&~m[779]&~m[780]&~m[781]&~m[805])|(~m[778]&m[779]&~m[780]&~m[781]&~m[805])|(~m[778]&~m[779]&m[780]&~m[781]&~m[805])|(m[778]&m[779]&~m[780]&m[781]&~m[805])|(m[778]&~m[779]&m[780]&m[781]&~m[805])|(~m[778]&m[779]&m[780]&m[781]&~m[805]))&BiasedRNG[709])|(((m[778]&~m[779]&~m[780]&~m[781]&m[805])|(~m[778]&m[779]&~m[780]&~m[781]&m[805])|(~m[778]&~m[779]&m[780]&~m[781]&m[805])|(m[778]&m[779]&~m[780]&m[781]&m[805])|(m[778]&~m[779]&m[780]&m[781]&m[805])|(~m[778]&m[779]&m[780]&m[781]&m[805]))&~BiasedRNG[709])|((m[778]&m[779]&~m[780]&~m[781]&~m[805])|(m[778]&~m[779]&m[780]&~m[781]&~m[805])|(~m[778]&m[779]&m[780]&~m[781]&~m[805])|(m[778]&m[779]&m[780]&~m[781]&~m[805])|(m[778]&m[779]&m[780]&m[781]&~m[805])|(m[778]&m[779]&~m[780]&~m[781]&m[805])|(m[778]&~m[779]&m[780]&~m[781]&m[805])|(~m[778]&m[779]&m[780]&~m[781]&m[805])|(m[778]&m[779]&m[780]&~m[781]&m[805])|(m[778]&m[779]&m[780]&m[781]&m[805]))):InitCond[1425];
    m[787] = run?((((m[783]&~m[784]&~m[785]&~m[786]&~m[810])|(~m[783]&m[784]&~m[785]&~m[786]&~m[810])|(~m[783]&~m[784]&m[785]&~m[786]&~m[810])|(m[783]&m[784]&~m[785]&m[786]&~m[810])|(m[783]&~m[784]&m[785]&m[786]&~m[810])|(~m[783]&m[784]&m[785]&m[786]&~m[810]))&BiasedRNG[710])|(((m[783]&~m[784]&~m[785]&~m[786]&m[810])|(~m[783]&m[784]&~m[785]&~m[786]&m[810])|(~m[783]&~m[784]&m[785]&~m[786]&m[810])|(m[783]&m[784]&~m[785]&m[786]&m[810])|(m[783]&~m[784]&m[785]&m[786]&m[810])|(~m[783]&m[784]&m[785]&m[786]&m[810]))&~BiasedRNG[710])|((m[783]&m[784]&~m[785]&~m[786]&~m[810])|(m[783]&~m[784]&m[785]&~m[786]&~m[810])|(~m[783]&m[784]&m[785]&~m[786]&~m[810])|(m[783]&m[784]&m[785]&~m[786]&~m[810])|(m[783]&m[784]&m[785]&m[786]&~m[810])|(m[783]&m[784]&~m[785]&~m[786]&m[810])|(m[783]&~m[784]&m[785]&~m[786]&m[810])|(~m[783]&m[784]&m[785]&~m[786]&m[810])|(m[783]&m[784]&m[785]&~m[786]&m[810])|(m[783]&m[784]&m[785]&m[786]&m[810]))):InitCond[1426];
    m[792] = run?((((m[788]&~m[789]&~m[790]&~m[791]&~m[815])|(~m[788]&m[789]&~m[790]&~m[791]&~m[815])|(~m[788]&~m[789]&m[790]&~m[791]&~m[815])|(m[788]&m[789]&~m[790]&m[791]&~m[815])|(m[788]&~m[789]&m[790]&m[791]&~m[815])|(~m[788]&m[789]&m[790]&m[791]&~m[815]))&BiasedRNG[711])|(((m[788]&~m[789]&~m[790]&~m[791]&m[815])|(~m[788]&m[789]&~m[790]&~m[791]&m[815])|(~m[788]&~m[789]&m[790]&~m[791]&m[815])|(m[788]&m[789]&~m[790]&m[791]&m[815])|(m[788]&~m[789]&m[790]&m[791]&m[815])|(~m[788]&m[789]&m[790]&m[791]&m[815]))&~BiasedRNG[711])|((m[788]&m[789]&~m[790]&~m[791]&~m[815])|(m[788]&~m[789]&m[790]&~m[791]&~m[815])|(~m[788]&m[789]&m[790]&~m[791]&~m[815])|(m[788]&m[789]&m[790]&~m[791]&~m[815])|(m[788]&m[789]&m[790]&m[791]&~m[815])|(m[788]&m[789]&~m[790]&~m[791]&m[815])|(m[788]&~m[789]&m[790]&~m[791]&m[815])|(~m[788]&m[789]&m[790]&~m[791]&m[815])|(m[788]&m[789]&m[790]&~m[791]&m[815])|(m[788]&m[789]&m[790]&m[791]&m[815]))):InitCond[1427];
    m[797] = run?((((m[793]&~m[794]&~m[795]&~m[796]&~m[820])|(~m[793]&m[794]&~m[795]&~m[796]&~m[820])|(~m[793]&~m[794]&m[795]&~m[796]&~m[820])|(m[793]&m[794]&~m[795]&m[796]&~m[820])|(m[793]&~m[794]&m[795]&m[796]&~m[820])|(~m[793]&m[794]&m[795]&m[796]&~m[820]))&BiasedRNG[712])|(((m[793]&~m[794]&~m[795]&~m[796]&m[820])|(~m[793]&m[794]&~m[795]&~m[796]&m[820])|(~m[793]&~m[794]&m[795]&~m[796]&m[820])|(m[793]&m[794]&~m[795]&m[796]&m[820])|(m[793]&~m[794]&m[795]&m[796]&m[820])|(~m[793]&m[794]&m[795]&m[796]&m[820]))&~BiasedRNG[712])|((m[793]&m[794]&~m[795]&~m[796]&~m[820])|(m[793]&~m[794]&m[795]&~m[796]&~m[820])|(~m[793]&m[794]&m[795]&~m[796]&~m[820])|(m[793]&m[794]&m[795]&~m[796]&~m[820])|(m[793]&m[794]&m[795]&m[796]&~m[820])|(m[793]&m[794]&~m[795]&~m[796]&m[820])|(m[793]&~m[794]&m[795]&~m[796]&m[820])|(~m[793]&m[794]&m[795]&~m[796]&m[820])|(m[793]&m[794]&m[795]&~m[796]&m[820])|(m[793]&m[794]&m[795]&m[796]&m[820]))):InitCond[1428];
    m[802] = run?((((m[798]&~m[799]&~m[800]&~m[801]&~m[825])|(~m[798]&m[799]&~m[800]&~m[801]&~m[825])|(~m[798]&~m[799]&m[800]&~m[801]&~m[825])|(m[798]&m[799]&~m[800]&m[801]&~m[825])|(m[798]&~m[799]&m[800]&m[801]&~m[825])|(~m[798]&m[799]&m[800]&m[801]&~m[825]))&BiasedRNG[713])|(((m[798]&~m[799]&~m[800]&~m[801]&m[825])|(~m[798]&m[799]&~m[800]&~m[801]&m[825])|(~m[798]&~m[799]&m[800]&~m[801]&m[825])|(m[798]&m[799]&~m[800]&m[801]&m[825])|(m[798]&~m[799]&m[800]&m[801]&m[825])|(~m[798]&m[799]&m[800]&m[801]&m[825]))&~BiasedRNG[713])|((m[798]&m[799]&~m[800]&~m[801]&~m[825])|(m[798]&~m[799]&m[800]&~m[801]&~m[825])|(~m[798]&m[799]&m[800]&~m[801]&~m[825])|(m[798]&m[799]&m[800]&~m[801]&~m[825])|(m[798]&m[799]&m[800]&m[801]&~m[825])|(m[798]&m[799]&~m[800]&~m[801]&m[825])|(m[798]&~m[799]&m[800]&~m[801]&m[825])|(~m[798]&m[799]&m[800]&~m[801]&m[825])|(m[798]&m[799]&m[800]&~m[801]&m[825])|(m[798]&m[799]&m[800]&m[801]&m[825]))):InitCond[1429];
    m[807] = run?((((m[803]&~m[804]&~m[805]&~m[806]&~m[835])|(~m[803]&m[804]&~m[805]&~m[806]&~m[835])|(~m[803]&~m[804]&m[805]&~m[806]&~m[835])|(m[803]&m[804]&~m[805]&m[806]&~m[835])|(m[803]&~m[804]&m[805]&m[806]&~m[835])|(~m[803]&m[804]&m[805]&m[806]&~m[835]))&BiasedRNG[714])|(((m[803]&~m[804]&~m[805]&~m[806]&m[835])|(~m[803]&m[804]&~m[805]&~m[806]&m[835])|(~m[803]&~m[804]&m[805]&~m[806]&m[835])|(m[803]&m[804]&~m[805]&m[806]&m[835])|(m[803]&~m[804]&m[805]&m[806]&m[835])|(~m[803]&m[804]&m[805]&m[806]&m[835]))&~BiasedRNG[714])|((m[803]&m[804]&~m[805]&~m[806]&~m[835])|(m[803]&~m[804]&m[805]&~m[806]&~m[835])|(~m[803]&m[804]&m[805]&~m[806]&~m[835])|(m[803]&m[804]&m[805]&~m[806]&~m[835])|(m[803]&m[804]&m[805]&m[806]&~m[835])|(m[803]&m[804]&~m[805]&~m[806]&m[835])|(m[803]&~m[804]&m[805]&~m[806]&m[835])|(~m[803]&m[804]&m[805]&~m[806]&m[835])|(m[803]&m[804]&m[805]&~m[806]&m[835])|(m[803]&m[804]&m[805]&m[806]&m[835]))):InitCond[1430];
    m[812] = run?((((m[808]&~m[809]&~m[810]&~m[811]&~m[840])|(~m[808]&m[809]&~m[810]&~m[811]&~m[840])|(~m[808]&~m[809]&m[810]&~m[811]&~m[840])|(m[808]&m[809]&~m[810]&m[811]&~m[840])|(m[808]&~m[809]&m[810]&m[811]&~m[840])|(~m[808]&m[809]&m[810]&m[811]&~m[840]))&BiasedRNG[715])|(((m[808]&~m[809]&~m[810]&~m[811]&m[840])|(~m[808]&m[809]&~m[810]&~m[811]&m[840])|(~m[808]&~m[809]&m[810]&~m[811]&m[840])|(m[808]&m[809]&~m[810]&m[811]&m[840])|(m[808]&~m[809]&m[810]&m[811]&m[840])|(~m[808]&m[809]&m[810]&m[811]&m[840]))&~BiasedRNG[715])|((m[808]&m[809]&~m[810]&~m[811]&~m[840])|(m[808]&~m[809]&m[810]&~m[811]&~m[840])|(~m[808]&m[809]&m[810]&~m[811]&~m[840])|(m[808]&m[809]&m[810]&~m[811]&~m[840])|(m[808]&m[809]&m[810]&m[811]&~m[840])|(m[808]&m[809]&~m[810]&~m[811]&m[840])|(m[808]&~m[809]&m[810]&~m[811]&m[840])|(~m[808]&m[809]&m[810]&~m[811]&m[840])|(m[808]&m[809]&m[810]&~m[811]&m[840])|(m[808]&m[809]&m[810]&m[811]&m[840]))):InitCond[1431];
    m[817] = run?((((m[813]&~m[814]&~m[815]&~m[816]&~m[845])|(~m[813]&m[814]&~m[815]&~m[816]&~m[845])|(~m[813]&~m[814]&m[815]&~m[816]&~m[845])|(m[813]&m[814]&~m[815]&m[816]&~m[845])|(m[813]&~m[814]&m[815]&m[816]&~m[845])|(~m[813]&m[814]&m[815]&m[816]&~m[845]))&BiasedRNG[716])|(((m[813]&~m[814]&~m[815]&~m[816]&m[845])|(~m[813]&m[814]&~m[815]&~m[816]&m[845])|(~m[813]&~m[814]&m[815]&~m[816]&m[845])|(m[813]&m[814]&~m[815]&m[816]&m[845])|(m[813]&~m[814]&m[815]&m[816]&m[845])|(~m[813]&m[814]&m[815]&m[816]&m[845]))&~BiasedRNG[716])|((m[813]&m[814]&~m[815]&~m[816]&~m[845])|(m[813]&~m[814]&m[815]&~m[816]&~m[845])|(~m[813]&m[814]&m[815]&~m[816]&~m[845])|(m[813]&m[814]&m[815]&~m[816]&~m[845])|(m[813]&m[814]&m[815]&m[816]&~m[845])|(m[813]&m[814]&~m[815]&~m[816]&m[845])|(m[813]&~m[814]&m[815]&~m[816]&m[845])|(~m[813]&m[814]&m[815]&~m[816]&m[845])|(m[813]&m[814]&m[815]&~m[816]&m[845])|(m[813]&m[814]&m[815]&m[816]&m[845]))):InitCond[1432];
    m[822] = run?((((m[818]&~m[819]&~m[820]&~m[821]&~m[850])|(~m[818]&m[819]&~m[820]&~m[821]&~m[850])|(~m[818]&~m[819]&m[820]&~m[821]&~m[850])|(m[818]&m[819]&~m[820]&m[821]&~m[850])|(m[818]&~m[819]&m[820]&m[821]&~m[850])|(~m[818]&m[819]&m[820]&m[821]&~m[850]))&BiasedRNG[717])|(((m[818]&~m[819]&~m[820]&~m[821]&m[850])|(~m[818]&m[819]&~m[820]&~m[821]&m[850])|(~m[818]&~m[819]&m[820]&~m[821]&m[850])|(m[818]&m[819]&~m[820]&m[821]&m[850])|(m[818]&~m[819]&m[820]&m[821]&m[850])|(~m[818]&m[819]&m[820]&m[821]&m[850]))&~BiasedRNG[717])|((m[818]&m[819]&~m[820]&~m[821]&~m[850])|(m[818]&~m[819]&m[820]&~m[821]&~m[850])|(~m[818]&m[819]&m[820]&~m[821]&~m[850])|(m[818]&m[819]&m[820]&~m[821]&~m[850])|(m[818]&m[819]&m[820]&m[821]&~m[850])|(m[818]&m[819]&~m[820]&~m[821]&m[850])|(m[818]&~m[819]&m[820]&~m[821]&m[850])|(~m[818]&m[819]&m[820]&~m[821]&m[850])|(m[818]&m[819]&m[820]&~m[821]&m[850])|(m[818]&m[819]&m[820]&m[821]&m[850]))):InitCond[1433];
    m[827] = run?((((m[823]&~m[824]&~m[825]&~m[826]&~m[855])|(~m[823]&m[824]&~m[825]&~m[826]&~m[855])|(~m[823]&~m[824]&m[825]&~m[826]&~m[855])|(m[823]&m[824]&~m[825]&m[826]&~m[855])|(m[823]&~m[824]&m[825]&m[826]&~m[855])|(~m[823]&m[824]&m[825]&m[826]&~m[855]))&BiasedRNG[718])|(((m[823]&~m[824]&~m[825]&~m[826]&m[855])|(~m[823]&m[824]&~m[825]&~m[826]&m[855])|(~m[823]&~m[824]&m[825]&~m[826]&m[855])|(m[823]&m[824]&~m[825]&m[826]&m[855])|(m[823]&~m[824]&m[825]&m[826]&m[855])|(~m[823]&m[824]&m[825]&m[826]&m[855]))&~BiasedRNG[718])|((m[823]&m[824]&~m[825]&~m[826]&~m[855])|(m[823]&~m[824]&m[825]&~m[826]&~m[855])|(~m[823]&m[824]&m[825]&~m[826]&~m[855])|(m[823]&m[824]&m[825]&~m[826]&~m[855])|(m[823]&m[824]&m[825]&m[826]&~m[855])|(m[823]&m[824]&~m[825]&~m[826]&m[855])|(m[823]&~m[824]&m[825]&~m[826]&m[855])|(~m[823]&m[824]&m[825]&~m[826]&m[855])|(m[823]&m[824]&m[825]&~m[826]&m[855])|(m[823]&m[824]&m[825]&m[826]&m[855]))):InitCond[1434];
    m[832] = run?((((m[828]&~m[829]&~m[830]&~m[831]&~m[860])|(~m[828]&m[829]&~m[830]&~m[831]&~m[860])|(~m[828]&~m[829]&m[830]&~m[831]&~m[860])|(m[828]&m[829]&~m[830]&m[831]&~m[860])|(m[828]&~m[829]&m[830]&m[831]&~m[860])|(~m[828]&m[829]&m[830]&m[831]&~m[860]))&BiasedRNG[719])|(((m[828]&~m[829]&~m[830]&~m[831]&m[860])|(~m[828]&m[829]&~m[830]&~m[831]&m[860])|(~m[828]&~m[829]&m[830]&~m[831]&m[860])|(m[828]&m[829]&~m[830]&m[831]&m[860])|(m[828]&~m[829]&m[830]&m[831]&m[860])|(~m[828]&m[829]&m[830]&m[831]&m[860]))&~BiasedRNG[719])|((m[828]&m[829]&~m[830]&~m[831]&~m[860])|(m[828]&~m[829]&m[830]&~m[831]&~m[860])|(~m[828]&m[829]&m[830]&~m[831]&~m[860])|(m[828]&m[829]&m[830]&~m[831]&~m[860])|(m[828]&m[829]&m[830]&m[831]&~m[860])|(m[828]&m[829]&~m[830]&~m[831]&m[860])|(m[828]&~m[829]&m[830]&~m[831]&m[860])|(~m[828]&m[829]&m[830]&~m[831]&m[860])|(m[828]&m[829]&m[830]&~m[831]&m[860])|(m[828]&m[829]&m[830]&m[831]&m[860]))):InitCond[1435];
    m[837] = run?((((m[833]&~m[834]&~m[835]&~m[836]&~m[870])|(~m[833]&m[834]&~m[835]&~m[836]&~m[870])|(~m[833]&~m[834]&m[835]&~m[836]&~m[870])|(m[833]&m[834]&~m[835]&m[836]&~m[870])|(m[833]&~m[834]&m[835]&m[836]&~m[870])|(~m[833]&m[834]&m[835]&m[836]&~m[870]))&BiasedRNG[720])|(((m[833]&~m[834]&~m[835]&~m[836]&m[870])|(~m[833]&m[834]&~m[835]&~m[836]&m[870])|(~m[833]&~m[834]&m[835]&~m[836]&m[870])|(m[833]&m[834]&~m[835]&m[836]&m[870])|(m[833]&~m[834]&m[835]&m[836]&m[870])|(~m[833]&m[834]&m[835]&m[836]&m[870]))&~BiasedRNG[720])|((m[833]&m[834]&~m[835]&~m[836]&~m[870])|(m[833]&~m[834]&m[835]&~m[836]&~m[870])|(~m[833]&m[834]&m[835]&~m[836]&~m[870])|(m[833]&m[834]&m[835]&~m[836]&~m[870])|(m[833]&m[834]&m[835]&m[836]&~m[870])|(m[833]&m[834]&~m[835]&~m[836]&m[870])|(m[833]&~m[834]&m[835]&~m[836]&m[870])|(~m[833]&m[834]&m[835]&~m[836]&m[870])|(m[833]&m[834]&m[835]&~m[836]&m[870])|(m[833]&m[834]&m[835]&m[836]&m[870]))):InitCond[1436];
    m[842] = run?((((m[838]&~m[839]&~m[840]&~m[841]&~m[875])|(~m[838]&m[839]&~m[840]&~m[841]&~m[875])|(~m[838]&~m[839]&m[840]&~m[841]&~m[875])|(m[838]&m[839]&~m[840]&m[841]&~m[875])|(m[838]&~m[839]&m[840]&m[841]&~m[875])|(~m[838]&m[839]&m[840]&m[841]&~m[875]))&BiasedRNG[721])|(((m[838]&~m[839]&~m[840]&~m[841]&m[875])|(~m[838]&m[839]&~m[840]&~m[841]&m[875])|(~m[838]&~m[839]&m[840]&~m[841]&m[875])|(m[838]&m[839]&~m[840]&m[841]&m[875])|(m[838]&~m[839]&m[840]&m[841]&m[875])|(~m[838]&m[839]&m[840]&m[841]&m[875]))&~BiasedRNG[721])|((m[838]&m[839]&~m[840]&~m[841]&~m[875])|(m[838]&~m[839]&m[840]&~m[841]&~m[875])|(~m[838]&m[839]&m[840]&~m[841]&~m[875])|(m[838]&m[839]&m[840]&~m[841]&~m[875])|(m[838]&m[839]&m[840]&m[841]&~m[875])|(m[838]&m[839]&~m[840]&~m[841]&m[875])|(m[838]&~m[839]&m[840]&~m[841]&m[875])|(~m[838]&m[839]&m[840]&~m[841]&m[875])|(m[838]&m[839]&m[840]&~m[841]&m[875])|(m[838]&m[839]&m[840]&m[841]&m[875]))):InitCond[1437];
    m[847] = run?((((m[843]&~m[844]&~m[845]&~m[846]&~m[880])|(~m[843]&m[844]&~m[845]&~m[846]&~m[880])|(~m[843]&~m[844]&m[845]&~m[846]&~m[880])|(m[843]&m[844]&~m[845]&m[846]&~m[880])|(m[843]&~m[844]&m[845]&m[846]&~m[880])|(~m[843]&m[844]&m[845]&m[846]&~m[880]))&BiasedRNG[722])|(((m[843]&~m[844]&~m[845]&~m[846]&m[880])|(~m[843]&m[844]&~m[845]&~m[846]&m[880])|(~m[843]&~m[844]&m[845]&~m[846]&m[880])|(m[843]&m[844]&~m[845]&m[846]&m[880])|(m[843]&~m[844]&m[845]&m[846]&m[880])|(~m[843]&m[844]&m[845]&m[846]&m[880]))&~BiasedRNG[722])|((m[843]&m[844]&~m[845]&~m[846]&~m[880])|(m[843]&~m[844]&m[845]&~m[846]&~m[880])|(~m[843]&m[844]&m[845]&~m[846]&~m[880])|(m[843]&m[844]&m[845]&~m[846]&~m[880])|(m[843]&m[844]&m[845]&m[846]&~m[880])|(m[843]&m[844]&~m[845]&~m[846]&m[880])|(m[843]&~m[844]&m[845]&~m[846]&m[880])|(~m[843]&m[844]&m[845]&~m[846]&m[880])|(m[843]&m[844]&m[845]&~m[846]&m[880])|(m[843]&m[844]&m[845]&m[846]&m[880]))):InitCond[1438];
    m[852] = run?((((m[848]&~m[849]&~m[850]&~m[851]&~m[885])|(~m[848]&m[849]&~m[850]&~m[851]&~m[885])|(~m[848]&~m[849]&m[850]&~m[851]&~m[885])|(m[848]&m[849]&~m[850]&m[851]&~m[885])|(m[848]&~m[849]&m[850]&m[851]&~m[885])|(~m[848]&m[849]&m[850]&m[851]&~m[885]))&BiasedRNG[723])|(((m[848]&~m[849]&~m[850]&~m[851]&m[885])|(~m[848]&m[849]&~m[850]&~m[851]&m[885])|(~m[848]&~m[849]&m[850]&~m[851]&m[885])|(m[848]&m[849]&~m[850]&m[851]&m[885])|(m[848]&~m[849]&m[850]&m[851]&m[885])|(~m[848]&m[849]&m[850]&m[851]&m[885]))&~BiasedRNG[723])|((m[848]&m[849]&~m[850]&~m[851]&~m[885])|(m[848]&~m[849]&m[850]&~m[851]&~m[885])|(~m[848]&m[849]&m[850]&~m[851]&~m[885])|(m[848]&m[849]&m[850]&~m[851]&~m[885])|(m[848]&m[849]&m[850]&m[851]&~m[885])|(m[848]&m[849]&~m[850]&~m[851]&m[885])|(m[848]&~m[849]&m[850]&~m[851]&m[885])|(~m[848]&m[849]&m[850]&~m[851]&m[885])|(m[848]&m[849]&m[850]&~m[851]&m[885])|(m[848]&m[849]&m[850]&m[851]&m[885]))):InitCond[1439];
    m[857] = run?((((m[853]&~m[854]&~m[855]&~m[856]&~m[890])|(~m[853]&m[854]&~m[855]&~m[856]&~m[890])|(~m[853]&~m[854]&m[855]&~m[856]&~m[890])|(m[853]&m[854]&~m[855]&m[856]&~m[890])|(m[853]&~m[854]&m[855]&m[856]&~m[890])|(~m[853]&m[854]&m[855]&m[856]&~m[890]))&BiasedRNG[724])|(((m[853]&~m[854]&~m[855]&~m[856]&m[890])|(~m[853]&m[854]&~m[855]&~m[856]&m[890])|(~m[853]&~m[854]&m[855]&~m[856]&m[890])|(m[853]&m[854]&~m[855]&m[856]&m[890])|(m[853]&~m[854]&m[855]&m[856]&m[890])|(~m[853]&m[854]&m[855]&m[856]&m[890]))&~BiasedRNG[724])|((m[853]&m[854]&~m[855]&~m[856]&~m[890])|(m[853]&~m[854]&m[855]&~m[856]&~m[890])|(~m[853]&m[854]&m[855]&~m[856]&~m[890])|(m[853]&m[854]&m[855]&~m[856]&~m[890])|(m[853]&m[854]&m[855]&m[856]&~m[890])|(m[853]&m[854]&~m[855]&~m[856]&m[890])|(m[853]&~m[854]&m[855]&~m[856]&m[890])|(~m[853]&m[854]&m[855]&~m[856]&m[890])|(m[853]&m[854]&m[855]&~m[856]&m[890])|(m[853]&m[854]&m[855]&m[856]&m[890]))):InitCond[1440];
    m[862] = run?((((m[858]&~m[859]&~m[860]&~m[861]&~m[895])|(~m[858]&m[859]&~m[860]&~m[861]&~m[895])|(~m[858]&~m[859]&m[860]&~m[861]&~m[895])|(m[858]&m[859]&~m[860]&m[861]&~m[895])|(m[858]&~m[859]&m[860]&m[861]&~m[895])|(~m[858]&m[859]&m[860]&m[861]&~m[895]))&BiasedRNG[725])|(((m[858]&~m[859]&~m[860]&~m[861]&m[895])|(~m[858]&m[859]&~m[860]&~m[861]&m[895])|(~m[858]&~m[859]&m[860]&~m[861]&m[895])|(m[858]&m[859]&~m[860]&m[861]&m[895])|(m[858]&~m[859]&m[860]&m[861]&m[895])|(~m[858]&m[859]&m[860]&m[861]&m[895]))&~BiasedRNG[725])|((m[858]&m[859]&~m[860]&~m[861]&~m[895])|(m[858]&~m[859]&m[860]&~m[861]&~m[895])|(~m[858]&m[859]&m[860]&~m[861]&~m[895])|(m[858]&m[859]&m[860]&~m[861]&~m[895])|(m[858]&m[859]&m[860]&m[861]&~m[895])|(m[858]&m[859]&~m[860]&~m[861]&m[895])|(m[858]&~m[859]&m[860]&~m[861]&m[895])|(~m[858]&m[859]&m[860]&~m[861]&m[895])|(m[858]&m[859]&m[860]&~m[861]&m[895])|(m[858]&m[859]&m[860]&m[861]&m[895]))):InitCond[1441];
    m[867] = run?((((m[863]&~m[864]&~m[865]&~m[866]&~m[900])|(~m[863]&m[864]&~m[865]&~m[866]&~m[900])|(~m[863]&~m[864]&m[865]&~m[866]&~m[900])|(m[863]&m[864]&~m[865]&m[866]&~m[900])|(m[863]&~m[864]&m[865]&m[866]&~m[900])|(~m[863]&m[864]&m[865]&m[866]&~m[900]))&BiasedRNG[726])|(((m[863]&~m[864]&~m[865]&~m[866]&m[900])|(~m[863]&m[864]&~m[865]&~m[866]&m[900])|(~m[863]&~m[864]&m[865]&~m[866]&m[900])|(m[863]&m[864]&~m[865]&m[866]&m[900])|(m[863]&~m[864]&m[865]&m[866]&m[900])|(~m[863]&m[864]&m[865]&m[866]&m[900]))&~BiasedRNG[726])|((m[863]&m[864]&~m[865]&~m[866]&~m[900])|(m[863]&~m[864]&m[865]&~m[866]&~m[900])|(~m[863]&m[864]&m[865]&~m[866]&~m[900])|(m[863]&m[864]&m[865]&~m[866]&~m[900])|(m[863]&m[864]&m[865]&m[866]&~m[900])|(m[863]&m[864]&~m[865]&~m[866]&m[900])|(m[863]&~m[864]&m[865]&~m[866]&m[900])|(~m[863]&m[864]&m[865]&~m[866]&m[900])|(m[863]&m[864]&m[865]&~m[866]&m[900])|(m[863]&m[864]&m[865]&m[866]&m[900]))):InitCond[1442];
    m[872] = run?((((m[868]&~m[869]&~m[870]&~m[871]&~m[910])|(~m[868]&m[869]&~m[870]&~m[871]&~m[910])|(~m[868]&~m[869]&m[870]&~m[871]&~m[910])|(m[868]&m[869]&~m[870]&m[871]&~m[910])|(m[868]&~m[869]&m[870]&m[871]&~m[910])|(~m[868]&m[869]&m[870]&m[871]&~m[910]))&BiasedRNG[727])|(((m[868]&~m[869]&~m[870]&~m[871]&m[910])|(~m[868]&m[869]&~m[870]&~m[871]&m[910])|(~m[868]&~m[869]&m[870]&~m[871]&m[910])|(m[868]&m[869]&~m[870]&m[871]&m[910])|(m[868]&~m[869]&m[870]&m[871]&m[910])|(~m[868]&m[869]&m[870]&m[871]&m[910]))&~BiasedRNG[727])|((m[868]&m[869]&~m[870]&~m[871]&~m[910])|(m[868]&~m[869]&m[870]&~m[871]&~m[910])|(~m[868]&m[869]&m[870]&~m[871]&~m[910])|(m[868]&m[869]&m[870]&~m[871]&~m[910])|(m[868]&m[869]&m[870]&m[871]&~m[910])|(m[868]&m[869]&~m[870]&~m[871]&m[910])|(m[868]&~m[869]&m[870]&~m[871]&m[910])|(~m[868]&m[869]&m[870]&~m[871]&m[910])|(m[868]&m[869]&m[870]&~m[871]&m[910])|(m[868]&m[869]&m[870]&m[871]&m[910]))):InitCond[1443];
    m[877] = run?((((m[873]&~m[874]&~m[875]&~m[876]&~m[915])|(~m[873]&m[874]&~m[875]&~m[876]&~m[915])|(~m[873]&~m[874]&m[875]&~m[876]&~m[915])|(m[873]&m[874]&~m[875]&m[876]&~m[915])|(m[873]&~m[874]&m[875]&m[876]&~m[915])|(~m[873]&m[874]&m[875]&m[876]&~m[915]))&BiasedRNG[728])|(((m[873]&~m[874]&~m[875]&~m[876]&m[915])|(~m[873]&m[874]&~m[875]&~m[876]&m[915])|(~m[873]&~m[874]&m[875]&~m[876]&m[915])|(m[873]&m[874]&~m[875]&m[876]&m[915])|(m[873]&~m[874]&m[875]&m[876]&m[915])|(~m[873]&m[874]&m[875]&m[876]&m[915]))&~BiasedRNG[728])|((m[873]&m[874]&~m[875]&~m[876]&~m[915])|(m[873]&~m[874]&m[875]&~m[876]&~m[915])|(~m[873]&m[874]&m[875]&~m[876]&~m[915])|(m[873]&m[874]&m[875]&~m[876]&~m[915])|(m[873]&m[874]&m[875]&m[876]&~m[915])|(m[873]&m[874]&~m[875]&~m[876]&m[915])|(m[873]&~m[874]&m[875]&~m[876]&m[915])|(~m[873]&m[874]&m[875]&~m[876]&m[915])|(m[873]&m[874]&m[875]&~m[876]&m[915])|(m[873]&m[874]&m[875]&m[876]&m[915]))):InitCond[1444];
    m[882] = run?((((m[878]&~m[879]&~m[880]&~m[881]&~m[920])|(~m[878]&m[879]&~m[880]&~m[881]&~m[920])|(~m[878]&~m[879]&m[880]&~m[881]&~m[920])|(m[878]&m[879]&~m[880]&m[881]&~m[920])|(m[878]&~m[879]&m[880]&m[881]&~m[920])|(~m[878]&m[879]&m[880]&m[881]&~m[920]))&BiasedRNG[729])|(((m[878]&~m[879]&~m[880]&~m[881]&m[920])|(~m[878]&m[879]&~m[880]&~m[881]&m[920])|(~m[878]&~m[879]&m[880]&~m[881]&m[920])|(m[878]&m[879]&~m[880]&m[881]&m[920])|(m[878]&~m[879]&m[880]&m[881]&m[920])|(~m[878]&m[879]&m[880]&m[881]&m[920]))&~BiasedRNG[729])|((m[878]&m[879]&~m[880]&~m[881]&~m[920])|(m[878]&~m[879]&m[880]&~m[881]&~m[920])|(~m[878]&m[879]&m[880]&~m[881]&~m[920])|(m[878]&m[879]&m[880]&~m[881]&~m[920])|(m[878]&m[879]&m[880]&m[881]&~m[920])|(m[878]&m[879]&~m[880]&~m[881]&m[920])|(m[878]&~m[879]&m[880]&~m[881]&m[920])|(~m[878]&m[879]&m[880]&~m[881]&m[920])|(m[878]&m[879]&m[880]&~m[881]&m[920])|(m[878]&m[879]&m[880]&m[881]&m[920]))):InitCond[1445];
    m[887] = run?((((m[883]&~m[884]&~m[885]&~m[886]&~m[925])|(~m[883]&m[884]&~m[885]&~m[886]&~m[925])|(~m[883]&~m[884]&m[885]&~m[886]&~m[925])|(m[883]&m[884]&~m[885]&m[886]&~m[925])|(m[883]&~m[884]&m[885]&m[886]&~m[925])|(~m[883]&m[884]&m[885]&m[886]&~m[925]))&BiasedRNG[730])|(((m[883]&~m[884]&~m[885]&~m[886]&m[925])|(~m[883]&m[884]&~m[885]&~m[886]&m[925])|(~m[883]&~m[884]&m[885]&~m[886]&m[925])|(m[883]&m[884]&~m[885]&m[886]&m[925])|(m[883]&~m[884]&m[885]&m[886]&m[925])|(~m[883]&m[884]&m[885]&m[886]&m[925]))&~BiasedRNG[730])|((m[883]&m[884]&~m[885]&~m[886]&~m[925])|(m[883]&~m[884]&m[885]&~m[886]&~m[925])|(~m[883]&m[884]&m[885]&~m[886]&~m[925])|(m[883]&m[884]&m[885]&~m[886]&~m[925])|(m[883]&m[884]&m[885]&m[886]&~m[925])|(m[883]&m[884]&~m[885]&~m[886]&m[925])|(m[883]&~m[884]&m[885]&~m[886]&m[925])|(~m[883]&m[884]&m[885]&~m[886]&m[925])|(m[883]&m[884]&m[885]&~m[886]&m[925])|(m[883]&m[884]&m[885]&m[886]&m[925]))):InitCond[1446];
    m[892] = run?((((m[888]&~m[889]&~m[890]&~m[891]&~m[930])|(~m[888]&m[889]&~m[890]&~m[891]&~m[930])|(~m[888]&~m[889]&m[890]&~m[891]&~m[930])|(m[888]&m[889]&~m[890]&m[891]&~m[930])|(m[888]&~m[889]&m[890]&m[891]&~m[930])|(~m[888]&m[889]&m[890]&m[891]&~m[930]))&BiasedRNG[731])|(((m[888]&~m[889]&~m[890]&~m[891]&m[930])|(~m[888]&m[889]&~m[890]&~m[891]&m[930])|(~m[888]&~m[889]&m[890]&~m[891]&m[930])|(m[888]&m[889]&~m[890]&m[891]&m[930])|(m[888]&~m[889]&m[890]&m[891]&m[930])|(~m[888]&m[889]&m[890]&m[891]&m[930]))&~BiasedRNG[731])|((m[888]&m[889]&~m[890]&~m[891]&~m[930])|(m[888]&~m[889]&m[890]&~m[891]&~m[930])|(~m[888]&m[889]&m[890]&~m[891]&~m[930])|(m[888]&m[889]&m[890]&~m[891]&~m[930])|(m[888]&m[889]&m[890]&m[891]&~m[930])|(m[888]&m[889]&~m[890]&~m[891]&m[930])|(m[888]&~m[889]&m[890]&~m[891]&m[930])|(~m[888]&m[889]&m[890]&~m[891]&m[930])|(m[888]&m[889]&m[890]&~m[891]&m[930])|(m[888]&m[889]&m[890]&m[891]&m[930]))):InitCond[1447];
    m[897] = run?((((m[893]&~m[894]&~m[895]&~m[896]&~m[935])|(~m[893]&m[894]&~m[895]&~m[896]&~m[935])|(~m[893]&~m[894]&m[895]&~m[896]&~m[935])|(m[893]&m[894]&~m[895]&m[896]&~m[935])|(m[893]&~m[894]&m[895]&m[896]&~m[935])|(~m[893]&m[894]&m[895]&m[896]&~m[935]))&BiasedRNG[732])|(((m[893]&~m[894]&~m[895]&~m[896]&m[935])|(~m[893]&m[894]&~m[895]&~m[896]&m[935])|(~m[893]&~m[894]&m[895]&~m[896]&m[935])|(m[893]&m[894]&~m[895]&m[896]&m[935])|(m[893]&~m[894]&m[895]&m[896]&m[935])|(~m[893]&m[894]&m[895]&m[896]&m[935]))&~BiasedRNG[732])|((m[893]&m[894]&~m[895]&~m[896]&~m[935])|(m[893]&~m[894]&m[895]&~m[896]&~m[935])|(~m[893]&m[894]&m[895]&~m[896]&~m[935])|(m[893]&m[894]&m[895]&~m[896]&~m[935])|(m[893]&m[894]&m[895]&m[896]&~m[935])|(m[893]&m[894]&~m[895]&~m[896]&m[935])|(m[893]&~m[894]&m[895]&~m[896]&m[935])|(~m[893]&m[894]&m[895]&~m[896]&m[935])|(m[893]&m[894]&m[895]&~m[896]&m[935])|(m[893]&m[894]&m[895]&m[896]&m[935]))):InitCond[1448];
    m[902] = run?((((m[898]&~m[899]&~m[900]&~m[901]&~m[940])|(~m[898]&m[899]&~m[900]&~m[901]&~m[940])|(~m[898]&~m[899]&m[900]&~m[901]&~m[940])|(m[898]&m[899]&~m[900]&m[901]&~m[940])|(m[898]&~m[899]&m[900]&m[901]&~m[940])|(~m[898]&m[899]&m[900]&m[901]&~m[940]))&BiasedRNG[733])|(((m[898]&~m[899]&~m[900]&~m[901]&m[940])|(~m[898]&m[899]&~m[900]&~m[901]&m[940])|(~m[898]&~m[899]&m[900]&~m[901]&m[940])|(m[898]&m[899]&~m[900]&m[901]&m[940])|(m[898]&~m[899]&m[900]&m[901]&m[940])|(~m[898]&m[899]&m[900]&m[901]&m[940]))&~BiasedRNG[733])|((m[898]&m[899]&~m[900]&~m[901]&~m[940])|(m[898]&~m[899]&m[900]&~m[901]&~m[940])|(~m[898]&m[899]&m[900]&~m[901]&~m[940])|(m[898]&m[899]&m[900]&~m[901]&~m[940])|(m[898]&m[899]&m[900]&m[901]&~m[940])|(m[898]&m[899]&~m[900]&~m[901]&m[940])|(m[898]&~m[899]&m[900]&~m[901]&m[940])|(~m[898]&m[899]&m[900]&~m[901]&m[940])|(m[898]&m[899]&m[900]&~m[901]&m[940])|(m[898]&m[899]&m[900]&m[901]&m[940]))):InitCond[1449];
    m[907] = run?((((m[903]&~m[904]&~m[905]&~m[906]&~m[945])|(~m[903]&m[904]&~m[905]&~m[906]&~m[945])|(~m[903]&~m[904]&m[905]&~m[906]&~m[945])|(m[903]&m[904]&~m[905]&m[906]&~m[945])|(m[903]&~m[904]&m[905]&m[906]&~m[945])|(~m[903]&m[904]&m[905]&m[906]&~m[945]))&BiasedRNG[734])|(((m[903]&~m[904]&~m[905]&~m[906]&m[945])|(~m[903]&m[904]&~m[905]&~m[906]&m[945])|(~m[903]&~m[904]&m[905]&~m[906]&m[945])|(m[903]&m[904]&~m[905]&m[906]&m[945])|(m[903]&~m[904]&m[905]&m[906]&m[945])|(~m[903]&m[904]&m[905]&m[906]&m[945]))&~BiasedRNG[734])|((m[903]&m[904]&~m[905]&~m[906]&~m[945])|(m[903]&~m[904]&m[905]&~m[906]&~m[945])|(~m[903]&m[904]&m[905]&~m[906]&~m[945])|(m[903]&m[904]&m[905]&~m[906]&~m[945])|(m[903]&m[904]&m[905]&m[906]&~m[945])|(m[903]&m[904]&~m[905]&~m[906]&m[945])|(m[903]&~m[904]&m[905]&~m[906]&m[945])|(~m[903]&m[904]&m[905]&~m[906]&m[945])|(m[903]&m[904]&m[905]&~m[906]&m[945])|(m[903]&m[904]&m[905]&m[906]&m[945]))):InitCond[1450];
    m[912] = run?((((m[908]&~m[909]&~m[910]&~m[911]&~m[955])|(~m[908]&m[909]&~m[910]&~m[911]&~m[955])|(~m[908]&~m[909]&m[910]&~m[911]&~m[955])|(m[908]&m[909]&~m[910]&m[911]&~m[955])|(m[908]&~m[909]&m[910]&m[911]&~m[955])|(~m[908]&m[909]&m[910]&m[911]&~m[955]))&BiasedRNG[735])|(((m[908]&~m[909]&~m[910]&~m[911]&m[955])|(~m[908]&m[909]&~m[910]&~m[911]&m[955])|(~m[908]&~m[909]&m[910]&~m[911]&m[955])|(m[908]&m[909]&~m[910]&m[911]&m[955])|(m[908]&~m[909]&m[910]&m[911]&m[955])|(~m[908]&m[909]&m[910]&m[911]&m[955]))&~BiasedRNG[735])|((m[908]&m[909]&~m[910]&~m[911]&~m[955])|(m[908]&~m[909]&m[910]&~m[911]&~m[955])|(~m[908]&m[909]&m[910]&~m[911]&~m[955])|(m[908]&m[909]&m[910]&~m[911]&~m[955])|(m[908]&m[909]&m[910]&m[911]&~m[955])|(m[908]&m[909]&~m[910]&~m[911]&m[955])|(m[908]&~m[909]&m[910]&~m[911]&m[955])|(~m[908]&m[909]&m[910]&~m[911]&m[955])|(m[908]&m[909]&m[910]&~m[911]&m[955])|(m[908]&m[909]&m[910]&m[911]&m[955]))):InitCond[1451];
    m[917] = run?((((m[913]&~m[914]&~m[915]&~m[916]&~m[960])|(~m[913]&m[914]&~m[915]&~m[916]&~m[960])|(~m[913]&~m[914]&m[915]&~m[916]&~m[960])|(m[913]&m[914]&~m[915]&m[916]&~m[960])|(m[913]&~m[914]&m[915]&m[916]&~m[960])|(~m[913]&m[914]&m[915]&m[916]&~m[960]))&BiasedRNG[736])|(((m[913]&~m[914]&~m[915]&~m[916]&m[960])|(~m[913]&m[914]&~m[915]&~m[916]&m[960])|(~m[913]&~m[914]&m[915]&~m[916]&m[960])|(m[913]&m[914]&~m[915]&m[916]&m[960])|(m[913]&~m[914]&m[915]&m[916]&m[960])|(~m[913]&m[914]&m[915]&m[916]&m[960]))&~BiasedRNG[736])|((m[913]&m[914]&~m[915]&~m[916]&~m[960])|(m[913]&~m[914]&m[915]&~m[916]&~m[960])|(~m[913]&m[914]&m[915]&~m[916]&~m[960])|(m[913]&m[914]&m[915]&~m[916]&~m[960])|(m[913]&m[914]&m[915]&m[916]&~m[960])|(m[913]&m[914]&~m[915]&~m[916]&m[960])|(m[913]&~m[914]&m[915]&~m[916]&m[960])|(~m[913]&m[914]&m[915]&~m[916]&m[960])|(m[913]&m[914]&m[915]&~m[916]&m[960])|(m[913]&m[914]&m[915]&m[916]&m[960]))):InitCond[1452];
    m[922] = run?((((m[918]&~m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&~m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&~m[920]&m[921]&~m[965])|(m[918]&~m[919]&m[920]&m[921]&~m[965])|(~m[918]&m[919]&m[920]&m[921]&~m[965]))&BiasedRNG[737])|(((m[918]&~m[919]&~m[920]&~m[921]&m[965])|(~m[918]&m[919]&~m[920]&~m[921]&m[965])|(~m[918]&~m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&~m[920]&m[921]&m[965])|(m[918]&~m[919]&m[920]&m[921]&m[965])|(~m[918]&m[919]&m[920]&m[921]&m[965]))&~BiasedRNG[737])|((m[918]&m[919]&~m[920]&~m[921]&~m[965])|(m[918]&~m[919]&m[920]&~m[921]&~m[965])|(~m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&m[921]&~m[965])|(m[918]&m[919]&~m[920]&~m[921]&m[965])|(m[918]&~m[919]&m[920]&~m[921]&m[965])|(~m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&m[921]&m[965]))):InitCond[1453];
    m[927] = run?((((m[923]&~m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&~m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&~m[925]&m[926]&~m[970])|(m[923]&~m[924]&m[925]&m[926]&~m[970])|(~m[923]&m[924]&m[925]&m[926]&~m[970]))&BiasedRNG[738])|(((m[923]&~m[924]&~m[925]&~m[926]&m[970])|(~m[923]&m[924]&~m[925]&~m[926]&m[970])|(~m[923]&~m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&~m[925]&m[926]&m[970])|(m[923]&~m[924]&m[925]&m[926]&m[970])|(~m[923]&m[924]&m[925]&m[926]&m[970]))&~BiasedRNG[738])|((m[923]&m[924]&~m[925]&~m[926]&~m[970])|(m[923]&~m[924]&m[925]&~m[926]&~m[970])|(~m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&m[926]&~m[970])|(m[923]&m[924]&~m[925]&~m[926]&m[970])|(m[923]&~m[924]&m[925]&~m[926]&m[970])|(~m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&m[926]&m[970]))):InitCond[1454];
    m[932] = run?((((m[928]&~m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&~m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&~m[930]&m[931]&~m[975])|(m[928]&~m[929]&m[930]&m[931]&~m[975])|(~m[928]&m[929]&m[930]&m[931]&~m[975]))&BiasedRNG[739])|(((m[928]&~m[929]&~m[930]&~m[931]&m[975])|(~m[928]&m[929]&~m[930]&~m[931]&m[975])|(~m[928]&~m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&~m[930]&m[931]&m[975])|(m[928]&~m[929]&m[930]&m[931]&m[975])|(~m[928]&m[929]&m[930]&m[931]&m[975]))&~BiasedRNG[739])|((m[928]&m[929]&~m[930]&~m[931]&~m[975])|(m[928]&~m[929]&m[930]&~m[931]&~m[975])|(~m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&m[931]&~m[975])|(m[928]&m[929]&~m[930]&~m[931]&m[975])|(m[928]&~m[929]&m[930]&~m[931]&m[975])|(~m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&m[931]&m[975]))):InitCond[1455];
    m[937] = run?((((m[933]&~m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&~m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&~m[935]&m[936]&~m[980])|(m[933]&~m[934]&m[935]&m[936]&~m[980])|(~m[933]&m[934]&m[935]&m[936]&~m[980]))&BiasedRNG[740])|(((m[933]&~m[934]&~m[935]&~m[936]&m[980])|(~m[933]&m[934]&~m[935]&~m[936]&m[980])|(~m[933]&~m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&~m[935]&m[936]&m[980])|(m[933]&~m[934]&m[935]&m[936]&m[980])|(~m[933]&m[934]&m[935]&m[936]&m[980]))&~BiasedRNG[740])|((m[933]&m[934]&~m[935]&~m[936]&~m[980])|(m[933]&~m[934]&m[935]&~m[936]&~m[980])|(~m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&m[936]&~m[980])|(m[933]&m[934]&~m[935]&~m[936]&m[980])|(m[933]&~m[934]&m[935]&~m[936]&m[980])|(~m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&m[936]&m[980]))):InitCond[1456];
    m[942] = run?((((m[938]&~m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&~m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&~m[940]&m[941]&~m[985])|(m[938]&~m[939]&m[940]&m[941]&~m[985])|(~m[938]&m[939]&m[940]&m[941]&~m[985]))&BiasedRNG[741])|(((m[938]&~m[939]&~m[940]&~m[941]&m[985])|(~m[938]&m[939]&~m[940]&~m[941]&m[985])|(~m[938]&~m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&~m[940]&m[941]&m[985])|(m[938]&~m[939]&m[940]&m[941]&m[985])|(~m[938]&m[939]&m[940]&m[941]&m[985]))&~BiasedRNG[741])|((m[938]&m[939]&~m[940]&~m[941]&~m[985])|(m[938]&~m[939]&m[940]&~m[941]&~m[985])|(~m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&m[941]&~m[985])|(m[938]&m[939]&~m[940]&~m[941]&m[985])|(m[938]&~m[939]&m[940]&~m[941]&m[985])|(~m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&m[941]&m[985]))):InitCond[1457];
    m[947] = run?((((m[943]&~m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&~m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&~m[945]&m[946]&~m[990])|(m[943]&~m[944]&m[945]&m[946]&~m[990])|(~m[943]&m[944]&m[945]&m[946]&~m[990]))&BiasedRNG[742])|(((m[943]&~m[944]&~m[945]&~m[946]&m[990])|(~m[943]&m[944]&~m[945]&~m[946]&m[990])|(~m[943]&~m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&~m[945]&m[946]&m[990])|(m[943]&~m[944]&m[945]&m[946]&m[990])|(~m[943]&m[944]&m[945]&m[946]&m[990]))&~BiasedRNG[742])|((m[943]&m[944]&~m[945]&~m[946]&~m[990])|(m[943]&~m[944]&m[945]&~m[946]&~m[990])|(~m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&m[946]&~m[990])|(m[943]&m[944]&~m[945]&~m[946]&m[990])|(m[943]&~m[944]&m[945]&~m[946]&m[990])|(~m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&m[946]&m[990]))):InitCond[1458];
    m[952] = run?((((m[948]&~m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&~m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&~m[950]&m[951]&~m[995])|(m[948]&~m[949]&m[950]&m[951]&~m[995])|(~m[948]&m[949]&m[950]&m[951]&~m[995]))&BiasedRNG[743])|(((m[948]&~m[949]&~m[950]&~m[951]&m[995])|(~m[948]&m[949]&~m[950]&~m[951]&m[995])|(~m[948]&~m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&~m[950]&m[951]&m[995])|(m[948]&~m[949]&m[950]&m[951]&m[995])|(~m[948]&m[949]&m[950]&m[951]&m[995]))&~BiasedRNG[743])|((m[948]&m[949]&~m[950]&~m[951]&~m[995])|(m[948]&~m[949]&m[950]&~m[951]&~m[995])|(~m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&m[951]&~m[995])|(m[948]&m[949]&~m[950]&~m[951]&m[995])|(m[948]&~m[949]&m[950]&~m[951]&m[995])|(~m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&m[951]&m[995]))):InitCond[1459];
    m[957] = run?((((m[953]&~m[954]&~m[955]&~m[956]&~m[1005])|(~m[953]&m[954]&~m[955]&~m[956]&~m[1005])|(~m[953]&~m[954]&m[955]&~m[956]&~m[1005])|(m[953]&m[954]&~m[955]&m[956]&~m[1005])|(m[953]&~m[954]&m[955]&m[956]&~m[1005])|(~m[953]&m[954]&m[955]&m[956]&~m[1005]))&BiasedRNG[744])|(((m[953]&~m[954]&~m[955]&~m[956]&m[1005])|(~m[953]&m[954]&~m[955]&~m[956]&m[1005])|(~m[953]&~m[954]&m[955]&~m[956]&m[1005])|(m[953]&m[954]&~m[955]&m[956]&m[1005])|(m[953]&~m[954]&m[955]&m[956]&m[1005])|(~m[953]&m[954]&m[955]&m[956]&m[1005]))&~BiasedRNG[744])|((m[953]&m[954]&~m[955]&~m[956]&~m[1005])|(m[953]&~m[954]&m[955]&~m[956]&~m[1005])|(~m[953]&m[954]&m[955]&~m[956]&~m[1005])|(m[953]&m[954]&m[955]&~m[956]&~m[1005])|(m[953]&m[954]&m[955]&m[956]&~m[1005])|(m[953]&m[954]&~m[955]&~m[956]&m[1005])|(m[953]&~m[954]&m[955]&~m[956]&m[1005])|(~m[953]&m[954]&m[955]&~m[956]&m[1005])|(m[953]&m[954]&m[955]&~m[956]&m[1005])|(m[953]&m[954]&m[955]&m[956]&m[1005]))):InitCond[1460];
    m[962] = run?((((m[958]&~m[959]&~m[960]&~m[961]&~m[1010])|(~m[958]&m[959]&~m[960]&~m[961]&~m[1010])|(~m[958]&~m[959]&m[960]&~m[961]&~m[1010])|(m[958]&m[959]&~m[960]&m[961]&~m[1010])|(m[958]&~m[959]&m[960]&m[961]&~m[1010])|(~m[958]&m[959]&m[960]&m[961]&~m[1010]))&BiasedRNG[745])|(((m[958]&~m[959]&~m[960]&~m[961]&m[1010])|(~m[958]&m[959]&~m[960]&~m[961]&m[1010])|(~m[958]&~m[959]&m[960]&~m[961]&m[1010])|(m[958]&m[959]&~m[960]&m[961]&m[1010])|(m[958]&~m[959]&m[960]&m[961]&m[1010])|(~m[958]&m[959]&m[960]&m[961]&m[1010]))&~BiasedRNG[745])|((m[958]&m[959]&~m[960]&~m[961]&~m[1010])|(m[958]&~m[959]&m[960]&~m[961]&~m[1010])|(~m[958]&m[959]&m[960]&~m[961]&~m[1010])|(m[958]&m[959]&m[960]&~m[961]&~m[1010])|(m[958]&m[959]&m[960]&m[961]&~m[1010])|(m[958]&m[959]&~m[960]&~m[961]&m[1010])|(m[958]&~m[959]&m[960]&~m[961]&m[1010])|(~m[958]&m[959]&m[960]&~m[961]&m[1010])|(m[958]&m[959]&m[960]&~m[961]&m[1010])|(m[958]&m[959]&m[960]&m[961]&m[1010]))):InitCond[1461];
    m[967] = run?((((m[963]&~m[964]&~m[965]&~m[966]&~m[1015])|(~m[963]&m[964]&~m[965]&~m[966]&~m[1015])|(~m[963]&~m[964]&m[965]&~m[966]&~m[1015])|(m[963]&m[964]&~m[965]&m[966]&~m[1015])|(m[963]&~m[964]&m[965]&m[966]&~m[1015])|(~m[963]&m[964]&m[965]&m[966]&~m[1015]))&BiasedRNG[746])|(((m[963]&~m[964]&~m[965]&~m[966]&m[1015])|(~m[963]&m[964]&~m[965]&~m[966]&m[1015])|(~m[963]&~m[964]&m[965]&~m[966]&m[1015])|(m[963]&m[964]&~m[965]&m[966]&m[1015])|(m[963]&~m[964]&m[965]&m[966]&m[1015])|(~m[963]&m[964]&m[965]&m[966]&m[1015]))&~BiasedRNG[746])|((m[963]&m[964]&~m[965]&~m[966]&~m[1015])|(m[963]&~m[964]&m[965]&~m[966]&~m[1015])|(~m[963]&m[964]&m[965]&~m[966]&~m[1015])|(m[963]&m[964]&m[965]&~m[966]&~m[1015])|(m[963]&m[964]&m[965]&m[966]&~m[1015])|(m[963]&m[964]&~m[965]&~m[966]&m[1015])|(m[963]&~m[964]&m[965]&~m[966]&m[1015])|(~m[963]&m[964]&m[965]&~m[966]&m[1015])|(m[963]&m[964]&m[965]&~m[966]&m[1015])|(m[963]&m[964]&m[965]&m[966]&m[1015]))):InitCond[1462];
    m[972] = run?((((m[968]&~m[969]&~m[970]&~m[971]&~m[1020])|(~m[968]&m[969]&~m[970]&~m[971]&~m[1020])|(~m[968]&~m[969]&m[970]&~m[971]&~m[1020])|(m[968]&m[969]&~m[970]&m[971]&~m[1020])|(m[968]&~m[969]&m[970]&m[971]&~m[1020])|(~m[968]&m[969]&m[970]&m[971]&~m[1020]))&BiasedRNG[747])|(((m[968]&~m[969]&~m[970]&~m[971]&m[1020])|(~m[968]&m[969]&~m[970]&~m[971]&m[1020])|(~m[968]&~m[969]&m[970]&~m[971]&m[1020])|(m[968]&m[969]&~m[970]&m[971]&m[1020])|(m[968]&~m[969]&m[970]&m[971]&m[1020])|(~m[968]&m[969]&m[970]&m[971]&m[1020]))&~BiasedRNG[747])|((m[968]&m[969]&~m[970]&~m[971]&~m[1020])|(m[968]&~m[969]&m[970]&~m[971]&~m[1020])|(~m[968]&m[969]&m[970]&~m[971]&~m[1020])|(m[968]&m[969]&m[970]&~m[971]&~m[1020])|(m[968]&m[969]&m[970]&m[971]&~m[1020])|(m[968]&m[969]&~m[970]&~m[971]&m[1020])|(m[968]&~m[969]&m[970]&~m[971]&m[1020])|(~m[968]&m[969]&m[970]&~m[971]&m[1020])|(m[968]&m[969]&m[970]&~m[971]&m[1020])|(m[968]&m[969]&m[970]&m[971]&m[1020]))):InitCond[1463];
    m[977] = run?((((m[973]&~m[974]&~m[975]&~m[976]&~m[1025])|(~m[973]&m[974]&~m[975]&~m[976]&~m[1025])|(~m[973]&~m[974]&m[975]&~m[976]&~m[1025])|(m[973]&m[974]&~m[975]&m[976]&~m[1025])|(m[973]&~m[974]&m[975]&m[976]&~m[1025])|(~m[973]&m[974]&m[975]&m[976]&~m[1025]))&BiasedRNG[748])|(((m[973]&~m[974]&~m[975]&~m[976]&m[1025])|(~m[973]&m[974]&~m[975]&~m[976]&m[1025])|(~m[973]&~m[974]&m[975]&~m[976]&m[1025])|(m[973]&m[974]&~m[975]&m[976]&m[1025])|(m[973]&~m[974]&m[975]&m[976]&m[1025])|(~m[973]&m[974]&m[975]&m[976]&m[1025]))&~BiasedRNG[748])|((m[973]&m[974]&~m[975]&~m[976]&~m[1025])|(m[973]&~m[974]&m[975]&~m[976]&~m[1025])|(~m[973]&m[974]&m[975]&~m[976]&~m[1025])|(m[973]&m[974]&m[975]&~m[976]&~m[1025])|(m[973]&m[974]&m[975]&m[976]&~m[1025])|(m[973]&m[974]&~m[975]&~m[976]&m[1025])|(m[973]&~m[974]&m[975]&~m[976]&m[1025])|(~m[973]&m[974]&m[975]&~m[976]&m[1025])|(m[973]&m[974]&m[975]&~m[976]&m[1025])|(m[973]&m[974]&m[975]&m[976]&m[1025]))):InitCond[1464];
    m[982] = run?((((m[978]&~m[979]&~m[980]&~m[981]&~m[1030])|(~m[978]&m[979]&~m[980]&~m[981]&~m[1030])|(~m[978]&~m[979]&m[980]&~m[981]&~m[1030])|(m[978]&m[979]&~m[980]&m[981]&~m[1030])|(m[978]&~m[979]&m[980]&m[981]&~m[1030])|(~m[978]&m[979]&m[980]&m[981]&~m[1030]))&BiasedRNG[749])|(((m[978]&~m[979]&~m[980]&~m[981]&m[1030])|(~m[978]&m[979]&~m[980]&~m[981]&m[1030])|(~m[978]&~m[979]&m[980]&~m[981]&m[1030])|(m[978]&m[979]&~m[980]&m[981]&m[1030])|(m[978]&~m[979]&m[980]&m[981]&m[1030])|(~m[978]&m[979]&m[980]&m[981]&m[1030]))&~BiasedRNG[749])|((m[978]&m[979]&~m[980]&~m[981]&~m[1030])|(m[978]&~m[979]&m[980]&~m[981]&~m[1030])|(~m[978]&m[979]&m[980]&~m[981]&~m[1030])|(m[978]&m[979]&m[980]&~m[981]&~m[1030])|(m[978]&m[979]&m[980]&m[981]&~m[1030])|(m[978]&m[979]&~m[980]&~m[981]&m[1030])|(m[978]&~m[979]&m[980]&~m[981]&m[1030])|(~m[978]&m[979]&m[980]&~m[981]&m[1030])|(m[978]&m[979]&m[980]&~m[981]&m[1030])|(m[978]&m[979]&m[980]&m[981]&m[1030]))):InitCond[1465];
    m[987] = run?((((m[983]&~m[984]&~m[985]&~m[986]&~m[1035])|(~m[983]&m[984]&~m[985]&~m[986]&~m[1035])|(~m[983]&~m[984]&m[985]&~m[986]&~m[1035])|(m[983]&m[984]&~m[985]&m[986]&~m[1035])|(m[983]&~m[984]&m[985]&m[986]&~m[1035])|(~m[983]&m[984]&m[985]&m[986]&~m[1035]))&BiasedRNG[750])|(((m[983]&~m[984]&~m[985]&~m[986]&m[1035])|(~m[983]&m[984]&~m[985]&~m[986]&m[1035])|(~m[983]&~m[984]&m[985]&~m[986]&m[1035])|(m[983]&m[984]&~m[985]&m[986]&m[1035])|(m[983]&~m[984]&m[985]&m[986]&m[1035])|(~m[983]&m[984]&m[985]&m[986]&m[1035]))&~BiasedRNG[750])|((m[983]&m[984]&~m[985]&~m[986]&~m[1035])|(m[983]&~m[984]&m[985]&~m[986]&~m[1035])|(~m[983]&m[984]&m[985]&~m[986]&~m[1035])|(m[983]&m[984]&m[985]&~m[986]&~m[1035])|(m[983]&m[984]&m[985]&m[986]&~m[1035])|(m[983]&m[984]&~m[985]&~m[986]&m[1035])|(m[983]&~m[984]&m[985]&~m[986]&m[1035])|(~m[983]&m[984]&m[985]&~m[986]&m[1035])|(m[983]&m[984]&m[985]&~m[986]&m[1035])|(m[983]&m[984]&m[985]&m[986]&m[1035]))):InitCond[1466];
    m[992] = run?((((m[988]&~m[989]&~m[990]&~m[991]&~m[1040])|(~m[988]&m[989]&~m[990]&~m[991]&~m[1040])|(~m[988]&~m[989]&m[990]&~m[991]&~m[1040])|(m[988]&m[989]&~m[990]&m[991]&~m[1040])|(m[988]&~m[989]&m[990]&m[991]&~m[1040])|(~m[988]&m[989]&m[990]&m[991]&~m[1040]))&BiasedRNG[751])|(((m[988]&~m[989]&~m[990]&~m[991]&m[1040])|(~m[988]&m[989]&~m[990]&~m[991]&m[1040])|(~m[988]&~m[989]&m[990]&~m[991]&m[1040])|(m[988]&m[989]&~m[990]&m[991]&m[1040])|(m[988]&~m[989]&m[990]&m[991]&m[1040])|(~m[988]&m[989]&m[990]&m[991]&m[1040]))&~BiasedRNG[751])|((m[988]&m[989]&~m[990]&~m[991]&~m[1040])|(m[988]&~m[989]&m[990]&~m[991]&~m[1040])|(~m[988]&m[989]&m[990]&~m[991]&~m[1040])|(m[988]&m[989]&m[990]&~m[991]&~m[1040])|(m[988]&m[989]&m[990]&m[991]&~m[1040])|(m[988]&m[989]&~m[990]&~m[991]&m[1040])|(m[988]&~m[989]&m[990]&~m[991]&m[1040])|(~m[988]&m[989]&m[990]&~m[991]&m[1040])|(m[988]&m[989]&m[990]&~m[991]&m[1040])|(m[988]&m[989]&m[990]&m[991]&m[1040]))):InitCond[1467];
    m[997] = run?((((m[993]&~m[994]&~m[995]&~m[996]&~m[1045])|(~m[993]&m[994]&~m[995]&~m[996]&~m[1045])|(~m[993]&~m[994]&m[995]&~m[996]&~m[1045])|(m[993]&m[994]&~m[995]&m[996]&~m[1045])|(m[993]&~m[994]&m[995]&m[996]&~m[1045])|(~m[993]&m[994]&m[995]&m[996]&~m[1045]))&BiasedRNG[752])|(((m[993]&~m[994]&~m[995]&~m[996]&m[1045])|(~m[993]&m[994]&~m[995]&~m[996]&m[1045])|(~m[993]&~m[994]&m[995]&~m[996]&m[1045])|(m[993]&m[994]&~m[995]&m[996]&m[1045])|(m[993]&~m[994]&m[995]&m[996]&m[1045])|(~m[993]&m[994]&m[995]&m[996]&m[1045]))&~BiasedRNG[752])|((m[993]&m[994]&~m[995]&~m[996]&~m[1045])|(m[993]&~m[994]&m[995]&~m[996]&~m[1045])|(~m[993]&m[994]&m[995]&~m[996]&~m[1045])|(m[993]&m[994]&m[995]&~m[996]&~m[1045])|(m[993]&m[994]&m[995]&m[996]&~m[1045])|(m[993]&m[994]&~m[995]&~m[996]&m[1045])|(m[993]&~m[994]&m[995]&~m[996]&m[1045])|(~m[993]&m[994]&m[995]&~m[996]&m[1045])|(m[993]&m[994]&m[995]&~m[996]&m[1045])|(m[993]&m[994]&m[995]&m[996]&m[1045]))):InitCond[1468];
    m[1002] = run?((((m[998]&~m[999]&~m[1000]&~m[1001]&~m[1050])|(~m[998]&m[999]&~m[1000]&~m[1001]&~m[1050])|(~m[998]&~m[999]&m[1000]&~m[1001]&~m[1050])|(m[998]&m[999]&~m[1000]&m[1001]&~m[1050])|(m[998]&~m[999]&m[1000]&m[1001]&~m[1050])|(~m[998]&m[999]&m[1000]&m[1001]&~m[1050]))&BiasedRNG[753])|(((m[998]&~m[999]&~m[1000]&~m[1001]&m[1050])|(~m[998]&m[999]&~m[1000]&~m[1001]&m[1050])|(~m[998]&~m[999]&m[1000]&~m[1001]&m[1050])|(m[998]&m[999]&~m[1000]&m[1001]&m[1050])|(m[998]&~m[999]&m[1000]&m[1001]&m[1050])|(~m[998]&m[999]&m[1000]&m[1001]&m[1050]))&~BiasedRNG[753])|((m[998]&m[999]&~m[1000]&~m[1001]&~m[1050])|(m[998]&~m[999]&m[1000]&~m[1001]&~m[1050])|(~m[998]&m[999]&m[1000]&~m[1001]&~m[1050])|(m[998]&m[999]&m[1000]&~m[1001]&~m[1050])|(m[998]&m[999]&m[1000]&m[1001]&~m[1050])|(m[998]&m[999]&~m[1000]&~m[1001]&m[1050])|(m[998]&~m[999]&m[1000]&~m[1001]&m[1050])|(~m[998]&m[999]&m[1000]&~m[1001]&m[1050])|(m[998]&m[999]&m[1000]&~m[1001]&m[1050])|(m[998]&m[999]&m[1000]&m[1001]&m[1050]))):InitCond[1469];
    m[1007] = run?((((m[1003]&~m[1004]&~m[1005]&~m[1006]&~m[1060])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1060])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1060])|(m[1003]&m[1004]&~m[1005]&m[1006]&~m[1060])|(m[1003]&~m[1004]&m[1005]&m[1006]&~m[1060])|(~m[1003]&m[1004]&m[1005]&m[1006]&~m[1060]))&BiasedRNG[754])|(((m[1003]&~m[1004]&~m[1005]&~m[1006]&m[1060])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&m[1060])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&m[1060])|(m[1003]&m[1004]&~m[1005]&m[1006]&m[1060])|(m[1003]&~m[1004]&m[1005]&m[1006]&m[1060])|(~m[1003]&m[1004]&m[1005]&m[1006]&m[1060]))&~BiasedRNG[754])|((m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1060])|(m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1060])|(~m[1003]&m[1004]&m[1005]&~m[1006]&~m[1060])|(m[1003]&m[1004]&m[1005]&~m[1006]&~m[1060])|(m[1003]&m[1004]&m[1005]&m[1006]&~m[1060])|(m[1003]&m[1004]&~m[1005]&~m[1006]&m[1060])|(m[1003]&~m[1004]&m[1005]&~m[1006]&m[1060])|(~m[1003]&m[1004]&m[1005]&~m[1006]&m[1060])|(m[1003]&m[1004]&m[1005]&~m[1006]&m[1060])|(m[1003]&m[1004]&m[1005]&m[1006]&m[1060]))):InitCond[1470];
    m[1012] = run?((((m[1008]&~m[1009]&~m[1010]&~m[1011]&~m[1065])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1065])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1065])|(m[1008]&m[1009]&~m[1010]&m[1011]&~m[1065])|(m[1008]&~m[1009]&m[1010]&m[1011]&~m[1065])|(~m[1008]&m[1009]&m[1010]&m[1011]&~m[1065]))&BiasedRNG[755])|(((m[1008]&~m[1009]&~m[1010]&~m[1011]&m[1065])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&m[1065])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&m[1065])|(m[1008]&m[1009]&~m[1010]&m[1011]&m[1065])|(m[1008]&~m[1009]&m[1010]&m[1011]&m[1065])|(~m[1008]&m[1009]&m[1010]&m[1011]&m[1065]))&~BiasedRNG[755])|((m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1065])|(m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1065])|(~m[1008]&m[1009]&m[1010]&~m[1011]&~m[1065])|(m[1008]&m[1009]&m[1010]&~m[1011]&~m[1065])|(m[1008]&m[1009]&m[1010]&m[1011]&~m[1065])|(m[1008]&m[1009]&~m[1010]&~m[1011]&m[1065])|(m[1008]&~m[1009]&m[1010]&~m[1011]&m[1065])|(~m[1008]&m[1009]&m[1010]&~m[1011]&m[1065])|(m[1008]&m[1009]&m[1010]&~m[1011]&m[1065])|(m[1008]&m[1009]&m[1010]&m[1011]&m[1065]))):InitCond[1471];
    m[1017] = run?((((m[1013]&~m[1014]&~m[1015]&~m[1016]&~m[1070])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1070])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1070])|(m[1013]&m[1014]&~m[1015]&m[1016]&~m[1070])|(m[1013]&~m[1014]&m[1015]&m[1016]&~m[1070])|(~m[1013]&m[1014]&m[1015]&m[1016]&~m[1070]))&BiasedRNG[756])|(((m[1013]&~m[1014]&~m[1015]&~m[1016]&m[1070])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&m[1070])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&m[1070])|(m[1013]&m[1014]&~m[1015]&m[1016]&m[1070])|(m[1013]&~m[1014]&m[1015]&m[1016]&m[1070])|(~m[1013]&m[1014]&m[1015]&m[1016]&m[1070]))&~BiasedRNG[756])|((m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1070])|(m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1070])|(~m[1013]&m[1014]&m[1015]&~m[1016]&~m[1070])|(m[1013]&m[1014]&m[1015]&~m[1016]&~m[1070])|(m[1013]&m[1014]&m[1015]&m[1016]&~m[1070])|(m[1013]&m[1014]&~m[1015]&~m[1016]&m[1070])|(m[1013]&~m[1014]&m[1015]&~m[1016]&m[1070])|(~m[1013]&m[1014]&m[1015]&~m[1016]&m[1070])|(m[1013]&m[1014]&m[1015]&~m[1016]&m[1070])|(m[1013]&m[1014]&m[1015]&m[1016]&m[1070]))):InitCond[1472];
    m[1022] = run?((((m[1018]&~m[1019]&~m[1020]&~m[1021]&~m[1075])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1075])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1075])|(m[1018]&m[1019]&~m[1020]&m[1021]&~m[1075])|(m[1018]&~m[1019]&m[1020]&m[1021]&~m[1075])|(~m[1018]&m[1019]&m[1020]&m[1021]&~m[1075]))&BiasedRNG[757])|(((m[1018]&~m[1019]&~m[1020]&~m[1021]&m[1075])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&m[1075])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&m[1075])|(m[1018]&m[1019]&~m[1020]&m[1021]&m[1075])|(m[1018]&~m[1019]&m[1020]&m[1021]&m[1075])|(~m[1018]&m[1019]&m[1020]&m[1021]&m[1075]))&~BiasedRNG[757])|((m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1075])|(m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1075])|(~m[1018]&m[1019]&m[1020]&~m[1021]&~m[1075])|(m[1018]&m[1019]&m[1020]&~m[1021]&~m[1075])|(m[1018]&m[1019]&m[1020]&m[1021]&~m[1075])|(m[1018]&m[1019]&~m[1020]&~m[1021]&m[1075])|(m[1018]&~m[1019]&m[1020]&~m[1021]&m[1075])|(~m[1018]&m[1019]&m[1020]&~m[1021]&m[1075])|(m[1018]&m[1019]&m[1020]&~m[1021]&m[1075])|(m[1018]&m[1019]&m[1020]&m[1021]&m[1075]))):InitCond[1473];
    m[1027] = run?((((m[1023]&~m[1024]&~m[1025]&~m[1026]&~m[1080])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1080])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1080])|(m[1023]&m[1024]&~m[1025]&m[1026]&~m[1080])|(m[1023]&~m[1024]&m[1025]&m[1026]&~m[1080])|(~m[1023]&m[1024]&m[1025]&m[1026]&~m[1080]))&BiasedRNG[758])|(((m[1023]&~m[1024]&~m[1025]&~m[1026]&m[1080])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&m[1080])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&m[1080])|(m[1023]&m[1024]&~m[1025]&m[1026]&m[1080])|(m[1023]&~m[1024]&m[1025]&m[1026]&m[1080])|(~m[1023]&m[1024]&m[1025]&m[1026]&m[1080]))&~BiasedRNG[758])|((m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1080])|(m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1080])|(~m[1023]&m[1024]&m[1025]&~m[1026]&~m[1080])|(m[1023]&m[1024]&m[1025]&~m[1026]&~m[1080])|(m[1023]&m[1024]&m[1025]&m[1026]&~m[1080])|(m[1023]&m[1024]&~m[1025]&~m[1026]&m[1080])|(m[1023]&~m[1024]&m[1025]&~m[1026]&m[1080])|(~m[1023]&m[1024]&m[1025]&~m[1026]&m[1080])|(m[1023]&m[1024]&m[1025]&~m[1026]&m[1080])|(m[1023]&m[1024]&m[1025]&m[1026]&m[1080]))):InitCond[1474];
    m[1032] = run?((((m[1028]&~m[1029]&~m[1030]&~m[1031]&~m[1085])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1085])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1085])|(m[1028]&m[1029]&~m[1030]&m[1031]&~m[1085])|(m[1028]&~m[1029]&m[1030]&m[1031]&~m[1085])|(~m[1028]&m[1029]&m[1030]&m[1031]&~m[1085]))&BiasedRNG[759])|(((m[1028]&~m[1029]&~m[1030]&~m[1031]&m[1085])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&m[1085])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&m[1085])|(m[1028]&m[1029]&~m[1030]&m[1031]&m[1085])|(m[1028]&~m[1029]&m[1030]&m[1031]&m[1085])|(~m[1028]&m[1029]&m[1030]&m[1031]&m[1085]))&~BiasedRNG[759])|((m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1085])|(m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1085])|(~m[1028]&m[1029]&m[1030]&~m[1031]&~m[1085])|(m[1028]&m[1029]&m[1030]&~m[1031]&~m[1085])|(m[1028]&m[1029]&m[1030]&m[1031]&~m[1085])|(m[1028]&m[1029]&~m[1030]&~m[1031]&m[1085])|(m[1028]&~m[1029]&m[1030]&~m[1031]&m[1085])|(~m[1028]&m[1029]&m[1030]&~m[1031]&m[1085])|(m[1028]&m[1029]&m[1030]&~m[1031]&m[1085])|(m[1028]&m[1029]&m[1030]&m[1031]&m[1085]))):InitCond[1475];
    m[1037] = run?((((m[1033]&~m[1034]&~m[1035]&~m[1036]&~m[1090])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1090])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1090])|(m[1033]&m[1034]&~m[1035]&m[1036]&~m[1090])|(m[1033]&~m[1034]&m[1035]&m[1036]&~m[1090])|(~m[1033]&m[1034]&m[1035]&m[1036]&~m[1090]))&BiasedRNG[760])|(((m[1033]&~m[1034]&~m[1035]&~m[1036]&m[1090])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&m[1090])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&m[1090])|(m[1033]&m[1034]&~m[1035]&m[1036]&m[1090])|(m[1033]&~m[1034]&m[1035]&m[1036]&m[1090])|(~m[1033]&m[1034]&m[1035]&m[1036]&m[1090]))&~BiasedRNG[760])|((m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1090])|(m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1090])|(~m[1033]&m[1034]&m[1035]&~m[1036]&~m[1090])|(m[1033]&m[1034]&m[1035]&~m[1036]&~m[1090])|(m[1033]&m[1034]&m[1035]&m[1036]&~m[1090])|(m[1033]&m[1034]&~m[1035]&~m[1036]&m[1090])|(m[1033]&~m[1034]&m[1035]&~m[1036]&m[1090])|(~m[1033]&m[1034]&m[1035]&~m[1036]&m[1090])|(m[1033]&m[1034]&m[1035]&~m[1036]&m[1090])|(m[1033]&m[1034]&m[1035]&m[1036]&m[1090]))):InitCond[1476];
    m[1042] = run?((((m[1038]&~m[1039]&~m[1040]&~m[1041]&~m[1095])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1095])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1095])|(m[1038]&m[1039]&~m[1040]&m[1041]&~m[1095])|(m[1038]&~m[1039]&m[1040]&m[1041]&~m[1095])|(~m[1038]&m[1039]&m[1040]&m[1041]&~m[1095]))&BiasedRNG[761])|(((m[1038]&~m[1039]&~m[1040]&~m[1041]&m[1095])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&m[1095])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&m[1095])|(m[1038]&m[1039]&~m[1040]&m[1041]&m[1095])|(m[1038]&~m[1039]&m[1040]&m[1041]&m[1095])|(~m[1038]&m[1039]&m[1040]&m[1041]&m[1095]))&~BiasedRNG[761])|((m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1095])|(m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1095])|(~m[1038]&m[1039]&m[1040]&~m[1041]&~m[1095])|(m[1038]&m[1039]&m[1040]&~m[1041]&~m[1095])|(m[1038]&m[1039]&m[1040]&m[1041]&~m[1095])|(m[1038]&m[1039]&~m[1040]&~m[1041]&m[1095])|(m[1038]&~m[1039]&m[1040]&~m[1041]&m[1095])|(~m[1038]&m[1039]&m[1040]&~m[1041]&m[1095])|(m[1038]&m[1039]&m[1040]&~m[1041]&m[1095])|(m[1038]&m[1039]&m[1040]&m[1041]&m[1095]))):InitCond[1477];
    m[1047] = run?((((m[1043]&~m[1044]&~m[1045]&~m[1046]&~m[1100])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1100])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1100])|(m[1043]&m[1044]&~m[1045]&m[1046]&~m[1100])|(m[1043]&~m[1044]&m[1045]&m[1046]&~m[1100])|(~m[1043]&m[1044]&m[1045]&m[1046]&~m[1100]))&BiasedRNG[762])|(((m[1043]&~m[1044]&~m[1045]&~m[1046]&m[1100])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&m[1100])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&m[1100])|(m[1043]&m[1044]&~m[1045]&m[1046]&m[1100])|(m[1043]&~m[1044]&m[1045]&m[1046]&m[1100])|(~m[1043]&m[1044]&m[1045]&m[1046]&m[1100]))&~BiasedRNG[762])|((m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1100])|(m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1100])|(~m[1043]&m[1044]&m[1045]&~m[1046]&~m[1100])|(m[1043]&m[1044]&m[1045]&~m[1046]&~m[1100])|(m[1043]&m[1044]&m[1045]&m[1046]&~m[1100])|(m[1043]&m[1044]&~m[1045]&~m[1046]&m[1100])|(m[1043]&~m[1044]&m[1045]&~m[1046]&m[1100])|(~m[1043]&m[1044]&m[1045]&~m[1046]&m[1100])|(m[1043]&m[1044]&m[1045]&~m[1046]&m[1100])|(m[1043]&m[1044]&m[1045]&m[1046]&m[1100]))):InitCond[1478];
    m[1052] = run?((((m[1048]&~m[1049]&~m[1050]&~m[1051]&~m[1105])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1105])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1105])|(m[1048]&m[1049]&~m[1050]&m[1051]&~m[1105])|(m[1048]&~m[1049]&m[1050]&m[1051]&~m[1105])|(~m[1048]&m[1049]&m[1050]&m[1051]&~m[1105]))&BiasedRNG[763])|(((m[1048]&~m[1049]&~m[1050]&~m[1051]&m[1105])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&m[1105])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&m[1105])|(m[1048]&m[1049]&~m[1050]&m[1051]&m[1105])|(m[1048]&~m[1049]&m[1050]&m[1051]&m[1105])|(~m[1048]&m[1049]&m[1050]&m[1051]&m[1105]))&~BiasedRNG[763])|((m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1105])|(m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1105])|(~m[1048]&m[1049]&m[1050]&~m[1051]&~m[1105])|(m[1048]&m[1049]&m[1050]&~m[1051]&~m[1105])|(m[1048]&m[1049]&m[1050]&m[1051]&~m[1105])|(m[1048]&m[1049]&~m[1050]&~m[1051]&m[1105])|(m[1048]&~m[1049]&m[1050]&~m[1051]&m[1105])|(~m[1048]&m[1049]&m[1050]&~m[1051]&m[1105])|(m[1048]&m[1049]&m[1050]&~m[1051]&m[1105])|(m[1048]&m[1049]&m[1050]&m[1051]&m[1105]))):InitCond[1479];
    m[1057] = run?((((m[1053]&~m[1054]&~m[1055]&~m[1056]&~m[1110])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1110])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1110])|(m[1053]&m[1054]&~m[1055]&m[1056]&~m[1110])|(m[1053]&~m[1054]&m[1055]&m[1056]&~m[1110])|(~m[1053]&m[1054]&m[1055]&m[1056]&~m[1110]))&BiasedRNG[764])|(((m[1053]&~m[1054]&~m[1055]&~m[1056]&m[1110])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&m[1110])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&m[1110])|(m[1053]&m[1054]&~m[1055]&m[1056]&m[1110])|(m[1053]&~m[1054]&m[1055]&m[1056]&m[1110])|(~m[1053]&m[1054]&m[1055]&m[1056]&m[1110]))&~BiasedRNG[764])|((m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1110])|(m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1110])|(~m[1053]&m[1054]&m[1055]&~m[1056]&~m[1110])|(m[1053]&m[1054]&m[1055]&~m[1056]&~m[1110])|(m[1053]&m[1054]&m[1055]&m[1056]&~m[1110])|(m[1053]&m[1054]&~m[1055]&~m[1056]&m[1110])|(m[1053]&~m[1054]&m[1055]&~m[1056]&m[1110])|(~m[1053]&m[1054]&m[1055]&~m[1056]&m[1110])|(m[1053]&m[1054]&m[1055]&~m[1056]&m[1110])|(m[1053]&m[1054]&m[1055]&m[1056]&m[1110]))):InitCond[1480];
    m[1062] = run?((((m[1058]&~m[1059]&~m[1060]&~m[1061]&~m[1120])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1120])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1120])|(m[1058]&m[1059]&~m[1060]&m[1061]&~m[1120])|(m[1058]&~m[1059]&m[1060]&m[1061]&~m[1120])|(~m[1058]&m[1059]&m[1060]&m[1061]&~m[1120]))&BiasedRNG[765])|(((m[1058]&~m[1059]&~m[1060]&~m[1061]&m[1120])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&m[1120])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&m[1120])|(m[1058]&m[1059]&~m[1060]&m[1061]&m[1120])|(m[1058]&~m[1059]&m[1060]&m[1061]&m[1120])|(~m[1058]&m[1059]&m[1060]&m[1061]&m[1120]))&~BiasedRNG[765])|((m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1120])|(m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1120])|(~m[1058]&m[1059]&m[1060]&~m[1061]&~m[1120])|(m[1058]&m[1059]&m[1060]&~m[1061]&~m[1120])|(m[1058]&m[1059]&m[1060]&m[1061]&~m[1120])|(m[1058]&m[1059]&~m[1060]&~m[1061]&m[1120])|(m[1058]&~m[1059]&m[1060]&~m[1061]&m[1120])|(~m[1058]&m[1059]&m[1060]&~m[1061]&m[1120])|(m[1058]&m[1059]&m[1060]&~m[1061]&m[1120])|(m[1058]&m[1059]&m[1060]&m[1061]&m[1120]))):InitCond[1481];
    m[1067] = run?((((m[1063]&~m[1064]&~m[1065]&~m[1066]&~m[1125])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1125])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1125])|(m[1063]&m[1064]&~m[1065]&m[1066]&~m[1125])|(m[1063]&~m[1064]&m[1065]&m[1066]&~m[1125])|(~m[1063]&m[1064]&m[1065]&m[1066]&~m[1125]))&BiasedRNG[766])|(((m[1063]&~m[1064]&~m[1065]&~m[1066]&m[1125])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&m[1125])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&m[1125])|(m[1063]&m[1064]&~m[1065]&m[1066]&m[1125])|(m[1063]&~m[1064]&m[1065]&m[1066]&m[1125])|(~m[1063]&m[1064]&m[1065]&m[1066]&m[1125]))&~BiasedRNG[766])|((m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1125])|(m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1125])|(~m[1063]&m[1064]&m[1065]&~m[1066]&~m[1125])|(m[1063]&m[1064]&m[1065]&~m[1066]&~m[1125])|(m[1063]&m[1064]&m[1065]&m[1066]&~m[1125])|(m[1063]&m[1064]&~m[1065]&~m[1066]&m[1125])|(m[1063]&~m[1064]&m[1065]&~m[1066]&m[1125])|(~m[1063]&m[1064]&m[1065]&~m[1066]&m[1125])|(m[1063]&m[1064]&m[1065]&~m[1066]&m[1125])|(m[1063]&m[1064]&m[1065]&m[1066]&m[1125]))):InitCond[1482];
    m[1072] = run?((((m[1068]&~m[1069]&~m[1070]&~m[1071]&~m[1130])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1130])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1130])|(m[1068]&m[1069]&~m[1070]&m[1071]&~m[1130])|(m[1068]&~m[1069]&m[1070]&m[1071]&~m[1130])|(~m[1068]&m[1069]&m[1070]&m[1071]&~m[1130]))&BiasedRNG[767])|(((m[1068]&~m[1069]&~m[1070]&~m[1071]&m[1130])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&m[1130])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&m[1130])|(m[1068]&m[1069]&~m[1070]&m[1071]&m[1130])|(m[1068]&~m[1069]&m[1070]&m[1071]&m[1130])|(~m[1068]&m[1069]&m[1070]&m[1071]&m[1130]))&~BiasedRNG[767])|((m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1130])|(m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1130])|(~m[1068]&m[1069]&m[1070]&~m[1071]&~m[1130])|(m[1068]&m[1069]&m[1070]&~m[1071]&~m[1130])|(m[1068]&m[1069]&m[1070]&m[1071]&~m[1130])|(m[1068]&m[1069]&~m[1070]&~m[1071]&m[1130])|(m[1068]&~m[1069]&m[1070]&~m[1071]&m[1130])|(~m[1068]&m[1069]&m[1070]&~m[1071]&m[1130])|(m[1068]&m[1069]&m[1070]&~m[1071]&m[1130])|(m[1068]&m[1069]&m[1070]&m[1071]&m[1130]))):InitCond[1483];
    m[1077] = run?((((m[1073]&~m[1074]&~m[1075]&~m[1076]&~m[1135])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1135])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1135])|(m[1073]&m[1074]&~m[1075]&m[1076]&~m[1135])|(m[1073]&~m[1074]&m[1075]&m[1076]&~m[1135])|(~m[1073]&m[1074]&m[1075]&m[1076]&~m[1135]))&BiasedRNG[768])|(((m[1073]&~m[1074]&~m[1075]&~m[1076]&m[1135])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&m[1135])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&m[1135])|(m[1073]&m[1074]&~m[1075]&m[1076]&m[1135])|(m[1073]&~m[1074]&m[1075]&m[1076]&m[1135])|(~m[1073]&m[1074]&m[1075]&m[1076]&m[1135]))&~BiasedRNG[768])|((m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1135])|(m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1135])|(~m[1073]&m[1074]&m[1075]&~m[1076]&~m[1135])|(m[1073]&m[1074]&m[1075]&~m[1076]&~m[1135])|(m[1073]&m[1074]&m[1075]&m[1076]&~m[1135])|(m[1073]&m[1074]&~m[1075]&~m[1076]&m[1135])|(m[1073]&~m[1074]&m[1075]&~m[1076]&m[1135])|(~m[1073]&m[1074]&m[1075]&~m[1076]&m[1135])|(m[1073]&m[1074]&m[1075]&~m[1076]&m[1135])|(m[1073]&m[1074]&m[1075]&m[1076]&m[1135]))):InitCond[1484];
    m[1082] = run?((((m[1078]&~m[1079]&~m[1080]&~m[1081]&~m[1140])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1140])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1140])|(m[1078]&m[1079]&~m[1080]&m[1081]&~m[1140])|(m[1078]&~m[1079]&m[1080]&m[1081]&~m[1140])|(~m[1078]&m[1079]&m[1080]&m[1081]&~m[1140]))&BiasedRNG[769])|(((m[1078]&~m[1079]&~m[1080]&~m[1081]&m[1140])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&m[1140])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&m[1140])|(m[1078]&m[1079]&~m[1080]&m[1081]&m[1140])|(m[1078]&~m[1079]&m[1080]&m[1081]&m[1140])|(~m[1078]&m[1079]&m[1080]&m[1081]&m[1140]))&~BiasedRNG[769])|((m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1140])|(m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1140])|(~m[1078]&m[1079]&m[1080]&~m[1081]&~m[1140])|(m[1078]&m[1079]&m[1080]&~m[1081]&~m[1140])|(m[1078]&m[1079]&m[1080]&m[1081]&~m[1140])|(m[1078]&m[1079]&~m[1080]&~m[1081]&m[1140])|(m[1078]&~m[1079]&m[1080]&~m[1081]&m[1140])|(~m[1078]&m[1079]&m[1080]&~m[1081]&m[1140])|(m[1078]&m[1079]&m[1080]&~m[1081]&m[1140])|(m[1078]&m[1079]&m[1080]&m[1081]&m[1140]))):InitCond[1485];
    m[1087] = run?((((m[1083]&~m[1084]&~m[1085]&~m[1086]&~m[1145])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1145])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1145])|(m[1083]&m[1084]&~m[1085]&m[1086]&~m[1145])|(m[1083]&~m[1084]&m[1085]&m[1086]&~m[1145])|(~m[1083]&m[1084]&m[1085]&m[1086]&~m[1145]))&BiasedRNG[770])|(((m[1083]&~m[1084]&~m[1085]&~m[1086]&m[1145])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&m[1145])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&m[1145])|(m[1083]&m[1084]&~m[1085]&m[1086]&m[1145])|(m[1083]&~m[1084]&m[1085]&m[1086]&m[1145])|(~m[1083]&m[1084]&m[1085]&m[1086]&m[1145]))&~BiasedRNG[770])|((m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1145])|(m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1145])|(~m[1083]&m[1084]&m[1085]&~m[1086]&~m[1145])|(m[1083]&m[1084]&m[1085]&~m[1086]&~m[1145])|(m[1083]&m[1084]&m[1085]&m[1086]&~m[1145])|(m[1083]&m[1084]&~m[1085]&~m[1086]&m[1145])|(m[1083]&~m[1084]&m[1085]&~m[1086]&m[1145])|(~m[1083]&m[1084]&m[1085]&~m[1086]&m[1145])|(m[1083]&m[1084]&m[1085]&~m[1086]&m[1145])|(m[1083]&m[1084]&m[1085]&m[1086]&m[1145]))):InitCond[1486];
    m[1092] = run?((((m[1088]&~m[1089]&~m[1090]&~m[1091]&~m[1150])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1150])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1150])|(m[1088]&m[1089]&~m[1090]&m[1091]&~m[1150])|(m[1088]&~m[1089]&m[1090]&m[1091]&~m[1150])|(~m[1088]&m[1089]&m[1090]&m[1091]&~m[1150]))&BiasedRNG[771])|(((m[1088]&~m[1089]&~m[1090]&~m[1091]&m[1150])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&m[1150])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&m[1150])|(m[1088]&m[1089]&~m[1090]&m[1091]&m[1150])|(m[1088]&~m[1089]&m[1090]&m[1091]&m[1150])|(~m[1088]&m[1089]&m[1090]&m[1091]&m[1150]))&~BiasedRNG[771])|((m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1150])|(m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1150])|(~m[1088]&m[1089]&m[1090]&~m[1091]&~m[1150])|(m[1088]&m[1089]&m[1090]&~m[1091]&~m[1150])|(m[1088]&m[1089]&m[1090]&m[1091]&~m[1150])|(m[1088]&m[1089]&~m[1090]&~m[1091]&m[1150])|(m[1088]&~m[1089]&m[1090]&~m[1091]&m[1150])|(~m[1088]&m[1089]&m[1090]&~m[1091]&m[1150])|(m[1088]&m[1089]&m[1090]&~m[1091]&m[1150])|(m[1088]&m[1089]&m[1090]&m[1091]&m[1150]))):InitCond[1487];
    m[1097] = run?((((m[1093]&~m[1094]&~m[1095]&~m[1096]&~m[1155])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1155])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1155])|(m[1093]&m[1094]&~m[1095]&m[1096]&~m[1155])|(m[1093]&~m[1094]&m[1095]&m[1096]&~m[1155])|(~m[1093]&m[1094]&m[1095]&m[1096]&~m[1155]))&BiasedRNG[772])|(((m[1093]&~m[1094]&~m[1095]&~m[1096]&m[1155])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&m[1155])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&m[1155])|(m[1093]&m[1094]&~m[1095]&m[1096]&m[1155])|(m[1093]&~m[1094]&m[1095]&m[1096]&m[1155])|(~m[1093]&m[1094]&m[1095]&m[1096]&m[1155]))&~BiasedRNG[772])|((m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1155])|(m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1155])|(~m[1093]&m[1094]&m[1095]&~m[1096]&~m[1155])|(m[1093]&m[1094]&m[1095]&~m[1096]&~m[1155])|(m[1093]&m[1094]&m[1095]&m[1096]&~m[1155])|(m[1093]&m[1094]&~m[1095]&~m[1096]&m[1155])|(m[1093]&~m[1094]&m[1095]&~m[1096]&m[1155])|(~m[1093]&m[1094]&m[1095]&~m[1096]&m[1155])|(m[1093]&m[1094]&m[1095]&~m[1096]&m[1155])|(m[1093]&m[1094]&m[1095]&m[1096]&m[1155]))):InitCond[1488];
    m[1102] = run?((((m[1098]&~m[1099]&~m[1100]&~m[1101]&~m[1160])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1160])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1160])|(m[1098]&m[1099]&~m[1100]&m[1101]&~m[1160])|(m[1098]&~m[1099]&m[1100]&m[1101]&~m[1160])|(~m[1098]&m[1099]&m[1100]&m[1101]&~m[1160]))&BiasedRNG[773])|(((m[1098]&~m[1099]&~m[1100]&~m[1101]&m[1160])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&m[1160])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&m[1160])|(m[1098]&m[1099]&~m[1100]&m[1101]&m[1160])|(m[1098]&~m[1099]&m[1100]&m[1101]&m[1160])|(~m[1098]&m[1099]&m[1100]&m[1101]&m[1160]))&~BiasedRNG[773])|((m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1160])|(m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1160])|(~m[1098]&m[1099]&m[1100]&~m[1101]&~m[1160])|(m[1098]&m[1099]&m[1100]&~m[1101]&~m[1160])|(m[1098]&m[1099]&m[1100]&m[1101]&~m[1160])|(m[1098]&m[1099]&~m[1100]&~m[1101]&m[1160])|(m[1098]&~m[1099]&m[1100]&~m[1101]&m[1160])|(~m[1098]&m[1099]&m[1100]&~m[1101]&m[1160])|(m[1098]&m[1099]&m[1100]&~m[1101]&m[1160])|(m[1098]&m[1099]&m[1100]&m[1101]&m[1160]))):InitCond[1489];
    m[1107] = run?((((m[1103]&~m[1104]&~m[1105]&~m[1106]&~m[1165])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1165])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1165])|(m[1103]&m[1104]&~m[1105]&m[1106]&~m[1165])|(m[1103]&~m[1104]&m[1105]&m[1106]&~m[1165])|(~m[1103]&m[1104]&m[1105]&m[1106]&~m[1165]))&BiasedRNG[774])|(((m[1103]&~m[1104]&~m[1105]&~m[1106]&m[1165])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&m[1165])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&m[1165])|(m[1103]&m[1104]&~m[1105]&m[1106]&m[1165])|(m[1103]&~m[1104]&m[1105]&m[1106]&m[1165])|(~m[1103]&m[1104]&m[1105]&m[1106]&m[1165]))&~BiasedRNG[774])|((m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1165])|(m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1165])|(~m[1103]&m[1104]&m[1105]&~m[1106]&~m[1165])|(m[1103]&m[1104]&m[1105]&~m[1106]&~m[1165])|(m[1103]&m[1104]&m[1105]&m[1106]&~m[1165])|(m[1103]&m[1104]&~m[1105]&~m[1106]&m[1165])|(m[1103]&~m[1104]&m[1105]&~m[1106]&m[1165])|(~m[1103]&m[1104]&m[1105]&~m[1106]&m[1165])|(m[1103]&m[1104]&m[1105]&~m[1106]&m[1165])|(m[1103]&m[1104]&m[1105]&m[1106]&m[1165]))):InitCond[1490];
    m[1112] = run?((((m[1108]&~m[1109]&~m[1110]&~m[1111]&~m[1170])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1170])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1170])|(m[1108]&m[1109]&~m[1110]&m[1111]&~m[1170])|(m[1108]&~m[1109]&m[1110]&m[1111]&~m[1170])|(~m[1108]&m[1109]&m[1110]&m[1111]&~m[1170]))&BiasedRNG[775])|(((m[1108]&~m[1109]&~m[1110]&~m[1111]&m[1170])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&m[1170])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&m[1170])|(m[1108]&m[1109]&~m[1110]&m[1111]&m[1170])|(m[1108]&~m[1109]&m[1110]&m[1111]&m[1170])|(~m[1108]&m[1109]&m[1110]&m[1111]&m[1170]))&~BiasedRNG[775])|((m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1170])|(m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1170])|(~m[1108]&m[1109]&m[1110]&~m[1111]&~m[1170])|(m[1108]&m[1109]&m[1110]&~m[1111]&~m[1170])|(m[1108]&m[1109]&m[1110]&m[1111]&~m[1170])|(m[1108]&m[1109]&~m[1110]&~m[1111]&m[1170])|(m[1108]&~m[1109]&m[1110]&~m[1111]&m[1170])|(~m[1108]&m[1109]&m[1110]&~m[1111]&m[1170])|(m[1108]&m[1109]&m[1110]&~m[1111]&m[1170])|(m[1108]&m[1109]&m[1110]&m[1111]&m[1170]))):InitCond[1491];
    m[1117] = run?((((m[1113]&~m[1114]&~m[1115]&~m[1116]&~m[1175])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1175])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1175])|(m[1113]&m[1114]&~m[1115]&m[1116]&~m[1175])|(m[1113]&~m[1114]&m[1115]&m[1116]&~m[1175])|(~m[1113]&m[1114]&m[1115]&m[1116]&~m[1175]))&BiasedRNG[776])|(((m[1113]&~m[1114]&~m[1115]&~m[1116]&m[1175])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&m[1175])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&m[1175])|(m[1113]&m[1114]&~m[1115]&m[1116]&m[1175])|(m[1113]&~m[1114]&m[1115]&m[1116]&m[1175])|(~m[1113]&m[1114]&m[1115]&m[1116]&m[1175]))&~BiasedRNG[776])|((m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1175])|(m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1175])|(~m[1113]&m[1114]&m[1115]&~m[1116]&~m[1175])|(m[1113]&m[1114]&m[1115]&~m[1116]&~m[1175])|(m[1113]&m[1114]&m[1115]&m[1116]&~m[1175])|(m[1113]&m[1114]&~m[1115]&~m[1116]&m[1175])|(m[1113]&~m[1114]&m[1115]&~m[1116]&m[1175])|(~m[1113]&m[1114]&m[1115]&~m[1116]&m[1175])|(m[1113]&m[1114]&m[1115]&~m[1116]&m[1175])|(m[1113]&m[1114]&m[1115]&m[1116]&m[1175]))):InitCond[1492];
    m[1122] = run?((((m[1118]&~m[1119]&~m[1120]&~m[1121]&~m[1185])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1185])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1185])|(m[1118]&m[1119]&~m[1120]&m[1121]&~m[1185])|(m[1118]&~m[1119]&m[1120]&m[1121]&~m[1185])|(~m[1118]&m[1119]&m[1120]&m[1121]&~m[1185]))&BiasedRNG[777])|(((m[1118]&~m[1119]&~m[1120]&~m[1121]&m[1185])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&m[1185])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&m[1185])|(m[1118]&m[1119]&~m[1120]&m[1121]&m[1185])|(m[1118]&~m[1119]&m[1120]&m[1121]&m[1185])|(~m[1118]&m[1119]&m[1120]&m[1121]&m[1185]))&~BiasedRNG[777])|((m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1185])|(m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1185])|(~m[1118]&m[1119]&m[1120]&~m[1121]&~m[1185])|(m[1118]&m[1119]&m[1120]&~m[1121]&~m[1185])|(m[1118]&m[1119]&m[1120]&m[1121]&~m[1185])|(m[1118]&m[1119]&~m[1120]&~m[1121]&m[1185])|(m[1118]&~m[1119]&m[1120]&~m[1121]&m[1185])|(~m[1118]&m[1119]&m[1120]&~m[1121]&m[1185])|(m[1118]&m[1119]&m[1120]&~m[1121]&m[1185])|(m[1118]&m[1119]&m[1120]&m[1121]&m[1185]))):InitCond[1493];
    m[1127] = run?((((m[1123]&~m[1124]&~m[1125]&~m[1126]&~m[1190])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1190])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1190])|(m[1123]&m[1124]&~m[1125]&m[1126]&~m[1190])|(m[1123]&~m[1124]&m[1125]&m[1126]&~m[1190])|(~m[1123]&m[1124]&m[1125]&m[1126]&~m[1190]))&BiasedRNG[778])|(((m[1123]&~m[1124]&~m[1125]&~m[1126]&m[1190])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&m[1190])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&m[1190])|(m[1123]&m[1124]&~m[1125]&m[1126]&m[1190])|(m[1123]&~m[1124]&m[1125]&m[1126]&m[1190])|(~m[1123]&m[1124]&m[1125]&m[1126]&m[1190]))&~BiasedRNG[778])|((m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1190])|(m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1190])|(~m[1123]&m[1124]&m[1125]&~m[1126]&~m[1190])|(m[1123]&m[1124]&m[1125]&~m[1126]&~m[1190])|(m[1123]&m[1124]&m[1125]&m[1126]&~m[1190])|(m[1123]&m[1124]&~m[1125]&~m[1126]&m[1190])|(m[1123]&~m[1124]&m[1125]&~m[1126]&m[1190])|(~m[1123]&m[1124]&m[1125]&~m[1126]&m[1190])|(m[1123]&m[1124]&m[1125]&~m[1126]&m[1190])|(m[1123]&m[1124]&m[1125]&m[1126]&m[1190]))):InitCond[1494];
    m[1132] = run?((((m[1128]&~m[1129]&~m[1130]&~m[1131]&~m[1195])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1195])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1195])|(m[1128]&m[1129]&~m[1130]&m[1131]&~m[1195])|(m[1128]&~m[1129]&m[1130]&m[1131]&~m[1195])|(~m[1128]&m[1129]&m[1130]&m[1131]&~m[1195]))&BiasedRNG[779])|(((m[1128]&~m[1129]&~m[1130]&~m[1131]&m[1195])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&m[1195])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&m[1195])|(m[1128]&m[1129]&~m[1130]&m[1131]&m[1195])|(m[1128]&~m[1129]&m[1130]&m[1131]&m[1195])|(~m[1128]&m[1129]&m[1130]&m[1131]&m[1195]))&~BiasedRNG[779])|((m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1195])|(m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1195])|(~m[1128]&m[1129]&m[1130]&~m[1131]&~m[1195])|(m[1128]&m[1129]&m[1130]&~m[1131]&~m[1195])|(m[1128]&m[1129]&m[1130]&m[1131]&~m[1195])|(m[1128]&m[1129]&~m[1130]&~m[1131]&m[1195])|(m[1128]&~m[1129]&m[1130]&~m[1131]&m[1195])|(~m[1128]&m[1129]&m[1130]&~m[1131]&m[1195])|(m[1128]&m[1129]&m[1130]&~m[1131]&m[1195])|(m[1128]&m[1129]&m[1130]&m[1131]&m[1195]))):InitCond[1495];
    m[1137] = run?((((m[1133]&~m[1134]&~m[1135]&~m[1136]&~m[1200])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1200])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1200])|(m[1133]&m[1134]&~m[1135]&m[1136]&~m[1200])|(m[1133]&~m[1134]&m[1135]&m[1136]&~m[1200])|(~m[1133]&m[1134]&m[1135]&m[1136]&~m[1200]))&BiasedRNG[780])|(((m[1133]&~m[1134]&~m[1135]&~m[1136]&m[1200])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&m[1200])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&m[1200])|(m[1133]&m[1134]&~m[1135]&m[1136]&m[1200])|(m[1133]&~m[1134]&m[1135]&m[1136]&m[1200])|(~m[1133]&m[1134]&m[1135]&m[1136]&m[1200]))&~BiasedRNG[780])|((m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1200])|(m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1200])|(~m[1133]&m[1134]&m[1135]&~m[1136]&~m[1200])|(m[1133]&m[1134]&m[1135]&~m[1136]&~m[1200])|(m[1133]&m[1134]&m[1135]&m[1136]&~m[1200])|(m[1133]&m[1134]&~m[1135]&~m[1136]&m[1200])|(m[1133]&~m[1134]&m[1135]&~m[1136]&m[1200])|(~m[1133]&m[1134]&m[1135]&~m[1136]&m[1200])|(m[1133]&m[1134]&m[1135]&~m[1136]&m[1200])|(m[1133]&m[1134]&m[1135]&m[1136]&m[1200]))):InitCond[1496];
    m[1142] = run?((((m[1138]&~m[1139]&~m[1140]&~m[1141]&~m[1205])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1205])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1205])|(m[1138]&m[1139]&~m[1140]&m[1141]&~m[1205])|(m[1138]&~m[1139]&m[1140]&m[1141]&~m[1205])|(~m[1138]&m[1139]&m[1140]&m[1141]&~m[1205]))&BiasedRNG[781])|(((m[1138]&~m[1139]&~m[1140]&~m[1141]&m[1205])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&m[1205])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&m[1205])|(m[1138]&m[1139]&~m[1140]&m[1141]&m[1205])|(m[1138]&~m[1139]&m[1140]&m[1141]&m[1205])|(~m[1138]&m[1139]&m[1140]&m[1141]&m[1205]))&~BiasedRNG[781])|((m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1205])|(m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1205])|(~m[1138]&m[1139]&m[1140]&~m[1141]&~m[1205])|(m[1138]&m[1139]&m[1140]&~m[1141]&~m[1205])|(m[1138]&m[1139]&m[1140]&m[1141]&~m[1205])|(m[1138]&m[1139]&~m[1140]&~m[1141]&m[1205])|(m[1138]&~m[1139]&m[1140]&~m[1141]&m[1205])|(~m[1138]&m[1139]&m[1140]&~m[1141]&m[1205])|(m[1138]&m[1139]&m[1140]&~m[1141]&m[1205])|(m[1138]&m[1139]&m[1140]&m[1141]&m[1205]))):InitCond[1497];
    m[1147] = run?((((m[1143]&~m[1144]&~m[1145]&~m[1146]&~m[1210])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1210])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1210])|(m[1143]&m[1144]&~m[1145]&m[1146]&~m[1210])|(m[1143]&~m[1144]&m[1145]&m[1146]&~m[1210])|(~m[1143]&m[1144]&m[1145]&m[1146]&~m[1210]))&BiasedRNG[782])|(((m[1143]&~m[1144]&~m[1145]&~m[1146]&m[1210])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&m[1210])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&m[1210])|(m[1143]&m[1144]&~m[1145]&m[1146]&m[1210])|(m[1143]&~m[1144]&m[1145]&m[1146]&m[1210])|(~m[1143]&m[1144]&m[1145]&m[1146]&m[1210]))&~BiasedRNG[782])|((m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1210])|(m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1210])|(~m[1143]&m[1144]&m[1145]&~m[1146]&~m[1210])|(m[1143]&m[1144]&m[1145]&~m[1146]&~m[1210])|(m[1143]&m[1144]&m[1145]&m[1146]&~m[1210])|(m[1143]&m[1144]&~m[1145]&~m[1146]&m[1210])|(m[1143]&~m[1144]&m[1145]&~m[1146]&m[1210])|(~m[1143]&m[1144]&m[1145]&~m[1146]&m[1210])|(m[1143]&m[1144]&m[1145]&~m[1146]&m[1210])|(m[1143]&m[1144]&m[1145]&m[1146]&m[1210]))):InitCond[1498];
    m[1152] = run?((((m[1148]&~m[1149]&~m[1150]&~m[1151]&~m[1215])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1215])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1215])|(m[1148]&m[1149]&~m[1150]&m[1151]&~m[1215])|(m[1148]&~m[1149]&m[1150]&m[1151]&~m[1215])|(~m[1148]&m[1149]&m[1150]&m[1151]&~m[1215]))&BiasedRNG[783])|(((m[1148]&~m[1149]&~m[1150]&~m[1151]&m[1215])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&m[1215])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&m[1215])|(m[1148]&m[1149]&~m[1150]&m[1151]&m[1215])|(m[1148]&~m[1149]&m[1150]&m[1151]&m[1215])|(~m[1148]&m[1149]&m[1150]&m[1151]&m[1215]))&~BiasedRNG[783])|((m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1215])|(m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1215])|(~m[1148]&m[1149]&m[1150]&~m[1151]&~m[1215])|(m[1148]&m[1149]&m[1150]&~m[1151]&~m[1215])|(m[1148]&m[1149]&m[1150]&m[1151]&~m[1215])|(m[1148]&m[1149]&~m[1150]&~m[1151]&m[1215])|(m[1148]&~m[1149]&m[1150]&~m[1151]&m[1215])|(~m[1148]&m[1149]&m[1150]&~m[1151]&m[1215])|(m[1148]&m[1149]&m[1150]&~m[1151]&m[1215])|(m[1148]&m[1149]&m[1150]&m[1151]&m[1215]))):InitCond[1499];
    m[1157] = run?((((m[1153]&~m[1154]&~m[1155]&~m[1156]&~m[1220])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1220])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1220])|(m[1153]&m[1154]&~m[1155]&m[1156]&~m[1220])|(m[1153]&~m[1154]&m[1155]&m[1156]&~m[1220])|(~m[1153]&m[1154]&m[1155]&m[1156]&~m[1220]))&BiasedRNG[784])|(((m[1153]&~m[1154]&~m[1155]&~m[1156]&m[1220])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&m[1220])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&m[1220])|(m[1153]&m[1154]&~m[1155]&m[1156]&m[1220])|(m[1153]&~m[1154]&m[1155]&m[1156]&m[1220])|(~m[1153]&m[1154]&m[1155]&m[1156]&m[1220]))&~BiasedRNG[784])|((m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1220])|(m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1220])|(~m[1153]&m[1154]&m[1155]&~m[1156]&~m[1220])|(m[1153]&m[1154]&m[1155]&~m[1156]&~m[1220])|(m[1153]&m[1154]&m[1155]&m[1156]&~m[1220])|(m[1153]&m[1154]&~m[1155]&~m[1156]&m[1220])|(m[1153]&~m[1154]&m[1155]&~m[1156]&m[1220])|(~m[1153]&m[1154]&m[1155]&~m[1156]&m[1220])|(m[1153]&m[1154]&m[1155]&~m[1156]&m[1220])|(m[1153]&m[1154]&m[1155]&m[1156]&m[1220]))):InitCond[1500];
    m[1162] = run?((((m[1158]&~m[1159]&~m[1160]&~m[1161]&~m[1225])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1225])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1225])|(m[1158]&m[1159]&~m[1160]&m[1161]&~m[1225])|(m[1158]&~m[1159]&m[1160]&m[1161]&~m[1225])|(~m[1158]&m[1159]&m[1160]&m[1161]&~m[1225]))&BiasedRNG[785])|(((m[1158]&~m[1159]&~m[1160]&~m[1161]&m[1225])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&m[1225])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&m[1225])|(m[1158]&m[1159]&~m[1160]&m[1161]&m[1225])|(m[1158]&~m[1159]&m[1160]&m[1161]&m[1225])|(~m[1158]&m[1159]&m[1160]&m[1161]&m[1225]))&~BiasedRNG[785])|((m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1225])|(m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1225])|(~m[1158]&m[1159]&m[1160]&~m[1161]&~m[1225])|(m[1158]&m[1159]&m[1160]&~m[1161]&~m[1225])|(m[1158]&m[1159]&m[1160]&m[1161]&~m[1225])|(m[1158]&m[1159]&~m[1160]&~m[1161]&m[1225])|(m[1158]&~m[1159]&m[1160]&~m[1161]&m[1225])|(~m[1158]&m[1159]&m[1160]&~m[1161]&m[1225])|(m[1158]&m[1159]&m[1160]&~m[1161]&m[1225])|(m[1158]&m[1159]&m[1160]&m[1161]&m[1225]))):InitCond[1501];
    m[1167] = run?((((m[1163]&~m[1164]&~m[1165]&~m[1166]&~m[1230])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1230])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1230])|(m[1163]&m[1164]&~m[1165]&m[1166]&~m[1230])|(m[1163]&~m[1164]&m[1165]&m[1166]&~m[1230])|(~m[1163]&m[1164]&m[1165]&m[1166]&~m[1230]))&BiasedRNG[786])|(((m[1163]&~m[1164]&~m[1165]&~m[1166]&m[1230])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&m[1230])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&m[1230])|(m[1163]&m[1164]&~m[1165]&m[1166]&m[1230])|(m[1163]&~m[1164]&m[1165]&m[1166]&m[1230])|(~m[1163]&m[1164]&m[1165]&m[1166]&m[1230]))&~BiasedRNG[786])|((m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1230])|(m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1230])|(~m[1163]&m[1164]&m[1165]&~m[1166]&~m[1230])|(m[1163]&m[1164]&m[1165]&~m[1166]&~m[1230])|(m[1163]&m[1164]&m[1165]&m[1166]&~m[1230])|(m[1163]&m[1164]&~m[1165]&~m[1166]&m[1230])|(m[1163]&~m[1164]&m[1165]&~m[1166]&m[1230])|(~m[1163]&m[1164]&m[1165]&~m[1166]&m[1230])|(m[1163]&m[1164]&m[1165]&~m[1166]&m[1230])|(m[1163]&m[1164]&m[1165]&m[1166]&m[1230]))):InitCond[1502];
    m[1172] = run?((((m[1168]&~m[1169]&~m[1170]&~m[1171]&~m[1235])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1235])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1235])|(m[1168]&m[1169]&~m[1170]&m[1171]&~m[1235])|(m[1168]&~m[1169]&m[1170]&m[1171]&~m[1235])|(~m[1168]&m[1169]&m[1170]&m[1171]&~m[1235]))&BiasedRNG[787])|(((m[1168]&~m[1169]&~m[1170]&~m[1171]&m[1235])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&m[1235])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&m[1235])|(m[1168]&m[1169]&~m[1170]&m[1171]&m[1235])|(m[1168]&~m[1169]&m[1170]&m[1171]&m[1235])|(~m[1168]&m[1169]&m[1170]&m[1171]&m[1235]))&~BiasedRNG[787])|((m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1235])|(m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1235])|(~m[1168]&m[1169]&m[1170]&~m[1171]&~m[1235])|(m[1168]&m[1169]&m[1170]&~m[1171]&~m[1235])|(m[1168]&m[1169]&m[1170]&m[1171]&~m[1235])|(m[1168]&m[1169]&~m[1170]&~m[1171]&m[1235])|(m[1168]&~m[1169]&m[1170]&~m[1171]&m[1235])|(~m[1168]&m[1169]&m[1170]&~m[1171]&m[1235])|(m[1168]&m[1169]&m[1170]&~m[1171]&m[1235])|(m[1168]&m[1169]&m[1170]&m[1171]&m[1235]))):InitCond[1503];
    m[1177] = run?((((m[1173]&~m[1174]&~m[1175]&~m[1176]&~m[1240])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1240])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1240])|(m[1173]&m[1174]&~m[1175]&m[1176]&~m[1240])|(m[1173]&~m[1174]&m[1175]&m[1176]&~m[1240])|(~m[1173]&m[1174]&m[1175]&m[1176]&~m[1240]))&BiasedRNG[788])|(((m[1173]&~m[1174]&~m[1175]&~m[1176]&m[1240])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&m[1240])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&m[1240])|(m[1173]&m[1174]&~m[1175]&m[1176]&m[1240])|(m[1173]&~m[1174]&m[1175]&m[1176]&m[1240])|(~m[1173]&m[1174]&m[1175]&m[1176]&m[1240]))&~BiasedRNG[788])|((m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1240])|(m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1240])|(~m[1173]&m[1174]&m[1175]&~m[1176]&~m[1240])|(m[1173]&m[1174]&m[1175]&~m[1176]&~m[1240])|(m[1173]&m[1174]&m[1175]&m[1176]&~m[1240])|(m[1173]&m[1174]&~m[1175]&~m[1176]&m[1240])|(m[1173]&~m[1174]&m[1175]&~m[1176]&m[1240])|(~m[1173]&m[1174]&m[1175]&~m[1176]&m[1240])|(m[1173]&m[1174]&m[1175]&~m[1176]&m[1240])|(m[1173]&m[1174]&m[1175]&m[1176]&m[1240]))):InitCond[1504];
    m[1182] = run?((((m[1178]&~m[1179]&~m[1180]&~m[1181]&~m[1245])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1245])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1245])|(m[1178]&m[1179]&~m[1180]&m[1181]&~m[1245])|(m[1178]&~m[1179]&m[1180]&m[1181]&~m[1245])|(~m[1178]&m[1179]&m[1180]&m[1181]&~m[1245]))&BiasedRNG[789])|(((m[1178]&~m[1179]&~m[1180]&~m[1181]&m[1245])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&m[1245])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&m[1245])|(m[1178]&m[1179]&~m[1180]&m[1181]&m[1245])|(m[1178]&~m[1179]&m[1180]&m[1181]&m[1245])|(~m[1178]&m[1179]&m[1180]&m[1181]&m[1245]))&~BiasedRNG[789])|((m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1245])|(m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1245])|(~m[1178]&m[1179]&m[1180]&~m[1181]&~m[1245])|(m[1178]&m[1179]&m[1180]&~m[1181]&~m[1245])|(m[1178]&m[1179]&m[1180]&m[1181]&~m[1245])|(m[1178]&m[1179]&~m[1180]&~m[1181]&m[1245])|(m[1178]&~m[1179]&m[1180]&~m[1181]&m[1245])|(~m[1178]&m[1179]&m[1180]&~m[1181]&m[1245])|(m[1178]&m[1179]&m[1180]&~m[1181]&m[1245])|(m[1178]&m[1179]&m[1180]&m[1181]&m[1245]))):InitCond[1505];
    m[1187] = run?((((m[1183]&~m[1184]&~m[1185]&~m[1186]&~m[1248])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1248])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1248])|(m[1183]&m[1184]&~m[1185]&m[1186]&~m[1248])|(m[1183]&~m[1184]&m[1185]&m[1186]&~m[1248])|(~m[1183]&m[1184]&m[1185]&m[1186]&~m[1248]))&BiasedRNG[790])|(((m[1183]&~m[1184]&~m[1185]&~m[1186]&m[1248])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&m[1248])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&m[1248])|(m[1183]&m[1184]&~m[1185]&m[1186]&m[1248])|(m[1183]&~m[1184]&m[1185]&m[1186]&m[1248])|(~m[1183]&m[1184]&m[1185]&m[1186]&m[1248]))&~BiasedRNG[790])|((m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1248])|(m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1248])|(~m[1183]&m[1184]&m[1185]&~m[1186]&~m[1248])|(m[1183]&m[1184]&m[1185]&~m[1186]&~m[1248])|(m[1183]&m[1184]&m[1185]&m[1186]&~m[1248])|(m[1183]&m[1184]&~m[1185]&~m[1186]&m[1248])|(m[1183]&~m[1184]&m[1185]&~m[1186]&m[1248])|(~m[1183]&m[1184]&m[1185]&~m[1186]&m[1248])|(m[1183]&m[1184]&m[1185]&~m[1186]&m[1248])|(m[1183]&m[1184]&m[1185]&m[1186]&m[1248]))):InitCond[1506];
    m[1192] = run?((((m[1188]&~m[1189]&~m[1190]&~m[1191]&~m[1250])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1250])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1250])|(m[1188]&m[1189]&~m[1190]&m[1191]&~m[1250])|(m[1188]&~m[1189]&m[1190]&m[1191]&~m[1250])|(~m[1188]&m[1189]&m[1190]&m[1191]&~m[1250]))&BiasedRNG[791])|(((m[1188]&~m[1189]&~m[1190]&~m[1191]&m[1250])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&m[1250])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&m[1250])|(m[1188]&m[1189]&~m[1190]&m[1191]&m[1250])|(m[1188]&~m[1189]&m[1190]&m[1191]&m[1250])|(~m[1188]&m[1189]&m[1190]&m[1191]&m[1250]))&~BiasedRNG[791])|((m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1250])|(m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1250])|(~m[1188]&m[1189]&m[1190]&~m[1191]&~m[1250])|(m[1188]&m[1189]&m[1190]&~m[1191]&~m[1250])|(m[1188]&m[1189]&m[1190]&m[1191]&~m[1250])|(m[1188]&m[1189]&~m[1190]&~m[1191]&m[1250])|(m[1188]&~m[1189]&m[1190]&~m[1191]&m[1250])|(~m[1188]&m[1189]&m[1190]&~m[1191]&m[1250])|(m[1188]&m[1189]&m[1190]&~m[1191]&m[1250])|(m[1188]&m[1189]&m[1190]&m[1191]&m[1250]))):InitCond[1507];
    m[1197] = run?((((m[1193]&~m[1194]&~m[1195]&~m[1196]&~m[1255])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1255])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1255])|(m[1193]&m[1194]&~m[1195]&m[1196]&~m[1255])|(m[1193]&~m[1194]&m[1195]&m[1196]&~m[1255])|(~m[1193]&m[1194]&m[1195]&m[1196]&~m[1255]))&BiasedRNG[792])|(((m[1193]&~m[1194]&~m[1195]&~m[1196]&m[1255])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&m[1255])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&m[1255])|(m[1193]&m[1194]&~m[1195]&m[1196]&m[1255])|(m[1193]&~m[1194]&m[1195]&m[1196]&m[1255])|(~m[1193]&m[1194]&m[1195]&m[1196]&m[1255]))&~BiasedRNG[792])|((m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1255])|(m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1255])|(~m[1193]&m[1194]&m[1195]&~m[1196]&~m[1255])|(m[1193]&m[1194]&m[1195]&~m[1196]&~m[1255])|(m[1193]&m[1194]&m[1195]&m[1196]&~m[1255])|(m[1193]&m[1194]&~m[1195]&~m[1196]&m[1255])|(m[1193]&~m[1194]&m[1195]&~m[1196]&m[1255])|(~m[1193]&m[1194]&m[1195]&~m[1196]&m[1255])|(m[1193]&m[1194]&m[1195]&~m[1196]&m[1255])|(m[1193]&m[1194]&m[1195]&m[1196]&m[1255]))):InitCond[1508];
    m[1202] = run?((((m[1198]&~m[1199]&~m[1200]&~m[1201]&~m[1260])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1260])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1260])|(m[1198]&m[1199]&~m[1200]&m[1201]&~m[1260])|(m[1198]&~m[1199]&m[1200]&m[1201]&~m[1260])|(~m[1198]&m[1199]&m[1200]&m[1201]&~m[1260]))&BiasedRNG[793])|(((m[1198]&~m[1199]&~m[1200]&~m[1201]&m[1260])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&m[1260])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&m[1260])|(m[1198]&m[1199]&~m[1200]&m[1201]&m[1260])|(m[1198]&~m[1199]&m[1200]&m[1201]&m[1260])|(~m[1198]&m[1199]&m[1200]&m[1201]&m[1260]))&~BiasedRNG[793])|((m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1260])|(m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1260])|(~m[1198]&m[1199]&m[1200]&~m[1201]&~m[1260])|(m[1198]&m[1199]&m[1200]&~m[1201]&~m[1260])|(m[1198]&m[1199]&m[1200]&m[1201]&~m[1260])|(m[1198]&m[1199]&~m[1200]&~m[1201]&m[1260])|(m[1198]&~m[1199]&m[1200]&~m[1201]&m[1260])|(~m[1198]&m[1199]&m[1200]&~m[1201]&m[1260])|(m[1198]&m[1199]&m[1200]&~m[1201]&m[1260])|(m[1198]&m[1199]&m[1200]&m[1201]&m[1260]))):InitCond[1509];
    m[1207] = run?((((m[1203]&~m[1204]&~m[1205]&~m[1206]&~m[1265])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1265])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1265])|(m[1203]&m[1204]&~m[1205]&m[1206]&~m[1265])|(m[1203]&~m[1204]&m[1205]&m[1206]&~m[1265])|(~m[1203]&m[1204]&m[1205]&m[1206]&~m[1265]))&BiasedRNG[794])|(((m[1203]&~m[1204]&~m[1205]&~m[1206]&m[1265])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&m[1265])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&m[1265])|(m[1203]&m[1204]&~m[1205]&m[1206]&m[1265])|(m[1203]&~m[1204]&m[1205]&m[1206]&m[1265])|(~m[1203]&m[1204]&m[1205]&m[1206]&m[1265]))&~BiasedRNG[794])|((m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1265])|(m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1265])|(~m[1203]&m[1204]&m[1205]&~m[1206]&~m[1265])|(m[1203]&m[1204]&m[1205]&~m[1206]&~m[1265])|(m[1203]&m[1204]&m[1205]&m[1206]&~m[1265])|(m[1203]&m[1204]&~m[1205]&~m[1206]&m[1265])|(m[1203]&~m[1204]&m[1205]&~m[1206]&m[1265])|(~m[1203]&m[1204]&m[1205]&~m[1206]&m[1265])|(m[1203]&m[1204]&m[1205]&~m[1206]&m[1265])|(m[1203]&m[1204]&m[1205]&m[1206]&m[1265]))):InitCond[1510];
    m[1212] = run?((((m[1208]&~m[1209]&~m[1210]&~m[1211]&~m[1270])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1270])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1270])|(m[1208]&m[1209]&~m[1210]&m[1211]&~m[1270])|(m[1208]&~m[1209]&m[1210]&m[1211]&~m[1270])|(~m[1208]&m[1209]&m[1210]&m[1211]&~m[1270]))&BiasedRNG[795])|(((m[1208]&~m[1209]&~m[1210]&~m[1211]&m[1270])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&m[1270])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&m[1270])|(m[1208]&m[1209]&~m[1210]&m[1211]&m[1270])|(m[1208]&~m[1209]&m[1210]&m[1211]&m[1270])|(~m[1208]&m[1209]&m[1210]&m[1211]&m[1270]))&~BiasedRNG[795])|((m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1270])|(m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1270])|(~m[1208]&m[1209]&m[1210]&~m[1211]&~m[1270])|(m[1208]&m[1209]&m[1210]&~m[1211]&~m[1270])|(m[1208]&m[1209]&m[1210]&m[1211]&~m[1270])|(m[1208]&m[1209]&~m[1210]&~m[1211]&m[1270])|(m[1208]&~m[1209]&m[1210]&~m[1211]&m[1270])|(~m[1208]&m[1209]&m[1210]&~m[1211]&m[1270])|(m[1208]&m[1209]&m[1210]&~m[1211]&m[1270])|(m[1208]&m[1209]&m[1210]&m[1211]&m[1270]))):InitCond[1511];
    m[1217] = run?((((m[1213]&~m[1214]&~m[1215]&~m[1216]&~m[1275])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1275])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1275])|(m[1213]&m[1214]&~m[1215]&m[1216]&~m[1275])|(m[1213]&~m[1214]&m[1215]&m[1216]&~m[1275])|(~m[1213]&m[1214]&m[1215]&m[1216]&~m[1275]))&BiasedRNG[796])|(((m[1213]&~m[1214]&~m[1215]&~m[1216]&m[1275])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&m[1275])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&m[1275])|(m[1213]&m[1214]&~m[1215]&m[1216]&m[1275])|(m[1213]&~m[1214]&m[1215]&m[1216]&m[1275])|(~m[1213]&m[1214]&m[1215]&m[1216]&m[1275]))&~BiasedRNG[796])|((m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1275])|(m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1275])|(~m[1213]&m[1214]&m[1215]&~m[1216]&~m[1275])|(m[1213]&m[1214]&m[1215]&~m[1216]&~m[1275])|(m[1213]&m[1214]&m[1215]&m[1216]&~m[1275])|(m[1213]&m[1214]&~m[1215]&~m[1216]&m[1275])|(m[1213]&~m[1214]&m[1215]&~m[1216]&m[1275])|(~m[1213]&m[1214]&m[1215]&~m[1216]&m[1275])|(m[1213]&m[1214]&m[1215]&~m[1216]&m[1275])|(m[1213]&m[1214]&m[1215]&m[1216]&m[1275]))):InitCond[1512];
    m[1222] = run?((((m[1218]&~m[1219]&~m[1220]&~m[1221]&~m[1280])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1280])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1280])|(m[1218]&m[1219]&~m[1220]&m[1221]&~m[1280])|(m[1218]&~m[1219]&m[1220]&m[1221]&~m[1280])|(~m[1218]&m[1219]&m[1220]&m[1221]&~m[1280]))&BiasedRNG[797])|(((m[1218]&~m[1219]&~m[1220]&~m[1221]&m[1280])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&m[1280])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&m[1280])|(m[1218]&m[1219]&~m[1220]&m[1221]&m[1280])|(m[1218]&~m[1219]&m[1220]&m[1221]&m[1280])|(~m[1218]&m[1219]&m[1220]&m[1221]&m[1280]))&~BiasedRNG[797])|((m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1280])|(m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1280])|(~m[1218]&m[1219]&m[1220]&~m[1221]&~m[1280])|(m[1218]&m[1219]&m[1220]&~m[1221]&~m[1280])|(m[1218]&m[1219]&m[1220]&m[1221]&~m[1280])|(m[1218]&m[1219]&~m[1220]&~m[1221]&m[1280])|(m[1218]&~m[1219]&m[1220]&~m[1221]&m[1280])|(~m[1218]&m[1219]&m[1220]&~m[1221]&m[1280])|(m[1218]&m[1219]&m[1220]&~m[1221]&m[1280])|(m[1218]&m[1219]&m[1220]&m[1221]&m[1280]))):InitCond[1513];
    m[1227] = run?((((m[1223]&~m[1224]&~m[1225]&~m[1226]&~m[1285])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1285])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1285])|(m[1223]&m[1224]&~m[1225]&m[1226]&~m[1285])|(m[1223]&~m[1224]&m[1225]&m[1226]&~m[1285])|(~m[1223]&m[1224]&m[1225]&m[1226]&~m[1285]))&BiasedRNG[798])|(((m[1223]&~m[1224]&~m[1225]&~m[1226]&m[1285])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&m[1285])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&m[1285])|(m[1223]&m[1224]&~m[1225]&m[1226]&m[1285])|(m[1223]&~m[1224]&m[1225]&m[1226]&m[1285])|(~m[1223]&m[1224]&m[1225]&m[1226]&m[1285]))&~BiasedRNG[798])|((m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1285])|(m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1285])|(~m[1223]&m[1224]&m[1225]&~m[1226]&~m[1285])|(m[1223]&m[1224]&m[1225]&~m[1226]&~m[1285])|(m[1223]&m[1224]&m[1225]&m[1226]&~m[1285])|(m[1223]&m[1224]&~m[1225]&~m[1226]&m[1285])|(m[1223]&~m[1224]&m[1225]&~m[1226]&m[1285])|(~m[1223]&m[1224]&m[1225]&~m[1226]&m[1285])|(m[1223]&m[1224]&m[1225]&~m[1226]&m[1285])|(m[1223]&m[1224]&m[1225]&m[1226]&m[1285]))):InitCond[1514];
    m[1232] = run?((((m[1228]&~m[1229]&~m[1230]&~m[1231]&~m[1290])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1290])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1290])|(m[1228]&m[1229]&~m[1230]&m[1231]&~m[1290])|(m[1228]&~m[1229]&m[1230]&m[1231]&~m[1290])|(~m[1228]&m[1229]&m[1230]&m[1231]&~m[1290]))&BiasedRNG[799])|(((m[1228]&~m[1229]&~m[1230]&~m[1231]&m[1290])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&m[1290])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&m[1290])|(m[1228]&m[1229]&~m[1230]&m[1231]&m[1290])|(m[1228]&~m[1229]&m[1230]&m[1231]&m[1290])|(~m[1228]&m[1229]&m[1230]&m[1231]&m[1290]))&~BiasedRNG[799])|((m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1290])|(m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1290])|(~m[1228]&m[1229]&m[1230]&~m[1231]&~m[1290])|(m[1228]&m[1229]&m[1230]&~m[1231]&~m[1290])|(m[1228]&m[1229]&m[1230]&m[1231]&~m[1290])|(m[1228]&m[1229]&~m[1230]&~m[1231]&m[1290])|(m[1228]&~m[1229]&m[1230]&~m[1231]&m[1290])|(~m[1228]&m[1229]&m[1230]&~m[1231]&m[1290])|(m[1228]&m[1229]&m[1230]&~m[1231]&m[1290])|(m[1228]&m[1229]&m[1230]&m[1231]&m[1290]))):InitCond[1515];
    m[1237] = run?((((m[1233]&~m[1234]&~m[1235]&~m[1236]&~m[1295])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1295])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1295])|(m[1233]&m[1234]&~m[1235]&m[1236]&~m[1295])|(m[1233]&~m[1234]&m[1235]&m[1236]&~m[1295])|(~m[1233]&m[1234]&m[1235]&m[1236]&~m[1295]))&BiasedRNG[800])|(((m[1233]&~m[1234]&~m[1235]&~m[1236]&m[1295])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&m[1295])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&m[1295])|(m[1233]&m[1234]&~m[1235]&m[1236]&m[1295])|(m[1233]&~m[1234]&m[1235]&m[1236]&m[1295])|(~m[1233]&m[1234]&m[1235]&m[1236]&m[1295]))&~BiasedRNG[800])|((m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1295])|(m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1295])|(~m[1233]&m[1234]&m[1235]&~m[1236]&~m[1295])|(m[1233]&m[1234]&m[1235]&~m[1236]&~m[1295])|(m[1233]&m[1234]&m[1235]&m[1236]&~m[1295])|(m[1233]&m[1234]&~m[1235]&~m[1236]&m[1295])|(m[1233]&~m[1234]&m[1235]&~m[1236]&m[1295])|(~m[1233]&m[1234]&m[1235]&~m[1236]&m[1295])|(m[1233]&m[1234]&m[1235]&~m[1236]&m[1295])|(m[1233]&m[1234]&m[1235]&m[1236]&m[1295]))):InitCond[1516];
    m[1242] = run?((((m[1238]&~m[1239]&~m[1240]&~m[1241]&~m[1300])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1300])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1300])|(m[1238]&m[1239]&~m[1240]&m[1241]&~m[1300])|(m[1238]&~m[1239]&m[1240]&m[1241]&~m[1300])|(~m[1238]&m[1239]&m[1240]&m[1241]&~m[1300]))&BiasedRNG[801])|(((m[1238]&~m[1239]&~m[1240]&~m[1241]&m[1300])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&m[1300])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&m[1300])|(m[1238]&m[1239]&~m[1240]&m[1241]&m[1300])|(m[1238]&~m[1239]&m[1240]&m[1241]&m[1300])|(~m[1238]&m[1239]&m[1240]&m[1241]&m[1300]))&~BiasedRNG[801])|((m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1300])|(m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1300])|(~m[1238]&m[1239]&m[1240]&~m[1241]&~m[1300])|(m[1238]&m[1239]&m[1240]&~m[1241]&~m[1300])|(m[1238]&m[1239]&m[1240]&m[1241]&~m[1300])|(m[1238]&m[1239]&~m[1240]&~m[1241]&m[1300])|(m[1238]&~m[1239]&m[1240]&~m[1241]&m[1300])|(~m[1238]&m[1239]&m[1240]&~m[1241]&m[1300])|(m[1238]&m[1239]&m[1240]&~m[1241]&m[1300])|(m[1238]&m[1239]&m[1240]&m[1241]&m[1300]))):InitCond[1517];
    m[1247] = run?((((m[1243]&~m[1244]&~m[1245]&~m[1246]&~m[1305])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1305])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1305])|(m[1243]&m[1244]&~m[1245]&m[1246]&~m[1305])|(m[1243]&~m[1244]&m[1245]&m[1246]&~m[1305])|(~m[1243]&m[1244]&m[1245]&m[1246]&~m[1305]))&BiasedRNG[802])|(((m[1243]&~m[1244]&~m[1245]&~m[1246]&m[1305])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&m[1305])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&m[1305])|(m[1243]&m[1244]&~m[1245]&m[1246]&m[1305])|(m[1243]&~m[1244]&m[1245]&m[1246]&m[1305])|(~m[1243]&m[1244]&m[1245]&m[1246]&m[1305]))&~BiasedRNG[802])|((m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1305])|(m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1305])|(~m[1243]&m[1244]&m[1245]&~m[1246]&~m[1305])|(m[1243]&m[1244]&m[1245]&~m[1246]&~m[1305])|(m[1243]&m[1244]&m[1245]&m[1246]&~m[1305])|(m[1243]&m[1244]&~m[1245]&~m[1246]&m[1305])|(m[1243]&~m[1244]&m[1245]&~m[1246]&m[1305])|(~m[1243]&m[1244]&m[1245]&~m[1246]&m[1305])|(m[1243]&m[1244]&m[1245]&~m[1246]&m[1305])|(m[1243]&m[1244]&m[1245]&m[1246]&m[1305]))):InitCond[1518];
    m[1252] = run?((((m[1248]&~m[1249]&~m[1250]&~m[1251]&~m[1308])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1308])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1308])|(m[1248]&m[1249]&~m[1250]&m[1251]&~m[1308])|(m[1248]&~m[1249]&m[1250]&m[1251]&~m[1308])|(~m[1248]&m[1249]&m[1250]&m[1251]&~m[1308]))&BiasedRNG[803])|(((m[1248]&~m[1249]&~m[1250]&~m[1251]&m[1308])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&m[1308])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&m[1308])|(m[1248]&m[1249]&~m[1250]&m[1251]&m[1308])|(m[1248]&~m[1249]&m[1250]&m[1251]&m[1308])|(~m[1248]&m[1249]&m[1250]&m[1251]&m[1308]))&~BiasedRNG[803])|((m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1308])|(m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1308])|(~m[1248]&m[1249]&m[1250]&~m[1251]&~m[1308])|(m[1248]&m[1249]&m[1250]&~m[1251]&~m[1308])|(m[1248]&m[1249]&m[1250]&m[1251]&~m[1308])|(m[1248]&m[1249]&~m[1250]&~m[1251]&m[1308])|(m[1248]&~m[1249]&m[1250]&~m[1251]&m[1308])|(~m[1248]&m[1249]&m[1250]&~m[1251]&m[1308])|(m[1248]&m[1249]&m[1250]&~m[1251]&m[1308])|(m[1248]&m[1249]&m[1250]&m[1251]&m[1308]))):InitCond[1519];
    m[1257] = run?((((m[1253]&~m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&~m[1310]))&BiasedRNG[804])|(((m[1253]&~m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&m[1310]))&~BiasedRNG[804])|((m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&m[1310]))):InitCond[1520];
    m[1262] = run?((((m[1258]&~m[1259]&~m[1260]&~m[1261]&~m[1315])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1315])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1315])|(m[1258]&m[1259]&~m[1260]&m[1261]&~m[1315])|(m[1258]&~m[1259]&m[1260]&m[1261]&~m[1315])|(~m[1258]&m[1259]&m[1260]&m[1261]&~m[1315]))&BiasedRNG[805])|(((m[1258]&~m[1259]&~m[1260]&~m[1261]&m[1315])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&m[1315])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&m[1315])|(m[1258]&m[1259]&~m[1260]&m[1261]&m[1315])|(m[1258]&~m[1259]&m[1260]&m[1261]&m[1315])|(~m[1258]&m[1259]&m[1260]&m[1261]&m[1315]))&~BiasedRNG[805])|((m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1315])|(m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1315])|(~m[1258]&m[1259]&m[1260]&~m[1261]&~m[1315])|(m[1258]&m[1259]&m[1260]&~m[1261]&~m[1315])|(m[1258]&m[1259]&m[1260]&m[1261]&~m[1315])|(m[1258]&m[1259]&~m[1260]&~m[1261]&m[1315])|(m[1258]&~m[1259]&m[1260]&~m[1261]&m[1315])|(~m[1258]&m[1259]&m[1260]&~m[1261]&m[1315])|(m[1258]&m[1259]&m[1260]&~m[1261]&m[1315])|(m[1258]&m[1259]&m[1260]&m[1261]&m[1315]))):InitCond[1521];
    m[1267] = run?((((m[1263]&~m[1264]&~m[1265]&~m[1266]&~m[1320])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1320])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1320])|(m[1263]&m[1264]&~m[1265]&m[1266]&~m[1320])|(m[1263]&~m[1264]&m[1265]&m[1266]&~m[1320])|(~m[1263]&m[1264]&m[1265]&m[1266]&~m[1320]))&BiasedRNG[806])|(((m[1263]&~m[1264]&~m[1265]&~m[1266]&m[1320])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&m[1320])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&m[1320])|(m[1263]&m[1264]&~m[1265]&m[1266]&m[1320])|(m[1263]&~m[1264]&m[1265]&m[1266]&m[1320])|(~m[1263]&m[1264]&m[1265]&m[1266]&m[1320]))&~BiasedRNG[806])|((m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1320])|(m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1320])|(~m[1263]&m[1264]&m[1265]&~m[1266]&~m[1320])|(m[1263]&m[1264]&m[1265]&~m[1266]&~m[1320])|(m[1263]&m[1264]&m[1265]&m[1266]&~m[1320])|(m[1263]&m[1264]&~m[1265]&~m[1266]&m[1320])|(m[1263]&~m[1264]&m[1265]&~m[1266]&m[1320])|(~m[1263]&m[1264]&m[1265]&~m[1266]&m[1320])|(m[1263]&m[1264]&m[1265]&~m[1266]&m[1320])|(m[1263]&m[1264]&m[1265]&m[1266]&m[1320]))):InitCond[1522];
    m[1272] = run?((((m[1268]&~m[1269]&~m[1270]&~m[1271]&~m[1325])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1325])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1325])|(m[1268]&m[1269]&~m[1270]&m[1271]&~m[1325])|(m[1268]&~m[1269]&m[1270]&m[1271]&~m[1325])|(~m[1268]&m[1269]&m[1270]&m[1271]&~m[1325]))&BiasedRNG[807])|(((m[1268]&~m[1269]&~m[1270]&~m[1271]&m[1325])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&m[1325])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&m[1325])|(m[1268]&m[1269]&~m[1270]&m[1271]&m[1325])|(m[1268]&~m[1269]&m[1270]&m[1271]&m[1325])|(~m[1268]&m[1269]&m[1270]&m[1271]&m[1325]))&~BiasedRNG[807])|((m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1325])|(m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1325])|(~m[1268]&m[1269]&m[1270]&~m[1271]&~m[1325])|(m[1268]&m[1269]&m[1270]&~m[1271]&~m[1325])|(m[1268]&m[1269]&m[1270]&m[1271]&~m[1325])|(m[1268]&m[1269]&~m[1270]&~m[1271]&m[1325])|(m[1268]&~m[1269]&m[1270]&~m[1271]&m[1325])|(~m[1268]&m[1269]&m[1270]&~m[1271]&m[1325])|(m[1268]&m[1269]&m[1270]&~m[1271]&m[1325])|(m[1268]&m[1269]&m[1270]&m[1271]&m[1325]))):InitCond[1523];
    m[1277] = run?((((m[1273]&~m[1274]&~m[1275]&~m[1276]&~m[1330])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1330])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1330])|(m[1273]&m[1274]&~m[1275]&m[1276]&~m[1330])|(m[1273]&~m[1274]&m[1275]&m[1276]&~m[1330])|(~m[1273]&m[1274]&m[1275]&m[1276]&~m[1330]))&BiasedRNG[808])|(((m[1273]&~m[1274]&~m[1275]&~m[1276]&m[1330])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&m[1330])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&m[1330])|(m[1273]&m[1274]&~m[1275]&m[1276]&m[1330])|(m[1273]&~m[1274]&m[1275]&m[1276]&m[1330])|(~m[1273]&m[1274]&m[1275]&m[1276]&m[1330]))&~BiasedRNG[808])|((m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1330])|(m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1330])|(~m[1273]&m[1274]&m[1275]&~m[1276]&~m[1330])|(m[1273]&m[1274]&m[1275]&~m[1276]&~m[1330])|(m[1273]&m[1274]&m[1275]&m[1276]&~m[1330])|(m[1273]&m[1274]&~m[1275]&~m[1276]&m[1330])|(m[1273]&~m[1274]&m[1275]&~m[1276]&m[1330])|(~m[1273]&m[1274]&m[1275]&~m[1276]&m[1330])|(m[1273]&m[1274]&m[1275]&~m[1276]&m[1330])|(m[1273]&m[1274]&m[1275]&m[1276]&m[1330]))):InitCond[1524];
    m[1282] = run?((((m[1278]&~m[1279]&~m[1280]&~m[1281]&~m[1335])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1335])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1335])|(m[1278]&m[1279]&~m[1280]&m[1281]&~m[1335])|(m[1278]&~m[1279]&m[1280]&m[1281]&~m[1335])|(~m[1278]&m[1279]&m[1280]&m[1281]&~m[1335]))&BiasedRNG[809])|(((m[1278]&~m[1279]&~m[1280]&~m[1281]&m[1335])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&m[1335])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&m[1335])|(m[1278]&m[1279]&~m[1280]&m[1281]&m[1335])|(m[1278]&~m[1279]&m[1280]&m[1281]&m[1335])|(~m[1278]&m[1279]&m[1280]&m[1281]&m[1335]))&~BiasedRNG[809])|((m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1335])|(m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1335])|(~m[1278]&m[1279]&m[1280]&~m[1281]&~m[1335])|(m[1278]&m[1279]&m[1280]&~m[1281]&~m[1335])|(m[1278]&m[1279]&m[1280]&m[1281]&~m[1335])|(m[1278]&m[1279]&~m[1280]&~m[1281]&m[1335])|(m[1278]&~m[1279]&m[1280]&~m[1281]&m[1335])|(~m[1278]&m[1279]&m[1280]&~m[1281]&m[1335])|(m[1278]&m[1279]&m[1280]&~m[1281]&m[1335])|(m[1278]&m[1279]&m[1280]&m[1281]&m[1335]))):InitCond[1525];
    m[1287] = run?((((m[1283]&~m[1284]&~m[1285]&~m[1286]&~m[1340])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1340])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1340])|(m[1283]&m[1284]&~m[1285]&m[1286]&~m[1340])|(m[1283]&~m[1284]&m[1285]&m[1286]&~m[1340])|(~m[1283]&m[1284]&m[1285]&m[1286]&~m[1340]))&BiasedRNG[810])|(((m[1283]&~m[1284]&~m[1285]&~m[1286]&m[1340])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&m[1340])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&m[1340])|(m[1283]&m[1284]&~m[1285]&m[1286]&m[1340])|(m[1283]&~m[1284]&m[1285]&m[1286]&m[1340])|(~m[1283]&m[1284]&m[1285]&m[1286]&m[1340]))&~BiasedRNG[810])|((m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1340])|(m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1340])|(~m[1283]&m[1284]&m[1285]&~m[1286]&~m[1340])|(m[1283]&m[1284]&m[1285]&~m[1286]&~m[1340])|(m[1283]&m[1284]&m[1285]&m[1286]&~m[1340])|(m[1283]&m[1284]&~m[1285]&~m[1286]&m[1340])|(m[1283]&~m[1284]&m[1285]&~m[1286]&m[1340])|(~m[1283]&m[1284]&m[1285]&~m[1286]&m[1340])|(m[1283]&m[1284]&m[1285]&~m[1286]&m[1340])|(m[1283]&m[1284]&m[1285]&m[1286]&m[1340]))):InitCond[1526];
    m[1292] = run?((((m[1288]&~m[1289]&~m[1290]&~m[1291]&~m[1345])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1345])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1345])|(m[1288]&m[1289]&~m[1290]&m[1291]&~m[1345])|(m[1288]&~m[1289]&m[1290]&m[1291]&~m[1345])|(~m[1288]&m[1289]&m[1290]&m[1291]&~m[1345]))&BiasedRNG[811])|(((m[1288]&~m[1289]&~m[1290]&~m[1291]&m[1345])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&m[1345])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&m[1345])|(m[1288]&m[1289]&~m[1290]&m[1291]&m[1345])|(m[1288]&~m[1289]&m[1290]&m[1291]&m[1345])|(~m[1288]&m[1289]&m[1290]&m[1291]&m[1345]))&~BiasedRNG[811])|((m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1345])|(m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1345])|(~m[1288]&m[1289]&m[1290]&~m[1291]&~m[1345])|(m[1288]&m[1289]&m[1290]&~m[1291]&~m[1345])|(m[1288]&m[1289]&m[1290]&m[1291]&~m[1345])|(m[1288]&m[1289]&~m[1290]&~m[1291]&m[1345])|(m[1288]&~m[1289]&m[1290]&~m[1291]&m[1345])|(~m[1288]&m[1289]&m[1290]&~m[1291]&m[1345])|(m[1288]&m[1289]&m[1290]&~m[1291]&m[1345])|(m[1288]&m[1289]&m[1290]&m[1291]&m[1345]))):InitCond[1527];
    m[1297] = run?((((m[1293]&~m[1294]&~m[1295]&~m[1296]&~m[1350])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1350])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1350])|(m[1293]&m[1294]&~m[1295]&m[1296]&~m[1350])|(m[1293]&~m[1294]&m[1295]&m[1296]&~m[1350])|(~m[1293]&m[1294]&m[1295]&m[1296]&~m[1350]))&BiasedRNG[812])|(((m[1293]&~m[1294]&~m[1295]&~m[1296]&m[1350])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&m[1350])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&m[1350])|(m[1293]&m[1294]&~m[1295]&m[1296]&m[1350])|(m[1293]&~m[1294]&m[1295]&m[1296]&m[1350])|(~m[1293]&m[1294]&m[1295]&m[1296]&m[1350]))&~BiasedRNG[812])|((m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1350])|(m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1350])|(~m[1293]&m[1294]&m[1295]&~m[1296]&~m[1350])|(m[1293]&m[1294]&m[1295]&~m[1296]&~m[1350])|(m[1293]&m[1294]&m[1295]&m[1296]&~m[1350])|(m[1293]&m[1294]&~m[1295]&~m[1296]&m[1350])|(m[1293]&~m[1294]&m[1295]&~m[1296]&m[1350])|(~m[1293]&m[1294]&m[1295]&~m[1296]&m[1350])|(m[1293]&m[1294]&m[1295]&~m[1296]&m[1350])|(m[1293]&m[1294]&m[1295]&m[1296]&m[1350]))):InitCond[1528];
    m[1302] = run?((((m[1298]&~m[1299]&~m[1300]&~m[1301]&~m[1355])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1355])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1355])|(m[1298]&m[1299]&~m[1300]&m[1301]&~m[1355])|(m[1298]&~m[1299]&m[1300]&m[1301]&~m[1355])|(~m[1298]&m[1299]&m[1300]&m[1301]&~m[1355]))&BiasedRNG[813])|(((m[1298]&~m[1299]&~m[1300]&~m[1301]&m[1355])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&m[1355])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&m[1355])|(m[1298]&m[1299]&~m[1300]&m[1301]&m[1355])|(m[1298]&~m[1299]&m[1300]&m[1301]&m[1355])|(~m[1298]&m[1299]&m[1300]&m[1301]&m[1355]))&~BiasedRNG[813])|((m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1355])|(m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1355])|(~m[1298]&m[1299]&m[1300]&~m[1301]&~m[1355])|(m[1298]&m[1299]&m[1300]&~m[1301]&~m[1355])|(m[1298]&m[1299]&m[1300]&m[1301]&~m[1355])|(m[1298]&m[1299]&~m[1300]&~m[1301]&m[1355])|(m[1298]&~m[1299]&m[1300]&~m[1301]&m[1355])|(~m[1298]&m[1299]&m[1300]&~m[1301]&m[1355])|(m[1298]&m[1299]&m[1300]&~m[1301]&m[1355])|(m[1298]&m[1299]&m[1300]&m[1301]&m[1355]))):InitCond[1529];
    m[1307] = run?((((m[1303]&~m[1304]&~m[1305]&~m[1306]&~m[1360])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1360])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1360])|(m[1303]&m[1304]&~m[1305]&m[1306]&~m[1360])|(m[1303]&~m[1304]&m[1305]&m[1306]&~m[1360])|(~m[1303]&m[1304]&m[1305]&m[1306]&~m[1360]))&BiasedRNG[814])|(((m[1303]&~m[1304]&~m[1305]&~m[1306]&m[1360])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&m[1360])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&m[1360])|(m[1303]&m[1304]&~m[1305]&m[1306]&m[1360])|(m[1303]&~m[1304]&m[1305]&m[1306]&m[1360])|(~m[1303]&m[1304]&m[1305]&m[1306]&m[1360]))&~BiasedRNG[814])|((m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1360])|(m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1360])|(~m[1303]&m[1304]&m[1305]&~m[1306]&~m[1360])|(m[1303]&m[1304]&m[1305]&~m[1306]&~m[1360])|(m[1303]&m[1304]&m[1305]&m[1306]&~m[1360])|(m[1303]&m[1304]&~m[1305]&~m[1306]&m[1360])|(m[1303]&~m[1304]&m[1305]&~m[1306]&m[1360])|(~m[1303]&m[1304]&m[1305]&~m[1306]&m[1360])|(m[1303]&m[1304]&m[1305]&~m[1306]&m[1360])|(m[1303]&m[1304]&m[1305]&m[1306]&m[1360]))):InitCond[1530];
    m[1312] = run?((((m[1308]&~m[1309]&~m[1310]&~m[1311]&~m[1363])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1363])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1363])|(m[1308]&m[1309]&~m[1310]&m[1311]&~m[1363])|(m[1308]&~m[1309]&m[1310]&m[1311]&~m[1363])|(~m[1308]&m[1309]&m[1310]&m[1311]&~m[1363]))&BiasedRNG[815])|(((m[1308]&~m[1309]&~m[1310]&~m[1311]&m[1363])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&m[1363])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&m[1363])|(m[1308]&m[1309]&~m[1310]&m[1311]&m[1363])|(m[1308]&~m[1309]&m[1310]&m[1311]&m[1363])|(~m[1308]&m[1309]&m[1310]&m[1311]&m[1363]))&~BiasedRNG[815])|((m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1363])|(m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1363])|(~m[1308]&m[1309]&m[1310]&~m[1311]&~m[1363])|(m[1308]&m[1309]&m[1310]&~m[1311]&~m[1363])|(m[1308]&m[1309]&m[1310]&m[1311]&~m[1363])|(m[1308]&m[1309]&~m[1310]&~m[1311]&m[1363])|(m[1308]&~m[1309]&m[1310]&~m[1311]&m[1363])|(~m[1308]&m[1309]&m[1310]&~m[1311]&m[1363])|(m[1308]&m[1309]&m[1310]&~m[1311]&m[1363])|(m[1308]&m[1309]&m[1310]&m[1311]&m[1363]))):InitCond[1531];
    m[1317] = run?((((m[1313]&~m[1314]&~m[1315]&~m[1316]&~m[1365])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1365])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1365])|(m[1313]&m[1314]&~m[1315]&m[1316]&~m[1365])|(m[1313]&~m[1314]&m[1315]&m[1316]&~m[1365])|(~m[1313]&m[1314]&m[1315]&m[1316]&~m[1365]))&BiasedRNG[816])|(((m[1313]&~m[1314]&~m[1315]&~m[1316]&m[1365])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&m[1365])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&m[1365])|(m[1313]&m[1314]&~m[1315]&m[1316]&m[1365])|(m[1313]&~m[1314]&m[1315]&m[1316]&m[1365])|(~m[1313]&m[1314]&m[1315]&m[1316]&m[1365]))&~BiasedRNG[816])|((m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1365])|(m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1365])|(~m[1313]&m[1314]&m[1315]&~m[1316]&~m[1365])|(m[1313]&m[1314]&m[1315]&~m[1316]&~m[1365])|(m[1313]&m[1314]&m[1315]&m[1316]&~m[1365])|(m[1313]&m[1314]&~m[1315]&~m[1316]&m[1365])|(m[1313]&~m[1314]&m[1315]&~m[1316]&m[1365])|(~m[1313]&m[1314]&m[1315]&~m[1316]&m[1365])|(m[1313]&m[1314]&m[1315]&~m[1316]&m[1365])|(m[1313]&m[1314]&m[1315]&m[1316]&m[1365]))):InitCond[1532];
    m[1322] = run?((((m[1318]&~m[1319]&~m[1320]&~m[1321]&~m[1370])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1370])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1370])|(m[1318]&m[1319]&~m[1320]&m[1321]&~m[1370])|(m[1318]&~m[1319]&m[1320]&m[1321]&~m[1370])|(~m[1318]&m[1319]&m[1320]&m[1321]&~m[1370]))&BiasedRNG[817])|(((m[1318]&~m[1319]&~m[1320]&~m[1321]&m[1370])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&m[1370])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&m[1370])|(m[1318]&m[1319]&~m[1320]&m[1321]&m[1370])|(m[1318]&~m[1319]&m[1320]&m[1321]&m[1370])|(~m[1318]&m[1319]&m[1320]&m[1321]&m[1370]))&~BiasedRNG[817])|((m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1370])|(m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1370])|(~m[1318]&m[1319]&m[1320]&~m[1321]&~m[1370])|(m[1318]&m[1319]&m[1320]&~m[1321]&~m[1370])|(m[1318]&m[1319]&m[1320]&m[1321]&~m[1370])|(m[1318]&m[1319]&~m[1320]&~m[1321]&m[1370])|(m[1318]&~m[1319]&m[1320]&~m[1321]&m[1370])|(~m[1318]&m[1319]&m[1320]&~m[1321]&m[1370])|(m[1318]&m[1319]&m[1320]&~m[1321]&m[1370])|(m[1318]&m[1319]&m[1320]&m[1321]&m[1370]))):InitCond[1533];
    m[1327] = run?((((m[1323]&~m[1324]&~m[1325]&~m[1326]&~m[1375])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1375])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1375])|(m[1323]&m[1324]&~m[1325]&m[1326]&~m[1375])|(m[1323]&~m[1324]&m[1325]&m[1326]&~m[1375])|(~m[1323]&m[1324]&m[1325]&m[1326]&~m[1375]))&BiasedRNG[818])|(((m[1323]&~m[1324]&~m[1325]&~m[1326]&m[1375])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&m[1375])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&m[1375])|(m[1323]&m[1324]&~m[1325]&m[1326]&m[1375])|(m[1323]&~m[1324]&m[1325]&m[1326]&m[1375])|(~m[1323]&m[1324]&m[1325]&m[1326]&m[1375]))&~BiasedRNG[818])|((m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1375])|(m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1375])|(~m[1323]&m[1324]&m[1325]&~m[1326]&~m[1375])|(m[1323]&m[1324]&m[1325]&~m[1326]&~m[1375])|(m[1323]&m[1324]&m[1325]&m[1326]&~m[1375])|(m[1323]&m[1324]&~m[1325]&~m[1326]&m[1375])|(m[1323]&~m[1324]&m[1325]&~m[1326]&m[1375])|(~m[1323]&m[1324]&m[1325]&~m[1326]&m[1375])|(m[1323]&m[1324]&m[1325]&~m[1326]&m[1375])|(m[1323]&m[1324]&m[1325]&m[1326]&m[1375]))):InitCond[1534];
    m[1332] = run?((((m[1328]&~m[1329]&~m[1330]&~m[1331]&~m[1380])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1380])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1380])|(m[1328]&m[1329]&~m[1330]&m[1331]&~m[1380])|(m[1328]&~m[1329]&m[1330]&m[1331]&~m[1380])|(~m[1328]&m[1329]&m[1330]&m[1331]&~m[1380]))&BiasedRNG[819])|(((m[1328]&~m[1329]&~m[1330]&~m[1331]&m[1380])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&m[1380])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&m[1380])|(m[1328]&m[1329]&~m[1330]&m[1331]&m[1380])|(m[1328]&~m[1329]&m[1330]&m[1331]&m[1380])|(~m[1328]&m[1329]&m[1330]&m[1331]&m[1380]))&~BiasedRNG[819])|((m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1380])|(m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1380])|(~m[1328]&m[1329]&m[1330]&~m[1331]&~m[1380])|(m[1328]&m[1329]&m[1330]&~m[1331]&~m[1380])|(m[1328]&m[1329]&m[1330]&m[1331]&~m[1380])|(m[1328]&m[1329]&~m[1330]&~m[1331]&m[1380])|(m[1328]&~m[1329]&m[1330]&~m[1331]&m[1380])|(~m[1328]&m[1329]&m[1330]&~m[1331]&m[1380])|(m[1328]&m[1329]&m[1330]&~m[1331]&m[1380])|(m[1328]&m[1329]&m[1330]&m[1331]&m[1380]))):InitCond[1535];
    m[1337] = run?((((m[1333]&~m[1334]&~m[1335]&~m[1336]&~m[1385])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1385])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1385])|(m[1333]&m[1334]&~m[1335]&m[1336]&~m[1385])|(m[1333]&~m[1334]&m[1335]&m[1336]&~m[1385])|(~m[1333]&m[1334]&m[1335]&m[1336]&~m[1385]))&BiasedRNG[820])|(((m[1333]&~m[1334]&~m[1335]&~m[1336]&m[1385])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&m[1385])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&m[1385])|(m[1333]&m[1334]&~m[1335]&m[1336]&m[1385])|(m[1333]&~m[1334]&m[1335]&m[1336]&m[1385])|(~m[1333]&m[1334]&m[1335]&m[1336]&m[1385]))&~BiasedRNG[820])|((m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1385])|(m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1385])|(~m[1333]&m[1334]&m[1335]&~m[1336]&~m[1385])|(m[1333]&m[1334]&m[1335]&~m[1336]&~m[1385])|(m[1333]&m[1334]&m[1335]&m[1336]&~m[1385])|(m[1333]&m[1334]&~m[1335]&~m[1336]&m[1385])|(m[1333]&~m[1334]&m[1335]&~m[1336]&m[1385])|(~m[1333]&m[1334]&m[1335]&~m[1336]&m[1385])|(m[1333]&m[1334]&m[1335]&~m[1336]&m[1385])|(m[1333]&m[1334]&m[1335]&m[1336]&m[1385]))):InitCond[1536];
    m[1342] = run?((((m[1338]&~m[1339]&~m[1340]&~m[1341]&~m[1390])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1390])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1390])|(m[1338]&m[1339]&~m[1340]&m[1341]&~m[1390])|(m[1338]&~m[1339]&m[1340]&m[1341]&~m[1390])|(~m[1338]&m[1339]&m[1340]&m[1341]&~m[1390]))&BiasedRNG[821])|(((m[1338]&~m[1339]&~m[1340]&~m[1341]&m[1390])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&m[1390])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&m[1390])|(m[1338]&m[1339]&~m[1340]&m[1341]&m[1390])|(m[1338]&~m[1339]&m[1340]&m[1341]&m[1390])|(~m[1338]&m[1339]&m[1340]&m[1341]&m[1390]))&~BiasedRNG[821])|((m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1390])|(m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1390])|(~m[1338]&m[1339]&m[1340]&~m[1341]&~m[1390])|(m[1338]&m[1339]&m[1340]&~m[1341]&~m[1390])|(m[1338]&m[1339]&m[1340]&m[1341]&~m[1390])|(m[1338]&m[1339]&~m[1340]&~m[1341]&m[1390])|(m[1338]&~m[1339]&m[1340]&~m[1341]&m[1390])|(~m[1338]&m[1339]&m[1340]&~m[1341]&m[1390])|(m[1338]&m[1339]&m[1340]&~m[1341]&m[1390])|(m[1338]&m[1339]&m[1340]&m[1341]&m[1390]))):InitCond[1537];
    m[1347] = run?((((m[1343]&~m[1344]&~m[1345]&~m[1346]&~m[1395])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1395])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1395])|(m[1343]&m[1344]&~m[1345]&m[1346]&~m[1395])|(m[1343]&~m[1344]&m[1345]&m[1346]&~m[1395])|(~m[1343]&m[1344]&m[1345]&m[1346]&~m[1395]))&BiasedRNG[822])|(((m[1343]&~m[1344]&~m[1345]&~m[1346]&m[1395])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&m[1395])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&m[1395])|(m[1343]&m[1344]&~m[1345]&m[1346]&m[1395])|(m[1343]&~m[1344]&m[1345]&m[1346]&m[1395])|(~m[1343]&m[1344]&m[1345]&m[1346]&m[1395]))&~BiasedRNG[822])|((m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1395])|(m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1395])|(~m[1343]&m[1344]&m[1345]&~m[1346]&~m[1395])|(m[1343]&m[1344]&m[1345]&~m[1346]&~m[1395])|(m[1343]&m[1344]&m[1345]&m[1346]&~m[1395])|(m[1343]&m[1344]&~m[1345]&~m[1346]&m[1395])|(m[1343]&~m[1344]&m[1345]&~m[1346]&m[1395])|(~m[1343]&m[1344]&m[1345]&~m[1346]&m[1395])|(m[1343]&m[1344]&m[1345]&~m[1346]&m[1395])|(m[1343]&m[1344]&m[1345]&m[1346]&m[1395]))):InitCond[1538];
    m[1352] = run?((((m[1348]&~m[1349]&~m[1350]&~m[1351]&~m[1400])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1400])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1400])|(m[1348]&m[1349]&~m[1350]&m[1351]&~m[1400])|(m[1348]&~m[1349]&m[1350]&m[1351]&~m[1400])|(~m[1348]&m[1349]&m[1350]&m[1351]&~m[1400]))&BiasedRNG[823])|(((m[1348]&~m[1349]&~m[1350]&~m[1351]&m[1400])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&m[1400])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&m[1400])|(m[1348]&m[1349]&~m[1350]&m[1351]&m[1400])|(m[1348]&~m[1349]&m[1350]&m[1351]&m[1400])|(~m[1348]&m[1349]&m[1350]&m[1351]&m[1400]))&~BiasedRNG[823])|((m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1400])|(m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1400])|(~m[1348]&m[1349]&m[1350]&~m[1351]&~m[1400])|(m[1348]&m[1349]&m[1350]&~m[1351]&~m[1400])|(m[1348]&m[1349]&m[1350]&m[1351]&~m[1400])|(m[1348]&m[1349]&~m[1350]&~m[1351]&m[1400])|(m[1348]&~m[1349]&m[1350]&~m[1351]&m[1400])|(~m[1348]&m[1349]&m[1350]&~m[1351]&m[1400])|(m[1348]&m[1349]&m[1350]&~m[1351]&m[1400])|(m[1348]&m[1349]&m[1350]&m[1351]&m[1400]))):InitCond[1539];
    m[1357] = run?((((m[1353]&~m[1354]&~m[1355]&~m[1356]&~m[1405])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1405])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1405])|(m[1353]&m[1354]&~m[1355]&m[1356]&~m[1405])|(m[1353]&~m[1354]&m[1355]&m[1356]&~m[1405])|(~m[1353]&m[1354]&m[1355]&m[1356]&~m[1405]))&BiasedRNG[824])|(((m[1353]&~m[1354]&~m[1355]&~m[1356]&m[1405])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&m[1405])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&m[1405])|(m[1353]&m[1354]&~m[1355]&m[1356]&m[1405])|(m[1353]&~m[1354]&m[1355]&m[1356]&m[1405])|(~m[1353]&m[1354]&m[1355]&m[1356]&m[1405]))&~BiasedRNG[824])|((m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1405])|(m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1405])|(~m[1353]&m[1354]&m[1355]&~m[1356]&~m[1405])|(m[1353]&m[1354]&m[1355]&~m[1356]&~m[1405])|(m[1353]&m[1354]&m[1355]&m[1356]&~m[1405])|(m[1353]&m[1354]&~m[1355]&~m[1356]&m[1405])|(m[1353]&~m[1354]&m[1355]&~m[1356]&m[1405])|(~m[1353]&m[1354]&m[1355]&~m[1356]&m[1405])|(m[1353]&m[1354]&m[1355]&~m[1356]&m[1405])|(m[1353]&m[1354]&m[1355]&m[1356]&m[1405]))):InitCond[1540];
    m[1362] = run?((((m[1358]&~m[1359]&~m[1360]&~m[1361]&~m[1410])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1410])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1410])|(m[1358]&m[1359]&~m[1360]&m[1361]&~m[1410])|(m[1358]&~m[1359]&m[1360]&m[1361]&~m[1410])|(~m[1358]&m[1359]&m[1360]&m[1361]&~m[1410]))&BiasedRNG[825])|(((m[1358]&~m[1359]&~m[1360]&~m[1361]&m[1410])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&m[1410])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&m[1410])|(m[1358]&m[1359]&~m[1360]&m[1361]&m[1410])|(m[1358]&~m[1359]&m[1360]&m[1361]&m[1410])|(~m[1358]&m[1359]&m[1360]&m[1361]&m[1410]))&~BiasedRNG[825])|((m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1410])|(m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1410])|(~m[1358]&m[1359]&m[1360]&~m[1361]&~m[1410])|(m[1358]&m[1359]&m[1360]&~m[1361]&~m[1410])|(m[1358]&m[1359]&m[1360]&m[1361]&~m[1410])|(m[1358]&m[1359]&~m[1360]&~m[1361]&m[1410])|(m[1358]&~m[1359]&m[1360]&~m[1361]&m[1410])|(~m[1358]&m[1359]&m[1360]&~m[1361]&m[1410])|(m[1358]&m[1359]&m[1360]&~m[1361]&m[1410])|(m[1358]&m[1359]&m[1360]&m[1361]&m[1410]))):InitCond[1541];
    m[1367] = run?((((m[1363]&~m[1364]&~m[1365]&~m[1366]&~m[1413])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1413])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1413])|(m[1363]&m[1364]&~m[1365]&m[1366]&~m[1413])|(m[1363]&~m[1364]&m[1365]&m[1366]&~m[1413])|(~m[1363]&m[1364]&m[1365]&m[1366]&~m[1413]))&BiasedRNG[826])|(((m[1363]&~m[1364]&~m[1365]&~m[1366]&m[1413])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&m[1413])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&m[1413])|(m[1363]&m[1364]&~m[1365]&m[1366]&m[1413])|(m[1363]&~m[1364]&m[1365]&m[1366]&m[1413])|(~m[1363]&m[1364]&m[1365]&m[1366]&m[1413]))&~BiasedRNG[826])|((m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1413])|(m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1413])|(~m[1363]&m[1364]&m[1365]&~m[1366]&~m[1413])|(m[1363]&m[1364]&m[1365]&~m[1366]&~m[1413])|(m[1363]&m[1364]&m[1365]&m[1366]&~m[1413])|(m[1363]&m[1364]&~m[1365]&~m[1366]&m[1413])|(m[1363]&~m[1364]&m[1365]&~m[1366]&m[1413])|(~m[1363]&m[1364]&m[1365]&~m[1366]&m[1413])|(m[1363]&m[1364]&m[1365]&~m[1366]&m[1413])|(m[1363]&m[1364]&m[1365]&m[1366]&m[1413]))):InitCond[1542];
    m[1372] = run?((((m[1368]&~m[1369]&~m[1370]&~m[1371]&~m[1415])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1415])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1415])|(m[1368]&m[1369]&~m[1370]&m[1371]&~m[1415])|(m[1368]&~m[1369]&m[1370]&m[1371]&~m[1415])|(~m[1368]&m[1369]&m[1370]&m[1371]&~m[1415]))&BiasedRNG[827])|(((m[1368]&~m[1369]&~m[1370]&~m[1371]&m[1415])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&m[1415])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&m[1415])|(m[1368]&m[1369]&~m[1370]&m[1371]&m[1415])|(m[1368]&~m[1369]&m[1370]&m[1371]&m[1415])|(~m[1368]&m[1369]&m[1370]&m[1371]&m[1415]))&~BiasedRNG[827])|((m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1415])|(m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1415])|(~m[1368]&m[1369]&m[1370]&~m[1371]&~m[1415])|(m[1368]&m[1369]&m[1370]&~m[1371]&~m[1415])|(m[1368]&m[1369]&m[1370]&m[1371]&~m[1415])|(m[1368]&m[1369]&~m[1370]&~m[1371]&m[1415])|(m[1368]&~m[1369]&m[1370]&~m[1371]&m[1415])|(~m[1368]&m[1369]&m[1370]&~m[1371]&m[1415])|(m[1368]&m[1369]&m[1370]&~m[1371]&m[1415])|(m[1368]&m[1369]&m[1370]&m[1371]&m[1415]))):InitCond[1543];
    m[1377] = run?((((m[1373]&~m[1374]&~m[1375]&~m[1376]&~m[1420])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1420])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1420])|(m[1373]&m[1374]&~m[1375]&m[1376]&~m[1420])|(m[1373]&~m[1374]&m[1375]&m[1376]&~m[1420])|(~m[1373]&m[1374]&m[1375]&m[1376]&~m[1420]))&BiasedRNG[828])|(((m[1373]&~m[1374]&~m[1375]&~m[1376]&m[1420])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&m[1420])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&m[1420])|(m[1373]&m[1374]&~m[1375]&m[1376]&m[1420])|(m[1373]&~m[1374]&m[1375]&m[1376]&m[1420])|(~m[1373]&m[1374]&m[1375]&m[1376]&m[1420]))&~BiasedRNG[828])|((m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1420])|(m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1420])|(~m[1373]&m[1374]&m[1375]&~m[1376]&~m[1420])|(m[1373]&m[1374]&m[1375]&~m[1376]&~m[1420])|(m[1373]&m[1374]&m[1375]&m[1376]&~m[1420])|(m[1373]&m[1374]&~m[1375]&~m[1376]&m[1420])|(m[1373]&~m[1374]&m[1375]&~m[1376]&m[1420])|(~m[1373]&m[1374]&m[1375]&~m[1376]&m[1420])|(m[1373]&m[1374]&m[1375]&~m[1376]&m[1420])|(m[1373]&m[1374]&m[1375]&m[1376]&m[1420]))):InitCond[1544];
    m[1382] = run?((((m[1378]&~m[1379]&~m[1380]&~m[1381]&~m[1425])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1425])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1425])|(m[1378]&m[1379]&~m[1380]&m[1381]&~m[1425])|(m[1378]&~m[1379]&m[1380]&m[1381]&~m[1425])|(~m[1378]&m[1379]&m[1380]&m[1381]&~m[1425]))&BiasedRNG[829])|(((m[1378]&~m[1379]&~m[1380]&~m[1381]&m[1425])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&m[1425])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&m[1425])|(m[1378]&m[1379]&~m[1380]&m[1381]&m[1425])|(m[1378]&~m[1379]&m[1380]&m[1381]&m[1425])|(~m[1378]&m[1379]&m[1380]&m[1381]&m[1425]))&~BiasedRNG[829])|((m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1425])|(m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1425])|(~m[1378]&m[1379]&m[1380]&~m[1381]&~m[1425])|(m[1378]&m[1379]&m[1380]&~m[1381]&~m[1425])|(m[1378]&m[1379]&m[1380]&m[1381]&~m[1425])|(m[1378]&m[1379]&~m[1380]&~m[1381]&m[1425])|(m[1378]&~m[1379]&m[1380]&~m[1381]&m[1425])|(~m[1378]&m[1379]&m[1380]&~m[1381]&m[1425])|(m[1378]&m[1379]&m[1380]&~m[1381]&m[1425])|(m[1378]&m[1379]&m[1380]&m[1381]&m[1425]))):InitCond[1545];
    m[1387] = run?((((m[1383]&~m[1384]&~m[1385]&~m[1386]&~m[1430])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1430])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1430])|(m[1383]&m[1384]&~m[1385]&m[1386]&~m[1430])|(m[1383]&~m[1384]&m[1385]&m[1386]&~m[1430])|(~m[1383]&m[1384]&m[1385]&m[1386]&~m[1430]))&BiasedRNG[830])|(((m[1383]&~m[1384]&~m[1385]&~m[1386]&m[1430])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&m[1430])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&m[1430])|(m[1383]&m[1384]&~m[1385]&m[1386]&m[1430])|(m[1383]&~m[1384]&m[1385]&m[1386]&m[1430])|(~m[1383]&m[1384]&m[1385]&m[1386]&m[1430]))&~BiasedRNG[830])|((m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1430])|(m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1430])|(~m[1383]&m[1384]&m[1385]&~m[1386]&~m[1430])|(m[1383]&m[1384]&m[1385]&~m[1386]&~m[1430])|(m[1383]&m[1384]&m[1385]&m[1386]&~m[1430])|(m[1383]&m[1384]&~m[1385]&~m[1386]&m[1430])|(m[1383]&~m[1384]&m[1385]&~m[1386]&m[1430])|(~m[1383]&m[1384]&m[1385]&~m[1386]&m[1430])|(m[1383]&m[1384]&m[1385]&~m[1386]&m[1430])|(m[1383]&m[1384]&m[1385]&m[1386]&m[1430]))):InitCond[1546];
    m[1392] = run?((((m[1388]&~m[1389]&~m[1390]&~m[1391]&~m[1435])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1435])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1435])|(m[1388]&m[1389]&~m[1390]&m[1391]&~m[1435])|(m[1388]&~m[1389]&m[1390]&m[1391]&~m[1435])|(~m[1388]&m[1389]&m[1390]&m[1391]&~m[1435]))&BiasedRNG[831])|(((m[1388]&~m[1389]&~m[1390]&~m[1391]&m[1435])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&m[1435])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&m[1435])|(m[1388]&m[1389]&~m[1390]&m[1391]&m[1435])|(m[1388]&~m[1389]&m[1390]&m[1391]&m[1435])|(~m[1388]&m[1389]&m[1390]&m[1391]&m[1435]))&~BiasedRNG[831])|((m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1435])|(m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1435])|(~m[1388]&m[1389]&m[1390]&~m[1391]&~m[1435])|(m[1388]&m[1389]&m[1390]&~m[1391]&~m[1435])|(m[1388]&m[1389]&m[1390]&m[1391]&~m[1435])|(m[1388]&m[1389]&~m[1390]&~m[1391]&m[1435])|(m[1388]&~m[1389]&m[1390]&~m[1391]&m[1435])|(~m[1388]&m[1389]&m[1390]&~m[1391]&m[1435])|(m[1388]&m[1389]&m[1390]&~m[1391]&m[1435])|(m[1388]&m[1389]&m[1390]&m[1391]&m[1435]))):InitCond[1547];
    m[1397] = run?((((m[1393]&~m[1394]&~m[1395]&~m[1396]&~m[1440])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1440])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1440])|(m[1393]&m[1394]&~m[1395]&m[1396]&~m[1440])|(m[1393]&~m[1394]&m[1395]&m[1396]&~m[1440])|(~m[1393]&m[1394]&m[1395]&m[1396]&~m[1440]))&BiasedRNG[832])|(((m[1393]&~m[1394]&~m[1395]&~m[1396]&m[1440])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&m[1440])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&m[1440])|(m[1393]&m[1394]&~m[1395]&m[1396]&m[1440])|(m[1393]&~m[1394]&m[1395]&m[1396]&m[1440])|(~m[1393]&m[1394]&m[1395]&m[1396]&m[1440]))&~BiasedRNG[832])|((m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1440])|(m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1440])|(~m[1393]&m[1394]&m[1395]&~m[1396]&~m[1440])|(m[1393]&m[1394]&m[1395]&~m[1396]&~m[1440])|(m[1393]&m[1394]&m[1395]&m[1396]&~m[1440])|(m[1393]&m[1394]&~m[1395]&~m[1396]&m[1440])|(m[1393]&~m[1394]&m[1395]&~m[1396]&m[1440])|(~m[1393]&m[1394]&m[1395]&~m[1396]&m[1440])|(m[1393]&m[1394]&m[1395]&~m[1396]&m[1440])|(m[1393]&m[1394]&m[1395]&m[1396]&m[1440]))):InitCond[1548];
    m[1402] = run?((((m[1398]&~m[1399]&~m[1400]&~m[1401]&~m[1445])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1445])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1445])|(m[1398]&m[1399]&~m[1400]&m[1401]&~m[1445])|(m[1398]&~m[1399]&m[1400]&m[1401]&~m[1445])|(~m[1398]&m[1399]&m[1400]&m[1401]&~m[1445]))&BiasedRNG[833])|(((m[1398]&~m[1399]&~m[1400]&~m[1401]&m[1445])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&m[1445])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&m[1445])|(m[1398]&m[1399]&~m[1400]&m[1401]&m[1445])|(m[1398]&~m[1399]&m[1400]&m[1401]&m[1445])|(~m[1398]&m[1399]&m[1400]&m[1401]&m[1445]))&~BiasedRNG[833])|((m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1445])|(m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1445])|(~m[1398]&m[1399]&m[1400]&~m[1401]&~m[1445])|(m[1398]&m[1399]&m[1400]&~m[1401]&~m[1445])|(m[1398]&m[1399]&m[1400]&m[1401]&~m[1445])|(m[1398]&m[1399]&~m[1400]&~m[1401]&m[1445])|(m[1398]&~m[1399]&m[1400]&~m[1401]&m[1445])|(~m[1398]&m[1399]&m[1400]&~m[1401]&m[1445])|(m[1398]&m[1399]&m[1400]&~m[1401]&m[1445])|(m[1398]&m[1399]&m[1400]&m[1401]&m[1445]))):InitCond[1549];
    m[1407] = run?((((m[1403]&~m[1404]&~m[1405]&~m[1406]&~m[1450])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1450])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1450])|(m[1403]&m[1404]&~m[1405]&m[1406]&~m[1450])|(m[1403]&~m[1404]&m[1405]&m[1406]&~m[1450])|(~m[1403]&m[1404]&m[1405]&m[1406]&~m[1450]))&BiasedRNG[834])|(((m[1403]&~m[1404]&~m[1405]&~m[1406]&m[1450])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&m[1450])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&m[1450])|(m[1403]&m[1404]&~m[1405]&m[1406]&m[1450])|(m[1403]&~m[1404]&m[1405]&m[1406]&m[1450])|(~m[1403]&m[1404]&m[1405]&m[1406]&m[1450]))&~BiasedRNG[834])|((m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1450])|(m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1450])|(~m[1403]&m[1404]&m[1405]&~m[1406]&~m[1450])|(m[1403]&m[1404]&m[1405]&~m[1406]&~m[1450])|(m[1403]&m[1404]&m[1405]&m[1406]&~m[1450])|(m[1403]&m[1404]&~m[1405]&~m[1406]&m[1450])|(m[1403]&~m[1404]&m[1405]&~m[1406]&m[1450])|(~m[1403]&m[1404]&m[1405]&~m[1406]&m[1450])|(m[1403]&m[1404]&m[1405]&~m[1406]&m[1450])|(m[1403]&m[1404]&m[1405]&m[1406]&m[1450]))):InitCond[1550];
    m[1412] = run?((((m[1408]&~m[1409]&~m[1410]&~m[1411]&~m[1455])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1455])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1455])|(m[1408]&m[1409]&~m[1410]&m[1411]&~m[1455])|(m[1408]&~m[1409]&m[1410]&m[1411]&~m[1455])|(~m[1408]&m[1409]&m[1410]&m[1411]&~m[1455]))&BiasedRNG[835])|(((m[1408]&~m[1409]&~m[1410]&~m[1411]&m[1455])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&m[1455])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&m[1455])|(m[1408]&m[1409]&~m[1410]&m[1411]&m[1455])|(m[1408]&~m[1409]&m[1410]&m[1411]&m[1455])|(~m[1408]&m[1409]&m[1410]&m[1411]&m[1455]))&~BiasedRNG[835])|((m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1455])|(m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1455])|(~m[1408]&m[1409]&m[1410]&~m[1411]&~m[1455])|(m[1408]&m[1409]&m[1410]&~m[1411]&~m[1455])|(m[1408]&m[1409]&m[1410]&m[1411]&~m[1455])|(m[1408]&m[1409]&~m[1410]&~m[1411]&m[1455])|(m[1408]&~m[1409]&m[1410]&~m[1411]&m[1455])|(~m[1408]&m[1409]&m[1410]&~m[1411]&m[1455])|(m[1408]&m[1409]&m[1410]&~m[1411]&m[1455])|(m[1408]&m[1409]&m[1410]&m[1411]&m[1455]))):InitCond[1551];
    m[1417] = run?((((m[1413]&~m[1414]&~m[1415]&~m[1416]&~m[1458])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1458])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1458])|(m[1413]&m[1414]&~m[1415]&m[1416]&~m[1458])|(m[1413]&~m[1414]&m[1415]&m[1416]&~m[1458])|(~m[1413]&m[1414]&m[1415]&m[1416]&~m[1458]))&BiasedRNG[836])|(((m[1413]&~m[1414]&~m[1415]&~m[1416]&m[1458])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&m[1458])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&m[1458])|(m[1413]&m[1414]&~m[1415]&m[1416]&m[1458])|(m[1413]&~m[1414]&m[1415]&m[1416]&m[1458])|(~m[1413]&m[1414]&m[1415]&m[1416]&m[1458]))&~BiasedRNG[836])|((m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1458])|(m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1458])|(~m[1413]&m[1414]&m[1415]&~m[1416]&~m[1458])|(m[1413]&m[1414]&m[1415]&~m[1416]&~m[1458])|(m[1413]&m[1414]&m[1415]&m[1416]&~m[1458])|(m[1413]&m[1414]&~m[1415]&~m[1416]&m[1458])|(m[1413]&~m[1414]&m[1415]&~m[1416]&m[1458])|(~m[1413]&m[1414]&m[1415]&~m[1416]&m[1458])|(m[1413]&m[1414]&m[1415]&~m[1416]&m[1458])|(m[1413]&m[1414]&m[1415]&m[1416]&m[1458]))):InitCond[1552];
    m[1422] = run?((((m[1418]&~m[1419]&~m[1420]&~m[1421]&~m[1460])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1460])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1460])|(m[1418]&m[1419]&~m[1420]&m[1421]&~m[1460])|(m[1418]&~m[1419]&m[1420]&m[1421]&~m[1460])|(~m[1418]&m[1419]&m[1420]&m[1421]&~m[1460]))&BiasedRNG[837])|(((m[1418]&~m[1419]&~m[1420]&~m[1421]&m[1460])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&m[1460])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&m[1460])|(m[1418]&m[1419]&~m[1420]&m[1421]&m[1460])|(m[1418]&~m[1419]&m[1420]&m[1421]&m[1460])|(~m[1418]&m[1419]&m[1420]&m[1421]&m[1460]))&~BiasedRNG[837])|((m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1460])|(m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1460])|(~m[1418]&m[1419]&m[1420]&~m[1421]&~m[1460])|(m[1418]&m[1419]&m[1420]&~m[1421]&~m[1460])|(m[1418]&m[1419]&m[1420]&m[1421]&~m[1460])|(m[1418]&m[1419]&~m[1420]&~m[1421]&m[1460])|(m[1418]&~m[1419]&m[1420]&~m[1421]&m[1460])|(~m[1418]&m[1419]&m[1420]&~m[1421]&m[1460])|(m[1418]&m[1419]&m[1420]&~m[1421]&m[1460])|(m[1418]&m[1419]&m[1420]&m[1421]&m[1460]))):InitCond[1553];
    m[1427] = run?((((m[1423]&~m[1424]&~m[1425]&~m[1426]&~m[1465])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1465])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1465])|(m[1423]&m[1424]&~m[1425]&m[1426]&~m[1465])|(m[1423]&~m[1424]&m[1425]&m[1426]&~m[1465])|(~m[1423]&m[1424]&m[1425]&m[1426]&~m[1465]))&BiasedRNG[838])|(((m[1423]&~m[1424]&~m[1425]&~m[1426]&m[1465])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&m[1465])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&m[1465])|(m[1423]&m[1424]&~m[1425]&m[1426]&m[1465])|(m[1423]&~m[1424]&m[1425]&m[1426]&m[1465])|(~m[1423]&m[1424]&m[1425]&m[1426]&m[1465]))&~BiasedRNG[838])|((m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1465])|(m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1465])|(~m[1423]&m[1424]&m[1425]&~m[1426]&~m[1465])|(m[1423]&m[1424]&m[1425]&~m[1426]&~m[1465])|(m[1423]&m[1424]&m[1425]&m[1426]&~m[1465])|(m[1423]&m[1424]&~m[1425]&~m[1426]&m[1465])|(m[1423]&~m[1424]&m[1425]&~m[1426]&m[1465])|(~m[1423]&m[1424]&m[1425]&~m[1426]&m[1465])|(m[1423]&m[1424]&m[1425]&~m[1426]&m[1465])|(m[1423]&m[1424]&m[1425]&m[1426]&m[1465]))):InitCond[1554];
    m[1432] = run?((((m[1428]&~m[1429]&~m[1430]&~m[1431]&~m[1470])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1470])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1470])|(m[1428]&m[1429]&~m[1430]&m[1431]&~m[1470])|(m[1428]&~m[1429]&m[1430]&m[1431]&~m[1470])|(~m[1428]&m[1429]&m[1430]&m[1431]&~m[1470]))&BiasedRNG[839])|(((m[1428]&~m[1429]&~m[1430]&~m[1431]&m[1470])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&m[1470])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&m[1470])|(m[1428]&m[1429]&~m[1430]&m[1431]&m[1470])|(m[1428]&~m[1429]&m[1430]&m[1431]&m[1470])|(~m[1428]&m[1429]&m[1430]&m[1431]&m[1470]))&~BiasedRNG[839])|((m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1470])|(m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1470])|(~m[1428]&m[1429]&m[1430]&~m[1431]&~m[1470])|(m[1428]&m[1429]&m[1430]&~m[1431]&~m[1470])|(m[1428]&m[1429]&m[1430]&m[1431]&~m[1470])|(m[1428]&m[1429]&~m[1430]&~m[1431]&m[1470])|(m[1428]&~m[1429]&m[1430]&~m[1431]&m[1470])|(~m[1428]&m[1429]&m[1430]&~m[1431]&m[1470])|(m[1428]&m[1429]&m[1430]&~m[1431]&m[1470])|(m[1428]&m[1429]&m[1430]&m[1431]&m[1470]))):InitCond[1555];
    m[1437] = run?((((m[1433]&~m[1434]&~m[1435]&~m[1436]&~m[1475])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1475])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1475])|(m[1433]&m[1434]&~m[1435]&m[1436]&~m[1475])|(m[1433]&~m[1434]&m[1435]&m[1436]&~m[1475])|(~m[1433]&m[1434]&m[1435]&m[1436]&~m[1475]))&BiasedRNG[840])|(((m[1433]&~m[1434]&~m[1435]&~m[1436]&m[1475])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&m[1475])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&m[1475])|(m[1433]&m[1434]&~m[1435]&m[1436]&m[1475])|(m[1433]&~m[1434]&m[1435]&m[1436]&m[1475])|(~m[1433]&m[1434]&m[1435]&m[1436]&m[1475]))&~BiasedRNG[840])|((m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1475])|(m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1475])|(~m[1433]&m[1434]&m[1435]&~m[1436]&~m[1475])|(m[1433]&m[1434]&m[1435]&~m[1436]&~m[1475])|(m[1433]&m[1434]&m[1435]&m[1436]&~m[1475])|(m[1433]&m[1434]&~m[1435]&~m[1436]&m[1475])|(m[1433]&~m[1434]&m[1435]&~m[1436]&m[1475])|(~m[1433]&m[1434]&m[1435]&~m[1436]&m[1475])|(m[1433]&m[1434]&m[1435]&~m[1436]&m[1475])|(m[1433]&m[1434]&m[1435]&m[1436]&m[1475]))):InitCond[1556];
    m[1442] = run?((((m[1438]&~m[1439]&~m[1440]&~m[1441]&~m[1480])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1480])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1480])|(m[1438]&m[1439]&~m[1440]&m[1441]&~m[1480])|(m[1438]&~m[1439]&m[1440]&m[1441]&~m[1480])|(~m[1438]&m[1439]&m[1440]&m[1441]&~m[1480]))&BiasedRNG[841])|(((m[1438]&~m[1439]&~m[1440]&~m[1441]&m[1480])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&m[1480])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&m[1480])|(m[1438]&m[1439]&~m[1440]&m[1441]&m[1480])|(m[1438]&~m[1439]&m[1440]&m[1441]&m[1480])|(~m[1438]&m[1439]&m[1440]&m[1441]&m[1480]))&~BiasedRNG[841])|((m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1480])|(m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1480])|(~m[1438]&m[1439]&m[1440]&~m[1441]&~m[1480])|(m[1438]&m[1439]&m[1440]&~m[1441]&~m[1480])|(m[1438]&m[1439]&m[1440]&m[1441]&~m[1480])|(m[1438]&m[1439]&~m[1440]&~m[1441]&m[1480])|(m[1438]&~m[1439]&m[1440]&~m[1441]&m[1480])|(~m[1438]&m[1439]&m[1440]&~m[1441]&m[1480])|(m[1438]&m[1439]&m[1440]&~m[1441]&m[1480])|(m[1438]&m[1439]&m[1440]&m[1441]&m[1480]))):InitCond[1557];
    m[1447] = run?((((m[1443]&~m[1444]&~m[1445]&~m[1446]&~m[1485])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1485])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1485])|(m[1443]&m[1444]&~m[1445]&m[1446]&~m[1485])|(m[1443]&~m[1444]&m[1445]&m[1446]&~m[1485])|(~m[1443]&m[1444]&m[1445]&m[1446]&~m[1485]))&BiasedRNG[842])|(((m[1443]&~m[1444]&~m[1445]&~m[1446]&m[1485])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&m[1485])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&m[1485])|(m[1443]&m[1444]&~m[1445]&m[1446]&m[1485])|(m[1443]&~m[1444]&m[1445]&m[1446]&m[1485])|(~m[1443]&m[1444]&m[1445]&m[1446]&m[1485]))&~BiasedRNG[842])|((m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1485])|(m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1485])|(~m[1443]&m[1444]&m[1445]&~m[1446]&~m[1485])|(m[1443]&m[1444]&m[1445]&~m[1446]&~m[1485])|(m[1443]&m[1444]&m[1445]&m[1446]&~m[1485])|(m[1443]&m[1444]&~m[1445]&~m[1446]&m[1485])|(m[1443]&~m[1444]&m[1445]&~m[1446]&m[1485])|(~m[1443]&m[1444]&m[1445]&~m[1446]&m[1485])|(m[1443]&m[1444]&m[1445]&~m[1446]&m[1485])|(m[1443]&m[1444]&m[1445]&m[1446]&m[1485]))):InitCond[1558];
    m[1452] = run?((((m[1448]&~m[1449]&~m[1450]&~m[1451]&~m[1490])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1490])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1490])|(m[1448]&m[1449]&~m[1450]&m[1451]&~m[1490])|(m[1448]&~m[1449]&m[1450]&m[1451]&~m[1490])|(~m[1448]&m[1449]&m[1450]&m[1451]&~m[1490]))&BiasedRNG[843])|(((m[1448]&~m[1449]&~m[1450]&~m[1451]&m[1490])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&m[1490])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&m[1490])|(m[1448]&m[1449]&~m[1450]&m[1451]&m[1490])|(m[1448]&~m[1449]&m[1450]&m[1451]&m[1490])|(~m[1448]&m[1449]&m[1450]&m[1451]&m[1490]))&~BiasedRNG[843])|((m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1490])|(m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1490])|(~m[1448]&m[1449]&m[1450]&~m[1451]&~m[1490])|(m[1448]&m[1449]&m[1450]&~m[1451]&~m[1490])|(m[1448]&m[1449]&m[1450]&m[1451]&~m[1490])|(m[1448]&m[1449]&~m[1450]&~m[1451]&m[1490])|(m[1448]&~m[1449]&m[1450]&~m[1451]&m[1490])|(~m[1448]&m[1449]&m[1450]&~m[1451]&m[1490])|(m[1448]&m[1449]&m[1450]&~m[1451]&m[1490])|(m[1448]&m[1449]&m[1450]&m[1451]&m[1490]))):InitCond[1559];
    m[1457] = run?((((m[1453]&~m[1454]&~m[1455]&~m[1456]&~m[1495])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1495])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1495])|(m[1453]&m[1454]&~m[1455]&m[1456]&~m[1495])|(m[1453]&~m[1454]&m[1455]&m[1456]&~m[1495])|(~m[1453]&m[1454]&m[1455]&m[1456]&~m[1495]))&BiasedRNG[844])|(((m[1453]&~m[1454]&~m[1455]&~m[1456]&m[1495])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&m[1495])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&m[1495])|(m[1453]&m[1454]&~m[1455]&m[1456]&m[1495])|(m[1453]&~m[1454]&m[1455]&m[1456]&m[1495])|(~m[1453]&m[1454]&m[1455]&m[1456]&m[1495]))&~BiasedRNG[844])|((m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1495])|(m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1495])|(~m[1453]&m[1454]&m[1455]&~m[1456]&~m[1495])|(m[1453]&m[1454]&m[1455]&~m[1456]&~m[1495])|(m[1453]&m[1454]&m[1455]&m[1456]&~m[1495])|(m[1453]&m[1454]&~m[1455]&~m[1456]&m[1495])|(m[1453]&~m[1454]&m[1455]&~m[1456]&m[1495])|(~m[1453]&m[1454]&m[1455]&~m[1456]&m[1495])|(m[1453]&m[1454]&m[1455]&~m[1456]&m[1495])|(m[1453]&m[1454]&m[1455]&m[1456]&m[1495]))):InitCond[1560];
    m[1462] = run?((((m[1458]&~m[1459]&~m[1460]&~m[1461]&~m[1498])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1498])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1498])|(m[1458]&m[1459]&~m[1460]&m[1461]&~m[1498])|(m[1458]&~m[1459]&m[1460]&m[1461]&~m[1498])|(~m[1458]&m[1459]&m[1460]&m[1461]&~m[1498]))&BiasedRNG[845])|(((m[1458]&~m[1459]&~m[1460]&~m[1461]&m[1498])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&m[1498])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&m[1498])|(m[1458]&m[1459]&~m[1460]&m[1461]&m[1498])|(m[1458]&~m[1459]&m[1460]&m[1461]&m[1498])|(~m[1458]&m[1459]&m[1460]&m[1461]&m[1498]))&~BiasedRNG[845])|((m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1498])|(m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1498])|(~m[1458]&m[1459]&m[1460]&~m[1461]&~m[1498])|(m[1458]&m[1459]&m[1460]&~m[1461]&~m[1498])|(m[1458]&m[1459]&m[1460]&m[1461]&~m[1498])|(m[1458]&m[1459]&~m[1460]&~m[1461]&m[1498])|(m[1458]&~m[1459]&m[1460]&~m[1461]&m[1498])|(~m[1458]&m[1459]&m[1460]&~m[1461]&m[1498])|(m[1458]&m[1459]&m[1460]&~m[1461]&m[1498])|(m[1458]&m[1459]&m[1460]&m[1461]&m[1498]))):InitCond[1561];
    m[1467] = run?((((m[1463]&~m[1464]&~m[1465]&~m[1466]&~m[1500])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1500])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1500])|(m[1463]&m[1464]&~m[1465]&m[1466]&~m[1500])|(m[1463]&~m[1464]&m[1465]&m[1466]&~m[1500])|(~m[1463]&m[1464]&m[1465]&m[1466]&~m[1500]))&BiasedRNG[846])|(((m[1463]&~m[1464]&~m[1465]&~m[1466]&m[1500])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&m[1500])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&m[1500])|(m[1463]&m[1464]&~m[1465]&m[1466]&m[1500])|(m[1463]&~m[1464]&m[1465]&m[1466]&m[1500])|(~m[1463]&m[1464]&m[1465]&m[1466]&m[1500]))&~BiasedRNG[846])|((m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1500])|(m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1500])|(~m[1463]&m[1464]&m[1465]&~m[1466]&~m[1500])|(m[1463]&m[1464]&m[1465]&~m[1466]&~m[1500])|(m[1463]&m[1464]&m[1465]&m[1466]&~m[1500])|(m[1463]&m[1464]&~m[1465]&~m[1466]&m[1500])|(m[1463]&~m[1464]&m[1465]&~m[1466]&m[1500])|(~m[1463]&m[1464]&m[1465]&~m[1466]&m[1500])|(m[1463]&m[1464]&m[1465]&~m[1466]&m[1500])|(m[1463]&m[1464]&m[1465]&m[1466]&m[1500]))):InitCond[1562];
    m[1472] = run?((((m[1468]&~m[1469]&~m[1470]&~m[1471]&~m[1505])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1505])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1505])|(m[1468]&m[1469]&~m[1470]&m[1471]&~m[1505])|(m[1468]&~m[1469]&m[1470]&m[1471]&~m[1505])|(~m[1468]&m[1469]&m[1470]&m[1471]&~m[1505]))&BiasedRNG[847])|(((m[1468]&~m[1469]&~m[1470]&~m[1471]&m[1505])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&m[1505])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&m[1505])|(m[1468]&m[1469]&~m[1470]&m[1471]&m[1505])|(m[1468]&~m[1469]&m[1470]&m[1471]&m[1505])|(~m[1468]&m[1469]&m[1470]&m[1471]&m[1505]))&~BiasedRNG[847])|((m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1505])|(m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1505])|(~m[1468]&m[1469]&m[1470]&~m[1471]&~m[1505])|(m[1468]&m[1469]&m[1470]&~m[1471]&~m[1505])|(m[1468]&m[1469]&m[1470]&m[1471]&~m[1505])|(m[1468]&m[1469]&~m[1470]&~m[1471]&m[1505])|(m[1468]&~m[1469]&m[1470]&~m[1471]&m[1505])|(~m[1468]&m[1469]&m[1470]&~m[1471]&m[1505])|(m[1468]&m[1469]&m[1470]&~m[1471]&m[1505])|(m[1468]&m[1469]&m[1470]&m[1471]&m[1505]))):InitCond[1563];
    m[1477] = run?((((m[1473]&~m[1474]&~m[1475]&~m[1476]&~m[1510])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1510])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1510])|(m[1473]&m[1474]&~m[1475]&m[1476]&~m[1510])|(m[1473]&~m[1474]&m[1475]&m[1476]&~m[1510])|(~m[1473]&m[1474]&m[1475]&m[1476]&~m[1510]))&BiasedRNG[848])|(((m[1473]&~m[1474]&~m[1475]&~m[1476]&m[1510])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&m[1510])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&m[1510])|(m[1473]&m[1474]&~m[1475]&m[1476]&m[1510])|(m[1473]&~m[1474]&m[1475]&m[1476]&m[1510])|(~m[1473]&m[1474]&m[1475]&m[1476]&m[1510]))&~BiasedRNG[848])|((m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1510])|(m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1510])|(~m[1473]&m[1474]&m[1475]&~m[1476]&~m[1510])|(m[1473]&m[1474]&m[1475]&~m[1476]&~m[1510])|(m[1473]&m[1474]&m[1475]&m[1476]&~m[1510])|(m[1473]&m[1474]&~m[1475]&~m[1476]&m[1510])|(m[1473]&~m[1474]&m[1475]&~m[1476]&m[1510])|(~m[1473]&m[1474]&m[1475]&~m[1476]&m[1510])|(m[1473]&m[1474]&m[1475]&~m[1476]&m[1510])|(m[1473]&m[1474]&m[1475]&m[1476]&m[1510]))):InitCond[1564];
    m[1482] = run?((((m[1478]&~m[1479]&~m[1480]&~m[1481]&~m[1515])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1515])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1515])|(m[1478]&m[1479]&~m[1480]&m[1481]&~m[1515])|(m[1478]&~m[1479]&m[1480]&m[1481]&~m[1515])|(~m[1478]&m[1479]&m[1480]&m[1481]&~m[1515]))&BiasedRNG[849])|(((m[1478]&~m[1479]&~m[1480]&~m[1481]&m[1515])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&m[1515])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&m[1515])|(m[1478]&m[1479]&~m[1480]&m[1481]&m[1515])|(m[1478]&~m[1479]&m[1480]&m[1481]&m[1515])|(~m[1478]&m[1479]&m[1480]&m[1481]&m[1515]))&~BiasedRNG[849])|((m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1515])|(m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1515])|(~m[1478]&m[1479]&m[1480]&~m[1481]&~m[1515])|(m[1478]&m[1479]&m[1480]&~m[1481]&~m[1515])|(m[1478]&m[1479]&m[1480]&m[1481]&~m[1515])|(m[1478]&m[1479]&~m[1480]&~m[1481]&m[1515])|(m[1478]&~m[1479]&m[1480]&~m[1481]&m[1515])|(~m[1478]&m[1479]&m[1480]&~m[1481]&m[1515])|(m[1478]&m[1479]&m[1480]&~m[1481]&m[1515])|(m[1478]&m[1479]&m[1480]&m[1481]&m[1515]))):InitCond[1565];
    m[1487] = run?((((m[1483]&~m[1484]&~m[1485]&~m[1486]&~m[1520])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1520])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1520])|(m[1483]&m[1484]&~m[1485]&m[1486]&~m[1520])|(m[1483]&~m[1484]&m[1485]&m[1486]&~m[1520])|(~m[1483]&m[1484]&m[1485]&m[1486]&~m[1520]))&BiasedRNG[850])|(((m[1483]&~m[1484]&~m[1485]&~m[1486]&m[1520])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&m[1520])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&m[1520])|(m[1483]&m[1484]&~m[1485]&m[1486]&m[1520])|(m[1483]&~m[1484]&m[1485]&m[1486]&m[1520])|(~m[1483]&m[1484]&m[1485]&m[1486]&m[1520]))&~BiasedRNG[850])|((m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1520])|(m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1520])|(~m[1483]&m[1484]&m[1485]&~m[1486]&~m[1520])|(m[1483]&m[1484]&m[1485]&~m[1486]&~m[1520])|(m[1483]&m[1484]&m[1485]&m[1486]&~m[1520])|(m[1483]&m[1484]&~m[1485]&~m[1486]&m[1520])|(m[1483]&~m[1484]&m[1485]&~m[1486]&m[1520])|(~m[1483]&m[1484]&m[1485]&~m[1486]&m[1520])|(m[1483]&m[1484]&m[1485]&~m[1486]&m[1520])|(m[1483]&m[1484]&m[1485]&m[1486]&m[1520]))):InitCond[1566];
    m[1492] = run?((((m[1488]&~m[1489]&~m[1490]&~m[1491]&~m[1525])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1525])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1525])|(m[1488]&m[1489]&~m[1490]&m[1491]&~m[1525])|(m[1488]&~m[1489]&m[1490]&m[1491]&~m[1525])|(~m[1488]&m[1489]&m[1490]&m[1491]&~m[1525]))&BiasedRNG[851])|(((m[1488]&~m[1489]&~m[1490]&~m[1491]&m[1525])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&m[1525])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&m[1525])|(m[1488]&m[1489]&~m[1490]&m[1491]&m[1525])|(m[1488]&~m[1489]&m[1490]&m[1491]&m[1525])|(~m[1488]&m[1489]&m[1490]&m[1491]&m[1525]))&~BiasedRNG[851])|((m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1525])|(m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1525])|(~m[1488]&m[1489]&m[1490]&~m[1491]&~m[1525])|(m[1488]&m[1489]&m[1490]&~m[1491]&~m[1525])|(m[1488]&m[1489]&m[1490]&m[1491]&~m[1525])|(m[1488]&m[1489]&~m[1490]&~m[1491]&m[1525])|(m[1488]&~m[1489]&m[1490]&~m[1491]&m[1525])|(~m[1488]&m[1489]&m[1490]&~m[1491]&m[1525])|(m[1488]&m[1489]&m[1490]&~m[1491]&m[1525])|(m[1488]&m[1489]&m[1490]&m[1491]&m[1525]))):InitCond[1567];
    m[1497] = run?((((m[1493]&~m[1494]&~m[1495]&~m[1496]&~m[1530])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1530])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1530])|(m[1493]&m[1494]&~m[1495]&m[1496]&~m[1530])|(m[1493]&~m[1494]&m[1495]&m[1496]&~m[1530])|(~m[1493]&m[1494]&m[1495]&m[1496]&~m[1530]))&BiasedRNG[852])|(((m[1493]&~m[1494]&~m[1495]&~m[1496]&m[1530])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&m[1530])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&m[1530])|(m[1493]&m[1494]&~m[1495]&m[1496]&m[1530])|(m[1493]&~m[1494]&m[1495]&m[1496]&m[1530])|(~m[1493]&m[1494]&m[1495]&m[1496]&m[1530]))&~BiasedRNG[852])|((m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1530])|(m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1530])|(~m[1493]&m[1494]&m[1495]&~m[1496]&~m[1530])|(m[1493]&m[1494]&m[1495]&~m[1496]&~m[1530])|(m[1493]&m[1494]&m[1495]&m[1496]&~m[1530])|(m[1493]&m[1494]&~m[1495]&~m[1496]&m[1530])|(m[1493]&~m[1494]&m[1495]&~m[1496]&m[1530])|(~m[1493]&m[1494]&m[1495]&~m[1496]&m[1530])|(m[1493]&m[1494]&m[1495]&~m[1496]&m[1530])|(m[1493]&m[1494]&m[1495]&m[1496]&m[1530]))):InitCond[1568];
    m[1502] = run?((((m[1498]&~m[1499]&~m[1500]&~m[1501]&~m[1533])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1533])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1533])|(m[1498]&m[1499]&~m[1500]&m[1501]&~m[1533])|(m[1498]&~m[1499]&m[1500]&m[1501]&~m[1533])|(~m[1498]&m[1499]&m[1500]&m[1501]&~m[1533]))&BiasedRNG[853])|(((m[1498]&~m[1499]&~m[1500]&~m[1501]&m[1533])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&m[1533])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&m[1533])|(m[1498]&m[1499]&~m[1500]&m[1501]&m[1533])|(m[1498]&~m[1499]&m[1500]&m[1501]&m[1533])|(~m[1498]&m[1499]&m[1500]&m[1501]&m[1533]))&~BiasedRNG[853])|((m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1533])|(m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1533])|(~m[1498]&m[1499]&m[1500]&~m[1501]&~m[1533])|(m[1498]&m[1499]&m[1500]&~m[1501]&~m[1533])|(m[1498]&m[1499]&m[1500]&m[1501]&~m[1533])|(m[1498]&m[1499]&~m[1500]&~m[1501]&m[1533])|(m[1498]&~m[1499]&m[1500]&~m[1501]&m[1533])|(~m[1498]&m[1499]&m[1500]&~m[1501]&m[1533])|(m[1498]&m[1499]&m[1500]&~m[1501]&m[1533])|(m[1498]&m[1499]&m[1500]&m[1501]&m[1533]))):InitCond[1569];
    m[1507] = run?((((m[1503]&~m[1504]&~m[1505]&~m[1506]&~m[1535])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1535])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1535])|(m[1503]&m[1504]&~m[1505]&m[1506]&~m[1535])|(m[1503]&~m[1504]&m[1505]&m[1506]&~m[1535])|(~m[1503]&m[1504]&m[1505]&m[1506]&~m[1535]))&BiasedRNG[854])|(((m[1503]&~m[1504]&~m[1505]&~m[1506]&m[1535])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&m[1535])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&m[1535])|(m[1503]&m[1504]&~m[1505]&m[1506]&m[1535])|(m[1503]&~m[1504]&m[1505]&m[1506]&m[1535])|(~m[1503]&m[1504]&m[1505]&m[1506]&m[1535]))&~BiasedRNG[854])|((m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1535])|(m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1535])|(~m[1503]&m[1504]&m[1505]&~m[1506]&~m[1535])|(m[1503]&m[1504]&m[1505]&~m[1506]&~m[1535])|(m[1503]&m[1504]&m[1505]&m[1506]&~m[1535])|(m[1503]&m[1504]&~m[1505]&~m[1506]&m[1535])|(m[1503]&~m[1504]&m[1505]&~m[1506]&m[1535])|(~m[1503]&m[1504]&m[1505]&~m[1506]&m[1535])|(m[1503]&m[1504]&m[1505]&~m[1506]&m[1535])|(m[1503]&m[1504]&m[1505]&m[1506]&m[1535]))):InitCond[1570];
    m[1512] = run?((((m[1508]&~m[1509]&~m[1510]&~m[1511]&~m[1540])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1540])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1540])|(m[1508]&m[1509]&~m[1510]&m[1511]&~m[1540])|(m[1508]&~m[1509]&m[1510]&m[1511]&~m[1540])|(~m[1508]&m[1509]&m[1510]&m[1511]&~m[1540]))&BiasedRNG[855])|(((m[1508]&~m[1509]&~m[1510]&~m[1511]&m[1540])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&m[1540])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&m[1540])|(m[1508]&m[1509]&~m[1510]&m[1511]&m[1540])|(m[1508]&~m[1509]&m[1510]&m[1511]&m[1540])|(~m[1508]&m[1509]&m[1510]&m[1511]&m[1540]))&~BiasedRNG[855])|((m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1540])|(m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1540])|(~m[1508]&m[1509]&m[1510]&~m[1511]&~m[1540])|(m[1508]&m[1509]&m[1510]&~m[1511]&~m[1540])|(m[1508]&m[1509]&m[1510]&m[1511]&~m[1540])|(m[1508]&m[1509]&~m[1510]&~m[1511]&m[1540])|(m[1508]&~m[1509]&m[1510]&~m[1511]&m[1540])|(~m[1508]&m[1509]&m[1510]&~m[1511]&m[1540])|(m[1508]&m[1509]&m[1510]&~m[1511]&m[1540])|(m[1508]&m[1509]&m[1510]&m[1511]&m[1540]))):InitCond[1571];
    m[1517] = run?((((m[1513]&~m[1514]&~m[1515]&~m[1516]&~m[1545])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1545])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1545])|(m[1513]&m[1514]&~m[1515]&m[1516]&~m[1545])|(m[1513]&~m[1514]&m[1515]&m[1516]&~m[1545])|(~m[1513]&m[1514]&m[1515]&m[1516]&~m[1545]))&BiasedRNG[856])|(((m[1513]&~m[1514]&~m[1515]&~m[1516]&m[1545])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&m[1545])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&m[1545])|(m[1513]&m[1514]&~m[1515]&m[1516]&m[1545])|(m[1513]&~m[1514]&m[1515]&m[1516]&m[1545])|(~m[1513]&m[1514]&m[1515]&m[1516]&m[1545]))&~BiasedRNG[856])|((m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1545])|(m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1545])|(~m[1513]&m[1514]&m[1515]&~m[1516]&~m[1545])|(m[1513]&m[1514]&m[1515]&~m[1516]&~m[1545])|(m[1513]&m[1514]&m[1515]&m[1516]&~m[1545])|(m[1513]&m[1514]&~m[1515]&~m[1516]&m[1545])|(m[1513]&~m[1514]&m[1515]&~m[1516]&m[1545])|(~m[1513]&m[1514]&m[1515]&~m[1516]&m[1545])|(m[1513]&m[1514]&m[1515]&~m[1516]&m[1545])|(m[1513]&m[1514]&m[1515]&m[1516]&m[1545]))):InitCond[1572];
    m[1522] = run?((((m[1518]&~m[1519]&~m[1520]&~m[1521]&~m[1550])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1550])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1550])|(m[1518]&m[1519]&~m[1520]&m[1521]&~m[1550])|(m[1518]&~m[1519]&m[1520]&m[1521]&~m[1550])|(~m[1518]&m[1519]&m[1520]&m[1521]&~m[1550]))&BiasedRNG[857])|(((m[1518]&~m[1519]&~m[1520]&~m[1521]&m[1550])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&m[1550])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&m[1550])|(m[1518]&m[1519]&~m[1520]&m[1521]&m[1550])|(m[1518]&~m[1519]&m[1520]&m[1521]&m[1550])|(~m[1518]&m[1519]&m[1520]&m[1521]&m[1550]))&~BiasedRNG[857])|((m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1550])|(m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1550])|(~m[1518]&m[1519]&m[1520]&~m[1521]&~m[1550])|(m[1518]&m[1519]&m[1520]&~m[1521]&~m[1550])|(m[1518]&m[1519]&m[1520]&m[1521]&~m[1550])|(m[1518]&m[1519]&~m[1520]&~m[1521]&m[1550])|(m[1518]&~m[1519]&m[1520]&~m[1521]&m[1550])|(~m[1518]&m[1519]&m[1520]&~m[1521]&m[1550])|(m[1518]&m[1519]&m[1520]&~m[1521]&m[1550])|(m[1518]&m[1519]&m[1520]&m[1521]&m[1550]))):InitCond[1573];
    m[1527] = run?((((m[1523]&~m[1524]&~m[1525]&~m[1526]&~m[1555])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1555])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1555])|(m[1523]&m[1524]&~m[1525]&m[1526]&~m[1555])|(m[1523]&~m[1524]&m[1525]&m[1526]&~m[1555])|(~m[1523]&m[1524]&m[1525]&m[1526]&~m[1555]))&BiasedRNG[858])|(((m[1523]&~m[1524]&~m[1525]&~m[1526]&m[1555])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&m[1555])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&m[1555])|(m[1523]&m[1524]&~m[1525]&m[1526]&m[1555])|(m[1523]&~m[1524]&m[1525]&m[1526]&m[1555])|(~m[1523]&m[1524]&m[1525]&m[1526]&m[1555]))&~BiasedRNG[858])|((m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1555])|(m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1555])|(~m[1523]&m[1524]&m[1525]&~m[1526]&~m[1555])|(m[1523]&m[1524]&m[1525]&~m[1526]&~m[1555])|(m[1523]&m[1524]&m[1525]&m[1526]&~m[1555])|(m[1523]&m[1524]&~m[1525]&~m[1526]&m[1555])|(m[1523]&~m[1524]&m[1525]&~m[1526]&m[1555])|(~m[1523]&m[1524]&m[1525]&~m[1526]&m[1555])|(m[1523]&m[1524]&m[1525]&~m[1526]&m[1555])|(m[1523]&m[1524]&m[1525]&m[1526]&m[1555]))):InitCond[1574];
    m[1532] = run?((((m[1528]&~m[1529]&~m[1530]&~m[1531]&~m[1560])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1560])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1560])|(m[1528]&m[1529]&~m[1530]&m[1531]&~m[1560])|(m[1528]&~m[1529]&m[1530]&m[1531]&~m[1560])|(~m[1528]&m[1529]&m[1530]&m[1531]&~m[1560]))&BiasedRNG[859])|(((m[1528]&~m[1529]&~m[1530]&~m[1531]&m[1560])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&m[1560])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&m[1560])|(m[1528]&m[1529]&~m[1530]&m[1531]&m[1560])|(m[1528]&~m[1529]&m[1530]&m[1531]&m[1560])|(~m[1528]&m[1529]&m[1530]&m[1531]&m[1560]))&~BiasedRNG[859])|((m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1560])|(m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1560])|(~m[1528]&m[1529]&m[1530]&~m[1531]&~m[1560])|(m[1528]&m[1529]&m[1530]&~m[1531]&~m[1560])|(m[1528]&m[1529]&m[1530]&m[1531]&~m[1560])|(m[1528]&m[1529]&~m[1530]&~m[1531]&m[1560])|(m[1528]&~m[1529]&m[1530]&~m[1531]&m[1560])|(~m[1528]&m[1529]&m[1530]&~m[1531]&m[1560])|(m[1528]&m[1529]&m[1530]&~m[1531]&m[1560])|(m[1528]&m[1529]&m[1530]&m[1531]&m[1560]))):InitCond[1575];
    m[1537] = run?((((m[1533]&~m[1534]&~m[1535]&~m[1536]&~m[1563])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1563])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1563])|(m[1533]&m[1534]&~m[1535]&m[1536]&~m[1563])|(m[1533]&~m[1534]&m[1535]&m[1536]&~m[1563])|(~m[1533]&m[1534]&m[1535]&m[1536]&~m[1563]))&BiasedRNG[860])|(((m[1533]&~m[1534]&~m[1535]&~m[1536]&m[1563])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&m[1563])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&m[1563])|(m[1533]&m[1534]&~m[1535]&m[1536]&m[1563])|(m[1533]&~m[1534]&m[1535]&m[1536]&m[1563])|(~m[1533]&m[1534]&m[1535]&m[1536]&m[1563]))&~BiasedRNG[860])|((m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1563])|(m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1563])|(~m[1533]&m[1534]&m[1535]&~m[1536]&~m[1563])|(m[1533]&m[1534]&m[1535]&~m[1536]&~m[1563])|(m[1533]&m[1534]&m[1535]&m[1536]&~m[1563])|(m[1533]&m[1534]&~m[1535]&~m[1536]&m[1563])|(m[1533]&~m[1534]&m[1535]&~m[1536]&m[1563])|(~m[1533]&m[1534]&m[1535]&~m[1536]&m[1563])|(m[1533]&m[1534]&m[1535]&~m[1536]&m[1563])|(m[1533]&m[1534]&m[1535]&m[1536]&m[1563]))):InitCond[1576];
    m[1542] = run?((((m[1538]&~m[1539]&~m[1540]&~m[1541]&~m[1565])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1565])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1565])|(m[1538]&m[1539]&~m[1540]&m[1541]&~m[1565])|(m[1538]&~m[1539]&m[1540]&m[1541]&~m[1565])|(~m[1538]&m[1539]&m[1540]&m[1541]&~m[1565]))&BiasedRNG[861])|(((m[1538]&~m[1539]&~m[1540]&~m[1541]&m[1565])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&m[1565])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&m[1565])|(m[1538]&m[1539]&~m[1540]&m[1541]&m[1565])|(m[1538]&~m[1539]&m[1540]&m[1541]&m[1565])|(~m[1538]&m[1539]&m[1540]&m[1541]&m[1565]))&~BiasedRNG[861])|((m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1565])|(m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1565])|(~m[1538]&m[1539]&m[1540]&~m[1541]&~m[1565])|(m[1538]&m[1539]&m[1540]&~m[1541]&~m[1565])|(m[1538]&m[1539]&m[1540]&m[1541]&~m[1565])|(m[1538]&m[1539]&~m[1540]&~m[1541]&m[1565])|(m[1538]&~m[1539]&m[1540]&~m[1541]&m[1565])|(~m[1538]&m[1539]&m[1540]&~m[1541]&m[1565])|(m[1538]&m[1539]&m[1540]&~m[1541]&m[1565])|(m[1538]&m[1539]&m[1540]&m[1541]&m[1565]))):InitCond[1577];
    m[1547] = run?((((m[1543]&~m[1544]&~m[1545]&~m[1546]&~m[1570])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1570])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1570])|(m[1543]&m[1544]&~m[1545]&m[1546]&~m[1570])|(m[1543]&~m[1544]&m[1545]&m[1546]&~m[1570])|(~m[1543]&m[1544]&m[1545]&m[1546]&~m[1570]))&BiasedRNG[862])|(((m[1543]&~m[1544]&~m[1545]&~m[1546]&m[1570])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&m[1570])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&m[1570])|(m[1543]&m[1544]&~m[1545]&m[1546]&m[1570])|(m[1543]&~m[1544]&m[1545]&m[1546]&m[1570])|(~m[1543]&m[1544]&m[1545]&m[1546]&m[1570]))&~BiasedRNG[862])|((m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1570])|(m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1570])|(~m[1543]&m[1544]&m[1545]&~m[1546]&~m[1570])|(m[1543]&m[1544]&m[1545]&~m[1546]&~m[1570])|(m[1543]&m[1544]&m[1545]&m[1546]&~m[1570])|(m[1543]&m[1544]&~m[1545]&~m[1546]&m[1570])|(m[1543]&~m[1544]&m[1545]&~m[1546]&m[1570])|(~m[1543]&m[1544]&m[1545]&~m[1546]&m[1570])|(m[1543]&m[1544]&m[1545]&~m[1546]&m[1570])|(m[1543]&m[1544]&m[1545]&m[1546]&m[1570]))):InitCond[1578];
    m[1552] = run?((((m[1548]&~m[1549]&~m[1550]&~m[1551]&~m[1575])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1575])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1575])|(m[1548]&m[1549]&~m[1550]&m[1551]&~m[1575])|(m[1548]&~m[1549]&m[1550]&m[1551]&~m[1575])|(~m[1548]&m[1549]&m[1550]&m[1551]&~m[1575]))&BiasedRNG[863])|(((m[1548]&~m[1549]&~m[1550]&~m[1551]&m[1575])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&m[1575])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&m[1575])|(m[1548]&m[1549]&~m[1550]&m[1551]&m[1575])|(m[1548]&~m[1549]&m[1550]&m[1551]&m[1575])|(~m[1548]&m[1549]&m[1550]&m[1551]&m[1575]))&~BiasedRNG[863])|((m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1575])|(m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1575])|(~m[1548]&m[1549]&m[1550]&~m[1551]&~m[1575])|(m[1548]&m[1549]&m[1550]&~m[1551]&~m[1575])|(m[1548]&m[1549]&m[1550]&m[1551]&~m[1575])|(m[1548]&m[1549]&~m[1550]&~m[1551]&m[1575])|(m[1548]&~m[1549]&m[1550]&~m[1551]&m[1575])|(~m[1548]&m[1549]&m[1550]&~m[1551]&m[1575])|(m[1548]&m[1549]&m[1550]&~m[1551]&m[1575])|(m[1548]&m[1549]&m[1550]&m[1551]&m[1575]))):InitCond[1579];
    m[1557] = run?((((m[1553]&~m[1554]&~m[1555]&~m[1556]&~m[1580])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1580])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1580])|(m[1553]&m[1554]&~m[1555]&m[1556]&~m[1580])|(m[1553]&~m[1554]&m[1555]&m[1556]&~m[1580])|(~m[1553]&m[1554]&m[1555]&m[1556]&~m[1580]))&BiasedRNG[864])|(((m[1553]&~m[1554]&~m[1555]&~m[1556]&m[1580])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&m[1580])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&m[1580])|(m[1553]&m[1554]&~m[1555]&m[1556]&m[1580])|(m[1553]&~m[1554]&m[1555]&m[1556]&m[1580])|(~m[1553]&m[1554]&m[1555]&m[1556]&m[1580]))&~BiasedRNG[864])|((m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1580])|(m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1580])|(~m[1553]&m[1554]&m[1555]&~m[1556]&~m[1580])|(m[1553]&m[1554]&m[1555]&~m[1556]&~m[1580])|(m[1553]&m[1554]&m[1555]&m[1556]&~m[1580])|(m[1553]&m[1554]&~m[1555]&~m[1556]&m[1580])|(m[1553]&~m[1554]&m[1555]&~m[1556]&m[1580])|(~m[1553]&m[1554]&m[1555]&~m[1556]&m[1580])|(m[1553]&m[1554]&m[1555]&~m[1556]&m[1580])|(m[1553]&m[1554]&m[1555]&m[1556]&m[1580]))):InitCond[1580];
    m[1562] = run?((((m[1558]&~m[1559]&~m[1560]&~m[1561]&~m[1585])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1585])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1585])|(m[1558]&m[1559]&~m[1560]&m[1561]&~m[1585])|(m[1558]&~m[1559]&m[1560]&m[1561]&~m[1585])|(~m[1558]&m[1559]&m[1560]&m[1561]&~m[1585]))&BiasedRNG[865])|(((m[1558]&~m[1559]&~m[1560]&~m[1561]&m[1585])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&m[1585])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&m[1585])|(m[1558]&m[1559]&~m[1560]&m[1561]&m[1585])|(m[1558]&~m[1559]&m[1560]&m[1561]&m[1585])|(~m[1558]&m[1559]&m[1560]&m[1561]&m[1585]))&~BiasedRNG[865])|((m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1585])|(m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1585])|(~m[1558]&m[1559]&m[1560]&~m[1561]&~m[1585])|(m[1558]&m[1559]&m[1560]&~m[1561]&~m[1585])|(m[1558]&m[1559]&m[1560]&m[1561]&~m[1585])|(m[1558]&m[1559]&~m[1560]&~m[1561]&m[1585])|(m[1558]&~m[1559]&m[1560]&~m[1561]&m[1585])|(~m[1558]&m[1559]&m[1560]&~m[1561]&m[1585])|(m[1558]&m[1559]&m[1560]&~m[1561]&m[1585])|(m[1558]&m[1559]&m[1560]&m[1561]&m[1585]))):InitCond[1581];
    m[1567] = run?((((m[1563]&~m[1564]&~m[1565]&~m[1566]&~m[1588])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1588])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1588])|(m[1563]&m[1564]&~m[1565]&m[1566]&~m[1588])|(m[1563]&~m[1564]&m[1565]&m[1566]&~m[1588])|(~m[1563]&m[1564]&m[1565]&m[1566]&~m[1588]))&BiasedRNG[866])|(((m[1563]&~m[1564]&~m[1565]&~m[1566]&m[1588])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&m[1588])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&m[1588])|(m[1563]&m[1564]&~m[1565]&m[1566]&m[1588])|(m[1563]&~m[1564]&m[1565]&m[1566]&m[1588])|(~m[1563]&m[1564]&m[1565]&m[1566]&m[1588]))&~BiasedRNG[866])|((m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1588])|(m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1588])|(~m[1563]&m[1564]&m[1565]&~m[1566]&~m[1588])|(m[1563]&m[1564]&m[1565]&~m[1566]&~m[1588])|(m[1563]&m[1564]&m[1565]&m[1566]&~m[1588])|(m[1563]&m[1564]&~m[1565]&~m[1566]&m[1588])|(m[1563]&~m[1564]&m[1565]&~m[1566]&m[1588])|(~m[1563]&m[1564]&m[1565]&~m[1566]&m[1588])|(m[1563]&m[1564]&m[1565]&~m[1566]&m[1588])|(m[1563]&m[1564]&m[1565]&m[1566]&m[1588]))):InitCond[1582];
    m[1572] = run?((((m[1568]&~m[1569]&~m[1570]&~m[1571]&~m[1590])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1590])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1590])|(m[1568]&m[1569]&~m[1570]&m[1571]&~m[1590])|(m[1568]&~m[1569]&m[1570]&m[1571]&~m[1590])|(~m[1568]&m[1569]&m[1570]&m[1571]&~m[1590]))&BiasedRNG[867])|(((m[1568]&~m[1569]&~m[1570]&~m[1571]&m[1590])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&m[1590])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&m[1590])|(m[1568]&m[1569]&~m[1570]&m[1571]&m[1590])|(m[1568]&~m[1569]&m[1570]&m[1571]&m[1590])|(~m[1568]&m[1569]&m[1570]&m[1571]&m[1590]))&~BiasedRNG[867])|((m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1590])|(m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1590])|(~m[1568]&m[1569]&m[1570]&~m[1571]&~m[1590])|(m[1568]&m[1569]&m[1570]&~m[1571]&~m[1590])|(m[1568]&m[1569]&m[1570]&m[1571]&~m[1590])|(m[1568]&m[1569]&~m[1570]&~m[1571]&m[1590])|(m[1568]&~m[1569]&m[1570]&~m[1571]&m[1590])|(~m[1568]&m[1569]&m[1570]&~m[1571]&m[1590])|(m[1568]&m[1569]&m[1570]&~m[1571]&m[1590])|(m[1568]&m[1569]&m[1570]&m[1571]&m[1590]))):InitCond[1583];
    m[1577] = run?((((m[1573]&~m[1574]&~m[1575]&~m[1576]&~m[1595])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1595])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1595])|(m[1573]&m[1574]&~m[1575]&m[1576]&~m[1595])|(m[1573]&~m[1574]&m[1575]&m[1576]&~m[1595])|(~m[1573]&m[1574]&m[1575]&m[1576]&~m[1595]))&BiasedRNG[868])|(((m[1573]&~m[1574]&~m[1575]&~m[1576]&m[1595])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&m[1595])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&m[1595])|(m[1573]&m[1574]&~m[1575]&m[1576]&m[1595])|(m[1573]&~m[1574]&m[1575]&m[1576]&m[1595])|(~m[1573]&m[1574]&m[1575]&m[1576]&m[1595]))&~BiasedRNG[868])|((m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1595])|(m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1595])|(~m[1573]&m[1574]&m[1575]&~m[1576]&~m[1595])|(m[1573]&m[1574]&m[1575]&~m[1576]&~m[1595])|(m[1573]&m[1574]&m[1575]&m[1576]&~m[1595])|(m[1573]&m[1574]&~m[1575]&~m[1576]&m[1595])|(m[1573]&~m[1574]&m[1575]&~m[1576]&m[1595])|(~m[1573]&m[1574]&m[1575]&~m[1576]&m[1595])|(m[1573]&m[1574]&m[1575]&~m[1576]&m[1595])|(m[1573]&m[1574]&m[1575]&m[1576]&m[1595]))):InitCond[1584];
    m[1582] = run?((((m[1578]&~m[1579]&~m[1580]&~m[1581]&~m[1600])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1600])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1600])|(m[1578]&m[1579]&~m[1580]&m[1581]&~m[1600])|(m[1578]&~m[1579]&m[1580]&m[1581]&~m[1600])|(~m[1578]&m[1579]&m[1580]&m[1581]&~m[1600]))&BiasedRNG[869])|(((m[1578]&~m[1579]&~m[1580]&~m[1581]&m[1600])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&m[1600])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&m[1600])|(m[1578]&m[1579]&~m[1580]&m[1581]&m[1600])|(m[1578]&~m[1579]&m[1580]&m[1581]&m[1600])|(~m[1578]&m[1579]&m[1580]&m[1581]&m[1600]))&~BiasedRNG[869])|((m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1600])|(m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1600])|(~m[1578]&m[1579]&m[1580]&~m[1581]&~m[1600])|(m[1578]&m[1579]&m[1580]&~m[1581]&~m[1600])|(m[1578]&m[1579]&m[1580]&m[1581]&~m[1600])|(m[1578]&m[1579]&~m[1580]&~m[1581]&m[1600])|(m[1578]&~m[1579]&m[1580]&~m[1581]&m[1600])|(~m[1578]&m[1579]&m[1580]&~m[1581]&m[1600])|(m[1578]&m[1579]&m[1580]&~m[1581]&m[1600])|(m[1578]&m[1579]&m[1580]&m[1581]&m[1600]))):InitCond[1585];
    m[1587] = run?((((m[1583]&~m[1584]&~m[1585]&~m[1586]&~m[1605])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1605])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1605])|(m[1583]&m[1584]&~m[1585]&m[1586]&~m[1605])|(m[1583]&~m[1584]&m[1585]&m[1586]&~m[1605])|(~m[1583]&m[1584]&m[1585]&m[1586]&~m[1605]))&BiasedRNG[870])|(((m[1583]&~m[1584]&~m[1585]&~m[1586]&m[1605])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&m[1605])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&m[1605])|(m[1583]&m[1584]&~m[1585]&m[1586]&m[1605])|(m[1583]&~m[1584]&m[1585]&m[1586]&m[1605])|(~m[1583]&m[1584]&m[1585]&m[1586]&m[1605]))&~BiasedRNG[870])|((m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1605])|(m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1605])|(~m[1583]&m[1584]&m[1585]&~m[1586]&~m[1605])|(m[1583]&m[1584]&m[1585]&~m[1586]&~m[1605])|(m[1583]&m[1584]&m[1585]&m[1586]&~m[1605])|(m[1583]&m[1584]&~m[1585]&~m[1586]&m[1605])|(m[1583]&~m[1584]&m[1585]&~m[1586]&m[1605])|(~m[1583]&m[1584]&m[1585]&~m[1586]&m[1605])|(m[1583]&m[1584]&m[1585]&~m[1586]&m[1605])|(m[1583]&m[1584]&m[1585]&m[1586]&m[1605]))):InitCond[1586];
    m[1592] = run?((((m[1588]&~m[1589]&~m[1590]&~m[1591]&~m[1608])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1608])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1608])|(m[1588]&m[1589]&~m[1590]&m[1591]&~m[1608])|(m[1588]&~m[1589]&m[1590]&m[1591]&~m[1608])|(~m[1588]&m[1589]&m[1590]&m[1591]&~m[1608]))&BiasedRNG[871])|(((m[1588]&~m[1589]&~m[1590]&~m[1591]&m[1608])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&m[1608])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&m[1608])|(m[1588]&m[1589]&~m[1590]&m[1591]&m[1608])|(m[1588]&~m[1589]&m[1590]&m[1591]&m[1608])|(~m[1588]&m[1589]&m[1590]&m[1591]&m[1608]))&~BiasedRNG[871])|((m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1608])|(m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1608])|(~m[1588]&m[1589]&m[1590]&~m[1591]&~m[1608])|(m[1588]&m[1589]&m[1590]&~m[1591]&~m[1608])|(m[1588]&m[1589]&m[1590]&m[1591]&~m[1608])|(m[1588]&m[1589]&~m[1590]&~m[1591]&m[1608])|(m[1588]&~m[1589]&m[1590]&~m[1591]&m[1608])|(~m[1588]&m[1589]&m[1590]&~m[1591]&m[1608])|(m[1588]&m[1589]&m[1590]&~m[1591]&m[1608])|(m[1588]&m[1589]&m[1590]&m[1591]&m[1608]))):InitCond[1587];
    m[1597] = run?((((m[1593]&~m[1594]&~m[1595]&~m[1596]&~m[1610])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1610])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1610])|(m[1593]&m[1594]&~m[1595]&m[1596]&~m[1610])|(m[1593]&~m[1594]&m[1595]&m[1596]&~m[1610])|(~m[1593]&m[1594]&m[1595]&m[1596]&~m[1610]))&BiasedRNG[872])|(((m[1593]&~m[1594]&~m[1595]&~m[1596]&m[1610])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&m[1610])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&m[1610])|(m[1593]&m[1594]&~m[1595]&m[1596]&m[1610])|(m[1593]&~m[1594]&m[1595]&m[1596]&m[1610])|(~m[1593]&m[1594]&m[1595]&m[1596]&m[1610]))&~BiasedRNG[872])|((m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1610])|(m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1610])|(~m[1593]&m[1594]&m[1595]&~m[1596]&~m[1610])|(m[1593]&m[1594]&m[1595]&~m[1596]&~m[1610])|(m[1593]&m[1594]&m[1595]&m[1596]&~m[1610])|(m[1593]&m[1594]&~m[1595]&~m[1596]&m[1610])|(m[1593]&~m[1594]&m[1595]&~m[1596]&m[1610])|(~m[1593]&m[1594]&m[1595]&~m[1596]&m[1610])|(m[1593]&m[1594]&m[1595]&~m[1596]&m[1610])|(m[1593]&m[1594]&m[1595]&m[1596]&m[1610]))):InitCond[1588];
    m[1602] = run?((((m[1598]&~m[1599]&~m[1600]&~m[1601]&~m[1615])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1615])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1615])|(m[1598]&m[1599]&~m[1600]&m[1601]&~m[1615])|(m[1598]&~m[1599]&m[1600]&m[1601]&~m[1615])|(~m[1598]&m[1599]&m[1600]&m[1601]&~m[1615]))&BiasedRNG[873])|(((m[1598]&~m[1599]&~m[1600]&~m[1601]&m[1615])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&m[1615])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&m[1615])|(m[1598]&m[1599]&~m[1600]&m[1601]&m[1615])|(m[1598]&~m[1599]&m[1600]&m[1601]&m[1615])|(~m[1598]&m[1599]&m[1600]&m[1601]&m[1615]))&~BiasedRNG[873])|((m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1615])|(m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1615])|(~m[1598]&m[1599]&m[1600]&~m[1601]&~m[1615])|(m[1598]&m[1599]&m[1600]&~m[1601]&~m[1615])|(m[1598]&m[1599]&m[1600]&m[1601]&~m[1615])|(m[1598]&m[1599]&~m[1600]&~m[1601]&m[1615])|(m[1598]&~m[1599]&m[1600]&~m[1601]&m[1615])|(~m[1598]&m[1599]&m[1600]&~m[1601]&m[1615])|(m[1598]&m[1599]&m[1600]&~m[1601]&m[1615])|(m[1598]&m[1599]&m[1600]&m[1601]&m[1615]))):InitCond[1589];
    m[1607] = run?((((m[1603]&~m[1604]&~m[1605]&~m[1606]&~m[1620])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1620])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1620])|(m[1603]&m[1604]&~m[1605]&m[1606]&~m[1620])|(m[1603]&~m[1604]&m[1605]&m[1606]&~m[1620])|(~m[1603]&m[1604]&m[1605]&m[1606]&~m[1620]))&BiasedRNG[874])|(((m[1603]&~m[1604]&~m[1605]&~m[1606]&m[1620])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&m[1620])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&m[1620])|(m[1603]&m[1604]&~m[1605]&m[1606]&m[1620])|(m[1603]&~m[1604]&m[1605]&m[1606]&m[1620])|(~m[1603]&m[1604]&m[1605]&m[1606]&m[1620]))&~BiasedRNG[874])|((m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1620])|(m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1620])|(~m[1603]&m[1604]&m[1605]&~m[1606]&~m[1620])|(m[1603]&m[1604]&m[1605]&~m[1606]&~m[1620])|(m[1603]&m[1604]&m[1605]&m[1606]&~m[1620])|(m[1603]&m[1604]&~m[1605]&~m[1606]&m[1620])|(m[1603]&~m[1604]&m[1605]&~m[1606]&m[1620])|(~m[1603]&m[1604]&m[1605]&~m[1606]&m[1620])|(m[1603]&m[1604]&m[1605]&~m[1606]&m[1620])|(m[1603]&m[1604]&m[1605]&m[1606]&m[1620]))):InitCond[1590];
    m[1612] = run?((((m[1608]&~m[1609]&~m[1610]&~m[1611]&~m[1623])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1623])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1623])|(m[1608]&m[1609]&~m[1610]&m[1611]&~m[1623])|(m[1608]&~m[1609]&m[1610]&m[1611]&~m[1623])|(~m[1608]&m[1609]&m[1610]&m[1611]&~m[1623]))&BiasedRNG[875])|(((m[1608]&~m[1609]&~m[1610]&~m[1611]&m[1623])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&m[1623])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&m[1623])|(m[1608]&m[1609]&~m[1610]&m[1611]&m[1623])|(m[1608]&~m[1609]&m[1610]&m[1611]&m[1623])|(~m[1608]&m[1609]&m[1610]&m[1611]&m[1623]))&~BiasedRNG[875])|((m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1623])|(m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1623])|(~m[1608]&m[1609]&m[1610]&~m[1611]&~m[1623])|(m[1608]&m[1609]&m[1610]&~m[1611]&~m[1623])|(m[1608]&m[1609]&m[1610]&m[1611]&~m[1623])|(m[1608]&m[1609]&~m[1610]&~m[1611]&m[1623])|(m[1608]&~m[1609]&m[1610]&~m[1611]&m[1623])|(~m[1608]&m[1609]&m[1610]&~m[1611]&m[1623])|(m[1608]&m[1609]&m[1610]&~m[1611]&m[1623])|(m[1608]&m[1609]&m[1610]&m[1611]&m[1623]))):InitCond[1591];
    m[1617] = run?((((m[1613]&~m[1614]&~m[1615]&~m[1616]&~m[1625])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1625])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1625])|(m[1613]&m[1614]&~m[1615]&m[1616]&~m[1625])|(m[1613]&~m[1614]&m[1615]&m[1616]&~m[1625])|(~m[1613]&m[1614]&m[1615]&m[1616]&~m[1625]))&BiasedRNG[876])|(((m[1613]&~m[1614]&~m[1615]&~m[1616]&m[1625])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&m[1625])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&m[1625])|(m[1613]&m[1614]&~m[1615]&m[1616]&m[1625])|(m[1613]&~m[1614]&m[1615]&m[1616]&m[1625])|(~m[1613]&m[1614]&m[1615]&m[1616]&m[1625]))&~BiasedRNG[876])|((m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1625])|(m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1625])|(~m[1613]&m[1614]&m[1615]&~m[1616]&~m[1625])|(m[1613]&m[1614]&m[1615]&~m[1616]&~m[1625])|(m[1613]&m[1614]&m[1615]&m[1616]&~m[1625])|(m[1613]&m[1614]&~m[1615]&~m[1616]&m[1625])|(m[1613]&~m[1614]&m[1615]&~m[1616]&m[1625])|(~m[1613]&m[1614]&m[1615]&~m[1616]&m[1625])|(m[1613]&m[1614]&m[1615]&~m[1616]&m[1625])|(m[1613]&m[1614]&m[1615]&m[1616]&m[1625]))):InitCond[1592];
    m[1622] = run?((((m[1618]&~m[1619]&~m[1620]&~m[1621]&~m[1630])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1630])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1630])|(m[1618]&m[1619]&~m[1620]&m[1621]&~m[1630])|(m[1618]&~m[1619]&m[1620]&m[1621]&~m[1630])|(~m[1618]&m[1619]&m[1620]&m[1621]&~m[1630]))&BiasedRNG[877])|(((m[1618]&~m[1619]&~m[1620]&~m[1621]&m[1630])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&m[1630])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&m[1630])|(m[1618]&m[1619]&~m[1620]&m[1621]&m[1630])|(m[1618]&~m[1619]&m[1620]&m[1621]&m[1630])|(~m[1618]&m[1619]&m[1620]&m[1621]&m[1630]))&~BiasedRNG[877])|((m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1630])|(m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1630])|(~m[1618]&m[1619]&m[1620]&~m[1621]&~m[1630])|(m[1618]&m[1619]&m[1620]&~m[1621]&~m[1630])|(m[1618]&m[1619]&m[1620]&m[1621]&~m[1630])|(m[1618]&m[1619]&~m[1620]&~m[1621]&m[1630])|(m[1618]&~m[1619]&m[1620]&~m[1621]&m[1630])|(~m[1618]&m[1619]&m[1620]&~m[1621]&m[1630])|(m[1618]&m[1619]&m[1620]&~m[1621]&m[1630])|(m[1618]&m[1619]&m[1620]&m[1621]&m[1630]))):InitCond[1593];
    m[1627] = run?((((m[1623]&~m[1624]&~m[1625]&~m[1626]&~m[1633])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1633])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1633])|(m[1623]&m[1624]&~m[1625]&m[1626]&~m[1633])|(m[1623]&~m[1624]&m[1625]&m[1626]&~m[1633])|(~m[1623]&m[1624]&m[1625]&m[1626]&~m[1633]))&BiasedRNG[878])|(((m[1623]&~m[1624]&~m[1625]&~m[1626]&m[1633])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&m[1633])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&m[1633])|(m[1623]&m[1624]&~m[1625]&m[1626]&m[1633])|(m[1623]&~m[1624]&m[1625]&m[1626]&m[1633])|(~m[1623]&m[1624]&m[1625]&m[1626]&m[1633]))&~BiasedRNG[878])|((m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1633])|(m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1633])|(~m[1623]&m[1624]&m[1625]&~m[1626]&~m[1633])|(m[1623]&m[1624]&m[1625]&~m[1626]&~m[1633])|(m[1623]&m[1624]&m[1625]&m[1626]&~m[1633])|(m[1623]&m[1624]&~m[1625]&~m[1626]&m[1633])|(m[1623]&~m[1624]&m[1625]&~m[1626]&m[1633])|(~m[1623]&m[1624]&m[1625]&~m[1626]&m[1633])|(m[1623]&m[1624]&m[1625]&~m[1626]&m[1633])|(m[1623]&m[1624]&m[1625]&m[1626]&m[1633]))):InitCond[1594];
    m[1632] = run?((((m[1628]&~m[1629]&~m[1630]&~m[1631]&~m[1635])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1635])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1635])|(m[1628]&m[1629]&~m[1630]&m[1631]&~m[1635])|(m[1628]&~m[1629]&m[1630]&m[1631]&~m[1635])|(~m[1628]&m[1629]&m[1630]&m[1631]&~m[1635]))&BiasedRNG[879])|(((m[1628]&~m[1629]&~m[1630]&~m[1631]&m[1635])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&m[1635])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&m[1635])|(m[1628]&m[1629]&~m[1630]&m[1631]&m[1635])|(m[1628]&~m[1629]&m[1630]&m[1631]&m[1635])|(~m[1628]&m[1629]&m[1630]&m[1631]&m[1635]))&~BiasedRNG[879])|((m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1635])|(m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1635])|(~m[1628]&m[1629]&m[1630]&~m[1631]&~m[1635])|(m[1628]&m[1629]&m[1630]&~m[1631]&~m[1635])|(m[1628]&m[1629]&m[1630]&m[1631]&~m[1635])|(m[1628]&m[1629]&~m[1630]&~m[1631]&m[1635])|(m[1628]&~m[1629]&m[1630]&~m[1631]&m[1635])|(~m[1628]&m[1629]&m[1630]&~m[1631]&m[1635])|(m[1628]&m[1629]&m[1630]&~m[1631]&m[1635])|(m[1628]&m[1629]&m[1630]&m[1631]&m[1635]))):InitCond[1595];
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[372]&LFSRcolor0[13]&LFSRcolor0[170]);
    BiasedRNG[1] = (LFSRcolor0[550]&LFSRcolor0[182]&LFSRcolor0[367]);
    BiasedRNG[2] = (LFSRcolor0[52]&LFSRcolor0[30]&LFSRcolor0[570]);
    BiasedRNG[3] = (LFSRcolor0[621]&LFSRcolor0[807]&LFSRcolor0[181]);
    BiasedRNG[4] = (LFSRcolor0[836]&LFSRcolor0[652]&LFSRcolor0[571]);
    BiasedRNG[5] = (LFSRcolor0[881]&LFSRcolor0[513]&LFSRcolor0[515]);
    BiasedRNG[6] = (LFSRcolor0[943]&LFSRcolor0[289]&LFSRcolor0[284]);
    BiasedRNG[7] = (LFSRcolor0[299]&LFSRcolor0[551]&LFSRcolor0[555]);
    BiasedRNG[8] = (LFSRcolor0[199]&LFSRcolor0[257]&LFSRcolor0[882]);
    BiasedRNG[9] = (LFSRcolor0[940]&LFSRcolor0[748]&LFSRcolor0[417]);
    BiasedRNG[10] = (LFSRcolor0[378]&LFSRcolor0[957]&LFSRcolor0[922]);
    BiasedRNG[11] = (LFSRcolor0[60]&LFSRcolor0[485]&LFSRcolor0[581]);
    BiasedRNG[12] = (LFSRcolor0[118]&LFSRcolor0[675]&LFSRcolor0[519]);
    BiasedRNG[13] = (LFSRcolor0[270]&LFSRcolor0[802]&LFSRcolor0[632]);
    BiasedRNG[14] = (LFSRcolor0[308]&LFSRcolor0[885]&LFSRcolor0[587]);
    BiasedRNG[15] = (LFSRcolor0[639]&LFSRcolor0[189]&LFSRcolor0[577]);
    BiasedRNG[16] = (LFSRcolor0[559]&LFSRcolor0[563]&LFSRcolor0[791]);
    BiasedRNG[17] = (LFSRcolor0[301]&LFSRcolor0[100]&LFSRcolor0[116]);
    BiasedRNG[18] = (LFSRcolor0[1]&LFSRcolor0[668]&LFSRcolor0[593]);
    BiasedRNG[19] = (LFSRcolor0[685]&LFSRcolor0[520]&LFSRcolor0[67]);
    BiasedRNG[20] = (LFSRcolor0[202]&LFSRcolor0[124]&LFSRcolor0[127]);
    BiasedRNG[21] = (LFSRcolor0[919]&LFSRcolor0[723]&LFSRcolor0[37]);
    BiasedRNG[22] = (LFSRcolor0[19]&LFSRcolor0[841]&LFSRcolor0[963]);
    BiasedRNG[23] = (LFSRcolor0[868]&LFSRcolor0[512]&LFSRcolor0[365]);
    BiasedRNG[24] = (LFSRcolor0[869]&LFSRcolor0[822]&LFSRcolor0[6]);
    BiasedRNG[25] = (LFSRcolor0[696]&LFSRcolor0[751]&LFSRcolor0[197]);
    BiasedRNG[26] = (LFSRcolor0[656]&LFSRcolor0[695]&LFSRcolor0[400]);
    BiasedRNG[27] = (LFSRcolor0[106]&LFSRcolor0[566]&LFSRcolor0[15]);
    BiasedRNG[28] = (LFSRcolor0[401]&LFSRcolor0[902]&LFSRcolor0[915]);
    BiasedRNG[29] = (LFSRcolor0[392]&LFSRcolor0[853]&LFSRcolor0[797]);
    BiasedRNG[30] = (LFSRcolor0[851]&LFSRcolor0[917]&LFSRcolor0[153]);
    BiasedRNG[31] = (LFSRcolor0[762]&LFSRcolor0[521]&LFSRcolor0[645]);
    BiasedRNG[32] = (LFSRcolor0[716]&LFSRcolor0[612]&LFSRcolor0[833]);
    BiasedRNG[33] = (LFSRcolor0[418]&LFSRcolor0[55]&LFSRcolor0[745]);
    BiasedRNG[34] = (LFSRcolor0[901]&LFSRcolor0[364]&LFSRcolor0[561]);
    BiasedRNG[35] = (LFSRcolor0[862]&LFSRcolor0[474]&LFSRcolor0[429]);
    BiasedRNG[36] = (LFSRcolor0[912]&LFSRcolor0[863]&LFSRcolor0[595]);
    BiasedRNG[37] = (LFSRcolor0[768]&LFSRcolor0[375]&LFSRcolor0[380]);
    BiasedRNG[38] = (LFSRcolor0[923]&LFSRcolor0[196]&LFSRcolor0[205]);
    BiasedRNG[39] = (LFSRcolor0[133]&LFSRcolor0[921]&LFSRcolor0[247]);
    BiasedRNG[40] = (LFSRcolor0[201]&LFSRcolor0[91]&LFSRcolor0[450]);
    BiasedRNG[41] = (LFSRcolor0[204]&LFSRcolor0[221]&LFSRcolor0[918]);
    BiasedRNG[42] = (LFSRcolor0[88]&LFSRcolor0[283]&LFSRcolor0[362]);
    BiasedRNG[43] = (LFSRcolor0[459]&LFSRcolor0[423]&LFSRcolor0[140]);
    BiasedRNG[44] = (LFSRcolor0[461]&LFSRcolor0[298]&LFSRcolor0[729]);
    BiasedRNG[45] = (LFSRcolor0[897]&LFSRcolor0[416]&LFSRcolor0[71]);
    BiasedRNG[46] = (LFSRcolor0[800]&LFSRcolor0[737]&LFSRcolor0[906]);
    BiasedRNG[47] = (LFSRcolor0[277]&LFSRcolor0[691]&LFSRcolor0[161]);
    BiasedRNG[48] = (LFSRcolor0[425]&LFSRcolor0[354]&LFSRcolor0[61]);
    BiasedRNG[49] = (LFSRcolor0[180]&LFSRcolor0[49]&LFSRcolor0[143]);
    BiasedRNG[50] = (LFSRcolor0[821]&LFSRcolor0[647]&LFSRcolor0[340]);
    BiasedRNG[51] = (LFSRcolor0[329]&LFSRcolor0[847]&LFSRcolor0[216]);
    BiasedRNG[52] = (LFSRcolor0[498]&LFSRcolor0[774]&LFSRcolor0[145]);
    BiasedRNG[53] = (LFSRcolor0[648]&LFSRcolor0[245]&LFSRcolor0[516]);
    BiasedRNG[54] = (LFSRcolor0[872]&LFSRcolor0[763]&LFSRcolor0[112]);
    BiasedRNG[55] = (LFSRcolor0[237]&LFSRcolor0[813]&LFSRcolor0[235]);
    BiasedRNG[56] = (LFSRcolor0[252]&LFSRcolor0[939]&LFSRcolor0[321]);
    BiasedRNG[57] = (LFSRcolor0[74]&LFSRcolor0[345]&LFSRcolor0[928]);
    BiasedRNG[58] = (LFSRcolor0[481]&LFSRcolor0[892]&LFSRcolor0[908]);
    BiasedRNG[59] = (LFSRcolor0[435]&LFSRcolor0[231]&LFSRcolor0[782]);
    BiasedRNG[60] = (LFSRcolor0[441]&LFSRcolor0[219]&LFSRcolor0[315]);
    BiasedRNG[61] = (LFSRcolor0[524]&LFSRcolor0[402]&LFSRcolor0[738]);
    BiasedRNG[62] = (LFSRcolor0[809]&LFSRcolor0[295]&LFSRcolor0[488]);
    BiasedRNG[63] = (LFSRcolor0[925]&LFSRcolor0[630]&LFSRcolor0[360]);
    BiasedRNG[64] = (LFSRcolor0[383]&LFSRcolor0[73]&LFSRcolor0[828]);
    BiasedRNG[65] = (LFSRcolor0[350]&LFSRcolor0[523]&LFSRcolor0[569]);
    BiasedRNG[66] = (LFSRcolor0[709]&LFSRcolor0[280]&LFSRcolor0[290]);
    BiasedRNG[67] = (LFSRcolor0[195]&LFSRcolor0[602]&LFSRcolor0[394]);
    BiasedRNG[68] = (LFSRcolor0[522]&LFSRcolor0[547]&LFSRcolor0[431]);
    BiasedRNG[69] = (LFSRcolor0[164]&LFSRcolor0[733]&LFSRcolor0[784]);
    BiasedRNG[70] = (LFSRcolor0[878]&LFSRcolor0[677]&LFSRcolor0[776]);
    BiasedRNG[71] = (LFSRcolor0[369]&LFSRcolor0[646]&LFSRcolor0[880]);
    BiasedRNG[72] = (LFSRcolor0[568]&LFSRcolor0[533]&LFSRcolor0[110]);
    BiasedRNG[73] = (LFSRcolor0[671]&LFSRcolor0[309]&LFSRcolor0[410]);
    BiasedRNG[74] = (LFSRcolor0[597]&LFSRcolor0[444]&LFSRcolor0[198]);
    BiasedRNG[75] = (LFSRcolor0[338]&LFSRcolor0[495]&LFSRcolor0[333]);
    BiasedRNG[76] = (LFSRcolor0[149]&LFSRcolor0[82]&LFSRcolor0[653]);
    BiasedRNG[77] = (LFSRcolor0[777]&LFSRcolor0[109]&LFSRcolor0[104]);
    BiasedRNG[78] = (LFSRcolor0[306]&LFSRcolor0[689]&LFSRcolor0[871]);
    BiasedRNG[79] = (LFSRcolor0[59]&LFSRcolor0[148]&LFSRcolor0[508]);
    BiasedRNG[80] = (LFSRcolor0[398]&LFSRcolor0[891]&LFSRcolor0[108]);
    BiasedRNG[81] = (LFSRcolor0[669]&LFSRcolor0[141]&LFSRcolor0[185]);
    BiasedRNG[82] = (LFSRcolor0[883]&LFSRcolor0[837]&LFSRcolor0[773]);
    BiasedRNG[83] = (LFSRcolor0[25]&LFSRcolor0[764]&LFSRcolor0[334]);
    BiasedRNG[84] = (LFSRcolor0[889]&LFSRcolor0[496]&LFSRcolor0[85]);
    BiasedRNG[85] = (LFSRcolor0[759]&LFSRcolor0[83]&LFSRcolor0[941]);
    BiasedRNG[86] = (LFSRcolor0[905]&LFSRcolor0[128]&LFSRcolor0[749]);
    BiasedRNG[87] = (LFSRcolor0[663]&LFSRcolor0[86]&LFSRcolor0[62]);
    BiasedRNG[88] = (LFSRcolor0[212]&LFSRcolor0[31]&LFSRcolor0[420]);
    BiasedRNG[89] = (LFSRcolor0[436]&LFSRcolor0[553]&LFSRcolor0[795]);
    BiasedRNG[90] = (LFSRcolor0[35]&LFSRcolor0[379]&LFSRcolor0[105]);
    BiasedRNG[91] = (LFSRcolor0[576]&LFSRcolor0[278]&LFSRcolor0[497]);
    BiasedRNG[92] = (LFSRcolor0[714]&LFSRcolor0[552]&LFSRcolor0[599]);
    BiasedRNG[93] = (LFSRcolor0[491]&LFSRcolor0[772]&LFSRcolor0[303]);
    BiasedRNG[94] = (LFSRcolor0[603]&LFSRcolor0[403]&LFSRcolor0[363]);
    BiasedRNG[95] = (LFSRcolor0[704]&LFSRcolor0[582]&LFSRcolor0[598]);
    BiasedRNG[96] = (LFSRcolor0[279]&LFSRcolor0[692]&LFSRcolor0[705]);
    BiasedRNG[97] = (LFSRcolor0[610]&LFSRcolor0[910]&LFSRcolor0[535]);
    BiasedRNG[98] = (LFSRcolor0[664]&LFSRcolor0[830]&LFSRcolor0[744]);
    BiasedRNG[99] = (LFSRcolor0[625]&LFSRcolor0[433]&LFSRcolor0[766]);
    BiasedRNG[100] = (LFSRcolor0[788]&LFSRcolor0[586]&LFSRcolor0[954]);
    BiasedRNG[101] = (LFSRcolor0[534]&LFSRcolor0[328]&LFSRcolor0[893]);
    BiasedRNG[102] = (LFSRcolor0[34]&LFSRcolor0[193]&LFSRcolor0[938]);
    BiasedRNG[103] = (LFSRcolor0[792]&LFSRcolor0[574]&LFSRcolor0[734]);
    BiasedRNG[104] = (LFSRcolor0[820]&LFSRcolor0[405]&LFSRcolor0[810]);
    BiasedRNG[105] = (LFSRcolor0[57]&LFSRcolor0[210]&LFSRcolor0[335]);
    BiasedRNG[106] = (LFSRcolor0[5]&LFSRcolor0[838]&LFSRcolor0[952]);
    BiasedRNG[107] = (LFSRcolor0[679]&LFSRcolor0[448]&LFSRcolor0[786]);
    BiasedRNG[108] = (LFSRcolor0[251]&LFSRcolor0[846]&LFSRcolor0[752]);
    BiasedRNG[109] = (LFSRcolor0[23]&LFSRcolor0[457]&LFSRcolor0[961]);
    BiasedRNG[110] = (LFSRcolor0[53]&LFSRcolor0[68]&LFSRcolor0[680]);
    BiasedRNG[111] = (LFSRcolor0[913]&LFSRcolor0[440]&LFSRcolor0[850]);
    BiasedRNG[112] = (LFSRcolor0[747]&LFSRcolor0[655]&LFSRcolor0[658]);
    BiasedRNG[113] = (LFSRcolor0[113]&LFSRcolor0[617]&LFSRcolor0[408]);
    BiasedRNG[114] = (LFSRcolor0[578]&LFSRcolor0[200]&LFSRcolor0[89]);
    BiasedRNG[115] = (LFSRcolor0[152]&LFSRcolor0[702]&LFSRcolor0[717]);
    BiasedRNG[116] = (LFSRcolor0[536]&LFSRcolor0[812]&LFSRcolor0[638]);
    BiasedRNG[117] = (LFSRcolor0[565]&LFSRcolor0[793]&LFSRcolor0[213]);
    BiasedRNG[118] = (LFSRcolor0[359]&LFSRcolor0[866]&LFSRcolor0[864]);
    BiasedRNG[119] = (LFSRcolor0[860]&LFSRcolor0[890]&LFSRcolor0[471]);
    BiasedRNG[120] = (LFSRcolor0[226]&LFSRcolor0[827]&LFSRcolor0[722]);
    BiasedRNG[121] = (LFSRcolor0[310]&LFSRcolor0[946]&LFSRcolor0[510]);
    BiasedRNG[122] = (LFSRcolor0[190]&LFSRcolor0[628]&LFSRcolor0[421]);
    BiasedRNG[123] = (LFSRcolor0[909]&LFSRcolor0[583]&LFSRcolor0[843]);
    BiasedRNG[124] = (LFSRcolor0[783]&LFSRcolor0[7]&LFSRcolor0[622]);
    BiasedRNG[125] = (LFSRcolor0[160]&LFSRcolor0[166]&LFSRcolor0[899]);
    BiasedRNG[126] = (LFSRcolor0[234]&LFSRcolor0[564]&LFSRcolor0[958]);
    BiasedRNG[127] = (LFSRcolor0[944]&LFSRcolor0[93]&LFSRcolor0[607]);
    BiasedRNG[128] = (LFSRcolor0[227]&LFSRcolor0[805]&LFSRcolor0[824]);
    BiasedRNG[129] = (LFSRcolor0[4]&LFSRcolor0[456]&LFSRcolor0[81]);
    BiasedRNG[130] = (LFSRcolor0[490]&LFSRcolor0[546]&LFSRcolor0[765]);
    BiasedRNG[131] = (LFSRcolor0[514]&LFSRcolor0[343]&LFSRcolor0[604]);
    BiasedRNG[132] = (LFSRcolor0[511]&LFSRcolor0[275]&LFSRcolor0[609]);
    BiasedRNG[133] = (LFSRcolor0[469]&LFSRcolor0[718]&LFSRcolor0[888]);
    BiasedRNG[134] = (LFSRcolor0[554]&LFSRcolor0[665]&LFSRcolor0[895]);
    BiasedRNG[135] = (LFSRcolor0[253]&LFSRcolor0[320]&LFSRcolor0[114]);
    BiasedRNG[136] = (LFSRcolor0[518]&LFSRcolor0[951]&LFSRcolor0[102]);
    BiasedRNG[137] = (LFSRcolor0[179]&LFSRcolor0[690]&LFSRcolor0[248]);
    BiasedRNG[138] = (LFSRcolor0[817]&LFSRcolor0[590]&LFSRcolor0[312]);
    BiasedRNG[139] = (LFSRcolor0[56]&LFSRcolor0[344]&LFSRcolor0[556]);
    BiasedRNG[140] = (LFSRcolor0[374]&LFSRcolor0[428]&LFSRcolor0[949]);
    BiasedRNG[141] = (LFSRcolor0[386]&LFSRcolor0[567]&LFSRcolor0[264]);
    BiasedRNG[142] = (LFSRcolor0[845]&LFSRcolor0[483]&LFSRcolor0[588]);
    BiasedRNG[143] = (LFSRcolor0[20]&LFSRcolor0[287]&LFSRcolor0[477]);
    BiasedRNG[144] = (LFSRcolor0[69]&LFSRcolor0[760]&LFSRcolor0[135]);
    BiasedRNG[145] = (LFSRcolor0[727]&LFSRcolor0[541]&LFSRcolor0[94]);
    BiasedRNG[146] = (LFSRcolor0[162]&LFSRcolor0[318]&LFSRcolor0[686]);
    BiasedRNG[147] = (LFSRcolor0[472]&LFSRcolor0[507]&LFSRcolor0[530]);
    BiasedRNG[148] = (LFSRcolor0[904]&LFSRcolor0[780]&LFSRcolor0[107]);
    BiasedRNG[149] = (LFSRcolor0[389]&LFSRcolor0[214]&LFSRcolor0[808]);
    BiasedRNG[150] = (LFSRcolor0[14]&LFSRcolor0[463]&LFSRcolor0[156]);
    BiasedRNG[151] = (LFSRcolor0[644]&LFSRcolor0[549]&LFSRcolor0[740]);
    BiasedRNG[152] = (LFSRcolor0[76]&LFSRcolor0[684]&LFSRcolor0[194]);
    BiasedRNG[153] = (LFSRcolor0[623]&LFSRcolor0[47]&LFSRcolor0[711]);
    BiasedRNG[154] = (LFSRcolor0[385]&LFSRcolor0[529]&LFSRcolor0[325]);
    BiasedRNG[155] = (LFSRcolor0[70]&LFSRcolor0[84]&LFSRcolor0[771]);
    BiasedRNG[156] = (LFSRcolor0[580]&LFSRcolor0[482]&LFSRcolor0[464]);
    BiasedRNG[157] = (LFSRcolor0[624]&LFSRcolor0[606]&LFSRcolor0[256]);
    BiasedRNG[158] = (LFSRcolor0[388]&LFSRcolor0[393]&LFSRcolor0[540]);
    BiasedRNG[159] = (LFSRcolor0[42]&LFSRcolor0[122]&LFSRcolor0[942]);
    BiasedRNG[160] = (LFSRcolor0[215]&LFSRcolor0[538]&LFSRcolor0[132]);
    BiasedRNG[161] = (LFSRcolor0[649]&LFSRcolor0[137]&LFSRcolor0[302]);
    BiasedRNG[162] = (LFSRcolor0[176]&LFSRcolor0[503]&LFSRcolor0[144]);
    BiasedRNG[163] = (LFSRcolor0[694]&LFSRcolor0[470]&LFSRcolor0[693]);
    BiasedRNG[164] = (LFSRcolor0[356]&LFSRcolor0[673]&LFSRcolor0[300]);
    BiasedRNG[165] = (LFSRcolor0[304]&LFSRcolor0[351]&LFSRcolor0[858]);
    BiasedRNG[166] = (LFSRcolor0[948]&LFSRcolor0[442]&LFSRcolor0[29]);
    BiasedRNG[167] = (LFSRcolor0[806]&LFSRcolor0[798]&LFSRcolor0[594]);
    BiasedRNG[168] = (LFSRcolor0[614]&LFSRcolor0[676]&LFSRcolor0[449]);
    BiasedRNG[169] = (LFSRcolor0[90]&LFSRcolor0[111]&LFSRcolor0[8]);
    BiasedRNG[170] = (LFSRcolor0[674]&LFSRcolor0[840]&LFSRcolor0[382]);
    BiasedRNG[171] = (LFSRcolor0[377]&LFSRcolor0[120]&LFSRcolor0[842]);
    BiasedRNG[172] = (LFSRcolor0[557]&LFSRcolor0[58]&LFSRcolor0[672]);
    BiasedRNG[173] = (LFSRcolor0[80]&LFSRcolor0[51]&LFSRcolor0[907]);
    BiasedRNG[174] = (LFSRcolor0[217]&LFSRcolor0[454]&LFSRcolor0[266]);
    BiasedRNG[175] = (LFSRcolor0[79]&LFSRcolor0[713]&LFSRcolor0[123]);
    BiasedRNG[176] = (LFSRcolor0[670]&LFSRcolor0[430]&LFSRcolor0[870]);
    BiasedRNG[177] = (LFSRcolor0[155]&LFSRcolor0[361]&LFSRcolor0[710]);
    BiasedRNG[178] = (LFSRcolor0[504]&LFSRcolor0[206]&LFSRcolor0[475]);
    BiasedRNG[179] = (LFSRcolor0[285]&LFSRcolor0[426]&LFSRcolor0[924]);
    BiasedRNG[180] = (LFSRcolor0[236]&LFSRcolor0[131]&LFSRcolor0[172]);
    BiasedRNG[181] = (LFSRcolor0[78]&LFSRcolor0[801]&LFSRcolor0[125]);
    BiasedRNG[182] = (LFSRcolor0[165]&LFSRcolor0[916]&LFSRcolor0[397]);
    BiasedRNG[183] = (LFSRcolor0[758]&LFSRcolor0[92]&LFSRcolor0[434]);
    BiasedRNG[184] = (LFSRcolor0[856]&LFSRcolor0[778]&LFSRcolor0[307]);
    BiasedRNG[185] = (LFSRcolor0[825]&LFSRcolor0[151]&LFSRcolor0[158]);
    BiasedRNG[186] = (LFSRcolor0[332]&LFSRcolor0[451]&LFSRcolor0[532]);
    BiasedRNG[187] = (LFSRcolor0[558]&LFSRcolor0[965]&LFSRcolor0[683]);
    BiasedRNG[188] = (LFSRcolor0[712]&LFSRcolor0[101]&LFSRcolor0[815]);
    BiasedRNG[189] = (LFSRcolor0[687]&LFSRcolor0[500]&LFSRcolor0[666]);
    BiasedRNG[190] = (LFSRcolor0[579]&LFSRcolor0[2]&LFSRcolor0[715]);
    BiasedRNG[191] = (LFSRcolor0[501]&LFSRcolor0[947]&LFSRcolor0[272]);
    BiasedRNG[192] = (LFSRcolor0[467]&LFSRcolor0[187]&LFSRcolor0[753]);
    BiasedRNG[193] = (LFSRcolor0[208]&LFSRcolor0[616]&LFSRcolor0[831]);
    BiasedRNG[194] = (LFSRcolor0[844]&LFSRcolor0[281]&LFSRcolor0[494]);
    BiasedRNG[195] = (LFSRcolor0[404]&LFSRcolor0[409]&LFSRcolor0[146]);
    BiasedRNG[196] = (LFSRcolor0[834]&LFSRcolor0[415]&LFSRcolor0[169]);
    BiasedRNG[197] = (LFSRcolor0[0]&LFSRcolor0[316]&LFSRcolor0[626]);
    BiasedRNG[198] = (LFSRcolor0[543]&LFSRcolor0[119]&LFSRcolor0[867]);
    BiasedRNG[199] = (LFSRcolor0[211]&LFSRcolor0[407]&LFSRcolor0[32]);
    BiasedRNG[200] = (LFSRcolor0[238]&LFSRcolor0[874]&LFSRcolor0[667]);
    BiasedRNG[201] = (LFSRcolor0[258]&LFSRcolor0[537]&LFSRcolor0[373]);
    BiasedRNG[202] = (LFSRcolor0[886]&LFSRcolor0[260]&LFSRcolor0[241]);
    BiasedRNG[203] = (LFSRcolor0[634]&LFSRcolor0[896]&LFSRcolor0[964]);
    BiasedRNG[204] = (LFSRcolor0[54]&LFSRcolor0[803]&LFSRcolor0[139]);
    BiasedRNG[205] = (LFSRcolor0[349]&LFSRcolor0[453]&LFSRcolor0[641]);
    BiasedRNG[206] = (LFSRcolor0[313]&LFSRcolor0[28]&LFSRcolor0[134]);
    BiasedRNG[207] = (LFSRcolor0[473]&LFSRcolor0[887]&LFSRcolor0[631]);
    BiasedRNG[208] = (LFSRcolor0[900]&LFSRcolor0[750]&LFSRcolor0[953]);
    BiasedRNG[209] = (LFSRcolor0[240]&LFSRcolor0[412]&LFSRcolor0[384]);
    BiasedRNG[210] = (LFSRcolor0[615]&LFSRcolor0[422]&LFSRcolor0[159]);
    BiasedRNG[211] = (LFSRcolor0[959]&LFSRcolor0[255]&LFSRcolor0[572]);
    BiasedRNG[212] = (LFSRcolor0[36]&LFSRcolor0[296]&LFSRcolor0[274]);
    BiasedRNG[213] = (LFSRcolor0[589]&LFSRcolor0[794]&LFSRcolor0[562]);
    BiasedRNG[214] = (LFSRcolor0[835]&LFSRcolor0[873]&LFSRcolor0[613]);
    BiasedRNG[215] = (LFSRcolor0[732]&LFSRcolor0[642]&LFSRcolor0[305]);
    BiasedRNG[216] = (LFSRcolor0[232]&LFSRcolor0[445]&LFSRcolor0[218]);
    BiasedRNG[217] = (LFSRcolor0[936]&LFSRcolor0[357]&LFSRcolor0[643]);
    BiasedRNG[218] = (LFSRcolor0[884]&LFSRcolor0[12]&LFSRcolor0[592]);
    BiasedRNG[219] = (LFSRcolor0[950]&LFSRcolor0[17]&LFSRcolor0[781]);
    BiasedRNG[220] = (LFSRcolor0[743]&LFSRcolor0[353]&LFSRcolor0[955]);
    BiasedRNG[221] = (LFSRcolor0[291]&LFSRcolor0[811]&LFSRcolor0[339]);
    BiasedRNG[222] = (LFSRcolor0[761]&LFSRcolor0[292]&LFSRcolor0[697]);
    BiasedRNG[223] = (LFSRcolor0[854]&LFSRcolor0[848]&LFSRcolor0[87]);
    BiasedRNG[224] = (LFSRcolor0[250]&LFSRcolor0[50]&LFSRcolor0[115]);
    BiasedRNG[225] = (LFSRcolor0[506]&LFSRcolor0[573]&LFSRcolor0[911]);
    BiasedRNG[226] = (LFSRcolor0[330]&LFSRcolor0[230]&LFSRcolor0[468]);
    BiasedRNG[227] = (LFSRcolor0[935]&LFSRcolor0[254]&LFSRcolor0[505]);
    BiasedRNG[228] = (LFSRcolor0[167]&LFSRcolor0[929]&LFSRcolor0[424]);
    BiasedRNG[229] = (LFSRcolor0[861]&LFSRcolor0[117]&LFSRcolor0[142]);
    BiasedRNG[230] = (LFSRcolor0[486]&LFSRcolor0[228]&LFSRcolor0[591]);
    BiasedRNG[231] = (LFSRcolor0[183]&LFSRcolor0[138]&LFSRcolor0[242]);
    BiasedRNG[232] = (LFSRcolor0[527]&LFSRcolor0[605]&LFSRcolor0[229]);
    BiasedRNG[233] = (LFSRcolor0[97]&LFSRcolor0[787]&LFSRcolor0[186]);
    BiasedRNG[234] = (LFSRcolor0[739]&LFSRcolor0[432]&LFSRcolor0[376]);
    BiasedRNG[235] = (LFSRcolor0[163]&LFSRcolor0[45]&LFSRcolor0[269]);
    BiasedRNG[236] = (LFSRcolor0[823]&LFSRcolor0[462]&LFSRcolor0[203]);
    BiasedRNG[237] = (LFSRcolor0[493]&LFSRcolor0[154]&LFSRcolor0[742]);
    BiasedRNG[238] = (LFSRcolor0[77]&LFSRcolor0[832]&LFSRcolor0[682]);
    BiasedRNG[239] = (LFSRcolor0[756]&LFSRcolor0[620]&LFSRcolor0[728]);
    BiasedRNG[240] = (LFSRcolor0[39]&LFSRcolor0[95]&LFSRcolor0[927]);
    BiasedRNG[241] = (LFSRcolor0[438]&LFSRcolor0[849]&LFSRcolor0[171]);
    BiasedRNG[242] = (LFSRcolor0[790]&LFSRcolor0[64]&LFSRcolor0[446]);
    BiasedRNG[243] = (LFSRcolor0[366]&LFSRcolor0[724]&LFSRcolor0[476]);
    BiasedRNG[244] = (LFSRcolor0[157]&LFSRcolor0[926]&LFSRcolor0[129]);
    BiasedRNG[245] = (LFSRcolor0[352]&LFSRcolor0[528]&LFSRcolor0[10]);
    BiasedRNG[246] = (LFSRcolor0[348]&LFSRcolor0[627]&LFSRcolor0[26]);
    BiasedRNG[247] = (LFSRcolor0[103]&LFSRcolor0[509]&LFSRcolor0[539]);
    BiasedRNG[248] = (LFSRcolor0[611]&LFSRcolor0[323]&LFSRcolor0[178]);
    BiasedRNG[249] = (LFSRcolor0[41]&LFSRcolor0[324]&LFSRcolor0[222]);
    BiasedRNG[250] = (LFSRcolor0[826]&LFSRcolor0[314]&LFSRcolor0[703]);
    BiasedRNG[251] = (LFSRcolor0[544]&LFSRcolor0[730]&LFSRcolor0[931]);
    UnbiasedRNG[0] = LFSRcolor0[220];
    UnbiasedRNG[1] = LFSRcolor0[721];
    UnbiasedRNG[2] = LFSRcolor0[249];
    UnbiasedRNG[3] = LFSRcolor0[701];
    UnbiasedRNG[4] = LFSRcolor0[618];
    UnbiasedRNG[5] = LFSRcolor0[769];
    UnbiasedRNG[6] = LFSRcolor0[779];
    UnbiasedRNG[7] = LFSRcolor0[865];
    UnbiasedRNG[8] = LFSRcolor0[478];
    UnbiasedRNG[9] = LFSRcolor0[719];
    UnbiasedRNG[10] = LFSRcolor0[852];
    UnbiasedRNG[11] = LFSRcolor0[619];
    UnbiasedRNG[12] = LFSRcolor0[903];
    UnbiasedRNG[13] = LFSRcolor0[706];
    UnbiasedRNG[14] = LFSRcolor0[243];
    UnbiasedRNG[15] = LFSRcolor0[545];
    UnbiasedRNG[16] = LFSRcolor0[755];
    UnbiasedRNG[17] = LFSRcolor0[46];
    UnbiasedRNG[18] = LFSRcolor0[175];
    UnbiasedRNG[19] = LFSRcolor0[596];
    UnbiasedRNG[20] = LFSRcolor0[437];
    UnbiasedRNG[21] = LFSRcolor0[736];
    UnbiasedRNG[22] = LFSRcolor0[608];
    UnbiasedRNG[23] = LFSRcolor0[18];
    UnbiasedRNG[24] = LFSRcolor0[443];
    UnbiasedRNG[25] = LFSRcolor0[188];
    UnbiasedRNG[26] = LFSRcolor0[9];
    UnbiasedRNG[27] = LFSRcolor0[413];
    UnbiasedRNG[28] = LFSRcolor0[168];
    UnbiasedRNG[29] = LFSRcolor0[358];
    UnbiasedRNG[30] = LFSRcolor0[585];
    UnbiasedRNG[31] = LFSRcolor0[75];
    UnbiasedRNG[32] = LFSRcolor0[650];
    UnbiasedRNG[33] = LFSRcolor0[391];
    UnbiasedRNG[34] = LFSRcolor0[136];
    UnbiasedRNG[35] = LFSRcolor0[525];
    UnbiasedRNG[36] = LFSRcolor0[859];
    UnbiasedRNG[37] = LFSRcolor0[934];
    UnbiasedRNG[38] = LFSRcolor0[785];
    UnbiasedRNG[39] = LFSRcolor0[297];
    UnbiasedRNG[40] = LFSRcolor0[633];
    UnbiasedRNG[41] = LFSRcolor0[480];
    UnbiasedRNG[42] = LFSRcolor0[96];
    UnbiasedRNG[43] = LFSRcolor0[355];
    UnbiasedRNG[44] = LFSRcolor0[659];
    UnbiasedRNG[45] = LFSRcolor0[66];
    UnbiasedRNG[46] = LFSRcolor0[98];
    UnbiasedRNG[47] = LFSRcolor0[499];
    UnbiasedRNG[48] = LFSRcolor0[839];
    UnbiasedRNG[49] = LFSRcolor0[72];
    UnbiasedRNG[50] = LFSRcolor0[757];
    UnbiasedRNG[51] = LFSRcolor0[720];
    UnbiasedRNG[52] = LFSRcolor0[263];
    UnbiasedRNG[53] = LFSRcolor0[439];
    UnbiasedRNG[54] = LFSRcolor0[347];
    UnbiasedRNG[55] = LFSRcolor0[857];
    UnbiasedRNG[56] = LFSRcolor0[342];
    UnbiasedRNG[57] = LFSRcolor0[63];
    UnbiasedRNG[58] = LFSRcolor0[419];
    UnbiasedRNG[59] = LFSRcolor0[326];
    UnbiasedRNG[60] = LFSRcolor0[920];
    UnbiasedRNG[61] = LFSRcolor0[584];
    UnbiasedRNG[62] = LFSRcolor0[38];
    UnbiasedRNG[63] = LFSRcolor0[726];
    UnbiasedRNG[64] = LFSRcolor0[286];
    UnbiasedRNG[65] = LFSRcolor0[898];
    UnbiasedRNG[66] = LFSRcolor0[651];
    UnbiasedRNG[67] = LFSRcolor0[399];
    UnbiasedRNG[68] = LFSRcolor0[21];
    UnbiasedRNG[69] = LFSRcolor0[293];
    UnbiasedRNG[70] = LFSRcolor0[427];
    UnbiasedRNG[71] = LFSRcolor0[877];
    UnbiasedRNG[72] = LFSRcolor0[636];
    UnbiasedRNG[73] = LFSRcolor0[126];
    UnbiasedRNG[74] = LFSRcolor0[396];
    UnbiasedRNG[75] = LFSRcolor0[331];
    UnbiasedRNG[76] = LFSRcolor0[22];
    UnbiasedRNG[77] = LFSRcolor0[43];
    UnbiasedRNG[78] = LFSRcolor0[489];
    UnbiasedRNG[79] = LFSRcolor0[945];
    UnbiasedRNG[80] = LFSRcolor0[804];
    UnbiasedRNG[81] = LFSRcolor0[814];
    UnbiasedRNG[82] = LFSRcolor0[390];
    UnbiasedRNG[83] = LFSRcolor0[688];
    UnbiasedRNG[84] = LFSRcolor0[24];
    UnbiasedRNG[85] = LFSRcolor0[327];
    UnbiasedRNG[86] = LFSRcolor0[44];
    UnbiasedRNG[87] = LFSRcolor0[246];
    UnbiasedRNG[88] = LFSRcolor0[99];
    UnbiasedRNG[89] = LFSRcolor0[244];
    UnbiasedRNG[90] = LFSRcolor0[207];
    UnbiasedRNG[91] = LFSRcolor0[268];
    UnbiasedRNG[92] = LFSRcolor0[560];
    UnbiasedRNG[93] = LFSRcolor0[33];
    UnbiasedRNG[94] = LFSRcolor0[775];
    UnbiasedRNG[95] = LFSRcolor0[875];
    UnbiasedRNG[96] = LFSRcolor0[174];
    UnbiasedRNG[97] = LFSRcolor0[40];
    UnbiasedRNG[98] = LFSRcolor0[731];
    UnbiasedRNG[99] = LFSRcolor0[458];
    UnbiasedRNG[100] = LFSRcolor0[262];
    UnbiasedRNG[101] = LFSRcolor0[452];
    UnbiasedRNG[102] = LFSRcolor0[319];
    UnbiasedRNG[103] = LFSRcolor0[147];
    UnbiasedRNG[104] = LFSRcolor0[465];
    UnbiasedRNG[105] = LFSRcolor0[657];
    UnbiasedRNG[106] = LFSRcolor0[288];
    UnbiasedRNG[107] = LFSRcolor0[406];
    UnbiasedRNG[108] = LFSRcolor0[699];
    UnbiasedRNG[109] = LFSRcolor0[177];
    UnbiasedRNG[110] = LFSRcolor0[487];
    UnbiasedRNG[111] = LFSRcolor0[855];
    UnbiasedRNG[112] = LFSRcolor0[542];
    UnbiasedRNG[113] = LFSRcolor0[767];
    UnbiasedRNG[114] = LFSRcolor0[322];
    UnbiasedRNG[115] = LFSRcolor0[233];
    UnbiasedRNG[116] = LFSRcolor0[224];
    UnbiasedRNG[117] = LFSRcolor0[816];
    UnbiasedRNG[118] = LFSRcolor0[681];
    UnbiasedRNG[119] = LFSRcolor0[819];
    UnbiasedRNG[120] = LFSRcolor0[660];
    UnbiasedRNG[121] = LFSRcolor0[48];
    UnbiasedRNG[122] = LFSRcolor0[184];
    UnbiasedRNG[123] = LFSRcolor0[265];
    UnbiasedRNG[124] = LFSRcolor0[191];
    UnbiasedRNG[125] = LFSRcolor0[700];
    UnbiasedRNG[126] = LFSRcolor0[273];
    UnbiasedRNG[127] = LFSRcolor0[661];
    UnbiasedRNG[128] = LFSRcolor0[678];
    UnbiasedRNG[129] = LFSRcolor0[411];
    UnbiasedRNG[130] = LFSRcolor0[387];
    UnbiasedRNG[131] = LFSRcolor0[11];
    UnbiasedRNG[132] = LFSRcolor0[3];
    UnbiasedRNG[133] = LFSRcolor0[662];
    UnbiasedRNG[134] = LFSRcolor0[960];
    UnbiasedRNG[135] = LFSRcolor0[600];
    UnbiasedRNG[136] = LFSRcolor0[130];
    UnbiasedRNG[137] = LFSRcolor0[879];
    UnbiasedRNG[138] = LFSRcolor0[395];
    UnbiasedRNG[139] = LFSRcolor0[637];
    UnbiasedRNG[140] = LFSRcolor0[492];
    UnbiasedRNG[141] = LFSRcolor0[517];
    UnbiasedRNG[142] = LFSRcolor0[381];
    UnbiasedRNG[143] = LFSRcolor0[575];
    UnbiasedRNG[144] = LFSRcolor0[962];
    UnbiasedRNG[145] = LFSRcolor0[930];
    UnbiasedRNG[146] = LFSRcolor0[337];
    UnbiasedRNG[147] = LFSRcolor0[707];
    UnbiasedRNG[148] = LFSRcolor0[261];
    UnbiasedRNG[149] = LFSRcolor0[894];
    UnbiasedRNG[150] = LFSRcolor0[311];
    UnbiasedRNG[151] = LFSRcolor0[271];
    UnbiasedRNG[152] = LFSRcolor0[708];
    UnbiasedRNG[153] = LFSRcolor0[225];
    UnbiasedRNG[154] = LFSRcolor0[635];
    UnbiasedRNG[155] = LFSRcolor0[796];
    UnbiasedRNG[156] = LFSRcolor0[460];
    UnbiasedRNG[157] = LFSRcolor0[526];
    UnbiasedRNG[158] = LFSRcolor0[654];
    UnbiasedRNG[159] = LFSRcolor0[601];
    UnbiasedRNG[160] = LFSRcolor0[65];
    UnbiasedRNG[161] = LFSRcolor0[818];
    UnbiasedRNG[162] = LFSRcolor0[479];
    UnbiasedRNG[163] = LFSRcolor0[770];
    UnbiasedRNG[164] = LFSRcolor0[829];
    UnbiasedRNG[165] = LFSRcolor0[466];
    UnbiasedRNG[166] = LFSRcolor0[735];
    UnbiasedRNG[167] = LFSRcolor0[368];
    UnbiasedRNG[168] = LFSRcolor0[455];
    UnbiasedRNG[169] = LFSRcolor0[640];
    UnbiasedRNG[170] = LFSRcolor0[223];
    UnbiasedRNG[171] = LFSRcolor0[239];
    UnbiasedRNG[172] = LFSRcolor0[548];
    UnbiasedRNG[173] = LFSRcolor0[121];
    UnbiasedRNG[174] = LFSRcolor0[741];
    UnbiasedRNG[175] = LFSRcolor0[746];
    UnbiasedRNG[176] = LFSRcolor0[371];
    UnbiasedRNG[177] = LFSRcolor0[336];
    UnbiasedRNG[178] = LFSRcolor0[876];
    UnbiasedRNG[179] = LFSRcolor0[956];
    UnbiasedRNG[180] = LFSRcolor0[447];
    UnbiasedRNG[181] = LFSRcolor0[317];
    UnbiasedRNG[182] = LFSRcolor0[414];
    UnbiasedRNG[183] = LFSRcolor0[346];
    UnbiasedRNG[184] = LFSRcolor0[27];
    UnbiasedRNG[185] = LFSRcolor0[173];
    UnbiasedRNG[186] = LFSRcolor0[725];
    UnbiasedRNG[187] = LFSRcolor0[370];
    UnbiasedRNG[188] = LFSRcolor0[294];
    UnbiasedRNG[189] = LFSRcolor0[341];
    UnbiasedRNG[190] = LFSRcolor0[932];
    UnbiasedRNG[191] = LFSRcolor0[531];
    UnbiasedRNG[192] = LFSRcolor0[16];
    UnbiasedRNG[193] = LFSRcolor0[150];
    UnbiasedRNG[194] = LFSRcolor0[698];
    UnbiasedRNG[195] = LFSRcolor0[799];
    UnbiasedRNG[196] = LFSRcolor0[259];
    UnbiasedRNG[197] = LFSRcolor0[282];
    UnbiasedRNG[198] = LFSRcolor0[276];
    UnbiasedRNG[199] = LFSRcolor0[502];
    UnbiasedRNG[200] = LFSRcolor0[937];
    UnbiasedRNG[201] = LFSRcolor0[267];
    UnbiasedRNG[202] = LFSRcolor0[192];
    UnbiasedRNG[203] = LFSRcolor0[914];
    UnbiasedRNG[204] = LFSRcolor0[209];
    UnbiasedRNG[205] = LFSRcolor0[629];
    UnbiasedRNG[206] = LFSRcolor0[484];
    UnbiasedRNG[207] = LFSRcolor0[754];
    UnbiasedRNG[208] = LFSRcolor0[933];
end

always @(posedge color0_clk) begin
    BiasedRNG[252] = (LFSRcolor1[634]&LFSRcolor1[644]&LFSRcolor1[516]);
    BiasedRNG[253] = (LFSRcolor1[537]&LFSRcolor1[733]&LFSRcolor1[913]);
    BiasedRNG[254] = (LFSRcolor1[555]&LFSRcolor1[703]&LFSRcolor1[108]);
    BiasedRNG[255] = (LFSRcolor1[168]&LFSRcolor1[915]&LFSRcolor1[298]);
    BiasedRNG[256] = (LFSRcolor1[601]&LFSRcolor1[754]&LFSRcolor1[606]);
    BiasedRNG[257] = (LFSRcolor1[114]&LFSRcolor1[706]&LFSRcolor1[22]);
    BiasedRNG[258] = (LFSRcolor1[234]&LFSRcolor1[869]&LFSRcolor1[612]);
    BiasedRNG[259] = (LFSRcolor1[164]&LFSRcolor1[160]&LFSRcolor1[468]);
    BiasedRNG[260] = (LFSRcolor1[742]&LFSRcolor1[477]&LFSRcolor1[26]);
    BiasedRNG[261] = (LFSRcolor1[72]&LFSRcolor1[497]&LFSRcolor1[62]);
    BiasedRNG[262] = (LFSRcolor1[216]&LFSRcolor1[358]&LFSRcolor1[140]);
    BiasedRNG[263] = (LFSRcolor1[628]&LFSRcolor1[657]&LFSRcolor1[213]);
    BiasedRNG[264] = (LFSRcolor1[387]&LFSRcolor1[569]&LFSRcolor1[350]);
    BiasedRNG[265] = (LFSRcolor1[133]&LFSRcolor1[960]&LFSRcolor1[262]);
    BiasedRNG[266] = (LFSRcolor1[553]&LFSRcolor1[364]&LFSRcolor1[233]);
    BiasedRNG[267] = (LFSRcolor1[187]&LFSRcolor1[826]&LFSRcolor1[856]);
    BiasedRNG[268] = (LFSRcolor1[789]&LFSRcolor1[522]&LFSRcolor1[67]);
    BiasedRNG[269] = (LFSRcolor1[761]&LFSRcolor1[505]&LFSRcolor1[565]);
    BiasedRNG[270] = (LFSRcolor1[331]&LFSRcolor1[290]&LFSRcolor1[14]);
    BiasedRNG[271] = (LFSRcolor1[647]&LFSRcolor1[66]&LFSRcolor1[223]);
    BiasedRNG[272] = (LFSRcolor1[372]&LFSRcolor1[585]&LFSRcolor1[773]);
    BiasedRNG[273] = (LFSRcolor1[626]&LFSRcolor1[0]&LFSRcolor1[566]);
    BiasedRNG[274] = (LFSRcolor1[183]&LFSRcolor1[151]&LFSRcolor1[849]);
    BiasedRNG[275] = (LFSRcolor1[7]&LFSRcolor1[135]&LFSRcolor1[887]);
    BiasedRNG[276] = (LFSRcolor1[699]&LFSRcolor1[113]&LFSRcolor1[488]);
    BiasedRNG[277] = (LFSRcolor1[873]&LFSRcolor1[814]&LFSRcolor1[670]);
    BiasedRNG[278] = (LFSRcolor1[660]&LFSRcolor1[767]&LFSRcolor1[294]);
    BiasedRNG[279] = (LFSRcolor1[776]&LFSRcolor1[297]&LFSRcolor1[145]);
    BiasedRNG[280] = (LFSRcolor1[250]&LFSRcolor1[756]&LFSRcolor1[661]);
    BiasedRNG[281] = (LFSRcolor1[197]&LFSRcolor1[76]&LFSRcolor1[83]);
    BiasedRNG[282] = (LFSRcolor1[58]&LFSRcolor1[907]&LFSRcolor1[413]);
    BiasedRNG[283] = (LFSRcolor1[426]&LFSRcolor1[843]&LFSRcolor1[638]);
    BiasedRNG[284] = (LFSRcolor1[775]&LFSRcolor1[781]&LFSRcolor1[275]);
    BiasedRNG[285] = (LFSRcolor1[407]&LFSRcolor1[627]&LFSRcolor1[922]);
    BiasedRNG[286] = (LFSRcolor1[302]&LFSRcolor1[249]&LFSRcolor1[681]);
    BiasedRNG[287] = (LFSRcolor1[27]&LFSRcolor1[401]&LFSRcolor1[519]);
    BiasedRNG[288] = (LFSRcolor1[144]&LFSRcolor1[906]&LFSRcolor1[85]);
    BiasedRNG[289] = (LFSRcolor1[343]&LFSRcolor1[373]&LFSRcolor1[437]);
    BiasedRNG[290] = (LFSRcolor1[711]&LFSRcolor1[651]&LFSRcolor1[646]);
    BiasedRNG[291] = (LFSRcolor1[117]&LFSRcolor1[951]&LFSRcolor1[86]);
    BiasedRNG[292] = (LFSRcolor1[821]&LFSRcolor1[54]&LFSRcolor1[78]);
    BiasedRNG[293] = (LFSRcolor1[475]&LFSRcolor1[424]&LFSRcolor1[898]);
    BiasedRNG[294] = (LFSRcolor1[124]&LFSRcolor1[796]&LFSRcolor1[837]);
    BiasedRNG[295] = (LFSRcolor1[920]&LFSRcolor1[893]&LFSRcolor1[687]);
    BiasedRNG[296] = (LFSRcolor1[104]&LFSRcolor1[688]&LFSRcolor1[276]);
    BiasedRNG[297] = (LFSRcolor1[890]&LFSRcolor1[929]&LFSRcolor1[24]);
    BiasedRNG[298] = (LFSRcolor1[696]&LFSRcolor1[584]&LFSRcolor1[351]);
    BiasedRNG[299] = (LFSRcolor1[74]&LFSRcolor1[884]&LFSRcolor1[451]);
    BiasedRNG[300] = (LFSRcolor1[546]&LFSRcolor1[941]&LFSRcolor1[581]);
    BiasedRNG[301] = (LFSRcolor1[323]&LFSRcolor1[631]&LFSRcolor1[274]);
    BiasedRNG[302] = (LFSRcolor1[247]&LFSRcolor1[47]&LFSRcolor1[746]);
    BiasedRNG[303] = (LFSRcolor1[701]&LFSRcolor1[589]&LFSRcolor1[410]);
    BiasedRNG[304] = (LFSRcolor1[344]&LFSRcolor1[745]&LFSRcolor1[320]);
    BiasedRNG[305] = (LFSRcolor1[860]&LFSRcolor1[678]&LFSRcolor1[473]);
    BiasedRNG[306] = (LFSRcolor1[273]&LFSRcolor1[734]&LFSRcolor1[790]);
    BiasedRNG[307] = (LFSRcolor1[205]&LFSRcolor1[850]&LFSRcolor1[526]);
    BiasedRNG[308] = (LFSRcolor1[875]&LFSRcolor1[25]&LFSRcolor1[316]);
    BiasedRNG[309] = (LFSRcolor1[391]&LFSRcolor1[788]&LFSRcolor1[712]);
    BiasedRNG[310] = (LFSRcolor1[455]&LFSRcolor1[91]&LFSRcolor1[357]);
    BiasedRNG[311] = (LFSRcolor1[404]&LFSRcolor1[341]&LFSRcolor1[936]);
    BiasedRNG[312] = (LFSRcolor1[28]&LFSRcolor1[405]&LFSRcolor1[942]);
    BiasedRNG[313] = (LFSRcolor1[540]&LFSRcolor1[122]&LFSRcolor1[286]);
    BiasedRNG[314] = (LFSRcolor1[96]&LFSRcolor1[599]&LFSRcolor1[349]);
    BiasedRNG[315] = (LFSRcolor1[610]&LFSRcolor1[365]&LFSRcolor1[637]);
    BiasedRNG[316] = (LFSRcolor1[466]&LFSRcolor1[174]&LFSRcolor1[421]);
    BiasedRNG[317] = (LFSRcolor1[818]&LFSRcolor1[182]&LFSRcolor1[260]);
    BiasedRNG[318] = (LFSRcolor1[386]&LFSRcolor1[959]&LFSRcolor1[918]);
    BiasedRNG[319] = (LFSRcolor1[359]&LFSRcolor1[901]&LFSRcolor1[478]);
    BiasedRNG[320] = (LFSRcolor1[236]&LFSRcolor1[598]&LFSRcolor1[417]);
    BiasedRNG[321] = (LFSRcolor1[643]&LFSRcolor1[652]&LFSRcolor1[563]);
    BiasedRNG[322] = (LFSRcolor1[143]&LFSRcolor1[642]&LFSRcolor1[877]);
    BiasedRNG[323] = (LFSRcolor1[499]&LFSRcolor1[943]&LFSRcolor1[119]);
    BiasedRNG[324] = (LFSRcolor1[648]&LFSRcolor1[380]&LFSRcolor1[442]);
    BiasedRNG[325] = (LFSRcolor1[523]&LFSRcolor1[686]&LFSRcolor1[954]);
    BiasedRNG[326] = (LFSRcolor1[607]&LFSRcolor1[293]&LFSRcolor1[709]);
    BiasedRNG[327] = (LFSRcolor1[33]&LFSRcolor1[287]&LFSRcolor1[494]);
    BiasedRNG[328] = (LFSRcolor1[769]&LFSRcolor1[708]&LFSRcolor1[217]);
    BiasedRNG[329] = (LFSRcolor1[740]&LFSRcolor1[513]&LFSRcolor1[673]);
    BiasedRNG[330] = (LFSRcolor1[30]&LFSRcolor1[892]&LFSRcolor1[604]);
    BiasedRNG[331] = (LFSRcolor1[547]&LFSRcolor1[324]&LFSRcolor1[29]);
    BiasedRNG[332] = (LFSRcolor1[753]&LFSRcolor1[962]&LFSRcolor1[747]);
    BiasedRNG[333] = (LFSRcolor1[271]&LFSRcolor1[808]&LFSRcolor1[50]);
    BiasedRNG[334] = (LFSRcolor1[330]&LFSRcolor1[356]&LFSRcolor1[450]);
    BiasedRNG[335] = (LFSRcolor1[758]&LFSRcolor1[348]&LFSRcolor1[640]);
    BiasedRNG[336] = (LFSRcolor1[810]&LFSRcolor1[95]&LFSRcolor1[162]);
    BiasedRNG[337] = (LFSRcolor1[864]&LFSRcolor1[543]&LFSRcolor1[832]);
    BiasedRNG[338] = (LFSRcolor1[218]&LFSRcolor1[101]&LFSRcolor1[191]);
    BiasedRNG[339] = (LFSRcolor1[944]&LFSRcolor1[389]&LFSRcolor1[852]);
    BiasedRNG[340] = (LFSRcolor1[34]&LFSRcolor1[783]&LFSRcolor1[908]);
    BiasedRNG[341] = (LFSRcolor1[487]&LFSRcolor1[20]&LFSRcolor1[189]);
    BiasedRNG[342] = (LFSRcolor1[572]&LFSRcolor1[617]&LFSRcolor1[493]);
    BiasedRNG[343] = (LFSRcolor1[173]&LFSRcolor1[806]&LFSRcolor1[346]);
    BiasedRNG[344] = (LFSRcolor1[310]&LFSRcolor1[576]&LFSRcolor1[55]);
    BiasedRNG[345] = (LFSRcolor1[683]&LFSRcolor1[669]&LFSRcolor1[422]);
    BiasedRNG[346] = (LFSRcolor1[520]&LFSRcolor1[486]&LFSRcolor1[2]);
    BiasedRNG[347] = (LFSRcolor1[492]&LFSRcolor1[272]&LFSRcolor1[946]);
    BiasedRNG[348] = (LFSRcolor1[307]&LFSRcolor1[695]&LFSRcolor1[504]);
    BiasedRNG[349] = (LFSRcolor1[70]&LFSRcolor1[876]&LFSRcolor1[730]);
    BiasedRNG[350] = (LFSRcolor1[454]&LFSRcolor1[623]&LFSRcolor1[77]);
    BiasedRNG[351] = (LFSRcolor1[739]&LFSRcolor1[891]&LFSRcolor1[347]);
    BiasedRNG[352] = (LFSRcolor1[184]&LFSRcolor1[550]&LFSRcolor1[490]);
    BiasedRNG[353] = (LFSRcolor1[564]&LFSRcolor1[861]&LFSRcolor1[895]);
    BiasedRNG[354] = (LFSRcolor1[656]&LFSRcolor1[420]&LFSRcolor1[84]);
    BiasedRNG[355] = (LFSRcolor1[268]&LFSRcolor1[618]&LFSRcolor1[453]);
    BiasedRNG[356] = (LFSRcolor1[512]&LFSRcolor1[221]&LFSRcolor1[384]);
    BiasedRNG[357] = (LFSRcolor1[819]&LFSRcolor1[694]&LFSRcolor1[237]);
    BiasedRNG[358] = (LFSRcolor1[684]&LFSRcolor1[3]&LFSRcolor1[253]);
    BiasedRNG[359] = (LFSRcolor1[805]&LFSRcolor1[592]&LFSRcolor1[774]);
    BiasedRNG[360] = (LFSRcolor1[762]&LFSRcolor1[905]&LFSRcolor1[414]);
    BiasedRNG[361] = (LFSRcolor1[289]&LFSRcolor1[948]&LFSRcolor1[541]);
    BiasedRNG[362] = (LFSRcolor1[691]&LFSRcolor1[432]&LFSRcolor1[266]);
    BiasedRNG[363] = (LFSRcolor1[211]&LFSRcolor1[177]&LFSRcolor1[882]);
    BiasedRNG[364] = (LFSRcolor1[430]&LFSRcolor1[532]&LFSRcolor1[222]);
    BiasedRNG[365] = (LFSRcolor1[855]&LFSRcolor1[868]&LFSRcolor1[427]);
    BiasedRNG[366] = (LFSRcolor1[258]&LFSRcolor1[562]&LFSRcolor1[509]);
    BiasedRNG[367] = (LFSRcolor1[81]&LFSRcolor1[445]&LFSRcolor1[672]);
    BiasedRNG[368] = (LFSRcolor1[12]&LFSRcolor1[649]&LFSRcolor1[215]);
    BiasedRNG[369] = (LFSRcolor1[452]&LFSRcolor1[671]&LFSRcolor1[476]);
    BiasedRNG[370] = (LFSRcolor1[6]&LFSRcolor1[533]&LFSRcolor1[120]);
    BiasedRNG[371] = (LFSRcolor1[139]&LFSRcolor1[777]&LFSRcolor1[834]);
    BiasedRNG[372] = (LFSRcolor1[202]&LFSRcolor1[921]&LFSRcolor1[406]);
    BiasedRNG[373] = (LFSRcolor1[961]&LFSRcolor1[418]&LFSRcolor1[303]);
    BiasedRNG[374] = (LFSRcolor1[829]&LFSRcolor1[658]&LFSRcolor1[82]);
    BiasedRNG[375] = (LFSRcolor1[879]&LFSRcolor1[482]&LFSRcolor1[751]);
    BiasedRNG[376] = (LFSRcolor1[136]&LFSRcolor1[524]&LFSRcolor1[574]);
    BiasedRNG[377] = (LFSRcolor1[322]&LFSRcolor1[366]&LFSRcolor1[390]);
    BiasedRNG[378] = (LFSRcolor1[827]&LFSRcolor1[799]&LFSRcolor1[156]);
    BiasedRNG[379] = (LFSRcolor1[381]&LFSRcolor1[245]&LFSRcolor1[64]);
    BiasedRNG[380] = (LFSRcolor1[116]&LFSRcolor1[785]&LFSRcolor1[716]);
    BiasedRNG[381] = (LFSRcolor1[749]&LFSRcolor1[332]&LFSRcolor1[851]);
    BiasedRNG[382] = (LFSRcolor1[5]&LFSRcolor1[822]&LFSRcolor1[106]);
    BiasedRNG[383] = (LFSRcolor1[440]&LFSRcolor1[889]&LFSRcolor1[393]);
    BiasedRNG[384] = (LFSRcolor1[379]&LFSRcolor1[698]&LFSRcolor1[639]);
    BiasedRNG[385] = (LFSRcolor1[308]&LFSRcolor1[632]&LFSRcolor1[534]);
    BiasedRNG[386] = (LFSRcolor1[321]&LFSRcolor1[685]&LFSRcolor1[682]);
    BiasedRNG[387] = (LFSRcolor1[105]&LFSRcolor1[813]&LFSRcolor1[737]);
    BiasedRNG[388] = (LFSRcolor1[327]&LFSRcolor1[57]&LFSRcolor1[862]);
    BiasedRNG[389] = (LFSRcolor1[616]&LFSRcolor1[295]&LFSRcolor1[462]);
    BiasedRNG[390] = (LFSRcolor1[719]&LFSRcolor1[680]&LFSRcolor1[267]);
    BiasedRNG[391] = (LFSRcolor1[556]&LFSRcolor1[883]&LFSRcolor1[125]);
    BiasedRNG[392] = (LFSRcolor1[763]&LFSRcolor1[11]&LFSRcolor1[940]);
    BiasedRNG[393] = (LFSRcolor1[193]&LFSRcolor1[305]&LFSRcolor1[741]);
    BiasedRNG[394] = (LFSRcolor1[704]&LFSRcolor1[662]&LFSRcolor1[146]);
    BiasedRNG[395] = (LFSRcolor1[870]&LFSRcolor1[154]&LFSRcolor1[645]);
    BiasedRNG[396] = (LFSRcolor1[782]&LFSRcolor1[690]&LFSRcolor1[394]);
    BiasedRNG[397] = (LFSRcolor1[791]&LFSRcolor1[429]&LFSRcolor1[545]);
    BiasedRNG[398] = (LFSRcolor1[137]&LFSRcolor1[471]&LFSRcolor1[159]);
    BiasedRNG[399] = (LFSRcolor1[49]&LFSRcolor1[744]&LFSRcolor1[428]);
    BiasedRNG[400] = (LFSRcolor1[578]&LFSRcolor1[557]&LFSRcolor1[148]);
    BiasedRNG[401] = (LFSRcolor1[899]&LFSRcolor1[911]&LFSRcolor1[726]);
    BiasedRNG[402] = (LFSRcolor1[538]&LFSRcolor1[315]&LFSRcolor1[625]);
    BiasedRNG[403] = (LFSRcolor1[700]&LFSRcolor1[663]&LFSRcolor1[725]);
    BiasedRNG[404] = (LFSRcolor1[515]&LFSRcolor1[283]&LFSRcolor1[859]);
    BiasedRNG[405] = (LFSRcolor1[242]&LFSRcolor1[460]&LFSRcolor1[395]);
    BiasedRNG[406] = (LFSRcolor1[474]&LFSRcolor1[396]&LFSRcolor1[485]);
    BiasedRNG[407] = (LFSRcolor1[251]&LFSRcolor1[138]&LFSRcolor1[312]);
    BiasedRNG[408] = (LFSRcolor1[31]&LFSRcolor1[506]&LFSRcolor1[748]);
    BiasedRNG[409] = (LFSRcolor1[835]&LFSRcolor1[400]&LFSRcolor1[824]);
    BiasedRNG[410] = (LFSRcolor1[472]&LFSRcolor1[675]&LFSRcolor1[755]);
    BiasedRNG[411] = (LFSRcolor1[710]&LFSRcolor1[728]&LFSRcolor1[65]);
    BiasedRNG[412] = (LFSRcolor1[172]&LFSRcolor1[10]&LFSRcolor1[548]);
    BiasedRNG[413] = (LFSRcolor1[886]&LFSRcolor1[676]&LFSRcolor1[370]);
    BiasedRNG[414] = (LFSRcolor1[150]&LFSRcolor1[539]&LFSRcolor1[411]);
    BiasedRNG[415] = (LFSRcolor1[360]&LFSRcolor1[306]&LFSRcolor1[525]);
    BiasedRNG[416] = (LFSRcolor1[207]&LFSRcolor1[441]&LFSRcolor1[807]);
    BiasedRNG[417] = (LFSRcolor1[803]&LFSRcolor1[664]&LFSRcolor1[342]);
    BiasedRNG[418] = (LFSRcolor1[48]&LFSRcolor1[464]&LFSRcolor1[19]);
    BiasedRNG[419] = (LFSRcolor1[110]&LFSRcolor1[641]&LFSRcolor1[314]);
    BiasedRNG[420] = (LFSRcolor1[134]&LFSRcolor1[957]&LFSRcolor1[254]);
    BiasedRNG[421] = (LFSRcolor1[175]&LFSRcolor1[155]&LFSRcolor1[219]);
    BiasedRNG[422] = (LFSRcolor1[402]&LFSRcolor1[795]&LFSRcolor1[896]);
    BiasedRNG[423] = (LFSRcolor1[792]&LFSRcolor1[717]&LFSRcolor1[831]);
    BiasedRNG[424] = (LFSRcolor1[208]&LFSRcolor1[89]&LFSRcolor1[201]);
    BiasedRNG[425] = (LFSRcolor1[147]&LFSRcolor1[735]&LFSRcolor1[333]);
    BiasedRNG[426] = (LFSRcolor1[503]&LFSRcolor1[759]&LFSRcolor1[339]);
    BiasedRNG[427] = (LFSRcolor1[677]&LFSRcolor1[252]&LFSRcolor1[956]);
    BiasedRNG[428] = (LFSRcolor1[697]&LFSRcolor1[620]&LFSRcolor1[419]);
    BiasedRNG[429] = (LFSRcolor1[444]&LFSRcolor1[98]&LFSRcolor1[61]);
    BiasedRNG[430] = (LFSRcolor1[32]&LFSRcolor1[702]&LFSRcolor1[60]);
    BiasedRNG[431] = (LFSRcolor1[917]&LFSRcolor1[797]&LFSRcolor1[828]);
    BiasedRNG[432] = (LFSRcolor1[815]&LFSRcolor1[854]&LFSRcolor1[629]);
    BiasedRNG[433] = (LFSRcolor1[508]&LFSRcolor1[587]&LFSRcolor1[521]);
    BiasedRNG[434] = (LFSRcolor1[398]&LFSRcolor1[867]&LFSRcolor1[498]);
    BiasedRNG[435] = (LFSRcolor1[866]&LFSRcolor1[434]&LFSRcolor1[37]);
    BiasedRNG[436] = (LFSRcolor1[560]&LFSRcolor1[766]&LFSRcolor1[804]);
    BiasedRNG[437] = (LFSRcolor1[171]&LFSRcolor1[528]&LFSRcolor1[383]);
    BiasedRNG[438] = (LFSRcolor1[542]&LFSRcolor1[853]&LFSRcolor1[841]);
    BiasedRNG[439] = (LFSRcolor1[232]&LFSRcolor1[353]&LFSRcolor1[609]);
    BiasedRNG[440] = (LFSRcolor1[881]&LFSRcolor1[71]&LFSRcolor1[300]);
    BiasedRNG[441] = (LFSRcolor1[181]&LFSRcolor1[561]&LFSRcolor1[200]);
    BiasedRNG[442] = (LFSRcolor1[830]&LFSRcolor1[46]&LFSRcolor1[583]);
    BiasedRNG[443] = (LFSRcolor1[375]&LFSRcolor1[653]&LFSRcolor1[52]);
    BiasedRNG[444] = (LFSRcolor1[425]&LFSRcolor1[535]&LFSRcolor1[126]);
    BiasedRNG[445] = (LFSRcolor1[963]&LFSRcolor1[689]&LFSRcolor1[80]);
    BiasedRNG[446] = (LFSRcolor1[501]&LFSRcolor1[329]&LFSRcolor1[99]);
    BiasedRNG[447] = (LFSRcolor1[374]&LFSRcolor1[527]&LFSRcolor1[633]);
    BiasedRNG[448] = (LFSRcolor1[621]&LFSRcolor1[16]&LFSRcolor1[750]);
    BiasedRNG[449] = (LFSRcolor1[833]&LFSRcolor1[588]&LFSRcolor1[403]);
    BiasedRNG[450] = (LFSRcolor1[210]&LFSRcolor1[914]&LFSRcolor1[212]);
    BiasedRNG[451] = (LFSRcolor1[340]&LFSRcolor1[910]&LFSRcolor1[580]);
    BiasedRNG[452] = (LFSRcolor1[90]&LFSRcolor1[279]&LFSRcolor1[439]);
    BiasedRNG[453] = (LFSRcolor1[705]&LFSRcolor1[235]&LFSRcolor1[206]);
    BiasedRNG[454] = (LFSRcolor1[894]&LFSRcolor1[635]&LFSRcolor1[68]);
    BiasedRNG[455] = (LFSRcolor1[282]&LFSRcolor1[93]&LFSRcolor1[240]);
    BiasedRNG[456] = (LFSRcolor1[825]&LFSRcolor1[40]&LFSRcolor1[903]);
    BiasedRNG[457] = (LFSRcolor1[935]&LFSRcolor1[666]&LFSRcolor1[352]);
    BiasedRNG[458] = (LFSRcolor1[261]&LFSRcolor1[812]&LFSRcolor1[479]);
    BiasedRNG[459] = (LFSRcolor1[558]&LFSRcolor1[916]&LFSRcolor1[225]);
    BiasedRNG[460] = (LFSRcolor1[665]&LFSRcolor1[385]&LFSRcolor1[722]);
    BiasedRNG[461] = (LFSRcolor1[397]&LFSRcolor1[507]&LFSRcolor1[945]);
    BiasedRNG[462] = (LFSRcolor1[291]&LFSRcolor1[239]&LFSRcolor1[622]);
    BiasedRNG[463] = (LFSRcolor1[170]&LFSRcolor1[619]&LFSRcolor1[142]);
    BiasedRNG[464] = (LFSRcolor1[371]&LFSRcolor1[338]&LFSRcolor1[723]);
    BiasedRNG[465] = (LFSRcolor1[299]&LFSRcolor1[392]&LFSRcolor1[277]);
    BiasedRNG[466] = (LFSRcolor1[336]&LFSRcolor1[367]&LFSRcolor1[1]);
    BiasedRNG[467] = (LFSRcolor1[495]&LFSRcolor1[602]&LFSRcolor1[655]);
    BiasedRNG[468] = (LFSRcolor1[292]&LFSRcolor1[613]&LFSRcolor1[415]);
    BiasedRNG[469] = (LFSRcolor1[798]&LFSRcolor1[939]&LFSRcolor1[382]);
    BiasedRNG[470] = (LFSRcolor1[255]&LFSRcolor1[874]&LFSRcolor1[947]);
    BiasedRNG[471] = (LFSRcolor1[129]&LFSRcolor1[56]&LFSRcolor1[871]);
    BiasedRNG[472] = (LFSRcolor1[500]&LFSRcolor1[369]&LFSRcolor1[190]);
    BiasedRNG[473] = (LFSRcolor1[130]&LFSRcolor1[79]&LFSRcolor1[531]);
    BiasedRNG[474] = (LFSRcolor1[465]&LFSRcolor1[771]&LFSRcolor1[284]);
    BiasedRNG[475] = (LFSRcolor1[39]&LFSRcolor1[209]&LFSRcolor1[467]);
    BiasedRNG[476] = (LFSRcolor1[227]&LFSRcolor1[44]&LFSRcolor1[158]);
    BiasedRNG[477] = (LFSRcolor1[611]&LFSRcolor1[600]&LFSRcolor1[551]);
    BiasedRNG[478] = (LFSRcolor1[912]&LFSRcolor1[559]&LFSRcolor1[169]);
    BiasedRNG[479] = (LFSRcolor1[409]&LFSRcolor1[301]&LFSRcolor1[337]);
    BiasedRNG[480] = (LFSRcolor1[377]&LFSRcolor1[707]&LFSRcolor1[842]);
    BiasedRNG[481] = (LFSRcolor1[165]&LFSRcolor1[765]&LFSRcolor1[502]);
    BiasedRNG[482] = (LFSRcolor1[123]&LFSRcolor1[176]&LFSRcolor1[636]);
    BiasedRNG[483] = (LFSRcolor1[313]&LFSRcolor1[319]&LFSRcolor1[127]);
    BiasedRNG[484] = (LFSRcolor1[265]&LFSRcolor1[570]&LFSRcolor1[536]);
    BiasedRNG[485] = (LFSRcolor1[423]&LFSRcolor1[844]&LFSRcolor1[100]);
    BiasedRNG[486] = (LFSRcolor1[594]&LFSRcolor1[368]&LFSRcolor1[484]);
    BiasedRNG[487] = (LFSRcolor1[412]&LFSRcolor1[128]&LFSRcolor1[752]);
    BiasedRNG[488] = (LFSRcolor1[923]&LFSRcolor1[102]&LFSRcolor1[848]);
    BiasedRNG[489] = (LFSRcolor1[469]&LFSRcolor1[318]&LFSRcolor1[668]);
    BiasedRNG[490] = (LFSRcolor1[256]&LFSRcolor1[816]&LFSRcolor1[933]);
    BiasedRNG[491] = (LFSRcolor1[888]&LFSRcolor1[226]&LFSRcolor1[679]);
    BiasedRNG[492] = (LFSRcolor1[729]&LFSRcolor1[431]&LFSRcolor1[721]);
    BiasedRNG[493] = (LFSRcolor1[567]&LFSRcolor1[480]&LFSRcolor1[624]);
    BiasedRNG[494] = (LFSRcolor1[285]&LFSRcolor1[720]&LFSRcolor1[713]);
    BiasedRNG[495] = (LFSRcolor1[220]&LFSRcolor1[111]&LFSRcolor1[794]);
    BiasedRNG[496] = (LFSRcolor1[35]&LFSRcolor1[667]&LFSRcolor1[772]);
    BiasedRNG[497] = (LFSRcolor1[614]&LFSRcolor1[334]&LFSRcolor1[483]);
    BiasedRNG[498] = (LFSRcolor1[549]&LFSRcolor1[399]&LFSRcolor1[311]);
    BiasedRNG[499] = (LFSRcolor1[582]&LFSRcolor1[654]&LFSRcolor1[186]);
    BiasedRNG[500] = (LFSRcolor1[731]&LFSRcolor1[801]&LFSRcolor1[17]);
    BiasedRNG[501] = (LFSRcolor1[408]&LFSRcolor1[443]&LFSRcolor1[650]);
    BiasedRNG[502] = (LFSRcolor1[109]&LFSRcolor1[840]&LFSRcolor1[904]);
    UnbiasedRNG[209] = LFSRcolor1[857];
    UnbiasedRNG[210] = LFSRcolor1[764];
    UnbiasedRNG[211] = LFSRcolor1[244];
    UnbiasedRNG[212] = LFSRcolor1[4];
    UnbiasedRNG[213] = LFSRcolor1[309];
    UnbiasedRNG[214] = LFSRcolor1[180];
    UnbiasedRNG[215] = LFSRcolor1[447];
    UnbiasedRNG[216] = LFSRcolor1[304];
    UnbiasedRNG[217] = LFSRcolor1[161];
    UnbiasedRNG[218] = LFSRcolor1[579];
    UnbiasedRNG[219] = LFSRcolor1[38];
    UnbiasedRNG[220] = LFSRcolor1[264];
    UnbiasedRNG[221] = LFSRcolor1[597];
    UnbiasedRNG[222] = LFSRcolor1[97];
    UnbiasedRNG[223] = LFSRcolor1[446];
    UnbiasedRNG[224] = LFSRcolor1[388];
    UnbiasedRNG[225] = LFSRcolor1[470];
    UnbiasedRNG[226] = LFSRcolor1[902];
    UnbiasedRNG[227] = LFSRcolor1[811];
    UnbiasedRNG[228] = LFSRcolor1[107];
    UnbiasedRNG[229] = LFSRcolor1[928];
    UnbiasedRNG[230] = LFSRcolor1[328];
    UnbiasedRNG[231] = LFSRcolor1[511];
    UnbiasedRNG[232] = LFSRcolor1[885];
    UnbiasedRNG[233] = LFSRcolor1[94];
    UnbiasedRNG[234] = LFSRcolor1[934];
    UnbiasedRNG[235] = LFSRcolor1[489];
    UnbiasedRNG[236] = LFSRcolor1[768];
    UnbiasedRNG[237] = LFSRcolor1[214];
    UnbiasedRNG[238] = LFSRcolor1[88];
    UnbiasedRNG[239] = LFSRcolor1[897];
    UnbiasedRNG[240] = LFSRcolor1[839];
    UnbiasedRNG[241] = LFSRcolor1[593];
    UnbiasedRNG[242] = LFSRcolor1[456];
    UnbiasedRNG[243] = LFSRcolor1[438];
    UnbiasedRNG[244] = LFSRcolor1[296];
    UnbiasedRNG[245] = LFSRcolor1[378];
    UnbiasedRNG[246] = LFSRcolor1[778];
    UnbiasedRNG[247] = LFSRcolor1[952];
    UnbiasedRNG[248] = LFSRcolor1[836];
    UnbiasedRNG[249] = LFSRcolor1[760];
    UnbiasedRNG[250] = LFSRcolor1[577];
    UnbiasedRNG[251] = LFSRcolor1[457];
    UnbiasedRNG[252] = LFSRcolor1[847];
    UnbiasedRNG[253] = LFSRcolor1[463];
    UnbiasedRNG[254] = LFSRcolor1[163];
    UnbiasedRNG[255] = LFSRcolor1[15];
    UnbiasedRNG[256] = LFSRcolor1[800];
    UnbiasedRNG[257] = LFSRcolor1[288];
    UnbiasedRNG[258] = LFSRcolor1[416];
    UnbiasedRNG[259] = LFSRcolor1[802];
    UnbiasedRNG[260] = LFSRcolor1[121];
    UnbiasedRNG[261] = LFSRcolor1[779];
    UnbiasedRNG[262] = LFSRcolor1[529];
    UnbiasedRNG[263] = LFSRcolor1[518];
    UnbiasedRNG[264] = LFSRcolor1[263];
    UnbiasedRNG[265] = LFSRcolor1[909];
    UnbiasedRNG[266] = LFSRcolor1[153];
    UnbiasedRNG[267] = LFSRcolor1[59];
    UnbiasedRNG[268] = LFSRcolor1[727];
    UnbiasedRNG[269] = LFSRcolor1[591];
    UnbiasedRNG[270] = LFSRcolor1[693];
    UnbiasedRNG[271] = LFSRcolor1[793];
    UnbiasedRNG[272] = LFSRcolor1[937];
    UnbiasedRNG[273] = LFSRcolor1[198];
    UnbiasedRNG[274] = LFSRcolor1[132];
    UnbiasedRNG[275] = LFSRcolor1[448];
    UnbiasedRNG[276] = LFSRcolor1[157];
    UnbiasedRNG[277] = LFSRcolor1[517];
    UnbiasedRNG[278] = LFSRcolor1[491];
    UnbiasedRNG[279] = LFSRcolor1[953];
    UnbiasedRNG[280] = LFSRcolor1[166];
    UnbiasedRNG[281] = LFSRcolor1[45];
    UnbiasedRNG[282] = LFSRcolor1[112];
    UnbiasedRNG[283] = LFSRcolor1[335];
    UnbiasedRNG[284] = LFSRcolor1[13];
    UnbiasedRNG[285] = LFSRcolor1[732];
    UnbiasedRNG[286] = LFSRcolor1[595];
    UnbiasedRNG[287] = LFSRcolor1[362];
    UnbiasedRNG[288] = LFSRcolor1[141];
    UnbiasedRNG[289] = LFSRcolor1[436];
    UnbiasedRNG[290] = LFSRcolor1[243];
    UnbiasedRNG[291] = LFSRcolor1[51];
    UnbiasedRNG[292] = LFSRcolor1[586];
    UnbiasedRNG[293] = LFSRcolor1[780];
    UnbiasedRNG[294] = LFSRcolor1[281];
    UnbiasedRNG[295] = LFSRcolor1[568];
    UnbiasedRNG[296] = LFSRcolor1[269];
    UnbiasedRNG[297] = LFSRcolor1[18];
    UnbiasedRNG[298] = LFSRcolor1[9];
    UnbiasedRNG[299] = LFSRcolor1[194];
    UnbiasedRNG[300] = LFSRcolor1[715];
    UnbiasedRNG[301] = LFSRcolor1[554];
    UnbiasedRNG[302] = LFSRcolor1[192];
    UnbiasedRNG[303] = LFSRcolor1[103];
    UnbiasedRNG[304] = LFSRcolor1[964];
    UnbiasedRNG[305] = LFSRcolor1[858];
    UnbiasedRNG[306] = LFSRcolor1[8];
    UnbiasedRNG[307] = LFSRcolor1[195];
    UnbiasedRNG[308] = LFSRcolor1[927];
    UnbiasedRNG[309] = LFSRcolor1[757];
    UnbiasedRNG[310] = LFSRcolor1[573];
    UnbiasedRNG[311] = LFSRcolor1[196];
    UnbiasedRNG[312] = LFSRcolor1[496];
    UnbiasedRNG[313] = LFSRcolor1[544];
    UnbiasedRNG[314] = LFSRcolor1[204];
    UnbiasedRNG[315] = LFSRcolor1[270];
    UnbiasedRNG[316] = LFSRcolor1[965];
    UnbiasedRNG[317] = LFSRcolor1[185];
    UnbiasedRNG[318] = LFSRcolor1[552];
    UnbiasedRNG[319] = LFSRcolor1[743];
    UnbiasedRNG[320] = LFSRcolor1[92];
    UnbiasedRNG[321] = LFSRcolor1[229];
    UnbiasedRNG[322] = LFSRcolor1[530];
    UnbiasedRNG[323] = LFSRcolor1[458];
    UnbiasedRNG[324] = LFSRcolor1[510];
    UnbiasedRNG[325] = LFSRcolor1[930];
    UnbiasedRNG[326] = LFSRcolor1[949];
    UnbiasedRNG[327] = LFSRcolor1[846];
    UnbiasedRNG[328] = LFSRcolor1[900];
    UnbiasedRNG[329] = LFSRcolor1[43];
    UnbiasedRNG[330] = LFSRcolor1[188];
    UnbiasedRNG[331] = LFSRcolor1[257];
    UnbiasedRNG[332] = LFSRcolor1[231];
    UnbiasedRNG[333] = LFSRcolor1[199];
    UnbiasedRNG[334] = LFSRcolor1[924];
    UnbiasedRNG[335] = LFSRcolor1[809];
    UnbiasedRNG[336] = LFSRcolor1[958];
    UnbiasedRNG[337] = LFSRcolor1[354];
    UnbiasedRNG[338] = LFSRcolor1[931];
    UnbiasedRNG[339] = LFSRcolor1[230];
    UnbiasedRNG[340] = LFSRcolor1[21];
    UnbiasedRNG[341] = LFSRcolor1[75];
    UnbiasedRNG[342] = LFSRcolor1[838];
    UnbiasedRNG[343] = LFSRcolor1[178];
    UnbiasedRNG[344] = LFSRcolor1[596];
    UnbiasedRNG[345] = LFSRcolor1[575];
    UnbiasedRNG[346] = LFSRcolor1[325];
    UnbiasedRNG[347] = LFSRcolor1[42];
    UnbiasedRNG[348] = LFSRcolor1[770];
    UnbiasedRNG[349] = LFSRcolor1[73];
    UnbiasedRNG[350] = LFSRcolor1[674];
    UnbiasedRNG[351] = LFSRcolor1[692];
    UnbiasedRNG[352] = LFSRcolor1[149];
    UnbiasedRNG[353] = LFSRcolor1[820];
    UnbiasedRNG[354] = LFSRcolor1[87];
    UnbiasedRNG[355] = LFSRcolor1[326];
    UnbiasedRNG[356] = LFSRcolor1[317];
    UnbiasedRNG[357] = LFSRcolor1[784];
    UnbiasedRNG[358] = LFSRcolor1[152];
    UnbiasedRNG[359] = LFSRcolor1[817];
    UnbiasedRNG[360] = LFSRcolor1[926];
    UnbiasedRNG[361] = LFSRcolor1[938];
    UnbiasedRNG[362] = LFSRcolor1[872];
    UnbiasedRNG[363] = LFSRcolor1[241];
    UnbiasedRNG[364] = LFSRcolor1[608];
    UnbiasedRNG[365] = LFSRcolor1[514];
    UnbiasedRNG[366] = LFSRcolor1[228];
    UnbiasedRNG[367] = LFSRcolor1[449];
    UnbiasedRNG[368] = LFSRcolor1[615];
    UnbiasedRNG[369] = LFSRcolor1[53];
    UnbiasedRNG[370] = LFSRcolor1[361];
    UnbiasedRNG[371] = LFSRcolor1[955];
    UnbiasedRNG[372] = LFSRcolor1[481];
    UnbiasedRNG[373] = LFSRcolor1[659];
    UnbiasedRNG[374] = LFSRcolor1[603];
    UnbiasedRNG[375] = LFSRcolor1[714];
    UnbiasedRNG[376] = LFSRcolor1[238];
    UnbiasedRNG[377] = LFSRcolor1[863];
    UnbiasedRNG[378] = LFSRcolor1[259];
    UnbiasedRNG[379] = LFSRcolor1[167];
    UnbiasedRNG[380] = LFSRcolor1[919];
    UnbiasedRNG[381] = LFSRcolor1[69];
    UnbiasedRNG[382] = LFSRcolor1[932];
    UnbiasedRNG[383] = LFSRcolor1[131];
    UnbiasedRNG[384] = LFSRcolor1[845];
    UnbiasedRNG[385] = LFSRcolor1[724];
end

always @(posedge color1_clk) begin
    BiasedRNG[503] = (LFSRcolor2[422]&LFSRcolor2[591]&LFSRcolor2[421]);
    BiasedRNG[504] = (LFSRcolor2[543]&LFSRcolor2[760]&LFSRcolor2[607]);
    BiasedRNG[505] = (LFSRcolor2[62]&LFSRcolor2[181]&LFSRcolor2[114]);
    BiasedRNG[506] = (LFSRcolor2[465]&LFSRcolor2[358]&LFSRcolor2[140]);
    BiasedRNG[507] = (LFSRcolor2[538]&LFSRcolor2[96]&LFSRcolor2[341]);
    BiasedRNG[508] = (LFSRcolor2[729]&LFSRcolor2[228]&LFSRcolor2[582]);
    BiasedRNG[509] = (LFSRcolor2[342]&LFSRcolor2[734]&LFSRcolor2[605]);
    BiasedRNG[510] = (LFSRcolor2[454]&LFSRcolor2[630]&LFSRcolor2[455]);
    BiasedRNG[511] = (LFSRcolor2[268]&LFSRcolor2[541]&LFSRcolor2[484]);
    BiasedRNG[512] = (LFSRcolor2[537]&LFSRcolor2[194]&LFSRcolor2[709]);
    BiasedRNG[513] = (LFSRcolor2[731]&LFSRcolor2[450]&LFSRcolor2[104]);
    BiasedRNG[514] = (LFSRcolor2[409]&LFSRcolor2[156]&LFSRcolor2[755]);
    BiasedRNG[515] = (LFSRcolor2[256]&LFSRcolor2[386]&LFSRcolor2[74]);
    BiasedRNG[516] = (LFSRcolor2[631]&LFSRcolor2[395]&LFSRcolor2[171]);
    BiasedRNG[517] = (LFSRcolor2[456]&LFSRcolor2[553]&LFSRcolor2[135]);
    BiasedRNG[518] = (LFSRcolor2[682]&LFSRcolor2[602]&LFSRcolor2[469]);
    BiasedRNG[519] = (LFSRcolor2[671]&LFSRcolor2[153]&LFSRcolor2[761]);
    BiasedRNG[520] = (LFSRcolor2[38]&LFSRcolor2[511]&LFSRcolor2[776]);
    BiasedRNG[521] = (LFSRcolor2[752]&LFSRcolor2[252]&LFSRcolor2[661]);
    BiasedRNG[522] = (LFSRcolor2[740]&LFSRcolor2[41]&LFSRcolor2[416]);
    BiasedRNG[523] = (LFSRcolor2[133]&LFSRcolor2[245]&LFSRcolor2[247]);
    BiasedRNG[524] = (LFSRcolor2[64]&LFSRcolor2[467]&LFSRcolor2[647]);
    BiasedRNG[525] = (LFSRcolor2[211]&LFSRcolor2[2]&LFSRcolor2[372]);
    BiasedRNG[526] = (LFSRcolor2[585]&LFSRcolor2[684]&LFSRcolor2[498]);
    BiasedRNG[527] = (LFSRcolor2[219]&LFSRcolor2[446]&LFSRcolor2[54]);
    BiasedRNG[528] = (LFSRcolor2[218]&LFSRcolor2[183]&LFSRcolor2[21]);
    BiasedRNG[529] = (LFSRcolor2[435]&LFSRcolor2[102]&LFSRcolor2[742]);
    BiasedRNG[530] = (LFSRcolor2[284]&LFSRcolor2[390]&LFSRcolor2[5]);
    BiasedRNG[531] = (LFSRcolor2[509]&LFSRcolor2[559]&LFSRcolor2[632]);
    BiasedRNG[532] = (LFSRcolor2[733]&LFSRcolor2[115]&LFSRcolor2[549]);
    BiasedRNG[533] = (LFSRcolor2[70]&LFSRcolor2[65]&LFSRcolor2[300]);
    BiasedRNG[534] = (LFSRcolor2[657]&LFSRcolor2[376]&LFSRcolor2[656]);
    BiasedRNG[535] = (LFSRcolor2[52]&LFSRcolor2[578]&LFSRcolor2[72]);
    BiasedRNG[536] = (LFSRcolor2[556]&LFSRcolor2[448]&LFSRcolor2[179]);
    BiasedRNG[537] = (LFSRcolor2[151]&LFSRcolor2[606]&LFSRcolor2[637]);
    BiasedRNG[538] = (LFSRcolor2[46]&LFSRcolor2[476]&LFSRcolor2[127]);
    BiasedRNG[539] = (LFSRcolor2[173]&LFSRcolor2[583]&LFSRcolor2[109]);
    BiasedRNG[540] = (LFSRcolor2[59]&LFSRcolor2[536]&LFSRcolor2[379]);
    BiasedRNG[541] = (LFSRcolor2[233]&LFSRcolor2[191]&LFSRcolor2[562]);
    BiasedRNG[542] = (LFSRcolor2[380]&LFSRcolor2[333]&LFSRcolor2[285]);
    BiasedRNG[543] = (LFSRcolor2[6]&LFSRcolor2[43]&LFSRcolor2[129]);
    BiasedRNG[544] = (LFSRcolor2[419]&LFSRcolor2[719]&LFSRcolor2[569]);
    BiasedRNG[545] = (LFSRcolor2[311]&LFSRcolor2[576]&LFSRcolor2[236]);
    BiasedRNG[546] = (LFSRcolor2[126]&LFSRcolor2[44]&LFSRcolor2[551]);
    BiasedRNG[547] = (LFSRcolor2[113]&LFSRcolor2[330]&LFSRcolor2[513]);
    BiasedRNG[548] = (LFSRcolor2[616]&LFSRcolor2[753]&LFSRcolor2[77]);
    BiasedRNG[549] = (LFSRcolor2[525]&LFSRcolor2[257]&LFSRcolor2[94]);
    BiasedRNG[550] = (LFSRcolor2[778]&LFSRcolor2[370]&LFSRcolor2[739]);
    BiasedRNG[551] = (LFSRcolor2[462]&LFSRcolor2[651]&LFSRcolor2[519]);
    BiasedRNG[552] = (LFSRcolor2[499]&LFSRcolor2[720]&LFSRcolor2[442]);
    BiasedRNG[553] = (LFSRcolor2[410]&LFSRcolor2[412]&LFSRcolor2[779]);
    BiasedRNG[554] = (LFSRcolor2[222]&LFSRcolor2[666]&LFSRcolor2[33]);
    BiasedRNG[555] = (LFSRcolor2[565]&LFSRcolor2[327]&LFSRcolor2[526]);
    BiasedRNG[556] = (LFSRcolor2[600]&LFSRcolor2[401]&LFSRcolor2[706]);
    BiasedRNG[557] = (LFSRcolor2[320]&LFSRcolor2[533]&LFSRcolor2[107]);
    BiasedRNG[558] = (LFSRcolor2[482]&LFSRcolor2[662]&LFSRcolor2[348]);
    BiasedRNG[559] = (LFSRcolor2[571]&LFSRcolor2[491]&LFSRcolor2[237]);
    BiasedRNG[560] = (LFSRcolor2[717]&LFSRcolor2[766]&LFSRcolor2[80]);
    BiasedRNG[561] = (LFSRcolor2[26]&LFSRcolor2[564]&LFSRcolor2[627]);
    BiasedRNG[562] = (LFSRcolor2[30]&LFSRcolor2[449]&LFSRcolor2[681]);
    BiasedRNG[563] = (LFSRcolor2[404]&LFSRcolor2[580]&LFSRcolor2[28]);
    BiasedRNG[564] = (LFSRcolor2[172]&LFSRcolor2[293]&LFSRcolor2[638]);
    BiasedRNG[565] = (LFSRcolor2[770]&LFSRcolor2[396]&LFSRcolor2[481]);
    BiasedRNG[566] = (LFSRcolor2[203]&LFSRcolor2[433]&LFSRcolor2[597]);
    BiasedRNG[567] = (LFSRcolor2[636]&LFSRcolor2[303]&LFSRcolor2[741]);
    BiasedRNG[568] = (LFSRcolor2[346]&LFSRcolor2[88]&LFSRcolor2[366]);
    BiasedRNG[569] = (LFSRcolor2[712]&LFSRcolor2[275]&LFSRcolor2[383]);
    BiasedRNG[570] = (LFSRcolor2[425]&LFSRcolor2[313]&LFSRcolor2[8]);
    BiasedRNG[571] = (LFSRcolor2[361]&LFSRcolor2[276]&LFSRcolor2[360]);
    BiasedRNG[572] = (LFSRcolor2[686]&LFSRcolor2[633]&LFSRcolor2[305]);
    BiasedRNG[573] = (LFSRcolor2[110]&LFSRcolor2[216]&LFSRcolor2[772]);
    BiasedRNG[574] = (LFSRcolor2[66]&LFSRcolor2[163]&LFSRcolor2[234]);
    BiasedRNG[575] = (LFSRcolor2[326]&LFSRcolor2[150]&LFSRcolor2[232]);
    BiasedRNG[576] = (LFSRcolor2[208]&LFSRcolor2[590]&LFSRcolor2[321]);
    BiasedRNG[577] = (LFSRcolor2[47]&LFSRcolor2[773]&LFSRcolor2[267]);
    BiasedRNG[578] = (LFSRcolor2[375]&LFSRcolor2[458]&LFSRcolor2[318]);
    BiasedRNG[579] = (LFSRcolor2[78]&LFSRcolor2[473]&LFSRcolor2[13]);
    BiasedRNG[580] = (LFSRcolor2[143]&LFSRcolor2[501]&LFSRcolor2[197]);
    BiasedRNG[581] = (LFSRcolor2[418]&LFSRcolor2[642]&LFSRcolor2[122]);
    BiasedRNG[582] = (LFSRcolor2[653]&LFSRcolor2[413]&LFSRcolor2[92]);
    BiasedRNG[583] = (LFSRcolor2[302]&LFSRcolor2[75]&LFSRcolor2[25]);
    BiasedRNG[584] = (LFSRcolor2[148]&LFSRcolor2[215]&LFSRcolor2[459]);
    BiasedRNG[585] = (LFSRcolor2[601]&LFSRcolor2[356]&LFSRcolor2[699]);
    BiasedRNG[586] = (LFSRcolor2[161]&LFSRcolor2[20]&LFSRcolor2[744]);
    BiasedRNG[587] = (LFSRcolor2[394]&LFSRcolor2[166]&LFSRcolor2[673]);
    BiasedRNG[588] = (LFSRcolor2[202]&LFSRcolor2[587]&LFSRcolor2[29]);
    BiasedRNG[589] = (LFSRcolor2[334]&LFSRcolor2[730]&LFSRcolor2[344]);
    BiasedRNG[590] = (LFSRcolor2[725]&LFSRcolor2[175]&LFSRcolor2[497]);
    BiasedRNG[591] = (LFSRcolor2[97]&LFSRcolor2[679]&LFSRcolor2[596]);
    BiasedRNG[592] = (LFSRcolor2[472]&LFSRcolor2[286]&LFSRcolor2[138]);
    BiasedRNG[593] = (LFSRcolor2[746]&LFSRcolor2[69]&LFSRcolor2[735]);
    BiasedRNG[594] = (LFSRcolor2[242]&LFSRcolor2[613]&LFSRcolor2[121]);
    BiasedRNG[595] = (LFSRcolor2[243]&LFSRcolor2[468]&LFSRcolor2[437]);
    BiasedRNG[596] = (LFSRcolor2[475]&LFSRcolor2[728]&LFSRcolor2[40]);
    BiasedRNG[597] = (LFSRcolor2[521]&LFSRcolor2[354]&LFSRcolor2[518]);
    BiasedRNG[598] = (LFSRcolor2[81]&LFSRcolor2[178]&LFSRcolor2[301]);
    BiasedRNG[599] = (LFSRcolor2[750]&LFSRcolor2[137]&LFSRcolor2[263]);
    BiasedRNG[600] = (LFSRcolor2[598]&LFSRcolor2[480]&LFSRcolor2[406]);
    BiasedRNG[601] = (LFSRcolor2[101]&LFSRcolor2[781]&LFSRcolor2[723]);
    BiasedRNG[602] = (LFSRcolor2[169]&LFSRcolor2[447]&LFSRcolor2[620]);
    BiasedRNG[603] = (LFSRcolor2[507]&LFSRcolor2[331]&LFSRcolor2[603]);
    BiasedRNG[604] = (LFSRcolor2[7]&LFSRcolor2[309]&LFSRcolor2[540]);
    BiasedRNG[605] = (LFSRcolor2[697]&LFSRcolor2[691]&LFSRcolor2[160]);
    BiasedRNG[606] = (LFSRcolor2[748]&LFSRcolor2[665]&LFSRcolor2[639]);
    BiasedRNG[607] = (LFSRcolor2[307]&LFSRcolor2[550]&LFSRcolor2[758]);
    BiasedRNG[608] = (LFSRcolor2[512]&LFSRcolor2[223]&LFSRcolor2[106]);
    BiasedRNG[609] = (LFSRcolor2[369]&LFSRcolor2[310]&LFSRcolor2[705]);
    BiasedRNG[610] = (LFSRcolor2[235]&LFSRcolor2[572]&LFSRcolor2[438]);
    BiasedRNG[611] = (LFSRcolor2[349]&LFSRcolor2[269]&LFSRcolor2[58]);
    BiasedRNG[612] = (LFSRcolor2[198]&LFSRcolor2[83]&LFSRcolor2[124]);
    BiasedRNG[613] = (LFSRcolor2[643]&LFSRcolor2[316]&LFSRcolor2[288]);
    BiasedRNG[614] = (LFSRcolor2[514]&LFSRcolor2[677]&LFSRcolor2[402]);
    BiasedRNG[615] = (LFSRcolor2[589]&LFSRcolor2[60]&LFSRcolor2[534]);
    BiasedRNG[616] = (LFSRcolor2[152]&LFSRcolor2[251]&LFSRcolor2[667]);
    BiasedRNG[617] = (LFSRcolor2[299]&LFSRcolor2[420]&LFSRcolor2[11]);
    BiasedRNG[618] = (LFSRcolor2[707]&LFSRcolor2[767]&LFSRcolor2[452]);
    BiasedRNG[619] = (LFSRcolor2[339]&LFSRcolor2[362]&LFSRcolor2[12]);
    BiasedRNG[620] = (LFSRcolor2[350]&LFSRcolor2[424]&LFSRcolor2[176]);
    BiasedRNG[621] = (LFSRcolor2[756]&LFSRcolor2[737]&LFSRcolor2[692]);
    BiasedRNG[622] = (LFSRcolor2[205]&LFSRcolor2[649]&LFSRcolor2[485]);
    BiasedRNG[623] = (LFSRcolor2[586]&LFSRcolor2[486]&LFSRcolor2[204]);
    BiasedRNG[624] = (LFSRcolor2[86]&LFSRcolor2[471]&LFSRcolor2[68]);
    BiasedRNG[625] = (LFSRcolor2[611]&LFSRcolor2[105]&LFSRcolor2[608]);
    BiasedRNG[626] = (LFSRcolor2[199]&LFSRcolor2[340]&LFSRcolor2[3]);
    BiasedRNG[627] = (LFSRcolor2[296]&LFSRcolor2[426]&LFSRcolor2[646]);
    BiasedRNG[628] = (LFSRcolor2[690]&LFSRcolor2[575]&LFSRcolor2[272]);
    BiasedRNG[629] = (LFSRcolor2[196]&LFSRcolor2[241]&LFSRcolor2[239]);
    BiasedRNG[630] = (LFSRcolor2[494]&LFSRcolor2[214]&LFSRcolor2[95]);
    BiasedRNG[631] = (LFSRcolor2[568]&LFSRcolor2[200]&LFSRcolor2[689]);
    BiasedRNG[632] = (LFSRcolor2[255]&LFSRcolor2[365]&LFSRcolor2[592]);
    BiasedRNG[633] = (LFSRcolor2[736]&LFSRcolor2[280]&LFSRcolor2[641]);
    BiasedRNG[634] = (LFSRcolor2[281]&LFSRcolor2[314]&LFSRcolor2[308]);
    BiasedRNG[635] = (LFSRcolor2[530]&LFSRcolor2[338]&LFSRcolor2[381]);
    BiasedRNG[636] = (LFSRcolor2[273]&LFSRcolor2[570]&LFSRcolor2[253]);
    BiasedRNG[637] = (LFSRcolor2[89]&LFSRcolor2[738]&LFSRcolor2[144]);
    BiasedRNG[638] = (LFSRcolor2[187]&LFSRcolor2[711]&LFSRcolor2[283]);
    BiasedRNG[639] = (LFSRcolor2[125]&LFSRcolor2[154]&LFSRcolor2[444]);
    BiasedRNG[640] = (LFSRcolor2[158]&LFSRcolor2[388]&LFSRcolor2[22]);
    BiasedRNG[641] = (LFSRcolor2[130]&LFSRcolor2[713]&LFSRcolor2[35]);
    BiasedRNG[642] = (LFSRcolor2[520]&LFSRcolor2[317]&LFSRcolor2[382]);
    BiasedRNG[643] = (LFSRcolor2[10]&LFSRcolor2[702]&LFSRcolor2[775]);
    BiasedRNG[644] = (LFSRcolor2[19]&LFSRcolor2[668]&LFSRcolor2[14]);
    BiasedRNG[645] = (LFSRcolor2[61]&LFSRcolor2[626]&LFSRcolor2[618]);
    BiasedRNG[646] = (LFSRcolor2[116]&LFSRcolor2[563]&LFSRcolor2[282]);
    BiasedRNG[647] = (LFSRcolor2[168]&LFSRcolor2[71]&LFSRcolor2[474]);
    BiasedRNG[648] = (LFSRcolor2[451]&LFSRcolor2[431]&LFSRcolor2[57]);
    BiasedRNG[649] = (LFSRcolor2[265]&LFSRcolor2[374]&LFSRcolor2[660]);
    BiasedRNG[650] = (LFSRcolor2[323]&LFSRcolor2[249]&LFSRcolor2[294]);
    BiasedRNG[651] = (LFSRcolor2[696]&LFSRcolor2[581]&LFSRcolor2[769]);
    BiasedRNG[652] = (LFSRcolor2[434]&LFSRcolor2[397]&LFSRcolor2[93]);
    BiasedRNG[653] = (LFSRcolor2[15]&LFSRcolor2[617]&LFSRcolor2[654]);
    BiasedRNG[654] = (LFSRcolor2[652]&LFSRcolor2[192]&LFSRcolor2[546]);
    BiasedRNG[655] = (LFSRcolor2[120]&LFSRcolor2[466]&LFSRcolor2[392]);
    BiasedRNG[656] = (LFSRcolor2[49]&LFSRcolor2[230]&LFSRcolor2[554]);
    BiasedRNG[657] = (LFSRcolor2[182]&LFSRcolor2[644]&LFSRcolor2[700]);
    BiasedRNG[658] = (LFSRcolor2[510]&LFSRcolor2[609]&LFSRcolor2[377]);
    BiasedRNG[659] = (LFSRcolor2[221]&LFSRcolor2[542]&LFSRcolor2[427]);
    BiasedRNG[660] = (LFSRcolor2[145]&LFSRcolor2[48]&LFSRcolor2[428]);
    BiasedRNG[661] = (LFSRcolor2[261]&LFSRcolor2[1]&LFSRcolor2[31]);
    BiasedRNG[662] = (LFSRcolor2[378]&LFSRcolor2[264]&LFSRcolor2[774]);
    BiasedRNG[663] = (LFSRcolor2[371]&LFSRcolor2[577]&LFSRcolor2[343]);
    BiasedRNG[664] = (LFSRcolor2[493]&LFSRcolor2[297]&LFSRcolor2[610]);
    BiasedRNG[665] = (LFSRcolor2[329]&LFSRcolor2[159]&LFSRcolor2[529]);
    BiasedRNG[666] = (LFSRcolor2[108]&LFSRcolor2[703]&LFSRcolor2[506]);
    BiasedRNG[667] = (LFSRcolor2[439]&LFSRcolor2[209]&LFSRcolor2[274]);
    BiasedRNG[668] = (LFSRcolor2[672]&LFSRcolor2[306]&LFSRcolor2[415]);
    BiasedRNG[669] = (LFSRcolor2[53]&LFSRcolor2[754]&LFSRcolor2[669]);
    BiasedRNG[670] = (LFSRcolor2[763]&LFSRcolor2[164]&LFSRcolor2[634]);
    BiasedRNG[671] = (LFSRcolor2[27]&LFSRcolor2[683]&LFSRcolor2[443]);
    BiasedRNG[672] = (LFSRcolor2[487]&LFSRcolor2[492]&LFSRcolor2[99]);
    BiasedRNG[673] = (LFSRcolor2[185]&LFSRcolor2[405]&LFSRcolor2[111]);
    BiasedRNG[674] = (LFSRcolor2[277]&LFSRcolor2[685]&LFSRcolor2[387]);
    BiasedRNG[675] = (LFSRcolor2[566]&LFSRcolor2[732]&LFSRcolor2[400]);
    BiasedRNG[676] = (LFSRcolor2[759]&LFSRcolor2[36]&LFSRcolor2[670]);
    BiasedRNG[677] = (LFSRcolor2[694]&LFSRcolor2[212]&LFSRcolor2[403]);
    BiasedRNG[678] = (LFSRcolor2[260]&LFSRcolor2[42]&LFSRcolor2[523]);
    BiasedRNG[679] = (LFSRcolor2[56]&LFSRcolor2[118]&LFSRcolor2[368]);
    BiasedRNG[680] = (LFSRcolor2[655]&LFSRcolor2[278]&LFSRcolor2[573]);
    BiasedRNG[681] = (LFSRcolor2[240]&LFSRcolor2[688]&LFSRcolor2[622]);
    BiasedRNG[682] = (LFSRcolor2[210]&LFSRcolor2[429]&LFSRcolor2[279]);
    BiasedRNG[683] = (LFSRcolor2[747]&LFSRcolor2[220]&LFSRcolor2[103]);
    BiasedRNG[684] = (LFSRcolor2[579]&LFSRcolor2[355]&LFSRcolor2[478]);
    BiasedRNG[685] = (LFSRcolor2[157]&LFSRcolor2[112]&LFSRcolor2[687]);
    BiasedRNG[686] = (LFSRcolor2[254]&LFSRcolor2[535]&LFSRcolor2[207]);
    BiasedRNG[687] = (LFSRcolor2[398]&LFSRcolor2[532]&LFSRcolor2[547]);
    BiasedRNG[688] = (LFSRcolor2[132]&LFSRcolor2[248]&LFSRcolor2[751]);
    BiasedRNG[689] = (LFSRcolor2[117]&LFSRcolor2[718]&LFSRcolor2[271]);
    BiasedRNG[690] = (LFSRcolor2[364]&LFSRcolor2[704]&LFSRcolor2[663]);
    BiasedRNG[691] = (LFSRcolor2[229]&LFSRcolor2[332]&LFSRcolor2[246]);
    BiasedRNG[692] = (LFSRcolor2[457]&LFSRcolor2[777]&LFSRcolor2[295]);
    BiasedRNG[693] = (LFSRcolor2[162]&LFSRcolor2[353]&LFSRcolor2[213]);
    BiasedRNG[694] = (LFSRcolor2[545]&LFSRcolor2[714]&LFSRcolor2[134]);
    BiasedRNG[695] = (LFSRcolor2[224]&LFSRcolor2[0]&LFSRcolor2[464]);
    BiasedRNG[696] = (LFSRcolor2[594]&LFSRcolor2[658]&LFSRcolor2[414]);
    BiasedRNG[697] = (LFSRcolor2[325]&LFSRcolor2[724]&LFSRcolor2[259]);
    BiasedRNG[698] = (LFSRcolor2[165]&LFSRcolor2[73]&LFSRcolor2[619]);
    UnbiasedRNG[386] = LFSRcolor2[24];
    UnbiasedRNG[387] = LFSRcolor2[552];
    UnbiasedRNG[388] = LFSRcolor2[389];
    UnbiasedRNG[389] = LFSRcolor2[508];
    UnbiasedRNG[390] = LFSRcolor2[17];
    UnbiasedRNG[391] = LFSRcolor2[155];
    UnbiasedRNG[392] = LFSRcolor2[722];
    UnbiasedRNG[393] = LFSRcolor2[367];
    UnbiasedRNG[394] = LFSRcolor2[544];
    UnbiasedRNG[395] = LFSRcolor2[500];
    UnbiasedRNG[396] = LFSRcolor2[335];
    UnbiasedRNG[397] = LFSRcolor2[287];
    UnbiasedRNG[398] = LFSRcolor2[757];
    UnbiasedRNG[399] = LFSRcolor2[34];
    UnbiasedRNG[400] = LFSRcolor2[483];
    UnbiasedRNG[401] = LFSRcolor2[244];
    UnbiasedRNG[402] = LFSRcolor2[262];
    UnbiasedRNG[403] = LFSRcolor2[693];
    UnbiasedRNG[404] = LFSRcolor2[615];
    UnbiasedRNG[405] = LFSRcolor2[290];
    UnbiasedRNG[406] = LFSRcolor2[16];
    UnbiasedRNG[407] = LFSRcolor2[411];
    UnbiasedRNG[408] = LFSRcolor2[18];
    UnbiasedRNG[409] = LFSRcolor2[505];
    UnbiasedRNG[410] = LFSRcolor2[100];
    UnbiasedRNG[411] = LFSRcolor2[488];
    UnbiasedRNG[412] = LFSRcolor2[91];
    UnbiasedRNG[413] = LFSRcolor2[528];
    UnbiasedRNG[414] = LFSRcolor2[440];
    UnbiasedRNG[415] = LFSRcolor2[558];
    UnbiasedRNG[416] = LFSRcolor2[504];
    UnbiasedRNG[417] = LFSRcolor2[189];
    UnbiasedRNG[418] = LFSRcolor2[393];
    UnbiasedRNG[419] = LFSRcolor2[231];
    UnbiasedRNG[420] = LFSRcolor2[479];
    UnbiasedRNG[421] = LFSRcolor2[441];
    UnbiasedRNG[422] = LFSRcolor2[408];
    UnbiasedRNG[423] = LFSRcolor2[407];
    UnbiasedRNG[424] = LFSRcolor2[385];
    UnbiasedRNG[425] = LFSRcolor2[432];
    UnbiasedRNG[426] = LFSRcolor2[23];
    UnbiasedRNG[427] = LFSRcolor2[593];
    UnbiasedRNG[428] = LFSRcolor2[195];
    UnbiasedRNG[429] = LFSRcolor2[430];
    UnbiasedRNG[430] = LFSRcolor2[503];
    UnbiasedRNG[431] = LFSRcolor2[351];
    UnbiasedRNG[432] = LFSRcolor2[79];
    UnbiasedRNG[433] = LFSRcolor2[347];
    UnbiasedRNG[434] = LFSRcolor2[250];
    UnbiasedRNG[435] = LFSRcolor2[648];
    UnbiasedRNG[436] = LFSRcolor2[357];
    UnbiasedRNG[437] = LFSRcolor2[604];
    UnbiasedRNG[438] = LFSRcolor2[304];
    UnbiasedRNG[439] = LFSRcolor2[762];
    UnbiasedRNG[440] = LFSRcolor2[289];
    UnbiasedRNG[441] = LFSRcolor2[359];
    UnbiasedRNG[442] = LFSRcolor2[625];
    UnbiasedRNG[443] = LFSRcolor2[67];
    UnbiasedRNG[444] = LFSRcolor2[312];
    UnbiasedRNG[445] = LFSRcolor2[131];
    UnbiasedRNG[446] = LFSRcolor2[768];
    UnbiasedRNG[447] = LFSRcolor2[336];
    UnbiasedRNG[448] = LFSRcolor2[423];
    UnbiasedRNG[449] = LFSRcolor2[315];
    UnbiasedRNG[450] = LFSRcolor2[522];
    UnbiasedRNG[451] = LFSRcolor2[612];
    UnbiasedRNG[452] = LFSRcolor2[710];
    UnbiasedRNG[453] = LFSRcolor2[567];
    UnbiasedRNG[454] = LFSRcolor2[695];
    UnbiasedRNG[455] = LFSRcolor2[496];
    UnbiasedRNG[456] = LFSRcolor2[32];
    UnbiasedRNG[457] = LFSRcolor2[595];
    UnbiasedRNG[458] = LFSRcolor2[460];
    UnbiasedRNG[459] = LFSRcolor2[266];
    UnbiasedRNG[460] = LFSRcolor2[4];
    UnbiasedRNG[461] = LFSRcolor2[85];
    UnbiasedRNG[462] = LFSRcolor2[461];
    UnbiasedRNG[463] = LFSRcolor2[745];
    UnbiasedRNG[464] = LFSRcolor2[328];
    UnbiasedRNG[465] = LFSRcolor2[352];
    UnbiasedRNG[466] = LFSRcolor2[515];
    UnbiasedRNG[467] = LFSRcolor2[292];
    UnbiasedRNG[468] = LFSRcolor2[184];
    UnbiasedRNG[469] = LFSRcolor2[780];
    UnbiasedRNG[470] = LFSRcolor2[588];
    UnbiasedRNG[471] = LFSRcolor2[436];
    UnbiasedRNG[472] = LFSRcolor2[193];
    UnbiasedRNG[473] = LFSRcolor2[680];
    UnbiasedRNG[474] = LFSRcolor2[258];
    UnbiasedRNG[475] = LFSRcolor2[557];
    UnbiasedRNG[476] = LFSRcolor2[524];
    UnbiasedRNG[477] = LFSRcolor2[727];
    UnbiasedRNG[478] = LFSRcolor2[489];
    UnbiasedRNG[479] = LFSRcolor2[119];
    UnbiasedRNG[480] = LFSRcolor2[675];
    UnbiasedRNG[481] = LFSRcolor2[516];
    UnbiasedRNG[482] = LFSRcolor2[676];
    UnbiasedRNG[483] = LFSRcolor2[531];
    UnbiasedRNG[484] = LFSRcolor2[764];
    UnbiasedRNG[485] = LFSRcolor2[39];
    UnbiasedRNG[486] = LFSRcolor2[721];
    UnbiasedRNG[487] = LFSRcolor2[574];
    UnbiasedRNG[488] = LFSRcolor2[55];
    UnbiasedRNG[489] = LFSRcolor2[560];
    UnbiasedRNG[490] = LFSRcolor2[584];
    UnbiasedRNG[491] = LFSRcolor2[291];
    UnbiasedRNG[492] = LFSRcolor2[190];
    UnbiasedRNG[493] = LFSRcolor2[51];
    UnbiasedRNG[494] = LFSRcolor2[128];
    UnbiasedRNG[495] = LFSRcolor2[495];
    UnbiasedRNG[496] = LFSRcolor2[765];
    UnbiasedRNG[497] = LFSRcolor2[50];
    UnbiasedRNG[498] = LFSRcolor2[123];
    UnbiasedRNG[499] = LFSRcolor2[139];
    UnbiasedRNG[500] = LFSRcolor2[674];
    UnbiasedRNG[501] = LFSRcolor2[698];
    UnbiasedRNG[502] = LFSRcolor2[63];
    UnbiasedRNG[503] = LFSRcolor2[527];
    UnbiasedRNG[504] = LFSRcolor2[614];
    UnbiasedRNG[505] = LFSRcolor2[90];
    UnbiasedRNG[506] = LFSRcolor2[628];
    UnbiasedRNG[507] = LFSRcolor2[561];
    UnbiasedRNG[508] = LFSRcolor2[743];
    UnbiasedRNG[509] = LFSRcolor2[373];
    UnbiasedRNG[510] = LFSRcolor2[136];
    UnbiasedRNG[511] = LFSRcolor2[659];
    UnbiasedRNG[512] = LFSRcolor2[186];
    UnbiasedRNG[513] = LFSRcolor2[502];
    UnbiasedRNG[514] = LFSRcolor2[635];
    UnbiasedRNG[515] = LFSRcolor2[453];
    UnbiasedRNG[516] = LFSRcolor2[417];
    UnbiasedRNG[517] = LFSRcolor2[399];
    UnbiasedRNG[518] = LFSRcolor2[726];
    UnbiasedRNG[519] = LFSRcolor2[149];
    UnbiasedRNG[520] = LFSRcolor2[201];
    UnbiasedRNG[521] = LFSRcolor2[645];
    UnbiasedRNG[522] = LFSRcolor2[322];
    UnbiasedRNG[523] = LFSRcolor2[363];
    UnbiasedRNG[524] = LFSRcolor2[37];
    UnbiasedRNG[525] = LFSRcolor2[384];
    UnbiasedRNG[526] = LFSRcolor2[708];
    UnbiasedRNG[527] = LFSRcolor2[9];
    UnbiasedRNG[528] = LFSRcolor2[463];
    UnbiasedRNG[529] = LFSRcolor2[445];
    UnbiasedRNG[530] = LFSRcolor2[621];
    UnbiasedRNG[531] = LFSRcolor2[82];
    UnbiasedRNG[532] = LFSRcolor2[599];
    UnbiasedRNG[533] = LFSRcolor2[142];
    UnbiasedRNG[534] = LFSRcolor2[345];
    UnbiasedRNG[535] = LFSRcolor2[391];
    UnbiasedRNG[536] = LFSRcolor2[337];
    UnbiasedRNG[537] = LFSRcolor2[715];
    UnbiasedRNG[538] = LFSRcolor2[141];
    UnbiasedRNG[539] = LFSRcolor2[555];
    UnbiasedRNG[540] = LFSRcolor2[664];
    UnbiasedRNG[541] = LFSRcolor2[716];
    UnbiasedRNG[542] = LFSRcolor2[174];
    UnbiasedRNG[543] = LFSRcolor2[170];
    UnbiasedRNG[544] = LFSRcolor2[98];
    UnbiasedRNG[545] = LFSRcolor2[87];
    UnbiasedRNG[546] = LFSRcolor2[146];
    UnbiasedRNG[547] = LFSRcolor2[226];
    UnbiasedRNG[548] = LFSRcolor2[147];
    UnbiasedRNG[549] = LFSRcolor2[771];
    UnbiasedRNG[550] = LFSRcolor2[678];
    UnbiasedRNG[551] = LFSRcolor2[45];
    UnbiasedRNG[552] = LFSRcolor2[298];
    UnbiasedRNG[553] = LFSRcolor2[490];
    UnbiasedRNG[554] = LFSRcolor2[180];
    UnbiasedRNG[555] = LFSRcolor2[624];
    UnbiasedRNG[556] = LFSRcolor2[701];
    UnbiasedRNG[557] = LFSRcolor2[217];
    UnbiasedRNG[558] = LFSRcolor2[650];
    UnbiasedRNG[559] = LFSRcolor2[548];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[560] = LFSRcolor3[120];
    UnbiasedRNG[561] = LFSRcolor3[25];
    UnbiasedRNG[562] = LFSRcolor3[108];
    UnbiasedRNG[563] = LFSRcolor3[117];
    UnbiasedRNG[564] = LFSRcolor3[74];
    UnbiasedRNG[565] = LFSRcolor3[15];
    UnbiasedRNG[566] = LFSRcolor3[166];
    UnbiasedRNG[567] = LFSRcolor3[111];
    UnbiasedRNG[568] = LFSRcolor3[107];
    UnbiasedRNG[569] = LFSRcolor3[100];
    UnbiasedRNG[570] = LFSRcolor3[142];
    UnbiasedRNG[571] = LFSRcolor3[4];
    UnbiasedRNG[572] = LFSRcolor3[36];
    UnbiasedRNG[573] = LFSRcolor3[69];
    UnbiasedRNG[574] = LFSRcolor3[57];
    UnbiasedRNG[575] = LFSRcolor3[102];
    UnbiasedRNG[576] = LFSRcolor3[132];
    UnbiasedRNG[577] = LFSRcolor3[130];
    UnbiasedRNG[578] = LFSRcolor3[32];
    UnbiasedRNG[579] = LFSRcolor3[165];
    UnbiasedRNG[580] = LFSRcolor3[9];
    UnbiasedRNG[581] = LFSRcolor3[115];
    UnbiasedRNG[582] = LFSRcolor3[180];
    UnbiasedRNG[583] = LFSRcolor3[162];
    UnbiasedRNG[584] = LFSRcolor3[126];
    UnbiasedRNG[585] = LFSRcolor3[122];
    UnbiasedRNG[586] = LFSRcolor3[119];
    UnbiasedRNG[587] = LFSRcolor3[138];
    UnbiasedRNG[588] = LFSRcolor3[152];
    UnbiasedRNG[589] = LFSRcolor3[45];
    UnbiasedRNG[590] = LFSRcolor3[72];
    UnbiasedRNG[591] = LFSRcolor3[154];
    UnbiasedRNG[592] = LFSRcolor3[164];
    UnbiasedRNG[593] = LFSRcolor3[134];
    UnbiasedRNG[594] = LFSRcolor3[77];
    UnbiasedRNG[595] = LFSRcolor3[63];
    UnbiasedRNG[596] = LFSRcolor3[68];
    UnbiasedRNG[597] = LFSRcolor3[66];
    UnbiasedRNG[598] = LFSRcolor3[1];
    UnbiasedRNG[599] = LFSRcolor3[73];
    UnbiasedRNG[600] = LFSRcolor3[96];
    UnbiasedRNG[601] = LFSRcolor3[136];
    UnbiasedRNG[602] = LFSRcolor3[92];
    UnbiasedRNG[603] = LFSRcolor3[150];
    UnbiasedRNG[604] = LFSRcolor3[146];
    UnbiasedRNG[605] = LFSRcolor3[159];
    UnbiasedRNG[606] = LFSRcolor3[26];
    UnbiasedRNG[607] = LFSRcolor3[99];
    UnbiasedRNG[608] = LFSRcolor3[106];
    UnbiasedRNG[609] = LFSRcolor3[118];
    UnbiasedRNG[610] = LFSRcolor3[13];
    UnbiasedRNG[611] = LFSRcolor3[11];
    UnbiasedRNG[612] = LFSRcolor3[71];
    UnbiasedRNG[613] = LFSRcolor3[116];
    UnbiasedRNG[614] = LFSRcolor3[80];
    UnbiasedRNG[615] = LFSRcolor3[10];
    UnbiasedRNG[616] = LFSRcolor3[85];
    UnbiasedRNG[617] = LFSRcolor3[113];
    UnbiasedRNG[618] = LFSRcolor3[82];
    UnbiasedRNG[619] = LFSRcolor3[176];
    UnbiasedRNG[620] = LFSRcolor3[88];
    UnbiasedRNG[621] = LFSRcolor3[40];
    UnbiasedRNG[622] = LFSRcolor3[61];
    UnbiasedRNG[623] = LFSRcolor3[67];
    UnbiasedRNG[624] = LFSRcolor3[42];
    UnbiasedRNG[625] = LFSRcolor3[5];
    UnbiasedRNG[626] = LFSRcolor3[149];
    UnbiasedRNG[627] = LFSRcolor3[14];
    UnbiasedRNG[628] = LFSRcolor3[30];
    UnbiasedRNG[629] = LFSRcolor3[75];
    UnbiasedRNG[630] = LFSRcolor3[163];
    UnbiasedRNG[631] = LFSRcolor3[112];
    UnbiasedRNG[632] = LFSRcolor3[94];
    UnbiasedRNG[633] = LFSRcolor3[151];
    UnbiasedRNG[634] = LFSRcolor3[27];
    UnbiasedRNG[635] = LFSRcolor3[17];
    UnbiasedRNG[636] = LFSRcolor3[34];
    UnbiasedRNG[637] = LFSRcolor3[33];
    UnbiasedRNG[638] = LFSRcolor3[167];
    UnbiasedRNG[639] = LFSRcolor3[181];
    UnbiasedRNG[640] = LFSRcolor3[177];
    UnbiasedRNG[641] = LFSRcolor3[64];
    UnbiasedRNG[642] = LFSRcolor3[62];
    UnbiasedRNG[643] = LFSRcolor3[83];
    UnbiasedRNG[644] = LFSRcolor3[78];
    UnbiasedRNG[645] = LFSRcolor3[21];
    UnbiasedRNG[646] = LFSRcolor3[12];
    UnbiasedRNG[647] = LFSRcolor3[147];
    UnbiasedRNG[648] = LFSRcolor3[49];
    UnbiasedRNG[649] = LFSRcolor3[29];
    UnbiasedRNG[650] = LFSRcolor3[133];
    UnbiasedRNG[651] = LFSRcolor3[125];
    UnbiasedRNG[652] = LFSRcolor3[182];
    UnbiasedRNG[653] = LFSRcolor3[56];
    UnbiasedRNG[654] = LFSRcolor3[139];
    UnbiasedRNG[655] = LFSRcolor3[178];
    UnbiasedRNG[656] = LFSRcolor3[38];
    UnbiasedRNG[657] = LFSRcolor3[31];
    UnbiasedRNG[658] = LFSRcolor3[103];
    UnbiasedRNG[659] = LFSRcolor3[141];
    UnbiasedRNG[660] = LFSRcolor3[161];
    UnbiasedRNG[661] = LFSRcolor3[46];
    UnbiasedRNG[662] = LFSRcolor3[175];
    UnbiasedRNG[663] = LFSRcolor3[86];
    UnbiasedRNG[664] = LFSRcolor3[3];
    UnbiasedRNG[665] = LFSRcolor3[24];
    UnbiasedRNG[666] = LFSRcolor3[109];
    UnbiasedRNG[667] = LFSRcolor3[140];
    UnbiasedRNG[668] = LFSRcolor3[173];
    UnbiasedRNG[669] = LFSRcolor3[168];
    UnbiasedRNG[670] = LFSRcolor3[90];
    UnbiasedRNG[671] = LFSRcolor3[59];
    UnbiasedRNG[672] = LFSRcolor3[172];
    UnbiasedRNG[673] = LFSRcolor3[114];
    UnbiasedRNG[674] = LFSRcolor3[121];
    UnbiasedRNG[675] = LFSRcolor3[160];
    UnbiasedRNG[676] = LFSRcolor3[47];
    UnbiasedRNG[677] = LFSRcolor3[48];
    UnbiasedRNG[678] = LFSRcolor3[97];
    UnbiasedRNG[679] = LFSRcolor3[7];
    UnbiasedRNG[680] = LFSRcolor3[81];
    UnbiasedRNG[681] = LFSRcolor3[44];
    UnbiasedRNG[682] = LFSRcolor3[135];
    UnbiasedRNG[683] = LFSRcolor3[144];
    UnbiasedRNG[684] = LFSRcolor3[6];
    UnbiasedRNG[685] = LFSRcolor3[98];
    UnbiasedRNG[686] = LFSRcolor3[110];
    UnbiasedRNG[687] = LFSRcolor3[79];
    UnbiasedRNG[688] = LFSRcolor3[91];
    UnbiasedRNG[689] = LFSRcolor3[2];
    UnbiasedRNG[690] = LFSRcolor3[89];
    UnbiasedRNG[691] = LFSRcolor3[18];
    UnbiasedRNG[692] = LFSRcolor3[22];
    UnbiasedRNG[693] = LFSRcolor3[95];
    UnbiasedRNG[694] = LFSRcolor3[35];
    UnbiasedRNG[695] = LFSRcolor3[16];
    UnbiasedRNG[696] = LFSRcolor3[127];
    UnbiasedRNG[697] = LFSRcolor3[37];
    UnbiasedRNG[698] = LFSRcolor3[70];
    UnbiasedRNG[699] = LFSRcolor3[65];
    UnbiasedRNG[700] = LFSRcolor3[0];
    UnbiasedRNG[701] = LFSRcolor3[148];
    UnbiasedRNG[702] = LFSRcolor3[104];
    UnbiasedRNG[703] = LFSRcolor3[155];
    UnbiasedRNG[704] = LFSRcolor3[174];
    UnbiasedRNG[705] = LFSRcolor3[87];
    UnbiasedRNG[706] = LFSRcolor3[19];
    UnbiasedRNG[707] = LFSRcolor3[153];
    UnbiasedRNG[708] = LFSRcolor3[145];
    UnbiasedRNG[709] = LFSRcolor3[53];
    UnbiasedRNG[710] = LFSRcolor3[84];
    UnbiasedRNG[711] = LFSRcolor3[124];
    UnbiasedRNG[712] = LFSRcolor3[8];
    UnbiasedRNG[713] = LFSRcolor3[23];
    UnbiasedRNG[714] = LFSRcolor3[183];
    UnbiasedRNG[715] = LFSRcolor3[52];
end

always @(posedge color3_clk) begin
    BiasedRNG[699] = (LFSRcolor4[184]&LFSRcolor4[185]&LFSRcolor4[428]);
    BiasedRNG[700] = (LFSRcolor4[113]&LFSRcolor4[255]&LFSRcolor4[158]);
    BiasedRNG[701] = (LFSRcolor4[253]&LFSRcolor4[267]&LFSRcolor4[340]);
    BiasedRNG[702] = (LFSRcolor4[476]&LFSRcolor4[94]&LFSRcolor4[529]);
    BiasedRNG[703] = (LFSRcolor4[522]&LFSRcolor4[139]&LFSRcolor4[22]);
    BiasedRNG[704] = (LFSRcolor4[426]&LFSRcolor4[242]&LFSRcolor4[485]);
    BiasedRNG[705] = (LFSRcolor4[226]&LFSRcolor4[145]&LFSRcolor4[373]);
    BiasedRNG[706] = (LFSRcolor4[164]&LFSRcolor4[260]&LFSRcolor4[236]);
    BiasedRNG[707] = (LFSRcolor4[111]&LFSRcolor4[30]&LFSRcolor4[179]);
    BiasedRNG[708] = (LFSRcolor4[76]&LFSRcolor4[292]&LFSRcolor4[17]);
    BiasedRNG[709] = (LFSRcolor4[535]&LFSRcolor4[460]&LFSRcolor4[382]);
    BiasedRNG[710] = (LFSRcolor4[157]&LFSRcolor4[237]&LFSRcolor4[11]);
    BiasedRNG[711] = (LFSRcolor4[73]&LFSRcolor4[490]&LFSRcolor4[310]);
    BiasedRNG[712] = (LFSRcolor4[296]&LFSRcolor4[8]&LFSRcolor4[399]);
    BiasedRNG[713] = (LFSRcolor4[534]&LFSRcolor4[265]&LFSRcolor4[539]);
    BiasedRNG[714] = (LFSRcolor4[50]&LFSRcolor4[216]&LFSRcolor4[286]);
    BiasedRNG[715] = (LFSRcolor4[304]&LFSRcolor4[154]&LFSRcolor4[104]);
    BiasedRNG[716] = (LFSRcolor4[225]&LFSRcolor4[177]&LFSRcolor4[72]);
    BiasedRNG[717] = (LFSRcolor4[427]&LFSRcolor4[152]&LFSRcolor4[109]);
    BiasedRNG[718] = (LFSRcolor4[454]&LFSRcolor4[189]&LFSRcolor4[147]);
    BiasedRNG[719] = (LFSRcolor4[506]&LFSRcolor4[429]&LFSRcolor4[256]);
    BiasedRNG[720] = (LFSRcolor4[53]&LFSRcolor4[354]&LFSRcolor4[339]);
    BiasedRNG[721] = (LFSRcolor4[335]&LFSRcolor4[295]&LFSRcolor4[209]);
    BiasedRNG[722] = (LFSRcolor4[264]&LFSRcolor4[180]&LFSRcolor4[401]);
    BiasedRNG[723] = (LFSRcolor4[370]&LFSRcolor4[488]&LFSRcolor4[257]);
    BiasedRNG[724] = (LFSRcolor4[252]&LFSRcolor4[379]&LFSRcolor4[368]);
    BiasedRNG[725] = (LFSRcolor4[144]&LFSRcolor4[176]&LFSRcolor4[510]);
    BiasedRNG[726] = (LFSRcolor4[26]&LFSRcolor4[375]&LFSRcolor4[538]);
    BiasedRNG[727] = (LFSRcolor4[308]&LFSRcolor4[19]&LFSRcolor4[376]);
    BiasedRNG[728] = (LFSRcolor4[526]&LFSRcolor4[270]&LFSRcolor4[150]);
    BiasedRNG[729] = (LFSRcolor4[407]&LFSRcolor4[80]&LFSRcolor4[352]);
    BiasedRNG[730] = (LFSRcolor4[505]&LFSRcolor4[239]&LFSRcolor4[462]);
    BiasedRNG[731] = (LFSRcolor4[381]&LFSRcolor4[168]&LFSRcolor4[56]);
    BiasedRNG[732] = (LFSRcolor4[475]&LFSRcolor4[112]&LFSRcolor4[481]);
    BiasedRNG[733] = (LFSRcolor4[108]&LFSRcolor4[298]&LFSRcolor4[521]);
    BiasedRNG[734] = (LFSRcolor4[213]&LFSRcolor4[437]&LFSRcolor4[142]);
    BiasedRNG[735] = (LFSRcolor4[120]&LFSRcolor4[291]&LFSRcolor4[330]);
    BiasedRNG[736] = (LFSRcolor4[227]&LFSRcolor4[272]&LFSRcolor4[230]);
    BiasedRNG[737] = (LFSRcolor4[307]&LFSRcolor4[93]&LFSRcolor4[371]);
    BiasedRNG[738] = (LFSRcolor4[132]&LFSRcolor4[249]&LFSRcolor4[141]);
    BiasedRNG[739] = (LFSRcolor4[235]&LFSRcolor4[440]&LFSRcolor4[172]);
    BiasedRNG[740] = (LFSRcolor4[9]&LFSRcolor4[268]&LFSRcolor4[169]);
    BiasedRNG[741] = (LFSRcolor4[34]&LFSRcolor4[60]&LFSRcolor4[218]);
    BiasedRNG[742] = (LFSRcolor4[342]&LFSRcolor4[130]&LFSRcolor4[170]);
    BiasedRNG[743] = (LFSRcolor4[380]&LFSRcolor4[28]&LFSRcolor4[314]);
    BiasedRNG[744] = (LFSRcolor4[62]&LFSRcolor4[470]&LFSRcolor4[424]);
    BiasedRNG[745] = (LFSRcolor4[489]&LFSRcolor4[173]&LFSRcolor4[420]);
    BiasedRNG[746] = (LFSRcolor4[222]&LFSRcolor4[312]&LFSRcolor4[114]);
    BiasedRNG[747] = (LFSRcolor4[85]&LFSRcolor4[305]&LFSRcolor4[88]);
    BiasedRNG[748] = (LFSRcolor4[394]&LFSRcolor4[182]&LFSRcolor4[101]);
    BiasedRNG[749] = (LFSRcolor4[450]&LFSRcolor4[215]&LFSRcolor4[29]);
    BiasedRNG[750] = (LFSRcolor4[149]&LFSRcolor4[482]&LFSRcolor4[166]);
    BiasedRNG[751] = (LFSRcolor4[200]&LFSRcolor4[337]&LFSRcolor4[315]);
    BiasedRNG[752] = (LFSRcolor4[2]&LFSRcolor4[91]&LFSRcolor4[456]);
    BiasedRNG[753] = (LFSRcolor4[325]&LFSRcolor4[214]&LFSRcolor4[497]);
    BiasedRNG[754] = (LFSRcolor4[455]&LFSRcolor4[279]&LFSRcolor4[229]);
    BiasedRNG[755] = (LFSRcolor4[87]&LFSRcolor4[33]&LFSRcolor4[378]);
    BiasedRNG[756] = (LFSRcolor4[527]&LFSRcolor4[202]&LFSRcolor4[518]);
    BiasedRNG[757] = (LFSRcolor4[311]&LFSRcolor4[119]&LFSRcolor4[461]);
    BiasedRNG[758] = (LFSRcolor4[405]&LFSRcolor4[126]&LFSRcolor4[508]);
    BiasedRNG[759] = (LFSRcolor4[174]&LFSRcolor4[417]&LFSRcolor4[361]);
    BiasedRNG[760] = (LFSRcolor4[474]&LFSRcolor4[477]&LFSRcolor4[273]);
    BiasedRNG[761] = (LFSRcolor4[322]&LFSRcolor4[42]&LFSRcolor4[77]);
    BiasedRNG[762] = (LFSRcolor4[102]&LFSRcolor4[439]&LFSRcolor4[32]);
    BiasedRNG[763] = (LFSRcolor4[333]&LFSRcolor4[366]&LFSRcolor4[194]);
    BiasedRNG[764] = (LFSRcolor4[363]&LFSRcolor4[384]&LFSRcolor4[121]);
    BiasedRNG[765] = (LFSRcolor4[148]&LFSRcolor4[5]&LFSRcolor4[282]);
    BiasedRNG[766] = (LFSRcolor4[106]&LFSRcolor4[509]&LFSRcolor4[65]);
    BiasedRNG[767] = (LFSRcolor4[473]&LFSRcolor4[309]&LFSRcolor4[64]);
    BiasedRNG[768] = (LFSRcolor4[374]&LFSRcolor4[21]&LFSRcolor4[45]);
    BiasedRNG[769] = (LFSRcolor4[36]&LFSRcolor4[458]&LFSRcolor4[391]);
    BiasedRNG[770] = (LFSRcolor4[357]&LFSRcolor4[127]&LFSRcolor4[107]);
    BiasedRNG[771] = (LFSRcolor4[343]&LFSRcolor4[530]&LFSRcolor4[536]);
    BiasedRNG[772] = (LFSRcolor4[369]&LFSRcolor4[175]&LFSRcolor4[445]);
    BiasedRNG[773] = (LFSRcolor4[444]&LFSRcolor4[269]&LFSRcolor4[457]);
    BiasedRNG[774] = (LFSRcolor4[66]&LFSRcolor4[71]&LFSRcolor4[517]);
    BiasedRNG[775] = (LFSRcolor4[364]&LFSRcolor4[78]&LFSRcolor4[425]);
    BiasedRNG[776] = (LFSRcolor4[435]&LFSRcolor4[507]&LFSRcolor4[188]);
    BiasedRNG[777] = (LFSRcolor4[3]&LFSRcolor4[332]&LFSRcolor4[67]);
    BiasedRNG[778] = (LFSRcolor4[258]&LFSRcolor4[46]&LFSRcolor4[250]);
    BiasedRNG[779] = (LFSRcolor4[96]&LFSRcolor4[234]&LFSRcolor4[303]);
    BiasedRNG[780] = (LFSRcolor4[89]&LFSRcolor4[178]&LFSRcolor4[397]);
    BiasedRNG[781] = (LFSRcolor4[95]&LFSRcolor4[400]&LFSRcolor4[365]);
    BiasedRNG[782] = (LFSRcolor4[186]&LFSRcolor4[299]&LFSRcolor4[484]);
    BiasedRNG[783] = (LFSRcolor4[122]&LFSRcolor4[20]&LFSRcolor4[90]);
    BiasedRNG[784] = (LFSRcolor4[207]&LFSRcolor4[422]&LFSRcolor4[468]);
    BiasedRNG[785] = (LFSRcolor4[387]&LFSRcolor4[165]&LFSRcolor4[324]);
    BiasedRNG[786] = (LFSRcolor4[465]&LFSRcolor4[471]&LFSRcolor4[319]);
    BiasedRNG[787] = (LFSRcolor4[463]&LFSRcolor4[284]&LFSRcolor4[37]);
    BiasedRNG[788] = (LFSRcolor4[546]&LFSRcolor4[283]&LFSRcolor4[306]);
    BiasedRNG[789] = (LFSRcolor4[123]&LFSRcolor4[434]&LFSRcolor4[344]);
    BiasedRNG[790] = (LFSRcolor4[187]&LFSRcolor4[39]&LFSRcolor4[385]);
    BiasedRNG[791] = (LFSRcolor4[155]&LFSRcolor4[466]&LFSRcolor4[233]);
    BiasedRNG[792] = (LFSRcolor4[27]&LFSRcolor4[433]&LFSRcolor4[501]);
    BiasedRNG[793] = (LFSRcolor4[396]&LFSRcolor4[349]&LFSRcolor4[251]);
    BiasedRNG[794] = (LFSRcolor4[124]&LFSRcolor4[494]&LFSRcolor4[492]);
    BiasedRNG[795] = (LFSRcolor4[116]&LFSRcolor4[74]&LFSRcolor4[443]);
    BiasedRNG[796] = (LFSRcolor4[198]&LFSRcolor4[61]&LFSRcolor4[98]);
    BiasedRNG[797] = (LFSRcolor4[219]&LFSRcolor4[79]&LFSRcolor4[146]);
    BiasedRNG[798] = (LFSRcolor4[524]&LFSRcolor4[447]&LFSRcolor4[51]);
    BiasedRNG[799] = (LFSRcolor4[356]&LFSRcolor4[70]&LFSRcolor4[416]);
    BiasedRNG[800] = (LFSRcolor4[261]&LFSRcolor4[83]&LFSRcolor4[504]);
    BiasedRNG[801] = (LFSRcolor4[525]&LFSRcolor4[453]&LFSRcolor4[386]);
    BiasedRNG[802] = (LFSRcolor4[163]&LFSRcolor4[75]&LFSRcolor4[217]);
    BiasedRNG[803] = (LFSRcolor4[115]&LFSRcolor4[478]&LFSRcolor4[103]);
    BiasedRNG[804] = (LFSRcolor4[542]&LFSRcolor4[193]&LFSRcolor4[245]);
    BiasedRNG[805] = (LFSRcolor4[289]&LFSRcolor4[452]&LFSRcolor4[244]);
    BiasedRNG[806] = (LFSRcolor4[208]&LFSRcolor4[14]&LFSRcolor4[377]);
    BiasedRNG[807] = (LFSRcolor4[320]&LFSRcolor4[533]&LFSRcolor4[353]);
    BiasedRNG[808] = (LFSRcolor4[136]&LFSRcolor4[448]&LFSRcolor4[551]);
    BiasedRNG[809] = (LFSRcolor4[211]&LFSRcolor4[281]&LFSRcolor4[197]);
    BiasedRNG[810] = (LFSRcolor4[59]&LFSRcolor4[159]&LFSRcolor4[446]);
    BiasedRNG[811] = (LFSRcolor4[297]&LFSRcolor4[487]&LFSRcolor4[503]);
    BiasedRNG[812] = (LFSRcolor4[247]&LFSRcolor4[129]&LFSRcolor4[451]);
    BiasedRNG[813] = (LFSRcolor4[259]&LFSRcolor4[362]&LFSRcolor4[86]);
    BiasedRNG[814] = (LFSRcolor4[442]&LFSRcolor4[500]&LFSRcolor4[301]);
    BiasedRNG[815] = (LFSRcolor4[153]&LFSRcolor4[498]&LFSRcolor4[24]);
    BiasedRNG[816] = (LFSRcolor4[18]&LFSRcolor4[204]&LFSRcolor4[128]);
    BiasedRNG[817] = (LFSRcolor4[68]&LFSRcolor4[31]&LFSRcolor4[511]);
    BiasedRNG[818] = (LFSRcolor4[274]&LFSRcolor4[520]&LFSRcolor4[161]);
    BiasedRNG[819] = (LFSRcolor4[532]&LFSRcolor4[232]&LFSRcolor4[43]);
    BiasedRNG[820] = (LFSRcolor4[224]&LFSRcolor4[398]&LFSRcolor4[49]);
    BiasedRNG[821] = (LFSRcolor4[201]&LFSRcolor4[92]&LFSRcolor4[99]);
    BiasedRNG[822] = (LFSRcolor4[351]&LFSRcolor4[436]&LFSRcolor4[318]);
    BiasedRNG[823] = (LFSRcolor4[413]&LFSRcolor4[548]&LFSRcolor4[133]);
    BiasedRNG[824] = (LFSRcolor4[288]&LFSRcolor4[389]&LFSRcolor4[13]);
    BiasedRNG[825] = (LFSRcolor4[84]&LFSRcolor4[280]&LFSRcolor4[545]);
    BiasedRNG[826] = (LFSRcolor4[38]&LFSRcolor4[316]&LFSRcolor4[294]);
    BiasedRNG[827] = (LFSRcolor4[338]&LFSRcolor4[411]&LFSRcolor4[547]);
    BiasedRNG[828] = (LFSRcolor4[388]&LFSRcolor4[105]&LFSRcolor4[346]);
    BiasedRNG[829] = (LFSRcolor4[358]&LFSRcolor4[285]&LFSRcolor4[415]);
    BiasedRNG[830] = (LFSRcolor4[278]&LFSRcolor4[210]&LFSRcolor4[160]);
    BiasedRNG[831] = (LFSRcolor4[383]&LFSRcolor4[205]&LFSRcolor4[430]);
    BiasedRNG[832] = (LFSRcolor4[359]&LFSRcolor4[276]&LFSRcolor4[499]);
    BiasedRNG[833] = (LFSRcolor4[138]&LFSRcolor4[528]&LFSRcolor4[537]);
    BiasedRNG[834] = (LFSRcolor4[156]&LFSRcolor4[502]&LFSRcolor4[57]);
    BiasedRNG[835] = (LFSRcolor4[183]&LFSRcolor4[350]&LFSRcolor4[414]);
    BiasedRNG[836] = (LFSRcolor4[543]&LFSRcolor4[403]&LFSRcolor4[243]);
    BiasedRNG[837] = (LFSRcolor4[35]&LFSRcolor4[441]&LFSRcolor4[329]);
    BiasedRNG[838] = (LFSRcolor4[6]&LFSRcolor4[206]&LFSRcolor4[134]);
    BiasedRNG[839] = (LFSRcolor4[231]&LFSRcolor4[326]&LFSRcolor4[479]);
    BiasedRNG[840] = (LFSRcolor4[181]&LFSRcolor4[223]&LFSRcolor4[302]);
    BiasedRNG[841] = (LFSRcolor4[140]&LFSRcolor4[390]&LFSRcolor4[496]);
    BiasedRNG[842] = (LFSRcolor4[195]&LFSRcolor4[12]&LFSRcolor4[412]);
    BiasedRNG[843] = (LFSRcolor4[345]&LFSRcolor4[459]&LFSRcolor4[47]);
    BiasedRNG[844] = (LFSRcolor4[52]&LFSRcolor4[246]&LFSRcolor4[355]);
    BiasedRNG[845] = (LFSRcolor4[313]&LFSRcolor4[483]&LFSRcolor4[151]);
    BiasedRNG[846] = (LFSRcolor4[7]&LFSRcolor4[514]&LFSRcolor4[336]);
    BiasedRNG[847] = (LFSRcolor4[23]&LFSRcolor4[15]&LFSRcolor4[54]);
    BiasedRNG[848] = (LFSRcolor4[467]&LFSRcolor4[0]&LFSRcolor4[290]);
    BiasedRNG[849] = (LFSRcolor4[531]&LFSRcolor4[167]&LFSRcolor4[162]);
    BiasedRNG[850] = (LFSRcolor4[1]&LFSRcolor4[192]&LFSRcolor4[423]);
    BiasedRNG[851] = (LFSRcolor4[392]&LFSRcolor4[321]&LFSRcolor4[190]);
    BiasedRNG[852] = (LFSRcolor4[491]&LFSRcolor4[360]&LFSRcolor4[432]);
    BiasedRNG[853] = (LFSRcolor4[395]&LFSRcolor4[421]&LFSRcolor4[408]);
    BiasedRNG[854] = (LFSRcolor4[10]&LFSRcolor4[367]&LFSRcolor4[317]);
    BiasedRNG[855] = (LFSRcolor4[81]&LFSRcolor4[271]&LFSRcolor4[254]);
    BiasedRNG[856] = (LFSRcolor4[495]&LFSRcolor4[82]&LFSRcolor4[248]);
    BiasedRNG[857] = (LFSRcolor4[410]&LFSRcolor4[431]&LFSRcolor4[540]);
    BiasedRNG[858] = (LFSRcolor4[464]&LFSRcolor4[347]&LFSRcolor4[275]);
    BiasedRNG[859] = (LFSRcolor4[372]&LFSRcolor4[199]&LFSRcolor4[203]);
    BiasedRNG[860] = (LFSRcolor4[212]&LFSRcolor4[171]&LFSRcolor4[240]);
    BiasedRNG[861] = (LFSRcolor4[334]&LFSRcolor4[196]&LFSRcolor4[323]);
    BiasedRNG[862] = (LFSRcolor4[263]&LFSRcolor4[25]&LFSRcolor4[402]);
    BiasedRNG[863] = (LFSRcolor4[480]&LFSRcolor4[287]&LFSRcolor4[48]);
    BiasedRNG[864] = (LFSRcolor4[238]&LFSRcolor4[63]&LFSRcolor4[519]);
    BiasedRNG[865] = (LFSRcolor4[549]&LFSRcolor4[493]&LFSRcolor4[220]);
    BiasedRNG[866] = (LFSRcolor4[331]&LFSRcolor4[266]&LFSRcolor4[409]);
    BiasedRNG[867] = (LFSRcolor4[541]&LFSRcolor4[137]&LFSRcolor4[69]);
    BiasedRNG[868] = (LFSRcolor4[419]&LFSRcolor4[486]&LFSRcolor4[341]);
    BiasedRNG[869] = (LFSRcolor4[191]&LFSRcolor4[300]&LFSRcolor4[404]);
    BiasedRNG[870] = (LFSRcolor4[293]&LFSRcolor4[117]&LFSRcolor4[328]);
    BiasedRNG[871] = (LFSRcolor4[110]&LFSRcolor4[58]&LFSRcolor4[513]);
    BiasedRNG[872] = (LFSRcolor4[40]&LFSRcolor4[472]&LFSRcolor4[438]);
    BiasedRNG[873] = (LFSRcolor4[348]&LFSRcolor4[418]&LFSRcolor4[469]);
    BiasedRNG[874] = (LFSRcolor4[16]&LFSRcolor4[4]&LFSRcolor4[100]);
    BiasedRNG[875] = (LFSRcolor4[44]&LFSRcolor4[125]&LFSRcolor4[516]);
    BiasedRNG[876] = (LFSRcolor4[262]&LFSRcolor4[131]&LFSRcolor4[512]);
    BiasedRNG[877] = (LFSRcolor4[221]&LFSRcolor4[544]&LFSRcolor4[406]);
    BiasedRNG[878] = (LFSRcolor4[55]&LFSRcolor4[97]&LFSRcolor4[228]);
    BiasedRNG[879] = (LFSRcolor4[118]&LFSRcolor4[327]&LFSRcolor4[515]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

//Generate the ILA for data collection:
ila_0 ILAinst(.clk(sample_clk),.probe0(run),.probe1(solution_flag),.probe2(failure),.probe3(counter[37:0]));

//Instantiate VIO:
vio_0 VIOinst (.clk(sample_clk),.probe_out0(reset),.probe_out1(solution_set[27:0]));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule