//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [37:0] counter;
initial counter = 38'b0;
reg [31:0] solution;
reg [31:0] solution_check;
wire [31:0] solution_set;
initial solution_check = 32'b11101011101110010100001101010001;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
reg [0:2079] InitCond;
reg run;
wire [1333:0] LFSRcolor0;
wire [1793:0] LFSRcolor1;
wire [1287:0] LFSRcolor2;
wire [229:0] LFSRcolor3;
wire [965:0] LFSRcolor4;
reg [1133:0] BiasedRNG;       //For I=+/-1 cases
reg [945:0] UnbiasedRNG;   //For I=0 cases
reg [0:2127] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[672] = 1'b1;
initial m[931] = 1'b0;
initial m[941] = 1'b0;
initial m[956] = 1'b0;
initial m[976] = 1'b1;
initial m[1001] = 1'b0;
initial m[1031] = 1'b1;
initial m[1066] = 1'b0;
initial m[1106] = 1'b1;
initial m[1151] = 1'b1;
initial m[1201] = 1'b0;
initial m[1256] = 1'b0;
initial m[1316] = 1'b0;
initial m[1381] = 1'b0;
initial m[1451] = 1'b1;
initial m[1526] = 1'b0;
initial m[1601] = 1'b1;
initial m[1671] = 1'b0;
initial m[1736] = 1'b0;
initial m[1796] = 1'b1;
initial m[1851] = 1'b1;
initial m[1901] = 1'b1;
initial m[1946] = 1'b0;
initial m[1986] = 1'b1;
initial m[2021] = 1'b1;
initial m[2051] = 1'b1;
initial m[2076] = 1'b0;
initial m[2096] = 1'b1;
initial m[2111] = 1'b0;
initial m[2121] = 1'b1;
initial m[2126] = 1'b1;
initial m[2127] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[930] = 1'b0;
initial m[940] = 1'b0;
initial m[955] = 1'b0;
initial m[975] = 1'b0;
initial m[1000] = 1'b0;
initial m[1030] = 1'b0;
initial m[1065] = 1'b0;
initial m[1105] = 1'b0;
initial m[1150] = 1'b0;
initial m[1200] = 1'b0;
initial m[1255] = 1'b0;
initial m[1315] = 1'b0;
initial m[1380] = 1'b0;
initial m[1450] = 1'b0;
initial m[1525] = 1'b0;
initial m[1528] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR0_11(.LFSRregister(LFSRcolor0[551:506]),.clk(sample_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR0_12(.LFSRregister(LFSRcolor0[597:552]),.clk(sample_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR0_13(.LFSRregister(LFSRcolor0[643:598]),.clk(sample_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR0_14(.LFSRregister(LFSRcolor0[689:644]),.clk(sample_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR0_15(.LFSRregister(LFSRcolor0[735:690]),.clk(sample_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR0_16(.LFSRregister(LFSRcolor0[781:736]),.clk(sample_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR0_17(.LFSRregister(LFSRcolor0[827:782]),.clk(sample_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR0_18(.LFSRregister(LFSRcolor0[873:828]),.clk(sample_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR0_19(.LFSRregister(LFSRcolor0[919:874]),.clk(sample_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR0_20(.LFSRregister(LFSRcolor0[965:920]),.clk(sample_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR0_21(.LFSRregister(LFSRcolor0[1011:966]),.clk(sample_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR0_22(.LFSRregister(LFSRcolor0[1057:1012]),.clk(sample_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR0_23(.LFSRregister(LFSRcolor0[1103:1058]),.clk(sample_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR0_24(.LFSRregister(LFSRcolor0[1149:1104]),.clk(sample_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR0_25(.LFSRregister(LFSRcolor0[1195:1150]),.clk(sample_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR0_26(.LFSRregister(LFSRcolor0[1241:1196]),.clk(sample_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR0_27(.LFSRregister(LFSRcolor0[1287:1242]),.clk(sample_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR0_28(.LFSRregister(LFSRcolor0[1333:1288]),.clk(sample_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR1_15(.LFSRregister(LFSRcolor1[735:690]),.clk(color0_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR1_16(.LFSRregister(LFSRcolor1[781:736]),.clk(color0_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR1_17(.LFSRregister(LFSRcolor1[827:782]),.clk(color0_clk));
lfsr #(.seed(46'b0011001000010001001111001110101111011111000110)) LFSR1_18(.LFSRregister(LFSRcolor1[873:828]),.clk(color0_clk));
lfsr #(.seed(46'b0101000110100000010101001000010000101101100110)) LFSR1_19(.LFSRregister(LFSRcolor1[919:874]),.clk(color0_clk));
lfsr #(.seed(46'b1110011010010011001010111010100101111111100000)) LFSR1_20(.LFSRregister(LFSRcolor1[965:920]),.clk(color0_clk));
lfsr #(.seed(46'b1001111000010100100001100010110000001111101011)) LFSR1_21(.LFSRregister(LFSRcolor1[1011:966]),.clk(color0_clk));
lfsr #(.seed(46'b0011101001111100110111000000010000101100111110)) LFSR1_22(.LFSRregister(LFSRcolor1[1057:1012]),.clk(color0_clk));
lfsr #(.seed(46'b1010111010001100001100010110010011100100101100)) LFSR1_23(.LFSRregister(LFSRcolor1[1103:1058]),.clk(color0_clk));
lfsr #(.seed(46'b1101010000110001000001011010110100010000110101)) LFSR1_24(.LFSRregister(LFSRcolor1[1149:1104]),.clk(color0_clk));
lfsr #(.seed(46'b0111111000001001010001100011001110110101101001)) LFSR1_25(.LFSRregister(LFSRcolor1[1195:1150]),.clk(color0_clk));
lfsr #(.seed(46'b0111011110101100100001111000001001111001010010)) LFSR1_26(.LFSRregister(LFSRcolor1[1241:1196]),.clk(color0_clk));
lfsr #(.seed(46'b0110010001011011111100000000110011011110000100)) LFSR1_27(.LFSRregister(LFSRcolor1[1287:1242]),.clk(color0_clk));
lfsr #(.seed(46'b1100101101001001110010011101110000001110111111)) LFSR1_28(.LFSRregister(LFSRcolor1[1333:1288]),.clk(color0_clk));
lfsr #(.seed(46'b1110010100000011100111110011000001001000000101)) LFSR1_29(.LFSRregister(LFSRcolor1[1379:1334]),.clk(color0_clk));
lfsr #(.seed(46'b1100111110111110000101110101010111111010101000)) LFSR1_30(.LFSRregister(LFSRcolor1[1425:1380]),.clk(color0_clk));
lfsr #(.seed(46'b1101101000110111001110111111011011100011111101)) LFSR1_31(.LFSRregister(LFSRcolor1[1471:1426]),.clk(color0_clk));
lfsr #(.seed(46'b1011100111101011110000001101111100001111100011)) LFSR1_32(.LFSRregister(LFSRcolor1[1517:1472]),.clk(color0_clk));
lfsr #(.seed(46'b1000011101010100110111010000000111000111010111)) LFSR1_33(.LFSRregister(LFSRcolor1[1563:1518]),.clk(color0_clk));
lfsr #(.seed(46'b0011001001101100101110110001011100100100110000)) LFSR1_34(.LFSRregister(LFSRcolor1[1609:1564]),.clk(color0_clk));
lfsr #(.seed(46'b0011110010011101000111111110100110110100101000)) LFSR1_35(.LFSRregister(LFSRcolor1[1655:1610]),.clk(color0_clk));
lfsr #(.seed(46'b1100000100011100010111001011000000101100110100)) LFSR1_36(.LFSRregister(LFSRcolor1[1701:1656]),.clk(color0_clk));
lfsr #(.seed(46'b1001101001101101001001111001110100110001100010)) LFSR1_37(.LFSRregister(LFSRcolor1[1747:1702]),.clk(color0_clk));
lfsr #(.seed(46'b1000000000001101011011010100000001101001001111)) LFSR1_38(.LFSRregister(LFSRcolor1[1793:1748]),.clk(color0_clk));
lfsr #(.seed(46'b1000011000100000010011100100110100001010000001)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0101000011110010010110011011111101010101011010)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0011111001110010110000110100101000000000100010)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0011101001110100101101111100101010101100110000)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1100111100001111010111011100011110001010110011)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0101101111111000101111101010111101100011110011)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1100101101101111100100111011110111010010100100)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b0110001110010011010100101010010010100100011000)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b0010101111101011001110100001110011000100001001)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b0100110100101000110001000110101010001110100101)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b1111010011010001011111110011011111011111011010)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b0011000010001101011100101011111101010001010111)) LFSR2_11(.LFSRregister(LFSRcolor2[551:506]),.clk(color1_clk));
lfsr #(.seed(46'b0011010011011000100111011100010000001110001110)) LFSR2_12(.LFSRregister(LFSRcolor2[597:552]),.clk(color1_clk));
lfsr #(.seed(46'b0010110000011111111111101000111101111100101000)) LFSR2_13(.LFSRregister(LFSRcolor2[643:598]),.clk(color1_clk));
lfsr #(.seed(46'b1110000110010010100110000110010000011111100110)) LFSR2_14(.LFSRregister(LFSRcolor2[689:644]),.clk(color1_clk));
lfsr #(.seed(46'b0011101100010010111110000100001011000110001101)) LFSR2_15(.LFSRregister(LFSRcolor2[735:690]),.clk(color1_clk));
lfsr #(.seed(46'b0010001010111001000011110110110110100001001011)) LFSR2_16(.LFSRregister(LFSRcolor2[781:736]),.clk(color1_clk));
lfsr #(.seed(46'b1010111110010100100000100111111111101010101011)) LFSR2_17(.LFSRregister(LFSRcolor2[827:782]),.clk(color1_clk));
lfsr #(.seed(46'b0000001101010010101110010000001110111100000000)) LFSR2_18(.LFSRregister(LFSRcolor2[873:828]),.clk(color1_clk));
lfsr #(.seed(46'b0001101011110001101001101001111111011101001010)) LFSR2_19(.LFSRregister(LFSRcolor2[919:874]),.clk(color1_clk));
lfsr #(.seed(46'b1010111010011010101000111010001000010011110111)) LFSR2_20(.LFSRregister(LFSRcolor2[965:920]),.clk(color1_clk));
lfsr #(.seed(46'b0001100101111110101010111111100101111000000011)) LFSR2_21(.LFSRregister(LFSRcolor2[1011:966]),.clk(color1_clk));
lfsr #(.seed(46'b1110110011101111100000001011100011010010100101)) LFSR2_22(.LFSRregister(LFSRcolor2[1057:1012]),.clk(color1_clk));
lfsr #(.seed(46'b1110101011011010101011001110110110100100110110)) LFSR2_23(.LFSRregister(LFSRcolor2[1103:1058]),.clk(color1_clk));
lfsr #(.seed(46'b0011111111100000000000011101001000101110111011)) LFSR2_24(.LFSRregister(LFSRcolor2[1149:1104]),.clk(color1_clk));
lfsr #(.seed(46'b0111111111000000001010100101100111000000010111)) LFSR2_25(.LFSRregister(LFSRcolor2[1195:1150]),.clk(color1_clk));
lfsr #(.seed(46'b0010111000110010000000110100011011001101000000)) LFSR2_26(.LFSRregister(LFSRcolor2[1241:1196]),.clk(color1_clk));
lfsr #(.seed(46'b1101101011000110111100101001100011010100111001)) LFSR2_27(.LFSRregister(LFSRcolor2[1287:1242]),.clk(color1_clk));
lfsr #(.seed(46'b1111011111010000011011010110110000011100001001)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1111101011000001010101111101111100010010110011)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b0101100101110001001001001101011110111001010010)) LFSR3_2(.LFSRregister(LFSRcolor3[137:92]),.clk(color2_clk));
lfsr #(.seed(46'b1101101001111010000010010010000100111110010001)) LFSR3_3(.LFSRregister(LFSRcolor3[183:138]),.clk(color2_clk));
lfsr #(.seed(46'b1111000000101100101101011010011110000100110011)) LFSR3_4(.LFSRregister(LFSRcolor3[229:184]),.clk(color2_clk));
lfsr #(.seed(46'b1101010101111111011100011001110101100110111001)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1000011111100100101011011011111000001100000011)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1011001100010110101100000111011111101000010100)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0100111111000101011011111100100110100001010010)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b1000111010001010000011110001100111110100110110)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b1100000100111011010101010100011010010011010000)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b0101010110001011110100001010110111000011000110)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b0110100110100010111000101000100010110011001010)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));
lfsr #(.seed(46'b1101101011000111110111100100101001001000001000)) LFSR4_8(.LFSRregister(LFSRcolor4[413:368]),.clk(color3_clk));
lfsr #(.seed(46'b0100101010101111111110001111100100100100000010)) LFSR4_9(.LFSRregister(LFSRcolor4[459:414]),.clk(color3_clk));
lfsr #(.seed(46'b0000001011001111100011100101111110011111110011)) LFSR4_10(.LFSRregister(LFSRcolor4[505:460]),.clk(color3_clk));
lfsr #(.seed(46'b0000011001011000001100001011001111011010110000)) LFSR4_11(.LFSRregister(LFSRcolor4[551:506]),.clk(color3_clk));
lfsr #(.seed(46'b0011010001101000011011101101001100000111110001)) LFSR4_12(.LFSRregister(LFSRcolor4[597:552]),.clk(color3_clk));
lfsr #(.seed(46'b1110101010010001010111100100100011110001110111)) LFSR4_13(.LFSRregister(LFSRcolor4[643:598]),.clk(color3_clk));
lfsr #(.seed(46'b0000101001010111110000010011110000110111101011)) LFSR4_14(.LFSRregister(LFSRcolor4[689:644]),.clk(color3_clk));
lfsr #(.seed(46'b0000011110001011011000010010101101101001100100)) LFSR4_15(.LFSRregister(LFSRcolor4[735:690]),.clk(color3_clk));
lfsr #(.seed(46'b0011110010101101111001000000011110000111110110)) LFSR4_16(.LFSRregister(LFSRcolor4[781:736]),.clk(color3_clk));
lfsr #(.seed(46'b0001011110001010011011010001010011100001100111)) LFSR4_17(.LFSRregister(LFSRcolor4[827:782]),.clk(color3_clk));
lfsr #(.seed(46'b0010011001101010001000101001001010101010110000)) LFSR4_18(.LFSRregister(LFSRcolor4[873:828]),.clk(color3_clk));
lfsr #(.seed(46'b1010001011001110001110110010000010100011011000)) LFSR4_19(.LFSRregister(LFSRcolor4[919:874]),.clk(color3_clk));
lfsr #(.seed(46'b1001101010011110100011110100010110011001110001)) LFSR4_20(.LFSRregister(LFSRcolor4[965:920]),.clk(color3_clk));
//To control whether the system runs or resets using VIO and counter:
always @(posedge sample_clk) begin
    if (reset) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 32'b0;
        failure = 1'b0;
        solution_check = solution_set;
        m[672] = solution_set[0];
        m[931] = solution_set[1];
        m[941] = solution_set[2];
        m[956] = solution_set[3];
        m[976] = solution_set[4];
        m[1001] = solution_set[5];
        m[1031] = solution_set[6];
        m[1066] = solution_set[7];
        m[1106] = solution_set[8];
        m[1151] = solution_set[9];
        m[1201] = solution_set[10];
        m[1256] = solution_set[11];
        m[1316] = solution_set[12];
        m[1381] = solution_set[13];
        m[1451] = solution_set[14];
        m[1526] = solution_set[15];
        m[1601] = solution_set[16];
        m[1671] = solution_set[17];
        m[1736] = solution_set[18];
        m[1796] = solution_set[19];
        m[1851] = solution_set[20];
        m[1901] = solution_set[21];
        m[1946] = solution_set[22];
        m[1986] = solution_set[23];
        m[2021] = solution_set[24];
        m[2051] = solution_set[25];
        m[2076] = solution_set[26];
        m[2096] = solution_set[27];
        m[2111] = solution_set[28];
        m[2121] = solution_set[29];
        m[2126] = solution_set[30];
        m[2127] = solution_set[31];
    end else if (solution_flag) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 32'b0;
        failure = 1'b0;
    end else if (counter < 38'b11111111111111111111111111111111111111) begin
        if (counter == 1) begin
            InitCond[0] = UnbiasedRNG[0];
            InitCond[1] = UnbiasedRNG[1];
            InitCond[2] = UnbiasedRNG[2];
            InitCond[3] = UnbiasedRNG[3];
            InitCond[4] = UnbiasedRNG[4];
            InitCond[5] = UnbiasedRNG[5];
            InitCond[6] = UnbiasedRNG[6];
            InitCond[7] = UnbiasedRNG[7];
            InitCond[8] = UnbiasedRNG[8];
            InitCond[9] = UnbiasedRNG[9];
            InitCond[10] = UnbiasedRNG[10];
            InitCond[11] = UnbiasedRNG[11];
            InitCond[12] = UnbiasedRNG[12];
            InitCond[13] = UnbiasedRNG[13];
            InitCond[14] = UnbiasedRNG[14];
            InitCond[15] = UnbiasedRNG[15];
            InitCond[16] = UnbiasedRNG[16];
            InitCond[17] = UnbiasedRNG[17];
            InitCond[18] = UnbiasedRNG[18];
            InitCond[19] = UnbiasedRNG[19];
            InitCond[20] = UnbiasedRNG[20];
            InitCond[21] = UnbiasedRNG[21];
            InitCond[22] = UnbiasedRNG[22];
            InitCond[23] = UnbiasedRNG[23];
            InitCond[24] = UnbiasedRNG[24];
            InitCond[25] = UnbiasedRNG[25];
            InitCond[26] = UnbiasedRNG[26];
            InitCond[27] = UnbiasedRNG[27];
            InitCond[28] = UnbiasedRNG[28];
            InitCond[29] = UnbiasedRNG[29];
            InitCond[30] = UnbiasedRNG[30];
            InitCond[31] = UnbiasedRNG[31];
            InitCond[32] = UnbiasedRNG[32];
            InitCond[33] = UnbiasedRNG[33];
            InitCond[34] = UnbiasedRNG[34];
            InitCond[35] = UnbiasedRNG[35];
            InitCond[36] = UnbiasedRNG[36];
            InitCond[37] = UnbiasedRNG[37];
            InitCond[38] = UnbiasedRNG[38];
            InitCond[39] = UnbiasedRNG[39];
            InitCond[40] = UnbiasedRNG[40];
            InitCond[41] = UnbiasedRNG[41];
            InitCond[42] = UnbiasedRNG[42];
            InitCond[43] = UnbiasedRNG[43];
            InitCond[44] = UnbiasedRNG[44];
            InitCond[45] = UnbiasedRNG[45];
            InitCond[46] = UnbiasedRNG[46];
            InitCond[47] = UnbiasedRNG[47];
            InitCond[48] = UnbiasedRNG[48];
            InitCond[49] = UnbiasedRNG[49];
            InitCond[50] = UnbiasedRNG[50];
            InitCond[51] = UnbiasedRNG[51];
            InitCond[52] = UnbiasedRNG[52];
            InitCond[53] = UnbiasedRNG[53];
            InitCond[54] = UnbiasedRNG[54];
            InitCond[55] = UnbiasedRNG[55];
            InitCond[56] = UnbiasedRNG[56];
            InitCond[57] = UnbiasedRNG[57];
            InitCond[58] = UnbiasedRNG[58];
            InitCond[59] = UnbiasedRNG[59];
            InitCond[60] = UnbiasedRNG[60];
            InitCond[61] = UnbiasedRNG[61];
            InitCond[62] = UnbiasedRNG[62];
            InitCond[63] = UnbiasedRNG[63];
            InitCond[64] = UnbiasedRNG[64];
            InitCond[65] = UnbiasedRNG[65];
            InitCond[66] = UnbiasedRNG[66];
            InitCond[67] = UnbiasedRNG[67];
            InitCond[68] = UnbiasedRNG[68];
            InitCond[69] = UnbiasedRNG[69];
            InitCond[70] = UnbiasedRNG[70];
            InitCond[71] = UnbiasedRNG[71];
            InitCond[72] = UnbiasedRNG[72];
            InitCond[73] = UnbiasedRNG[73];
            InitCond[74] = UnbiasedRNG[74];
            InitCond[75] = UnbiasedRNG[75];
            InitCond[76] = UnbiasedRNG[76];
            InitCond[77] = UnbiasedRNG[77];
            InitCond[78] = UnbiasedRNG[78];
            InitCond[79] = UnbiasedRNG[79];
            InitCond[80] = UnbiasedRNG[80];
            InitCond[81] = UnbiasedRNG[81];
            InitCond[82] = UnbiasedRNG[82];
            InitCond[83] = UnbiasedRNG[83];
            InitCond[84] = UnbiasedRNG[84];
            InitCond[85] = UnbiasedRNG[85];
            InitCond[86] = UnbiasedRNG[86];
            InitCond[87] = UnbiasedRNG[87];
            InitCond[88] = UnbiasedRNG[88];
            InitCond[89] = UnbiasedRNG[89];
            InitCond[90] = UnbiasedRNG[90];
            InitCond[91] = UnbiasedRNG[91];
            InitCond[92] = UnbiasedRNG[92];
            InitCond[93] = UnbiasedRNG[93];
            InitCond[94] = UnbiasedRNG[94];
            InitCond[95] = UnbiasedRNG[95];
            InitCond[96] = UnbiasedRNG[96];
            InitCond[97] = UnbiasedRNG[97];
            InitCond[98] = UnbiasedRNG[98];
            InitCond[99] = UnbiasedRNG[99];
            InitCond[100] = UnbiasedRNG[100];
            InitCond[101] = UnbiasedRNG[101];
            InitCond[102] = UnbiasedRNG[102];
            InitCond[103] = UnbiasedRNG[103];
            InitCond[104] = UnbiasedRNG[104];
            InitCond[105] = UnbiasedRNG[105];
            InitCond[106] = UnbiasedRNG[106];
            InitCond[107] = UnbiasedRNG[107];
            InitCond[108] = UnbiasedRNG[108];
            InitCond[109] = UnbiasedRNG[109];
            InitCond[110] = UnbiasedRNG[110];
            InitCond[111] = UnbiasedRNG[111];
            InitCond[112] = UnbiasedRNG[112];
            InitCond[113] = UnbiasedRNG[113];
            InitCond[114] = UnbiasedRNG[114];
            InitCond[115] = UnbiasedRNG[115];
            InitCond[116] = UnbiasedRNG[116];
            InitCond[117] = UnbiasedRNG[117];
            InitCond[118] = UnbiasedRNG[118];
            InitCond[119] = UnbiasedRNG[119];
            InitCond[120] = UnbiasedRNG[120];
            InitCond[121] = UnbiasedRNG[121];
            InitCond[122] = UnbiasedRNG[122];
            InitCond[123] = UnbiasedRNG[123];
            InitCond[124] = UnbiasedRNG[124];
            InitCond[125] = UnbiasedRNG[125];
            InitCond[126] = UnbiasedRNG[126];
            InitCond[127] = UnbiasedRNG[127];
            InitCond[128] = UnbiasedRNG[128];
            InitCond[129] = UnbiasedRNG[129];
            InitCond[130] = UnbiasedRNG[130];
            InitCond[131] = UnbiasedRNG[131];
            InitCond[132] = UnbiasedRNG[132];
            InitCond[133] = UnbiasedRNG[133];
            InitCond[134] = UnbiasedRNG[134];
            InitCond[135] = UnbiasedRNG[135];
            InitCond[136] = UnbiasedRNG[136];
            InitCond[137] = UnbiasedRNG[137];
            InitCond[138] = UnbiasedRNG[138];
            InitCond[139] = UnbiasedRNG[139];
            InitCond[140] = UnbiasedRNG[140];
            InitCond[141] = UnbiasedRNG[141];
            InitCond[142] = UnbiasedRNG[142];
            InitCond[143] = UnbiasedRNG[143];
            InitCond[144] = UnbiasedRNG[144];
            InitCond[145] = UnbiasedRNG[145];
            InitCond[146] = UnbiasedRNG[146];
            InitCond[147] = UnbiasedRNG[147];
            InitCond[148] = UnbiasedRNG[148];
            InitCond[149] = UnbiasedRNG[149];
            InitCond[150] = UnbiasedRNG[150];
            InitCond[151] = UnbiasedRNG[151];
            InitCond[152] = UnbiasedRNG[152];
            InitCond[153] = UnbiasedRNG[153];
            InitCond[154] = UnbiasedRNG[154];
            InitCond[155] = UnbiasedRNG[155];
            InitCond[156] = UnbiasedRNG[156];
            InitCond[157] = UnbiasedRNG[157];
            InitCond[158] = UnbiasedRNG[158];
            InitCond[159] = UnbiasedRNG[159];
            InitCond[160] = UnbiasedRNG[160];
            InitCond[161] = UnbiasedRNG[161];
            InitCond[162] = UnbiasedRNG[162];
            InitCond[163] = UnbiasedRNG[163];
            InitCond[164] = UnbiasedRNG[164];
            InitCond[165] = UnbiasedRNG[165];
            InitCond[166] = UnbiasedRNG[166];
            InitCond[167] = UnbiasedRNG[167];
            InitCond[168] = UnbiasedRNG[168];
            InitCond[169] = UnbiasedRNG[169];
            InitCond[170] = UnbiasedRNG[170];
            InitCond[171] = UnbiasedRNG[171];
            InitCond[172] = UnbiasedRNG[172];
            InitCond[173] = UnbiasedRNG[173];
            InitCond[174] = UnbiasedRNG[174];
            InitCond[175] = UnbiasedRNG[175];
            InitCond[176] = UnbiasedRNG[176];
            InitCond[177] = UnbiasedRNG[177];
            InitCond[178] = UnbiasedRNG[178];
            InitCond[179] = UnbiasedRNG[179];
            InitCond[180] = UnbiasedRNG[180];
            InitCond[181] = UnbiasedRNG[181];
            InitCond[182] = UnbiasedRNG[182];
            InitCond[183] = UnbiasedRNG[183];
            InitCond[184] = UnbiasedRNG[184];
            InitCond[185] = UnbiasedRNG[185];
            InitCond[186] = UnbiasedRNG[186];
            InitCond[187] = UnbiasedRNG[187];
            InitCond[188] = UnbiasedRNG[188];
            InitCond[189] = UnbiasedRNG[189];
            InitCond[190] = UnbiasedRNG[190];
            InitCond[191] = UnbiasedRNG[191];
            InitCond[192] = UnbiasedRNG[192];
            InitCond[193] = UnbiasedRNG[193];
            InitCond[194] = UnbiasedRNG[194];
            InitCond[195] = UnbiasedRNG[195];
            InitCond[196] = UnbiasedRNG[196];
            InitCond[197] = UnbiasedRNG[197];
            InitCond[198] = UnbiasedRNG[198];
            InitCond[199] = UnbiasedRNG[199];
            InitCond[200] = UnbiasedRNG[200];
            InitCond[201] = UnbiasedRNG[201];
            InitCond[202] = UnbiasedRNG[202];
            InitCond[203] = UnbiasedRNG[203];
            InitCond[204] = UnbiasedRNG[204];
            InitCond[205] = UnbiasedRNG[205];
            InitCond[206] = UnbiasedRNG[206];
            InitCond[207] = UnbiasedRNG[207];
            InitCond[208] = UnbiasedRNG[208];
            InitCond[209] = UnbiasedRNG[209];
            InitCond[210] = UnbiasedRNG[210];
            InitCond[211] = UnbiasedRNG[211];
            InitCond[212] = UnbiasedRNG[212];
            InitCond[213] = UnbiasedRNG[213];
            InitCond[214] = UnbiasedRNG[214];
            InitCond[215] = UnbiasedRNG[215];
            InitCond[216] = UnbiasedRNG[216];
            InitCond[217] = UnbiasedRNG[217];
            InitCond[218] = UnbiasedRNG[218];
            InitCond[219] = UnbiasedRNG[219];
            InitCond[220] = UnbiasedRNG[220];
            InitCond[221] = UnbiasedRNG[221];
            InitCond[222] = UnbiasedRNG[222];
            InitCond[223] = UnbiasedRNG[223];
            InitCond[224] = UnbiasedRNG[224];
            InitCond[225] = UnbiasedRNG[225];
            InitCond[226] = UnbiasedRNG[226];
            InitCond[227] = UnbiasedRNG[227];
            InitCond[228] = UnbiasedRNG[228];
            InitCond[229] = UnbiasedRNG[229];
            InitCond[230] = UnbiasedRNG[230];
            InitCond[231] = UnbiasedRNG[231];
            InitCond[232] = UnbiasedRNG[232];
            InitCond[233] = UnbiasedRNG[233];
            InitCond[234] = UnbiasedRNG[234];
            InitCond[235] = UnbiasedRNG[235];
            InitCond[236] = UnbiasedRNG[236];
            InitCond[237] = UnbiasedRNG[237];
            InitCond[238] = UnbiasedRNG[238];
            InitCond[239] = UnbiasedRNG[239];
            InitCond[240] = UnbiasedRNG[240];
            InitCond[241] = UnbiasedRNG[241];
            InitCond[242] = UnbiasedRNG[242];
            InitCond[243] = UnbiasedRNG[243];
            InitCond[244] = UnbiasedRNG[244];
            InitCond[245] = UnbiasedRNG[245];
            InitCond[246] = UnbiasedRNG[246];
            InitCond[247] = UnbiasedRNG[247];
            InitCond[248] = UnbiasedRNG[248];
            InitCond[249] = UnbiasedRNG[249];
            InitCond[250] = UnbiasedRNG[250];
            InitCond[251] = UnbiasedRNG[251];
            InitCond[252] = UnbiasedRNG[252];
            InitCond[253] = UnbiasedRNG[253];
            InitCond[254] = UnbiasedRNG[254];
            InitCond[255] = UnbiasedRNG[255];
            InitCond[256] = UnbiasedRNG[256];
            InitCond[257] = UnbiasedRNG[257];
            InitCond[258] = UnbiasedRNG[258];
            InitCond[259] = UnbiasedRNG[259];
            InitCond[260] = UnbiasedRNG[260];
            InitCond[261] = UnbiasedRNG[261];
            InitCond[262] = UnbiasedRNG[262];
            InitCond[263] = UnbiasedRNG[263];
            InitCond[264] = UnbiasedRNG[264];
            InitCond[265] = UnbiasedRNG[265];
            InitCond[266] = UnbiasedRNG[266];
            InitCond[267] = UnbiasedRNG[267];
            InitCond[268] = UnbiasedRNG[268];
            InitCond[269] = UnbiasedRNG[269];
            InitCond[270] = UnbiasedRNG[270];
            InitCond[271] = UnbiasedRNG[271];
            InitCond[272] = UnbiasedRNG[272];
            InitCond[273] = UnbiasedRNG[273];
            InitCond[274] = UnbiasedRNG[274];
            InitCond[275] = UnbiasedRNG[275];
            InitCond[276] = UnbiasedRNG[276];
            InitCond[277] = UnbiasedRNG[277];
            InitCond[278] = UnbiasedRNG[278];
            InitCond[279] = UnbiasedRNG[279];
            InitCond[280] = UnbiasedRNG[280];
            InitCond[281] = UnbiasedRNG[281];
            InitCond[282] = UnbiasedRNG[282];
            InitCond[283] = UnbiasedRNG[283];
            InitCond[284] = UnbiasedRNG[284];
            InitCond[285] = UnbiasedRNG[285];
            InitCond[286] = UnbiasedRNG[286];
            InitCond[287] = UnbiasedRNG[287];
            InitCond[288] = UnbiasedRNG[288];
            InitCond[289] = UnbiasedRNG[289];
            InitCond[290] = UnbiasedRNG[290];
            InitCond[291] = UnbiasedRNG[291];
            InitCond[292] = UnbiasedRNG[292];
            InitCond[293] = UnbiasedRNG[293];
            InitCond[294] = UnbiasedRNG[294];
            InitCond[295] = UnbiasedRNG[295];
            InitCond[296] = UnbiasedRNG[296];
            InitCond[297] = UnbiasedRNG[297];
            InitCond[298] = UnbiasedRNG[298];
            InitCond[299] = UnbiasedRNG[299];
            InitCond[300] = UnbiasedRNG[300];
            InitCond[301] = UnbiasedRNG[301];
            InitCond[302] = UnbiasedRNG[302];
            InitCond[303] = UnbiasedRNG[303];
            InitCond[304] = UnbiasedRNG[304];
            InitCond[305] = UnbiasedRNG[305];
            InitCond[306] = UnbiasedRNG[306];
            InitCond[307] = UnbiasedRNG[307];
            InitCond[308] = UnbiasedRNG[308];
            InitCond[309] = UnbiasedRNG[309];
            InitCond[310] = UnbiasedRNG[310];
            InitCond[311] = UnbiasedRNG[311];
            InitCond[312] = UnbiasedRNG[312];
            InitCond[313] = UnbiasedRNG[313];
            InitCond[314] = UnbiasedRNG[314];
            InitCond[315] = UnbiasedRNG[315];
            InitCond[316] = UnbiasedRNG[316];
            InitCond[317] = UnbiasedRNG[317];
            InitCond[318] = UnbiasedRNG[318];
            InitCond[319] = UnbiasedRNG[319];
            InitCond[320] = UnbiasedRNG[320];
            InitCond[321] = UnbiasedRNG[321];
            InitCond[322] = UnbiasedRNG[322];
            InitCond[323] = UnbiasedRNG[323];
            InitCond[324] = UnbiasedRNG[324];
            InitCond[325] = UnbiasedRNG[325];
            InitCond[326] = UnbiasedRNG[326];
            InitCond[327] = UnbiasedRNG[327];
            InitCond[328] = UnbiasedRNG[328];
            InitCond[329] = UnbiasedRNG[329];
            InitCond[330] = UnbiasedRNG[330];
            InitCond[331] = UnbiasedRNG[331];
            InitCond[332] = UnbiasedRNG[332];
            InitCond[333] = UnbiasedRNG[333];
            InitCond[334] = UnbiasedRNG[334];
            InitCond[335] = UnbiasedRNG[335];
            InitCond[336] = UnbiasedRNG[336];
            InitCond[337] = UnbiasedRNG[337];
            InitCond[338] = UnbiasedRNG[338];
            InitCond[339] = UnbiasedRNG[339];
            InitCond[340] = UnbiasedRNG[340];
            InitCond[341] = UnbiasedRNG[341];
            InitCond[342] = UnbiasedRNG[342];
            InitCond[343] = UnbiasedRNG[343];
            InitCond[344] = UnbiasedRNG[344];
            InitCond[345] = UnbiasedRNG[345];
            InitCond[346] = UnbiasedRNG[346];
            InitCond[347] = UnbiasedRNG[347];
            InitCond[348] = UnbiasedRNG[348];
            InitCond[349] = UnbiasedRNG[349];
            InitCond[350] = UnbiasedRNG[350];
            InitCond[351] = UnbiasedRNG[351];
            InitCond[352] = UnbiasedRNG[352];
            InitCond[353] = UnbiasedRNG[353];
            InitCond[354] = UnbiasedRNG[354];
            InitCond[355] = UnbiasedRNG[355];
            InitCond[356] = UnbiasedRNG[356];
            InitCond[357] = UnbiasedRNG[357];
            InitCond[358] = UnbiasedRNG[358];
            InitCond[359] = UnbiasedRNG[359];
            InitCond[360] = UnbiasedRNG[360];
            InitCond[361] = UnbiasedRNG[361];
            InitCond[362] = UnbiasedRNG[362];
            InitCond[363] = UnbiasedRNG[363];
            InitCond[364] = UnbiasedRNG[364];
            InitCond[365] = UnbiasedRNG[365];
            InitCond[366] = UnbiasedRNG[366];
            InitCond[367] = UnbiasedRNG[367];
            InitCond[368] = UnbiasedRNG[368];
            InitCond[369] = UnbiasedRNG[369];
            InitCond[370] = UnbiasedRNG[370];
            InitCond[371] = UnbiasedRNG[371];
            InitCond[372] = UnbiasedRNG[372];
            InitCond[373] = UnbiasedRNG[373];
            InitCond[374] = UnbiasedRNG[374];
            InitCond[375] = UnbiasedRNG[375];
            InitCond[376] = UnbiasedRNG[376];
            InitCond[377] = UnbiasedRNG[377];
            InitCond[378] = UnbiasedRNG[378];
            InitCond[379] = UnbiasedRNG[379];
            InitCond[380] = UnbiasedRNG[380];
            InitCond[381] = UnbiasedRNG[381];
            InitCond[382] = UnbiasedRNG[382];
            InitCond[383] = UnbiasedRNG[383];
            InitCond[384] = UnbiasedRNG[384];
            InitCond[385] = UnbiasedRNG[385];
            InitCond[386] = UnbiasedRNG[386];
            InitCond[387] = UnbiasedRNG[387];
            InitCond[388] = UnbiasedRNG[388];
            InitCond[389] = UnbiasedRNG[389];
            InitCond[390] = UnbiasedRNG[390];
            InitCond[391] = UnbiasedRNG[391];
            InitCond[392] = UnbiasedRNG[392];
            InitCond[393] = UnbiasedRNG[393];
            InitCond[394] = UnbiasedRNG[394];
            InitCond[395] = UnbiasedRNG[395];
            InitCond[396] = UnbiasedRNG[396];
            InitCond[397] = UnbiasedRNG[397];
            InitCond[398] = UnbiasedRNG[398];
            InitCond[399] = UnbiasedRNG[399];
            InitCond[400] = UnbiasedRNG[400];
            InitCond[401] = UnbiasedRNG[401];
            InitCond[402] = UnbiasedRNG[402];
            InitCond[403] = UnbiasedRNG[403];
            InitCond[404] = UnbiasedRNG[404];
            InitCond[405] = UnbiasedRNG[405];
            InitCond[406] = UnbiasedRNG[406];
            InitCond[407] = UnbiasedRNG[407];
            InitCond[408] = UnbiasedRNG[408];
            InitCond[409] = UnbiasedRNG[409];
            InitCond[410] = UnbiasedRNG[410];
            InitCond[411] = UnbiasedRNG[411];
            InitCond[412] = UnbiasedRNG[412];
            InitCond[413] = UnbiasedRNG[413];
            InitCond[414] = UnbiasedRNG[414];
            InitCond[415] = UnbiasedRNG[415];
            InitCond[416] = UnbiasedRNG[416];
            InitCond[417] = UnbiasedRNG[417];
            InitCond[418] = UnbiasedRNG[418];
            InitCond[419] = UnbiasedRNG[419];
            InitCond[420] = UnbiasedRNG[420];
            InitCond[421] = UnbiasedRNG[421];
            InitCond[422] = UnbiasedRNG[422];
            InitCond[423] = UnbiasedRNG[423];
            InitCond[424] = UnbiasedRNG[424];
            InitCond[425] = UnbiasedRNG[425];
            InitCond[426] = UnbiasedRNG[426];
            InitCond[427] = UnbiasedRNG[427];
            InitCond[428] = UnbiasedRNG[428];
            InitCond[429] = UnbiasedRNG[429];
            InitCond[430] = UnbiasedRNG[430];
            InitCond[431] = UnbiasedRNG[431];
            InitCond[432] = UnbiasedRNG[432];
            InitCond[433] = UnbiasedRNG[433];
            InitCond[434] = UnbiasedRNG[434];
            InitCond[435] = UnbiasedRNG[435];
            InitCond[436] = UnbiasedRNG[436];
            InitCond[437] = UnbiasedRNG[437];
            InitCond[438] = UnbiasedRNG[438];
            InitCond[439] = UnbiasedRNG[439];
            InitCond[440] = UnbiasedRNG[440];
            InitCond[441] = UnbiasedRNG[441];
            InitCond[442] = UnbiasedRNG[442];
            InitCond[443] = UnbiasedRNG[443];
            InitCond[444] = UnbiasedRNG[444];
            InitCond[445] = UnbiasedRNG[445];
            InitCond[446] = UnbiasedRNG[446];
            InitCond[447] = UnbiasedRNG[447];
            InitCond[448] = UnbiasedRNG[448];
            InitCond[449] = UnbiasedRNG[449];
            InitCond[450] = UnbiasedRNG[450];
            InitCond[451] = UnbiasedRNG[451];
            InitCond[452] = UnbiasedRNG[452];
            InitCond[453] = UnbiasedRNG[453];
            InitCond[454] = UnbiasedRNG[454];
            InitCond[455] = UnbiasedRNG[455];
            InitCond[456] = UnbiasedRNG[456];
            InitCond[457] = UnbiasedRNG[457];
            InitCond[458] = UnbiasedRNG[458];
            InitCond[459] = UnbiasedRNG[459];
            InitCond[460] = UnbiasedRNG[460];
            InitCond[461] = UnbiasedRNG[461];
            InitCond[462] = UnbiasedRNG[462];
            InitCond[463] = UnbiasedRNG[463];
            InitCond[464] = UnbiasedRNG[464];
            InitCond[465] = UnbiasedRNG[465];
            InitCond[466] = UnbiasedRNG[466];
            InitCond[467] = UnbiasedRNG[467];
            InitCond[468] = UnbiasedRNG[468];
            InitCond[469] = UnbiasedRNG[469];
            InitCond[470] = UnbiasedRNG[470];
            InitCond[471] = UnbiasedRNG[471];
            InitCond[472] = UnbiasedRNG[472];
            InitCond[473] = UnbiasedRNG[473];
            InitCond[474] = UnbiasedRNG[474];
            InitCond[475] = UnbiasedRNG[475];
            InitCond[476] = UnbiasedRNG[476];
            InitCond[477] = UnbiasedRNG[477];
            InitCond[478] = UnbiasedRNG[478];
            InitCond[479] = UnbiasedRNG[479];
            InitCond[480] = UnbiasedRNG[480];
            InitCond[481] = UnbiasedRNG[481];
            InitCond[482] = UnbiasedRNG[482];
            InitCond[483] = UnbiasedRNG[483];
            InitCond[484] = UnbiasedRNG[484];
            InitCond[485] = UnbiasedRNG[485];
            InitCond[486] = UnbiasedRNG[486];
            InitCond[487] = UnbiasedRNG[487];
            InitCond[488] = UnbiasedRNG[488];
            InitCond[489] = UnbiasedRNG[489];
            InitCond[490] = UnbiasedRNG[490];
            InitCond[491] = UnbiasedRNG[491];
            InitCond[492] = UnbiasedRNG[492];
            InitCond[493] = UnbiasedRNG[493];
            InitCond[494] = UnbiasedRNG[494];
            InitCond[495] = UnbiasedRNG[495];
            InitCond[496] = UnbiasedRNG[496];
            InitCond[497] = UnbiasedRNG[497];
            InitCond[498] = UnbiasedRNG[498];
            InitCond[499] = UnbiasedRNG[499];
            InitCond[500] = UnbiasedRNG[500];
            InitCond[501] = UnbiasedRNG[501];
            InitCond[502] = UnbiasedRNG[502];
            InitCond[503] = UnbiasedRNG[503];
            InitCond[504] = UnbiasedRNG[504];
            InitCond[505] = UnbiasedRNG[505];
            InitCond[506] = UnbiasedRNG[506];
            InitCond[507] = UnbiasedRNG[507];
            InitCond[508] = UnbiasedRNG[508];
            InitCond[509] = UnbiasedRNG[509];
            InitCond[510] = UnbiasedRNG[510];
            InitCond[511] = UnbiasedRNG[511];
            InitCond[512] = UnbiasedRNG[512];
            InitCond[513] = UnbiasedRNG[513];
            InitCond[514] = UnbiasedRNG[514];
            InitCond[515] = UnbiasedRNG[515];
            InitCond[516] = UnbiasedRNG[516];
            InitCond[517] = UnbiasedRNG[517];
            InitCond[518] = UnbiasedRNG[518];
            InitCond[519] = UnbiasedRNG[519];
            InitCond[520] = UnbiasedRNG[520];
            InitCond[521] = UnbiasedRNG[521];
            InitCond[522] = UnbiasedRNG[522];
            InitCond[523] = UnbiasedRNG[523];
            InitCond[524] = UnbiasedRNG[524];
            InitCond[525] = UnbiasedRNG[525];
            InitCond[526] = UnbiasedRNG[526];
            InitCond[527] = UnbiasedRNG[527];
            InitCond[528] = UnbiasedRNG[528];
            InitCond[529] = UnbiasedRNG[529];
            InitCond[530] = UnbiasedRNG[530];
            InitCond[531] = UnbiasedRNG[531];
            InitCond[532] = UnbiasedRNG[532];
            InitCond[533] = UnbiasedRNG[533];
            InitCond[534] = UnbiasedRNG[534];
            InitCond[535] = UnbiasedRNG[535];
            InitCond[536] = UnbiasedRNG[536];
            InitCond[537] = UnbiasedRNG[537];
            InitCond[538] = UnbiasedRNG[538];
            InitCond[539] = UnbiasedRNG[539];
            InitCond[540] = UnbiasedRNG[540];
            InitCond[541] = UnbiasedRNG[541];
            InitCond[542] = UnbiasedRNG[542];
            InitCond[543] = UnbiasedRNG[543];
            InitCond[544] = UnbiasedRNG[544];
            InitCond[545] = UnbiasedRNG[545];
            InitCond[546] = UnbiasedRNG[546];
            InitCond[547] = UnbiasedRNG[547];
            InitCond[548] = UnbiasedRNG[548];
            InitCond[549] = UnbiasedRNG[549];
            InitCond[550] = UnbiasedRNG[550];
            InitCond[551] = UnbiasedRNG[551];
            InitCond[552] = UnbiasedRNG[552];
            InitCond[553] = UnbiasedRNG[553];
            InitCond[554] = UnbiasedRNG[554];
            InitCond[555] = UnbiasedRNG[555];
            InitCond[556] = UnbiasedRNG[556];
            InitCond[557] = UnbiasedRNG[557];
            InitCond[558] = UnbiasedRNG[558];
            InitCond[559] = UnbiasedRNG[559];
            InitCond[560] = UnbiasedRNG[560];
            InitCond[561] = UnbiasedRNG[561];
            InitCond[562] = UnbiasedRNG[562];
            InitCond[563] = UnbiasedRNG[563];
            InitCond[564] = UnbiasedRNG[564];
            InitCond[565] = UnbiasedRNG[565];
            InitCond[566] = UnbiasedRNG[566];
            InitCond[567] = UnbiasedRNG[567];
            InitCond[568] = UnbiasedRNG[568];
            InitCond[569] = UnbiasedRNG[569];
            InitCond[570] = UnbiasedRNG[570];
            InitCond[571] = UnbiasedRNG[571];
            InitCond[572] = UnbiasedRNG[572];
            InitCond[573] = UnbiasedRNG[573];
            InitCond[574] = UnbiasedRNG[574];
            InitCond[575] = UnbiasedRNG[575];
            InitCond[576] = UnbiasedRNG[576];
            InitCond[577] = UnbiasedRNG[577];
            InitCond[578] = UnbiasedRNG[578];
            InitCond[579] = UnbiasedRNG[579];
            InitCond[580] = UnbiasedRNG[580];
            InitCond[581] = UnbiasedRNG[581];
            InitCond[582] = UnbiasedRNG[582];
            InitCond[583] = UnbiasedRNG[583];
            InitCond[584] = UnbiasedRNG[584];
            InitCond[585] = UnbiasedRNG[585];
            InitCond[586] = UnbiasedRNG[586];
            InitCond[587] = UnbiasedRNG[587];
            InitCond[588] = UnbiasedRNG[588];
            InitCond[589] = UnbiasedRNG[589];
            InitCond[590] = UnbiasedRNG[590];
            InitCond[591] = UnbiasedRNG[591];
            InitCond[592] = UnbiasedRNG[592];
            InitCond[593] = UnbiasedRNG[593];
            InitCond[594] = UnbiasedRNG[594];
            InitCond[595] = UnbiasedRNG[595];
            InitCond[596] = UnbiasedRNG[596];
            InitCond[597] = UnbiasedRNG[597];
            InitCond[598] = UnbiasedRNG[598];
            InitCond[599] = UnbiasedRNG[599];
            InitCond[600] = UnbiasedRNG[600];
            InitCond[601] = UnbiasedRNG[601];
            InitCond[602] = UnbiasedRNG[602];
            InitCond[603] = UnbiasedRNG[603];
            InitCond[604] = UnbiasedRNG[604];
            InitCond[605] = UnbiasedRNG[605];
            InitCond[606] = UnbiasedRNG[606];
            InitCond[607] = UnbiasedRNG[607];
            InitCond[608] = UnbiasedRNG[608];
            InitCond[609] = UnbiasedRNG[609];
            InitCond[610] = UnbiasedRNG[610];
            InitCond[611] = UnbiasedRNG[611];
            InitCond[612] = UnbiasedRNG[612];
            InitCond[613] = UnbiasedRNG[613];
            InitCond[614] = UnbiasedRNG[614];
            InitCond[615] = UnbiasedRNG[615];
            InitCond[616] = UnbiasedRNG[616];
            InitCond[617] = UnbiasedRNG[617];
            InitCond[618] = UnbiasedRNG[618];
            InitCond[619] = UnbiasedRNG[619];
            InitCond[620] = UnbiasedRNG[620];
            InitCond[621] = UnbiasedRNG[621];
            InitCond[622] = UnbiasedRNG[622];
            InitCond[623] = UnbiasedRNG[623];
            InitCond[624] = UnbiasedRNG[624];
            InitCond[625] = UnbiasedRNG[625];
            InitCond[626] = UnbiasedRNG[626];
            InitCond[627] = UnbiasedRNG[627];
            InitCond[628] = UnbiasedRNG[628];
            InitCond[629] = UnbiasedRNG[629];
            InitCond[630] = UnbiasedRNG[630];
            InitCond[631] = UnbiasedRNG[631];
            InitCond[632] = UnbiasedRNG[632];
            InitCond[633] = UnbiasedRNG[633];
            InitCond[634] = UnbiasedRNG[634];
            InitCond[635] = UnbiasedRNG[635];
            InitCond[636] = UnbiasedRNG[636];
            InitCond[637] = UnbiasedRNG[637];
            InitCond[638] = UnbiasedRNG[638];
            InitCond[639] = UnbiasedRNG[639];
            InitCond[640] = UnbiasedRNG[640];
            InitCond[641] = UnbiasedRNG[641];
            InitCond[642] = UnbiasedRNG[642];
            InitCond[643] = UnbiasedRNG[643];
            InitCond[644] = UnbiasedRNG[644];
            InitCond[645] = UnbiasedRNG[645];
            InitCond[646] = UnbiasedRNG[646];
            InitCond[647] = UnbiasedRNG[647];
            InitCond[648] = UnbiasedRNG[648];
            InitCond[649] = UnbiasedRNG[649];
            InitCond[650] = UnbiasedRNG[650];
            InitCond[651] = UnbiasedRNG[651];
            InitCond[652] = UnbiasedRNG[652];
            InitCond[653] = UnbiasedRNG[653];
            InitCond[654] = UnbiasedRNG[654];
            InitCond[655] = UnbiasedRNG[655];
            InitCond[656] = UnbiasedRNG[656];
            InitCond[657] = UnbiasedRNG[657];
            InitCond[658] = UnbiasedRNG[658];
            InitCond[659] = UnbiasedRNG[659];
            InitCond[660] = UnbiasedRNG[660];
            InitCond[661] = UnbiasedRNG[661];
            InitCond[662] = UnbiasedRNG[662];
            InitCond[663] = UnbiasedRNG[663];
            InitCond[664] = UnbiasedRNG[664];
            InitCond[665] = UnbiasedRNG[665];
            InitCond[666] = UnbiasedRNG[666];
            InitCond[667] = UnbiasedRNG[667];
            InitCond[668] = UnbiasedRNG[668];
            InitCond[669] = UnbiasedRNG[669];
            InitCond[670] = UnbiasedRNG[670];
            InitCond[671] = UnbiasedRNG[671];
            InitCond[672] = UnbiasedRNG[672];
            InitCond[673] = UnbiasedRNG[673];
            InitCond[674] = UnbiasedRNG[674];
            InitCond[675] = UnbiasedRNG[675];
            InitCond[676] = UnbiasedRNG[676];
            InitCond[677] = UnbiasedRNG[677];
            InitCond[678] = UnbiasedRNG[678];
            InitCond[679] = UnbiasedRNG[679];
            InitCond[680] = UnbiasedRNG[680];
            InitCond[681] = UnbiasedRNG[681];
            InitCond[682] = UnbiasedRNG[682];
            InitCond[683] = UnbiasedRNG[683];
            InitCond[684] = UnbiasedRNG[684];
            InitCond[685] = UnbiasedRNG[685];
            InitCond[686] = UnbiasedRNG[686];
            InitCond[687] = UnbiasedRNG[687];
            InitCond[688] = UnbiasedRNG[688];
            InitCond[689] = UnbiasedRNG[689];
            InitCond[690] = UnbiasedRNG[690];
            InitCond[691] = UnbiasedRNG[691];
            InitCond[692] = UnbiasedRNG[692];
            InitCond[693] = UnbiasedRNG[693];
            InitCond[694] = UnbiasedRNG[694];
            InitCond[695] = UnbiasedRNG[695];
            InitCond[696] = UnbiasedRNG[696];
            InitCond[697] = UnbiasedRNG[697];
            InitCond[698] = UnbiasedRNG[698];
            InitCond[699] = UnbiasedRNG[699];
            InitCond[700] = UnbiasedRNG[700];
            InitCond[701] = UnbiasedRNG[701];
            InitCond[702] = UnbiasedRNG[702];
            InitCond[703] = UnbiasedRNG[703];
            InitCond[704] = UnbiasedRNG[704];
            InitCond[705] = UnbiasedRNG[705];
            InitCond[706] = UnbiasedRNG[706];
            InitCond[707] = UnbiasedRNG[707];
            InitCond[708] = UnbiasedRNG[708];
            InitCond[709] = UnbiasedRNG[709];
            InitCond[710] = UnbiasedRNG[710];
            InitCond[711] = UnbiasedRNG[711];
            InitCond[712] = UnbiasedRNG[712];
            InitCond[713] = UnbiasedRNG[713];
            InitCond[714] = UnbiasedRNG[714];
            InitCond[715] = UnbiasedRNG[715];
            InitCond[716] = UnbiasedRNG[716];
            InitCond[717] = UnbiasedRNG[717];
            InitCond[718] = UnbiasedRNG[718];
            InitCond[719] = UnbiasedRNG[719];
            InitCond[720] = UnbiasedRNG[720];
            InitCond[721] = UnbiasedRNG[721];
            InitCond[722] = UnbiasedRNG[722];
            InitCond[723] = UnbiasedRNG[723];
            InitCond[724] = UnbiasedRNG[724];
            InitCond[725] = UnbiasedRNG[725];
            InitCond[726] = UnbiasedRNG[726];
            InitCond[727] = UnbiasedRNG[727];
            InitCond[728] = UnbiasedRNG[728];
            InitCond[729] = UnbiasedRNG[729];
            InitCond[730] = UnbiasedRNG[730];
            InitCond[731] = UnbiasedRNG[731];
            InitCond[732] = UnbiasedRNG[732];
            InitCond[733] = UnbiasedRNG[733];
            InitCond[734] = UnbiasedRNG[734];
            InitCond[735] = UnbiasedRNG[735];
            InitCond[736] = UnbiasedRNG[736];
            InitCond[737] = UnbiasedRNG[737];
            InitCond[738] = UnbiasedRNG[738];
            InitCond[739] = UnbiasedRNG[739];
            InitCond[740] = UnbiasedRNG[740];
            InitCond[741] = UnbiasedRNG[741];
            InitCond[742] = UnbiasedRNG[742];
            InitCond[743] = UnbiasedRNG[743];
            InitCond[744] = UnbiasedRNG[744];
            InitCond[745] = UnbiasedRNG[745];
            InitCond[746] = UnbiasedRNG[746];
            InitCond[747] = UnbiasedRNG[747];
            InitCond[748] = UnbiasedRNG[748];
            InitCond[749] = UnbiasedRNG[749];
            InitCond[750] = UnbiasedRNG[750];
            InitCond[751] = UnbiasedRNG[751];
            InitCond[752] = UnbiasedRNG[752];
            InitCond[753] = UnbiasedRNG[753];
            InitCond[754] = UnbiasedRNG[754];
            InitCond[755] = UnbiasedRNG[755];
            InitCond[756] = UnbiasedRNG[756];
            InitCond[757] = UnbiasedRNG[757];
            InitCond[758] = UnbiasedRNG[758];
            InitCond[759] = UnbiasedRNG[759];
            InitCond[760] = UnbiasedRNG[760];
            InitCond[761] = UnbiasedRNG[761];
            InitCond[762] = UnbiasedRNG[762];
            InitCond[763] = UnbiasedRNG[763];
            InitCond[764] = UnbiasedRNG[764];
            InitCond[765] = UnbiasedRNG[765];
            InitCond[766] = UnbiasedRNG[766];
            InitCond[767] = UnbiasedRNG[767];
            InitCond[768] = UnbiasedRNG[768];
            InitCond[769] = UnbiasedRNG[769];
            InitCond[770] = UnbiasedRNG[770];
            InitCond[771] = UnbiasedRNG[771];
            InitCond[772] = UnbiasedRNG[772];
            InitCond[773] = UnbiasedRNG[773];
            InitCond[774] = UnbiasedRNG[774];
            InitCond[775] = UnbiasedRNG[775];
            InitCond[776] = UnbiasedRNG[776];
            InitCond[777] = UnbiasedRNG[777];
            InitCond[778] = UnbiasedRNG[778];
            InitCond[779] = UnbiasedRNG[779];
            InitCond[780] = UnbiasedRNG[780];
            InitCond[781] = UnbiasedRNG[781];
            InitCond[782] = UnbiasedRNG[782];
            InitCond[783] = UnbiasedRNG[783];
            InitCond[784] = UnbiasedRNG[784];
            InitCond[785] = UnbiasedRNG[785];
            InitCond[786] = UnbiasedRNG[786];
            InitCond[787] = UnbiasedRNG[787];
            InitCond[788] = UnbiasedRNG[788];
            InitCond[789] = UnbiasedRNG[789];
            InitCond[790] = UnbiasedRNG[790];
            InitCond[791] = UnbiasedRNG[791];
            InitCond[792] = UnbiasedRNG[792];
            InitCond[793] = UnbiasedRNG[793];
            InitCond[794] = UnbiasedRNG[794];
            InitCond[795] = UnbiasedRNG[795];
            InitCond[796] = UnbiasedRNG[796];
            InitCond[797] = UnbiasedRNG[797];
            InitCond[798] = UnbiasedRNG[798];
            InitCond[799] = UnbiasedRNG[799];
            InitCond[800] = UnbiasedRNG[800];
            InitCond[801] = UnbiasedRNG[801];
            InitCond[802] = UnbiasedRNG[802];
            InitCond[803] = UnbiasedRNG[803];
            InitCond[804] = UnbiasedRNG[804];
            InitCond[805] = UnbiasedRNG[805];
            InitCond[806] = UnbiasedRNG[806];
            InitCond[807] = UnbiasedRNG[807];
            InitCond[808] = UnbiasedRNG[808];
            InitCond[809] = UnbiasedRNG[809];
            InitCond[810] = UnbiasedRNG[810];
            InitCond[811] = UnbiasedRNG[811];
            InitCond[812] = UnbiasedRNG[812];
            InitCond[813] = UnbiasedRNG[813];
            InitCond[814] = UnbiasedRNG[814];
            InitCond[815] = UnbiasedRNG[815];
            InitCond[816] = UnbiasedRNG[816];
            InitCond[817] = UnbiasedRNG[817];
            InitCond[818] = UnbiasedRNG[818];
            InitCond[819] = UnbiasedRNG[819];
            InitCond[820] = UnbiasedRNG[820];
            InitCond[821] = UnbiasedRNG[821];
            InitCond[822] = UnbiasedRNG[822];
            InitCond[823] = UnbiasedRNG[823];
            InitCond[824] = UnbiasedRNG[824];
            InitCond[825] = UnbiasedRNG[825];
            InitCond[826] = UnbiasedRNG[826];
            InitCond[827] = UnbiasedRNG[827];
            InitCond[828] = UnbiasedRNG[828];
            InitCond[829] = UnbiasedRNG[829];
            InitCond[830] = UnbiasedRNG[830];
            InitCond[831] = UnbiasedRNG[831];
            InitCond[832] = UnbiasedRNG[832];
            InitCond[833] = UnbiasedRNG[833];
            InitCond[834] = UnbiasedRNG[834];
            InitCond[835] = UnbiasedRNG[835];
            InitCond[836] = UnbiasedRNG[836];
            InitCond[837] = UnbiasedRNG[837];
            InitCond[838] = UnbiasedRNG[838];
            InitCond[839] = UnbiasedRNG[839];
            InitCond[840] = UnbiasedRNG[840];
            InitCond[841] = UnbiasedRNG[841];
            InitCond[842] = UnbiasedRNG[842];
            InitCond[843] = UnbiasedRNG[843];
            InitCond[844] = UnbiasedRNG[844];
            InitCond[845] = UnbiasedRNG[845];
            InitCond[846] = UnbiasedRNG[846];
            InitCond[847] = UnbiasedRNG[847];
            InitCond[848] = UnbiasedRNG[848];
            InitCond[849] = UnbiasedRNG[849];
            InitCond[850] = UnbiasedRNG[850];
            InitCond[851] = UnbiasedRNG[851];
            InitCond[852] = UnbiasedRNG[852];
            InitCond[853] = UnbiasedRNG[853];
            InitCond[854] = UnbiasedRNG[854];
            InitCond[855] = UnbiasedRNG[855];
            InitCond[856] = UnbiasedRNG[856];
            InitCond[857] = UnbiasedRNG[857];
            InitCond[858] = UnbiasedRNG[858];
            InitCond[859] = UnbiasedRNG[859];
            InitCond[860] = UnbiasedRNG[860];
            InitCond[861] = UnbiasedRNG[861];
            InitCond[862] = UnbiasedRNG[862];
            InitCond[863] = UnbiasedRNG[863];
            InitCond[864] = UnbiasedRNG[864];
            InitCond[865] = UnbiasedRNG[865];
            InitCond[866] = UnbiasedRNG[866];
            InitCond[867] = UnbiasedRNG[867];
            InitCond[868] = UnbiasedRNG[868];
            InitCond[869] = UnbiasedRNG[869];
            InitCond[870] = UnbiasedRNG[870];
            InitCond[871] = UnbiasedRNG[871];
            InitCond[872] = UnbiasedRNG[872];
            InitCond[873] = UnbiasedRNG[873];
            InitCond[874] = UnbiasedRNG[874];
            InitCond[875] = UnbiasedRNG[875];
            InitCond[876] = UnbiasedRNG[876];
            InitCond[877] = UnbiasedRNG[877];
            InitCond[878] = UnbiasedRNG[878];
            InitCond[879] = UnbiasedRNG[879];
            InitCond[880] = UnbiasedRNG[880];
            InitCond[881] = UnbiasedRNG[881];
            InitCond[882] = UnbiasedRNG[882];
            InitCond[883] = UnbiasedRNG[883];
            InitCond[884] = UnbiasedRNG[884];
            InitCond[885] = UnbiasedRNG[885];
            InitCond[886] = UnbiasedRNG[886];
            InitCond[887] = UnbiasedRNG[887];
            InitCond[888] = UnbiasedRNG[888];
            InitCond[889] = UnbiasedRNG[889];
            InitCond[890] = UnbiasedRNG[890];
            InitCond[891] = UnbiasedRNG[891];
            InitCond[892] = UnbiasedRNG[892];
            InitCond[893] = UnbiasedRNG[893];
            InitCond[894] = UnbiasedRNG[894];
            InitCond[895] = UnbiasedRNG[895];
            InitCond[896] = UnbiasedRNG[896];
            InitCond[897] = UnbiasedRNG[897];
            InitCond[898] = UnbiasedRNG[898];
            InitCond[899] = UnbiasedRNG[899];
            InitCond[900] = UnbiasedRNG[900];
            InitCond[901] = UnbiasedRNG[901];
            InitCond[902] = UnbiasedRNG[902];
            InitCond[903] = UnbiasedRNG[903];
            InitCond[904] = UnbiasedRNG[904];
            InitCond[905] = UnbiasedRNG[905];
            InitCond[906] = UnbiasedRNG[906];
            InitCond[907] = UnbiasedRNG[907];
            InitCond[908] = UnbiasedRNG[908];
            InitCond[909] = UnbiasedRNG[909];
            InitCond[910] = UnbiasedRNG[910];
            InitCond[911] = UnbiasedRNG[911];
            InitCond[912] = UnbiasedRNG[912];
            InitCond[913] = UnbiasedRNG[913];
            InitCond[914] = UnbiasedRNG[914];
            InitCond[915] = UnbiasedRNG[915];
            InitCond[916] = UnbiasedRNG[916];
            InitCond[917] = UnbiasedRNG[917];
            InitCond[918] = UnbiasedRNG[918];
            InitCond[919] = UnbiasedRNG[919];
            InitCond[920] = UnbiasedRNG[920];
            InitCond[921] = UnbiasedRNG[921];
            InitCond[922] = UnbiasedRNG[922];
            InitCond[923] = UnbiasedRNG[923];
            InitCond[924] = UnbiasedRNG[924];
            InitCond[925] = UnbiasedRNG[925];
            InitCond[926] = UnbiasedRNG[926];
            InitCond[927] = UnbiasedRNG[927];
            InitCond[928] = UnbiasedRNG[928];
            InitCond[929] = UnbiasedRNG[929];
            InitCond[930] = UnbiasedRNG[930];
            InitCond[931] = UnbiasedRNG[931];
            InitCond[932] = UnbiasedRNG[932];
            InitCond[933] = UnbiasedRNG[933];
            InitCond[934] = UnbiasedRNG[934];
            InitCond[935] = UnbiasedRNG[935];
            InitCond[936] = UnbiasedRNG[936];
            InitCond[937] = UnbiasedRNG[937];
            InitCond[938] = UnbiasedRNG[938];
            InitCond[939] = UnbiasedRNG[939];
            InitCond[940] = UnbiasedRNG[940];
            InitCond[941] = UnbiasedRNG[941];
            InitCond[942] = UnbiasedRNG[942];
            InitCond[943] = UnbiasedRNG[943];
            InitCond[944] = UnbiasedRNG[944];
            InitCond[945] = UnbiasedRNG[945];
        end
        else if (counter == 2) begin
            InitCond[946] = UnbiasedRNG[0];
            InitCond[947] = UnbiasedRNG[1];
            InitCond[948] = UnbiasedRNG[2];
            InitCond[949] = UnbiasedRNG[3];
            InitCond[950] = UnbiasedRNG[4];
            InitCond[951] = UnbiasedRNG[5];
            InitCond[952] = UnbiasedRNG[6];
            InitCond[953] = UnbiasedRNG[7];
            InitCond[954] = UnbiasedRNG[8];
            InitCond[955] = UnbiasedRNG[9];
            InitCond[956] = UnbiasedRNG[10];
            InitCond[957] = UnbiasedRNG[11];
            InitCond[958] = UnbiasedRNG[12];
            InitCond[959] = UnbiasedRNG[13];
            InitCond[960] = UnbiasedRNG[14];
            InitCond[961] = UnbiasedRNG[15];
            InitCond[962] = UnbiasedRNG[16];
            InitCond[963] = UnbiasedRNG[17];
            InitCond[964] = UnbiasedRNG[18];
            InitCond[965] = UnbiasedRNG[19];
            InitCond[966] = UnbiasedRNG[20];
            InitCond[967] = UnbiasedRNG[21];
            InitCond[968] = UnbiasedRNG[22];
            InitCond[969] = UnbiasedRNG[23];
            InitCond[970] = UnbiasedRNG[24];
            InitCond[971] = UnbiasedRNG[25];
            InitCond[972] = UnbiasedRNG[26];
            InitCond[973] = UnbiasedRNG[27];
            InitCond[974] = UnbiasedRNG[28];
            InitCond[975] = UnbiasedRNG[29];
            InitCond[976] = UnbiasedRNG[30];
            InitCond[977] = UnbiasedRNG[31];
            InitCond[978] = UnbiasedRNG[32];
            InitCond[979] = UnbiasedRNG[33];
            InitCond[980] = UnbiasedRNG[34];
            InitCond[981] = UnbiasedRNG[35];
            InitCond[982] = UnbiasedRNG[36];
            InitCond[983] = UnbiasedRNG[37];
            InitCond[984] = UnbiasedRNG[38];
            InitCond[985] = UnbiasedRNG[39];
            InitCond[986] = UnbiasedRNG[40];
            InitCond[987] = UnbiasedRNG[41];
            InitCond[988] = UnbiasedRNG[42];
            InitCond[989] = UnbiasedRNG[43];
            InitCond[990] = UnbiasedRNG[44];
            InitCond[991] = UnbiasedRNG[45];
            InitCond[992] = UnbiasedRNG[46];
            InitCond[993] = UnbiasedRNG[47];
            InitCond[994] = UnbiasedRNG[48];
            InitCond[995] = UnbiasedRNG[49];
            InitCond[996] = UnbiasedRNG[50];
            InitCond[997] = UnbiasedRNG[51];
            InitCond[998] = UnbiasedRNG[52];
            InitCond[999] = UnbiasedRNG[53];
            InitCond[1000] = UnbiasedRNG[54];
            InitCond[1001] = UnbiasedRNG[55];
            InitCond[1002] = UnbiasedRNG[56];
            InitCond[1003] = UnbiasedRNG[57];
            InitCond[1004] = UnbiasedRNG[58];
            InitCond[1005] = UnbiasedRNG[59];
            InitCond[1006] = UnbiasedRNG[60];
            InitCond[1007] = UnbiasedRNG[61];
            InitCond[1008] = UnbiasedRNG[62];
            InitCond[1009] = UnbiasedRNG[63];
            InitCond[1010] = UnbiasedRNG[64];
            InitCond[1011] = UnbiasedRNG[65];
            InitCond[1012] = UnbiasedRNG[66];
            InitCond[1013] = UnbiasedRNG[67];
            InitCond[1014] = UnbiasedRNG[68];
            InitCond[1015] = UnbiasedRNG[69];
            InitCond[1016] = UnbiasedRNG[70];
            InitCond[1017] = UnbiasedRNG[71];
            InitCond[1018] = UnbiasedRNG[72];
            InitCond[1019] = UnbiasedRNG[73];
            InitCond[1020] = UnbiasedRNG[74];
            InitCond[1021] = UnbiasedRNG[75];
            InitCond[1022] = UnbiasedRNG[76];
            InitCond[1023] = UnbiasedRNG[77];
            InitCond[1024] = UnbiasedRNG[78];
            InitCond[1025] = UnbiasedRNG[79];
            InitCond[1026] = UnbiasedRNG[80];
            InitCond[1027] = UnbiasedRNG[81];
            InitCond[1028] = UnbiasedRNG[82];
            InitCond[1029] = UnbiasedRNG[83];
            InitCond[1030] = UnbiasedRNG[84];
            InitCond[1031] = UnbiasedRNG[85];
            InitCond[1032] = UnbiasedRNG[86];
            InitCond[1033] = UnbiasedRNG[87];
            InitCond[1034] = UnbiasedRNG[88];
            InitCond[1035] = UnbiasedRNG[89];
            InitCond[1036] = UnbiasedRNG[90];
            InitCond[1037] = UnbiasedRNG[91];
            InitCond[1038] = UnbiasedRNG[92];
            InitCond[1039] = UnbiasedRNG[93];
            InitCond[1040] = UnbiasedRNG[94];
            InitCond[1041] = UnbiasedRNG[95];
            InitCond[1042] = UnbiasedRNG[96];
            InitCond[1043] = UnbiasedRNG[97];
            InitCond[1044] = UnbiasedRNG[98];
            InitCond[1045] = UnbiasedRNG[99];
            InitCond[1046] = UnbiasedRNG[100];
            InitCond[1047] = UnbiasedRNG[101];
            InitCond[1048] = UnbiasedRNG[102];
            InitCond[1049] = UnbiasedRNG[103];
            InitCond[1050] = UnbiasedRNG[104];
            InitCond[1051] = UnbiasedRNG[105];
            InitCond[1052] = UnbiasedRNG[106];
            InitCond[1053] = UnbiasedRNG[107];
            InitCond[1054] = UnbiasedRNG[108];
            InitCond[1055] = UnbiasedRNG[109];
            InitCond[1056] = UnbiasedRNG[110];
            InitCond[1057] = UnbiasedRNG[111];
            InitCond[1058] = UnbiasedRNG[112];
            InitCond[1059] = UnbiasedRNG[113];
            InitCond[1060] = UnbiasedRNG[114];
            InitCond[1061] = UnbiasedRNG[115];
            InitCond[1062] = UnbiasedRNG[116];
            InitCond[1063] = UnbiasedRNG[117];
            InitCond[1064] = UnbiasedRNG[118];
            InitCond[1065] = UnbiasedRNG[119];
            InitCond[1066] = UnbiasedRNG[120];
            InitCond[1067] = UnbiasedRNG[121];
            InitCond[1068] = UnbiasedRNG[122];
            InitCond[1069] = UnbiasedRNG[123];
            InitCond[1070] = UnbiasedRNG[124];
            InitCond[1071] = UnbiasedRNG[125];
            InitCond[1072] = UnbiasedRNG[126];
            InitCond[1073] = UnbiasedRNG[127];
            InitCond[1074] = UnbiasedRNG[128];
            InitCond[1075] = UnbiasedRNG[129];
            InitCond[1076] = UnbiasedRNG[130];
            InitCond[1077] = UnbiasedRNG[131];
            InitCond[1078] = UnbiasedRNG[132];
            InitCond[1079] = UnbiasedRNG[133];
            InitCond[1080] = UnbiasedRNG[134];
            InitCond[1081] = UnbiasedRNG[135];
            InitCond[1082] = UnbiasedRNG[136];
            InitCond[1083] = UnbiasedRNG[137];
            InitCond[1084] = UnbiasedRNG[138];
            InitCond[1085] = UnbiasedRNG[139];
            InitCond[1086] = UnbiasedRNG[140];
            InitCond[1087] = UnbiasedRNG[141];
            InitCond[1088] = UnbiasedRNG[142];
            InitCond[1089] = UnbiasedRNG[143];
            InitCond[1090] = UnbiasedRNG[144];
            InitCond[1091] = UnbiasedRNG[145];
            InitCond[1092] = UnbiasedRNG[146];
            InitCond[1093] = UnbiasedRNG[147];
            InitCond[1094] = UnbiasedRNG[148];
            InitCond[1095] = UnbiasedRNG[149];
            InitCond[1096] = UnbiasedRNG[150];
            InitCond[1097] = UnbiasedRNG[151];
            InitCond[1098] = UnbiasedRNG[152];
            InitCond[1099] = UnbiasedRNG[153];
            InitCond[1100] = UnbiasedRNG[154];
            InitCond[1101] = UnbiasedRNG[155];
            InitCond[1102] = UnbiasedRNG[156];
            InitCond[1103] = UnbiasedRNG[157];
            InitCond[1104] = UnbiasedRNG[158];
            InitCond[1105] = UnbiasedRNG[159];
            InitCond[1106] = UnbiasedRNG[160];
            InitCond[1107] = UnbiasedRNG[161];
            InitCond[1108] = UnbiasedRNG[162];
            InitCond[1109] = UnbiasedRNG[163];
            InitCond[1110] = UnbiasedRNG[164];
            InitCond[1111] = UnbiasedRNG[165];
            InitCond[1112] = UnbiasedRNG[166];
            InitCond[1113] = UnbiasedRNG[167];
            InitCond[1114] = UnbiasedRNG[168];
            InitCond[1115] = UnbiasedRNG[169];
            InitCond[1116] = UnbiasedRNG[170];
            InitCond[1117] = UnbiasedRNG[171];
            InitCond[1118] = UnbiasedRNG[172];
            InitCond[1119] = UnbiasedRNG[173];
            InitCond[1120] = UnbiasedRNG[174];
            InitCond[1121] = UnbiasedRNG[175];
            InitCond[1122] = UnbiasedRNG[176];
            InitCond[1123] = UnbiasedRNG[177];
            InitCond[1124] = UnbiasedRNG[178];
            InitCond[1125] = UnbiasedRNG[179];
            InitCond[1126] = UnbiasedRNG[180];
            InitCond[1127] = UnbiasedRNG[181];
            InitCond[1128] = UnbiasedRNG[182];
            InitCond[1129] = UnbiasedRNG[183];
            InitCond[1130] = UnbiasedRNG[184];
            InitCond[1131] = UnbiasedRNG[185];
            InitCond[1132] = UnbiasedRNG[186];
            InitCond[1133] = UnbiasedRNG[187];
            InitCond[1134] = UnbiasedRNG[188];
            InitCond[1135] = UnbiasedRNG[189];
            InitCond[1136] = UnbiasedRNG[190];
            InitCond[1137] = UnbiasedRNG[191];
            InitCond[1138] = UnbiasedRNG[192];
            InitCond[1139] = UnbiasedRNG[193];
            InitCond[1140] = UnbiasedRNG[194];
            InitCond[1141] = UnbiasedRNG[195];
            InitCond[1142] = UnbiasedRNG[196];
            InitCond[1143] = UnbiasedRNG[197];
            InitCond[1144] = UnbiasedRNG[198];
            InitCond[1145] = UnbiasedRNG[199];
            InitCond[1146] = UnbiasedRNG[200];
            InitCond[1147] = UnbiasedRNG[201];
            InitCond[1148] = UnbiasedRNG[202];
            InitCond[1149] = UnbiasedRNG[203];
            InitCond[1150] = UnbiasedRNG[204];
            InitCond[1151] = UnbiasedRNG[205];
            InitCond[1152] = UnbiasedRNG[206];
            InitCond[1153] = UnbiasedRNG[207];
            InitCond[1154] = UnbiasedRNG[208];
            InitCond[1155] = UnbiasedRNG[209];
            InitCond[1156] = UnbiasedRNG[210];
            InitCond[1157] = UnbiasedRNG[211];
            InitCond[1158] = UnbiasedRNG[212];
            InitCond[1159] = UnbiasedRNG[213];
            InitCond[1160] = UnbiasedRNG[214];
            InitCond[1161] = UnbiasedRNG[215];
            InitCond[1162] = UnbiasedRNG[216];
            InitCond[1163] = UnbiasedRNG[217];
            InitCond[1164] = UnbiasedRNG[218];
            InitCond[1165] = UnbiasedRNG[219];
            InitCond[1166] = UnbiasedRNG[220];
            InitCond[1167] = UnbiasedRNG[221];
            InitCond[1168] = UnbiasedRNG[222];
            InitCond[1169] = UnbiasedRNG[223];
            InitCond[1170] = UnbiasedRNG[224];
            InitCond[1171] = UnbiasedRNG[225];
            InitCond[1172] = UnbiasedRNG[226];
            InitCond[1173] = UnbiasedRNG[227];
            InitCond[1174] = UnbiasedRNG[228];
            InitCond[1175] = UnbiasedRNG[229];
            InitCond[1176] = UnbiasedRNG[230];
            InitCond[1177] = UnbiasedRNG[231];
            InitCond[1178] = UnbiasedRNG[232];
            InitCond[1179] = UnbiasedRNG[233];
            InitCond[1180] = UnbiasedRNG[234];
            InitCond[1181] = UnbiasedRNG[235];
            InitCond[1182] = UnbiasedRNG[236];
            InitCond[1183] = UnbiasedRNG[237];
            InitCond[1184] = UnbiasedRNG[238];
            InitCond[1185] = UnbiasedRNG[239];
            InitCond[1186] = UnbiasedRNG[240];
            InitCond[1187] = UnbiasedRNG[241];
            InitCond[1188] = UnbiasedRNG[242];
            InitCond[1189] = UnbiasedRNG[243];
            InitCond[1190] = UnbiasedRNG[244];
            InitCond[1191] = UnbiasedRNG[245];
            InitCond[1192] = UnbiasedRNG[246];
            InitCond[1193] = UnbiasedRNG[247];
            InitCond[1194] = UnbiasedRNG[248];
            InitCond[1195] = UnbiasedRNG[249];
            InitCond[1196] = UnbiasedRNG[250];
            InitCond[1197] = UnbiasedRNG[251];
            InitCond[1198] = UnbiasedRNG[252];
            InitCond[1199] = UnbiasedRNG[253];
            InitCond[1200] = UnbiasedRNG[254];
            InitCond[1201] = UnbiasedRNG[255];
            InitCond[1202] = UnbiasedRNG[256];
            InitCond[1203] = UnbiasedRNG[257];
            InitCond[1204] = UnbiasedRNG[258];
            InitCond[1205] = UnbiasedRNG[259];
            InitCond[1206] = UnbiasedRNG[260];
            InitCond[1207] = UnbiasedRNG[261];
            InitCond[1208] = UnbiasedRNG[262];
            InitCond[1209] = UnbiasedRNG[263];
            InitCond[1210] = UnbiasedRNG[264];
            InitCond[1211] = UnbiasedRNG[265];
            InitCond[1212] = UnbiasedRNG[266];
            InitCond[1213] = UnbiasedRNG[267];
            InitCond[1214] = UnbiasedRNG[268];
            InitCond[1215] = UnbiasedRNG[269];
            InitCond[1216] = UnbiasedRNG[270];
            InitCond[1217] = UnbiasedRNG[271];
            InitCond[1218] = UnbiasedRNG[272];
            InitCond[1219] = UnbiasedRNG[273];
            InitCond[1220] = UnbiasedRNG[274];
            InitCond[1221] = UnbiasedRNG[275];
            InitCond[1222] = UnbiasedRNG[276];
            InitCond[1223] = UnbiasedRNG[277];
            InitCond[1224] = UnbiasedRNG[278];
            InitCond[1225] = UnbiasedRNG[279];
            InitCond[1226] = UnbiasedRNG[280];
            InitCond[1227] = UnbiasedRNG[281];
            InitCond[1228] = UnbiasedRNG[282];
            InitCond[1229] = UnbiasedRNG[283];
            InitCond[1230] = UnbiasedRNG[284];
            InitCond[1231] = UnbiasedRNG[285];
            InitCond[1232] = UnbiasedRNG[286];
            InitCond[1233] = UnbiasedRNG[287];
            InitCond[1234] = UnbiasedRNG[288];
            InitCond[1235] = UnbiasedRNG[289];
            InitCond[1236] = UnbiasedRNG[290];
            InitCond[1237] = UnbiasedRNG[291];
            InitCond[1238] = UnbiasedRNG[292];
            InitCond[1239] = UnbiasedRNG[293];
            InitCond[1240] = UnbiasedRNG[294];
            InitCond[1241] = UnbiasedRNG[295];
            InitCond[1242] = UnbiasedRNG[296];
            InitCond[1243] = UnbiasedRNG[297];
            InitCond[1244] = UnbiasedRNG[298];
            InitCond[1245] = UnbiasedRNG[299];
            InitCond[1246] = UnbiasedRNG[300];
            InitCond[1247] = UnbiasedRNG[301];
            InitCond[1248] = UnbiasedRNG[302];
            InitCond[1249] = UnbiasedRNG[303];
            InitCond[1250] = UnbiasedRNG[304];
            InitCond[1251] = UnbiasedRNG[305];
            InitCond[1252] = UnbiasedRNG[306];
            InitCond[1253] = UnbiasedRNG[307];
            InitCond[1254] = UnbiasedRNG[308];
            InitCond[1255] = UnbiasedRNG[309];
            InitCond[1256] = UnbiasedRNG[310];
            InitCond[1257] = UnbiasedRNG[311];
            InitCond[1258] = UnbiasedRNG[312];
            InitCond[1259] = UnbiasedRNG[313];
            InitCond[1260] = UnbiasedRNG[314];
            InitCond[1261] = UnbiasedRNG[315];
            InitCond[1262] = UnbiasedRNG[316];
            InitCond[1263] = UnbiasedRNG[317];
            InitCond[1264] = UnbiasedRNG[318];
            InitCond[1265] = UnbiasedRNG[319];
            InitCond[1266] = UnbiasedRNG[320];
            InitCond[1267] = UnbiasedRNG[321];
            InitCond[1268] = UnbiasedRNG[322];
            InitCond[1269] = UnbiasedRNG[323];
            InitCond[1270] = UnbiasedRNG[324];
            InitCond[1271] = UnbiasedRNG[325];
            InitCond[1272] = UnbiasedRNG[326];
            InitCond[1273] = UnbiasedRNG[327];
            InitCond[1274] = UnbiasedRNG[328];
            InitCond[1275] = UnbiasedRNG[329];
            InitCond[1276] = UnbiasedRNG[330];
            InitCond[1277] = UnbiasedRNG[331];
            InitCond[1278] = UnbiasedRNG[332];
            InitCond[1279] = UnbiasedRNG[333];
            InitCond[1280] = UnbiasedRNG[334];
            InitCond[1281] = UnbiasedRNG[335];
            InitCond[1282] = UnbiasedRNG[336];
            InitCond[1283] = UnbiasedRNG[337];
            InitCond[1284] = UnbiasedRNG[338];
            InitCond[1285] = UnbiasedRNG[339];
            InitCond[1286] = UnbiasedRNG[340];
            InitCond[1287] = UnbiasedRNG[341];
            InitCond[1288] = UnbiasedRNG[342];
            InitCond[1289] = UnbiasedRNG[343];
            InitCond[1290] = UnbiasedRNG[344];
            InitCond[1291] = UnbiasedRNG[345];
            InitCond[1292] = UnbiasedRNG[346];
            InitCond[1293] = UnbiasedRNG[347];
            InitCond[1294] = UnbiasedRNG[348];
            InitCond[1295] = UnbiasedRNG[349];
            InitCond[1296] = UnbiasedRNG[350];
            InitCond[1297] = UnbiasedRNG[351];
            InitCond[1298] = UnbiasedRNG[352];
            InitCond[1299] = UnbiasedRNG[353];
            InitCond[1300] = UnbiasedRNG[354];
            InitCond[1301] = UnbiasedRNG[355];
            InitCond[1302] = UnbiasedRNG[356];
            InitCond[1303] = UnbiasedRNG[357];
            InitCond[1304] = UnbiasedRNG[358];
            InitCond[1305] = UnbiasedRNG[359];
            InitCond[1306] = UnbiasedRNG[360];
            InitCond[1307] = UnbiasedRNG[361];
            InitCond[1308] = UnbiasedRNG[362];
            InitCond[1309] = UnbiasedRNG[363];
            InitCond[1310] = UnbiasedRNG[364];
            InitCond[1311] = UnbiasedRNG[365];
            InitCond[1312] = UnbiasedRNG[366];
            InitCond[1313] = UnbiasedRNG[367];
            InitCond[1314] = UnbiasedRNG[368];
            InitCond[1315] = UnbiasedRNG[369];
            InitCond[1316] = UnbiasedRNG[370];
            InitCond[1317] = UnbiasedRNG[371];
            InitCond[1318] = UnbiasedRNG[372];
            InitCond[1319] = UnbiasedRNG[373];
            InitCond[1320] = UnbiasedRNG[374];
            InitCond[1321] = UnbiasedRNG[375];
            InitCond[1322] = UnbiasedRNG[376];
            InitCond[1323] = UnbiasedRNG[377];
            InitCond[1324] = UnbiasedRNG[378];
            InitCond[1325] = UnbiasedRNG[379];
            InitCond[1326] = UnbiasedRNG[380];
            InitCond[1327] = UnbiasedRNG[381];
            InitCond[1328] = UnbiasedRNG[382];
            InitCond[1329] = UnbiasedRNG[383];
            InitCond[1330] = UnbiasedRNG[384];
            InitCond[1331] = UnbiasedRNG[385];
            InitCond[1332] = UnbiasedRNG[386];
            InitCond[1333] = UnbiasedRNG[387];
            InitCond[1334] = UnbiasedRNG[388];
            InitCond[1335] = UnbiasedRNG[389];
            InitCond[1336] = UnbiasedRNG[390];
            InitCond[1337] = UnbiasedRNG[391];
            InitCond[1338] = UnbiasedRNG[392];
            InitCond[1339] = UnbiasedRNG[393];
            InitCond[1340] = UnbiasedRNG[394];
            InitCond[1341] = UnbiasedRNG[395];
            InitCond[1342] = UnbiasedRNG[396];
            InitCond[1343] = UnbiasedRNG[397];
            InitCond[1344] = UnbiasedRNG[398];
            InitCond[1345] = UnbiasedRNG[399];
            InitCond[1346] = UnbiasedRNG[400];
            InitCond[1347] = UnbiasedRNG[401];
            InitCond[1348] = UnbiasedRNG[402];
            InitCond[1349] = UnbiasedRNG[403];
            InitCond[1350] = UnbiasedRNG[404];
            InitCond[1351] = UnbiasedRNG[405];
            InitCond[1352] = UnbiasedRNG[406];
            InitCond[1353] = UnbiasedRNG[407];
            InitCond[1354] = UnbiasedRNG[408];
            InitCond[1355] = UnbiasedRNG[409];
            InitCond[1356] = UnbiasedRNG[410];
            InitCond[1357] = UnbiasedRNG[411];
            InitCond[1358] = UnbiasedRNG[412];
            InitCond[1359] = UnbiasedRNG[413];
            InitCond[1360] = UnbiasedRNG[414];
            InitCond[1361] = UnbiasedRNG[415];
            InitCond[1362] = UnbiasedRNG[416];
            InitCond[1363] = UnbiasedRNG[417];
            InitCond[1364] = UnbiasedRNG[418];
            InitCond[1365] = UnbiasedRNG[419];
            InitCond[1366] = UnbiasedRNG[420];
            InitCond[1367] = UnbiasedRNG[421];
            InitCond[1368] = UnbiasedRNG[422];
            InitCond[1369] = UnbiasedRNG[423];
            InitCond[1370] = UnbiasedRNG[424];
            InitCond[1371] = UnbiasedRNG[425];
            InitCond[1372] = UnbiasedRNG[426];
            InitCond[1373] = UnbiasedRNG[427];
            InitCond[1374] = UnbiasedRNG[428];
            InitCond[1375] = UnbiasedRNG[429];
            InitCond[1376] = UnbiasedRNG[430];
            InitCond[1377] = UnbiasedRNG[431];
            InitCond[1378] = UnbiasedRNG[432];
            InitCond[1379] = UnbiasedRNG[433];
            InitCond[1380] = UnbiasedRNG[434];
            InitCond[1381] = UnbiasedRNG[435];
            InitCond[1382] = UnbiasedRNG[436];
            InitCond[1383] = UnbiasedRNG[437];
            InitCond[1384] = UnbiasedRNG[438];
            InitCond[1385] = UnbiasedRNG[439];
            InitCond[1386] = UnbiasedRNG[440];
            InitCond[1387] = UnbiasedRNG[441];
            InitCond[1388] = UnbiasedRNG[442];
            InitCond[1389] = UnbiasedRNG[443];
            InitCond[1390] = UnbiasedRNG[444];
            InitCond[1391] = UnbiasedRNG[445];
            InitCond[1392] = UnbiasedRNG[446];
            InitCond[1393] = UnbiasedRNG[447];
            InitCond[1394] = UnbiasedRNG[448];
            InitCond[1395] = UnbiasedRNG[449];
            InitCond[1396] = UnbiasedRNG[450];
            InitCond[1397] = UnbiasedRNG[451];
            InitCond[1398] = UnbiasedRNG[452];
            InitCond[1399] = UnbiasedRNG[453];
            InitCond[1400] = UnbiasedRNG[454];
            InitCond[1401] = UnbiasedRNG[455];
            InitCond[1402] = UnbiasedRNG[456];
            InitCond[1403] = UnbiasedRNG[457];
            InitCond[1404] = UnbiasedRNG[458];
            InitCond[1405] = UnbiasedRNG[459];
            InitCond[1406] = UnbiasedRNG[460];
            InitCond[1407] = UnbiasedRNG[461];
            InitCond[1408] = UnbiasedRNG[462];
            InitCond[1409] = UnbiasedRNG[463];
            InitCond[1410] = UnbiasedRNG[464];
            InitCond[1411] = UnbiasedRNG[465];
            InitCond[1412] = UnbiasedRNG[466];
            InitCond[1413] = UnbiasedRNG[467];
            InitCond[1414] = UnbiasedRNG[468];
            InitCond[1415] = UnbiasedRNG[469];
            InitCond[1416] = UnbiasedRNG[470];
            InitCond[1417] = UnbiasedRNG[471];
            InitCond[1418] = UnbiasedRNG[472];
            InitCond[1419] = UnbiasedRNG[473];
            InitCond[1420] = UnbiasedRNG[474];
            InitCond[1421] = UnbiasedRNG[475];
            InitCond[1422] = UnbiasedRNG[476];
            InitCond[1423] = UnbiasedRNG[477];
            InitCond[1424] = UnbiasedRNG[478];
            InitCond[1425] = UnbiasedRNG[479];
            InitCond[1426] = UnbiasedRNG[480];
            InitCond[1427] = UnbiasedRNG[481];
            InitCond[1428] = UnbiasedRNG[482];
            InitCond[1429] = UnbiasedRNG[483];
            InitCond[1430] = UnbiasedRNG[484];
            InitCond[1431] = UnbiasedRNG[485];
            InitCond[1432] = UnbiasedRNG[486];
            InitCond[1433] = UnbiasedRNG[487];
            InitCond[1434] = UnbiasedRNG[488];
            InitCond[1435] = UnbiasedRNG[489];
            InitCond[1436] = UnbiasedRNG[490];
            InitCond[1437] = UnbiasedRNG[491];
            InitCond[1438] = UnbiasedRNG[492];
            InitCond[1439] = UnbiasedRNG[493];
            InitCond[1440] = UnbiasedRNG[494];
            InitCond[1441] = UnbiasedRNG[495];
            InitCond[1442] = UnbiasedRNG[496];
            InitCond[1443] = UnbiasedRNG[497];
            InitCond[1444] = UnbiasedRNG[498];
            InitCond[1445] = UnbiasedRNG[499];
            InitCond[1446] = UnbiasedRNG[500];
            InitCond[1447] = UnbiasedRNG[501];
            InitCond[1448] = UnbiasedRNG[502];
            InitCond[1449] = UnbiasedRNG[503];
            InitCond[1450] = UnbiasedRNG[504];
            InitCond[1451] = UnbiasedRNG[505];
            InitCond[1452] = UnbiasedRNG[506];
            InitCond[1453] = UnbiasedRNG[507];
            InitCond[1454] = UnbiasedRNG[508];
            InitCond[1455] = UnbiasedRNG[509];
            InitCond[1456] = UnbiasedRNG[510];
            InitCond[1457] = UnbiasedRNG[511];
            InitCond[1458] = UnbiasedRNG[512];
            InitCond[1459] = UnbiasedRNG[513];
            InitCond[1460] = UnbiasedRNG[514];
            InitCond[1461] = UnbiasedRNG[515];
            InitCond[1462] = UnbiasedRNG[516];
            InitCond[1463] = UnbiasedRNG[517];
            InitCond[1464] = UnbiasedRNG[518];
            InitCond[1465] = UnbiasedRNG[519];
            InitCond[1466] = UnbiasedRNG[520];
            InitCond[1467] = UnbiasedRNG[521];
            InitCond[1468] = UnbiasedRNG[522];
            InitCond[1469] = UnbiasedRNG[523];
            InitCond[1470] = UnbiasedRNG[524];
            InitCond[1471] = UnbiasedRNG[525];
            InitCond[1472] = UnbiasedRNG[526];
            InitCond[1473] = UnbiasedRNG[527];
            InitCond[1474] = UnbiasedRNG[528];
            InitCond[1475] = UnbiasedRNG[529];
            InitCond[1476] = UnbiasedRNG[530];
            InitCond[1477] = UnbiasedRNG[531];
            InitCond[1478] = UnbiasedRNG[532];
            InitCond[1479] = UnbiasedRNG[533];
            InitCond[1480] = UnbiasedRNG[534];
            InitCond[1481] = UnbiasedRNG[535];
            InitCond[1482] = UnbiasedRNG[536];
            InitCond[1483] = UnbiasedRNG[537];
            InitCond[1484] = UnbiasedRNG[538];
            InitCond[1485] = UnbiasedRNG[539];
            InitCond[1486] = UnbiasedRNG[540];
            InitCond[1487] = UnbiasedRNG[541];
            InitCond[1488] = UnbiasedRNG[542];
            InitCond[1489] = UnbiasedRNG[543];
            InitCond[1490] = UnbiasedRNG[544];
            InitCond[1491] = UnbiasedRNG[545];
            InitCond[1492] = UnbiasedRNG[546];
            InitCond[1493] = UnbiasedRNG[547];
            InitCond[1494] = UnbiasedRNG[548];
            InitCond[1495] = UnbiasedRNG[549];
            InitCond[1496] = UnbiasedRNG[550];
            InitCond[1497] = UnbiasedRNG[551];
            InitCond[1498] = UnbiasedRNG[552];
            InitCond[1499] = UnbiasedRNG[553];
            InitCond[1500] = UnbiasedRNG[554];
            InitCond[1501] = UnbiasedRNG[555];
            InitCond[1502] = UnbiasedRNG[556];
            InitCond[1503] = UnbiasedRNG[557];
            InitCond[1504] = UnbiasedRNG[558];
            InitCond[1505] = UnbiasedRNG[559];
            InitCond[1506] = UnbiasedRNG[560];
            InitCond[1507] = UnbiasedRNG[561];
            InitCond[1508] = UnbiasedRNG[562];
            InitCond[1509] = UnbiasedRNG[563];
            InitCond[1510] = UnbiasedRNG[564];
            InitCond[1511] = UnbiasedRNG[565];
            InitCond[1512] = UnbiasedRNG[566];
            InitCond[1513] = UnbiasedRNG[567];
            InitCond[1514] = UnbiasedRNG[568];
            InitCond[1515] = UnbiasedRNG[569];
            InitCond[1516] = UnbiasedRNG[570];
            InitCond[1517] = UnbiasedRNG[571];
            InitCond[1518] = UnbiasedRNG[572];
            InitCond[1519] = UnbiasedRNG[573];
            InitCond[1520] = UnbiasedRNG[574];
            InitCond[1521] = UnbiasedRNG[575];
            InitCond[1522] = UnbiasedRNG[576];
            InitCond[1523] = UnbiasedRNG[577];
            InitCond[1524] = UnbiasedRNG[578];
            InitCond[1525] = UnbiasedRNG[579];
            InitCond[1526] = UnbiasedRNG[580];
            InitCond[1527] = UnbiasedRNG[581];
            InitCond[1528] = UnbiasedRNG[582];
            InitCond[1529] = UnbiasedRNG[583];
            InitCond[1530] = UnbiasedRNG[584];
            InitCond[1531] = UnbiasedRNG[585];
            InitCond[1532] = UnbiasedRNG[586];
            InitCond[1533] = UnbiasedRNG[587];
            InitCond[1534] = UnbiasedRNG[588];
            InitCond[1535] = UnbiasedRNG[589];
            InitCond[1536] = UnbiasedRNG[590];
            InitCond[1537] = UnbiasedRNG[591];
            InitCond[1538] = UnbiasedRNG[592];
            InitCond[1539] = UnbiasedRNG[593];
            InitCond[1540] = UnbiasedRNG[594];
            InitCond[1541] = UnbiasedRNG[595];
            InitCond[1542] = UnbiasedRNG[596];
            InitCond[1543] = UnbiasedRNG[597];
            InitCond[1544] = UnbiasedRNG[598];
            InitCond[1545] = UnbiasedRNG[599];
            InitCond[1546] = UnbiasedRNG[600];
            InitCond[1547] = UnbiasedRNG[601];
            InitCond[1548] = UnbiasedRNG[602];
            InitCond[1549] = UnbiasedRNG[603];
            InitCond[1550] = UnbiasedRNG[604];
            InitCond[1551] = UnbiasedRNG[605];
            InitCond[1552] = UnbiasedRNG[606];
            InitCond[1553] = UnbiasedRNG[607];
            InitCond[1554] = UnbiasedRNG[608];
            InitCond[1555] = UnbiasedRNG[609];
            InitCond[1556] = UnbiasedRNG[610];
            InitCond[1557] = UnbiasedRNG[611];
            InitCond[1558] = UnbiasedRNG[612];
            InitCond[1559] = UnbiasedRNG[613];
            InitCond[1560] = UnbiasedRNG[614];
            InitCond[1561] = UnbiasedRNG[615];
            InitCond[1562] = UnbiasedRNG[616];
            InitCond[1563] = UnbiasedRNG[617];
            InitCond[1564] = UnbiasedRNG[618];
            InitCond[1565] = UnbiasedRNG[619];
            InitCond[1566] = UnbiasedRNG[620];
            InitCond[1567] = UnbiasedRNG[621];
            InitCond[1568] = UnbiasedRNG[622];
            InitCond[1569] = UnbiasedRNG[623];
            InitCond[1570] = UnbiasedRNG[624];
            InitCond[1571] = UnbiasedRNG[625];
            InitCond[1572] = UnbiasedRNG[626];
            InitCond[1573] = UnbiasedRNG[627];
            InitCond[1574] = UnbiasedRNG[628];
            InitCond[1575] = UnbiasedRNG[629];
            InitCond[1576] = UnbiasedRNG[630];
            InitCond[1577] = UnbiasedRNG[631];
            InitCond[1578] = UnbiasedRNG[632];
            InitCond[1579] = UnbiasedRNG[633];
            InitCond[1580] = UnbiasedRNG[634];
            InitCond[1581] = UnbiasedRNG[635];
            InitCond[1582] = UnbiasedRNG[636];
            InitCond[1583] = UnbiasedRNG[637];
            InitCond[1584] = UnbiasedRNG[638];
            InitCond[1585] = UnbiasedRNG[639];
            InitCond[1586] = UnbiasedRNG[640];
            InitCond[1587] = UnbiasedRNG[641];
            InitCond[1588] = UnbiasedRNG[642];
            InitCond[1589] = UnbiasedRNG[643];
            InitCond[1590] = UnbiasedRNG[644];
            InitCond[1591] = UnbiasedRNG[645];
            InitCond[1592] = UnbiasedRNG[646];
            InitCond[1593] = UnbiasedRNG[647];
            InitCond[1594] = UnbiasedRNG[648];
            InitCond[1595] = UnbiasedRNG[649];
            InitCond[1596] = UnbiasedRNG[650];
            InitCond[1597] = UnbiasedRNG[651];
            InitCond[1598] = UnbiasedRNG[652];
            InitCond[1599] = UnbiasedRNG[653];
            InitCond[1600] = UnbiasedRNG[654];
            InitCond[1601] = UnbiasedRNG[655];
            InitCond[1602] = UnbiasedRNG[656];
            InitCond[1603] = UnbiasedRNG[657];
            InitCond[1604] = UnbiasedRNG[658];
            InitCond[1605] = UnbiasedRNG[659];
            InitCond[1606] = UnbiasedRNG[660];
            InitCond[1607] = UnbiasedRNG[661];
            InitCond[1608] = UnbiasedRNG[662];
            InitCond[1609] = UnbiasedRNG[663];
            InitCond[1610] = UnbiasedRNG[664];
            InitCond[1611] = UnbiasedRNG[665];
            InitCond[1612] = UnbiasedRNG[666];
            InitCond[1613] = UnbiasedRNG[667];
            InitCond[1614] = UnbiasedRNG[668];
            InitCond[1615] = UnbiasedRNG[669];
            InitCond[1616] = UnbiasedRNG[670];
            InitCond[1617] = UnbiasedRNG[671];
            InitCond[1618] = UnbiasedRNG[672];
            InitCond[1619] = UnbiasedRNG[673];
            InitCond[1620] = UnbiasedRNG[674];
            InitCond[1621] = UnbiasedRNG[675];
            InitCond[1622] = UnbiasedRNG[676];
            InitCond[1623] = UnbiasedRNG[677];
            InitCond[1624] = UnbiasedRNG[678];
            InitCond[1625] = UnbiasedRNG[679];
            InitCond[1626] = UnbiasedRNG[680];
            InitCond[1627] = UnbiasedRNG[681];
            InitCond[1628] = UnbiasedRNG[682];
            InitCond[1629] = UnbiasedRNG[683];
            InitCond[1630] = UnbiasedRNG[684];
            InitCond[1631] = UnbiasedRNG[685];
            InitCond[1632] = UnbiasedRNG[686];
            InitCond[1633] = UnbiasedRNG[687];
            InitCond[1634] = UnbiasedRNG[688];
            InitCond[1635] = UnbiasedRNG[689];
            InitCond[1636] = UnbiasedRNG[690];
            InitCond[1637] = UnbiasedRNG[691];
            InitCond[1638] = UnbiasedRNG[692];
            InitCond[1639] = UnbiasedRNG[693];
            InitCond[1640] = UnbiasedRNG[694];
            InitCond[1641] = UnbiasedRNG[695];
            InitCond[1642] = UnbiasedRNG[696];
            InitCond[1643] = UnbiasedRNG[697];
            InitCond[1644] = UnbiasedRNG[698];
            InitCond[1645] = UnbiasedRNG[699];
            InitCond[1646] = UnbiasedRNG[700];
            InitCond[1647] = UnbiasedRNG[701];
            InitCond[1648] = UnbiasedRNG[702];
            InitCond[1649] = UnbiasedRNG[703];
            InitCond[1650] = UnbiasedRNG[704];
            InitCond[1651] = UnbiasedRNG[705];
            InitCond[1652] = UnbiasedRNG[706];
            InitCond[1653] = UnbiasedRNG[707];
            InitCond[1654] = UnbiasedRNG[708];
            InitCond[1655] = UnbiasedRNG[709];
            InitCond[1656] = UnbiasedRNG[710];
            InitCond[1657] = UnbiasedRNG[711];
            InitCond[1658] = UnbiasedRNG[712];
            InitCond[1659] = UnbiasedRNG[713];
            InitCond[1660] = UnbiasedRNG[714];
            InitCond[1661] = UnbiasedRNG[715];
            InitCond[1662] = UnbiasedRNG[716];
            InitCond[1663] = UnbiasedRNG[717];
            InitCond[1664] = UnbiasedRNG[718];
            InitCond[1665] = UnbiasedRNG[719];
            InitCond[1666] = UnbiasedRNG[720];
            InitCond[1667] = UnbiasedRNG[721];
            InitCond[1668] = UnbiasedRNG[722];
            InitCond[1669] = UnbiasedRNG[723];
            InitCond[1670] = UnbiasedRNG[724];
            InitCond[1671] = UnbiasedRNG[725];
            InitCond[1672] = UnbiasedRNG[726];
            InitCond[1673] = UnbiasedRNG[727];
            InitCond[1674] = UnbiasedRNG[728];
            InitCond[1675] = UnbiasedRNG[729];
            InitCond[1676] = UnbiasedRNG[730];
            InitCond[1677] = UnbiasedRNG[731];
            InitCond[1678] = UnbiasedRNG[732];
            InitCond[1679] = UnbiasedRNG[733];
            InitCond[1680] = UnbiasedRNG[734];
            InitCond[1681] = UnbiasedRNG[735];
            InitCond[1682] = UnbiasedRNG[736];
            InitCond[1683] = UnbiasedRNG[737];
            InitCond[1684] = UnbiasedRNG[738];
            InitCond[1685] = UnbiasedRNG[739];
            InitCond[1686] = UnbiasedRNG[740];
            InitCond[1687] = UnbiasedRNG[741];
            InitCond[1688] = UnbiasedRNG[742];
            InitCond[1689] = UnbiasedRNG[743];
            InitCond[1690] = UnbiasedRNG[744];
            InitCond[1691] = UnbiasedRNG[745];
            InitCond[1692] = UnbiasedRNG[746];
            InitCond[1693] = UnbiasedRNG[747];
            InitCond[1694] = UnbiasedRNG[748];
            InitCond[1695] = UnbiasedRNG[749];
            InitCond[1696] = UnbiasedRNG[750];
            InitCond[1697] = UnbiasedRNG[751];
            InitCond[1698] = UnbiasedRNG[752];
            InitCond[1699] = UnbiasedRNG[753];
            InitCond[1700] = UnbiasedRNG[754];
            InitCond[1701] = UnbiasedRNG[755];
            InitCond[1702] = UnbiasedRNG[756];
            InitCond[1703] = UnbiasedRNG[757];
            InitCond[1704] = UnbiasedRNG[758];
            InitCond[1705] = UnbiasedRNG[759];
            InitCond[1706] = UnbiasedRNG[760];
            InitCond[1707] = UnbiasedRNG[761];
            InitCond[1708] = UnbiasedRNG[762];
            InitCond[1709] = UnbiasedRNG[763];
            InitCond[1710] = UnbiasedRNG[764];
            InitCond[1711] = UnbiasedRNG[765];
            InitCond[1712] = UnbiasedRNG[766];
            InitCond[1713] = UnbiasedRNG[767];
            InitCond[1714] = UnbiasedRNG[768];
            InitCond[1715] = UnbiasedRNG[769];
            InitCond[1716] = UnbiasedRNG[770];
            InitCond[1717] = UnbiasedRNG[771];
            InitCond[1718] = UnbiasedRNG[772];
            InitCond[1719] = UnbiasedRNG[773];
            InitCond[1720] = UnbiasedRNG[774];
            InitCond[1721] = UnbiasedRNG[775];
            InitCond[1722] = UnbiasedRNG[776];
            InitCond[1723] = UnbiasedRNG[777];
            InitCond[1724] = UnbiasedRNG[778];
            InitCond[1725] = UnbiasedRNG[779];
            InitCond[1726] = UnbiasedRNG[780];
            InitCond[1727] = UnbiasedRNG[781];
            InitCond[1728] = UnbiasedRNG[782];
            InitCond[1729] = UnbiasedRNG[783];
            InitCond[1730] = UnbiasedRNG[784];
            InitCond[1731] = UnbiasedRNG[785];
            InitCond[1732] = UnbiasedRNG[786];
            InitCond[1733] = UnbiasedRNG[787];
            InitCond[1734] = UnbiasedRNG[788];
            InitCond[1735] = UnbiasedRNG[789];
            InitCond[1736] = UnbiasedRNG[790];
            InitCond[1737] = UnbiasedRNG[791];
            InitCond[1738] = UnbiasedRNG[792];
            InitCond[1739] = UnbiasedRNG[793];
            InitCond[1740] = UnbiasedRNG[794];
            InitCond[1741] = UnbiasedRNG[795];
            InitCond[1742] = UnbiasedRNG[796];
            InitCond[1743] = UnbiasedRNG[797];
            InitCond[1744] = UnbiasedRNG[798];
            InitCond[1745] = UnbiasedRNG[799];
            InitCond[1746] = UnbiasedRNG[800];
            InitCond[1747] = UnbiasedRNG[801];
            InitCond[1748] = UnbiasedRNG[802];
            InitCond[1749] = UnbiasedRNG[803];
            InitCond[1750] = UnbiasedRNG[804];
            InitCond[1751] = UnbiasedRNG[805];
            InitCond[1752] = UnbiasedRNG[806];
            InitCond[1753] = UnbiasedRNG[807];
            InitCond[1754] = UnbiasedRNG[808];
            InitCond[1755] = UnbiasedRNG[809];
            InitCond[1756] = UnbiasedRNG[810];
            InitCond[1757] = UnbiasedRNG[811];
            InitCond[1758] = UnbiasedRNG[812];
            InitCond[1759] = UnbiasedRNG[813];
            InitCond[1760] = UnbiasedRNG[814];
            InitCond[1761] = UnbiasedRNG[815];
            InitCond[1762] = UnbiasedRNG[816];
            InitCond[1763] = UnbiasedRNG[817];
            InitCond[1764] = UnbiasedRNG[818];
            InitCond[1765] = UnbiasedRNG[819];
            InitCond[1766] = UnbiasedRNG[820];
            InitCond[1767] = UnbiasedRNG[821];
            InitCond[1768] = UnbiasedRNG[822];
            InitCond[1769] = UnbiasedRNG[823];
            InitCond[1770] = UnbiasedRNG[824];
            InitCond[1771] = UnbiasedRNG[825];
            InitCond[1772] = UnbiasedRNG[826];
            InitCond[1773] = UnbiasedRNG[827];
            InitCond[1774] = UnbiasedRNG[828];
            InitCond[1775] = UnbiasedRNG[829];
            InitCond[1776] = UnbiasedRNG[830];
            InitCond[1777] = UnbiasedRNG[831];
            InitCond[1778] = UnbiasedRNG[832];
            InitCond[1779] = UnbiasedRNG[833];
            InitCond[1780] = UnbiasedRNG[834];
            InitCond[1781] = UnbiasedRNG[835];
            InitCond[1782] = UnbiasedRNG[836];
            InitCond[1783] = UnbiasedRNG[837];
            InitCond[1784] = UnbiasedRNG[838];
            InitCond[1785] = UnbiasedRNG[839];
            InitCond[1786] = UnbiasedRNG[840];
            InitCond[1787] = UnbiasedRNG[841];
            InitCond[1788] = UnbiasedRNG[842];
            InitCond[1789] = UnbiasedRNG[843];
            InitCond[1790] = UnbiasedRNG[844];
            InitCond[1791] = UnbiasedRNG[845];
            InitCond[1792] = UnbiasedRNG[846];
            InitCond[1793] = UnbiasedRNG[847];
            InitCond[1794] = UnbiasedRNG[848];
            InitCond[1795] = UnbiasedRNG[849];
            InitCond[1796] = UnbiasedRNG[850];
            InitCond[1797] = UnbiasedRNG[851];
            InitCond[1798] = UnbiasedRNG[852];
            InitCond[1799] = UnbiasedRNG[853];
            InitCond[1800] = UnbiasedRNG[854];
            InitCond[1801] = UnbiasedRNG[855];
            InitCond[1802] = UnbiasedRNG[856];
            InitCond[1803] = UnbiasedRNG[857];
            InitCond[1804] = UnbiasedRNG[858];
            InitCond[1805] = UnbiasedRNG[859];
            InitCond[1806] = UnbiasedRNG[860];
            InitCond[1807] = UnbiasedRNG[861];
            InitCond[1808] = UnbiasedRNG[862];
            InitCond[1809] = UnbiasedRNG[863];
            InitCond[1810] = UnbiasedRNG[864];
            InitCond[1811] = UnbiasedRNG[865];
            InitCond[1812] = UnbiasedRNG[866];
            InitCond[1813] = UnbiasedRNG[867];
            InitCond[1814] = UnbiasedRNG[868];
            InitCond[1815] = UnbiasedRNG[869];
            InitCond[1816] = UnbiasedRNG[870];
            InitCond[1817] = UnbiasedRNG[871];
            InitCond[1818] = UnbiasedRNG[872];
            InitCond[1819] = UnbiasedRNG[873];
            InitCond[1820] = UnbiasedRNG[874];
            InitCond[1821] = UnbiasedRNG[875];
            InitCond[1822] = UnbiasedRNG[876];
            InitCond[1823] = UnbiasedRNG[877];
            InitCond[1824] = UnbiasedRNG[878];
            InitCond[1825] = UnbiasedRNG[879];
            InitCond[1826] = UnbiasedRNG[880];
            InitCond[1827] = UnbiasedRNG[881];
            InitCond[1828] = UnbiasedRNG[882];
            InitCond[1829] = UnbiasedRNG[883];
            InitCond[1830] = UnbiasedRNG[884];
            InitCond[1831] = UnbiasedRNG[885];
            InitCond[1832] = UnbiasedRNG[886];
            InitCond[1833] = UnbiasedRNG[887];
            InitCond[1834] = UnbiasedRNG[888];
            InitCond[1835] = UnbiasedRNG[889];
            InitCond[1836] = UnbiasedRNG[890];
            InitCond[1837] = UnbiasedRNG[891];
            InitCond[1838] = UnbiasedRNG[892];
            InitCond[1839] = UnbiasedRNG[893];
            InitCond[1840] = UnbiasedRNG[894];
            InitCond[1841] = UnbiasedRNG[895];
            InitCond[1842] = UnbiasedRNG[896];
            InitCond[1843] = UnbiasedRNG[897];
            InitCond[1844] = UnbiasedRNG[898];
            InitCond[1845] = UnbiasedRNG[899];
            InitCond[1846] = UnbiasedRNG[900];
            InitCond[1847] = UnbiasedRNG[901];
            InitCond[1848] = UnbiasedRNG[902];
            InitCond[1849] = UnbiasedRNG[903];
            InitCond[1850] = UnbiasedRNG[904];
            InitCond[1851] = UnbiasedRNG[905];
            InitCond[1852] = UnbiasedRNG[906];
            InitCond[1853] = UnbiasedRNG[907];
            InitCond[1854] = UnbiasedRNG[908];
            InitCond[1855] = UnbiasedRNG[909];
            InitCond[1856] = UnbiasedRNG[910];
            InitCond[1857] = UnbiasedRNG[911];
            InitCond[1858] = UnbiasedRNG[912];
            InitCond[1859] = UnbiasedRNG[913];
            InitCond[1860] = UnbiasedRNG[914];
            InitCond[1861] = UnbiasedRNG[915];
            InitCond[1862] = UnbiasedRNG[916];
            InitCond[1863] = UnbiasedRNG[917];
            InitCond[1864] = UnbiasedRNG[918];
            InitCond[1865] = UnbiasedRNG[919];
            InitCond[1866] = UnbiasedRNG[920];
            InitCond[1867] = UnbiasedRNG[921];
            InitCond[1868] = UnbiasedRNG[922];
            InitCond[1869] = UnbiasedRNG[923];
            InitCond[1870] = UnbiasedRNG[924];
            InitCond[1871] = UnbiasedRNG[925];
            InitCond[1872] = UnbiasedRNG[926];
            InitCond[1873] = UnbiasedRNG[927];
            InitCond[1874] = UnbiasedRNG[928];
            InitCond[1875] = UnbiasedRNG[929];
            InitCond[1876] = UnbiasedRNG[930];
            InitCond[1877] = UnbiasedRNG[931];
            InitCond[1878] = UnbiasedRNG[932];
            InitCond[1879] = UnbiasedRNG[933];
            InitCond[1880] = UnbiasedRNG[934];
            InitCond[1881] = UnbiasedRNG[935];
            InitCond[1882] = UnbiasedRNG[936];
            InitCond[1883] = UnbiasedRNG[937];
            InitCond[1884] = UnbiasedRNG[938];
            InitCond[1885] = UnbiasedRNG[939];
            InitCond[1886] = UnbiasedRNG[940];
            InitCond[1887] = UnbiasedRNG[941];
            InitCond[1888] = UnbiasedRNG[942];
            InitCond[1889] = UnbiasedRNG[943];
            InitCond[1890] = UnbiasedRNG[944];
            InitCond[1891] = UnbiasedRNG[945];
        end
        else if (counter == 3) begin
            InitCond[1892] = UnbiasedRNG[0];
            InitCond[1893] = UnbiasedRNG[1];
            InitCond[1894] = UnbiasedRNG[2];
            InitCond[1895] = UnbiasedRNG[3];
            InitCond[1896] = UnbiasedRNG[4];
            InitCond[1897] = UnbiasedRNG[5];
            InitCond[1898] = UnbiasedRNG[6];
            InitCond[1899] = UnbiasedRNG[7];
            InitCond[1900] = UnbiasedRNG[8];
            InitCond[1901] = UnbiasedRNG[9];
            InitCond[1902] = UnbiasedRNG[10];
            InitCond[1903] = UnbiasedRNG[11];
            InitCond[1904] = UnbiasedRNG[12];
            InitCond[1905] = UnbiasedRNG[13];
            InitCond[1906] = UnbiasedRNG[14];
            InitCond[1907] = UnbiasedRNG[15];
            InitCond[1908] = UnbiasedRNG[16];
            InitCond[1909] = UnbiasedRNG[17];
            InitCond[1910] = UnbiasedRNG[18];
            InitCond[1911] = UnbiasedRNG[19];
            InitCond[1912] = UnbiasedRNG[20];
            InitCond[1913] = UnbiasedRNG[21];
            InitCond[1914] = UnbiasedRNG[22];
            InitCond[1915] = UnbiasedRNG[23];
            InitCond[1916] = UnbiasedRNG[24];
            InitCond[1917] = UnbiasedRNG[25];
            InitCond[1918] = UnbiasedRNG[26];
            InitCond[1919] = UnbiasedRNG[27];
            InitCond[1920] = UnbiasedRNG[28];
            InitCond[1921] = UnbiasedRNG[29];
            InitCond[1922] = UnbiasedRNG[30];
            InitCond[1923] = UnbiasedRNG[31];
            InitCond[1924] = UnbiasedRNG[32];
            InitCond[1925] = UnbiasedRNG[33];
            InitCond[1926] = UnbiasedRNG[34];
            InitCond[1927] = UnbiasedRNG[35];
            InitCond[1928] = UnbiasedRNG[36];
            InitCond[1929] = UnbiasedRNG[37];
            InitCond[1930] = UnbiasedRNG[38];
            InitCond[1931] = UnbiasedRNG[39];
            InitCond[1932] = UnbiasedRNG[40];
            InitCond[1933] = UnbiasedRNG[41];
            InitCond[1934] = UnbiasedRNG[42];
            InitCond[1935] = UnbiasedRNG[43];
            InitCond[1936] = UnbiasedRNG[44];
            InitCond[1937] = UnbiasedRNG[45];
            InitCond[1938] = UnbiasedRNG[46];
            InitCond[1939] = UnbiasedRNG[47];
            InitCond[1940] = UnbiasedRNG[48];
            InitCond[1941] = UnbiasedRNG[49];
            InitCond[1942] = UnbiasedRNG[50];
            InitCond[1943] = UnbiasedRNG[51];
            InitCond[1944] = UnbiasedRNG[52];
            InitCond[1945] = UnbiasedRNG[53];
            InitCond[1946] = UnbiasedRNG[54];
            InitCond[1947] = UnbiasedRNG[55];
            InitCond[1948] = UnbiasedRNG[56];
            InitCond[1949] = UnbiasedRNG[57];
            InitCond[1950] = UnbiasedRNG[58];
            InitCond[1951] = UnbiasedRNG[59];
            InitCond[1952] = UnbiasedRNG[60];
            InitCond[1953] = UnbiasedRNG[61];
            InitCond[1954] = UnbiasedRNG[62];
            InitCond[1955] = UnbiasedRNG[63];
            InitCond[1956] = UnbiasedRNG[64];
            InitCond[1957] = UnbiasedRNG[65];
            InitCond[1958] = UnbiasedRNG[66];
            InitCond[1959] = UnbiasedRNG[67];
            InitCond[1960] = UnbiasedRNG[68];
            InitCond[1961] = UnbiasedRNG[69];
            InitCond[1962] = UnbiasedRNG[70];
            InitCond[1963] = UnbiasedRNG[71];
            InitCond[1964] = UnbiasedRNG[72];
            InitCond[1965] = UnbiasedRNG[73];
            InitCond[1966] = UnbiasedRNG[74];
            InitCond[1967] = UnbiasedRNG[75];
            InitCond[1968] = UnbiasedRNG[76];
            InitCond[1969] = UnbiasedRNG[77];
            InitCond[1970] = UnbiasedRNG[78];
            InitCond[1971] = UnbiasedRNG[79];
            InitCond[1972] = UnbiasedRNG[80];
            InitCond[1973] = UnbiasedRNG[81];
            InitCond[1974] = UnbiasedRNG[82];
            InitCond[1975] = UnbiasedRNG[83];
            InitCond[1976] = UnbiasedRNG[84];
            InitCond[1977] = UnbiasedRNG[85];
            InitCond[1978] = UnbiasedRNG[86];
            InitCond[1979] = UnbiasedRNG[87];
            InitCond[1980] = UnbiasedRNG[88];
            InitCond[1981] = UnbiasedRNG[89];
            InitCond[1982] = UnbiasedRNG[90];
            InitCond[1983] = UnbiasedRNG[91];
            InitCond[1984] = UnbiasedRNG[92];
            InitCond[1985] = UnbiasedRNG[93];
            InitCond[1986] = UnbiasedRNG[94];
            InitCond[1987] = UnbiasedRNG[95];
            InitCond[1988] = UnbiasedRNG[96];
            InitCond[1989] = UnbiasedRNG[97];
            InitCond[1990] = UnbiasedRNG[98];
            InitCond[1991] = UnbiasedRNG[99];
            InitCond[1992] = UnbiasedRNG[100];
            InitCond[1993] = UnbiasedRNG[101];
            InitCond[1994] = UnbiasedRNG[102];
            InitCond[1995] = UnbiasedRNG[103];
            InitCond[1996] = UnbiasedRNG[104];
            InitCond[1997] = UnbiasedRNG[105];
            InitCond[1998] = UnbiasedRNG[106];
            InitCond[1999] = UnbiasedRNG[107];
            InitCond[2000] = UnbiasedRNG[108];
            InitCond[2001] = UnbiasedRNG[109];
            InitCond[2002] = UnbiasedRNG[110];
            InitCond[2003] = UnbiasedRNG[111];
            InitCond[2004] = UnbiasedRNG[112];
            InitCond[2005] = UnbiasedRNG[113];
            InitCond[2006] = UnbiasedRNG[114];
            InitCond[2007] = UnbiasedRNG[115];
            InitCond[2008] = UnbiasedRNG[116];
            InitCond[2009] = UnbiasedRNG[117];
            InitCond[2010] = UnbiasedRNG[118];
            InitCond[2011] = UnbiasedRNG[119];
            InitCond[2012] = UnbiasedRNG[120];
            InitCond[2013] = UnbiasedRNG[121];
            InitCond[2014] = UnbiasedRNG[122];
            InitCond[2015] = UnbiasedRNG[123];
            InitCond[2016] = UnbiasedRNG[124];
            InitCond[2017] = UnbiasedRNG[125];
            InitCond[2018] = UnbiasedRNG[126];
            InitCond[2019] = UnbiasedRNG[127];
            InitCond[2020] = UnbiasedRNG[128];
            InitCond[2021] = UnbiasedRNG[129];
            InitCond[2022] = UnbiasedRNG[130];
            InitCond[2023] = UnbiasedRNG[131];
            InitCond[2024] = UnbiasedRNG[132];
            InitCond[2025] = UnbiasedRNG[133];
            InitCond[2026] = UnbiasedRNG[134];
            InitCond[2027] = UnbiasedRNG[135];
            InitCond[2028] = UnbiasedRNG[136];
            InitCond[2029] = UnbiasedRNG[137];
            InitCond[2030] = UnbiasedRNG[138];
            InitCond[2031] = UnbiasedRNG[139];
            InitCond[2032] = UnbiasedRNG[140];
            InitCond[2033] = UnbiasedRNG[141];
            InitCond[2034] = UnbiasedRNG[142];
            InitCond[2035] = UnbiasedRNG[143];
            InitCond[2036] = UnbiasedRNG[144];
            InitCond[2037] = UnbiasedRNG[145];
            InitCond[2038] = UnbiasedRNG[146];
            InitCond[2039] = UnbiasedRNG[147];
            InitCond[2040] = UnbiasedRNG[148];
            InitCond[2041] = UnbiasedRNG[149];
            InitCond[2042] = UnbiasedRNG[150];
            InitCond[2043] = UnbiasedRNG[151];
            InitCond[2044] = UnbiasedRNG[152];
            InitCond[2045] = UnbiasedRNG[153];
            InitCond[2046] = UnbiasedRNG[154];
            InitCond[2047] = UnbiasedRNG[155];
            InitCond[2048] = UnbiasedRNG[156];
            InitCond[2049] = UnbiasedRNG[157];
            InitCond[2050] = UnbiasedRNG[158];
            InitCond[2051] = UnbiasedRNG[159];
            InitCond[2052] = UnbiasedRNG[160];
            InitCond[2053] = UnbiasedRNG[161];
            InitCond[2054] = UnbiasedRNG[162];
            InitCond[2055] = UnbiasedRNG[163];
            InitCond[2056] = UnbiasedRNG[164];
            InitCond[2057] = UnbiasedRNG[165];
            InitCond[2058] = UnbiasedRNG[166];
            InitCond[2059] = UnbiasedRNG[167];
            InitCond[2060] = UnbiasedRNG[168];
            InitCond[2061] = UnbiasedRNG[169];
            InitCond[2062] = UnbiasedRNG[170];
            InitCond[2063] = UnbiasedRNG[171];
            InitCond[2064] = UnbiasedRNG[172];
            InitCond[2065] = UnbiasedRNG[173];
            InitCond[2066] = UnbiasedRNG[174];
            InitCond[2067] = UnbiasedRNG[175];
            InitCond[2068] = UnbiasedRNG[176];
            InitCond[2069] = UnbiasedRNG[177];
            InitCond[2070] = UnbiasedRNG[178];
            InitCond[2071] = UnbiasedRNG[179];
            InitCond[2072] = UnbiasedRNG[180];
            InitCond[2073] = UnbiasedRNG[181];
            InitCond[2074] = UnbiasedRNG[182];
            InitCond[2075] = UnbiasedRNG[183];
            InitCond[2076] = UnbiasedRNG[184];
            InitCond[2077] = UnbiasedRNG[185];
            InitCond[2078] = UnbiasedRNG[186];
            InitCond[2079] = UnbiasedRNG[187];
        end
        else if (counter==5)
            run = 1'b1;
        counter = counter+38'b1;
        solution = {m[15],m[14],m[13],m[12],m[11],m[10],m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[31],m[30],m[29],m[28],m[27],m[26],m[25],m[24],m[23],m[22],m[21],m[20],m[19],m[18],m[17],m[16]};
    end else begin 
        counter = 38'b0;
        failure = 1'b1;
        run = 1'b0;
    end
end

//To measure on only the last step using ILA:
always @(negedge sample_clk) begin
    if (solution_flag)
        solution_flag = 1'b0;
    else if ((run & (solution == solution_check)) | failure)
        solution_flag = 1'b1;
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = run?((((m[32]&m[33]&~m[34]&~m[35])|(m[32]&~m[33]&m[34]&~m[35])|(~m[32]&m[33]&m[34]&~m[35])|(m[32]&~m[33]&~m[34]&m[35])|(~m[32]&m[33]&~m[34]&m[35])|(~m[32]&~m[33]&m[34]&m[35]))&UnbiasedRNG[0])|((m[32]&m[33]&m[34]&~m[35])|(m[32]&m[33]&~m[34]&m[35])|(m[32]&~m[33]&m[34]&m[35])|(~m[32]&m[33]&m[34]&m[35])|(m[32]&m[33]&m[34]&m[35]))):InitCond[0];
    m[1] = run?((((m[36]&m[37]&~m[38]&~m[39])|(m[36]&~m[37]&m[38]&~m[39])|(~m[36]&m[37]&m[38]&~m[39])|(m[36]&~m[37]&~m[38]&m[39])|(~m[36]&m[37]&~m[38]&m[39])|(~m[36]&~m[37]&m[38]&m[39]))&UnbiasedRNG[1])|((m[36]&m[37]&m[38]&~m[39])|(m[36]&m[37]&~m[38]&m[39])|(m[36]&~m[37]&m[38]&m[39])|(~m[36]&m[37]&m[38]&m[39])|(m[36]&m[37]&m[38]&m[39]))):InitCond[1];
    m[2] = run?((((m[40]&m[41]&~m[42]&~m[43])|(m[40]&~m[41]&m[42]&~m[43])|(~m[40]&m[41]&m[42]&~m[43])|(m[40]&~m[41]&~m[42]&m[43])|(~m[40]&m[41]&~m[42]&m[43])|(~m[40]&~m[41]&m[42]&m[43]))&UnbiasedRNG[2])|((m[40]&m[41]&m[42]&~m[43])|(m[40]&m[41]&~m[42]&m[43])|(m[40]&~m[41]&m[42]&m[43])|(~m[40]&m[41]&m[42]&m[43])|(m[40]&m[41]&m[42]&m[43]))):InitCond[2];
    m[3] = run?((((m[44]&m[45]&~m[46]&~m[47])|(m[44]&~m[45]&m[46]&~m[47])|(~m[44]&m[45]&m[46]&~m[47])|(m[44]&~m[45]&~m[46]&m[47])|(~m[44]&m[45]&~m[46]&m[47])|(~m[44]&~m[45]&m[46]&m[47]))&UnbiasedRNG[3])|((m[44]&m[45]&m[46]&~m[47])|(m[44]&m[45]&~m[46]&m[47])|(m[44]&~m[45]&m[46]&m[47])|(~m[44]&m[45]&m[46]&m[47])|(m[44]&m[45]&m[46]&m[47]))):InitCond[3];
    m[4] = run?((((m[48]&m[49]&~m[50]&~m[51])|(m[48]&~m[49]&m[50]&~m[51])|(~m[48]&m[49]&m[50]&~m[51])|(m[48]&~m[49]&~m[50]&m[51])|(~m[48]&m[49]&~m[50]&m[51])|(~m[48]&~m[49]&m[50]&m[51]))&UnbiasedRNG[4])|((m[48]&m[49]&m[50]&~m[51])|(m[48]&m[49]&~m[50]&m[51])|(m[48]&~m[49]&m[50]&m[51])|(~m[48]&m[49]&m[50]&m[51])|(m[48]&m[49]&m[50]&m[51]))):InitCond[4];
    m[5] = run?((((m[52]&m[53]&~m[54]&~m[55])|(m[52]&~m[53]&m[54]&~m[55])|(~m[52]&m[53]&m[54]&~m[55])|(m[52]&~m[53]&~m[54]&m[55])|(~m[52]&m[53]&~m[54]&m[55])|(~m[52]&~m[53]&m[54]&m[55]))&UnbiasedRNG[5])|((m[52]&m[53]&m[54]&~m[55])|(m[52]&m[53]&~m[54]&m[55])|(m[52]&~m[53]&m[54]&m[55])|(~m[52]&m[53]&m[54]&m[55])|(m[52]&m[53]&m[54]&m[55]))):InitCond[5];
    m[6] = run?((((m[56]&m[57]&~m[58]&~m[59])|(m[56]&~m[57]&m[58]&~m[59])|(~m[56]&m[57]&m[58]&~m[59])|(m[56]&~m[57]&~m[58]&m[59])|(~m[56]&m[57]&~m[58]&m[59])|(~m[56]&~m[57]&m[58]&m[59]))&UnbiasedRNG[6])|((m[56]&m[57]&m[58]&~m[59])|(m[56]&m[57]&~m[58]&m[59])|(m[56]&~m[57]&m[58]&m[59])|(~m[56]&m[57]&m[58]&m[59])|(m[56]&m[57]&m[58]&m[59]))):InitCond[6];
    m[7] = run?((((m[60]&m[61]&~m[62]&~m[63])|(m[60]&~m[61]&m[62]&~m[63])|(~m[60]&m[61]&m[62]&~m[63])|(m[60]&~m[61]&~m[62]&m[63])|(~m[60]&m[61]&~m[62]&m[63])|(~m[60]&~m[61]&m[62]&m[63]))&UnbiasedRNG[7])|((m[60]&m[61]&m[62]&~m[63])|(m[60]&m[61]&~m[62]&m[63])|(m[60]&~m[61]&m[62]&m[63])|(~m[60]&m[61]&m[62]&m[63])|(m[60]&m[61]&m[62]&m[63]))):InitCond[7];
    m[8] = run?((((m[64]&m[65]&~m[66]&~m[67])|(m[64]&~m[65]&m[66]&~m[67])|(~m[64]&m[65]&m[66]&~m[67])|(m[64]&~m[65]&~m[66]&m[67])|(~m[64]&m[65]&~m[66]&m[67])|(~m[64]&~m[65]&m[66]&m[67]))&UnbiasedRNG[8])|((m[64]&m[65]&m[66]&~m[67])|(m[64]&m[65]&~m[66]&m[67])|(m[64]&~m[65]&m[66]&m[67])|(~m[64]&m[65]&m[66]&m[67])|(m[64]&m[65]&m[66]&m[67]))):InitCond[8];
    m[9] = run?((((m[68]&m[69]&~m[70]&~m[71])|(m[68]&~m[69]&m[70]&~m[71])|(~m[68]&m[69]&m[70]&~m[71])|(m[68]&~m[69]&~m[70]&m[71])|(~m[68]&m[69]&~m[70]&m[71])|(~m[68]&~m[69]&m[70]&m[71]))&UnbiasedRNG[9])|((m[68]&m[69]&m[70]&~m[71])|(m[68]&m[69]&~m[70]&m[71])|(m[68]&~m[69]&m[70]&m[71])|(~m[68]&m[69]&m[70]&m[71])|(m[68]&m[69]&m[70]&m[71]))):InitCond[9];
    m[10] = run?((((m[72]&m[73]&~m[74]&~m[75])|(m[72]&~m[73]&m[74]&~m[75])|(~m[72]&m[73]&m[74]&~m[75])|(m[72]&~m[73]&~m[74]&m[75])|(~m[72]&m[73]&~m[74]&m[75])|(~m[72]&~m[73]&m[74]&m[75]))&UnbiasedRNG[10])|((m[72]&m[73]&m[74]&~m[75])|(m[72]&m[73]&~m[74]&m[75])|(m[72]&~m[73]&m[74]&m[75])|(~m[72]&m[73]&m[74]&m[75])|(m[72]&m[73]&m[74]&m[75]))):InitCond[10];
    m[11] = run?((((m[76]&m[77]&~m[78]&~m[79])|(m[76]&~m[77]&m[78]&~m[79])|(~m[76]&m[77]&m[78]&~m[79])|(m[76]&~m[77]&~m[78]&m[79])|(~m[76]&m[77]&~m[78]&m[79])|(~m[76]&~m[77]&m[78]&m[79]))&UnbiasedRNG[11])|((m[76]&m[77]&m[78]&~m[79])|(m[76]&m[77]&~m[78]&m[79])|(m[76]&~m[77]&m[78]&m[79])|(~m[76]&m[77]&m[78]&m[79])|(m[76]&m[77]&m[78]&m[79]))):InitCond[11];
    m[12] = run?((((m[80]&m[81]&~m[82]&~m[83])|(m[80]&~m[81]&m[82]&~m[83])|(~m[80]&m[81]&m[82]&~m[83])|(m[80]&~m[81]&~m[82]&m[83])|(~m[80]&m[81]&~m[82]&m[83])|(~m[80]&~m[81]&m[82]&m[83]))&UnbiasedRNG[12])|((m[80]&m[81]&m[82]&~m[83])|(m[80]&m[81]&~m[82]&m[83])|(m[80]&~m[81]&m[82]&m[83])|(~m[80]&m[81]&m[82]&m[83])|(m[80]&m[81]&m[82]&m[83]))):InitCond[12];
    m[13] = run?((((m[84]&m[85]&~m[86]&~m[87])|(m[84]&~m[85]&m[86]&~m[87])|(~m[84]&m[85]&m[86]&~m[87])|(m[84]&~m[85]&~m[86]&m[87])|(~m[84]&m[85]&~m[86]&m[87])|(~m[84]&~m[85]&m[86]&m[87]))&UnbiasedRNG[13])|((m[84]&m[85]&m[86]&~m[87])|(m[84]&m[85]&~m[86]&m[87])|(m[84]&~m[85]&m[86]&m[87])|(~m[84]&m[85]&m[86]&m[87])|(m[84]&m[85]&m[86]&m[87]))):InitCond[13];
    m[14] = run?((((m[88]&m[89]&~m[90]&~m[91])|(m[88]&~m[89]&m[90]&~m[91])|(~m[88]&m[89]&m[90]&~m[91])|(m[88]&~m[89]&~m[90]&m[91])|(~m[88]&m[89]&~m[90]&m[91])|(~m[88]&~m[89]&m[90]&m[91]))&UnbiasedRNG[14])|((m[88]&m[89]&m[90]&~m[91])|(m[88]&m[89]&~m[90]&m[91])|(m[88]&~m[89]&m[90]&m[91])|(~m[88]&m[89]&m[90]&m[91])|(m[88]&m[89]&m[90]&m[91]))):InitCond[14];
    m[15] = run?((((m[92]&m[93]&~m[94]&~m[95])|(m[92]&~m[93]&m[94]&~m[95])|(~m[92]&m[93]&m[94]&~m[95])|(m[92]&~m[93]&~m[94]&m[95])|(~m[92]&m[93]&~m[94]&m[95])|(~m[92]&~m[93]&m[94]&m[95]))&UnbiasedRNG[15])|((m[92]&m[93]&m[94]&~m[95])|(m[92]&m[93]&~m[94]&m[95])|(m[92]&~m[93]&m[94]&m[95])|(~m[92]&m[93]&m[94]&m[95])|(m[92]&m[93]&m[94]&m[95]))):InitCond[15];
    m[16] = run?((((m[96]&m[97]&~m[98]&~m[99])|(m[96]&~m[97]&m[98]&~m[99])|(~m[96]&m[97]&m[98]&~m[99])|(m[96]&~m[97]&~m[98]&m[99])|(~m[96]&m[97]&~m[98]&m[99])|(~m[96]&~m[97]&m[98]&m[99]))&UnbiasedRNG[16])|((m[96]&m[97]&m[98]&~m[99])|(m[96]&m[97]&~m[98]&m[99])|(m[96]&~m[97]&m[98]&m[99])|(~m[96]&m[97]&m[98]&m[99])|(m[96]&m[97]&m[98]&m[99]))):InitCond[16];
    m[17] = run?((((m[100]&m[101]&~m[102]&~m[103])|(m[100]&~m[101]&m[102]&~m[103])|(~m[100]&m[101]&m[102]&~m[103])|(m[100]&~m[101]&~m[102]&m[103])|(~m[100]&m[101]&~m[102]&m[103])|(~m[100]&~m[101]&m[102]&m[103]))&UnbiasedRNG[17])|((m[100]&m[101]&m[102]&~m[103])|(m[100]&m[101]&~m[102]&m[103])|(m[100]&~m[101]&m[102]&m[103])|(~m[100]&m[101]&m[102]&m[103])|(m[100]&m[101]&m[102]&m[103]))):InitCond[17];
    m[18] = run?((((m[104]&m[105]&~m[106]&~m[107])|(m[104]&~m[105]&m[106]&~m[107])|(~m[104]&m[105]&m[106]&~m[107])|(m[104]&~m[105]&~m[106]&m[107])|(~m[104]&m[105]&~m[106]&m[107])|(~m[104]&~m[105]&m[106]&m[107]))&UnbiasedRNG[18])|((m[104]&m[105]&m[106]&~m[107])|(m[104]&m[105]&~m[106]&m[107])|(m[104]&~m[105]&m[106]&m[107])|(~m[104]&m[105]&m[106]&m[107])|(m[104]&m[105]&m[106]&m[107]))):InitCond[18];
    m[19] = run?((((m[108]&m[109]&~m[110]&~m[111])|(m[108]&~m[109]&m[110]&~m[111])|(~m[108]&m[109]&m[110]&~m[111])|(m[108]&~m[109]&~m[110]&m[111])|(~m[108]&m[109]&~m[110]&m[111])|(~m[108]&~m[109]&m[110]&m[111]))&UnbiasedRNG[19])|((m[108]&m[109]&m[110]&~m[111])|(m[108]&m[109]&~m[110]&m[111])|(m[108]&~m[109]&m[110]&m[111])|(~m[108]&m[109]&m[110]&m[111])|(m[108]&m[109]&m[110]&m[111]))):InitCond[19];
    m[20] = run?((((m[112]&m[113]&~m[114]&~m[115])|(m[112]&~m[113]&m[114]&~m[115])|(~m[112]&m[113]&m[114]&~m[115])|(m[112]&~m[113]&~m[114]&m[115])|(~m[112]&m[113]&~m[114]&m[115])|(~m[112]&~m[113]&m[114]&m[115]))&UnbiasedRNG[20])|((m[112]&m[113]&m[114]&~m[115])|(m[112]&m[113]&~m[114]&m[115])|(m[112]&~m[113]&m[114]&m[115])|(~m[112]&m[113]&m[114]&m[115])|(m[112]&m[113]&m[114]&m[115]))):InitCond[20];
    m[21] = run?((((m[116]&m[117]&~m[118]&~m[119])|(m[116]&~m[117]&m[118]&~m[119])|(~m[116]&m[117]&m[118]&~m[119])|(m[116]&~m[117]&~m[118]&m[119])|(~m[116]&m[117]&~m[118]&m[119])|(~m[116]&~m[117]&m[118]&m[119]))&UnbiasedRNG[21])|((m[116]&m[117]&m[118]&~m[119])|(m[116]&m[117]&~m[118]&m[119])|(m[116]&~m[117]&m[118]&m[119])|(~m[116]&m[117]&m[118]&m[119])|(m[116]&m[117]&m[118]&m[119]))):InitCond[21];
    m[22] = run?((((m[120]&m[121]&~m[122]&~m[123])|(m[120]&~m[121]&m[122]&~m[123])|(~m[120]&m[121]&m[122]&~m[123])|(m[120]&~m[121]&~m[122]&m[123])|(~m[120]&m[121]&~m[122]&m[123])|(~m[120]&~m[121]&m[122]&m[123]))&UnbiasedRNG[22])|((m[120]&m[121]&m[122]&~m[123])|(m[120]&m[121]&~m[122]&m[123])|(m[120]&~m[121]&m[122]&m[123])|(~m[120]&m[121]&m[122]&m[123])|(m[120]&m[121]&m[122]&m[123]))):InitCond[22];
    m[23] = run?((((m[124]&m[125]&~m[126]&~m[127])|(m[124]&~m[125]&m[126]&~m[127])|(~m[124]&m[125]&m[126]&~m[127])|(m[124]&~m[125]&~m[126]&m[127])|(~m[124]&m[125]&~m[126]&m[127])|(~m[124]&~m[125]&m[126]&m[127]))&UnbiasedRNG[23])|((m[124]&m[125]&m[126]&~m[127])|(m[124]&m[125]&~m[126]&m[127])|(m[124]&~m[125]&m[126]&m[127])|(~m[124]&m[125]&m[126]&m[127])|(m[124]&m[125]&m[126]&m[127]))):InitCond[23];
    m[24] = run?((((m[128]&m[129]&~m[130]&~m[131])|(m[128]&~m[129]&m[130]&~m[131])|(~m[128]&m[129]&m[130]&~m[131])|(m[128]&~m[129]&~m[130]&m[131])|(~m[128]&m[129]&~m[130]&m[131])|(~m[128]&~m[129]&m[130]&m[131]))&UnbiasedRNG[24])|((m[128]&m[129]&m[130]&~m[131])|(m[128]&m[129]&~m[130]&m[131])|(m[128]&~m[129]&m[130]&m[131])|(~m[128]&m[129]&m[130]&m[131])|(m[128]&m[129]&m[130]&m[131]))):InitCond[24];
    m[25] = run?((((m[132]&m[133]&~m[134]&~m[135])|(m[132]&~m[133]&m[134]&~m[135])|(~m[132]&m[133]&m[134]&~m[135])|(m[132]&~m[133]&~m[134]&m[135])|(~m[132]&m[133]&~m[134]&m[135])|(~m[132]&~m[133]&m[134]&m[135]))&UnbiasedRNG[25])|((m[132]&m[133]&m[134]&~m[135])|(m[132]&m[133]&~m[134]&m[135])|(m[132]&~m[133]&m[134]&m[135])|(~m[132]&m[133]&m[134]&m[135])|(m[132]&m[133]&m[134]&m[135]))):InitCond[25];
    m[26] = run?((((m[136]&m[137]&~m[138]&~m[139])|(m[136]&~m[137]&m[138]&~m[139])|(~m[136]&m[137]&m[138]&~m[139])|(m[136]&~m[137]&~m[138]&m[139])|(~m[136]&m[137]&~m[138]&m[139])|(~m[136]&~m[137]&m[138]&m[139]))&UnbiasedRNG[26])|((m[136]&m[137]&m[138]&~m[139])|(m[136]&m[137]&~m[138]&m[139])|(m[136]&~m[137]&m[138]&m[139])|(~m[136]&m[137]&m[138]&m[139])|(m[136]&m[137]&m[138]&m[139]))):InitCond[26];
    m[27] = run?((((m[140]&m[141]&~m[142]&~m[143])|(m[140]&~m[141]&m[142]&~m[143])|(~m[140]&m[141]&m[142]&~m[143])|(m[140]&~m[141]&~m[142]&m[143])|(~m[140]&m[141]&~m[142]&m[143])|(~m[140]&~m[141]&m[142]&m[143]))&UnbiasedRNG[27])|((m[140]&m[141]&m[142]&~m[143])|(m[140]&m[141]&~m[142]&m[143])|(m[140]&~m[141]&m[142]&m[143])|(~m[140]&m[141]&m[142]&m[143])|(m[140]&m[141]&m[142]&m[143]))):InitCond[27];
    m[28] = run?((((m[144]&m[145]&~m[146]&~m[147])|(m[144]&~m[145]&m[146]&~m[147])|(~m[144]&m[145]&m[146]&~m[147])|(m[144]&~m[145]&~m[146]&m[147])|(~m[144]&m[145]&~m[146]&m[147])|(~m[144]&~m[145]&m[146]&m[147]))&UnbiasedRNG[28])|((m[144]&m[145]&m[146]&~m[147])|(m[144]&m[145]&~m[146]&m[147])|(m[144]&~m[145]&m[146]&m[147])|(~m[144]&m[145]&m[146]&m[147])|(m[144]&m[145]&m[146]&m[147]))):InitCond[28];
    m[29] = run?((((m[148]&m[149]&~m[150]&~m[151])|(m[148]&~m[149]&m[150]&~m[151])|(~m[148]&m[149]&m[150]&~m[151])|(m[148]&~m[149]&~m[150]&m[151])|(~m[148]&m[149]&~m[150]&m[151])|(~m[148]&~m[149]&m[150]&m[151]))&UnbiasedRNG[29])|((m[148]&m[149]&m[150]&~m[151])|(m[148]&m[149]&~m[150]&m[151])|(m[148]&~m[149]&m[150]&m[151])|(~m[148]&m[149]&m[150]&m[151])|(m[148]&m[149]&m[150]&m[151]))):InitCond[29];
    m[30] = run?((((m[152]&m[153]&~m[154]&~m[155])|(m[152]&~m[153]&m[154]&~m[155])|(~m[152]&m[153]&m[154]&~m[155])|(m[152]&~m[153]&~m[154]&m[155])|(~m[152]&m[153]&~m[154]&m[155])|(~m[152]&~m[153]&m[154]&m[155]))&UnbiasedRNG[30])|((m[152]&m[153]&m[154]&~m[155])|(m[152]&m[153]&~m[154]&m[155])|(m[152]&~m[153]&m[154]&m[155])|(~m[152]&m[153]&m[154]&m[155])|(m[152]&m[153]&m[154]&m[155]))):InitCond[30];
    m[31] = run?((((m[156]&m[157]&~m[158]&~m[159])|(m[156]&~m[157]&m[158]&~m[159])|(~m[156]&m[157]&m[158]&~m[159])|(m[156]&~m[157]&~m[158]&m[159])|(~m[156]&m[157]&~m[158]&m[159])|(~m[156]&~m[157]&m[158]&m[159]))&UnbiasedRNG[31])|((m[156]&m[157]&m[158]&~m[159])|(m[156]&m[157]&~m[158]&m[159])|(m[156]&~m[157]&m[158]&m[159])|(~m[156]&m[157]&m[158]&m[159])|(m[156]&m[157]&m[158]&m[159]))):InitCond[31];
    m[160] = run?((((~m[32]&~m[416]&~m[672])|(m[32]&m[416]&~m[672]))&BiasedRNG[0])|(((m[32]&~m[416]&~m[672])|(~m[32]&m[416]&m[672]))&~BiasedRNG[0])|((~m[32]&~m[416]&m[672])|(m[32]&~m[416]&m[672])|(m[32]&m[416]&m[672]))):InitCond[32];
    m[161] = run?((((~m[32]&~m[432]&~m[688])|(m[32]&m[432]&~m[688]))&BiasedRNG[1])|(((m[32]&~m[432]&~m[688])|(~m[32]&m[432]&m[688]))&~BiasedRNG[1])|((~m[32]&~m[432]&m[688])|(m[32]&~m[432]&m[688])|(m[32]&m[432]&m[688]))):InitCond[33];
    m[162] = run?((((~m[32]&~m[448]&~m[704])|(m[32]&m[448]&~m[704]))&BiasedRNG[2])|(((m[32]&~m[448]&~m[704])|(~m[32]&m[448]&m[704]))&~BiasedRNG[2])|((~m[32]&~m[448]&m[704])|(m[32]&~m[448]&m[704])|(m[32]&m[448]&m[704]))):InitCond[34];
    m[163] = run?((((~m[32]&~m[464]&~m[720])|(m[32]&m[464]&~m[720]))&BiasedRNG[3])|(((m[32]&~m[464]&~m[720])|(~m[32]&m[464]&m[720]))&~BiasedRNG[3])|((~m[32]&~m[464]&m[720])|(m[32]&~m[464]&m[720])|(m[32]&m[464]&m[720]))):InitCond[35];
    m[164] = run?((((~m[33]&~m[480]&~m[736])|(m[33]&m[480]&~m[736]))&BiasedRNG[4])|(((m[33]&~m[480]&~m[736])|(~m[33]&m[480]&m[736]))&~BiasedRNG[4])|((~m[33]&~m[480]&m[736])|(m[33]&~m[480]&m[736])|(m[33]&m[480]&m[736]))):InitCond[36];
    m[165] = run?((((~m[33]&~m[496]&~m[752])|(m[33]&m[496]&~m[752]))&BiasedRNG[5])|(((m[33]&~m[496]&~m[752])|(~m[33]&m[496]&m[752]))&~BiasedRNG[5])|((~m[33]&~m[496]&m[752])|(m[33]&~m[496]&m[752])|(m[33]&m[496]&m[752]))):InitCond[37];
    m[166] = run?((((~m[33]&~m[512]&~m[768])|(m[33]&m[512]&~m[768]))&BiasedRNG[6])|(((m[33]&~m[512]&~m[768])|(~m[33]&m[512]&m[768]))&~BiasedRNG[6])|((~m[33]&~m[512]&m[768])|(m[33]&~m[512]&m[768])|(m[33]&m[512]&m[768]))):InitCond[38];
    m[167] = run?((((~m[33]&~m[528]&~m[784])|(m[33]&m[528]&~m[784]))&BiasedRNG[7])|(((m[33]&~m[528]&~m[784])|(~m[33]&m[528]&m[784]))&~BiasedRNG[7])|((~m[33]&~m[528]&m[784])|(m[33]&~m[528]&m[784])|(m[33]&m[528]&m[784]))):InitCond[39];
    m[168] = run?((((~m[34]&~m[544]&~m[800])|(m[34]&m[544]&~m[800]))&BiasedRNG[8])|(((m[34]&~m[544]&~m[800])|(~m[34]&m[544]&m[800]))&~BiasedRNG[8])|((~m[34]&~m[544]&m[800])|(m[34]&~m[544]&m[800])|(m[34]&m[544]&m[800]))):InitCond[40];
    m[169] = run?((((~m[34]&~m[560]&~m[816])|(m[34]&m[560]&~m[816]))&BiasedRNG[9])|(((m[34]&~m[560]&~m[816])|(~m[34]&m[560]&m[816]))&~BiasedRNG[9])|((~m[34]&~m[560]&m[816])|(m[34]&~m[560]&m[816])|(m[34]&m[560]&m[816]))):InitCond[41];
    m[170] = run?((((~m[34]&~m[576]&~m[832])|(m[34]&m[576]&~m[832]))&BiasedRNG[10])|(((m[34]&~m[576]&~m[832])|(~m[34]&m[576]&m[832]))&~BiasedRNG[10])|((~m[34]&~m[576]&m[832])|(m[34]&~m[576]&m[832])|(m[34]&m[576]&m[832]))):InitCond[42];
    m[171] = run?((((~m[34]&~m[592]&~m[848])|(m[34]&m[592]&~m[848]))&BiasedRNG[11])|(((m[34]&~m[592]&~m[848])|(~m[34]&m[592]&m[848]))&~BiasedRNG[11])|((~m[34]&~m[592]&m[848])|(m[34]&~m[592]&m[848])|(m[34]&m[592]&m[848]))):InitCond[43];
    m[172] = run?((((~m[35]&~m[608]&~m[864])|(m[35]&m[608]&~m[864]))&BiasedRNG[12])|(((m[35]&~m[608]&~m[864])|(~m[35]&m[608]&m[864]))&~BiasedRNG[12])|((~m[35]&~m[608]&m[864])|(m[35]&~m[608]&m[864])|(m[35]&m[608]&m[864]))):InitCond[44];
    m[173] = run?((((~m[35]&~m[624]&~m[880])|(m[35]&m[624]&~m[880]))&BiasedRNG[13])|(((m[35]&~m[624]&~m[880])|(~m[35]&m[624]&m[880]))&~BiasedRNG[13])|((~m[35]&~m[624]&m[880])|(m[35]&~m[624]&m[880])|(m[35]&m[624]&m[880]))):InitCond[45];
    m[174] = run?((((~m[35]&~m[640]&~m[896])|(m[35]&m[640]&~m[896]))&BiasedRNG[14])|(((m[35]&~m[640]&~m[896])|(~m[35]&m[640]&m[896]))&~BiasedRNG[14])|((~m[35]&~m[640]&m[896])|(m[35]&~m[640]&m[896])|(m[35]&m[640]&m[896]))):InitCond[46];
    m[175] = run?((((~m[35]&~m[656]&~m[912])|(m[35]&m[656]&~m[912]))&BiasedRNG[15])|(((m[35]&~m[656]&~m[912])|(~m[35]&m[656]&m[912]))&~BiasedRNG[15])|((~m[35]&~m[656]&m[912])|(m[35]&~m[656]&m[912])|(m[35]&m[656]&m[912]))):InitCond[47];
    m[176] = run?((((~m[36]&~m[417]&~m[673])|(m[36]&m[417]&~m[673]))&BiasedRNG[16])|(((m[36]&~m[417]&~m[673])|(~m[36]&m[417]&m[673]))&~BiasedRNG[16])|((~m[36]&~m[417]&m[673])|(m[36]&~m[417]&m[673])|(m[36]&m[417]&m[673]))):InitCond[48];
    m[177] = run?((((~m[36]&~m[433]&~m[689])|(m[36]&m[433]&~m[689]))&BiasedRNG[17])|(((m[36]&~m[433]&~m[689])|(~m[36]&m[433]&m[689]))&~BiasedRNG[17])|((~m[36]&~m[433]&m[689])|(m[36]&~m[433]&m[689])|(m[36]&m[433]&m[689]))):InitCond[49];
    m[178] = run?((((~m[36]&~m[449]&~m[705])|(m[36]&m[449]&~m[705]))&BiasedRNG[18])|(((m[36]&~m[449]&~m[705])|(~m[36]&m[449]&m[705]))&~BiasedRNG[18])|((~m[36]&~m[449]&m[705])|(m[36]&~m[449]&m[705])|(m[36]&m[449]&m[705]))):InitCond[50];
    m[179] = run?((((~m[36]&~m[465]&~m[721])|(m[36]&m[465]&~m[721]))&BiasedRNG[19])|(((m[36]&~m[465]&~m[721])|(~m[36]&m[465]&m[721]))&~BiasedRNG[19])|((~m[36]&~m[465]&m[721])|(m[36]&~m[465]&m[721])|(m[36]&m[465]&m[721]))):InitCond[51];
    m[180] = run?((((~m[37]&~m[481]&~m[737])|(m[37]&m[481]&~m[737]))&BiasedRNG[20])|(((m[37]&~m[481]&~m[737])|(~m[37]&m[481]&m[737]))&~BiasedRNG[20])|((~m[37]&~m[481]&m[737])|(m[37]&~m[481]&m[737])|(m[37]&m[481]&m[737]))):InitCond[52];
    m[181] = run?((((~m[37]&~m[497]&~m[753])|(m[37]&m[497]&~m[753]))&BiasedRNG[21])|(((m[37]&~m[497]&~m[753])|(~m[37]&m[497]&m[753]))&~BiasedRNG[21])|((~m[37]&~m[497]&m[753])|(m[37]&~m[497]&m[753])|(m[37]&m[497]&m[753]))):InitCond[53];
    m[182] = run?((((~m[37]&~m[513]&~m[769])|(m[37]&m[513]&~m[769]))&BiasedRNG[22])|(((m[37]&~m[513]&~m[769])|(~m[37]&m[513]&m[769]))&~BiasedRNG[22])|((~m[37]&~m[513]&m[769])|(m[37]&~m[513]&m[769])|(m[37]&m[513]&m[769]))):InitCond[54];
    m[183] = run?((((~m[37]&~m[529]&~m[785])|(m[37]&m[529]&~m[785]))&BiasedRNG[23])|(((m[37]&~m[529]&~m[785])|(~m[37]&m[529]&m[785]))&~BiasedRNG[23])|((~m[37]&~m[529]&m[785])|(m[37]&~m[529]&m[785])|(m[37]&m[529]&m[785]))):InitCond[55];
    m[184] = run?((((~m[38]&~m[545]&~m[801])|(m[38]&m[545]&~m[801]))&BiasedRNG[24])|(((m[38]&~m[545]&~m[801])|(~m[38]&m[545]&m[801]))&~BiasedRNG[24])|((~m[38]&~m[545]&m[801])|(m[38]&~m[545]&m[801])|(m[38]&m[545]&m[801]))):InitCond[56];
    m[185] = run?((((~m[38]&~m[561]&~m[817])|(m[38]&m[561]&~m[817]))&BiasedRNG[25])|(((m[38]&~m[561]&~m[817])|(~m[38]&m[561]&m[817]))&~BiasedRNG[25])|((~m[38]&~m[561]&m[817])|(m[38]&~m[561]&m[817])|(m[38]&m[561]&m[817]))):InitCond[57];
    m[186] = run?((((~m[38]&~m[577]&~m[833])|(m[38]&m[577]&~m[833]))&BiasedRNG[26])|(((m[38]&~m[577]&~m[833])|(~m[38]&m[577]&m[833]))&~BiasedRNG[26])|((~m[38]&~m[577]&m[833])|(m[38]&~m[577]&m[833])|(m[38]&m[577]&m[833]))):InitCond[58];
    m[187] = run?((((~m[38]&~m[593]&~m[849])|(m[38]&m[593]&~m[849]))&BiasedRNG[27])|(((m[38]&~m[593]&~m[849])|(~m[38]&m[593]&m[849]))&~BiasedRNG[27])|((~m[38]&~m[593]&m[849])|(m[38]&~m[593]&m[849])|(m[38]&m[593]&m[849]))):InitCond[59];
    m[188] = run?((((~m[39]&~m[609]&~m[865])|(m[39]&m[609]&~m[865]))&BiasedRNG[28])|(((m[39]&~m[609]&~m[865])|(~m[39]&m[609]&m[865]))&~BiasedRNG[28])|((~m[39]&~m[609]&m[865])|(m[39]&~m[609]&m[865])|(m[39]&m[609]&m[865]))):InitCond[60];
    m[189] = run?((((~m[39]&~m[625]&~m[881])|(m[39]&m[625]&~m[881]))&BiasedRNG[29])|(((m[39]&~m[625]&~m[881])|(~m[39]&m[625]&m[881]))&~BiasedRNG[29])|((~m[39]&~m[625]&m[881])|(m[39]&~m[625]&m[881])|(m[39]&m[625]&m[881]))):InitCond[61];
    m[190] = run?((((~m[39]&~m[641]&~m[897])|(m[39]&m[641]&~m[897]))&BiasedRNG[30])|(((m[39]&~m[641]&~m[897])|(~m[39]&m[641]&m[897]))&~BiasedRNG[30])|((~m[39]&~m[641]&m[897])|(m[39]&~m[641]&m[897])|(m[39]&m[641]&m[897]))):InitCond[62];
    m[191] = run?((((~m[39]&~m[657]&~m[913])|(m[39]&m[657]&~m[913]))&BiasedRNG[31])|(((m[39]&~m[657]&~m[913])|(~m[39]&m[657]&m[913]))&~BiasedRNG[31])|((~m[39]&~m[657]&m[913])|(m[39]&~m[657]&m[913])|(m[39]&m[657]&m[913]))):InitCond[63];
    m[192] = run?((((~m[40]&~m[418]&~m[674])|(m[40]&m[418]&~m[674]))&BiasedRNG[32])|(((m[40]&~m[418]&~m[674])|(~m[40]&m[418]&m[674]))&~BiasedRNG[32])|((~m[40]&~m[418]&m[674])|(m[40]&~m[418]&m[674])|(m[40]&m[418]&m[674]))):InitCond[64];
    m[193] = run?((((~m[40]&~m[434]&~m[690])|(m[40]&m[434]&~m[690]))&BiasedRNG[33])|(((m[40]&~m[434]&~m[690])|(~m[40]&m[434]&m[690]))&~BiasedRNG[33])|((~m[40]&~m[434]&m[690])|(m[40]&~m[434]&m[690])|(m[40]&m[434]&m[690]))):InitCond[65];
    m[194] = run?((((~m[40]&~m[450]&~m[706])|(m[40]&m[450]&~m[706]))&BiasedRNG[34])|(((m[40]&~m[450]&~m[706])|(~m[40]&m[450]&m[706]))&~BiasedRNG[34])|((~m[40]&~m[450]&m[706])|(m[40]&~m[450]&m[706])|(m[40]&m[450]&m[706]))):InitCond[66];
    m[195] = run?((((~m[40]&~m[466]&~m[722])|(m[40]&m[466]&~m[722]))&BiasedRNG[35])|(((m[40]&~m[466]&~m[722])|(~m[40]&m[466]&m[722]))&~BiasedRNG[35])|((~m[40]&~m[466]&m[722])|(m[40]&~m[466]&m[722])|(m[40]&m[466]&m[722]))):InitCond[67];
    m[196] = run?((((~m[41]&~m[482]&~m[738])|(m[41]&m[482]&~m[738]))&BiasedRNG[36])|(((m[41]&~m[482]&~m[738])|(~m[41]&m[482]&m[738]))&~BiasedRNG[36])|((~m[41]&~m[482]&m[738])|(m[41]&~m[482]&m[738])|(m[41]&m[482]&m[738]))):InitCond[68];
    m[197] = run?((((~m[41]&~m[498]&~m[754])|(m[41]&m[498]&~m[754]))&BiasedRNG[37])|(((m[41]&~m[498]&~m[754])|(~m[41]&m[498]&m[754]))&~BiasedRNG[37])|((~m[41]&~m[498]&m[754])|(m[41]&~m[498]&m[754])|(m[41]&m[498]&m[754]))):InitCond[69];
    m[198] = run?((((~m[41]&~m[514]&~m[770])|(m[41]&m[514]&~m[770]))&BiasedRNG[38])|(((m[41]&~m[514]&~m[770])|(~m[41]&m[514]&m[770]))&~BiasedRNG[38])|((~m[41]&~m[514]&m[770])|(m[41]&~m[514]&m[770])|(m[41]&m[514]&m[770]))):InitCond[70];
    m[199] = run?((((~m[41]&~m[530]&~m[786])|(m[41]&m[530]&~m[786]))&BiasedRNG[39])|(((m[41]&~m[530]&~m[786])|(~m[41]&m[530]&m[786]))&~BiasedRNG[39])|((~m[41]&~m[530]&m[786])|(m[41]&~m[530]&m[786])|(m[41]&m[530]&m[786]))):InitCond[71];
    m[200] = run?((((~m[42]&~m[546]&~m[802])|(m[42]&m[546]&~m[802]))&BiasedRNG[40])|(((m[42]&~m[546]&~m[802])|(~m[42]&m[546]&m[802]))&~BiasedRNG[40])|((~m[42]&~m[546]&m[802])|(m[42]&~m[546]&m[802])|(m[42]&m[546]&m[802]))):InitCond[72];
    m[201] = run?((((~m[42]&~m[562]&~m[818])|(m[42]&m[562]&~m[818]))&BiasedRNG[41])|(((m[42]&~m[562]&~m[818])|(~m[42]&m[562]&m[818]))&~BiasedRNG[41])|((~m[42]&~m[562]&m[818])|(m[42]&~m[562]&m[818])|(m[42]&m[562]&m[818]))):InitCond[73];
    m[202] = run?((((~m[42]&~m[578]&~m[834])|(m[42]&m[578]&~m[834]))&BiasedRNG[42])|(((m[42]&~m[578]&~m[834])|(~m[42]&m[578]&m[834]))&~BiasedRNG[42])|((~m[42]&~m[578]&m[834])|(m[42]&~m[578]&m[834])|(m[42]&m[578]&m[834]))):InitCond[74];
    m[203] = run?((((~m[42]&~m[594]&~m[850])|(m[42]&m[594]&~m[850]))&BiasedRNG[43])|(((m[42]&~m[594]&~m[850])|(~m[42]&m[594]&m[850]))&~BiasedRNG[43])|((~m[42]&~m[594]&m[850])|(m[42]&~m[594]&m[850])|(m[42]&m[594]&m[850]))):InitCond[75];
    m[204] = run?((((~m[43]&~m[610]&~m[866])|(m[43]&m[610]&~m[866]))&BiasedRNG[44])|(((m[43]&~m[610]&~m[866])|(~m[43]&m[610]&m[866]))&~BiasedRNG[44])|((~m[43]&~m[610]&m[866])|(m[43]&~m[610]&m[866])|(m[43]&m[610]&m[866]))):InitCond[76];
    m[205] = run?((((~m[43]&~m[626]&~m[882])|(m[43]&m[626]&~m[882]))&BiasedRNG[45])|(((m[43]&~m[626]&~m[882])|(~m[43]&m[626]&m[882]))&~BiasedRNG[45])|((~m[43]&~m[626]&m[882])|(m[43]&~m[626]&m[882])|(m[43]&m[626]&m[882]))):InitCond[77];
    m[206] = run?((((~m[43]&~m[642]&~m[898])|(m[43]&m[642]&~m[898]))&BiasedRNG[46])|(((m[43]&~m[642]&~m[898])|(~m[43]&m[642]&m[898]))&~BiasedRNG[46])|((~m[43]&~m[642]&m[898])|(m[43]&~m[642]&m[898])|(m[43]&m[642]&m[898]))):InitCond[78];
    m[207] = run?((((~m[43]&~m[658]&~m[914])|(m[43]&m[658]&~m[914]))&BiasedRNG[47])|(((m[43]&~m[658]&~m[914])|(~m[43]&m[658]&m[914]))&~BiasedRNG[47])|((~m[43]&~m[658]&m[914])|(m[43]&~m[658]&m[914])|(m[43]&m[658]&m[914]))):InitCond[79];
    m[208] = run?((((~m[44]&~m[419]&~m[675])|(m[44]&m[419]&~m[675]))&BiasedRNG[48])|(((m[44]&~m[419]&~m[675])|(~m[44]&m[419]&m[675]))&~BiasedRNG[48])|((~m[44]&~m[419]&m[675])|(m[44]&~m[419]&m[675])|(m[44]&m[419]&m[675]))):InitCond[80];
    m[209] = run?((((~m[44]&~m[435]&~m[691])|(m[44]&m[435]&~m[691]))&BiasedRNG[49])|(((m[44]&~m[435]&~m[691])|(~m[44]&m[435]&m[691]))&~BiasedRNG[49])|((~m[44]&~m[435]&m[691])|(m[44]&~m[435]&m[691])|(m[44]&m[435]&m[691]))):InitCond[81];
    m[210] = run?((((~m[44]&~m[451]&~m[707])|(m[44]&m[451]&~m[707]))&BiasedRNG[50])|(((m[44]&~m[451]&~m[707])|(~m[44]&m[451]&m[707]))&~BiasedRNG[50])|((~m[44]&~m[451]&m[707])|(m[44]&~m[451]&m[707])|(m[44]&m[451]&m[707]))):InitCond[82];
    m[211] = run?((((~m[44]&~m[467]&~m[723])|(m[44]&m[467]&~m[723]))&BiasedRNG[51])|(((m[44]&~m[467]&~m[723])|(~m[44]&m[467]&m[723]))&~BiasedRNG[51])|((~m[44]&~m[467]&m[723])|(m[44]&~m[467]&m[723])|(m[44]&m[467]&m[723]))):InitCond[83];
    m[212] = run?((((~m[45]&~m[483]&~m[739])|(m[45]&m[483]&~m[739]))&BiasedRNG[52])|(((m[45]&~m[483]&~m[739])|(~m[45]&m[483]&m[739]))&~BiasedRNG[52])|((~m[45]&~m[483]&m[739])|(m[45]&~m[483]&m[739])|(m[45]&m[483]&m[739]))):InitCond[84];
    m[213] = run?((((~m[45]&~m[499]&~m[755])|(m[45]&m[499]&~m[755]))&BiasedRNG[53])|(((m[45]&~m[499]&~m[755])|(~m[45]&m[499]&m[755]))&~BiasedRNG[53])|((~m[45]&~m[499]&m[755])|(m[45]&~m[499]&m[755])|(m[45]&m[499]&m[755]))):InitCond[85];
    m[214] = run?((((~m[45]&~m[515]&~m[771])|(m[45]&m[515]&~m[771]))&BiasedRNG[54])|(((m[45]&~m[515]&~m[771])|(~m[45]&m[515]&m[771]))&~BiasedRNG[54])|((~m[45]&~m[515]&m[771])|(m[45]&~m[515]&m[771])|(m[45]&m[515]&m[771]))):InitCond[86];
    m[215] = run?((((~m[45]&~m[531]&~m[787])|(m[45]&m[531]&~m[787]))&BiasedRNG[55])|(((m[45]&~m[531]&~m[787])|(~m[45]&m[531]&m[787]))&~BiasedRNG[55])|((~m[45]&~m[531]&m[787])|(m[45]&~m[531]&m[787])|(m[45]&m[531]&m[787]))):InitCond[87];
    m[216] = run?((((~m[46]&~m[547]&~m[803])|(m[46]&m[547]&~m[803]))&BiasedRNG[56])|(((m[46]&~m[547]&~m[803])|(~m[46]&m[547]&m[803]))&~BiasedRNG[56])|((~m[46]&~m[547]&m[803])|(m[46]&~m[547]&m[803])|(m[46]&m[547]&m[803]))):InitCond[88];
    m[217] = run?((((~m[46]&~m[563]&~m[819])|(m[46]&m[563]&~m[819]))&BiasedRNG[57])|(((m[46]&~m[563]&~m[819])|(~m[46]&m[563]&m[819]))&~BiasedRNG[57])|((~m[46]&~m[563]&m[819])|(m[46]&~m[563]&m[819])|(m[46]&m[563]&m[819]))):InitCond[89];
    m[218] = run?((((~m[46]&~m[579]&~m[835])|(m[46]&m[579]&~m[835]))&BiasedRNG[58])|(((m[46]&~m[579]&~m[835])|(~m[46]&m[579]&m[835]))&~BiasedRNG[58])|((~m[46]&~m[579]&m[835])|(m[46]&~m[579]&m[835])|(m[46]&m[579]&m[835]))):InitCond[90];
    m[219] = run?((((~m[46]&~m[595]&~m[851])|(m[46]&m[595]&~m[851]))&BiasedRNG[59])|(((m[46]&~m[595]&~m[851])|(~m[46]&m[595]&m[851]))&~BiasedRNG[59])|((~m[46]&~m[595]&m[851])|(m[46]&~m[595]&m[851])|(m[46]&m[595]&m[851]))):InitCond[91];
    m[220] = run?((((~m[47]&~m[611]&~m[867])|(m[47]&m[611]&~m[867]))&BiasedRNG[60])|(((m[47]&~m[611]&~m[867])|(~m[47]&m[611]&m[867]))&~BiasedRNG[60])|((~m[47]&~m[611]&m[867])|(m[47]&~m[611]&m[867])|(m[47]&m[611]&m[867]))):InitCond[92];
    m[221] = run?((((~m[47]&~m[627]&~m[883])|(m[47]&m[627]&~m[883]))&BiasedRNG[61])|(((m[47]&~m[627]&~m[883])|(~m[47]&m[627]&m[883]))&~BiasedRNG[61])|((~m[47]&~m[627]&m[883])|(m[47]&~m[627]&m[883])|(m[47]&m[627]&m[883]))):InitCond[93];
    m[222] = run?((((~m[47]&~m[643]&~m[899])|(m[47]&m[643]&~m[899]))&BiasedRNG[62])|(((m[47]&~m[643]&~m[899])|(~m[47]&m[643]&m[899]))&~BiasedRNG[62])|((~m[47]&~m[643]&m[899])|(m[47]&~m[643]&m[899])|(m[47]&m[643]&m[899]))):InitCond[94];
    m[223] = run?((((~m[47]&~m[659]&~m[915])|(m[47]&m[659]&~m[915]))&BiasedRNG[63])|(((m[47]&~m[659]&~m[915])|(~m[47]&m[659]&m[915]))&~BiasedRNG[63])|((~m[47]&~m[659]&m[915])|(m[47]&~m[659]&m[915])|(m[47]&m[659]&m[915]))):InitCond[95];
    m[224] = run?((((~m[48]&~m[420]&~m[676])|(m[48]&m[420]&~m[676]))&BiasedRNG[64])|(((m[48]&~m[420]&~m[676])|(~m[48]&m[420]&m[676]))&~BiasedRNG[64])|((~m[48]&~m[420]&m[676])|(m[48]&~m[420]&m[676])|(m[48]&m[420]&m[676]))):InitCond[96];
    m[225] = run?((((~m[48]&~m[436]&~m[692])|(m[48]&m[436]&~m[692]))&BiasedRNG[65])|(((m[48]&~m[436]&~m[692])|(~m[48]&m[436]&m[692]))&~BiasedRNG[65])|((~m[48]&~m[436]&m[692])|(m[48]&~m[436]&m[692])|(m[48]&m[436]&m[692]))):InitCond[97];
    m[226] = run?((((~m[48]&~m[452]&~m[708])|(m[48]&m[452]&~m[708]))&BiasedRNG[66])|(((m[48]&~m[452]&~m[708])|(~m[48]&m[452]&m[708]))&~BiasedRNG[66])|((~m[48]&~m[452]&m[708])|(m[48]&~m[452]&m[708])|(m[48]&m[452]&m[708]))):InitCond[98];
    m[227] = run?((((~m[48]&~m[468]&~m[724])|(m[48]&m[468]&~m[724]))&BiasedRNG[67])|(((m[48]&~m[468]&~m[724])|(~m[48]&m[468]&m[724]))&~BiasedRNG[67])|((~m[48]&~m[468]&m[724])|(m[48]&~m[468]&m[724])|(m[48]&m[468]&m[724]))):InitCond[99];
    m[228] = run?((((~m[49]&~m[484]&~m[740])|(m[49]&m[484]&~m[740]))&BiasedRNG[68])|(((m[49]&~m[484]&~m[740])|(~m[49]&m[484]&m[740]))&~BiasedRNG[68])|((~m[49]&~m[484]&m[740])|(m[49]&~m[484]&m[740])|(m[49]&m[484]&m[740]))):InitCond[100];
    m[229] = run?((((~m[49]&~m[500]&~m[756])|(m[49]&m[500]&~m[756]))&BiasedRNG[69])|(((m[49]&~m[500]&~m[756])|(~m[49]&m[500]&m[756]))&~BiasedRNG[69])|((~m[49]&~m[500]&m[756])|(m[49]&~m[500]&m[756])|(m[49]&m[500]&m[756]))):InitCond[101];
    m[230] = run?((((~m[49]&~m[516]&~m[772])|(m[49]&m[516]&~m[772]))&BiasedRNG[70])|(((m[49]&~m[516]&~m[772])|(~m[49]&m[516]&m[772]))&~BiasedRNG[70])|((~m[49]&~m[516]&m[772])|(m[49]&~m[516]&m[772])|(m[49]&m[516]&m[772]))):InitCond[102];
    m[231] = run?((((~m[49]&~m[532]&~m[788])|(m[49]&m[532]&~m[788]))&BiasedRNG[71])|(((m[49]&~m[532]&~m[788])|(~m[49]&m[532]&m[788]))&~BiasedRNG[71])|((~m[49]&~m[532]&m[788])|(m[49]&~m[532]&m[788])|(m[49]&m[532]&m[788]))):InitCond[103];
    m[232] = run?((((~m[50]&~m[548]&~m[804])|(m[50]&m[548]&~m[804]))&BiasedRNG[72])|(((m[50]&~m[548]&~m[804])|(~m[50]&m[548]&m[804]))&~BiasedRNG[72])|((~m[50]&~m[548]&m[804])|(m[50]&~m[548]&m[804])|(m[50]&m[548]&m[804]))):InitCond[104];
    m[233] = run?((((~m[50]&~m[564]&~m[820])|(m[50]&m[564]&~m[820]))&BiasedRNG[73])|(((m[50]&~m[564]&~m[820])|(~m[50]&m[564]&m[820]))&~BiasedRNG[73])|((~m[50]&~m[564]&m[820])|(m[50]&~m[564]&m[820])|(m[50]&m[564]&m[820]))):InitCond[105];
    m[234] = run?((((~m[50]&~m[580]&~m[836])|(m[50]&m[580]&~m[836]))&BiasedRNG[74])|(((m[50]&~m[580]&~m[836])|(~m[50]&m[580]&m[836]))&~BiasedRNG[74])|((~m[50]&~m[580]&m[836])|(m[50]&~m[580]&m[836])|(m[50]&m[580]&m[836]))):InitCond[106];
    m[235] = run?((((~m[50]&~m[596]&~m[852])|(m[50]&m[596]&~m[852]))&BiasedRNG[75])|(((m[50]&~m[596]&~m[852])|(~m[50]&m[596]&m[852]))&~BiasedRNG[75])|((~m[50]&~m[596]&m[852])|(m[50]&~m[596]&m[852])|(m[50]&m[596]&m[852]))):InitCond[107];
    m[236] = run?((((~m[51]&~m[612]&~m[868])|(m[51]&m[612]&~m[868]))&BiasedRNG[76])|(((m[51]&~m[612]&~m[868])|(~m[51]&m[612]&m[868]))&~BiasedRNG[76])|((~m[51]&~m[612]&m[868])|(m[51]&~m[612]&m[868])|(m[51]&m[612]&m[868]))):InitCond[108];
    m[237] = run?((((~m[51]&~m[628]&~m[884])|(m[51]&m[628]&~m[884]))&BiasedRNG[77])|(((m[51]&~m[628]&~m[884])|(~m[51]&m[628]&m[884]))&~BiasedRNG[77])|((~m[51]&~m[628]&m[884])|(m[51]&~m[628]&m[884])|(m[51]&m[628]&m[884]))):InitCond[109];
    m[238] = run?((((~m[51]&~m[644]&~m[900])|(m[51]&m[644]&~m[900]))&BiasedRNG[78])|(((m[51]&~m[644]&~m[900])|(~m[51]&m[644]&m[900]))&~BiasedRNG[78])|((~m[51]&~m[644]&m[900])|(m[51]&~m[644]&m[900])|(m[51]&m[644]&m[900]))):InitCond[110];
    m[239] = run?((((~m[51]&~m[660]&~m[916])|(m[51]&m[660]&~m[916]))&BiasedRNG[79])|(((m[51]&~m[660]&~m[916])|(~m[51]&m[660]&m[916]))&~BiasedRNG[79])|((~m[51]&~m[660]&m[916])|(m[51]&~m[660]&m[916])|(m[51]&m[660]&m[916]))):InitCond[111];
    m[240] = run?((((~m[52]&~m[421]&~m[677])|(m[52]&m[421]&~m[677]))&BiasedRNG[80])|(((m[52]&~m[421]&~m[677])|(~m[52]&m[421]&m[677]))&~BiasedRNG[80])|((~m[52]&~m[421]&m[677])|(m[52]&~m[421]&m[677])|(m[52]&m[421]&m[677]))):InitCond[112];
    m[241] = run?((((~m[52]&~m[437]&~m[693])|(m[52]&m[437]&~m[693]))&BiasedRNG[81])|(((m[52]&~m[437]&~m[693])|(~m[52]&m[437]&m[693]))&~BiasedRNG[81])|((~m[52]&~m[437]&m[693])|(m[52]&~m[437]&m[693])|(m[52]&m[437]&m[693]))):InitCond[113];
    m[242] = run?((((~m[52]&~m[453]&~m[709])|(m[52]&m[453]&~m[709]))&BiasedRNG[82])|(((m[52]&~m[453]&~m[709])|(~m[52]&m[453]&m[709]))&~BiasedRNG[82])|((~m[52]&~m[453]&m[709])|(m[52]&~m[453]&m[709])|(m[52]&m[453]&m[709]))):InitCond[114];
    m[243] = run?((((~m[52]&~m[469]&~m[725])|(m[52]&m[469]&~m[725]))&BiasedRNG[83])|(((m[52]&~m[469]&~m[725])|(~m[52]&m[469]&m[725]))&~BiasedRNG[83])|((~m[52]&~m[469]&m[725])|(m[52]&~m[469]&m[725])|(m[52]&m[469]&m[725]))):InitCond[115];
    m[244] = run?((((~m[53]&~m[485]&~m[741])|(m[53]&m[485]&~m[741]))&BiasedRNG[84])|(((m[53]&~m[485]&~m[741])|(~m[53]&m[485]&m[741]))&~BiasedRNG[84])|((~m[53]&~m[485]&m[741])|(m[53]&~m[485]&m[741])|(m[53]&m[485]&m[741]))):InitCond[116];
    m[245] = run?((((~m[53]&~m[501]&~m[757])|(m[53]&m[501]&~m[757]))&BiasedRNG[85])|(((m[53]&~m[501]&~m[757])|(~m[53]&m[501]&m[757]))&~BiasedRNG[85])|((~m[53]&~m[501]&m[757])|(m[53]&~m[501]&m[757])|(m[53]&m[501]&m[757]))):InitCond[117];
    m[246] = run?((((~m[53]&~m[517]&~m[773])|(m[53]&m[517]&~m[773]))&BiasedRNG[86])|(((m[53]&~m[517]&~m[773])|(~m[53]&m[517]&m[773]))&~BiasedRNG[86])|((~m[53]&~m[517]&m[773])|(m[53]&~m[517]&m[773])|(m[53]&m[517]&m[773]))):InitCond[118];
    m[247] = run?((((~m[53]&~m[533]&~m[789])|(m[53]&m[533]&~m[789]))&BiasedRNG[87])|(((m[53]&~m[533]&~m[789])|(~m[53]&m[533]&m[789]))&~BiasedRNG[87])|((~m[53]&~m[533]&m[789])|(m[53]&~m[533]&m[789])|(m[53]&m[533]&m[789]))):InitCond[119];
    m[248] = run?((((~m[54]&~m[549]&~m[805])|(m[54]&m[549]&~m[805]))&BiasedRNG[88])|(((m[54]&~m[549]&~m[805])|(~m[54]&m[549]&m[805]))&~BiasedRNG[88])|((~m[54]&~m[549]&m[805])|(m[54]&~m[549]&m[805])|(m[54]&m[549]&m[805]))):InitCond[120];
    m[249] = run?((((~m[54]&~m[565]&~m[821])|(m[54]&m[565]&~m[821]))&BiasedRNG[89])|(((m[54]&~m[565]&~m[821])|(~m[54]&m[565]&m[821]))&~BiasedRNG[89])|((~m[54]&~m[565]&m[821])|(m[54]&~m[565]&m[821])|(m[54]&m[565]&m[821]))):InitCond[121];
    m[250] = run?((((~m[54]&~m[581]&~m[837])|(m[54]&m[581]&~m[837]))&BiasedRNG[90])|(((m[54]&~m[581]&~m[837])|(~m[54]&m[581]&m[837]))&~BiasedRNG[90])|((~m[54]&~m[581]&m[837])|(m[54]&~m[581]&m[837])|(m[54]&m[581]&m[837]))):InitCond[122];
    m[251] = run?((((~m[54]&~m[597]&~m[853])|(m[54]&m[597]&~m[853]))&BiasedRNG[91])|(((m[54]&~m[597]&~m[853])|(~m[54]&m[597]&m[853]))&~BiasedRNG[91])|((~m[54]&~m[597]&m[853])|(m[54]&~m[597]&m[853])|(m[54]&m[597]&m[853]))):InitCond[123];
    m[252] = run?((((~m[55]&~m[613]&~m[869])|(m[55]&m[613]&~m[869]))&BiasedRNG[92])|(((m[55]&~m[613]&~m[869])|(~m[55]&m[613]&m[869]))&~BiasedRNG[92])|((~m[55]&~m[613]&m[869])|(m[55]&~m[613]&m[869])|(m[55]&m[613]&m[869]))):InitCond[124];
    m[253] = run?((((~m[55]&~m[629]&~m[885])|(m[55]&m[629]&~m[885]))&BiasedRNG[93])|(((m[55]&~m[629]&~m[885])|(~m[55]&m[629]&m[885]))&~BiasedRNG[93])|((~m[55]&~m[629]&m[885])|(m[55]&~m[629]&m[885])|(m[55]&m[629]&m[885]))):InitCond[125];
    m[254] = run?((((~m[55]&~m[645]&~m[901])|(m[55]&m[645]&~m[901]))&BiasedRNG[94])|(((m[55]&~m[645]&~m[901])|(~m[55]&m[645]&m[901]))&~BiasedRNG[94])|((~m[55]&~m[645]&m[901])|(m[55]&~m[645]&m[901])|(m[55]&m[645]&m[901]))):InitCond[126];
    m[255] = run?((((~m[55]&~m[661]&~m[917])|(m[55]&m[661]&~m[917]))&BiasedRNG[95])|(((m[55]&~m[661]&~m[917])|(~m[55]&m[661]&m[917]))&~BiasedRNG[95])|((~m[55]&~m[661]&m[917])|(m[55]&~m[661]&m[917])|(m[55]&m[661]&m[917]))):InitCond[127];
    m[256] = run?((((~m[56]&~m[422]&~m[678])|(m[56]&m[422]&~m[678]))&BiasedRNG[96])|(((m[56]&~m[422]&~m[678])|(~m[56]&m[422]&m[678]))&~BiasedRNG[96])|((~m[56]&~m[422]&m[678])|(m[56]&~m[422]&m[678])|(m[56]&m[422]&m[678]))):InitCond[128];
    m[257] = run?((((~m[56]&~m[438]&~m[694])|(m[56]&m[438]&~m[694]))&BiasedRNG[97])|(((m[56]&~m[438]&~m[694])|(~m[56]&m[438]&m[694]))&~BiasedRNG[97])|((~m[56]&~m[438]&m[694])|(m[56]&~m[438]&m[694])|(m[56]&m[438]&m[694]))):InitCond[129];
    m[258] = run?((((~m[56]&~m[454]&~m[710])|(m[56]&m[454]&~m[710]))&BiasedRNG[98])|(((m[56]&~m[454]&~m[710])|(~m[56]&m[454]&m[710]))&~BiasedRNG[98])|((~m[56]&~m[454]&m[710])|(m[56]&~m[454]&m[710])|(m[56]&m[454]&m[710]))):InitCond[130];
    m[259] = run?((((~m[56]&~m[470]&~m[726])|(m[56]&m[470]&~m[726]))&BiasedRNG[99])|(((m[56]&~m[470]&~m[726])|(~m[56]&m[470]&m[726]))&~BiasedRNG[99])|((~m[56]&~m[470]&m[726])|(m[56]&~m[470]&m[726])|(m[56]&m[470]&m[726]))):InitCond[131];
    m[260] = run?((((~m[57]&~m[486]&~m[742])|(m[57]&m[486]&~m[742]))&BiasedRNG[100])|(((m[57]&~m[486]&~m[742])|(~m[57]&m[486]&m[742]))&~BiasedRNG[100])|((~m[57]&~m[486]&m[742])|(m[57]&~m[486]&m[742])|(m[57]&m[486]&m[742]))):InitCond[132];
    m[261] = run?((((~m[57]&~m[502]&~m[758])|(m[57]&m[502]&~m[758]))&BiasedRNG[101])|(((m[57]&~m[502]&~m[758])|(~m[57]&m[502]&m[758]))&~BiasedRNG[101])|((~m[57]&~m[502]&m[758])|(m[57]&~m[502]&m[758])|(m[57]&m[502]&m[758]))):InitCond[133];
    m[262] = run?((((~m[57]&~m[518]&~m[774])|(m[57]&m[518]&~m[774]))&BiasedRNG[102])|(((m[57]&~m[518]&~m[774])|(~m[57]&m[518]&m[774]))&~BiasedRNG[102])|((~m[57]&~m[518]&m[774])|(m[57]&~m[518]&m[774])|(m[57]&m[518]&m[774]))):InitCond[134];
    m[263] = run?((((~m[57]&~m[534]&~m[790])|(m[57]&m[534]&~m[790]))&BiasedRNG[103])|(((m[57]&~m[534]&~m[790])|(~m[57]&m[534]&m[790]))&~BiasedRNG[103])|((~m[57]&~m[534]&m[790])|(m[57]&~m[534]&m[790])|(m[57]&m[534]&m[790]))):InitCond[135];
    m[264] = run?((((~m[58]&~m[550]&~m[806])|(m[58]&m[550]&~m[806]))&BiasedRNG[104])|(((m[58]&~m[550]&~m[806])|(~m[58]&m[550]&m[806]))&~BiasedRNG[104])|((~m[58]&~m[550]&m[806])|(m[58]&~m[550]&m[806])|(m[58]&m[550]&m[806]))):InitCond[136];
    m[265] = run?((((~m[58]&~m[566]&~m[822])|(m[58]&m[566]&~m[822]))&BiasedRNG[105])|(((m[58]&~m[566]&~m[822])|(~m[58]&m[566]&m[822]))&~BiasedRNG[105])|((~m[58]&~m[566]&m[822])|(m[58]&~m[566]&m[822])|(m[58]&m[566]&m[822]))):InitCond[137];
    m[266] = run?((((~m[58]&~m[582]&~m[838])|(m[58]&m[582]&~m[838]))&BiasedRNG[106])|(((m[58]&~m[582]&~m[838])|(~m[58]&m[582]&m[838]))&~BiasedRNG[106])|((~m[58]&~m[582]&m[838])|(m[58]&~m[582]&m[838])|(m[58]&m[582]&m[838]))):InitCond[138];
    m[267] = run?((((~m[58]&~m[598]&~m[854])|(m[58]&m[598]&~m[854]))&BiasedRNG[107])|(((m[58]&~m[598]&~m[854])|(~m[58]&m[598]&m[854]))&~BiasedRNG[107])|((~m[58]&~m[598]&m[854])|(m[58]&~m[598]&m[854])|(m[58]&m[598]&m[854]))):InitCond[139];
    m[268] = run?((((~m[59]&~m[614]&~m[870])|(m[59]&m[614]&~m[870]))&BiasedRNG[108])|(((m[59]&~m[614]&~m[870])|(~m[59]&m[614]&m[870]))&~BiasedRNG[108])|((~m[59]&~m[614]&m[870])|(m[59]&~m[614]&m[870])|(m[59]&m[614]&m[870]))):InitCond[140];
    m[269] = run?((((~m[59]&~m[630]&~m[886])|(m[59]&m[630]&~m[886]))&BiasedRNG[109])|(((m[59]&~m[630]&~m[886])|(~m[59]&m[630]&m[886]))&~BiasedRNG[109])|((~m[59]&~m[630]&m[886])|(m[59]&~m[630]&m[886])|(m[59]&m[630]&m[886]))):InitCond[141];
    m[270] = run?((((~m[59]&~m[646]&~m[902])|(m[59]&m[646]&~m[902]))&BiasedRNG[110])|(((m[59]&~m[646]&~m[902])|(~m[59]&m[646]&m[902]))&~BiasedRNG[110])|((~m[59]&~m[646]&m[902])|(m[59]&~m[646]&m[902])|(m[59]&m[646]&m[902]))):InitCond[142];
    m[271] = run?((((~m[59]&~m[662]&~m[918])|(m[59]&m[662]&~m[918]))&BiasedRNG[111])|(((m[59]&~m[662]&~m[918])|(~m[59]&m[662]&m[918]))&~BiasedRNG[111])|((~m[59]&~m[662]&m[918])|(m[59]&~m[662]&m[918])|(m[59]&m[662]&m[918]))):InitCond[143];
    m[272] = run?((((~m[60]&~m[423]&~m[679])|(m[60]&m[423]&~m[679]))&BiasedRNG[112])|(((m[60]&~m[423]&~m[679])|(~m[60]&m[423]&m[679]))&~BiasedRNG[112])|((~m[60]&~m[423]&m[679])|(m[60]&~m[423]&m[679])|(m[60]&m[423]&m[679]))):InitCond[144];
    m[273] = run?((((~m[60]&~m[439]&~m[695])|(m[60]&m[439]&~m[695]))&BiasedRNG[113])|(((m[60]&~m[439]&~m[695])|(~m[60]&m[439]&m[695]))&~BiasedRNG[113])|((~m[60]&~m[439]&m[695])|(m[60]&~m[439]&m[695])|(m[60]&m[439]&m[695]))):InitCond[145];
    m[274] = run?((((~m[60]&~m[455]&~m[711])|(m[60]&m[455]&~m[711]))&BiasedRNG[114])|(((m[60]&~m[455]&~m[711])|(~m[60]&m[455]&m[711]))&~BiasedRNG[114])|((~m[60]&~m[455]&m[711])|(m[60]&~m[455]&m[711])|(m[60]&m[455]&m[711]))):InitCond[146];
    m[275] = run?((((~m[60]&~m[471]&~m[727])|(m[60]&m[471]&~m[727]))&BiasedRNG[115])|(((m[60]&~m[471]&~m[727])|(~m[60]&m[471]&m[727]))&~BiasedRNG[115])|((~m[60]&~m[471]&m[727])|(m[60]&~m[471]&m[727])|(m[60]&m[471]&m[727]))):InitCond[147];
    m[276] = run?((((~m[61]&~m[487]&~m[743])|(m[61]&m[487]&~m[743]))&BiasedRNG[116])|(((m[61]&~m[487]&~m[743])|(~m[61]&m[487]&m[743]))&~BiasedRNG[116])|((~m[61]&~m[487]&m[743])|(m[61]&~m[487]&m[743])|(m[61]&m[487]&m[743]))):InitCond[148];
    m[277] = run?((((~m[61]&~m[503]&~m[759])|(m[61]&m[503]&~m[759]))&BiasedRNG[117])|(((m[61]&~m[503]&~m[759])|(~m[61]&m[503]&m[759]))&~BiasedRNG[117])|((~m[61]&~m[503]&m[759])|(m[61]&~m[503]&m[759])|(m[61]&m[503]&m[759]))):InitCond[149];
    m[278] = run?((((~m[61]&~m[519]&~m[775])|(m[61]&m[519]&~m[775]))&BiasedRNG[118])|(((m[61]&~m[519]&~m[775])|(~m[61]&m[519]&m[775]))&~BiasedRNG[118])|((~m[61]&~m[519]&m[775])|(m[61]&~m[519]&m[775])|(m[61]&m[519]&m[775]))):InitCond[150];
    m[279] = run?((((~m[61]&~m[535]&~m[791])|(m[61]&m[535]&~m[791]))&BiasedRNG[119])|(((m[61]&~m[535]&~m[791])|(~m[61]&m[535]&m[791]))&~BiasedRNG[119])|((~m[61]&~m[535]&m[791])|(m[61]&~m[535]&m[791])|(m[61]&m[535]&m[791]))):InitCond[151];
    m[280] = run?((((~m[62]&~m[551]&~m[807])|(m[62]&m[551]&~m[807]))&BiasedRNG[120])|(((m[62]&~m[551]&~m[807])|(~m[62]&m[551]&m[807]))&~BiasedRNG[120])|((~m[62]&~m[551]&m[807])|(m[62]&~m[551]&m[807])|(m[62]&m[551]&m[807]))):InitCond[152];
    m[281] = run?((((~m[62]&~m[567]&~m[823])|(m[62]&m[567]&~m[823]))&BiasedRNG[121])|(((m[62]&~m[567]&~m[823])|(~m[62]&m[567]&m[823]))&~BiasedRNG[121])|((~m[62]&~m[567]&m[823])|(m[62]&~m[567]&m[823])|(m[62]&m[567]&m[823]))):InitCond[153];
    m[282] = run?((((~m[62]&~m[583]&~m[839])|(m[62]&m[583]&~m[839]))&BiasedRNG[122])|(((m[62]&~m[583]&~m[839])|(~m[62]&m[583]&m[839]))&~BiasedRNG[122])|((~m[62]&~m[583]&m[839])|(m[62]&~m[583]&m[839])|(m[62]&m[583]&m[839]))):InitCond[154];
    m[283] = run?((((~m[62]&~m[599]&~m[855])|(m[62]&m[599]&~m[855]))&BiasedRNG[123])|(((m[62]&~m[599]&~m[855])|(~m[62]&m[599]&m[855]))&~BiasedRNG[123])|((~m[62]&~m[599]&m[855])|(m[62]&~m[599]&m[855])|(m[62]&m[599]&m[855]))):InitCond[155];
    m[284] = run?((((~m[63]&~m[615]&~m[871])|(m[63]&m[615]&~m[871]))&BiasedRNG[124])|(((m[63]&~m[615]&~m[871])|(~m[63]&m[615]&m[871]))&~BiasedRNG[124])|((~m[63]&~m[615]&m[871])|(m[63]&~m[615]&m[871])|(m[63]&m[615]&m[871]))):InitCond[156];
    m[285] = run?((((~m[63]&~m[631]&~m[887])|(m[63]&m[631]&~m[887]))&BiasedRNG[125])|(((m[63]&~m[631]&~m[887])|(~m[63]&m[631]&m[887]))&~BiasedRNG[125])|((~m[63]&~m[631]&m[887])|(m[63]&~m[631]&m[887])|(m[63]&m[631]&m[887]))):InitCond[157];
    m[286] = run?((((~m[63]&~m[647]&~m[903])|(m[63]&m[647]&~m[903]))&BiasedRNG[126])|(((m[63]&~m[647]&~m[903])|(~m[63]&m[647]&m[903]))&~BiasedRNG[126])|((~m[63]&~m[647]&m[903])|(m[63]&~m[647]&m[903])|(m[63]&m[647]&m[903]))):InitCond[158];
    m[287] = run?((((~m[63]&~m[663]&~m[919])|(m[63]&m[663]&~m[919]))&BiasedRNG[127])|(((m[63]&~m[663]&~m[919])|(~m[63]&m[663]&m[919]))&~BiasedRNG[127])|((~m[63]&~m[663]&m[919])|(m[63]&~m[663]&m[919])|(m[63]&m[663]&m[919]))):InitCond[159];
    m[288] = run?((((~m[64]&~m[424]&~m[680])|(m[64]&m[424]&~m[680]))&BiasedRNG[128])|(((m[64]&~m[424]&~m[680])|(~m[64]&m[424]&m[680]))&~BiasedRNG[128])|((~m[64]&~m[424]&m[680])|(m[64]&~m[424]&m[680])|(m[64]&m[424]&m[680]))):InitCond[160];
    m[289] = run?((((~m[64]&~m[440]&~m[696])|(m[64]&m[440]&~m[696]))&BiasedRNG[129])|(((m[64]&~m[440]&~m[696])|(~m[64]&m[440]&m[696]))&~BiasedRNG[129])|((~m[64]&~m[440]&m[696])|(m[64]&~m[440]&m[696])|(m[64]&m[440]&m[696]))):InitCond[161];
    m[290] = run?((((~m[64]&~m[456]&~m[712])|(m[64]&m[456]&~m[712]))&BiasedRNG[130])|(((m[64]&~m[456]&~m[712])|(~m[64]&m[456]&m[712]))&~BiasedRNG[130])|((~m[64]&~m[456]&m[712])|(m[64]&~m[456]&m[712])|(m[64]&m[456]&m[712]))):InitCond[162];
    m[291] = run?((((~m[64]&~m[472]&~m[728])|(m[64]&m[472]&~m[728]))&BiasedRNG[131])|(((m[64]&~m[472]&~m[728])|(~m[64]&m[472]&m[728]))&~BiasedRNG[131])|((~m[64]&~m[472]&m[728])|(m[64]&~m[472]&m[728])|(m[64]&m[472]&m[728]))):InitCond[163];
    m[292] = run?((((~m[65]&~m[488]&~m[744])|(m[65]&m[488]&~m[744]))&BiasedRNG[132])|(((m[65]&~m[488]&~m[744])|(~m[65]&m[488]&m[744]))&~BiasedRNG[132])|((~m[65]&~m[488]&m[744])|(m[65]&~m[488]&m[744])|(m[65]&m[488]&m[744]))):InitCond[164];
    m[293] = run?((((~m[65]&~m[504]&~m[760])|(m[65]&m[504]&~m[760]))&BiasedRNG[133])|(((m[65]&~m[504]&~m[760])|(~m[65]&m[504]&m[760]))&~BiasedRNG[133])|((~m[65]&~m[504]&m[760])|(m[65]&~m[504]&m[760])|(m[65]&m[504]&m[760]))):InitCond[165];
    m[294] = run?((((~m[65]&~m[520]&~m[776])|(m[65]&m[520]&~m[776]))&BiasedRNG[134])|(((m[65]&~m[520]&~m[776])|(~m[65]&m[520]&m[776]))&~BiasedRNG[134])|((~m[65]&~m[520]&m[776])|(m[65]&~m[520]&m[776])|(m[65]&m[520]&m[776]))):InitCond[166];
    m[295] = run?((((~m[65]&~m[536]&~m[792])|(m[65]&m[536]&~m[792]))&BiasedRNG[135])|(((m[65]&~m[536]&~m[792])|(~m[65]&m[536]&m[792]))&~BiasedRNG[135])|((~m[65]&~m[536]&m[792])|(m[65]&~m[536]&m[792])|(m[65]&m[536]&m[792]))):InitCond[167];
    m[296] = run?((((~m[66]&~m[552]&~m[808])|(m[66]&m[552]&~m[808]))&BiasedRNG[136])|(((m[66]&~m[552]&~m[808])|(~m[66]&m[552]&m[808]))&~BiasedRNG[136])|((~m[66]&~m[552]&m[808])|(m[66]&~m[552]&m[808])|(m[66]&m[552]&m[808]))):InitCond[168];
    m[297] = run?((((~m[66]&~m[568]&~m[824])|(m[66]&m[568]&~m[824]))&BiasedRNG[137])|(((m[66]&~m[568]&~m[824])|(~m[66]&m[568]&m[824]))&~BiasedRNG[137])|((~m[66]&~m[568]&m[824])|(m[66]&~m[568]&m[824])|(m[66]&m[568]&m[824]))):InitCond[169];
    m[298] = run?((((~m[66]&~m[584]&~m[840])|(m[66]&m[584]&~m[840]))&BiasedRNG[138])|(((m[66]&~m[584]&~m[840])|(~m[66]&m[584]&m[840]))&~BiasedRNG[138])|((~m[66]&~m[584]&m[840])|(m[66]&~m[584]&m[840])|(m[66]&m[584]&m[840]))):InitCond[170];
    m[299] = run?((((~m[66]&~m[600]&~m[856])|(m[66]&m[600]&~m[856]))&BiasedRNG[139])|(((m[66]&~m[600]&~m[856])|(~m[66]&m[600]&m[856]))&~BiasedRNG[139])|((~m[66]&~m[600]&m[856])|(m[66]&~m[600]&m[856])|(m[66]&m[600]&m[856]))):InitCond[171];
    m[300] = run?((((~m[67]&~m[616]&~m[872])|(m[67]&m[616]&~m[872]))&BiasedRNG[140])|(((m[67]&~m[616]&~m[872])|(~m[67]&m[616]&m[872]))&~BiasedRNG[140])|((~m[67]&~m[616]&m[872])|(m[67]&~m[616]&m[872])|(m[67]&m[616]&m[872]))):InitCond[172];
    m[301] = run?((((~m[67]&~m[632]&~m[888])|(m[67]&m[632]&~m[888]))&BiasedRNG[141])|(((m[67]&~m[632]&~m[888])|(~m[67]&m[632]&m[888]))&~BiasedRNG[141])|((~m[67]&~m[632]&m[888])|(m[67]&~m[632]&m[888])|(m[67]&m[632]&m[888]))):InitCond[173];
    m[302] = run?((((~m[67]&~m[648]&~m[904])|(m[67]&m[648]&~m[904]))&BiasedRNG[142])|(((m[67]&~m[648]&~m[904])|(~m[67]&m[648]&m[904]))&~BiasedRNG[142])|((~m[67]&~m[648]&m[904])|(m[67]&~m[648]&m[904])|(m[67]&m[648]&m[904]))):InitCond[174];
    m[303] = run?((((~m[67]&~m[664]&~m[920])|(m[67]&m[664]&~m[920]))&BiasedRNG[143])|(((m[67]&~m[664]&~m[920])|(~m[67]&m[664]&m[920]))&~BiasedRNG[143])|((~m[67]&~m[664]&m[920])|(m[67]&~m[664]&m[920])|(m[67]&m[664]&m[920]))):InitCond[175];
    m[304] = run?((((~m[68]&~m[425]&~m[681])|(m[68]&m[425]&~m[681]))&BiasedRNG[144])|(((m[68]&~m[425]&~m[681])|(~m[68]&m[425]&m[681]))&~BiasedRNG[144])|((~m[68]&~m[425]&m[681])|(m[68]&~m[425]&m[681])|(m[68]&m[425]&m[681]))):InitCond[176];
    m[305] = run?((((~m[68]&~m[441]&~m[697])|(m[68]&m[441]&~m[697]))&BiasedRNG[145])|(((m[68]&~m[441]&~m[697])|(~m[68]&m[441]&m[697]))&~BiasedRNG[145])|((~m[68]&~m[441]&m[697])|(m[68]&~m[441]&m[697])|(m[68]&m[441]&m[697]))):InitCond[177];
    m[306] = run?((((~m[68]&~m[457]&~m[713])|(m[68]&m[457]&~m[713]))&BiasedRNG[146])|(((m[68]&~m[457]&~m[713])|(~m[68]&m[457]&m[713]))&~BiasedRNG[146])|((~m[68]&~m[457]&m[713])|(m[68]&~m[457]&m[713])|(m[68]&m[457]&m[713]))):InitCond[178];
    m[307] = run?((((~m[68]&~m[473]&~m[729])|(m[68]&m[473]&~m[729]))&BiasedRNG[147])|(((m[68]&~m[473]&~m[729])|(~m[68]&m[473]&m[729]))&~BiasedRNG[147])|((~m[68]&~m[473]&m[729])|(m[68]&~m[473]&m[729])|(m[68]&m[473]&m[729]))):InitCond[179];
    m[308] = run?((((~m[69]&~m[489]&~m[745])|(m[69]&m[489]&~m[745]))&BiasedRNG[148])|(((m[69]&~m[489]&~m[745])|(~m[69]&m[489]&m[745]))&~BiasedRNG[148])|((~m[69]&~m[489]&m[745])|(m[69]&~m[489]&m[745])|(m[69]&m[489]&m[745]))):InitCond[180];
    m[309] = run?((((~m[69]&~m[505]&~m[761])|(m[69]&m[505]&~m[761]))&BiasedRNG[149])|(((m[69]&~m[505]&~m[761])|(~m[69]&m[505]&m[761]))&~BiasedRNG[149])|((~m[69]&~m[505]&m[761])|(m[69]&~m[505]&m[761])|(m[69]&m[505]&m[761]))):InitCond[181];
    m[310] = run?((((~m[69]&~m[521]&~m[777])|(m[69]&m[521]&~m[777]))&BiasedRNG[150])|(((m[69]&~m[521]&~m[777])|(~m[69]&m[521]&m[777]))&~BiasedRNG[150])|((~m[69]&~m[521]&m[777])|(m[69]&~m[521]&m[777])|(m[69]&m[521]&m[777]))):InitCond[182];
    m[311] = run?((((~m[69]&~m[537]&~m[793])|(m[69]&m[537]&~m[793]))&BiasedRNG[151])|(((m[69]&~m[537]&~m[793])|(~m[69]&m[537]&m[793]))&~BiasedRNG[151])|((~m[69]&~m[537]&m[793])|(m[69]&~m[537]&m[793])|(m[69]&m[537]&m[793]))):InitCond[183];
    m[312] = run?((((~m[70]&~m[553]&~m[809])|(m[70]&m[553]&~m[809]))&BiasedRNG[152])|(((m[70]&~m[553]&~m[809])|(~m[70]&m[553]&m[809]))&~BiasedRNG[152])|((~m[70]&~m[553]&m[809])|(m[70]&~m[553]&m[809])|(m[70]&m[553]&m[809]))):InitCond[184];
    m[313] = run?((((~m[70]&~m[569]&~m[825])|(m[70]&m[569]&~m[825]))&BiasedRNG[153])|(((m[70]&~m[569]&~m[825])|(~m[70]&m[569]&m[825]))&~BiasedRNG[153])|((~m[70]&~m[569]&m[825])|(m[70]&~m[569]&m[825])|(m[70]&m[569]&m[825]))):InitCond[185];
    m[314] = run?((((~m[70]&~m[585]&~m[841])|(m[70]&m[585]&~m[841]))&BiasedRNG[154])|(((m[70]&~m[585]&~m[841])|(~m[70]&m[585]&m[841]))&~BiasedRNG[154])|((~m[70]&~m[585]&m[841])|(m[70]&~m[585]&m[841])|(m[70]&m[585]&m[841]))):InitCond[186];
    m[315] = run?((((~m[70]&~m[601]&~m[857])|(m[70]&m[601]&~m[857]))&BiasedRNG[155])|(((m[70]&~m[601]&~m[857])|(~m[70]&m[601]&m[857]))&~BiasedRNG[155])|((~m[70]&~m[601]&m[857])|(m[70]&~m[601]&m[857])|(m[70]&m[601]&m[857]))):InitCond[187];
    m[316] = run?((((~m[71]&~m[617]&~m[873])|(m[71]&m[617]&~m[873]))&BiasedRNG[156])|(((m[71]&~m[617]&~m[873])|(~m[71]&m[617]&m[873]))&~BiasedRNG[156])|((~m[71]&~m[617]&m[873])|(m[71]&~m[617]&m[873])|(m[71]&m[617]&m[873]))):InitCond[188];
    m[317] = run?((((~m[71]&~m[633]&~m[889])|(m[71]&m[633]&~m[889]))&BiasedRNG[157])|(((m[71]&~m[633]&~m[889])|(~m[71]&m[633]&m[889]))&~BiasedRNG[157])|((~m[71]&~m[633]&m[889])|(m[71]&~m[633]&m[889])|(m[71]&m[633]&m[889]))):InitCond[189];
    m[318] = run?((((~m[71]&~m[649]&~m[905])|(m[71]&m[649]&~m[905]))&BiasedRNG[158])|(((m[71]&~m[649]&~m[905])|(~m[71]&m[649]&m[905]))&~BiasedRNG[158])|((~m[71]&~m[649]&m[905])|(m[71]&~m[649]&m[905])|(m[71]&m[649]&m[905]))):InitCond[190];
    m[319] = run?((((~m[71]&~m[665]&~m[921])|(m[71]&m[665]&~m[921]))&BiasedRNG[159])|(((m[71]&~m[665]&~m[921])|(~m[71]&m[665]&m[921]))&~BiasedRNG[159])|((~m[71]&~m[665]&m[921])|(m[71]&~m[665]&m[921])|(m[71]&m[665]&m[921]))):InitCond[191];
    m[320] = run?((((~m[72]&~m[426]&~m[682])|(m[72]&m[426]&~m[682]))&BiasedRNG[160])|(((m[72]&~m[426]&~m[682])|(~m[72]&m[426]&m[682]))&~BiasedRNG[160])|((~m[72]&~m[426]&m[682])|(m[72]&~m[426]&m[682])|(m[72]&m[426]&m[682]))):InitCond[192];
    m[321] = run?((((~m[72]&~m[442]&~m[698])|(m[72]&m[442]&~m[698]))&BiasedRNG[161])|(((m[72]&~m[442]&~m[698])|(~m[72]&m[442]&m[698]))&~BiasedRNG[161])|((~m[72]&~m[442]&m[698])|(m[72]&~m[442]&m[698])|(m[72]&m[442]&m[698]))):InitCond[193];
    m[322] = run?((((~m[72]&~m[458]&~m[714])|(m[72]&m[458]&~m[714]))&BiasedRNG[162])|(((m[72]&~m[458]&~m[714])|(~m[72]&m[458]&m[714]))&~BiasedRNG[162])|((~m[72]&~m[458]&m[714])|(m[72]&~m[458]&m[714])|(m[72]&m[458]&m[714]))):InitCond[194];
    m[323] = run?((((~m[72]&~m[474]&~m[730])|(m[72]&m[474]&~m[730]))&BiasedRNG[163])|(((m[72]&~m[474]&~m[730])|(~m[72]&m[474]&m[730]))&~BiasedRNG[163])|((~m[72]&~m[474]&m[730])|(m[72]&~m[474]&m[730])|(m[72]&m[474]&m[730]))):InitCond[195];
    m[324] = run?((((~m[73]&~m[490]&~m[746])|(m[73]&m[490]&~m[746]))&BiasedRNG[164])|(((m[73]&~m[490]&~m[746])|(~m[73]&m[490]&m[746]))&~BiasedRNG[164])|((~m[73]&~m[490]&m[746])|(m[73]&~m[490]&m[746])|(m[73]&m[490]&m[746]))):InitCond[196];
    m[325] = run?((((~m[73]&~m[506]&~m[762])|(m[73]&m[506]&~m[762]))&BiasedRNG[165])|(((m[73]&~m[506]&~m[762])|(~m[73]&m[506]&m[762]))&~BiasedRNG[165])|((~m[73]&~m[506]&m[762])|(m[73]&~m[506]&m[762])|(m[73]&m[506]&m[762]))):InitCond[197];
    m[326] = run?((((~m[73]&~m[522]&~m[778])|(m[73]&m[522]&~m[778]))&BiasedRNG[166])|(((m[73]&~m[522]&~m[778])|(~m[73]&m[522]&m[778]))&~BiasedRNG[166])|((~m[73]&~m[522]&m[778])|(m[73]&~m[522]&m[778])|(m[73]&m[522]&m[778]))):InitCond[198];
    m[327] = run?((((~m[73]&~m[538]&~m[794])|(m[73]&m[538]&~m[794]))&BiasedRNG[167])|(((m[73]&~m[538]&~m[794])|(~m[73]&m[538]&m[794]))&~BiasedRNG[167])|((~m[73]&~m[538]&m[794])|(m[73]&~m[538]&m[794])|(m[73]&m[538]&m[794]))):InitCond[199];
    m[328] = run?((((~m[74]&~m[554]&~m[810])|(m[74]&m[554]&~m[810]))&BiasedRNG[168])|(((m[74]&~m[554]&~m[810])|(~m[74]&m[554]&m[810]))&~BiasedRNG[168])|((~m[74]&~m[554]&m[810])|(m[74]&~m[554]&m[810])|(m[74]&m[554]&m[810]))):InitCond[200];
    m[329] = run?((((~m[74]&~m[570]&~m[826])|(m[74]&m[570]&~m[826]))&BiasedRNG[169])|(((m[74]&~m[570]&~m[826])|(~m[74]&m[570]&m[826]))&~BiasedRNG[169])|((~m[74]&~m[570]&m[826])|(m[74]&~m[570]&m[826])|(m[74]&m[570]&m[826]))):InitCond[201];
    m[330] = run?((((~m[74]&~m[586]&~m[842])|(m[74]&m[586]&~m[842]))&BiasedRNG[170])|(((m[74]&~m[586]&~m[842])|(~m[74]&m[586]&m[842]))&~BiasedRNG[170])|((~m[74]&~m[586]&m[842])|(m[74]&~m[586]&m[842])|(m[74]&m[586]&m[842]))):InitCond[202];
    m[331] = run?((((~m[74]&~m[602]&~m[858])|(m[74]&m[602]&~m[858]))&BiasedRNG[171])|(((m[74]&~m[602]&~m[858])|(~m[74]&m[602]&m[858]))&~BiasedRNG[171])|((~m[74]&~m[602]&m[858])|(m[74]&~m[602]&m[858])|(m[74]&m[602]&m[858]))):InitCond[203];
    m[332] = run?((((~m[75]&~m[618]&~m[874])|(m[75]&m[618]&~m[874]))&BiasedRNG[172])|(((m[75]&~m[618]&~m[874])|(~m[75]&m[618]&m[874]))&~BiasedRNG[172])|((~m[75]&~m[618]&m[874])|(m[75]&~m[618]&m[874])|(m[75]&m[618]&m[874]))):InitCond[204];
    m[333] = run?((((~m[75]&~m[634]&~m[890])|(m[75]&m[634]&~m[890]))&BiasedRNG[173])|(((m[75]&~m[634]&~m[890])|(~m[75]&m[634]&m[890]))&~BiasedRNG[173])|((~m[75]&~m[634]&m[890])|(m[75]&~m[634]&m[890])|(m[75]&m[634]&m[890]))):InitCond[205];
    m[334] = run?((((~m[75]&~m[650]&~m[906])|(m[75]&m[650]&~m[906]))&BiasedRNG[174])|(((m[75]&~m[650]&~m[906])|(~m[75]&m[650]&m[906]))&~BiasedRNG[174])|((~m[75]&~m[650]&m[906])|(m[75]&~m[650]&m[906])|(m[75]&m[650]&m[906]))):InitCond[206];
    m[335] = run?((((~m[75]&~m[666]&~m[922])|(m[75]&m[666]&~m[922]))&BiasedRNG[175])|(((m[75]&~m[666]&~m[922])|(~m[75]&m[666]&m[922]))&~BiasedRNG[175])|((~m[75]&~m[666]&m[922])|(m[75]&~m[666]&m[922])|(m[75]&m[666]&m[922]))):InitCond[207];
    m[336] = run?((((~m[76]&~m[427]&~m[683])|(m[76]&m[427]&~m[683]))&BiasedRNG[176])|(((m[76]&~m[427]&~m[683])|(~m[76]&m[427]&m[683]))&~BiasedRNG[176])|((~m[76]&~m[427]&m[683])|(m[76]&~m[427]&m[683])|(m[76]&m[427]&m[683]))):InitCond[208];
    m[337] = run?((((~m[76]&~m[443]&~m[699])|(m[76]&m[443]&~m[699]))&BiasedRNG[177])|(((m[76]&~m[443]&~m[699])|(~m[76]&m[443]&m[699]))&~BiasedRNG[177])|((~m[76]&~m[443]&m[699])|(m[76]&~m[443]&m[699])|(m[76]&m[443]&m[699]))):InitCond[209];
    m[338] = run?((((~m[76]&~m[459]&~m[715])|(m[76]&m[459]&~m[715]))&BiasedRNG[178])|(((m[76]&~m[459]&~m[715])|(~m[76]&m[459]&m[715]))&~BiasedRNG[178])|((~m[76]&~m[459]&m[715])|(m[76]&~m[459]&m[715])|(m[76]&m[459]&m[715]))):InitCond[210];
    m[339] = run?((((~m[76]&~m[475]&~m[731])|(m[76]&m[475]&~m[731]))&BiasedRNG[179])|(((m[76]&~m[475]&~m[731])|(~m[76]&m[475]&m[731]))&~BiasedRNG[179])|((~m[76]&~m[475]&m[731])|(m[76]&~m[475]&m[731])|(m[76]&m[475]&m[731]))):InitCond[211];
    m[340] = run?((((~m[77]&~m[491]&~m[747])|(m[77]&m[491]&~m[747]))&BiasedRNG[180])|(((m[77]&~m[491]&~m[747])|(~m[77]&m[491]&m[747]))&~BiasedRNG[180])|((~m[77]&~m[491]&m[747])|(m[77]&~m[491]&m[747])|(m[77]&m[491]&m[747]))):InitCond[212];
    m[341] = run?((((~m[77]&~m[507]&~m[763])|(m[77]&m[507]&~m[763]))&BiasedRNG[181])|(((m[77]&~m[507]&~m[763])|(~m[77]&m[507]&m[763]))&~BiasedRNG[181])|((~m[77]&~m[507]&m[763])|(m[77]&~m[507]&m[763])|(m[77]&m[507]&m[763]))):InitCond[213];
    m[342] = run?((((~m[77]&~m[523]&~m[779])|(m[77]&m[523]&~m[779]))&BiasedRNG[182])|(((m[77]&~m[523]&~m[779])|(~m[77]&m[523]&m[779]))&~BiasedRNG[182])|((~m[77]&~m[523]&m[779])|(m[77]&~m[523]&m[779])|(m[77]&m[523]&m[779]))):InitCond[214];
    m[343] = run?((((~m[77]&~m[539]&~m[795])|(m[77]&m[539]&~m[795]))&BiasedRNG[183])|(((m[77]&~m[539]&~m[795])|(~m[77]&m[539]&m[795]))&~BiasedRNG[183])|((~m[77]&~m[539]&m[795])|(m[77]&~m[539]&m[795])|(m[77]&m[539]&m[795]))):InitCond[215];
    m[344] = run?((((~m[78]&~m[555]&~m[811])|(m[78]&m[555]&~m[811]))&BiasedRNG[184])|(((m[78]&~m[555]&~m[811])|(~m[78]&m[555]&m[811]))&~BiasedRNG[184])|((~m[78]&~m[555]&m[811])|(m[78]&~m[555]&m[811])|(m[78]&m[555]&m[811]))):InitCond[216];
    m[345] = run?((((~m[78]&~m[571]&~m[827])|(m[78]&m[571]&~m[827]))&BiasedRNG[185])|(((m[78]&~m[571]&~m[827])|(~m[78]&m[571]&m[827]))&~BiasedRNG[185])|((~m[78]&~m[571]&m[827])|(m[78]&~m[571]&m[827])|(m[78]&m[571]&m[827]))):InitCond[217];
    m[346] = run?((((~m[78]&~m[587]&~m[843])|(m[78]&m[587]&~m[843]))&BiasedRNG[186])|(((m[78]&~m[587]&~m[843])|(~m[78]&m[587]&m[843]))&~BiasedRNG[186])|((~m[78]&~m[587]&m[843])|(m[78]&~m[587]&m[843])|(m[78]&m[587]&m[843]))):InitCond[218];
    m[347] = run?((((~m[78]&~m[603]&~m[859])|(m[78]&m[603]&~m[859]))&BiasedRNG[187])|(((m[78]&~m[603]&~m[859])|(~m[78]&m[603]&m[859]))&~BiasedRNG[187])|((~m[78]&~m[603]&m[859])|(m[78]&~m[603]&m[859])|(m[78]&m[603]&m[859]))):InitCond[219];
    m[348] = run?((((~m[79]&~m[619]&~m[875])|(m[79]&m[619]&~m[875]))&BiasedRNG[188])|(((m[79]&~m[619]&~m[875])|(~m[79]&m[619]&m[875]))&~BiasedRNG[188])|((~m[79]&~m[619]&m[875])|(m[79]&~m[619]&m[875])|(m[79]&m[619]&m[875]))):InitCond[220];
    m[349] = run?((((~m[79]&~m[635]&~m[891])|(m[79]&m[635]&~m[891]))&BiasedRNG[189])|(((m[79]&~m[635]&~m[891])|(~m[79]&m[635]&m[891]))&~BiasedRNG[189])|((~m[79]&~m[635]&m[891])|(m[79]&~m[635]&m[891])|(m[79]&m[635]&m[891]))):InitCond[221];
    m[350] = run?((((~m[79]&~m[651]&~m[907])|(m[79]&m[651]&~m[907]))&BiasedRNG[190])|(((m[79]&~m[651]&~m[907])|(~m[79]&m[651]&m[907]))&~BiasedRNG[190])|((~m[79]&~m[651]&m[907])|(m[79]&~m[651]&m[907])|(m[79]&m[651]&m[907]))):InitCond[222];
    m[351] = run?((((~m[79]&~m[667]&~m[923])|(m[79]&m[667]&~m[923]))&BiasedRNG[191])|(((m[79]&~m[667]&~m[923])|(~m[79]&m[667]&m[923]))&~BiasedRNG[191])|((~m[79]&~m[667]&m[923])|(m[79]&~m[667]&m[923])|(m[79]&m[667]&m[923]))):InitCond[223];
    m[352] = run?((((~m[80]&~m[428]&~m[684])|(m[80]&m[428]&~m[684]))&BiasedRNG[192])|(((m[80]&~m[428]&~m[684])|(~m[80]&m[428]&m[684]))&~BiasedRNG[192])|((~m[80]&~m[428]&m[684])|(m[80]&~m[428]&m[684])|(m[80]&m[428]&m[684]))):InitCond[224];
    m[353] = run?((((~m[80]&~m[444]&~m[700])|(m[80]&m[444]&~m[700]))&BiasedRNG[193])|(((m[80]&~m[444]&~m[700])|(~m[80]&m[444]&m[700]))&~BiasedRNG[193])|((~m[80]&~m[444]&m[700])|(m[80]&~m[444]&m[700])|(m[80]&m[444]&m[700]))):InitCond[225];
    m[354] = run?((((~m[80]&~m[460]&~m[716])|(m[80]&m[460]&~m[716]))&BiasedRNG[194])|(((m[80]&~m[460]&~m[716])|(~m[80]&m[460]&m[716]))&~BiasedRNG[194])|((~m[80]&~m[460]&m[716])|(m[80]&~m[460]&m[716])|(m[80]&m[460]&m[716]))):InitCond[226];
    m[355] = run?((((~m[80]&~m[476]&~m[732])|(m[80]&m[476]&~m[732]))&BiasedRNG[195])|(((m[80]&~m[476]&~m[732])|(~m[80]&m[476]&m[732]))&~BiasedRNG[195])|((~m[80]&~m[476]&m[732])|(m[80]&~m[476]&m[732])|(m[80]&m[476]&m[732]))):InitCond[227];
    m[356] = run?((((~m[81]&~m[492]&~m[748])|(m[81]&m[492]&~m[748]))&BiasedRNG[196])|(((m[81]&~m[492]&~m[748])|(~m[81]&m[492]&m[748]))&~BiasedRNG[196])|((~m[81]&~m[492]&m[748])|(m[81]&~m[492]&m[748])|(m[81]&m[492]&m[748]))):InitCond[228];
    m[357] = run?((((~m[81]&~m[508]&~m[764])|(m[81]&m[508]&~m[764]))&BiasedRNG[197])|(((m[81]&~m[508]&~m[764])|(~m[81]&m[508]&m[764]))&~BiasedRNG[197])|((~m[81]&~m[508]&m[764])|(m[81]&~m[508]&m[764])|(m[81]&m[508]&m[764]))):InitCond[229];
    m[358] = run?((((~m[81]&~m[524]&~m[780])|(m[81]&m[524]&~m[780]))&BiasedRNG[198])|(((m[81]&~m[524]&~m[780])|(~m[81]&m[524]&m[780]))&~BiasedRNG[198])|((~m[81]&~m[524]&m[780])|(m[81]&~m[524]&m[780])|(m[81]&m[524]&m[780]))):InitCond[230];
    m[359] = run?((((~m[81]&~m[540]&~m[796])|(m[81]&m[540]&~m[796]))&BiasedRNG[199])|(((m[81]&~m[540]&~m[796])|(~m[81]&m[540]&m[796]))&~BiasedRNG[199])|((~m[81]&~m[540]&m[796])|(m[81]&~m[540]&m[796])|(m[81]&m[540]&m[796]))):InitCond[231];
    m[360] = run?((((~m[82]&~m[556]&~m[812])|(m[82]&m[556]&~m[812]))&BiasedRNG[200])|(((m[82]&~m[556]&~m[812])|(~m[82]&m[556]&m[812]))&~BiasedRNG[200])|((~m[82]&~m[556]&m[812])|(m[82]&~m[556]&m[812])|(m[82]&m[556]&m[812]))):InitCond[232];
    m[361] = run?((((~m[82]&~m[572]&~m[828])|(m[82]&m[572]&~m[828]))&BiasedRNG[201])|(((m[82]&~m[572]&~m[828])|(~m[82]&m[572]&m[828]))&~BiasedRNG[201])|((~m[82]&~m[572]&m[828])|(m[82]&~m[572]&m[828])|(m[82]&m[572]&m[828]))):InitCond[233];
    m[362] = run?((((~m[82]&~m[588]&~m[844])|(m[82]&m[588]&~m[844]))&BiasedRNG[202])|(((m[82]&~m[588]&~m[844])|(~m[82]&m[588]&m[844]))&~BiasedRNG[202])|((~m[82]&~m[588]&m[844])|(m[82]&~m[588]&m[844])|(m[82]&m[588]&m[844]))):InitCond[234];
    m[363] = run?((((~m[82]&~m[604]&~m[860])|(m[82]&m[604]&~m[860]))&BiasedRNG[203])|(((m[82]&~m[604]&~m[860])|(~m[82]&m[604]&m[860]))&~BiasedRNG[203])|((~m[82]&~m[604]&m[860])|(m[82]&~m[604]&m[860])|(m[82]&m[604]&m[860]))):InitCond[235];
    m[364] = run?((((~m[83]&~m[620]&~m[876])|(m[83]&m[620]&~m[876]))&BiasedRNG[204])|(((m[83]&~m[620]&~m[876])|(~m[83]&m[620]&m[876]))&~BiasedRNG[204])|((~m[83]&~m[620]&m[876])|(m[83]&~m[620]&m[876])|(m[83]&m[620]&m[876]))):InitCond[236];
    m[365] = run?((((~m[83]&~m[636]&~m[892])|(m[83]&m[636]&~m[892]))&BiasedRNG[205])|(((m[83]&~m[636]&~m[892])|(~m[83]&m[636]&m[892]))&~BiasedRNG[205])|((~m[83]&~m[636]&m[892])|(m[83]&~m[636]&m[892])|(m[83]&m[636]&m[892]))):InitCond[237];
    m[366] = run?((((~m[83]&~m[652]&~m[908])|(m[83]&m[652]&~m[908]))&BiasedRNG[206])|(((m[83]&~m[652]&~m[908])|(~m[83]&m[652]&m[908]))&~BiasedRNG[206])|((~m[83]&~m[652]&m[908])|(m[83]&~m[652]&m[908])|(m[83]&m[652]&m[908]))):InitCond[238];
    m[367] = run?((((~m[83]&~m[668]&~m[924])|(m[83]&m[668]&~m[924]))&BiasedRNG[207])|(((m[83]&~m[668]&~m[924])|(~m[83]&m[668]&m[924]))&~BiasedRNG[207])|((~m[83]&~m[668]&m[924])|(m[83]&~m[668]&m[924])|(m[83]&m[668]&m[924]))):InitCond[239];
    m[368] = run?((((~m[84]&~m[429]&~m[685])|(m[84]&m[429]&~m[685]))&BiasedRNG[208])|(((m[84]&~m[429]&~m[685])|(~m[84]&m[429]&m[685]))&~BiasedRNG[208])|((~m[84]&~m[429]&m[685])|(m[84]&~m[429]&m[685])|(m[84]&m[429]&m[685]))):InitCond[240];
    m[369] = run?((((~m[84]&~m[445]&~m[701])|(m[84]&m[445]&~m[701]))&BiasedRNG[209])|(((m[84]&~m[445]&~m[701])|(~m[84]&m[445]&m[701]))&~BiasedRNG[209])|((~m[84]&~m[445]&m[701])|(m[84]&~m[445]&m[701])|(m[84]&m[445]&m[701]))):InitCond[241];
    m[370] = run?((((~m[84]&~m[461]&~m[717])|(m[84]&m[461]&~m[717]))&BiasedRNG[210])|(((m[84]&~m[461]&~m[717])|(~m[84]&m[461]&m[717]))&~BiasedRNG[210])|((~m[84]&~m[461]&m[717])|(m[84]&~m[461]&m[717])|(m[84]&m[461]&m[717]))):InitCond[242];
    m[371] = run?((((~m[84]&~m[477]&~m[733])|(m[84]&m[477]&~m[733]))&BiasedRNG[211])|(((m[84]&~m[477]&~m[733])|(~m[84]&m[477]&m[733]))&~BiasedRNG[211])|((~m[84]&~m[477]&m[733])|(m[84]&~m[477]&m[733])|(m[84]&m[477]&m[733]))):InitCond[243];
    m[372] = run?((((~m[85]&~m[493]&~m[749])|(m[85]&m[493]&~m[749]))&BiasedRNG[212])|(((m[85]&~m[493]&~m[749])|(~m[85]&m[493]&m[749]))&~BiasedRNG[212])|((~m[85]&~m[493]&m[749])|(m[85]&~m[493]&m[749])|(m[85]&m[493]&m[749]))):InitCond[244];
    m[373] = run?((((~m[85]&~m[509]&~m[765])|(m[85]&m[509]&~m[765]))&BiasedRNG[213])|(((m[85]&~m[509]&~m[765])|(~m[85]&m[509]&m[765]))&~BiasedRNG[213])|((~m[85]&~m[509]&m[765])|(m[85]&~m[509]&m[765])|(m[85]&m[509]&m[765]))):InitCond[245];
    m[374] = run?((((~m[85]&~m[525]&~m[781])|(m[85]&m[525]&~m[781]))&BiasedRNG[214])|(((m[85]&~m[525]&~m[781])|(~m[85]&m[525]&m[781]))&~BiasedRNG[214])|((~m[85]&~m[525]&m[781])|(m[85]&~m[525]&m[781])|(m[85]&m[525]&m[781]))):InitCond[246];
    m[375] = run?((((~m[85]&~m[541]&~m[797])|(m[85]&m[541]&~m[797]))&BiasedRNG[215])|(((m[85]&~m[541]&~m[797])|(~m[85]&m[541]&m[797]))&~BiasedRNG[215])|((~m[85]&~m[541]&m[797])|(m[85]&~m[541]&m[797])|(m[85]&m[541]&m[797]))):InitCond[247];
    m[376] = run?((((~m[86]&~m[557]&~m[813])|(m[86]&m[557]&~m[813]))&BiasedRNG[216])|(((m[86]&~m[557]&~m[813])|(~m[86]&m[557]&m[813]))&~BiasedRNG[216])|((~m[86]&~m[557]&m[813])|(m[86]&~m[557]&m[813])|(m[86]&m[557]&m[813]))):InitCond[248];
    m[377] = run?((((~m[86]&~m[573]&~m[829])|(m[86]&m[573]&~m[829]))&BiasedRNG[217])|(((m[86]&~m[573]&~m[829])|(~m[86]&m[573]&m[829]))&~BiasedRNG[217])|((~m[86]&~m[573]&m[829])|(m[86]&~m[573]&m[829])|(m[86]&m[573]&m[829]))):InitCond[249];
    m[378] = run?((((~m[86]&~m[589]&~m[845])|(m[86]&m[589]&~m[845]))&BiasedRNG[218])|(((m[86]&~m[589]&~m[845])|(~m[86]&m[589]&m[845]))&~BiasedRNG[218])|((~m[86]&~m[589]&m[845])|(m[86]&~m[589]&m[845])|(m[86]&m[589]&m[845]))):InitCond[250];
    m[379] = run?((((~m[86]&~m[605]&~m[861])|(m[86]&m[605]&~m[861]))&BiasedRNG[219])|(((m[86]&~m[605]&~m[861])|(~m[86]&m[605]&m[861]))&~BiasedRNG[219])|((~m[86]&~m[605]&m[861])|(m[86]&~m[605]&m[861])|(m[86]&m[605]&m[861]))):InitCond[251];
    m[380] = run?((((~m[87]&~m[621]&~m[877])|(m[87]&m[621]&~m[877]))&BiasedRNG[220])|(((m[87]&~m[621]&~m[877])|(~m[87]&m[621]&m[877]))&~BiasedRNG[220])|((~m[87]&~m[621]&m[877])|(m[87]&~m[621]&m[877])|(m[87]&m[621]&m[877]))):InitCond[252];
    m[381] = run?((((~m[87]&~m[637]&~m[893])|(m[87]&m[637]&~m[893]))&BiasedRNG[221])|(((m[87]&~m[637]&~m[893])|(~m[87]&m[637]&m[893]))&~BiasedRNG[221])|((~m[87]&~m[637]&m[893])|(m[87]&~m[637]&m[893])|(m[87]&m[637]&m[893]))):InitCond[253];
    m[382] = run?((((~m[87]&~m[653]&~m[909])|(m[87]&m[653]&~m[909]))&BiasedRNG[222])|(((m[87]&~m[653]&~m[909])|(~m[87]&m[653]&m[909]))&~BiasedRNG[222])|((~m[87]&~m[653]&m[909])|(m[87]&~m[653]&m[909])|(m[87]&m[653]&m[909]))):InitCond[254];
    m[383] = run?((((~m[87]&~m[669]&~m[925])|(m[87]&m[669]&~m[925]))&BiasedRNG[223])|(((m[87]&~m[669]&~m[925])|(~m[87]&m[669]&m[925]))&~BiasedRNG[223])|((~m[87]&~m[669]&m[925])|(m[87]&~m[669]&m[925])|(m[87]&m[669]&m[925]))):InitCond[255];
    m[384] = run?((((~m[88]&~m[430]&~m[686])|(m[88]&m[430]&~m[686]))&BiasedRNG[224])|(((m[88]&~m[430]&~m[686])|(~m[88]&m[430]&m[686]))&~BiasedRNG[224])|((~m[88]&~m[430]&m[686])|(m[88]&~m[430]&m[686])|(m[88]&m[430]&m[686]))):InitCond[256];
    m[385] = run?((((~m[88]&~m[446]&~m[702])|(m[88]&m[446]&~m[702]))&BiasedRNG[225])|(((m[88]&~m[446]&~m[702])|(~m[88]&m[446]&m[702]))&~BiasedRNG[225])|((~m[88]&~m[446]&m[702])|(m[88]&~m[446]&m[702])|(m[88]&m[446]&m[702]))):InitCond[257];
    m[386] = run?((((~m[88]&~m[462]&~m[718])|(m[88]&m[462]&~m[718]))&BiasedRNG[226])|(((m[88]&~m[462]&~m[718])|(~m[88]&m[462]&m[718]))&~BiasedRNG[226])|((~m[88]&~m[462]&m[718])|(m[88]&~m[462]&m[718])|(m[88]&m[462]&m[718]))):InitCond[258];
    m[387] = run?((((~m[88]&~m[478]&~m[734])|(m[88]&m[478]&~m[734]))&BiasedRNG[227])|(((m[88]&~m[478]&~m[734])|(~m[88]&m[478]&m[734]))&~BiasedRNG[227])|((~m[88]&~m[478]&m[734])|(m[88]&~m[478]&m[734])|(m[88]&m[478]&m[734]))):InitCond[259];
    m[388] = run?((((~m[89]&~m[494]&~m[750])|(m[89]&m[494]&~m[750]))&BiasedRNG[228])|(((m[89]&~m[494]&~m[750])|(~m[89]&m[494]&m[750]))&~BiasedRNG[228])|((~m[89]&~m[494]&m[750])|(m[89]&~m[494]&m[750])|(m[89]&m[494]&m[750]))):InitCond[260];
    m[389] = run?((((~m[89]&~m[510]&~m[766])|(m[89]&m[510]&~m[766]))&BiasedRNG[229])|(((m[89]&~m[510]&~m[766])|(~m[89]&m[510]&m[766]))&~BiasedRNG[229])|((~m[89]&~m[510]&m[766])|(m[89]&~m[510]&m[766])|(m[89]&m[510]&m[766]))):InitCond[261];
    m[390] = run?((((~m[89]&~m[526]&~m[782])|(m[89]&m[526]&~m[782]))&BiasedRNG[230])|(((m[89]&~m[526]&~m[782])|(~m[89]&m[526]&m[782]))&~BiasedRNG[230])|((~m[89]&~m[526]&m[782])|(m[89]&~m[526]&m[782])|(m[89]&m[526]&m[782]))):InitCond[262];
    m[391] = run?((((~m[89]&~m[542]&~m[798])|(m[89]&m[542]&~m[798]))&BiasedRNG[231])|(((m[89]&~m[542]&~m[798])|(~m[89]&m[542]&m[798]))&~BiasedRNG[231])|((~m[89]&~m[542]&m[798])|(m[89]&~m[542]&m[798])|(m[89]&m[542]&m[798]))):InitCond[263];
    m[392] = run?((((~m[90]&~m[558]&~m[814])|(m[90]&m[558]&~m[814]))&BiasedRNG[232])|(((m[90]&~m[558]&~m[814])|(~m[90]&m[558]&m[814]))&~BiasedRNG[232])|((~m[90]&~m[558]&m[814])|(m[90]&~m[558]&m[814])|(m[90]&m[558]&m[814]))):InitCond[264];
    m[393] = run?((((~m[90]&~m[574]&~m[830])|(m[90]&m[574]&~m[830]))&BiasedRNG[233])|(((m[90]&~m[574]&~m[830])|(~m[90]&m[574]&m[830]))&~BiasedRNG[233])|((~m[90]&~m[574]&m[830])|(m[90]&~m[574]&m[830])|(m[90]&m[574]&m[830]))):InitCond[265];
    m[394] = run?((((~m[90]&~m[590]&~m[846])|(m[90]&m[590]&~m[846]))&BiasedRNG[234])|(((m[90]&~m[590]&~m[846])|(~m[90]&m[590]&m[846]))&~BiasedRNG[234])|((~m[90]&~m[590]&m[846])|(m[90]&~m[590]&m[846])|(m[90]&m[590]&m[846]))):InitCond[266];
    m[395] = run?((((~m[90]&~m[606]&~m[862])|(m[90]&m[606]&~m[862]))&BiasedRNG[235])|(((m[90]&~m[606]&~m[862])|(~m[90]&m[606]&m[862]))&~BiasedRNG[235])|((~m[90]&~m[606]&m[862])|(m[90]&~m[606]&m[862])|(m[90]&m[606]&m[862]))):InitCond[267];
    m[396] = run?((((~m[91]&~m[622]&~m[878])|(m[91]&m[622]&~m[878]))&BiasedRNG[236])|(((m[91]&~m[622]&~m[878])|(~m[91]&m[622]&m[878]))&~BiasedRNG[236])|((~m[91]&~m[622]&m[878])|(m[91]&~m[622]&m[878])|(m[91]&m[622]&m[878]))):InitCond[268];
    m[397] = run?((((~m[91]&~m[638]&~m[894])|(m[91]&m[638]&~m[894]))&BiasedRNG[237])|(((m[91]&~m[638]&~m[894])|(~m[91]&m[638]&m[894]))&~BiasedRNG[237])|((~m[91]&~m[638]&m[894])|(m[91]&~m[638]&m[894])|(m[91]&m[638]&m[894]))):InitCond[269];
    m[398] = run?((((~m[91]&~m[654]&~m[910])|(m[91]&m[654]&~m[910]))&BiasedRNG[238])|(((m[91]&~m[654]&~m[910])|(~m[91]&m[654]&m[910]))&~BiasedRNG[238])|((~m[91]&~m[654]&m[910])|(m[91]&~m[654]&m[910])|(m[91]&m[654]&m[910]))):InitCond[270];
    m[399] = run?((((~m[91]&~m[670]&~m[926])|(m[91]&m[670]&~m[926]))&BiasedRNG[239])|(((m[91]&~m[670]&~m[926])|(~m[91]&m[670]&m[926]))&~BiasedRNG[239])|((~m[91]&~m[670]&m[926])|(m[91]&~m[670]&m[926])|(m[91]&m[670]&m[926]))):InitCond[271];
    m[400] = run?((((~m[92]&~m[431]&~m[687])|(m[92]&m[431]&~m[687]))&BiasedRNG[240])|(((m[92]&~m[431]&~m[687])|(~m[92]&m[431]&m[687]))&~BiasedRNG[240])|((~m[92]&~m[431]&m[687])|(m[92]&~m[431]&m[687])|(m[92]&m[431]&m[687]))):InitCond[272];
    m[401] = run?((((~m[92]&~m[447]&~m[703])|(m[92]&m[447]&~m[703]))&BiasedRNG[241])|(((m[92]&~m[447]&~m[703])|(~m[92]&m[447]&m[703]))&~BiasedRNG[241])|((~m[92]&~m[447]&m[703])|(m[92]&~m[447]&m[703])|(m[92]&m[447]&m[703]))):InitCond[273];
    m[402] = run?((((~m[92]&~m[463]&~m[719])|(m[92]&m[463]&~m[719]))&BiasedRNG[242])|(((m[92]&~m[463]&~m[719])|(~m[92]&m[463]&m[719]))&~BiasedRNG[242])|((~m[92]&~m[463]&m[719])|(m[92]&~m[463]&m[719])|(m[92]&m[463]&m[719]))):InitCond[274];
    m[403] = run?((((~m[92]&~m[479]&~m[735])|(m[92]&m[479]&~m[735]))&BiasedRNG[243])|(((m[92]&~m[479]&~m[735])|(~m[92]&m[479]&m[735]))&~BiasedRNG[243])|((~m[92]&~m[479]&m[735])|(m[92]&~m[479]&m[735])|(m[92]&m[479]&m[735]))):InitCond[275];
    m[404] = run?((((~m[93]&~m[495]&~m[751])|(m[93]&m[495]&~m[751]))&BiasedRNG[244])|(((m[93]&~m[495]&~m[751])|(~m[93]&m[495]&m[751]))&~BiasedRNG[244])|((~m[93]&~m[495]&m[751])|(m[93]&~m[495]&m[751])|(m[93]&m[495]&m[751]))):InitCond[276];
    m[405] = run?((((~m[93]&~m[511]&~m[767])|(m[93]&m[511]&~m[767]))&BiasedRNG[245])|(((m[93]&~m[511]&~m[767])|(~m[93]&m[511]&m[767]))&~BiasedRNG[245])|((~m[93]&~m[511]&m[767])|(m[93]&~m[511]&m[767])|(m[93]&m[511]&m[767]))):InitCond[277];
    m[406] = run?((((~m[93]&~m[527]&~m[783])|(m[93]&m[527]&~m[783]))&BiasedRNG[246])|(((m[93]&~m[527]&~m[783])|(~m[93]&m[527]&m[783]))&~BiasedRNG[246])|((~m[93]&~m[527]&m[783])|(m[93]&~m[527]&m[783])|(m[93]&m[527]&m[783]))):InitCond[278];
    m[407] = run?((((~m[93]&~m[543]&~m[799])|(m[93]&m[543]&~m[799]))&BiasedRNG[247])|(((m[93]&~m[543]&~m[799])|(~m[93]&m[543]&m[799]))&~BiasedRNG[247])|((~m[93]&~m[543]&m[799])|(m[93]&~m[543]&m[799])|(m[93]&m[543]&m[799]))):InitCond[279];
    m[408] = run?((((~m[94]&~m[559]&~m[815])|(m[94]&m[559]&~m[815]))&BiasedRNG[248])|(((m[94]&~m[559]&~m[815])|(~m[94]&m[559]&m[815]))&~BiasedRNG[248])|((~m[94]&~m[559]&m[815])|(m[94]&~m[559]&m[815])|(m[94]&m[559]&m[815]))):InitCond[280];
    m[409] = run?((((~m[94]&~m[575]&~m[831])|(m[94]&m[575]&~m[831]))&BiasedRNG[249])|(((m[94]&~m[575]&~m[831])|(~m[94]&m[575]&m[831]))&~BiasedRNG[249])|((~m[94]&~m[575]&m[831])|(m[94]&~m[575]&m[831])|(m[94]&m[575]&m[831]))):InitCond[281];
    m[410] = run?((((~m[94]&~m[591]&~m[847])|(m[94]&m[591]&~m[847]))&BiasedRNG[250])|(((m[94]&~m[591]&~m[847])|(~m[94]&m[591]&m[847]))&~BiasedRNG[250])|((~m[94]&~m[591]&m[847])|(m[94]&~m[591]&m[847])|(m[94]&m[591]&m[847]))):InitCond[282];
    m[411] = run?((((~m[94]&~m[607]&~m[863])|(m[94]&m[607]&~m[863]))&BiasedRNG[251])|(((m[94]&~m[607]&~m[863])|(~m[94]&m[607]&m[863]))&~BiasedRNG[251])|((~m[94]&~m[607]&m[863])|(m[94]&~m[607]&m[863])|(m[94]&m[607]&m[863]))):InitCond[283];
    m[412] = run?((((~m[95]&~m[623]&~m[879])|(m[95]&m[623]&~m[879]))&BiasedRNG[252])|(((m[95]&~m[623]&~m[879])|(~m[95]&m[623]&m[879]))&~BiasedRNG[252])|((~m[95]&~m[623]&m[879])|(m[95]&~m[623]&m[879])|(m[95]&m[623]&m[879]))):InitCond[284];
    m[413] = run?((((~m[95]&~m[639]&~m[895])|(m[95]&m[639]&~m[895]))&BiasedRNG[253])|(((m[95]&~m[639]&~m[895])|(~m[95]&m[639]&m[895]))&~BiasedRNG[253])|((~m[95]&~m[639]&m[895])|(m[95]&~m[639]&m[895])|(m[95]&m[639]&m[895]))):InitCond[285];
    m[414] = run?((((~m[95]&~m[655]&~m[911])|(m[95]&m[655]&~m[911]))&BiasedRNG[254])|(((m[95]&~m[655]&~m[911])|(~m[95]&m[655]&m[911]))&~BiasedRNG[254])|((~m[95]&~m[655]&m[911])|(m[95]&~m[655]&m[911])|(m[95]&m[655]&m[911]))):InitCond[286];
    m[415] = run?((((~m[95]&~m[671]&~m[927])|(m[95]&m[671]&~m[927]))&BiasedRNG[255])|(((m[95]&~m[671]&~m[927])|(~m[95]&m[671]&m[927]))&~BiasedRNG[255])|((~m[95]&~m[671]&m[927])|(m[95]&~m[671]&m[927])|(m[95]&m[671]&m[927]))):InitCond[287];
    m[928] = run?((((m[673]&~m[929]&~m[930]&~m[931]&~m[932])|(~m[673]&~m[929]&~m[930]&m[931]&~m[932])|(m[673]&m[929]&~m[930]&m[931]&~m[932])|(m[673]&~m[929]&m[930]&m[931]&~m[932])|(~m[673]&m[929]&~m[930]&~m[931]&m[932])|(~m[673]&~m[929]&m[930]&~m[931]&m[932])|(m[673]&m[929]&m[930]&~m[931]&m[932])|(~m[673]&m[929]&m[930]&m[931]&m[932]))&UnbiasedRNG[32])|((m[673]&~m[929]&~m[930]&m[931]&~m[932])|(~m[673]&~m[929]&~m[930]&~m[931]&m[932])|(m[673]&~m[929]&~m[930]&~m[931]&m[932])|(m[673]&m[929]&~m[930]&~m[931]&m[932])|(m[673]&~m[929]&m[930]&~m[931]&m[932])|(~m[673]&~m[929]&~m[930]&m[931]&m[932])|(m[673]&~m[929]&~m[930]&m[931]&m[932])|(~m[673]&m[929]&~m[930]&m[931]&m[932])|(m[673]&m[929]&~m[930]&m[931]&m[932])|(~m[673]&~m[929]&m[930]&m[931]&m[932])|(m[673]&~m[929]&m[930]&m[931]&m[932])|(m[673]&m[929]&m[930]&m[931]&m[932]))):InitCond[288];
    m[933] = run?((((m[674]&~m[934]&~m[935]&~m[936]&~m[937])|(~m[674]&~m[934]&~m[935]&m[936]&~m[937])|(m[674]&m[934]&~m[935]&m[936]&~m[937])|(m[674]&~m[934]&m[935]&m[936]&~m[937])|(~m[674]&m[934]&~m[935]&~m[936]&m[937])|(~m[674]&~m[934]&m[935]&~m[936]&m[937])|(m[674]&m[934]&m[935]&~m[936]&m[937])|(~m[674]&m[934]&m[935]&m[936]&m[937]))&UnbiasedRNG[33])|((m[674]&~m[934]&~m[935]&m[936]&~m[937])|(~m[674]&~m[934]&~m[935]&~m[936]&m[937])|(m[674]&~m[934]&~m[935]&~m[936]&m[937])|(m[674]&m[934]&~m[935]&~m[936]&m[937])|(m[674]&~m[934]&m[935]&~m[936]&m[937])|(~m[674]&~m[934]&~m[935]&m[936]&m[937])|(m[674]&~m[934]&~m[935]&m[936]&m[937])|(~m[674]&m[934]&~m[935]&m[936]&m[937])|(m[674]&m[934]&~m[935]&m[936]&m[937])|(~m[674]&~m[934]&m[935]&m[936]&m[937])|(m[674]&~m[934]&m[935]&m[936]&m[937])|(m[674]&m[934]&m[935]&m[936]&m[937]))):InitCond[289];
    m[938] = run?((((m[936]&~m[939]&~m[940]&~m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&m[941]&~m[942])|(m[936]&m[939]&~m[940]&m[941]&~m[942])|(m[936]&~m[939]&m[940]&m[941]&~m[942])|(~m[936]&m[939]&~m[940]&~m[941]&m[942])|(~m[936]&~m[939]&m[940]&~m[941]&m[942])|(m[936]&m[939]&m[940]&~m[941]&m[942])|(~m[936]&m[939]&m[940]&m[941]&m[942]))&UnbiasedRNG[34])|((m[936]&~m[939]&~m[940]&m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&m[940]&~m[941]&m[942])|(~m[936]&~m[939]&~m[940]&m[941]&m[942])|(m[936]&~m[939]&~m[940]&m[941]&m[942])|(~m[936]&m[939]&~m[940]&m[941]&m[942])|(m[936]&m[939]&~m[940]&m[941]&m[942])|(~m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&m[939]&m[940]&m[941]&m[942]))):InitCond[290];
    m[943] = run?((((m[675]&~m[944]&~m[945]&~m[946]&~m[947])|(~m[675]&~m[944]&~m[945]&m[946]&~m[947])|(m[675]&m[944]&~m[945]&m[946]&~m[947])|(m[675]&~m[944]&m[945]&m[946]&~m[947])|(~m[675]&m[944]&~m[945]&~m[946]&m[947])|(~m[675]&~m[944]&m[945]&~m[946]&m[947])|(m[675]&m[944]&m[945]&~m[946]&m[947])|(~m[675]&m[944]&m[945]&m[946]&m[947]))&UnbiasedRNG[35])|((m[675]&~m[944]&~m[945]&m[946]&~m[947])|(~m[675]&~m[944]&~m[945]&~m[946]&m[947])|(m[675]&~m[944]&~m[945]&~m[946]&m[947])|(m[675]&m[944]&~m[945]&~m[946]&m[947])|(m[675]&~m[944]&m[945]&~m[946]&m[947])|(~m[675]&~m[944]&~m[945]&m[946]&m[947])|(m[675]&~m[944]&~m[945]&m[946]&m[947])|(~m[675]&m[944]&~m[945]&m[946]&m[947])|(m[675]&m[944]&~m[945]&m[946]&m[947])|(~m[675]&~m[944]&m[945]&m[946]&m[947])|(m[675]&~m[944]&m[945]&m[946]&m[947])|(m[675]&m[944]&m[945]&m[946]&m[947]))):InitCond[291];
    m[948] = run?((((m[946]&~m[949]&~m[950]&~m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&m[951]&~m[952])|(m[946]&m[949]&~m[950]&m[951]&~m[952])|(m[946]&~m[949]&m[950]&m[951]&~m[952])|(~m[946]&m[949]&~m[950]&~m[951]&m[952])|(~m[946]&~m[949]&m[950]&~m[951]&m[952])|(m[946]&m[949]&m[950]&~m[951]&m[952])|(~m[946]&m[949]&m[950]&m[951]&m[952]))&UnbiasedRNG[36])|((m[946]&~m[949]&~m[950]&m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&m[950]&~m[951]&m[952])|(~m[946]&~m[949]&~m[950]&m[951]&m[952])|(m[946]&~m[949]&~m[950]&m[951]&m[952])|(~m[946]&m[949]&~m[950]&m[951]&m[952])|(m[946]&m[949]&~m[950]&m[951]&m[952])|(~m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&m[949]&m[950]&m[951]&m[952]))):InitCond[292];
    m[953] = run?((((m[951]&~m[954]&~m[955]&~m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&m[956]&~m[957])|(m[951]&m[954]&~m[955]&m[956]&~m[957])|(m[951]&~m[954]&m[955]&m[956]&~m[957])|(~m[951]&m[954]&~m[955]&~m[956]&m[957])|(~m[951]&~m[954]&m[955]&~m[956]&m[957])|(m[951]&m[954]&m[955]&~m[956]&m[957])|(~m[951]&m[954]&m[955]&m[956]&m[957]))&UnbiasedRNG[37])|((m[951]&~m[954]&~m[955]&m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&m[955]&~m[956]&m[957])|(~m[951]&~m[954]&~m[955]&m[956]&m[957])|(m[951]&~m[954]&~m[955]&m[956]&m[957])|(~m[951]&m[954]&~m[955]&m[956]&m[957])|(m[951]&m[954]&~m[955]&m[956]&m[957])|(~m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&m[954]&m[955]&m[956]&m[957]))):InitCond[293];
    m[958] = run?((((m[676]&~m[959]&~m[960]&~m[961]&~m[962])|(~m[676]&~m[959]&~m[960]&m[961]&~m[962])|(m[676]&m[959]&~m[960]&m[961]&~m[962])|(m[676]&~m[959]&m[960]&m[961]&~m[962])|(~m[676]&m[959]&~m[960]&~m[961]&m[962])|(~m[676]&~m[959]&m[960]&~m[961]&m[962])|(m[676]&m[959]&m[960]&~m[961]&m[962])|(~m[676]&m[959]&m[960]&m[961]&m[962]))&UnbiasedRNG[38])|((m[676]&~m[959]&~m[960]&m[961]&~m[962])|(~m[676]&~m[959]&~m[960]&~m[961]&m[962])|(m[676]&~m[959]&~m[960]&~m[961]&m[962])|(m[676]&m[959]&~m[960]&~m[961]&m[962])|(m[676]&~m[959]&m[960]&~m[961]&m[962])|(~m[676]&~m[959]&~m[960]&m[961]&m[962])|(m[676]&~m[959]&~m[960]&m[961]&m[962])|(~m[676]&m[959]&~m[960]&m[961]&m[962])|(m[676]&m[959]&~m[960]&m[961]&m[962])|(~m[676]&~m[959]&m[960]&m[961]&m[962])|(m[676]&~m[959]&m[960]&m[961]&m[962])|(m[676]&m[959]&m[960]&m[961]&m[962]))):InitCond[294];
    m[963] = run?((((m[961]&~m[964]&~m[965]&~m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&m[966]&~m[967])|(m[961]&m[964]&~m[965]&m[966]&~m[967])|(m[961]&~m[964]&m[965]&m[966]&~m[967])|(~m[961]&m[964]&~m[965]&~m[966]&m[967])|(~m[961]&~m[964]&m[965]&~m[966]&m[967])|(m[961]&m[964]&m[965]&~m[966]&m[967])|(~m[961]&m[964]&m[965]&m[966]&m[967]))&UnbiasedRNG[39])|((m[961]&~m[964]&~m[965]&m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&m[965]&~m[966]&m[967])|(~m[961]&~m[964]&~m[965]&m[966]&m[967])|(m[961]&~m[964]&~m[965]&m[966]&m[967])|(~m[961]&m[964]&~m[965]&m[966]&m[967])|(m[961]&m[964]&~m[965]&m[966]&m[967])|(~m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&m[964]&m[965]&m[966]&m[967]))):InitCond[295];
    m[968] = run?((((m[966]&~m[969]&~m[970]&~m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&m[971]&~m[972])|(m[966]&m[969]&~m[970]&m[971]&~m[972])|(m[966]&~m[969]&m[970]&m[971]&~m[972])|(~m[966]&m[969]&~m[970]&~m[971]&m[972])|(~m[966]&~m[969]&m[970]&~m[971]&m[972])|(m[966]&m[969]&m[970]&~m[971]&m[972])|(~m[966]&m[969]&m[970]&m[971]&m[972]))&UnbiasedRNG[40])|((m[966]&~m[969]&~m[970]&m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&m[970]&~m[971]&m[972])|(~m[966]&~m[969]&~m[970]&m[971]&m[972])|(m[966]&~m[969]&~m[970]&m[971]&m[972])|(~m[966]&m[969]&~m[970]&m[971]&m[972])|(m[966]&m[969]&~m[970]&m[971]&m[972])|(~m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&m[969]&m[970]&m[971]&m[972]))):InitCond[296];
    m[973] = run?((((m[971]&~m[974]&~m[975]&~m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&m[976]&~m[977])|(m[971]&m[974]&~m[975]&m[976]&~m[977])|(m[971]&~m[974]&m[975]&m[976]&~m[977])|(~m[971]&m[974]&~m[975]&~m[976]&m[977])|(~m[971]&~m[974]&m[975]&~m[976]&m[977])|(m[971]&m[974]&m[975]&~m[976]&m[977])|(~m[971]&m[974]&m[975]&m[976]&m[977]))&UnbiasedRNG[41])|((m[971]&~m[974]&~m[975]&m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&m[975]&~m[976]&m[977])|(~m[971]&~m[974]&~m[975]&m[976]&m[977])|(m[971]&~m[974]&~m[975]&m[976]&m[977])|(~m[971]&m[974]&~m[975]&m[976]&m[977])|(m[971]&m[974]&~m[975]&m[976]&m[977])|(~m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&m[974]&m[975]&m[976]&m[977]))):InitCond[297];
    m[978] = run?((((m[677]&~m[979]&~m[980]&~m[981]&~m[982])|(~m[677]&~m[979]&~m[980]&m[981]&~m[982])|(m[677]&m[979]&~m[980]&m[981]&~m[982])|(m[677]&~m[979]&m[980]&m[981]&~m[982])|(~m[677]&m[979]&~m[980]&~m[981]&m[982])|(~m[677]&~m[979]&m[980]&~m[981]&m[982])|(m[677]&m[979]&m[980]&~m[981]&m[982])|(~m[677]&m[979]&m[980]&m[981]&m[982]))&UnbiasedRNG[42])|((m[677]&~m[979]&~m[980]&m[981]&~m[982])|(~m[677]&~m[979]&~m[980]&~m[981]&m[982])|(m[677]&~m[979]&~m[980]&~m[981]&m[982])|(m[677]&m[979]&~m[980]&~m[981]&m[982])|(m[677]&~m[979]&m[980]&~m[981]&m[982])|(~m[677]&~m[979]&~m[980]&m[981]&m[982])|(m[677]&~m[979]&~m[980]&m[981]&m[982])|(~m[677]&m[979]&~m[980]&m[981]&m[982])|(m[677]&m[979]&~m[980]&m[981]&m[982])|(~m[677]&~m[979]&m[980]&m[981]&m[982])|(m[677]&~m[979]&m[980]&m[981]&m[982])|(m[677]&m[979]&m[980]&m[981]&m[982]))):InitCond[298];
    m[983] = run?((((m[981]&~m[984]&~m[985]&~m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&m[986]&~m[987])|(m[981]&m[984]&~m[985]&m[986]&~m[987])|(m[981]&~m[984]&m[985]&m[986]&~m[987])|(~m[981]&m[984]&~m[985]&~m[986]&m[987])|(~m[981]&~m[984]&m[985]&~m[986]&m[987])|(m[981]&m[984]&m[985]&~m[986]&m[987])|(~m[981]&m[984]&m[985]&m[986]&m[987]))&UnbiasedRNG[43])|((m[981]&~m[984]&~m[985]&m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&m[985]&~m[986]&m[987])|(~m[981]&~m[984]&~m[985]&m[986]&m[987])|(m[981]&~m[984]&~m[985]&m[986]&m[987])|(~m[981]&m[984]&~m[985]&m[986]&m[987])|(m[981]&m[984]&~m[985]&m[986]&m[987])|(~m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&m[984]&m[985]&m[986]&m[987]))):InitCond[299];
    m[988] = run?((((m[986]&~m[989]&~m[990]&~m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&m[991]&~m[992])|(m[986]&m[989]&~m[990]&m[991]&~m[992])|(m[986]&~m[989]&m[990]&m[991]&~m[992])|(~m[986]&m[989]&~m[990]&~m[991]&m[992])|(~m[986]&~m[989]&m[990]&~m[991]&m[992])|(m[986]&m[989]&m[990]&~m[991]&m[992])|(~m[986]&m[989]&m[990]&m[991]&m[992]))&UnbiasedRNG[44])|((m[986]&~m[989]&~m[990]&m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&m[990]&~m[991]&m[992])|(~m[986]&~m[989]&~m[990]&m[991]&m[992])|(m[986]&~m[989]&~m[990]&m[991]&m[992])|(~m[986]&m[989]&~m[990]&m[991]&m[992])|(m[986]&m[989]&~m[990]&m[991]&m[992])|(~m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&m[989]&m[990]&m[991]&m[992]))):InitCond[300];
    m[993] = run?((((m[991]&~m[994]&~m[995]&~m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&m[996]&~m[997])|(m[991]&m[994]&~m[995]&m[996]&~m[997])|(m[991]&~m[994]&m[995]&m[996]&~m[997])|(~m[991]&m[994]&~m[995]&~m[996]&m[997])|(~m[991]&~m[994]&m[995]&~m[996]&m[997])|(m[991]&m[994]&m[995]&~m[996]&m[997])|(~m[991]&m[994]&m[995]&m[996]&m[997]))&UnbiasedRNG[45])|((m[991]&~m[994]&~m[995]&m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&m[995]&~m[996]&m[997])|(~m[991]&~m[994]&~m[995]&m[996]&m[997])|(m[991]&~m[994]&~m[995]&m[996]&m[997])|(~m[991]&m[994]&~m[995]&m[996]&m[997])|(m[991]&m[994]&~m[995]&m[996]&m[997])|(~m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&m[994]&m[995]&m[996]&m[997]))):InitCond[301];
    m[998] = run?((((m[996]&~m[999]&~m[1000]&~m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&~m[1002])|(~m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&m[999]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[46])|((m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&m[999]&m[1000]&m[1001]&m[1002]))):InitCond[302];
    m[1003] = run?((((m[678]&~m[1004]&~m[1005]&~m[1006]&~m[1007])|(~m[678]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(m[678]&m[1004]&~m[1005]&m[1006]&~m[1007])|(m[678]&~m[1004]&m[1005]&m[1006]&~m[1007])|(~m[678]&m[1004]&~m[1005]&~m[1006]&m[1007])|(~m[678]&~m[1004]&m[1005]&~m[1006]&m[1007])|(m[678]&m[1004]&m[1005]&~m[1006]&m[1007])|(~m[678]&m[1004]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[47])|((m[678]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(~m[678]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[678]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[678]&m[1004]&~m[1005]&~m[1006]&m[1007])|(m[678]&~m[1004]&m[1005]&~m[1006]&m[1007])|(~m[678]&~m[1004]&~m[1005]&m[1006]&m[1007])|(m[678]&~m[1004]&~m[1005]&m[1006]&m[1007])|(~m[678]&m[1004]&~m[1005]&m[1006]&m[1007])|(m[678]&m[1004]&~m[1005]&m[1006]&m[1007])|(~m[678]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[678]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[678]&m[1004]&m[1005]&m[1006]&m[1007]))):InitCond[303];
    m[1008] = run?((((m[1006]&~m[1009]&~m[1010]&~m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&~m[1012])|(~m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&m[1009]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[48])|((m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&m[1011]&m[1012]))):InitCond[304];
    m[1013] = run?((((m[1011]&~m[1014]&~m[1015]&~m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&~m[1017])|(~m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[49])|((m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))):InitCond[305];
    m[1018] = run?((((m[1016]&~m[1019]&~m[1020]&~m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&~m[1022])|(~m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[50])|((m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))):InitCond[306];
    m[1023] = run?((((m[1021]&~m[1024]&~m[1025]&~m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&~m[1027])|(~m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[51])|((m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))):InitCond[307];
    m[1028] = run?((((m[1026]&~m[1029]&~m[1030]&~m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&~m[1032])|(~m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[52])|((m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))):InitCond[308];
    m[1033] = run?((((m[679]&~m[1034]&~m[1035]&~m[1036]&~m[1037])|(~m[679]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(m[679]&m[1034]&~m[1035]&m[1036]&~m[1037])|(m[679]&~m[1034]&m[1035]&m[1036]&~m[1037])|(~m[679]&m[1034]&~m[1035]&~m[1036]&m[1037])|(~m[679]&~m[1034]&m[1035]&~m[1036]&m[1037])|(m[679]&m[1034]&m[1035]&~m[1036]&m[1037])|(~m[679]&m[1034]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[53])|((m[679]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(~m[679]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[679]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[679]&m[1034]&~m[1035]&~m[1036]&m[1037])|(m[679]&~m[1034]&m[1035]&~m[1036]&m[1037])|(~m[679]&~m[1034]&~m[1035]&m[1036]&m[1037])|(m[679]&~m[1034]&~m[1035]&m[1036]&m[1037])|(~m[679]&m[1034]&~m[1035]&m[1036]&m[1037])|(m[679]&m[1034]&~m[1035]&m[1036]&m[1037])|(~m[679]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[679]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[679]&m[1034]&m[1035]&m[1036]&m[1037]))):InitCond[309];
    m[1038] = run?((((m[1036]&~m[1039]&~m[1040]&~m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&~m[1042])|(~m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[54])|((m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))):InitCond[310];
    m[1043] = run?((((m[1041]&~m[1044]&~m[1045]&~m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&~m[1047])|(~m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[55])|((m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))):InitCond[311];
    m[1048] = run?((((m[1046]&~m[1049]&~m[1050]&~m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&~m[1052])|(~m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&m[1049]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[56])|((m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&m[1051]&m[1052]))):InitCond[312];
    m[1053] = run?((((m[1051]&~m[1054]&~m[1055]&~m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&~m[1057])|(~m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[57])|((m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))):InitCond[313];
    m[1058] = run?((((m[1056]&~m[1059]&~m[1060]&~m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&~m[1062])|(~m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&m[1059]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[58])|((m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&m[1061]&m[1062]))):InitCond[314];
    m[1063] = run?((((m[1061]&~m[1064]&~m[1065]&~m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&~m[1067])|(~m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[59])|((m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))):InitCond[315];
    m[1068] = run?((((m[680]&~m[1069]&~m[1070]&~m[1071]&~m[1072])|(~m[680]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(m[680]&m[1069]&~m[1070]&m[1071]&~m[1072])|(m[680]&~m[1069]&m[1070]&m[1071]&~m[1072])|(~m[680]&m[1069]&~m[1070]&~m[1071]&m[1072])|(~m[680]&~m[1069]&m[1070]&~m[1071]&m[1072])|(m[680]&m[1069]&m[1070]&~m[1071]&m[1072])|(~m[680]&m[1069]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[60])|((m[680]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(~m[680]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[680]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[680]&m[1069]&~m[1070]&~m[1071]&m[1072])|(m[680]&~m[1069]&m[1070]&~m[1071]&m[1072])|(~m[680]&~m[1069]&~m[1070]&m[1071]&m[1072])|(m[680]&~m[1069]&~m[1070]&m[1071]&m[1072])|(~m[680]&m[1069]&~m[1070]&m[1071]&m[1072])|(m[680]&m[1069]&~m[1070]&m[1071]&m[1072])|(~m[680]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[680]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[680]&m[1069]&m[1070]&m[1071]&m[1072]))):InitCond[316];
    m[1073] = run?((((m[1071]&~m[1074]&~m[1075]&~m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&~m[1077])|(~m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[61])|((m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))):InitCond[317];
    m[1078] = run?((((m[1076]&~m[1079]&~m[1080]&~m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&~m[1082])|(~m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[62])|((m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))):InitCond[318];
    m[1083] = run?((((m[1081]&~m[1084]&~m[1085]&~m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&~m[1087])|(~m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&m[1084]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[63])|((m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&m[1086]&m[1087]))):InitCond[319];
    m[1088] = run?((((m[1086]&~m[1089]&~m[1090]&~m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&~m[1092])|(~m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[64])|((m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))):InitCond[320];
    m[1093] = run?((((m[1091]&~m[1094]&~m[1095]&~m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&~m[1097])|(~m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[65])|((m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))):InitCond[321];
    m[1098] = run?((((m[1096]&~m[1099]&~m[1100]&~m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&~m[1102])|(~m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[66])|((m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))):InitCond[322];
    m[1103] = run?((((m[1101]&~m[1104]&~m[1105]&~m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&~m[1107])|(~m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[67])|((m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))):InitCond[323];
    m[1108] = run?((((m[681]&~m[1109]&~m[1110]&~m[1111]&~m[1112])|(~m[681]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(m[681]&m[1109]&~m[1110]&m[1111]&~m[1112])|(m[681]&~m[1109]&m[1110]&m[1111]&~m[1112])|(~m[681]&m[1109]&~m[1110]&~m[1111]&m[1112])|(~m[681]&~m[1109]&m[1110]&~m[1111]&m[1112])|(m[681]&m[1109]&m[1110]&~m[1111]&m[1112])|(~m[681]&m[1109]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[68])|((m[681]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(~m[681]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[681]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[681]&m[1109]&~m[1110]&~m[1111]&m[1112])|(m[681]&~m[1109]&m[1110]&~m[1111]&m[1112])|(~m[681]&~m[1109]&~m[1110]&m[1111]&m[1112])|(m[681]&~m[1109]&~m[1110]&m[1111]&m[1112])|(~m[681]&m[1109]&~m[1110]&m[1111]&m[1112])|(m[681]&m[1109]&~m[1110]&m[1111]&m[1112])|(~m[681]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[681]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[681]&m[1109]&m[1110]&m[1111]&m[1112]))):InitCond[324];
    m[1113] = run?((((m[1111]&~m[1114]&~m[1115]&~m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&~m[1117])|(~m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&m[1114]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[69])|((m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&m[1116]&m[1117]))):InitCond[325];
    m[1118] = run?((((m[1116]&~m[1119]&~m[1120]&~m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&~m[1122])|(~m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&m[1119]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[70])|((m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&m[1121]&m[1122]))):InitCond[326];
    m[1123] = run?((((m[1121]&~m[1124]&~m[1125]&~m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&~m[1127])|(~m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[71])|((m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))):InitCond[327];
    m[1128] = run?((((m[1126]&~m[1129]&~m[1130]&~m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&~m[1132])|(~m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[72])|((m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))):InitCond[328];
    m[1133] = run?((((m[1131]&~m[1134]&~m[1135]&~m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&~m[1137])|(~m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[73])|((m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))):InitCond[329];
    m[1138] = run?((((m[1136]&~m[1139]&~m[1140]&~m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&~m[1142])|(~m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&m[1139]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[74])|((m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&m[1141]&m[1142]))):InitCond[330];
    m[1143] = run?((((m[1141]&~m[1144]&~m[1145]&~m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&~m[1147])|(~m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[75])|((m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))):InitCond[331];
    m[1148] = run?((((m[1146]&~m[1149]&~m[1150]&~m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&~m[1152])|(~m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[76])|((m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))):InitCond[332];
    m[1153] = run?((((m[682]&~m[1154]&~m[1155]&~m[1156]&~m[1157])|(~m[682]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(m[682]&m[1154]&~m[1155]&m[1156]&~m[1157])|(m[682]&~m[1154]&m[1155]&m[1156]&~m[1157])|(~m[682]&m[1154]&~m[1155]&~m[1156]&m[1157])|(~m[682]&~m[1154]&m[1155]&~m[1156]&m[1157])|(m[682]&m[1154]&m[1155]&~m[1156]&m[1157])|(~m[682]&m[1154]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[77])|((m[682]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(~m[682]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[682]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[682]&m[1154]&~m[1155]&~m[1156]&m[1157])|(m[682]&~m[1154]&m[1155]&~m[1156]&m[1157])|(~m[682]&~m[1154]&~m[1155]&m[1156]&m[1157])|(m[682]&~m[1154]&~m[1155]&m[1156]&m[1157])|(~m[682]&m[1154]&~m[1155]&m[1156]&m[1157])|(m[682]&m[1154]&~m[1155]&m[1156]&m[1157])|(~m[682]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[682]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[682]&m[1154]&m[1155]&m[1156]&m[1157]))):InitCond[333];
    m[1158] = run?((((m[1156]&~m[1159]&~m[1160]&~m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&~m[1162])|(~m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&m[1159]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[78])|((m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&m[1161]&m[1162]))):InitCond[334];
    m[1163] = run?((((m[1161]&~m[1164]&~m[1165]&~m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&~m[1167])|(~m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[79])|((m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))):InitCond[335];
    m[1168] = run?((((m[1166]&~m[1169]&~m[1170]&~m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&~m[1172])|(~m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[80])|((m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))):InitCond[336];
    m[1173] = run?((((m[1171]&~m[1174]&~m[1175]&~m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&~m[1177])|(~m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&m[1174]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[81])|((m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&m[1176]&m[1177]))):InitCond[337];
    m[1178] = run?((((m[1176]&~m[1179]&~m[1180]&~m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&~m[1182])|(~m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[82])|((m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))):InitCond[338];
    m[1183] = run?((((m[1181]&~m[1184]&~m[1185]&~m[1186]&~m[1187])|(~m[1181]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1181]&m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1181]&~m[1184]&m[1185]&m[1186]&~m[1187])|(~m[1181]&m[1184]&~m[1185]&~m[1186]&m[1187])|(~m[1181]&~m[1184]&m[1185]&~m[1186]&m[1187])|(m[1181]&m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1181]&m[1184]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[83])|((m[1181]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(~m[1181]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1181]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1181]&m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1181]&~m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1181]&~m[1184]&~m[1185]&m[1186]&m[1187])|(m[1181]&~m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1181]&m[1184]&~m[1185]&m[1186]&m[1187])|(m[1181]&m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1181]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1181]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1181]&m[1184]&m[1185]&m[1186]&m[1187]))):InitCond[339];
    m[1188] = run?((((m[1186]&~m[1189]&~m[1190]&~m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&~m[1192])|(~m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&m[1189]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[84])|((m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&m[1191]&m[1192]))):InitCond[340];
    m[1193] = run?((((m[1191]&~m[1194]&~m[1195]&~m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&~m[1197])|(~m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&m[1194]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[85])|((m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&m[1196]&m[1197]))):InitCond[341];
    m[1198] = run?((((m[1196]&~m[1199]&~m[1200]&~m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&~m[1202])|(~m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&m[1199]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[86])|((m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&m[1201]&m[1202]))):InitCond[342];
    m[1203] = run?((((m[683]&~m[1204]&~m[1205]&~m[1206]&~m[1207])|(~m[683]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(m[683]&m[1204]&~m[1205]&m[1206]&~m[1207])|(m[683]&~m[1204]&m[1205]&m[1206]&~m[1207])|(~m[683]&m[1204]&~m[1205]&~m[1206]&m[1207])|(~m[683]&~m[1204]&m[1205]&~m[1206]&m[1207])|(m[683]&m[1204]&m[1205]&~m[1206]&m[1207])|(~m[683]&m[1204]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[87])|((m[683]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(~m[683]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[683]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[683]&m[1204]&~m[1205]&~m[1206]&m[1207])|(m[683]&~m[1204]&m[1205]&~m[1206]&m[1207])|(~m[683]&~m[1204]&~m[1205]&m[1206]&m[1207])|(m[683]&~m[1204]&~m[1205]&m[1206]&m[1207])|(~m[683]&m[1204]&~m[1205]&m[1206]&m[1207])|(m[683]&m[1204]&~m[1205]&m[1206]&m[1207])|(~m[683]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[683]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[683]&m[1204]&m[1205]&m[1206]&m[1207]))):InitCond[343];
    m[1208] = run?((((m[1206]&~m[1209]&~m[1210]&~m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&~m[1212])|(~m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&m[1209]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[88])|((m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&m[1211]&m[1212]))):InitCond[344];
    m[1213] = run?((((m[1211]&~m[1214]&~m[1215]&~m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&~m[1217])|(~m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&m[1214]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[89])|((m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&m[1216]&m[1217]))):InitCond[345];
    m[1218] = run?((((m[1216]&~m[1219]&~m[1220]&~m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&~m[1222])|(~m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&m[1219]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[90])|((m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&m[1221]&m[1222]))):InitCond[346];
    m[1223] = run?((((m[1221]&~m[1224]&~m[1225]&~m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&~m[1227])|(~m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&m[1224]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[91])|((m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&m[1226]&m[1227]))):InitCond[347];
    m[1228] = run?((((m[1226]&~m[1229]&~m[1230]&~m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&~m[1232])|(~m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&m[1229]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[92])|((m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&m[1231]&m[1232]))):InitCond[348];
    m[1233] = run?((((m[1231]&~m[1234]&~m[1235]&~m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&~m[1237])|(~m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&m[1234]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[93])|((m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&m[1236]&m[1237]))):InitCond[349];
    m[1238] = run?((((m[1236]&~m[1239]&~m[1240]&~m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&~m[1242])|(~m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&m[1239]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[94])|((m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&m[1241]&m[1242]))):InitCond[350];
    m[1243] = run?((((m[1241]&~m[1244]&~m[1245]&~m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&~m[1247])|(~m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&m[1244]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[95])|((m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&m[1246]&m[1247]))):InitCond[351];
    m[1248] = run?((((m[1246]&~m[1249]&~m[1250]&~m[1251]&~m[1252])|(~m[1246]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1246]&m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1246]&~m[1249]&m[1250]&m[1251]&~m[1252])|(~m[1246]&m[1249]&~m[1250]&~m[1251]&m[1252])|(~m[1246]&~m[1249]&m[1250]&~m[1251]&m[1252])|(m[1246]&m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1246]&m[1249]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[96])|((m[1246]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(~m[1246]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1246]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1246]&m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1246]&~m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1246]&~m[1249]&~m[1250]&m[1251]&m[1252])|(m[1246]&~m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1246]&m[1249]&~m[1250]&m[1251]&m[1252])|(m[1246]&m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1246]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1246]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1246]&m[1249]&m[1250]&m[1251]&m[1252]))):InitCond[352];
    m[1253] = run?((((m[1251]&~m[1254]&~m[1255]&~m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&~m[1257])|(~m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&m[1254]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[97])|((m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&m[1256]&m[1257]))):InitCond[353];
    m[1258] = run?((((m[684]&~m[1259]&~m[1260]&~m[1261]&~m[1262])|(~m[684]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(m[684]&m[1259]&~m[1260]&m[1261]&~m[1262])|(m[684]&~m[1259]&m[1260]&m[1261]&~m[1262])|(~m[684]&m[1259]&~m[1260]&~m[1261]&m[1262])|(~m[684]&~m[1259]&m[1260]&~m[1261]&m[1262])|(m[684]&m[1259]&m[1260]&~m[1261]&m[1262])|(~m[684]&m[1259]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[98])|((m[684]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(~m[684]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[684]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[684]&m[1259]&~m[1260]&~m[1261]&m[1262])|(m[684]&~m[1259]&m[1260]&~m[1261]&m[1262])|(~m[684]&~m[1259]&~m[1260]&m[1261]&m[1262])|(m[684]&~m[1259]&~m[1260]&m[1261]&m[1262])|(~m[684]&m[1259]&~m[1260]&m[1261]&m[1262])|(m[684]&m[1259]&~m[1260]&m[1261]&m[1262])|(~m[684]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[684]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[684]&m[1259]&m[1260]&m[1261]&m[1262]))):InitCond[354];
    m[1263] = run?((((m[1261]&~m[1264]&~m[1265]&~m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&~m[1267])|(~m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&m[1264]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[99])|((m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&m[1266]&m[1267]))):InitCond[355];
    m[1268] = run?((((m[1266]&~m[1269]&~m[1270]&~m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&~m[1272])|(~m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&m[1269]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[100])|((m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&m[1271]&m[1272]))):InitCond[356];
    m[1273] = run?((((m[1271]&~m[1274]&~m[1275]&~m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&~m[1277])|(~m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&m[1274]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[101])|((m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&m[1276]&m[1277]))):InitCond[357];
    m[1278] = run?((((m[1276]&~m[1279]&~m[1280]&~m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&~m[1282])|(~m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&m[1279]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[102])|((m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&m[1281]&m[1282]))):InitCond[358];
    m[1283] = run?((((m[1281]&~m[1284]&~m[1285]&~m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&~m[1287])|(~m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&m[1284]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[103])|((m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&m[1286]&m[1287]))):InitCond[359];
    m[1288] = run?((((m[1286]&~m[1289]&~m[1290]&~m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&~m[1292])|(~m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&m[1289]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[104])|((m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&m[1291]&m[1292]))):InitCond[360];
    m[1293] = run?((((m[1291]&~m[1294]&~m[1295]&~m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&~m[1297])|(~m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&m[1294]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[105])|((m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&m[1296]&m[1297]))):InitCond[361];
    m[1298] = run?((((m[1296]&~m[1299]&~m[1300]&~m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&~m[1302])|(~m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&m[1299]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[106])|((m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&m[1301]&m[1302]))):InitCond[362];
    m[1303] = run?((((m[1301]&~m[1304]&~m[1305]&~m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&~m[1307])|(~m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&m[1304]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[107])|((m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&m[1306]&m[1307]))):InitCond[363];
    m[1308] = run?((((m[1306]&~m[1309]&~m[1310]&~m[1311]&~m[1312])|(~m[1306]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1306]&m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1306]&~m[1309]&m[1310]&m[1311]&~m[1312])|(~m[1306]&m[1309]&~m[1310]&~m[1311]&m[1312])|(~m[1306]&~m[1309]&m[1310]&~m[1311]&m[1312])|(m[1306]&m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1306]&m[1309]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[108])|((m[1306]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(~m[1306]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1306]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1306]&m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1306]&~m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1306]&~m[1309]&~m[1310]&m[1311]&m[1312])|(m[1306]&~m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1306]&m[1309]&~m[1310]&m[1311]&m[1312])|(m[1306]&m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1306]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1306]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1306]&m[1309]&m[1310]&m[1311]&m[1312]))):InitCond[364];
    m[1313] = run?((((m[1311]&~m[1314]&~m[1315]&~m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&~m[1317])|(~m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&m[1314]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[109])|((m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&m[1316]&m[1317]))):InitCond[365];
    m[1318] = run?((((m[685]&~m[1319]&~m[1320]&~m[1321]&~m[1322])|(~m[685]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(m[685]&m[1319]&~m[1320]&m[1321]&~m[1322])|(m[685]&~m[1319]&m[1320]&m[1321]&~m[1322])|(~m[685]&m[1319]&~m[1320]&~m[1321]&m[1322])|(~m[685]&~m[1319]&m[1320]&~m[1321]&m[1322])|(m[685]&m[1319]&m[1320]&~m[1321]&m[1322])|(~m[685]&m[1319]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[110])|((m[685]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(~m[685]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[685]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[685]&m[1319]&~m[1320]&~m[1321]&m[1322])|(m[685]&~m[1319]&m[1320]&~m[1321]&m[1322])|(~m[685]&~m[1319]&~m[1320]&m[1321]&m[1322])|(m[685]&~m[1319]&~m[1320]&m[1321]&m[1322])|(~m[685]&m[1319]&~m[1320]&m[1321]&m[1322])|(m[685]&m[1319]&~m[1320]&m[1321]&m[1322])|(~m[685]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[685]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[685]&m[1319]&m[1320]&m[1321]&m[1322]))):InitCond[366];
    m[1323] = run?((((m[1321]&~m[1324]&~m[1325]&~m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&~m[1327])|(~m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&m[1324]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[111])|((m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&m[1326]&m[1327]))):InitCond[367];
    m[1328] = run?((((m[1326]&~m[1329]&~m[1330]&~m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&~m[1332])|(~m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&m[1329]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[112])|((m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&m[1331]&m[1332]))):InitCond[368];
    m[1333] = run?((((m[1331]&~m[1334]&~m[1335]&~m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&~m[1337])|(~m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&m[1334]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[113])|((m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&m[1336]&m[1337]))):InitCond[369];
    m[1338] = run?((((m[1336]&~m[1339]&~m[1340]&~m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&~m[1342])|(~m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&m[1339]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[114])|((m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&m[1341]&m[1342]))):InitCond[370];
    m[1343] = run?((((m[1341]&~m[1344]&~m[1345]&~m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&~m[1347])|(~m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&m[1344]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[115])|((m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&m[1346]&m[1347]))):InitCond[371];
    m[1348] = run?((((m[1346]&~m[1349]&~m[1350]&~m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&~m[1352])|(~m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&m[1349]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[116])|((m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&m[1351]&m[1352]))):InitCond[372];
    m[1353] = run?((((m[1351]&~m[1354]&~m[1355]&~m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&~m[1357])|(~m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&m[1354]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[117])|((m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&m[1356]&m[1357]))):InitCond[373];
    m[1358] = run?((((m[1356]&~m[1359]&~m[1360]&~m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&~m[1362])|(~m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&m[1359]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[118])|((m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&m[1361]&m[1362]))):InitCond[374];
    m[1363] = run?((((m[1361]&~m[1364]&~m[1365]&~m[1366]&~m[1367])|(~m[1361]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1361]&m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1361]&~m[1364]&m[1365]&m[1366]&~m[1367])|(~m[1361]&m[1364]&~m[1365]&~m[1366]&m[1367])|(~m[1361]&~m[1364]&m[1365]&~m[1366]&m[1367])|(m[1361]&m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1361]&m[1364]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[119])|((m[1361]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(~m[1361]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1361]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1361]&m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1361]&~m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1361]&~m[1364]&~m[1365]&m[1366]&m[1367])|(m[1361]&~m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1361]&m[1364]&~m[1365]&m[1366]&m[1367])|(m[1361]&m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1361]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1361]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1361]&m[1364]&m[1365]&m[1366]&m[1367]))):InitCond[375];
    m[1368] = run?((((m[1366]&~m[1369]&~m[1370]&~m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&~m[1372])|(~m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&m[1369]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[120])|((m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&m[1371]&m[1372]))):InitCond[376];
    m[1373] = run?((((m[1371]&~m[1374]&~m[1375]&~m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&~m[1377])|(~m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&m[1374]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[121])|((m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&m[1376]&m[1377]))):InitCond[377];
    m[1378] = run?((((m[1376]&~m[1379]&~m[1380]&~m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&~m[1382])|(~m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&m[1379]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[122])|((m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&m[1381]&m[1382]))):InitCond[378];
    m[1383] = run?((((m[686]&~m[1384]&~m[1385]&~m[1386]&~m[1387])|(~m[686]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(m[686]&m[1384]&~m[1385]&m[1386]&~m[1387])|(m[686]&~m[1384]&m[1385]&m[1386]&~m[1387])|(~m[686]&m[1384]&~m[1385]&~m[1386]&m[1387])|(~m[686]&~m[1384]&m[1385]&~m[1386]&m[1387])|(m[686]&m[1384]&m[1385]&~m[1386]&m[1387])|(~m[686]&m[1384]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[123])|((m[686]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(~m[686]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[686]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[686]&m[1384]&~m[1385]&~m[1386]&m[1387])|(m[686]&~m[1384]&m[1385]&~m[1386]&m[1387])|(~m[686]&~m[1384]&~m[1385]&m[1386]&m[1387])|(m[686]&~m[1384]&~m[1385]&m[1386]&m[1387])|(~m[686]&m[1384]&~m[1385]&m[1386]&m[1387])|(m[686]&m[1384]&~m[1385]&m[1386]&m[1387])|(~m[686]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[686]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[686]&m[1384]&m[1385]&m[1386]&m[1387]))):InitCond[379];
    m[1388] = run?((((m[1386]&~m[1389]&~m[1390]&~m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&~m[1392])|(~m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&m[1389]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[124])|((m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&m[1391]&m[1392]))):InitCond[380];
    m[1393] = run?((((m[1391]&~m[1394]&~m[1395]&~m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&~m[1397])|(~m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&m[1394]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[125])|((m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&m[1396]&m[1397]))):InitCond[381];
    m[1398] = run?((((m[1396]&~m[1399]&~m[1400]&~m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&~m[1402])|(~m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&m[1399]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[126])|((m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&m[1401]&m[1402]))):InitCond[382];
    m[1403] = run?((((m[1401]&~m[1404]&~m[1405]&~m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&~m[1407])|(~m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&m[1404]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[127])|((m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&m[1406]&m[1407]))):InitCond[383];
    m[1408] = run?((((m[1406]&~m[1409]&~m[1410]&~m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&~m[1412])|(~m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&m[1409]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[128])|((m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&m[1411]&m[1412]))):InitCond[384];
    m[1413] = run?((((m[1411]&~m[1414]&~m[1415]&~m[1416]&~m[1417])|(~m[1411]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1411]&m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1411]&~m[1414]&m[1415]&m[1416]&~m[1417])|(~m[1411]&m[1414]&~m[1415]&~m[1416]&m[1417])|(~m[1411]&~m[1414]&m[1415]&~m[1416]&m[1417])|(m[1411]&m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1411]&m[1414]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[129])|((m[1411]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(~m[1411]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1411]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1411]&m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1411]&~m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1411]&~m[1414]&~m[1415]&m[1416]&m[1417])|(m[1411]&~m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1411]&m[1414]&~m[1415]&m[1416]&m[1417])|(m[1411]&m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1411]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1411]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1411]&m[1414]&m[1415]&m[1416]&m[1417]))):InitCond[385];
    m[1418] = run?((((m[1416]&~m[1419]&~m[1420]&~m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&~m[1422])|(~m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&m[1419]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[130])|((m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&m[1421]&m[1422]))):InitCond[386];
    m[1423] = run?((((m[1421]&~m[1424]&~m[1425]&~m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&~m[1427])|(~m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&m[1424]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[131])|((m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&m[1426]&m[1427]))):InitCond[387];
    m[1428] = run?((((m[1426]&~m[1429]&~m[1430]&~m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&~m[1432])|(~m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&m[1429]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[132])|((m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&m[1431]&m[1432]))):InitCond[388];
    m[1433] = run?((((m[1431]&~m[1434]&~m[1435]&~m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&~m[1437])|(~m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&m[1434]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[133])|((m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&m[1436]&m[1437]))):InitCond[389];
    m[1438] = run?((((m[1436]&~m[1439]&~m[1440]&~m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&~m[1442])|(~m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&m[1439]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[134])|((m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&m[1441]&m[1442]))):InitCond[390];
    m[1443] = run?((((m[1441]&~m[1444]&~m[1445]&~m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&~m[1447])|(~m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&m[1444]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[135])|((m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&m[1446]&m[1447]))):InitCond[391];
    m[1448] = run?((((m[1446]&~m[1449]&~m[1450]&~m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&~m[1452])|(~m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&m[1449]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[136])|((m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&m[1451]&m[1452]))):InitCond[392];
    m[1453] = run?((((m[687]&~m[1454]&~m[1455]&~m[1456]&~m[1457])|(~m[687]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(m[687]&m[1454]&~m[1455]&m[1456]&~m[1457])|(m[687]&~m[1454]&m[1455]&m[1456]&~m[1457])|(~m[687]&m[1454]&~m[1455]&~m[1456]&m[1457])|(~m[687]&~m[1454]&m[1455]&~m[1456]&m[1457])|(m[687]&m[1454]&m[1455]&~m[1456]&m[1457])|(~m[687]&m[1454]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[137])|((m[687]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(~m[687]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[687]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[687]&m[1454]&~m[1455]&~m[1456]&m[1457])|(m[687]&~m[1454]&m[1455]&~m[1456]&m[1457])|(~m[687]&~m[1454]&~m[1455]&m[1456]&m[1457])|(m[687]&~m[1454]&~m[1455]&m[1456]&m[1457])|(~m[687]&m[1454]&~m[1455]&m[1456]&m[1457])|(m[687]&m[1454]&~m[1455]&m[1456]&m[1457])|(~m[687]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[687]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[687]&m[1454]&m[1455]&m[1456]&m[1457]))):InitCond[393];
    m[1458] = run?((((m[1456]&~m[1459]&~m[1460]&~m[1461]&~m[1462])|(~m[1456]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1456]&m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1456]&~m[1459]&m[1460]&m[1461]&~m[1462])|(~m[1456]&m[1459]&~m[1460]&~m[1461]&m[1462])|(~m[1456]&~m[1459]&m[1460]&~m[1461]&m[1462])|(m[1456]&m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1456]&m[1459]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[138])|((m[1456]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(~m[1456]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1456]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1456]&m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1456]&~m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1456]&~m[1459]&~m[1460]&m[1461]&m[1462])|(m[1456]&~m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1456]&m[1459]&~m[1460]&m[1461]&m[1462])|(m[1456]&m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1456]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1456]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1456]&m[1459]&m[1460]&m[1461]&m[1462]))):InitCond[394];
    m[1463] = run?((((m[1461]&~m[1464]&~m[1465]&~m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&~m[1467])|(~m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&m[1464]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[139])|((m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&m[1466]&m[1467]))):InitCond[395];
    m[1468] = run?((((m[1466]&~m[1469]&~m[1470]&~m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&~m[1472])|(~m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&m[1469]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[140])|((m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&m[1471]&m[1472]))):InitCond[396];
    m[1473] = run?((((m[1471]&~m[1474]&~m[1475]&~m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&~m[1477])|(~m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&m[1474]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[141])|((m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&m[1476]&m[1477]))):InitCond[397];
    m[1478] = run?((((m[1476]&~m[1479]&~m[1480]&~m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&~m[1482])|(~m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&m[1479]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[142])|((m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&m[1481]&m[1482]))):InitCond[398];
    m[1483] = run?((((m[1481]&~m[1484]&~m[1485]&~m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&~m[1487])|(~m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&m[1484]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[143])|((m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&m[1486]&m[1487]))):InitCond[399];
    m[1488] = run?((((m[1486]&~m[1489]&~m[1490]&~m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&~m[1492])|(~m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&m[1489]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[144])|((m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&m[1491]&m[1492]))):InitCond[400];
    m[1493] = run?((((m[1491]&~m[1494]&~m[1495]&~m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&~m[1497])|(~m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&m[1494]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[145])|((m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&m[1496]&m[1497]))):InitCond[401];
    m[1498] = run?((((m[1496]&~m[1499]&~m[1500]&~m[1501]&~m[1502])|(~m[1496]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1496]&m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1496]&~m[1499]&m[1500]&m[1501]&~m[1502])|(~m[1496]&m[1499]&~m[1500]&~m[1501]&m[1502])|(~m[1496]&~m[1499]&m[1500]&~m[1501]&m[1502])|(m[1496]&m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1496]&m[1499]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[146])|((m[1496]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(~m[1496]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1496]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1496]&m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1496]&~m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1496]&~m[1499]&~m[1500]&m[1501]&m[1502])|(m[1496]&~m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1496]&m[1499]&~m[1500]&m[1501]&m[1502])|(m[1496]&m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1496]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1496]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1496]&m[1499]&m[1500]&m[1501]&m[1502]))):InitCond[402];
    m[1503] = run?((((m[1501]&~m[1504]&~m[1505]&~m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&~m[1507])|(~m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&m[1504]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[147])|((m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&m[1506]&m[1507]))):InitCond[403];
    m[1508] = run?((((m[1506]&~m[1509]&~m[1510]&~m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&~m[1512])|(~m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&m[1509]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[148])|((m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&m[1511]&m[1512]))):InitCond[404];
    m[1513] = run?((((m[1511]&~m[1514]&~m[1515]&~m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&~m[1517])|(~m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&m[1514]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[149])|((m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&m[1516]&m[1517]))):InitCond[405];
    m[1518] = run?((((m[1516]&~m[1519]&~m[1520]&~m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&~m[1522])|(~m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&m[1519]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[150])|((m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&m[1521]&m[1522]))):InitCond[406];
    m[1523] = run?((((m[1521]&~m[1524]&~m[1525]&~m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&~m[1527])|(~m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&m[1524]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[151])|((m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&m[1526]&m[1527]))):InitCond[407];
    m[1533] = run?((((m[1531]&~m[1534]&~m[1535]&~m[1536]&~m[1537])|(~m[1531]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1531]&m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1531]&~m[1534]&m[1535]&m[1536]&~m[1537])|(~m[1531]&m[1534]&~m[1535]&~m[1536]&m[1537])|(~m[1531]&~m[1534]&m[1535]&~m[1536]&m[1537])|(m[1531]&m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1531]&m[1534]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[152])|((m[1531]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(~m[1531]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1531]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1531]&m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1531]&~m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1531]&~m[1534]&~m[1535]&m[1536]&m[1537])|(m[1531]&~m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1531]&m[1534]&~m[1535]&m[1536]&m[1537])|(m[1531]&m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1531]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1531]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1531]&m[1534]&m[1535]&m[1536]&m[1537]))):InitCond[408];
    m[1538] = run?((((m[1536]&~m[1539]&~m[1540]&~m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&~m[1542])|(~m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&m[1539]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[153])|((m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&m[1541]&m[1542]))):InitCond[409];
    m[1543] = run?((((m[1541]&~m[1544]&~m[1545]&~m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&~m[1547])|(~m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&m[1544]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[154])|((m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&m[1546]&m[1547]))):InitCond[410];
    m[1548] = run?((((m[1546]&~m[1549]&~m[1550]&~m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&~m[1552])|(~m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&m[1549]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[155])|((m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&m[1551]&m[1552]))):InitCond[411];
    m[1553] = run?((((m[1551]&~m[1554]&~m[1555]&~m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&~m[1557])|(~m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&m[1554]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[156])|((m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&m[1556]&m[1557]))):InitCond[412];
    m[1558] = run?((((m[1556]&~m[1559]&~m[1560]&~m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&~m[1562])|(~m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&m[1559]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[157])|((m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&m[1561]&m[1562]))):InitCond[413];
    m[1563] = run?((((m[1561]&~m[1564]&~m[1565]&~m[1566]&~m[1567])|(~m[1561]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1561]&m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1561]&~m[1564]&m[1565]&m[1566]&~m[1567])|(~m[1561]&m[1564]&~m[1565]&~m[1566]&m[1567])|(~m[1561]&~m[1564]&m[1565]&~m[1566]&m[1567])|(m[1561]&m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1561]&m[1564]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[158])|((m[1561]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(~m[1561]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1561]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1561]&m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1561]&~m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1561]&~m[1564]&~m[1565]&m[1566]&m[1567])|(m[1561]&~m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1561]&m[1564]&~m[1565]&m[1566]&m[1567])|(m[1561]&m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1561]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1561]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1561]&m[1564]&m[1565]&m[1566]&m[1567]))):InitCond[414];
    m[1568] = run?((((m[1566]&~m[1569]&~m[1570]&~m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&~m[1572])|(~m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&m[1569]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[159])|((m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&m[1571]&m[1572]))):InitCond[415];
    m[1573] = run?((((m[1571]&~m[1574]&~m[1575]&~m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&~m[1577])|(~m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&m[1574]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[160])|((m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&m[1576]&m[1577]))):InitCond[416];
    m[1578] = run?((((m[1576]&~m[1579]&~m[1580]&~m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&~m[1582])|(~m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&m[1579]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[161])|((m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&m[1581]&m[1582]))):InitCond[417];
    m[1583] = run?((((m[1581]&~m[1584]&~m[1585]&~m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&~m[1587])|(~m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&m[1584]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[162])|((m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&m[1586]&m[1587]))):InitCond[418];
    m[1588] = run?((((m[1586]&~m[1589]&~m[1590]&~m[1591]&~m[1592])|(~m[1586]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1586]&m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1586]&~m[1589]&m[1590]&m[1591]&~m[1592])|(~m[1586]&m[1589]&~m[1590]&~m[1591]&m[1592])|(~m[1586]&~m[1589]&m[1590]&~m[1591]&m[1592])|(m[1586]&m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1586]&m[1589]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[163])|((m[1586]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(~m[1586]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1586]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1586]&m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1586]&~m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1586]&~m[1589]&~m[1590]&m[1591]&m[1592])|(m[1586]&~m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1586]&m[1589]&~m[1590]&m[1591]&m[1592])|(m[1586]&m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1586]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1586]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1586]&m[1589]&m[1590]&m[1591]&m[1592]))):InitCond[419];
    m[1593] = run?((((m[1591]&~m[1594]&~m[1595]&~m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&~m[1597])|(~m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&m[1594]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[164])|((m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&m[1596]&m[1597]))):InitCond[420];
    m[1598] = run?((((m[1596]&~m[1599]&~m[1600]&~m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&~m[1602])|(~m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&m[1599]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[165])|((m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&m[1601]&m[1602]))):InitCond[421];
    m[1603] = run?((((m[1532]&~m[1604]&~m[1605]&~m[1606]&~m[1607])|(~m[1532]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1532]&m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1532]&~m[1604]&m[1605]&m[1606]&~m[1607])|(~m[1532]&m[1604]&~m[1605]&~m[1606]&m[1607])|(~m[1532]&~m[1604]&m[1605]&~m[1606]&m[1607])|(m[1532]&m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1532]&m[1604]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[166])|((m[1532]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(~m[1532]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1532]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1532]&m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1532]&~m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1532]&~m[1604]&~m[1605]&m[1606]&m[1607])|(m[1532]&~m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1532]&m[1604]&~m[1605]&m[1606]&m[1607])|(m[1532]&m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1532]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1532]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1532]&m[1604]&m[1605]&m[1606]&m[1607]))):InitCond[422];
    m[1608] = run?((((m[1606]&~m[1609]&~m[1610]&~m[1611]&~m[1612])|(~m[1606]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1606]&m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1606]&~m[1609]&m[1610]&m[1611]&~m[1612])|(~m[1606]&m[1609]&~m[1610]&~m[1611]&m[1612])|(~m[1606]&~m[1609]&m[1610]&~m[1611]&m[1612])|(m[1606]&m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1606]&m[1609]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[167])|((m[1606]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(~m[1606]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1606]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1606]&m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1606]&~m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1606]&~m[1609]&~m[1610]&m[1611]&m[1612])|(m[1606]&~m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1606]&m[1609]&~m[1610]&m[1611]&m[1612])|(m[1606]&m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1606]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1606]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1606]&m[1609]&m[1610]&m[1611]&m[1612]))):InitCond[423];
    m[1613] = run?((((m[1611]&~m[1614]&~m[1615]&~m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&~m[1617])|(~m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&m[1614]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[168])|((m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&m[1616]&m[1617]))):InitCond[424];
    m[1618] = run?((((m[1616]&~m[1619]&~m[1620]&~m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&~m[1622])|(~m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&m[1619]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[169])|((m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&m[1621]&m[1622]))):InitCond[425];
    m[1623] = run?((((m[1621]&~m[1624]&~m[1625]&~m[1626]&~m[1627])|(~m[1621]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1621]&m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1621]&~m[1624]&m[1625]&m[1626]&~m[1627])|(~m[1621]&m[1624]&~m[1625]&~m[1626]&m[1627])|(~m[1621]&~m[1624]&m[1625]&~m[1626]&m[1627])|(m[1621]&m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1621]&m[1624]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[170])|((m[1621]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(~m[1621]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1621]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1621]&m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1621]&~m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1621]&~m[1624]&~m[1625]&m[1626]&m[1627])|(m[1621]&~m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1621]&m[1624]&~m[1625]&m[1626]&m[1627])|(m[1621]&m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1621]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1621]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1621]&m[1624]&m[1625]&m[1626]&m[1627]))):InitCond[426];
    m[1628] = run?((((m[1626]&~m[1629]&~m[1630]&~m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&~m[1632])|(~m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&m[1629]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[171])|((m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&m[1631]&m[1632]))):InitCond[427];
    m[1633] = run?((((m[1631]&~m[1634]&~m[1635]&~m[1636]&~m[1637])|(~m[1631]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1631]&m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1631]&~m[1634]&m[1635]&m[1636]&~m[1637])|(~m[1631]&m[1634]&~m[1635]&~m[1636]&m[1637])|(~m[1631]&~m[1634]&m[1635]&~m[1636]&m[1637])|(m[1631]&m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1631]&m[1634]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[172])|((m[1631]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(~m[1631]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1631]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1631]&m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1631]&~m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1631]&~m[1634]&~m[1635]&m[1636]&m[1637])|(m[1631]&~m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1631]&m[1634]&~m[1635]&m[1636]&m[1637])|(m[1631]&m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1631]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1631]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1631]&m[1634]&m[1635]&m[1636]&m[1637]))):InitCond[428];
    m[1638] = run?((((m[1636]&~m[1639]&~m[1640]&~m[1641]&~m[1642])|(~m[1636]&~m[1639]&~m[1640]&m[1641]&~m[1642])|(m[1636]&m[1639]&~m[1640]&m[1641]&~m[1642])|(m[1636]&~m[1639]&m[1640]&m[1641]&~m[1642])|(~m[1636]&m[1639]&~m[1640]&~m[1641]&m[1642])|(~m[1636]&~m[1639]&m[1640]&~m[1641]&m[1642])|(m[1636]&m[1639]&m[1640]&~m[1641]&m[1642])|(~m[1636]&m[1639]&m[1640]&m[1641]&m[1642]))&UnbiasedRNG[173])|((m[1636]&~m[1639]&~m[1640]&m[1641]&~m[1642])|(~m[1636]&~m[1639]&~m[1640]&~m[1641]&m[1642])|(m[1636]&~m[1639]&~m[1640]&~m[1641]&m[1642])|(m[1636]&m[1639]&~m[1640]&~m[1641]&m[1642])|(m[1636]&~m[1639]&m[1640]&~m[1641]&m[1642])|(~m[1636]&~m[1639]&~m[1640]&m[1641]&m[1642])|(m[1636]&~m[1639]&~m[1640]&m[1641]&m[1642])|(~m[1636]&m[1639]&~m[1640]&m[1641]&m[1642])|(m[1636]&m[1639]&~m[1640]&m[1641]&m[1642])|(~m[1636]&~m[1639]&m[1640]&m[1641]&m[1642])|(m[1636]&~m[1639]&m[1640]&m[1641]&m[1642])|(m[1636]&m[1639]&m[1640]&m[1641]&m[1642]))):InitCond[429];
    m[1643] = run?((((m[1641]&~m[1644]&~m[1645]&~m[1646]&~m[1647])|(~m[1641]&~m[1644]&~m[1645]&m[1646]&~m[1647])|(m[1641]&m[1644]&~m[1645]&m[1646]&~m[1647])|(m[1641]&~m[1644]&m[1645]&m[1646]&~m[1647])|(~m[1641]&m[1644]&~m[1645]&~m[1646]&m[1647])|(~m[1641]&~m[1644]&m[1645]&~m[1646]&m[1647])|(m[1641]&m[1644]&m[1645]&~m[1646]&m[1647])|(~m[1641]&m[1644]&m[1645]&m[1646]&m[1647]))&UnbiasedRNG[174])|((m[1641]&~m[1644]&~m[1645]&m[1646]&~m[1647])|(~m[1641]&~m[1644]&~m[1645]&~m[1646]&m[1647])|(m[1641]&~m[1644]&~m[1645]&~m[1646]&m[1647])|(m[1641]&m[1644]&~m[1645]&~m[1646]&m[1647])|(m[1641]&~m[1644]&m[1645]&~m[1646]&m[1647])|(~m[1641]&~m[1644]&~m[1645]&m[1646]&m[1647])|(m[1641]&~m[1644]&~m[1645]&m[1646]&m[1647])|(~m[1641]&m[1644]&~m[1645]&m[1646]&m[1647])|(m[1641]&m[1644]&~m[1645]&m[1646]&m[1647])|(~m[1641]&~m[1644]&m[1645]&m[1646]&m[1647])|(m[1641]&~m[1644]&m[1645]&m[1646]&m[1647])|(m[1641]&m[1644]&m[1645]&m[1646]&m[1647]))):InitCond[430];
    m[1648] = run?((((m[1646]&~m[1649]&~m[1650]&~m[1651]&~m[1652])|(~m[1646]&~m[1649]&~m[1650]&m[1651]&~m[1652])|(m[1646]&m[1649]&~m[1650]&m[1651]&~m[1652])|(m[1646]&~m[1649]&m[1650]&m[1651]&~m[1652])|(~m[1646]&m[1649]&~m[1650]&~m[1651]&m[1652])|(~m[1646]&~m[1649]&m[1650]&~m[1651]&m[1652])|(m[1646]&m[1649]&m[1650]&~m[1651]&m[1652])|(~m[1646]&m[1649]&m[1650]&m[1651]&m[1652]))&UnbiasedRNG[175])|((m[1646]&~m[1649]&~m[1650]&m[1651]&~m[1652])|(~m[1646]&~m[1649]&~m[1650]&~m[1651]&m[1652])|(m[1646]&~m[1649]&~m[1650]&~m[1651]&m[1652])|(m[1646]&m[1649]&~m[1650]&~m[1651]&m[1652])|(m[1646]&~m[1649]&m[1650]&~m[1651]&m[1652])|(~m[1646]&~m[1649]&~m[1650]&m[1651]&m[1652])|(m[1646]&~m[1649]&~m[1650]&m[1651]&m[1652])|(~m[1646]&m[1649]&~m[1650]&m[1651]&m[1652])|(m[1646]&m[1649]&~m[1650]&m[1651]&m[1652])|(~m[1646]&~m[1649]&m[1650]&m[1651]&m[1652])|(m[1646]&~m[1649]&m[1650]&m[1651]&m[1652])|(m[1646]&m[1649]&m[1650]&m[1651]&m[1652]))):InitCond[431];
    m[1653] = run?((((m[1651]&~m[1654]&~m[1655]&~m[1656]&~m[1657])|(~m[1651]&~m[1654]&~m[1655]&m[1656]&~m[1657])|(m[1651]&m[1654]&~m[1655]&m[1656]&~m[1657])|(m[1651]&~m[1654]&m[1655]&m[1656]&~m[1657])|(~m[1651]&m[1654]&~m[1655]&~m[1656]&m[1657])|(~m[1651]&~m[1654]&m[1655]&~m[1656]&m[1657])|(m[1651]&m[1654]&m[1655]&~m[1656]&m[1657])|(~m[1651]&m[1654]&m[1655]&m[1656]&m[1657]))&UnbiasedRNG[176])|((m[1651]&~m[1654]&~m[1655]&m[1656]&~m[1657])|(~m[1651]&~m[1654]&~m[1655]&~m[1656]&m[1657])|(m[1651]&~m[1654]&~m[1655]&~m[1656]&m[1657])|(m[1651]&m[1654]&~m[1655]&~m[1656]&m[1657])|(m[1651]&~m[1654]&m[1655]&~m[1656]&m[1657])|(~m[1651]&~m[1654]&~m[1655]&m[1656]&m[1657])|(m[1651]&~m[1654]&~m[1655]&m[1656]&m[1657])|(~m[1651]&m[1654]&~m[1655]&m[1656]&m[1657])|(m[1651]&m[1654]&~m[1655]&m[1656]&m[1657])|(~m[1651]&~m[1654]&m[1655]&m[1656]&m[1657])|(m[1651]&~m[1654]&m[1655]&m[1656]&m[1657])|(m[1651]&m[1654]&m[1655]&m[1656]&m[1657]))):InitCond[432];
    m[1658] = run?((((m[1656]&~m[1659]&~m[1660]&~m[1661]&~m[1662])|(~m[1656]&~m[1659]&~m[1660]&m[1661]&~m[1662])|(m[1656]&m[1659]&~m[1660]&m[1661]&~m[1662])|(m[1656]&~m[1659]&m[1660]&m[1661]&~m[1662])|(~m[1656]&m[1659]&~m[1660]&~m[1661]&m[1662])|(~m[1656]&~m[1659]&m[1660]&~m[1661]&m[1662])|(m[1656]&m[1659]&m[1660]&~m[1661]&m[1662])|(~m[1656]&m[1659]&m[1660]&m[1661]&m[1662]))&UnbiasedRNG[177])|((m[1656]&~m[1659]&~m[1660]&m[1661]&~m[1662])|(~m[1656]&~m[1659]&~m[1660]&~m[1661]&m[1662])|(m[1656]&~m[1659]&~m[1660]&~m[1661]&m[1662])|(m[1656]&m[1659]&~m[1660]&~m[1661]&m[1662])|(m[1656]&~m[1659]&m[1660]&~m[1661]&m[1662])|(~m[1656]&~m[1659]&~m[1660]&m[1661]&m[1662])|(m[1656]&~m[1659]&~m[1660]&m[1661]&m[1662])|(~m[1656]&m[1659]&~m[1660]&m[1661]&m[1662])|(m[1656]&m[1659]&~m[1660]&m[1661]&m[1662])|(~m[1656]&~m[1659]&m[1660]&m[1661]&m[1662])|(m[1656]&~m[1659]&m[1660]&m[1661]&m[1662])|(m[1656]&m[1659]&m[1660]&m[1661]&m[1662]))):InitCond[433];
    m[1663] = run?((((m[1661]&~m[1664]&~m[1665]&~m[1666]&~m[1667])|(~m[1661]&~m[1664]&~m[1665]&m[1666]&~m[1667])|(m[1661]&m[1664]&~m[1665]&m[1666]&~m[1667])|(m[1661]&~m[1664]&m[1665]&m[1666]&~m[1667])|(~m[1661]&m[1664]&~m[1665]&~m[1666]&m[1667])|(~m[1661]&~m[1664]&m[1665]&~m[1666]&m[1667])|(m[1661]&m[1664]&m[1665]&~m[1666]&m[1667])|(~m[1661]&m[1664]&m[1665]&m[1666]&m[1667]))&UnbiasedRNG[178])|((m[1661]&~m[1664]&~m[1665]&m[1666]&~m[1667])|(~m[1661]&~m[1664]&~m[1665]&~m[1666]&m[1667])|(m[1661]&~m[1664]&~m[1665]&~m[1666]&m[1667])|(m[1661]&m[1664]&~m[1665]&~m[1666]&m[1667])|(m[1661]&~m[1664]&m[1665]&~m[1666]&m[1667])|(~m[1661]&~m[1664]&~m[1665]&m[1666]&m[1667])|(m[1661]&~m[1664]&~m[1665]&m[1666]&m[1667])|(~m[1661]&m[1664]&~m[1665]&m[1666]&m[1667])|(m[1661]&m[1664]&~m[1665]&m[1666]&m[1667])|(~m[1661]&~m[1664]&m[1665]&m[1666]&m[1667])|(m[1661]&~m[1664]&m[1665]&m[1666]&m[1667])|(m[1661]&m[1664]&m[1665]&m[1666]&m[1667]))):InitCond[434];
    m[1668] = run?((((m[1666]&~m[1669]&~m[1670]&~m[1671]&~m[1672])|(~m[1666]&~m[1669]&~m[1670]&m[1671]&~m[1672])|(m[1666]&m[1669]&~m[1670]&m[1671]&~m[1672])|(m[1666]&~m[1669]&m[1670]&m[1671]&~m[1672])|(~m[1666]&m[1669]&~m[1670]&~m[1671]&m[1672])|(~m[1666]&~m[1669]&m[1670]&~m[1671]&m[1672])|(m[1666]&m[1669]&m[1670]&~m[1671]&m[1672])|(~m[1666]&m[1669]&m[1670]&m[1671]&m[1672]))&UnbiasedRNG[179])|((m[1666]&~m[1669]&~m[1670]&m[1671]&~m[1672])|(~m[1666]&~m[1669]&~m[1670]&~m[1671]&m[1672])|(m[1666]&~m[1669]&~m[1670]&~m[1671]&m[1672])|(m[1666]&m[1669]&~m[1670]&~m[1671]&m[1672])|(m[1666]&~m[1669]&m[1670]&~m[1671]&m[1672])|(~m[1666]&~m[1669]&~m[1670]&m[1671]&m[1672])|(m[1666]&~m[1669]&~m[1670]&m[1671]&m[1672])|(~m[1666]&m[1669]&~m[1670]&m[1671]&m[1672])|(m[1666]&m[1669]&~m[1670]&m[1671]&m[1672])|(~m[1666]&~m[1669]&m[1670]&m[1671]&m[1672])|(m[1666]&~m[1669]&m[1670]&m[1671]&m[1672])|(m[1666]&m[1669]&m[1670]&m[1671]&m[1672]))):InitCond[435];
    m[1673] = run?((((m[1607]&~m[1674]&~m[1675]&~m[1676]&~m[1677])|(~m[1607]&~m[1674]&~m[1675]&m[1676]&~m[1677])|(m[1607]&m[1674]&~m[1675]&m[1676]&~m[1677])|(m[1607]&~m[1674]&m[1675]&m[1676]&~m[1677])|(~m[1607]&m[1674]&~m[1675]&~m[1676]&m[1677])|(~m[1607]&~m[1674]&m[1675]&~m[1676]&m[1677])|(m[1607]&m[1674]&m[1675]&~m[1676]&m[1677])|(~m[1607]&m[1674]&m[1675]&m[1676]&m[1677]))&UnbiasedRNG[180])|((m[1607]&~m[1674]&~m[1675]&m[1676]&~m[1677])|(~m[1607]&~m[1674]&~m[1675]&~m[1676]&m[1677])|(m[1607]&~m[1674]&~m[1675]&~m[1676]&m[1677])|(m[1607]&m[1674]&~m[1675]&~m[1676]&m[1677])|(m[1607]&~m[1674]&m[1675]&~m[1676]&m[1677])|(~m[1607]&~m[1674]&~m[1675]&m[1676]&m[1677])|(m[1607]&~m[1674]&~m[1675]&m[1676]&m[1677])|(~m[1607]&m[1674]&~m[1675]&m[1676]&m[1677])|(m[1607]&m[1674]&~m[1675]&m[1676]&m[1677])|(~m[1607]&~m[1674]&m[1675]&m[1676]&m[1677])|(m[1607]&~m[1674]&m[1675]&m[1676]&m[1677])|(m[1607]&m[1674]&m[1675]&m[1676]&m[1677]))):InitCond[436];
    m[1678] = run?((((m[1676]&~m[1679]&~m[1680]&~m[1681]&~m[1682])|(~m[1676]&~m[1679]&~m[1680]&m[1681]&~m[1682])|(m[1676]&m[1679]&~m[1680]&m[1681]&~m[1682])|(m[1676]&~m[1679]&m[1680]&m[1681]&~m[1682])|(~m[1676]&m[1679]&~m[1680]&~m[1681]&m[1682])|(~m[1676]&~m[1679]&m[1680]&~m[1681]&m[1682])|(m[1676]&m[1679]&m[1680]&~m[1681]&m[1682])|(~m[1676]&m[1679]&m[1680]&m[1681]&m[1682]))&UnbiasedRNG[181])|((m[1676]&~m[1679]&~m[1680]&m[1681]&~m[1682])|(~m[1676]&~m[1679]&~m[1680]&~m[1681]&m[1682])|(m[1676]&~m[1679]&~m[1680]&~m[1681]&m[1682])|(m[1676]&m[1679]&~m[1680]&~m[1681]&m[1682])|(m[1676]&~m[1679]&m[1680]&~m[1681]&m[1682])|(~m[1676]&~m[1679]&~m[1680]&m[1681]&m[1682])|(m[1676]&~m[1679]&~m[1680]&m[1681]&m[1682])|(~m[1676]&m[1679]&~m[1680]&m[1681]&m[1682])|(m[1676]&m[1679]&~m[1680]&m[1681]&m[1682])|(~m[1676]&~m[1679]&m[1680]&m[1681]&m[1682])|(m[1676]&~m[1679]&m[1680]&m[1681]&m[1682])|(m[1676]&m[1679]&m[1680]&m[1681]&m[1682]))):InitCond[437];
    m[1683] = run?((((m[1681]&~m[1684]&~m[1685]&~m[1686]&~m[1687])|(~m[1681]&~m[1684]&~m[1685]&m[1686]&~m[1687])|(m[1681]&m[1684]&~m[1685]&m[1686]&~m[1687])|(m[1681]&~m[1684]&m[1685]&m[1686]&~m[1687])|(~m[1681]&m[1684]&~m[1685]&~m[1686]&m[1687])|(~m[1681]&~m[1684]&m[1685]&~m[1686]&m[1687])|(m[1681]&m[1684]&m[1685]&~m[1686]&m[1687])|(~m[1681]&m[1684]&m[1685]&m[1686]&m[1687]))&UnbiasedRNG[182])|((m[1681]&~m[1684]&~m[1685]&m[1686]&~m[1687])|(~m[1681]&~m[1684]&~m[1685]&~m[1686]&m[1687])|(m[1681]&~m[1684]&~m[1685]&~m[1686]&m[1687])|(m[1681]&m[1684]&~m[1685]&~m[1686]&m[1687])|(m[1681]&~m[1684]&m[1685]&~m[1686]&m[1687])|(~m[1681]&~m[1684]&~m[1685]&m[1686]&m[1687])|(m[1681]&~m[1684]&~m[1685]&m[1686]&m[1687])|(~m[1681]&m[1684]&~m[1685]&m[1686]&m[1687])|(m[1681]&m[1684]&~m[1685]&m[1686]&m[1687])|(~m[1681]&~m[1684]&m[1685]&m[1686]&m[1687])|(m[1681]&~m[1684]&m[1685]&m[1686]&m[1687])|(m[1681]&m[1684]&m[1685]&m[1686]&m[1687]))):InitCond[438];
    m[1688] = run?((((m[1686]&~m[1689]&~m[1690]&~m[1691]&~m[1692])|(~m[1686]&~m[1689]&~m[1690]&m[1691]&~m[1692])|(m[1686]&m[1689]&~m[1690]&m[1691]&~m[1692])|(m[1686]&~m[1689]&m[1690]&m[1691]&~m[1692])|(~m[1686]&m[1689]&~m[1690]&~m[1691]&m[1692])|(~m[1686]&~m[1689]&m[1690]&~m[1691]&m[1692])|(m[1686]&m[1689]&m[1690]&~m[1691]&m[1692])|(~m[1686]&m[1689]&m[1690]&m[1691]&m[1692]))&UnbiasedRNG[183])|((m[1686]&~m[1689]&~m[1690]&m[1691]&~m[1692])|(~m[1686]&~m[1689]&~m[1690]&~m[1691]&m[1692])|(m[1686]&~m[1689]&~m[1690]&~m[1691]&m[1692])|(m[1686]&m[1689]&~m[1690]&~m[1691]&m[1692])|(m[1686]&~m[1689]&m[1690]&~m[1691]&m[1692])|(~m[1686]&~m[1689]&~m[1690]&m[1691]&m[1692])|(m[1686]&~m[1689]&~m[1690]&m[1691]&m[1692])|(~m[1686]&m[1689]&~m[1690]&m[1691]&m[1692])|(m[1686]&m[1689]&~m[1690]&m[1691]&m[1692])|(~m[1686]&~m[1689]&m[1690]&m[1691]&m[1692])|(m[1686]&~m[1689]&m[1690]&m[1691]&m[1692])|(m[1686]&m[1689]&m[1690]&m[1691]&m[1692]))):InitCond[439];
    m[1693] = run?((((m[1691]&~m[1694]&~m[1695]&~m[1696]&~m[1697])|(~m[1691]&~m[1694]&~m[1695]&m[1696]&~m[1697])|(m[1691]&m[1694]&~m[1695]&m[1696]&~m[1697])|(m[1691]&~m[1694]&m[1695]&m[1696]&~m[1697])|(~m[1691]&m[1694]&~m[1695]&~m[1696]&m[1697])|(~m[1691]&~m[1694]&m[1695]&~m[1696]&m[1697])|(m[1691]&m[1694]&m[1695]&~m[1696]&m[1697])|(~m[1691]&m[1694]&m[1695]&m[1696]&m[1697]))&UnbiasedRNG[184])|((m[1691]&~m[1694]&~m[1695]&m[1696]&~m[1697])|(~m[1691]&~m[1694]&~m[1695]&~m[1696]&m[1697])|(m[1691]&~m[1694]&~m[1695]&~m[1696]&m[1697])|(m[1691]&m[1694]&~m[1695]&~m[1696]&m[1697])|(m[1691]&~m[1694]&m[1695]&~m[1696]&m[1697])|(~m[1691]&~m[1694]&~m[1695]&m[1696]&m[1697])|(m[1691]&~m[1694]&~m[1695]&m[1696]&m[1697])|(~m[1691]&m[1694]&~m[1695]&m[1696]&m[1697])|(m[1691]&m[1694]&~m[1695]&m[1696]&m[1697])|(~m[1691]&~m[1694]&m[1695]&m[1696]&m[1697])|(m[1691]&~m[1694]&m[1695]&m[1696]&m[1697])|(m[1691]&m[1694]&m[1695]&m[1696]&m[1697]))):InitCond[440];
    m[1698] = run?((((m[1696]&~m[1699]&~m[1700]&~m[1701]&~m[1702])|(~m[1696]&~m[1699]&~m[1700]&m[1701]&~m[1702])|(m[1696]&m[1699]&~m[1700]&m[1701]&~m[1702])|(m[1696]&~m[1699]&m[1700]&m[1701]&~m[1702])|(~m[1696]&m[1699]&~m[1700]&~m[1701]&m[1702])|(~m[1696]&~m[1699]&m[1700]&~m[1701]&m[1702])|(m[1696]&m[1699]&m[1700]&~m[1701]&m[1702])|(~m[1696]&m[1699]&m[1700]&m[1701]&m[1702]))&UnbiasedRNG[185])|((m[1696]&~m[1699]&~m[1700]&m[1701]&~m[1702])|(~m[1696]&~m[1699]&~m[1700]&~m[1701]&m[1702])|(m[1696]&~m[1699]&~m[1700]&~m[1701]&m[1702])|(m[1696]&m[1699]&~m[1700]&~m[1701]&m[1702])|(m[1696]&~m[1699]&m[1700]&~m[1701]&m[1702])|(~m[1696]&~m[1699]&~m[1700]&m[1701]&m[1702])|(m[1696]&~m[1699]&~m[1700]&m[1701]&m[1702])|(~m[1696]&m[1699]&~m[1700]&m[1701]&m[1702])|(m[1696]&m[1699]&~m[1700]&m[1701]&m[1702])|(~m[1696]&~m[1699]&m[1700]&m[1701]&m[1702])|(m[1696]&~m[1699]&m[1700]&m[1701]&m[1702])|(m[1696]&m[1699]&m[1700]&m[1701]&m[1702]))):InitCond[441];
    m[1703] = run?((((m[1701]&~m[1704]&~m[1705]&~m[1706]&~m[1707])|(~m[1701]&~m[1704]&~m[1705]&m[1706]&~m[1707])|(m[1701]&m[1704]&~m[1705]&m[1706]&~m[1707])|(m[1701]&~m[1704]&m[1705]&m[1706]&~m[1707])|(~m[1701]&m[1704]&~m[1705]&~m[1706]&m[1707])|(~m[1701]&~m[1704]&m[1705]&~m[1706]&m[1707])|(m[1701]&m[1704]&m[1705]&~m[1706]&m[1707])|(~m[1701]&m[1704]&m[1705]&m[1706]&m[1707]))&UnbiasedRNG[186])|((m[1701]&~m[1704]&~m[1705]&m[1706]&~m[1707])|(~m[1701]&~m[1704]&~m[1705]&~m[1706]&m[1707])|(m[1701]&~m[1704]&~m[1705]&~m[1706]&m[1707])|(m[1701]&m[1704]&~m[1705]&~m[1706]&m[1707])|(m[1701]&~m[1704]&m[1705]&~m[1706]&m[1707])|(~m[1701]&~m[1704]&~m[1705]&m[1706]&m[1707])|(m[1701]&~m[1704]&~m[1705]&m[1706]&m[1707])|(~m[1701]&m[1704]&~m[1705]&m[1706]&m[1707])|(m[1701]&m[1704]&~m[1705]&m[1706]&m[1707])|(~m[1701]&~m[1704]&m[1705]&m[1706]&m[1707])|(m[1701]&~m[1704]&m[1705]&m[1706]&m[1707])|(m[1701]&m[1704]&m[1705]&m[1706]&m[1707]))):InitCond[442];
    m[1708] = run?((((m[1706]&~m[1709]&~m[1710]&~m[1711]&~m[1712])|(~m[1706]&~m[1709]&~m[1710]&m[1711]&~m[1712])|(m[1706]&m[1709]&~m[1710]&m[1711]&~m[1712])|(m[1706]&~m[1709]&m[1710]&m[1711]&~m[1712])|(~m[1706]&m[1709]&~m[1710]&~m[1711]&m[1712])|(~m[1706]&~m[1709]&m[1710]&~m[1711]&m[1712])|(m[1706]&m[1709]&m[1710]&~m[1711]&m[1712])|(~m[1706]&m[1709]&m[1710]&m[1711]&m[1712]))&UnbiasedRNG[187])|((m[1706]&~m[1709]&~m[1710]&m[1711]&~m[1712])|(~m[1706]&~m[1709]&~m[1710]&~m[1711]&m[1712])|(m[1706]&~m[1709]&~m[1710]&~m[1711]&m[1712])|(m[1706]&m[1709]&~m[1710]&~m[1711]&m[1712])|(m[1706]&~m[1709]&m[1710]&~m[1711]&m[1712])|(~m[1706]&~m[1709]&~m[1710]&m[1711]&m[1712])|(m[1706]&~m[1709]&~m[1710]&m[1711]&m[1712])|(~m[1706]&m[1709]&~m[1710]&m[1711]&m[1712])|(m[1706]&m[1709]&~m[1710]&m[1711]&m[1712])|(~m[1706]&~m[1709]&m[1710]&m[1711]&m[1712])|(m[1706]&~m[1709]&m[1710]&m[1711]&m[1712])|(m[1706]&m[1709]&m[1710]&m[1711]&m[1712]))):InitCond[443];
    m[1713] = run?((((m[1711]&~m[1714]&~m[1715]&~m[1716]&~m[1717])|(~m[1711]&~m[1714]&~m[1715]&m[1716]&~m[1717])|(m[1711]&m[1714]&~m[1715]&m[1716]&~m[1717])|(m[1711]&~m[1714]&m[1715]&m[1716]&~m[1717])|(~m[1711]&m[1714]&~m[1715]&~m[1716]&m[1717])|(~m[1711]&~m[1714]&m[1715]&~m[1716]&m[1717])|(m[1711]&m[1714]&m[1715]&~m[1716]&m[1717])|(~m[1711]&m[1714]&m[1715]&m[1716]&m[1717]))&UnbiasedRNG[188])|((m[1711]&~m[1714]&~m[1715]&m[1716]&~m[1717])|(~m[1711]&~m[1714]&~m[1715]&~m[1716]&m[1717])|(m[1711]&~m[1714]&~m[1715]&~m[1716]&m[1717])|(m[1711]&m[1714]&~m[1715]&~m[1716]&m[1717])|(m[1711]&~m[1714]&m[1715]&~m[1716]&m[1717])|(~m[1711]&~m[1714]&~m[1715]&m[1716]&m[1717])|(m[1711]&~m[1714]&~m[1715]&m[1716]&m[1717])|(~m[1711]&m[1714]&~m[1715]&m[1716]&m[1717])|(m[1711]&m[1714]&~m[1715]&m[1716]&m[1717])|(~m[1711]&~m[1714]&m[1715]&m[1716]&m[1717])|(m[1711]&~m[1714]&m[1715]&m[1716]&m[1717])|(m[1711]&m[1714]&m[1715]&m[1716]&m[1717]))):InitCond[444];
    m[1718] = run?((((m[1716]&~m[1719]&~m[1720]&~m[1721]&~m[1722])|(~m[1716]&~m[1719]&~m[1720]&m[1721]&~m[1722])|(m[1716]&m[1719]&~m[1720]&m[1721]&~m[1722])|(m[1716]&~m[1719]&m[1720]&m[1721]&~m[1722])|(~m[1716]&m[1719]&~m[1720]&~m[1721]&m[1722])|(~m[1716]&~m[1719]&m[1720]&~m[1721]&m[1722])|(m[1716]&m[1719]&m[1720]&~m[1721]&m[1722])|(~m[1716]&m[1719]&m[1720]&m[1721]&m[1722]))&UnbiasedRNG[189])|((m[1716]&~m[1719]&~m[1720]&m[1721]&~m[1722])|(~m[1716]&~m[1719]&~m[1720]&~m[1721]&m[1722])|(m[1716]&~m[1719]&~m[1720]&~m[1721]&m[1722])|(m[1716]&m[1719]&~m[1720]&~m[1721]&m[1722])|(m[1716]&~m[1719]&m[1720]&~m[1721]&m[1722])|(~m[1716]&~m[1719]&~m[1720]&m[1721]&m[1722])|(m[1716]&~m[1719]&~m[1720]&m[1721]&m[1722])|(~m[1716]&m[1719]&~m[1720]&m[1721]&m[1722])|(m[1716]&m[1719]&~m[1720]&m[1721]&m[1722])|(~m[1716]&~m[1719]&m[1720]&m[1721]&m[1722])|(m[1716]&~m[1719]&m[1720]&m[1721]&m[1722])|(m[1716]&m[1719]&m[1720]&m[1721]&m[1722]))):InitCond[445];
    m[1723] = run?((((m[1721]&~m[1724]&~m[1725]&~m[1726]&~m[1727])|(~m[1721]&~m[1724]&~m[1725]&m[1726]&~m[1727])|(m[1721]&m[1724]&~m[1725]&m[1726]&~m[1727])|(m[1721]&~m[1724]&m[1725]&m[1726]&~m[1727])|(~m[1721]&m[1724]&~m[1725]&~m[1726]&m[1727])|(~m[1721]&~m[1724]&m[1725]&~m[1726]&m[1727])|(m[1721]&m[1724]&m[1725]&~m[1726]&m[1727])|(~m[1721]&m[1724]&m[1725]&m[1726]&m[1727]))&UnbiasedRNG[190])|((m[1721]&~m[1724]&~m[1725]&m[1726]&~m[1727])|(~m[1721]&~m[1724]&~m[1725]&~m[1726]&m[1727])|(m[1721]&~m[1724]&~m[1725]&~m[1726]&m[1727])|(m[1721]&m[1724]&~m[1725]&~m[1726]&m[1727])|(m[1721]&~m[1724]&m[1725]&~m[1726]&m[1727])|(~m[1721]&~m[1724]&~m[1725]&m[1726]&m[1727])|(m[1721]&~m[1724]&~m[1725]&m[1726]&m[1727])|(~m[1721]&m[1724]&~m[1725]&m[1726]&m[1727])|(m[1721]&m[1724]&~m[1725]&m[1726]&m[1727])|(~m[1721]&~m[1724]&m[1725]&m[1726]&m[1727])|(m[1721]&~m[1724]&m[1725]&m[1726]&m[1727])|(m[1721]&m[1724]&m[1725]&m[1726]&m[1727]))):InitCond[446];
    m[1728] = run?((((m[1726]&~m[1729]&~m[1730]&~m[1731]&~m[1732])|(~m[1726]&~m[1729]&~m[1730]&m[1731]&~m[1732])|(m[1726]&m[1729]&~m[1730]&m[1731]&~m[1732])|(m[1726]&~m[1729]&m[1730]&m[1731]&~m[1732])|(~m[1726]&m[1729]&~m[1730]&~m[1731]&m[1732])|(~m[1726]&~m[1729]&m[1730]&~m[1731]&m[1732])|(m[1726]&m[1729]&m[1730]&~m[1731]&m[1732])|(~m[1726]&m[1729]&m[1730]&m[1731]&m[1732]))&UnbiasedRNG[191])|((m[1726]&~m[1729]&~m[1730]&m[1731]&~m[1732])|(~m[1726]&~m[1729]&~m[1730]&~m[1731]&m[1732])|(m[1726]&~m[1729]&~m[1730]&~m[1731]&m[1732])|(m[1726]&m[1729]&~m[1730]&~m[1731]&m[1732])|(m[1726]&~m[1729]&m[1730]&~m[1731]&m[1732])|(~m[1726]&~m[1729]&~m[1730]&m[1731]&m[1732])|(m[1726]&~m[1729]&~m[1730]&m[1731]&m[1732])|(~m[1726]&m[1729]&~m[1730]&m[1731]&m[1732])|(m[1726]&m[1729]&~m[1730]&m[1731]&m[1732])|(~m[1726]&~m[1729]&m[1730]&m[1731]&m[1732])|(m[1726]&~m[1729]&m[1730]&m[1731]&m[1732])|(m[1726]&m[1729]&m[1730]&m[1731]&m[1732]))):InitCond[447];
    m[1733] = run?((((m[1731]&~m[1734]&~m[1735]&~m[1736]&~m[1737])|(~m[1731]&~m[1734]&~m[1735]&m[1736]&~m[1737])|(m[1731]&m[1734]&~m[1735]&m[1736]&~m[1737])|(m[1731]&~m[1734]&m[1735]&m[1736]&~m[1737])|(~m[1731]&m[1734]&~m[1735]&~m[1736]&m[1737])|(~m[1731]&~m[1734]&m[1735]&~m[1736]&m[1737])|(m[1731]&m[1734]&m[1735]&~m[1736]&m[1737])|(~m[1731]&m[1734]&m[1735]&m[1736]&m[1737]))&UnbiasedRNG[192])|((m[1731]&~m[1734]&~m[1735]&m[1736]&~m[1737])|(~m[1731]&~m[1734]&~m[1735]&~m[1736]&m[1737])|(m[1731]&~m[1734]&~m[1735]&~m[1736]&m[1737])|(m[1731]&m[1734]&~m[1735]&~m[1736]&m[1737])|(m[1731]&~m[1734]&m[1735]&~m[1736]&m[1737])|(~m[1731]&~m[1734]&~m[1735]&m[1736]&m[1737])|(m[1731]&~m[1734]&~m[1735]&m[1736]&m[1737])|(~m[1731]&m[1734]&~m[1735]&m[1736]&m[1737])|(m[1731]&m[1734]&~m[1735]&m[1736]&m[1737])|(~m[1731]&~m[1734]&m[1735]&m[1736]&m[1737])|(m[1731]&~m[1734]&m[1735]&m[1736]&m[1737])|(m[1731]&m[1734]&m[1735]&m[1736]&m[1737]))):InitCond[448];
    m[1738] = run?((((m[1677]&~m[1739]&~m[1740]&~m[1741]&~m[1742])|(~m[1677]&~m[1739]&~m[1740]&m[1741]&~m[1742])|(m[1677]&m[1739]&~m[1740]&m[1741]&~m[1742])|(m[1677]&~m[1739]&m[1740]&m[1741]&~m[1742])|(~m[1677]&m[1739]&~m[1740]&~m[1741]&m[1742])|(~m[1677]&~m[1739]&m[1740]&~m[1741]&m[1742])|(m[1677]&m[1739]&m[1740]&~m[1741]&m[1742])|(~m[1677]&m[1739]&m[1740]&m[1741]&m[1742]))&UnbiasedRNG[193])|((m[1677]&~m[1739]&~m[1740]&m[1741]&~m[1742])|(~m[1677]&~m[1739]&~m[1740]&~m[1741]&m[1742])|(m[1677]&~m[1739]&~m[1740]&~m[1741]&m[1742])|(m[1677]&m[1739]&~m[1740]&~m[1741]&m[1742])|(m[1677]&~m[1739]&m[1740]&~m[1741]&m[1742])|(~m[1677]&~m[1739]&~m[1740]&m[1741]&m[1742])|(m[1677]&~m[1739]&~m[1740]&m[1741]&m[1742])|(~m[1677]&m[1739]&~m[1740]&m[1741]&m[1742])|(m[1677]&m[1739]&~m[1740]&m[1741]&m[1742])|(~m[1677]&~m[1739]&m[1740]&m[1741]&m[1742])|(m[1677]&~m[1739]&m[1740]&m[1741]&m[1742])|(m[1677]&m[1739]&m[1740]&m[1741]&m[1742]))):InitCond[449];
    m[1743] = run?((((m[1741]&~m[1744]&~m[1745]&~m[1746]&~m[1747])|(~m[1741]&~m[1744]&~m[1745]&m[1746]&~m[1747])|(m[1741]&m[1744]&~m[1745]&m[1746]&~m[1747])|(m[1741]&~m[1744]&m[1745]&m[1746]&~m[1747])|(~m[1741]&m[1744]&~m[1745]&~m[1746]&m[1747])|(~m[1741]&~m[1744]&m[1745]&~m[1746]&m[1747])|(m[1741]&m[1744]&m[1745]&~m[1746]&m[1747])|(~m[1741]&m[1744]&m[1745]&m[1746]&m[1747]))&UnbiasedRNG[194])|((m[1741]&~m[1744]&~m[1745]&m[1746]&~m[1747])|(~m[1741]&~m[1744]&~m[1745]&~m[1746]&m[1747])|(m[1741]&~m[1744]&~m[1745]&~m[1746]&m[1747])|(m[1741]&m[1744]&~m[1745]&~m[1746]&m[1747])|(m[1741]&~m[1744]&m[1745]&~m[1746]&m[1747])|(~m[1741]&~m[1744]&~m[1745]&m[1746]&m[1747])|(m[1741]&~m[1744]&~m[1745]&m[1746]&m[1747])|(~m[1741]&m[1744]&~m[1745]&m[1746]&m[1747])|(m[1741]&m[1744]&~m[1745]&m[1746]&m[1747])|(~m[1741]&~m[1744]&m[1745]&m[1746]&m[1747])|(m[1741]&~m[1744]&m[1745]&m[1746]&m[1747])|(m[1741]&m[1744]&m[1745]&m[1746]&m[1747]))):InitCond[450];
    m[1748] = run?((((m[1746]&~m[1749]&~m[1750]&~m[1751]&~m[1752])|(~m[1746]&~m[1749]&~m[1750]&m[1751]&~m[1752])|(m[1746]&m[1749]&~m[1750]&m[1751]&~m[1752])|(m[1746]&~m[1749]&m[1750]&m[1751]&~m[1752])|(~m[1746]&m[1749]&~m[1750]&~m[1751]&m[1752])|(~m[1746]&~m[1749]&m[1750]&~m[1751]&m[1752])|(m[1746]&m[1749]&m[1750]&~m[1751]&m[1752])|(~m[1746]&m[1749]&m[1750]&m[1751]&m[1752]))&UnbiasedRNG[195])|((m[1746]&~m[1749]&~m[1750]&m[1751]&~m[1752])|(~m[1746]&~m[1749]&~m[1750]&~m[1751]&m[1752])|(m[1746]&~m[1749]&~m[1750]&~m[1751]&m[1752])|(m[1746]&m[1749]&~m[1750]&~m[1751]&m[1752])|(m[1746]&~m[1749]&m[1750]&~m[1751]&m[1752])|(~m[1746]&~m[1749]&~m[1750]&m[1751]&m[1752])|(m[1746]&~m[1749]&~m[1750]&m[1751]&m[1752])|(~m[1746]&m[1749]&~m[1750]&m[1751]&m[1752])|(m[1746]&m[1749]&~m[1750]&m[1751]&m[1752])|(~m[1746]&~m[1749]&m[1750]&m[1751]&m[1752])|(m[1746]&~m[1749]&m[1750]&m[1751]&m[1752])|(m[1746]&m[1749]&m[1750]&m[1751]&m[1752]))):InitCond[451];
    m[1753] = run?((((m[1751]&~m[1754]&~m[1755]&~m[1756]&~m[1757])|(~m[1751]&~m[1754]&~m[1755]&m[1756]&~m[1757])|(m[1751]&m[1754]&~m[1755]&m[1756]&~m[1757])|(m[1751]&~m[1754]&m[1755]&m[1756]&~m[1757])|(~m[1751]&m[1754]&~m[1755]&~m[1756]&m[1757])|(~m[1751]&~m[1754]&m[1755]&~m[1756]&m[1757])|(m[1751]&m[1754]&m[1755]&~m[1756]&m[1757])|(~m[1751]&m[1754]&m[1755]&m[1756]&m[1757]))&UnbiasedRNG[196])|((m[1751]&~m[1754]&~m[1755]&m[1756]&~m[1757])|(~m[1751]&~m[1754]&~m[1755]&~m[1756]&m[1757])|(m[1751]&~m[1754]&~m[1755]&~m[1756]&m[1757])|(m[1751]&m[1754]&~m[1755]&~m[1756]&m[1757])|(m[1751]&~m[1754]&m[1755]&~m[1756]&m[1757])|(~m[1751]&~m[1754]&~m[1755]&m[1756]&m[1757])|(m[1751]&~m[1754]&~m[1755]&m[1756]&m[1757])|(~m[1751]&m[1754]&~m[1755]&m[1756]&m[1757])|(m[1751]&m[1754]&~m[1755]&m[1756]&m[1757])|(~m[1751]&~m[1754]&m[1755]&m[1756]&m[1757])|(m[1751]&~m[1754]&m[1755]&m[1756]&m[1757])|(m[1751]&m[1754]&m[1755]&m[1756]&m[1757]))):InitCond[452];
    m[1758] = run?((((m[1756]&~m[1759]&~m[1760]&~m[1761]&~m[1762])|(~m[1756]&~m[1759]&~m[1760]&m[1761]&~m[1762])|(m[1756]&m[1759]&~m[1760]&m[1761]&~m[1762])|(m[1756]&~m[1759]&m[1760]&m[1761]&~m[1762])|(~m[1756]&m[1759]&~m[1760]&~m[1761]&m[1762])|(~m[1756]&~m[1759]&m[1760]&~m[1761]&m[1762])|(m[1756]&m[1759]&m[1760]&~m[1761]&m[1762])|(~m[1756]&m[1759]&m[1760]&m[1761]&m[1762]))&UnbiasedRNG[197])|((m[1756]&~m[1759]&~m[1760]&m[1761]&~m[1762])|(~m[1756]&~m[1759]&~m[1760]&~m[1761]&m[1762])|(m[1756]&~m[1759]&~m[1760]&~m[1761]&m[1762])|(m[1756]&m[1759]&~m[1760]&~m[1761]&m[1762])|(m[1756]&~m[1759]&m[1760]&~m[1761]&m[1762])|(~m[1756]&~m[1759]&~m[1760]&m[1761]&m[1762])|(m[1756]&~m[1759]&~m[1760]&m[1761]&m[1762])|(~m[1756]&m[1759]&~m[1760]&m[1761]&m[1762])|(m[1756]&m[1759]&~m[1760]&m[1761]&m[1762])|(~m[1756]&~m[1759]&m[1760]&m[1761]&m[1762])|(m[1756]&~m[1759]&m[1760]&m[1761]&m[1762])|(m[1756]&m[1759]&m[1760]&m[1761]&m[1762]))):InitCond[453];
    m[1763] = run?((((m[1761]&~m[1764]&~m[1765]&~m[1766]&~m[1767])|(~m[1761]&~m[1764]&~m[1765]&m[1766]&~m[1767])|(m[1761]&m[1764]&~m[1765]&m[1766]&~m[1767])|(m[1761]&~m[1764]&m[1765]&m[1766]&~m[1767])|(~m[1761]&m[1764]&~m[1765]&~m[1766]&m[1767])|(~m[1761]&~m[1764]&m[1765]&~m[1766]&m[1767])|(m[1761]&m[1764]&m[1765]&~m[1766]&m[1767])|(~m[1761]&m[1764]&m[1765]&m[1766]&m[1767]))&UnbiasedRNG[198])|((m[1761]&~m[1764]&~m[1765]&m[1766]&~m[1767])|(~m[1761]&~m[1764]&~m[1765]&~m[1766]&m[1767])|(m[1761]&~m[1764]&~m[1765]&~m[1766]&m[1767])|(m[1761]&m[1764]&~m[1765]&~m[1766]&m[1767])|(m[1761]&~m[1764]&m[1765]&~m[1766]&m[1767])|(~m[1761]&~m[1764]&~m[1765]&m[1766]&m[1767])|(m[1761]&~m[1764]&~m[1765]&m[1766]&m[1767])|(~m[1761]&m[1764]&~m[1765]&m[1766]&m[1767])|(m[1761]&m[1764]&~m[1765]&m[1766]&m[1767])|(~m[1761]&~m[1764]&m[1765]&m[1766]&m[1767])|(m[1761]&~m[1764]&m[1765]&m[1766]&m[1767])|(m[1761]&m[1764]&m[1765]&m[1766]&m[1767]))):InitCond[454];
    m[1768] = run?((((m[1766]&~m[1769]&~m[1770]&~m[1771]&~m[1772])|(~m[1766]&~m[1769]&~m[1770]&m[1771]&~m[1772])|(m[1766]&m[1769]&~m[1770]&m[1771]&~m[1772])|(m[1766]&~m[1769]&m[1770]&m[1771]&~m[1772])|(~m[1766]&m[1769]&~m[1770]&~m[1771]&m[1772])|(~m[1766]&~m[1769]&m[1770]&~m[1771]&m[1772])|(m[1766]&m[1769]&m[1770]&~m[1771]&m[1772])|(~m[1766]&m[1769]&m[1770]&m[1771]&m[1772]))&UnbiasedRNG[199])|((m[1766]&~m[1769]&~m[1770]&m[1771]&~m[1772])|(~m[1766]&~m[1769]&~m[1770]&~m[1771]&m[1772])|(m[1766]&~m[1769]&~m[1770]&~m[1771]&m[1772])|(m[1766]&m[1769]&~m[1770]&~m[1771]&m[1772])|(m[1766]&~m[1769]&m[1770]&~m[1771]&m[1772])|(~m[1766]&~m[1769]&~m[1770]&m[1771]&m[1772])|(m[1766]&~m[1769]&~m[1770]&m[1771]&m[1772])|(~m[1766]&m[1769]&~m[1770]&m[1771]&m[1772])|(m[1766]&m[1769]&~m[1770]&m[1771]&m[1772])|(~m[1766]&~m[1769]&m[1770]&m[1771]&m[1772])|(m[1766]&~m[1769]&m[1770]&m[1771]&m[1772])|(m[1766]&m[1769]&m[1770]&m[1771]&m[1772]))):InitCond[455];
    m[1773] = run?((((m[1771]&~m[1774]&~m[1775]&~m[1776]&~m[1777])|(~m[1771]&~m[1774]&~m[1775]&m[1776]&~m[1777])|(m[1771]&m[1774]&~m[1775]&m[1776]&~m[1777])|(m[1771]&~m[1774]&m[1775]&m[1776]&~m[1777])|(~m[1771]&m[1774]&~m[1775]&~m[1776]&m[1777])|(~m[1771]&~m[1774]&m[1775]&~m[1776]&m[1777])|(m[1771]&m[1774]&m[1775]&~m[1776]&m[1777])|(~m[1771]&m[1774]&m[1775]&m[1776]&m[1777]))&UnbiasedRNG[200])|((m[1771]&~m[1774]&~m[1775]&m[1776]&~m[1777])|(~m[1771]&~m[1774]&~m[1775]&~m[1776]&m[1777])|(m[1771]&~m[1774]&~m[1775]&~m[1776]&m[1777])|(m[1771]&m[1774]&~m[1775]&~m[1776]&m[1777])|(m[1771]&~m[1774]&m[1775]&~m[1776]&m[1777])|(~m[1771]&~m[1774]&~m[1775]&m[1776]&m[1777])|(m[1771]&~m[1774]&~m[1775]&m[1776]&m[1777])|(~m[1771]&m[1774]&~m[1775]&m[1776]&m[1777])|(m[1771]&m[1774]&~m[1775]&m[1776]&m[1777])|(~m[1771]&~m[1774]&m[1775]&m[1776]&m[1777])|(m[1771]&~m[1774]&m[1775]&m[1776]&m[1777])|(m[1771]&m[1774]&m[1775]&m[1776]&m[1777]))):InitCond[456];
    m[1778] = run?((((m[1776]&~m[1779]&~m[1780]&~m[1781]&~m[1782])|(~m[1776]&~m[1779]&~m[1780]&m[1781]&~m[1782])|(m[1776]&m[1779]&~m[1780]&m[1781]&~m[1782])|(m[1776]&~m[1779]&m[1780]&m[1781]&~m[1782])|(~m[1776]&m[1779]&~m[1780]&~m[1781]&m[1782])|(~m[1776]&~m[1779]&m[1780]&~m[1781]&m[1782])|(m[1776]&m[1779]&m[1780]&~m[1781]&m[1782])|(~m[1776]&m[1779]&m[1780]&m[1781]&m[1782]))&UnbiasedRNG[201])|((m[1776]&~m[1779]&~m[1780]&m[1781]&~m[1782])|(~m[1776]&~m[1779]&~m[1780]&~m[1781]&m[1782])|(m[1776]&~m[1779]&~m[1780]&~m[1781]&m[1782])|(m[1776]&m[1779]&~m[1780]&~m[1781]&m[1782])|(m[1776]&~m[1779]&m[1780]&~m[1781]&m[1782])|(~m[1776]&~m[1779]&~m[1780]&m[1781]&m[1782])|(m[1776]&~m[1779]&~m[1780]&m[1781]&m[1782])|(~m[1776]&m[1779]&~m[1780]&m[1781]&m[1782])|(m[1776]&m[1779]&~m[1780]&m[1781]&m[1782])|(~m[1776]&~m[1779]&m[1780]&m[1781]&m[1782])|(m[1776]&~m[1779]&m[1780]&m[1781]&m[1782])|(m[1776]&m[1779]&m[1780]&m[1781]&m[1782]))):InitCond[457];
    m[1783] = run?((((m[1781]&~m[1784]&~m[1785]&~m[1786]&~m[1787])|(~m[1781]&~m[1784]&~m[1785]&m[1786]&~m[1787])|(m[1781]&m[1784]&~m[1785]&m[1786]&~m[1787])|(m[1781]&~m[1784]&m[1785]&m[1786]&~m[1787])|(~m[1781]&m[1784]&~m[1785]&~m[1786]&m[1787])|(~m[1781]&~m[1784]&m[1785]&~m[1786]&m[1787])|(m[1781]&m[1784]&m[1785]&~m[1786]&m[1787])|(~m[1781]&m[1784]&m[1785]&m[1786]&m[1787]))&UnbiasedRNG[202])|((m[1781]&~m[1784]&~m[1785]&m[1786]&~m[1787])|(~m[1781]&~m[1784]&~m[1785]&~m[1786]&m[1787])|(m[1781]&~m[1784]&~m[1785]&~m[1786]&m[1787])|(m[1781]&m[1784]&~m[1785]&~m[1786]&m[1787])|(m[1781]&~m[1784]&m[1785]&~m[1786]&m[1787])|(~m[1781]&~m[1784]&~m[1785]&m[1786]&m[1787])|(m[1781]&~m[1784]&~m[1785]&m[1786]&m[1787])|(~m[1781]&m[1784]&~m[1785]&m[1786]&m[1787])|(m[1781]&m[1784]&~m[1785]&m[1786]&m[1787])|(~m[1781]&~m[1784]&m[1785]&m[1786]&m[1787])|(m[1781]&~m[1784]&m[1785]&m[1786]&m[1787])|(m[1781]&m[1784]&m[1785]&m[1786]&m[1787]))):InitCond[458];
    m[1788] = run?((((m[1786]&~m[1789]&~m[1790]&~m[1791]&~m[1792])|(~m[1786]&~m[1789]&~m[1790]&m[1791]&~m[1792])|(m[1786]&m[1789]&~m[1790]&m[1791]&~m[1792])|(m[1786]&~m[1789]&m[1790]&m[1791]&~m[1792])|(~m[1786]&m[1789]&~m[1790]&~m[1791]&m[1792])|(~m[1786]&~m[1789]&m[1790]&~m[1791]&m[1792])|(m[1786]&m[1789]&m[1790]&~m[1791]&m[1792])|(~m[1786]&m[1789]&m[1790]&m[1791]&m[1792]))&UnbiasedRNG[203])|((m[1786]&~m[1789]&~m[1790]&m[1791]&~m[1792])|(~m[1786]&~m[1789]&~m[1790]&~m[1791]&m[1792])|(m[1786]&~m[1789]&~m[1790]&~m[1791]&m[1792])|(m[1786]&m[1789]&~m[1790]&~m[1791]&m[1792])|(m[1786]&~m[1789]&m[1790]&~m[1791]&m[1792])|(~m[1786]&~m[1789]&~m[1790]&m[1791]&m[1792])|(m[1786]&~m[1789]&~m[1790]&m[1791]&m[1792])|(~m[1786]&m[1789]&~m[1790]&m[1791]&m[1792])|(m[1786]&m[1789]&~m[1790]&m[1791]&m[1792])|(~m[1786]&~m[1789]&m[1790]&m[1791]&m[1792])|(m[1786]&~m[1789]&m[1790]&m[1791]&m[1792])|(m[1786]&m[1789]&m[1790]&m[1791]&m[1792]))):InitCond[459];
    m[1793] = run?((((m[1791]&~m[1794]&~m[1795]&~m[1796]&~m[1797])|(~m[1791]&~m[1794]&~m[1795]&m[1796]&~m[1797])|(m[1791]&m[1794]&~m[1795]&m[1796]&~m[1797])|(m[1791]&~m[1794]&m[1795]&m[1796]&~m[1797])|(~m[1791]&m[1794]&~m[1795]&~m[1796]&m[1797])|(~m[1791]&~m[1794]&m[1795]&~m[1796]&m[1797])|(m[1791]&m[1794]&m[1795]&~m[1796]&m[1797])|(~m[1791]&m[1794]&m[1795]&m[1796]&m[1797]))&UnbiasedRNG[204])|((m[1791]&~m[1794]&~m[1795]&m[1796]&~m[1797])|(~m[1791]&~m[1794]&~m[1795]&~m[1796]&m[1797])|(m[1791]&~m[1794]&~m[1795]&~m[1796]&m[1797])|(m[1791]&m[1794]&~m[1795]&~m[1796]&m[1797])|(m[1791]&~m[1794]&m[1795]&~m[1796]&m[1797])|(~m[1791]&~m[1794]&~m[1795]&m[1796]&m[1797])|(m[1791]&~m[1794]&~m[1795]&m[1796]&m[1797])|(~m[1791]&m[1794]&~m[1795]&m[1796]&m[1797])|(m[1791]&m[1794]&~m[1795]&m[1796]&m[1797])|(~m[1791]&~m[1794]&m[1795]&m[1796]&m[1797])|(m[1791]&~m[1794]&m[1795]&m[1796]&m[1797])|(m[1791]&m[1794]&m[1795]&m[1796]&m[1797]))):InitCond[460];
    m[1798] = run?((((m[1742]&~m[1799]&~m[1800]&~m[1801]&~m[1802])|(~m[1742]&~m[1799]&~m[1800]&m[1801]&~m[1802])|(m[1742]&m[1799]&~m[1800]&m[1801]&~m[1802])|(m[1742]&~m[1799]&m[1800]&m[1801]&~m[1802])|(~m[1742]&m[1799]&~m[1800]&~m[1801]&m[1802])|(~m[1742]&~m[1799]&m[1800]&~m[1801]&m[1802])|(m[1742]&m[1799]&m[1800]&~m[1801]&m[1802])|(~m[1742]&m[1799]&m[1800]&m[1801]&m[1802]))&UnbiasedRNG[205])|((m[1742]&~m[1799]&~m[1800]&m[1801]&~m[1802])|(~m[1742]&~m[1799]&~m[1800]&~m[1801]&m[1802])|(m[1742]&~m[1799]&~m[1800]&~m[1801]&m[1802])|(m[1742]&m[1799]&~m[1800]&~m[1801]&m[1802])|(m[1742]&~m[1799]&m[1800]&~m[1801]&m[1802])|(~m[1742]&~m[1799]&~m[1800]&m[1801]&m[1802])|(m[1742]&~m[1799]&~m[1800]&m[1801]&m[1802])|(~m[1742]&m[1799]&~m[1800]&m[1801]&m[1802])|(m[1742]&m[1799]&~m[1800]&m[1801]&m[1802])|(~m[1742]&~m[1799]&m[1800]&m[1801]&m[1802])|(m[1742]&~m[1799]&m[1800]&m[1801]&m[1802])|(m[1742]&m[1799]&m[1800]&m[1801]&m[1802]))):InitCond[461];
    m[1803] = run?((((m[1801]&~m[1804]&~m[1805]&~m[1806]&~m[1807])|(~m[1801]&~m[1804]&~m[1805]&m[1806]&~m[1807])|(m[1801]&m[1804]&~m[1805]&m[1806]&~m[1807])|(m[1801]&~m[1804]&m[1805]&m[1806]&~m[1807])|(~m[1801]&m[1804]&~m[1805]&~m[1806]&m[1807])|(~m[1801]&~m[1804]&m[1805]&~m[1806]&m[1807])|(m[1801]&m[1804]&m[1805]&~m[1806]&m[1807])|(~m[1801]&m[1804]&m[1805]&m[1806]&m[1807]))&UnbiasedRNG[206])|((m[1801]&~m[1804]&~m[1805]&m[1806]&~m[1807])|(~m[1801]&~m[1804]&~m[1805]&~m[1806]&m[1807])|(m[1801]&~m[1804]&~m[1805]&~m[1806]&m[1807])|(m[1801]&m[1804]&~m[1805]&~m[1806]&m[1807])|(m[1801]&~m[1804]&m[1805]&~m[1806]&m[1807])|(~m[1801]&~m[1804]&~m[1805]&m[1806]&m[1807])|(m[1801]&~m[1804]&~m[1805]&m[1806]&m[1807])|(~m[1801]&m[1804]&~m[1805]&m[1806]&m[1807])|(m[1801]&m[1804]&~m[1805]&m[1806]&m[1807])|(~m[1801]&~m[1804]&m[1805]&m[1806]&m[1807])|(m[1801]&~m[1804]&m[1805]&m[1806]&m[1807])|(m[1801]&m[1804]&m[1805]&m[1806]&m[1807]))):InitCond[462];
    m[1808] = run?((((m[1806]&~m[1809]&~m[1810]&~m[1811]&~m[1812])|(~m[1806]&~m[1809]&~m[1810]&m[1811]&~m[1812])|(m[1806]&m[1809]&~m[1810]&m[1811]&~m[1812])|(m[1806]&~m[1809]&m[1810]&m[1811]&~m[1812])|(~m[1806]&m[1809]&~m[1810]&~m[1811]&m[1812])|(~m[1806]&~m[1809]&m[1810]&~m[1811]&m[1812])|(m[1806]&m[1809]&m[1810]&~m[1811]&m[1812])|(~m[1806]&m[1809]&m[1810]&m[1811]&m[1812]))&UnbiasedRNG[207])|((m[1806]&~m[1809]&~m[1810]&m[1811]&~m[1812])|(~m[1806]&~m[1809]&~m[1810]&~m[1811]&m[1812])|(m[1806]&~m[1809]&~m[1810]&~m[1811]&m[1812])|(m[1806]&m[1809]&~m[1810]&~m[1811]&m[1812])|(m[1806]&~m[1809]&m[1810]&~m[1811]&m[1812])|(~m[1806]&~m[1809]&~m[1810]&m[1811]&m[1812])|(m[1806]&~m[1809]&~m[1810]&m[1811]&m[1812])|(~m[1806]&m[1809]&~m[1810]&m[1811]&m[1812])|(m[1806]&m[1809]&~m[1810]&m[1811]&m[1812])|(~m[1806]&~m[1809]&m[1810]&m[1811]&m[1812])|(m[1806]&~m[1809]&m[1810]&m[1811]&m[1812])|(m[1806]&m[1809]&m[1810]&m[1811]&m[1812]))):InitCond[463];
    m[1813] = run?((((m[1811]&~m[1814]&~m[1815]&~m[1816]&~m[1817])|(~m[1811]&~m[1814]&~m[1815]&m[1816]&~m[1817])|(m[1811]&m[1814]&~m[1815]&m[1816]&~m[1817])|(m[1811]&~m[1814]&m[1815]&m[1816]&~m[1817])|(~m[1811]&m[1814]&~m[1815]&~m[1816]&m[1817])|(~m[1811]&~m[1814]&m[1815]&~m[1816]&m[1817])|(m[1811]&m[1814]&m[1815]&~m[1816]&m[1817])|(~m[1811]&m[1814]&m[1815]&m[1816]&m[1817]))&UnbiasedRNG[208])|((m[1811]&~m[1814]&~m[1815]&m[1816]&~m[1817])|(~m[1811]&~m[1814]&~m[1815]&~m[1816]&m[1817])|(m[1811]&~m[1814]&~m[1815]&~m[1816]&m[1817])|(m[1811]&m[1814]&~m[1815]&~m[1816]&m[1817])|(m[1811]&~m[1814]&m[1815]&~m[1816]&m[1817])|(~m[1811]&~m[1814]&~m[1815]&m[1816]&m[1817])|(m[1811]&~m[1814]&~m[1815]&m[1816]&m[1817])|(~m[1811]&m[1814]&~m[1815]&m[1816]&m[1817])|(m[1811]&m[1814]&~m[1815]&m[1816]&m[1817])|(~m[1811]&~m[1814]&m[1815]&m[1816]&m[1817])|(m[1811]&~m[1814]&m[1815]&m[1816]&m[1817])|(m[1811]&m[1814]&m[1815]&m[1816]&m[1817]))):InitCond[464];
    m[1818] = run?((((m[1816]&~m[1819]&~m[1820]&~m[1821]&~m[1822])|(~m[1816]&~m[1819]&~m[1820]&m[1821]&~m[1822])|(m[1816]&m[1819]&~m[1820]&m[1821]&~m[1822])|(m[1816]&~m[1819]&m[1820]&m[1821]&~m[1822])|(~m[1816]&m[1819]&~m[1820]&~m[1821]&m[1822])|(~m[1816]&~m[1819]&m[1820]&~m[1821]&m[1822])|(m[1816]&m[1819]&m[1820]&~m[1821]&m[1822])|(~m[1816]&m[1819]&m[1820]&m[1821]&m[1822]))&UnbiasedRNG[209])|((m[1816]&~m[1819]&~m[1820]&m[1821]&~m[1822])|(~m[1816]&~m[1819]&~m[1820]&~m[1821]&m[1822])|(m[1816]&~m[1819]&~m[1820]&~m[1821]&m[1822])|(m[1816]&m[1819]&~m[1820]&~m[1821]&m[1822])|(m[1816]&~m[1819]&m[1820]&~m[1821]&m[1822])|(~m[1816]&~m[1819]&~m[1820]&m[1821]&m[1822])|(m[1816]&~m[1819]&~m[1820]&m[1821]&m[1822])|(~m[1816]&m[1819]&~m[1820]&m[1821]&m[1822])|(m[1816]&m[1819]&~m[1820]&m[1821]&m[1822])|(~m[1816]&~m[1819]&m[1820]&m[1821]&m[1822])|(m[1816]&~m[1819]&m[1820]&m[1821]&m[1822])|(m[1816]&m[1819]&m[1820]&m[1821]&m[1822]))):InitCond[465];
    m[1823] = run?((((m[1821]&~m[1824]&~m[1825]&~m[1826]&~m[1827])|(~m[1821]&~m[1824]&~m[1825]&m[1826]&~m[1827])|(m[1821]&m[1824]&~m[1825]&m[1826]&~m[1827])|(m[1821]&~m[1824]&m[1825]&m[1826]&~m[1827])|(~m[1821]&m[1824]&~m[1825]&~m[1826]&m[1827])|(~m[1821]&~m[1824]&m[1825]&~m[1826]&m[1827])|(m[1821]&m[1824]&m[1825]&~m[1826]&m[1827])|(~m[1821]&m[1824]&m[1825]&m[1826]&m[1827]))&UnbiasedRNG[210])|((m[1821]&~m[1824]&~m[1825]&m[1826]&~m[1827])|(~m[1821]&~m[1824]&~m[1825]&~m[1826]&m[1827])|(m[1821]&~m[1824]&~m[1825]&~m[1826]&m[1827])|(m[1821]&m[1824]&~m[1825]&~m[1826]&m[1827])|(m[1821]&~m[1824]&m[1825]&~m[1826]&m[1827])|(~m[1821]&~m[1824]&~m[1825]&m[1826]&m[1827])|(m[1821]&~m[1824]&~m[1825]&m[1826]&m[1827])|(~m[1821]&m[1824]&~m[1825]&m[1826]&m[1827])|(m[1821]&m[1824]&~m[1825]&m[1826]&m[1827])|(~m[1821]&~m[1824]&m[1825]&m[1826]&m[1827])|(m[1821]&~m[1824]&m[1825]&m[1826]&m[1827])|(m[1821]&m[1824]&m[1825]&m[1826]&m[1827]))):InitCond[466];
    m[1828] = run?((((m[1826]&~m[1829]&~m[1830]&~m[1831]&~m[1832])|(~m[1826]&~m[1829]&~m[1830]&m[1831]&~m[1832])|(m[1826]&m[1829]&~m[1830]&m[1831]&~m[1832])|(m[1826]&~m[1829]&m[1830]&m[1831]&~m[1832])|(~m[1826]&m[1829]&~m[1830]&~m[1831]&m[1832])|(~m[1826]&~m[1829]&m[1830]&~m[1831]&m[1832])|(m[1826]&m[1829]&m[1830]&~m[1831]&m[1832])|(~m[1826]&m[1829]&m[1830]&m[1831]&m[1832]))&UnbiasedRNG[211])|((m[1826]&~m[1829]&~m[1830]&m[1831]&~m[1832])|(~m[1826]&~m[1829]&~m[1830]&~m[1831]&m[1832])|(m[1826]&~m[1829]&~m[1830]&~m[1831]&m[1832])|(m[1826]&m[1829]&~m[1830]&~m[1831]&m[1832])|(m[1826]&~m[1829]&m[1830]&~m[1831]&m[1832])|(~m[1826]&~m[1829]&~m[1830]&m[1831]&m[1832])|(m[1826]&~m[1829]&~m[1830]&m[1831]&m[1832])|(~m[1826]&m[1829]&~m[1830]&m[1831]&m[1832])|(m[1826]&m[1829]&~m[1830]&m[1831]&m[1832])|(~m[1826]&~m[1829]&m[1830]&m[1831]&m[1832])|(m[1826]&~m[1829]&m[1830]&m[1831]&m[1832])|(m[1826]&m[1829]&m[1830]&m[1831]&m[1832]))):InitCond[467];
    m[1833] = run?((((m[1831]&~m[1834]&~m[1835]&~m[1836]&~m[1837])|(~m[1831]&~m[1834]&~m[1835]&m[1836]&~m[1837])|(m[1831]&m[1834]&~m[1835]&m[1836]&~m[1837])|(m[1831]&~m[1834]&m[1835]&m[1836]&~m[1837])|(~m[1831]&m[1834]&~m[1835]&~m[1836]&m[1837])|(~m[1831]&~m[1834]&m[1835]&~m[1836]&m[1837])|(m[1831]&m[1834]&m[1835]&~m[1836]&m[1837])|(~m[1831]&m[1834]&m[1835]&m[1836]&m[1837]))&UnbiasedRNG[212])|((m[1831]&~m[1834]&~m[1835]&m[1836]&~m[1837])|(~m[1831]&~m[1834]&~m[1835]&~m[1836]&m[1837])|(m[1831]&~m[1834]&~m[1835]&~m[1836]&m[1837])|(m[1831]&m[1834]&~m[1835]&~m[1836]&m[1837])|(m[1831]&~m[1834]&m[1835]&~m[1836]&m[1837])|(~m[1831]&~m[1834]&~m[1835]&m[1836]&m[1837])|(m[1831]&~m[1834]&~m[1835]&m[1836]&m[1837])|(~m[1831]&m[1834]&~m[1835]&m[1836]&m[1837])|(m[1831]&m[1834]&~m[1835]&m[1836]&m[1837])|(~m[1831]&~m[1834]&m[1835]&m[1836]&m[1837])|(m[1831]&~m[1834]&m[1835]&m[1836]&m[1837])|(m[1831]&m[1834]&m[1835]&m[1836]&m[1837]))):InitCond[468];
    m[1838] = run?((((m[1836]&~m[1839]&~m[1840]&~m[1841]&~m[1842])|(~m[1836]&~m[1839]&~m[1840]&m[1841]&~m[1842])|(m[1836]&m[1839]&~m[1840]&m[1841]&~m[1842])|(m[1836]&~m[1839]&m[1840]&m[1841]&~m[1842])|(~m[1836]&m[1839]&~m[1840]&~m[1841]&m[1842])|(~m[1836]&~m[1839]&m[1840]&~m[1841]&m[1842])|(m[1836]&m[1839]&m[1840]&~m[1841]&m[1842])|(~m[1836]&m[1839]&m[1840]&m[1841]&m[1842]))&UnbiasedRNG[213])|((m[1836]&~m[1839]&~m[1840]&m[1841]&~m[1842])|(~m[1836]&~m[1839]&~m[1840]&~m[1841]&m[1842])|(m[1836]&~m[1839]&~m[1840]&~m[1841]&m[1842])|(m[1836]&m[1839]&~m[1840]&~m[1841]&m[1842])|(m[1836]&~m[1839]&m[1840]&~m[1841]&m[1842])|(~m[1836]&~m[1839]&~m[1840]&m[1841]&m[1842])|(m[1836]&~m[1839]&~m[1840]&m[1841]&m[1842])|(~m[1836]&m[1839]&~m[1840]&m[1841]&m[1842])|(m[1836]&m[1839]&~m[1840]&m[1841]&m[1842])|(~m[1836]&~m[1839]&m[1840]&m[1841]&m[1842])|(m[1836]&~m[1839]&m[1840]&m[1841]&m[1842])|(m[1836]&m[1839]&m[1840]&m[1841]&m[1842]))):InitCond[469];
    m[1843] = run?((((m[1841]&~m[1844]&~m[1845]&~m[1846]&~m[1847])|(~m[1841]&~m[1844]&~m[1845]&m[1846]&~m[1847])|(m[1841]&m[1844]&~m[1845]&m[1846]&~m[1847])|(m[1841]&~m[1844]&m[1845]&m[1846]&~m[1847])|(~m[1841]&m[1844]&~m[1845]&~m[1846]&m[1847])|(~m[1841]&~m[1844]&m[1845]&~m[1846]&m[1847])|(m[1841]&m[1844]&m[1845]&~m[1846]&m[1847])|(~m[1841]&m[1844]&m[1845]&m[1846]&m[1847]))&UnbiasedRNG[214])|((m[1841]&~m[1844]&~m[1845]&m[1846]&~m[1847])|(~m[1841]&~m[1844]&~m[1845]&~m[1846]&m[1847])|(m[1841]&~m[1844]&~m[1845]&~m[1846]&m[1847])|(m[1841]&m[1844]&~m[1845]&~m[1846]&m[1847])|(m[1841]&~m[1844]&m[1845]&~m[1846]&m[1847])|(~m[1841]&~m[1844]&~m[1845]&m[1846]&m[1847])|(m[1841]&~m[1844]&~m[1845]&m[1846]&m[1847])|(~m[1841]&m[1844]&~m[1845]&m[1846]&m[1847])|(m[1841]&m[1844]&~m[1845]&m[1846]&m[1847])|(~m[1841]&~m[1844]&m[1845]&m[1846]&m[1847])|(m[1841]&~m[1844]&m[1845]&m[1846]&m[1847])|(m[1841]&m[1844]&m[1845]&m[1846]&m[1847]))):InitCond[470];
    m[1848] = run?((((m[1846]&~m[1849]&~m[1850]&~m[1851]&~m[1852])|(~m[1846]&~m[1849]&~m[1850]&m[1851]&~m[1852])|(m[1846]&m[1849]&~m[1850]&m[1851]&~m[1852])|(m[1846]&~m[1849]&m[1850]&m[1851]&~m[1852])|(~m[1846]&m[1849]&~m[1850]&~m[1851]&m[1852])|(~m[1846]&~m[1849]&m[1850]&~m[1851]&m[1852])|(m[1846]&m[1849]&m[1850]&~m[1851]&m[1852])|(~m[1846]&m[1849]&m[1850]&m[1851]&m[1852]))&UnbiasedRNG[215])|((m[1846]&~m[1849]&~m[1850]&m[1851]&~m[1852])|(~m[1846]&~m[1849]&~m[1850]&~m[1851]&m[1852])|(m[1846]&~m[1849]&~m[1850]&~m[1851]&m[1852])|(m[1846]&m[1849]&~m[1850]&~m[1851]&m[1852])|(m[1846]&~m[1849]&m[1850]&~m[1851]&m[1852])|(~m[1846]&~m[1849]&~m[1850]&m[1851]&m[1852])|(m[1846]&~m[1849]&~m[1850]&m[1851]&m[1852])|(~m[1846]&m[1849]&~m[1850]&m[1851]&m[1852])|(m[1846]&m[1849]&~m[1850]&m[1851]&m[1852])|(~m[1846]&~m[1849]&m[1850]&m[1851]&m[1852])|(m[1846]&~m[1849]&m[1850]&m[1851]&m[1852])|(m[1846]&m[1849]&m[1850]&m[1851]&m[1852]))):InitCond[471];
    m[1853] = run?((((m[1802]&~m[1854]&~m[1855]&~m[1856]&~m[1857])|(~m[1802]&~m[1854]&~m[1855]&m[1856]&~m[1857])|(m[1802]&m[1854]&~m[1855]&m[1856]&~m[1857])|(m[1802]&~m[1854]&m[1855]&m[1856]&~m[1857])|(~m[1802]&m[1854]&~m[1855]&~m[1856]&m[1857])|(~m[1802]&~m[1854]&m[1855]&~m[1856]&m[1857])|(m[1802]&m[1854]&m[1855]&~m[1856]&m[1857])|(~m[1802]&m[1854]&m[1855]&m[1856]&m[1857]))&UnbiasedRNG[216])|((m[1802]&~m[1854]&~m[1855]&m[1856]&~m[1857])|(~m[1802]&~m[1854]&~m[1855]&~m[1856]&m[1857])|(m[1802]&~m[1854]&~m[1855]&~m[1856]&m[1857])|(m[1802]&m[1854]&~m[1855]&~m[1856]&m[1857])|(m[1802]&~m[1854]&m[1855]&~m[1856]&m[1857])|(~m[1802]&~m[1854]&~m[1855]&m[1856]&m[1857])|(m[1802]&~m[1854]&~m[1855]&m[1856]&m[1857])|(~m[1802]&m[1854]&~m[1855]&m[1856]&m[1857])|(m[1802]&m[1854]&~m[1855]&m[1856]&m[1857])|(~m[1802]&~m[1854]&m[1855]&m[1856]&m[1857])|(m[1802]&~m[1854]&m[1855]&m[1856]&m[1857])|(m[1802]&m[1854]&m[1855]&m[1856]&m[1857]))):InitCond[472];
    m[1858] = run?((((m[1856]&~m[1859]&~m[1860]&~m[1861]&~m[1862])|(~m[1856]&~m[1859]&~m[1860]&m[1861]&~m[1862])|(m[1856]&m[1859]&~m[1860]&m[1861]&~m[1862])|(m[1856]&~m[1859]&m[1860]&m[1861]&~m[1862])|(~m[1856]&m[1859]&~m[1860]&~m[1861]&m[1862])|(~m[1856]&~m[1859]&m[1860]&~m[1861]&m[1862])|(m[1856]&m[1859]&m[1860]&~m[1861]&m[1862])|(~m[1856]&m[1859]&m[1860]&m[1861]&m[1862]))&UnbiasedRNG[217])|((m[1856]&~m[1859]&~m[1860]&m[1861]&~m[1862])|(~m[1856]&~m[1859]&~m[1860]&~m[1861]&m[1862])|(m[1856]&~m[1859]&~m[1860]&~m[1861]&m[1862])|(m[1856]&m[1859]&~m[1860]&~m[1861]&m[1862])|(m[1856]&~m[1859]&m[1860]&~m[1861]&m[1862])|(~m[1856]&~m[1859]&~m[1860]&m[1861]&m[1862])|(m[1856]&~m[1859]&~m[1860]&m[1861]&m[1862])|(~m[1856]&m[1859]&~m[1860]&m[1861]&m[1862])|(m[1856]&m[1859]&~m[1860]&m[1861]&m[1862])|(~m[1856]&~m[1859]&m[1860]&m[1861]&m[1862])|(m[1856]&~m[1859]&m[1860]&m[1861]&m[1862])|(m[1856]&m[1859]&m[1860]&m[1861]&m[1862]))):InitCond[473];
    m[1863] = run?((((m[1861]&~m[1864]&~m[1865]&~m[1866]&~m[1867])|(~m[1861]&~m[1864]&~m[1865]&m[1866]&~m[1867])|(m[1861]&m[1864]&~m[1865]&m[1866]&~m[1867])|(m[1861]&~m[1864]&m[1865]&m[1866]&~m[1867])|(~m[1861]&m[1864]&~m[1865]&~m[1866]&m[1867])|(~m[1861]&~m[1864]&m[1865]&~m[1866]&m[1867])|(m[1861]&m[1864]&m[1865]&~m[1866]&m[1867])|(~m[1861]&m[1864]&m[1865]&m[1866]&m[1867]))&UnbiasedRNG[218])|((m[1861]&~m[1864]&~m[1865]&m[1866]&~m[1867])|(~m[1861]&~m[1864]&~m[1865]&~m[1866]&m[1867])|(m[1861]&~m[1864]&~m[1865]&~m[1866]&m[1867])|(m[1861]&m[1864]&~m[1865]&~m[1866]&m[1867])|(m[1861]&~m[1864]&m[1865]&~m[1866]&m[1867])|(~m[1861]&~m[1864]&~m[1865]&m[1866]&m[1867])|(m[1861]&~m[1864]&~m[1865]&m[1866]&m[1867])|(~m[1861]&m[1864]&~m[1865]&m[1866]&m[1867])|(m[1861]&m[1864]&~m[1865]&m[1866]&m[1867])|(~m[1861]&~m[1864]&m[1865]&m[1866]&m[1867])|(m[1861]&~m[1864]&m[1865]&m[1866]&m[1867])|(m[1861]&m[1864]&m[1865]&m[1866]&m[1867]))):InitCond[474];
    m[1868] = run?((((m[1866]&~m[1869]&~m[1870]&~m[1871]&~m[1872])|(~m[1866]&~m[1869]&~m[1870]&m[1871]&~m[1872])|(m[1866]&m[1869]&~m[1870]&m[1871]&~m[1872])|(m[1866]&~m[1869]&m[1870]&m[1871]&~m[1872])|(~m[1866]&m[1869]&~m[1870]&~m[1871]&m[1872])|(~m[1866]&~m[1869]&m[1870]&~m[1871]&m[1872])|(m[1866]&m[1869]&m[1870]&~m[1871]&m[1872])|(~m[1866]&m[1869]&m[1870]&m[1871]&m[1872]))&UnbiasedRNG[219])|((m[1866]&~m[1869]&~m[1870]&m[1871]&~m[1872])|(~m[1866]&~m[1869]&~m[1870]&~m[1871]&m[1872])|(m[1866]&~m[1869]&~m[1870]&~m[1871]&m[1872])|(m[1866]&m[1869]&~m[1870]&~m[1871]&m[1872])|(m[1866]&~m[1869]&m[1870]&~m[1871]&m[1872])|(~m[1866]&~m[1869]&~m[1870]&m[1871]&m[1872])|(m[1866]&~m[1869]&~m[1870]&m[1871]&m[1872])|(~m[1866]&m[1869]&~m[1870]&m[1871]&m[1872])|(m[1866]&m[1869]&~m[1870]&m[1871]&m[1872])|(~m[1866]&~m[1869]&m[1870]&m[1871]&m[1872])|(m[1866]&~m[1869]&m[1870]&m[1871]&m[1872])|(m[1866]&m[1869]&m[1870]&m[1871]&m[1872]))):InitCond[475];
    m[1873] = run?((((m[1871]&~m[1874]&~m[1875]&~m[1876]&~m[1877])|(~m[1871]&~m[1874]&~m[1875]&m[1876]&~m[1877])|(m[1871]&m[1874]&~m[1875]&m[1876]&~m[1877])|(m[1871]&~m[1874]&m[1875]&m[1876]&~m[1877])|(~m[1871]&m[1874]&~m[1875]&~m[1876]&m[1877])|(~m[1871]&~m[1874]&m[1875]&~m[1876]&m[1877])|(m[1871]&m[1874]&m[1875]&~m[1876]&m[1877])|(~m[1871]&m[1874]&m[1875]&m[1876]&m[1877]))&UnbiasedRNG[220])|((m[1871]&~m[1874]&~m[1875]&m[1876]&~m[1877])|(~m[1871]&~m[1874]&~m[1875]&~m[1876]&m[1877])|(m[1871]&~m[1874]&~m[1875]&~m[1876]&m[1877])|(m[1871]&m[1874]&~m[1875]&~m[1876]&m[1877])|(m[1871]&~m[1874]&m[1875]&~m[1876]&m[1877])|(~m[1871]&~m[1874]&~m[1875]&m[1876]&m[1877])|(m[1871]&~m[1874]&~m[1875]&m[1876]&m[1877])|(~m[1871]&m[1874]&~m[1875]&m[1876]&m[1877])|(m[1871]&m[1874]&~m[1875]&m[1876]&m[1877])|(~m[1871]&~m[1874]&m[1875]&m[1876]&m[1877])|(m[1871]&~m[1874]&m[1875]&m[1876]&m[1877])|(m[1871]&m[1874]&m[1875]&m[1876]&m[1877]))):InitCond[476];
    m[1878] = run?((((m[1876]&~m[1879]&~m[1880]&~m[1881]&~m[1882])|(~m[1876]&~m[1879]&~m[1880]&m[1881]&~m[1882])|(m[1876]&m[1879]&~m[1880]&m[1881]&~m[1882])|(m[1876]&~m[1879]&m[1880]&m[1881]&~m[1882])|(~m[1876]&m[1879]&~m[1880]&~m[1881]&m[1882])|(~m[1876]&~m[1879]&m[1880]&~m[1881]&m[1882])|(m[1876]&m[1879]&m[1880]&~m[1881]&m[1882])|(~m[1876]&m[1879]&m[1880]&m[1881]&m[1882]))&UnbiasedRNG[221])|((m[1876]&~m[1879]&~m[1880]&m[1881]&~m[1882])|(~m[1876]&~m[1879]&~m[1880]&~m[1881]&m[1882])|(m[1876]&~m[1879]&~m[1880]&~m[1881]&m[1882])|(m[1876]&m[1879]&~m[1880]&~m[1881]&m[1882])|(m[1876]&~m[1879]&m[1880]&~m[1881]&m[1882])|(~m[1876]&~m[1879]&~m[1880]&m[1881]&m[1882])|(m[1876]&~m[1879]&~m[1880]&m[1881]&m[1882])|(~m[1876]&m[1879]&~m[1880]&m[1881]&m[1882])|(m[1876]&m[1879]&~m[1880]&m[1881]&m[1882])|(~m[1876]&~m[1879]&m[1880]&m[1881]&m[1882])|(m[1876]&~m[1879]&m[1880]&m[1881]&m[1882])|(m[1876]&m[1879]&m[1880]&m[1881]&m[1882]))):InitCond[477];
    m[1883] = run?((((m[1881]&~m[1884]&~m[1885]&~m[1886]&~m[1887])|(~m[1881]&~m[1884]&~m[1885]&m[1886]&~m[1887])|(m[1881]&m[1884]&~m[1885]&m[1886]&~m[1887])|(m[1881]&~m[1884]&m[1885]&m[1886]&~m[1887])|(~m[1881]&m[1884]&~m[1885]&~m[1886]&m[1887])|(~m[1881]&~m[1884]&m[1885]&~m[1886]&m[1887])|(m[1881]&m[1884]&m[1885]&~m[1886]&m[1887])|(~m[1881]&m[1884]&m[1885]&m[1886]&m[1887]))&UnbiasedRNG[222])|((m[1881]&~m[1884]&~m[1885]&m[1886]&~m[1887])|(~m[1881]&~m[1884]&~m[1885]&~m[1886]&m[1887])|(m[1881]&~m[1884]&~m[1885]&~m[1886]&m[1887])|(m[1881]&m[1884]&~m[1885]&~m[1886]&m[1887])|(m[1881]&~m[1884]&m[1885]&~m[1886]&m[1887])|(~m[1881]&~m[1884]&~m[1885]&m[1886]&m[1887])|(m[1881]&~m[1884]&~m[1885]&m[1886]&m[1887])|(~m[1881]&m[1884]&~m[1885]&m[1886]&m[1887])|(m[1881]&m[1884]&~m[1885]&m[1886]&m[1887])|(~m[1881]&~m[1884]&m[1885]&m[1886]&m[1887])|(m[1881]&~m[1884]&m[1885]&m[1886]&m[1887])|(m[1881]&m[1884]&m[1885]&m[1886]&m[1887]))):InitCond[478];
    m[1888] = run?((((m[1886]&~m[1889]&~m[1890]&~m[1891]&~m[1892])|(~m[1886]&~m[1889]&~m[1890]&m[1891]&~m[1892])|(m[1886]&m[1889]&~m[1890]&m[1891]&~m[1892])|(m[1886]&~m[1889]&m[1890]&m[1891]&~m[1892])|(~m[1886]&m[1889]&~m[1890]&~m[1891]&m[1892])|(~m[1886]&~m[1889]&m[1890]&~m[1891]&m[1892])|(m[1886]&m[1889]&m[1890]&~m[1891]&m[1892])|(~m[1886]&m[1889]&m[1890]&m[1891]&m[1892]))&UnbiasedRNG[223])|((m[1886]&~m[1889]&~m[1890]&m[1891]&~m[1892])|(~m[1886]&~m[1889]&~m[1890]&~m[1891]&m[1892])|(m[1886]&~m[1889]&~m[1890]&~m[1891]&m[1892])|(m[1886]&m[1889]&~m[1890]&~m[1891]&m[1892])|(m[1886]&~m[1889]&m[1890]&~m[1891]&m[1892])|(~m[1886]&~m[1889]&~m[1890]&m[1891]&m[1892])|(m[1886]&~m[1889]&~m[1890]&m[1891]&m[1892])|(~m[1886]&m[1889]&~m[1890]&m[1891]&m[1892])|(m[1886]&m[1889]&~m[1890]&m[1891]&m[1892])|(~m[1886]&~m[1889]&m[1890]&m[1891]&m[1892])|(m[1886]&~m[1889]&m[1890]&m[1891]&m[1892])|(m[1886]&m[1889]&m[1890]&m[1891]&m[1892]))):InitCond[479];
    m[1893] = run?((((m[1891]&~m[1894]&~m[1895]&~m[1896]&~m[1897])|(~m[1891]&~m[1894]&~m[1895]&m[1896]&~m[1897])|(m[1891]&m[1894]&~m[1895]&m[1896]&~m[1897])|(m[1891]&~m[1894]&m[1895]&m[1896]&~m[1897])|(~m[1891]&m[1894]&~m[1895]&~m[1896]&m[1897])|(~m[1891]&~m[1894]&m[1895]&~m[1896]&m[1897])|(m[1891]&m[1894]&m[1895]&~m[1896]&m[1897])|(~m[1891]&m[1894]&m[1895]&m[1896]&m[1897]))&UnbiasedRNG[224])|((m[1891]&~m[1894]&~m[1895]&m[1896]&~m[1897])|(~m[1891]&~m[1894]&~m[1895]&~m[1896]&m[1897])|(m[1891]&~m[1894]&~m[1895]&~m[1896]&m[1897])|(m[1891]&m[1894]&~m[1895]&~m[1896]&m[1897])|(m[1891]&~m[1894]&m[1895]&~m[1896]&m[1897])|(~m[1891]&~m[1894]&~m[1895]&m[1896]&m[1897])|(m[1891]&~m[1894]&~m[1895]&m[1896]&m[1897])|(~m[1891]&m[1894]&~m[1895]&m[1896]&m[1897])|(m[1891]&m[1894]&~m[1895]&m[1896]&m[1897])|(~m[1891]&~m[1894]&m[1895]&m[1896]&m[1897])|(m[1891]&~m[1894]&m[1895]&m[1896]&m[1897])|(m[1891]&m[1894]&m[1895]&m[1896]&m[1897]))):InitCond[480];
    m[1898] = run?((((m[1896]&~m[1899]&~m[1900]&~m[1901]&~m[1902])|(~m[1896]&~m[1899]&~m[1900]&m[1901]&~m[1902])|(m[1896]&m[1899]&~m[1900]&m[1901]&~m[1902])|(m[1896]&~m[1899]&m[1900]&m[1901]&~m[1902])|(~m[1896]&m[1899]&~m[1900]&~m[1901]&m[1902])|(~m[1896]&~m[1899]&m[1900]&~m[1901]&m[1902])|(m[1896]&m[1899]&m[1900]&~m[1901]&m[1902])|(~m[1896]&m[1899]&m[1900]&m[1901]&m[1902]))&UnbiasedRNG[225])|((m[1896]&~m[1899]&~m[1900]&m[1901]&~m[1902])|(~m[1896]&~m[1899]&~m[1900]&~m[1901]&m[1902])|(m[1896]&~m[1899]&~m[1900]&~m[1901]&m[1902])|(m[1896]&m[1899]&~m[1900]&~m[1901]&m[1902])|(m[1896]&~m[1899]&m[1900]&~m[1901]&m[1902])|(~m[1896]&~m[1899]&~m[1900]&m[1901]&m[1902])|(m[1896]&~m[1899]&~m[1900]&m[1901]&m[1902])|(~m[1896]&m[1899]&~m[1900]&m[1901]&m[1902])|(m[1896]&m[1899]&~m[1900]&m[1901]&m[1902])|(~m[1896]&~m[1899]&m[1900]&m[1901]&m[1902])|(m[1896]&~m[1899]&m[1900]&m[1901]&m[1902])|(m[1896]&m[1899]&m[1900]&m[1901]&m[1902]))):InitCond[481];
    m[1903] = run?((((m[1857]&~m[1904]&~m[1905]&~m[1906]&~m[1907])|(~m[1857]&~m[1904]&~m[1905]&m[1906]&~m[1907])|(m[1857]&m[1904]&~m[1905]&m[1906]&~m[1907])|(m[1857]&~m[1904]&m[1905]&m[1906]&~m[1907])|(~m[1857]&m[1904]&~m[1905]&~m[1906]&m[1907])|(~m[1857]&~m[1904]&m[1905]&~m[1906]&m[1907])|(m[1857]&m[1904]&m[1905]&~m[1906]&m[1907])|(~m[1857]&m[1904]&m[1905]&m[1906]&m[1907]))&UnbiasedRNG[226])|((m[1857]&~m[1904]&~m[1905]&m[1906]&~m[1907])|(~m[1857]&~m[1904]&~m[1905]&~m[1906]&m[1907])|(m[1857]&~m[1904]&~m[1905]&~m[1906]&m[1907])|(m[1857]&m[1904]&~m[1905]&~m[1906]&m[1907])|(m[1857]&~m[1904]&m[1905]&~m[1906]&m[1907])|(~m[1857]&~m[1904]&~m[1905]&m[1906]&m[1907])|(m[1857]&~m[1904]&~m[1905]&m[1906]&m[1907])|(~m[1857]&m[1904]&~m[1905]&m[1906]&m[1907])|(m[1857]&m[1904]&~m[1905]&m[1906]&m[1907])|(~m[1857]&~m[1904]&m[1905]&m[1906]&m[1907])|(m[1857]&~m[1904]&m[1905]&m[1906]&m[1907])|(m[1857]&m[1904]&m[1905]&m[1906]&m[1907]))):InitCond[482];
    m[1908] = run?((((m[1906]&~m[1909]&~m[1910]&~m[1911]&~m[1912])|(~m[1906]&~m[1909]&~m[1910]&m[1911]&~m[1912])|(m[1906]&m[1909]&~m[1910]&m[1911]&~m[1912])|(m[1906]&~m[1909]&m[1910]&m[1911]&~m[1912])|(~m[1906]&m[1909]&~m[1910]&~m[1911]&m[1912])|(~m[1906]&~m[1909]&m[1910]&~m[1911]&m[1912])|(m[1906]&m[1909]&m[1910]&~m[1911]&m[1912])|(~m[1906]&m[1909]&m[1910]&m[1911]&m[1912]))&UnbiasedRNG[227])|((m[1906]&~m[1909]&~m[1910]&m[1911]&~m[1912])|(~m[1906]&~m[1909]&~m[1910]&~m[1911]&m[1912])|(m[1906]&~m[1909]&~m[1910]&~m[1911]&m[1912])|(m[1906]&m[1909]&~m[1910]&~m[1911]&m[1912])|(m[1906]&~m[1909]&m[1910]&~m[1911]&m[1912])|(~m[1906]&~m[1909]&~m[1910]&m[1911]&m[1912])|(m[1906]&~m[1909]&~m[1910]&m[1911]&m[1912])|(~m[1906]&m[1909]&~m[1910]&m[1911]&m[1912])|(m[1906]&m[1909]&~m[1910]&m[1911]&m[1912])|(~m[1906]&~m[1909]&m[1910]&m[1911]&m[1912])|(m[1906]&~m[1909]&m[1910]&m[1911]&m[1912])|(m[1906]&m[1909]&m[1910]&m[1911]&m[1912]))):InitCond[483];
    m[1913] = run?((((m[1911]&~m[1914]&~m[1915]&~m[1916]&~m[1917])|(~m[1911]&~m[1914]&~m[1915]&m[1916]&~m[1917])|(m[1911]&m[1914]&~m[1915]&m[1916]&~m[1917])|(m[1911]&~m[1914]&m[1915]&m[1916]&~m[1917])|(~m[1911]&m[1914]&~m[1915]&~m[1916]&m[1917])|(~m[1911]&~m[1914]&m[1915]&~m[1916]&m[1917])|(m[1911]&m[1914]&m[1915]&~m[1916]&m[1917])|(~m[1911]&m[1914]&m[1915]&m[1916]&m[1917]))&UnbiasedRNG[228])|((m[1911]&~m[1914]&~m[1915]&m[1916]&~m[1917])|(~m[1911]&~m[1914]&~m[1915]&~m[1916]&m[1917])|(m[1911]&~m[1914]&~m[1915]&~m[1916]&m[1917])|(m[1911]&m[1914]&~m[1915]&~m[1916]&m[1917])|(m[1911]&~m[1914]&m[1915]&~m[1916]&m[1917])|(~m[1911]&~m[1914]&~m[1915]&m[1916]&m[1917])|(m[1911]&~m[1914]&~m[1915]&m[1916]&m[1917])|(~m[1911]&m[1914]&~m[1915]&m[1916]&m[1917])|(m[1911]&m[1914]&~m[1915]&m[1916]&m[1917])|(~m[1911]&~m[1914]&m[1915]&m[1916]&m[1917])|(m[1911]&~m[1914]&m[1915]&m[1916]&m[1917])|(m[1911]&m[1914]&m[1915]&m[1916]&m[1917]))):InitCond[484];
    m[1918] = run?((((m[1916]&~m[1919]&~m[1920]&~m[1921]&~m[1922])|(~m[1916]&~m[1919]&~m[1920]&m[1921]&~m[1922])|(m[1916]&m[1919]&~m[1920]&m[1921]&~m[1922])|(m[1916]&~m[1919]&m[1920]&m[1921]&~m[1922])|(~m[1916]&m[1919]&~m[1920]&~m[1921]&m[1922])|(~m[1916]&~m[1919]&m[1920]&~m[1921]&m[1922])|(m[1916]&m[1919]&m[1920]&~m[1921]&m[1922])|(~m[1916]&m[1919]&m[1920]&m[1921]&m[1922]))&UnbiasedRNG[229])|((m[1916]&~m[1919]&~m[1920]&m[1921]&~m[1922])|(~m[1916]&~m[1919]&~m[1920]&~m[1921]&m[1922])|(m[1916]&~m[1919]&~m[1920]&~m[1921]&m[1922])|(m[1916]&m[1919]&~m[1920]&~m[1921]&m[1922])|(m[1916]&~m[1919]&m[1920]&~m[1921]&m[1922])|(~m[1916]&~m[1919]&~m[1920]&m[1921]&m[1922])|(m[1916]&~m[1919]&~m[1920]&m[1921]&m[1922])|(~m[1916]&m[1919]&~m[1920]&m[1921]&m[1922])|(m[1916]&m[1919]&~m[1920]&m[1921]&m[1922])|(~m[1916]&~m[1919]&m[1920]&m[1921]&m[1922])|(m[1916]&~m[1919]&m[1920]&m[1921]&m[1922])|(m[1916]&m[1919]&m[1920]&m[1921]&m[1922]))):InitCond[485];
    m[1923] = run?((((m[1921]&~m[1924]&~m[1925]&~m[1926]&~m[1927])|(~m[1921]&~m[1924]&~m[1925]&m[1926]&~m[1927])|(m[1921]&m[1924]&~m[1925]&m[1926]&~m[1927])|(m[1921]&~m[1924]&m[1925]&m[1926]&~m[1927])|(~m[1921]&m[1924]&~m[1925]&~m[1926]&m[1927])|(~m[1921]&~m[1924]&m[1925]&~m[1926]&m[1927])|(m[1921]&m[1924]&m[1925]&~m[1926]&m[1927])|(~m[1921]&m[1924]&m[1925]&m[1926]&m[1927]))&UnbiasedRNG[230])|((m[1921]&~m[1924]&~m[1925]&m[1926]&~m[1927])|(~m[1921]&~m[1924]&~m[1925]&~m[1926]&m[1927])|(m[1921]&~m[1924]&~m[1925]&~m[1926]&m[1927])|(m[1921]&m[1924]&~m[1925]&~m[1926]&m[1927])|(m[1921]&~m[1924]&m[1925]&~m[1926]&m[1927])|(~m[1921]&~m[1924]&~m[1925]&m[1926]&m[1927])|(m[1921]&~m[1924]&~m[1925]&m[1926]&m[1927])|(~m[1921]&m[1924]&~m[1925]&m[1926]&m[1927])|(m[1921]&m[1924]&~m[1925]&m[1926]&m[1927])|(~m[1921]&~m[1924]&m[1925]&m[1926]&m[1927])|(m[1921]&~m[1924]&m[1925]&m[1926]&m[1927])|(m[1921]&m[1924]&m[1925]&m[1926]&m[1927]))):InitCond[486];
    m[1928] = run?((((m[1926]&~m[1929]&~m[1930]&~m[1931]&~m[1932])|(~m[1926]&~m[1929]&~m[1930]&m[1931]&~m[1932])|(m[1926]&m[1929]&~m[1930]&m[1931]&~m[1932])|(m[1926]&~m[1929]&m[1930]&m[1931]&~m[1932])|(~m[1926]&m[1929]&~m[1930]&~m[1931]&m[1932])|(~m[1926]&~m[1929]&m[1930]&~m[1931]&m[1932])|(m[1926]&m[1929]&m[1930]&~m[1931]&m[1932])|(~m[1926]&m[1929]&m[1930]&m[1931]&m[1932]))&UnbiasedRNG[231])|((m[1926]&~m[1929]&~m[1930]&m[1931]&~m[1932])|(~m[1926]&~m[1929]&~m[1930]&~m[1931]&m[1932])|(m[1926]&~m[1929]&~m[1930]&~m[1931]&m[1932])|(m[1926]&m[1929]&~m[1930]&~m[1931]&m[1932])|(m[1926]&~m[1929]&m[1930]&~m[1931]&m[1932])|(~m[1926]&~m[1929]&~m[1930]&m[1931]&m[1932])|(m[1926]&~m[1929]&~m[1930]&m[1931]&m[1932])|(~m[1926]&m[1929]&~m[1930]&m[1931]&m[1932])|(m[1926]&m[1929]&~m[1930]&m[1931]&m[1932])|(~m[1926]&~m[1929]&m[1930]&m[1931]&m[1932])|(m[1926]&~m[1929]&m[1930]&m[1931]&m[1932])|(m[1926]&m[1929]&m[1930]&m[1931]&m[1932]))):InitCond[487];
    m[1933] = run?((((m[1931]&~m[1934]&~m[1935]&~m[1936]&~m[1937])|(~m[1931]&~m[1934]&~m[1935]&m[1936]&~m[1937])|(m[1931]&m[1934]&~m[1935]&m[1936]&~m[1937])|(m[1931]&~m[1934]&m[1935]&m[1936]&~m[1937])|(~m[1931]&m[1934]&~m[1935]&~m[1936]&m[1937])|(~m[1931]&~m[1934]&m[1935]&~m[1936]&m[1937])|(m[1931]&m[1934]&m[1935]&~m[1936]&m[1937])|(~m[1931]&m[1934]&m[1935]&m[1936]&m[1937]))&UnbiasedRNG[232])|((m[1931]&~m[1934]&~m[1935]&m[1936]&~m[1937])|(~m[1931]&~m[1934]&~m[1935]&~m[1936]&m[1937])|(m[1931]&~m[1934]&~m[1935]&~m[1936]&m[1937])|(m[1931]&m[1934]&~m[1935]&~m[1936]&m[1937])|(m[1931]&~m[1934]&m[1935]&~m[1936]&m[1937])|(~m[1931]&~m[1934]&~m[1935]&m[1936]&m[1937])|(m[1931]&~m[1934]&~m[1935]&m[1936]&m[1937])|(~m[1931]&m[1934]&~m[1935]&m[1936]&m[1937])|(m[1931]&m[1934]&~m[1935]&m[1936]&m[1937])|(~m[1931]&~m[1934]&m[1935]&m[1936]&m[1937])|(m[1931]&~m[1934]&m[1935]&m[1936]&m[1937])|(m[1931]&m[1934]&m[1935]&m[1936]&m[1937]))):InitCond[488];
    m[1938] = run?((((m[1936]&~m[1939]&~m[1940]&~m[1941]&~m[1942])|(~m[1936]&~m[1939]&~m[1940]&m[1941]&~m[1942])|(m[1936]&m[1939]&~m[1940]&m[1941]&~m[1942])|(m[1936]&~m[1939]&m[1940]&m[1941]&~m[1942])|(~m[1936]&m[1939]&~m[1940]&~m[1941]&m[1942])|(~m[1936]&~m[1939]&m[1940]&~m[1941]&m[1942])|(m[1936]&m[1939]&m[1940]&~m[1941]&m[1942])|(~m[1936]&m[1939]&m[1940]&m[1941]&m[1942]))&UnbiasedRNG[233])|((m[1936]&~m[1939]&~m[1940]&m[1941]&~m[1942])|(~m[1936]&~m[1939]&~m[1940]&~m[1941]&m[1942])|(m[1936]&~m[1939]&~m[1940]&~m[1941]&m[1942])|(m[1936]&m[1939]&~m[1940]&~m[1941]&m[1942])|(m[1936]&~m[1939]&m[1940]&~m[1941]&m[1942])|(~m[1936]&~m[1939]&~m[1940]&m[1941]&m[1942])|(m[1936]&~m[1939]&~m[1940]&m[1941]&m[1942])|(~m[1936]&m[1939]&~m[1940]&m[1941]&m[1942])|(m[1936]&m[1939]&~m[1940]&m[1941]&m[1942])|(~m[1936]&~m[1939]&m[1940]&m[1941]&m[1942])|(m[1936]&~m[1939]&m[1940]&m[1941]&m[1942])|(m[1936]&m[1939]&m[1940]&m[1941]&m[1942]))):InitCond[489];
    m[1943] = run?((((m[1941]&~m[1944]&~m[1945]&~m[1946]&~m[1947])|(~m[1941]&~m[1944]&~m[1945]&m[1946]&~m[1947])|(m[1941]&m[1944]&~m[1945]&m[1946]&~m[1947])|(m[1941]&~m[1944]&m[1945]&m[1946]&~m[1947])|(~m[1941]&m[1944]&~m[1945]&~m[1946]&m[1947])|(~m[1941]&~m[1944]&m[1945]&~m[1946]&m[1947])|(m[1941]&m[1944]&m[1945]&~m[1946]&m[1947])|(~m[1941]&m[1944]&m[1945]&m[1946]&m[1947]))&UnbiasedRNG[234])|((m[1941]&~m[1944]&~m[1945]&m[1946]&~m[1947])|(~m[1941]&~m[1944]&~m[1945]&~m[1946]&m[1947])|(m[1941]&~m[1944]&~m[1945]&~m[1946]&m[1947])|(m[1941]&m[1944]&~m[1945]&~m[1946]&m[1947])|(m[1941]&~m[1944]&m[1945]&~m[1946]&m[1947])|(~m[1941]&~m[1944]&~m[1945]&m[1946]&m[1947])|(m[1941]&~m[1944]&~m[1945]&m[1946]&m[1947])|(~m[1941]&m[1944]&~m[1945]&m[1946]&m[1947])|(m[1941]&m[1944]&~m[1945]&m[1946]&m[1947])|(~m[1941]&~m[1944]&m[1945]&m[1946]&m[1947])|(m[1941]&~m[1944]&m[1945]&m[1946]&m[1947])|(m[1941]&m[1944]&m[1945]&m[1946]&m[1947]))):InitCond[490];
    m[1948] = run?((((m[1907]&~m[1949]&~m[1950]&~m[1951]&~m[1952])|(~m[1907]&~m[1949]&~m[1950]&m[1951]&~m[1952])|(m[1907]&m[1949]&~m[1950]&m[1951]&~m[1952])|(m[1907]&~m[1949]&m[1950]&m[1951]&~m[1952])|(~m[1907]&m[1949]&~m[1950]&~m[1951]&m[1952])|(~m[1907]&~m[1949]&m[1950]&~m[1951]&m[1952])|(m[1907]&m[1949]&m[1950]&~m[1951]&m[1952])|(~m[1907]&m[1949]&m[1950]&m[1951]&m[1952]))&UnbiasedRNG[235])|((m[1907]&~m[1949]&~m[1950]&m[1951]&~m[1952])|(~m[1907]&~m[1949]&~m[1950]&~m[1951]&m[1952])|(m[1907]&~m[1949]&~m[1950]&~m[1951]&m[1952])|(m[1907]&m[1949]&~m[1950]&~m[1951]&m[1952])|(m[1907]&~m[1949]&m[1950]&~m[1951]&m[1952])|(~m[1907]&~m[1949]&~m[1950]&m[1951]&m[1952])|(m[1907]&~m[1949]&~m[1950]&m[1951]&m[1952])|(~m[1907]&m[1949]&~m[1950]&m[1951]&m[1952])|(m[1907]&m[1949]&~m[1950]&m[1951]&m[1952])|(~m[1907]&~m[1949]&m[1950]&m[1951]&m[1952])|(m[1907]&~m[1949]&m[1950]&m[1951]&m[1952])|(m[1907]&m[1949]&m[1950]&m[1951]&m[1952]))):InitCond[491];
    m[1953] = run?((((m[1951]&~m[1954]&~m[1955]&~m[1956]&~m[1957])|(~m[1951]&~m[1954]&~m[1955]&m[1956]&~m[1957])|(m[1951]&m[1954]&~m[1955]&m[1956]&~m[1957])|(m[1951]&~m[1954]&m[1955]&m[1956]&~m[1957])|(~m[1951]&m[1954]&~m[1955]&~m[1956]&m[1957])|(~m[1951]&~m[1954]&m[1955]&~m[1956]&m[1957])|(m[1951]&m[1954]&m[1955]&~m[1956]&m[1957])|(~m[1951]&m[1954]&m[1955]&m[1956]&m[1957]))&UnbiasedRNG[236])|((m[1951]&~m[1954]&~m[1955]&m[1956]&~m[1957])|(~m[1951]&~m[1954]&~m[1955]&~m[1956]&m[1957])|(m[1951]&~m[1954]&~m[1955]&~m[1956]&m[1957])|(m[1951]&m[1954]&~m[1955]&~m[1956]&m[1957])|(m[1951]&~m[1954]&m[1955]&~m[1956]&m[1957])|(~m[1951]&~m[1954]&~m[1955]&m[1956]&m[1957])|(m[1951]&~m[1954]&~m[1955]&m[1956]&m[1957])|(~m[1951]&m[1954]&~m[1955]&m[1956]&m[1957])|(m[1951]&m[1954]&~m[1955]&m[1956]&m[1957])|(~m[1951]&~m[1954]&m[1955]&m[1956]&m[1957])|(m[1951]&~m[1954]&m[1955]&m[1956]&m[1957])|(m[1951]&m[1954]&m[1955]&m[1956]&m[1957]))):InitCond[492];
    m[1958] = run?((((m[1956]&~m[1959]&~m[1960]&~m[1961]&~m[1962])|(~m[1956]&~m[1959]&~m[1960]&m[1961]&~m[1962])|(m[1956]&m[1959]&~m[1960]&m[1961]&~m[1962])|(m[1956]&~m[1959]&m[1960]&m[1961]&~m[1962])|(~m[1956]&m[1959]&~m[1960]&~m[1961]&m[1962])|(~m[1956]&~m[1959]&m[1960]&~m[1961]&m[1962])|(m[1956]&m[1959]&m[1960]&~m[1961]&m[1962])|(~m[1956]&m[1959]&m[1960]&m[1961]&m[1962]))&UnbiasedRNG[237])|((m[1956]&~m[1959]&~m[1960]&m[1961]&~m[1962])|(~m[1956]&~m[1959]&~m[1960]&~m[1961]&m[1962])|(m[1956]&~m[1959]&~m[1960]&~m[1961]&m[1962])|(m[1956]&m[1959]&~m[1960]&~m[1961]&m[1962])|(m[1956]&~m[1959]&m[1960]&~m[1961]&m[1962])|(~m[1956]&~m[1959]&~m[1960]&m[1961]&m[1962])|(m[1956]&~m[1959]&~m[1960]&m[1961]&m[1962])|(~m[1956]&m[1959]&~m[1960]&m[1961]&m[1962])|(m[1956]&m[1959]&~m[1960]&m[1961]&m[1962])|(~m[1956]&~m[1959]&m[1960]&m[1961]&m[1962])|(m[1956]&~m[1959]&m[1960]&m[1961]&m[1962])|(m[1956]&m[1959]&m[1960]&m[1961]&m[1962]))):InitCond[493];
    m[1963] = run?((((m[1961]&~m[1964]&~m[1965]&~m[1966]&~m[1967])|(~m[1961]&~m[1964]&~m[1965]&m[1966]&~m[1967])|(m[1961]&m[1964]&~m[1965]&m[1966]&~m[1967])|(m[1961]&~m[1964]&m[1965]&m[1966]&~m[1967])|(~m[1961]&m[1964]&~m[1965]&~m[1966]&m[1967])|(~m[1961]&~m[1964]&m[1965]&~m[1966]&m[1967])|(m[1961]&m[1964]&m[1965]&~m[1966]&m[1967])|(~m[1961]&m[1964]&m[1965]&m[1966]&m[1967]))&UnbiasedRNG[238])|((m[1961]&~m[1964]&~m[1965]&m[1966]&~m[1967])|(~m[1961]&~m[1964]&~m[1965]&~m[1966]&m[1967])|(m[1961]&~m[1964]&~m[1965]&~m[1966]&m[1967])|(m[1961]&m[1964]&~m[1965]&~m[1966]&m[1967])|(m[1961]&~m[1964]&m[1965]&~m[1966]&m[1967])|(~m[1961]&~m[1964]&~m[1965]&m[1966]&m[1967])|(m[1961]&~m[1964]&~m[1965]&m[1966]&m[1967])|(~m[1961]&m[1964]&~m[1965]&m[1966]&m[1967])|(m[1961]&m[1964]&~m[1965]&m[1966]&m[1967])|(~m[1961]&~m[1964]&m[1965]&m[1966]&m[1967])|(m[1961]&~m[1964]&m[1965]&m[1966]&m[1967])|(m[1961]&m[1964]&m[1965]&m[1966]&m[1967]))):InitCond[494];
    m[1968] = run?((((m[1966]&~m[1969]&~m[1970]&~m[1971]&~m[1972])|(~m[1966]&~m[1969]&~m[1970]&m[1971]&~m[1972])|(m[1966]&m[1969]&~m[1970]&m[1971]&~m[1972])|(m[1966]&~m[1969]&m[1970]&m[1971]&~m[1972])|(~m[1966]&m[1969]&~m[1970]&~m[1971]&m[1972])|(~m[1966]&~m[1969]&m[1970]&~m[1971]&m[1972])|(m[1966]&m[1969]&m[1970]&~m[1971]&m[1972])|(~m[1966]&m[1969]&m[1970]&m[1971]&m[1972]))&UnbiasedRNG[239])|((m[1966]&~m[1969]&~m[1970]&m[1971]&~m[1972])|(~m[1966]&~m[1969]&~m[1970]&~m[1971]&m[1972])|(m[1966]&~m[1969]&~m[1970]&~m[1971]&m[1972])|(m[1966]&m[1969]&~m[1970]&~m[1971]&m[1972])|(m[1966]&~m[1969]&m[1970]&~m[1971]&m[1972])|(~m[1966]&~m[1969]&~m[1970]&m[1971]&m[1972])|(m[1966]&~m[1969]&~m[1970]&m[1971]&m[1972])|(~m[1966]&m[1969]&~m[1970]&m[1971]&m[1972])|(m[1966]&m[1969]&~m[1970]&m[1971]&m[1972])|(~m[1966]&~m[1969]&m[1970]&m[1971]&m[1972])|(m[1966]&~m[1969]&m[1970]&m[1971]&m[1972])|(m[1966]&m[1969]&m[1970]&m[1971]&m[1972]))):InitCond[495];
    m[1973] = run?((((m[1971]&~m[1974]&~m[1975]&~m[1976]&~m[1977])|(~m[1971]&~m[1974]&~m[1975]&m[1976]&~m[1977])|(m[1971]&m[1974]&~m[1975]&m[1976]&~m[1977])|(m[1971]&~m[1974]&m[1975]&m[1976]&~m[1977])|(~m[1971]&m[1974]&~m[1975]&~m[1976]&m[1977])|(~m[1971]&~m[1974]&m[1975]&~m[1976]&m[1977])|(m[1971]&m[1974]&m[1975]&~m[1976]&m[1977])|(~m[1971]&m[1974]&m[1975]&m[1976]&m[1977]))&UnbiasedRNG[240])|((m[1971]&~m[1974]&~m[1975]&m[1976]&~m[1977])|(~m[1971]&~m[1974]&~m[1975]&~m[1976]&m[1977])|(m[1971]&~m[1974]&~m[1975]&~m[1976]&m[1977])|(m[1971]&m[1974]&~m[1975]&~m[1976]&m[1977])|(m[1971]&~m[1974]&m[1975]&~m[1976]&m[1977])|(~m[1971]&~m[1974]&~m[1975]&m[1976]&m[1977])|(m[1971]&~m[1974]&~m[1975]&m[1976]&m[1977])|(~m[1971]&m[1974]&~m[1975]&m[1976]&m[1977])|(m[1971]&m[1974]&~m[1975]&m[1976]&m[1977])|(~m[1971]&~m[1974]&m[1975]&m[1976]&m[1977])|(m[1971]&~m[1974]&m[1975]&m[1976]&m[1977])|(m[1971]&m[1974]&m[1975]&m[1976]&m[1977]))):InitCond[496];
    m[1978] = run?((((m[1976]&~m[1979]&~m[1980]&~m[1981]&~m[1982])|(~m[1976]&~m[1979]&~m[1980]&m[1981]&~m[1982])|(m[1976]&m[1979]&~m[1980]&m[1981]&~m[1982])|(m[1976]&~m[1979]&m[1980]&m[1981]&~m[1982])|(~m[1976]&m[1979]&~m[1980]&~m[1981]&m[1982])|(~m[1976]&~m[1979]&m[1980]&~m[1981]&m[1982])|(m[1976]&m[1979]&m[1980]&~m[1981]&m[1982])|(~m[1976]&m[1979]&m[1980]&m[1981]&m[1982]))&UnbiasedRNG[241])|((m[1976]&~m[1979]&~m[1980]&m[1981]&~m[1982])|(~m[1976]&~m[1979]&~m[1980]&~m[1981]&m[1982])|(m[1976]&~m[1979]&~m[1980]&~m[1981]&m[1982])|(m[1976]&m[1979]&~m[1980]&~m[1981]&m[1982])|(m[1976]&~m[1979]&m[1980]&~m[1981]&m[1982])|(~m[1976]&~m[1979]&~m[1980]&m[1981]&m[1982])|(m[1976]&~m[1979]&~m[1980]&m[1981]&m[1982])|(~m[1976]&m[1979]&~m[1980]&m[1981]&m[1982])|(m[1976]&m[1979]&~m[1980]&m[1981]&m[1982])|(~m[1976]&~m[1979]&m[1980]&m[1981]&m[1982])|(m[1976]&~m[1979]&m[1980]&m[1981]&m[1982])|(m[1976]&m[1979]&m[1980]&m[1981]&m[1982]))):InitCond[497];
    m[1983] = run?((((m[1981]&~m[1984]&~m[1985]&~m[1986]&~m[1987])|(~m[1981]&~m[1984]&~m[1985]&m[1986]&~m[1987])|(m[1981]&m[1984]&~m[1985]&m[1986]&~m[1987])|(m[1981]&~m[1984]&m[1985]&m[1986]&~m[1987])|(~m[1981]&m[1984]&~m[1985]&~m[1986]&m[1987])|(~m[1981]&~m[1984]&m[1985]&~m[1986]&m[1987])|(m[1981]&m[1984]&m[1985]&~m[1986]&m[1987])|(~m[1981]&m[1984]&m[1985]&m[1986]&m[1987]))&UnbiasedRNG[242])|((m[1981]&~m[1984]&~m[1985]&m[1986]&~m[1987])|(~m[1981]&~m[1984]&~m[1985]&~m[1986]&m[1987])|(m[1981]&~m[1984]&~m[1985]&~m[1986]&m[1987])|(m[1981]&m[1984]&~m[1985]&~m[1986]&m[1987])|(m[1981]&~m[1984]&m[1985]&~m[1986]&m[1987])|(~m[1981]&~m[1984]&~m[1985]&m[1986]&m[1987])|(m[1981]&~m[1984]&~m[1985]&m[1986]&m[1987])|(~m[1981]&m[1984]&~m[1985]&m[1986]&m[1987])|(m[1981]&m[1984]&~m[1985]&m[1986]&m[1987])|(~m[1981]&~m[1984]&m[1985]&m[1986]&m[1987])|(m[1981]&~m[1984]&m[1985]&m[1986]&m[1987])|(m[1981]&m[1984]&m[1985]&m[1986]&m[1987]))):InitCond[498];
    m[1988] = run?((((m[1952]&~m[1989]&~m[1990]&~m[1991]&~m[1992])|(~m[1952]&~m[1989]&~m[1990]&m[1991]&~m[1992])|(m[1952]&m[1989]&~m[1990]&m[1991]&~m[1992])|(m[1952]&~m[1989]&m[1990]&m[1991]&~m[1992])|(~m[1952]&m[1989]&~m[1990]&~m[1991]&m[1992])|(~m[1952]&~m[1989]&m[1990]&~m[1991]&m[1992])|(m[1952]&m[1989]&m[1990]&~m[1991]&m[1992])|(~m[1952]&m[1989]&m[1990]&m[1991]&m[1992]))&UnbiasedRNG[243])|((m[1952]&~m[1989]&~m[1990]&m[1991]&~m[1992])|(~m[1952]&~m[1989]&~m[1990]&~m[1991]&m[1992])|(m[1952]&~m[1989]&~m[1990]&~m[1991]&m[1992])|(m[1952]&m[1989]&~m[1990]&~m[1991]&m[1992])|(m[1952]&~m[1989]&m[1990]&~m[1991]&m[1992])|(~m[1952]&~m[1989]&~m[1990]&m[1991]&m[1992])|(m[1952]&~m[1989]&~m[1990]&m[1991]&m[1992])|(~m[1952]&m[1989]&~m[1990]&m[1991]&m[1992])|(m[1952]&m[1989]&~m[1990]&m[1991]&m[1992])|(~m[1952]&~m[1989]&m[1990]&m[1991]&m[1992])|(m[1952]&~m[1989]&m[1990]&m[1991]&m[1992])|(m[1952]&m[1989]&m[1990]&m[1991]&m[1992]))):InitCond[499];
    m[1993] = run?((((m[1991]&~m[1994]&~m[1995]&~m[1996]&~m[1997])|(~m[1991]&~m[1994]&~m[1995]&m[1996]&~m[1997])|(m[1991]&m[1994]&~m[1995]&m[1996]&~m[1997])|(m[1991]&~m[1994]&m[1995]&m[1996]&~m[1997])|(~m[1991]&m[1994]&~m[1995]&~m[1996]&m[1997])|(~m[1991]&~m[1994]&m[1995]&~m[1996]&m[1997])|(m[1991]&m[1994]&m[1995]&~m[1996]&m[1997])|(~m[1991]&m[1994]&m[1995]&m[1996]&m[1997]))&UnbiasedRNG[244])|((m[1991]&~m[1994]&~m[1995]&m[1996]&~m[1997])|(~m[1991]&~m[1994]&~m[1995]&~m[1996]&m[1997])|(m[1991]&~m[1994]&~m[1995]&~m[1996]&m[1997])|(m[1991]&m[1994]&~m[1995]&~m[1996]&m[1997])|(m[1991]&~m[1994]&m[1995]&~m[1996]&m[1997])|(~m[1991]&~m[1994]&~m[1995]&m[1996]&m[1997])|(m[1991]&~m[1994]&~m[1995]&m[1996]&m[1997])|(~m[1991]&m[1994]&~m[1995]&m[1996]&m[1997])|(m[1991]&m[1994]&~m[1995]&m[1996]&m[1997])|(~m[1991]&~m[1994]&m[1995]&m[1996]&m[1997])|(m[1991]&~m[1994]&m[1995]&m[1996]&m[1997])|(m[1991]&m[1994]&m[1995]&m[1996]&m[1997]))):InitCond[500];
    m[1998] = run?((((m[1996]&~m[1999]&~m[2000]&~m[2001]&~m[2002])|(~m[1996]&~m[1999]&~m[2000]&m[2001]&~m[2002])|(m[1996]&m[1999]&~m[2000]&m[2001]&~m[2002])|(m[1996]&~m[1999]&m[2000]&m[2001]&~m[2002])|(~m[1996]&m[1999]&~m[2000]&~m[2001]&m[2002])|(~m[1996]&~m[1999]&m[2000]&~m[2001]&m[2002])|(m[1996]&m[1999]&m[2000]&~m[2001]&m[2002])|(~m[1996]&m[1999]&m[2000]&m[2001]&m[2002]))&UnbiasedRNG[245])|((m[1996]&~m[1999]&~m[2000]&m[2001]&~m[2002])|(~m[1996]&~m[1999]&~m[2000]&~m[2001]&m[2002])|(m[1996]&~m[1999]&~m[2000]&~m[2001]&m[2002])|(m[1996]&m[1999]&~m[2000]&~m[2001]&m[2002])|(m[1996]&~m[1999]&m[2000]&~m[2001]&m[2002])|(~m[1996]&~m[1999]&~m[2000]&m[2001]&m[2002])|(m[1996]&~m[1999]&~m[2000]&m[2001]&m[2002])|(~m[1996]&m[1999]&~m[2000]&m[2001]&m[2002])|(m[1996]&m[1999]&~m[2000]&m[2001]&m[2002])|(~m[1996]&~m[1999]&m[2000]&m[2001]&m[2002])|(m[1996]&~m[1999]&m[2000]&m[2001]&m[2002])|(m[1996]&m[1999]&m[2000]&m[2001]&m[2002]))):InitCond[501];
    m[2003] = run?((((m[2001]&~m[2004]&~m[2005]&~m[2006]&~m[2007])|(~m[2001]&~m[2004]&~m[2005]&m[2006]&~m[2007])|(m[2001]&m[2004]&~m[2005]&m[2006]&~m[2007])|(m[2001]&~m[2004]&m[2005]&m[2006]&~m[2007])|(~m[2001]&m[2004]&~m[2005]&~m[2006]&m[2007])|(~m[2001]&~m[2004]&m[2005]&~m[2006]&m[2007])|(m[2001]&m[2004]&m[2005]&~m[2006]&m[2007])|(~m[2001]&m[2004]&m[2005]&m[2006]&m[2007]))&UnbiasedRNG[246])|((m[2001]&~m[2004]&~m[2005]&m[2006]&~m[2007])|(~m[2001]&~m[2004]&~m[2005]&~m[2006]&m[2007])|(m[2001]&~m[2004]&~m[2005]&~m[2006]&m[2007])|(m[2001]&m[2004]&~m[2005]&~m[2006]&m[2007])|(m[2001]&~m[2004]&m[2005]&~m[2006]&m[2007])|(~m[2001]&~m[2004]&~m[2005]&m[2006]&m[2007])|(m[2001]&~m[2004]&~m[2005]&m[2006]&m[2007])|(~m[2001]&m[2004]&~m[2005]&m[2006]&m[2007])|(m[2001]&m[2004]&~m[2005]&m[2006]&m[2007])|(~m[2001]&~m[2004]&m[2005]&m[2006]&m[2007])|(m[2001]&~m[2004]&m[2005]&m[2006]&m[2007])|(m[2001]&m[2004]&m[2005]&m[2006]&m[2007]))):InitCond[502];
    m[2008] = run?((((m[2006]&~m[2009]&~m[2010]&~m[2011]&~m[2012])|(~m[2006]&~m[2009]&~m[2010]&m[2011]&~m[2012])|(m[2006]&m[2009]&~m[2010]&m[2011]&~m[2012])|(m[2006]&~m[2009]&m[2010]&m[2011]&~m[2012])|(~m[2006]&m[2009]&~m[2010]&~m[2011]&m[2012])|(~m[2006]&~m[2009]&m[2010]&~m[2011]&m[2012])|(m[2006]&m[2009]&m[2010]&~m[2011]&m[2012])|(~m[2006]&m[2009]&m[2010]&m[2011]&m[2012]))&UnbiasedRNG[247])|((m[2006]&~m[2009]&~m[2010]&m[2011]&~m[2012])|(~m[2006]&~m[2009]&~m[2010]&~m[2011]&m[2012])|(m[2006]&~m[2009]&~m[2010]&~m[2011]&m[2012])|(m[2006]&m[2009]&~m[2010]&~m[2011]&m[2012])|(m[2006]&~m[2009]&m[2010]&~m[2011]&m[2012])|(~m[2006]&~m[2009]&~m[2010]&m[2011]&m[2012])|(m[2006]&~m[2009]&~m[2010]&m[2011]&m[2012])|(~m[2006]&m[2009]&~m[2010]&m[2011]&m[2012])|(m[2006]&m[2009]&~m[2010]&m[2011]&m[2012])|(~m[2006]&~m[2009]&m[2010]&m[2011]&m[2012])|(m[2006]&~m[2009]&m[2010]&m[2011]&m[2012])|(m[2006]&m[2009]&m[2010]&m[2011]&m[2012]))):InitCond[503];
    m[2013] = run?((((m[2011]&~m[2014]&~m[2015]&~m[2016]&~m[2017])|(~m[2011]&~m[2014]&~m[2015]&m[2016]&~m[2017])|(m[2011]&m[2014]&~m[2015]&m[2016]&~m[2017])|(m[2011]&~m[2014]&m[2015]&m[2016]&~m[2017])|(~m[2011]&m[2014]&~m[2015]&~m[2016]&m[2017])|(~m[2011]&~m[2014]&m[2015]&~m[2016]&m[2017])|(m[2011]&m[2014]&m[2015]&~m[2016]&m[2017])|(~m[2011]&m[2014]&m[2015]&m[2016]&m[2017]))&UnbiasedRNG[248])|((m[2011]&~m[2014]&~m[2015]&m[2016]&~m[2017])|(~m[2011]&~m[2014]&~m[2015]&~m[2016]&m[2017])|(m[2011]&~m[2014]&~m[2015]&~m[2016]&m[2017])|(m[2011]&m[2014]&~m[2015]&~m[2016]&m[2017])|(m[2011]&~m[2014]&m[2015]&~m[2016]&m[2017])|(~m[2011]&~m[2014]&~m[2015]&m[2016]&m[2017])|(m[2011]&~m[2014]&~m[2015]&m[2016]&m[2017])|(~m[2011]&m[2014]&~m[2015]&m[2016]&m[2017])|(m[2011]&m[2014]&~m[2015]&m[2016]&m[2017])|(~m[2011]&~m[2014]&m[2015]&m[2016]&m[2017])|(m[2011]&~m[2014]&m[2015]&m[2016]&m[2017])|(m[2011]&m[2014]&m[2015]&m[2016]&m[2017]))):InitCond[504];
    m[2018] = run?((((m[2016]&~m[2019]&~m[2020]&~m[2021]&~m[2022])|(~m[2016]&~m[2019]&~m[2020]&m[2021]&~m[2022])|(m[2016]&m[2019]&~m[2020]&m[2021]&~m[2022])|(m[2016]&~m[2019]&m[2020]&m[2021]&~m[2022])|(~m[2016]&m[2019]&~m[2020]&~m[2021]&m[2022])|(~m[2016]&~m[2019]&m[2020]&~m[2021]&m[2022])|(m[2016]&m[2019]&m[2020]&~m[2021]&m[2022])|(~m[2016]&m[2019]&m[2020]&m[2021]&m[2022]))&UnbiasedRNG[249])|((m[2016]&~m[2019]&~m[2020]&m[2021]&~m[2022])|(~m[2016]&~m[2019]&~m[2020]&~m[2021]&m[2022])|(m[2016]&~m[2019]&~m[2020]&~m[2021]&m[2022])|(m[2016]&m[2019]&~m[2020]&~m[2021]&m[2022])|(m[2016]&~m[2019]&m[2020]&~m[2021]&m[2022])|(~m[2016]&~m[2019]&~m[2020]&m[2021]&m[2022])|(m[2016]&~m[2019]&~m[2020]&m[2021]&m[2022])|(~m[2016]&m[2019]&~m[2020]&m[2021]&m[2022])|(m[2016]&m[2019]&~m[2020]&m[2021]&m[2022])|(~m[2016]&~m[2019]&m[2020]&m[2021]&m[2022])|(m[2016]&~m[2019]&m[2020]&m[2021]&m[2022])|(m[2016]&m[2019]&m[2020]&m[2021]&m[2022]))):InitCond[505];
    m[2023] = run?((((m[1992]&~m[2024]&~m[2025]&~m[2026]&~m[2027])|(~m[1992]&~m[2024]&~m[2025]&m[2026]&~m[2027])|(m[1992]&m[2024]&~m[2025]&m[2026]&~m[2027])|(m[1992]&~m[2024]&m[2025]&m[2026]&~m[2027])|(~m[1992]&m[2024]&~m[2025]&~m[2026]&m[2027])|(~m[1992]&~m[2024]&m[2025]&~m[2026]&m[2027])|(m[1992]&m[2024]&m[2025]&~m[2026]&m[2027])|(~m[1992]&m[2024]&m[2025]&m[2026]&m[2027]))&UnbiasedRNG[250])|((m[1992]&~m[2024]&~m[2025]&m[2026]&~m[2027])|(~m[1992]&~m[2024]&~m[2025]&~m[2026]&m[2027])|(m[1992]&~m[2024]&~m[2025]&~m[2026]&m[2027])|(m[1992]&m[2024]&~m[2025]&~m[2026]&m[2027])|(m[1992]&~m[2024]&m[2025]&~m[2026]&m[2027])|(~m[1992]&~m[2024]&~m[2025]&m[2026]&m[2027])|(m[1992]&~m[2024]&~m[2025]&m[2026]&m[2027])|(~m[1992]&m[2024]&~m[2025]&m[2026]&m[2027])|(m[1992]&m[2024]&~m[2025]&m[2026]&m[2027])|(~m[1992]&~m[2024]&m[2025]&m[2026]&m[2027])|(m[1992]&~m[2024]&m[2025]&m[2026]&m[2027])|(m[1992]&m[2024]&m[2025]&m[2026]&m[2027]))):InitCond[506];
    m[2028] = run?((((m[2026]&~m[2029]&~m[2030]&~m[2031]&~m[2032])|(~m[2026]&~m[2029]&~m[2030]&m[2031]&~m[2032])|(m[2026]&m[2029]&~m[2030]&m[2031]&~m[2032])|(m[2026]&~m[2029]&m[2030]&m[2031]&~m[2032])|(~m[2026]&m[2029]&~m[2030]&~m[2031]&m[2032])|(~m[2026]&~m[2029]&m[2030]&~m[2031]&m[2032])|(m[2026]&m[2029]&m[2030]&~m[2031]&m[2032])|(~m[2026]&m[2029]&m[2030]&m[2031]&m[2032]))&UnbiasedRNG[251])|((m[2026]&~m[2029]&~m[2030]&m[2031]&~m[2032])|(~m[2026]&~m[2029]&~m[2030]&~m[2031]&m[2032])|(m[2026]&~m[2029]&~m[2030]&~m[2031]&m[2032])|(m[2026]&m[2029]&~m[2030]&~m[2031]&m[2032])|(m[2026]&~m[2029]&m[2030]&~m[2031]&m[2032])|(~m[2026]&~m[2029]&~m[2030]&m[2031]&m[2032])|(m[2026]&~m[2029]&~m[2030]&m[2031]&m[2032])|(~m[2026]&m[2029]&~m[2030]&m[2031]&m[2032])|(m[2026]&m[2029]&~m[2030]&m[2031]&m[2032])|(~m[2026]&~m[2029]&m[2030]&m[2031]&m[2032])|(m[2026]&~m[2029]&m[2030]&m[2031]&m[2032])|(m[2026]&m[2029]&m[2030]&m[2031]&m[2032]))):InitCond[507];
    m[2033] = run?((((m[2031]&~m[2034]&~m[2035]&~m[2036]&~m[2037])|(~m[2031]&~m[2034]&~m[2035]&m[2036]&~m[2037])|(m[2031]&m[2034]&~m[2035]&m[2036]&~m[2037])|(m[2031]&~m[2034]&m[2035]&m[2036]&~m[2037])|(~m[2031]&m[2034]&~m[2035]&~m[2036]&m[2037])|(~m[2031]&~m[2034]&m[2035]&~m[2036]&m[2037])|(m[2031]&m[2034]&m[2035]&~m[2036]&m[2037])|(~m[2031]&m[2034]&m[2035]&m[2036]&m[2037]))&UnbiasedRNG[252])|((m[2031]&~m[2034]&~m[2035]&m[2036]&~m[2037])|(~m[2031]&~m[2034]&~m[2035]&~m[2036]&m[2037])|(m[2031]&~m[2034]&~m[2035]&~m[2036]&m[2037])|(m[2031]&m[2034]&~m[2035]&~m[2036]&m[2037])|(m[2031]&~m[2034]&m[2035]&~m[2036]&m[2037])|(~m[2031]&~m[2034]&~m[2035]&m[2036]&m[2037])|(m[2031]&~m[2034]&~m[2035]&m[2036]&m[2037])|(~m[2031]&m[2034]&~m[2035]&m[2036]&m[2037])|(m[2031]&m[2034]&~m[2035]&m[2036]&m[2037])|(~m[2031]&~m[2034]&m[2035]&m[2036]&m[2037])|(m[2031]&~m[2034]&m[2035]&m[2036]&m[2037])|(m[2031]&m[2034]&m[2035]&m[2036]&m[2037]))):InitCond[508];
    m[2038] = run?((((m[2036]&~m[2039]&~m[2040]&~m[2041]&~m[2042])|(~m[2036]&~m[2039]&~m[2040]&m[2041]&~m[2042])|(m[2036]&m[2039]&~m[2040]&m[2041]&~m[2042])|(m[2036]&~m[2039]&m[2040]&m[2041]&~m[2042])|(~m[2036]&m[2039]&~m[2040]&~m[2041]&m[2042])|(~m[2036]&~m[2039]&m[2040]&~m[2041]&m[2042])|(m[2036]&m[2039]&m[2040]&~m[2041]&m[2042])|(~m[2036]&m[2039]&m[2040]&m[2041]&m[2042]))&UnbiasedRNG[253])|((m[2036]&~m[2039]&~m[2040]&m[2041]&~m[2042])|(~m[2036]&~m[2039]&~m[2040]&~m[2041]&m[2042])|(m[2036]&~m[2039]&~m[2040]&~m[2041]&m[2042])|(m[2036]&m[2039]&~m[2040]&~m[2041]&m[2042])|(m[2036]&~m[2039]&m[2040]&~m[2041]&m[2042])|(~m[2036]&~m[2039]&~m[2040]&m[2041]&m[2042])|(m[2036]&~m[2039]&~m[2040]&m[2041]&m[2042])|(~m[2036]&m[2039]&~m[2040]&m[2041]&m[2042])|(m[2036]&m[2039]&~m[2040]&m[2041]&m[2042])|(~m[2036]&~m[2039]&m[2040]&m[2041]&m[2042])|(m[2036]&~m[2039]&m[2040]&m[2041]&m[2042])|(m[2036]&m[2039]&m[2040]&m[2041]&m[2042]))):InitCond[509];
    m[2043] = run?((((m[2041]&~m[2044]&~m[2045]&~m[2046]&~m[2047])|(~m[2041]&~m[2044]&~m[2045]&m[2046]&~m[2047])|(m[2041]&m[2044]&~m[2045]&m[2046]&~m[2047])|(m[2041]&~m[2044]&m[2045]&m[2046]&~m[2047])|(~m[2041]&m[2044]&~m[2045]&~m[2046]&m[2047])|(~m[2041]&~m[2044]&m[2045]&~m[2046]&m[2047])|(m[2041]&m[2044]&m[2045]&~m[2046]&m[2047])|(~m[2041]&m[2044]&m[2045]&m[2046]&m[2047]))&UnbiasedRNG[254])|((m[2041]&~m[2044]&~m[2045]&m[2046]&~m[2047])|(~m[2041]&~m[2044]&~m[2045]&~m[2046]&m[2047])|(m[2041]&~m[2044]&~m[2045]&~m[2046]&m[2047])|(m[2041]&m[2044]&~m[2045]&~m[2046]&m[2047])|(m[2041]&~m[2044]&m[2045]&~m[2046]&m[2047])|(~m[2041]&~m[2044]&~m[2045]&m[2046]&m[2047])|(m[2041]&~m[2044]&~m[2045]&m[2046]&m[2047])|(~m[2041]&m[2044]&~m[2045]&m[2046]&m[2047])|(m[2041]&m[2044]&~m[2045]&m[2046]&m[2047])|(~m[2041]&~m[2044]&m[2045]&m[2046]&m[2047])|(m[2041]&~m[2044]&m[2045]&m[2046]&m[2047])|(m[2041]&m[2044]&m[2045]&m[2046]&m[2047]))):InitCond[510];
    m[2048] = run?((((m[2046]&~m[2049]&~m[2050]&~m[2051]&~m[2052])|(~m[2046]&~m[2049]&~m[2050]&m[2051]&~m[2052])|(m[2046]&m[2049]&~m[2050]&m[2051]&~m[2052])|(m[2046]&~m[2049]&m[2050]&m[2051]&~m[2052])|(~m[2046]&m[2049]&~m[2050]&~m[2051]&m[2052])|(~m[2046]&~m[2049]&m[2050]&~m[2051]&m[2052])|(m[2046]&m[2049]&m[2050]&~m[2051]&m[2052])|(~m[2046]&m[2049]&m[2050]&m[2051]&m[2052]))&UnbiasedRNG[255])|((m[2046]&~m[2049]&~m[2050]&m[2051]&~m[2052])|(~m[2046]&~m[2049]&~m[2050]&~m[2051]&m[2052])|(m[2046]&~m[2049]&~m[2050]&~m[2051]&m[2052])|(m[2046]&m[2049]&~m[2050]&~m[2051]&m[2052])|(m[2046]&~m[2049]&m[2050]&~m[2051]&m[2052])|(~m[2046]&~m[2049]&~m[2050]&m[2051]&m[2052])|(m[2046]&~m[2049]&~m[2050]&m[2051]&m[2052])|(~m[2046]&m[2049]&~m[2050]&m[2051]&m[2052])|(m[2046]&m[2049]&~m[2050]&m[2051]&m[2052])|(~m[2046]&~m[2049]&m[2050]&m[2051]&m[2052])|(m[2046]&~m[2049]&m[2050]&m[2051]&m[2052])|(m[2046]&m[2049]&m[2050]&m[2051]&m[2052]))):InitCond[511];
    m[2053] = run?((((m[2027]&~m[2054]&~m[2055]&~m[2056]&~m[2057])|(~m[2027]&~m[2054]&~m[2055]&m[2056]&~m[2057])|(m[2027]&m[2054]&~m[2055]&m[2056]&~m[2057])|(m[2027]&~m[2054]&m[2055]&m[2056]&~m[2057])|(~m[2027]&m[2054]&~m[2055]&~m[2056]&m[2057])|(~m[2027]&~m[2054]&m[2055]&~m[2056]&m[2057])|(m[2027]&m[2054]&m[2055]&~m[2056]&m[2057])|(~m[2027]&m[2054]&m[2055]&m[2056]&m[2057]))&UnbiasedRNG[256])|((m[2027]&~m[2054]&~m[2055]&m[2056]&~m[2057])|(~m[2027]&~m[2054]&~m[2055]&~m[2056]&m[2057])|(m[2027]&~m[2054]&~m[2055]&~m[2056]&m[2057])|(m[2027]&m[2054]&~m[2055]&~m[2056]&m[2057])|(m[2027]&~m[2054]&m[2055]&~m[2056]&m[2057])|(~m[2027]&~m[2054]&~m[2055]&m[2056]&m[2057])|(m[2027]&~m[2054]&~m[2055]&m[2056]&m[2057])|(~m[2027]&m[2054]&~m[2055]&m[2056]&m[2057])|(m[2027]&m[2054]&~m[2055]&m[2056]&m[2057])|(~m[2027]&~m[2054]&m[2055]&m[2056]&m[2057])|(m[2027]&~m[2054]&m[2055]&m[2056]&m[2057])|(m[2027]&m[2054]&m[2055]&m[2056]&m[2057]))):InitCond[512];
    m[2058] = run?((((m[2056]&~m[2059]&~m[2060]&~m[2061]&~m[2062])|(~m[2056]&~m[2059]&~m[2060]&m[2061]&~m[2062])|(m[2056]&m[2059]&~m[2060]&m[2061]&~m[2062])|(m[2056]&~m[2059]&m[2060]&m[2061]&~m[2062])|(~m[2056]&m[2059]&~m[2060]&~m[2061]&m[2062])|(~m[2056]&~m[2059]&m[2060]&~m[2061]&m[2062])|(m[2056]&m[2059]&m[2060]&~m[2061]&m[2062])|(~m[2056]&m[2059]&m[2060]&m[2061]&m[2062]))&UnbiasedRNG[257])|((m[2056]&~m[2059]&~m[2060]&m[2061]&~m[2062])|(~m[2056]&~m[2059]&~m[2060]&~m[2061]&m[2062])|(m[2056]&~m[2059]&~m[2060]&~m[2061]&m[2062])|(m[2056]&m[2059]&~m[2060]&~m[2061]&m[2062])|(m[2056]&~m[2059]&m[2060]&~m[2061]&m[2062])|(~m[2056]&~m[2059]&~m[2060]&m[2061]&m[2062])|(m[2056]&~m[2059]&~m[2060]&m[2061]&m[2062])|(~m[2056]&m[2059]&~m[2060]&m[2061]&m[2062])|(m[2056]&m[2059]&~m[2060]&m[2061]&m[2062])|(~m[2056]&~m[2059]&m[2060]&m[2061]&m[2062])|(m[2056]&~m[2059]&m[2060]&m[2061]&m[2062])|(m[2056]&m[2059]&m[2060]&m[2061]&m[2062]))):InitCond[513];
    m[2063] = run?((((m[2061]&~m[2064]&~m[2065]&~m[2066]&~m[2067])|(~m[2061]&~m[2064]&~m[2065]&m[2066]&~m[2067])|(m[2061]&m[2064]&~m[2065]&m[2066]&~m[2067])|(m[2061]&~m[2064]&m[2065]&m[2066]&~m[2067])|(~m[2061]&m[2064]&~m[2065]&~m[2066]&m[2067])|(~m[2061]&~m[2064]&m[2065]&~m[2066]&m[2067])|(m[2061]&m[2064]&m[2065]&~m[2066]&m[2067])|(~m[2061]&m[2064]&m[2065]&m[2066]&m[2067]))&UnbiasedRNG[258])|((m[2061]&~m[2064]&~m[2065]&m[2066]&~m[2067])|(~m[2061]&~m[2064]&~m[2065]&~m[2066]&m[2067])|(m[2061]&~m[2064]&~m[2065]&~m[2066]&m[2067])|(m[2061]&m[2064]&~m[2065]&~m[2066]&m[2067])|(m[2061]&~m[2064]&m[2065]&~m[2066]&m[2067])|(~m[2061]&~m[2064]&~m[2065]&m[2066]&m[2067])|(m[2061]&~m[2064]&~m[2065]&m[2066]&m[2067])|(~m[2061]&m[2064]&~m[2065]&m[2066]&m[2067])|(m[2061]&m[2064]&~m[2065]&m[2066]&m[2067])|(~m[2061]&~m[2064]&m[2065]&m[2066]&m[2067])|(m[2061]&~m[2064]&m[2065]&m[2066]&m[2067])|(m[2061]&m[2064]&m[2065]&m[2066]&m[2067]))):InitCond[514];
    m[2068] = run?((((m[2066]&~m[2069]&~m[2070]&~m[2071]&~m[2072])|(~m[2066]&~m[2069]&~m[2070]&m[2071]&~m[2072])|(m[2066]&m[2069]&~m[2070]&m[2071]&~m[2072])|(m[2066]&~m[2069]&m[2070]&m[2071]&~m[2072])|(~m[2066]&m[2069]&~m[2070]&~m[2071]&m[2072])|(~m[2066]&~m[2069]&m[2070]&~m[2071]&m[2072])|(m[2066]&m[2069]&m[2070]&~m[2071]&m[2072])|(~m[2066]&m[2069]&m[2070]&m[2071]&m[2072]))&UnbiasedRNG[259])|((m[2066]&~m[2069]&~m[2070]&m[2071]&~m[2072])|(~m[2066]&~m[2069]&~m[2070]&~m[2071]&m[2072])|(m[2066]&~m[2069]&~m[2070]&~m[2071]&m[2072])|(m[2066]&m[2069]&~m[2070]&~m[2071]&m[2072])|(m[2066]&~m[2069]&m[2070]&~m[2071]&m[2072])|(~m[2066]&~m[2069]&~m[2070]&m[2071]&m[2072])|(m[2066]&~m[2069]&~m[2070]&m[2071]&m[2072])|(~m[2066]&m[2069]&~m[2070]&m[2071]&m[2072])|(m[2066]&m[2069]&~m[2070]&m[2071]&m[2072])|(~m[2066]&~m[2069]&m[2070]&m[2071]&m[2072])|(m[2066]&~m[2069]&m[2070]&m[2071]&m[2072])|(m[2066]&m[2069]&m[2070]&m[2071]&m[2072]))):InitCond[515];
    m[2073] = run?((((m[2071]&~m[2074]&~m[2075]&~m[2076]&~m[2077])|(~m[2071]&~m[2074]&~m[2075]&m[2076]&~m[2077])|(m[2071]&m[2074]&~m[2075]&m[2076]&~m[2077])|(m[2071]&~m[2074]&m[2075]&m[2076]&~m[2077])|(~m[2071]&m[2074]&~m[2075]&~m[2076]&m[2077])|(~m[2071]&~m[2074]&m[2075]&~m[2076]&m[2077])|(m[2071]&m[2074]&m[2075]&~m[2076]&m[2077])|(~m[2071]&m[2074]&m[2075]&m[2076]&m[2077]))&UnbiasedRNG[260])|((m[2071]&~m[2074]&~m[2075]&m[2076]&~m[2077])|(~m[2071]&~m[2074]&~m[2075]&~m[2076]&m[2077])|(m[2071]&~m[2074]&~m[2075]&~m[2076]&m[2077])|(m[2071]&m[2074]&~m[2075]&~m[2076]&m[2077])|(m[2071]&~m[2074]&m[2075]&~m[2076]&m[2077])|(~m[2071]&~m[2074]&~m[2075]&m[2076]&m[2077])|(m[2071]&~m[2074]&~m[2075]&m[2076]&m[2077])|(~m[2071]&m[2074]&~m[2075]&m[2076]&m[2077])|(m[2071]&m[2074]&~m[2075]&m[2076]&m[2077])|(~m[2071]&~m[2074]&m[2075]&m[2076]&m[2077])|(m[2071]&~m[2074]&m[2075]&m[2076]&m[2077])|(m[2071]&m[2074]&m[2075]&m[2076]&m[2077]))):InitCond[516];
    m[2078] = run?((((m[2057]&~m[2079]&~m[2080]&~m[2081]&~m[2082])|(~m[2057]&~m[2079]&~m[2080]&m[2081]&~m[2082])|(m[2057]&m[2079]&~m[2080]&m[2081]&~m[2082])|(m[2057]&~m[2079]&m[2080]&m[2081]&~m[2082])|(~m[2057]&m[2079]&~m[2080]&~m[2081]&m[2082])|(~m[2057]&~m[2079]&m[2080]&~m[2081]&m[2082])|(m[2057]&m[2079]&m[2080]&~m[2081]&m[2082])|(~m[2057]&m[2079]&m[2080]&m[2081]&m[2082]))&UnbiasedRNG[261])|((m[2057]&~m[2079]&~m[2080]&m[2081]&~m[2082])|(~m[2057]&~m[2079]&~m[2080]&~m[2081]&m[2082])|(m[2057]&~m[2079]&~m[2080]&~m[2081]&m[2082])|(m[2057]&m[2079]&~m[2080]&~m[2081]&m[2082])|(m[2057]&~m[2079]&m[2080]&~m[2081]&m[2082])|(~m[2057]&~m[2079]&~m[2080]&m[2081]&m[2082])|(m[2057]&~m[2079]&~m[2080]&m[2081]&m[2082])|(~m[2057]&m[2079]&~m[2080]&m[2081]&m[2082])|(m[2057]&m[2079]&~m[2080]&m[2081]&m[2082])|(~m[2057]&~m[2079]&m[2080]&m[2081]&m[2082])|(m[2057]&~m[2079]&m[2080]&m[2081]&m[2082])|(m[2057]&m[2079]&m[2080]&m[2081]&m[2082]))):InitCond[517];
    m[2083] = run?((((m[2081]&~m[2084]&~m[2085]&~m[2086]&~m[2087])|(~m[2081]&~m[2084]&~m[2085]&m[2086]&~m[2087])|(m[2081]&m[2084]&~m[2085]&m[2086]&~m[2087])|(m[2081]&~m[2084]&m[2085]&m[2086]&~m[2087])|(~m[2081]&m[2084]&~m[2085]&~m[2086]&m[2087])|(~m[2081]&~m[2084]&m[2085]&~m[2086]&m[2087])|(m[2081]&m[2084]&m[2085]&~m[2086]&m[2087])|(~m[2081]&m[2084]&m[2085]&m[2086]&m[2087]))&UnbiasedRNG[262])|((m[2081]&~m[2084]&~m[2085]&m[2086]&~m[2087])|(~m[2081]&~m[2084]&~m[2085]&~m[2086]&m[2087])|(m[2081]&~m[2084]&~m[2085]&~m[2086]&m[2087])|(m[2081]&m[2084]&~m[2085]&~m[2086]&m[2087])|(m[2081]&~m[2084]&m[2085]&~m[2086]&m[2087])|(~m[2081]&~m[2084]&~m[2085]&m[2086]&m[2087])|(m[2081]&~m[2084]&~m[2085]&m[2086]&m[2087])|(~m[2081]&m[2084]&~m[2085]&m[2086]&m[2087])|(m[2081]&m[2084]&~m[2085]&m[2086]&m[2087])|(~m[2081]&~m[2084]&m[2085]&m[2086]&m[2087])|(m[2081]&~m[2084]&m[2085]&m[2086]&m[2087])|(m[2081]&m[2084]&m[2085]&m[2086]&m[2087]))):InitCond[518];
    m[2088] = run?((((m[2086]&~m[2089]&~m[2090]&~m[2091]&~m[2092])|(~m[2086]&~m[2089]&~m[2090]&m[2091]&~m[2092])|(m[2086]&m[2089]&~m[2090]&m[2091]&~m[2092])|(m[2086]&~m[2089]&m[2090]&m[2091]&~m[2092])|(~m[2086]&m[2089]&~m[2090]&~m[2091]&m[2092])|(~m[2086]&~m[2089]&m[2090]&~m[2091]&m[2092])|(m[2086]&m[2089]&m[2090]&~m[2091]&m[2092])|(~m[2086]&m[2089]&m[2090]&m[2091]&m[2092]))&UnbiasedRNG[263])|((m[2086]&~m[2089]&~m[2090]&m[2091]&~m[2092])|(~m[2086]&~m[2089]&~m[2090]&~m[2091]&m[2092])|(m[2086]&~m[2089]&~m[2090]&~m[2091]&m[2092])|(m[2086]&m[2089]&~m[2090]&~m[2091]&m[2092])|(m[2086]&~m[2089]&m[2090]&~m[2091]&m[2092])|(~m[2086]&~m[2089]&~m[2090]&m[2091]&m[2092])|(m[2086]&~m[2089]&~m[2090]&m[2091]&m[2092])|(~m[2086]&m[2089]&~m[2090]&m[2091]&m[2092])|(m[2086]&m[2089]&~m[2090]&m[2091]&m[2092])|(~m[2086]&~m[2089]&m[2090]&m[2091]&m[2092])|(m[2086]&~m[2089]&m[2090]&m[2091]&m[2092])|(m[2086]&m[2089]&m[2090]&m[2091]&m[2092]))):InitCond[519];
    m[2093] = run?((((m[2091]&~m[2094]&~m[2095]&~m[2096]&~m[2097])|(~m[2091]&~m[2094]&~m[2095]&m[2096]&~m[2097])|(m[2091]&m[2094]&~m[2095]&m[2096]&~m[2097])|(m[2091]&~m[2094]&m[2095]&m[2096]&~m[2097])|(~m[2091]&m[2094]&~m[2095]&~m[2096]&m[2097])|(~m[2091]&~m[2094]&m[2095]&~m[2096]&m[2097])|(m[2091]&m[2094]&m[2095]&~m[2096]&m[2097])|(~m[2091]&m[2094]&m[2095]&m[2096]&m[2097]))&UnbiasedRNG[264])|((m[2091]&~m[2094]&~m[2095]&m[2096]&~m[2097])|(~m[2091]&~m[2094]&~m[2095]&~m[2096]&m[2097])|(m[2091]&~m[2094]&~m[2095]&~m[2096]&m[2097])|(m[2091]&m[2094]&~m[2095]&~m[2096]&m[2097])|(m[2091]&~m[2094]&m[2095]&~m[2096]&m[2097])|(~m[2091]&~m[2094]&~m[2095]&m[2096]&m[2097])|(m[2091]&~m[2094]&~m[2095]&m[2096]&m[2097])|(~m[2091]&m[2094]&~m[2095]&m[2096]&m[2097])|(m[2091]&m[2094]&~m[2095]&m[2096]&m[2097])|(~m[2091]&~m[2094]&m[2095]&m[2096]&m[2097])|(m[2091]&~m[2094]&m[2095]&m[2096]&m[2097])|(m[2091]&m[2094]&m[2095]&m[2096]&m[2097]))):InitCond[520];
    m[2098] = run?((((m[2082]&~m[2099]&~m[2100]&~m[2101]&~m[2102])|(~m[2082]&~m[2099]&~m[2100]&m[2101]&~m[2102])|(m[2082]&m[2099]&~m[2100]&m[2101]&~m[2102])|(m[2082]&~m[2099]&m[2100]&m[2101]&~m[2102])|(~m[2082]&m[2099]&~m[2100]&~m[2101]&m[2102])|(~m[2082]&~m[2099]&m[2100]&~m[2101]&m[2102])|(m[2082]&m[2099]&m[2100]&~m[2101]&m[2102])|(~m[2082]&m[2099]&m[2100]&m[2101]&m[2102]))&UnbiasedRNG[265])|((m[2082]&~m[2099]&~m[2100]&m[2101]&~m[2102])|(~m[2082]&~m[2099]&~m[2100]&~m[2101]&m[2102])|(m[2082]&~m[2099]&~m[2100]&~m[2101]&m[2102])|(m[2082]&m[2099]&~m[2100]&~m[2101]&m[2102])|(m[2082]&~m[2099]&m[2100]&~m[2101]&m[2102])|(~m[2082]&~m[2099]&~m[2100]&m[2101]&m[2102])|(m[2082]&~m[2099]&~m[2100]&m[2101]&m[2102])|(~m[2082]&m[2099]&~m[2100]&m[2101]&m[2102])|(m[2082]&m[2099]&~m[2100]&m[2101]&m[2102])|(~m[2082]&~m[2099]&m[2100]&m[2101]&m[2102])|(m[2082]&~m[2099]&m[2100]&m[2101]&m[2102])|(m[2082]&m[2099]&m[2100]&m[2101]&m[2102]))):InitCond[521];
    m[2103] = run?((((m[2101]&~m[2104]&~m[2105]&~m[2106]&~m[2107])|(~m[2101]&~m[2104]&~m[2105]&m[2106]&~m[2107])|(m[2101]&m[2104]&~m[2105]&m[2106]&~m[2107])|(m[2101]&~m[2104]&m[2105]&m[2106]&~m[2107])|(~m[2101]&m[2104]&~m[2105]&~m[2106]&m[2107])|(~m[2101]&~m[2104]&m[2105]&~m[2106]&m[2107])|(m[2101]&m[2104]&m[2105]&~m[2106]&m[2107])|(~m[2101]&m[2104]&m[2105]&m[2106]&m[2107]))&UnbiasedRNG[266])|((m[2101]&~m[2104]&~m[2105]&m[2106]&~m[2107])|(~m[2101]&~m[2104]&~m[2105]&~m[2106]&m[2107])|(m[2101]&~m[2104]&~m[2105]&~m[2106]&m[2107])|(m[2101]&m[2104]&~m[2105]&~m[2106]&m[2107])|(m[2101]&~m[2104]&m[2105]&~m[2106]&m[2107])|(~m[2101]&~m[2104]&~m[2105]&m[2106]&m[2107])|(m[2101]&~m[2104]&~m[2105]&m[2106]&m[2107])|(~m[2101]&m[2104]&~m[2105]&m[2106]&m[2107])|(m[2101]&m[2104]&~m[2105]&m[2106]&m[2107])|(~m[2101]&~m[2104]&m[2105]&m[2106]&m[2107])|(m[2101]&~m[2104]&m[2105]&m[2106]&m[2107])|(m[2101]&m[2104]&m[2105]&m[2106]&m[2107]))):InitCond[522];
    m[2108] = run?((((m[2106]&~m[2109]&~m[2110]&~m[2111]&~m[2112])|(~m[2106]&~m[2109]&~m[2110]&m[2111]&~m[2112])|(m[2106]&m[2109]&~m[2110]&m[2111]&~m[2112])|(m[2106]&~m[2109]&m[2110]&m[2111]&~m[2112])|(~m[2106]&m[2109]&~m[2110]&~m[2111]&m[2112])|(~m[2106]&~m[2109]&m[2110]&~m[2111]&m[2112])|(m[2106]&m[2109]&m[2110]&~m[2111]&m[2112])|(~m[2106]&m[2109]&m[2110]&m[2111]&m[2112]))&UnbiasedRNG[267])|((m[2106]&~m[2109]&~m[2110]&m[2111]&~m[2112])|(~m[2106]&~m[2109]&~m[2110]&~m[2111]&m[2112])|(m[2106]&~m[2109]&~m[2110]&~m[2111]&m[2112])|(m[2106]&m[2109]&~m[2110]&~m[2111]&m[2112])|(m[2106]&~m[2109]&m[2110]&~m[2111]&m[2112])|(~m[2106]&~m[2109]&~m[2110]&m[2111]&m[2112])|(m[2106]&~m[2109]&~m[2110]&m[2111]&m[2112])|(~m[2106]&m[2109]&~m[2110]&m[2111]&m[2112])|(m[2106]&m[2109]&~m[2110]&m[2111]&m[2112])|(~m[2106]&~m[2109]&m[2110]&m[2111]&m[2112])|(m[2106]&~m[2109]&m[2110]&m[2111]&m[2112])|(m[2106]&m[2109]&m[2110]&m[2111]&m[2112]))):InitCond[523];
    m[2113] = run?((((m[2102]&~m[2114]&~m[2115]&~m[2116]&~m[2117])|(~m[2102]&~m[2114]&~m[2115]&m[2116]&~m[2117])|(m[2102]&m[2114]&~m[2115]&m[2116]&~m[2117])|(m[2102]&~m[2114]&m[2115]&m[2116]&~m[2117])|(~m[2102]&m[2114]&~m[2115]&~m[2116]&m[2117])|(~m[2102]&~m[2114]&m[2115]&~m[2116]&m[2117])|(m[2102]&m[2114]&m[2115]&~m[2116]&m[2117])|(~m[2102]&m[2114]&m[2115]&m[2116]&m[2117]))&UnbiasedRNG[268])|((m[2102]&~m[2114]&~m[2115]&m[2116]&~m[2117])|(~m[2102]&~m[2114]&~m[2115]&~m[2116]&m[2117])|(m[2102]&~m[2114]&~m[2115]&~m[2116]&m[2117])|(m[2102]&m[2114]&~m[2115]&~m[2116]&m[2117])|(m[2102]&~m[2114]&m[2115]&~m[2116]&m[2117])|(~m[2102]&~m[2114]&~m[2115]&m[2116]&m[2117])|(m[2102]&~m[2114]&~m[2115]&m[2116]&m[2117])|(~m[2102]&m[2114]&~m[2115]&m[2116]&m[2117])|(m[2102]&m[2114]&~m[2115]&m[2116]&m[2117])|(~m[2102]&~m[2114]&m[2115]&m[2116]&m[2117])|(m[2102]&~m[2114]&m[2115]&m[2116]&m[2117])|(m[2102]&m[2114]&m[2115]&m[2116]&m[2117]))):InitCond[524];
    m[2118] = run?((((m[2116]&~m[2119]&~m[2120]&~m[2121]&~m[2122])|(~m[2116]&~m[2119]&~m[2120]&m[2121]&~m[2122])|(m[2116]&m[2119]&~m[2120]&m[2121]&~m[2122])|(m[2116]&~m[2119]&m[2120]&m[2121]&~m[2122])|(~m[2116]&m[2119]&~m[2120]&~m[2121]&m[2122])|(~m[2116]&~m[2119]&m[2120]&~m[2121]&m[2122])|(m[2116]&m[2119]&m[2120]&~m[2121]&m[2122])|(~m[2116]&m[2119]&m[2120]&m[2121]&m[2122]))&UnbiasedRNG[269])|((m[2116]&~m[2119]&~m[2120]&m[2121]&~m[2122])|(~m[2116]&~m[2119]&~m[2120]&~m[2121]&m[2122])|(m[2116]&~m[2119]&~m[2120]&~m[2121]&m[2122])|(m[2116]&m[2119]&~m[2120]&~m[2121]&m[2122])|(m[2116]&~m[2119]&m[2120]&~m[2121]&m[2122])|(~m[2116]&~m[2119]&~m[2120]&m[2121]&m[2122])|(m[2116]&~m[2119]&~m[2120]&m[2121]&m[2122])|(~m[2116]&m[2119]&~m[2120]&m[2121]&m[2122])|(m[2116]&m[2119]&~m[2120]&m[2121]&m[2122])|(~m[2116]&~m[2119]&m[2120]&m[2121]&m[2122])|(m[2116]&~m[2119]&m[2120]&m[2121]&m[2122])|(m[2116]&m[2119]&m[2120]&m[2121]&m[2122]))):InitCond[525];
    m[2123] = run?((((m[2117]&~m[2124]&~m[2125]&~m[2126]&~m[2127])|(~m[2117]&~m[2124]&~m[2125]&m[2126]&~m[2127])|(m[2117]&m[2124]&~m[2125]&m[2126]&~m[2127])|(m[2117]&~m[2124]&m[2125]&m[2126]&~m[2127])|(~m[2117]&m[2124]&~m[2125]&~m[2126]&m[2127])|(~m[2117]&~m[2124]&m[2125]&~m[2126]&m[2127])|(m[2117]&m[2124]&m[2125]&~m[2126]&m[2127])|(~m[2117]&m[2124]&m[2125]&m[2126]&m[2127]))&UnbiasedRNG[270])|((m[2117]&~m[2124]&~m[2125]&m[2126]&~m[2127])|(~m[2117]&~m[2124]&~m[2125]&~m[2126]&m[2127])|(m[2117]&~m[2124]&~m[2125]&~m[2126]&m[2127])|(m[2117]&m[2124]&~m[2125]&~m[2126]&m[2127])|(m[2117]&~m[2124]&m[2125]&~m[2126]&m[2127])|(~m[2117]&~m[2124]&~m[2125]&m[2126]&m[2127])|(m[2117]&~m[2124]&~m[2125]&m[2126]&m[2127])|(~m[2117]&m[2124]&~m[2125]&m[2126]&m[2127])|(m[2117]&m[2124]&~m[2125]&m[2126]&m[2127])|(~m[2117]&~m[2124]&m[2125]&m[2126]&m[2127])|(m[2117]&~m[2124]&m[2125]&m[2126]&m[2127])|(m[2117]&m[2124]&m[2125]&m[2126]&m[2127]))):InitCond[526];
end

always @(posedge color1_clk) begin
    m[32] = run?((((m[0]&m[160]&~m[161]&~m[162]&~m[163])|(m[0]&~m[160]&m[161]&~m[162]&~m[163])|(~m[0]&m[160]&m[161]&~m[162]&~m[163])|(m[0]&~m[160]&~m[161]&m[162]&~m[163])|(~m[0]&m[160]&~m[161]&m[162]&~m[163])|(~m[0]&~m[160]&m[161]&m[162]&~m[163])|(m[0]&~m[160]&~m[161]&~m[162]&m[163])|(~m[0]&m[160]&~m[161]&~m[162]&m[163])|(~m[0]&~m[160]&m[161]&~m[162]&m[163])|(~m[0]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[256])|(((m[0]&m[160]&m[161]&~m[162]&~m[163])|(m[0]&m[160]&~m[161]&m[162]&~m[163])|(m[0]&~m[160]&m[161]&m[162]&~m[163])|(~m[0]&m[160]&m[161]&m[162]&~m[163])|(m[0]&m[160]&~m[161]&~m[162]&m[163])|(m[0]&~m[160]&m[161]&~m[162]&m[163])|(~m[0]&m[160]&m[161]&~m[162]&m[163])|(m[0]&~m[160]&~m[161]&m[162]&m[163])|(~m[0]&m[160]&~m[161]&m[162]&m[163])|(~m[0]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[256])|((m[0]&m[160]&m[161]&m[162]&~m[163])|(m[0]&m[160]&m[161]&~m[162]&m[163])|(m[0]&m[160]&~m[161]&m[162]&m[163])|(m[0]&~m[160]&m[161]&m[162]&m[163])|(~m[0]&m[160]&m[161]&m[162]&m[163])|(m[0]&m[160]&m[161]&m[162]&m[163]))):InitCond[527];
    m[33] = run?((((m[0]&m[164]&~m[165]&~m[166]&~m[167])|(m[0]&~m[164]&m[165]&~m[166]&~m[167])|(~m[0]&m[164]&m[165]&~m[166]&~m[167])|(m[0]&~m[164]&~m[165]&m[166]&~m[167])|(~m[0]&m[164]&~m[165]&m[166]&~m[167])|(~m[0]&~m[164]&m[165]&m[166]&~m[167])|(m[0]&~m[164]&~m[165]&~m[166]&m[167])|(~m[0]&m[164]&~m[165]&~m[166]&m[167])|(~m[0]&~m[164]&m[165]&~m[166]&m[167])|(~m[0]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[257])|(((m[0]&m[164]&m[165]&~m[166]&~m[167])|(m[0]&m[164]&~m[165]&m[166]&~m[167])|(m[0]&~m[164]&m[165]&m[166]&~m[167])|(~m[0]&m[164]&m[165]&m[166]&~m[167])|(m[0]&m[164]&~m[165]&~m[166]&m[167])|(m[0]&~m[164]&m[165]&~m[166]&m[167])|(~m[0]&m[164]&m[165]&~m[166]&m[167])|(m[0]&~m[164]&~m[165]&m[166]&m[167])|(~m[0]&m[164]&~m[165]&m[166]&m[167])|(~m[0]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[257])|((m[0]&m[164]&m[165]&m[166]&~m[167])|(m[0]&m[164]&m[165]&~m[166]&m[167])|(m[0]&m[164]&~m[165]&m[166]&m[167])|(m[0]&~m[164]&m[165]&m[166]&m[167])|(~m[0]&m[164]&m[165]&m[166]&m[167])|(m[0]&m[164]&m[165]&m[166]&m[167]))):InitCond[528];
    m[34] = run?((((m[0]&m[168]&~m[169]&~m[170]&~m[171])|(m[0]&~m[168]&m[169]&~m[170]&~m[171])|(~m[0]&m[168]&m[169]&~m[170]&~m[171])|(m[0]&~m[168]&~m[169]&m[170]&~m[171])|(~m[0]&m[168]&~m[169]&m[170]&~m[171])|(~m[0]&~m[168]&m[169]&m[170]&~m[171])|(m[0]&~m[168]&~m[169]&~m[170]&m[171])|(~m[0]&m[168]&~m[169]&~m[170]&m[171])|(~m[0]&~m[168]&m[169]&~m[170]&m[171])|(~m[0]&~m[168]&~m[169]&m[170]&m[171]))&BiasedRNG[258])|(((m[0]&m[168]&m[169]&~m[170]&~m[171])|(m[0]&m[168]&~m[169]&m[170]&~m[171])|(m[0]&~m[168]&m[169]&m[170]&~m[171])|(~m[0]&m[168]&m[169]&m[170]&~m[171])|(m[0]&m[168]&~m[169]&~m[170]&m[171])|(m[0]&~m[168]&m[169]&~m[170]&m[171])|(~m[0]&m[168]&m[169]&~m[170]&m[171])|(m[0]&~m[168]&~m[169]&m[170]&m[171])|(~m[0]&m[168]&~m[169]&m[170]&m[171])|(~m[0]&~m[168]&m[169]&m[170]&m[171]))&~BiasedRNG[258])|((m[0]&m[168]&m[169]&m[170]&~m[171])|(m[0]&m[168]&m[169]&~m[170]&m[171])|(m[0]&m[168]&~m[169]&m[170]&m[171])|(m[0]&~m[168]&m[169]&m[170]&m[171])|(~m[0]&m[168]&m[169]&m[170]&m[171])|(m[0]&m[168]&m[169]&m[170]&m[171]))):InitCond[529];
    m[35] = run?((((m[0]&m[172]&~m[173]&~m[174]&~m[175])|(m[0]&~m[172]&m[173]&~m[174]&~m[175])|(~m[0]&m[172]&m[173]&~m[174]&~m[175])|(m[0]&~m[172]&~m[173]&m[174]&~m[175])|(~m[0]&m[172]&~m[173]&m[174]&~m[175])|(~m[0]&~m[172]&m[173]&m[174]&~m[175])|(m[0]&~m[172]&~m[173]&~m[174]&m[175])|(~m[0]&m[172]&~m[173]&~m[174]&m[175])|(~m[0]&~m[172]&m[173]&~m[174]&m[175])|(~m[0]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[259])|(((m[0]&m[172]&m[173]&~m[174]&~m[175])|(m[0]&m[172]&~m[173]&m[174]&~m[175])|(m[0]&~m[172]&m[173]&m[174]&~m[175])|(~m[0]&m[172]&m[173]&m[174]&~m[175])|(m[0]&m[172]&~m[173]&~m[174]&m[175])|(m[0]&~m[172]&m[173]&~m[174]&m[175])|(~m[0]&m[172]&m[173]&~m[174]&m[175])|(m[0]&~m[172]&~m[173]&m[174]&m[175])|(~m[0]&m[172]&~m[173]&m[174]&m[175])|(~m[0]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[259])|((m[0]&m[172]&m[173]&m[174]&~m[175])|(m[0]&m[172]&m[173]&~m[174]&m[175])|(m[0]&m[172]&~m[173]&m[174]&m[175])|(m[0]&~m[172]&m[173]&m[174]&m[175])|(~m[0]&m[172]&m[173]&m[174]&m[175])|(m[0]&m[172]&m[173]&m[174]&m[175]))):InitCond[530];
    m[36] = run?((((m[1]&m[176]&~m[177]&~m[178]&~m[179])|(m[1]&~m[176]&m[177]&~m[178]&~m[179])|(~m[1]&m[176]&m[177]&~m[178]&~m[179])|(m[1]&~m[176]&~m[177]&m[178]&~m[179])|(~m[1]&m[176]&~m[177]&m[178]&~m[179])|(~m[1]&~m[176]&m[177]&m[178]&~m[179])|(m[1]&~m[176]&~m[177]&~m[178]&m[179])|(~m[1]&m[176]&~m[177]&~m[178]&m[179])|(~m[1]&~m[176]&m[177]&~m[178]&m[179])|(~m[1]&~m[176]&~m[177]&m[178]&m[179]))&BiasedRNG[260])|(((m[1]&m[176]&m[177]&~m[178]&~m[179])|(m[1]&m[176]&~m[177]&m[178]&~m[179])|(m[1]&~m[176]&m[177]&m[178]&~m[179])|(~m[1]&m[176]&m[177]&m[178]&~m[179])|(m[1]&m[176]&~m[177]&~m[178]&m[179])|(m[1]&~m[176]&m[177]&~m[178]&m[179])|(~m[1]&m[176]&m[177]&~m[178]&m[179])|(m[1]&~m[176]&~m[177]&m[178]&m[179])|(~m[1]&m[176]&~m[177]&m[178]&m[179])|(~m[1]&~m[176]&m[177]&m[178]&m[179]))&~BiasedRNG[260])|((m[1]&m[176]&m[177]&m[178]&~m[179])|(m[1]&m[176]&m[177]&~m[178]&m[179])|(m[1]&m[176]&~m[177]&m[178]&m[179])|(m[1]&~m[176]&m[177]&m[178]&m[179])|(~m[1]&m[176]&m[177]&m[178]&m[179])|(m[1]&m[176]&m[177]&m[178]&m[179]))):InitCond[531];
    m[37] = run?((((m[1]&m[180]&~m[181]&~m[182]&~m[183])|(m[1]&~m[180]&m[181]&~m[182]&~m[183])|(~m[1]&m[180]&m[181]&~m[182]&~m[183])|(m[1]&~m[180]&~m[181]&m[182]&~m[183])|(~m[1]&m[180]&~m[181]&m[182]&~m[183])|(~m[1]&~m[180]&m[181]&m[182]&~m[183])|(m[1]&~m[180]&~m[181]&~m[182]&m[183])|(~m[1]&m[180]&~m[181]&~m[182]&m[183])|(~m[1]&~m[180]&m[181]&~m[182]&m[183])|(~m[1]&~m[180]&~m[181]&m[182]&m[183]))&BiasedRNG[261])|(((m[1]&m[180]&m[181]&~m[182]&~m[183])|(m[1]&m[180]&~m[181]&m[182]&~m[183])|(m[1]&~m[180]&m[181]&m[182]&~m[183])|(~m[1]&m[180]&m[181]&m[182]&~m[183])|(m[1]&m[180]&~m[181]&~m[182]&m[183])|(m[1]&~m[180]&m[181]&~m[182]&m[183])|(~m[1]&m[180]&m[181]&~m[182]&m[183])|(m[1]&~m[180]&~m[181]&m[182]&m[183])|(~m[1]&m[180]&~m[181]&m[182]&m[183])|(~m[1]&~m[180]&m[181]&m[182]&m[183]))&~BiasedRNG[261])|((m[1]&m[180]&m[181]&m[182]&~m[183])|(m[1]&m[180]&m[181]&~m[182]&m[183])|(m[1]&m[180]&~m[181]&m[182]&m[183])|(m[1]&~m[180]&m[181]&m[182]&m[183])|(~m[1]&m[180]&m[181]&m[182]&m[183])|(m[1]&m[180]&m[181]&m[182]&m[183]))):InitCond[532];
    m[38] = run?((((m[1]&m[184]&~m[185]&~m[186]&~m[187])|(m[1]&~m[184]&m[185]&~m[186]&~m[187])|(~m[1]&m[184]&m[185]&~m[186]&~m[187])|(m[1]&~m[184]&~m[185]&m[186]&~m[187])|(~m[1]&m[184]&~m[185]&m[186]&~m[187])|(~m[1]&~m[184]&m[185]&m[186]&~m[187])|(m[1]&~m[184]&~m[185]&~m[186]&m[187])|(~m[1]&m[184]&~m[185]&~m[186]&m[187])|(~m[1]&~m[184]&m[185]&~m[186]&m[187])|(~m[1]&~m[184]&~m[185]&m[186]&m[187]))&BiasedRNG[262])|(((m[1]&m[184]&m[185]&~m[186]&~m[187])|(m[1]&m[184]&~m[185]&m[186]&~m[187])|(m[1]&~m[184]&m[185]&m[186]&~m[187])|(~m[1]&m[184]&m[185]&m[186]&~m[187])|(m[1]&m[184]&~m[185]&~m[186]&m[187])|(m[1]&~m[184]&m[185]&~m[186]&m[187])|(~m[1]&m[184]&m[185]&~m[186]&m[187])|(m[1]&~m[184]&~m[185]&m[186]&m[187])|(~m[1]&m[184]&~m[185]&m[186]&m[187])|(~m[1]&~m[184]&m[185]&m[186]&m[187]))&~BiasedRNG[262])|((m[1]&m[184]&m[185]&m[186]&~m[187])|(m[1]&m[184]&m[185]&~m[186]&m[187])|(m[1]&m[184]&~m[185]&m[186]&m[187])|(m[1]&~m[184]&m[185]&m[186]&m[187])|(~m[1]&m[184]&m[185]&m[186]&m[187])|(m[1]&m[184]&m[185]&m[186]&m[187]))):InitCond[533];
    m[39] = run?((((m[1]&m[188]&~m[189]&~m[190]&~m[191])|(m[1]&~m[188]&m[189]&~m[190]&~m[191])|(~m[1]&m[188]&m[189]&~m[190]&~m[191])|(m[1]&~m[188]&~m[189]&m[190]&~m[191])|(~m[1]&m[188]&~m[189]&m[190]&~m[191])|(~m[1]&~m[188]&m[189]&m[190]&~m[191])|(m[1]&~m[188]&~m[189]&~m[190]&m[191])|(~m[1]&m[188]&~m[189]&~m[190]&m[191])|(~m[1]&~m[188]&m[189]&~m[190]&m[191])|(~m[1]&~m[188]&~m[189]&m[190]&m[191]))&BiasedRNG[263])|(((m[1]&m[188]&m[189]&~m[190]&~m[191])|(m[1]&m[188]&~m[189]&m[190]&~m[191])|(m[1]&~m[188]&m[189]&m[190]&~m[191])|(~m[1]&m[188]&m[189]&m[190]&~m[191])|(m[1]&m[188]&~m[189]&~m[190]&m[191])|(m[1]&~m[188]&m[189]&~m[190]&m[191])|(~m[1]&m[188]&m[189]&~m[190]&m[191])|(m[1]&~m[188]&~m[189]&m[190]&m[191])|(~m[1]&m[188]&~m[189]&m[190]&m[191])|(~m[1]&~m[188]&m[189]&m[190]&m[191]))&~BiasedRNG[263])|((m[1]&m[188]&m[189]&m[190]&~m[191])|(m[1]&m[188]&m[189]&~m[190]&m[191])|(m[1]&m[188]&~m[189]&m[190]&m[191])|(m[1]&~m[188]&m[189]&m[190]&m[191])|(~m[1]&m[188]&m[189]&m[190]&m[191])|(m[1]&m[188]&m[189]&m[190]&m[191]))):InitCond[534];
    m[40] = run?((((m[2]&m[192]&~m[193]&~m[194]&~m[195])|(m[2]&~m[192]&m[193]&~m[194]&~m[195])|(~m[2]&m[192]&m[193]&~m[194]&~m[195])|(m[2]&~m[192]&~m[193]&m[194]&~m[195])|(~m[2]&m[192]&~m[193]&m[194]&~m[195])|(~m[2]&~m[192]&m[193]&m[194]&~m[195])|(m[2]&~m[192]&~m[193]&~m[194]&m[195])|(~m[2]&m[192]&~m[193]&~m[194]&m[195])|(~m[2]&~m[192]&m[193]&~m[194]&m[195])|(~m[2]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[264])|(((m[2]&m[192]&m[193]&~m[194]&~m[195])|(m[2]&m[192]&~m[193]&m[194]&~m[195])|(m[2]&~m[192]&m[193]&m[194]&~m[195])|(~m[2]&m[192]&m[193]&m[194]&~m[195])|(m[2]&m[192]&~m[193]&~m[194]&m[195])|(m[2]&~m[192]&m[193]&~m[194]&m[195])|(~m[2]&m[192]&m[193]&~m[194]&m[195])|(m[2]&~m[192]&~m[193]&m[194]&m[195])|(~m[2]&m[192]&~m[193]&m[194]&m[195])|(~m[2]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[264])|((m[2]&m[192]&m[193]&m[194]&~m[195])|(m[2]&m[192]&m[193]&~m[194]&m[195])|(m[2]&m[192]&~m[193]&m[194]&m[195])|(m[2]&~m[192]&m[193]&m[194]&m[195])|(~m[2]&m[192]&m[193]&m[194]&m[195])|(m[2]&m[192]&m[193]&m[194]&m[195]))):InitCond[535];
    m[41] = run?((((m[2]&m[196]&~m[197]&~m[198]&~m[199])|(m[2]&~m[196]&m[197]&~m[198]&~m[199])|(~m[2]&m[196]&m[197]&~m[198]&~m[199])|(m[2]&~m[196]&~m[197]&m[198]&~m[199])|(~m[2]&m[196]&~m[197]&m[198]&~m[199])|(~m[2]&~m[196]&m[197]&m[198]&~m[199])|(m[2]&~m[196]&~m[197]&~m[198]&m[199])|(~m[2]&m[196]&~m[197]&~m[198]&m[199])|(~m[2]&~m[196]&m[197]&~m[198]&m[199])|(~m[2]&~m[196]&~m[197]&m[198]&m[199]))&BiasedRNG[265])|(((m[2]&m[196]&m[197]&~m[198]&~m[199])|(m[2]&m[196]&~m[197]&m[198]&~m[199])|(m[2]&~m[196]&m[197]&m[198]&~m[199])|(~m[2]&m[196]&m[197]&m[198]&~m[199])|(m[2]&m[196]&~m[197]&~m[198]&m[199])|(m[2]&~m[196]&m[197]&~m[198]&m[199])|(~m[2]&m[196]&m[197]&~m[198]&m[199])|(m[2]&~m[196]&~m[197]&m[198]&m[199])|(~m[2]&m[196]&~m[197]&m[198]&m[199])|(~m[2]&~m[196]&m[197]&m[198]&m[199]))&~BiasedRNG[265])|((m[2]&m[196]&m[197]&m[198]&~m[199])|(m[2]&m[196]&m[197]&~m[198]&m[199])|(m[2]&m[196]&~m[197]&m[198]&m[199])|(m[2]&~m[196]&m[197]&m[198]&m[199])|(~m[2]&m[196]&m[197]&m[198]&m[199])|(m[2]&m[196]&m[197]&m[198]&m[199]))):InitCond[536];
    m[42] = run?((((m[2]&m[200]&~m[201]&~m[202]&~m[203])|(m[2]&~m[200]&m[201]&~m[202]&~m[203])|(~m[2]&m[200]&m[201]&~m[202]&~m[203])|(m[2]&~m[200]&~m[201]&m[202]&~m[203])|(~m[2]&m[200]&~m[201]&m[202]&~m[203])|(~m[2]&~m[200]&m[201]&m[202]&~m[203])|(m[2]&~m[200]&~m[201]&~m[202]&m[203])|(~m[2]&m[200]&~m[201]&~m[202]&m[203])|(~m[2]&~m[200]&m[201]&~m[202]&m[203])|(~m[2]&~m[200]&~m[201]&m[202]&m[203]))&BiasedRNG[266])|(((m[2]&m[200]&m[201]&~m[202]&~m[203])|(m[2]&m[200]&~m[201]&m[202]&~m[203])|(m[2]&~m[200]&m[201]&m[202]&~m[203])|(~m[2]&m[200]&m[201]&m[202]&~m[203])|(m[2]&m[200]&~m[201]&~m[202]&m[203])|(m[2]&~m[200]&m[201]&~m[202]&m[203])|(~m[2]&m[200]&m[201]&~m[202]&m[203])|(m[2]&~m[200]&~m[201]&m[202]&m[203])|(~m[2]&m[200]&~m[201]&m[202]&m[203])|(~m[2]&~m[200]&m[201]&m[202]&m[203]))&~BiasedRNG[266])|((m[2]&m[200]&m[201]&m[202]&~m[203])|(m[2]&m[200]&m[201]&~m[202]&m[203])|(m[2]&m[200]&~m[201]&m[202]&m[203])|(m[2]&~m[200]&m[201]&m[202]&m[203])|(~m[2]&m[200]&m[201]&m[202]&m[203])|(m[2]&m[200]&m[201]&m[202]&m[203]))):InitCond[537];
    m[43] = run?((((m[2]&m[204]&~m[205]&~m[206]&~m[207])|(m[2]&~m[204]&m[205]&~m[206]&~m[207])|(~m[2]&m[204]&m[205]&~m[206]&~m[207])|(m[2]&~m[204]&~m[205]&m[206]&~m[207])|(~m[2]&m[204]&~m[205]&m[206]&~m[207])|(~m[2]&~m[204]&m[205]&m[206]&~m[207])|(m[2]&~m[204]&~m[205]&~m[206]&m[207])|(~m[2]&m[204]&~m[205]&~m[206]&m[207])|(~m[2]&~m[204]&m[205]&~m[206]&m[207])|(~m[2]&~m[204]&~m[205]&m[206]&m[207]))&BiasedRNG[267])|(((m[2]&m[204]&m[205]&~m[206]&~m[207])|(m[2]&m[204]&~m[205]&m[206]&~m[207])|(m[2]&~m[204]&m[205]&m[206]&~m[207])|(~m[2]&m[204]&m[205]&m[206]&~m[207])|(m[2]&m[204]&~m[205]&~m[206]&m[207])|(m[2]&~m[204]&m[205]&~m[206]&m[207])|(~m[2]&m[204]&m[205]&~m[206]&m[207])|(m[2]&~m[204]&~m[205]&m[206]&m[207])|(~m[2]&m[204]&~m[205]&m[206]&m[207])|(~m[2]&~m[204]&m[205]&m[206]&m[207]))&~BiasedRNG[267])|((m[2]&m[204]&m[205]&m[206]&~m[207])|(m[2]&m[204]&m[205]&~m[206]&m[207])|(m[2]&m[204]&~m[205]&m[206]&m[207])|(m[2]&~m[204]&m[205]&m[206]&m[207])|(~m[2]&m[204]&m[205]&m[206]&m[207])|(m[2]&m[204]&m[205]&m[206]&m[207]))):InitCond[538];
    m[44] = run?((((m[3]&m[208]&~m[209]&~m[210]&~m[211])|(m[3]&~m[208]&m[209]&~m[210]&~m[211])|(~m[3]&m[208]&m[209]&~m[210]&~m[211])|(m[3]&~m[208]&~m[209]&m[210]&~m[211])|(~m[3]&m[208]&~m[209]&m[210]&~m[211])|(~m[3]&~m[208]&m[209]&m[210]&~m[211])|(m[3]&~m[208]&~m[209]&~m[210]&m[211])|(~m[3]&m[208]&~m[209]&~m[210]&m[211])|(~m[3]&~m[208]&m[209]&~m[210]&m[211])|(~m[3]&~m[208]&~m[209]&m[210]&m[211]))&BiasedRNG[268])|(((m[3]&m[208]&m[209]&~m[210]&~m[211])|(m[3]&m[208]&~m[209]&m[210]&~m[211])|(m[3]&~m[208]&m[209]&m[210]&~m[211])|(~m[3]&m[208]&m[209]&m[210]&~m[211])|(m[3]&m[208]&~m[209]&~m[210]&m[211])|(m[3]&~m[208]&m[209]&~m[210]&m[211])|(~m[3]&m[208]&m[209]&~m[210]&m[211])|(m[3]&~m[208]&~m[209]&m[210]&m[211])|(~m[3]&m[208]&~m[209]&m[210]&m[211])|(~m[3]&~m[208]&m[209]&m[210]&m[211]))&~BiasedRNG[268])|((m[3]&m[208]&m[209]&m[210]&~m[211])|(m[3]&m[208]&m[209]&~m[210]&m[211])|(m[3]&m[208]&~m[209]&m[210]&m[211])|(m[3]&~m[208]&m[209]&m[210]&m[211])|(~m[3]&m[208]&m[209]&m[210]&m[211])|(m[3]&m[208]&m[209]&m[210]&m[211]))):InitCond[539];
    m[45] = run?((((m[3]&m[212]&~m[213]&~m[214]&~m[215])|(m[3]&~m[212]&m[213]&~m[214]&~m[215])|(~m[3]&m[212]&m[213]&~m[214]&~m[215])|(m[3]&~m[212]&~m[213]&m[214]&~m[215])|(~m[3]&m[212]&~m[213]&m[214]&~m[215])|(~m[3]&~m[212]&m[213]&m[214]&~m[215])|(m[3]&~m[212]&~m[213]&~m[214]&m[215])|(~m[3]&m[212]&~m[213]&~m[214]&m[215])|(~m[3]&~m[212]&m[213]&~m[214]&m[215])|(~m[3]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[269])|(((m[3]&m[212]&m[213]&~m[214]&~m[215])|(m[3]&m[212]&~m[213]&m[214]&~m[215])|(m[3]&~m[212]&m[213]&m[214]&~m[215])|(~m[3]&m[212]&m[213]&m[214]&~m[215])|(m[3]&m[212]&~m[213]&~m[214]&m[215])|(m[3]&~m[212]&m[213]&~m[214]&m[215])|(~m[3]&m[212]&m[213]&~m[214]&m[215])|(m[3]&~m[212]&~m[213]&m[214]&m[215])|(~m[3]&m[212]&~m[213]&m[214]&m[215])|(~m[3]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[269])|((m[3]&m[212]&m[213]&m[214]&~m[215])|(m[3]&m[212]&m[213]&~m[214]&m[215])|(m[3]&m[212]&~m[213]&m[214]&m[215])|(m[3]&~m[212]&m[213]&m[214]&m[215])|(~m[3]&m[212]&m[213]&m[214]&m[215])|(m[3]&m[212]&m[213]&m[214]&m[215]))):InitCond[540];
    m[46] = run?((((m[3]&m[216]&~m[217]&~m[218]&~m[219])|(m[3]&~m[216]&m[217]&~m[218]&~m[219])|(~m[3]&m[216]&m[217]&~m[218]&~m[219])|(m[3]&~m[216]&~m[217]&m[218]&~m[219])|(~m[3]&m[216]&~m[217]&m[218]&~m[219])|(~m[3]&~m[216]&m[217]&m[218]&~m[219])|(m[3]&~m[216]&~m[217]&~m[218]&m[219])|(~m[3]&m[216]&~m[217]&~m[218]&m[219])|(~m[3]&~m[216]&m[217]&~m[218]&m[219])|(~m[3]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[270])|(((m[3]&m[216]&m[217]&~m[218]&~m[219])|(m[3]&m[216]&~m[217]&m[218]&~m[219])|(m[3]&~m[216]&m[217]&m[218]&~m[219])|(~m[3]&m[216]&m[217]&m[218]&~m[219])|(m[3]&m[216]&~m[217]&~m[218]&m[219])|(m[3]&~m[216]&m[217]&~m[218]&m[219])|(~m[3]&m[216]&m[217]&~m[218]&m[219])|(m[3]&~m[216]&~m[217]&m[218]&m[219])|(~m[3]&m[216]&~m[217]&m[218]&m[219])|(~m[3]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[270])|((m[3]&m[216]&m[217]&m[218]&~m[219])|(m[3]&m[216]&m[217]&~m[218]&m[219])|(m[3]&m[216]&~m[217]&m[218]&m[219])|(m[3]&~m[216]&m[217]&m[218]&m[219])|(~m[3]&m[216]&m[217]&m[218]&m[219])|(m[3]&m[216]&m[217]&m[218]&m[219]))):InitCond[541];
    m[47] = run?((((m[3]&m[220]&~m[221]&~m[222]&~m[223])|(m[3]&~m[220]&m[221]&~m[222]&~m[223])|(~m[3]&m[220]&m[221]&~m[222]&~m[223])|(m[3]&~m[220]&~m[221]&m[222]&~m[223])|(~m[3]&m[220]&~m[221]&m[222]&~m[223])|(~m[3]&~m[220]&m[221]&m[222]&~m[223])|(m[3]&~m[220]&~m[221]&~m[222]&m[223])|(~m[3]&m[220]&~m[221]&~m[222]&m[223])|(~m[3]&~m[220]&m[221]&~m[222]&m[223])|(~m[3]&~m[220]&~m[221]&m[222]&m[223]))&BiasedRNG[271])|(((m[3]&m[220]&m[221]&~m[222]&~m[223])|(m[3]&m[220]&~m[221]&m[222]&~m[223])|(m[3]&~m[220]&m[221]&m[222]&~m[223])|(~m[3]&m[220]&m[221]&m[222]&~m[223])|(m[3]&m[220]&~m[221]&~m[222]&m[223])|(m[3]&~m[220]&m[221]&~m[222]&m[223])|(~m[3]&m[220]&m[221]&~m[222]&m[223])|(m[3]&~m[220]&~m[221]&m[222]&m[223])|(~m[3]&m[220]&~m[221]&m[222]&m[223])|(~m[3]&~m[220]&m[221]&m[222]&m[223]))&~BiasedRNG[271])|((m[3]&m[220]&m[221]&m[222]&~m[223])|(m[3]&m[220]&m[221]&~m[222]&m[223])|(m[3]&m[220]&~m[221]&m[222]&m[223])|(m[3]&~m[220]&m[221]&m[222]&m[223])|(~m[3]&m[220]&m[221]&m[222]&m[223])|(m[3]&m[220]&m[221]&m[222]&m[223]))):InitCond[542];
    m[48] = run?((((m[4]&m[224]&~m[225]&~m[226]&~m[227])|(m[4]&~m[224]&m[225]&~m[226]&~m[227])|(~m[4]&m[224]&m[225]&~m[226]&~m[227])|(m[4]&~m[224]&~m[225]&m[226]&~m[227])|(~m[4]&m[224]&~m[225]&m[226]&~m[227])|(~m[4]&~m[224]&m[225]&m[226]&~m[227])|(m[4]&~m[224]&~m[225]&~m[226]&m[227])|(~m[4]&m[224]&~m[225]&~m[226]&m[227])|(~m[4]&~m[224]&m[225]&~m[226]&m[227])|(~m[4]&~m[224]&~m[225]&m[226]&m[227]))&BiasedRNG[272])|(((m[4]&m[224]&m[225]&~m[226]&~m[227])|(m[4]&m[224]&~m[225]&m[226]&~m[227])|(m[4]&~m[224]&m[225]&m[226]&~m[227])|(~m[4]&m[224]&m[225]&m[226]&~m[227])|(m[4]&m[224]&~m[225]&~m[226]&m[227])|(m[4]&~m[224]&m[225]&~m[226]&m[227])|(~m[4]&m[224]&m[225]&~m[226]&m[227])|(m[4]&~m[224]&~m[225]&m[226]&m[227])|(~m[4]&m[224]&~m[225]&m[226]&m[227])|(~m[4]&~m[224]&m[225]&m[226]&m[227]))&~BiasedRNG[272])|((m[4]&m[224]&m[225]&m[226]&~m[227])|(m[4]&m[224]&m[225]&~m[226]&m[227])|(m[4]&m[224]&~m[225]&m[226]&m[227])|(m[4]&~m[224]&m[225]&m[226]&m[227])|(~m[4]&m[224]&m[225]&m[226]&m[227])|(m[4]&m[224]&m[225]&m[226]&m[227]))):InitCond[543];
    m[49] = run?((((m[4]&m[228]&~m[229]&~m[230]&~m[231])|(m[4]&~m[228]&m[229]&~m[230]&~m[231])|(~m[4]&m[228]&m[229]&~m[230]&~m[231])|(m[4]&~m[228]&~m[229]&m[230]&~m[231])|(~m[4]&m[228]&~m[229]&m[230]&~m[231])|(~m[4]&~m[228]&m[229]&m[230]&~m[231])|(m[4]&~m[228]&~m[229]&~m[230]&m[231])|(~m[4]&m[228]&~m[229]&~m[230]&m[231])|(~m[4]&~m[228]&m[229]&~m[230]&m[231])|(~m[4]&~m[228]&~m[229]&m[230]&m[231]))&BiasedRNG[273])|(((m[4]&m[228]&m[229]&~m[230]&~m[231])|(m[4]&m[228]&~m[229]&m[230]&~m[231])|(m[4]&~m[228]&m[229]&m[230]&~m[231])|(~m[4]&m[228]&m[229]&m[230]&~m[231])|(m[4]&m[228]&~m[229]&~m[230]&m[231])|(m[4]&~m[228]&m[229]&~m[230]&m[231])|(~m[4]&m[228]&m[229]&~m[230]&m[231])|(m[4]&~m[228]&~m[229]&m[230]&m[231])|(~m[4]&m[228]&~m[229]&m[230]&m[231])|(~m[4]&~m[228]&m[229]&m[230]&m[231]))&~BiasedRNG[273])|((m[4]&m[228]&m[229]&m[230]&~m[231])|(m[4]&m[228]&m[229]&~m[230]&m[231])|(m[4]&m[228]&~m[229]&m[230]&m[231])|(m[4]&~m[228]&m[229]&m[230]&m[231])|(~m[4]&m[228]&m[229]&m[230]&m[231])|(m[4]&m[228]&m[229]&m[230]&m[231]))):InitCond[544];
    m[50] = run?((((m[4]&m[232]&~m[233]&~m[234]&~m[235])|(m[4]&~m[232]&m[233]&~m[234]&~m[235])|(~m[4]&m[232]&m[233]&~m[234]&~m[235])|(m[4]&~m[232]&~m[233]&m[234]&~m[235])|(~m[4]&m[232]&~m[233]&m[234]&~m[235])|(~m[4]&~m[232]&m[233]&m[234]&~m[235])|(m[4]&~m[232]&~m[233]&~m[234]&m[235])|(~m[4]&m[232]&~m[233]&~m[234]&m[235])|(~m[4]&~m[232]&m[233]&~m[234]&m[235])|(~m[4]&~m[232]&~m[233]&m[234]&m[235]))&BiasedRNG[274])|(((m[4]&m[232]&m[233]&~m[234]&~m[235])|(m[4]&m[232]&~m[233]&m[234]&~m[235])|(m[4]&~m[232]&m[233]&m[234]&~m[235])|(~m[4]&m[232]&m[233]&m[234]&~m[235])|(m[4]&m[232]&~m[233]&~m[234]&m[235])|(m[4]&~m[232]&m[233]&~m[234]&m[235])|(~m[4]&m[232]&m[233]&~m[234]&m[235])|(m[4]&~m[232]&~m[233]&m[234]&m[235])|(~m[4]&m[232]&~m[233]&m[234]&m[235])|(~m[4]&~m[232]&m[233]&m[234]&m[235]))&~BiasedRNG[274])|((m[4]&m[232]&m[233]&m[234]&~m[235])|(m[4]&m[232]&m[233]&~m[234]&m[235])|(m[4]&m[232]&~m[233]&m[234]&m[235])|(m[4]&~m[232]&m[233]&m[234]&m[235])|(~m[4]&m[232]&m[233]&m[234]&m[235])|(m[4]&m[232]&m[233]&m[234]&m[235]))):InitCond[545];
    m[51] = run?((((m[4]&m[236]&~m[237]&~m[238]&~m[239])|(m[4]&~m[236]&m[237]&~m[238]&~m[239])|(~m[4]&m[236]&m[237]&~m[238]&~m[239])|(m[4]&~m[236]&~m[237]&m[238]&~m[239])|(~m[4]&m[236]&~m[237]&m[238]&~m[239])|(~m[4]&~m[236]&m[237]&m[238]&~m[239])|(m[4]&~m[236]&~m[237]&~m[238]&m[239])|(~m[4]&m[236]&~m[237]&~m[238]&m[239])|(~m[4]&~m[236]&m[237]&~m[238]&m[239])|(~m[4]&~m[236]&~m[237]&m[238]&m[239]))&BiasedRNG[275])|(((m[4]&m[236]&m[237]&~m[238]&~m[239])|(m[4]&m[236]&~m[237]&m[238]&~m[239])|(m[4]&~m[236]&m[237]&m[238]&~m[239])|(~m[4]&m[236]&m[237]&m[238]&~m[239])|(m[4]&m[236]&~m[237]&~m[238]&m[239])|(m[4]&~m[236]&m[237]&~m[238]&m[239])|(~m[4]&m[236]&m[237]&~m[238]&m[239])|(m[4]&~m[236]&~m[237]&m[238]&m[239])|(~m[4]&m[236]&~m[237]&m[238]&m[239])|(~m[4]&~m[236]&m[237]&m[238]&m[239]))&~BiasedRNG[275])|((m[4]&m[236]&m[237]&m[238]&~m[239])|(m[4]&m[236]&m[237]&~m[238]&m[239])|(m[4]&m[236]&~m[237]&m[238]&m[239])|(m[4]&~m[236]&m[237]&m[238]&m[239])|(~m[4]&m[236]&m[237]&m[238]&m[239])|(m[4]&m[236]&m[237]&m[238]&m[239]))):InitCond[546];
    m[52] = run?((((m[5]&m[240]&~m[241]&~m[242]&~m[243])|(m[5]&~m[240]&m[241]&~m[242]&~m[243])|(~m[5]&m[240]&m[241]&~m[242]&~m[243])|(m[5]&~m[240]&~m[241]&m[242]&~m[243])|(~m[5]&m[240]&~m[241]&m[242]&~m[243])|(~m[5]&~m[240]&m[241]&m[242]&~m[243])|(m[5]&~m[240]&~m[241]&~m[242]&m[243])|(~m[5]&m[240]&~m[241]&~m[242]&m[243])|(~m[5]&~m[240]&m[241]&~m[242]&m[243])|(~m[5]&~m[240]&~m[241]&m[242]&m[243]))&BiasedRNG[276])|(((m[5]&m[240]&m[241]&~m[242]&~m[243])|(m[5]&m[240]&~m[241]&m[242]&~m[243])|(m[5]&~m[240]&m[241]&m[242]&~m[243])|(~m[5]&m[240]&m[241]&m[242]&~m[243])|(m[5]&m[240]&~m[241]&~m[242]&m[243])|(m[5]&~m[240]&m[241]&~m[242]&m[243])|(~m[5]&m[240]&m[241]&~m[242]&m[243])|(m[5]&~m[240]&~m[241]&m[242]&m[243])|(~m[5]&m[240]&~m[241]&m[242]&m[243])|(~m[5]&~m[240]&m[241]&m[242]&m[243]))&~BiasedRNG[276])|((m[5]&m[240]&m[241]&m[242]&~m[243])|(m[5]&m[240]&m[241]&~m[242]&m[243])|(m[5]&m[240]&~m[241]&m[242]&m[243])|(m[5]&~m[240]&m[241]&m[242]&m[243])|(~m[5]&m[240]&m[241]&m[242]&m[243])|(m[5]&m[240]&m[241]&m[242]&m[243]))):InitCond[547];
    m[53] = run?((((m[5]&m[244]&~m[245]&~m[246]&~m[247])|(m[5]&~m[244]&m[245]&~m[246]&~m[247])|(~m[5]&m[244]&m[245]&~m[246]&~m[247])|(m[5]&~m[244]&~m[245]&m[246]&~m[247])|(~m[5]&m[244]&~m[245]&m[246]&~m[247])|(~m[5]&~m[244]&m[245]&m[246]&~m[247])|(m[5]&~m[244]&~m[245]&~m[246]&m[247])|(~m[5]&m[244]&~m[245]&~m[246]&m[247])|(~m[5]&~m[244]&m[245]&~m[246]&m[247])|(~m[5]&~m[244]&~m[245]&m[246]&m[247]))&BiasedRNG[277])|(((m[5]&m[244]&m[245]&~m[246]&~m[247])|(m[5]&m[244]&~m[245]&m[246]&~m[247])|(m[5]&~m[244]&m[245]&m[246]&~m[247])|(~m[5]&m[244]&m[245]&m[246]&~m[247])|(m[5]&m[244]&~m[245]&~m[246]&m[247])|(m[5]&~m[244]&m[245]&~m[246]&m[247])|(~m[5]&m[244]&m[245]&~m[246]&m[247])|(m[5]&~m[244]&~m[245]&m[246]&m[247])|(~m[5]&m[244]&~m[245]&m[246]&m[247])|(~m[5]&~m[244]&m[245]&m[246]&m[247]))&~BiasedRNG[277])|((m[5]&m[244]&m[245]&m[246]&~m[247])|(m[5]&m[244]&m[245]&~m[246]&m[247])|(m[5]&m[244]&~m[245]&m[246]&m[247])|(m[5]&~m[244]&m[245]&m[246]&m[247])|(~m[5]&m[244]&m[245]&m[246]&m[247])|(m[5]&m[244]&m[245]&m[246]&m[247]))):InitCond[548];
    m[54] = run?((((m[5]&m[248]&~m[249]&~m[250]&~m[251])|(m[5]&~m[248]&m[249]&~m[250]&~m[251])|(~m[5]&m[248]&m[249]&~m[250]&~m[251])|(m[5]&~m[248]&~m[249]&m[250]&~m[251])|(~m[5]&m[248]&~m[249]&m[250]&~m[251])|(~m[5]&~m[248]&m[249]&m[250]&~m[251])|(m[5]&~m[248]&~m[249]&~m[250]&m[251])|(~m[5]&m[248]&~m[249]&~m[250]&m[251])|(~m[5]&~m[248]&m[249]&~m[250]&m[251])|(~m[5]&~m[248]&~m[249]&m[250]&m[251]))&BiasedRNG[278])|(((m[5]&m[248]&m[249]&~m[250]&~m[251])|(m[5]&m[248]&~m[249]&m[250]&~m[251])|(m[5]&~m[248]&m[249]&m[250]&~m[251])|(~m[5]&m[248]&m[249]&m[250]&~m[251])|(m[5]&m[248]&~m[249]&~m[250]&m[251])|(m[5]&~m[248]&m[249]&~m[250]&m[251])|(~m[5]&m[248]&m[249]&~m[250]&m[251])|(m[5]&~m[248]&~m[249]&m[250]&m[251])|(~m[5]&m[248]&~m[249]&m[250]&m[251])|(~m[5]&~m[248]&m[249]&m[250]&m[251]))&~BiasedRNG[278])|((m[5]&m[248]&m[249]&m[250]&~m[251])|(m[5]&m[248]&m[249]&~m[250]&m[251])|(m[5]&m[248]&~m[249]&m[250]&m[251])|(m[5]&~m[248]&m[249]&m[250]&m[251])|(~m[5]&m[248]&m[249]&m[250]&m[251])|(m[5]&m[248]&m[249]&m[250]&m[251]))):InitCond[549];
    m[55] = run?((((m[5]&m[252]&~m[253]&~m[254]&~m[255])|(m[5]&~m[252]&m[253]&~m[254]&~m[255])|(~m[5]&m[252]&m[253]&~m[254]&~m[255])|(m[5]&~m[252]&~m[253]&m[254]&~m[255])|(~m[5]&m[252]&~m[253]&m[254]&~m[255])|(~m[5]&~m[252]&m[253]&m[254]&~m[255])|(m[5]&~m[252]&~m[253]&~m[254]&m[255])|(~m[5]&m[252]&~m[253]&~m[254]&m[255])|(~m[5]&~m[252]&m[253]&~m[254]&m[255])|(~m[5]&~m[252]&~m[253]&m[254]&m[255]))&BiasedRNG[279])|(((m[5]&m[252]&m[253]&~m[254]&~m[255])|(m[5]&m[252]&~m[253]&m[254]&~m[255])|(m[5]&~m[252]&m[253]&m[254]&~m[255])|(~m[5]&m[252]&m[253]&m[254]&~m[255])|(m[5]&m[252]&~m[253]&~m[254]&m[255])|(m[5]&~m[252]&m[253]&~m[254]&m[255])|(~m[5]&m[252]&m[253]&~m[254]&m[255])|(m[5]&~m[252]&~m[253]&m[254]&m[255])|(~m[5]&m[252]&~m[253]&m[254]&m[255])|(~m[5]&~m[252]&m[253]&m[254]&m[255]))&~BiasedRNG[279])|((m[5]&m[252]&m[253]&m[254]&~m[255])|(m[5]&m[252]&m[253]&~m[254]&m[255])|(m[5]&m[252]&~m[253]&m[254]&m[255])|(m[5]&~m[252]&m[253]&m[254]&m[255])|(~m[5]&m[252]&m[253]&m[254]&m[255])|(m[5]&m[252]&m[253]&m[254]&m[255]))):InitCond[550];
    m[56] = run?((((m[6]&m[256]&~m[257]&~m[258]&~m[259])|(m[6]&~m[256]&m[257]&~m[258]&~m[259])|(~m[6]&m[256]&m[257]&~m[258]&~m[259])|(m[6]&~m[256]&~m[257]&m[258]&~m[259])|(~m[6]&m[256]&~m[257]&m[258]&~m[259])|(~m[6]&~m[256]&m[257]&m[258]&~m[259])|(m[6]&~m[256]&~m[257]&~m[258]&m[259])|(~m[6]&m[256]&~m[257]&~m[258]&m[259])|(~m[6]&~m[256]&m[257]&~m[258]&m[259])|(~m[6]&~m[256]&~m[257]&m[258]&m[259]))&BiasedRNG[280])|(((m[6]&m[256]&m[257]&~m[258]&~m[259])|(m[6]&m[256]&~m[257]&m[258]&~m[259])|(m[6]&~m[256]&m[257]&m[258]&~m[259])|(~m[6]&m[256]&m[257]&m[258]&~m[259])|(m[6]&m[256]&~m[257]&~m[258]&m[259])|(m[6]&~m[256]&m[257]&~m[258]&m[259])|(~m[6]&m[256]&m[257]&~m[258]&m[259])|(m[6]&~m[256]&~m[257]&m[258]&m[259])|(~m[6]&m[256]&~m[257]&m[258]&m[259])|(~m[6]&~m[256]&m[257]&m[258]&m[259]))&~BiasedRNG[280])|((m[6]&m[256]&m[257]&m[258]&~m[259])|(m[6]&m[256]&m[257]&~m[258]&m[259])|(m[6]&m[256]&~m[257]&m[258]&m[259])|(m[6]&~m[256]&m[257]&m[258]&m[259])|(~m[6]&m[256]&m[257]&m[258]&m[259])|(m[6]&m[256]&m[257]&m[258]&m[259]))):InitCond[551];
    m[57] = run?((((m[6]&m[260]&~m[261]&~m[262]&~m[263])|(m[6]&~m[260]&m[261]&~m[262]&~m[263])|(~m[6]&m[260]&m[261]&~m[262]&~m[263])|(m[6]&~m[260]&~m[261]&m[262]&~m[263])|(~m[6]&m[260]&~m[261]&m[262]&~m[263])|(~m[6]&~m[260]&m[261]&m[262]&~m[263])|(m[6]&~m[260]&~m[261]&~m[262]&m[263])|(~m[6]&m[260]&~m[261]&~m[262]&m[263])|(~m[6]&~m[260]&m[261]&~m[262]&m[263])|(~m[6]&~m[260]&~m[261]&m[262]&m[263]))&BiasedRNG[281])|(((m[6]&m[260]&m[261]&~m[262]&~m[263])|(m[6]&m[260]&~m[261]&m[262]&~m[263])|(m[6]&~m[260]&m[261]&m[262]&~m[263])|(~m[6]&m[260]&m[261]&m[262]&~m[263])|(m[6]&m[260]&~m[261]&~m[262]&m[263])|(m[6]&~m[260]&m[261]&~m[262]&m[263])|(~m[6]&m[260]&m[261]&~m[262]&m[263])|(m[6]&~m[260]&~m[261]&m[262]&m[263])|(~m[6]&m[260]&~m[261]&m[262]&m[263])|(~m[6]&~m[260]&m[261]&m[262]&m[263]))&~BiasedRNG[281])|((m[6]&m[260]&m[261]&m[262]&~m[263])|(m[6]&m[260]&m[261]&~m[262]&m[263])|(m[6]&m[260]&~m[261]&m[262]&m[263])|(m[6]&~m[260]&m[261]&m[262]&m[263])|(~m[6]&m[260]&m[261]&m[262]&m[263])|(m[6]&m[260]&m[261]&m[262]&m[263]))):InitCond[552];
    m[58] = run?((((m[6]&m[264]&~m[265]&~m[266]&~m[267])|(m[6]&~m[264]&m[265]&~m[266]&~m[267])|(~m[6]&m[264]&m[265]&~m[266]&~m[267])|(m[6]&~m[264]&~m[265]&m[266]&~m[267])|(~m[6]&m[264]&~m[265]&m[266]&~m[267])|(~m[6]&~m[264]&m[265]&m[266]&~m[267])|(m[6]&~m[264]&~m[265]&~m[266]&m[267])|(~m[6]&m[264]&~m[265]&~m[266]&m[267])|(~m[6]&~m[264]&m[265]&~m[266]&m[267])|(~m[6]&~m[264]&~m[265]&m[266]&m[267]))&BiasedRNG[282])|(((m[6]&m[264]&m[265]&~m[266]&~m[267])|(m[6]&m[264]&~m[265]&m[266]&~m[267])|(m[6]&~m[264]&m[265]&m[266]&~m[267])|(~m[6]&m[264]&m[265]&m[266]&~m[267])|(m[6]&m[264]&~m[265]&~m[266]&m[267])|(m[6]&~m[264]&m[265]&~m[266]&m[267])|(~m[6]&m[264]&m[265]&~m[266]&m[267])|(m[6]&~m[264]&~m[265]&m[266]&m[267])|(~m[6]&m[264]&~m[265]&m[266]&m[267])|(~m[6]&~m[264]&m[265]&m[266]&m[267]))&~BiasedRNG[282])|((m[6]&m[264]&m[265]&m[266]&~m[267])|(m[6]&m[264]&m[265]&~m[266]&m[267])|(m[6]&m[264]&~m[265]&m[266]&m[267])|(m[6]&~m[264]&m[265]&m[266]&m[267])|(~m[6]&m[264]&m[265]&m[266]&m[267])|(m[6]&m[264]&m[265]&m[266]&m[267]))):InitCond[553];
    m[59] = run?((((m[6]&m[268]&~m[269]&~m[270]&~m[271])|(m[6]&~m[268]&m[269]&~m[270]&~m[271])|(~m[6]&m[268]&m[269]&~m[270]&~m[271])|(m[6]&~m[268]&~m[269]&m[270]&~m[271])|(~m[6]&m[268]&~m[269]&m[270]&~m[271])|(~m[6]&~m[268]&m[269]&m[270]&~m[271])|(m[6]&~m[268]&~m[269]&~m[270]&m[271])|(~m[6]&m[268]&~m[269]&~m[270]&m[271])|(~m[6]&~m[268]&m[269]&~m[270]&m[271])|(~m[6]&~m[268]&~m[269]&m[270]&m[271]))&BiasedRNG[283])|(((m[6]&m[268]&m[269]&~m[270]&~m[271])|(m[6]&m[268]&~m[269]&m[270]&~m[271])|(m[6]&~m[268]&m[269]&m[270]&~m[271])|(~m[6]&m[268]&m[269]&m[270]&~m[271])|(m[6]&m[268]&~m[269]&~m[270]&m[271])|(m[6]&~m[268]&m[269]&~m[270]&m[271])|(~m[6]&m[268]&m[269]&~m[270]&m[271])|(m[6]&~m[268]&~m[269]&m[270]&m[271])|(~m[6]&m[268]&~m[269]&m[270]&m[271])|(~m[6]&~m[268]&m[269]&m[270]&m[271]))&~BiasedRNG[283])|((m[6]&m[268]&m[269]&m[270]&~m[271])|(m[6]&m[268]&m[269]&~m[270]&m[271])|(m[6]&m[268]&~m[269]&m[270]&m[271])|(m[6]&~m[268]&m[269]&m[270]&m[271])|(~m[6]&m[268]&m[269]&m[270]&m[271])|(m[6]&m[268]&m[269]&m[270]&m[271]))):InitCond[554];
    m[60] = run?((((m[7]&m[272]&~m[273]&~m[274]&~m[275])|(m[7]&~m[272]&m[273]&~m[274]&~m[275])|(~m[7]&m[272]&m[273]&~m[274]&~m[275])|(m[7]&~m[272]&~m[273]&m[274]&~m[275])|(~m[7]&m[272]&~m[273]&m[274]&~m[275])|(~m[7]&~m[272]&m[273]&m[274]&~m[275])|(m[7]&~m[272]&~m[273]&~m[274]&m[275])|(~m[7]&m[272]&~m[273]&~m[274]&m[275])|(~m[7]&~m[272]&m[273]&~m[274]&m[275])|(~m[7]&~m[272]&~m[273]&m[274]&m[275]))&BiasedRNG[284])|(((m[7]&m[272]&m[273]&~m[274]&~m[275])|(m[7]&m[272]&~m[273]&m[274]&~m[275])|(m[7]&~m[272]&m[273]&m[274]&~m[275])|(~m[7]&m[272]&m[273]&m[274]&~m[275])|(m[7]&m[272]&~m[273]&~m[274]&m[275])|(m[7]&~m[272]&m[273]&~m[274]&m[275])|(~m[7]&m[272]&m[273]&~m[274]&m[275])|(m[7]&~m[272]&~m[273]&m[274]&m[275])|(~m[7]&m[272]&~m[273]&m[274]&m[275])|(~m[7]&~m[272]&m[273]&m[274]&m[275]))&~BiasedRNG[284])|((m[7]&m[272]&m[273]&m[274]&~m[275])|(m[7]&m[272]&m[273]&~m[274]&m[275])|(m[7]&m[272]&~m[273]&m[274]&m[275])|(m[7]&~m[272]&m[273]&m[274]&m[275])|(~m[7]&m[272]&m[273]&m[274]&m[275])|(m[7]&m[272]&m[273]&m[274]&m[275]))):InitCond[555];
    m[61] = run?((((m[7]&m[276]&~m[277]&~m[278]&~m[279])|(m[7]&~m[276]&m[277]&~m[278]&~m[279])|(~m[7]&m[276]&m[277]&~m[278]&~m[279])|(m[7]&~m[276]&~m[277]&m[278]&~m[279])|(~m[7]&m[276]&~m[277]&m[278]&~m[279])|(~m[7]&~m[276]&m[277]&m[278]&~m[279])|(m[7]&~m[276]&~m[277]&~m[278]&m[279])|(~m[7]&m[276]&~m[277]&~m[278]&m[279])|(~m[7]&~m[276]&m[277]&~m[278]&m[279])|(~m[7]&~m[276]&~m[277]&m[278]&m[279]))&BiasedRNG[285])|(((m[7]&m[276]&m[277]&~m[278]&~m[279])|(m[7]&m[276]&~m[277]&m[278]&~m[279])|(m[7]&~m[276]&m[277]&m[278]&~m[279])|(~m[7]&m[276]&m[277]&m[278]&~m[279])|(m[7]&m[276]&~m[277]&~m[278]&m[279])|(m[7]&~m[276]&m[277]&~m[278]&m[279])|(~m[7]&m[276]&m[277]&~m[278]&m[279])|(m[7]&~m[276]&~m[277]&m[278]&m[279])|(~m[7]&m[276]&~m[277]&m[278]&m[279])|(~m[7]&~m[276]&m[277]&m[278]&m[279]))&~BiasedRNG[285])|((m[7]&m[276]&m[277]&m[278]&~m[279])|(m[7]&m[276]&m[277]&~m[278]&m[279])|(m[7]&m[276]&~m[277]&m[278]&m[279])|(m[7]&~m[276]&m[277]&m[278]&m[279])|(~m[7]&m[276]&m[277]&m[278]&m[279])|(m[7]&m[276]&m[277]&m[278]&m[279]))):InitCond[556];
    m[62] = run?((((m[7]&m[280]&~m[281]&~m[282]&~m[283])|(m[7]&~m[280]&m[281]&~m[282]&~m[283])|(~m[7]&m[280]&m[281]&~m[282]&~m[283])|(m[7]&~m[280]&~m[281]&m[282]&~m[283])|(~m[7]&m[280]&~m[281]&m[282]&~m[283])|(~m[7]&~m[280]&m[281]&m[282]&~m[283])|(m[7]&~m[280]&~m[281]&~m[282]&m[283])|(~m[7]&m[280]&~m[281]&~m[282]&m[283])|(~m[7]&~m[280]&m[281]&~m[282]&m[283])|(~m[7]&~m[280]&~m[281]&m[282]&m[283]))&BiasedRNG[286])|(((m[7]&m[280]&m[281]&~m[282]&~m[283])|(m[7]&m[280]&~m[281]&m[282]&~m[283])|(m[7]&~m[280]&m[281]&m[282]&~m[283])|(~m[7]&m[280]&m[281]&m[282]&~m[283])|(m[7]&m[280]&~m[281]&~m[282]&m[283])|(m[7]&~m[280]&m[281]&~m[282]&m[283])|(~m[7]&m[280]&m[281]&~m[282]&m[283])|(m[7]&~m[280]&~m[281]&m[282]&m[283])|(~m[7]&m[280]&~m[281]&m[282]&m[283])|(~m[7]&~m[280]&m[281]&m[282]&m[283]))&~BiasedRNG[286])|((m[7]&m[280]&m[281]&m[282]&~m[283])|(m[7]&m[280]&m[281]&~m[282]&m[283])|(m[7]&m[280]&~m[281]&m[282]&m[283])|(m[7]&~m[280]&m[281]&m[282]&m[283])|(~m[7]&m[280]&m[281]&m[282]&m[283])|(m[7]&m[280]&m[281]&m[282]&m[283]))):InitCond[557];
    m[63] = run?((((m[7]&m[284]&~m[285]&~m[286]&~m[287])|(m[7]&~m[284]&m[285]&~m[286]&~m[287])|(~m[7]&m[284]&m[285]&~m[286]&~m[287])|(m[7]&~m[284]&~m[285]&m[286]&~m[287])|(~m[7]&m[284]&~m[285]&m[286]&~m[287])|(~m[7]&~m[284]&m[285]&m[286]&~m[287])|(m[7]&~m[284]&~m[285]&~m[286]&m[287])|(~m[7]&m[284]&~m[285]&~m[286]&m[287])|(~m[7]&~m[284]&m[285]&~m[286]&m[287])|(~m[7]&~m[284]&~m[285]&m[286]&m[287]))&BiasedRNG[287])|(((m[7]&m[284]&m[285]&~m[286]&~m[287])|(m[7]&m[284]&~m[285]&m[286]&~m[287])|(m[7]&~m[284]&m[285]&m[286]&~m[287])|(~m[7]&m[284]&m[285]&m[286]&~m[287])|(m[7]&m[284]&~m[285]&~m[286]&m[287])|(m[7]&~m[284]&m[285]&~m[286]&m[287])|(~m[7]&m[284]&m[285]&~m[286]&m[287])|(m[7]&~m[284]&~m[285]&m[286]&m[287])|(~m[7]&m[284]&~m[285]&m[286]&m[287])|(~m[7]&~m[284]&m[285]&m[286]&m[287]))&~BiasedRNG[287])|((m[7]&m[284]&m[285]&m[286]&~m[287])|(m[7]&m[284]&m[285]&~m[286]&m[287])|(m[7]&m[284]&~m[285]&m[286]&m[287])|(m[7]&~m[284]&m[285]&m[286]&m[287])|(~m[7]&m[284]&m[285]&m[286]&m[287])|(m[7]&m[284]&m[285]&m[286]&m[287]))):InitCond[558];
    m[64] = run?((((m[8]&m[288]&~m[289]&~m[290]&~m[291])|(m[8]&~m[288]&m[289]&~m[290]&~m[291])|(~m[8]&m[288]&m[289]&~m[290]&~m[291])|(m[8]&~m[288]&~m[289]&m[290]&~m[291])|(~m[8]&m[288]&~m[289]&m[290]&~m[291])|(~m[8]&~m[288]&m[289]&m[290]&~m[291])|(m[8]&~m[288]&~m[289]&~m[290]&m[291])|(~m[8]&m[288]&~m[289]&~m[290]&m[291])|(~m[8]&~m[288]&m[289]&~m[290]&m[291])|(~m[8]&~m[288]&~m[289]&m[290]&m[291]))&BiasedRNG[288])|(((m[8]&m[288]&m[289]&~m[290]&~m[291])|(m[8]&m[288]&~m[289]&m[290]&~m[291])|(m[8]&~m[288]&m[289]&m[290]&~m[291])|(~m[8]&m[288]&m[289]&m[290]&~m[291])|(m[8]&m[288]&~m[289]&~m[290]&m[291])|(m[8]&~m[288]&m[289]&~m[290]&m[291])|(~m[8]&m[288]&m[289]&~m[290]&m[291])|(m[8]&~m[288]&~m[289]&m[290]&m[291])|(~m[8]&m[288]&~m[289]&m[290]&m[291])|(~m[8]&~m[288]&m[289]&m[290]&m[291]))&~BiasedRNG[288])|((m[8]&m[288]&m[289]&m[290]&~m[291])|(m[8]&m[288]&m[289]&~m[290]&m[291])|(m[8]&m[288]&~m[289]&m[290]&m[291])|(m[8]&~m[288]&m[289]&m[290]&m[291])|(~m[8]&m[288]&m[289]&m[290]&m[291])|(m[8]&m[288]&m[289]&m[290]&m[291]))):InitCond[559];
    m[65] = run?((((m[8]&m[292]&~m[293]&~m[294]&~m[295])|(m[8]&~m[292]&m[293]&~m[294]&~m[295])|(~m[8]&m[292]&m[293]&~m[294]&~m[295])|(m[8]&~m[292]&~m[293]&m[294]&~m[295])|(~m[8]&m[292]&~m[293]&m[294]&~m[295])|(~m[8]&~m[292]&m[293]&m[294]&~m[295])|(m[8]&~m[292]&~m[293]&~m[294]&m[295])|(~m[8]&m[292]&~m[293]&~m[294]&m[295])|(~m[8]&~m[292]&m[293]&~m[294]&m[295])|(~m[8]&~m[292]&~m[293]&m[294]&m[295]))&BiasedRNG[289])|(((m[8]&m[292]&m[293]&~m[294]&~m[295])|(m[8]&m[292]&~m[293]&m[294]&~m[295])|(m[8]&~m[292]&m[293]&m[294]&~m[295])|(~m[8]&m[292]&m[293]&m[294]&~m[295])|(m[8]&m[292]&~m[293]&~m[294]&m[295])|(m[8]&~m[292]&m[293]&~m[294]&m[295])|(~m[8]&m[292]&m[293]&~m[294]&m[295])|(m[8]&~m[292]&~m[293]&m[294]&m[295])|(~m[8]&m[292]&~m[293]&m[294]&m[295])|(~m[8]&~m[292]&m[293]&m[294]&m[295]))&~BiasedRNG[289])|((m[8]&m[292]&m[293]&m[294]&~m[295])|(m[8]&m[292]&m[293]&~m[294]&m[295])|(m[8]&m[292]&~m[293]&m[294]&m[295])|(m[8]&~m[292]&m[293]&m[294]&m[295])|(~m[8]&m[292]&m[293]&m[294]&m[295])|(m[8]&m[292]&m[293]&m[294]&m[295]))):InitCond[560];
    m[66] = run?((((m[8]&m[296]&~m[297]&~m[298]&~m[299])|(m[8]&~m[296]&m[297]&~m[298]&~m[299])|(~m[8]&m[296]&m[297]&~m[298]&~m[299])|(m[8]&~m[296]&~m[297]&m[298]&~m[299])|(~m[8]&m[296]&~m[297]&m[298]&~m[299])|(~m[8]&~m[296]&m[297]&m[298]&~m[299])|(m[8]&~m[296]&~m[297]&~m[298]&m[299])|(~m[8]&m[296]&~m[297]&~m[298]&m[299])|(~m[8]&~m[296]&m[297]&~m[298]&m[299])|(~m[8]&~m[296]&~m[297]&m[298]&m[299]))&BiasedRNG[290])|(((m[8]&m[296]&m[297]&~m[298]&~m[299])|(m[8]&m[296]&~m[297]&m[298]&~m[299])|(m[8]&~m[296]&m[297]&m[298]&~m[299])|(~m[8]&m[296]&m[297]&m[298]&~m[299])|(m[8]&m[296]&~m[297]&~m[298]&m[299])|(m[8]&~m[296]&m[297]&~m[298]&m[299])|(~m[8]&m[296]&m[297]&~m[298]&m[299])|(m[8]&~m[296]&~m[297]&m[298]&m[299])|(~m[8]&m[296]&~m[297]&m[298]&m[299])|(~m[8]&~m[296]&m[297]&m[298]&m[299]))&~BiasedRNG[290])|((m[8]&m[296]&m[297]&m[298]&~m[299])|(m[8]&m[296]&m[297]&~m[298]&m[299])|(m[8]&m[296]&~m[297]&m[298]&m[299])|(m[8]&~m[296]&m[297]&m[298]&m[299])|(~m[8]&m[296]&m[297]&m[298]&m[299])|(m[8]&m[296]&m[297]&m[298]&m[299]))):InitCond[561];
    m[67] = run?((((m[8]&m[300]&~m[301]&~m[302]&~m[303])|(m[8]&~m[300]&m[301]&~m[302]&~m[303])|(~m[8]&m[300]&m[301]&~m[302]&~m[303])|(m[8]&~m[300]&~m[301]&m[302]&~m[303])|(~m[8]&m[300]&~m[301]&m[302]&~m[303])|(~m[8]&~m[300]&m[301]&m[302]&~m[303])|(m[8]&~m[300]&~m[301]&~m[302]&m[303])|(~m[8]&m[300]&~m[301]&~m[302]&m[303])|(~m[8]&~m[300]&m[301]&~m[302]&m[303])|(~m[8]&~m[300]&~m[301]&m[302]&m[303]))&BiasedRNG[291])|(((m[8]&m[300]&m[301]&~m[302]&~m[303])|(m[8]&m[300]&~m[301]&m[302]&~m[303])|(m[8]&~m[300]&m[301]&m[302]&~m[303])|(~m[8]&m[300]&m[301]&m[302]&~m[303])|(m[8]&m[300]&~m[301]&~m[302]&m[303])|(m[8]&~m[300]&m[301]&~m[302]&m[303])|(~m[8]&m[300]&m[301]&~m[302]&m[303])|(m[8]&~m[300]&~m[301]&m[302]&m[303])|(~m[8]&m[300]&~m[301]&m[302]&m[303])|(~m[8]&~m[300]&m[301]&m[302]&m[303]))&~BiasedRNG[291])|((m[8]&m[300]&m[301]&m[302]&~m[303])|(m[8]&m[300]&m[301]&~m[302]&m[303])|(m[8]&m[300]&~m[301]&m[302]&m[303])|(m[8]&~m[300]&m[301]&m[302]&m[303])|(~m[8]&m[300]&m[301]&m[302]&m[303])|(m[8]&m[300]&m[301]&m[302]&m[303]))):InitCond[562];
    m[68] = run?((((m[9]&m[304]&~m[305]&~m[306]&~m[307])|(m[9]&~m[304]&m[305]&~m[306]&~m[307])|(~m[9]&m[304]&m[305]&~m[306]&~m[307])|(m[9]&~m[304]&~m[305]&m[306]&~m[307])|(~m[9]&m[304]&~m[305]&m[306]&~m[307])|(~m[9]&~m[304]&m[305]&m[306]&~m[307])|(m[9]&~m[304]&~m[305]&~m[306]&m[307])|(~m[9]&m[304]&~m[305]&~m[306]&m[307])|(~m[9]&~m[304]&m[305]&~m[306]&m[307])|(~m[9]&~m[304]&~m[305]&m[306]&m[307]))&BiasedRNG[292])|(((m[9]&m[304]&m[305]&~m[306]&~m[307])|(m[9]&m[304]&~m[305]&m[306]&~m[307])|(m[9]&~m[304]&m[305]&m[306]&~m[307])|(~m[9]&m[304]&m[305]&m[306]&~m[307])|(m[9]&m[304]&~m[305]&~m[306]&m[307])|(m[9]&~m[304]&m[305]&~m[306]&m[307])|(~m[9]&m[304]&m[305]&~m[306]&m[307])|(m[9]&~m[304]&~m[305]&m[306]&m[307])|(~m[9]&m[304]&~m[305]&m[306]&m[307])|(~m[9]&~m[304]&m[305]&m[306]&m[307]))&~BiasedRNG[292])|((m[9]&m[304]&m[305]&m[306]&~m[307])|(m[9]&m[304]&m[305]&~m[306]&m[307])|(m[9]&m[304]&~m[305]&m[306]&m[307])|(m[9]&~m[304]&m[305]&m[306]&m[307])|(~m[9]&m[304]&m[305]&m[306]&m[307])|(m[9]&m[304]&m[305]&m[306]&m[307]))):InitCond[563];
    m[69] = run?((((m[9]&m[308]&~m[309]&~m[310]&~m[311])|(m[9]&~m[308]&m[309]&~m[310]&~m[311])|(~m[9]&m[308]&m[309]&~m[310]&~m[311])|(m[9]&~m[308]&~m[309]&m[310]&~m[311])|(~m[9]&m[308]&~m[309]&m[310]&~m[311])|(~m[9]&~m[308]&m[309]&m[310]&~m[311])|(m[9]&~m[308]&~m[309]&~m[310]&m[311])|(~m[9]&m[308]&~m[309]&~m[310]&m[311])|(~m[9]&~m[308]&m[309]&~m[310]&m[311])|(~m[9]&~m[308]&~m[309]&m[310]&m[311]))&BiasedRNG[293])|(((m[9]&m[308]&m[309]&~m[310]&~m[311])|(m[9]&m[308]&~m[309]&m[310]&~m[311])|(m[9]&~m[308]&m[309]&m[310]&~m[311])|(~m[9]&m[308]&m[309]&m[310]&~m[311])|(m[9]&m[308]&~m[309]&~m[310]&m[311])|(m[9]&~m[308]&m[309]&~m[310]&m[311])|(~m[9]&m[308]&m[309]&~m[310]&m[311])|(m[9]&~m[308]&~m[309]&m[310]&m[311])|(~m[9]&m[308]&~m[309]&m[310]&m[311])|(~m[9]&~m[308]&m[309]&m[310]&m[311]))&~BiasedRNG[293])|((m[9]&m[308]&m[309]&m[310]&~m[311])|(m[9]&m[308]&m[309]&~m[310]&m[311])|(m[9]&m[308]&~m[309]&m[310]&m[311])|(m[9]&~m[308]&m[309]&m[310]&m[311])|(~m[9]&m[308]&m[309]&m[310]&m[311])|(m[9]&m[308]&m[309]&m[310]&m[311]))):InitCond[564];
    m[70] = run?((((m[9]&m[312]&~m[313]&~m[314]&~m[315])|(m[9]&~m[312]&m[313]&~m[314]&~m[315])|(~m[9]&m[312]&m[313]&~m[314]&~m[315])|(m[9]&~m[312]&~m[313]&m[314]&~m[315])|(~m[9]&m[312]&~m[313]&m[314]&~m[315])|(~m[9]&~m[312]&m[313]&m[314]&~m[315])|(m[9]&~m[312]&~m[313]&~m[314]&m[315])|(~m[9]&m[312]&~m[313]&~m[314]&m[315])|(~m[9]&~m[312]&m[313]&~m[314]&m[315])|(~m[9]&~m[312]&~m[313]&m[314]&m[315]))&BiasedRNG[294])|(((m[9]&m[312]&m[313]&~m[314]&~m[315])|(m[9]&m[312]&~m[313]&m[314]&~m[315])|(m[9]&~m[312]&m[313]&m[314]&~m[315])|(~m[9]&m[312]&m[313]&m[314]&~m[315])|(m[9]&m[312]&~m[313]&~m[314]&m[315])|(m[9]&~m[312]&m[313]&~m[314]&m[315])|(~m[9]&m[312]&m[313]&~m[314]&m[315])|(m[9]&~m[312]&~m[313]&m[314]&m[315])|(~m[9]&m[312]&~m[313]&m[314]&m[315])|(~m[9]&~m[312]&m[313]&m[314]&m[315]))&~BiasedRNG[294])|((m[9]&m[312]&m[313]&m[314]&~m[315])|(m[9]&m[312]&m[313]&~m[314]&m[315])|(m[9]&m[312]&~m[313]&m[314]&m[315])|(m[9]&~m[312]&m[313]&m[314]&m[315])|(~m[9]&m[312]&m[313]&m[314]&m[315])|(m[9]&m[312]&m[313]&m[314]&m[315]))):InitCond[565];
    m[71] = run?((((m[9]&m[316]&~m[317]&~m[318]&~m[319])|(m[9]&~m[316]&m[317]&~m[318]&~m[319])|(~m[9]&m[316]&m[317]&~m[318]&~m[319])|(m[9]&~m[316]&~m[317]&m[318]&~m[319])|(~m[9]&m[316]&~m[317]&m[318]&~m[319])|(~m[9]&~m[316]&m[317]&m[318]&~m[319])|(m[9]&~m[316]&~m[317]&~m[318]&m[319])|(~m[9]&m[316]&~m[317]&~m[318]&m[319])|(~m[9]&~m[316]&m[317]&~m[318]&m[319])|(~m[9]&~m[316]&~m[317]&m[318]&m[319]))&BiasedRNG[295])|(((m[9]&m[316]&m[317]&~m[318]&~m[319])|(m[9]&m[316]&~m[317]&m[318]&~m[319])|(m[9]&~m[316]&m[317]&m[318]&~m[319])|(~m[9]&m[316]&m[317]&m[318]&~m[319])|(m[9]&m[316]&~m[317]&~m[318]&m[319])|(m[9]&~m[316]&m[317]&~m[318]&m[319])|(~m[9]&m[316]&m[317]&~m[318]&m[319])|(m[9]&~m[316]&~m[317]&m[318]&m[319])|(~m[9]&m[316]&~m[317]&m[318]&m[319])|(~m[9]&~m[316]&m[317]&m[318]&m[319]))&~BiasedRNG[295])|((m[9]&m[316]&m[317]&m[318]&~m[319])|(m[9]&m[316]&m[317]&~m[318]&m[319])|(m[9]&m[316]&~m[317]&m[318]&m[319])|(m[9]&~m[316]&m[317]&m[318]&m[319])|(~m[9]&m[316]&m[317]&m[318]&m[319])|(m[9]&m[316]&m[317]&m[318]&m[319]))):InitCond[566];
    m[72] = run?((((m[10]&m[320]&~m[321]&~m[322]&~m[323])|(m[10]&~m[320]&m[321]&~m[322]&~m[323])|(~m[10]&m[320]&m[321]&~m[322]&~m[323])|(m[10]&~m[320]&~m[321]&m[322]&~m[323])|(~m[10]&m[320]&~m[321]&m[322]&~m[323])|(~m[10]&~m[320]&m[321]&m[322]&~m[323])|(m[10]&~m[320]&~m[321]&~m[322]&m[323])|(~m[10]&m[320]&~m[321]&~m[322]&m[323])|(~m[10]&~m[320]&m[321]&~m[322]&m[323])|(~m[10]&~m[320]&~m[321]&m[322]&m[323]))&BiasedRNG[296])|(((m[10]&m[320]&m[321]&~m[322]&~m[323])|(m[10]&m[320]&~m[321]&m[322]&~m[323])|(m[10]&~m[320]&m[321]&m[322]&~m[323])|(~m[10]&m[320]&m[321]&m[322]&~m[323])|(m[10]&m[320]&~m[321]&~m[322]&m[323])|(m[10]&~m[320]&m[321]&~m[322]&m[323])|(~m[10]&m[320]&m[321]&~m[322]&m[323])|(m[10]&~m[320]&~m[321]&m[322]&m[323])|(~m[10]&m[320]&~m[321]&m[322]&m[323])|(~m[10]&~m[320]&m[321]&m[322]&m[323]))&~BiasedRNG[296])|((m[10]&m[320]&m[321]&m[322]&~m[323])|(m[10]&m[320]&m[321]&~m[322]&m[323])|(m[10]&m[320]&~m[321]&m[322]&m[323])|(m[10]&~m[320]&m[321]&m[322]&m[323])|(~m[10]&m[320]&m[321]&m[322]&m[323])|(m[10]&m[320]&m[321]&m[322]&m[323]))):InitCond[567];
    m[73] = run?((((m[10]&m[324]&~m[325]&~m[326]&~m[327])|(m[10]&~m[324]&m[325]&~m[326]&~m[327])|(~m[10]&m[324]&m[325]&~m[326]&~m[327])|(m[10]&~m[324]&~m[325]&m[326]&~m[327])|(~m[10]&m[324]&~m[325]&m[326]&~m[327])|(~m[10]&~m[324]&m[325]&m[326]&~m[327])|(m[10]&~m[324]&~m[325]&~m[326]&m[327])|(~m[10]&m[324]&~m[325]&~m[326]&m[327])|(~m[10]&~m[324]&m[325]&~m[326]&m[327])|(~m[10]&~m[324]&~m[325]&m[326]&m[327]))&BiasedRNG[297])|(((m[10]&m[324]&m[325]&~m[326]&~m[327])|(m[10]&m[324]&~m[325]&m[326]&~m[327])|(m[10]&~m[324]&m[325]&m[326]&~m[327])|(~m[10]&m[324]&m[325]&m[326]&~m[327])|(m[10]&m[324]&~m[325]&~m[326]&m[327])|(m[10]&~m[324]&m[325]&~m[326]&m[327])|(~m[10]&m[324]&m[325]&~m[326]&m[327])|(m[10]&~m[324]&~m[325]&m[326]&m[327])|(~m[10]&m[324]&~m[325]&m[326]&m[327])|(~m[10]&~m[324]&m[325]&m[326]&m[327]))&~BiasedRNG[297])|((m[10]&m[324]&m[325]&m[326]&~m[327])|(m[10]&m[324]&m[325]&~m[326]&m[327])|(m[10]&m[324]&~m[325]&m[326]&m[327])|(m[10]&~m[324]&m[325]&m[326]&m[327])|(~m[10]&m[324]&m[325]&m[326]&m[327])|(m[10]&m[324]&m[325]&m[326]&m[327]))):InitCond[568];
    m[74] = run?((((m[10]&m[328]&~m[329]&~m[330]&~m[331])|(m[10]&~m[328]&m[329]&~m[330]&~m[331])|(~m[10]&m[328]&m[329]&~m[330]&~m[331])|(m[10]&~m[328]&~m[329]&m[330]&~m[331])|(~m[10]&m[328]&~m[329]&m[330]&~m[331])|(~m[10]&~m[328]&m[329]&m[330]&~m[331])|(m[10]&~m[328]&~m[329]&~m[330]&m[331])|(~m[10]&m[328]&~m[329]&~m[330]&m[331])|(~m[10]&~m[328]&m[329]&~m[330]&m[331])|(~m[10]&~m[328]&~m[329]&m[330]&m[331]))&BiasedRNG[298])|(((m[10]&m[328]&m[329]&~m[330]&~m[331])|(m[10]&m[328]&~m[329]&m[330]&~m[331])|(m[10]&~m[328]&m[329]&m[330]&~m[331])|(~m[10]&m[328]&m[329]&m[330]&~m[331])|(m[10]&m[328]&~m[329]&~m[330]&m[331])|(m[10]&~m[328]&m[329]&~m[330]&m[331])|(~m[10]&m[328]&m[329]&~m[330]&m[331])|(m[10]&~m[328]&~m[329]&m[330]&m[331])|(~m[10]&m[328]&~m[329]&m[330]&m[331])|(~m[10]&~m[328]&m[329]&m[330]&m[331]))&~BiasedRNG[298])|((m[10]&m[328]&m[329]&m[330]&~m[331])|(m[10]&m[328]&m[329]&~m[330]&m[331])|(m[10]&m[328]&~m[329]&m[330]&m[331])|(m[10]&~m[328]&m[329]&m[330]&m[331])|(~m[10]&m[328]&m[329]&m[330]&m[331])|(m[10]&m[328]&m[329]&m[330]&m[331]))):InitCond[569];
    m[75] = run?((((m[10]&m[332]&~m[333]&~m[334]&~m[335])|(m[10]&~m[332]&m[333]&~m[334]&~m[335])|(~m[10]&m[332]&m[333]&~m[334]&~m[335])|(m[10]&~m[332]&~m[333]&m[334]&~m[335])|(~m[10]&m[332]&~m[333]&m[334]&~m[335])|(~m[10]&~m[332]&m[333]&m[334]&~m[335])|(m[10]&~m[332]&~m[333]&~m[334]&m[335])|(~m[10]&m[332]&~m[333]&~m[334]&m[335])|(~m[10]&~m[332]&m[333]&~m[334]&m[335])|(~m[10]&~m[332]&~m[333]&m[334]&m[335]))&BiasedRNG[299])|(((m[10]&m[332]&m[333]&~m[334]&~m[335])|(m[10]&m[332]&~m[333]&m[334]&~m[335])|(m[10]&~m[332]&m[333]&m[334]&~m[335])|(~m[10]&m[332]&m[333]&m[334]&~m[335])|(m[10]&m[332]&~m[333]&~m[334]&m[335])|(m[10]&~m[332]&m[333]&~m[334]&m[335])|(~m[10]&m[332]&m[333]&~m[334]&m[335])|(m[10]&~m[332]&~m[333]&m[334]&m[335])|(~m[10]&m[332]&~m[333]&m[334]&m[335])|(~m[10]&~m[332]&m[333]&m[334]&m[335]))&~BiasedRNG[299])|((m[10]&m[332]&m[333]&m[334]&~m[335])|(m[10]&m[332]&m[333]&~m[334]&m[335])|(m[10]&m[332]&~m[333]&m[334]&m[335])|(m[10]&~m[332]&m[333]&m[334]&m[335])|(~m[10]&m[332]&m[333]&m[334]&m[335])|(m[10]&m[332]&m[333]&m[334]&m[335]))):InitCond[570];
    m[76] = run?((((m[11]&m[336]&~m[337]&~m[338]&~m[339])|(m[11]&~m[336]&m[337]&~m[338]&~m[339])|(~m[11]&m[336]&m[337]&~m[338]&~m[339])|(m[11]&~m[336]&~m[337]&m[338]&~m[339])|(~m[11]&m[336]&~m[337]&m[338]&~m[339])|(~m[11]&~m[336]&m[337]&m[338]&~m[339])|(m[11]&~m[336]&~m[337]&~m[338]&m[339])|(~m[11]&m[336]&~m[337]&~m[338]&m[339])|(~m[11]&~m[336]&m[337]&~m[338]&m[339])|(~m[11]&~m[336]&~m[337]&m[338]&m[339]))&BiasedRNG[300])|(((m[11]&m[336]&m[337]&~m[338]&~m[339])|(m[11]&m[336]&~m[337]&m[338]&~m[339])|(m[11]&~m[336]&m[337]&m[338]&~m[339])|(~m[11]&m[336]&m[337]&m[338]&~m[339])|(m[11]&m[336]&~m[337]&~m[338]&m[339])|(m[11]&~m[336]&m[337]&~m[338]&m[339])|(~m[11]&m[336]&m[337]&~m[338]&m[339])|(m[11]&~m[336]&~m[337]&m[338]&m[339])|(~m[11]&m[336]&~m[337]&m[338]&m[339])|(~m[11]&~m[336]&m[337]&m[338]&m[339]))&~BiasedRNG[300])|((m[11]&m[336]&m[337]&m[338]&~m[339])|(m[11]&m[336]&m[337]&~m[338]&m[339])|(m[11]&m[336]&~m[337]&m[338]&m[339])|(m[11]&~m[336]&m[337]&m[338]&m[339])|(~m[11]&m[336]&m[337]&m[338]&m[339])|(m[11]&m[336]&m[337]&m[338]&m[339]))):InitCond[571];
    m[77] = run?((((m[11]&m[340]&~m[341]&~m[342]&~m[343])|(m[11]&~m[340]&m[341]&~m[342]&~m[343])|(~m[11]&m[340]&m[341]&~m[342]&~m[343])|(m[11]&~m[340]&~m[341]&m[342]&~m[343])|(~m[11]&m[340]&~m[341]&m[342]&~m[343])|(~m[11]&~m[340]&m[341]&m[342]&~m[343])|(m[11]&~m[340]&~m[341]&~m[342]&m[343])|(~m[11]&m[340]&~m[341]&~m[342]&m[343])|(~m[11]&~m[340]&m[341]&~m[342]&m[343])|(~m[11]&~m[340]&~m[341]&m[342]&m[343]))&BiasedRNG[301])|(((m[11]&m[340]&m[341]&~m[342]&~m[343])|(m[11]&m[340]&~m[341]&m[342]&~m[343])|(m[11]&~m[340]&m[341]&m[342]&~m[343])|(~m[11]&m[340]&m[341]&m[342]&~m[343])|(m[11]&m[340]&~m[341]&~m[342]&m[343])|(m[11]&~m[340]&m[341]&~m[342]&m[343])|(~m[11]&m[340]&m[341]&~m[342]&m[343])|(m[11]&~m[340]&~m[341]&m[342]&m[343])|(~m[11]&m[340]&~m[341]&m[342]&m[343])|(~m[11]&~m[340]&m[341]&m[342]&m[343]))&~BiasedRNG[301])|((m[11]&m[340]&m[341]&m[342]&~m[343])|(m[11]&m[340]&m[341]&~m[342]&m[343])|(m[11]&m[340]&~m[341]&m[342]&m[343])|(m[11]&~m[340]&m[341]&m[342]&m[343])|(~m[11]&m[340]&m[341]&m[342]&m[343])|(m[11]&m[340]&m[341]&m[342]&m[343]))):InitCond[572];
    m[78] = run?((((m[11]&m[344]&~m[345]&~m[346]&~m[347])|(m[11]&~m[344]&m[345]&~m[346]&~m[347])|(~m[11]&m[344]&m[345]&~m[346]&~m[347])|(m[11]&~m[344]&~m[345]&m[346]&~m[347])|(~m[11]&m[344]&~m[345]&m[346]&~m[347])|(~m[11]&~m[344]&m[345]&m[346]&~m[347])|(m[11]&~m[344]&~m[345]&~m[346]&m[347])|(~m[11]&m[344]&~m[345]&~m[346]&m[347])|(~m[11]&~m[344]&m[345]&~m[346]&m[347])|(~m[11]&~m[344]&~m[345]&m[346]&m[347]))&BiasedRNG[302])|(((m[11]&m[344]&m[345]&~m[346]&~m[347])|(m[11]&m[344]&~m[345]&m[346]&~m[347])|(m[11]&~m[344]&m[345]&m[346]&~m[347])|(~m[11]&m[344]&m[345]&m[346]&~m[347])|(m[11]&m[344]&~m[345]&~m[346]&m[347])|(m[11]&~m[344]&m[345]&~m[346]&m[347])|(~m[11]&m[344]&m[345]&~m[346]&m[347])|(m[11]&~m[344]&~m[345]&m[346]&m[347])|(~m[11]&m[344]&~m[345]&m[346]&m[347])|(~m[11]&~m[344]&m[345]&m[346]&m[347]))&~BiasedRNG[302])|((m[11]&m[344]&m[345]&m[346]&~m[347])|(m[11]&m[344]&m[345]&~m[346]&m[347])|(m[11]&m[344]&~m[345]&m[346]&m[347])|(m[11]&~m[344]&m[345]&m[346]&m[347])|(~m[11]&m[344]&m[345]&m[346]&m[347])|(m[11]&m[344]&m[345]&m[346]&m[347]))):InitCond[573];
    m[79] = run?((((m[11]&m[348]&~m[349]&~m[350]&~m[351])|(m[11]&~m[348]&m[349]&~m[350]&~m[351])|(~m[11]&m[348]&m[349]&~m[350]&~m[351])|(m[11]&~m[348]&~m[349]&m[350]&~m[351])|(~m[11]&m[348]&~m[349]&m[350]&~m[351])|(~m[11]&~m[348]&m[349]&m[350]&~m[351])|(m[11]&~m[348]&~m[349]&~m[350]&m[351])|(~m[11]&m[348]&~m[349]&~m[350]&m[351])|(~m[11]&~m[348]&m[349]&~m[350]&m[351])|(~m[11]&~m[348]&~m[349]&m[350]&m[351]))&BiasedRNG[303])|(((m[11]&m[348]&m[349]&~m[350]&~m[351])|(m[11]&m[348]&~m[349]&m[350]&~m[351])|(m[11]&~m[348]&m[349]&m[350]&~m[351])|(~m[11]&m[348]&m[349]&m[350]&~m[351])|(m[11]&m[348]&~m[349]&~m[350]&m[351])|(m[11]&~m[348]&m[349]&~m[350]&m[351])|(~m[11]&m[348]&m[349]&~m[350]&m[351])|(m[11]&~m[348]&~m[349]&m[350]&m[351])|(~m[11]&m[348]&~m[349]&m[350]&m[351])|(~m[11]&~m[348]&m[349]&m[350]&m[351]))&~BiasedRNG[303])|((m[11]&m[348]&m[349]&m[350]&~m[351])|(m[11]&m[348]&m[349]&~m[350]&m[351])|(m[11]&m[348]&~m[349]&m[350]&m[351])|(m[11]&~m[348]&m[349]&m[350]&m[351])|(~m[11]&m[348]&m[349]&m[350]&m[351])|(m[11]&m[348]&m[349]&m[350]&m[351]))):InitCond[574];
    m[80] = run?((((m[12]&m[352]&~m[353]&~m[354]&~m[355])|(m[12]&~m[352]&m[353]&~m[354]&~m[355])|(~m[12]&m[352]&m[353]&~m[354]&~m[355])|(m[12]&~m[352]&~m[353]&m[354]&~m[355])|(~m[12]&m[352]&~m[353]&m[354]&~m[355])|(~m[12]&~m[352]&m[353]&m[354]&~m[355])|(m[12]&~m[352]&~m[353]&~m[354]&m[355])|(~m[12]&m[352]&~m[353]&~m[354]&m[355])|(~m[12]&~m[352]&m[353]&~m[354]&m[355])|(~m[12]&~m[352]&~m[353]&m[354]&m[355]))&BiasedRNG[304])|(((m[12]&m[352]&m[353]&~m[354]&~m[355])|(m[12]&m[352]&~m[353]&m[354]&~m[355])|(m[12]&~m[352]&m[353]&m[354]&~m[355])|(~m[12]&m[352]&m[353]&m[354]&~m[355])|(m[12]&m[352]&~m[353]&~m[354]&m[355])|(m[12]&~m[352]&m[353]&~m[354]&m[355])|(~m[12]&m[352]&m[353]&~m[354]&m[355])|(m[12]&~m[352]&~m[353]&m[354]&m[355])|(~m[12]&m[352]&~m[353]&m[354]&m[355])|(~m[12]&~m[352]&m[353]&m[354]&m[355]))&~BiasedRNG[304])|((m[12]&m[352]&m[353]&m[354]&~m[355])|(m[12]&m[352]&m[353]&~m[354]&m[355])|(m[12]&m[352]&~m[353]&m[354]&m[355])|(m[12]&~m[352]&m[353]&m[354]&m[355])|(~m[12]&m[352]&m[353]&m[354]&m[355])|(m[12]&m[352]&m[353]&m[354]&m[355]))):InitCond[575];
    m[81] = run?((((m[12]&m[356]&~m[357]&~m[358]&~m[359])|(m[12]&~m[356]&m[357]&~m[358]&~m[359])|(~m[12]&m[356]&m[357]&~m[358]&~m[359])|(m[12]&~m[356]&~m[357]&m[358]&~m[359])|(~m[12]&m[356]&~m[357]&m[358]&~m[359])|(~m[12]&~m[356]&m[357]&m[358]&~m[359])|(m[12]&~m[356]&~m[357]&~m[358]&m[359])|(~m[12]&m[356]&~m[357]&~m[358]&m[359])|(~m[12]&~m[356]&m[357]&~m[358]&m[359])|(~m[12]&~m[356]&~m[357]&m[358]&m[359]))&BiasedRNG[305])|(((m[12]&m[356]&m[357]&~m[358]&~m[359])|(m[12]&m[356]&~m[357]&m[358]&~m[359])|(m[12]&~m[356]&m[357]&m[358]&~m[359])|(~m[12]&m[356]&m[357]&m[358]&~m[359])|(m[12]&m[356]&~m[357]&~m[358]&m[359])|(m[12]&~m[356]&m[357]&~m[358]&m[359])|(~m[12]&m[356]&m[357]&~m[358]&m[359])|(m[12]&~m[356]&~m[357]&m[358]&m[359])|(~m[12]&m[356]&~m[357]&m[358]&m[359])|(~m[12]&~m[356]&m[357]&m[358]&m[359]))&~BiasedRNG[305])|((m[12]&m[356]&m[357]&m[358]&~m[359])|(m[12]&m[356]&m[357]&~m[358]&m[359])|(m[12]&m[356]&~m[357]&m[358]&m[359])|(m[12]&~m[356]&m[357]&m[358]&m[359])|(~m[12]&m[356]&m[357]&m[358]&m[359])|(m[12]&m[356]&m[357]&m[358]&m[359]))):InitCond[576];
    m[82] = run?((((m[12]&m[360]&~m[361]&~m[362]&~m[363])|(m[12]&~m[360]&m[361]&~m[362]&~m[363])|(~m[12]&m[360]&m[361]&~m[362]&~m[363])|(m[12]&~m[360]&~m[361]&m[362]&~m[363])|(~m[12]&m[360]&~m[361]&m[362]&~m[363])|(~m[12]&~m[360]&m[361]&m[362]&~m[363])|(m[12]&~m[360]&~m[361]&~m[362]&m[363])|(~m[12]&m[360]&~m[361]&~m[362]&m[363])|(~m[12]&~m[360]&m[361]&~m[362]&m[363])|(~m[12]&~m[360]&~m[361]&m[362]&m[363]))&BiasedRNG[306])|(((m[12]&m[360]&m[361]&~m[362]&~m[363])|(m[12]&m[360]&~m[361]&m[362]&~m[363])|(m[12]&~m[360]&m[361]&m[362]&~m[363])|(~m[12]&m[360]&m[361]&m[362]&~m[363])|(m[12]&m[360]&~m[361]&~m[362]&m[363])|(m[12]&~m[360]&m[361]&~m[362]&m[363])|(~m[12]&m[360]&m[361]&~m[362]&m[363])|(m[12]&~m[360]&~m[361]&m[362]&m[363])|(~m[12]&m[360]&~m[361]&m[362]&m[363])|(~m[12]&~m[360]&m[361]&m[362]&m[363]))&~BiasedRNG[306])|((m[12]&m[360]&m[361]&m[362]&~m[363])|(m[12]&m[360]&m[361]&~m[362]&m[363])|(m[12]&m[360]&~m[361]&m[362]&m[363])|(m[12]&~m[360]&m[361]&m[362]&m[363])|(~m[12]&m[360]&m[361]&m[362]&m[363])|(m[12]&m[360]&m[361]&m[362]&m[363]))):InitCond[577];
    m[83] = run?((((m[12]&m[364]&~m[365]&~m[366]&~m[367])|(m[12]&~m[364]&m[365]&~m[366]&~m[367])|(~m[12]&m[364]&m[365]&~m[366]&~m[367])|(m[12]&~m[364]&~m[365]&m[366]&~m[367])|(~m[12]&m[364]&~m[365]&m[366]&~m[367])|(~m[12]&~m[364]&m[365]&m[366]&~m[367])|(m[12]&~m[364]&~m[365]&~m[366]&m[367])|(~m[12]&m[364]&~m[365]&~m[366]&m[367])|(~m[12]&~m[364]&m[365]&~m[366]&m[367])|(~m[12]&~m[364]&~m[365]&m[366]&m[367]))&BiasedRNG[307])|(((m[12]&m[364]&m[365]&~m[366]&~m[367])|(m[12]&m[364]&~m[365]&m[366]&~m[367])|(m[12]&~m[364]&m[365]&m[366]&~m[367])|(~m[12]&m[364]&m[365]&m[366]&~m[367])|(m[12]&m[364]&~m[365]&~m[366]&m[367])|(m[12]&~m[364]&m[365]&~m[366]&m[367])|(~m[12]&m[364]&m[365]&~m[366]&m[367])|(m[12]&~m[364]&~m[365]&m[366]&m[367])|(~m[12]&m[364]&~m[365]&m[366]&m[367])|(~m[12]&~m[364]&m[365]&m[366]&m[367]))&~BiasedRNG[307])|((m[12]&m[364]&m[365]&m[366]&~m[367])|(m[12]&m[364]&m[365]&~m[366]&m[367])|(m[12]&m[364]&~m[365]&m[366]&m[367])|(m[12]&~m[364]&m[365]&m[366]&m[367])|(~m[12]&m[364]&m[365]&m[366]&m[367])|(m[12]&m[364]&m[365]&m[366]&m[367]))):InitCond[578];
    m[84] = run?((((m[13]&m[368]&~m[369]&~m[370]&~m[371])|(m[13]&~m[368]&m[369]&~m[370]&~m[371])|(~m[13]&m[368]&m[369]&~m[370]&~m[371])|(m[13]&~m[368]&~m[369]&m[370]&~m[371])|(~m[13]&m[368]&~m[369]&m[370]&~m[371])|(~m[13]&~m[368]&m[369]&m[370]&~m[371])|(m[13]&~m[368]&~m[369]&~m[370]&m[371])|(~m[13]&m[368]&~m[369]&~m[370]&m[371])|(~m[13]&~m[368]&m[369]&~m[370]&m[371])|(~m[13]&~m[368]&~m[369]&m[370]&m[371]))&BiasedRNG[308])|(((m[13]&m[368]&m[369]&~m[370]&~m[371])|(m[13]&m[368]&~m[369]&m[370]&~m[371])|(m[13]&~m[368]&m[369]&m[370]&~m[371])|(~m[13]&m[368]&m[369]&m[370]&~m[371])|(m[13]&m[368]&~m[369]&~m[370]&m[371])|(m[13]&~m[368]&m[369]&~m[370]&m[371])|(~m[13]&m[368]&m[369]&~m[370]&m[371])|(m[13]&~m[368]&~m[369]&m[370]&m[371])|(~m[13]&m[368]&~m[369]&m[370]&m[371])|(~m[13]&~m[368]&m[369]&m[370]&m[371]))&~BiasedRNG[308])|((m[13]&m[368]&m[369]&m[370]&~m[371])|(m[13]&m[368]&m[369]&~m[370]&m[371])|(m[13]&m[368]&~m[369]&m[370]&m[371])|(m[13]&~m[368]&m[369]&m[370]&m[371])|(~m[13]&m[368]&m[369]&m[370]&m[371])|(m[13]&m[368]&m[369]&m[370]&m[371]))):InitCond[579];
    m[85] = run?((((m[13]&m[372]&~m[373]&~m[374]&~m[375])|(m[13]&~m[372]&m[373]&~m[374]&~m[375])|(~m[13]&m[372]&m[373]&~m[374]&~m[375])|(m[13]&~m[372]&~m[373]&m[374]&~m[375])|(~m[13]&m[372]&~m[373]&m[374]&~m[375])|(~m[13]&~m[372]&m[373]&m[374]&~m[375])|(m[13]&~m[372]&~m[373]&~m[374]&m[375])|(~m[13]&m[372]&~m[373]&~m[374]&m[375])|(~m[13]&~m[372]&m[373]&~m[374]&m[375])|(~m[13]&~m[372]&~m[373]&m[374]&m[375]))&BiasedRNG[309])|(((m[13]&m[372]&m[373]&~m[374]&~m[375])|(m[13]&m[372]&~m[373]&m[374]&~m[375])|(m[13]&~m[372]&m[373]&m[374]&~m[375])|(~m[13]&m[372]&m[373]&m[374]&~m[375])|(m[13]&m[372]&~m[373]&~m[374]&m[375])|(m[13]&~m[372]&m[373]&~m[374]&m[375])|(~m[13]&m[372]&m[373]&~m[374]&m[375])|(m[13]&~m[372]&~m[373]&m[374]&m[375])|(~m[13]&m[372]&~m[373]&m[374]&m[375])|(~m[13]&~m[372]&m[373]&m[374]&m[375]))&~BiasedRNG[309])|((m[13]&m[372]&m[373]&m[374]&~m[375])|(m[13]&m[372]&m[373]&~m[374]&m[375])|(m[13]&m[372]&~m[373]&m[374]&m[375])|(m[13]&~m[372]&m[373]&m[374]&m[375])|(~m[13]&m[372]&m[373]&m[374]&m[375])|(m[13]&m[372]&m[373]&m[374]&m[375]))):InitCond[580];
    m[86] = run?((((m[13]&m[376]&~m[377]&~m[378]&~m[379])|(m[13]&~m[376]&m[377]&~m[378]&~m[379])|(~m[13]&m[376]&m[377]&~m[378]&~m[379])|(m[13]&~m[376]&~m[377]&m[378]&~m[379])|(~m[13]&m[376]&~m[377]&m[378]&~m[379])|(~m[13]&~m[376]&m[377]&m[378]&~m[379])|(m[13]&~m[376]&~m[377]&~m[378]&m[379])|(~m[13]&m[376]&~m[377]&~m[378]&m[379])|(~m[13]&~m[376]&m[377]&~m[378]&m[379])|(~m[13]&~m[376]&~m[377]&m[378]&m[379]))&BiasedRNG[310])|(((m[13]&m[376]&m[377]&~m[378]&~m[379])|(m[13]&m[376]&~m[377]&m[378]&~m[379])|(m[13]&~m[376]&m[377]&m[378]&~m[379])|(~m[13]&m[376]&m[377]&m[378]&~m[379])|(m[13]&m[376]&~m[377]&~m[378]&m[379])|(m[13]&~m[376]&m[377]&~m[378]&m[379])|(~m[13]&m[376]&m[377]&~m[378]&m[379])|(m[13]&~m[376]&~m[377]&m[378]&m[379])|(~m[13]&m[376]&~m[377]&m[378]&m[379])|(~m[13]&~m[376]&m[377]&m[378]&m[379]))&~BiasedRNG[310])|((m[13]&m[376]&m[377]&m[378]&~m[379])|(m[13]&m[376]&m[377]&~m[378]&m[379])|(m[13]&m[376]&~m[377]&m[378]&m[379])|(m[13]&~m[376]&m[377]&m[378]&m[379])|(~m[13]&m[376]&m[377]&m[378]&m[379])|(m[13]&m[376]&m[377]&m[378]&m[379]))):InitCond[581];
    m[87] = run?((((m[13]&m[380]&~m[381]&~m[382]&~m[383])|(m[13]&~m[380]&m[381]&~m[382]&~m[383])|(~m[13]&m[380]&m[381]&~m[382]&~m[383])|(m[13]&~m[380]&~m[381]&m[382]&~m[383])|(~m[13]&m[380]&~m[381]&m[382]&~m[383])|(~m[13]&~m[380]&m[381]&m[382]&~m[383])|(m[13]&~m[380]&~m[381]&~m[382]&m[383])|(~m[13]&m[380]&~m[381]&~m[382]&m[383])|(~m[13]&~m[380]&m[381]&~m[382]&m[383])|(~m[13]&~m[380]&~m[381]&m[382]&m[383]))&BiasedRNG[311])|(((m[13]&m[380]&m[381]&~m[382]&~m[383])|(m[13]&m[380]&~m[381]&m[382]&~m[383])|(m[13]&~m[380]&m[381]&m[382]&~m[383])|(~m[13]&m[380]&m[381]&m[382]&~m[383])|(m[13]&m[380]&~m[381]&~m[382]&m[383])|(m[13]&~m[380]&m[381]&~m[382]&m[383])|(~m[13]&m[380]&m[381]&~m[382]&m[383])|(m[13]&~m[380]&~m[381]&m[382]&m[383])|(~m[13]&m[380]&~m[381]&m[382]&m[383])|(~m[13]&~m[380]&m[381]&m[382]&m[383]))&~BiasedRNG[311])|((m[13]&m[380]&m[381]&m[382]&~m[383])|(m[13]&m[380]&m[381]&~m[382]&m[383])|(m[13]&m[380]&~m[381]&m[382]&m[383])|(m[13]&~m[380]&m[381]&m[382]&m[383])|(~m[13]&m[380]&m[381]&m[382]&m[383])|(m[13]&m[380]&m[381]&m[382]&m[383]))):InitCond[582];
    m[88] = run?((((m[14]&m[384]&~m[385]&~m[386]&~m[387])|(m[14]&~m[384]&m[385]&~m[386]&~m[387])|(~m[14]&m[384]&m[385]&~m[386]&~m[387])|(m[14]&~m[384]&~m[385]&m[386]&~m[387])|(~m[14]&m[384]&~m[385]&m[386]&~m[387])|(~m[14]&~m[384]&m[385]&m[386]&~m[387])|(m[14]&~m[384]&~m[385]&~m[386]&m[387])|(~m[14]&m[384]&~m[385]&~m[386]&m[387])|(~m[14]&~m[384]&m[385]&~m[386]&m[387])|(~m[14]&~m[384]&~m[385]&m[386]&m[387]))&BiasedRNG[312])|(((m[14]&m[384]&m[385]&~m[386]&~m[387])|(m[14]&m[384]&~m[385]&m[386]&~m[387])|(m[14]&~m[384]&m[385]&m[386]&~m[387])|(~m[14]&m[384]&m[385]&m[386]&~m[387])|(m[14]&m[384]&~m[385]&~m[386]&m[387])|(m[14]&~m[384]&m[385]&~m[386]&m[387])|(~m[14]&m[384]&m[385]&~m[386]&m[387])|(m[14]&~m[384]&~m[385]&m[386]&m[387])|(~m[14]&m[384]&~m[385]&m[386]&m[387])|(~m[14]&~m[384]&m[385]&m[386]&m[387]))&~BiasedRNG[312])|((m[14]&m[384]&m[385]&m[386]&~m[387])|(m[14]&m[384]&m[385]&~m[386]&m[387])|(m[14]&m[384]&~m[385]&m[386]&m[387])|(m[14]&~m[384]&m[385]&m[386]&m[387])|(~m[14]&m[384]&m[385]&m[386]&m[387])|(m[14]&m[384]&m[385]&m[386]&m[387]))):InitCond[583];
    m[89] = run?((((m[14]&m[388]&~m[389]&~m[390]&~m[391])|(m[14]&~m[388]&m[389]&~m[390]&~m[391])|(~m[14]&m[388]&m[389]&~m[390]&~m[391])|(m[14]&~m[388]&~m[389]&m[390]&~m[391])|(~m[14]&m[388]&~m[389]&m[390]&~m[391])|(~m[14]&~m[388]&m[389]&m[390]&~m[391])|(m[14]&~m[388]&~m[389]&~m[390]&m[391])|(~m[14]&m[388]&~m[389]&~m[390]&m[391])|(~m[14]&~m[388]&m[389]&~m[390]&m[391])|(~m[14]&~m[388]&~m[389]&m[390]&m[391]))&BiasedRNG[313])|(((m[14]&m[388]&m[389]&~m[390]&~m[391])|(m[14]&m[388]&~m[389]&m[390]&~m[391])|(m[14]&~m[388]&m[389]&m[390]&~m[391])|(~m[14]&m[388]&m[389]&m[390]&~m[391])|(m[14]&m[388]&~m[389]&~m[390]&m[391])|(m[14]&~m[388]&m[389]&~m[390]&m[391])|(~m[14]&m[388]&m[389]&~m[390]&m[391])|(m[14]&~m[388]&~m[389]&m[390]&m[391])|(~m[14]&m[388]&~m[389]&m[390]&m[391])|(~m[14]&~m[388]&m[389]&m[390]&m[391]))&~BiasedRNG[313])|((m[14]&m[388]&m[389]&m[390]&~m[391])|(m[14]&m[388]&m[389]&~m[390]&m[391])|(m[14]&m[388]&~m[389]&m[390]&m[391])|(m[14]&~m[388]&m[389]&m[390]&m[391])|(~m[14]&m[388]&m[389]&m[390]&m[391])|(m[14]&m[388]&m[389]&m[390]&m[391]))):InitCond[584];
    m[90] = run?((((m[14]&m[392]&~m[393]&~m[394]&~m[395])|(m[14]&~m[392]&m[393]&~m[394]&~m[395])|(~m[14]&m[392]&m[393]&~m[394]&~m[395])|(m[14]&~m[392]&~m[393]&m[394]&~m[395])|(~m[14]&m[392]&~m[393]&m[394]&~m[395])|(~m[14]&~m[392]&m[393]&m[394]&~m[395])|(m[14]&~m[392]&~m[393]&~m[394]&m[395])|(~m[14]&m[392]&~m[393]&~m[394]&m[395])|(~m[14]&~m[392]&m[393]&~m[394]&m[395])|(~m[14]&~m[392]&~m[393]&m[394]&m[395]))&BiasedRNG[314])|(((m[14]&m[392]&m[393]&~m[394]&~m[395])|(m[14]&m[392]&~m[393]&m[394]&~m[395])|(m[14]&~m[392]&m[393]&m[394]&~m[395])|(~m[14]&m[392]&m[393]&m[394]&~m[395])|(m[14]&m[392]&~m[393]&~m[394]&m[395])|(m[14]&~m[392]&m[393]&~m[394]&m[395])|(~m[14]&m[392]&m[393]&~m[394]&m[395])|(m[14]&~m[392]&~m[393]&m[394]&m[395])|(~m[14]&m[392]&~m[393]&m[394]&m[395])|(~m[14]&~m[392]&m[393]&m[394]&m[395]))&~BiasedRNG[314])|((m[14]&m[392]&m[393]&m[394]&~m[395])|(m[14]&m[392]&m[393]&~m[394]&m[395])|(m[14]&m[392]&~m[393]&m[394]&m[395])|(m[14]&~m[392]&m[393]&m[394]&m[395])|(~m[14]&m[392]&m[393]&m[394]&m[395])|(m[14]&m[392]&m[393]&m[394]&m[395]))):InitCond[585];
    m[91] = run?((((m[14]&m[396]&~m[397]&~m[398]&~m[399])|(m[14]&~m[396]&m[397]&~m[398]&~m[399])|(~m[14]&m[396]&m[397]&~m[398]&~m[399])|(m[14]&~m[396]&~m[397]&m[398]&~m[399])|(~m[14]&m[396]&~m[397]&m[398]&~m[399])|(~m[14]&~m[396]&m[397]&m[398]&~m[399])|(m[14]&~m[396]&~m[397]&~m[398]&m[399])|(~m[14]&m[396]&~m[397]&~m[398]&m[399])|(~m[14]&~m[396]&m[397]&~m[398]&m[399])|(~m[14]&~m[396]&~m[397]&m[398]&m[399]))&BiasedRNG[315])|(((m[14]&m[396]&m[397]&~m[398]&~m[399])|(m[14]&m[396]&~m[397]&m[398]&~m[399])|(m[14]&~m[396]&m[397]&m[398]&~m[399])|(~m[14]&m[396]&m[397]&m[398]&~m[399])|(m[14]&m[396]&~m[397]&~m[398]&m[399])|(m[14]&~m[396]&m[397]&~m[398]&m[399])|(~m[14]&m[396]&m[397]&~m[398]&m[399])|(m[14]&~m[396]&~m[397]&m[398]&m[399])|(~m[14]&m[396]&~m[397]&m[398]&m[399])|(~m[14]&~m[396]&m[397]&m[398]&m[399]))&~BiasedRNG[315])|((m[14]&m[396]&m[397]&m[398]&~m[399])|(m[14]&m[396]&m[397]&~m[398]&m[399])|(m[14]&m[396]&~m[397]&m[398]&m[399])|(m[14]&~m[396]&m[397]&m[398]&m[399])|(~m[14]&m[396]&m[397]&m[398]&m[399])|(m[14]&m[396]&m[397]&m[398]&m[399]))):InitCond[586];
    m[92] = run?((((m[15]&m[400]&~m[401]&~m[402]&~m[403])|(m[15]&~m[400]&m[401]&~m[402]&~m[403])|(~m[15]&m[400]&m[401]&~m[402]&~m[403])|(m[15]&~m[400]&~m[401]&m[402]&~m[403])|(~m[15]&m[400]&~m[401]&m[402]&~m[403])|(~m[15]&~m[400]&m[401]&m[402]&~m[403])|(m[15]&~m[400]&~m[401]&~m[402]&m[403])|(~m[15]&m[400]&~m[401]&~m[402]&m[403])|(~m[15]&~m[400]&m[401]&~m[402]&m[403])|(~m[15]&~m[400]&~m[401]&m[402]&m[403]))&BiasedRNG[316])|(((m[15]&m[400]&m[401]&~m[402]&~m[403])|(m[15]&m[400]&~m[401]&m[402]&~m[403])|(m[15]&~m[400]&m[401]&m[402]&~m[403])|(~m[15]&m[400]&m[401]&m[402]&~m[403])|(m[15]&m[400]&~m[401]&~m[402]&m[403])|(m[15]&~m[400]&m[401]&~m[402]&m[403])|(~m[15]&m[400]&m[401]&~m[402]&m[403])|(m[15]&~m[400]&~m[401]&m[402]&m[403])|(~m[15]&m[400]&~m[401]&m[402]&m[403])|(~m[15]&~m[400]&m[401]&m[402]&m[403]))&~BiasedRNG[316])|((m[15]&m[400]&m[401]&m[402]&~m[403])|(m[15]&m[400]&m[401]&~m[402]&m[403])|(m[15]&m[400]&~m[401]&m[402]&m[403])|(m[15]&~m[400]&m[401]&m[402]&m[403])|(~m[15]&m[400]&m[401]&m[402]&m[403])|(m[15]&m[400]&m[401]&m[402]&m[403]))):InitCond[587];
    m[93] = run?((((m[15]&m[404]&~m[405]&~m[406]&~m[407])|(m[15]&~m[404]&m[405]&~m[406]&~m[407])|(~m[15]&m[404]&m[405]&~m[406]&~m[407])|(m[15]&~m[404]&~m[405]&m[406]&~m[407])|(~m[15]&m[404]&~m[405]&m[406]&~m[407])|(~m[15]&~m[404]&m[405]&m[406]&~m[407])|(m[15]&~m[404]&~m[405]&~m[406]&m[407])|(~m[15]&m[404]&~m[405]&~m[406]&m[407])|(~m[15]&~m[404]&m[405]&~m[406]&m[407])|(~m[15]&~m[404]&~m[405]&m[406]&m[407]))&BiasedRNG[317])|(((m[15]&m[404]&m[405]&~m[406]&~m[407])|(m[15]&m[404]&~m[405]&m[406]&~m[407])|(m[15]&~m[404]&m[405]&m[406]&~m[407])|(~m[15]&m[404]&m[405]&m[406]&~m[407])|(m[15]&m[404]&~m[405]&~m[406]&m[407])|(m[15]&~m[404]&m[405]&~m[406]&m[407])|(~m[15]&m[404]&m[405]&~m[406]&m[407])|(m[15]&~m[404]&~m[405]&m[406]&m[407])|(~m[15]&m[404]&~m[405]&m[406]&m[407])|(~m[15]&~m[404]&m[405]&m[406]&m[407]))&~BiasedRNG[317])|((m[15]&m[404]&m[405]&m[406]&~m[407])|(m[15]&m[404]&m[405]&~m[406]&m[407])|(m[15]&m[404]&~m[405]&m[406]&m[407])|(m[15]&~m[404]&m[405]&m[406]&m[407])|(~m[15]&m[404]&m[405]&m[406]&m[407])|(m[15]&m[404]&m[405]&m[406]&m[407]))):InitCond[588];
    m[94] = run?((((m[15]&m[408]&~m[409]&~m[410]&~m[411])|(m[15]&~m[408]&m[409]&~m[410]&~m[411])|(~m[15]&m[408]&m[409]&~m[410]&~m[411])|(m[15]&~m[408]&~m[409]&m[410]&~m[411])|(~m[15]&m[408]&~m[409]&m[410]&~m[411])|(~m[15]&~m[408]&m[409]&m[410]&~m[411])|(m[15]&~m[408]&~m[409]&~m[410]&m[411])|(~m[15]&m[408]&~m[409]&~m[410]&m[411])|(~m[15]&~m[408]&m[409]&~m[410]&m[411])|(~m[15]&~m[408]&~m[409]&m[410]&m[411]))&BiasedRNG[318])|(((m[15]&m[408]&m[409]&~m[410]&~m[411])|(m[15]&m[408]&~m[409]&m[410]&~m[411])|(m[15]&~m[408]&m[409]&m[410]&~m[411])|(~m[15]&m[408]&m[409]&m[410]&~m[411])|(m[15]&m[408]&~m[409]&~m[410]&m[411])|(m[15]&~m[408]&m[409]&~m[410]&m[411])|(~m[15]&m[408]&m[409]&~m[410]&m[411])|(m[15]&~m[408]&~m[409]&m[410]&m[411])|(~m[15]&m[408]&~m[409]&m[410]&m[411])|(~m[15]&~m[408]&m[409]&m[410]&m[411]))&~BiasedRNG[318])|((m[15]&m[408]&m[409]&m[410]&~m[411])|(m[15]&m[408]&m[409]&~m[410]&m[411])|(m[15]&m[408]&~m[409]&m[410]&m[411])|(m[15]&~m[408]&m[409]&m[410]&m[411])|(~m[15]&m[408]&m[409]&m[410]&m[411])|(m[15]&m[408]&m[409]&m[410]&m[411]))):InitCond[589];
    m[95] = run?((((m[15]&m[412]&~m[413]&~m[414]&~m[415])|(m[15]&~m[412]&m[413]&~m[414]&~m[415])|(~m[15]&m[412]&m[413]&~m[414]&~m[415])|(m[15]&~m[412]&~m[413]&m[414]&~m[415])|(~m[15]&m[412]&~m[413]&m[414]&~m[415])|(~m[15]&~m[412]&m[413]&m[414]&~m[415])|(m[15]&~m[412]&~m[413]&~m[414]&m[415])|(~m[15]&m[412]&~m[413]&~m[414]&m[415])|(~m[15]&~m[412]&m[413]&~m[414]&m[415])|(~m[15]&~m[412]&~m[413]&m[414]&m[415]))&BiasedRNG[319])|(((m[15]&m[412]&m[413]&~m[414]&~m[415])|(m[15]&m[412]&~m[413]&m[414]&~m[415])|(m[15]&~m[412]&m[413]&m[414]&~m[415])|(~m[15]&m[412]&m[413]&m[414]&~m[415])|(m[15]&m[412]&~m[413]&~m[414]&m[415])|(m[15]&~m[412]&m[413]&~m[414]&m[415])|(~m[15]&m[412]&m[413]&~m[414]&m[415])|(m[15]&~m[412]&~m[413]&m[414]&m[415])|(~m[15]&m[412]&~m[413]&m[414]&m[415])|(~m[15]&~m[412]&m[413]&m[414]&m[415]))&~BiasedRNG[319])|((m[15]&m[412]&m[413]&m[414]&~m[415])|(m[15]&m[412]&m[413]&~m[414]&m[415])|(m[15]&m[412]&~m[413]&m[414]&m[415])|(m[15]&~m[412]&m[413]&m[414]&m[415])|(~m[15]&m[412]&m[413]&m[414]&m[415])|(m[15]&m[412]&m[413]&m[414]&m[415]))):InitCond[590];
    m[96] = run?((((m[16]&m[416]&~m[417]&~m[418]&~m[419])|(m[16]&~m[416]&m[417]&~m[418]&~m[419])|(~m[16]&m[416]&m[417]&~m[418]&~m[419])|(m[16]&~m[416]&~m[417]&m[418]&~m[419])|(~m[16]&m[416]&~m[417]&m[418]&~m[419])|(~m[16]&~m[416]&m[417]&m[418]&~m[419])|(m[16]&~m[416]&~m[417]&~m[418]&m[419])|(~m[16]&m[416]&~m[417]&~m[418]&m[419])|(~m[16]&~m[416]&m[417]&~m[418]&m[419])|(~m[16]&~m[416]&~m[417]&m[418]&m[419]))&BiasedRNG[320])|(((m[16]&m[416]&m[417]&~m[418]&~m[419])|(m[16]&m[416]&~m[417]&m[418]&~m[419])|(m[16]&~m[416]&m[417]&m[418]&~m[419])|(~m[16]&m[416]&m[417]&m[418]&~m[419])|(m[16]&m[416]&~m[417]&~m[418]&m[419])|(m[16]&~m[416]&m[417]&~m[418]&m[419])|(~m[16]&m[416]&m[417]&~m[418]&m[419])|(m[16]&~m[416]&~m[417]&m[418]&m[419])|(~m[16]&m[416]&~m[417]&m[418]&m[419])|(~m[16]&~m[416]&m[417]&m[418]&m[419]))&~BiasedRNG[320])|((m[16]&m[416]&m[417]&m[418]&~m[419])|(m[16]&m[416]&m[417]&~m[418]&m[419])|(m[16]&m[416]&~m[417]&m[418]&m[419])|(m[16]&~m[416]&m[417]&m[418]&m[419])|(~m[16]&m[416]&m[417]&m[418]&m[419])|(m[16]&m[416]&m[417]&m[418]&m[419]))):InitCond[591];
    m[97] = run?((((m[16]&m[420]&~m[421]&~m[422]&~m[423])|(m[16]&~m[420]&m[421]&~m[422]&~m[423])|(~m[16]&m[420]&m[421]&~m[422]&~m[423])|(m[16]&~m[420]&~m[421]&m[422]&~m[423])|(~m[16]&m[420]&~m[421]&m[422]&~m[423])|(~m[16]&~m[420]&m[421]&m[422]&~m[423])|(m[16]&~m[420]&~m[421]&~m[422]&m[423])|(~m[16]&m[420]&~m[421]&~m[422]&m[423])|(~m[16]&~m[420]&m[421]&~m[422]&m[423])|(~m[16]&~m[420]&~m[421]&m[422]&m[423]))&BiasedRNG[321])|(((m[16]&m[420]&m[421]&~m[422]&~m[423])|(m[16]&m[420]&~m[421]&m[422]&~m[423])|(m[16]&~m[420]&m[421]&m[422]&~m[423])|(~m[16]&m[420]&m[421]&m[422]&~m[423])|(m[16]&m[420]&~m[421]&~m[422]&m[423])|(m[16]&~m[420]&m[421]&~m[422]&m[423])|(~m[16]&m[420]&m[421]&~m[422]&m[423])|(m[16]&~m[420]&~m[421]&m[422]&m[423])|(~m[16]&m[420]&~m[421]&m[422]&m[423])|(~m[16]&~m[420]&m[421]&m[422]&m[423]))&~BiasedRNG[321])|((m[16]&m[420]&m[421]&m[422]&~m[423])|(m[16]&m[420]&m[421]&~m[422]&m[423])|(m[16]&m[420]&~m[421]&m[422]&m[423])|(m[16]&~m[420]&m[421]&m[422]&m[423])|(~m[16]&m[420]&m[421]&m[422]&m[423])|(m[16]&m[420]&m[421]&m[422]&m[423]))):InitCond[592];
    m[98] = run?((((m[16]&m[424]&~m[425]&~m[426]&~m[427])|(m[16]&~m[424]&m[425]&~m[426]&~m[427])|(~m[16]&m[424]&m[425]&~m[426]&~m[427])|(m[16]&~m[424]&~m[425]&m[426]&~m[427])|(~m[16]&m[424]&~m[425]&m[426]&~m[427])|(~m[16]&~m[424]&m[425]&m[426]&~m[427])|(m[16]&~m[424]&~m[425]&~m[426]&m[427])|(~m[16]&m[424]&~m[425]&~m[426]&m[427])|(~m[16]&~m[424]&m[425]&~m[426]&m[427])|(~m[16]&~m[424]&~m[425]&m[426]&m[427]))&BiasedRNG[322])|(((m[16]&m[424]&m[425]&~m[426]&~m[427])|(m[16]&m[424]&~m[425]&m[426]&~m[427])|(m[16]&~m[424]&m[425]&m[426]&~m[427])|(~m[16]&m[424]&m[425]&m[426]&~m[427])|(m[16]&m[424]&~m[425]&~m[426]&m[427])|(m[16]&~m[424]&m[425]&~m[426]&m[427])|(~m[16]&m[424]&m[425]&~m[426]&m[427])|(m[16]&~m[424]&~m[425]&m[426]&m[427])|(~m[16]&m[424]&~m[425]&m[426]&m[427])|(~m[16]&~m[424]&m[425]&m[426]&m[427]))&~BiasedRNG[322])|((m[16]&m[424]&m[425]&m[426]&~m[427])|(m[16]&m[424]&m[425]&~m[426]&m[427])|(m[16]&m[424]&~m[425]&m[426]&m[427])|(m[16]&~m[424]&m[425]&m[426]&m[427])|(~m[16]&m[424]&m[425]&m[426]&m[427])|(m[16]&m[424]&m[425]&m[426]&m[427]))):InitCond[593];
    m[99] = run?((((m[16]&m[428]&~m[429]&~m[430]&~m[431])|(m[16]&~m[428]&m[429]&~m[430]&~m[431])|(~m[16]&m[428]&m[429]&~m[430]&~m[431])|(m[16]&~m[428]&~m[429]&m[430]&~m[431])|(~m[16]&m[428]&~m[429]&m[430]&~m[431])|(~m[16]&~m[428]&m[429]&m[430]&~m[431])|(m[16]&~m[428]&~m[429]&~m[430]&m[431])|(~m[16]&m[428]&~m[429]&~m[430]&m[431])|(~m[16]&~m[428]&m[429]&~m[430]&m[431])|(~m[16]&~m[428]&~m[429]&m[430]&m[431]))&BiasedRNG[323])|(((m[16]&m[428]&m[429]&~m[430]&~m[431])|(m[16]&m[428]&~m[429]&m[430]&~m[431])|(m[16]&~m[428]&m[429]&m[430]&~m[431])|(~m[16]&m[428]&m[429]&m[430]&~m[431])|(m[16]&m[428]&~m[429]&~m[430]&m[431])|(m[16]&~m[428]&m[429]&~m[430]&m[431])|(~m[16]&m[428]&m[429]&~m[430]&m[431])|(m[16]&~m[428]&~m[429]&m[430]&m[431])|(~m[16]&m[428]&~m[429]&m[430]&m[431])|(~m[16]&~m[428]&m[429]&m[430]&m[431]))&~BiasedRNG[323])|((m[16]&m[428]&m[429]&m[430]&~m[431])|(m[16]&m[428]&m[429]&~m[430]&m[431])|(m[16]&m[428]&~m[429]&m[430]&m[431])|(m[16]&~m[428]&m[429]&m[430]&m[431])|(~m[16]&m[428]&m[429]&m[430]&m[431])|(m[16]&m[428]&m[429]&m[430]&m[431]))):InitCond[594];
    m[100] = run?((((m[17]&m[432]&~m[433]&~m[434]&~m[435])|(m[17]&~m[432]&m[433]&~m[434]&~m[435])|(~m[17]&m[432]&m[433]&~m[434]&~m[435])|(m[17]&~m[432]&~m[433]&m[434]&~m[435])|(~m[17]&m[432]&~m[433]&m[434]&~m[435])|(~m[17]&~m[432]&m[433]&m[434]&~m[435])|(m[17]&~m[432]&~m[433]&~m[434]&m[435])|(~m[17]&m[432]&~m[433]&~m[434]&m[435])|(~m[17]&~m[432]&m[433]&~m[434]&m[435])|(~m[17]&~m[432]&~m[433]&m[434]&m[435]))&BiasedRNG[324])|(((m[17]&m[432]&m[433]&~m[434]&~m[435])|(m[17]&m[432]&~m[433]&m[434]&~m[435])|(m[17]&~m[432]&m[433]&m[434]&~m[435])|(~m[17]&m[432]&m[433]&m[434]&~m[435])|(m[17]&m[432]&~m[433]&~m[434]&m[435])|(m[17]&~m[432]&m[433]&~m[434]&m[435])|(~m[17]&m[432]&m[433]&~m[434]&m[435])|(m[17]&~m[432]&~m[433]&m[434]&m[435])|(~m[17]&m[432]&~m[433]&m[434]&m[435])|(~m[17]&~m[432]&m[433]&m[434]&m[435]))&~BiasedRNG[324])|((m[17]&m[432]&m[433]&m[434]&~m[435])|(m[17]&m[432]&m[433]&~m[434]&m[435])|(m[17]&m[432]&~m[433]&m[434]&m[435])|(m[17]&~m[432]&m[433]&m[434]&m[435])|(~m[17]&m[432]&m[433]&m[434]&m[435])|(m[17]&m[432]&m[433]&m[434]&m[435]))):InitCond[595];
    m[101] = run?((((m[17]&m[436]&~m[437]&~m[438]&~m[439])|(m[17]&~m[436]&m[437]&~m[438]&~m[439])|(~m[17]&m[436]&m[437]&~m[438]&~m[439])|(m[17]&~m[436]&~m[437]&m[438]&~m[439])|(~m[17]&m[436]&~m[437]&m[438]&~m[439])|(~m[17]&~m[436]&m[437]&m[438]&~m[439])|(m[17]&~m[436]&~m[437]&~m[438]&m[439])|(~m[17]&m[436]&~m[437]&~m[438]&m[439])|(~m[17]&~m[436]&m[437]&~m[438]&m[439])|(~m[17]&~m[436]&~m[437]&m[438]&m[439]))&BiasedRNG[325])|(((m[17]&m[436]&m[437]&~m[438]&~m[439])|(m[17]&m[436]&~m[437]&m[438]&~m[439])|(m[17]&~m[436]&m[437]&m[438]&~m[439])|(~m[17]&m[436]&m[437]&m[438]&~m[439])|(m[17]&m[436]&~m[437]&~m[438]&m[439])|(m[17]&~m[436]&m[437]&~m[438]&m[439])|(~m[17]&m[436]&m[437]&~m[438]&m[439])|(m[17]&~m[436]&~m[437]&m[438]&m[439])|(~m[17]&m[436]&~m[437]&m[438]&m[439])|(~m[17]&~m[436]&m[437]&m[438]&m[439]))&~BiasedRNG[325])|((m[17]&m[436]&m[437]&m[438]&~m[439])|(m[17]&m[436]&m[437]&~m[438]&m[439])|(m[17]&m[436]&~m[437]&m[438]&m[439])|(m[17]&~m[436]&m[437]&m[438]&m[439])|(~m[17]&m[436]&m[437]&m[438]&m[439])|(m[17]&m[436]&m[437]&m[438]&m[439]))):InitCond[596];
    m[102] = run?((((m[17]&m[440]&~m[441]&~m[442]&~m[443])|(m[17]&~m[440]&m[441]&~m[442]&~m[443])|(~m[17]&m[440]&m[441]&~m[442]&~m[443])|(m[17]&~m[440]&~m[441]&m[442]&~m[443])|(~m[17]&m[440]&~m[441]&m[442]&~m[443])|(~m[17]&~m[440]&m[441]&m[442]&~m[443])|(m[17]&~m[440]&~m[441]&~m[442]&m[443])|(~m[17]&m[440]&~m[441]&~m[442]&m[443])|(~m[17]&~m[440]&m[441]&~m[442]&m[443])|(~m[17]&~m[440]&~m[441]&m[442]&m[443]))&BiasedRNG[326])|(((m[17]&m[440]&m[441]&~m[442]&~m[443])|(m[17]&m[440]&~m[441]&m[442]&~m[443])|(m[17]&~m[440]&m[441]&m[442]&~m[443])|(~m[17]&m[440]&m[441]&m[442]&~m[443])|(m[17]&m[440]&~m[441]&~m[442]&m[443])|(m[17]&~m[440]&m[441]&~m[442]&m[443])|(~m[17]&m[440]&m[441]&~m[442]&m[443])|(m[17]&~m[440]&~m[441]&m[442]&m[443])|(~m[17]&m[440]&~m[441]&m[442]&m[443])|(~m[17]&~m[440]&m[441]&m[442]&m[443]))&~BiasedRNG[326])|((m[17]&m[440]&m[441]&m[442]&~m[443])|(m[17]&m[440]&m[441]&~m[442]&m[443])|(m[17]&m[440]&~m[441]&m[442]&m[443])|(m[17]&~m[440]&m[441]&m[442]&m[443])|(~m[17]&m[440]&m[441]&m[442]&m[443])|(m[17]&m[440]&m[441]&m[442]&m[443]))):InitCond[597];
    m[103] = run?((((m[17]&m[444]&~m[445]&~m[446]&~m[447])|(m[17]&~m[444]&m[445]&~m[446]&~m[447])|(~m[17]&m[444]&m[445]&~m[446]&~m[447])|(m[17]&~m[444]&~m[445]&m[446]&~m[447])|(~m[17]&m[444]&~m[445]&m[446]&~m[447])|(~m[17]&~m[444]&m[445]&m[446]&~m[447])|(m[17]&~m[444]&~m[445]&~m[446]&m[447])|(~m[17]&m[444]&~m[445]&~m[446]&m[447])|(~m[17]&~m[444]&m[445]&~m[446]&m[447])|(~m[17]&~m[444]&~m[445]&m[446]&m[447]))&BiasedRNG[327])|(((m[17]&m[444]&m[445]&~m[446]&~m[447])|(m[17]&m[444]&~m[445]&m[446]&~m[447])|(m[17]&~m[444]&m[445]&m[446]&~m[447])|(~m[17]&m[444]&m[445]&m[446]&~m[447])|(m[17]&m[444]&~m[445]&~m[446]&m[447])|(m[17]&~m[444]&m[445]&~m[446]&m[447])|(~m[17]&m[444]&m[445]&~m[446]&m[447])|(m[17]&~m[444]&~m[445]&m[446]&m[447])|(~m[17]&m[444]&~m[445]&m[446]&m[447])|(~m[17]&~m[444]&m[445]&m[446]&m[447]))&~BiasedRNG[327])|((m[17]&m[444]&m[445]&m[446]&~m[447])|(m[17]&m[444]&m[445]&~m[446]&m[447])|(m[17]&m[444]&~m[445]&m[446]&m[447])|(m[17]&~m[444]&m[445]&m[446]&m[447])|(~m[17]&m[444]&m[445]&m[446]&m[447])|(m[17]&m[444]&m[445]&m[446]&m[447]))):InitCond[598];
    m[104] = run?((((m[18]&m[448]&~m[449]&~m[450]&~m[451])|(m[18]&~m[448]&m[449]&~m[450]&~m[451])|(~m[18]&m[448]&m[449]&~m[450]&~m[451])|(m[18]&~m[448]&~m[449]&m[450]&~m[451])|(~m[18]&m[448]&~m[449]&m[450]&~m[451])|(~m[18]&~m[448]&m[449]&m[450]&~m[451])|(m[18]&~m[448]&~m[449]&~m[450]&m[451])|(~m[18]&m[448]&~m[449]&~m[450]&m[451])|(~m[18]&~m[448]&m[449]&~m[450]&m[451])|(~m[18]&~m[448]&~m[449]&m[450]&m[451]))&BiasedRNG[328])|(((m[18]&m[448]&m[449]&~m[450]&~m[451])|(m[18]&m[448]&~m[449]&m[450]&~m[451])|(m[18]&~m[448]&m[449]&m[450]&~m[451])|(~m[18]&m[448]&m[449]&m[450]&~m[451])|(m[18]&m[448]&~m[449]&~m[450]&m[451])|(m[18]&~m[448]&m[449]&~m[450]&m[451])|(~m[18]&m[448]&m[449]&~m[450]&m[451])|(m[18]&~m[448]&~m[449]&m[450]&m[451])|(~m[18]&m[448]&~m[449]&m[450]&m[451])|(~m[18]&~m[448]&m[449]&m[450]&m[451]))&~BiasedRNG[328])|((m[18]&m[448]&m[449]&m[450]&~m[451])|(m[18]&m[448]&m[449]&~m[450]&m[451])|(m[18]&m[448]&~m[449]&m[450]&m[451])|(m[18]&~m[448]&m[449]&m[450]&m[451])|(~m[18]&m[448]&m[449]&m[450]&m[451])|(m[18]&m[448]&m[449]&m[450]&m[451]))):InitCond[599];
    m[105] = run?((((m[18]&m[452]&~m[453]&~m[454]&~m[455])|(m[18]&~m[452]&m[453]&~m[454]&~m[455])|(~m[18]&m[452]&m[453]&~m[454]&~m[455])|(m[18]&~m[452]&~m[453]&m[454]&~m[455])|(~m[18]&m[452]&~m[453]&m[454]&~m[455])|(~m[18]&~m[452]&m[453]&m[454]&~m[455])|(m[18]&~m[452]&~m[453]&~m[454]&m[455])|(~m[18]&m[452]&~m[453]&~m[454]&m[455])|(~m[18]&~m[452]&m[453]&~m[454]&m[455])|(~m[18]&~m[452]&~m[453]&m[454]&m[455]))&BiasedRNG[329])|(((m[18]&m[452]&m[453]&~m[454]&~m[455])|(m[18]&m[452]&~m[453]&m[454]&~m[455])|(m[18]&~m[452]&m[453]&m[454]&~m[455])|(~m[18]&m[452]&m[453]&m[454]&~m[455])|(m[18]&m[452]&~m[453]&~m[454]&m[455])|(m[18]&~m[452]&m[453]&~m[454]&m[455])|(~m[18]&m[452]&m[453]&~m[454]&m[455])|(m[18]&~m[452]&~m[453]&m[454]&m[455])|(~m[18]&m[452]&~m[453]&m[454]&m[455])|(~m[18]&~m[452]&m[453]&m[454]&m[455]))&~BiasedRNG[329])|((m[18]&m[452]&m[453]&m[454]&~m[455])|(m[18]&m[452]&m[453]&~m[454]&m[455])|(m[18]&m[452]&~m[453]&m[454]&m[455])|(m[18]&~m[452]&m[453]&m[454]&m[455])|(~m[18]&m[452]&m[453]&m[454]&m[455])|(m[18]&m[452]&m[453]&m[454]&m[455]))):InitCond[600];
    m[106] = run?((((m[18]&m[456]&~m[457]&~m[458]&~m[459])|(m[18]&~m[456]&m[457]&~m[458]&~m[459])|(~m[18]&m[456]&m[457]&~m[458]&~m[459])|(m[18]&~m[456]&~m[457]&m[458]&~m[459])|(~m[18]&m[456]&~m[457]&m[458]&~m[459])|(~m[18]&~m[456]&m[457]&m[458]&~m[459])|(m[18]&~m[456]&~m[457]&~m[458]&m[459])|(~m[18]&m[456]&~m[457]&~m[458]&m[459])|(~m[18]&~m[456]&m[457]&~m[458]&m[459])|(~m[18]&~m[456]&~m[457]&m[458]&m[459]))&BiasedRNG[330])|(((m[18]&m[456]&m[457]&~m[458]&~m[459])|(m[18]&m[456]&~m[457]&m[458]&~m[459])|(m[18]&~m[456]&m[457]&m[458]&~m[459])|(~m[18]&m[456]&m[457]&m[458]&~m[459])|(m[18]&m[456]&~m[457]&~m[458]&m[459])|(m[18]&~m[456]&m[457]&~m[458]&m[459])|(~m[18]&m[456]&m[457]&~m[458]&m[459])|(m[18]&~m[456]&~m[457]&m[458]&m[459])|(~m[18]&m[456]&~m[457]&m[458]&m[459])|(~m[18]&~m[456]&m[457]&m[458]&m[459]))&~BiasedRNG[330])|((m[18]&m[456]&m[457]&m[458]&~m[459])|(m[18]&m[456]&m[457]&~m[458]&m[459])|(m[18]&m[456]&~m[457]&m[458]&m[459])|(m[18]&~m[456]&m[457]&m[458]&m[459])|(~m[18]&m[456]&m[457]&m[458]&m[459])|(m[18]&m[456]&m[457]&m[458]&m[459]))):InitCond[601];
    m[107] = run?((((m[18]&m[460]&~m[461]&~m[462]&~m[463])|(m[18]&~m[460]&m[461]&~m[462]&~m[463])|(~m[18]&m[460]&m[461]&~m[462]&~m[463])|(m[18]&~m[460]&~m[461]&m[462]&~m[463])|(~m[18]&m[460]&~m[461]&m[462]&~m[463])|(~m[18]&~m[460]&m[461]&m[462]&~m[463])|(m[18]&~m[460]&~m[461]&~m[462]&m[463])|(~m[18]&m[460]&~m[461]&~m[462]&m[463])|(~m[18]&~m[460]&m[461]&~m[462]&m[463])|(~m[18]&~m[460]&~m[461]&m[462]&m[463]))&BiasedRNG[331])|(((m[18]&m[460]&m[461]&~m[462]&~m[463])|(m[18]&m[460]&~m[461]&m[462]&~m[463])|(m[18]&~m[460]&m[461]&m[462]&~m[463])|(~m[18]&m[460]&m[461]&m[462]&~m[463])|(m[18]&m[460]&~m[461]&~m[462]&m[463])|(m[18]&~m[460]&m[461]&~m[462]&m[463])|(~m[18]&m[460]&m[461]&~m[462]&m[463])|(m[18]&~m[460]&~m[461]&m[462]&m[463])|(~m[18]&m[460]&~m[461]&m[462]&m[463])|(~m[18]&~m[460]&m[461]&m[462]&m[463]))&~BiasedRNG[331])|((m[18]&m[460]&m[461]&m[462]&~m[463])|(m[18]&m[460]&m[461]&~m[462]&m[463])|(m[18]&m[460]&~m[461]&m[462]&m[463])|(m[18]&~m[460]&m[461]&m[462]&m[463])|(~m[18]&m[460]&m[461]&m[462]&m[463])|(m[18]&m[460]&m[461]&m[462]&m[463]))):InitCond[602];
    m[108] = run?((((m[19]&m[464]&~m[465]&~m[466]&~m[467])|(m[19]&~m[464]&m[465]&~m[466]&~m[467])|(~m[19]&m[464]&m[465]&~m[466]&~m[467])|(m[19]&~m[464]&~m[465]&m[466]&~m[467])|(~m[19]&m[464]&~m[465]&m[466]&~m[467])|(~m[19]&~m[464]&m[465]&m[466]&~m[467])|(m[19]&~m[464]&~m[465]&~m[466]&m[467])|(~m[19]&m[464]&~m[465]&~m[466]&m[467])|(~m[19]&~m[464]&m[465]&~m[466]&m[467])|(~m[19]&~m[464]&~m[465]&m[466]&m[467]))&BiasedRNG[332])|(((m[19]&m[464]&m[465]&~m[466]&~m[467])|(m[19]&m[464]&~m[465]&m[466]&~m[467])|(m[19]&~m[464]&m[465]&m[466]&~m[467])|(~m[19]&m[464]&m[465]&m[466]&~m[467])|(m[19]&m[464]&~m[465]&~m[466]&m[467])|(m[19]&~m[464]&m[465]&~m[466]&m[467])|(~m[19]&m[464]&m[465]&~m[466]&m[467])|(m[19]&~m[464]&~m[465]&m[466]&m[467])|(~m[19]&m[464]&~m[465]&m[466]&m[467])|(~m[19]&~m[464]&m[465]&m[466]&m[467]))&~BiasedRNG[332])|((m[19]&m[464]&m[465]&m[466]&~m[467])|(m[19]&m[464]&m[465]&~m[466]&m[467])|(m[19]&m[464]&~m[465]&m[466]&m[467])|(m[19]&~m[464]&m[465]&m[466]&m[467])|(~m[19]&m[464]&m[465]&m[466]&m[467])|(m[19]&m[464]&m[465]&m[466]&m[467]))):InitCond[603];
    m[109] = run?((((m[19]&m[468]&~m[469]&~m[470]&~m[471])|(m[19]&~m[468]&m[469]&~m[470]&~m[471])|(~m[19]&m[468]&m[469]&~m[470]&~m[471])|(m[19]&~m[468]&~m[469]&m[470]&~m[471])|(~m[19]&m[468]&~m[469]&m[470]&~m[471])|(~m[19]&~m[468]&m[469]&m[470]&~m[471])|(m[19]&~m[468]&~m[469]&~m[470]&m[471])|(~m[19]&m[468]&~m[469]&~m[470]&m[471])|(~m[19]&~m[468]&m[469]&~m[470]&m[471])|(~m[19]&~m[468]&~m[469]&m[470]&m[471]))&BiasedRNG[333])|(((m[19]&m[468]&m[469]&~m[470]&~m[471])|(m[19]&m[468]&~m[469]&m[470]&~m[471])|(m[19]&~m[468]&m[469]&m[470]&~m[471])|(~m[19]&m[468]&m[469]&m[470]&~m[471])|(m[19]&m[468]&~m[469]&~m[470]&m[471])|(m[19]&~m[468]&m[469]&~m[470]&m[471])|(~m[19]&m[468]&m[469]&~m[470]&m[471])|(m[19]&~m[468]&~m[469]&m[470]&m[471])|(~m[19]&m[468]&~m[469]&m[470]&m[471])|(~m[19]&~m[468]&m[469]&m[470]&m[471]))&~BiasedRNG[333])|((m[19]&m[468]&m[469]&m[470]&~m[471])|(m[19]&m[468]&m[469]&~m[470]&m[471])|(m[19]&m[468]&~m[469]&m[470]&m[471])|(m[19]&~m[468]&m[469]&m[470]&m[471])|(~m[19]&m[468]&m[469]&m[470]&m[471])|(m[19]&m[468]&m[469]&m[470]&m[471]))):InitCond[604];
    m[110] = run?((((m[19]&m[472]&~m[473]&~m[474]&~m[475])|(m[19]&~m[472]&m[473]&~m[474]&~m[475])|(~m[19]&m[472]&m[473]&~m[474]&~m[475])|(m[19]&~m[472]&~m[473]&m[474]&~m[475])|(~m[19]&m[472]&~m[473]&m[474]&~m[475])|(~m[19]&~m[472]&m[473]&m[474]&~m[475])|(m[19]&~m[472]&~m[473]&~m[474]&m[475])|(~m[19]&m[472]&~m[473]&~m[474]&m[475])|(~m[19]&~m[472]&m[473]&~m[474]&m[475])|(~m[19]&~m[472]&~m[473]&m[474]&m[475]))&BiasedRNG[334])|(((m[19]&m[472]&m[473]&~m[474]&~m[475])|(m[19]&m[472]&~m[473]&m[474]&~m[475])|(m[19]&~m[472]&m[473]&m[474]&~m[475])|(~m[19]&m[472]&m[473]&m[474]&~m[475])|(m[19]&m[472]&~m[473]&~m[474]&m[475])|(m[19]&~m[472]&m[473]&~m[474]&m[475])|(~m[19]&m[472]&m[473]&~m[474]&m[475])|(m[19]&~m[472]&~m[473]&m[474]&m[475])|(~m[19]&m[472]&~m[473]&m[474]&m[475])|(~m[19]&~m[472]&m[473]&m[474]&m[475]))&~BiasedRNG[334])|((m[19]&m[472]&m[473]&m[474]&~m[475])|(m[19]&m[472]&m[473]&~m[474]&m[475])|(m[19]&m[472]&~m[473]&m[474]&m[475])|(m[19]&~m[472]&m[473]&m[474]&m[475])|(~m[19]&m[472]&m[473]&m[474]&m[475])|(m[19]&m[472]&m[473]&m[474]&m[475]))):InitCond[605];
    m[111] = run?((((m[19]&m[476]&~m[477]&~m[478]&~m[479])|(m[19]&~m[476]&m[477]&~m[478]&~m[479])|(~m[19]&m[476]&m[477]&~m[478]&~m[479])|(m[19]&~m[476]&~m[477]&m[478]&~m[479])|(~m[19]&m[476]&~m[477]&m[478]&~m[479])|(~m[19]&~m[476]&m[477]&m[478]&~m[479])|(m[19]&~m[476]&~m[477]&~m[478]&m[479])|(~m[19]&m[476]&~m[477]&~m[478]&m[479])|(~m[19]&~m[476]&m[477]&~m[478]&m[479])|(~m[19]&~m[476]&~m[477]&m[478]&m[479]))&BiasedRNG[335])|(((m[19]&m[476]&m[477]&~m[478]&~m[479])|(m[19]&m[476]&~m[477]&m[478]&~m[479])|(m[19]&~m[476]&m[477]&m[478]&~m[479])|(~m[19]&m[476]&m[477]&m[478]&~m[479])|(m[19]&m[476]&~m[477]&~m[478]&m[479])|(m[19]&~m[476]&m[477]&~m[478]&m[479])|(~m[19]&m[476]&m[477]&~m[478]&m[479])|(m[19]&~m[476]&~m[477]&m[478]&m[479])|(~m[19]&m[476]&~m[477]&m[478]&m[479])|(~m[19]&~m[476]&m[477]&m[478]&m[479]))&~BiasedRNG[335])|((m[19]&m[476]&m[477]&m[478]&~m[479])|(m[19]&m[476]&m[477]&~m[478]&m[479])|(m[19]&m[476]&~m[477]&m[478]&m[479])|(m[19]&~m[476]&m[477]&m[478]&m[479])|(~m[19]&m[476]&m[477]&m[478]&m[479])|(m[19]&m[476]&m[477]&m[478]&m[479]))):InitCond[606];
    m[112] = run?((((m[20]&m[480]&~m[481]&~m[482]&~m[483])|(m[20]&~m[480]&m[481]&~m[482]&~m[483])|(~m[20]&m[480]&m[481]&~m[482]&~m[483])|(m[20]&~m[480]&~m[481]&m[482]&~m[483])|(~m[20]&m[480]&~m[481]&m[482]&~m[483])|(~m[20]&~m[480]&m[481]&m[482]&~m[483])|(m[20]&~m[480]&~m[481]&~m[482]&m[483])|(~m[20]&m[480]&~m[481]&~m[482]&m[483])|(~m[20]&~m[480]&m[481]&~m[482]&m[483])|(~m[20]&~m[480]&~m[481]&m[482]&m[483]))&BiasedRNG[336])|(((m[20]&m[480]&m[481]&~m[482]&~m[483])|(m[20]&m[480]&~m[481]&m[482]&~m[483])|(m[20]&~m[480]&m[481]&m[482]&~m[483])|(~m[20]&m[480]&m[481]&m[482]&~m[483])|(m[20]&m[480]&~m[481]&~m[482]&m[483])|(m[20]&~m[480]&m[481]&~m[482]&m[483])|(~m[20]&m[480]&m[481]&~m[482]&m[483])|(m[20]&~m[480]&~m[481]&m[482]&m[483])|(~m[20]&m[480]&~m[481]&m[482]&m[483])|(~m[20]&~m[480]&m[481]&m[482]&m[483]))&~BiasedRNG[336])|((m[20]&m[480]&m[481]&m[482]&~m[483])|(m[20]&m[480]&m[481]&~m[482]&m[483])|(m[20]&m[480]&~m[481]&m[482]&m[483])|(m[20]&~m[480]&m[481]&m[482]&m[483])|(~m[20]&m[480]&m[481]&m[482]&m[483])|(m[20]&m[480]&m[481]&m[482]&m[483]))):InitCond[607];
    m[113] = run?((((m[20]&m[484]&~m[485]&~m[486]&~m[487])|(m[20]&~m[484]&m[485]&~m[486]&~m[487])|(~m[20]&m[484]&m[485]&~m[486]&~m[487])|(m[20]&~m[484]&~m[485]&m[486]&~m[487])|(~m[20]&m[484]&~m[485]&m[486]&~m[487])|(~m[20]&~m[484]&m[485]&m[486]&~m[487])|(m[20]&~m[484]&~m[485]&~m[486]&m[487])|(~m[20]&m[484]&~m[485]&~m[486]&m[487])|(~m[20]&~m[484]&m[485]&~m[486]&m[487])|(~m[20]&~m[484]&~m[485]&m[486]&m[487]))&BiasedRNG[337])|(((m[20]&m[484]&m[485]&~m[486]&~m[487])|(m[20]&m[484]&~m[485]&m[486]&~m[487])|(m[20]&~m[484]&m[485]&m[486]&~m[487])|(~m[20]&m[484]&m[485]&m[486]&~m[487])|(m[20]&m[484]&~m[485]&~m[486]&m[487])|(m[20]&~m[484]&m[485]&~m[486]&m[487])|(~m[20]&m[484]&m[485]&~m[486]&m[487])|(m[20]&~m[484]&~m[485]&m[486]&m[487])|(~m[20]&m[484]&~m[485]&m[486]&m[487])|(~m[20]&~m[484]&m[485]&m[486]&m[487]))&~BiasedRNG[337])|((m[20]&m[484]&m[485]&m[486]&~m[487])|(m[20]&m[484]&m[485]&~m[486]&m[487])|(m[20]&m[484]&~m[485]&m[486]&m[487])|(m[20]&~m[484]&m[485]&m[486]&m[487])|(~m[20]&m[484]&m[485]&m[486]&m[487])|(m[20]&m[484]&m[485]&m[486]&m[487]))):InitCond[608];
    m[114] = run?((((m[20]&m[488]&~m[489]&~m[490]&~m[491])|(m[20]&~m[488]&m[489]&~m[490]&~m[491])|(~m[20]&m[488]&m[489]&~m[490]&~m[491])|(m[20]&~m[488]&~m[489]&m[490]&~m[491])|(~m[20]&m[488]&~m[489]&m[490]&~m[491])|(~m[20]&~m[488]&m[489]&m[490]&~m[491])|(m[20]&~m[488]&~m[489]&~m[490]&m[491])|(~m[20]&m[488]&~m[489]&~m[490]&m[491])|(~m[20]&~m[488]&m[489]&~m[490]&m[491])|(~m[20]&~m[488]&~m[489]&m[490]&m[491]))&BiasedRNG[338])|(((m[20]&m[488]&m[489]&~m[490]&~m[491])|(m[20]&m[488]&~m[489]&m[490]&~m[491])|(m[20]&~m[488]&m[489]&m[490]&~m[491])|(~m[20]&m[488]&m[489]&m[490]&~m[491])|(m[20]&m[488]&~m[489]&~m[490]&m[491])|(m[20]&~m[488]&m[489]&~m[490]&m[491])|(~m[20]&m[488]&m[489]&~m[490]&m[491])|(m[20]&~m[488]&~m[489]&m[490]&m[491])|(~m[20]&m[488]&~m[489]&m[490]&m[491])|(~m[20]&~m[488]&m[489]&m[490]&m[491]))&~BiasedRNG[338])|((m[20]&m[488]&m[489]&m[490]&~m[491])|(m[20]&m[488]&m[489]&~m[490]&m[491])|(m[20]&m[488]&~m[489]&m[490]&m[491])|(m[20]&~m[488]&m[489]&m[490]&m[491])|(~m[20]&m[488]&m[489]&m[490]&m[491])|(m[20]&m[488]&m[489]&m[490]&m[491]))):InitCond[609];
    m[115] = run?((((m[20]&m[492]&~m[493]&~m[494]&~m[495])|(m[20]&~m[492]&m[493]&~m[494]&~m[495])|(~m[20]&m[492]&m[493]&~m[494]&~m[495])|(m[20]&~m[492]&~m[493]&m[494]&~m[495])|(~m[20]&m[492]&~m[493]&m[494]&~m[495])|(~m[20]&~m[492]&m[493]&m[494]&~m[495])|(m[20]&~m[492]&~m[493]&~m[494]&m[495])|(~m[20]&m[492]&~m[493]&~m[494]&m[495])|(~m[20]&~m[492]&m[493]&~m[494]&m[495])|(~m[20]&~m[492]&~m[493]&m[494]&m[495]))&BiasedRNG[339])|(((m[20]&m[492]&m[493]&~m[494]&~m[495])|(m[20]&m[492]&~m[493]&m[494]&~m[495])|(m[20]&~m[492]&m[493]&m[494]&~m[495])|(~m[20]&m[492]&m[493]&m[494]&~m[495])|(m[20]&m[492]&~m[493]&~m[494]&m[495])|(m[20]&~m[492]&m[493]&~m[494]&m[495])|(~m[20]&m[492]&m[493]&~m[494]&m[495])|(m[20]&~m[492]&~m[493]&m[494]&m[495])|(~m[20]&m[492]&~m[493]&m[494]&m[495])|(~m[20]&~m[492]&m[493]&m[494]&m[495]))&~BiasedRNG[339])|((m[20]&m[492]&m[493]&m[494]&~m[495])|(m[20]&m[492]&m[493]&~m[494]&m[495])|(m[20]&m[492]&~m[493]&m[494]&m[495])|(m[20]&~m[492]&m[493]&m[494]&m[495])|(~m[20]&m[492]&m[493]&m[494]&m[495])|(m[20]&m[492]&m[493]&m[494]&m[495]))):InitCond[610];
    m[116] = run?((((m[21]&m[496]&~m[497]&~m[498]&~m[499])|(m[21]&~m[496]&m[497]&~m[498]&~m[499])|(~m[21]&m[496]&m[497]&~m[498]&~m[499])|(m[21]&~m[496]&~m[497]&m[498]&~m[499])|(~m[21]&m[496]&~m[497]&m[498]&~m[499])|(~m[21]&~m[496]&m[497]&m[498]&~m[499])|(m[21]&~m[496]&~m[497]&~m[498]&m[499])|(~m[21]&m[496]&~m[497]&~m[498]&m[499])|(~m[21]&~m[496]&m[497]&~m[498]&m[499])|(~m[21]&~m[496]&~m[497]&m[498]&m[499]))&BiasedRNG[340])|(((m[21]&m[496]&m[497]&~m[498]&~m[499])|(m[21]&m[496]&~m[497]&m[498]&~m[499])|(m[21]&~m[496]&m[497]&m[498]&~m[499])|(~m[21]&m[496]&m[497]&m[498]&~m[499])|(m[21]&m[496]&~m[497]&~m[498]&m[499])|(m[21]&~m[496]&m[497]&~m[498]&m[499])|(~m[21]&m[496]&m[497]&~m[498]&m[499])|(m[21]&~m[496]&~m[497]&m[498]&m[499])|(~m[21]&m[496]&~m[497]&m[498]&m[499])|(~m[21]&~m[496]&m[497]&m[498]&m[499]))&~BiasedRNG[340])|((m[21]&m[496]&m[497]&m[498]&~m[499])|(m[21]&m[496]&m[497]&~m[498]&m[499])|(m[21]&m[496]&~m[497]&m[498]&m[499])|(m[21]&~m[496]&m[497]&m[498]&m[499])|(~m[21]&m[496]&m[497]&m[498]&m[499])|(m[21]&m[496]&m[497]&m[498]&m[499]))):InitCond[611];
    m[117] = run?((((m[21]&m[500]&~m[501]&~m[502]&~m[503])|(m[21]&~m[500]&m[501]&~m[502]&~m[503])|(~m[21]&m[500]&m[501]&~m[502]&~m[503])|(m[21]&~m[500]&~m[501]&m[502]&~m[503])|(~m[21]&m[500]&~m[501]&m[502]&~m[503])|(~m[21]&~m[500]&m[501]&m[502]&~m[503])|(m[21]&~m[500]&~m[501]&~m[502]&m[503])|(~m[21]&m[500]&~m[501]&~m[502]&m[503])|(~m[21]&~m[500]&m[501]&~m[502]&m[503])|(~m[21]&~m[500]&~m[501]&m[502]&m[503]))&BiasedRNG[341])|(((m[21]&m[500]&m[501]&~m[502]&~m[503])|(m[21]&m[500]&~m[501]&m[502]&~m[503])|(m[21]&~m[500]&m[501]&m[502]&~m[503])|(~m[21]&m[500]&m[501]&m[502]&~m[503])|(m[21]&m[500]&~m[501]&~m[502]&m[503])|(m[21]&~m[500]&m[501]&~m[502]&m[503])|(~m[21]&m[500]&m[501]&~m[502]&m[503])|(m[21]&~m[500]&~m[501]&m[502]&m[503])|(~m[21]&m[500]&~m[501]&m[502]&m[503])|(~m[21]&~m[500]&m[501]&m[502]&m[503]))&~BiasedRNG[341])|((m[21]&m[500]&m[501]&m[502]&~m[503])|(m[21]&m[500]&m[501]&~m[502]&m[503])|(m[21]&m[500]&~m[501]&m[502]&m[503])|(m[21]&~m[500]&m[501]&m[502]&m[503])|(~m[21]&m[500]&m[501]&m[502]&m[503])|(m[21]&m[500]&m[501]&m[502]&m[503]))):InitCond[612];
    m[118] = run?((((m[21]&m[504]&~m[505]&~m[506]&~m[507])|(m[21]&~m[504]&m[505]&~m[506]&~m[507])|(~m[21]&m[504]&m[505]&~m[506]&~m[507])|(m[21]&~m[504]&~m[505]&m[506]&~m[507])|(~m[21]&m[504]&~m[505]&m[506]&~m[507])|(~m[21]&~m[504]&m[505]&m[506]&~m[507])|(m[21]&~m[504]&~m[505]&~m[506]&m[507])|(~m[21]&m[504]&~m[505]&~m[506]&m[507])|(~m[21]&~m[504]&m[505]&~m[506]&m[507])|(~m[21]&~m[504]&~m[505]&m[506]&m[507]))&BiasedRNG[342])|(((m[21]&m[504]&m[505]&~m[506]&~m[507])|(m[21]&m[504]&~m[505]&m[506]&~m[507])|(m[21]&~m[504]&m[505]&m[506]&~m[507])|(~m[21]&m[504]&m[505]&m[506]&~m[507])|(m[21]&m[504]&~m[505]&~m[506]&m[507])|(m[21]&~m[504]&m[505]&~m[506]&m[507])|(~m[21]&m[504]&m[505]&~m[506]&m[507])|(m[21]&~m[504]&~m[505]&m[506]&m[507])|(~m[21]&m[504]&~m[505]&m[506]&m[507])|(~m[21]&~m[504]&m[505]&m[506]&m[507]))&~BiasedRNG[342])|((m[21]&m[504]&m[505]&m[506]&~m[507])|(m[21]&m[504]&m[505]&~m[506]&m[507])|(m[21]&m[504]&~m[505]&m[506]&m[507])|(m[21]&~m[504]&m[505]&m[506]&m[507])|(~m[21]&m[504]&m[505]&m[506]&m[507])|(m[21]&m[504]&m[505]&m[506]&m[507]))):InitCond[613];
    m[119] = run?((((m[21]&m[508]&~m[509]&~m[510]&~m[511])|(m[21]&~m[508]&m[509]&~m[510]&~m[511])|(~m[21]&m[508]&m[509]&~m[510]&~m[511])|(m[21]&~m[508]&~m[509]&m[510]&~m[511])|(~m[21]&m[508]&~m[509]&m[510]&~m[511])|(~m[21]&~m[508]&m[509]&m[510]&~m[511])|(m[21]&~m[508]&~m[509]&~m[510]&m[511])|(~m[21]&m[508]&~m[509]&~m[510]&m[511])|(~m[21]&~m[508]&m[509]&~m[510]&m[511])|(~m[21]&~m[508]&~m[509]&m[510]&m[511]))&BiasedRNG[343])|(((m[21]&m[508]&m[509]&~m[510]&~m[511])|(m[21]&m[508]&~m[509]&m[510]&~m[511])|(m[21]&~m[508]&m[509]&m[510]&~m[511])|(~m[21]&m[508]&m[509]&m[510]&~m[511])|(m[21]&m[508]&~m[509]&~m[510]&m[511])|(m[21]&~m[508]&m[509]&~m[510]&m[511])|(~m[21]&m[508]&m[509]&~m[510]&m[511])|(m[21]&~m[508]&~m[509]&m[510]&m[511])|(~m[21]&m[508]&~m[509]&m[510]&m[511])|(~m[21]&~m[508]&m[509]&m[510]&m[511]))&~BiasedRNG[343])|((m[21]&m[508]&m[509]&m[510]&~m[511])|(m[21]&m[508]&m[509]&~m[510]&m[511])|(m[21]&m[508]&~m[509]&m[510]&m[511])|(m[21]&~m[508]&m[509]&m[510]&m[511])|(~m[21]&m[508]&m[509]&m[510]&m[511])|(m[21]&m[508]&m[509]&m[510]&m[511]))):InitCond[614];
    m[120] = run?((((m[22]&m[512]&~m[513]&~m[514]&~m[515])|(m[22]&~m[512]&m[513]&~m[514]&~m[515])|(~m[22]&m[512]&m[513]&~m[514]&~m[515])|(m[22]&~m[512]&~m[513]&m[514]&~m[515])|(~m[22]&m[512]&~m[513]&m[514]&~m[515])|(~m[22]&~m[512]&m[513]&m[514]&~m[515])|(m[22]&~m[512]&~m[513]&~m[514]&m[515])|(~m[22]&m[512]&~m[513]&~m[514]&m[515])|(~m[22]&~m[512]&m[513]&~m[514]&m[515])|(~m[22]&~m[512]&~m[513]&m[514]&m[515]))&BiasedRNG[344])|(((m[22]&m[512]&m[513]&~m[514]&~m[515])|(m[22]&m[512]&~m[513]&m[514]&~m[515])|(m[22]&~m[512]&m[513]&m[514]&~m[515])|(~m[22]&m[512]&m[513]&m[514]&~m[515])|(m[22]&m[512]&~m[513]&~m[514]&m[515])|(m[22]&~m[512]&m[513]&~m[514]&m[515])|(~m[22]&m[512]&m[513]&~m[514]&m[515])|(m[22]&~m[512]&~m[513]&m[514]&m[515])|(~m[22]&m[512]&~m[513]&m[514]&m[515])|(~m[22]&~m[512]&m[513]&m[514]&m[515]))&~BiasedRNG[344])|((m[22]&m[512]&m[513]&m[514]&~m[515])|(m[22]&m[512]&m[513]&~m[514]&m[515])|(m[22]&m[512]&~m[513]&m[514]&m[515])|(m[22]&~m[512]&m[513]&m[514]&m[515])|(~m[22]&m[512]&m[513]&m[514]&m[515])|(m[22]&m[512]&m[513]&m[514]&m[515]))):InitCond[615];
    m[121] = run?((((m[22]&m[516]&~m[517]&~m[518]&~m[519])|(m[22]&~m[516]&m[517]&~m[518]&~m[519])|(~m[22]&m[516]&m[517]&~m[518]&~m[519])|(m[22]&~m[516]&~m[517]&m[518]&~m[519])|(~m[22]&m[516]&~m[517]&m[518]&~m[519])|(~m[22]&~m[516]&m[517]&m[518]&~m[519])|(m[22]&~m[516]&~m[517]&~m[518]&m[519])|(~m[22]&m[516]&~m[517]&~m[518]&m[519])|(~m[22]&~m[516]&m[517]&~m[518]&m[519])|(~m[22]&~m[516]&~m[517]&m[518]&m[519]))&BiasedRNG[345])|(((m[22]&m[516]&m[517]&~m[518]&~m[519])|(m[22]&m[516]&~m[517]&m[518]&~m[519])|(m[22]&~m[516]&m[517]&m[518]&~m[519])|(~m[22]&m[516]&m[517]&m[518]&~m[519])|(m[22]&m[516]&~m[517]&~m[518]&m[519])|(m[22]&~m[516]&m[517]&~m[518]&m[519])|(~m[22]&m[516]&m[517]&~m[518]&m[519])|(m[22]&~m[516]&~m[517]&m[518]&m[519])|(~m[22]&m[516]&~m[517]&m[518]&m[519])|(~m[22]&~m[516]&m[517]&m[518]&m[519]))&~BiasedRNG[345])|((m[22]&m[516]&m[517]&m[518]&~m[519])|(m[22]&m[516]&m[517]&~m[518]&m[519])|(m[22]&m[516]&~m[517]&m[518]&m[519])|(m[22]&~m[516]&m[517]&m[518]&m[519])|(~m[22]&m[516]&m[517]&m[518]&m[519])|(m[22]&m[516]&m[517]&m[518]&m[519]))):InitCond[616];
    m[122] = run?((((m[22]&m[520]&~m[521]&~m[522]&~m[523])|(m[22]&~m[520]&m[521]&~m[522]&~m[523])|(~m[22]&m[520]&m[521]&~m[522]&~m[523])|(m[22]&~m[520]&~m[521]&m[522]&~m[523])|(~m[22]&m[520]&~m[521]&m[522]&~m[523])|(~m[22]&~m[520]&m[521]&m[522]&~m[523])|(m[22]&~m[520]&~m[521]&~m[522]&m[523])|(~m[22]&m[520]&~m[521]&~m[522]&m[523])|(~m[22]&~m[520]&m[521]&~m[522]&m[523])|(~m[22]&~m[520]&~m[521]&m[522]&m[523]))&BiasedRNG[346])|(((m[22]&m[520]&m[521]&~m[522]&~m[523])|(m[22]&m[520]&~m[521]&m[522]&~m[523])|(m[22]&~m[520]&m[521]&m[522]&~m[523])|(~m[22]&m[520]&m[521]&m[522]&~m[523])|(m[22]&m[520]&~m[521]&~m[522]&m[523])|(m[22]&~m[520]&m[521]&~m[522]&m[523])|(~m[22]&m[520]&m[521]&~m[522]&m[523])|(m[22]&~m[520]&~m[521]&m[522]&m[523])|(~m[22]&m[520]&~m[521]&m[522]&m[523])|(~m[22]&~m[520]&m[521]&m[522]&m[523]))&~BiasedRNG[346])|((m[22]&m[520]&m[521]&m[522]&~m[523])|(m[22]&m[520]&m[521]&~m[522]&m[523])|(m[22]&m[520]&~m[521]&m[522]&m[523])|(m[22]&~m[520]&m[521]&m[522]&m[523])|(~m[22]&m[520]&m[521]&m[522]&m[523])|(m[22]&m[520]&m[521]&m[522]&m[523]))):InitCond[617];
    m[123] = run?((((m[22]&m[524]&~m[525]&~m[526]&~m[527])|(m[22]&~m[524]&m[525]&~m[526]&~m[527])|(~m[22]&m[524]&m[525]&~m[526]&~m[527])|(m[22]&~m[524]&~m[525]&m[526]&~m[527])|(~m[22]&m[524]&~m[525]&m[526]&~m[527])|(~m[22]&~m[524]&m[525]&m[526]&~m[527])|(m[22]&~m[524]&~m[525]&~m[526]&m[527])|(~m[22]&m[524]&~m[525]&~m[526]&m[527])|(~m[22]&~m[524]&m[525]&~m[526]&m[527])|(~m[22]&~m[524]&~m[525]&m[526]&m[527]))&BiasedRNG[347])|(((m[22]&m[524]&m[525]&~m[526]&~m[527])|(m[22]&m[524]&~m[525]&m[526]&~m[527])|(m[22]&~m[524]&m[525]&m[526]&~m[527])|(~m[22]&m[524]&m[525]&m[526]&~m[527])|(m[22]&m[524]&~m[525]&~m[526]&m[527])|(m[22]&~m[524]&m[525]&~m[526]&m[527])|(~m[22]&m[524]&m[525]&~m[526]&m[527])|(m[22]&~m[524]&~m[525]&m[526]&m[527])|(~m[22]&m[524]&~m[525]&m[526]&m[527])|(~m[22]&~m[524]&m[525]&m[526]&m[527]))&~BiasedRNG[347])|((m[22]&m[524]&m[525]&m[526]&~m[527])|(m[22]&m[524]&m[525]&~m[526]&m[527])|(m[22]&m[524]&~m[525]&m[526]&m[527])|(m[22]&~m[524]&m[525]&m[526]&m[527])|(~m[22]&m[524]&m[525]&m[526]&m[527])|(m[22]&m[524]&m[525]&m[526]&m[527]))):InitCond[618];
    m[124] = run?((((m[23]&m[528]&~m[529]&~m[530]&~m[531])|(m[23]&~m[528]&m[529]&~m[530]&~m[531])|(~m[23]&m[528]&m[529]&~m[530]&~m[531])|(m[23]&~m[528]&~m[529]&m[530]&~m[531])|(~m[23]&m[528]&~m[529]&m[530]&~m[531])|(~m[23]&~m[528]&m[529]&m[530]&~m[531])|(m[23]&~m[528]&~m[529]&~m[530]&m[531])|(~m[23]&m[528]&~m[529]&~m[530]&m[531])|(~m[23]&~m[528]&m[529]&~m[530]&m[531])|(~m[23]&~m[528]&~m[529]&m[530]&m[531]))&BiasedRNG[348])|(((m[23]&m[528]&m[529]&~m[530]&~m[531])|(m[23]&m[528]&~m[529]&m[530]&~m[531])|(m[23]&~m[528]&m[529]&m[530]&~m[531])|(~m[23]&m[528]&m[529]&m[530]&~m[531])|(m[23]&m[528]&~m[529]&~m[530]&m[531])|(m[23]&~m[528]&m[529]&~m[530]&m[531])|(~m[23]&m[528]&m[529]&~m[530]&m[531])|(m[23]&~m[528]&~m[529]&m[530]&m[531])|(~m[23]&m[528]&~m[529]&m[530]&m[531])|(~m[23]&~m[528]&m[529]&m[530]&m[531]))&~BiasedRNG[348])|((m[23]&m[528]&m[529]&m[530]&~m[531])|(m[23]&m[528]&m[529]&~m[530]&m[531])|(m[23]&m[528]&~m[529]&m[530]&m[531])|(m[23]&~m[528]&m[529]&m[530]&m[531])|(~m[23]&m[528]&m[529]&m[530]&m[531])|(m[23]&m[528]&m[529]&m[530]&m[531]))):InitCond[619];
    m[125] = run?((((m[23]&m[532]&~m[533]&~m[534]&~m[535])|(m[23]&~m[532]&m[533]&~m[534]&~m[535])|(~m[23]&m[532]&m[533]&~m[534]&~m[535])|(m[23]&~m[532]&~m[533]&m[534]&~m[535])|(~m[23]&m[532]&~m[533]&m[534]&~m[535])|(~m[23]&~m[532]&m[533]&m[534]&~m[535])|(m[23]&~m[532]&~m[533]&~m[534]&m[535])|(~m[23]&m[532]&~m[533]&~m[534]&m[535])|(~m[23]&~m[532]&m[533]&~m[534]&m[535])|(~m[23]&~m[532]&~m[533]&m[534]&m[535]))&BiasedRNG[349])|(((m[23]&m[532]&m[533]&~m[534]&~m[535])|(m[23]&m[532]&~m[533]&m[534]&~m[535])|(m[23]&~m[532]&m[533]&m[534]&~m[535])|(~m[23]&m[532]&m[533]&m[534]&~m[535])|(m[23]&m[532]&~m[533]&~m[534]&m[535])|(m[23]&~m[532]&m[533]&~m[534]&m[535])|(~m[23]&m[532]&m[533]&~m[534]&m[535])|(m[23]&~m[532]&~m[533]&m[534]&m[535])|(~m[23]&m[532]&~m[533]&m[534]&m[535])|(~m[23]&~m[532]&m[533]&m[534]&m[535]))&~BiasedRNG[349])|((m[23]&m[532]&m[533]&m[534]&~m[535])|(m[23]&m[532]&m[533]&~m[534]&m[535])|(m[23]&m[532]&~m[533]&m[534]&m[535])|(m[23]&~m[532]&m[533]&m[534]&m[535])|(~m[23]&m[532]&m[533]&m[534]&m[535])|(m[23]&m[532]&m[533]&m[534]&m[535]))):InitCond[620];
    m[126] = run?((((m[23]&m[536]&~m[537]&~m[538]&~m[539])|(m[23]&~m[536]&m[537]&~m[538]&~m[539])|(~m[23]&m[536]&m[537]&~m[538]&~m[539])|(m[23]&~m[536]&~m[537]&m[538]&~m[539])|(~m[23]&m[536]&~m[537]&m[538]&~m[539])|(~m[23]&~m[536]&m[537]&m[538]&~m[539])|(m[23]&~m[536]&~m[537]&~m[538]&m[539])|(~m[23]&m[536]&~m[537]&~m[538]&m[539])|(~m[23]&~m[536]&m[537]&~m[538]&m[539])|(~m[23]&~m[536]&~m[537]&m[538]&m[539]))&BiasedRNG[350])|(((m[23]&m[536]&m[537]&~m[538]&~m[539])|(m[23]&m[536]&~m[537]&m[538]&~m[539])|(m[23]&~m[536]&m[537]&m[538]&~m[539])|(~m[23]&m[536]&m[537]&m[538]&~m[539])|(m[23]&m[536]&~m[537]&~m[538]&m[539])|(m[23]&~m[536]&m[537]&~m[538]&m[539])|(~m[23]&m[536]&m[537]&~m[538]&m[539])|(m[23]&~m[536]&~m[537]&m[538]&m[539])|(~m[23]&m[536]&~m[537]&m[538]&m[539])|(~m[23]&~m[536]&m[537]&m[538]&m[539]))&~BiasedRNG[350])|((m[23]&m[536]&m[537]&m[538]&~m[539])|(m[23]&m[536]&m[537]&~m[538]&m[539])|(m[23]&m[536]&~m[537]&m[538]&m[539])|(m[23]&~m[536]&m[537]&m[538]&m[539])|(~m[23]&m[536]&m[537]&m[538]&m[539])|(m[23]&m[536]&m[537]&m[538]&m[539]))):InitCond[621];
    m[127] = run?((((m[23]&m[540]&~m[541]&~m[542]&~m[543])|(m[23]&~m[540]&m[541]&~m[542]&~m[543])|(~m[23]&m[540]&m[541]&~m[542]&~m[543])|(m[23]&~m[540]&~m[541]&m[542]&~m[543])|(~m[23]&m[540]&~m[541]&m[542]&~m[543])|(~m[23]&~m[540]&m[541]&m[542]&~m[543])|(m[23]&~m[540]&~m[541]&~m[542]&m[543])|(~m[23]&m[540]&~m[541]&~m[542]&m[543])|(~m[23]&~m[540]&m[541]&~m[542]&m[543])|(~m[23]&~m[540]&~m[541]&m[542]&m[543]))&BiasedRNG[351])|(((m[23]&m[540]&m[541]&~m[542]&~m[543])|(m[23]&m[540]&~m[541]&m[542]&~m[543])|(m[23]&~m[540]&m[541]&m[542]&~m[543])|(~m[23]&m[540]&m[541]&m[542]&~m[543])|(m[23]&m[540]&~m[541]&~m[542]&m[543])|(m[23]&~m[540]&m[541]&~m[542]&m[543])|(~m[23]&m[540]&m[541]&~m[542]&m[543])|(m[23]&~m[540]&~m[541]&m[542]&m[543])|(~m[23]&m[540]&~m[541]&m[542]&m[543])|(~m[23]&~m[540]&m[541]&m[542]&m[543]))&~BiasedRNG[351])|((m[23]&m[540]&m[541]&m[542]&~m[543])|(m[23]&m[540]&m[541]&~m[542]&m[543])|(m[23]&m[540]&~m[541]&m[542]&m[543])|(m[23]&~m[540]&m[541]&m[542]&m[543])|(~m[23]&m[540]&m[541]&m[542]&m[543])|(m[23]&m[540]&m[541]&m[542]&m[543]))):InitCond[622];
    m[128] = run?((((m[24]&m[544]&~m[545]&~m[546]&~m[547])|(m[24]&~m[544]&m[545]&~m[546]&~m[547])|(~m[24]&m[544]&m[545]&~m[546]&~m[547])|(m[24]&~m[544]&~m[545]&m[546]&~m[547])|(~m[24]&m[544]&~m[545]&m[546]&~m[547])|(~m[24]&~m[544]&m[545]&m[546]&~m[547])|(m[24]&~m[544]&~m[545]&~m[546]&m[547])|(~m[24]&m[544]&~m[545]&~m[546]&m[547])|(~m[24]&~m[544]&m[545]&~m[546]&m[547])|(~m[24]&~m[544]&~m[545]&m[546]&m[547]))&BiasedRNG[352])|(((m[24]&m[544]&m[545]&~m[546]&~m[547])|(m[24]&m[544]&~m[545]&m[546]&~m[547])|(m[24]&~m[544]&m[545]&m[546]&~m[547])|(~m[24]&m[544]&m[545]&m[546]&~m[547])|(m[24]&m[544]&~m[545]&~m[546]&m[547])|(m[24]&~m[544]&m[545]&~m[546]&m[547])|(~m[24]&m[544]&m[545]&~m[546]&m[547])|(m[24]&~m[544]&~m[545]&m[546]&m[547])|(~m[24]&m[544]&~m[545]&m[546]&m[547])|(~m[24]&~m[544]&m[545]&m[546]&m[547]))&~BiasedRNG[352])|((m[24]&m[544]&m[545]&m[546]&~m[547])|(m[24]&m[544]&m[545]&~m[546]&m[547])|(m[24]&m[544]&~m[545]&m[546]&m[547])|(m[24]&~m[544]&m[545]&m[546]&m[547])|(~m[24]&m[544]&m[545]&m[546]&m[547])|(m[24]&m[544]&m[545]&m[546]&m[547]))):InitCond[623];
    m[129] = run?((((m[24]&m[548]&~m[549]&~m[550]&~m[551])|(m[24]&~m[548]&m[549]&~m[550]&~m[551])|(~m[24]&m[548]&m[549]&~m[550]&~m[551])|(m[24]&~m[548]&~m[549]&m[550]&~m[551])|(~m[24]&m[548]&~m[549]&m[550]&~m[551])|(~m[24]&~m[548]&m[549]&m[550]&~m[551])|(m[24]&~m[548]&~m[549]&~m[550]&m[551])|(~m[24]&m[548]&~m[549]&~m[550]&m[551])|(~m[24]&~m[548]&m[549]&~m[550]&m[551])|(~m[24]&~m[548]&~m[549]&m[550]&m[551]))&BiasedRNG[353])|(((m[24]&m[548]&m[549]&~m[550]&~m[551])|(m[24]&m[548]&~m[549]&m[550]&~m[551])|(m[24]&~m[548]&m[549]&m[550]&~m[551])|(~m[24]&m[548]&m[549]&m[550]&~m[551])|(m[24]&m[548]&~m[549]&~m[550]&m[551])|(m[24]&~m[548]&m[549]&~m[550]&m[551])|(~m[24]&m[548]&m[549]&~m[550]&m[551])|(m[24]&~m[548]&~m[549]&m[550]&m[551])|(~m[24]&m[548]&~m[549]&m[550]&m[551])|(~m[24]&~m[548]&m[549]&m[550]&m[551]))&~BiasedRNG[353])|((m[24]&m[548]&m[549]&m[550]&~m[551])|(m[24]&m[548]&m[549]&~m[550]&m[551])|(m[24]&m[548]&~m[549]&m[550]&m[551])|(m[24]&~m[548]&m[549]&m[550]&m[551])|(~m[24]&m[548]&m[549]&m[550]&m[551])|(m[24]&m[548]&m[549]&m[550]&m[551]))):InitCond[624];
    m[130] = run?((((m[24]&m[552]&~m[553]&~m[554]&~m[555])|(m[24]&~m[552]&m[553]&~m[554]&~m[555])|(~m[24]&m[552]&m[553]&~m[554]&~m[555])|(m[24]&~m[552]&~m[553]&m[554]&~m[555])|(~m[24]&m[552]&~m[553]&m[554]&~m[555])|(~m[24]&~m[552]&m[553]&m[554]&~m[555])|(m[24]&~m[552]&~m[553]&~m[554]&m[555])|(~m[24]&m[552]&~m[553]&~m[554]&m[555])|(~m[24]&~m[552]&m[553]&~m[554]&m[555])|(~m[24]&~m[552]&~m[553]&m[554]&m[555]))&BiasedRNG[354])|(((m[24]&m[552]&m[553]&~m[554]&~m[555])|(m[24]&m[552]&~m[553]&m[554]&~m[555])|(m[24]&~m[552]&m[553]&m[554]&~m[555])|(~m[24]&m[552]&m[553]&m[554]&~m[555])|(m[24]&m[552]&~m[553]&~m[554]&m[555])|(m[24]&~m[552]&m[553]&~m[554]&m[555])|(~m[24]&m[552]&m[553]&~m[554]&m[555])|(m[24]&~m[552]&~m[553]&m[554]&m[555])|(~m[24]&m[552]&~m[553]&m[554]&m[555])|(~m[24]&~m[552]&m[553]&m[554]&m[555]))&~BiasedRNG[354])|((m[24]&m[552]&m[553]&m[554]&~m[555])|(m[24]&m[552]&m[553]&~m[554]&m[555])|(m[24]&m[552]&~m[553]&m[554]&m[555])|(m[24]&~m[552]&m[553]&m[554]&m[555])|(~m[24]&m[552]&m[553]&m[554]&m[555])|(m[24]&m[552]&m[553]&m[554]&m[555]))):InitCond[625];
    m[131] = run?((((m[24]&m[556]&~m[557]&~m[558]&~m[559])|(m[24]&~m[556]&m[557]&~m[558]&~m[559])|(~m[24]&m[556]&m[557]&~m[558]&~m[559])|(m[24]&~m[556]&~m[557]&m[558]&~m[559])|(~m[24]&m[556]&~m[557]&m[558]&~m[559])|(~m[24]&~m[556]&m[557]&m[558]&~m[559])|(m[24]&~m[556]&~m[557]&~m[558]&m[559])|(~m[24]&m[556]&~m[557]&~m[558]&m[559])|(~m[24]&~m[556]&m[557]&~m[558]&m[559])|(~m[24]&~m[556]&~m[557]&m[558]&m[559]))&BiasedRNG[355])|(((m[24]&m[556]&m[557]&~m[558]&~m[559])|(m[24]&m[556]&~m[557]&m[558]&~m[559])|(m[24]&~m[556]&m[557]&m[558]&~m[559])|(~m[24]&m[556]&m[557]&m[558]&~m[559])|(m[24]&m[556]&~m[557]&~m[558]&m[559])|(m[24]&~m[556]&m[557]&~m[558]&m[559])|(~m[24]&m[556]&m[557]&~m[558]&m[559])|(m[24]&~m[556]&~m[557]&m[558]&m[559])|(~m[24]&m[556]&~m[557]&m[558]&m[559])|(~m[24]&~m[556]&m[557]&m[558]&m[559]))&~BiasedRNG[355])|((m[24]&m[556]&m[557]&m[558]&~m[559])|(m[24]&m[556]&m[557]&~m[558]&m[559])|(m[24]&m[556]&~m[557]&m[558]&m[559])|(m[24]&~m[556]&m[557]&m[558]&m[559])|(~m[24]&m[556]&m[557]&m[558]&m[559])|(m[24]&m[556]&m[557]&m[558]&m[559]))):InitCond[626];
    m[132] = run?((((m[25]&m[560]&~m[561]&~m[562]&~m[563])|(m[25]&~m[560]&m[561]&~m[562]&~m[563])|(~m[25]&m[560]&m[561]&~m[562]&~m[563])|(m[25]&~m[560]&~m[561]&m[562]&~m[563])|(~m[25]&m[560]&~m[561]&m[562]&~m[563])|(~m[25]&~m[560]&m[561]&m[562]&~m[563])|(m[25]&~m[560]&~m[561]&~m[562]&m[563])|(~m[25]&m[560]&~m[561]&~m[562]&m[563])|(~m[25]&~m[560]&m[561]&~m[562]&m[563])|(~m[25]&~m[560]&~m[561]&m[562]&m[563]))&BiasedRNG[356])|(((m[25]&m[560]&m[561]&~m[562]&~m[563])|(m[25]&m[560]&~m[561]&m[562]&~m[563])|(m[25]&~m[560]&m[561]&m[562]&~m[563])|(~m[25]&m[560]&m[561]&m[562]&~m[563])|(m[25]&m[560]&~m[561]&~m[562]&m[563])|(m[25]&~m[560]&m[561]&~m[562]&m[563])|(~m[25]&m[560]&m[561]&~m[562]&m[563])|(m[25]&~m[560]&~m[561]&m[562]&m[563])|(~m[25]&m[560]&~m[561]&m[562]&m[563])|(~m[25]&~m[560]&m[561]&m[562]&m[563]))&~BiasedRNG[356])|((m[25]&m[560]&m[561]&m[562]&~m[563])|(m[25]&m[560]&m[561]&~m[562]&m[563])|(m[25]&m[560]&~m[561]&m[562]&m[563])|(m[25]&~m[560]&m[561]&m[562]&m[563])|(~m[25]&m[560]&m[561]&m[562]&m[563])|(m[25]&m[560]&m[561]&m[562]&m[563]))):InitCond[627];
    m[133] = run?((((m[25]&m[564]&~m[565]&~m[566]&~m[567])|(m[25]&~m[564]&m[565]&~m[566]&~m[567])|(~m[25]&m[564]&m[565]&~m[566]&~m[567])|(m[25]&~m[564]&~m[565]&m[566]&~m[567])|(~m[25]&m[564]&~m[565]&m[566]&~m[567])|(~m[25]&~m[564]&m[565]&m[566]&~m[567])|(m[25]&~m[564]&~m[565]&~m[566]&m[567])|(~m[25]&m[564]&~m[565]&~m[566]&m[567])|(~m[25]&~m[564]&m[565]&~m[566]&m[567])|(~m[25]&~m[564]&~m[565]&m[566]&m[567]))&BiasedRNG[357])|(((m[25]&m[564]&m[565]&~m[566]&~m[567])|(m[25]&m[564]&~m[565]&m[566]&~m[567])|(m[25]&~m[564]&m[565]&m[566]&~m[567])|(~m[25]&m[564]&m[565]&m[566]&~m[567])|(m[25]&m[564]&~m[565]&~m[566]&m[567])|(m[25]&~m[564]&m[565]&~m[566]&m[567])|(~m[25]&m[564]&m[565]&~m[566]&m[567])|(m[25]&~m[564]&~m[565]&m[566]&m[567])|(~m[25]&m[564]&~m[565]&m[566]&m[567])|(~m[25]&~m[564]&m[565]&m[566]&m[567]))&~BiasedRNG[357])|((m[25]&m[564]&m[565]&m[566]&~m[567])|(m[25]&m[564]&m[565]&~m[566]&m[567])|(m[25]&m[564]&~m[565]&m[566]&m[567])|(m[25]&~m[564]&m[565]&m[566]&m[567])|(~m[25]&m[564]&m[565]&m[566]&m[567])|(m[25]&m[564]&m[565]&m[566]&m[567]))):InitCond[628];
    m[134] = run?((((m[25]&m[568]&~m[569]&~m[570]&~m[571])|(m[25]&~m[568]&m[569]&~m[570]&~m[571])|(~m[25]&m[568]&m[569]&~m[570]&~m[571])|(m[25]&~m[568]&~m[569]&m[570]&~m[571])|(~m[25]&m[568]&~m[569]&m[570]&~m[571])|(~m[25]&~m[568]&m[569]&m[570]&~m[571])|(m[25]&~m[568]&~m[569]&~m[570]&m[571])|(~m[25]&m[568]&~m[569]&~m[570]&m[571])|(~m[25]&~m[568]&m[569]&~m[570]&m[571])|(~m[25]&~m[568]&~m[569]&m[570]&m[571]))&BiasedRNG[358])|(((m[25]&m[568]&m[569]&~m[570]&~m[571])|(m[25]&m[568]&~m[569]&m[570]&~m[571])|(m[25]&~m[568]&m[569]&m[570]&~m[571])|(~m[25]&m[568]&m[569]&m[570]&~m[571])|(m[25]&m[568]&~m[569]&~m[570]&m[571])|(m[25]&~m[568]&m[569]&~m[570]&m[571])|(~m[25]&m[568]&m[569]&~m[570]&m[571])|(m[25]&~m[568]&~m[569]&m[570]&m[571])|(~m[25]&m[568]&~m[569]&m[570]&m[571])|(~m[25]&~m[568]&m[569]&m[570]&m[571]))&~BiasedRNG[358])|((m[25]&m[568]&m[569]&m[570]&~m[571])|(m[25]&m[568]&m[569]&~m[570]&m[571])|(m[25]&m[568]&~m[569]&m[570]&m[571])|(m[25]&~m[568]&m[569]&m[570]&m[571])|(~m[25]&m[568]&m[569]&m[570]&m[571])|(m[25]&m[568]&m[569]&m[570]&m[571]))):InitCond[629];
    m[135] = run?((((m[25]&m[572]&~m[573]&~m[574]&~m[575])|(m[25]&~m[572]&m[573]&~m[574]&~m[575])|(~m[25]&m[572]&m[573]&~m[574]&~m[575])|(m[25]&~m[572]&~m[573]&m[574]&~m[575])|(~m[25]&m[572]&~m[573]&m[574]&~m[575])|(~m[25]&~m[572]&m[573]&m[574]&~m[575])|(m[25]&~m[572]&~m[573]&~m[574]&m[575])|(~m[25]&m[572]&~m[573]&~m[574]&m[575])|(~m[25]&~m[572]&m[573]&~m[574]&m[575])|(~m[25]&~m[572]&~m[573]&m[574]&m[575]))&BiasedRNG[359])|(((m[25]&m[572]&m[573]&~m[574]&~m[575])|(m[25]&m[572]&~m[573]&m[574]&~m[575])|(m[25]&~m[572]&m[573]&m[574]&~m[575])|(~m[25]&m[572]&m[573]&m[574]&~m[575])|(m[25]&m[572]&~m[573]&~m[574]&m[575])|(m[25]&~m[572]&m[573]&~m[574]&m[575])|(~m[25]&m[572]&m[573]&~m[574]&m[575])|(m[25]&~m[572]&~m[573]&m[574]&m[575])|(~m[25]&m[572]&~m[573]&m[574]&m[575])|(~m[25]&~m[572]&m[573]&m[574]&m[575]))&~BiasedRNG[359])|((m[25]&m[572]&m[573]&m[574]&~m[575])|(m[25]&m[572]&m[573]&~m[574]&m[575])|(m[25]&m[572]&~m[573]&m[574]&m[575])|(m[25]&~m[572]&m[573]&m[574]&m[575])|(~m[25]&m[572]&m[573]&m[574]&m[575])|(m[25]&m[572]&m[573]&m[574]&m[575]))):InitCond[630];
    m[136] = run?((((m[26]&m[576]&~m[577]&~m[578]&~m[579])|(m[26]&~m[576]&m[577]&~m[578]&~m[579])|(~m[26]&m[576]&m[577]&~m[578]&~m[579])|(m[26]&~m[576]&~m[577]&m[578]&~m[579])|(~m[26]&m[576]&~m[577]&m[578]&~m[579])|(~m[26]&~m[576]&m[577]&m[578]&~m[579])|(m[26]&~m[576]&~m[577]&~m[578]&m[579])|(~m[26]&m[576]&~m[577]&~m[578]&m[579])|(~m[26]&~m[576]&m[577]&~m[578]&m[579])|(~m[26]&~m[576]&~m[577]&m[578]&m[579]))&BiasedRNG[360])|(((m[26]&m[576]&m[577]&~m[578]&~m[579])|(m[26]&m[576]&~m[577]&m[578]&~m[579])|(m[26]&~m[576]&m[577]&m[578]&~m[579])|(~m[26]&m[576]&m[577]&m[578]&~m[579])|(m[26]&m[576]&~m[577]&~m[578]&m[579])|(m[26]&~m[576]&m[577]&~m[578]&m[579])|(~m[26]&m[576]&m[577]&~m[578]&m[579])|(m[26]&~m[576]&~m[577]&m[578]&m[579])|(~m[26]&m[576]&~m[577]&m[578]&m[579])|(~m[26]&~m[576]&m[577]&m[578]&m[579]))&~BiasedRNG[360])|((m[26]&m[576]&m[577]&m[578]&~m[579])|(m[26]&m[576]&m[577]&~m[578]&m[579])|(m[26]&m[576]&~m[577]&m[578]&m[579])|(m[26]&~m[576]&m[577]&m[578]&m[579])|(~m[26]&m[576]&m[577]&m[578]&m[579])|(m[26]&m[576]&m[577]&m[578]&m[579]))):InitCond[631];
    m[137] = run?((((m[26]&m[580]&~m[581]&~m[582]&~m[583])|(m[26]&~m[580]&m[581]&~m[582]&~m[583])|(~m[26]&m[580]&m[581]&~m[582]&~m[583])|(m[26]&~m[580]&~m[581]&m[582]&~m[583])|(~m[26]&m[580]&~m[581]&m[582]&~m[583])|(~m[26]&~m[580]&m[581]&m[582]&~m[583])|(m[26]&~m[580]&~m[581]&~m[582]&m[583])|(~m[26]&m[580]&~m[581]&~m[582]&m[583])|(~m[26]&~m[580]&m[581]&~m[582]&m[583])|(~m[26]&~m[580]&~m[581]&m[582]&m[583]))&BiasedRNG[361])|(((m[26]&m[580]&m[581]&~m[582]&~m[583])|(m[26]&m[580]&~m[581]&m[582]&~m[583])|(m[26]&~m[580]&m[581]&m[582]&~m[583])|(~m[26]&m[580]&m[581]&m[582]&~m[583])|(m[26]&m[580]&~m[581]&~m[582]&m[583])|(m[26]&~m[580]&m[581]&~m[582]&m[583])|(~m[26]&m[580]&m[581]&~m[582]&m[583])|(m[26]&~m[580]&~m[581]&m[582]&m[583])|(~m[26]&m[580]&~m[581]&m[582]&m[583])|(~m[26]&~m[580]&m[581]&m[582]&m[583]))&~BiasedRNG[361])|((m[26]&m[580]&m[581]&m[582]&~m[583])|(m[26]&m[580]&m[581]&~m[582]&m[583])|(m[26]&m[580]&~m[581]&m[582]&m[583])|(m[26]&~m[580]&m[581]&m[582]&m[583])|(~m[26]&m[580]&m[581]&m[582]&m[583])|(m[26]&m[580]&m[581]&m[582]&m[583]))):InitCond[632];
    m[138] = run?((((m[26]&m[584]&~m[585]&~m[586]&~m[587])|(m[26]&~m[584]&m[585]&~m[586]&~m[587])|(~m[26]&m[584]&m[585]&~m[586]&~m[587])|(m[26]&~m[584]&~m[585]&m[586]&~m[587])|(~m[26]&m[584]&~m[585]&m[586]&~m[587])|(~m[26]&~m[584]&m[585]&m[586]&~m[587])|(m[26]&~m[584]&~m[585]&~m[586]&m[587])|(~m[26]&m[584]&~m[585]&~m[586]&m[587])|(~m[26]&~m[584]&m[585]&~m[586]&m[587])|(~m[26]&~m[584]&~m[585]&m[586]&m[587]))&BiasedRNG[362])|(((m[26]&m[584]&m[585]&~m[586]&~m[587])|(m[26]&m[584]&~m[585]&m[586]&~m[587])|(m[26]&~m[584]&m[585]&m[586]&~m[587])|(~m[26]&m[584]&m[585]&m[586]&~m[587])|(m[26]&m[584]&~m[585]&~m[586]&m[587])|(m[26]&~m[584]&m[585]&~m[586]&m[587])|(~m[26]&m[584]&m[585]&~m[586]&m[587])|(m[26]&~m[584]&~m[585]&m[586]&m[587])|(~m[26]&m[584]&~m[585]&m[586]&m[587])|(~m[26]&~m[584]&m[585]&m[586]&m[587]))&~BiasedRNG[362])|((m[26]&m[584]&m[585]&m[586]&~m[587])|(m[26]&m[584]&m[585]&~m[586]&m[587])|(m[26]&m[584]&~m[585]&m[586]&m[587])|(m[26]&~m[584]&m[585]&m[586]&m[587])|(~m[26]&m[584]&m[585]&m[586]&m[587])|(m[26]&m[584]&m[585]&m[586]&m[587]))):InitCond[633];
    m[139] = run?((((m[26]&m[588]&~m[589]&~m[590]&~m[591])|(m[26]&~m[588]&m[589]&~m[590]&~m[591])|(~m[26]&m[588]&m[589]&~m[590]&~m[591])|(m[26]&~m[588]&~m[589]&m[590]&~m[591])|(~m[26]&m[588]&~m[589]&m[590]&~m[591])|(~m[26]&~m[588]&m[589]&m[590]&~m[591])|(m[26]&~m[588]&~m[589]&~m[590]&m[591])|(~m[26]&m[588]&~m[589]&~m[590]&m[591])|(~m[26]&~m[588]&m[589]&~m[590]&m[591])|(~m[26]&~m[588]&~m[589]&m[590]&m[591]))&BiasedRNG[363])|(((m[26]&m[588]&m[589]&~m[590]&~m[591])|(m[26]&m[588]&~m[589]&m[590]&~m[591])|(m[26]&~m[588]&m[589]&m[590]&~m[591])|(~m[26]&m[588]&m[589]&m[590]&~m[591])|(m[26]&m[588]&~m[589]&~m[590]&m[591])|(m[26]&~m[588]&m[589]&~m[590]&m[591])|(~m[26]&m[588]&m[589]&~m[590]&m[591])|(m[26]&~m[588]&~m[589]&m[590]&m[591])|(~m[26]&m[588]&~m[589]&m[590]&m[591])|(~m[26]&~m[588]&m[589]&m[590]&m[591]))&~BiasedRNG[363])|((m[26]&m[588]&m[589]&m[590]&~m[591])|(m[26]&m[588]&m[589]&~m[590]&m[591])|(m[26]&m[588]&~m[589]&m[590]&m[591])|(m[26]&~m[588]&m[589]&m[590]&m[591])|(~m[26]&m[588]&m[589]&m[590]&m[591])|(m[26]&m[588]&m[589]&m[590]&m[591]))):InitCond[634];
    m[140] = run?((((m[27]&m[592]&~m[593]&~m[594]&~m[595])|(m[27]&~m[592]&m[593]&~m[594]&~m[595])|(~m[27]&m[592]&m[593]&~m[594]&~m[595])|(m[27]&~m[592]&~m[593]&m[594]&~m[595])|(~m[27]&m[592]&~m[593]&m[594]&~m[595])|(~m[27]&~m[592]&m[593]&m[594]&~m[595])|(m[27]&~m[592]&~m[593]&~m[594]&m[595])|(~m[27]&m[592]&~m[593]&~m[594]&m[595])|(~m[27]&~m[592]&m[593]&~m[594]&m[595])|(~m[27]&~m[592]&~m[593]&m[594]&m[595]))&BiasedRNG[364])|(((m[27]&m[592]&m[593]&~m[594]&~m[595])|(m[27]&m[592]&~m[593]&m[594]&~m[595])|(m[27]&~m[592]&m[593]&m[594]&~m[595])|(~m[27]&m[592]&m[593]&m[594]&~m[595])|(m[27]&m[592]&~m[593]&~m[594]&m[595])|(m[27]&~m[592]&m[593]&~m[594]&m[595])|(~m[27]&m[592]&m[593]&~m[594]&m[595])|(m[27]&~m[592]&~m[593]&m[594]&m[595])|(~m[27]&m[592]&~m[593]&m[594]&m[595])|(~m[27]&~m[592]&m[593]&m[594]&m[595]))&~BiasedRNG[364])|((m[27]&m[592]&m[593]&m[594]&~m[595])|(m[27]&m[592]&m[593]&~m[594]&m[595])|(m[27]&m[592]&~m[593]&m[594]&m[595])|(m[27]&~m[592]&m[593]&m[594]&m[595])|(~m[27]&m[592]&m[593]&m[594]&m[595])|(m[27]&m[592]&m[593]&m[594]&m[595]))):InitCond[635];
    m[141] = run?((((m[27]&m[596]&~m[597]&~m[598]&~m[599])|(m[27]&~m[596]&m[597]&~m[598]&~m[599])|(~m[27]&m[596]&m[597]&~m[598]&~m[599])|(m[27]&~m[596]&~m[597]&m[598]&~m[599])|(~m[27]&m[596]&~m[597]&m[598]&~m[599])|(~m[27]&~m[596]&m[597]&m[598]&~m[599])|(m[27]&~m[596]&~m[597]&~m[598]&m[599])|(~m[27]&m[596]&~m[597]&~m[598]&m[599])|(~m[27]&~m[596]&m[597]&~m[598]&m[599])|(~m[27]&~m[596]&~m[597]&m[598]&m[599]))&BiasedRNG[365])|(((m[27]&m[596]&m[597]&~m[598]&~m[599])|(m[27]&m[596]&~m[597]&m[598]&~m[599])|(m[27]&~m[596]&m[597]&m[598]&~m[599])|(~m[27]&m[596]&m[597]&m[598]&~m[599])|(m[27]&m[596]&~m[597]&~m[598]&m[599])|(m[27]&~m[596]&m[597]&~m[598]&m[599])|(~m[27]&m[596]&m[597]&~m[598]&m[599])|(m[27]&~m[596]&~m[597]&m[598]&m[599])|(~m[27]&m[596]&~m[597]&m[598]&m[599])|(~m[27]&~m[596]&m[597]&m[598]&m[599]))&~BiasedRNG[365])|((m[27]&m[596]&m[597]&m[598]&~m[599])|(m[27]&m[596]&m[597]&~m[598]&m[599])|(m[27]&m[596]&~m[597]&m[598]&m[599])|(m[27]&~m[596]&m[597]&m[598]&m[599])|(~m[27]&m[596]&m[597]&m[598]&m[599])|(m[27]&m[596]&m[597]&m[598]&m[599]))):InitCond[636];
    m[142] = run?((((m[27]&m[600]&~m[601]&~m[602]&~m[603])|(m[27]&~m[600]&m[601]&~m[602]&~m[603])|(~m[27]&m[600]&m[601]&~m[602]&~m[603])|(m[27]&~m[600]&~m[601]&m[602]&~m[603])|(~m[27]&m[600]&~m[601]&m[602]&~m[603])|(~m[27]&~m[600]&m[601]&m[602]&~m[603])|(m[27]&~m[600]&~m[601]&~m[602]&m[603])|(~m[27]&m[600]&~m[601]&~m[602]&m[603])|(~m[27]&~m[600]&m[601]&~m[602]&m[603])|(~m[27]&~m[600]&~m[601]&m[602]&m[603]))&BiasedRNG[366])|(((m[27]&m[600]&m[601]&~m[602]&~m[603])|(m[27]&m[600]&~m[601]&m[602]&~m[603])|(m[27]&~m[600]&m[601]&m[602]&~m[603])|(~m[27]&m[600]&m[601]&m[602]&~m[603])|(m[27]&m[600]&~m[601]&~m[602]&m[603])|(m[27]&~m[600]&m[601]&~m[602]&m[603])|(~m[27]&m[600]&m[601]&~m[602]&m[603])|(m[27]&~m[600]&~m[601]&m[602]&m[603])|(~m[27]&m[600]&~m[601]&m[602]&m[603])|(~m[27]&~m[600]&m[601]&m[602]&m[603]))&~BiasedRNG[366])|((m[27]&m[600]&m[601]&m[602]&~m[603])|(m[27]&m[600]&m[601]&~m[602]&m[603])|(m[27]&m[600]&~m[601]&m[602]&m[603])|(m[27]&~m[600]&m[601]&m[602]&m[603])|(~m[27]&m[600]&m[601]&m[602]&m[603])|(m[27]&m[600]&m[601]&m[602]&m[603]))):InitCond[637];
    m[143] = run?((((m[27]&m[604]&~m[605]&~m[606]&~m[607])|(m[27]&~m[604]&m[605]&~m[606]&~m[607])|(~m[27]&m[604]&m[605]&~m[606]&~m[607])|(m[27]&~m[604]&~m[605]&m[606]&~m[607])|(~m[27]&m[604]&~m[605]&m[606]&~m[607])|(~m[27]&~m[604]&m[605]&m[606]&~m[607])|(m[27]&~m[604]&~m[605]&~m[606]&m[607])|(~m[27]&m[604]&~m[605]&~m[606]&m[607])|(~m[27]&~m[604]&m[605]&~m[606]&m[607])|(~m[27]&~m[604]&~m[605]&m[606]&m[607]))&BiasedRNG[367])|(((m[27]&m[604]&m[605]&~m[606]&~m[607])|(m[27]&m[604]&~m[605]&m[606]&~m[607])|(m[27]&~m[604]&m[605]&m[606]&~m[607])|(~m[27]&m[604]&m[605]&m[606]&~m[607])|(m[27]&m[604]&~m[605]&~m[606]&m[607])|(m[27]&~m[604]&m[605]&~m[606]&m[607])|(~m[27]&m[604]&m[605]&~m[606]&m[607])|(m[27]&~m[604]&~m[605]&m[606]&m[607])|(~m[27]&m[604]&~m[605]&m[606]&m[607])|(~m[27]&~m[604]&m[605]&m[606]&m[607]))&~BiasedRNG[367])|((m[27]&m[604]&m[605]&m[606]&~m[607])|(m[27]&m[604]&m[605]&~m[606]&m[607])|(m[27]&m[604]&~m[605]&m[606]&m[607])|(m[27]&~m[604]&m[605]&m[606]&m[607])|(~m[27]&m[604]&m[605]&m[606]&m[607])|(m[27]&m[604]&m[605]&m[606]&m[607]))):InitCond[638];
    m[144] = run?((((m[28]&m[608]&~m[609]&~m[610]&~m[611])|(m[28]&~m[608]&m[609]&~m[610]&~m[611])|(~m[28]&m[608]&m[609]&~m[610]&~m[611])|(m[28]&~m[608]&~m[609]&m[610]&~m[611])|(~m[28]&m[608]&~m[609]&m[610]&~m[611])|(~m[28]&~m[608]&m[609]&m[610]&~m[611])|(m[28]&~m[608]&~m[609]&~m[610]&m[611])|(~m[28]&m[608]&~m[609]&~m[610]&m[611])|(~m[28]&~m[608]&m[609]&~m[610]&m[611])|(~m[28]&~m[608]&~m[609]&m[610]&m[611]))&BiasedRNG[368])|(((m[28]&m[608]&m[609]&~m[610]&~m[611])|(m[28]&m[608]&~m[609]&m[610]&~m[611])|(m[28]&~m[608]&m[609]&m[610]&~m[611])|(~m[28]&m[608]&m[609]&m[610]&~m[611])|(m[28]&m[608]&~m[609]&~m[610]&m[611])|(m[28]&~m[608]&m[609]&~m[610]&m[611])|(~m[28]&m[608]&m[609]&~m[610]&m[611])|(m[28]&~m[608]&~m[609]&m[610]&m[611])|(~m[28]&m[608]&~m[609]&m[610]&m[611])|(~m[28]&~m[608]&m[609]&m[610]&m[611]))&~BiasedRNG[368])|((m[28]&m[608]&m[609]&m[610]&~m[611])|(m[28]&m[608]&m[609]&~m[610]&m[611])|(m[28]&m[608]&~m[609]&m[610]&m[611])|(m[28]&~m[608]&m[609]&m[610]&m[611])|(~m[28]&m[608]&m[609]&m[610]&m[611])|(m[28]&m[608]&m[609]&m[610]&m[611]))):InitCond[639];
    m[145] = run?((((m[28]&m[612]&~m[613]&~m[614]&~m[615])|(m[28]&~m[612]&m[613]&~m[614]&~m[615])|(~m[28]&m[612]&m[613]&~m[614]&~m[615])|(m[28]&~m[612]&~m[613]&m[614]&~m[615])|(~m[28]&m[612]&~m[613]&m[614]&~m[615])|(~m[28]&~m[612]&m[613]&m[614]&~m[615])|(m[28]&~m[612]&~m[613]&~m[614]&m[615])|(~m[28]&m[612]&~m[613]&~m[614]&m[615])|(~m[28]&~m[612]&m[613]&~m[614]&m[615])|(~m[28]&~m[612]&~m[613]&m[614]&m[615]))&BiasedRNG[369])|(((m[28]&m[612]&m[613]&~m[614]&~m[615])|(m[28]&m[612]&~m[613]&m[614]&~m[615])|(m[28]&~m[612]&m[613]&m[614]&~m[615])|(~m[28]&m[612]&m[613]&m[614]&~m[615])|(m[28]&m[612]&~m[613]&~m[614]&m[615])|(m[28]&~m[612]&m[613]&~m[614]&m[615])|(~m[28]&m[612]&m[613]&~m[614]&m[615])|(m[28]&~m[612]&~m[613]&m[614]&m[615])|(~m[28]&m[612]&~m[613]&m[614]&m[615])|(~m[28]&~m[612]&m[613]&m[614]&m[615]))&~BiasedRNG[369])|((m[28]&m[612]&m[613]&m[614]&~m[615])|(m[28]&m[612]&m[613]&~m[614]&m[615])|(m[28]&m[612]&~m[613]&m[614]&m[615])|(m[28]&~m[612]&m[613]&m[614]&m[615])|(~m[28]&m[612]&m[613]&m[614]&m[615])|(m[28]&m[612]&m[613]&m[614]&m[615]))):InitCond[640];
    m[146] = run?((((m[28]&m[616]&~m[617]&~m[618]&~m[619])|(m[28]&~m[616]&m[617]&~m[618]&~m[619])|(~m[28]&m[616]&m[617]&~m[618]&~m[619])|(m[28]&~m[616]&~m[617]&m[618]&~m[619])|(~m[28]&m[616]&~m[617]&m[618]&~m[619])|(~m[28]&~m[616]&m[617]&m[618]&~m[619])|(m[28]&~m[616]&~m[617]&~m[618]&m[619])|(~m[28]&m[616]&~m[617]&~m[618]&m[619])|(~m[28]&~m[616]&m[617]&~m[618]&m[619])|(~m[28]&~m[616]&~m[617]&m[618]&m[619]))&BiasedRNG[370])|(((m[28]&m[616]&m[617]&~m[618]&~m[619])|(m[28]&m[616]&~m[617]&m[618]&~m[619])|(m[28]&~m[616]&m[617]&m[618]&~m[619])|(~m[28]&m[616]&m[617]&m[618]&~m[619])|(m[28]&m[616]&~m[617]&~m[618]&m[619])|(m[28]&~m[616]&m[617]&~m[618]&m[619])|(~m[28]&m[616]&m[617]&~m[618]&m[619])|(m[28]&~m[616]&~m[617]&m[618]&m[619])|(~m[28]&m[616]&~m[617]&m[618]&m[619])|(~m[28]&~m[616]&m[617]&m[618]&m[619]))&~BiasedRNG[370])|((m[28]&m[616]&m[617]&m[618]&~m[619])|(m[28]&m[616]&m[617]&~m[618]&m[619])|(m[28]&m[616]&~m[617]&m[618]&m[619])|(m[28]&~m[616]&m[617]&m[618]&m[619])|(~m[28]&m[616]&m[617]&m[618]&m[619])|(m[28]&m[616]&m[617]&m[618]&m[619]))):InitCond[641];
    m[147] = run?((((m[28]&m[620]&~m[621]&~m[622]&~m[623])|(m[28]&~m[620]&m[621]&~m[622]&~m[623])|(~m[28]&m[620]&m[621]&~m[622]&~m[623])|(m[28]&~m[620]&~m[621]&m[622]&~m[623])|(~m[28]&m[620]&~m[621]&m[622]&~m[623])|(~m[28]&~m[620]&m[621]&m[622]&~m[623])|(m[28]&~m[620]&~m[621]&~m[622]&m[623])|(~m[28]&m[620]&~m[621]&~m[622]&m[623])|(~m[28]&~m[620]&m[621]&~m[622]&m[623])|(~m[28]&~m[620]&~m[621]&m[622]&m[623]))&BiasedRNG[371])|(((m[28]&m[620]&m[621]&~m[622]&~m[623])|(m[28]&m[620]&~m[621]&m[622]&~m[623])|(m[28]&~m[620]&m[621]&m[622]&~m[623])|(~m[28]&m[620]&m[621]&m[622]&~m[623])|(m[28]&m[620]&~m[621]&~m[622]&m[623])|(m[28]&~m[620]&m[621]&~m[622]&m[623])|(~m[28]&m[620]&m[621]&~m[622]&m[623])|(m[28]&~m[620]&~m[621]&m[622]&m[623])|(~m[28]&m[620]&~m[621]&m[622]&m[623])|(~m[28]&~m[620]&m[621]&m[622]&m[623]))&~BiasedRNG[371])|((m[28]&m[620]&m[621]&m[622]&~m[623])|(m[28]&m[620]&m[621]&~m[622]&m[623])|(m[28]&m[620]&~m[621]&m[622]&m[623])|(m[28]&~m[620]&m[621]&m[622]&m[623])|(~m[28]&m[620]&m[621]&m[622]&m[623])|(m[28]&m[620]&m[621]&m[622]&m[623]))):InitCond[642];
    m[148] = run?((((m[29]&m[624]&~m[625]&~m[626]&~m[627])|(m[29]&~m[624]&m[625]&~m[626]&~m[627])|(~m[29]&m[624]&m[625]&~m[626]&~m[627])|(m[29]&~m[624]&~m[625]&m[626]&~m[627])|(~m[29]&m[624]&~m[625]&m[626]&~m[627])|(~m[29]&~m[624]&m[625]&m[626]&~m[627])|(m[29]&~m[624]&~m[625]&~m[626]&m[627])|(~m[29]&m[624]&~m[625]&~m[626]&m[627])|(~m[29]&~m[624]&m[625]&~m[626]&m[627])|(~m[29]&~m[624]&~m[625]&m[626]&m[627]))&BiasedRNG[372])|(((m[29]&m[624]&m[625]&~m[626]&~m[627])|(m[29]&m[624]&~m[625]&m[626]&~m[627])|(m[29]&~m[624]&m[625]&m[626]&~m[627])|(~m[29]&m[624]&m[625]&m[626]&~m[627])|(m[29]&m[624]&~m[625]&~m[626]&m[627])|(m[29]&~m[624]&m[625]&~m[626]&m[627])|(~m[29]&m[624]&m[625]&~m[626]&m[627])|(m[29]&~m[624]&~m[625]&m[626]&m[627])|(~m[29]&m[624]&~m[625]&m[626]&m[627])|(~m[29]&~m[624]&m[625]&m[626]&m[627]))&~BiasedRNG[372])|((m[29]&m[624]&m[625]&m[626]&~m[627])|(m[29]&m[624]&m[625]&~m[626]&m[627])|(m[29]&m[624]&~m[625]&m[626]&m[627])|(m[29]&~m[624]&m[625]&m[626]&m[627])|(~m[29]&m[624]&m[625]&m[626]&m[627])|(m[29]&m[624]&m[625]&m[626]&m[627]))):InitCond[643];
    m[149] = run?((((m[29]&m[628]&~m[629]&~m[630]&~m[631])|(m[29]&~m[628]&m[629]&~m[630]&~m[631])|(~m[29]&m[628]&m[629]&~m[630]&~m[631])|(m[29]&~m[628]&~m[629]&m[630]&~m[631])|(~m[29]&m[628]&~m[629]&m[630]&~m[631])|(~m[29]&~m[628]&m[629]&m[630]&~m[631])|(m[29]&~m[628]&~m[629]&~m[630]&m[631])|(~m[29]&m[628]&~m[629]&~m[630]&m[631])|(~m[29]&~m[628]&m[629]&~m[630]&m[631])|(~m[29]&~m[628]&~m[629]&m[630]&m[631]))&BiasedRNG[373])|(((m[29]&m[628]&m[629]&~m[630]&~m[631])|(m[29]&m[628]&~m[629]&m[630]&~m[631])|(m[29]&~m[628]&m[629]&m[630]&~m[631])|(~m[29]&m[628]&m[629]&m[630]&~m[631])|(m[29]&m[628]&~m[629]&~m[630]&m[631])|(m[29]&~m[628]&m[629]&~m[630]&m[631])|(~m[29]&m[628]&m[629]&~m[630]&m[631])|(m[29]&~m[628]&~m[629]&m[630]&m[631])|(~m[29]&m[628]&~m[629]&m[630]&m[631])|(~m[29]&~m[628]&m[629]&m[630]&m[631]))&~BiasedRNG[373])|((m[29]&m[628]&m[629]&m[630]&~m[631])|(m[29]&m[628]&m[629]&~m[630]&m[631])|(m[29]&m[628]&~m[629]&m[630]&m[631])|(m[29]&~m[628]&m[629]&m[630]&m[631])|(~m[29]&m[628]&m[629]&m[630]&m[631])|(m[29]&m[628]&m[629]&m[630]&m[631]))):InitCond[644];
    m[150] = run?((((m[29]&m[632]&~m[633]&~m[634]&~m[635])|(m[29]&~m[632]&m[633]&~m[634]&~m[635])|(~m[29]&m[632]&m[633]&~m[634]&~m[635])|(m[29]&~m[632]&~m[633]&m[634]&~m[635])|(~m[29]&m[632]&~m[633]&m[634]&~m[635])|(~m[29]&~m[632]&m[633]&m[634]&~m[635])|(m[29]&~m[632]&~m[633]&~m[634]&m[635])|(~m[29]&m[632]&~m[633]&~m[634]&m[635])|(~m[29]&~m[632]&m[633]&~m[634]&m[635])|(~m[29]&~m[632]&~m[633]&m[634]&m[635]))&BiasedRNG[374])|(((m[29]&m[632]&m[633]&~m[634]&~m[635])|(m[29]&m[632]&~m[633]&m[634]&~m[635])|(m[29]&~m[632]&m[633]&m[634]&~m[635])|(~m[29]&m[632]&m[633]&m[634]&~m[635])|(m[29]&m[632]&~m[633]&~m[634]&m[635])|(m[29]&~m[632]&m[633]&~m[634]&m[635])|(~m[29]&m[632]&m[633]&~m[634]&m[635])|(m[29]&~m[632]&~m[633]&m[634]&m[635])|(~m[29]&m[632]&~m[633]&m[634]&m[635])|(~m[29]&~m[632]&m[633]&m[634]&m[635]))&~BiasedRNG[374])|((m[29]&m[632]&m[633]&m[634]&~m[635])|(m[29]&m[632]&m[633]&~m[634]&m[635])|(m[29]&m[632]&~m[633]&m[634]&m[635])|(m[29]&~m[632]&m[633]&m[634]&m[635])|(~m[29]&m[632]&m[633]&m[634]&m[635])|(m[29]&m[632]&m[633]&m[634]&m[635]))):InitCond[645];
    m[151] = run?((((m[29]&m[636]&~m[637]&~m[638]&~m[639])|(m[29]&~m[636]&m[637]&~m[638]&~m[639])|(~m[29]&m[636]&m[637]&~m[638]&~m[639])|(m[29]&~m[636]&~m[637]&m[638]&~m[639])|(~m[29]&m[636]&~m[637]&m[638]&~m[639])|(~m[29]&~m[636]&m[637]&m[638]&~m[639])|(m[29]&~m[636]&~m[637]&~m[638]&m[639])|(~m[29]&m[636]&~m[637]&~m[638]&m[639])|(~m[29]&~m[636]&m[637]&~m[638]&m[639])|(~m[29]&~m[636]&~m[637]&m[638]&m[639]))&BiasedRNG[375])|(((m[29]&m[636]&m[637]&~m[638]&~m[639])|(m[29]&m[636]&~m[637]&m[638]&~m[639])|(m[29]&~m[636]&m[637]&m[638]&~m[639])|(~m[29]&m[636]&m[637]&m[638]&~m[639])|(m[29]&m[636]&~m[637]&~m[638]&m[639])|(m[29]&~m[636]&m[637]&~m[638]&m[639])|(~m[29]&m[636]&m[637]&~m[638]&m[639])|(m[29]&~m[636]&~m[637]&m[638]&m[639])|(~m[29]&m[636]&~m[637]&m[638]&m[639])|(~m[29]&~m[636]&m[637]&m[638]&m[639]))&~BiasedRNG[375])|((m[29]&m[636]&m[637]&m[638]&~m[639])|(m[29]&m[636]&m[637]&~m[638]&m[639])|(m[29]&m[636]&~m[637]&m[638]&m[639])|(m[29]&~m[636]&m[637]&m[638]&m[639])|(~m[29]&m[636]&m[637]&m[638]&m[639])|(m[29]&m[636]&m[637]&m[638]&m[639]))):InitCond[646];
    m[152] = run?((((m[30]&m[640]&~m[641]&~m[642]&~m[643])|(m[30]&~m[640]&m[641]&~m[642]&~m[643])|(~m[30]&m[640]&m[641]&~m[642]&~m[643])|(m[30]&~m[640]&~m[641]&m[642]&~m[643])|(~m[30]&m[640]&~m[641]&m[642]&~m[643])|(~m[30]&~m[640]&m[641]&m[642]&~m[643])|(m[30]&~m[640]&~m[641]&~m[642]&m[643])|(~m[30]&m[640]&~m[641]&~m[642]&m[643])|(~m[30]&~m[640]&m[641]&~m[642]&m[643])|(~m[30]&~m[640]&~m[641]&m[642]&m[643]))&BiasedRNG[376])|(((m[30]&m[640]&m[641]&~m[642]&~m[643])|(m[30]&m[640]&~m[641]&m[642]&~m[643])|(m[30]&~m[640]&m[641]&m[642]&~m[643])|(~m[30]&m[640]&m[641]&m[642]&~m[643])|(m[30]&m[640]&~m[641]&~m[642]&m[643])|(m[30]&~m[640]&m[641]&~m[642]&m[643])|(~m[30]&m[640]&m[641]&~m[642]&m[643])|(m[30]&~m[640]&~m[641]&m[642]&m[643])|(~m[30]&m[640]&~m[641]&m[642]&m[643])|(~m[30]&~m[640]&m[641]&m[642]&m[643]))&~BiasedRNG[376])|((m[30]&m[640]&m[641]&m[642]&~m[643])|(m[30]&m[640]&m[641]&~m[642]&m[643])|(m[30]&m[640]&~m[641]&m[642]&m[643])|(m[30]&~m[640]&m[641]&m[642]&m[643])|(~m[30]&m[640]&m[641]&m[642]&m[643])|(m[30]&m[640]&m[641]&m[642]&m[643]))):InitCond[647];
    m[153] = run?((((m[30]&m[644]&~m[645]&~m[646]&~m[647])|(m[30]&~m[644]&m[645]&~m[646]&~m[647])|(~m[30]&m[644]&m[645]&~m[646]&~m[647])|(m[30]&~m[644]&~m[645]&m[646]&~m[647])|(~m[30]&m[644]&~m[645]&m[646]&~m[647])|(~m[30]&~m[644]&m[645]&m[646]&~m[647])|(m[30]&~m[644]&~m[645]&~m[646]&m[647])|(~m[30]&m[644]&~m[645]&~m[646]&m[647])|(~m[30]&~m[644]&m[645]&~m[646]&m[647])|(~m[30]&~m[644]&~m[645]&m[646]&m[647]))&BiasedRNG[377])|(((m[30]&m[644]&m[645]&~m[646]&~m[647])|(m[30]&m[644]&~m[645]&m[646]&~m[647])|(m[30]&~m[644]&m[645]&m[646]&~m[647])|(~m[30]&m[644]&m[645]&m[646]&~m[647])|(m[30]&m[644]&~m[645]&~m[646]&m[647])|(m[30]&~m[644]&m[645]&~m[646]&m[647])|(~m[30]&m[644]&m[645]&~m[646]&m[647])|(m[30]&~m[644]&~m[645]&m[646]&m[647])|(~m[30]&m[644]&~m[645]&m[646]&m[647])|(~m[30]&~m[644]&m[645]&m[646]&m[647]))&~BiasedRNG[377])|((m[30]&m[644]&m[645]&m[646]&~m[647])|(m[30]&m[644]&m[645]&~m[646]&m[647])|(m[30]&m[644]&~m[645]&m[646]&m[647])|(m[30]&~m[644]&m[645]&m[646]&m[647])|(~m[30]&m[644]&m[645]&m[646]&m[647])|(m[30]&m[644]&m[645]&m[646]&m[647]))):InitCond[648];
    m[154] = run?((((m[30]&m[648]&~m[649]&~m[650]&~m[651])|(m[30]&~m[648]&m[649]&~m[650]&~m[651])|(~m[30]&m[648]&m[649]&~m[650]&~m[651])|(m[30]&~m[648]&~m[649]&m[650]&~m[651])|(~m[30]&m[648]&~m[649]&m[650]&~m[651])|(~m[30]&~m[648]&m[649]&m[650]&~m[651])|(m[30]&~m[648]&~m[649]&~m[650]&m[651])|(~m[30]&m[648]&~m[649]&~m[650]&m[651])|(~m[30]&~m[648]&m[649]&~m[650]&m[651])|(~m[30]&~m[648]&~m[649]&m[650]&m[651]))&BiasedRNG[378])|(((m[30]&m[648]&m[649]&~m[650]&~m[651])|(m[30]&m[648]&~m[649]&m[650]&~m[651])|(m[30]&~m[648]&m[649]&m[650]&~m[651])|(~m[30]&m[648]&m[649]&m[650]&~m[651])|(m[30]&m[648]&~m[649]&~m[650]&m[651])|(m[30]&~m[648]&m[649]&~m[650]&m[651])|(~m[30]&m[648]&m[649]&~m[650]&m[651])|(m[30]&~m[648]&~m[649]&m[650]&m[651])|(~m[30]&m[648]&~m[649]&m[650]&m[651])|(~m[30]&~m[648]&m[649]&m[650]&m[651]))&~BiasedRNG[378])|((m[30]&m[648]&m[649]&m[650]&~m[651])|(m[30]&m[648]&m[649]&~m[650]&m[651])|(m[30]&m[648]&~m[649]&m[650]&m[651])|(m[30]&~m[648]&m[649]&m[650]&m[651])|(~m[30]&m[648]&m[649]&m[650]&m[651])|(m[30]&m[648]&m[649]&m[650]&m[651]))):InitCond[649];
    m[155] = run?((((m[30]&m[652]&~m[653]&~m[654]&~m[655])|(m[30]&~m[652]&m[653]&~m[654]&~m[655])|(~m[30]&m[652]&m[653]&~m[654]&~m[655])|(m[30]&~m[652]&~m[653]&m[654]&~m[655])|(~m[30]&m[652]&~m[653]&m[654]&~m[655])|(~m[30]&~m[652]&m[653]&m[654]&~m[655])|(m[30]&~m[652]&~m[653]&~m[654]&m[655])|(~m[30]&m[652]&~m[653]&~m[654]&m[655])|(~m[30]&~m[652]&m[653]&~m[654]&m[655])|(~m[30]&~m[652]&~m[653]&m[654]&m[655]))&BiasedRNG[379])|(((m[30]&m[652]&m[653]&~m[654]&~m[655])|(m[30]&m[652]&~m[653]&m[654]&~m[655])|(m[30]&~m[652]&m[653]&m[654]&~m[655])|(~m[30]&m[652]&m[653]&m[654]&~m[655])|(m[30]&m[652]&~m[653]&~m[654]&m[655])|(m[30]&~m[652]&m[653]&~m[654]&m[655])|(~m[30]&m[652]&m[653]&~m[654]&m[655])|(m[30]&~m[652]&~m[653]&m[654]&m[655])|(~m[30]&m[652]&~m[653]&m[654]&m[655])|(~m[30]&~m[652]&m[653]&m[654]&m[655]))&~BiasedRNG[379])|((m[30]&m[652]&m[653]&m[654]&~m[655])|(m[30]&m[652]&m[653]&~m[654]&m[655])|(m[30]&m[652]&~m[653]&m[654]&m[655])|(m[30]&~m[652]&m[653]&m[654]&m[655])|(~m[30]&m[652]&m[653]&m[654]&m[655])|(m[30]&m[652]&m[653]&m[654]&m[655]))):InitCond[650];
    m[156] = run?((((m[31]&m[656]&~m[657]&~m[658]&~m[659])|(m[31]&~m[656]&m[657]&~m[658]&~m[659])|(~m[31]&m[656]&m[657]&~m[658]&~m[659])|(m[31]&~m[656]&~m[657]&m[658]&~m[659])|(~m[31]&m[656]&~m[657]&m[658]&~m[659])|(~m[31]&~m[656]&m[657]&m[658]&~m[659])|(m[31]&~m[656]&~m[657]&~m[658]&m[659])|(~m[31]&m[656]&~m[657]&~m[658]&m[659])|(~m[31]&~m[656]&m[657]&~m[658]&m[659])|(~m[31]&~m[656]&~m[657]&m[658]&m[659]))&BiasedRNG[380])|(((m[31]&m[656]&m[657]&~m[658]&~m[659])|(m[31]&m[656]&~m[657]&m[658]&~m[659])|(m[31]&~m[656]&m[657]&m[658]&~m[659])|(~m[31]&m[656]&m[657]&m[658]&~m[659])|(m[31]&m[656]&~m[657]&~m[658]&m[659])|(m[31]&~m[656]&m[657]&~m[658]&m[659])|(~m[31]&m[656]&m[657]&~m[658]&m[659])|(m[31]&~m[656]&~m[657]&m[658]&m[659])|(~m[31]&m[656]&~m[657]&m[658]&m[659])|(~m[31]&~m[656]&m[657]&m[658]&m[659]))&~BiasedRNG[380])|((m[31]&m[656]&m[657]&m[658]&~m[659])|(m[31]&m[656]&m[657]&~m[658]&m[659])|(m[31]&m[656]&~m[657]&m[658]&m[659])|(m[31]&~m[656]&m[657]&m[658]&m[659])|(~m[31]&m[656]&m[657]&m[658]&m[659])|(m[31]&m[656]&m[657]&m[658]&m[659]))):InitCond[651];
    m[157] = run?((((m[31]&m[660]&~m[661]&~m[662]&~m[663])|(m[31]&~m[660]&m[661]&~m[662]&~m[663])|(~m[31]&m[660]&m[661]&~m[662]&~m[663])|(m[31]&~m[660]&~m[661]&m[662]&~m[663])|(~m[31]&m[660]&~m[661]&m[662]&~m[663])|(~m[31]&~m[660]&m[661]&m[662]&~m[663])|(m[31]&~m[660]&~m[661]&~m[662]&m[663])|(~m[31]&m[660]&~m[661]&~m[662]&m[663])|(~m[31]&~m[660]&m[661]&~m[662]&m[663])|(~m[31]&~m[660]&~m[661]&m[662]&m[663]))&BiasedRNG[381])|(((m[31]&m[660]&m[661]&~m[662]&~m[663])|(m[31]&m[660]&~m[661]&m[662]&~m[663])|(m[31]&~m[660]&m[661]&m[662]&~m[663])|(~m[31]&m[660]&m[661]&m[662]&~m[663])|(m[31]&m[660]&~m[661]&~m[662]&m[663])|(m[31]&~m[660]&m[661]&~m[662]&m[663])|(~m[31]&m[660]&m[661]&~m[662]&m[663])|(m[31]&~m[660]&~m[661]&m[662]&m[663])|(~m[31]&m[660]&~m[661]&m[662]&m[663])|(~m[31]&~m[660]&m[661]&m[662]&m[663]))&~BiasedRNG[381])|((m[31]&m[660]&m[661]&m[662]&~m[663])|(m[31]&m[660]&m[661]&~m[662]&m[663])|(m[31]&m[660]&~m[661]&m[662]&m[663])|(m[31]&~m[660]&m[661]&m[662]&m[663])|(~m[31]&m[660]&m[661]&m[662]&m[663])|(m[31]&m[660]&m[661]&m[662]&m[663]))):InitCond[652];
    m[158] = run?((((m[31]&m[664]&~m[665]&~m[666]&~m[667])|(m[31]&~m[664]&m[665]&~m[666]&~m[667])|(~m[31]&m[664]&m[665]&~m[666]&~m[667])|(m[31]&~m[664]&~m[665]&m[666]&~m[667])|(~m[31]&m[664]&~m[665]&m[666]&~m[667])|(~m[31]&~m[664]&m[665]&m[666]&~m[667])|(m[31]&~m[664]&~m[665]&~m[666]&m[667])|(~m[31]&m[664]&~m[665]&~m[666]&m[667])|(~m[31]&~m[664]&m[665]&~m[666]&m[667])|(~m[31]&~m[664]&~m[665]&m[666]&m[667]))&BiasedRNG[382])|(((m[31]&m[664]&m[665]&~m[666]&~m[667])|(m[31]&m[664]&~m[665]&m[666]&~m[667])|(m[31]&~m[664]&m[665]&m[666]&~m[667])|(~m[31]&m[664]&m[665]&m[666]&~m[667])|(m[31]&m[664]&~m[665]&~m[666]&m[667])|(m[31]&~m[664]&m[665]&~m[666]&m[667])|(~m[31]&m[664]&m[665]&~m[666]&m[667])|(m[31]&~m[664]&~m[665]&m[666]&m[667])|(~m[31]&m[664]&~m[665]&m[666]&m[667])|(~m[31]&~m[664]&m[665]&m[666]&m[667]))&~BiasedRNG[382])|((m[31]&m[664]&m[665]&m[666]&~m[667])|(m[31]&m[664]&m[665]&~m[666]&m[667])|(m[31]&m[664]&~m[665]&m[666]&m[667])|(m[31]&~m[664]&m[665]&m[666]&m[667])|(~m[31]&m[664]&m[665]&m[666]&m[667])|(m[31]&m[664]&m[665]&m[666]&m[667]))):InitCond[653];
    m[159] = run?((((m[31]&m[668]&~m[669]&~m[670]&~m[671])|(m[31]&~m[668]&m[669]&~m[670]&~m[671])|(~m[31]&m[668]&m[669]&~m[670]&~m[671])|(m[31]&~m[668]&~m[669]&m[670]&~m[671])|(~m[31]&m[668]&~m[669]&m[670]&~m[671])|(~m[31]&~m[668]&m[669]&m[670]&~m[671])|(m[31]&~m[668]&~m[669]&~m[670]&m[671])|(~m[31]&m[668]&~m[669]&~m[670]&m[671])|(~m[31]&~m[668]&m[669]&~m[670]&m[671])|(~m[31]&~m[668]&~m[669]&m[670]&m[671]))&BiasedRNG[383])|(((m[31]&m[668]&m[669]&~m[670]&~m[671])|(m[31]&m[668]&~m[669]&m[670]&~m[671])|(m[31]&~m[668]&m[669]&m[670]&~m[671])|(~m[31]&m[668]&m[669]&m[670]&~m[671])|(m[31]&m[668]&~m[669]&~m[670]&m[671])|(m[31]&~m[668]&m[669]&~m[670]&m[671])|(~m[31]&m[668]&m[669]&~m[670]&m[671])|(m[31]&~m[668]&~m[669]&m[670]&m[671])|(~m[31]&m[668]&~m[669]&m[670]&m[671])|(~m[31]&~m[668]&m[669]&m[670]&m[671]))&~BiasedRNG[383])|((m[31]&m[668]&m[669]&m[670]&~m[671])|(m[31]&m[668]&m[669]&~m[670]&m[671])|(m[31]&m[668]&~m[669]&m[670]&m[671])|(m[31]&~m[668]&m[669]&m[670]&m[671])|(~m[31]&m[668]&m[669]&m[670]&m[671])|(m[31]&m[668]&m[669]&m[670]&m[671]))):InitCond[654];
    m[673] = run?((((m[176]&~m[417]&m[928])|(~m[176]&m[417]&m[928]))&BiasedRNG[384])|(((m[176]&m[417]&~m[928]))&~BiasedRNG[384])|((m[176]&m[417]&m[928]))):InitCond[655];
    m[674] = run?((((m[192]&~m[418]&m[933])|(~m[192]&m[418]&m[933]))&BiasedRNG[385])|(((m[192]&m[418]&~m[933]))&~BiasedRNG[385])|((m[192]&m[418]&m[933]))):InitCond[656];
    m[675] = run?((((m[208]&~m[419]&m[943])|(~m[208]&m[419]&m[943]))&BiasedRNG[386])|(((m[208]&m[419]&~m[943]))&~BiasedRNG[386])|((m[208]&m[419]&m[943]))):InitCond[657];
    m[676] = run?((((m[224]&~m[420]&m[958])|(~m[224]&m[420]&m[958]))&BiasedRNG[387])|(((m[224]&m[420]&~m[958]))&~BiasedRNG[387])|((m[224]&m[420]&m[958]))):InitCond[658];
    m[677] = run?((((m[240]&~m[421]&m[978])|(~m[240]&m[421]&m[978]))&BiasedRNG[388])|(((m[240]&m[421]&~m[978]))&~BiasedRNG[388])|((m[240]&m[421]&m[978]))):InitCond[659];
    m[678] = run?((((m[256]&~m[422]&m[1003])|(~m[256]&m[422]&m[1003]))&BiasedRNG[389])|(((m[256]&m[422]&~m[1003]))&~BiasedRNG[389])|((m[256]&m[422]&m[1003]))):InitCond[660];
    m[679] = run?((((m[272]&~m[423]&m[1033])|(~m[272]&m[423]&m[1033]))&BiasedRNG[390])|(((m[272]&m[423]&~m[1033]))&~BiasedRNG[390])|((m[272]&m[423]&m[1033]))):InitCond[661];
    m[680] = run?((((m[288]&~m[424]&m[1068])|(~m[288]&m[424]&m[1068]))&BiasedRNG[391])|(((m[288]&m[424]&~m[1068]))&~BiasedRNG[391])|((m[288]&m[424]&m[1068]))):InitCond[662];
    m[681] = run?((((m[304]&~m[425]&m[1108])|(~m[304]&m[425]&m[1108]))&BiasedRNG[392])|(((m[304]&m[425]&~m[1108]))&~BiasedRNG[392])|((m[304]&m[425]&m[1108]))):InitCond[663];
    m[682] = run?((((m[320]&~m[426]&m[1153])|(~m[320]&m[426]&m[1153]))&BiasedRNG[393])|(((m[320]&m[426]&~m[1153]))&~BiasedRNG[393])|((m[320]&m[426]&m[1153]))):InitCond[664];
    m[683] = run?((((m[336]&~m[427]&m[1203])|(~m[336]&m[427]&m[1203]))&BiasedRNG[394])|(((m[336]&m[427]&~m[1203]))&~BiasedRNG[394])|((m[336]&m[427]&m[1203]))):InitCond[665];
    m[684] = run?((((m[352]&~m[428]&m[1258])|(~m[352]&m[428]&m[1258]))&BiasedRNG[395])|(((m[352]&m[428]&~m[1258]))&~BiasedRNG[395])|((m[352]&m[428]&m[1258]))):InitCond[666];
    m[685] = run?((((m[368]&~m[429]&m[1318])|(~m[368]&m[429]&m[1318]))&BiasedRNG[396])|(((m[368]&m[429]&~m[1318]))&~BiasedRNG[396])|((m[368]&m[429]&m[1318]))):InitCond[667];
    m[686] = run?((((m[384]&~m[430]&m[1383])|(~m[384]&m[430]&m[1383]))&BiasedRNG[397])|(((m[384]&m[430]&~m[1383]))&~BiasedRNG[397])|((m[384]&m[430]&m[1383]))):InitCond[668];
    m[687] = run?((((m[400]&~m[431]&m[1453])|(~m[400]&m[431]&m[1453]))&BiasedRNG[398])|(((m[400]&m[431]&~m[1453]))&~BiasedRNG[398])|((m[400]&m[431]&m[1453]))):InitCond[669];
    m[688] = run?((((m[161]&~m[432]&m[929])|(~m[161]&m[432]&m[929]))&BiasedRNG[399])|(((m[161]&m[432]&~m[929]))&~BiasedRNG[399])|((m[161]&m[432]&m[929]))):InitCond[670];
    m[689] = run?((((m[177]&~m[433]&m[934])|(~m[177]&m[433]&m[934]))&BiasedRNG[400])|(((m[177]&m[433]&~m[934]))&~BiasedRNG[400])|((m[177]&m[433]&m[934]))):InitCond[671];
    m[690] = run?((((m[193]&~m[434]&m[944])|(~m[193]&m[434]&m[944]))&BiasedRNG[401])|(((m[193]&m[434]&~m[944]))&~BiasedRNG[401])|((m[193]&m[434]&m[944]))):InitCond[672];
    m[691] = run?((((m[209]&~m[435]&m[959])|(~m[209]&m[435]&m[959]))&BiasedRNG[402])|(((m[209]&m[435]&~m[959]))&~BiasedRNG[402])|((m[209]&m[435]&m[959]))):InitCond[673];
    m[692] = run?((((m[225]&~m[436]&m[979])|(~m[225]&m[436]&m[979]))&BiasedRNG[403])|(((m[225]&m[436]&~m[979]))&~BiasedRNG[403])|((m[225]&m[436]&m[979]))):InitCond[674];
    m[693] = run?((((m[241]&~m[437]&m[1004])|(~m[241]&m[437]&m[1004]))&BiasedRNG[404])|(((m[241]&m[437]&~m[1004]))&~BiasedRNG[404])|((m[241]&m[437]&m[1004]))):InitCond[675];
    m[694] = run?((((m[257]&~m[438]&m[1034])|(~m[257]&m[438]&m[1034]))&BiasedRNG[405])|(((m[257]&m[438]&~m[1034]))&~BiasedRNG[405])|((m[257]&m[438]&m[1034]))):InitCond[676];
    m[695] = run?((((m[273]&~m[439]&m[1069])|(~m[273]&m[439]&m[1069]))&BiasedRNG[406])|(((m[273]&m[439]&~m[1069]))&~BiasedRNG[406])|((m[273]&m[439]&m[1069]))):InitCond[677];
    m[696] = run?((((m[289]&~m[440]&m[1109])|(~m[289]&m[440]&m[1109]))&BiasedRNG[407])|(((m[289]&m[440]&~m[1109]))&~BiasedRNG[407])|((m[289]&m[440]&m[1109]))):InitCond[678];
    m[697] = run?((((m[305]&~m[441]&m[1154])|(~m[305]&m[441]&m[1154]))&BiasedRNG[408])|(((m[305]&m[441]&~m[1154]))&~BiasedRNG[408])|((m[305]&m[441]&m[1154]))):InitCond[679];
    m[698] = run?((((m[321]&~m[442]&m[1204])|(~m[321]&m[442]&m[1204]))&BiasedRNG[409])|(((m[321]&m[442]&~m[1204]))&~BiasedRNG[409])|((m[321]&m[442]&m[1204]))):InitCond[680];
    m[699] = run?((((m[337]&~m[443]&m[1259])|(~m[337]&m[443]&m[1259]))&BiasedRNG[410])|(((m[337]&m[443]&~m[1259]))&~BiasedRNG[410])|((m[337]&m[443]&m[1259]))):InitCond[681];
    m[700] = run?((((m[353]&~m[444]&m[1319])|(~m[353]&m[444]&m[1319]))&BiasedRNG[411])|(((m[353]&m[444]&~m[1319]))&~BiasedRNG[411])|((m[353]&m[444]&m[1319]))):InitCond[682];
    m[701] = run?((((m[369]&~m[445]&m[1384])|(~m[369]&m[445]&m[1384]))&BiasedRNG[412])|(((m[369]&m[445]&~m[1384]))&~BiasedRNG[412])|((m[369]&m[445]&m[1384]))):InitCond[683];
    m[702] = run?((((m[385]&~m[446]&m[1454])|(~m[385]&m[446]&m[1454]))&BiasedRNG[413])|(((m[385]&m[446]&~m[1454]))&~BiasedRNG[413])|((m[385]&m[446]&m[1454]))):InitCond[684];
    m[703] = run?((((m[401]&~m[447]&m[1529])|(~m[401]&m[447]&m[1529]))&BiasedRNG[414])|(((m[401]&m[447]&~m[1529]))&~BiasedRNG[414])|((m[401]&m[447]&m[1529]))):InitCond[685];
    m[704] = run?((((m[162]&~m[448]&m[939])|(~m[162]&m[448]&m[939]))&BiasedRNG[415])|(((m[162]&m[448]&~m[939]))&~BiasedRNG[415])|((m[162]&m[448]&m[939]))):InitCond[686];
    m[705] = run?((((m[178]&~m[449]&m[949])|(~m[178]&m[449]&m[949]))&BiasedRNG[416])|(((m[178]&m[449]&~m[949]))&~BiasedRNG[416])|((m[178]&m[449]&m[949]))):InitCond[687];
    m[706] = run?((((m[194]&~m[450]&m[964])|(~m[194]&m[450]&m[964]))&BiasedRNG[417])|(((m[194]&m[450]&~m[964]))&~BiasedRNG[417])|((m[194]&m[450]&m[964]))):InitCond[688];
    m[707] = run?((((m[210]&~m[451]&m[984])|(~m[210]&m[451]&m[984]))&BiasedRNG[418])|(((m[210]&m[451]&~m[984]))&~BiasedRNG[418])|((m[210]&m[451]&m[984]))):InitCond[689];
    m[708] = run?((((m[226]&~m[452]&m[1009])|(~m[226]&m[452]&m[1009]))&BiasedRNG[419])|(((m[226]&m[452]&~m[1009]))&~BiasedRNG[419])|((m[226]&m[452]&m[1009]))):InitCond[690];
    m[709] = run?((((m[242]&~m[453]&m[1039])|(~m[242]&m[453]&m[1039]))&BiasedRNG[420])|(((m[242]&m[453]&~m[1039]))&~BiasedRNG[420])|((m[242]&m[453]&m[1039]))):InitCond[691];
    m[710] = run?((((m[258]&~m[454]&m[1074])|(~m[258]&m[454]&m[1074]))&BiasedRNG[421])|(((m[258]&m[454]&~m[1074]))&~BiasedRNG[421])|((m[258]&m[454]&m[1074]))):InitCond[692];
    m[711] = run?((((m[274]&~m[455]&m[1114])|(~m[274]&m[455]&m[1114]))&BiasedRNG[422])|(((m[274]&m[455]&~m[1114]))&~BiasedRNG[422])|((m[274]&m[455]&m[1114]))):InitCond[693];
    m[712] = run?((((m[290]&~m[456]&m[1159])|(~m[290]&m[456]&m[1159]))&BiasedRNG[423])|(((m[290]&m[456]&~m[1159]))&~BiasedRNG[423])|((m[290]&m[456]&m[1159]))):InitCond[694];
    m[713] = run?((((m[306]&~m[457]&m[1209])|(~m[306]&m[457]&m[1209]))&BiasedRNG[424])|(((m[306]&m[457]&~m[1209]))&~BiasedRNG[424])|((m[306]&m[457]&m[1209]))):InitCond[695];
    m[714] = run?((((m[322]&~m[458]&m[1264])|(~m[322]&m[458]&m[1264]))&BiasedRNG[425])|(((m[322]&m[458]&~m[1264]))&~BiasedRNG[425])|((m[322]&m[458]&m[1264]))):InitCond[696];
    m[715] = run?((((m[338]&~m[459]&m[1324])|(~m[338]&m[459]&m[1324]))&BiasedRNG[426])|(((m[338]&m[459]&~m[1324]))&~BiasedRNG[426])|((m[338]&m[459]&m[1324]))):InitCond[697];
    m[716] = run?((((m[354]&~m[460]&m[1389])|(~m[354]&m[460]&m[1389]))&BiasedRNG[427])|(((m[354]&m[460]&~m[1389]))&~BiasedRNG[427])|((m[354]&m[460]&m[1389]))):InitCond[698];
    m[717] = run?((((m[370]&~m[461]&m[1459])|(~m[370]&m[461]&m[1459]))&BiasedRNG[428])|(((m[370]&m[461]&~m[1459]))&~BiasedRNG[428])|((m[370]&m[461]&m[1459]))):InitCond[699];
    m[718] = run?((((m[386]&~m[462]&m[1534])|(~m[386]&m[462]&m[1534]))&BiasedRNG[429])|(((m[386]&m[462]&~m[1534]))&~BiasedRNG[429])|((m[386]&m[462]&m[1534]))):InitCond[700];
    m[719] = run?((((m[402]&~m[463]&m[1604])|(~m[402]&m[463]&m[1604]))&BiasedRNG[430])|(((m[402]&m[463]&~m[1604]))&~BiasedRNG[430])|((m[402]&m[463]&m[1604]))):InitCond[701];
    m[720] = run?((((m[163]&~m[464]&m[954])|(~m[163]&m[464]&m[954]))&BiasedRNG[431])|(((m[163]&m[464]&~m[954]))&~BiasedRNG[431])|((m[163]&m[464]&m[954]))):InitCond[702];
    m[721] = run?((((m[179]&~m[465]&m[969])|(~m[179]&m[465]&m[969]))&BiasedRNG[432])|(((m[179]&m[465]&~m[969]))&~BiasedRNG[432])|((m[179]&m[465]&m[969]))):InitCond[703];
    m[722] = run?((((m[195]&~m[466]&m[989])|(~m[195]&m[466]&m[989]))&BiasedRNG[433])|(((m[195]&m[466]&~m[989]))&~BiasedRNG[433])|((m[195]&m[466]&m[989]))):InitCond[704];
    m[723] = run?((((m[211]&~m[467]&m[1014])|(~m[211]&m[467]&m[1014]))&BiasedRNG[434])|(((m[211]&m[467]&~m[1014]))&~BiasedRNG[434])|((m[211]&m[467]&m[1014]))):InitCond[705];
    m[724] = run?((((m[227]&~m[468]&m[1044])|(~m[227]&m[468]&m[1044]))&BiasedRNG[435])|(((m[227]&m[468]&~m[1044]))&~BiasedRNG[435])|((m[227]&m[468]&m[1044]))):InitCond[706];
    m[725] = run?((((m[243]&~m[469]&m[1079])|(~m[243]&m[469]&m[1079]))&BiasedRNG[436])|(((m[243]&m[469]&~m[1079]))&~BiasedRNG[436])|((m[243]&m[469]&m[1079]))):InitCond[707];
    m[726] = run?((((m[259]&~m[470]&m[1119])|(~m[259]&m[470]&m[1119]))&BiasedRNG[437])|(((m[259]&m[470]&~m[1119]))&~BiasedRNG[437])|((m[259]&m[470]&m[1119]))):InitCond[708];
    m[727] = run?((((m[275]&~m[471]&m[1164])|(~m[275]&m[471]&m[1164]))&BiasedRNG[438])|(((m[275]&m[471]&~m[1164]))&~BiasedRNG[438])|((m[275]&m[471]&m[1164]))):InitCond[709];
    m[728] = run?((((m[291]&~m[472]&m[1214])|(~m[291]&m[472]&m[1214]))&BiasedRNG[439])|(((m[291]&m[472]&~m[1214]))&~BiasedRNG[439])|((m[291]&m[472]&m[1214]))):InitCond[710];
    m[729] = run?((((m[307]&~m[473]&m[1269])|(~m[307]&m[473]&m[1269]))&BiasedRNG[440])|(((m[307]&m[473]&~m[1269]))&~BiasedRNG[440])|((m[307]&m[473]&m[1269]))):InitCond[711];
    m[730] = run?((((m[323]&~m[474]&m[1329])|(~m[323]&m[474]&m[1329]))&BiasedRNG[441])|(((m[323]&m[474]&~m[1329]))&~BiasedRNG[441])|((m[323]&m[474]&m[1329]))):InitCond[712];
    m[731] = run?((((m[339]&~m[475]&m[1394])|(~m[339]&m[475]&m[1394]))&BiasedRNG[442])|(((m[339]&m[475]&~m[1394]))&~BiasedRNG[442])|((m[339]&m[475]&m[1394]))):InitCond[713];
    m[732] = run?((((m[355]&~m[476]&m[1464])|(~m[355]&m[476]&m[1464]))&BiasedRNG[443])|(((m[355]&m[476]&~m[1464]))&~BiasedRNG[443])|((m[355]&m[476]&m[1464]))):InitCond[714];
    m[733] = run?((((m[371]&~m[477]&m[1539])|(~m[371]&m[477]&m[1539]))&BiasedRNG[444])|(((m[371]&m[477]&~m[1539]))&~BiasedRNG[444])|((m[371]&m[477]&m[1539]))):InitCond[715];
    m[734] = run?((((m[387]&~m[478]&m[1609])|(~m[387]&m[478]&m[1609]))&BiasedRNG[445])|(((m[387]&m[478]&~m[1609]))&~BiasedRNG[445])|((m[387]&m[478]&m[1609]))):InitCond[716];
    m[735] = run?((((m[403]&~m[479]&m[1674])|(~m[403]&m[479]&m[1674]))&BiasedRNG[446])|(((m[403]&m[479]&~m[1674]))&~BiasedRNG[446])|((m[403]&m[479]&m[1674]))):InitCond[717];
    m[736] = run?((((m[164]&~m[480]&m[974])|(~m[164]&m[480]&m[974]))&BiasedRNG[447])|(((m[164]&m[480]&~m[974]))&~BiasedRNG[447])|((m[164]&m[480]&m[974]))):InitCond[718];
    m[737] = run?((((m[180]&~m[481]&m[994])|(~m[180]&m[481]&m[994]))&BiasedRNG[448])|(((m[180]&m[481]&~m[994]))&~BiasedRNG[448])|((m[180]&m[481]&m[994]))):InitCond[719];
    m[738] = run?((((m[196]&~m[482]&m[1019])|(~m[196]&m[482]&m[1019]))&BiasedRNG[449])|(((m[196]&m[482]&~m[1019]))&~BiasedRNG[449])|((m[196]&m[482]&m[1019]))):InitCond[720];
    m[739] = run?((((m[212]&~m[483]&m[1049])|(~m[212]&m[483]&m[1049]))&BiasedRNG[450])|(((m[212]&m[483]&~m[1049]))&~BiasedRNG[450])|((m[212]&m[483]&m[1049]))):InitCond[721];
    m[740] = run?((((m[228]&~m[484]&m[1084])|(~m[228]&m[484]&m[1084]))&BiasedRNG[451])|(((m[228]&m[484]&~m[1084]))&~BiasedRNG[451])|((m[228]&m[484]&m[1084]))):InitCond[722];
    m[741] = run?((((m[244]&~m[485]&m[1124])|(~m[244]&m[485]&m[1124]))&BiasedRNG[452])|(((m[244]&m[485]&~m[1124]))&~BiasedRNG[452])|((m[244]&m[485]&m[1124]))):InitCond[723];
    m[742] = run?((((m[260]&~m[486]&m[1169])|(~m[260]&m[486]&m[1169]))&BiasedRNG[453])|(((m[260]&m[486]&~m[1169]))&~BiasedRNG[453])|((m[260]&m[486]&m[1169]))):InitCond[724];
    m[743] = run?((((m[276]&~m[487]&m[1219])|(~m[276]&m[487]&m[1219]))&BiasedRNG[454])|(((m[276]&m[487]&~m[1219]))&~BiasedRNG[454])|((m[276]&m[487]&m[1219]))):InitCond[725];
    m[744] = run?((((m[292]&~m[488]&m[1274])|(~m[292]&m[488]&m[1274]))&BiasedRNG[455])|(((m[292]&m[488]&~m[1274]))&~BiasedRNG[455])|((m[292]&m[488]&m[1274]))):InitCond[726];
    m[745] = run?((((m[308]&~m[489]&m[1334])|(~m[308]&m[489]&m[1334]))&BiasedRNG[456])|(((m[308]&m[489]&~m[1334]))&~BiasedRNG[456])|((m[308]&m[489]&m[1334]))):InitCond[727];
    m[746] = run?((((m[324]&~m[490]&m[1399])|(~m[324]&m[490]&m[1399]))&BiasedRNG[457])|(((m[324]&m[490]&~m[1399]))&~BiasedRNG[457])|((m[324]&m[490]&m[1399]))):InitCond[728];
    m[747] = run?((((m[340]&~m[491]&m[1469])|(~m[340]&m[491]&m[1469]))&BiasedRNG[458])|(((m[340]&m[491]&~m[1469]))&~BiasedRNG[458])|((m[340]&m[491]&m[1469]))):InitCond[729];
    m[748] = run?((((m[356]&~m[492]&m[1544])|(~m[356]&m[492]&m[1544]))&BiasedRNG[459])|(((m[356]&m[492]&~m[1544]))&~BiasedRNG[459])|((m[356]&m[492]&m[1544]))):InitCond[730];
    m[749] = run?((((m[372]&~m[493]&m[1614])|(~m[372]&m[493]&m[1614]))&BiasedRNG[460])|(((m[372]&m[493]&~m[1614]))&~BiasedRNG[460])|((m[372]&m[493]&m[1614]))):InitCond[731];
    m[750] = run?((((m[388]&~m[494]&m[1679])|(~m[388]&m[494]&m[1679]))&BiasedRNG[461])|(((m[388]&m[494]&~m[1679]))&~BiasedRNG[461])|((m[388]&m[494]&m[1679]))):InitCond[732];
    m[751] = run?((((m[404]&~m[495]&m[1739])|(~m[404]&m[495]&m[1739]))&BiasedRNG[462])|(((m[404]&m[495]&~m[1739]))&~BiasedRNG[462])|((m[404]&m[495]&m[1739]))):InitCond[733];
    m[752] = run?((((m[165]&~m[496]&m[999])|(~m[165]&m[496]&m[999]))&BiasedRNG[463])|(((m[165]&m[496]&~m[999]))&~BiasedRNG[463])|((m[165]&m[496]&m[999]))):InitCond[734];
    m[753] = run?((((m[181]&~m[497]&m[1024])|(~m[181]&m[497]&m[1024]))&BiasedRNG[464])|(((m[181]&m[497]&~m[1024]))&~BiasedRNG[464])|((m[181]&m[497]&m[1024]))):InitCond[735];
    m[754] = run?((((m[197]&~m[498]&m[1054])|(~m[197]&m[498]&m[1054]))&BiasedRNG[465])|(((m[197]&m[498]&~m[1054]))&~BiasedRNG[465])|((m[197]&m[498]&m[1054]))):InitCond[736];
    m[755] = run?((((m[213]&~m[499]&m[1089])|(~m[213]&m[499]&m[1089]))&BiasedRNG[466])|(((m[213]&m[499]&~m[1089]))&~BiasedRNG[466])|((m[213]&m[499]&m[1089]))):InitCond[737];
    m[756] = run?((((m[229]&~m[500]&m[1129])|(~m[229]&m[500]&m[1129]))&BiasedRNG[467])|(((m[229]&m[500]&~m[1129]))&~BiasedRNG[467])|((m[229]&m[500]&m[1129]))):InitCond[738];
    m[757] = run?((((m[245]&~m[501]&m[1174])|(~m[245]&m[501]&m[1174]))&BiasedRNG[468])|(((m[245]&m[501]&~m[1174]))&~BiasedRNG[468])|((m[245]&m[501]&m[1174]))):InitCond[739];
    m[758] = run?((((m[261]&~m[502]&m[1224])|(~m[261]&m[502]&m[1224]))&BiasedRNG[469])|(((m[261]&m[502]&~m[1224]))&~BiasedRNG[469])|((m[261]&m[502]&m[1224]))):InitCond[740];
    m[759] = run?((((m[277]&~m[503]&m[1279])|(~m[277]&m[503]&m[1279]))&BiasedRNG[470])|(((m[277]&m[503]&~m[1279]))&~BiasedRNG[470])|((m[277]&m[503]&m[1279]))):InitCond[741];
    m[760] = run?((((m[293]&~m[504]&m[1339])|(~m[293]&m[504]&m[1339]))&BiasedRNG[471])|(((m[293]&m[504]&~m[1339]))&~BiasedRNG[471])|((m[293]&m[504]&m[1339]))):InitCond[742];
    m[761] = run?((((m[309]&~m[505]&m[1404])|(~m[309]&m[505]&m[1404]))&BiasedRNG[472])|(((m[309]&m[505]&~m[1404]))&~BiasedRNG[472])|((m[309]&m[505]&m[1404]))):InitCond[743];
    m[762] = run?((((m[325]&~m[506]&m[1474])|(~m[325]&m[506]&m[1474]))&BiasedRNG[473])|(((m[325]&m[506]&~m[1474]))&~BiasedRNG[473])|((m[325]&m[506]&m[1474]))):InitCond[744];
    m[763] = run?((((m[341]&~m[507]&m[1549])|(~m[341]&m[507]&m[1549]))&BiasedRNG[474])|(((m[341]&m[507]&~m[1549]))&~BiasedRNG[474])|((m[341]&m[507]&m[1549]))):InitCond[745];
    m[764] = run?((((m[357]&~m[508]&m[1619])|(~m[357]&m[508]&m[1619]))&BiasedRNG[475])|(((m[357]&m[508]&~m[1619]))&~BiasedRNG[475])|((m[357]&m[508]&m[1619]))):InitCond[746];
    m[765] = run?((((m[373]&~m[509]&m[1684])|(~m[373]&m[509]&m[1684]))&BiasedRNG[476])|(((m[373]&m[509]&~m[1684]))&~BiasedRNG[476])|((m[373]&m[509]&m[1684]))):InitCond[747];
    m[766] = run?((((m[389]&~m[510]&m[1744])|(~m[389]&m[510]&m[1744]))&BiasedRNG[477])|(((m[389]&m[510]&~m[1744]))&~BiasedRNG[477])|((m[389]&m[510]&m[1744]))):InitCond[748];
    m[767] = run?((((m[405]&~m[511]&m[1799])|(~m[405]&m[511]&m[1799]))&BiasedRNG[478])|(((m[405]&m[511]&~m[1799]))&~BiasedRNG[478])|((m[405]&m[511]&m[1799]))):InitCond[749];
    m[768] = run?((((m[166]&~m[512]&m[1029])|(~m[166]&m[512]&m[1029]))&BiasedRNG[479])|(((m[166]&m[512]&~m[1029]))&~BiasedRNG[479])|((m[166]&m[512]&m[1029]))):InitCond[750];
    m[769] = run?((((m[182]&~m[513]&m[1059])|(~m[182]&m[513]&m[1059]))&BiasedRNG[480])|(((m[182]&m[513]&~m[1059]))&~BiasedRNG[480])|((m[182]&m[513]&m[1059]))):InitCond[751];
    m[770] = run?((((m[198]&~m[514]&m[1094])|(~m[198]&m[514]&m[1094]))&BiasedRNG[481])|(((m[198]&m[514]&~m[1094]))&~BiasedRNG[481])|((m[198]&m[514]&m[1094]))):InitCond[752];
    m[771] = run?((((m[214]&~m[515]&m[1134])|(~m[214]&m[515]&m[1134]))&BiasedRNG[482])|(((m[214]&m[515]&~m[1134]))&~BiasedRNG[482])|((m[214]&m[515]&m[1134]))):InitCond[753];
    m[772] = run?((((m[230]&~m[516]&m[1179])|(~m[230]&m[516]&m[1179]))&BiasedRNG[483])|(((m[230]&m[516]&~m[1179]))&~BiasedRNG[483])|((m[230]&m[516]&m[1179]))):InitCond[754];
    m[773] = run?((((m[246]&~m[517]&m[1229])|(~m[246]&m[517]&m[1229]))&BiasedRNG[484])|(((m[246]&m[517]&~m[1229]))&~BiasedRNG[484])|((m[246]&m[517]&m[1229]))):InitCond[755];
    m[774] = run?((((m[262]&~m[518]&m[1284])|(~m[262]&m[518]&m[1284]))&BiasedRNG[485])|(((m[262]&m[518]&~m[1284]))&~BiasedRNG[485])|((m[262]&m[518]&m[1284]))):InitCond[756];
    m[775] = run?((((m[278]&~m[519]&m[1344])|(~m[278]&m[519]&m[1344]))&BiasedRNG[486])|(((m[278]&m[519]&~m[1344]))&~BiasedRNG[486])|((m[278]&m[519]&m[1344]))):InitCond[757];
    m[776] = run?((((m[294]&~m[520]&m[1409])|(~m[294]&m[520]&m[1409]))&BiasedRNG[487])|(((m[294]&m[520]&~m[1409]))&~BiasedRNG[487])|((m[294]&m[520]&m[1409]))):InitCond[758];
    m[777] = run?((((m[310]&~m[521]&m[1479])|(~m[310]&m[521]&m[1479]))&BiasedRNG[488])|(((m[310]&m[521]&~m[1479]))&~BiasedRNG[488])|((m[310]&m[521]&m[1479]))):InitCond[759];
    m[778] = run?((((m[326]&~m[522]&m[1554])|(~m[326]&m[522]&m[1554]))&BiasedRNG[489])|(((m[326]&m[522]&~m[1554]))&~BiasedRNG[489])|((m[326]&m[522]&m[1554]))):InitCond[760];
    m[779] = run?((((m[342]&~m[523]&m[1624])|(~m[342]&m[523]&m[1624]))&BiasedRNG[490])|(((m[342]&m[523]&~m[1624]))&~BiasedRNG[490])|((m[342]&m[523]&m[1624]))):InitCond[761];
    m[780] = run?((((m[358]&~m[524]&m[1689])|(~m[358]&m[524]&m[1689]))&BiasedRNG[491])|(((m[358]&m[524]&~m[1689]))&~BiasedRNG[491])|((m[358]&m[524]&m[1689]))):InitCond[762];
    m[781] = run?((((m[374]&~m[525]&m[1749])|(~m[374]&m[525]&m[1749]))&BiasedRNG[492])|(((m[374]&m[525]&~m[1749]))&~BiasedRNG[492])|((m[374]&m[525]&m[1749]))):InitCond[763];
    m[782] = run?((((m[390]&~m[526]&m[1804])|(~m[390]&m[526]&m[1804]))&BiasedRNG[493])|(((m[390]&m[526]&~m[1804]))&~BiasedRNG[493])|((m[390]&m[526]&m[1804]))):InitCond[764];
    m[783] = run?((((m[406]&~m[527]&m[1854])|(~m[406]&m[527]&m[1854]))&BiasedRNG[494])|(((m[406]&m[527]&~m[1854]))&~BiasedRNG[494])|((m[406]&m[527]&m[1854]))):InitCond[765];
    m[784] = run?((((m[167]&~m[528]&m[1064])|(~m[167]&m[528]&m[1064]))&BiasedRNG[495])|(((m[167]&m[528]&~m[1064]))&~BiasedRNG[495])|((m[167]&m[528]&m[1064]))):InitCond[766];
    m[785] = run?((((m[183]&~m[529]&m[1099])|(~m[183]&m[529]&m[1099]))&BiasedRNG[496])|(((m[183]&m[529]&~m[1099]))&~BiasedRNG[496])|((m[183]&m[529]&m[1099]))):InitCond[767];
    m[786] = run?((((m[199]&~m[530]&m[1139])|(~m[199]&m[530]&m[1139]))&BiasedRNG[497])|(((m[199]&m[530]&~m[1139]))&~BiasedRNG[497])|((m[199]&m[530]&m[1139]))):InitCond[768];
    m[787] = run?((((m[215]&~m[531]&m[1184])|(~m[215]&m[531]&m[1184]))&BiasedRNG[498])|(((m[215]&m[531]&~m[1184]))&~BiasedRNG[498])|((m[215]&m[531]&m[1184]))):InitCond[769];
    m[788] = run?((((m[231]&~m[532]&m[1234])|(~m[231]&m[532]&m[1234]))&BiasedRNG[499])|(((m[231]&m[532]&~m[1234]))&~BiasedRNG[499])|((m[231]&m[532]&m[1234]))):InitCond[770];
    m[789] = run?((((m[247]&~m[533]&m[1289])|(~m[247]&m[533]&m[1289]))&BiasedRNG[500])|(((m[247]&m[533]&~m[1289]))&~BiasedRNG[500])|((m[247]&m[533]&m[1289]))):InitCond[771];
    m[790] = run?((((m[263]&~m[534]&m[1349])|(~m[263]&m[534]&m[1349]))&BiasedRNG[501])|(((m[263]&m[534]&~m[1349]))&~BiasedRNG[501])|((m[263]&m[534]&m[1349]))):InitCond[772];
    m[791] = run?((((m[279]&~m[535]&m[1414])|(~m[279]&m[535]&m[1414]))&BiasedRNG[502])|(((m[279]&m[535]&~m[1414]))&~BiasedRNG[502])|((m[279]&m[535]&m[1414]))):InitCond[773];
    m[792] = run?((((m[295]&~m[536]&m[1484])|(~m[295]&m[536]&m[1484]))&BiasedRNG[503])|(((m[295]&m[536]&~m[1484]))&~BiasedRNG[503])|((m[295]&m[536]&m[1484]))):InitCond[774];
    m[793] = run?((((m[311]&~m[537]&m[1559])|(~m[311]&m[537]&m[1559]))&BiasedRNG[504])|(((m[311]&m[537]&~m[1559]))&~BiasedRNG[504])|((m[311]&m[537]&m[1559]))):InitCond[775];
    m[794] = run?((((m[327]&~m[538]&m[1629])|(~m[327]&m[538]&m[1629]))&BiasedRNG[505])|(((m[327]&m[538]&~m[1629]))&~BiasedRNG[505])|((m[327]&m[538]&m[1629]))):InitCond[776];
    m[795] = run?((((m[343]&~m[539]&m[1694])|(~m[343]&m[539]&m[1694]))&BiasedRNG[506])|(((m[343]&m[539]&~m[1694]))&~BiasedRNG[506])|((m[343]&m[539]&m[1694]))):InitCond[777];
    m[796] = run?((((m[359]&~m[540]&m[1754])|(~m[359]&m[540]&m[1754]))&BiasedRNG[507])|(((m[359]&m[540]&~m[1754]))&~BiasedRNG[507])|((m[359]&m[540]&m[1754]))):InitCond[778];
    m[797] = run?((((m[375]&~m[541]&m[1809])|(~m[375]&m[541]&m[1809]))&BiasedRNG[508])|(((m[375]&m[541]&~m[1809]))&~BiasedRNG[508])|((m[375]&m[541]&m[1809]))):InitCond[779];
    m[798] = run?((((m[391]&~m[542]&m[1859])|(~m[391]&m[542]&m[1859]))&BiasedRNG[509])|(((m[391]&m[542]&~m[1859]))&~BiasedRNG[509])|((m[391]&m[542]&m[1859]))):InitCond[780];
    m[799] = run?((((m[407]&~m[543]&m[1904])|(~m[407]&m[543]&m[1904]))&BiasedRNG[510])|(((m[407]&m[543]&~m[1904]))&~BiasedRNG[510])|((m[407]&m[543]&m[1904]))):InitCond[781];
    m[800] = run?((((m[168]&~m[544]&m[1104])|(~m[168]&m[544]&m[1104]))&BiasedRNG[511])|(((m[168]&m[544]&~m[1104]))&~BiasedRNG[511])|((m[168]&m[544]&m[1104]))):InitCond[782];
    m[801] = run?((((m[184]&~m[545]&m[1144])|(~m[184]&m[545]&m[1144]))&BiasedRNG[512])|(((m[184]&m[545]&~m[1144]))&~BiasedRNG[512])|((m[184]&m[545]&m[1144]))):InitCond[783];
    m[802] = run?((((m[200]&~m[546]&m[1189])|(~m[200]&m[546]&m[1189]))&BiasedRNG[513])|(((m[200]&m[546]&~m[1189]))&~BiasedRNG[513])|((m[200]&m[546]&m[1189]))):InitCond[784];
    m[803] = run?((((m[216]&~m[547]&m[1239])|(~m[216]&m[547]&m[1239]))&BiasedRNG[514])|(((m[216]&m[547]&~m[1239]))&~BiasedRNG[514])|((m[216]&m[547]&m[1239]))):InitCond[785];
    m[804] = run?((((m[232]&~m[548]&m[1294])|(~m[232]&m[548]&m[1294]))&BiasedRNG[515])|(((m[232]&m[548]&~m[1294]))&~BiasedRNG[515])|((m[232]&m[548]&m[1294]))):InitCond[786];
    m[805] = run?((((m[248]&~m[549]&m[1354])|(~m[248]&m[549]&m[1354]))&BiasedRNG[516])|(((m[248]&m[549]&~m[1354]))&~BiasedRNG[516])|((m[248]&m[549]&m[1354]))):InitCond[787];
    m[806] = run?((((m[264]&~m[550]&m[1419])|(~m[264]&m[550]&m[1419]))&BiasedRNG[517])|(((m[264]&m[550]&~m[1419]))&~BiasedRNG[517])|((m[264]&m[550]&m[1419]))):InitCond[788];
    m[807] = run?((((m[280]&~m[551]&m[1489])|(~m[280]&m[551]&m[1489]))&BiasedRNG[518])|(((m[280]&m[551]&~m[1489]))&~BiasedRNG[518])|((m[280]&m[551]&m[1489]))):InitCond[789];
    m[808] = run?((((m[296]&~m[552]&m[1564])|(~m[296]&m[552]&m[1564]))&BiasedRNG[519])|(((m[296]&m[552]&~m[1564]))&~BiasedRNG[519])|((m[296]&m[552]&m[1564]))):InitCond[790];
    m[809] = run?((((m[312]&~m[553]&m[1634])|(~m[312]&m[553]&m[1634]))&BiasedRNG[520])|(((m[312]&m[553]&~m[1634]))&~BiasedRNG[520])|((m[312]&m[553]&m[1634]))):InitCond[791];
    m[810] = run?((((m[328]&~m[554]&m[1699])|(~m[328]&m[554]&m[1699]))&BiasedRNG[521])|(((m[328]&m[554]&~m[1699]))&~BiasedRNG[521])|((m[328]&m[554]&m[1699]))):InitCond[792];
    m[811] = run?((((m[344]&~m[555]&m[1759])|(~m[344]&m[555]&m[1759]))&BiasedRNG[522])|(((m[344]&m[555]&~m[1759]))&~BiasedRNG[522])|((m[344]&m[555]&m[1759]))):InitCond[793];
    m[812] = run?((((m[360]&~m[556]&m[1814])|(~m[360]&m[556]&m[1814]))&BiasedRNG[523])|(((m[360]&m[556]&~m[1814]))&~BiasedRNG[523])|((m[360]&m[556]&m[1814]))):InitCond[794];
    m[813] = run?((((m[376]&~m[557]&m[1864])|(~m[376]&m[557]&m[1864]))&BiasedRNG[524])|(((m[376]&m[557]&~m[1864]))&~BiasedRNG[524])|((m[376]&m[557]&m[1864]))):InitCond[795];
    m[814] = run?((((m[392]&~m[558]&m[1909])|(~m[392]&m[558]&m[1909]))&BiasedRNG[525])|(((m[392]&m[558]&~m[1909]))&~BiasedRNG[525])|((m[392]&m[558]&m[1909]))):InitCond[796];
    m[815] = run?((((m[408]&~m[559]&m[1949])|(~m[408]&m[559]&m[1949]))&BiasedRNG[526])|(((m[408]&m[559]&~m[1949]))&~BiasedRNG[526])|((m[408]&m[559]&m[1949]))):InitCond[797];
    m[816] = run?((((m[169]&~m[560]&m[1149])|(~m[169]&m[560]&m[1149]))&BiasedRNG[527])|(((m[169]&m[560]&~m[1149]))&~BiasedRNG[527])|((m[169]&m[560]&m[1149]))):InitCond[798];
    m[817] = run?((((m[185]&~m[561]&m[1194])|(~m[185]&m[561]&m[1194]))&BiasedRNG[528])|(((m[185]&m[561]&~m[1194]))&~BiasedRNG[528])|((m[185]&m[561]&m[1194]))):InitCond[799];
    m[818] = run?((((m[201]&~m[562]&m[1244])|(~m[201]&m[562]&m[1244]))&BiasedRNG[529])|(((m[201]&m[562]&~m[1244]))&~BiasedRNG[529])|((m[201]&m[562]&m[1244]))):InitCond[800];
    m[819] = run?((((m[217]&~m[563]&m[1299])|(~m[217]&m[563]&m[1299]))&BiasedRNG[530])|(((m[217]&m[563]&~m[1299]))&~BiasedRNG[530])|((m[217]&m[563]&m[1299]))):InitCond[801];
    m[820] = run?((((m[233]&~m[564]&m[1359])|(~m[233]&m[564]&m[1359]))&BiasedRNG[531])|(((m[233]&m[564]&~m[1359]))&~BiasedRNG[531])|((m[233]&m[564]&m[1359]))):InitCond[802];
    m[821] = run?((((m[249]&~m[565]&m[1424])|(~m[249]&m[565]&m[1424]))&BiasedRNG[532])|(((m[249]&m[565]&~m[1424]))&~BiasedRNG[532])|((m[249]&m[565]&m[1424]))):InitCond[803];
    m[822] = run?((((m[265]&~m[566]&m[1494])|(~m[265]&m[566]&m[1494]))&BiasedRNG[533])|(((m[265]&m[566]&~m[1494]))&~BiasedRNG[533])|((m[265]&m[566]&m[1494]))):InitCond[804];
    m[823] = run?((((m[281]&~m[567]&m[1569])|(~m[281]&m[567]&m[1569]))&BiasedRNG[534])|(((m[281]&m[567]&~m[1569]))&~BiasedRNG[534])|((m[281]&m[567]&m[1569]))):InitCond[805];
    m[824] = run?((((m[297]&~m[568]&m[1639])|(~m[297]&m[568]&m[1639]))&BiasedRNG[535])|(((m[297]&m[568]&~m[1639]))&~BiasedRNG[535])|((m[297]&m[568]&m[1639]))):InitCond[806];
    m[825] = run?((((m[313]&~m[569]&m[1704])|(~m[313]&m[569]&m[1704]))&BiasedRNG[536])|(((m[313]&m[569]&~m[1704]))&~BiasedRNG[536])|((m[313]&m[569]&m[1704]))):InitCond[807];
    m[826] = run?((((m[329]&~m[570]&m[1764])|(~m[329]&m[570]&m[1764]))&BiasedRNG[537])|(((m[329]&m[570]&~m[1764]))&~BiasedRNG[537])|((m[329]&m[570]&m[1764]))):InitCond[808];
    m[827] = run?((((m[345]&~m[571]&m[1819])|(~m[345]&m[571]&m[1819]))&BiasedRNG[538])|(((m[345]&m[571]&~m[1819]))&~BiasedRNG[538])|((m[345]&m[571]&m[1819]))):InitCond[809];
    m[828] = run?((((m[361]&~m[572]&m[1869])|(~m[361]&m[572]&m[1869]))&BiasedRNG[539])|(((m[361]&m[572]&~m[1869]))&~BiasedRNG[539])|((m[361]&m[572]&m[1869]))):InitCond[810];
    m[829] = run?((((m[377]&~m[573]&m[1914])|(~m[377]&m[573]&m[1914]))&BiasedRNG[540])|(((m[377]&m[573]&~m[1914]))&~BiasedRNG[540])|((m[377]&m[573]&m[1914]))):InitCond[811];
    m[830] = run?((((m[393]&~m[574]&m[1954])|(~m[393]&m[574]&m[1954]))&BiasedRNG[541])|(((m[393]&m[574]&~m[1954]))&~BiasedRNG[541])|((m[393]&m[574]&m[1954]))):InitCond[812];
    m[831] = run?((((m[409]&~m[575]&m[1989])|(~m[409]&m[575]&m[1989]))&BiasedRNG[542])|(((m[409]&m[575]&~m[1989]))&~BiasedRNG[542])|((m[409]&m[575]&m[1989]))):InitCond[813];
    m[832] = run?((((m[170]&~m[576]&m[1199])|(~m[170]&m[576]&m[1199]))&BiasedRNG[543])|(((m[170]&m[576]&~m[1199]))&~BiasedRNG[543])|((m[170]&m[576]&m[1199]))):InitCond[814];
    m[833] = run?((((m[186]&~m[577]&m[1249])|(~m[186]&m[577]&m[1249]))&BiasedRNG[544])|(((m[186]&m[577]&~m[1249]))&~BiasedRNG[544])|((m[186]&m[577]&m[1249]))):InitCond[815];
    m[834] = run?((((m[202]&~m[578]&m[1304])|(~m[202]&m[578]&m[1304]))&BiasedRNG[545])|(((m[202]&m[578]&~m[1304]))&~BiasedRNG[545])|((m[202]&m[578]&m[1304]))):InitCond[816];
    m[835] = run?((((m[218]&~m[579]&m[1364])|(~m[218]&m[579]&m[1364]))&BiasedRNG[546])|(((m[218]&m[579]&~m[1364]))&~BiasedRNG[546])|((m[218]&m[579]&m[1364]))):InitCond[817];
    m[836] = run?((((m[234]&~m[580]&m[1429])|(~m[234]&m[580]&m[1429]))&BiasedRNG[547])|(((m[234]&m[580]&~m[1429]))&~BiasedRNG[547])|((m[234]&m[580]&m[1429]))):InitCond[818];
    m[837] = run?((((m[250]&~m[581]&m[1499])|(~m[250]&m[581]&m[1499]))&BiasedRNG[548])|(((m[250]&m[581]&~m[1499]))&~BiasedRNG[548])|((m[250]&m[581]&m[1499]))):InitCond[819];
    m[838] = run?((((m[266]&~m[582]&m[1574])|(~m[266]&m[582]&m[1574]))&BiasedRNG[549])|(((m[266]&m[582]&~m[1574]))&~BiasedRNG[549])|((m[266]&m[582]&m[1574]))):InitCond[820];
    m[839] = run?((((m[282]&~m[583]&m[1644])|(~m[282]&m[583]&m[1644]))&BiasedRNG[550])|(((m[282]&m[583]&~m[1644]))&~BiasedRNG[550])|((m[282]&m[583]&m[1644]))):InitCond[821];
    m[840] = run?((((m[298]&~m[584]&m[1709])|(~m[298]&m[584]&m[1709]))&BiasedRNG[551])|(((m[298]&m[584]&~m[1709]))&~BiasedRNG[551])|((m[298]&m[584]&m[1709]))):InitCond[822];
    m[841] = run?((((m[314]&~m[585]&m[1769])|(~m[314]&m[585]&m[1769]))&BiasedRNG[552])|(((m[314]&m[585]&~m[1769]))&~BiasedRNG[552])|((m[314]&m[585]&m[1769]))):InitCond[823];
    m[842] = run?((((m[330]&~m[586]&m[1824])|(~m[330]&m[586]&m[1824]))&BiasedRNG[553])|(((m[330]&m[586]&~m[1824]))&~BiasedRNG[553])|((m[330]&m[586]&m[1824]))):InitCond[824];
    m[843] = run?((((m[346]&~m[587]&m[1874])|(~m[346]&m[587]&m[1874]))&BiasedRNG[554])|(((m[346]&m[587]&~m[1874]))&~BiasedRNG[554])|((m[346]&m[587]&m[1874]))):InitCond[825];
    m[844] = run?((((m[362]&~m[588]&m[1919])|(~m[362]&m[588]&m[1919]))&BiasedRNG[555])|(((m[362]&m[588]&~m[1919]))&~BiasedRNG[555])|((m[362]&m[588]&m[1919]))):InitCond[826];
    m[845] = run?((((m[378]&~m[589]&m[1959])|(~m[378]&m[589]&m[1959]))&BiasedRNG[556])|(((m[378]&m[589]&~m[1959]))&~BiasedRNG[556])|((m[378]&m[589]&m[1959]))):InitCond[827];
    m[846] = run?((((m[394]&~m[590]&m[1994])|(~m[394]&m[590]&m[1994]))&BiasedRNG[557])|(((m[394]&m[590]&~m[1994]))&~BiasedRNG[557])|((m[394]&m[590]&m[1994]))):InitCond[828];
    m[847] = run?((((m[410]&~m[591]&m[2024])|(~m[410]&m[591]&m[2024]))&BiasedRNG[558])|(((m[410]&m[591]&~m[2024]))&~BiasedRNG[558])|((m[410]&m[591]&m[2024]))):InitCond[829];
    m[848] = run?((((m[171]&~m[592]&m[1254])|(~m[171]&m[592]&m[1254]))&BiasedRNG[559])|(((m[171]&m[592]&~m[1254]))&~BiasedRNG[559])|((m[171]&m[592]&m[1254]))):InitCond[830];
    m[849] = run?((((m[187]&~m[593]&m[1309])|(~m[187]&m[593]&m[1309]))&BiasedRNG[560])|(((m[187]&m[593]&~m[1309]))&~BiasedRNG[560])|((m[187]&m[593]&m[1309]))):InitCond[831];
    m[850] = run?((((m[203]&~m[594]&m[1369])|(~m[203]&m[594]&m[1369]))&BiasedRNG[561])|(((m[203]&m[594]&~m[1369]))&~BiasedRNG[561])|((m[203]&m[594]&m[1369]))):InitCond[832];
    m[851] = run?((((m[219]&~m[595]&m[1434])|(~m[219]&m[595]&m[1434]))&BiasedRNG[562])|(((m[219]&m[595]&~m[1434]))&~BiasedRNG[562])|((m[219]&m[595]&m[1434]))):InitCond[833];
    m[852] = run?((((m[235]&~m[596]&m[1504])|(~m[235]&m[596]&m[1504]))&BiasedRNG[563])|(((m[235]&m[596]&~m[1504]))&~BiasedRNG[563])|((m[235]&m[596]&m[1504]))):InitCond[834];
    m[853] = run?((((m[251]&~m[597]&m[1579])|(~m[251]&m[597]&m[1579]))&BiasedRNG[564])|(((m[251]&m[597]&~m[1579]))&~BiasedRNG[564])|((m[251]&m[597]&m[1579]))):InitCond[835];
    m[854] = run?((((m[267]&~m[598]&m[1649])|(~m[267]&m[598]&m[1649]))&BiasedRNG[565])|(((m[267]&m[598]&~m[1649]))&~BiasedRNG[565])|((m[267]&m[598]&m[1649]))):InitCond[836];
    m[855] = run?((((m[283]&~m[599]&m[1714])|(~m[283]&m[599]&m[1714]))&BiasedRNG[566])|(((m[283]&m[599]&~m[1714]))&~BiasedRNG[566])|((m[283]&m[599]&m[1714]))):InitCond[837];
    m[856] = run?((((m[299]&~m[600]&m[1774])|(~m[299]&m[600]&m[1774]))&BiasedRNG[567])|(((m[299]&m[600]&~m[1774]))&~BiasedRNG[567])|((m[299]&m[600]&m[1774]))):InitCond[838];
    m[857] = run?((((m[315]&~m[601]&m[1829])|(~m[315]&m[601]&m[1829]))&BiasedRNG[568])|(((m[315]&m[601]&~m[1829]))&~BiasedRNG[568])|((m[315]&m[601]&m[1829]))):InitCond[839];
    m[858] = run?((((m[331]&~m[602]&m[1879])|(~m[331]&m[602]&m[1879]))&BiasedRNG[569])|(((m[331]&m[602]&~m[1879]))&~BiasedRNG[569])|((m[331]&m[602]&m[1879]))):InitCond[840];
    m[859] = run?((((m[347]&~m[603]&m[1924])|(~m[347]&m[603]&m[1924]))&BiasedRNG[570])|(((m[347]&m[603]&~m[1924]))&~BiasedRNG[570])|((m[347]&m[603]&m[1924]))):InitCond[841];
    m[860] = run?((((m[363]&~m[604]&m[1964])|(~m[363]&m[604]&m[1964]))&BiasedRNG[571])|(((m[363]&m[604]&~m[1964]))&~BiasedRNG[571])|((m[363]&m[604]&m[1964]))):InitCond[842];
    m[861] = run?((((m[379]&~m[605]&m[1999])|(~m[379]&m[605]&m[1999]))&BiasedRNG[572])|(((m[379]&m[605]&~m[1999]))&~BiasedRNG[572])|((m[379]&m[605]&m[1999]))):InitCond[843];
    m[862] = run?((((m[395]&~m[606]&m[2029])|(~m[395]&m[606]&m[2029]))&BiasedRNG[573])|(((m[395]&m[606]&~m[2029]))&~BiasedRNG[573])|((m[395]&m[606]&m[2029]))):InitCond[844];
    m[863] = run?((((m[411]&~m[607]&m[2054])|(~m[411]&m[607]&m[2054]))&BiasedRNG[574])|(((m[411]&m[607]&~m[2054]))&~BiasedRNG[574])|((m[411]&m[607]&m[2054]))):InitCond[845];
    m[864] = run?((((m[172]&~m[608]&m[1314])|(~m[172]&m[608]&m[1314]))&BiasedRNG[575])|(((m[172]&m[608]&~m[1314]))&~BiasedRNG[575])|((m[172]&m[608]&m[1314]))):InitCond[846];
    m[865] = run?((((m[188]&~m[609]&m[1374])|(~m[188]&m[609]&m[1374]))&BiasedRNG[576])|(((m[188]&m[609]&~m[1374]))&~BiasedRNG[576])|((m[188]&m[609]&m[1374]))):InitCond[847];
    m[866] = run?((((m[204]&~m[610]&m[1439])|(~m[204]&m[610]&m[1439]))&BiasedRNG[577])|(((m[204]&m[610]&~m[1439]))&~BiasedRNG[577])|((m[204]&m[610]&m[1439]))):InitCond[848];
    m[867] = run?((((m[220]&~m[611]&m[1509])|(~m[220]&m[611]&m[1509]))&BiasedRNG[578])|(((m[220]&m[611]&~m[1509]))&~BiasedRNG[578])|((m[220]&m[611]&m[1509]))):InitCond[849];
    m[868] = run?((((m[236]&~m[612]&m[1584])|(~m[236]&m[612]&m[1584]))&BiasedRNG[579])|(((m[236]&m[612]&~m[1584]))&~BiasedRNG[579])|((m[236]&m[612]&m[1584]))):InitCond[850];
    m[869] = run?((((m[252]&~m[613]&m[1654])|(~m[252]&m[613]&m[1654]))&BiasedRNG[580])|(((m[252]&m[613]&~m[1654]))&~BiasedRNG[580])|((m[252]&m[613]&m[1654]))):InitCond[851];
    m[870] = run?((((m[268]&~m[614]&m[1719])|(~m[268]&m[614]&m[1719]))&BiasedRNG[581])|(((m[268]&m[614]&~m[1719]))&~BiasedRNG[581])|((m[268]&m[614]&m[1719]))):InitCond[852];
    m[871] = run?((((m[284]&~m[615]&m[1779])|(~m[284]&m[615]&m[1779]))&BiasedRNG[582])|(((m[284]&m[615]&~m[1779]))&~BiasedRNG[582])|((m[284]&m[615]&m[1779]))):InitCond[853];
    m[872] = run?((((m[300]&~m[616]&m[1834])|(~m[300]&m[616]&m[1834]))&BiasedRNG[583])|(((m[300]&m[616]&~m[1834]))&~BiasedRNG[583])|((m[300]&m[616]&m[1834]))):InitCond[854];
    m[873] = run?((((m[316]&~m[617]&m[1884])|(~m[316]&m[617]&m[1884]))&BiasedRNG[584])|(((m[316]&m[617]&~m[1884]))&~BiasedRNG[584])|((m[316]&m[617]&m[1884]))):InitCond[855];
    m[874] = run?((((m[332]&~m[618]&m[1929])|(~m[332]&m[618]&m[1929]))&BiasedRNG[585])|(((m[332]&m[618]&~m[1929]))&~BiasedRNG[585])|((m[332]&m[618]&m[1929]))):InitCond[856];
    m[875] = run?((((m[348]&~m[619]&m[1969])|(~m[348]&m[619]&m[1969]))&BiasedRNG[586])|(((m[348]&m[619]&~m[1969]))&~BiasedRNG[586])|((m[348]&m[619]&m[1969]))):InitCond[857];
    m[876] = run?((((m[364]&~m[620]&m[2004])|(~m[364]&m[620]&m[2004]))&BiasedRNG[587])|(((m[364]&m[620]&~m[2004]))&~BiasedRNG[587])|((m[364]&m[620]&m[2004]))):InitCond[858];
    m[877] = run?((((m[380]&~m[621]&m[2034])|(~m[380]&m[621]&m[2034]))&BiasedRNG[588])|(((m[380]&m[621]&~m[2034]))&~BiasedRNG[588])|((m[380]&m[621]&m[2034]))):InitCond[859];
    m[878] = run?((((m[396]&~m[622]&m[2059])|(~m[396]&m[622]&m[2059]))&BiasedRNG[589])|(((m[396]&m[622]&~m[2059]))&~BiasedRNG[589])|((m[396]&m[622]&m[2059]))):InitCond[860];
    m[879] = run?((((m[412]&~m[623]&m[2079])|(~m[412]&m[623]&m[2079]))&BiasedRNG[590])|(((m[412]&m[623]&~m[2079]))&~BiasedRNG[590])|((m[412]&m[623]&m[2079]))):InitCond[861];
    m[880] = run?((((m[173]&~m[624]&m[1379])|(~m[173]&m[624]&m[1379]))&BiasedRNG[591])|(((m[173]&m[624]&~m[1379]))&~BiasedRNG[591])|((m[173]&m[624]&m[1379]))):InitCond[862];
    m[881] = run?((((m[189]&~m[625]&m[1444])|(~m[189]&m[625]&m[1444]))&BiasedRNG[592])|(((m[189]&m[625]&~m[1444]))&~BiasedRNG[592])|((m[189]&m[625]&m[1444]))):InitCond[863];
    m[882] = run?((((m[205]&~m[626]&m[1514])|(~m[205]&m[626]&m[1514]))&BiasedRNG[593])|(((m[205]&m[626]&~m[1514]))&~BiasedRNG[593])|((m[205]&m[626]&m[1514]))):InitCond[864];
    m[883] = run?((((m[221]&~m[627]&m[1589])|(~m[221]&m[627]&m[1589]))&BiasedRNG[594])|(((m[221]&m[627]&~m[1589]))&~BiasedRNG[594])|((m[221]&m[627]&m[1589]))):InitCond[865];
    m[884] = run?((((m[237]&~m[628]&m[1659])|(~m[237]&m[628]&m[1659]))&BiasedRNG[595])|(((m[237]&m[628]&~m[1659]))&~BiasedRNG[595])|((m[237]&m[628]&m[1659]))):InitCond[866];
    m[885] = run?((((m[253]&~m[629]&m[1724])|(~m[253]&m[629]&m[1724]))&BiasedRNG[596])|(((m[253]&m[629]&~m[1724]))&~BiasedRNG[596])|((m[253]&m[629]&m[1724]))):InitCond[867];
    m[886] = run?((((m[269]&~m[630]&m[1784])|(~m[269]&m[630]&m[1784]))&BiasedRNG[597])|(((m[269]&m[630]&~m[1784]))&~BiasedRNG[597])|((m[269]&m[630]&m[1784]))):InitCond[868];
    m[887] = run?((((m[285]&~m[631]&m[1839])|(~m[285]&m[631]&m[1839]))&BiasedRNG[598])|(((m[285]&m[631]&~m[1839]))&~BiasedRNG[598])|((m[285]&m[631]&m[1839]))):InitCond[869];
    m[888] = run?((((m[301]&~m[632]&m[1889])|(~m[301]&m[632]&m[1889]))&BiasedRNG[599])|(((m[301]&m[632]&~m[1889]))&~BiasedRNG[599])|((m[301]&m[632]&m[1889]))):InitCond[870];
    m[889] = run?((((m[317]&~m[633]&m[1934])|(~m[317]&m[633]&m[1934]))&BiasedRNG[600])|(((m[317]&m[633]&~m[1934]))&~BiasedRNG[600])|((m[317]&m[633]&m[1934]))):InitCond[871];
    m[890] = run?((((m[333]&~m[634]&m[1974])|(~m[333]&m[634]&m[1974]))&BiasedRNG[601])|(((m[333]&m[634]&~m[1974]))&~BiasedRNG[601])|((m[333]&m[634]&m[1974]))):InitCond[872];
    m[891] = run?((((m[349]&~m[635]&m[2009])|(~m[349]&m[635]&m[2009]))&BiasedRNG[602])|(((m[349]&m[635]&~m[2009]))&~BiasedRNG[602])|((m[349]&m[635]&m[2009]))):InitCond[873];
    m[892] = run?((((m[365]&~m[636]&m[2039])|(~m[365]&m[636]&m[2039]))&BiasedRNG[603])|(((m[365]&m[636]&~m[2039]))&~BiasedRNG[603])|((m[365]&m[636]&m[2039]))):InitCond[874];
    m[893] = run?((((m[381]&~m[637]&m[2064])|(~m[381]&m[637]&m[2064]))&BiasedRNG[604])|(((m[381]&m[637]&~m[2064]))&~BiasedRNG[604])|((m[381]&m[637]&m[2064]))):InitCond[875];
    m[894] = run?((((m[397]&~m[638]&m[2084])|(~m[397]&m[638]&m[2084]))&BiasedRNG[605])|(((m[397]&m[638]&~m[2084]))&~BiasedRNG[605])|((m[397]&m[638]&m[2084]))):InitCond[876];
    m[895] = run?((((m[413]&~m[639]&m[2099])|(~m[413]&m[639]&m[2099]))&BiasedRNG[606])|(((m[413]&m[639]&~m[2099]))&~BiasedRNG[606])|((m[413]&m[639]&m[2099]))):InitCond[877];
    m[896] = run?((((m[174]&~m[640]&m[1449])|(~m[174]&m[640]&m[1449]))&BiasedRNG[607])|(((m[174]&m[640]&~m[1449]))&~BiasedRNG[607])|((m[174]&m[640]&m[1449]))):InitCond[878];
    m[897] = run?((((m[190]&~m[641]&m[1519])|(~m[190]&m[641]&m[1519]))&BiasedRNG[608])|(((m[190]&m[641]&~m[1519]))&~BiasedRNG[608])|((m[190]&m[641]&m[1519]))):InitCond[879];
    m[898] = run?((((m[206]&~m[642]&m[1594])|(~m[206]&m[642]&m[1594]))&BiasedRNG[609])|(((m[206]&m[642]&~m[1594]))&~BiasedRNG[609])|((m[206]&m[642]&m[1594]))):InitCond[880];
    m[899] = run?((((m[222]&~m[643]&m[1664])|(~m[222]&m[643]&m[1664]))&BiasedRNG[610])|(((m[222]&m[643]&~m[1664]))&~BiasedRNG[610])|((m[222]&m[643]&m[1664]))):InitCond[881];
    m[900] = run?((((m[238]&~m[644]&m[1729])|(~m[238]&m[644]&m[1729]))&BiasedRNG[611])|(((m[238]&m[644]&~m[1729]))&~BiasedRNG[611])|((m[238]&m[644]&m[1729]))):InitCond[882];
    m[901] = run?((((m[254]&~m[645]&m[1789])|(~m[254]&m[645]&m[1789]))&BiasedRNG[612])|(((m[254]&m[645]&~m[1789]))&~BiasedRNG[612])|((m[254]&m[645]&m[1789]))):InitCond[883];
    m[902] = run?((((m[270]&~m[646]&m[1844])|(~m[270]&m[646]&m[1844]))&BiasedRNG[613])|(((m[270]&m[646]&~m[1844]))&~BiasedRNG[613])|((m[270]&m[646]&m[1844]))):InitCond[884];
    m[903] = run?((((m[286]&~m[647]&m[1894])|(~m[286]&m[647]&m[1894]))&BiasedRNG[614])|(((m[286]&m[647]&~m[1894]))&~BiasedRNG[614])|((m[286]&m[647]&m[1894]))):InitCond[885];
    m[904] = run?((((m[302]&~m[648]&m[1939])|(~m[302]&m[648]&m[1939]))&BiasedRNG[615])|(((m[302]&m[648]&~m[1939]))&~BiasedRNG[615])|((m[302]&m[648]&m[1939]))):InitCond[886];
    m[905] = run?((((m[318]&~m[649]&m[1979])|(~m[318]&m[649]&m[1979]))&BiasedRNG[616])|(((m[318]&m[649]&~m[1979]))&~BiasedRNG[616])|((m[318]&m[649]&m[1979]))):InitCond[887];
    m[906] = run?((((m[334]&~m[650]&m[2014])|(~m[334]&m[650]&m[2014]))&BiasedRNG[617])|(((m[334]&m[650]&~m[2014]))&~BiasedRNG[617])|((m[334]&m[650]&m[2014]))):InitCond[888];
    m[907] = run?((((m[350]&~m[651]&m[2044])|(~m[350]&m[651]&m[2044]))&BiasedRNG[618])|(((m[350]&m[651]&~m[2044]))&~BiasedRNG[618])|((m[350]&m[651]&m[2044]))):InitCond[889];
    m[908] = run?((((m[366]&~m[652]&m[2069])|(~m[366]&m[652]&m[2069]))&BiasedRNG[619])|(((m[366]&m[652]&~m[2069]))&~BiasedRNG[619])|((m[366]&m[652]&m[2069]))):InitCond[890];
    m[909] = run?((((m[382]&~m[653]&m[2089])|(~m[382]&m[653]&m[2089]))&BiasedRNG[620])|(((m[382]&m[653]&~m[2089]))&~BiasedRNG[620])|((m[382]&m[653]&m[2089]))):InitCond[891];
    m[910] = run?((((m[398]&~m[654]&m[2104])|(~m[398]&m[654]&m[2104]))&BiasedRNG[621])|(((m[398]&m[654]&~m[2104]))&~BiasedRNG[621])|((m[398]&m[654]&m[2104]))):InitCond[892];
    m[911] = run?((((m[414]&~m[655]&m[2114])|(~m[414]&m[655]&m[2114]))&BiasedRNG[622])|(((m[414]&m[655]&~m[2114]))&~BiasedRNG[622])|((m[414]&m[655]&m[2114]))):InitCond[893];
    m[912] = run?((((m[175]&~m[656]&m[1524])|(~m[175]&m[656]&m[1524]))&BiasedRNG[623])|(((m[175]&m[656]&~m[1524]))&~BiasedRNG[623])|((m[175]&m[656]&m[1524]))):InitCond[894];
    m[913] = run?((((m[191]&~m[657]&m[1599])|(~m[191]&m[657]&m[1599]))&BiasedRNG[624])|(((m[191]&m[657]&~m[1599]))&~BiasedRNG[624])|((m[191]&m[657]&m[1599]))):InitCond[895];
    m[914] = run?((((m[207]&~m[658]&m[1669])|(~m[207]&m[658]&m[1669]))&BiasedRNG[625])|(((m[207]&m[658]&~m[1669]))&~BiasedRNG[625])|((m[207]&m[658]&m[1669]))):InitCond[896];
    m[915] = run?((((m[223]&~m[659]&m[1734])|(~m[223]&m[659]&m[1734]))&BiasedRNG[626])|(((m[223]&m[659]&~m[1734]))&~BiasedRNG[626])|((m[223]&m[659]&m[1734]))):InitCond[897];
    m[916] = run?((((m[239]&~m[660]&m[1794])|(~m[239]&m[660]&m[1794]))&BiasedRNG[627])|(((m[239]&m[660]&~m[1794]))&~BiasedRNG[627])|((m[239]&m[660]&m[1794]))):InitCond[898];
    m[917] = run?((((m[255]&~m[661]&m[1849])|(~m[255]&m[661]&m[1849]))&BiasedRNG[628])|(((m[255]&m[661]&~m[1849]))&~BiasedRNG[628])|((m[255]&m[661]&m[1849]))):InitCond[899];
    m[918] = run?((((m[271]&~m[662]&m[1899])|(~m[271]&m[662]&m[1899]))&BiasedRNG[629])|(((m[271]&m[662]&~m[1899]))&~BiasedRNG[629])|((m[271]&m[662]&m[1899]))):InitCond[900];
    m[919] = run?((((m[287]&~m[663]&m[1944])|(~m[287]&m[663]&m[1944]))&BiasedRNG[630])|(((m[287]&m[663]&~m[1944]))&~BiasedRNG[630])|((m[287]&m[663]&m[1944]))):InitCond[901];
    m[920] = run?((((m[303]&~m[664]&m[1984])|(~m[303]&m[664]&m[1984]))&BiasedRNG[631])|(((m[303]&m[664]&~m[1984]))&~BiasedRNG[631])|((m[303]&m[664]&m[1984]))):InitCond[902];
    m[921] = run?((((m[319]&~m[665]&m[2019])|(~m[319]&m[665]&m[2019]))&BiasedRNG[632])|(((m[319]&m[665]&~m[2019]))&~BiasedRNG[632])|((m[319]&m[665]&m[2019]))):InitCond[903];
    m[922] = run?((((m[335]&~m[666]&m[2049])|(~m[335]&m[666]&m[2049]))&BiasedRNG[633])|(((m[335]&m[666]&~m[2049]))&~BiasedRNG[633])|((m[335]&m[666]&m[2049]))):InitCond[904];
    m[923] = run?((((m[351]&~m[667]&m[2074])|(~m[351]&m[667]&m[2074]))&BiasedRNG[634])|(((m[351]&m[667]&~m[2074]))&~BiasedRNG[634])|((m[351]&m[667]&m[2074]))):InitCond[905];
    m[924] = run?((((m[367]&~m[668]&m[2094])|(~m[367]&m[668]&m[2094]))&BiasedRNG[635])|(((m[367]&m[668]&~m[2094]))&~BiasedRNG[635])|((m[367]&m[668]&m[2094]))):InitCond[906];
    m[925] = run?((((m[383]&~m[669]&m[2109])|(~m[383]&m[669]&m[2109]))&BiasedRNG[636])|(((m[383]&m[669]&~m[2109]))&~BiasedRNG[636])|((m[383]&m[669]&m[2109]))):InitCond[907];
    m[926] = run?((((m[399]&~m[670]&m[2119])|(~m[399]&m[670]&m[2119]))&BiasedRNG[637])|(((m[399]&m[670]&~m[2119]))&~BiasedRNG[637])|((m[399]&m[670]&m[2119]))):InitCond[908];
    m[927] = run?((((m[415]&~m[671]&m[2124])|(~m[415]&m[671]&m[2124]))&BiasedRNG[638])|(((m[415]&m[671]&~m[2124]))&~BiasedRNG[638])|((m[415]&m[671]&m[2124]))):InitCond[909];
    m[935] = run?((((m[932]&~m[933]&~m[934]&~m[936]&~m[937])|(~m[932]&~m[933]&~m[934]&m[936]&~m[937])|(m[932]&m[933]&~m[934]&m[936]&~m[937])|(m[932]&~m[933]&m[934]&m[936]&~m[937])|(~m[932]&m[933]&~m[934]&~m[936]&m[937])|(~m[932]&~m[933]&m[934]&~m[936]&m[937])|(m[932]&m[933]&m[934]&~m[936]&m[937])|(~m[932]&m[933]&m[934]&m[936]&m[937]))&UnbiasedRNG[271])|((m[932]&~m[933]&~m[934]&m[936]&~m[937])|(~m[932]&~m[933]&~m[934]&~m[936]&m[937])|(m[932]&~m[933]&~m[934]&~m[936]&m[937])|(m[932]&m[933]&~m[934]&~m[936]&m[937])|(m[932]&~m[933]&m[934]&~m[936]&m[937])|(~m[932]&~m[933]&~m[934]&m[936]&m[937])|(m[932]&~m[933]&~m[934]&m[936]&m[937])|(~m[932]&m[933]&~m[934]&m[936]&m[937])|(m[932]&m[933]&~m[934]&m[936]&m[937])|(~m[932]&~m[933]&m[934]&m[936]&m[937])|(m[932]&~m[933]&m[934]&m[936]&m[937])|(m[932]&m[933]&m[934]&m[936]&m[937]))):InitCond[910];
    m[945] = run?((((m[937]&~m[943]&~m[944]&~m[946]&~m[947])|(~m[937]&~m[943]&~m[944]&m[946]&~m[947])|(m[937]&m[943]&~m[944]&m[946]&~m[947])|(m[937]&~m[943]&m[944]&m[946]&~m[947])|(~m[937]&m[943]&~m[944]&~m[946]&m[947])|(~m[937]&~m[943]&m[944]&~m[946]&m[947])|(m[937]&m[943]&m[944]&~m[946]&m[947])|(~m[937]&m[943]&m[944]&m[946]&m[947]))&UnbiasedRNG[272])|((m[937]&~m[943]&~m[944]&m[946]&~m[947])|(~m[937]&~m[943]&~m[944]&~m[946]&m[947])|(m[937]&~m[943]&~m[944]&~m[946]&m[947])|(m[937]&m[943]&~m[944]&~m[946]&m[947])|(m[937]&~m[943]&m[944]&~m[946]&m[947])|(~m[937]&~m[943]&~m[944]&m[946]&m[947])|(m[937]&~m[943]&~m[944]&m[946]&m[947])|(~m[937]&m[943]&~m[944]&m[946]&m[947])|(m[937]&m[943]&~m[944]&m[946]&m[947])|(~m[937]&~m[943]&m[944]&m[946]&m[947])|(m[937]&~m[943]&m[944]&m[946]&m[947])|(m[937]&m[943]&m[944]&m[946]&m[947]))):InitCond[911];
    m[950] = run?((((m[942]&~m[948]&~m[949]&~m[951]&~m[952])|(~m[942]&~m[948]&~m[949]&m[951]&~m[952])|(m[942]&m[948]&~m[949]&m[951]&~m[952])|(m[942]&~m[948]&m[949]&m[951]&~m[952])|(~m[942]&m[948]&~m[949]&~m[951]&m[952])|(~m[942]&~m[948]&m[949]&~m[951]&m[952])|(m[942]&m[948]&m[949]&~m[951]&m[952])|(~m[942]&m[948]&m[949]&m[951]&m[952]))&UnbiasedRNG[273])|((m[942]&~m[948]&~m[949]&m[951]&~m[952])|(~m[942]&~m[948]&~m[949]&~m[951]&m[952])|(m[942]&~m[948]&~m[949]&~m[951]&m[952])|(m[942]&m[948]&~m[949]&~m[951]&m[952])|(m[942]&~m[948]&m[949]&~m[951]&m[952])|(~m[942]&~m[948]&~m[949]&m[951]&m[952])|(m[942]&~m[948]&~m[949]&m[951]&m[952])|(~m[942]&m[948]&~m[949]&m[951]&m[952])|(m[942]&m[948]&~m[949]&m[951]&m[952])|(~m[942]&~m[948]&m[949]&m[951]&m[952])|(m[942]&~m[948]&m[949]&m[951]&m[952])|(m[942]&m[948]&m[949]&m[951]&m[952]))):InitCond[912];
    m[960] = run?((((m[947]&~m[958]&~m[959]&~m[961]&~m[962])|(~m[947]&~m[958]&~m[959]&m[961]&~m[962])|(m[947]&m[958]&~m[959]&m[961]&~m[962])|(m[947]&~m[958]&m[959]&m[961]&~m[962])|(~m[947]&m[958]&~m[959]&~m[961]&m[962])|(~m[947]&~m[958]&m[959]&~m[961]&m[962])|(m[947]&m[958]&m[959]&~m[961]&m[962])|(~m[947]&m[958]&m[959]&m[961]&m[962]))&UnbiasedRNG[274])|((m[947]&~m[958]&~m[959]&m[961]&~m[962])|(~m[947]&~m[958]&~m[959]&~m[961]&m[962])|(m[947]&~m[958]&~m[959]&~m[961]&m[962])|(m[947]&m[958]&~m[959]&~m[961]&m[962])|(m[947]&~m[958]&m[959]&~m[961]&m[962])|(~m[947]&~m[958]&~m[959]&m[961]&m[962])|(m[947]&~m[958]&~m[959]&m[961]&m[962])|(~m[947]&m[958]&~m[959]&m[961]&m[962])|(m[947]&m[958]&~m[959]&m[961]&m[962])|(~m[947]&~m[958]&m[959]&m[961]&m[962])|(m[947]&~m[958]&m[959]&m[961]&m[962])|(m[947]&m[958]&m[959]&m[961]&m[962]))):InitCond[913];
    m[965] = run?((((m[952]&~m[963]&~m[964]&~m[966]&~m[967])|(~m[952]&~m[963]&~m[964]&m[966]&~m[967])|(m[952]&m[963]&~m[964]&m[966]&~m[967])|(m[952]&~m[963]&m[964]&m[966]&~m[967])|(~m[952]&m[963]&~m[964]&~m[966]&m[967])|(~m[952]&~m[963]&m[964]&~m[966]&m[967])|(m[952]&m[963]&m[964]&~m[966]&m[967])|(~m[952]&m[963]&m[964]&m[966]&m[967]))&UnbiasedRNG[275])|((m[952]&~m[963]&~m[964]&m[966]&~m[967])|(~m[952]&~m[963]&~m[964]&~m[966]&m[967])|(m[952]&~m[963]&~m[964]&~m[966]&m[967])|(m[952]&m[963]&~m[964]&~m[966]&m[967])|(m[952]&~m[963]&m[964]&~m[966]&m[967])|(~m[952]&~m[963]&~m[964]&m[966]&m[967])|(m[952]&~m[963]&~m[964]&m[966]&m[967])|(~m[952]&m[963]&~m[964]&m[966]&m[967])|(m[952]&m[963]&~m[964]&m[966]&m[967])|(~m[952]&~m[963]&m[964]&m[966]&m[967])|(m[952]&~m[963]&m[964]&m[966]&m[967])|(m[952]&m[963]&m[964]&m[966]&m[967]))):InitCond[914];
    m[970] = run?((((m[957]&~m[968]&~m[969]&~m[971]&~m[972])|(~m[957]&~m[968]&~m[969]&m[971]&~m[972])|(m[957]&m[968]&~m[969]&m[971]&~m[972])|(m[957]&~m[968]&m[969]&m[971]&~m[972])|(~m[957]&m[968]&~m[969]&~m[971]&m[972])|(~m[957]&~m[968]&m[969]&~m[971]&m[972])|(m[957]&m[968]&m[969]&~m[971]&m[972])|(~m[957]&m[968]&m[969]&m[971]&m[972]))&UnbiasedRNG[276])|((m[957]&~m[968]&~m[969]&m[971]&~m[972])|(~m[957]&~m[968]&~m[969]&~m[971]&m[972])|(m[957]&~m[968]&~m[969]&~m[971]&m[972])|(m[957]&m[968]&~m[969]&~m[971]&m[972])|(m[957]&~m[968]&m[969]&~m[971]&m[972])|(~m[957]&~m[968]&~m[969]&m[971]&m[972])|(m[957]&~m[968]&~m[969]&m[971]&m[972])|(~m[957]&m[968]&~m[969]&m[971]&m[972])|(m[957]&m[968]&~m[969]&m[971]&m[972])|(~m[957]&~m[968]&m[969]&m[971]&m[972])|(m[957]&~m[968]&m[969]&m[971]&m[972])|(m[957]&m[968]&m[969]&m[971]&m[972]))):InitCond[915];
    m[980] = run?((((m[962]&~m[978]&~m[979]&~m[981]&~m[982])|(~m[962]&~m[978]&~m[979]&m[981]&~m[982])|(m[962]&m[978]&~m[979]&m[981]&~m[982])|(m[962]&~m[978]&m[979]&m[981]&~m[982])|(~m[962]&m[978]&~m[979]&~m[981]&m[982])|(~m[962]&~m[978]&m[979]&~m[981]&m[982])|(m[962]&m[978]&m[979]&~m[981]&m[982])|(~m[962]&m[978]&m[979]&m[981]&m[982]))&UnbiasedRNG[277])|((m[962]&~m[978]&~m[979]&m[981]&~m[982])|(~m[962]&~m[978]&~m[979]&~m[981]&m[982])|(m[962]&~m[978]&~m[979]&~m[981]&m[982])|(m[962]&m[978]&~m[979]&~m[981]&m[982])|(m[962]&~m[978]&m[979]&~m[981]&m[982])|(~m[962]&~m[978]&~m[979]&m[981]&m[982])|(m[962]&~m[978]&~m[979]&m[981]&m[982])|(~m[962]&m[978]&~m[979]&m[981]&m[982])|(m[962]&m[978]&~m[979]&m[981]&m[982])|(~m[962]&~m[978]&m[979]&m[981]&m[982])|(m[962]&~m[978]&m[979]&m[981]&m[982])|(m[962]&m[978]&m[979]&m[981]&m[982]))):InitCond[916];
    m[985] = run?((((m[967]&~m[983]&~m[984]&~m[986]&~m[987])|(~m[967]&~m[983]&~m[984]&m[986]&~m[987])|(m[967]&m[983]&~m[984]&m[986]&~m[987])|(m[967]&~m[983]&m[984]&m[986]&~m[987])|(~m[967]&m[983]&~m[984]&~m[986]&m[987])|(~m[967]&~m[983]&m[984]&~m[986]&m[987])|(m[967]&m[983]&m[984]&~m[986]&m[987])|(~m[967]&m[983]&m[984]&m[986]&m[987]))&UnbiasedRNG[278])|((m[967]&~m[983]&~m[984]&m[986]&~m[987])|(~m[967]&~m[983]&~m[984]&~m[986]&m[987])|(m[967]&~m[983]&~m[984]&~m[986]&m[987])|(m[967]&m[983]&~m[984]&~m[986]&m[987])|(m[967]&~m[983]&m[984]&~m[986]&m[987])|(~m[967]&~m[983]&~m[984]&m[986]&m[987])|(m[967]&~m[983]&~m[984]&m[986]&m[987])|(~m[967]&m[983]&~m[984]&m[986]&m[987])|(m[967]&m[983]&~m[984]&m[986]&m[987])|(~m[967]&~m[983]&m[984]&m[986]&m[987])|(m[967]&~m[983]&m[984]&m[986]&m[987])|(m[967]&m[983]&m[984]&m[986]&m[987]))):InitCond[917];
    m[990] = run?((((m[972]&~m[988]&~m[989]&~m[991]&~m[992])|(~m[972]&~m[988]&~m[989]&m[991]&~m[992])|(m[972]&m[988]&~m[989]&m[991]&~m[992])|(m[972]&~m[988]&m[989]&m[991]&~m[992])|(~m[972]&m[988]&~m[989]&~m[991]&m[992])|(~m[972]&~m[988]&m[989]&~m[991]&m[992])|(m[972]&m[988]&m[989]&~m[991]&m[992])|(~m[972]&m[988]&m[989]&m[991]&m[992]))&UnbiasedRNG[279])|((m[972]&~m[988]&~m[989]&m[991]&~m[992])|(~m[972]&~m[988]&~m[989]&~m[991]&m[992])|(m[972]&~m[988]&~m[989]&~m[991]&m[992])|(m[972]&m[988]&~m[989]&~m[991]&m[992])|(m[972]&~m[988]&m[989]&~m[991]&m[992])|(~m[972]&~m[988]&~m[989]&m[991]&m[992])|(m[972]&~m[988]&~m[989]&m[991]&m[992])|(~m[972]&m[988]&~m[989]&m[991]&m[992])|(m[972]&m[988]&~m[989]&m[991]&m[992])|(~m[972]&~m[988]&m[989]&m[991]&m[992])|(m[972]&~m[988]&m[989]&m[991]&m[992])|(m[972]&m[988]&m[989]&m[991]&m[992]))):InitCond[918];
    m[995] = run?((((m[977]&~m[993]&~m[994]&~m[996]&~m[997])|(~m[977]&~m[993]&~m[994]&m[996]&~m[997])|(m[977]&m[993]&~m[994]&m[996]&~m[997])|(m[977]&~m[993]&m[994]&m[996]&~m[997])|(~m[977]&m[993]&~m[994]&~m[996]&m[997])|(~m[977]&~m[993]&m[994]&~m[996]&m[997])|(m[977]&m[993]&m[994]&~m[996]&m[997])|(~m[977]&m[993]&m[994]&m[996]&m[997]))&UnbiasedRNG[280])|((m[977]&~m[993]&~m[994]&m[996]&~m[997])|(~m[977]&~m[993]&~m[994]&~m[996]&m[997])|(m[977]&~m[993]&~m[994]&~m[996]&m[997])|(m[977]&m[993]&~m[994]&~m[996]&m[997])|(m[977]&~m[993]&m[994]&~m[996]&m[997])|(~m[977]&~m[993]&~m[994]&m[996]&m[997])|(m[977]&~m[993]&~m[994]&m[996]&m[997])|(~m[977]&m[993]&~m[994]&m[996]&m[997])|(m[977]&m[993]&~m[994]&m[996]&m[997])|(~m[977]&~m[993]&m[994]&m[996]&m[997])|(m[977]&~m[993]&m[994]&m[996]&m[997])|(m[977]&m[993]&m[994]&m[996]&m[997]))):InitCond[919];
    m[1005] = run?((((m[982]&~m[1003]&~m[1004]&~m[1006]&~m[1007])|(~m[982]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(m[982]&m[1003]&~m[1004]&m[1006]&~m[1007])|(m[982]&~m[1003]&m[1004]&m[1006]&~m[1007])|(~m[982]&m[1003]&~m[1004]&~m[1006]&m[1007])|(~m[982]&~m[1003]&m[1004]&~m[1006]&m[1007])|(m[982]&m[1003]&m[1004]&~m[1006]&m[1007])|(~m[982]&m[1003]&m[1004]&m[1006]&m[1007]))&UnbiasedRNG[281])|((m[982]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(~m[982]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[982]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[982]&m[1003]&~m[1004]&~m[1006]&m[1007])|(m[982]&~m[1003]&m[1004]&~m[1006]&m[1007])|(~m[982]&~m[1003]&~m[1004]&m[1006]&m[1007])|(m[982]&~m[1003]&~m[1004]&m[1006]&m[1007])|(~m[982]&m[1003]&~m[1004]&m[1006]&m[1007])|(m[982]&m[1003]&~m[1004]&m[1006]&m[1007])|(~m[982]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[982]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[982]&m[1003]&m[1004]&m[1006]&m[1007]))):InitCond[920];
    m[1010] = run?((((m[987]&~m[1008]&~m[1009]&~m[1011]&~m[1012])|(~m[987]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(m[987]&m[1008]&~m[1009]&m[1011]&~m[1012])|(m[987]&~m[1008]&m[1009]&m[1011]&~m[1012])|(~m[987]&m[1008]&~m[1009]&~m[1011]&m[1012])|(~m[987]&~m[1008]&m[1009]&~m[1011]&m[1012])|(m[987]&m[1008]&m[1009]&~m[1011]&m[1012])|(~m[987]&m[1008]&m[1009]&m[1011]&m[1012]))&UnbiasedRNG[282])|((m[987]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(~m[987]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[987]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[987]&m[1008]&~m[1009]&~m[1011]&m[1012])|(m[987]&~m[1008]&m[1009]&~m[1011]&m[1012])|(~m[987]&~m[1008]&~m[1009]&m[1011]&m[1012])|(m[987]&~m[1008]&~m[1009]&m[1011]&m[1012])|(~m[987]&m[1008]&~m[1009]&m[1011]&m[1012])|(m[987]&m[1008]&~m[1009]&m[1011]&m[1012])|(~m[987]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[987]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[987]&m[1008]&m[1009]&m[1011]&m[1012]))):InitCond[921];
    m[1015] = run?((((m[992]&~m[1013]&~m[1014]&~m[1016]&~m[1017])|(~m[992]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(m[992]&m[1013]&~m[1014]&m[1016]&~m[1017])|(m[992]&~m[1013]&m[1014]&m[1016]&~m[1017])|(~m[992]&m[1013]&~m[1014]&~m[1016]&m[1017])|(~m[992]&~m[1013]&m[1014]&~m[1016]&m[1017])|(m[992]&m[1013]&m[1014]&~m[1016]&m[1017])|(~m[992]&m[1013]&m[1014]&m[1016]&m[1017]))&UnbiasedRNG[283])|((m[992]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(~m[992]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[992]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[992]&m[1013]&~m[1014]&~m[1016]&m[1017])|(m[992]&~m[1013]&m[1014]&~m[1016]&m[1017])|(~m[992]&~m[1013]&~m[1014]&m[1016]&m[1017])|(m[992]&~m[1013]&~m[1014]&m[1016]&m[1017])|(~m[992]&m[1013]&~m[1014]&m[1016]&m[1017])|(m[992]&m[1013]&~m[1014]&m[1016]&m[1017])|(~m[992]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[992]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[992]&m[1013]&m[1014]&m[1016]&m[1017]))):InitCond[922];
    m[1020] = run?((((m[997]&~m[1018]&~m[1019]&~m[1021]&~m[1022])|(~m[997]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(m[997]&m[1018]&~m[1019]&m[1021]&~m[1022])|(m[997]&~m[1018]&m[1019]&m[1021]&~m[1022])|(~m[997]&m[1018]&~m[1019]&~m[1021]&m[1022])|(~m[997]&~m[1018]&m[1019]&~m[1021]&m[1022])|(m[997]&m[1018]&m[1019]&~m[1021]&m[1022])|(~m[997]&m[1018]&m[1019]&m[1021]&m[1022]))&UnbiasedRNG[284])|((m[997]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(~m[997]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[997]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[997]&m[1018]&~m[1019]&~m[1021]&m[1022])|(m[997]&~m[1018]&m[1019]&~m[1021]&m[1022])|(~m[997]&~m[1018]&~m[1019]&m[1021]&m[1022])|(m[997]&~m[1018]&~m[1019]&m[1021]&m[1022])|(~m[997]&m[1018]&~m[1019]&m[1021]&m[1022])|(m[997]&m[1018]&~m[1019]&m[1021]&m[1022])|(~m[997]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[997]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[997]&m[1018]&m[1019]&m[1021]&m[1022]))):InitCond[923];
    m[1025] = run?((((m[1002]&~m[1023]&~m[1024]&~m[1026]&~m[1027])|(~m[1002]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(m[1002]&m[1023]&~m[1024]&m[1026]&~m[1027])|(m[1002]&~m[1023]&m[1024]&m[1026]&~m[1027])|(~m[1002]&m[1023]&~m[1024]&~m[1026]&m[1027])|(~m[1002]&~m[1023]&m[1024]&~m[1026]&m[1027])|(m[1002]&m[1023]&m[1024]&~m[1026]&m[1027])|(~m[1002]&m[1023]&m[1024]&m[1026]&m[1027]))&UnbiasedRNG[285])|((m[1002]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(~m[1002]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[1002]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[1002]&m[1023]&~m[1024]&~m[1026]&m[1027])|(m[1002]&~m[1023]&m[1024]&~m[1026]&m[1027])|(~m[1002]&~m[1023]&~m[1024]&m[1026]&m[1027])|(m[1002]&~m[1023]&~m[1024]&m[1026]&m[1027])|(~m[1002]&m[1023]&~m[1024]&m[1026]&m[1027])|(m[1002]&m[1023]&~m[1024]&m[1026]&m[1027])|(~m[1002]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[1002]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[1002]&m[1023]&m[1024]&m[1026]&m[1027]))):InitCond[924];
    m[1035] = run?((((m[1007]&~m[1033]&~m[1034]&~m[1036]&~m[1037])|(~m[1007]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(m[1007]&m[1033]&~m[1034]&m[1036]&~m[1037])|(m[1007]&~m[1033]&m[1034]&m[1036]&~m[1037])|(~m[1007]&m[1033]&~m[1034]&~m[1036]&m[1037])|(~m[1007]&~m[1033]&m[1034]&~m[1036]&m[1037])|(m[1007]&m[1033]&m[1034]&~m[1036]&m[1037])|(~m[1007]&m[1033]&m[1034]&m[1036]&m[1037]))&UnbiasedRNG[286])|((m[1007]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(~m[1007]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[1007]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[1007]&m[1033]&~m[1034]&~m[1036]&m[1037])|(m[1007]&~m[1033]&m[1034]&~m[1036]&m[1037])|(~m[1007]&~m[1033]&~m[1034]&m[1036]&m[1037])|(m[1007]&~m[1033]&~m[1034]&m[1036]&m[1037])|(~m[1007]&m[1033]&~m[1034]&m[1036]&m[1037])|(m[1007]&m[1033]&~m[1034]&m[1036]&m[1037])|(~m[1007]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[1007]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[1007]&m[1033]&m[1034]&m[1036]&m[1037]))):InitCond[925];
    m[1040] = run?((((m[1012]&~m[1038]&~m[1039]&~m[1041]&~m[1042])|(~m[1012]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1012]&m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1012]&~m[1038]&m[1039]&m[1041]&~m[1042])|(~m[1012]&m[1038]&~m[1039]&~m[1041]&m[1042])|(~m[1012]&~m[1038]&m[1039]&~m[1041]&m[1042])|(m[1012]&m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1012]&m[1038]&m[1039]&m[1041]&m[1042]))&UnbiasedRNG[287])|((m[1012]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(~m[1012]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1012]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1012]&m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1012]&~m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1012]&~m[1038]&~m[1039]&m[1041]&m[1042])|(m[1012]&~m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1012]&m[1038]&~m[1039]&m[1041]&m[1042])|(m[1012]&m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1012]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1012]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1012]&m[1038]&m[1039]&m[1041]&m[1042]))):InitCond[926];
    m[1045] = run?((((m[1017]&~m[1043]&~m[1044]&~m[1046]&~m[1047])|(~m[1017]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1017]&m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1017]&~m[1043]&m[1044]&m[1046]&~m[1047])|(~m[1017]&m[1043]&~m[1044]&~m[1046]&m[1047])|(~m[1017]&~m[1043]&m[1044]&~m[1046]&m[1047])|(m[1017]&m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1017]&m[1043]&m[1044]&m[1046]&m[1047]))&UnbiasedRNG[288])|((m[1017]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(~m[1017]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1017]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1017]&m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1017]&~m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1017]&~m[1043]&~m[1044]&m[1046]&m[1047])|(m[1017]&~m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1017]&m[1043]&~m[1044]&m[1046]&m[1047])|(m[1017]&m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1017]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1017]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1017]&m[1043]&m[1044]&m[1046]&m[1047]))):InitCond[927];
    m[1050] = run?((((m[1022]&~m[1048]&~m[1049]&~m[1051]&~m[1052])|(~m[1022]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1022]&m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1022]&~m[1048]&m[1049]&m[1051]&~m[1052])|(~m[1022]&m[1048]&~m[1049]&~m[1051]&m[1052])|(~m[1022]&~m[1048]&m[1049]&~m[1051]&m[1052])|(m[1022]&m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1022]&m[1048]&m[1049]&m[1051]&m[1052]))&UnbiasedRNG[289])|((m[1022]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(~m[1022]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1022]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1022]&m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1022]&~m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1022]&~m[1048]&~m[1049]&m[1051]&m[1052])|(m[1022]&~m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1022]&m[1048]&~m[1049]&m[1051]&m[1052])|(m[1022]&m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1022]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1022]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1022]&m[1048]&m[1049]&m[1051]&m[1052]))):InitCond[928];
    m[1055] = run?((((m[1027]&~m[1053]&~m[1054]&~m[1056]&~m[1057])|(~m[1027]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1027]&m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1027]&~m[1053]&m[1054]&m[1056]&~m[1057])|(~m[1027]&m[1053]&~m[1054]&~m[1056]&m[1057])|(~m[1027]&~m[1053]&m[1054]&~m[1056]&m[1057])|(m[1027]&m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1027]&m[1053]&m[1054]&m[1056]&m[1057]))&UnbiasedRNG[290])|((m[1027]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(~m[1027]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1027]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1027]&m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1027]&~m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1027]&~m[1053]&~m[1054]&m[1056]&m[1057])|(m[1027]&~m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1027]&m[1053]&~m[1054]&m[1056]&m[1057])|(m[1027]&m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1027]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1027]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1027]&m[1053]&m[1054]&m[1056]&m[1057]))):InitCond[929];
    m[1060] = run?((((m[1032]&~m[1058]&~m[1059]&~m[1061]&~m[1062])|(~m[1032]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1032]&m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1032]&~m[1058]&m[1059]&m[1061]&~m[1062])|(~m[1032]&m[1058]&~m[1059]&~m[1061]&m[1062])|(~m[1032]&~m[1058]&m[1059]&~m[1061]&m[1062])|(m[1032]&m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1032]&m[1058]&m[1059]&m[1061]&m[1062]))&UnbiasedRNG[291])|((m[1032]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(~m[1032]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1032]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1032]&m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1032]&~m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1032]&~m[1058]&~m[1059]&m[1061]&m[1062])|(m[1032]&~m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1032]&m[1058]&~m[1059]&m[1061]&m[1062])|(m[1032]&m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1032]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1032]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1032]&m[1058]&m[1059]&m[1061]&m[1062]))):InitCond[930];
    m[1070] = run?((((m[1037]&~m[1068]&~m[1069]&~m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&~m[1072])|(~m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&m[1068]&m[1069]&m[1071]&m[1072]))&UnbiasedRNG[292])|((m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&m[1071]&m[1072]))):InitCond[931];
    m[1075] = run?((((m[1042]&~m[1073]&~m[1074]&~m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&~m[1077])|(~m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&m[1073]&m[1074]&m[1076]&m[1077]))&UnbiasedRNG[293])|((m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&m[1076]&m[1077]))):InitCond[932];
    m[1080] = run?((((m[1047]&~m[1078]&~m[1079]&~m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&~m[1082])|(~m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&m[1078]&m[1079]&m[1081]&m[1082]))&UnbiasedRNG[294])|((m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&m[1081]&m[1082]))):InitCond[933];
    m[1085] = run?((((m[1052]&~m[1083]&~m[1084]&~m[1086]&~m[1087])|(~m[1052]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1052]&m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1052]&~m[1083]&m[1084]&m[1086]&~m[1087])|(~m[1052]&m[1083]&~m[1084]&~m[1086]&m[1087])|(~m[1052]&~m[1083]&m[1084]&~m[1086]&m[1087])|(m[1052]&m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1052]&m[1083]&m[1084]&m[1086]&m[1087]))&UnbiasedRNG[295])|((m[1052]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(~m[1052]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1052]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1052]&m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1052]&~m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1052]&~m[1083]&~m[1084]&m[1086]&m[1087])|(m[1052]&~m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1052]&m[1083]&~m[1084]&m[1086]&m[1087])|(m[1052]&m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1052]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1052]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1052]&m[1083]&m[1084]&m[1086]&m[1087]))):InitCond[934];
    m[1090] = run?((((m[1057]&~m[1088]&~m[1089]&~m[1091]&~m[1092])|(~m[1057]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1057]&m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1057]&~m[1088]&m[1089]&m[1091]&~m[1092])|(~m[1057]&m[1088]&~m[1089]&~m[1091]&m[1092])|(~m[1057]&~m[1088]&m[1089]&~m[1091]&m[1092])|(m[1057]&m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1057]&m[1088]&m[1089]&m[1091]&m[1092]))&UnbiasedRNG[296])|((m[1057]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(~m[1057]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1057]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1057]&m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1057]&~m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1057]&~m[1088]&~m[1089]&m[1091]&m[1092])|(m[1057]&~m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1057]&m[1088]&~m[1089]&m[1091]&m[1092])|(m[1057]&m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1057]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1057]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1057]&m[1088]&m[1089]&m[1091]&m[1092]))):InitCond[935];
    m[1095] = run?((((m[1062]&~m[1093]&~m[1094]&~m[1096]&~m[1097])|(~m[1062]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1062]&m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1062]&~m[1093]&m[1094]&m[1096]&~m[1097])|(~m[1062]&m[1093]&~m[1094]&~m[1096]&m[1097])|(~m[1062]&~m[1093]&m[1094]&~m[1096]&m[1097])|(m[1062]&m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1062]&m[1093]&m[1094]&m[1096]&m[1097]))&UnbiasedRNG[297])|((m[1062]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(~m[1062]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1062]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1062]&m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1062]&~m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1062]&~m[1093]&~m[1094]&m[1096]&m[1097])|(m[1062]&~m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1062]&m[1093]&~m[1094]&m[1096]&m[1097])|(m[1062]&m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1062]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1062]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1062]&m[1093]&m[1094]&m[1096]&m[1097]))):InitCond[936];
    m[1100] = run?((((m[1067]&~m[1098]&~m[1099]&~m[1101]&~m[1102])|(~m[1067]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1067]&m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1067]&~m[1098]&m[1099]&m[1101]&~m[1102])|(~m[1067]&m[1098]&~m[1099]&~m[1101]&m[1102])|(~m[1067]&~m[1098]&m[1099]&~m[1101]&m[1102])|(m[1067]&m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1067]&m[1098]&m[1099]&m[1101]&m[1102]))&UnbiasedRNG[298])|((m[1067]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(~m[1067]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1067]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1067]&m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1067]&~m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1067]&~m[1098]&~m[1099]&m[1101]&m[1102])|(m[1067]&~m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1067]&m[1098]&~m[1099]&m[1101]&m[1102])|(m[1067]&m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1067]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1067]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1067]&m[1098]&m[1099]&m[1101]&m[1102]))):InitCond[937];
    m[1110] = run?((((m[1072]&~m[1108]&~m[1109]&~m[1111]&~m[1112])|(~m[1072]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1072]&m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1072]&~m[1108]&m[1109]&m[1111]&~m[1112])|(~m[1072]&m[1108]&~m[1109]&~m[1111]&m[1112])|(~m[1072]&~m[1108]&m[1109]&~m[1111]&m[1112])|(m[1072]&m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1072]&m[1108]&m[1109]&m[1111]&m[1112]))&UnbiasedRNG[299])|((m[1072]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(~m[1072]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1072]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1072]&m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1072]&~m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1072]&~m[1108]&~m[1109]&m[1111]&m[1112])|(m[1072]&~m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1072]&m[1108]&~m[1109]&m[1111]&m[1112])|(m[1072]&m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1072]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1072]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1072]&m[1108]&m[1109]&m[1111]&m[1112]))):InitCond[938];
    m[1115] = run?((((m[1077]&~m[1113]&~m[1114]&~m[1116]&~m[1117])|(~m[1077]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1077]&m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1077]&~m[1113]&m[1114]&m[1116]&~m[1117])|(~m[1077]&m[1113]&~m[1114]&~m[1116]&m[1117])|(~m[1077]&~m[1113]&m[1114]&~m[1116]&m[1117])|(m[1077]&m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1077]&m[1113]&m[1114]&m[1116]&m[1117]))&UnbiasedRNG[300])|((m[1077]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(~m[1077]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1077]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1077]&m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1077]&~m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1077]&~m[1113]&~m[1114]&m[1116]&m[1117])|(m[1077]&~m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1077]&m[1113]&~m[1114]&m[1116]&m[1117])|(m[1077]&m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1077]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1077]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1077]&m[1113]&m[1114]&m[1116]&m[1117]))):InitCond[939];
    m[1120] = run?((((m[1082]&~m[1118]&~m[1119]&~m[1121]&~m[1122])|(~m[1082]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1082]&m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1082]&~m[1118]&m[1119]&m[1121]&~m[1122])|(~m[1082]&m[1118]&~m[1119]&~m[1121]&m[1122])|(~m[1082]&~m[1118]&m[1119]&~m[1121]&m[1122])|(m[1082]&m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1082]&m[1118]&m[1119]&m[1121]&m[1122]))&UnbiasedRNG[301])|((m[1082]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(~m[1082]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1082]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1082]&m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1082]&~m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1082]&~m[1118]&~m[1119]&m[1121]&m[1122])|(m[1082]&~m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1082]&m[1118]&~m[1119]&m[1121]&m[1122])|(m[1082]&m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1082]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1082]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1082]&m[1118]&m[1119]&m[1121]&m[1122]))):InitCond[940];
    m[1125] = run?((((m[1087]&~m[1123]&~m[1124]&~m[1126]&~m[1127])|(~m[1087]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1087]&m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1087]&~m[1123]&m[1124]&m[1126]&~m[1127])|(~m[1087]&m[1123]&~m[1124]&~m[1126]&m[1127])|(~m[1087]&~m[1123]&m[1124]&~m[1126]&m[1127])|(m[1087]&m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1087]&m[1123]&m[1124]&m[1126]&m[1127]))&UnbiasedRNG[302])|((m[1087]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(~m[1087]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1087]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1087]&m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1087]&~m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1087]&~m[1123]&~m[1124]&m[1126]&m[1127])|(m[1087]&~m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1087]&m[1123]&~m[1124]&m[1126]&m[1127])|(m[1087]&m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1087]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1087]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1087]&m[1123]&m[1124]&m[1126]&m[1127]))):InitCond[941];
    m[1130] = run?((((m[1092]&~m[1128]&~m[1129]&~m[1131]&~m[1132])|(~m[1092]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1092]&m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1092]&~m[1128]&m[1129]&m[1131]&~m[1132])|(~m[1092]&m[1128]&~m[1129]&~m[1131]&m[1132])|(~m[1092]&~m[1128]&m[1129]&~m[1131]&m[1132])|(m[1092]&m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1092]&m[1128]&m[1129]&m[1131]&m[1132]))&UnbiasedRNG[303])|((m[1092]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(~m[1092]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1092]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1092]&m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1092]&~m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1092]&~m[1128]&~m[1129]&m[1131]&m[1132])|(m[1092]&~m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1092]&m[1128]&~m[1129]&m[1131]&m[1132])|(m[1092]&m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1092]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1092]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1092]&m[1128]&m[1129]&m[1131]&m[1132]))):InitCond[942];
    m[1135] = run?((((m[1097]&~m[1133]&~m[1134]&~m[1136]&~m[1137])|(~m[1097]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1097]&m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1097]&~m[1133]&m[1134]&m[1136]&~m[1137])|(~m[1097]&m[1133]&~m[1134]&~m[1136]&m[1137])|(~m[1097]&~m[1133]&m[1134]&~m[1136]&m[1137])|(m[1097]&m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1097]&m[1133]&m[1134]&m[1136]&m[1137]))&UnbiasedRNG[304])|((m[1097]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(~m[1097]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1097]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1097]&m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1097]&~m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1097]&~m[1133]&~m[1134]&m[1136]&m[1137])|(m[1097]&~m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1097]&m[1133]&~m[1134]&m[1136]&m[1137])|(m[1097]&m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1097]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1097]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1097]&m[1133]&m[1134]&m[1136]&m[1137]))):InitCond[943];
    m[1140] = run?((((m[1102]&~m[1138]&~m[1139]&~m[1141]&~m[1142])|(~m[1102]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1102]&m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1102]&~m[1138]&m[1139]&m[1141]&~m[1142])|(~m[1102]&m[1138]&~m[1139]&~m[1141]&m[1142])|(~m[1102]&~m[1138]&m[1139]&~m[1141]&m[1142])|(m[1102]&m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1102]&m[1138]&m[1139]&m[1141]&m[1142]))&UnbiasedRNG[305])|((m[1102]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(~m[1102]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1102]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1102]&m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1102]&~m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1102]&~m[1138]&~m[1139]&m[1141]&m[1142])|(m[1102]&~m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1102]&m[1138]&~m[1139]&m[1141]&m[1142])|(m[1102]&m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1102]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1102]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1102]&m[1138]&m[1139]&m[1141]&m[1142]))):InitCond[944];
    m[1145] = run?((((m[1107]&~m[1143]&~m[1144]&~m[1146]&~m[1147])|(~m[1107]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1107]&m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1107]&~m[1143]&m[1144]&m[1146]&~m[1147])|(~m[1107]&m[1143]&~m[1144]&~m[1146]&m[1147])|(~m[1107]&~m[1143]&m[1144]&~m[1146]&m[1147])|(m[1107]&m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1107]&m[1143]&m[1144]&m[1146]&m[1147]))&UnbiasedRNG[306])|((m[1107]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(~m[1107]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1107]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1107]&m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1107]&~m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1107]&~m[1143]&~m[1144]&m[1146]&m[1147])|(m[1107]&~m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1107]&m[1143]&~m[1144]&m[1146]&m[1147])|(m[1107]&m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1107]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1107]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1107]&m[1143]&m[1144]&m[1146]&m[1147]))):InitCond[945];
    m[1155] = run?((((m[1112]&~m[1153]&~m[1154]&~m[1156]&~m[1157])|(~m[1112]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1112]&m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1112]&~m[1153]&m[1154]&m[1156]&~m[1157])|(~m[1112]&m[1153]&~m[1154]&~m[1156]&m[1157])|(~m[1112]&~m[1153]&m[1154]&~m[1156]&m[1157])|(m[1112]&m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1112]&m[1153]&m[1154]&m[1156]&m[1157]))&UnbiasedRNG[307])|((m[1112]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(~m[1112]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1112]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1112]&m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1112]&~m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1112]&~m[1153]&~m[1154]&m[1156]&m[1157])|(m[1112]&~m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1112]&m[1153]&~m[1154]&m[1156]&m[1157])|(m[1112]&m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1112]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1112]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1112]&m[1153]&m[1154]&m[1156]&m[1157]))):InitCond[946];
    m[1160] = run?((((m[1117]&~m[1158]&~m[1159]&~m[1161]&~m[1162])|(~m[1117]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1117]&m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1117]&~m[1158]&m[1159]&m[1161]&~m[1162])|(~m[1117]&m[1158]&~m[1159]&~m[1161]&m[1162])|(~m[1117]&~m[1158]&m[1159]&~m[1161]&m[1162])|(m[1117]&m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1117]&m[1158]&m[1159]&m[1161]&m[1162]))&UnbiasedRNG[308])|((m[1117]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(~m[1117]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1117]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1117]&m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1117]&~m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1117]&~m[1158]&~m[1159]&m[1161]&m[1162])|(m[1117]&~m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1117]&m[1158]&~m[1159]&m[1161]&m[1162])|(m[1117]&m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1117]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1117]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1117]&m[1158]&m[1159]&m[1161]&m[1162]))):InitCond[947];
    m[1165] = run?((((m[1122]&~m[1163]&~m[1164]&~m[1166]&~m[1167])|(~m[1122]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1122]&m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1122]&~m[1163]&m[1164]&m[1166]&~m[1167])|(~m[1122]&m[1163]&~m[1164]&~m[1166]&m[1167])|(~m[1122]&~m[1163]&m[1164]&~m[1166]&m[1167])|(m[1122]&m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1122]&m[1163]&m[1164]&m[1166]&m[1167]))&UnbiasedRNG[309])|((m[1122]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(~m[1122]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1122]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1122]&m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1122]&~m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1122]&~m[1163]&~m[1164]&m[1166]&m[1167])|(m[1122]&~m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1122]&m[1163]&~m[1164]&m[1166]&m[1167])|(m[1122]&m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1122]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1122]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1122]&m[1163]&m[1164]&m[1166]&m[1167]))):InitCond[948];
    m[1170] = run?((((m[1127]&~m[1168]&~m[1169]&~m[1171]&~m[1172])|(~m[1127]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1127]&m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1127]&~m[1168]&m[1169]&m[1171]&~m[1172])|(~m[1127]&m[1168]&~m[1169]&~m[1171]&m[1172])|(~m[1127]&~m[1168]&m[1169]&~m[1171]&m[1172])|(m[1127]&m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1127]&m[1168]&m[1169]&m[1171]&m[1172]))&UnbiasedRNG[310])|((m[1127]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(~m[1127]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1127]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1127]&m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1127]&~m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1127]&~m[1168]&~m[1169]&m[1171]&m[1172])|(m[1127]&~m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1127]&m[1168]&~m[1169]&m[1171]&m[1172])|(m[1127]&m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1127]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1127]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1127]&m[1168]&m[1169]&m[1171]&m[1172]))):InitCond[949];
    m[1175] = run?((((m[1132]&~m[1173]&~m[1174]&~m[1176]&~m[1177])|(~m[1132]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1132]&m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1132]&~m[1173]&m[1174]&m[1176]&~m[1177])|(~m[1132]&m[1173]&~m[1174]&~m[1176]&m[1177])|(~m[1132]&~m[1173]&m[1174]&~m[1176]&m[1177])|(m[1132]&m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1132]&m[1173]&m[1174]&m[1176]&m[1177]))&UnbiasedRNG[311])|((m[1132]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(~m[1132]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1132]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1132]&m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1132]&~m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1132]&~m[1173]&~m[1174]&m[1176]&m[1177])|(m[1132]&~m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1132]&m[1173]&~m[1174]&m[1176]&m[1177])|(m[1132]&m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1132]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1132]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1132]&m[1173]&m[1174]&m[1176]&m[1177]))):InitCond[950];
    m[1180] = run?((((m[1137]&~m[1178]&~m[1179]&~m[1181]&~m[1182])|(~m[1137]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1137]&m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1137]&~m[1178]&m[1179]&m[1181]&~m[1182])|(~m[1137]&m[1178]&~m[1179]&~m[1181]&m[1182])|(~m[1137]&~m[1178]&m[1179]&~m[1181]&m[1182])|(m[1137]&m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1137]&m[1178]&m[1179]&m[1181]&m[1182]))&UnbiasedRNG[312])|((m[1137]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(~m[1137]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1137]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1137]&m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1137]&~m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1137]&~m[1178]&~m[1179]&m[1181]&m[1182])|(m[1137]&~m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1137]&m[1178]&~m[1179]&m[1181]&m[1182])|(m[1137]&m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1137]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1137]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1137]&m[1178]&m[1179]&m[1181]&m[1182]))):InitCond[951];
    m[1185] = run?((((m[1142]&~m[1183]&~m[1184]&~m[1186]&~m[1187])|(~m[1142]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1142]&m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1142]&~m[1183]&m[1184]&m[1186]&~m[1187])|(~m[1142]&m[1183]&~m[1184]&~m[1186]&m[1187])|(~m[1142]&~m[1183]&m[1184]&~m[1186]&m[1187])|(m[1142]&m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1142]&m[1183]&m[1184]&m[1186]&m[1187]))&UnbiasedRNG[313])|((m[1142]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(~m[1142]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1142]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1142]&m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1142]&~m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1142]&~m[1183]&~m[1184]&m[1186]&m[1187])|(m[1142]&~m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1142]&m[1183]&~m[1184]&m[1186]&m[1187])|(m[1142]&m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1142]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1142]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1142]&m[1183]&m[1184]&m[1186]&m[1187]))):InitCond[952];
    m[1190] = run?((((m[1147]&~m[1188]&~m[1189]&~m[1191]&~m[1192])|(~m[1147]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1147]&m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1147]&~m[1188]&m[1189]&m[1191]&~m[1192])|(~m[1147]&m[1188]&~m[1189]&~m[1191]&m[1192])|(~m[1147]&~m[1188]&m[1189]&~m[1191]&m[1192])|(m[1147]&m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1147]&m[1188]&m[1189]&m[1191]&m[1192]))&UnbiasedRNG[314])|((m[1147]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(~m[1147]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1147]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1147]&m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1147]&~m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1147]&~m[1188]&~m[1189]&m[1191]&m[1192])|(m[1147]&~m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1147]&m[1188]&~m[1189]&m[1191]&m[1192])|(m[1147]&m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1147]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1147]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1147]&m[1188]&m[1189]&m[1191]&m[1192]))):InitCond[953];
    m[1195] = run?((((m[1152]&~m[1193]&~m[1194]&~m[1196]&~m[1197])|(~m[1152]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1152]&m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1152]&~m[1193]&m[1194]&m[1196]&~m[1197])|(~m[1152]&m[1193]&~m[1194]&~m[1196]&m[1197])|(~m[1152]&~m[1193]&m[1194]&~m[1196]&m[1197])|(m[1152]&m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1152]&m[1193]&m[1194]&m[1196]&m[1197]))&UnbiasedRNG[315])|((m[1152]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(~m[1152]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1152]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1152]&m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1152]&~m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1152]&~m[1193]&~m[1194]&m[1196]&m[1197])|(m[1152]&~m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1152]&m[1193]&~m[1194]&m[1196]&m[1197])|(m[1152]&m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1152]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1152]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1152]&m[1193]&m[1194]&m[1196]&m[1197]))):InitCond[954];
    m[1205] = run?((((m[1157]&~m[1203]&~m[1204]&~m[1206]&~m[1207])|(~m[1157]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1157]&m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1157]&~m[1203]&m[1204]&m[1206]&~m[1207])|(~m[1157]&m[1203]&~m[1204]&~m[1206]&m[1207])|(~m[1157]&~m[1203]&m[1204]&~m[1206]&m[1207])|(m[1157]&m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1157]&m[1203]&m[1204]&m[1206]&m[1207]))&UnbiasedRNG[316])|((m[1157]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(~m[1157]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1157]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1157]&m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1157]&~m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1157]&~m[1203]&~m[1204]&m[1206]&m[1207])|(m[1157]&~m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1157]&m[1203]&~m[1204]&m[1206]&m[1207])|(m[1157]&m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1157]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1157]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1157]&m[1203]&m[1204]&m[1206]&m[1207]))):InitCond[955];
    m[1210] = run?((((m[1162]&~m[1208]&~m[1209]&~m[1211]&~m[1212])|(~m[1162]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1162]&m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1162]&~m[1208]&m[1209]&m[1211]&~m[1212])|(~m[1162]&m[1208]&~m[1209]&~m[1211]&m[1212])|(~m[1162]&~m[1208]&m[1209]&~m[1211]&m[1212])|(m[1162]&m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1162]&m[1208]&m[1209]&m[1211]&m[1212]))&UnbiasedRNG[317])|((m[1162]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(~m[1162]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1162]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1162]&m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1162]&~m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1162]&~m[1208]&~m[1209]&m[1211]&m[1212])|(m[1162]&~m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1162]&m[1208]&~m[1209]&m[1211]&m[1212])|(m[1162]&m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1162]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1162]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1162]&m[1208]&m[1209]&m[1211]&m[1212]))):InitCond[956];
    m[1215] = run?((((m[1167]&~m[1213]&~m[1214]&~m[1216]&~m[1217])|(~m[1167]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1167]&m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1167]&~m[1213]&m[1214]&m[1216]&~m[1217])|(~m[1167]&m[1213]&~m[1214]&~m[1216]&m[1217])|(~m[1167]&~m[1213]&m[1214]&~m[1216]&m[1217])|(m[1167]&m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1167]&m[1213]&m[1214]&m[1216]&m[1217]))&UnbiasedRNG[318])|((m[1167]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(~m[1167]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1167]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1167]&m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1167]&~m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1167]&~m[1213]&~m[1214]&m[1216]&m[1217])|(m[1167]&~m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1167]&m[1213]&~m[1214]&m[1216]&m[1217])|(m[1167]&m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1167]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1167]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1167]&m[1213]&m[1214]&m[1216]&m[1217]))):InitCond[957];
    m[1220] = run?((((m[1172]&~m[1218]&~m[1219]&~m[1221]&~m[1222])|(~m[1172]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1172]&m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1172]&~m[1218]&m[1219]&m[1221]&~m[1222])|(~m[1172]&m[1218]&~m[1219]&~m[1221]&m[1222])|(~m[1172]&~m[1218]&m[1219]&~m[1221]&m[1222])|(m[1172]&m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1172]&m[1218]&m[1219]&m[1221]&m[1222]))&UnbiasedRNG[319])|((m[1172]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(~m[1172]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1172]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1172]&m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1172]&~m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1172]&~m[1218]&~m[1219]&m[1221]&m[1222])|(m[1172]&~m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1172]&m[1218]&~m[1219]&m[1221]&m[1222])|(m[1172]&m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1172]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1172]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1172]&m[1218]&m[1219]&m[1221]&m[1222]))):InitCond[958];
    m[1225] = run?((((m[1177]&~m[1223]&~m[1224]&~m[1226]&~m[1227])|(~m[1177]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1177]&m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1177]&~m[1223]&m[1224]&m[1226]&~m[1227])|(~m[1177]&m[1223]&~m[1224]&~m[1226]&m[1227])|(~m[1177]&~m[1223]&m[1224]&~m[1226]&m[1227])|(m[1177]&m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1177]&m[1223]&m[1224]&m[1226]&m[1227]))&UnbiasedRNG[320])|((m[1177]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(~m[1177]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1177]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1177]&m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1177]&~m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1177]&~m[1223]&~m[1224]&m[1226]&m[1227])|(m[1177]&~m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1177]&m[1223]&~m[1224]&m[1226]&m[1227])|(m[1177]&m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1177]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1177]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1177]&m[1223]&m[1224]&m[1226]&m[1227]))):InitCond[959];
    m[1230] = run?((((m[1182]&~m[1228]&~m[1229]&~m[1231]&~m[1232])|(~m[1182]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1182]&m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1182]&~m[1228]&m[1229]&m[1231]&~m[1232])|(~m[1182]&m[1228]&~m[1229]&~m[1231]&m[1232])|(~m[1182]&~m[1228]&m[1229]&~m[1231]&m[1232])|(m[1182]&m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1182]&m[1228]&m[1229]&m[1231]&m[1232]))&UnbiasedRNG[321])|((m[1182]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(~m[1182]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1182]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1182]&m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1182]&~m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1182]&~m[1228]&~m[1229]&m[1231]&m[1232])|(m[1182]&~m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1182]&m[1228]&~m[1229]&m[1231]&m[1232])|(m[1182]&m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1182]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1182]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1182]&m[1228]&m[1229]&m[1231]&m[1232]))):InitCond[960];
    m[1235] = run?((((m[1187]&~m[1233]&~m[1234]&~m[1236]&~m[1237])|(~m[1187]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1187]&m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1187]&~m[1233]&m[1234]&m[1236]&~m[1237])|(~m[1187]&m[1233]&~m[1234]&~m[1236]&m[1237])|(~m[1187]&~m[1233]&m[1234]&~m[1236]&m[1237])|(m[1187]&m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1187]&m[1233]&m[1234]&m[1236]&m[1237]))&UnbiasedRNG[322])|((m[1187]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(~m[1187]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1187]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1187]&m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1187]&~m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1187]&~m[1233]&~m[1234]&m[1236]&m[1237])|(m[1187]&~m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1187]&m[1233]&~m[1234]&m[1236]&m[1237])|(m[1187]&m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1187]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1187]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1187]&m[1233]&m[1234]&m[1236]&m[1237]))):InitCond[961];
    m[1240] = run?((((m[1192]&~m[1238]&~m[1239]&~m[1241]&~m[1242])|(~m[1192]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1192]&m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1192]&~m[1238]&m[1239]&m[1241]&~m[1242])|(~m[1192]&m[1238]&~m[1239]&~m[1241]&m[1242])|(~m[1192]&~m[1238]&m[1239]&~m[1241]&m[1242])|(m[1192]&m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1192]&m[1238]&m[1239]&m[1241]&m[1242]))&UnbiasedRNG[323])|((m[1192]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(~m[1192]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1192]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1192]&m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1192]&~m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1192]&~m[1238]&~m[1239]&m[1241]&m[1242])|(m[1192]&~m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1192]&m[1238]&~m[1239]&m[1241]&m[1242])|(m[1192]&m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1192]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1192]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1192]&m[1238]&m[1239]&m[1241]&m[1242]))):InitCond[962];
    m[1245] = run?((((m[1197]&~m[1243]&~m[1244]&~m[1246]&~m[1247])|(~m[1197]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1197]&m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1197]&~m[1243]&m[1244]&m[1246]&~m[1247])|(~m[1197]&m[1243]&~m[1244]&~m[1246]&m[1247])|(~m[1197]&~m[1243]&m[1244]&~m[1246]&m[1247])|(m[1197]&m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1197]&m[1243]&m[1244]&m[1246]&m[1247]))&UnbiasedRNG[324])|((m[1197]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(~m[1197]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1197]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1197]&m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1197]&~m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1197]&~m[1243]&~m[1244]&m[1246]&m[1247])|(m[1197]&~m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1197]&m[1243]&~m[1244]&m[1246]&m[1247])|(m[1197]&m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1197]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1197]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1197]&m[1243]&m[1244]&m[1246]&m[1247]))):InitCond[963];
    m[1250] = run?((((m[1202]&~m[1248]&~m[1249]&~m[1251]&~m[1252])|(~m[1202]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1202]&m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1202]&~m[1248]&m[1249]&m[1251]&~m[1252])|(~m[1202]&m[1248]&~m[1249]&~m[1251]&m[1252])|(~m[1202]&~m[1248]&m[1249]&~m[1251]&m[1252])|(m[1202]&m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1202]&m[1248]&m[1249]&m[1251]&m[1252]))&UnbiasedRNG[325])|((m[1202]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(~m[1202]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1202]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1202]&m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1202]&~m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1202]&~m[1248]&~m[1249]&m[1251]&m[1252])|(m[1202]&~m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1202]&m[1248]&~m[1249]&m[1251]&m[1252])|(m[1202]&m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1202]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1202]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1202]&m[1248]&m[1249]&m[1251]&m[1252]))):InitCond[964];
    m[1260] = run?((((m[1207]&~m[1258]&~m[1259]&~m[1261]&~m[1262])|(~m[1207]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1207]&m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1207]&~m[1258]&m[1259]&m[1261]&~m[1262])|(~m[1207]&m[1258]&~m[1259]&~m[1261]&m[1262])|(~m[1207]&~m[1258]&m[1259]&~m[1261]&m[1262])|(m[1207]&m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1207]&m[1258]&m[1259]&m[1261]&m[1262]))&UnbiasedRNG[326])|((m[1207]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(~m[1207]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1207]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1207]&m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1207]&~m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1207]&~m[1258]&~m[1259]&m[1261]&m[1262])|(m[1207]&~m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1207]&m[1258]&~m[1259]&m[1261]&m[1262])|(m[1207]&m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1207]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1207]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1207]&m[1258]&m[1259]&m[1261]&m[1262]))):InitCond[965];
    m[1265] = run?((((m[1212]&~m[1263]&~m[1264]&~m[1266]&~m[1267])|(~m[1212]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1212]&m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1212]&~m[1263]&m[1264]&m[1266]&~m[1267])|(~m[1212]&m[1263]&~m[1264]&~m[1266]&m[1267])|(~m[1212]&~m[1263]&m[1264]&~m[1266]&m[1267])|(m[1212]&m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1212]&m[1263]&m[1264]&m[1266]&m[1267]))&UnbiasedRNG[327])|((m[1212]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(~m[1212]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1212]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1212]&m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1212]&~m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1212]&~m[1263]&~m[1264]&m[1266]&m[1267])|(m[1212]&~m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1212]&m[1263]&~m[1264]&m[1266]&m[1267])|(m[1212]&m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1212]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1212]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1212]&m[1263]&m[1264]&m[1266]&m[1267]))):InitCond[966];
    m[1270] = run?((((m[1217]&~m[1268]&~m[1269]&~m[1271]&~m[1272])|(~m[1217]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1217]&m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1217]&~m[1268]&m[1269]&m[1271]&~m[1272])|(~m[1217]&m[1268]&~m[1269]&~m[1271]&m[1272])|(~m[1217]&~m[1268]&m[1269]&~m[1271]&m[1272])|(m[1217]&m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1217]&m[1268]&m[1269]&m[1271]&m[1272]))&UnbiasedRNG[328])|((m[1217]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(~m[1217]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1217]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1217]&m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1217]&~m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1217]&~m[1268]&~m[1269]&m[1271]&m[1272])|(m[1217]&~m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1217]&m[1268]&~m[1269]&m[1271]&m[1272])|(m[1217]&m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1217]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1217]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1217]&m[1268]&m[1269]&m[1271]&m[1272]))):InitCond[967];
    m[1275] = run?((((m[1222]&~m[1273]&~m[1274]&~m[1276]&~m[1277])|(~m[1222]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1222]&m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1222]&~m[1273]&m[1274]&m[1276]&~m[1277])|(~m[1222]&m[1273]&~m[1274]&~m[1276]&m[1277])|(~m[1222]&~m[1273]&m[1274]&~m[1276]&m[1277])|(m[1222]&m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1222]&m[1273]&m[1274]&m[1276]&m[1277]))&UnbiasedRNG[329])|((m[1222]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(~m[1222]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1222]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1222]&m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1222]&~m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1222]&~m[1273]&~m[1274]&m[1276]&m[1277])|(m[1222]&~m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1222]&m[1273]&~m[1274]&m[1276]&m[1277])|(m[1222]&m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1222]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1222]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1222]&m[1273]&m[1274]&m[1276]&m[1277]))):InitCond[968];
    m[1280] = run?((((m[1227]&~m[1278]&~m[1279]&~m[1281]&~m[1282])|(~m[1227]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1227]&m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1227]&~m[1278]&m[1279]&m[1281]&~m[1282])|(~m[1227]&m[1278]&~m[1279]&~m[1281]&m[1282])|(~m[1227]&~m[1278]&m[1279]&~m[1281]&m[1282])|(m[1227]&m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1227]&m[1278]&m[1279]&m[1281]&m[1282]))&UnbiasedRNG[330])|((m[1227]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(~m[1227]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1227]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1227]&m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1227]&~m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1227]&~m[1278]&~m[1279]&m[1281]&m[1282])|(m[1227]&~m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1227]&m[1278]&~m[1279]&m[1281]&m[1282])|(m[1227]&m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1227]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1227]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1227]&m[1278]&m[1279]&m[1281]&m[1282]))):InitCond[969];
    m[1285] = run?((((m[1232]&~m[1283]&~m[1284]&~m[1286]&~m[1287])|(~m[1232]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1232]&m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1232]&~m[1283]&m[1284]&m[1286]&~m[1287])|(~m[1232]&m[1283]&~m[1284]&~m[1286]&m[1287])|(~m[1232]&~m[1283]&m[1284]&~m[1286]&m[1287])|(m[1232]&m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1232]&m[1283]&m[1284]&m[1286]&m[1287]))&UnbiasedRNG[331])|((m[1232]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(~m[1232]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1232]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1232]&m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1232]&~m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1232]&~m[1283]&~m[1284]&m[1286]&m[1287])|(m[1232]&~m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1232]&m[1283]&~m[1284]&m[1286]&m[1287])|(m[1232]&m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1232]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1232]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1232]&m[1283]&m[1284]&m[1286]&m[1287]))):InitCond[970];
    m[1290] = run?((((m[1237]&~m[1288]&~m[1289]&~m[1291]&~m[1292])|(~m[1237]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1237]&m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1237]&~m[1288]&m[1289]&m[1291]&~m[1292])|(~m[1237]&m[1288]&~m[1289]&~m[1291]&m[1292])|(~m[1237]&~m[1288]&m[1289]&~m[1291]&m[1292])|(m[1237]&m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1237]&m[1288]&m[1289]&m[1291]&m[1292]))&UnbiasedRNG[332])|((m[1237]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(~m[1237]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1237]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1237]&m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1237]&~m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1237]&~m[1288]&~m[1289]&m[1291]&m[1292])|(m[1237]&~m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1237]&m[1288]&~m[1289]&m[1291]&m[1292])|(m[1237]&m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1237]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1237]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1237]&m[1288]&m[1289]&m[1291]&m[1292]))):InitCond[971];
    m[1295] = run?((((m[1242]&~m[1293]&~m[1294]&~m[1296]&~m[1297])|(~m[1242]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1242]&m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1242]&~m[1293]&m[1294]&m[1296]&~m[1297])|(~m[1242]&m[1293]&~m[1294]&~m[1296]&m[1297])|(~m[1242]&~m[1293]&m[1294]&~m[1296]&m[1297])|(m[1242]&m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1242]&m[1293]&m[1294]&m[1296]&m[1297]))&UnbiasedRNG[333])|((m[1242]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(~m[1242]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1242]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1242]&m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1242]&~m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1242]&~m[1293]&~m[1294]&m[1296]&m[1297])|(m[1242]&~m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1242]&m[1293]&~m[1294]&m[1296]&m[1297])|(m[1242]&m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1242]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1242]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1242]&m[1293]&m[1294]&m[1296]&m[1297]))):InitCond[972];
    m[1300] = run?((((m[1247]&~m[1298]&~m[1299]&~m[1301]&~m[1302])|(~m[1247]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1247]&m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1247]&~m[1298]&m[1299]&m[1301]&~m[1302])|(~m[1247]&m[1298]&~m[1299]&~m[1301]&m[1302])|(~m[1247]&~m[1298]&m[1299]&~m[1301]&m[1302])|(m[1247]&m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1247]&m[1298]&m[1299]&m[1301]&m[1302]))&UnbiasedRNG[334])|((m[1247]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(~m[1247]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1247]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1247]&m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1247]&~m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1247]&~m[1298]&~m[1299]&m[1301]&m[1302])|(m[1247]&~m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1247]&m[1298]&~m[1299]&m[1301]&m[1302])|(m[1247]&m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1247]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1247]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1247]&m[1298]&m[1299]&m[1301]&m[1302]))):InitCond[973];
    m[1305] = run?((((m[1252]&~m[1303]&~m[1304]&~m[1306]&~m[1307])|(~m[1252]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1252]&m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1252]&~m[1303]&m[1304]&m[1306]&~m[1307])|(~m[1252]&m[1303]&~m[1304]&~m[1306]&m[1307])|(~m[1252]&~m[1303]&m[1304]&~m[1306]&m[1307])|(m[1252]&m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1252]&m[1303]&m[1304]&m[1306]&m[1307]))&UnbiasedRNG[335])|((m[1252]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(~m[1252]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1252]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1252]&m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1252]&~m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1252]&~m[1303]&~m[1304]&m[1306]&m[1307])|(m[1252]&~m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1252]&m[1303]&~m[1304]&m[1306]&m[1307])|(m[1252]&m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1252]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1252]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1252]&m[1303]&m[1304]&m[1306]&m[1307]))):InitCond[974];
    m[1310] = run?((((m[1257]&~m[1308]&~m[1309]&~m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&~m[1312])|(~m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&m[1308]&m[1309]&m[1311]&m[1312]))&UnbiasedRNG[336])|((m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&m[1311]&m[1312]))):InitCond[975];
    m[1320] = run?((((m[1262]&~m[1318]&~m[1319]&~m[1321]&~m[1322])|(~m[1262]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1262]&m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1262]&~m[1318]&m[1319]&m[1321]&~m[1322])|(~m[1262]&m[1318]&~m[1319]&~m[1321]&m[1322])|(~m[1262]&~m[1318]&m[1319]&~m[1321]&m[1322])|(m[1262]&m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1262]&m[1318]&m[1319]&m[1321]&m[1322]))&UnbiasedRNG[337])|((m[1262]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(~m[1262]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1262]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1262]&m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1262]&~m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1262]&~m[1318]&~m[1319]&m[1321]&m[1322])|(m[1262]&~m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1262]&m[1318]&~m[1319]&m[1321]&m[1322])|(m[1262]&m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1262]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1262]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1262]&m[1318]&m[1319]&m[1321]&m[1322]))):InitCond[976];
    m[1325] = run?((((m[1267]&~m[1323]&~m[1324]&~m[1326]&~m[1327])|(~m[1267]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1267]&m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1267]&~m[1323]&m[1324]&m[1326]&~m[1327])|(~m[1267]&m[1323]&~m[1324]&~m[1326]&m[1327])|(~m[1267]&~m[1323]&m[1324]&~m[1326]&m[1327])|(m[1267]&m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1267]&m[1323]&m[1324]&m[1326]&m[1327]))&UnbiasedRNG[338])|((m[1267]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(~m[1267]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1267]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1267]&m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1267]&~m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1267]&~m[1323]&~m[1324]&m[1326]&m[1327])|(m[1267]&~m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1267]&m[1323]&~m[1324]&m[1326]&m[1327])|(m[1267]&m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1267]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1267]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1267]&m[1323]&m[1324]&m[1326]&m[1327]))):InitCond[977];
    m[1330] = run?((((m[1272]&~m[1328]&~m[1329]&~m[1331]&~m[1332])|(~m[1272]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1272]&m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1272]&~m[1328]&m[1329]&m[1331]&~m[1332])|(~m[1272]&m[1328]&~m[1329]&~m[1331]&m[1332])|(~m[1272]&~m[1328]&m[1329]&~m[1331]&m[1332])|(m[1272]&m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1272]&m[1328]&m[1329]&m[1331]&m[1332]))&UnbiasedRNG[339])|((m[1272]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(~m[1272]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1272]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1272]&m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1272]&~m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1272]&~m[1328]&~m[1329]&m[1331]&m[1332])|(m[1272]&~m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1272]&m[1328]&~m[1329]&m[1331]&m[1332])|(m[1272]&m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1272]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1272]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1272]&m[1328]&m[1329]&m[1331]&m[1332]))):InitCond[978];
    m[1335] = run?((((m[1277]&~m[1333]&~m[1334]&~m[1336]&~m[1337])|(~m[1277]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1277]&m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1277]&~m[1333]&m[1334]&m[1336]&~m[1337])|(~m[1277]&m[1333]&~m[1334]&~m[1336]&m[1337])|(~m[1277]&~m[1333]&m[1334]&~m[1336]&m[1337])|(m[1277]&m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1277]&m[1333]&m[1334]&m[1336]&m[1337]))&UnbiasedRNG[340])|((m[1277]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(~m[1277]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1277]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1277]&m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1277]&~m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1277]&~m[1333]&~m[1334]&m[1336]&m[1337])|(m[1277]&~m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1277]&m[1333]&~m[1334]&m[1336]&m[1337])|(m[1277]&m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1277]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1277]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1277]&m[1333]&m[1334]&m[1336]&m[1337]))):InitCond[979];
    m[1340] = run?((((m[1282]&~m[1338]&~m[1339]&~m[1341]&~m[1342])|(~m[1282]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1282]&m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1282]&~m[1338]&m[1339]&m[1341]&~m[1342])|(~m[1282]&m[1338]&~m[1339]&~m[1341]&m[1342])|(~m[1282]&~m[1338]&m[1339]&~m[1341]&m[1342])|(m[1282]&m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1282]&m[1338]&m[1339]&m[1341]&m[1342]))&UnbiasedRNG[341])|((m[1282]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(~m[1282]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1282]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1282]&m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1282]&~m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1282]&~m[1338]&~m[1339]&m[1341]&m[1342])|(m[1282]&~m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1282]&m[1338]&~m[1339]&m[1341]&m[1342])|(m[1282]&m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1282]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1282]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1282]&m[1338]&m[1339]&m[1341]&m[1342]))):InitCond[980];
    m[1345] = run?((((m[1287]&~m[1343]&~m[1344]&~m[1346]&~m[1347])|(~m[1287]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1287]&m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1287]&~m[1343]&m[1344]&m[1346]&~m[1347])|(~m[1287]&m[1343]&~m[1344]&~m[1346]&m[1347])|(~m[1287]&~m[1343]&m[1344]&~m[1346]&m[1347])|(m[1287]&m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1287]&m[1343]&m[1344]&m[1346]&m[1347]))&UnbiasedRNG[342])|((m[1287]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(~m[1287]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1287]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1287]&m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1287]&~m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1287]&~m[1343]&~m[1344]&m[1346]&m[1347])|(m[1287]&~m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1287]&m[1343]&~m[1344]&m[1346]&m[1347])|(m[1287]&m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1287]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1287]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1287]&m[1343]&m[1344]&m[1346]&m[1347]))):InitCond[981];
    m[1350] = run?((((m[1292]&~m[1348]&~m[1349]&~m[1351]&~m[1352])|(~m[1292]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1292]&m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1292]&~m[1348]&m[1349]&m[1351]&~m[1352])|(~m[1292]&m[1348]&~m[1349]&~m[1351]&m[1352])|(~m[1292]&~m[1348]&m[1349]&~m[1351]&m[1352])|(m[1292]&m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1292]&m[1348]&m[1349]&m[1351]&m[1352]))&UnbiasedRNG[343])|((m[1292]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(~m[1292]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1292]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1292]&m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1292]&~m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1292]&~m[1348]&~m[1349]&m[1351]&m[1352])|(m[1292]&~m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1292]&m[1348]&~m[1349]&m[1351]&m[1352])|(m[1292]&m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1292]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1292]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1292]&m[1348]&m[1349]&m[1351]&m[1352]))):InitCond[982];
    m[1355] = run?((((m[1297]&~m[1353]&~m[1354]&~m[1356]&~m[1357])|(~m[1297]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1297]&m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1297]&~m[1353]&m[1354]&m[1356]&~m[1357])|(~m[1297]&m[1353]&~m[1354]&~m[1356]&m[1357])|(~m[1297]&~m[1353]&m[1354]&~m[1356]&m[1357])|(m[1297]&m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1297]&m[1353]&m[1354]&m[1356]&m[1357]))&UnbiasedRNG[344])|((m[1297]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(~m[1297]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1297]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1297]&m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1297]&~m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1297]&~m[1353]&~m[1354]&m[1356]&m[1357])|(m[1297]&~m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1297]&m[1353]&~m[1354]&m[1356]&m[1357])|(m[1297]&m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1297]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1297]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1297]&m[1353]&m[1354]&m[1356]&m[1357]))):InitCond[983];
    m[1360] = run?((((m[1302]&~m[1358]&~m[1359]&~m[1361]&~m[1362])|(~m[1302]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1302]&m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1302]&~m[1358]&m[1359]&m[1361]&~m[1362])|(~m[1302]&m[1358]&~m[1359]&~m[1361]&m[1362])|(~m[1302]&~m[1358]&m[1359]&~m[1361]&m[1362])|(m[1302]&m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1302]&m[1358]&m[1359]&m[1361]&m[1362]))&UnbiasedRNG[345])|((m[1302]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(~m[1302]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1302]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1302]&m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1302]&~m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1302]&~m[1358]&~m[1359]&m[1361]&m[1362])|(m[1302]&~m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1302]&m[1358]&~m[1359]&m[1361]&m[1362])|(m[1302]&m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1302]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1302]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1302]&m[1358]&m[1359]&m[1361]&m[1362]))):InitCond[984];
    m[1365] = run?((((m[1307]&~m[1363]&~m[1364]&~m[1366]&~m[1367])|(~m[1307]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1307]&m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1307]&~m[1363]&m[1364]&m[1366]&~m[1367])|(~m[1307]&m[1363]&~m[1364]&~m[1366]&m[1367])|(~m[1307]&~m[1363]&m[1364]&~m[1366]&m[1367])|(m[1307]&m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1307]&m[1363]&m[1364]&m[1366]&m[1367]))&UnbiasedRNG[346])|((m[1307]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(~m[1307]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1307]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1307]&m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1307]&~m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1307]&~m[1363]&~m[1364]&m[1366]&m[1367])|(m[1307]&~m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1307]&m[1363]&~m[1364]&m[1366]&m[1367])|(m[1307]&m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1307]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1307]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1307]&m[1363]&m[1364]&m[1366]&m[1367]))):InitCond[985];
    m[1370] = run?((((m[1312]&~m[1368]&~m[1369]&~m[1371]&~m[1372])|(~m[1312]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1312]&m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1312]&~m[1368]&m[1369]&m[1371]&~m[1372])|(~m[1312]&m[1368]&~m[1369]&~m[1371]&m[1372])|(~m[1312]&~m[1368]&m[1369]&~m[1371]&m[1372])|(m[1312]&m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1312]&m[1368]&m[1369]&m[1371]&m[1372]))&UnbiasedRNG[347])|((m[1312]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(~m[1312]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1312]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1312]&m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1312]&~m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1312]&~m[1368]&~m[1369]&m[1371]&m[1372])|(m[1312]&~m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1312]&m[1368]&~m[1369]&m[1371]&m[1372])|(m[1312]&m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1312]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1312]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1312]&m[1368]&m[1369]&m[1371]&m[1372]))):InitCond[986];
    m[1375] = run?((((m[1317]&~m[1373]&~m[1374]&~m[1376]&~m[1377])|(~m[1317]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1317]&m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1317]&~m[1373]&m[1374]&m[1376]&~m[1377])|(~m[1317]&m[1373]&~m[1374]&~m[1376]&m[1377])|(~m[1317]&~m[1373]&m[1374]&~m[1376]&m[1377])|(m[1317]&m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1317]&m[1373]&m[1374]&m[1376]&m[1377]))&UnbiasedRNG[348])|((m[1317]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(~m[1317]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1317]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1317]&m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1317]&~m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1317]&~m[1373]&~m[1374]&m[1376]&m[1377])|(m[1317]&~m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1317]&m[1373]&~m[1374]&m[1376]&m[1377])|(m[1317]&m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1317]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1317]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1317]&m[1373]&m[1374]&m[1376]&m[1377]))):InitCond[987];
    m[1385] = run?((((m[1322]&~m[1383]&~m[1384]&~m[1386]&~m[1387])|(~m[1322]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1322]&m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1322]&~m[1383]&m[1384]&m[1386]&~m[1387])|(~m[1322]&m[1383]&~m[1384]&~m[1386]&m[1387])|(~m[1322]&~m[1383]&m[1384]&~m[1386]&m[1387])|(m[1322]&m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1322]&m[1383]&m[1384]&m[1386]&m[1387]))&UnbiasedRNG[349])|((m[1322]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(~m[1322]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1322]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1322]&m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1322]&~m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1322]&~m[1383]&~m[1384]&m[1386]&m[1387])|(m[1322]&~m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1322]&m[1383]&~m[1384]&m[1386]&m[1387])|(m[1322]&m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1322]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1322]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1322]&m[1383]&m[1384]&m[1386]&m[1387]))):InitCond[988];
    m[1390] = run?((((m[1327]&~m[1388]&~m[1389]&~m[1391]&~m[1392])|(~m[1327]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1327]&m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1327]&~m[1388]&m[1389]&m[1391]&~m[1392])|(~m[1327]&m[1388]&~m[1389]&~m[1391]&m[1392])|(~m[1327]&~m[1388]&m[1389]&~m[1391]&m[1392])|(m[1327]&m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1327]&m[1388]&m[1389]&m[1391]&m[1392]))&UnbiasedRNG[350])|((m[1327]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(~m[1327]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1327]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1327]&m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1327]&~m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1327]&~m[1388]&~m[1389]&m[1391]&m[1392])|(m[1327]&~m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1327]&m[1388]&~m[1389]&m[1391]&m[1392])|(m[1327]&m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1327]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1327]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1327]&m[1388]&m[1389]&m[1391]&m[1392]))):InitCond[989];
    m[1395] = run?((((m[1332]&~m[1393]&~m[1394]&~m[1396]&~m[1397])|(~m[1332]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1332]&m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1332]&~m[1393]&m[1394]&m[1396]&~m[1397])|(~m[1332]&m[1393]&~m[1394]&~m[1396]&m[1397])|(~m[1332]&~m[1393]&m[1394]&~m[1396]&m[1397])|(m[1332]&m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1332]&m[1393]&m[1394]&m[1396]&m[1397]))&UnbiasedRNG[351])|((m[1332]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(~m[1332]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1332]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1332]&m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1332]&~m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1332]&~m[1393]&~m[1394]&m[1396]&m[1397])|(m[1332]&~m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1332]&m[1393]&~m[1394]&m[1396]&m[1397])|(m[1332]&m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1332]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1332]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1332]&m[1393]&m[1394]&m[1396]&m[1397]))):InitCond[990];
    m[1400] = run?((((m[1337]&~m[1398]&~m[1399]&~m[1401]&~m[1402])|(~m[1337]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1337]&m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1337]&~m[1398]&m[1399]&m[1401]&~m[1402])|(~m[1337]&m[1398]&~m[1399]&~m[1401]&m[1402])|(~m[1337]&~m[1398]&m[1399]&~m[1401]&m[1402])|(m[1337]&m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1337]&m[1398]&m[1399]&m[1401]&m[1402]))&UnbiasedRNG[352])|((m[1337]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(~m[1337]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1337]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1337]&m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1337]&~m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1337]&~m[1398]&~m[1399]&m[1401]&m[1402])|(m[1337]&~m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1337]&m[1398]&~m[1399]&m[1401]&m[1402])|(m[1337]&m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1337]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1337]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1337]&m[1398]&m[1399]&m[1401]&m[1402]))):InitCond[991];
    m[1405] = run?((((m[1342]&~m[1403]&~m[1404]&~m[1406]&~m[1407])|(~m[1342]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1342]&m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1342]&~m[1403]&m[1404]&m[1406]&~m[1407])|(~m[1342]&m[1403]&~m[1404]&~m[1406]&m[1407])|(~m[1342]&~m[1403]&m[1404]&~m[1406]&m[1407])|(m[1342]&m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1342]&m[1403]&m[1404]&m[1406]&m[1407]))&UnbiasedRNG[353])|((m[1342]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(~m[1342]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1342]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1342]&m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1342]&~m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1342]&~m[1403]&~m[1404]&m[1406]&m[1407])|(m[1342]&~m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1342]&m[1403]&~m[1404]&m[1406]&m[1407])|(m[1342]&m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1342]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1342]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1342]&m[1403]&m[1404]&m[1406]&m[1407]))):InitCond[992];
    m[1410] = run?((((m[1347]&~m[1408]&~m[1409]&~m[1411]&~m[1412])|(~m[1347]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1347]&m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1347]&~m[1408]&m[1409]&m[1411]&~m[1412])|(~m[1347]&m[1408]&~m[1409]&~m[1411]&m[1412])|(~m[1347]&~m[1408]&m[1409]&~m[1411]&m[1412])|(m[1347]&m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1347]&m[1408]&m[1409]&m[1411]&m[1412]))&UnbiasedRNG[354])|((m[1347]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(~m[1347]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1347]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1347]&m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1347]&~m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1347]&~m[1408]&~m[1409]&m[1411]&m[1412])|(m[1347]&~m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1347]&m[1408]&~m[1409]&m[1411]&m[1412])|(m[1347]&m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1347]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1347]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1347]&m[1408]&m[1409]&m[1411]&m[1412]))):InitCond[993];
    m[1415] = run?((((m[1352]&~m[1413]&~m[1414]&~m[1416]&~m[1417])|(~m[1352]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1352]&m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1352]&~m[1413]&m[1414]&m[1416]&~m[1417])|(~m[1352]&m[1413]&~m[1414]&~m[1416]&m[1417])|(~m[1352]&~m[1413]&m[1414]&~m[1416]&m[1417])|(m[1352]&m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1352]&m[1413]&m[1414]&m[1416]&m[1417]))&UnbiasedRNG[355])|((m[1352]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(~m[1352]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1352]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1352]&m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1352]&~m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1352]&~m[1413]&~m[1414]&m[1416]&m[1417])|(m[1352]&~m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1352]&m[1413]&~m[1414]&m[1416]&m[1417])|(m[1352]&m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1352]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1352]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1352]&m[1413]&m[1414]&m[1416]&m[1417]))):InitCond[994];
    m[1420] = run?((((m[1357]&~m[1418]&~m[1419]&~m[1421]&~m[1422])|(~m[1357]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1357]&m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1357]&~m[1418]&m[1419]&m[1421]&~m[1422])|(~m[1357]&m[1418]&~m[1419]&~m[1421]&m[1422])|(~m[1357]&~m[1418]&m[1419]&~m[1421]&m[1422])|(m[1357]&m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1357]&m[1418]&m[1419]&m[1421]&m[1422]))&UnbiasedRNG[356])|((m[1357]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(~m[1357]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1357]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1357]&m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1357]&~m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1357]&~m[1418]&~m[1419]&m[1421]&m[1422])|(m[1357]&~m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1357]&m[1418]&~m[1419]&m[1421]&m[1422])|(m[1357]&m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1357]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1357]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1357]&m[1418]&m[1419]&m[1421]&m[1422]))):InitCond[995];
    m[1425] = run?((((m[1362]&~m[1423]&~m[1424]&~m[1426]&~m[1427])|(~m[1362]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1362]&m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1362]&~m[1423]&m[1424]&m[1426]&~m[1427])|(~m[1362]&m[1423]&~m[1424]&~m[1426]&m[1427])|(~m[1362]&~m[1423]&m[1424]&~m[1426]&m[1427])|(m[1362]&m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1362]&m[1423]&m[1424]&m[1426]&m[1427]))&UnbiasedRNG[357])|((m[1362]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(~m[1362]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1362]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1362]&m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1362]&~m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1362]&~m[1423]&~m[1424]&m[1426]&m[1427])|(m[1362]&~m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1362]&m[1423]&~m[1424]&m[1426]&m[1427])|(m[1362]&m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1362]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1362]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1362]&m[1423]&m[1424]&m[1426]&m[1427]))):InitCond[996];
    m[1430] = run?((((m[1367]&~m[1428]&~m[1429]&~m[1431]&~m[1432])|(~m[1367]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1367]&m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1367]&~m[1428]&m[1429]&m[1431]&~m[1432])|(~m[1367]&m[1428]&~m[1429]&~m[1431]&m[1432])|(~m[1367]&~m[1428]&m[1429]&~m[1431]&m[1432])|(m[1367]&m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1367]&m[1428]&m[1429]&m[1431]&m[1432]))&UnbiasedRNG[358])|((m[1367]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(~m[1367]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1367]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1367]&m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1367]&~m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1367]&~m[1428]&~m[1429]&m[1431]&m[1432])|(m[1367]&~m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1367]&m[1428]&~m[1429]&m[1431]&m[1432])|(m[1367]&m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1367]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1367]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1367]&m[1428]&m[1429]&m[1431]&m[1432]))):InitCond[997];
    m[1435] = run?((((m[1372]&~m[1433]&~m[1434]&~m[1436]&~m[1437])|(~m[1372]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1372]&m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1372]&~m[1433]&m[1434]&m[1436]&~m[1437])|(~m[1372]&m[1433]&~m[1434]&~m[1436]&m[1437])|(~m[1372]&~m[1433]&m[1434]&~m[1436]&m[1437])|(m[1372]&m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1372]&m[1433]&m[1434]&m[1436]&m[1437]))&UnbiasedRNG[359])|((m[1372]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(~m[1372]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1372]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1372]&m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1372]&~m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1372]&~m[1433]&~m[1434]&m[1436]&m[1437])|(m[1372]&~m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1372]&m[1433]&~m[1434]&m[1436]&m[1437])|(m[1372]&m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1372]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1372]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1372]&m[1433]&m[1434]&m[1436]&m[1437]))):InitCond[998];
    m[1440] = run?((((m[1377]&~m[1438]&~m[1439]&~m[1441]&~m[1442])|(~m[1377]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1377]&m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1377]&~m[1438]&m[1439]&m[1441]&~m[1442])|(~m[1377]&m[1438]&~m[1439]&~m[1441]&m[1442])|(~m[1377]&~m[1438]&m[1439]&~m[1441]&m[1442])|(m[1377]&m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1377]&m[1438]&m[1439]&m[1441]&m[1442]))&UnbiasedRNG[360])|((m[1377]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(~m[1377]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1377]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1377]&m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1377]&~m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1377]&~m[1438]&~m[1439]&m[1441]&m[1442])|(m[1377]&~m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1377]&m[1438]&~m[1439]&m[1441]&m[1442])|(m[1377]&m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1377]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1377]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1377]&m[1438]&m[1439]&m[1441]&m[1442]))):InitCond[999];
    m[1445] = run?((((m[1382]&~m[1443]&~m[1444]&~m[1446]&~m[1447])|(~m[1382]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1382]&m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1382]&~m[1443]&m[1444]&m[1446]&~m[1447])|(~m[1382]&m[1443]&~m[1444]&~m[1446]&m[1447])|(~m[1382]&~m[1443]&m[1444]&~m[1446]&m[1447])|(m[1382]&m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1382]&m[1443]&m[1444]&m[1446]&m[1447]))&UnbiasedRNG[361])|((m[1382]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(~m[1382]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1382]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1382]&m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1382]&~m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1382]&~m[1443]&~m[1444]&m[1446]&m[1447])|(m[1382]&~m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1382]&m[1443]&~m[1444]&m[1446]&m[1447])|(m[1382]&m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1382]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1382]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1382]&m[1443]&m[1444]&m[1446]&m[1447]))):InitCond[1000];
    m[1455] = run?((((m[1387]&~m[1453]&~m[1454]&~m[1456]&~m[1457])|(~m[1387]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1387]&m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1387]&~m[1453]&m[1454]&m[1456]&~m[1457])|(~m[1387]&m[1453]&~m[1454]&~m[1456]&m[1457])|(~m[1387]&~m[1453]&m[1454]&~m[1456]&m[1457])|(m[1387]&m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1387]&m[1453]&m[1454]&m[1456]&m[1457]))&UnbiasedRNG[362])|((m[1387]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(~m[1387]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1387]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1387]&m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1387]&~m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1387]&~m[1453]&~m[1454]&m[1456]&m[1457])|(m[1387]&~m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1387]&m[1453]&~m[1454]&m[1456]&m[1457])|(m[1387]&m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1387]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1387]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1387]&m[1453]&m[1454]&m[1456]&m[1457]))):InitCond[1001];
    m[1460] = run?((((m[1392]&~m[1458]&~m[1459]&~m[1461]&~m[1462])|(~m[1392]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1392]&m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1392]&~m[1458]&m[1459]&m[1461]&~m[1462])|(~m[1392]&m[1458]&~m[1459]&~m[1461]&m[1462])|(~m[1392]&~m[1458]&m[1459]&~m[1461]&m[1462])|(m[1392]&m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1392]&m[1458]&m[1459]&m[1461]&m[1462]))&UnbiasedRNG[363])|((m[1392]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(~m[1392]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1392]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1392]&m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1392]&~m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1392]&~m[1458]&~m[1459]&m[1461]&m[1462])|(m[1392]&~m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1392]&m[1458]&~m[1459]&m[1461]&m[1462])|(m[1392]&m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1392]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1392]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1392]&m[1458]&m[1459]&m[1461]&m[1462]))):InitCond[1002];
    m[1465] = run?((((m[1397]&~m[1463]&~m[1464]&~m[1466]&~m[1467])|(~m[1397]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1397]&m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1397]&~m[1463]&m[1464]&m[1466]&~m[1467])|(~m[1397]&m[1463]&~m[1464]&~m[1466]&m[1467])|(~m[1397]&~m[1463]&m[1464]&~m[1466]&m[1467])|(m[1397]&m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1397]&m[1463]&m[1464]&m[1466]&m[1467]))&UnbiasedRNG[364])|((m[1397]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(~m[1397]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1397]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1397]&m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1397]&~m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1397]&~m[1463]&~m[1464]&m[1466]&m[1467])|(m[1397]&~m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1397]&m[1463]&~m[1464]&m[1466]&m[1467])|(m[1397]&m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1397]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1397]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1397]&m[1463]&m[1464]&m[1466]&m[1467]))):InitCond[1003];
    m[1470] = run?((((m[1402]&~m[1468]&~m[1469]&~m[1471]&~m[1472])|(~m[1402]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1402]&m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1402]&~m[1468]&m[1469]&m[1471]&~m[1472])|(~m[1402]&m[1468]&~m[1469]&~m[1471]&m[1472])|(~m[1402]&~m[1468]&m[1469]&~m[1471]&m[1472])|(m[1402]&m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1402]&m[1468]&m[1469]&m[1471]&m[1472]))&UnbiasedRNG[365])|((m[1402]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(~m[1402]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1402]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1402]&m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1402]&~m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1402]&~m[1468]&~m[1469]&m[1471]&m[1472])|(m[1402]&~m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1402]&m[1468]&~m[1469]&m[1471]&m[1472])|(m[1402]&m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1402]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1402]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1402]&m[1468]&m[1469]&m[1471]&m[1472]))):InitCond[1004];
    m[1475] = run?((((m[1407]&~m[1473]&~m[1474]&~m[1476]&~m[1477])|(~m[1407]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1407]&m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1407]&~m[1473]&m[1474]&m[1476]&~m[1477])|(~m[1407]&m[1473]&~m[1474]&~m[1476]&m[1477])|(~m[1407]&~m[1473]&m[1474]&~m[1476]&m[1477])|(m[1407]&m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1407]&m[1473]&m[1474]&m[1476]&m[1477]))&UnbiasedRNG[366])|((m[1407]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(~m[1407]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1407]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1407]&m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1407]&~m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1407]&~m[1473]&~m[1474]&m[1476]&m[1477])|(m[1407]&~m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1407]&m[1473]&~m[1474]&m[1476]&m[1477])|(m[1407]&m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1407]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1407]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1407]&m[1473]&m[1474]&m[1476]&m[1477]))):InitCond[1005];
    m[1480] = run?((((m[1412]&~m[1478]&~m[1479]&~m[1481]&~m[1482])|(~m[1412]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1412]&m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1412]&~m[1478]&m[1479]&m[1481]&~m[1482])|(~m[1412]&m[1478]&~m[1479]&~m[1481]&m[1482])|(~m[1412]&~m[1478]&m[1479]&~m[1481]&m[1482])|(m[1412]&m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1412]&m[1478]&m[1479]&m[1481]&m[1482]))&UnbiasedRNG[367])|((m[1412]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(~m[1412]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1412]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1412]&m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1412]&~m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1412]&~m[1478]&~m[1479]&m[1481]&m[1482])|(m[1412]&~m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1412]&m[1478]&~m[1479]&m[1481]&m[1482])|(m[1412]&m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1412]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1412]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1412]&m[1478]&m[1479]&m[1481]&m[1482]))):InitCond[1006];
    m[1485] = run?((((m[1417]&~m[1483]&~m[1484]&~m[1486]&~m[1487])|(~m[1417]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1417]&m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1417]&~m[1483]&m[1484]&m[1486]&~m[1487])|(~m[1417]&m[1483]&~m[1484]&~m[1486]&m[1487])|(~m[1417]&~m[1483]&m[1484]&~m[1486]&m[1487])|(m[1417]&m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1417]&m[1483]&m[1484]&m[1486]&m[1487]))&UnbiasedRNG[368])|((m[1417]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(~m[1417]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1417]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1417]&m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1417]&~m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1417]&~m[1483]&~m[1484]&m[1486]&m[1487])|(m[1417]&~m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1417]&m[1483]&~m[1484]&m[1486]&m[1487])|(m[1417]&m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1417]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1417]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1417]&m[1483]&m[1484]&m[1486]&m[1487]))):InitCond[1007];
    m[1490] = run?((((m[1422]&~m[1488]&~m[1489]&~m[1491]&~m[1492])|(~m[1422]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1422]&m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1422]&~m[1488]&m[1489]&m[1491]&~m[1492])|(~m[1422]&m[1488]&~m[1489]&~m[1491]&m[1492])|(~m[1422]&~m[1488]&m[1489]&~m[1491]&m[1492])|(m[1422]&m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1422]&m[1488]&m[1489]&m[1491]&m[1492]))&UnbiasedRNG[369])|((m[1422]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(~m[1422]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1422]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1422]&m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1422]&~m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1422]&~m[1488]&~m[1489]&m[1491]&m[1492])|(m[1422]&~m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1422]&m[1488]&~m[1489]&m[1491]&m[1492])|(m[1422]&m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1422]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1422]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1422]&m[1488]&m[1489]&m[1491]&m[1492]))):InitCond[1008];
    m[1495] = run?((((m[1427]&~m[1493]&~m[1494]&~m[1496]&~m[1497])|(~m[1427]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1427]&m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1427]&~m[1493]&m[1494]&m[1496]&~m[1497])|(~m[1427]&m[1493]&~m[1494]&~m[1496]&m[1497])|(~m[1427]&~m[1493]&m[1494]&~m[1496]&m[1497])|(m[1427]&m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1427]&m[1493]&m[1494]&m[1496]&m[1497]))&UnbiasedRNG[370])|((m[1427]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(~m[1427]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1427]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1427]&m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1427]&~m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1427]&~m[1493]&~m[1494]&m[1496]&m[1497])|(m[1427]&~m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1427]&m[1493]&~m[1494]&m[1496]&m[1497])|(m[1427]&m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1427]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1427]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1427]&m[1493]&m[1494]&m[1496]&m[1497]))):InitCond[1009];
    m[1500] = run?((((m[1432]&~m[1498]&~m[1499]&~m[1501]&~m[1502])|(~m[1432]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1432]&m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1432]&~m[1498]&m[1499]&m[1501]&~m[1502])|(~m[1432]&m[1498]&~m[1499]&~m[1501]&m[1502])|(~m[1432]&~m[1498]&m[1499]&~m[1501]&m[1502])|(m[1432]&m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1432]&m[1498]&m[1499]&m[1501]&m[1502]))&UnbiasedRNG[371])|((m[1432]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(~m[1432]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1432]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1432]&m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1432]&~m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1432]&~m[1498]&~m[1499]&m[1501]&m[1502])|(m[1432]&~m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1432]&m[1498]&~m[1499]&m[1501]&m[1502])|(m[1432]&m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1432]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1432]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1432]&m[1498]&m[1499]&m[1501]&m[1502]))):InitCond[1010];
    m[1505] = run?((((m[1437]&~m[1503]&~m[1504]&~m[1506]&~m[1507])|(~m[1437]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1437]&m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1437]&~m[1503]&m[1504]&m[1506]&~m[1507])|(~m[1437]&m[1503]&~m[1504]&~m[1506]&m[1507])|(~m[1437]&~m[1503]&m[1504]&~m[1506]&m[1507])|(m[1437]&m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1437]&m[1503]&m[1504]&m[1506]&m[1507]))&UnbiasedRNG[372])|((m[1437]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(~m[1437]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1437]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1437]&m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1437]&~m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1437]&~m[1503]&~m[1504]&m[1506]&m[1507])|(m[1437]&~m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1437]&m[1503]&~m[1504]&m[1506]&m[1507])|(m[1437]&m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1437]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1437]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1437]&m[1503]&m[1504]&m[1506]&m[1507]))):InitCond[1011];
    m[1510] = run?((((m[1442]&~m[1508]&~m[1509]&~m[1511]&~m[1512])|(~m[1442]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1442]&m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1442]&~m[1508]&m[1509]&m[1511]&~m[1512])|(~m[1442]&m[1508]&~m[1509]&~m[1511]&m[1512])|(~m[1442]&~m[1508]&m[1509]&~m[1511]&m[1512])|(m[1442]&m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1442]&m[1508]&m[1509]&m[1511]&m[1512]))&UnbiasedRNG[373])|((m[1442]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(~m[1442]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1442]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1442]&m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1442]&~m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1442]&~m[1508]&~m[1509]&m[1511]&m[1512])|(m[1442]&~m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1442]&m[1508]&~m[1509]&m[1511]&m[1512])|(m[1442]&m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1442]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1442]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1442]&m[1508]&m[1509]&m[1511]&m[1512]))):InitCond[1012];
    m[1515] = run?((((m[1447]&~m[1513]&~m[1514]&~m[1516]&~m[1517])|(~m[1447]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1447]&m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1447]&~m[1513]&m[1514]&m[1516]&~m[1517])|(~m[1447]&m[1513]&~m[1514]&~m[1516]&m[1517])|(~m[1447]&~m[1513]&m[1514]&~m[1516]&m[1517])|(m[1447]&m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1447]&m[1513]&m[1514]&m[1516]&m[1517]))&UnbiasedRNG[374])|((m[1447]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(~m[1447]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1447]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1447]&m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1447]&~m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1447]&~m[1513]&~m[1514]&m[1516]&m[1517])|(m[1447]&~m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1447]&m[1513]&~m[1514]&m[1516]&m[1517])|(m[1447]&m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1447]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1447]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1447]&m[1513]&m[1514]&m[1516]&m[1517]))):InitCond[1013];
    m[1520] = run?((((m[1452]&~m[1518]&~m[1519]&~m[1521]&~m[1522])|(~m[1452]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1452]&m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1452]&~m[1518]&m[1519]&m[1521]&~m[1522])|(~m[1452]&m[1518]&~m[1519]&~m[1521]&m[1522])|(~m[1452]&~m[1518]&m[1519]&~m[1521]&m[1522])|(m[1452]&m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1452]&m[1518]&m[1519]&m[1521]&m[1522]))&UnbiasedRNG[375])|((m[1452]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(~m[1452]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1452]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1452]&m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1452]&~m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1452]&~m[1518]&~m[1519]&m[1521]&m[1522])|(m[1452]&~m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1452]&m[1518]&~m[1519]&m[1521]&m[1522])|(m[1452]&m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1452]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1452]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1452]&m[1518]&m[1519]&m[1521]&m[1522]))):InitCond[1014];
    m[1530] = run?((((m[1457]&~m[1528]&~m[1529]&~m[1531]&~m[1532])|(~m[1457]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1457]&m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1457]&~m[1528]&m[1529]&m[1531]&~m[1532])|(~m[1457]&m[1528]&~m[1529]&~m[1531]&m[1532])|(~m[1457]&~m[1528]&m[1529]&~m[1531]&m[1532])|(m[1457]&m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1457]&m[1528]&m[1529]&m[1531]&m[1532]))&UnbiasedRNG[376])|((m[1457]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(~m[1457]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1457]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1457]&m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1457]&~m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1457]&~m[1528]&~m[1529]&m[1531]&m[1532])|(m[1457]&~m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1457]&m[1528]&~m[1529]&m[1531]&m[1532])|(m[1457]&m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1457]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1457]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1457]&m[1528]&m[1529]&m[1531]&m[1532]))):InitCond[1015];
    m[1535] = run?((((m[1462]&~m[1533]&~m[1534]&~m[1536]&~m[1537])|(~m[1462]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1462]&m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1462]&~m[1533]&m[1534]&m[1536]&~m[1537])|(~m[1462]&m[1533]&~m[1534]&~m[1536]&m[1537])|(~m[1462]&~m[1533]&m[1534]&~m[1536]&m[1537])|(m[1462]&m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1462]&m[1533]&m[1534]&m[1536]&m[1537]))&UnbiasedRNG[377])|((m[1462]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(~m[1462]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1462]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1462]&m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1462]&~m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1462]&~m[1533]&~m[1534]&m[1536]&m[1537])|(m[1462]&~m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1462]&m[1533]&~m[1534]&m[1536]&m[1537])|(m[1462]&m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1462]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1462]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1462]&m[1533]&m[1534]&m[1536]&m[1537]))):InitCond[1016];
    m[1540] = run?((((m[1467]&~m[1538]&~m[1539]&~m[1541]&~m[1542])|(~m[1467]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1467]&m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1467]&~m[1538]&m[1539]&m[1541]&~m[1542])|(~m[1467]&m[1538]&~m[1539]&~m[1541]&m[1542])|(~m[1467]&~m[1538]&m[1539]&~m[1541]&m[1542])|(m[1467]&m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1467]&m[1538]&m[1539]&m[1541]&m[1542]))&UnbiasedRNG[378])|((m[1467]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(~m[1467]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1467]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1467]&m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1467]&~m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1467]&~m[1538]&~m[1539]&m[1541]&m[1542])|(m[1467]&~m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1467]&m[1538]&~m[1539]&m[1541]&m[1542])|(m[1467]&m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1467]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1467]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1467]&m[1538]&m[1539]&m[1541]&m[1542]))):InitCond[1017];
    m[1545] = run?((((m[1472]&~m[1543]&~m[1544]&~m[1546]&~m[1547])|(~m[1472]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1472]&m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1472]&~m[1543]&m[1544]&m[1546]&~m[1547])|(~m[1472]&m[1543]&~m[1544]&~m[1546]&m[1547])|(~m[1472]&~m[1543]&m[1544]&~m[1546]&m[1547])|(m[1472]&m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1472]&m[1543]&m[1544]&m[1546]&m[1547]))&UnbiasedRNG[379])|((m[1472]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(~m[1472]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1472]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1472]&m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1472]&~m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1472]&~m[1543]&~m[1544]&m[1546]&m[1547])|(m[1472]&~m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1472]&m[1543]&~m[1544]&m[1546]&m[1547])|(m[1472]&m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1472]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1472]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1472]&m[1543]&m[1544]&m[1546]&m[1547]))):InitCond[1018];
    m[1550] = run?((((m[1477]&~m[1548]&~m[1549]&~m[1551]&~m[1552])|(~m[1477]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1477]&m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1477]&~m[1548]&m[1549]&m[1551]&~m[1552])|(~m[1477]&m[1548]&~m[1549]&~m[1551]&m[1552])|(~m[1477]&~m[1548]&m[1549]&~m[1551]&m[1552])|(m[1477]&m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1477]&m[1548]&m[1549]&m[1551]&m[1552]))&UnbiasedRNG[380])|((m[1477]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(~m[1477]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1477]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1477]&m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1477]&~m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1477]&~m[1548]&~m[1549]&m[1551]&m[1552])|(m[1477]&~m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1477]&m[1548]&~m[1549]&m[1551]&m[1552])|(m[1477]&m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1477]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1477]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1477]&m[1548]&m[1549]&m[1551]&m[1552]))):InitCond[1019];
    m[1555] = run?((((m[1482]&~m[1553]&~m[1554]&~m[1556]&~m[1557])|(~m[1482]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1482]&m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1482]&~m[1553]&m[1554]&m[1556]&~m[1557])|(~m[1482]&m[1553]&~m[1554]&~m[1556]&m[1557])|(~m[1482]&~m[1553]&m[1554]&~m[1556]&m[1557])|(m[1482]&m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1482]&m[1553]&m[1554]&m[1556]&m[1557]))&UnbiasedRNG[381])|((m[1482]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(~m[1482]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1482]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1482]&m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1482]&~m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1482]&~m[1553]&~m[1554]&m[1556]&m[1557])|(m[1482]&~m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1482]&m[1553]&~m[1554]&m[1556]&m[1557])|(m[1482]&m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1482]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1482]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1482]&m[1553]&m[1554]&m[1556]&m[1557]))):InitCond[1020];
    m[1560] = run?((((m[1487]&~m[1558]&~m[1559]&~m[1561]&~m[1562])|(~m[1487]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1487]&m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1487]&~m[1558]&m[1559]&m[1561]&~m[1562])|(~m[1487]&m[1558]&~m[1559]&~m[1561]&m[1562])|(~m[1487]&~m[1558]&m[1559]&~m[1561]&m[1562])|(m[1487]&m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1487]&m[1558]&m[1559]&m[1561]&m[1562]))&UnbiasedRNG[382])|((m[1487]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(~m[1487]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1487]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1487]&m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1487]&~m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1487]&~m[1558]&~m[1559]&m[1561]&m[1562])|(m[1487]&~m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1487]&m[1558]&~m[1559]&m[1561]&m[1562])|(m[1487]&m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1487]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1487]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1487]&m[1558]&m[1559]&m[1561]&m[1562]))):InitCond[1021];
    m[1565] = run?((((m[1492]&~m[1563]&~m[1564]&~m[1566]&~m[1567])|(~m[1492]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1492]&m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1492]&~m[1563]&m[1564]&m[1566]&~m[1567])|(~m[1492]&m[1563]&~m[1564]&~m[1566]&m[1567])|(~m[1492]&~m[1563]&m[1564]&~m[1566]&m[1567])|(m[1492]&m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1492]&m[1563]&m[1564]&m[1566]&m[1567]))&UnbiasedRNG[383])|((m[1492]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(~m[1492]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1492]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1492]&m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1492]&~m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1492]&~m[1563]&~m[1564]&m[1566]&m[1567])|(m[1492]&~m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1492]&m[1563]&~m[1564]&m[1566]&m[1567])|(m[1492]&m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1492]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1492]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1492]&m[1563]&m[1564]&m[1566]&m[1567]))):InitCond[1022];
    m[1570] = run?((((m[1497]&~m[1568]&~m[1569]&~m[1571]&~m[1572])|(~m[1497]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1497]&m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1497]&~m[1568]&m[1569]&m[1571]&~m[1572])|(~m[1497]&m[1568]&~m[1569]&~m[1571]&m[1572])|(~m[1497]&~m[1568]&m[1569]&~m[1571]&m[1572])|(m[1497]&m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1497]&m[1568]&m[1569]&m[1571]&m[1572]))&UnbiasedRNG[384])|((m[1497]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(~m[1497]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1497]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1497]&m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1497]&~m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1497]&~m[1568]&~m[1569]&m[1571]&m[1572])|(m[1497]&~m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1497]&m[1568]&~m[1569]&m[1571]&m[1572])|(m[1497]&m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1497]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1497]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1497]&m[1568]&m[1569]&m[1571]&m[1572]))):InitCond[1023];
    m[1575] = run?((((m[1502]&~m[1573]&~m[1574]&~m[1576]&~m[1577])|(~m[1502]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1502]&m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1502]&~m[1573]&m[1574]&m[1576]&~m[1577])|(~m[1502]&m[1573]&~m[1574]&~m[1576]&m[1577])|(~m[1502]&~m[1573]&m[1574]&~m[1576]&m[1577])|(m[1502]&m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1502]&m[1573]&m[1574]&m[1576]&m[1577]))&UnbiasedRNG[385])|((m[1502]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(~m[1502]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1502]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1502]&m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1502]&~m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1502]&~m[1573]&~m[1574]&m[1576]&m[1577])|(m[1502]&~m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1502]&m[1573]&~m[1574]&m[1576]&m[1577])|(m[1502]&m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1502]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1502]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1502]&m[1573]&m[1574]&m[1576]&m[1577]))):InitCond[1024];
    m[1580] = run?((((m[1507]&~m[1578]&~m[1579]&~m[1581]&~m[1582])|(~m[1507]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1507]&m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1507]&~m[1578]&m[1579]&m[1581]&~m[1582])|(~m[1507]&m[1578]&~m[1579]&~m[1581]&m[1582])|(~m[1507]&~m[1578]&m[1579]&~m[1581]&m[1582])|(m[1507]&m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1507]&m[1578]&m[1579]&m[1581]&m[1582]))&UnbiasedRNG[386])|((m[1507]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(~m[1507]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1507]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1507]&m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1507]&~m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1507]&~m[1578]&~m[1579]&m[1581]&m[1582])|(m[1507]&~m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1507]&m[1578]&~m[1579]&m[1581]&m[1582])|(m[1507]&m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1507]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1507]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1507]&m[1578]&m[1579]&m[1581]&m[1582]))):InitCond[1025];
    m[1585] = run?((((m[1512]&~m[1583]&~m[1584]&~m[1586]&~m[1587])|(~m[1512]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1512]&m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1512]&~m[1583]&m[1584]&m[1586]&~m[1587])|(~m[1512]&m[1583]&~m[1584]&~m[1586]&m[1587])|(~m[1512]&~m[1583]&m[1584]&~m[1586]&m[1587])|(m[1512]&m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1512]&m[1583]&m[1584]&m[1586]&m[1587]))&UnbiasedRNG[387])|((m[1512]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(~m[1512]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1512]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1512]&m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1512]&~m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1512]&~m[1583]&~m[1584]&m[1586]&m[1587])|(m[1512]&~m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1512]&m[1583]&~m[1584]&m[1586]&m[1587])|(m[1512]&m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1512]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1512]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1512]&m[1583]&m[1584]&m[1586]&m[1587]))):InitCond[1026];
    m[1590] = run?((((m[1517]&~m[1588]&~m[1589]&~m[1591]&~m[1592])|(~m[1517]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1517]&m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1517]&~m[1588]&m[1589]&m[1591]&~m[1592])|(~m[1517]&m[1588]&~m[1589]&~m[1591]&m[1592])|(~m[1517]&~m[1588]&m[1589]&~m[1591]&m[1592])|(m[1517]&m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1517]&m[1588]&m[1589]&m[1591]&m[1592]))&UnbiasedRNG[388])|((m[1517]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(~m[1517]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1517]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1517]&m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1517]&~m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1517]&~m[1588]&~m[1589]&m[1591]&m[1592])|(m[1517]&~m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1517]&m[1588]&~m[1589]&m[1591]&m[1592])|(m[1517]&m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1517]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1517]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1517]&m[1588]&m[1589]&m[1591]&m[1592]))):InitCond[1027];
    m[1595] = run?((((m[1522]&~m[1593]&~m[1594]&~m[1596]&~m[1597])|(~m[1522]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1522]&m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1522]&~m[1593]&m[1594]&m[1596]&~m[1597])|(~m[1522]&m[1593]&~m[1594]&~m[1596]&m[1597])|(~m[1522]&~m[1593]&m[1594]&~m[1596]&m[1597])|(m[1522]&m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1522]&m[1593]&m[1594]&m[1596]&m[1597]))&UnbiasedRNG[389])|((m[1522]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(~m[1522]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1522]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1522]&m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1522]&~m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1522]&~m[1593]&~m[1594]&m[1596]&m[1597])|(m[1522]&~m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1522]&m[1593]&~m[1594]&m[1596]&m[1597])|(m[1522]&m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1522]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1522]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1522]&m[1593]&m[1594]&m[1596]&m[1597]))):InitCond[1028];
    m[1600] = run?((((m[1527]&~m[1598]&~m[1599]&~m[1601]&~m[1602])|(~m[1527]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1527]&m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1527]&~m[1598]&m[1599]&m[1601]&~m[1602])|(~m[1527]&m[1598]&~m[1599]&~m[1601]&m[1602])|(~m[1527]&~m[1598]&m[1599]&~m[1601]&m[1602])|(m[1527]&m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1527]&m[1598]&m[1599]&m[1601]&m[1602]))&UnbiasedRNG[390])|((m[1527]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(~m[1527]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1527]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1527]&m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1527]&~m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1527]&~m[1598]&~m[1599]&m[1601]&m[1602])|(m[1527]&~m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1527]&m[1598]&~m[1599]&m[1601]&m[1602])|(m[1527]&m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1527]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1527]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1527]&m[1598]&m[1599]&m[1601]&m[1602]))):InitCond[1029];
    m[1605] = run?((((m[1537]&~m[1603]&~m[1604]&~m[1606]&~m[1607])|(~m[1537]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1537]&m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1537]&~m[1603]&m[1604]&m[1606]&~m[1607])|(~m[1537]&m[1603]&~m[1604]&~m[1606]&m[1607])|(~m[1537]&~m[1603]&m[1604]&~m[1606]&m[1607])|(m[1537]&m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1537]&m[1603]&m[1604]&m[1606]&m[1607]))&UnbiasedRNG[391])|((m[1537]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(~m[1537]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1537]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1537]&m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1537]&~m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1537]&~m[1603]&~m[1604]&m[1606]&m[1607])|(m[1537]&~m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1537]&m[1603]&~m[1604]&m[1606]&m[1607])|(m[1537]&m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1537]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1537]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1537]&m[1603]&m[1604]&m[1606]&m[1607]))):InitCond[1030];
    m[1610] = run?((((m[1542]&~m[1608]&~m[1609]&~m[1611]&~m[1612])|(~m[1542]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1542]&m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1542]&~m[1608]&m[1609]&m[1611]&~m[1612])|(~m[1542]&m[1608]&~m[1609]&~m[1611]&m[1612])|(~m[1542]&~m[1608]&m[1609]&~m[1611]&m[1612])|(m[1542]&m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1542]&m[1608]&m[1609]&m[1611]&m[1612]))&UnbiasedRNG[392])|((m[1542]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(~m[1542]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1542]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1542]&m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1542]&~m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1542]&~m[1608]&~m[1609]&m[1611]&m[1612])|(m[1542]&~m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1542]&m[1608]&~m[1609]&m[1611]&m[1612])|(m[1542]&m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1542]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1542]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1542]&m[1608]&m[1609]&m[1611]&m[1612]))):InitCond[1031];
    m[1615] = run?((((m[1547]&~m[1613]&~m[1614]&~m[1616]&~m[1617])|(~m[1547]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1547]&m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1547]&~m[1613]&m[1614]&m[1616]&~m[1617])|(~m[1547]&m[1613]&~m[1614]&~m[1616]&m[1617])|(~m[1547]&~m[1613]&m[1614]&~m[1616]&m[1617])|(m[1547]&m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1547]&m[1613]&m[1614]&m[1616]&m[1617]))&UnbiasedRNG[393])|((m[1547]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(~m[1547]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1547]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1547]&m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1547]&~m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1547]&~m[1613]&~m[1614]&m[1616]&m[1617])|(m[1547]&~m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1547]&m[1613]&~m[1614]&m[1616]&m[1617])|(m[1547]&m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1547]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1547]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1547]&m[1613]&m[1614]&m[1616]&m[1617]))):InitCond[1032];
    m[1620] = run?((((m[1552]&~m[1618]&~m[1619]&~m[1621]&~m[1622])|(~m[1552]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1552]&m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1552]&~m[1618]&m[1619]&m[1621]&~m[1622])|(~m[1552]&m[1618]&~m[1619]&~m[1621]&m[1622])|(~m[1552]&~m[1618]&m[1619]&~m[1621]&m[1622])|(m[1552]&m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1552]&m[1618]&m[1619]&m[1621]&m[1622]))&UnbiasedRNG[394])|((m[1552]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(~m[1552]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1552]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1552]&m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1552]&~m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1552]&~m[1618]&~m[1619]&m[1621]&m[1622])|(m[1552]&~m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1552]&m[1618]&~m[1619]&m[1621]&m[1622])|(m[1552]&m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1552]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1552]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1552]&m[1618]&m[1619]&m[1621]&m[1622]))):InitCond[1033];
    m[1625] = run?((((m[1557]&~m[1623]&~m[1624]&~m[1626]&~m[1627])|(~m[1557]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1557]&m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1557]&~m[1623]&m[1624]&m[1626]&~m[1627])|(~m[1557]&m[1623]&~m[1624]&~m[1626]&m[1627])|(~m[1557]&~m[1623]&m[1624]&~m[1626]&m[1627])|(m[1557]&m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1557]&m[1623]&m[1624]&m[1626]&m[1627]))&UnbiasedRNG[395])|((m[1557]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(~m[1557]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1557]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1557]&m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1557]&~m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1557]&~m[1623]&~m[1624]&m[1626]&m[1627])|(m[1557]&~m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1557]&m[1623]&~m[1624]&m[1626]&m[1627])|(m[1557]&m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1557]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1557]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1557]&m[1623]&m[1624]&m[1626]&m[1627]))):InitCond[1034];
    m[1630] = run?((((m[1562]&~m[1628]&~m[1629]&~m[1631]&~m[1632])|(~m[1562]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1562]&m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1562]&~m[1628]&m[1629]&m[1631]&~m[1632])|(~m[1562]&m[1628]&~m[1629]&~m[1631]&m[1632])|(~m[1562]&~m[1628]&m[1629]&~m[1631]&m[1632])|(m[1562]&m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1562]&m[1628]&m[1629]&m[1631]&m[1632]))&UnbiasedRNG[396])|((m[1562]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(~m[1562]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1562]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1562]&m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1562]&~m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1562]&~m[1628]&~m[1629]&m[1631]&m[1632])|(m[1562]&~m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1562]&m[1628]&~m[1629]&m[1631]&m[1632])|(m[1562]&m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1562]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1562]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1562]&m[1628]&m[1629]&m[1631]&m[1632]))):InitCond[1035];
    m[1635] = run?((((m[1567]&~m[1633]&~m[1634]&~m[1636]&~m[1637])|(~m[1567]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1567]&m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1567]&~m[1633]&m[1634]&m[1636]&~m[1637])|(~m[1567]&m[1633]&~m[1634]&~m[1636]&m[1637])|(~m[1567]&~m[1633]&m[1634]&~m[1636]&m[1637])|(m[1567]&m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1567]&m[1633]&m[1634]&m[1636]&m[1637]))&UnbiasedRNG[397])|((m[1567]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(~m[1567]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1567]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1567]&m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1567]&~m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1567]&~m[1633]&~m[1634]&m[1636]&m[1637])|(m[1567]&~m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1567]&m[1633]&~m[1634]&m[1636]&m[1637])|(m[1567]&m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1567]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1567]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1567]&m[1633]&m[1634]&m[1636]&m[1637]))):InitCond[1036];
    m[1640] = run?((((m[1572]&~m[1638]&~m[1639]&~m[1641]&~m[1642])|(~m[1572]&~m[1638]&~m[1639]&m[1641]&~m[1642])|(m[1572]&m[1638]&~m[1639]&m[1641]&~m[1642])|(m[1572]&~m[1638]&m[1639]&m[1641]&~m[1642])|(~m[1572]&m[1638]&~m[1639]&~m[1641]&m[1642])|(~m[1572]&~m[1638]&m[1639]&~m[1641]&m[1642])|(m[1572]&m[1638]&m[1639]&~m[1641]&m[1642])|(~m[1572]&m[1638]&m[1639]&m[1641]&m[1642]))&UnbiasedRNG[398])|((m[1572]&~m[1638]&~m[1639]&m[1641]&~m[1642])|(~m[1572]&~m[1638]&~m[1639]&~m[1641]&m[1642])|(m[1572]&~m[1638]&~m[1639]&~m[1641]&m[1642])|(m[1572]&m[1638]&~m[1639]&~m[1641]&m[1642])|(m[1572]&~m[1638]&m[1639]&~m[1641]&m[1642])|(~m[1572]&~m[1638]&~m[1639]&m[1641]&m[1642])|(m[1572]&~m[1638]&~m[1639]&m[1641]&m[1642])|(~m[1572]&m[1638]&~m[1639]&m[1641]&m[1642])|(m[1572]&m[1638]&~m[1639]&m[1641]&m[1642])|(~m[1572]&~m[1638]&m[1639]&m[1641]&m[1642])|(m[1572]&~m[1638]&m[1639]&m[1641]&m[1642])|(m[1572]&m[1638]&m[1639]&m[1641]&m[1642]))):InitCond[1037];
    m[1645] = run?((((m[1577]&~m[1643]&~m[1644]&~m[1646]&~m[1647])|(~m[1577]&~m[1643]&~m[1644]&m[1646]&~m[1647])|(m[1577]&m[1643]&~m[1644]&m[1646]&~m[1647])|(m[1577]&~m[1643]&m[1644]&m[1646]&~m[1647])|(~m[1577]&m[1643]&~m[1644]&~m[1646]&m[1647])|(~m[1577]&~m[1643]&m[1644]&~m[1646]&m[1647])|(m[1577]&m[1643]&m[1644]&~m[1646]&m[1647])|(~m[1577]&m[1643]&m[1644]&m[1646]&m[1647]))&UnbiasedRNG[399])|((m[1577]&~m[1643]&~m[1644]&m[1646]&~m[1647])|(~m[1577]&~m[1643]&~m[1644]&~m[1646]&m[1647])|(m[1577]&~m[1643]&~m[1644]&~m[1646]&m[1647])|(m[1577]&m[1643]&~m[1644]&~m[1646]&m[1647])|(m[1577]&~m[1643]&m[1644]&~m[1646]&m[1647])|(~m[1577]&~m[1643]&~m[1644]&m[1646]&m[1647])|(m[1577]&~m[1643]&~m[1644]&m[1646]&m[1647])|(~m[1577]&m[1643]&~m[1644]&m[1646]&m[1647])|(m[1577]&m[1643]&~m[1644]&m[1646]&m[1647])|(~m[1577]&~m[1643]&m[1644]&m[1646]&m[1647])|(m[1577]&~m[1643]&m[1644]&m[1646]&m[1647])|(m[1577]&m[1643]&m[1644]&m[1646]&m[1647]))):InitCond[1038];
    m[1650] = run?((((m[1582]&~m[1648]&~m[1649]&~m[1651]&~m[1652])|(~m[1582]&~m[1648]&~m[1649]&m[1651]&~m[1652])|(m[1582]&m[1648]&~m[1649]&m[1651]&~m[1652])|(m[1582]&~m[1648]&m[1649]&m[1651]&~m[1652])|(~m[1582]&m[1648]&~m[1649]&~m[1651]&m[1652])|(~m[1582]&~m[1648]&m[1649]&~m[1651]&m[1652])|(m[1582]&m[1648]&m[1649]&~m[1651]&m[1652])|(~m[1582]&m[1648]&m[1649]&m[1651]&m[1652]))&UnbiasedRNG[400])|((m[1582]&~m[1648]&~m[1649]&m[1651]&~m[1652])|(~m[1582]&~m[1648]&~m[1649]&~m[1651]&m[1652])|(m[1582]&~m[1648]&~m[1649]&~m[1651]&m[1652])|(m[1582]&m[1648]&~m[1649]&~m[1651]&m[1652])|(m[1582]&~m[1648]&m[1649]&~m[1651]&m[1652])|(~m[1582]&~m[1648]&~m[1649]&m[1651]&m[1652])|(m[1582]&~m[1648]&~m[1649]&m[1651]&m[1652])|(~m[1582]&m[1648]&~m[1649]&m[1651]&m[1652])|(m[1582]&m[1648]&~m[1649]&m[1651]&m[1652])|(~m[1582]&~m[1648]&m[1649]&m[1651]&m[1652])|(m[1582]&~m[1648]&m[1649]&m[1651]&m[1652])|(m[1582]&m[1648]&m[1649]&m[1651]&m[1652]))):InitCond[1039];
    m[1655] = run?((((m[1587]&~m[1653]&~m[1654]&~m[1656]&~m[1657])|(~m[1587]&~m[1653]&~m[1654]&m[1656]&~m[1657])|(m[1587]&m[1653]&~m[1654]&m[1656]&~m[1657])|(m[1587]&~m[1653]&m[1654]&m[1656]&~m[1657])|(~m[1587]&m[1653]&~m[1654]&~m[1656]&m[1657])|(~m[1587]&~m[1653]&m[1654]&~m[1656]&m[1657])|(m[1587]&m[1653]&m[1654]&~m[1656]&m[1657])|(~m[1587]&m[1653]&m[1654]&m[1656]&m[1657]))&UnbiasedRNG[401])|((m[1587]&~m[1653]&~m[1654]&m[1656]&~m[1657])|(~m[1587]&~m[1653]&~m[1654]&~m[1656]&m[1657])|(m[1587]&~m[1653]&~m[1654]&~m[1656]&m[1657])|(m[1587]&m[1653]&~m[1654]&~m[1656]&m[1657])|(m[1587]&~m[1653]&m[1654]&~m[1656]&m[1657])|(~m[1587]&~m[1653]&~m[1654]&m[1656]&m[1657])|(m[1587]&~m[1653]&~m[1654]&m[1656]&m[1657])|(~m[1587]&m[1653]&~m[1654]&m[1656]&m[1657])|(m[1587]&m[1653]&~m[1654]&m[1656]&m[1657])|(~m[1587]&~m[1653]&m[1654]&m[1656]&m[1657])|(m[1587]&~m[1653]&m[1654]&m[1656]&m[1657])|(m[1587]&m[1653]&m[1654]&m[1656]&m[1657]))):InitCond[1040];
    m[1660] = run?((((m[1592]&~m[1658]&~m[1659]&~m[1661]&~m[1662])|(~m[1592]&~m[1658]&~m[1659]&m[1661]&~m[1662])|(m[1592]&m[1658]&~m[1659]&m[1661]&~m[1662])|(m[1592]&~m[1658]&m[1659]&m[1661]&~m[1662])|(~m[1592]&m[1658]&~m[1659]&~m[1661]&m[1662])|(~m[1592]&~m[1658]&m[1659]&~m[1661]&m[1662])|(m[1592]&m[1658]&m[1659]&~m[1661]&m[1662])|(~m[1592]&m[1658]&m[1659]&m[1661]&m[1662]))&UnbiasedRNG[402])|((m[1592]&~m[1658]&~m[1659]&m[1661]&~m[1662])|(~m[1592]&~m[1658]&~m[1659]&~m[1661]&m[1662])|(m[1592]&~m[1658]&~m[1659]&~m[1661]&m[1662])|(m[1592]&m[1658]&~m[1659]&~m[1661]&m[1662])|(m[1592]&~m[1658]&m[1659]&~m[1661]&m[1662])|(~m[1592]&~m[1658]&~m[1659]&m[1661]&m[1662])|(m[1592]&~m[1658]&~m[1659]&m[1661]&m[1662])|(~m[1592]&m[1658]&~m[1659]&m[1661]&m[1662])|(m[1592]&m[1658]&~m[1659]&m[1661]&m[1662])|(~m[1592]&~m[1658]&m[1659]&m[1661]&m[1662])|(m[1592]&~m[1658]&m[1659]&m[1661]&m[1662])|(m[1592]&m[1658]&m[1659]&m[1661]&m[1662]))):InitCond[1041];
    m[1665] = run?((((m[1597]&~m[1663]&~m[1664]&~m[1666]&~m[1667])|(~m[1597]&~m[1663]&~m[1664]&m[1666]&~m[1667])|(m[1597]&m[1663]&~m[1664]&m[1666]&~m[1667])|(m[1597]&~m[1663]&m[1664]&m[1666]&~m[1667])|(~m[1597]&m[1663]&~m[1664]&~m[1666]&m[1667])|(~m[1597]&~m[1663]&m[1664]&~m[1666]&m[1667])|(m[1597]&m[1663]&m[1664]&~m[1666]&m[1667])|(~m[1597]&m[1663]&m[1664]&m[1666]&m[1667]))&UnbiasedRNG[403])|((m[1597]&~m[1663]&~m[1664]&m[1666]&~m[1667])|(~m[1597]&~m[1663]&~m[1664]&~m[1666]&m[1667])|(m[1597]&~m[1663]&~m[1664]&~m[1666]&m[1667])|(m[1597]&m[1663]&~m[1664]&~m[1666]&m[1667])|(m[1597]&~m[1663]&m[1664]&~m[1666]&m[1667])|(~m[1597]&~m[1663]&~m[1664]&m[1666]&m[1667])|(m[1597]&~m[1663]&~m[1664]&m[1666]&m[1667])|(~m[1597]&m[1663]&~m[1664]&m[1666]&m[1667])|(m[1597]&m[1663]&~m[1664]&m[1666]&m[1667])|(~m[1597]&~m[1663]&m[1664]&m[1666]&m[1667])|(m[1597]&~m[1663]&m[1664]&m[1666]&m[1667])|(m[1597]&m[1663]&m[1664]&m[1666]&m[1667]))):InitCond[1042];
    m[1670] = run?((((m[1602]&~m[1668]&~m[1669]&~m[1671]&~m[1672])|(~m[1602]&~m[1668]&~m[1669]&m[1671]&~m[1672])|(m[1602]&m[1668]&~m[1669]&m[1671]&~m[1672])|(m[1602]&~m[1668]&m[1669]&m[1671]&~m[1672])|(~m[1602]&m[1668]&~m[1669]&~m[1671]&m[1672])|(~m[1602]&~m[1668]&m[1669]&~m[1671]&m[1672])|(m[1602]&m[1668]&m[1669]&~m[1671]&m[1672])|(~m[1602]&m[1668]&m[1669]&m[1671]&m[1672]))&UnbiasedRNG[404])|((m[1602]&~m[1668]&~m[1669]&m[1671]&~m[1672])|(~m[1602]&~m[1668]&~m[1669]&~m[1671]&m[1672])|(m[1602]&~m[1668]&~m[1669]&~m[1671]&m[1672])|(m[1602]&m[1668]&~m[1669]&~m[1671]&m[1672])|(m[1602]&~m[1668]&m[1669]&~m[1671]&m[1672])|(~m[1602]&~m[1668]&~m[1669]&m[1671]&m[1672])|(m[1602]&~m[1668]&~m[1669]&m[1671]&m[1672])|(~m[1602]&m[1668]&~m[1669]&m[1671]&m[1672])|(m[1602]&m[1668]&~m[1669]&m[1671]&m[1672])|(~m[1602]&~m[1668]&m[1669]&m[1671]&m[1672])|(m[1602]&~m[1668]&m[1669]&m[1671]&m[1672])|(m[1602]&m[1668]&m[1669]&m[1671]&m[1672]))):InitCond[1043];
    m[1675] = run?((((m[1612]&~m[1673]&~m[1674]&~m[1676]&~m[1677])|(~m[1612]&~m[1673]&~m[1674]&m[1676]&~m[1677])|(m[1612]&m[1673]&~m[1674]&m[1676]&~m[1677])|(m[1612]&~m[1673]&m[1674]&m[1676]&~m[1677])|(~m[1612]&m[1673]&~m[1674]&~m[1676]&m[1677])|(~m[1612]&~m[1673]&m[1674]&~m[1676]&m[1677])|(m[1612]&m[1673]&m[1674]&~m[1676]&m[1677])|(~m[1612]&m[1673]&m[1674]&m[1676]&m[1677]))&UnbiasedRNG[405])|((m[1612]&~m[1673]&~m[1674]&m[1676]&~m[1677])|(~m[1612]&~m[1673]&~m[1674]&~m[1676]&m[1677])|(m[1612]&~m[1673]&~m[1674]&~m[1676]&m[1677])|(m[1612]&m[1673]&~m[1674]&~m[1676]&m[1677])|(m[1612]&~m[1673]&m[1674]&~m[1676]&m[1677])|(~m[1612]&~m[1673]&~m[1674]&m[1676]&m[1677])|(m[1612]&~m[1673]&~m[1674]&m[1676]&m[1677])|(~m[1612]&m[1673]&~m[1674]&m[1676]&m[1677])|(m[1612]&m[1673]&~m[1674]&m[1676]&m[1677])|(~m[1612]&~m[1673]&m[1674]&m[1676]&m[1677])|(m[1612]&~m[1673]&m[1674]&m[1676]&m[1677])|(m[1612]&m[1673]&m[1674]&m[1676]&m[1677]))):InitCond[1044];
    m[1680] = run?((((m[1617]&~m[1678]&~m[1679]&~m[1681]&~m[1682])|(~m[1617]&~m[1678]&~m[1679]&m[1681]&~m[1682])|(m[1617]&m[1678]&~m[1679]&m[1681]&~m[1682])|(m[1617]&~m[1678]&m[1679]&m[1681]&~m[1682])|(~m[1617]&m[1678]&~m[1679]&~m[1681]&m[1682])|(~m[1617]&~m[1678]&m[1679]&~m[1681]&m[1682])|(m[1617]&m[1678]&m[1679]&~m[1681]&m[1682])|(~m[1617]&m[1678]&m[1679]&m[1681]&m[1682]))&UnbiasedRNG[406])|((m[1617]&~m[1678]&~m[1679]&m[1681]&~m[1682])|(~m[1617]&~m[1678]&~m[1679]&~m[1681]&m[1682])|(m[1617]&~m[1678]&~m[1679]&~m[1681]&m[1682])|(m[1617]&m[1678]&~m[1679]&~m[1681]&m[1682])|(m[1617]&~m[1678]&m[1679]&~m[1681]&m[1682])|(~m[1617]&~m[1678]&~m[1679]&m[1681]&m[1682])|(m[1617]&~m[1678]&~m[1679]&m[1681]&m[1682])|(~m[1617]&m[1678]&~m[1679]&m[1681]&m[1682])|(m[1617]&m[1678]&~m[1679]&m[1681]&m[1682])|(~m[1617]&~m[1678]&m[1679]&m[1681]&m[1682])|(m[1617]&~m[1678]&m[1679]&m[1681]&m[1682])|(m[1617]&m[1678]&m[1679]&m[1681]&m[1682]))):InitCond[1045];
    m[1685] = run?((((m[1622]&~m[1683]&~m[1684]&~m[1686]&~m[1687])|(~m[1622]&~m[1683]&~m[1684]&m[1686]&~m[1687])|(m[1622]&m[1683]&~m[1684]&m[1686]&~m[1687])|(m[1622]&~m[1683]&m[1684]&m[1686]&~m[1687])|(~m[1622]&m[1683]&~m[1684]&~m[1686]&m[1687])|(~m[1622]&~m[1683]&m[1684]&~m[1686]&m[1687])|(m[1622]&m[1683]&m[1684]&~m[1686]&m[1687])|(~m[1622]&m[1683]&m[1684]&m[1686]&m[1687]))&UnbiasedRNG[407])|((m[1622]&~m[1683]&~m[1684]&m[1686]&~m[1687])|(~m[1622]&~m[1683]&~m[1684]&~m[1686]&m[1687])|(m[1622]&~m[1683]&~m[1684]&~m[1686]&m[1687])|(m[1622]&m[1683]&~m[1684]&~m[1686]&m[1687])|(m[1622]&~m[1683]&m[1684]&~m[1686]&m[1687])|(~m[1622]&~m[1683]&~m[1684]&m[1686]&m[1687])|(m[1622]&~m[1683]&~m[1684]&m[1686]&m[1687])|(~m[1622]&m[1683]&~m[1684]&m[1686]&m[1687])|(m[1622]&m[1683]&~m[1684]&m[1686]&m[1687])|(~m[1622]&~m[1683]&m[1684]&m[1686]&m[1687])|(m[1622]&~m[1683]&m[1684]&m[1686]&m[1687])|(m[1622]&m[1683]&m[1684]&m[1686]&m[1687]))):InitCond[1046];
    m[1690] = run?((((m[1627]&~m[1688]&~m[1689]&~m[1691]&~m[1692])|(~m[1627]&~m[1688]&~m[1689]&m[1691]&~m[1692])|(m[1627]&m[1688]&~m[1689]&m[1691]&~m[1692])|(m[1627]&~m[1688]&m[1689]&m[1691]&~m[1692])|(~m[1627]&m[1688]&~m[1689]&~m[1691]&m[1692])|(~m[1627]&~m[1688]&m[1689]&~m[1691]&m[1692])|(m[1627]&m[1688]&m[1689]&~m[1691]&m[1692])|(~m[1627]&m[1688]&m[1689]&m[1691]&m[1692]))&UnbiasedRNG[408])|((m[1627]&~m[1688]&~m[1689]&m[1691]&~m[1692])|(~m[1627]&~m[1688]&~m[1689]&~m[1691]&m[1692])|(m[1627]&~m[1688]&~m[1689]&~m[1691]&m[1692])|(m[1627]&m[1688]&~m[1689]&~m[1691]&m[1692])|(m[1627]&~m[1688]&m[1689]&~m[1691]&m[1692])|(~m[1627]&~m[1688]&~m[1689]&m[1691]&m[1692])|(m[1627]&~m[1688]&~m[1689]&m[1691]&m[1692])|(~m[1627]&m[1688]&~m[1689]&m[1691]&m[1692])|(m[1627]&m[1688]&~m[1689]&m[1691]&m[1692])|(~m[1627]&~m[1688]&m[1689]&m[1691]&m[1692])|(m[1627]&~m[1688]&m[1689]&m[1691]&m[1692])|(m[1627]&m[1688]&m[1689]&m[1691]&m[1692]))):InitCond[1047];
    m[1695] = run?((((m[1632]&~m[1693]&~m[1694]&~m[1696]&~m[1697])|(~m[1632]&~m[1693]&~m[1694]&m[1696]&~m[1697])|(m[1632]&m[1693]&~m[1694]&m[1696]&~m[1697])|(m[1632]&~m[1693]&m[1694]&m[1696]&~m[1697])|(~m[1632]&m[1693]&~m[1694]&~m[1696]&m[1697])|(~m[1632]&~m[1693]&m[1694]&~m[1696]&m[1697])|(m[1632]&m[1693]&m[1694]&~m[1696]&m[1697])|(~m[1632]&m[1693]&m[1694]&m[1696]&m[1697]))&UnbiasedRNG[409])|((m[1632]&~m[1693]&~m[1694]&m[1696]&~m[1697])|(~m[1632]&~m[1693]&~m[1694]&~m[1696]&m[1697])|(m[1632]&~m[1693]&~m[1694]&~m[1696]&m[1697])|(m[1632]&m[1693]&~m[1694]&~m[1696]&m[1697])|(m[1632]&~m[1693]&m[1694]&~m[1696]&m[1697])|(~m[1632]&~m[1693]&~m[1694]&m[1696]&m[1697])|(m[1632]&~m[1693]&~m[1694]&m[1696]&m[1697])|(~m[1632]&m[1693]&~m[1694]&m[1696]&m[1697])|(m[1632]&m[1693]&~m[1694]&m[1696]&m[1697])|(~m[1632]&~m[1693]&m[1694]&m[1696]&m[1697])|(m[1632]&~m[1693]&m[1694]&m[1696]&m[1697])|(m[1632]&m[1693]&m[1694]&m[1696]&m[1697]))):InitCond[1048];
    m[1700] = run?((((m[1637]&~m[1698]&~m[1699]&~m[1701]&~m[1702])|(~m[1637]&~m[1698]&~m[1699]&m[1701]&~m[1702])|(m[1637]&m[1698]&~m[1699]&m[1701]&~m[1702])|(m[1637]&~m[1698]&m[1699]&m[1701]&~m[1702])|(~m[1637]&m[1698]&~m[1699]&~m[1701]&m[1702])|(~m[1637]&~m[1698]&m[1699]&~m[1701]&m[1702])|(m[1637]&m[1698]&m[1699]&~m[1701]&m[1702])|(~m[1637]&m[1698]&m[1699]&m[1701]&m[1702]))&UnbiasedRNG[410])|((m[1637]&~m[1698]&~m[1699]&m[1701]&~m[1702])|(~m[1637]&~m[1698]&~m[1699]&~m[1701]&m[1702])|(m[1637]&~m[1698]&~m[1699]&~m[1701]&m[1702])|(m[1637]&m[1698]&~m[1699]&~m[1701]&m[1702])|(m[1637]&~m[1698]&m[1699]&~m[1701]&m[1702])|(~m[1637]&~m[1698]&~m[1699]&m[1701]&m[1702])|(m[1637]&~m[1698]&~m[1699]&m[1701]&m[1702])|(~m[1637]&m[1698]&~m[1699]&m[1701]&m[1702])|(m[1637]&m[1698]&~m[1699]&m[1701]&m[1702])|(~m[1637]&~m[1698]&m[1699]&m[1701]&m[1702])|(m[1637]&~m[1698]&m[1699]&m[1701]&m[1702])|(m[1637]&m[1698]&m[1699]&m[1701]&m[1702]))):InitCond[1049];
    m[1705] = run?((((m[1642]&~m[1703]&~m[1704]&~m[1706]&~m[1707])|(~m[1642]&~m[1703]&~m[1704]&m[1706]&~m[1707])|(m[1642]&m[1703]&~m[1704]&m[1706]&~m[1707])|(m[1642]&~m[1703]&m[1704]&m[1706]&~m[1707])|(~m[1642]&m[1703]&~m[1704]&~m[1706]&m[1707])|(~m[1642]&~m[1703]&m[1704]&~m[1706]&m[1707])|(m[1642]&m[1703]&m[1704]&~m[1706]&m[1707])|(~m[1642]&m[1703]&m[1704]&m[1706]&m[1707]))&UnbiasedRNG[411])|((m[1642]&~m[1703]&~m[1704]&m[1706]&~m[1707])|(~m[1642]&~m[1703]&~m[1704]&~m[1706]&m[1707])|(m[1642]&~m[1703]&~m[1704]&~m[1706]&m[1707])|(m[1642]&m[1703]&~m[1704]&~m[1706]&m[1707])|(m[1642]&~m[1703]&m[1704]&~m[1706]&m[1707])|(~m[1642]&~m[1703]&~m[1704]&m[1706]&m[1707])|(m[1642]&~m[1703]&~m[1704]&m[1706]&m[1707])|(~m[1642]&m[1703]&~m[1704]&m[1706]&m[1707])|(m[1642]&m[1703]&~m[1704]&m[1706]&m[1707])|(~m[1642]&~m[1703]&m[1704]&m[1706]&m[1707])|(m[1642]&~m[1703]&m[1704]&m[1706]&m[1707])|(m[1642]&m[1703]&m[1704]&m[1706]&m[1707]))):InitCond[1050];
    m[1710] = run?((((m[1647]&~m[1708]&~m[1709]&~m[1711]&~m[1712])|(~m[1647]&~m[1708]&~m[1709]&m[1711]&~m[1712])|(m[1647]&m[1708]&~m[1709]&m[1711]&~m[1712])|(m[1647]&~m[1708]&m[1709]&m[1711]&~m[1712])|(~m[1647]&m[1708]&~m[1709]&~m[1711]&m[1712])|(~m[1647]&~m[1708]&m[1709]&~m[1711]&m[1712])|(m[1647]&m[1708]&m[1709]&~m[1711]&m[1712])|(~m[1647]&m[1708]&m[1709]&m[1711]&m[1712]))&UnbiasedRNG[412])|((m[1647]&~m[1708]&~m[1709]&m[1711]&~m[1712])|(~m[1647]&~m[1708]&~m[1709]&~m[1711]&m[1712])|(m[1647]&~m[1708]&~m[1709]&~m[1711]&m[1712])|(m[1647]&m[1708]&~m[1709]&~m[1711]&m[1712])|(m[1647]&~m[1708]&m[1709]&~m[1711]&m[1712])|(~m[1647]&~m[1708]&~m[1709]&m[1711]&m[1712])|(m[1647]&~m[1708]&~m[1709]&m[1711]&m[1712])|(~m[1647]&m[1708]&~m[1709]&m[1711]&m[1712])|(m[1647]&m[1708]&~m[1709]&m[1711]&m[1712])|(~m[1647]&~m[1708]&m[1709]&m[1711]&m[1712])|(m[1647]&~m[1708]&m[1709]&m[1711]&m[1712])|(m[1647]&m[1708]&m[1709]&m[1711]&m[1712]))):InitCond[1051];
    m[1715] = run?((((m[1652]&~m[1713]&~m[1714]&~m[1716]&~m[1717])|(~m[1652]&~m[1713]&~m[1714]&m[1716]&~m[1717])|(m[1652]&m[1713]&~m[1714]&m[1716]&~m[1717])|(m[1652]&~m[1713]&m[1714]&m[1716]&~m[1717])|(~m[1652]&m[1713]&~m[1714]&~m[1716]&m[1717])|(~m[1652]&~m[1713]&m[1714]&~m[1716]&m[1717])|(m[1652]&m[1713]&m[1714]&~m[1716]&m[1717])|(~m[1652]&m[1713]&m[1714]&m[1716]&m[1717]))&UnbiasedRNG[413])|((m[1652]&~m[1713]&~m[1714]&m[1716]&~m[1717])|(~m[1652]&~m[1713]&~m[1714]&~m[1716]&m[1717])|(m[1652]&~m[1713]&~m[1714]&~m[1716]&m[1717])|(m[1652]&m[1713]&~m[1714]&~m[1716]&m[1717])|(m[1652]&~m[1713]&m[1714]&~m[1716]&m[1717])|(~m[1652]&~m[1713]&~m[1714]&m[1716]&m[1717])|(m[1652]&~m[1713]&~m[1714]&m[1716]&m[1717])|(~m[1652]&m[1713]&~m[1714]&m[1716]&m[1717])|(m[1652]&m[1713]&~m[1714]&m[1716]&m[1717])|(~m[1652]&~m[1713]&m[1714]&m[1716]&m[1717])|(m[1652]&~m[1713]&m[1714]&m[1716]&m[1717])|(m[1652]&m[1713]&m[1714]&m[1716]&m[1717]))):InitCond[1052];
    m[1720] = run?((((m[1657]&~m[1718]&~m[1719]&~m[1721]&~m[1722])|(~m[1657]&~m[1718]&~m[1719]&m[1721]&~m[1722])|(m[1657]&m[1718]&~m[1719]&m[1721]&~m[1722])|(m[1657]&~m[1718]&m[1719]&m[1721]&~m[1722])|(~m[1657]&m[1718]&~m[1719]&~m[1721]&m[1722])|(~m[1657]&~m[1718]&m[1719]&~m[1721]&m[1722])|(m[1657]&m[1718]&m[1719]&~m[1721]&m[1722])|(~m[1657]&m[1718]&m[1719]&m[1721]&m[1722]))&UnbiasedRNG[414])|((m[1657]&~m[1718]&~m[1719]&m[1721]&~m[1722])|(~m[1657]&~m[1718]&~m[1719]&~m[1721]&m[1722])|(m[1657]&~m[1718]&~m[1719]&~m[1721]&m[1722])|(m[1657]&m[1718]&~m[1719]&~m[1721]&m[1722])|(m[1657]&~m[1718]&m[1719]&~m[1721]&m[1722])|(~m[1657]&~m[1718]&~m[1719]&m[1721]&m[1722])|(m[1657]&~m[1718]&~m[1719]&m[1721]&m[1722])|(~m[1657]&m[1718]&~m[1719]&m[1721]&m[1722])|(m[1657]&m[1718]&~m[1719]&m[1721]&m[1722])|(~m[1657]&~m[1718]&m[1719]&m[1721]&m[1722])|(m[1657]&~m[1718]&m[1719]&m[1721]&m[1722])|(m[1657]&m[1718]&m[1719]&m[1721]&m[1722]))):InitCond[1053];
    m[1725] = run?((((m[1662]&~m[1723]&~m[1724]&~m[1726]&~m[1727])|(~m[1662]&~m[1723]&~m[1724]&m[1726]&~m[1727])|(m[1662]&m[1723]&~m[1724]&m[1726]&~m[1727])|(m[1662]&~m[1723]&m[1724]&m[1726]&~m[1727])|(~m[1662]&m[1723]&~m[1724]&~m[1726]&m[1727])|(~m[1662]&~m[1723]&m[1724]&~m[1726]&m[1727])|(m[1662]&m[1723]&m[1724]&~m[1726]&m[1727])|(~m[1662]&m[1723]&m[1724]&m[1726]&m[1727]))&UnbiasedRNG[415])|((m[1662]&~m[1723]&~m[1724]&m[1726]&~m[1727])|(~m[1662]&~m[1723]&~m[1724]&~m[1726]&m[1727])|(m[1662]&~m[1723]&~m[1724]&~m[1726]&m[1727])|(m[1662]&m[1723]&~m[1724]&~m[1726]&m[1727])|(m[1662]&~m[1723]&m[1724]&~m[1726]&m[1727])|(~m[1662]&~m[1723]&~m[1724]&m[1726]&m[1727])|(m[1662]&~m[1723]&~m[1724]&m[1726]&m[1727])|(~m[1662]&m[1723]&~m[1724]&m[1726]&m[1727])|(m[1662]&m[1723]&~m[1724]&m[1726]&m[1727])|(~m[1662]&~m[1723]&m[1724]&m[1726]&m[1727])|(m[1662]&~m[1723]&m[1724]&m[1726]&m[1727])|(m[1662]&m[1723]&m[1724]&m[1726]&m[1727]))):InitCond[1054];
    m[1730] = run?((((m[1667]&~m[1728]&~m[1729]&~m[1731]&~m[1732])|(~m[1667]&~m[1728]&~m[1729]&m[1731]&~m[1732])|(m[1667]&m[1728]&~m[1729]&m[1731]&~m[1732])|(m[1667]&~m[1728]&m[1729]&m[1731]&~m[1732])|(~m[1667]&m[1728]&~m[1729]&~m[1731]&m[1732])|(~m[1667]&~m[1728]&m[1729]&~m[1731]&m[1732])|(m[1667]&m[1728]&m[1729]&~m[1731]&m[1732])|(~m[1667]&m[1728]&m[1729]&m[1731]&m[1732]))&UnbiasedRNG[416])|((m[1667]&~m[1728]&~m[1729]&m[1731]&~m[1732])|(~m[1667]&~m[1728]&~m[1729]&~m[1731]&m[1732])|(m[1667]&~m[1728]&~m[1729]&~m[1731]&m[1732])|(m[1667]&m[1728]&~m[1729]&~m[1731]&m[1732])|(m[1667]&~m[1728]&m[1729]&~m[1731]&m[1732])|(~m[1667]&~m[1728]&~m[1729]&m[1731]&m[1732])|(m[1667]&~m[1728]&~m[1729]&m[1731]&m[1732])|(~m[1667]&m[1728]&~m[1729]&m[1731]&m[1732])|(m[1667]&m[1728]&~m[1729]&m[1731]&m[1732])|(~m[1667]&~m[1728]&m[1729]&m[1731]&m[1732])|(m[1667]&~m[1728]&m[1729]&m[1731]&m[1732])|(m[1667]&m[1728]&m[1729]&m[1731]&m[1732]))):InitCond[1055];
    m[1735] = run?((((m[1672]&~m[1733]&~m[1734]&~m[1736]&~m[1737])|(~m[1672]&~m[1733]&~m[1734]&m[1736]&~m[1737])|(m[1672]&m[1733]&~m[1734]&m[1736]&~m[1737])|(m[1672]&~m[1733]&m[1734]&m[1736]&~m[1737])|(~m[1672]&m[1733]&~m[1734]&~m[1736]&m[1737])|(~m[1672]&~m[1733]&m[1734]&~m[1736]&m[1737])|(m[1672]&m[1733]&m[1734]&~m[1736]&m[1737])|(~m[1672]&m[1733]&m[1734]&m[1736]&m[1737]))&UnbiasedRNG[417])|((m[1672]&~m[1733]&~m[1734]&m[1736]&~m[1737])|(~m[1672]&~m[1733]&~m[1734]&~m[1736]&m[1737])|(m[1672]&~m[1733]&~m[1734]&~m[1736]&m[1737])|(m[1672]&m[1733]&~m[1734]&~m[1736]&m[1737])|(m[1672]&~m[1733]&m[1734]&~m[1736]&m[1737])|(~m[1672]&~m[1733]&~m[1734]&m[1736]&m[1737])|(m[1672]&~m[1733]&~m[1734]&m[1736]&m[1737])|(~m[1672]&m[1733]&~m[1734]&m[1736]&m[1737])|(m[1672]&m[1733]&~m[1734]&m[1736]&m[1737])|(~m[1672]&~m[1733]&m[1734]&m[1736]&m[1737])|(m[1672]&~m[1733]&m[1734]&m[1736]&m[1737])|(m[1672]&m[1733]&m[1734]&m[1736]&m[1737]))):InitCond[1056];
    m[1740] = run?((((m[1682]&~m[1738]&~m[1739]&~m[1741]&~m[1742])|(~m[1682]&~m[1738]&~m[1739]&m[1741]&~m[1742])|(m[1682]&m[1738]&~m[1739]&m[1741]&~m[1742])|(m[1682]&~m[1738]&m[1739]&m[1741]&~m[1742])|(~m[1682]&m[1738]&~m[1739]&~m[1741]&m[1742])|(~m[1682]&~m[1738]&m[1739]&~m[1741]&m[1742])|(m[1682]&m[1738]&m[1739]&~m[1741]&m[1742])|(~m[1682]&m[1738]&m[1739]&m[1741]&m[1742]))&UnbiasedRNG[418])|((m[1682]&~m[1738]&~m[1739]&m[1741]&~m[1742])|(~m[1682]&~m[1738]&~m[1739]&~m[1741]&m[1742])|(m[1682]&~m[1738]&~m[1739]&~m[1741]&m[1742])|(m[1682]&m[1738]&~m[1739]&~m[1741]&m[1742])|(m[1682]&~m[1738]&m[1739]&~m[1741]&m[1742])|(~m[1682]&~m[1738]&~m[1739]&m[1741]&m[1742])|(m[1682]&~m[1738]&~m[1739]&m[1741]&m[1742])|(~m[1682]&m[1738]&~m[1739]&m[1741]&m[1742])|(m[1682]&m[1738]&~m[1739]&m[1741]&m[1742])|(~m[1682]&~m[1738]&m[1739]&m[1741]&m[1742])|(m[1682]&~m[1738]&m[1739]&m[1741]&m[1742])|(m[1682]&m[1738]&m[1739]&m[1741]&m[1742]))):InitCond[1057];
    m[1745] = run?((((m[1687]&~m[1743]&~m[1744]&~m[1746]&~m[1747])|(~m[1687]&~m[1743]&~m[1744]&m[1746]&~m[1747])|(m[1687]&m[1743]&~m[1744]&m[1746]&~m[1747])|(m[1687]&~m[1743]&m[1744]&m[1746]&~m[1747])|(~m[1687]&m[1743]&~m[1744]&~m[1746]&m[1747])|(~m[1687]&~m[1743]&m[1744]&~m[1746]&m[1747])|(m[1687]&m[1743]&m[1744]&~m[1746]&m[1747])|(~m[1687]&m[1743]&m[1744]&m[1746]&m[1747]))&UnbiasedRNG[419])|((m[1687]&~m[1743]&~m[1744]&m[1746]&~m[1747])|(~m[1687]&~m[1743]&~m[1744]&~m[1746]&m[1747])|(m[1687]&~m[1743]&~m[1744]&~m[1746]&m[1747])|(m[1687]&m[1743]&~m[1744]&~m[1746]&m[1747])|(m[1687]&~m[1743]&m[1744]&~m[1746]&m[1747])|(~m[1687]&~m[1743]&~m[1744]&m[1746]&m[1747])|(m[1687]&~m[1743]&~m[1744]&m[1746]&m[1747])|(~m[1687]&m[1743]&~m[1744]&m[1746]&m[1747])|(m[1687]&m[1743]&~m[1744]&m[1746]&m[1747])|(~m[1687]&~m[1743]&m[1744]&m[1746]&m[1747])|(m[1687]&~m[1743]&m[1744]&m[1746]&m[1747])|(m[1687]&m[1743]&m[1744]&m[1746]&m[1747]))):InitCond[1058];
    m[1750] = run?((((m[1692]&~m[1748]&~m[1749]&~m[1751]&~m[1752])|(~m[1692]&~m[1748]&~m[1749]&m[1751]&~m[1752])|(m[1692]&m[1748]&~m[1749]&m[1751]&~m[1752])|(m[1692]&~m[1748]&m[1749]&m[1751]&~m[1752])|(~m[1692]&m[1748]&~m[1749]&~m[1751]&m[1752])|(~m[1692]&~m[1748]&m[1749]&~m[1751]&m[1752])|(m[1692]&m[1748]&m[1749]&~m[1751]&m[1752])|(~m[1692]&m[1748]&m[1749]&m[1751]&m[1752]))&UnbiasedRNG[420])|((m[1692]&~m[1748]&~m[1749]&m[1751]&~m[1752])|(~m[1692]&~m[1748]&~m[1749]&~m[1751]&m[1752])|(m[1692]&~m[1748]&~m[1749]&~m[1751]&m[1752])|(m[1692]&m[1748]&~m[1749]&~m[1751]&m[1752])|(m[1692]&~m[1748]&m[1749]&~m[1751]&m[1752])|(~m[1692]&~m[1748]&~m[1749]&m[1751]&m[1752])|(m[1692]&~m[1748]&~m[1749]&m[1751]&m[1752])|(~m[1692]&m[1748]&~m[1749]&m[1751]&m[1752])|(m[1692]&m[1748]&~m[1749]&m[1751]&m[1752])|(~m[1692]&~m[1748]&m[1749]&m[1751]&m[1752])|(m[1692]&~m[1748]&m[1749]&m[1751]&m[1752])|(m[1692]&m[1748]&m[1749]&m[1751]&m[1752]))):InitCond[1059];
    m[1755] = run?((((m[1697]&~m[1753]&~m[1754]&~m[1756]&~m[1757])|(~m[1697]&~m[1753]&~m[1754]&m[1756]&~m[1757])|(m[1697]&m[1753]&~m[1754]&m[1756]&~m[1757])|(m[1697]&~m[1753]&m[1754]&m[1756]&~m[1757])|(~m[1697]&m[1753]&~m[1754]&~m[1756]&m[1757])|(~m[1697]&~m[1753]&m[1754]&~m[1756]&m[1757])|(m[1697]&m[1753]&m[1754]&~m[1756]&m[1757])|(~m[1697]&m[1753]&m[1754]&m[1756]&m[1757]))&UnbiasedRNG[421])|((m[1697]&~m[1753]&~m[1754]&m[1756]&~m[1757])|(~m[1697]&~m[1753]&~m[1754]&~m[1756]&m[1757])|(m[1697]&~m[1753]&~m[1754]&~m[1756]&m[1757])|(m[1697]&m[1753]&~m[1754]&~m[1756]&m[1757])|(m[1697]&~m[1753]&m[1754]&~m[1756]&m[1757])|(~m[1697]&~m[1753]&~m[1754]&m[1756]&m[1757])|(m[1697]&~m[1753]&~m[1754]&m[1756]&m[1757])|(~m[1697]&m[1753]&~m[1754]&m[1756]&m[1757])|(m[1697]&m[1753]&~m[1754]&m[1756]&m[1757])|(~m[1697]&~m[1753]&m[1754]&m[1756]&m[1757])|(m[1697]&~m[1753]&m[1754]&m[1756]&m[1757])|(m[1697]&m[1753]&m[1754]&m[1756]&m[1757]))):InitCond[1060];
    m[1760] = run?((((m[1702]&~m[1758]&~m[1759]&~m[1761]&~m[1762])|(~m[1702]&~m[1758]&~m[1759]&m[1761]&~m[1762])|(m[1702]&m[1758]&~m[1759]&m[1761]&~m[1762])|(m[1702]&~m[1758]&m[1759]&m[1761]&~m[1762])|(~m[1702]&m[1758]&~m[1759]&~m[1761]&m[1762])|(~m[1702]&~m[1758]&m[1759]&~m[1761]&m[1762])|(m[1702]&m[1758]&m[1759]&~m[1761]&m[1762])|(~m[1702]&m[1758]&m[1759]&m[1761]&m[1762]))&UnbiasedRNG[422])|((m[1702]&~m[1758]&~m[1759]&m[1761]&~m[1762])|(~m[1702]&~m[1758]&~m[1759]&~m[1761]&m[1762])|(m[1702]&~m[1758]&~m[1759]&~m[1761]&m[1762])|(m[1702]&m[1758]&~m[1759]&~m[1761]&m[1762])|(m[1702]&~m[1758]&m[1759]&~m[1761]&m[1762])|(~m[1702]&~m[1758]&~m[1759]&m[1761]&m[1762])|(m[1702]&~m[1758]&~m[1759]&m[1761]&m[1762])|(~m[1702]&m[1758]&~m[1759]&m[1761]&m[1762])|(m[1702]&m[1758]&~m[1759]&m[1761]&m[1762])|(~m[1702]&~m[1758]&m[1759]&m[1761]&m[1762])|(m[1702]&~m[1758]&m[1759]&m[1761]&m[1762])|(m[1702]&m[1758]&m[1759]&m[1761]&m[1762]))):InitCond[1061];
    m[1765] = run?((((m[1707]&~m[1763]&~m[1764]&~m[1766]&~m[1767])|(~m[1707]&~m[1763]&~m[1764]&m[1766]&~m[1767])|(m[1707]&m[1763]&~m[1764]&m[1766]&~m[1767])|(m[1707]&~m[1763]&m[1764]&m[1766]&~m[1767])|(~m[1707]&m[1763]&~m[1764]&~m[1766]&m[1767])|(~m[1707]&~m[1763]&m[1764]&~m[1766]&m[1767])|(m[1707]&m[1763]&m[1764]&~m[1766]&m[1767])|(~m[1707]&m[1763]&m[1764]&m[1766]&m[1767]))&UnbiasedRNG[423])|((m[1707]&~m[1763]&~m[1764]&m[1766]&~m[1767])|(~m[1707]&~m[1763]&~m[1764]&~m[1766]&m[1767])|(m[1707]&~m[1763]&~m[1764]&~m[1766]&m[1767])|(m[1707]&m[1763]&~m[1764]&~m[1766]&m[1767])|(m[1707]&~m[1763]&m[1764]&~m[1766]&m[1767])|(~m[1707]&~m[1763]&~m[1764]&m[1766]&m[1767])|(m[1707]&~m[1763]&~m[1764]&m[1766]&m[1767])|(~m[1707]&m[1763]&~m[1764]&m[1766]&m[1767])|(m[1707]&m[1763]&~m[1764]&m[1766]&m[1767])|(~m[1707]&~m[1763]&m[1764]&m[1766]&m[1767])|(m[1707]&~m[1763]&m[1764]&m[1766]&m[1767])|(m[1707]&m[1763]&m[1764]&m[1766]&m[1767]))):InitCond[1062];
    m[1770] = run?((((m[1712]&~m[1768]&~m[1769]&~m[1771]&~m[1772])|(~m[1712]&~m[1768]&~m[1769]&m[1771]&~m[1772])|(m[1712]&m[1768]&~m[1769]&m[1771]&~m[1772])|(m[1712]&~m[1768]&m[1769]&m[1771]&~m[1772])|(~m[1712]&m[1768]&~m[1769]&~m[1771]&m[1772])|(~m[1712]&~m[1768]&m[1769]&~m[1771]&m[1772])|(m[1712]&m[1768]&m[1769]&~m[1771]&m[1772])|(~m[1712]&m[1768]&m[1769]&m[1771]&m[1772]))&UnbiasedRNG[424])|((m[1712]&~m[1768]&~m[1769]&m[1771]&~m[1772])|(~m[1712]&~m[1768]&~m[1769]&~m[1771]&m[1772])|(m[1712]&~m[1768]&~m[1769]&~m[1771]&m[1772])|(m[1712]&m[1768]&~m[1769]&~m[1771]&m[1772])|(m[1712]&~m[1768]&m[1769]&~m[1771]&m[1772])|(~m[1712]&~m[1768]&~m[1769]&m[1771]&m[1772])|(m[1712]&~m[1768]&~m[1769]&m[1771]&m[1772])|(~m[1712]&m[1768]&~m[1769]&m[1771]&m[1772])|(m[1712]&m[1768]&~m[1769]&m[1771]&m[1772])|(~m[1712]&~m[1768]&m[1769]&m[1771]&m[1772])|(m[1712]&~m[1768]&m[1769]&m[1771]&m[1772])|(m[1712]&m[1768]&m[1769]&m[1771]&m[1772]))):InitCond[1063];
    m[1775] = run?((((m[1717]&~m[1773]&~m[1774]&~m[1776]&~m[1777])|(~m[1717]&~m[1773]&~m[1774]&m[1776]&~m[1777])|(m[1717]&m[1773]&~m[1774]&m[1776]&~m[1777])|(m[1717]&~m[1773]&m[1774]&m[1776]&~m[1777])|(~m[1717]&m[1773]&~m[1774]&~m[1776]&m[1777])|(~m[1717]&~m[1773]&m[1774]&~m[1776]&m[1777])|(m[1717]&m[1773]&m[1774]&~m[1776]&m[1777])|(~m[1717]&m[1773]&m[1774]&m[1776]&m[1777]))&UnbiasedRNG[425])|((m[1717]&~m[1773]&~m[1774]&m[1776]&~m[1777])|(~m[1717]&~m[1773]&~m[1774]&~m[1776]&m[1777])|(m[1717]&~m[1773]&~m[1774]&~m[1776]&m[1777])|(m[1717]&m[1773]&~m[1774]&~m[1776]&m[1777])|(m[1717]&~m[1773]&m[1774]&~m[1776]&m[1777])|(~m[1717]&~m[1773]&~m[1774]&m[1776]&m[1777])|(m[1717]&~m[1773]&~m[1774]&m[1776]&m[1777])|(~m[1717]&m[1773]&~m[1774]&m[1776]&m[1777])|(m[1717]&m[1773]&~m[1774]&m[1776]&m[1777])|(~m[1717]&~m[1773]&m[1774]&m[1776]&m[1777])|(m[1717]&~m[1773]&m[1774]&m[1776]&m[1777])|(m[1717]&m[1773]&m[1774]&m[1776]&m[1777]))):InitCond[1064];
    m[1780] = run?((((m[1722]&~m[1778]&~m[1779]&~m[1781]&~m[1782])|(~m[1722]&~m[1778]&~m[1779]&m[1781]&~m[1782])|(m[1722]&m[1778]&~m[1779]&m[1781]&~m[1782])|(m[1722]&~m[1778]&m[1779]&m[1781]&~m[1782])|(~m[1722]&m[1778]&~m[1779]&~m[1781]&m[1782])|(~m[1722]&~m[1778]&m[1779]&~m[1781]&m[1782])|(m[1722]&m[1778]&m[1779]&~m[1781]&m[1782])|(~m[1722]&m[1778]&m[1779]&m[1781]&m[1782]))&UnbiasedRNG[426])|((m[1722]&~m[1778]&~m[1779]&m[1781]&~m[1782])|(~m[1722]&~m[1778]&~m[1779]&~m[1781]&m[1782])|(m[1722]&~m[1778]&~m[1779]&~m[1781]&m[1782])|(m[1722]&m[1778]&~m[1779]&~m[1781]&m[1782])|(m[1722]&~m[1778]&m[1779]&~m[1781]&m[1782])|(~m[1722]&~m[1778]&~m[1779]&m[1781]&m[1782])|(m[1722]&~m[1778]&~m[1779]&m[1781]&m[1782])|(~m[1722]&m[1778]&~m[1779]&m[1781]&m[1782])|(m[1722]&m[1778]&~m[1779]&m[1781]&m[1782])|(~m[1722]&~m[1778]&m[1779]&m[1781]&m[1782])|(m[1722]&~m[1778]&m[1779]&m[1781]&m[1782])|(m[1722]&m[1778]&m[1779]&m[1781]&m[1782]))):InitCond[1065];
    m[1785] = run?((((m[1727]&~m[1783]&~m[1784]&~m[1786]&~m[1787])|(~m[1727]&~m[1783]&~m[1784]&m[1786]&~m[1787])|(m[1727]&m[1783]&~m[1784]&m[1786]&~m[1787])|(m[1727]&~m[1783]&m[1784]&m[1786]&~m[1787])|(~m[1727]&m[1783]&~m[1784]&~m[1786]&m[1787])|(~m[1727]&~m[1783]&m[1784]&~m[1786]&m[1787])|(m[1727]&m[1783]&m[1784]&~m[1786]&m[1787])|(~m[1727]&m[1783]&m[1784]&m[1786]&m[1787]))&UnbiasedRNG[427])|((m[1727]&~m[1783]&~m[1784]&m[1786]&~m[1787])|(~m[1727]&~m[1783]&~m[1784]&~m[1786]&m[1787])|(m[1727]&~m[1783]&~m[1784]&~m[1786]&m[1787])|(m[1727]&m[1783]&~m[1784]&~m[1786]&m[1787])|(m[1727]&~m[1783]&m[1784]&~m[1786]&m[1787])|(~m[1727]&~m[1783]&~m[1784]&m[1786]&m[1787])|(m[1727]&~m[1783]&~m[1784]&m[1786]&m[1787])|(~m[1727]&m[1783]&~m[1784]&m[1786]&m[1787])|(m[1727]&m[1783]&~m[1784]&m[1786]&m[1787])|(~m[1727]&~m[1783]&m[1784]&m[1786]&m[1787])|(m[1727]&~m[1783]&m[1784]&m[1786]&m[1787])|(m[1727]&m[1783]&m[1784]&m[1786]&m[1787]))):InitCond[1066];
    m[1790] = run?((((m[1732]&~m[1788]&~m[1789]&~m[1791]&~m[1792])|(~m[1732]&~m[1788]&~m[1789]&m[1791]&~m[1792])|(m[1732]&m[1788]&~m[1789]&m[1791]&~m[1792])|(m[1732]&~m[1788]&m[1789]&m[1791]&~m[1792])|(~m[1732]&m[1788]&~m[1789]&~m[1791]&m[1792])|(~m[1732]&~m[1788]&m[1789]&~m[1791]&m[1792])|(m[1732]&m[1788]&m[1789]&~m[1791]&m[1792])|(~m[1732]&m[1788]&m[1789]&m[1791]&m[1792]))&UnbiasedRNG[428])|((m[1732]&~m[1788]&~m[1789]&m[1791]&~m[1792])|(~m[1732]&~m[1788]&~m[1789]&~m[1791]&m[1792])|(m[1732]&~m[1788]&~m[1789]&~m[1791]&m[1792])|(m[1732]&m[1788]&~m[1789]&~m[1791]&m[1792])|(m[1732]&~m[1788]&m[1789]&~m[1791]&m[1792])|(~m[1732]&~m[1788]&~m[1789]&m[1791]&m[1792])|(m[1732]&~m[1788]&~m[1789]&m[1791]&m[1792])|(~m[1732]&m[1788]&~m[1789]&m[1791]&m[1792])|(m[1732]&m[1788]&~m[1789]&m[1791]&m[1792])|(~m[1732]&~m[1788]&m[1789]&m[1791]&m[1792])|(m[1732]&~m[1788]&m[1789]&m[1791]&m[1792])|(m[1732]&m[1788]&m[1789]&m[1791]&m[1792]))):InitCond[1067];
    m[1795] = run?((((m[1737]&~m[1793]&~m[1794]&~m[1796]&~m[1797])|(~m[1737]&~m[1793]&~m[1794]&m[1796]&~m[1797])|(m[1737]&m[1793]&~m[1794]&m[1796]&~m[1797])|(m[1737]&~m[1793]&m[1794]&m[1796]&~m[1797])|(~m[1737]&m[1793]&~m[1794]&~m[1796]&m[1797])|(~m[1737]&~m[1793]&m[1794]&~m[1796]&m[1797])|(m[1737]&m[1793]&m[1794]&~m[1796]&m[1797])|(~m[1737]&m[1793]&m[1794]&m[1796]&m[1797]))&UnbiasedRNG[429])|((m[1737]&~m[1793]&~m[1794]&m[1796]&~m[1797])|(~m[1737]&~m[1793]&~m[1794]&~m[1796]&m[1797])|(m[1737]&~m[1793]&~m[1794]&~m[1796]&m[1797])|(m[1737]&m[1793]&~m[1794]&~m[1796]&m[1797])|(m[1737]&~m[1793]&m[1794]&~m[1796]&m[1797])|(~m[1737]&~m[1793]&~m[1794]&m[1796]&m[1797])|(m[1737]&~m[1793]&~m[1794]&m[1796]&m[1797])|(~m[1737]&m[1793]&~m[1794]&m[1796]&m[1797])|(m[1737]&m[1793]&~m[1794]&m[1796]&m[1797])|(~m[1737]&~m[1793]&m[1794]&m[1796]&m[1797])|(m[1737]&~m[1793]&m[1794]&m[1796]&m[1797])|(m[1737]&m[1793]&m[1794]&m[1796]&m[1797]))):InitCond[1068];
    m[1800] = run?((((m[1747]&~m[1798]&~m[1799]&~m[1801]&~m[1802])|(~m[1747]&~m[1798]&~m[1799]&m[1801]&~m[1802])|(m[1747]&m[1798]&~m[1799]&m[1801]&~m[1802])|(m[1747]&~m[1798]&m[1799]&m[1801]&~m[1802])|(~m[1747]&m[1798]&~m[1799]&~m[1801]&m[1802])|(~m[1747]&~m[1798]&m[1799]&~m[1801]&m[1802])|(m[1747]&m[1798]&m[1799]&~m[1801]&m[1802])|(~m[1747]&m[1798]&m[1799]&m[1801]&m[1802]))&UnbiasedRNG[430])|((m[1747]&~m[1798]&~m[1799]&m[1801]&~m[1802])|(~m[1747]&~m[1798]&~m[1799]&~m[1801]&m[1802])|(m[1747]&~m[1798]&~m[1799]&~m[1801]&m[1802])|(m[1747]&m[1798]&~m[1799]&~m[1801]&m[1802])|(m[1747]&~m[1798]&m[1799]&~m[1801]&m[1802])|(~m[1747]&~m[1798]&~m[1799]&m[1801]&m[1802])|(m[1747]&~m[1798]&~m[1799]&m[1801]&m[1802])|(~m[1747]&m[1798]&~m[1799]&m[1801]&m[1802])|(m[1747]&m[1798]&~m[1799]&m[1801]&m[1802])|(~m[1747]&~m[1798]&m[1799]&m[1801]&m[1802])|(m[1747]&~m[1798]&m[1799]&m[1801]&m[1802])|(m[1747]&m[1798]&m[1799]&m[1801]&m[1802]))):InitCond[1069];
    m[1805] = run?((((m[1752]&~m[1803]&~m[1804]&~m[1806]&~m[1807])|(~m[1752]&~m[1803]&~m[1804]&m[1806]&~m[1807])|(m[1752]&m[1803]&~m[1804]&m[1806]&~m[1807])|(m[1752]&~m[1803]&m[1804]&m[1806]&~m[1807])|(~m[1752]&m[1803]&~m[1804]&~m[1806]&m[1807])|(~m[1752]&~m[1803]&m[1804]&~m[1806]&m[1807])|(m[1752]&m[1803]&m[1804]&~m[1806]&m[1807])|(~m[1752]&m[1803]&m[1804]&m[1806]&m[1807]))&UnbiasedRNG[431])|((m[1752]&~m[1803]&~m[1804]&m[1806]&~m[1807])|(~m[1752]&~m[1803]&~m[1804]&~m[1806]&m[1807])|(m[1752]&~m[1803]&~m[1804]&~m[1806]&m[1807])|(m[1752]&m[1803]&~m[1804]&~m[1806]&m[1807])|(m[1752]&~m[1803]&m[1804]&~m[1806]&m[1807])|(~m[1752]&~m[1803]&~m[1804]&m[1806]&m[1807])|(m[1752]&~m[1803]&~m[1804]&m[1806]&m[1807])|(~m[1752]&m[1803]&~m[1804]&m[1806]&m[1807])|(m[1752]&m[1803]&~m[1804]&m[1806]&m[1807])|(~m[1752]&~m[1803]&m[1804]&m[1806]&m[1807])|(m[1752]&~m[1803]&m[1804]&m[1806]&m[1807])|(m[1752]&m[1803]&m[1804]&m[1806]&m[1807]))):InitCond[1070];
    m[1810] = run?((((m[1757]&~m[1808]&~m[1809]&~m[1811]&~m[1812])|(~m[1757]&~m[1808]&~m[1809]&m[1811]&~m[1812])|(m[1757]&m[1808]&~m[1809]&m[1811]&~m[1812])|(m[1757]&~m[1808]&m[1809]&m[1811]&~m[1812])|(~m[1757]&m[1808]&~m[1809]&~m[1811]&m[1812])|(~m[1757]&~m[1808]&m[1809]&~m[1811]&m[1812])|(m[1757]&m[1808]&m[1809]&~m[1811]&m[1812])|(~m[1757]&m[1808]&m[1809]&m[1811]&m[1812]))&UnbiasedRNG[432])|((m[1757]&~m[1808]&~m[1809]&m[1811]&~m[1812])|(~m[1757]&~m[1808]&~m[1809]&~m[1811]&m[1812])|(m[1757]&~m[1808]&~m[1809]&~m[1811]&m[1812])|(m[1757]&m[1808]&~m[1809]&~m[1811]&m[1812])|(m[1757]&~m[1808]&m[1809]&~m[1811]&m[1812])|(~m[1757]&~m[1808]&~m[1809]&m[1811]&m[1812])|(m[1757]&~m[1808]&~m[1809]&m[1811]&m[1812])|(~m[1757]&m[1808]&~m[1809]&m[1811]&m[1812])|(m[1757]&m[1808]&~m[1809]&m[1811]&m[1812])|(~m[1757]&~m[1808]&m[1809]&m[1811]&m[1812])|(m[1757]&~m[1808]&m[1809]&m[1811]&m[1812])|(m[1757]&m[1808]&m[1809]&m[1811]&m[1812]))):InitCond[1071];
    m[1815] = run?((((m[1762]&~m[1813]&~m[1814]&~m[1816]&~m[1817])|(~m[1762]&~m[1813]&~m[1814]&m[1816]&~m[1817])|(m[1762]&m[1813]&~m[1814]&m[1816]&~m[1817])|(m[1762]&~m[1813]&m[1814]&m[1816]&~m[1817])|(~m[1762]&m[1813]&~m[1814]&~m[1816]&m[1817])|(~m[1762]&~m[1813]&m[1814]&~m[1816]&m[1817])|(m[1762]&m[1813]&m[1814]&~m[1816]&m[1817])|(~m[1762]&m[1813]&m[1814]&m[1816]&m[1817]))&UnbiasedRNG[433])|((m[1762]&~m[1813]&~m[1814]&m[1816]&~m[1817])|(~m[1762]&~m[1813]&~m[1814]&~m[1816]&m[1817])|(m[1762]&~m[1813]&~m[1814]&~m[1816]&m[1817])|(m[1762]&m[1813]&~m[1814]&~m[1816]&m[1817])|(m[1762]&~m[1813]&m[1814]&~m[1816]&m[1817])|(~m[1762]&~m[1813]&~m[1814]&m[1816]&m[1817])|(m[1762]&~m[1813]&~m[1814]&m[1816]&m[1817])|(~m[1762]&m[1813]&~m[1814]&m[1816]&m[1817])|(m[1762]&m[1813]&~m[1814]&m[1816]&m[1817])|(~m[1762]&~m[1813]&m[1814]&m[1816]&m[1817])|(m[1762]&~m[1813]&m[1814]&m[1816]&m[1817])|(m[1762]&m[1813]&m[1814]&m[1816]&m[1817]))):InitCond[1072];
    m[1820] = run?((((m[1767]&~m[1818]&~m[1819]&~m[1821]&~m[1822])|(~m[1767]&~m[1818]&~m[1819]&m[1821]&~m[1822])|(m[1767]&m[1818]&~m[1819]&m[1821]&~m[1822])|(m[1767]&~m[1818]&m[1819]&m[1821]&~m[1822])|(~m[1767]&m[1818]&~m[1819]&~m[1821]&m[1822])|(~m[1767]&~m[1818]&m[1819]&~m[1821]&m[1822])|(m[1767]&m[1818]&m[1819]&~m[1821]&m[1822])|(~m[1767]&m[1818]&m[1819]&m[1821]&m[1822]))&UnbiasedRNG[434])|((m[1767]&~m[1818]&~m[1819]&m[1821]&~m[1822])|(~m[1767]&~m[1818]&~m[1819]&~m[1821]&m[1822])|(m[1767]&~m[1818]&~m[1819]&~m[1821]&m[1822])|(m[1767]&m[1818]&~m[1819]&~m[1821]&m[1822])|(m[1767]&~m[1818]&m[1819]&~m[1821]&m[1822])|(~m[1767]&~m[1818]&~m[1819]&m[1821]&m[1822])|(m[1767]&~m[1818]&~m[1819]&m[1821]&m[1822])|(~m[1767]&m[1818]&~m[1819]&m[1821]&m[1822])|(m[1767]&m[1818]&~m[1819]&m[1821]&m[1822])|(~m[1767]&~m[1818]&m[1819]&m[1821]&m[1822])|(m[1767]&~m[1818]&m[1819]&m[1821]&m[1822])|(m[1767]&m[1818]&m[1819]&m[1821]&m[1822]))):InitCond[1073];
    m[1825] = run?((((m[1772]&~m[1823]&~m[1824]&~m[1826]&~m[1827])|(~m[1772]&~m[1823]&~m[1824]&m[1826]&~m[1827])|(m[1772]&m[1823]&~m[1824]&m[1826]&~m[1827])|(m[1772]&~m[1823]&m[1824]&m[1826]&~m[1827])|(~m[1772]&m[1823]&~m[1824]&~m[1826]&m[1827])|(~m[1772]&~m[1823]&m[1824]&~m[1826]&m[1827])|(m[1772]&m[1823]&m[1824]&~m[1826]&m[1827])|(~m[1772]&m[1823]&m[1824]&m[1826]&m[1827]))&UnbiasedRNG[435])|((m[1772]&~m[1823]&~m[1824]&m[1826]&~m[1827])|(~m[1772]&~m[1823]&~m[1824]&~m[1826]&m[1827])|(m[1772]&~m[1823]&~m[1824]&~m[1826]&m[1827])|(m[1772]&m[1823]&~m[1824]&~m[1826]&m[1827])|(m[1772]&~m[1823]&m[1824]&~m[1826]&m[1827])|(~m[1772]&~m[1823]&~m[1824]&m[1826]&m[1827])|(m[1772]&~m[1823]&~m[1824]&m[1826]&m[1827])|(~m[1772]&m[1823]&~m[1824]&m[1826]&m[1827])|(m[1772]&m[1823]&~m[1824]&m[1826]&m[1827])|(~m[1772]&~m[1823]&m[1824]&m[1826]&m[1827])|(m[1772]&~m[1823]&m[1824]&m[1826]&m[1827])|(m[1772]&m[1823]&m[1824]&m[1826]&m[1827]))):InitCond[1074];
    m[1830] = run?((((m[1777]&~m[1828]&~m[1829]&~m[1831]&~m[1832])|(~m[1777]&~m[1828]&~m[1829]&m[1831]&~m[1832])|(m[1777]&m[1828]&~m[1829]&m[1831]&~m[1832])|(m[1777]&~m[1828]&m[1829]&m[1831]&~m[1832])|(~m[1777]&m[1828]&~m[1829]&~m[1831]&m[1832])|(~m[1777]&~m[1828]&m[1829]&~m[1831]&m[1832])|(m[1777]&m[1828]&m[1829]&~m[1831]&m[1832])|(~m[1777]&m[1828]&m[1829]&m[1831]&m[1832]))&UnbiasedRNG[436])|((m[1777]&~m[1828]&~m[1829]&m[1831]&~m[1832])|(~m[1777]&~m[1828]&~m[1829]&~m[1831]&m[1832])|(m[1777]&~m[1828]&~m[1829]&~m[1831]&m[1832])|(m[1777]&m[1828]&~m[1829]&~m[1831]&m[1832])|(m[1777]&~m[1828]&m[1829]&~m[1831]&m[1832])|(~m[1777]&~m[1828]&~m[1829]&m[1831]&m[1832])|(m[1777]&~m[1828]&~m[1829]&m[1831]&m[1832])|(~m[1777]&m[1828]&~m[1829]&m[1831]&m[1832])|(m[1777]&m[1828]&~m[1829]&m[1831]&m[1832])|(~m[1777]&~m[1828]&m[1829]&m[1831]&m[1832])|(m[1777]&~m[1828]&m[1829]&m[1831]&m[1832])|(m[1777]&m[1828]&m[1829]&m[1831]&m[1832]))):InitCond[1075];
    m[1835] = run?((((m[1782]&~m[1833]&~m[1834]&~m[1836]&~m[1837])|(~m[1782]&~m[1833]&~m[1834]&m[1836]&~m[1837])|(m[1782]&m[1833]&~m[1834]&m[1836]&~m[1837])|(m[1782]&~m[1833]&m[1834]&m[1836]&~m[1837])|(~m[1782]&m[1833]&~m[1834]&~m[1836]&m[1837])|(~m[1782]&~m[1833]&m[1834]&~m[1836]&m[1837])|(m[1782]&m[1833]&m[1834]&~m[1836]&m[1837])|(~m[1782]&m[1833]&m[1834]&m[1836]&m[1837]))&UnbiasedRNG[437])|((m[1782]&~m[1833]&~m[1834]&m[1836]&~m[1837])|(~m[1782]&~m[1833]&~m[1834]&~m[1836]&m[1837])|(m[1782]&~m[1833]&~m[1834]&~m[1836]&m[1837])|(m[1782]&m[1833]&~m[1834]&~m[1836]&m[1837])|(m[1782]&~m[1833]&m[1834]&~m[1836]&m[1837])|(~m[1782]&~m[1833]&~m[1834]&m[1836]&m[1837])|(m[1782]&~m[1833]&~m[1834]&m[1836]&m[1837])|(~m[1782]&m[1833]&~m[1834]&m[1836]&m[1837])|(m[1782]&m[1833]&~m[1834]&m[1836]&m[1837])|(~m[1782]&~m[1833]&m[1834]&m[1836]&m[1837])|(m[1782]&~m[1833]&m[1834]&m[1836]&m[1837])|(m[1782]&m[1833]&m[1834]&m[1836]&m[1837]))):InitCond[1076];
    m[1840] = run?((((m[1787]&~m[1838]&~m[1839]&~m[1841]&~m[1842])|(~m[1787]&~m[1838]&~m[1839]&m[1841]&~m[1842])|(m[1787]&m[1838]&~m[1839]&m[1841]&~m[1842])|(m[1787]&~m[1838]&m[1839]&m[1841]&~m[1842])|(~m[1787]&m[1838]&~m[1839]&~m[1841]&m[1842])|(~m[1787]&~m[1838]&m[1839]&~m[1841]&m[1842])|(m[1787]&m[1838]&m[1839]&~m[1841]&m[1842])|(~m[1787]&m[1838]&m[1839]&m[1841]&m[1842]))&UnbiasedRNG[438])|((m[1787]&~m[1838]&~m[1839]&m[1841]&~m[1842])|(~m[1787]&~m[1838]&~m[1839]&~m[1841]&m[1842])|(m[1787]&~m[1838]&~m[1839]&~m[1841]&m[1842])|(m[1787]&m[1838]&~m[1839]&~m[1841]&m[1842])|(m[1787]&~m[1838]&m[1839]&~m[1841]&m[1842])|(~m[1787]&~m[1838]&~m[1839]&m[1841]&m[1842])|(m[1787]&~m[1838]&~m[1839]&m[1841]&m[1842])|(~m[1787]&m[1838]&~m[1839]&m[1841]&m[1842])|(m[1787]&m[1838]&~m[1839]&m[1841]&m[1842])|(~m[1787]&~m[1838]&m[1839]&m[1841]&m[1842])|(m[1787]&~m[1838]&m[1839]&m[1841]&m[1842])|(m[1787]&m[1838]&m[1839]&m[1841]&m[1842]))):InitCond[1077];
    m[1845] = run?((((m[1792]&~m[1843]&~m[1844]&~m[1846]&~m[1847])|(~m[1792]&~m[1843]&~m[1844]&m[1846]&~m[1847])|(m[1792]&m[1843]&~m[1844]&m[1846]&~m[1847])|(m[1792]&~m[1843]&m[1844]&m[1846]&~m[1847])|(~m[1792]&m[1843]&~m[1844]&~m[1846]&m[1847])|(~m[1792]&~m[1843]&m[1844]&~m[1846]&m[1847])|(m[1792]&m[1843]&m[1844]&~m[1846]&m[1847])|(~m[1792]&m[1843]&m[1844]&m[1846]&m[1847]))&UnbiasedRNG[439])|((m[1792]&~m[1843]&~m[1844]&m[1846]&~m[1847])|(~m[1792]&~m[1843]&~m[1844]&~m[1846]&m[1847])|(m[1792]&~m[1843]&~m[1844]&~m[1846]&m[1847])|(m[1792]&m[1843]&~m[1844]&~m[1846]&m[1847])|(m[1792]&~m[1843]&m[1844]&~m[1846]&m[1847])|(~m[1792]&~m[1843]&~m[1844]&m[1846]&m[1847])|(m[1792]&~m[1843]&~m[1844]&m[1846]&m[1847])|(~m[1792]&m[1843]&~m[1844]&m[1846]&m[1847])|(m[1792]&m[1843]&~m[1844]&m[1846]&m[1847])|(~m[1792]&~m[1843]&m[1844]&m[1846]&m[1847])|(m[1792]&~m[1843]&m[1844]&m[1846]&m[1847])|(m[1792]&m[1843]&m[1844]&m[1846]&m[1847]))):InitCond[1078];
    m[1850] = run?((((m[1797]&~m[1848]&~m[1849]&~m[1851]&~m[1852])|(~m[1797]&~m[1848]&~m[1849]&m[1851]&~m[1852])|(m[1797]&m[1848]&~m[1849]&m[1851]&~m[1852])|(m[1797]&~m[1848]&m[1849]&m[1851]&~m[1852])|(~m[1797]&m[1848]&~m[1849]&~m[1851]&m[1852])|(~m[1797]&~m[1848]&m[1849]&~m[1851]&m[1852])|(m[1797]&m[1848]&m[1849]&~m[1851]&m[1852])|(~m[1797]&m[1848]&m[1849]&m[1851]&m[1852]))&UnbiasedRNG[440])|((m[1797]&~m[1848]&~m[1849]&m[1851]&~m[1852])|(~m[1797]&~m[1848]&~m[1849]&~m[1851]&m[1852])|(m[1797]&~m[1848]&~m[1849]&~m[1851]&m[1852])|(m[1797]&m[1848]&~m[1849]&~m[1851]&m[1852])|(m[1797]&~m[1848]&m[1849]&~m[1851]&m[1852])|(~m[1797]&~m[1848]&~m[1849]&m[1851]&m[1852])|(m[1797]&~m[1848]&~m[1849]&m[1851]&m[1852])|(~m[1797]&m[1848]&~m[1849]&m[1851]&m[1852])|(m[1797]&m[1848]&~m[1849]&m[1851]&m[1852])|(~m[1797]&~m[1848]&m[1849]&m[1851]&m[1852])|(m[1797]&~m[1848]&m[1849]&m[1851]&m[1852])|(m[1797]&m[1848]&m[1849]&m[1851]&m[1852]))):InitCond[1079];
    m[1855] = run?((((m[1807]&~m[1853]&~m[1854]&~m[1856]&~m[1857])|(~m[1807]&~m[1853]&~m[1854]&m[1856]&~m[1857])|(m[1807]&m[1853]&~m[1854]&m[1856]&~m[1857])|(m[1807]&~m[1853]&m[1854]&m[1856]&~m[1857])|(~m[1807]&m[1853]&~m[1854]&~m[1856]&m[1857])|(~m[1807]&~m[1853]&m[1854]&~m[1856]&m[1857])|(m[1807]&m[1853]&m[1854]&~m[1856]&m[1857])|(~m[1807]&m[1853]&m[1854]&m[1856]&m[1857]))&UnbiasedRNG[441])|((m[1807]&~m[1853]&~m[1854]&m[1856]&~m[1857])|(~m[1807]&~m[1853]&~m[1854]&~m[1856]&m[1857])|(m[1807]&~m[1853]&~m[1854]&~m[1856]&m[1857])|(m[1807]&m[1853]&~m[1854]&~m[1856]&m[1857])|(m[1807]&~m[1853]&m[1854]&~m[1856]&m[1857])|(~m[1807]&~m[1853]&~m[1854]&m[1856]&m[1857])|(m[1807]&~m[1853]&~m[1854]&m[1856]&m[1857])|(~m[1807]&m[1853]&~m[1854]&m[1856]&m[1857])|(m[1807]&m[1853]&~m[1854]&m[1856]&m[1857])|(~m[1807]&~m[1853]&m[1854]&m[1856]&m[1857])|(m[1807]&~m[1853]&m[1854]&m[1856]&m[1857])|(m[1807]&m[1853]&m[1854]&m[1856]&m[1857]))):InitCond[1080];
    m[1860] = run?((((m[1812]&~m[1858]&~m[1859]&~m[1861]&~m[1862])|(~m[1812]&~m[1858]&~m[1859]&m[1861]&~m[1862])|(m[1812]&m[1858]&~m[1859]&m[1861]&~m[1862])|(m[1812]&~m[1858]&m[1859]&m[1861]&~m[1862])|(~m[1812]&m[1858]&~m[1859]&~m[1861]&m[1862])|(~m[1812]&~m[1858]&m[1859]&~m[1861]&m[1862])|(m[1812]&m[1858]&m[1859]&~m[1861]&m[1862])|(~m[1812]&m[1858]&m[1859]&m[1861]&m[1862]))&UnbiasedRNG[442])|((m[1812]&~m[1858]&~m[1859]&m[1861]&~m[1862])|(~m[1812]&~m[1858]&~m[1859]&~m[1861]&m[1862])|(m[1812]&~m[1858]&~m[1859]&~m[1861]&m[1862])|(m[1812]&m[1858]&~m[1859]&~m[1861]&m[1862])|(m[1812]&~m[1858]&m[1859]&~m[1861]&m[1862])|(~m[1812]&~m[1858]&~m[1859]&m[1861]&m[1862])|(m[1812]&~m[1858]&~m[1859]&m[1861]&m[1862])|(~m[1812]&m[1858]&~m[1859]&m[1861]&m[1862])|(m[1812]&m[1858]&~m[1859]&m[1861]&m[1862])|(~m[1812]&~m[1858]&m[1859]&m[1861]&m[1862])|(m[1812]&~m[1858]&m[1859]&m[1861]&m[1862])|(m[1812]&m[1858]&m[1859]&m[1861]&m[1862]))):InitCond[1081];
    m[1865] = run?((((m[1817]&~m[1863]&~m[1864]&~m[1866]&~m[1867])|(~m[1817]&~m[1863]&~m[1864]&m[1866]&~m[1867])|(m[1817]&m[1863]&~m[1864]&m[1866]&~m[1867])|(m[1817]&~m[1863]&m[1864]&m[1866]&~m[1867])|(~m[1817]&m[1863]&~m[1864]&~m[1866]&m[1867])|(~m[1817]&~m[1863]&m[1864]&~m[1866]&m[1867])|(m[1817]&m[1863]&m[1864]&~m[1866]&m[1867])|(~m[1817]&m[1863]&m[1864]&m[1866]&m[1867]))&UnbiasedRNG[443])|((m[1817]&~m[1863]&~m[1864]&m[1866]&~m[1867])|(~m[1817]&~m[1863]&~m[1864]&~m[1866]&m[1867])|(m[1817]&~m[1863]&~m[1864]&~m[1866]&m[1867])|(m[1817]&m[1863]&~m[1864]&~m[1866]&m[1867])|(m[1817]&~m[1863]&m[1864]&~m[1866]&m[1867])|(~m[1817]&~m[1863]&~m[1864]&m[1866]&m[1867])|(m[1817]&~m[1863]&~m[1864]&m[1866]&m[1867])|(~m[1817]&m[1863]&~m[1864]&m[1866]&m[1867])|(m[1817]&m[1863]&~m[1864]&m[1866]&m[1867])|(~m[1817]&~m[1863]&m[1864]&m[1866]&m[1867])|(m[1817]&~m[1863]&m[1864]&m[1866]&m[1867])|(m[1817]&m[1863]&m[1864]&m[1866]&m[1867]))):InitCond[1082];
    m[1870] = run?((((m[1822]&~m[1868]&~m[1869]&~m[1871]&~m[1872])|(~m[1822]&~m[1868]&~m[1869]&m[1871]&~m[1872])|(m[1822]&m[1868]&~m[1869]&m[1871]&~m[1872])|(m[1822]&~m[1868]&m[1869]&m[1871]&~m[1872])|(~m[1822]&m[1868]&~m[1869]&~m[1871]&m[1872])|(~m[1822]&~m[1868]&m[1869]&~m[1871]&m[1872])|(m[1822]&m[1868]&m[1869]&~m[1871]&m[1872])|(~m[1822]&m[1868]&m[1869]&m[1871]&m[1872]))&UnbiasedRNG[444])|((m[1822]&~m[1868]&~m[1869]&m[1871]&~m[1872])|(~m[1822]&~m[1868]&~m[1869]&~m[1871]&m[1872])|(m[1822]&~m[1868]&~m[1869]&~m[1871]&m[1872])|(m[1822]&m[1868]&~m[1869]&~m[1871]&m[1872])|(m[1822]&~m[1868]&m[1869]&~m[1871]&m[1872])|(~m[1822]&~m[1868]&~m[1869]&m[1871]&m[1872])|(m[1822]&~m[1868]&~m[1869]&m[1871]&m[1872])|(~m[1822]&m[1868]&~m[1869]&m[1871]&m[1872])|(m[1822]&m[1868]&~m[1869]&m[1871]&m[1872])|(~m[1822]&~m[1868]&m[1869]&m[1871]&m[1872])|(m[1822]&~m[1868]&m[1869]&m[1871]&m[1872])|(m[1822]&m[1868]&m[1869]&m[1871]&m[1872]))):InitCond[1083];
    m[1875] = run?((((m[1827]&~m[1873]&~m[1874]&~m[1876]&~m[1877])|(~m[1827]&~m[1873]&~m[1874]&m[1876]&~m[1877])|(m[1827]&m[1873]&~m[1874]&m[1876]&~m[1877])|(m[1827]&~m[1873]&m[1874]&m[1876]&~m[1877])|(~m[1827]&m[1873]&~m[1874]&~m[1876]&m[1877])|(~m[1827]&~m[1873]&m[1874]&~m[1876]&m[1877])|(m[1827]&m[1873]&m[1874]&~m[1876]&m[1877])|(~m[1827]&m[1873]&m[1874]&m[1876]&m[1877]))&UnbiasedRNG[445])|((m[1827]&~m[1873]&~m[1874]&m[1876]&~m[1877])|(~m[1827]&~m[1873]&~m[1874]&~m[1876]&m[1877])|(m[1827]&~m[1873]&~m[1874]&~m[1876]&m[1877])|(m[1827]&m[1873]&~m[1874]&~m[1876]&m[1877])|(m[1827]&~m[1873]&m[1874]&~m[1876]&m[1877])|(~m[1827]&~m[1873]&~m[1874]&m[1876]&m[1877])|(m[1827]&~m[1873]&~m[1874]&m[1876]&m[1877])|(~m[1827]&m[1873]&~m[1874]&m[1876]&m[1877])|(m[1827]&m[1873]&~m[1874]&m[1876]&m[1877])|(~m[1827]&~m[1873]&m[1874]&m[1876]&m[1877])|(m[1827]&~m[1873]&m[1874]&m[1876]&m[1877])|(m[1827]&m[1873]&m[1874]&m[1876]&m[1877]))):InitCond[1084];
    m[1880] = run?((((m[1832]&~m[1878]&~m[1879]&~m[1881]&~m[1882])|(~m[1832]&~m[1878]&~m[1879]&m[1881]&~m[1882])|(m[1832]&m[1878]&~m[1879]&m[1881]&~m[1882])|(m[1832]&~m[1878]&m[1879]&m[1881]&~m[1882])|(~m[1832]&m[1878]&~m[1879]&~m[1881]&m[1882])|(~m[1832]&~m[1878]&m[1879]&~m[1881]&m[1882])|(m[1832]&m[1878]&m[1879]&~m[1881]&m[1882])|(~m[1832]&m[1878]&m[1879]&m[1881]&m[1882]))&UnbiasedRNG[446])|((m[1832]&~m[1878]&~m[1879]&m[1881]&~m[1882])|(~m[1832]&~m[1878]&~m[1879]&~m[1881]&m[1882])|(m[1832]&~m[1878]&~m[1879]&~m[1881]&m[1882])|(m[1832]&m[1878]&~m[1879]&~m[1881]&m[1882])|(m[1832]&~m[1878]&m[1879]&~m[1881]&m[1882])|(~m[1832]&~m[1878]&~m[1879]&m[1881]&m[1882])|(m[1832]&~m[1878]&~m[1879]&m[1881]&m[1882])|(~m[1832]&m[1878]&~m[1879]&m[1881]&m[1882])|(m[1832]&m[1878]&~m[1879]&m[1881]&m[1882])|(~m[1832]&~m[1878]&m[1879]&m[1881]&m[1882])|(m[1832]&~m[1878]&m[1879]&m[1881]&m[1882])|(m[1832]&m[1878]&m[1879]&m[1881]&m[1882]))):InitCond[1085];
    m[1885] = run?((((m[1837]&~m[1883]&~m[1884]&~m[1886]&~m[1887])|(~m[1837]&~m[1883]&~m[1884]&m[1886]&~m[1887])|(m[1837]&m[1883]&~m[1884]&m[1886]&~m[1887])|(m[1837]&~m[1883]&m[1884]&m[1886]&~m[1887])|(~m[1837]&m[1883]&~m[1884]&~m[1886]&m[1887])|(~m[1837]&~m[1883]&m[1884]&~m[1886]&m[1887])|(m[1837]&m[1883]&m[1884]&~m[1886]&m[1887])|(~m[1837]&m[1883]&m[1884]&m[1886]&m[1887]))&UnbiasedRNG[447])|((m[1837]&~m[1883]&~m[1884]&m[1886]&~m[1887])|(~m[1837]&~m[1883]&~m[1884]&~m[1886]&m[1887])|(m[1837]&~m[1883]&~m[1884]&~m[1886]&m[1887])|(m[1837]&m[1883]&~m[1884]&~m[1886]&m[1887])|(m[1837]&~m[1883]&m[1884]&~m[1886]&m[1887])|(~m[1837]&~m[1883]&~m[1884]&m[1886]&m[1887])|(m[1837]&~m[1883]&~m[1884]&m[1886]&m[1887])|(~m[1837]&m[1883]&~m[1884]&m[1886]&m[1887])|(m[1837]&m[1883]&~m[1884]&m[1886]&m[1887])|(~m[1837]&~m[1883]&m[1884]&m[1886]&m[1887])|(m[1837]&~m[1883]&m[1884]&m[1886]&m[1887])|(m[1837]&m[1883]&m[1884]&m[1886]&m[1887]))):InitCond[1086];
    m[1890] = run?((((m[1842]&~m[1888]&~m[1889]&~m[1891]&~m[1892])|(~m[1842]&~m[1888]&~m[1889]&m[1891]&~m[1892])|(m[1842]&m[1888]&~m[1889]&m[1891]&~m[1892])|(m[1842]&~m[1888]&m[1889]&m[1891]&~m[1892])|(~m[1842]&m[1888]&~m[1889]&~m[1891]&m[1892])|(~m[1842]&~m[1888]&m[1889]&~m[1891]&m[1892])|(m[1842]&m[1888]&m[1889]&~m[1891]&m[1892])|(~m[1842]&m[1888]&m[1889]&m[1891]&m[1892]))&UnbiasedRNG[448])|((m[1842]&~m[1888]&~m[1889]&m[1891]&~m[1892])|(~m[1842]&~m[1888]&~m[1889]&~m[1891]&m[1892])|(m[1842]&~m[1888]&~m[1889]&~m[1891]&m[1892])|(m[1842]&m[1888]&~m[1889]&~m[1891]&m[1892])|(m[1842]&~m[1888]&m[1889]&~m[1891]&m[1892])|(~m[1842]&~m[1888]&~m[1889]&m[1891]&m[1892])|(m[1842]&~m[1888]&~m[1889]&m[1891]&m[1892])|(~m[1842]&m[1888]&~m[1889]&m[1891]&m[1892])|(m[1842]&m[1888]&~m[1889]&m[1891]&m[1892])|(~m[1842]&~m[1888]&m[1889]&m[1891]&m[1892])|(m[1842]&~m[1888]&m[1889]&m[1891]&m[1892])|(m[1842]&m[1888]&m[1889]&m[1891]&m[1892]))):InitCond[1087];
    m[1895] = run?((((m[1847]&~m[1893]&~m[1894]&~m[1896]&~m[1897])|(~m[1847]&~m[1893]&~m[1894]&m[1896]&~m[1897])|(m[1847]&m[1893]&~m[1894]&m[1896]&~m[1897])|(m[1847]&~m[1893]&m[1894]&m[1896]&~m[1897])|(~m[1847]&m[1893]&~m[1894]&~m[1896]&m[1897])|(~m[1847]&~m[1893]&m[1894]&~m[1896]&m[1897])|(m[1847]&m[1893]&m[1894]&~m[1896]&m[1897])|(~m[1847]&m[1893]&m[1894]&m[1896]&m[1897]))&UnbiasedRNG[449])|((m[1847]&~m[1893]&~m[1894]&m[1896]&~m[1897])|(~m[1847]&~m[1893]&~m[1894]&~m[1896]&m[1897])|(m[1847]&~m[1893]&~m[1894]&~m[1896]&m[1897])|(m[1847]&m[1893]&~m[1894]&~m[1896]&m[1897])|(m[1847]&~m[1893]&m[1894]&~m[1896]&m[1897])|(~m[1847]&~m[1893]&~m[1894]&m[1896]&m[1897])|(m[1847]&~m[1893]&~m[1894]&m[1896]&m[1897])|(~m[1847]&m[1893]&~m[1894]&m[1896]&m[1897])|(m[1847]&m[1893]&~m[1894]&m[1896]&m[1897])|(~m[1847]&~m[1893]&m[1894]&m[1896]&m[1897])|(m[1847]&~m[1893]&m[1894]&m[1896]&m[1897])|(m[1847]&m[1893]&m[1894]&m[1896]&m[1897]))):InitCond[1088];
    m[1900] = run?((((m[1852]&~m[1898]&~m[1899]&~m[1901]&~m[1902])|(~m[1852]&~m[1898]&~m[1899]&m[1901]&~m[1902])|(m[1852]&m[1898]&~m[1899]&m[1901]&~m[1902])|(m[1852]&~m[1898]&m[1899]&m[1901]&~m[1902])|(~m[1852]&m[1898]&~m[1899]&~m[1901]&m[1902])|(~m[1852]&~m[1898]&m[1899]&~m[1901]&m[1902])|(m[1852]&m[1898]&m[1899]&~m[1901]&m[1902])|(~m[1852]&m[1898]&m[1899]&m[1901]&m[1902]))&UnbiasedRNG[450])|((m[1852]&~m[1898]&~m[1899]&m[1901]&~m[1902])|(~m[1852]&~m[1898]&~m[1899]&~m[1901]&m[1902])|(m[1852]&~m[1898]&~m[1899]&~m[1901]&m[1902])|(m[1852]&m[1898]&~m[1899]&~m[1901]&m[1902])|(m[1852]&~m[1898]&m[1899]&~m[1901]&m[1902])|(~m[1852]&~m[1898]&~m[1899]&m[1901]&m[1902])|(m[1852]&~m[1898]&~m[1899]&m[1901]&m[1902])|(~m[1852]&m[1898]&~m[1899]&m[1901]&m[1902])|(m[1852]&m[1898]&~m[1899]&m[1901]&m[1902])|(~m[1852]&~m[1898]&m[1899]&m[1901]&m[1902])|(m[1852]&~m[1898]&m[1899]&m[1901]&m[1902])|(m[1852]&m[1898]&m[1899]&m[1901]&m[1902]))):InitCond[1089];
    m[1905] = run?((((m[1862]&~m[1903]&~m[1904]&~m[1906]&~m[1907])|(~m[1862]&~m[1903]&~m[1904]&m[1906]&~m[1907])|(m[1862]&m[1903]&~m[1904]&m[1906]&~m[1907])|(m[1862]&~m[1903]&m[1904]&m[1906]&~m[1907])|(~m[1862]&m[1903]&~m[1904]&~m[1906]&m[1907])|(~m[1862]&~m[1903]&m[1904]&~m[1906]&m[1907])|(m[1862]&m[1903]&m[1904]&~m[1906]&m[1907])|(~m[1862]&m[1903]&m[1904]&m[1906]&m[1907]))&UnbiasedRNG[451])|((m[1862]&~m[1903]&~m[1904]&m[1906]&~m[1907])|(~m[1862]&~m[1903]&~m[1904]&~m[1906]&m[1907])|(m[1862]&~m[1903]&~m[1904]&~m[1906]&m[1907])|(m[1862]&m[1903]&~m[1904]&~m[1906]&m[1907])|(m[1862]&~m[1903]&m[1904]&~m[1906]&m[1907])|(~m[1862]&~m[1903]&~m[1904]&m[1906]&m[1907])|(m[1862]&~m[1903]&~m[1904]&m[1906]&m[1907])|(~m[1862]&m[1903]&~m[1904]&m[1906]&m[1907])|(m[1862]&m[1903]&~m[1904]&m[1906]&m[1907])|(~m[1862]&~m[1903]&m[1904]&m[1906]&m[1907])|(m[1862]&~m[1903]&m[1904]&m[1906]&m[1907])|(m[1862]&m[1903]&m[1904]&m[1906]&m[1907]))):InitCond[1090];
    m[1910] = run?((((m[1867]&~m[1908]&~m[1909]&~m[1911]&~m[1912])|(~m[1867]&~m[1908]&~m[1909]&m[1911]&~m[1912])|(m[1867]&m[1908]&~m[1909]&m[1911]&~m[1912])|(m[1867]&~m[1908]&m[1909]&m[1911]&~m[1912])|(~m[1867]&m[1908]&~m[1909]&~m[1911]&m[1912])|(~m[1867]&~m[1908]&m[1909]&~m[1911]&m[1912])|(m[1867]&m[1908]&m[1909]&~m[1911]&m[1912])|(~m[1867]&m[1908]&m[1909]&m[1911]&m[1912]))&UnbiasedRNG[452])|((m[1867]&~m[1908]&~m[1909]&m[1911]&~m[1912])|(~m[1867]&~m[1908]&~m[1909]&~m[1911]&m[1912])|(m[1867]&~m[1908]&~m[1909]&~m[1911]&m[1912])|(m[1867]&m[1908]&~m[1909]&~m[1911]&m[1912])|(m[1867]&~m[1908]&m[1909]&~m[1911]&m[1912])|(~m[1867]&~m[1908]&~m[1909]&m[1911]&m[1912])|(m[1867]&~m[1908]&~m[1909]&m[1911]&m[1912])|(~m[1867]&m[1908]&~m[1909]&m[1911]&m[1912])|(m[1867]&m[1908]&~m[1909]&m[1911]&m[1912])|(~m[1867]&~m[1908]&m[1909]&m[1911]&m[1912])|(m[1867]&~m[1908]&m[1909]&m[1911]&m[1912])|(m[1867]&m[1908]&m[1909]&m[1911]&m[1912]))):InitCond[1091];
    m[1915] = run?((((m[1872]&~m[1913]&~m[1914]&~m[1916]&~m[1917])|(~m[1872]&~m[1913]&~m[1914]&m[1916]&~m[1917])|(m[1872]&m[1913]&~m[1914]&m[1916]&~m[1917])|(m[1872]&~m[1913]&m[1914]&m[1916]&~m[1917])|(~m[1872]&m[1913]&~m[1914]&~m[1916]&m[1917])|(~m[1872]&~m[1913]&m[1914]&~m[1916]&m[1917])|(m[1872]&m[1913]&m[1914]&~m[1916]&m[1917])|(~m[1872]&m[1913]&m[1914]&m[1916]&m[1917]))&UnbiasedRNG[453])|((m[1872]&~m[1913]&~m[1914]&m[1916]&~m[1917])|(~m[1872]&~m[1913]&~m[1914]&~m[1916]&m[1917])|(m[1872]&~m[1913]&~m[1914]&~m[1916]&m[1917])|(m[1872]&m[1913]&~m[1914]&~m[1916]&m[1917])|(m[1872]&~m[1913]&m[1914]&~m[1916]&m[1917])|(~m[1872]&~m[1913]&~m[1914]&m[1916]&m[1917])|(m[1872]&~m[1913]&~m[1914]&m[1916]&m[1917])|(~m[1872]&m[1913]&~m[1914]&m[1916]&m[1917])|(m[1872]&m[1913]&~m[1914]&m[1916]&m[1917])|(~m[1872]&~m[1913]&m[1914]&m[1916]&m[1917])|(m[1872]&~m[1913]&m[1914]&m[1916]&m[1917])|(m[1872]&m[1913]&m[1914]&m[1916]&m[1917]))):InitCond[1092];
    m[1920] = run?((((m[1877]&~m[1918]&~m[1919]&~m[1921]&~m[1922])|(~m[1877]&~m[1918]&~m[1919]&m[1921]&~m[1922])|(m[1877]&m[1918]&~m[1919]&m[1921]&~m[1922])|(m[1877]&~m[1918]&m[1919]&m[1921]&~m[1922])|(~m[1877]&m[1918]&~m[1919]&~m[1921]&m[1922])|(~m[1877]&~m[1918]&m[1919]&~m[1921]&m[1922])|(m[1877]&m[1918]&m[1919]&~m[1921]&m[1922])|(~m[1877]&m[1918]&m[1919]&m[1921]&m[1922]))&UnbiasedRNG[454])|((m[1877]&~m[1918]&~m[1919]&m[1921]&~m[1922])|(~m[1877]&~m[1918]&~m[1919]&~m[1921]&m[1922])|(m[1877]&~m[1918]&~m[1919]&~m[1921]&m[1922])|(m[1877]&m[1918]&~m[1919]&~m[1921]&m[1922])|(m[1877]&~m[1918]&m[1919]&~m[1921]&m[1922])|(~m[1877]&~m[1918]&~m[1919]&m[1921]&m[1922])|(m[1877]&~m[1918]&~m[1919]&m[1921]&m[1922])|(~m[1877]&m[1918]&~m[1919]&m[1921]&m[1922])|(m[1877]&m[1918]&~m[1919]&m[1921]&m[1922])|(~m[1877]&~m[1918]&m[1919]&m[1921]&m[1922])|(m[1877]&~m[1918]&m[1919]&m[1921]&m[1922])|(m[1877]&m[1918]&m[1919]&m[1921]&m[1922]))):InitCond[1093];
    m[1925] = run?((((m[1882]&~m[1923]&~m[1924]&~m[1926]&~m[1927])|(~m[1882]&~m[1923]&~m[1924]&m[1926]&~m[1927])|(m[1882]&m[1923]&~m[1924]&m[1926]&~m[1927])|(m[1882]&~m[1923]&m[1924]&m[1926]&~m[1927])|(~m[1882]&m[1923]&~m[1924]&~m[1926]&m[1927])|(~m[1882]&~m[1923]&m[1924]&~m[1926]&m[1927])|(m[1882]&m[1923]&m[1924]&~m[1926]&m[1927])|(~m[1882]&m[1923]&m[1924]&m[1926]&m[1927]))&UnbiasedRNG[455])|((m[1882]&~m[1923]&~m[1924]&m[1926]&~m[1927])|(~m[1882]&~m[1923]&~m[1924]&~m[1926]&m[1927])|(m[1882]&~m[1923]&~m[1924]&~m[1926]&m[1927])|(m[1882]&m[1923]&~m[1924]&~m[1926]&m[1927])|(m[1882]&~m[1923]&m[1924]&~m[1926]&m[1927])|(~m[1882]&~m[1923]&~m[1924]&m[1926]&m[1927])|(m[1882]&~m[1923]&~m[1924]&m[1926]&m[1927])|(~m[1882]&m[1923]&~m[1924]&m[1926]&m[1927])|(m[1882]&m[1923]&~m[1924]&m[1926]&m[1927])|(~m[1882]&~m[1923]&m[1924]&m[1926]&m[1927])|(m[1882]&~m[1923]&m[1924]&m[1926]&m[1927])|(m[1882]&m[1923]&m[1924]&m[1926]&m[1927]))):InitCond[1094];
    m[1930] = run?((((m[1887]&~m[1928]&~m[1929]&~m[1931]&~m[1932])|(~m[1887]&~m[1928]&~m[1929]&m[1931]&~m[1932])|(m[1887]&m[1928]&~m[1929]&m[1931]&~m[1932])|(m[1887]&~m[1928]&m[1929]&m[1931]&~m[1932])|(~m[1887]&m[1928]&~m[1929]&~m[1931]&m[1932])|(~m[1887]&~m[1928]&m[1929]&~m[1931]&m[1932])|(m[1887]&m[1928]&m[1929]&~m[1931]&m[1932])|(~m[1887]&m[1928]&m[1929]&m[1931]&m[1932]))&UnbiasedRNG[456])|((m[1887]&~m[1928]&~m[1929]&m[1931]&~m[1932])|(~m[1887]&~m[1928]&~m[1929]&~m[1931]&m[1932])|(m[1887]&~m[1928]&~m[1929]&~m[1931]&m[1932])|(m[1887]&m[1928]&~m[1929]&~m[1931]&m[1932])|(m[1887]&~m[1928]&m[1929]&~m[1931]&m[1932])|(~m[1887]&~m[1928]&~m[1929]&m[1931]&m[1932])|(m[1887]&~m[1928]&~m[1929]&m[1931]&m[1932])|(~m[1887]&m[1928]&~m[1929]&m[1931]&m[1932])|(m[1887]&m[1928]&~m[1929]&m[1931]&m[1932])|(~m[1887]&~m[1928]&m[1929]&m[1931]&m[1932])|(m[1887]&~m[1928]&m[1929]&m[1931]&m[1932])|(m[1887]&m[1928]&m[1929]&m[1931]&m[1932]))):InitCond[1095];
    m[1935] = run?((((m[1892]&~m[1933]&~m[1934]&~m[1936]&~m[1937])|(~m[1892]&~m[1933]&~m[1934]&m[1936]&~m[1937])|(m[1892]&m[1933]&~m[1934]&m[1936]&~m[1937])|(m[1892]&~m[1933]&m[1934]&m[1936]&~m[1937])|(~m[1892]&m[1933]&~m[1934]&~m[1936]&m[1937])|(~m[1892]&~m[1933]&m[1934]&~m[1936]&m[1937])|(m[1892]&m[1933]&m[1934]&~m[1936]&m[1937])|(~m[1892]&m[1933]&m[1934]&m[1936]&m[1937]))&UnbiasedRNG[457])|((m[1892]&~m[1933]&~m[1934]&m[1936]&~m[1937])|(~m[1892]&~m[1933]&~m[1934]&~m[1936]&m[1937])|(m[1892]&~m[1933]&~m[1934]&~m[1936]&m[1937])|(m[1892]&m[1933]&~m[1934]&~m[1936]&m[1937])|(m[1892]&~m[1933]&m[1934]&~m[1936]&m[1937])|(~m[1892]&~m[1933]&~m[1934]&m[1936]&m[1937])|(m[1892]&~m[1933]&~m[1934]&m[1936]&m[1937])|(~m[1892]&m[1933]&~m[1934]&m[1936]&m[1937])|(m[1892]&m[1933]&~m[1934]&m[1936]&m[1937])|(~m[1892]&~m[1933]&m[1934]&m[1936]&m[1937])|(m[1892]&~m[1933]&m[1934]&m[1936]&m[1937])|(m[1892]&m[1933]&m[1934]&m[1936]&m[1937]))):InitCond[1096];
    m[1940] = run?((((m[1897]&~m[1938]&~m[1939]&~m[1941]&~m[1942])|(~m[1897]&~m[1938]&~m[1939]&m[1941]&~m[1942])|(m[1897]&m[1938]&~m[1939]&m[1941]&~m[1942])|(m[1897]&~m[1938]&m[1939]&m[1941]&~m[1942])|(~m[1897]&m[1938]&~m[1939]&~m[1941]&m[1942])|(~m[1897]&~m[1938]&m[1939]&~m[1941]&m[1942])|(m[1897]&m[1938]&m[1939]&~m[1941]&m[1942])|(~m[1897]&m[1938]&m[1939]&m[1941]&m[1942]))&UnbiasedRNG[458])|((m[1897]&~m[1938]&~m[1939]&m[1941]&~m[1942])|(~m[1897]&~m[1938]&~m[1939]&~m[1941]&m[1942])|(m[1897]&~m[1938]&~m[1939]&~m[1941]&m[1942])|(m[1897]&m[1938]&~m[1939]&~m[1941]&m[1942])|(m[1897]&~m[1938]&m[1939]&~m[1941]&m[1942])|(~m[1897]&~m[1938]&~m[1939]&m[1941]&m[1942])|(m[1897]&~m[1938]&~m[1939]&m[1941]&m[1942])|(~m[1897]&m[1938]&~m[1939]&m[1941]&m[1942])|(m[1897]&m[1938]&~m[1939]&m[1941]&m[1942])|(~m[1897]&~m[1938]&m[1939]&m[1941]&m[1942])|(m[1897]&~m[1938]&m[1939]&m[1941]&m[1942])|(m[1897]&m[1938]&m[1939]&m[1941]&m[1942]))):InitCond[1097];
    m[1945] = run?((((m[1902]&~m[1943]&~m[1944]&~m[1946]&~m[1947])|(~m[1902]&~m[1943]&~m[1944]&m[1946]&~m[1947])|(m[1902]&m[1943]&~m[1944]&m[1946]&~m[1947])|(m[1902]&~m[1943]&m[1944]&m[1946]&~m[1947])|(~m[1902]&m[1943]&~m[1944]&~m[1946]&m[1947])|(~m[1902]&~m[1943]&m[1944]&~m[1946]&m[1947])|(m[1902]&m[1943]&m[1944]&~m[1946]&m[1947])|(~m[1902]&m[1943]&m[1944]&m[1946]&m[1947]))&UnbiasedRNG[459])|((m[1902]&~m[1943]&~m[1944]&m[1946]&~m[1947])|(~m[1902]&~m[1943]&~m[1944]&~m[1946]&m[1947])|(m[1902]&~m[1943]&~m[1944]&~m[1946]&m[1947])|(m[1902]&m[1943]&~m[1944]&~m[1946]&m[1947])|(m[1902]&~m[1943]&m[1944]&~m[1946]&m[1947])|(~m[1902]&~m[1943]&~m[1944]&m[1946]&m[1947])|(m[1902]&~m[1943]&~m[1944]&m[1946]&m[1947])|(~m[1902]&m[1943]&~m[1944]&m[1946]&m[1947])|(m[1902]&m[1943]&~m[1944]&m[1946]&m[1947])|(~m[1902]&~m[1943]&m[1944]&m[1946]&m[1947])|(m[1902]&~m[1943]&m[1944]&m[1946]&m[1947])|(m[1902]&m[1943]&m[1944]&m[1946]&m[1947]))):InitCond[1098];
    m[1950] = run?((((m[1912]&~m[1948]&~m[1949]&~m[1951]&~m[1952])|(~m[1912]&~m[1948]&~m[1949]&m[1951]&~m[1952])|(m[1912]&m[1948]&~m[1949]&m[1951]&~m[1952])|(m[1912]&~m[1948]&m[1949]&m[1951]&~m[1952])|(~m[1912]&m[1948]&~m[1949]&~m[1951]&m[1952])|(~m[1912]&~m[1948]&m[1949]&~m[1951]&m[1952])|(m[1912]&m[1948]&m[1949]&~m[1951]&m[1952])|(~m[1912]&m[1948]&m[1949]&m[1951]&m[1952]))&UnbiasedRNG[460])|((m[1912]&~m[1948]&~m[1949]&m[1951]&~m[1952])|(~m[1912]&~m[1948]&~m[1949]&~m[1951]&m[1952])|(m[1912]&~m[1948]&~m[1949]&~m[1951]&m[1952])|(m[1912]&m[1948]&~m[1949]&~m[1951]&m[1952])|(m[1912]&~m[1948]&m[1949]&~m[1951]&m[1952])|(~m[1912]&~m[1948]&~m[1949]&m[1951]&m[1952])|(m[1912]&~m[1948]&~m[1949]&m[1951]&m[1952])|(~m[1912]&m[1948]&~m[1949]&m[1951]&m[1952])|(m[1912]&m[1948]&~m[1949]&m[1951]&m[1952])|(~m[1912]&~m[1948]&m[1949]&m[1951]&m[1952])|(m[1912]&~m[1948]&m[1949]&m[1951]&m[1952])|(m[1912]&m[1948]&m[1949]&m[1951]&m[1952]))):InitCond[1099];
    m[1955] = run?((((m[1917]&~m[1953]&~m[1954]&~m[1956]&~m[1957])|(~m[1917]&~m[1953]&~m[1954]&m[1956]&~m[1957])|(m[1917]&m[1953]&~m[1954]&m[1956]&~m[1957])|(m[1917]&~m[1953]&m[1954]&m[1956]&~m[1957])|(~m[1917]&m[1953]&~m[1954]&~m[1956]&m[1957])|(~m[1917]&~m[1953]&m[1954]&~m[1956]&m[1957])|(m[1917]&m[1953]&m[1954]&~m[1956]&m[1957])|(~m[1917]&m[1953]&m[1954]&m[1956]&m[1957]))&UnbiasedRNG[461])|((m[1917]&~m[1953]&~m[1954]&m[1956]&~m[1957])|(~m[1917]&~m[1953]&~m[1954]&~m[1956]&m[1957])|(m[1917]&~m[1953]&~m[1954]&~m[1956]&m[1957])|(m[1917]&m[1953]&~m[1954]&~m[1956]&m[1957])|(m[1917]&~m[1953]&m[1954]&~m[1956]&m[1957])|(~m[1917]&~m[1953]&~m[1954]&m[1956]&m[1957])|(m[1917]&~m[1953]&~m[1954]&m[1956]&m[1957])|(~m[1917]&m[1953]&~m[1954]&m[1956]&m[1957])|(m[1917]&m[1953]&~m[1954]&m[1956]&m[1957])|(~m[1917]&~m[1953]&m[1954]&m[1956]&m[1957])|(m[1917]&~m[1953]&m[1954]&m[1956]&m[1957])|(m[1917]&m[1953]&m[1954]&m[1956]&m[1957]))):InitCond[1100];
    m[1960] = run?((((m[1922]&~m[1958]&~m[1959]&~m[1961]&~m[1962])|(~m[1922]&~m[1958]&~m[1959]&m[1961]&~m[1962])|(m[1922]&m[1958]&~m[1959]&m[1961]&~m[1962])|(m[1922]&~m[1958]&m[1959]&m[1961]&~m[1962])|(~m[1922]&m[1958]&~m[1959]&~m[1961]&m[1962])|(~m[1922]&~m[1958]&m[1959]&~m[1961]&m[1962])|(m[1922]&m[1958]&m[1959]&~m[1961]&m[1962])|(~m[1922]&m[1958]&m[1959]&m[1961]&m[1962]))&UnbiasedRNG[462])|((m[1922]&~m[1958]&~m[1959]&m[1961]&~m[1962])|(~m[1922]&~m[1958]&~m[1959]&~m[1961]&m[1962])|(m[1922]&~m[1958]&~m[1959]&~m[1961]&m[1962])|(m[1922]&m[1958]&~m[1959]&~m[1961]&m[1962])|(m[1922]&~m[1958]&m[1959]&~m[1961]&m[1962])|(~m[1922]&~m[1958]&~m[1959]&m[1961]&m[1962])|(m[1922]&~m[1958]&~m[1959]&m[1961]&m[1962])|(~m[1922]&m[1958]&~m[1959]&m[1961]&m[1962])|(m[1922]&m[1958]&~m[1959]&m[1961]&m[1962])|(~m[1922]&~m[1958]&m[1959]&m[1961]&m[1962])|(m[1922]&~m[1958]&m[1959]&m[1961]&m[1962])|(m[1922]&m[1958]&m[1959]&m[1961]&m[1962]))):InitCond[1101];
    m[1965] = run?((((m[1927]&~m[1963]&~m[1964]&~m[1966]&~m[1967])|(~m[1927]&~m[1963]&~m[1964]&m[1966]&~m[1967])|(m[1927]&m[1963]&~m[1964]&m[1966]&~m[1967])|(m[1927]&~m[1963]&m[1964]&m[1966]&~m[1967])|(~m[1927]&m[1963]&~m[1964]&~m[1966]&m[1967])|(~m[1927]&~m[1963]&m[1964]&~m[1966]&m[1967])|(m[1927]&m[1963]&m[1964]&~m[1966]&m[1967])|(~m[1927]&m[1963]&m[1964]&m[1966]&m[1967]))&UnbiasedRNG[463])|((m[1927]&~m[1963]&~m[1964]&m[1966]&~m[1967])|(~m[1927]&~m[1963]&~m[1964]&~m[1966]&m[1967])|(m[1927]&~m[1963]&~m[1964]&~m[1966]&m[1967])|(m[1927]&m[1963]&~m[1964]&~m[1966]&m[1967])|(m[1927]&~m[1963]&m[1964]&~m[1966]&m[1967])|(~m[1927]&~m[1963]&~m[1964]&m[1966]&m[1967])|(m[1927]&~m[1963]&~m[1964]&m[1966]&m[1967])|(~m[1927]&m[1963]&~m[1964]&m[1966]&m[1967])|(m[1927]&m[1963]&~m[1964]&m[1966]&m[1967])|(~m[1927]&~m[1963]&m[1964]&m[1966]&m[1967])|(m[1927]&~m[1963]&m[1964]&m[1966]&m[1967])|(m[1927]&m[1963]&m[1964]&m[1966]&m[1967]))):InitCond[1102];
    m[1970] = run?((((m[1932]&~m[1968]&~m[1969]&~m[1971]&~m[1972])|(~m[1932]&~m[1968]&~m[1969]&m[1971]&~m[1972])|(m[1932]&m[1968]&~m[1969]&m[1971]&~m[1972])|(m[1932]&~m[1968]&m[1969]&m[1971]&~m[1972])|(~m[1932]&m[1968]&~m[1969]&~m[1971]&m[1972])|(~m[1932]&~m[1968]&m[1969]&~m[1971]&m[1972])|(m[1932]&m[1968]&m[1969]&~m[1971]&m[1972])|(~m[1932]&m[1968]&m[1969]&m[1971]&m[1972]))&UnbiasedRNG[464])|((m[1932]&~m[1968]&~m[1969]&m[1971]&~m[1972])|(~m[1932]&~m[1968]&~m[1969]&~m[1971]&m[1972])|(m[1932]&~m[1968]&~m[1969]&~m[1971]&m[1972])|(m[1932]&m[1968]&~m[1969]&~m[1971]&m[1972])|(m[1932]&~m[1968]&m[1969]&~m[1971]&m[1972])|(~m[1932]&~m[1968]&~m[1969]&m[1971]&m[1972])|(m[1932]&~m[1968]&~m[1969]&m[1971]&m[1972])|(~m[1932]&m[1968]&~m[1969]&m[1971]&m[1972])|(m[1932]&m[1968]&~m[1969]&m[1971]&m[1972])|(~m[1932]&~m[1968]&m[1969]&m[1971]&m[1972])|(m[1932]&~m[1968]&m[1969]&m[1971]&m[1972])|(m[1932]&m[1968]&m[1969]&m[1971]&m[1972]))):InitCond[1103];
    m[1975] = run?((((m[1937]&~m[1973]&~m[1974]&~m[1976]&~m[1977])|(~m[1937]&~m[1973]&~m[1974]&m[1976]&~m[1977])|(m[1937]&m[1973]&~m[1974]&m[1976]&~m[1977])|(m[1937]&~m[1973]&m[1974]&m[1976]&~m[1977])|(~m[1937]&m[1973]&~m[1974]&~m[1976]&m[1977])|(~m[1937]&~m[1973]&m[1974]&~m[1976]&m[1977])|(m[1937]&m[1973]&m[1974]&~m[1976]&m[1977])|(~m[1937]&m[1973]&m[1974]&m[1976]&m[1977]))&UnbiasedRNG[465])|((m[1937]&~m[1973]&~m[1974]&m[1976]&~m[1977])|(~m[1937]&~m[1973]&~m[1974]&~m[1976]&m[1977])|(m[1937]&~m[1973]&~m[1974]&~m[1976]&m[1977])|(m[1937]&m[1973]&~m[1974]&~m[1976]&m[1977])|(m[1937]&~m[1973]&m[1974]&~m[1976]&m[1977])|(~m[1937]&~m[1973]&~m[1974]&m[1976]&m[1977])|(m[1937]&~m[1973]&~m[1974]&m[1976]&m[1977])|(~m[1937]&m[1973]&~m[1974]&m[1976]&m[1977])|(m[1937]&m[1973]&~m[1974]&m[1976]&m[1977])|(~m[1937]&~m[1973]&m[1974]&m[1976]&m[1977])|(m[1937]&~m[1973]&m[1974]&m[1976]&m[1977])|(m[1937]&m[1973]&m[1974]&m[1976]&m[1977]))):InitCond[1104];
    m[1980] = run?((((m[1942]&~m[1978]&~m[1979]&~m[1981]&~m[1982])|(~m[1942]&~m[1978]&~m[1979]&m[1981]&~m[1982])|(m[1942]&m[1978]&~m[1979]&m[1981]&~m[1982])|(m[1942]&~m[1978]&m[1979]&m[1981]&~m[1982])|(~m[1942]&m[1978]&~m[1979]&~m[1981]&m[1982])|(~m[1942]&~m[1978]&m[1979]&~m[1981]&m[1982])|(m[1942]&m[1978]&m[1979]&~m[1981]&m[1982])|(~m[1942]&m[1978]&m[1979]&m[1981]&m[1982]))&UnbiasedRNG[466])|((m[1942]&~m[1978]&~m[1979]&m[1981]&~m[1982])|(~m[1942]&~m[1978]&~m[1979]&~m[1981]&m[1982])|(m[1942]&~m[1978]&~m[1979]&~m[1981]&m[1982])|(m[1942]&m[1978]&~m[1979]&~m[1981]&m[1982])|(m[1942]&~m[1978]&m[1979]&~m[1981]&m[1982])|(~m[1942]&~m[1978]&~m[1979]&m[1981]&m[1982])|(m[1942]&~m[1978]&~m[1979]&m[1981]&m[1982])|(~m[1942]&m[1978]&~m[1979]&m[1981]&m[1982])|(m[1942]&m[1978]&~m[1979]&m[1981]&m[1982])|(~m[1942]&~m[1978]&m[1979]&m[1981]&m[1982])|(m[1942]&~m[1978]&m[1979]&m[1981]&m[1982])|(m[1942]&m[1978]&m[1979]&m[1981]&m[1982]))):InitCond[1105];
    m[1985] = run?((((m[1947]&~m[1983]&~m[1984]&~m[1986]&~m[1987])|(~m[1947]&~m[1983]&~m[1984]&m[1986]&~m[1987])|(m[1947]&m[1983]&~m[1984]&m[1986]&~m[1987])|(m[1947]&~m[1983]&m[1984]&m[1986]&~m[1987])|(~m[1947]&m[1983]&~m[1984]&~m[1986]&m[1987])|(~m[1947]&~m[1983]&m[1984]&~m[1986]&m[1987])|(m[1947]&m[1983]&m[1984]&~m[1986]&m[1987])|(~m[1947]&m[1983]&m[1984]&m[1986]&m[1987]))&UnbiasedRNG[467])|((m[1947]&~m[1983]&~m[1984]&m[1986]&~m[1987])|(~m[1947]&~m[1983]&~m[1984]&~m[1986]&m[1987])|(m[1947]&~m[1983]&~m[1984]&~m[1986]&m[1987])|(m[1947]&m[1983]&~m[1984]&~m[1986]&m[1987])|(m[1947]&~m[1983]&m[1984]&~m[1986]&m[1987])|(~m[1947]&~m[1983]&~m[1984]&m[1986]&m[1987])|(m[1947]&~m[1983]&~m[1984]&m[1986]&m[1987])|(~m[1947]&m[1983]&~m[1984]&m[1986]&m[1987])|(m[1947]&m[1983]&~m[1984]&m[1986]&m[1987])|(~m[1947]&~m[1983]&m[1984]&m[1986]&m[1987])|(m[1947]&~m[1983]&m[1984]&m[1986]&m[1987])|(m[1947]&m[1983]&m[1984]&m[1986]&m[1987]))):InitCond[1106];
    m[1990] = run?((((m[1957]&~m[1988]&~m[1989]&~m[1991]&~m[1992])|(~m[1957]&~m[1988]&~m[1989]&m[1991]&~m[1992])|(m[1957]&m[1988]&~m[1989]&m[1991]&~m[1992])|(m[1957]&~m[1988]&m[1989]&m[1991]&~m[1992])|(~m[1957]&m[1988]&~m[1989]&~m[1991]&m[1992])|(~m[1957]&~m[1988]&m[1989]&~m[1991]&m[1992])|(m[1957]&m[1988]&m[1989]&~m[1991]&m[1992])|(~m[1957]&m[1988]&m[1989]&m[1991]&m[1992]))&UnbiasedRNG[468])|((m[1957]&~m[1988]&~m[1989]&m[1991]&~m[1992])|(~m[1957]&~m[1988]&~m[1989]&~m[1991]&m[1992])|(m[1957]&~m[1988]&~m[1989]&~m[1991]&m[1992])|(m[1957]&m[1988]&~m[1989]&~m[1991]&m[1992])|(m[1957]&~m[1988]&m[1989]&~m[1991]&m[1992])|(~m[1957]&~m[1988]&~m[1989]&m[1991]&m[1992])|(m[1957]&~m[1988]&~m[1989]&m[1991]&m[1992])|(~m[1957]&m[1988]&~m[1989]&m[1991]&m[1992])|(m[1957]&m[1988]&~m[1989]&m[1991]&m[1992])|(~m[1957]&~m[1988]&m[1989]&m[1991]&m[1992])|(m[1957]&~m[1988]&m[1989]&m[1991]&m[1992])|(m[1957]&m[1988]&m[1989]&m[1991]&m[1992]))):InitCond[1107];
    m[1995] = run?((((m[1962]&~m[1993]&~m[1994]&~m[1996]&~m[1997])|(~m[1962]&~m[1993]&~m[1994]&m[1996]&~m[1997])|(m[1962]&m[1993]&~m[1994]&m[1996]&~m[1997])|(m[1962]&~m[1993]&m[1994]&m[1996]&~m[1997])|(~m[1962]&m[1993]&~m[1994]&~m[1996]&m[1997])|(~m[1962]&~m[1993]&m[1994]&~m[1996]&m[1997])|(m[1962]&m[1993]&m[1994]&~m[1996]&m[1997])|(~m[1962]&m[1993]&m[1994]&m[1996]&m[1997]))&UnbiasedRNG[469])|((m[1962]&~m[1993]&~m[1994]&m[1996]&~m[1997])|(~m[1962]&~m[1993]&~m[1994]&~m[1996]&m[1997])|(m[1962]&~m[1993]&~m[1994]&~m[1996]&m[1997])|(m[1962]&m[1993]&~m[1994]&~m[1996]&m[1997])|(m[1962]&~m[1993]&m[1994]&~m[1996]&m[1997])|(~m[1962]&~m[1993]&~m[1994]&m[1996]&m[1997])|(m[1962]&~m[1993]&~m[1994]&m[1996]&m[1997])|(~m[1962]&m[1993]&~m[1994]&m[1996]&m[1997])|(m[1962]&m[1993]&~m[1994]&m[1996]&m[1997])|(~m[1962]&~m[1993]&m[1994]&m[1996]&m[1997])|(m[1962]&~m[1993]&m[1994]&m[1996]&m[1997])|(m[1962]&m[1993]&m[1994]&m[1996]&m[1997]))):InitCond[1108];
    m[2000] = run?((((m[1967]&~m[1998]&~m[1999]&~m[2001]&~m[2002])|(~m[1967]&~m[1998]&~m[1999]&m[2001]&~m[2002])|(m[1967]&m[1998]&~m[1999]&m[2001]&~m[2002])|(m[1967]&~m[1998]&m[1999]&m[2001]&~m[2002])|(~m[1967]&m[1998]&~m[1999]&~m[2001]&m[2002])|(~m[1967]&~m[1998]&m[1999]&~m[2001]&m[2002])|(m[1967]&m[1998]&m[1999]&~m[2001]&m[2002])|(~m[1967]&m[1998]&m[1999]&m[2001]&m[2002]))&UnbiasedRNG[470])|((m[1967]&~m[1998]&~m[1999]&m[2001]&~m[2002])|(~m[1967]&~m[1998]&~m[1999]&~m[2001]&m[2002])|(m[1967]&~m[1998]&~m[1999]&~m[2001]&m[2002])|(m[1967]&m[1998]&~m[1999]&~m[2001]&m[2002])|(m[1967]&~m[1998]&m[1999]&~m[2001]&m[2002])|(~m[1967]&~m[1998]&~m[1999]&m[2001]&m[2002])|(m[1967]&~m[1998]&~m[1999]&m[2001]&m[2002])|(~m[1967]&m[1998]&~m[1999]&m[2001]&m[2002])|(m[1967]&m[1998]&~m[1999]&m[2001]&m[2002])|(~m[1967]&~m[1998]&m[1999]&m[2001]&m[2002])|(m[1967]&~m[1998]&m[1999]&m[2001]&m[2002])|(m[1967]&m[1998]&m[1999]&m[2001]&m[2002]))):InitCond[1109];
    m[2005] = run?((((m[1972]&~m[2003]&~m[2004]&~m[2006]&~m[2007])|(~m[1972]&~m[2003]&~m[2004]&m[2006]&~m[2007])|(m[1972]&m[2003]&~m[2004]&m[2006]&~m[2007])|(m[1972]&~m[2003]&m[2004]&m[2006]&~m[2007])|(~m[1972]&m[2003]&~m[2004]&~m[2006]&m[2007])|(~m[1972]&~m[2003]&m[2004]&~m[2006]&m[2007])|(m[1972]&m[2003]&m[2004]&~m[2006]&m[2007])|(~m[1972]&m[2003]&m[2004]&m[2006]&m[2007]))&UnbiasedRNG[471])|((m[1972]&~m[2003]&~m[2004]&m[2006]&~m[2007])|(~m[1972]&~m[2003]&~m[2004]&~m[2006]&m[2007])|(m[1972]&~m[2003]&~m[2004]&~m[2006]&m[2007])|(m[1972]&m[2003]&~m[2004]&~m[2006]&m[2007])|(m[1972]&~m[2003]&m[2004]&~m[2006]&m[2007])|(~m[1972]&~m[2003]&~m[2004]&m[2006]&m[2007])|(m[1972]&~m[2003]&~m[2004]&m[2006]&m[2007])|(~m[1972]&m[2003]&~m[2004]&m[2006]&m[2007])|(m[1972]&m[2003]&~m[2004]&m[2006]&m[2007])|(~m[1972]&~m[2003]&m[2004]&m[2006]&m[2007])|(m[1972]&~m[2003]&m[2004]&m[2006]&m[2007])|(m[1972]&m[2003]&m[2004]&m[2006]&m[2007]))):InitCond[1110];
    m[2010] = run?((((m[1977]&~m[2008]&~m[2009]&~m[2011]&~m[2012])|(~m[1977]&~m[2008]&~m[2009]&m[2011]&~m[2012])|(m[1977]&m[2008]&~m[2009]&m[2011]&~m[2012])|(m[1977]&~m[2008]&m[2009]&m[2011]&~m[2012])|(~m[1977]&m[2008]&~m[2009]&~m[2011]&m[2012])|(~m[1977]&~m[2008]&m[2009]&~m[2011]&m[2012])|(m[1977]&m[2008]&m[2009]&~m[2011]&m[2012])|(~m[1977]&m[2008]&m[2009]&m[2011]&m[2012]))&UnbiasedRNG[472])|((m[1977]&~m[2008]&~m[2009]&m[2011]&~m[2012])|(~m[1977]&~m[2008]&~m[2009]&~m[2011]&m[2012])|(m[1977]&~m[2008]&~m[2009]&~m[2011]&m[2012])|(m[1977]&m[2008]&~m[2009]&~m[2011]&m[2012])|(m[1977]&~m[2008]&m[2009]&~m[2011]&m[2012])|(~m[1977]&~m[2008]&~m[2009]&m[2011]&m[2012])|(m[1977]&~m[2008]&~m[2009]&m[2011]&m[2012])|(~m[1977]&m[2008]&~m[2009]&m[2011]&m[2012])|(m[1977]&m[2008]&~m[2009]&m[2011]&m[2012])|(~m[1977]&~m[2008]&m[2009]&m[2011]&m[2012])|(m[1977]&~m[2008]&m[2009]&m[2011]&m[2012])|(m[1977]&m[2008]&m[2009]&m[2011]&m[2012]))):InitCond[1111];
    m[2015] = run?((((m[1982]&~m[2013]&~m[2014]&~m[2016]&~m[2017])|(~m[1982]&~m[2013]&~m[2014]&m[2016]&~m[2017])|(m[1982]&m[2013]&~m[2014]&m[2016]&~m[2017])|(m[1982]&~m[2013]&m[2014]&m[2016]&~m[2017])|(~m[1982]&m[2013]&~m[2014]&~m[2016]&m[2017])|(~m[1982]&~m[2013]&m[2014]&~m[2016]&m[2017])|(m[1982]&m[2013]&m[2014]&~m[2016]&m[2017])|(~m[1982]&m[2013]&m[2014]&m[2016]&m[2017]))&UnbiasedRNG[473])|((m[1982]&~m[2013]&~m[2014]&m[2016]&~m[2017])|(~m[1982]&~m[2013]&~m[2014]&~m[2016]&m[2017])|(m[1982]&~m[2013]&~m[2014]&~m[2016]&m[2017])|(m[1982]&m[2013]&~m[2014]&~m[2016]&m[2017])|(m[1982]&~m[2013]&m[2014]&~m[2016]&m[2017])|(~m[1982]&~m[2013]&~m[2014]&m[2016]&m[2017])|(m[1982]&~m[2013]&~m[2014]&m[2016]&m[2017])|(~m[1982]&m[2013]&~m[2014]&m[2016]&m[2017])|(m[1982]&m[2013]&~m[2014]&m[2016]&m[2017])|(~m[1982]&~m[2013]&m[2014]&m[2016]&m[2017])|(m[1982]&~m[2013]&m[2014]&m[2016]&m[2017])|(m[1982]&m[2013]&m[2014]&m[2016]&m[2017]))):InitCond[1112];
    m[2020] = run?((((m[1987]&~m[2018]&~m[2019]&~m[2021]&~m[2022])|(~m[1987]&~m[2018]&~m[2019]&m[2021]&~m[2022])|(m[1987]&m[2018]&~m[2019]&m[2021]&~m[2022])|(m[1987]&~m[2018]&m[2019]&m[2021]&~m[2022])|(~m[1987]&m[2018]&~m[2019]&~m[2021]&m[2022])|(~m[1987]&~m[2018]&m[2019]&~m[2021]&m[2022])|(m[1987]&m[2018]&m[2019]&~m[2021]&m[2022])|(~m[1987]&m[2018]&m[2019]&m[2021]&m[2022]))&UnbiasedRNG[474])|((m[1987]&~m[2018]&~m[2019]&m[2021]&~m[2022])|(~m[1987]&~m[2018]&~m[2019]&~m[2021]&m[2022])|(m[1987]&~m[2018]&~m[2019]&~m[2021]&m[2022])|(m[1987]&m[2018]&~m[2019]&~m[2021]&m[2022])|(m[1987]&~m[2018]&m[2019]&~m[2021]&m[2022])|(~m[1987]&~m[2018]&~m[2019]&m[2021]&m[2022])|(m[1987]&~m[2018]&~m[2019]&m[2021]&m[2022])|(~m[1987]&m[2018]&~m[2019]&m[2021]&m[2022])|(m[1987]&m[2018]&~m[2019]&m[2021]&m[2022])|(~m[1987]&~m[2018]&m[2019]&m[2021]&m[2022])|(m[1987]&~m[2018]&m[2019]&m[2021]&m[2022])|(m[1987]&m[2018]&m[2019]&m[2021]&m[2022]))):InitCond[1113];
    m[2025] = run?((((m[1997]&~m[2023]&~m[2024]&~m[2026]&~m[2027])|(~m[1997]&~m[2023]&~m[2024]&m[2026]&~m[2027])|(m[1997]&m[2023]&~m[2024]&m[2026]&~m[2027])|(m[1997]&~m[2023]&m[2024]&m[2026]&~m[2027])|(~m[1997]&m[2023]&~m[2024]&~m[2026]&m[2027])|(~m[1997]&~m[2023]&m[2024]&~m[2026]&m[2027])|(m[1997]&m[2023]&m[2024]&~m[2026]&m[2027])|(~m[1997]&m[2023]&m[2024]&m[2026]&m[2027]))&UnbiasedRNG[475])|((m[1997]&~m[2023]&~m[2024]&m[2026]&~m[2027])|(~m[1997]&~m[2023]&~m[2024]&~m[2026]&m[2027])|(m[1997]&~m[2023]&~m[2024]&~m[2026]&m[2027])|(m[1997]&m[2023]&~m[2024]&~m[2026]&m[2027])|(m[1997]&~m[2023]&m[2024]&~m[2026]&m[2027])|(~m[1997]&~m[2023]&~m[2024]&m[2026]&m[2027])|(m[1997]&~m[2023]&~m[2024]&m[2026]&m[2027])|(~m[1997]&m[2023]&~m[2024]&m[2026]&m[2027])|(m[1997]&m[2023]&~m[2024]&m[2026]&m[2027])|(~m[1997]&~m[2023]&m[2024]&m[2026]&m[2027])|(m[1997]&~m[2023]&m[2024]&m[2026]&m[2027])|(m[1997]&m[2023]&m[2024]&m[2026]&m[2027]))):InitCond[1114];
    m[2030] = run?((((m[2002]&~m[2028]&~m[2029]&~m[2031]&~m[2032])|(~m[2002]&~m[2028]&~m[2029]&m[2031]&~m[2032])|(m[2002]&m[2028]&~m[2029]&m[2031]&~m[2032])|(m[2002]&~m[2028]&m[2029]&m[2031]&~m[2032])|(~m[2002]&m[2028]&~m[2029]&~m[2031]&m[2032])|(~m[2002]&~m[2028]&m[2029]&~m[2031]&m[2032])|(m[2002]&m[2028]&m[2029]&~m[2031]&m[2032])|(~m[2002]&m[2028]&m[2029]&m[2031]&m[2032]))&UnbiasedRNG[476])|((m[2002]&~m[2028]&~m[2029]&m[2031]&~m[2032])|(~m[2002]&~m[2028]&~m[2029]&~m[2031]&m[2032])|(m[2002]&~m[2028]&~m[2029]&~m[2031]&m[2032])|(m[2002]&m[2028]&~m[2029]&~m[2031]&m[2032])|(m[2002]&~m[2028]&m[2029]&~m[2031]&m[2032])|(~m[2002]&~m[2028]&~m[2029]&m[2031]&m[2032])|(m[2002]&~m[2028]&~m[2029]&m[2031]&m[2032])|(~m[2002]&m[2028]&~m[2029]&m[2031]&m[2032])|(m[2002]&m[2028]&~m[2029]&m[2031]&m[2032])|(~m[2002]&~m[2028]&m[2029]&m[2031]&m[2032])|(m[2002]&~m[2028]&m[2029]&m[2031]&m[2032])|(m[2002]&m[2028]&m[2029]&m[2031]&m[2032]))):InitCond[1115];
    m[2035] = run?((((m[2007]&~m[2033]&~m[2034]&~m[2036]&~m[2037])|(~m[2007]&~m[2033]&~m[2034]&m[2036]&~m[2037])|(m[2007]&m[2033]&~m[2034]&m[2036]&~m[2037])|(m[2007]&~m[2033]&m[2034]&m[2036]&~m[2037])|(~m[2007]&m[2033]&~m[2034]&~m[2036]&m[2037])|(~m[2007]&~m[2033]&m[2034]&~m[2036]&m[2037])|(m[2007]&m[2033]&m[2034]&~m[2036]&m[2037])|(~m[2007]&m[2033]&m[2034]&m[2036]&m[2037]))&UnbiasedRNG[477])|((m[2007]&~m[2033]&~m[2034]&m[2036]&~m[2037])|(~m[2007]&~m[2033]&~m[2034]&~m[2036]&m[2037])|(m[2007]&~m[2033]&~m[2034]&~m[2036]&m[2037])|(m[2007]&m[2033]&~m[2034]&~m[2036]&m[2037])|(m[2007]&~m[2033]&m[2034]&~m[2036]&m[2037])|(~m[2007]&~m[2033]&~m[2034]&m[2036]&m[2037])|(m[2007]&~m[2033]&~m[2034]&m[2036]&m[2037])|(~m[2007]&m[2033]&~m[2034]&m[2036]&m[2037])|(m[2007]&m[2033]&~m[2034]&m[2036]&m[2037])|(~m[2007]&~m[2033]&m[2034]&m[2036]&m[2037])|(m[2007]&~m[2033]&m[2034]&m[2036]&m[2037])|(m[2007]&m[2033]&m[2034]&m[2036]&m[2037]))):InitCond[1116];
    m[2040] = run?((((m[2012]&~m[2038]&~m[2039]&~m[2041]&~m[2042])|(~m[2012]&~m[2038]&~m[2039]&m[2041]&~m[2042])|(m[2012]&m[2038]&~m[2039]&m[2041]&~m[2042])|(m[2012]&~m[2038]&m[2039]&m[2041]&~m[2042])|(~m[2012]&m[2038]&~m[2039]&~m[2041]&m[2042])|(~m[2012]&~m[2038]&m[2039]&~m[2041]&m[2042])|(m[2012]&m[2038]&m[2039]&~m[2041]&m[2042])|(~m[2012]&m[2038]&m[2039]&m[2041]&m[2042]))&UnbiasedRNG[478])|((m[2012]&~m[2038]&~m[2039]&m[2041]&~m[2042])|(~m[2012]&~m[2038]&~m[2039]&~m[2041]&m[2042])|(m[2012]&~m[2038]&~m[2039]&~m[2041]&m[2042])|(m[2012]&m[2038]&~m[2039]&~m[2041]&m[2042])|(m[2012]&~m[2038]&m[2039]&~m[2041]&m[2042])|(~m[2012]&~m[2038]&~m[2039]&m[2041]&m[2042])|(m[2012]&~m[2038]&~m[2039]&m[2041]&m[2042])|(~m[2012]&m[2038]&~m[2039]&m[2041]&m[2042])|(m[2012]&m[2038]&~m[2039]&m[2041]&m[2042])|(~m[2012]&~m[2038]&m[2039]&m[2041]&m[2042])|(m[2012]&~m[2038]&m[2039]&m[2041]&m[2042])|(m[2012]&m[2038]&m[2039]&m[2041]&m[2042]))):InitCond[1117];
    m[2045] = run?((((m[2017]&~m[2043]&~m[2044]&~m[2046]&~m[2047])|(~m[2017]&~m[2043]&~m[2044]&m[2046]&~m[2047])|(m[2017]&m[2043]&~m[2044]&m[2046]&~m[2047])|(m[2017]&~m[2043]&m[2044]&m[2046]&~m[2047])|(~m[2017]&m[2043]&~m[2044]&~m[2046]&m[2047])|(~m[2017]&~m[2043]&m[2044]&~m[2046]&m[2047])|(m[2017]&m[2043]&m[2044]&~m[2046]&m[2047])|(~m[2017]&m[2043]&m[2044]&m[2046]&m[2047]))&UnbiasedRNG[479])|((m[2017]&~m[2043]&~m[2044]&m[2046]&~m[2047])|(~m[2017]&~m[2043]&~m[2044]&~m[2046]&m[2047])|(m[2017]&~m[2043]&~m[2044]&~m[2046]&m[2047])|(m[2017]&m[2043]&~m[2044]&~m[2046]&m[2047])|(m[2017]&~m[2043]&m[2044]&~m[2046]&m[2047])|(~m[2017]&~m[2043]&~m[2044]&m[2046]&m[2047])|(m[2017]&~m[2043]&~m[2044]&m[2046]&m[2047])|(~m[2017]&m[2043]&~m[2044]&m[2046]&m[2047])|(m[2017]&m[2043]&~m[2044]&m[2046]&m[2047])|(~m[2017]&~m[2043]&m[2044]&m[2046]&m[2047])|(m[2017]&~m[2043]&m[2044]&m[2046]&m[2047])|(m[2017]&m[2043]&m[2044]&m[2046]&m[2047]))):InitCond[1118];
    m[2050] = run?((((m[2022]&~m[2048]&~m[2049]&~m[2051]&~m[2052])|(~m[2022]&~m[2048]&~m[2049]&m[2051]&~m[2052])|(m[2022]&m[2048]&~m[2049]&m[2051]&~m[2052])|(m[2022]&~m[2048]&m[2049]&m[2051]&~m[2052])|(~m[2022]&m[2048]&~m[2049]&~m[2051]&m[2052])|(~m[2022]&~m[2048]&m[2049]&~m[2051]&m[2052])|(m[2022]&m[2048]&m[2049]&~m[2051]&m[2052])|(~m[2022]&m[2048]&m[2049]&m[2051]&m[2052]))&UnbiasedRNG[480])|((m[2022]&~m[2048]&~m[2049]&m[2051]&~m[2052])|(~m[2022]&~m[2048]&~m[2049]&~m[2051]&m[2052])|(m[2022]&~m[2048]&~m[2049]&~m[2051]&m[2052])|(m[2022]&m[2048]&~m[2049]&~m[2051]&m[2052])|(m[2022]&~m[2048]&m[2049]&~m[2051]&m[2052])|(~m[2022]&~m[2048]&~m[2049]&m[2051]&m[2052])|(m[2022]&~m[2048]&~m[2049]&m[2051]&m[2052])|(~m[2022]&m[2048]&~m[2049]&m[2051]&m[2052])|(m[2022]&m[2048]&~m[2049]&m[2051]&m[2052])|(~m[2022]&~m[2048]&m[2049]&m[2051]&m[2052])|(m[2022]&~m[2048]&m[2049]&m[2051]&m[2052])|(m[2022]&m[2048]&m[2049]&m[2051]&m[2052]))):InitCond[1119];
    m[2055] = run?((((m[2032]&~m[2053]&~m[2054]&~m[2056]&~m[2057])|(~m[2032]&~m[2053]&~m[2054]&m[2056]&~m[2057])|(m[2032]&m[2053]&~m[2054]&m[2056]&~m[2057])|(m[2032]&~m[2053]&m[2054]&m[2056]&~m[2057])|(~m[2032]&m[2053]&~m[2054]&~m[2056]&m[2057])|(~m[2032]&~m[2053]&m[2054]&~m[2056]&m[2057])|(m[2032]&m[2053]&m[2054]&~m[2056]&m[2057])|(~m[2032]&m[2053]&m[2054]&m[2056]&m[2057]))&UnbiasedRNG[481])|((m[2032]&~m[2053]&~m[2054]&m[2056]&~m[2057])|(~m[2032]&~m[2053]&~m[2054]&~m[2056]&m[2057])|(m[2032]&~m[2053]&~m[2054]&~m[2056]&m[2057])|(m[2032]&m[2053]&~m[2054]&~m[2056]&m[2057])|(m[2032]&~m[2053]&m[2054]&~m[2056]&m[2057])|(~m[2032]&~m[2053]&~m[2054]&m[2056]&m[2057])|(m[2032]&~m[2053]&~m[2054]&m[2056]&m[2057])|(~m[2032]&m[2053]&~m[2054]&m[2056]&m[2057])|(m[2032]&m[2053]&~m[2054]&m[2056]&m[2057])|(~m[2032]&~m[2053]&m[2054]&m[2056]&m[2057])|(m[2032]&~m[2053]&m[2054]&m[2056]&m[2057])|(m[2032]&m[2053]&m[2054]&m[2056]&m[2057]))):InitCond[1120];
    m[2060] = run?((((m[2037]&~m[2058]&~m[2059]&~m[2061]&~m[2062])|(~m[2037]&~m[2058]&~m[2059]&m[2061]&~m[2062])|(m[2037]&m[2058]&~m[2059]&m[2061]&~m[2062])|(m[2037]&~m[2058]&m[2059]&m[2061]&~m[2062])|(~m[2037]&m[2058]&~m[2059]&~m[2061]&m[2062])|(~m[2037]&~m[2058]&m[2059]&~m[2061]&m[2062])|(m[2037]&m[2058]&m[2059]&~m[2061]&m[2062])|(~m[2037]&m[2058]&m[2059]&m[2061]&m[2062]))&UnbiasedRNG[482])|((m[2037]&~m[2058]&~m[2059]&m[2061]&~m[2062])|(~m[2037]&~m[2058]&~m[2059]&~m[2061]&m[2062])|(m[2037]&~m[2058]&~m[2059]&~m[2061]&m[2062])|(m[2037]&m[2058]&~m[2059]&~m[2061]&m[2062])|(m[2037]&~m[2058]&m[2059]&~m[2061]&m[2062])|(~m[2037]&~m[2058]&~m[2059]&m[2061]&m[2062])|(m[2037]&~m[2058]&~m[2059]&m[2061]&m[2062])|(~m[2037]&m[2058]&~m[2059]&m[2061]&m[2062])|(m[2037]&m[2058]&~m[2059]&m[2061]&m[2062])|(~m[2037]&~m[2058]&m[2059]&m[2061]&m[2062])|(m[2037]&~m[2058]&m[2059]&m[2061]&m[2062])|(m[2037]&m[2058]&m[2059]&m[2061]&m[2062]))):InitCond[1121];
    m[2065] = run?((((m[2042]&~m[2063]&~m[2064]&~m[2066]&~m[2067])|(~m[2042]&~m[2063]&~m[2064]&m[2066]&~m[2067])|(m[2042]&m[2063]&~m[2064]&m[2066]&~m[2067])|(m[2042]&~m[2063]&m[2064]&m[2066]&~m[2067])|(~m[2042]&m[2063]&~m[2064]&~m[2066]&m[2067])|(~m[2042]&~m[2063]&m[2064]&~m[2066]&m[2067])|(m[2042]&m[2063]&m[2064]&~m[2066]&m[2067])|(~m[2042]&m[2063]&m[2064]&m[2066]&m[2067]))&UnbiasedRNG[483])|((m[2042]&~m[2063]&~m[2064]&m[2066]&~m[2067])|(~m[2042]&~m[2063]&~m[2064]&~m[2066]&m[2067])|(m[2042]&~m[2063]&~m[2064]&~m[2066]&m[2067])|(m[2042]&m[2063]&~m[2064]&~m[2066]&m[2067])|(m[2042]&~m[2063]&m[2064]&~m[2066]&m[2067])|(~m[2042]&~m[2063]&~m[2064]&m[2066]&m[2067])|(m[2042]&~m[2063]&~m[2064]&m[2066]&m[2067])|(~m[2042]&m[2063]&~m[2064]&m[2066]&m[2067])|(m[2042]&m[2063]&~m[2064]&m[2066]&m[2067])|(~m[2042]&~m[2063]&m[2064]&m[2066]&m[2067])|(m[2042]&~m[2063]&m[2064]&m[2066]&m[2067])|(m[2042]&m[2063]&m[2064]&m[2066]&m[2067]))):InitCond[1122];
    m[2070] = run?((((m[2047]&~m[2068]&~m[2069]&~m[2071]&~m[2072])|(~m[2047]&~m[2068]&~m[2069]&m[2071]&~m[2072])|(m[2047]&m[2068]&~m[2069]&m[2071]&~m[2072])|(m[2047]&~m[2068]&m[2069]&m[2071]&~m[2072])|(~m[2047]&m[2068]&~m[2069]&~m[2071]&m[2072])|(~m[2047]&~m[2068]&m[2069]&~m[2071]&m[2072])|(m[2047]&m[2068]&m[2069]&~m[2071]&m[2072])|(~m[2047]&m[2068]&m[2069]&m[2071]&m[2072]))&UnbiasedRNG[484])|((m[2047]&~m[2068]&~m[2069]&m[2071]&~m[2072])|(~m[2047]&~m[2068]&~m[2069]&~m[2071]&m[2072])|(m[2047]&~m[2068]&~m[2069]&~m[2071]&m[2072])|(m[2047]&m[2068]&~m[2069]&~m[2071]&m[2072])|(m[2047]&~m[2068]&m[2069]&~m[2071]&m[2072])|(~m[2047]&~m[2068]&~m[2069]&m[2071]&m[2072])|(m[2047]&~m[2068]&~m[2069]&m[2071]&m[2072])|(~m[2047]&m[2068]&~m[2069]&m[2071]&m[2072])|(m[2047]&m[2068]&~m[2069]&m[2071]&m[2072])|(~m[2047]&~m[2068]&m[2069]&m[2071]&m[2072])|(m[2047]&~m[2068]&m[2069]&m[2071]&m[2072])|(m[2047]&m[2068]&m[2069]&m[2071]&m[2072]))):InitCond[1123];
    m[2075] = run?((((m[2052]&~m[2073]&~m[2074]&~m[2076]&~m[2077])|(~m[2052]&~m[2073]&~m[2074]&m[2076]&~m[2077])|(m[2052]&m[2073]&~m[2074]&m[2076]&~m[2077])|(m[2052]&~m[2073]&m[2074]&m[2076]&~m[2077])|(~m[2052]&m[2073]&~m[2074]&~m[2076]&m[2077])|(~m[2052]&~m[2073]&m[2074]&~m[2076]&m[2077])|(m[2052]&m[2073]&m[2074]&~m[2076]&m[2077])|(~m[2052]&m[2073]&m[2074]&m[2076]&m[2077]))&UnbiasedRNG[485])|((m[2052]&~m[2073]&~m[2074]&m[2076]&~m[2077])|(~m[2052]&~m[2073]&~m[2074]&~m[2076]&m[2077])|(m[2052]&~m[2073]&~m[2074]&~m[2076]&m[2077])|(m[2052]&m[2073]&~m[2074]&~m[2076]&m[2077])|(m[2052]&~m[2073]&m[2074]&~m[2076]&m[2077])|(~m[2052]&~m[2073]&~m[2074]&m[2076]&m[2077])|(m[2052]&~m[2073]&~m[2074]&m[2076]&m[2077])|(~m[2052]&m[2073]&~m[2074]&m[2076]&m[2077])|(m[2052]&m[2073]&~m[2074]&m[2076]&m[2077])|(~m[2052]&~m[2073]&m[2074]&m[2076]&m[2077])|(m[2052]&~m[2073]&m[2074]&m[2076]&m[2077])|(m[2052]&m[2073]&m[2074]&m[2076]&m[2077]))):InitCond[1124];
    m[2080] = run?((((m[2062]&~m[2078]&~m[2079]&~m[2081]&~m[2082])|(~m[2062]&~m[2078]&~m[2079]&m[2081]&~m[2082])|(m[2062]&m[2078]&~m[2079]&m[2081]&~m[2082])|(m[2062]&~m[2078]&m[2079]&m[2081]&~m[2082])|(~m[2062]&m[2078]&~m[2079]&~m[2081]&m[2082])|(~m[2062]&~m[2078]&m[2079]&~m[2081]&m[2082])|(m[2062]&m[2078]&m[2079]&~m[2081]&m[2082])|(~m[2062]&m[2078]&m[2079]&m[2081]&m[2082]))&UnbiasedRNG[486])|((m[2062]&~m[2078]&~m[2079]&m[2081]&~m[2082])|(~m[2062]&~m[2078]&~m[2079]&~m[2081]&m[2082])|(m[2062]&~m[2078]&~m[2079]&~m[2081]&m[2082])|(m[2062]&m[2078]&~m[2079]&~m[2081]&m[2082])|(m[2062]&~m[2078]&m[2079]&~m[2081]&m[2082])|(~m[2062]&~m[2078]&~m[2079]&m[2081]&m[2082])|(m[2062]&~m[2078]&~m[2079]&m[2081]&m[2082])|(~m[2062]&m[2078]&~m[2079]&m[2081]&m[2082])|(m[2062]&m[2078]&~m[2079]&m[2081]&m[2082])|(~m[2062]&~m[2078]&m[2079]&m[2081]&m[2082])|(m[2062]&~m[2078]&m[2079]&m[2081]&m[2082])|(m[2062]&m[2078]&m[2079]&m[2081]&m[2082]))):InitCond[1125];
    m[2085] = run?((((m[2067]&~m[2083]&~m[2084]&~m[2086]&~m[2087])|(~m[2067]&~m[2083]&~m[2084]&m[2086]&~m[2087])|(m[2067]&m[2083]&~m[2084]&m[2086]&~m[2087])|(m[2067]&~m[2083]&m[2084]&m[2086]&~m[2087])|(~m[2067]&m[2083]&~m[2084]&~m[2086]&m[2087])|(~m[2067]&~m[2083]&m[2084]&~m[2086]&m[2087])|(m[2067]&m[2083]&m[2084]&~m[2086]&m[2087])|(~m[2067]&m[2083]&m[2084]&m[2086]&m[2087]))&UnbiasedRNG[487])|((m[2067]&~m[2083]&~m[2084]&m[2086]&~m[2087])|(~m[2067]&~m[2083]&~m[2084]&~m[2086]&m[2087])|(m[2067]&~m[2083]&~m[2084]&~m[2086]&m[2087])|(m[2067]&m[2083]&~m[2084]&~m[2086]&m[2087])|(m[2067]&~m[2083]&m[2084]&~m[2086]&m[2087])|(~m[2067]&~m[2083]&~m[2084]&m[2086]&m[2087])|(m[2067]&~m[2083]&~m[2084]&m[2086]&m[2087])|(~m[2067]&m[2083]&~m[2084]&m[2086]&m[2087])|(m[2067]&m[2083]&~m[2084]&m[2086]&m[2087])|(~m[2067]&~m[2083]&m[2084]&m[2086]&m[2087])|(m[2067]&~m[2083]&m[2084]&m[2086]&m[2087])|(m[2067]&m[2083]&m[2084]&m[2086]&m[2087]))):InitCond[1126];
    m[2090] = run?((((m[2072]&~m[2088]&~m[2089]&~m[2091]&~m[2092])|(~m[2072]&~m[2088]&~m[2089]&m[2091]&~m[2092])|(m[2072]&m[2088]&~m[2089]&m[2091]&~m[2092])|(m[2072]&~m[2088]&m[2089]&m[2091]&~m[2092])|(~m[2072]&m[2088]&~m[2089]&~m[2091]&m[2092])|(~m[2072]&~m[2088]&m[2089]&~m[2091]&m[2092])|(m[2072]&m[2088]&m[2089]&~m[2091]&m[2092])|(~m[2072]&m[2088]&m[2089]&m[2091]&m[2092]))&UnbiasedRNG[488])|((m[2072]&~m[2088]&~m[2089]&m[2091]&~m[2092])|(~m[2072]&~m[2088]&~m[2089]&~m[2091]&m[2092])|(m[2072]&~m[2088]&~m[2089]&~m[2091]&m[2092])|(m[2072]&m[2088]&~m[2089]&~m[2091]&m[2092])|(m[2072]&~m[2088]&m[2089]&~m[2091]&m[2092])|(~m[2072]&~m[2088]&~m[2089]&m[2091]&m[2092])|(m[2072]&~m[2088]&~m[2089]&m[2091]&m[2092])|(~m[2072]&m[2088]&~m[2089]&m[2091]&m[2092])|(m[2072]&m[2088]&~m[2089]&m[2091]&m[2092])|(~m[2072]&~m[2088]&m[2089]&m[2091]&m[2092])|(m[2072]&~m[2088]&m[2089]&m[2091]&m[2092])|(m[2072]&m[2088]&m[2089]&m[2091]&m[2092]))):InitCond[1127];
    m[2095] = run?((((m[2077]&~m[2093]&~m[2094]&~m[2096]&~m[2097])|(~m[2077]&~m[2093]&~m[2094]&m[2096]&~m[2097])|(m[2077]&m[2093]&~m[2094]&m[2096]&~m[2097])|(m[2077]&~m[2093]&m[2094]&m[2096]&~m[2097])|(~m[2077]&m[2093]&~m[2094]&~m[2096]&m[2097])|(~m[2077]&~m[2093]&m[2094]&~m[2096]&m[2097])|(m[2077]&m[2093]&m[2094]&~m[2096]&m[2097])|(~m[2077]&m[2093]&m[2094]&m[2096]&m[2097]))&UnbiasedRNG[489])|((m[2077]&~m[2093]&~m[2094]&m[2096]&~m[2097])|(~m[2077]&~m[2093]&~m[2094]&~m[2096]&m[2097])|(m[2077]&~m[2093]&~m[2094]&~m[2096]&m[2097])|(m[2077]&m[2093]&~m[2094]&~m[2096]&m[2097])|(m[2077]&~m[2093]&m[2094]&~m[2096]&m[2097])|(~m[2077]&~m[2093]&~m[2094]&m[2096]&m[2097])|(m[2077]&~m[2093]&~m[2094]&m[2096]&m[2097])|(~m[2077]&m[2093]&~m[2094]&m[2096]&m[2097])|(m[2077]&m[2093]&~m[2094]&m[2096]&m[2097])|(~m[2077]&~m[2093]&m[2094]&m[2096]&m[2097])|(m[2077]&~m[2093]&m[2094]&m[2096]&m[2097])|(m[2077]&m[2093]&m[2094]&m[2096]&m[2097]))):InitCond[1128];
    m[2100] = run?((((m[2087]&~m[2098]&~m[2099]&~m[2101]&~m[2102])|(~m[2087]&~m[2098]&~m[2099]&m[2101]&~m[2102])|(m[2087]&m[2098]&~m[2099]&m[2101]&~m[2102])|(m[2087]&~m[2098]&m[2099]&m[2101]&~m[2102])|(~m[2087]&m[2098]&~m[2099]&~m[2101]&m[2102])|(~m[2087]&~m[2098]&m[2099]&~m[2101]&m[2102])|(m[2087]&m[2098]&m[2099]&~m[2101]&m[2102])|(~m[2087]&m[2098]&m[2099]&m[2101]&m[2102]))&UnbiasedRNG[490])|((m[2087]&~m[2098]&~m[2099]&m[2101]&~m[2102])|(~m[2087]&~m[2098]&~m[2099]&~m[2101]&m[2102])|(m[2087]&~m[2098]&~m[2099]&~m[2101]&m[2102])|(m[2087]&m[2098]&~m[2099]&~m[2101]&m[2102])|(m[2087]&~m[2098]&m[2099]&~m[2101]&m[2102])|(~m[2087]&~m[2098]&~m[2099]&m[2101]&m[2102])|(m[2087]&~m[2098]&~m[2099]&m[2101]&m[2102])|(~m[2087]&m[2098]&~m[2099]&m[2101]&m[2102])|(m[2087]&m[2098]&~m[2099]&m[2101]&m[2102])|(~m[2087]&~m[2098]&m[2099]&m[2101]&m[2102])|(m[2087]&~m[2098]&m[2099]&m[2101]&m[2102])|(m[2087]&m[2098]&m[2099]&m[2101]&m[2102]))):InitCond[1129];
    m[2105] = run?((((m[2092]&~m[2103]&~m[2104]&~m[2106]&~m[2107])|(~m[2092]&~m[2103]&~m[2104]&m[2106]&~m[2107])|(m[2092]&m[2103]&~m[2104]&m[2106]&~m[2107])|(m[2092]&~m[2103]&m[2104]&m[2106]&~m[2107])|(~m[2092]&m[2103]&~m[2104]&~m[2106]&m[2107])|(~m[2092]&~m[2103]&m[2104]&~m[2106]&m[2107])|(m[2092]&m[2103]&m[2104]&~m[2106]&m[2107])|(~m[2092]&m[2103]&m[2104]&m[2106]&m[2107]))&UnbiasedRNG[491])|((m[2092]&~m[2103]&~m[2104]&m[2106]&~m[2107])|(~m[2092]&~m[2103]&~m[2104]&~m[2106]&m[2107])|(m[2092]&~m[2103]&~m[2104]&~m[2106]&m[2107])|(m[2092]&m[2103]&~m[2104]&~m[2106]&m[2107])|(m[2092]&~m[2103]&m[2104]&~m[2106]&m[2107])|(~m[2092]&~m[2103]&~m[2104]&m[2106]&m[2107])|(m[2092]&~m[2103]&~m[2104]&m[2106]&m[2107])|(~m[2092]&m[2103]&~m[2104]&m[2106]&m[2107])|(m[2092]&m[2103]&~m[2104]&m[2106]&m[2107])|(~m[2092]&~m[2103]&m[2104]&m[2106]&m[2107])|(m[2092]&~m[2103]&m[2104]&m[2106]&m[2107])|(m[2092]&m[2103]&m[2104]&m[2106]&m[2107]))):InitCond[1130];
    m[2110] = run?((((m[2097]&~m[2108]&~m[2109]&~m[2111]&~m[2112])|(~m[2097]&~m[2108]&~m[2109]&m[2111]&~m[2112])|(m[2097]&m[2108]&~m[2109]&m[2111]&~m[2112])|(m[2097]&~m[2108]&m[2109]&m[2111]&~m[2112])|(~m[2097]&m[2108]&~m[2109]&~m[2111]&m[2112])|(~m[2097]&~m[2108]&m[2109]&~m[2111]&m[2112])|(m[2097]&m[2108]&m[2109]&~m[2111]&m[2112])|(~m[2097]&m[2108]&m[2109]&m[2111]&m[2112]))&UnbiasedRNG[492])|((m[2097]&~m[2108]&~m[2109]&m[2111]&~m[2112])|(~m[2097]&~m[2108]&~m[2109]&~m[2111]&m[2112])|(m[2097]&~m[2108]&~m[2109]&~m[2111]&m[2112])|(m[2097]&m[2108]&~m[2109]&~m[2111]&m[2112])|(m[2097]&~m[2108]&m[2109]&~m[2111]&m[2112])|(~m[2097]&~m[2108]&~m[2109]&m[2111]&m[2112])|(m[2097]&~m[2108]&~m[2109]&m[2111]&m[2112])|(~m[2097]&m[2108]&~m[2109]&m[2111]&m[2112])|(m[2097]&m[2108]&~m[2109]&m[2111]&m[2112])|(~m[2097]&~m[2108]&m[2109]&m[2111]&m[2112])|(m[2097]&~m[2108]&m[2109]&m[2111]&m[2112])|(m[2097]&m[2108]&m[2109]&m[2111]&m[2112]))):InitCond[1131];
    m[2115] = run?((((m[2107]&~m[2113]&~m[2114]&~m[2116]&~m[2117])|(~m[2107]&~m[2113]&~m[2114]&m[2116]&~m[2117])|(m[2107]&m[2113]&~m[2114]&m[2116]&~m[2117])|(m[2107]&~m[2113]&m[2114]&m[2116]&~m[2117])|(~m[2107]&m[2113]&~m[2114]&~m[2116]&m[2117])|(~m[2107]&~m[2113]&m[2114]&~m[2116]&m[2117])|(m[2107]&m[2113]&m[2114]&~m[2116]&m[2117])|(~m[2107]&m[2113]&m[2114]&m[2116]&m[2117]))&UnbiasedRNG[493])|((m[2107]&~m[2113]&~m[2114]&m[2116]&~m[2117])|(~m[2107]&~m[2113]&~m[2114]&~m[2116]&m[2117])|(m[2107]&~m[2113]&~m[2114]&~m[2116]&m[2117])|(m[2107]&m[2113]&~m[2114]&~m[2116]&m[2117])|(m[2107]&~m[2113]&m[2114]&~m[2116]&m[2117])|(~m[2107]&~m[2113]&~m[2114]&m[2116]&m[2117])|(m[2107]&~m[2113]&~m[2114]&m[2116]&m[2117])|(~m[2107]&m[2113]&~m[2114]&m[2116]&m[2117])|(m[2107]&m[2113]&~m[2114]&m[2116]&m[2117])|(~m[2107]&~m[2113]&m[2114]&m[2116]&m[2117])|(m[2107]&~m[2113]&m[2114]&m[2116]&m[2117])|(m[2107]&m[2113]&m[2114]&m[2116]&m[2117]))):InitCond[1132];
    m[2120] = run?((((m[2112]&~m[2118]&~m[2119]&~m[2121]&~m[2122])|(~m[2112]&~m[2118]&~m[2119]&m[2121]&~m[2122])|(m[2112]&m[2118]&~m[2119]&m[2121]&~m[2122])|(m[2112]&~m[2118]&m[2119]&m[2121]&~m[2122])|(~m[2112]&m[2118]&~m[2119]&~m[2121]&m[2122])|(~m[2112]&~m[2118]&m[2119]&~m[2121]&m[2122])|(m[2112]&m[2118]&m[2119]&~m[2121]&m[2122])|(~m[2112]&m[2118]&m[2119]&m[2121]&m[2122]))&UnbiasedRNG[494])|((m[2112]&~m[2118]&~m[2119]&m[2121]&~m[2122])|(~m[2112]&~m[2118]&~m[2119]&~m[2121]&m[2122])|(m[2112]&~m[2118]&~m[2119]&~m[2121]&m[2122])|(m[2112]&m[2118]&~m[2119]&~m[2121]&m[2122])|(m[2112]&~m[2118]&m[2119]&~m[2121]&m[2122])|(~m[2112]&~m[2118]&~m[2119]&m[2121]&m[2122])|(m[2112]&~m[2118]&~m[2119]&m[2121]&m[2122])|(~m[2112]&m[2118]&~m[2119]&m[2121]&m[2122])|(m[2112]&m[2118]&~m[2119]&m[2121]&m[2122])|(~m[2112]&~m[2118]&m[2119]&m[2121]&m[2122])|(m[2112]&~m[2118]&m[2119]&m[2121]&m[2122])|(m[2112]&m[2118]&m[2119]&m[2121]&m[2122]))):InitCond[1133];
    m[2125] = run?((((m[2122]&~m[2123]&~m[2124]&~m[2126]&~m[2127])|(~m[2122]&~m[2123]&~m[2124]&m[2126]&~m[2127])|(m[2122]&m[2123]&~m[2124]&m[2126]&~m[2127])|(m[2122]&~m[2123]&m[2124]&m[2126]&~m[2127])|(~m[2122]&m[2123]&~m[2124]&~m[2126]&m[2127])|(~m[2122]&~m[2123]&m[2124]&~m[2126]&m[2127])|(m[2122]&m[2123]&m[2124]&~m[2126]&m[2127])|(~m[2122]&m[2123]&m[2124]&m[2126]&m[2127]))&UnbiasedRNG[495])|((m[2122]&~m[2123]&~m[2124]&m[2126]&~m[2127])|(~m[2122]&~m[2123]&~m[2124]&~m[2126]&m[2127])|(m[2122]&~m[2123]&~m[2124]&~m[2126]&m[2127])|(m[2122]&m[2123]&~m[2124]&~m[2126]&m[2127])|(m[2122]&~m[2123]&m[2124]&~m[2126]&m[2127])|(~m[2122]&~m[2123]&~m[2124]&m[2126]&m[2127])|(m[2122]&~m[2123]&~m[2124]&m[2126]&m[2127])|(~m[2122]&m[2123]&~m[2124]&m[2126]&m[2127])|(m[2122]&m[2123]&~m[2124]&m[2126]&m[2127])|(~m[2122]&~m[2123]&m[2124]&m[2126]&m[2127])|(m[2122]&~m[2123]&m[2124]&m[2126]&m[2127])|(m[2122]&m[2123]&m[2124]&m[2126]&m[2127]))):InitCond[1134];
end

always @(posedge color2_clk) begin
    m[416] = run?((((~m[96]&~m[160]&~m[672])|(m[96]&m[160]&~m[672]))&BiasedRNG[639])|(((m[96]&~m[160]&~m[672])|(~m[96]&m[160]&m[672]))&~BiasedRNG[639])|((~m[96]&~m[160]&m[672])|(m[96]&~m[160]&m[672])|(m[96]&m[160]&m[672]))):InitCond[1135];
    m[417] = run?((((~m[96]&~m[176]&~m[673])|(m[96]&m[176]&~m[673]))&BiasedRNG[640])|(((m[96]&~m[176]&~m[673])|(~m[96]&m[176]&m[673]))&~BiasedRNG[640])|((~m[96]&~m[176]&m[673])|(m[96]&~m[176]&m[673])|(m[96]&m[176]&m[673]))):InitCond[1136];
    m[418] = run?((((~m[96]&~m[192]&~m[674])|(m[96]&m[192]&~m[674]))&BiasedRNG[641])|(((m[96]&~m[192]&~m[674])|(~m[96]&m[192]&m[674]))&~BiasedRNG[641])|((~m[96]&~m[192]&m[674])|(m[96]&~m[192]&m[674])|(m[96]&m[192]&m[674]))):InitCond[1137];
    m[419] = run?((((~m[96]&~m[208]&~m[675])|(m[96]&m[208]&~m[675]))&BiasedRNG[642])|(((m[96]&~m[208]&~m[675])|(~m[96]&m[208]&m[675]))&~BiasedRNG[642])|((~m[96]&~m[208]&m[675])|(m[96]&~m[208]&m[675])|(m[96]&m[208]&m[675]))):InitCond[1138];
    m[420] = run?((((~m[97]&~m[224]&~m[676])|(m[97]&m[224]&~m[676]))&BiasedRNG[643])|(((m[97]&~m[224]&~m[676])|(~m[97]&m[224]&m[676]))&~BiasedRNG[643])|((~m[97]&~m[224]&m[676])|(m[97]&~m[224]&m[676])|(m[97]&m[224]&m[676]))):InitCond[1139];
    m[421] = run?((((~m[97]&~m[240]&~m[677])|(m[97]&m[240]&~m[677]))&BiasedRNG[644])|(((m[97]&~m[240]&~m[677])|(~m[97]&m[240]&m[677]))&~BiasedRNG[644])|((~m[97]&~m[240]&m[677])|(m[97]&~m[240]&m[677])|(m[97]&m[240]&m[677]))):InitCond[1140];
    m[422] = run?((((~m[97]&~m[256]&~m[678])|(m[97]&m[256]&~m[678]))&BiasedRNG[645])|(((m[97]&~m[256]&~m[678])|(~m[97]&m[256]&m[678]))&~BiasedRNG[645])|((~m[97]&~m[256]&m[678])|(m[97]&~m[256]&m[678])|(m[97]&m[256]&m[678]))):InitCond[1141];
    m[423] = run?((((~m[97]&~m[272]&~m[679])|(m[97]&m[272]&~m[679]))&BiasedRNG[646])|(((m[97]&~m[272]&~m[679])|(~m[97]&m[272]&m[679]))&~BiasedRNG[646])|((~m[97]&~m[272]&m[679])|(m[97]&~m[272]&m[679])|(m[97]&m[272]&m[679]))):InitCond[1142];
    m[424] = run?((((~m[98]&~m[288]&~m[680])|(m[98]&m[288]&~m[680]))&BiasedRNG[647])|(((m[98]&~m[288]&~m[680])|(~m[98]&m[288]&m[680]))&~BiasedRNG[647])|((~m[98]&~m[288]&m[680])|(m[98]&~m[288]&m[680])|(m[98]&m[288]&m[680]))):InitCond[1143];
    m[425] = run?((((~m[98]&~m[304]&~m[681])|(m[98]&m[304]&~m[681]))&BiasedRNG[648])|(((m[98]&~m[304]&~m[681])|(~m[98]&m[304]&m[681]))&~BiasedRNG[648])|((~m[98]&~m[304]&m[681])|(m[98]&~m[304]&m[681])|(m[98]&m[304]&m[681]))):InitCond[1144];
    m[426] = run?((((~m[98]&~m[320]&~m[682])|(m[98]&m[320]&~m[682]))&BiasedRNG[649])|(((m[98]&~m[320]&~m[682])|(~m[98]&m[320]&m[682]))&~BiasedRNG[649])|((~m[98]&~m[320]&m[682])|(m[98]&~m[320]&m[682])|(m[98]&m[320]&m[682]))):InitCond[1145];
    m[427] = run?((((~m[98]&~m[336]&~m[683])|(m[98]&m[336]&~m[683]))&BiasedRNG[650])|(((m[98]&~m[336]&~m[683])|(~m[98]&m[336]&m[683]))&~BiasedRNG[650])|((~m[98]&~m[336]&m[683])|(m[98]&~m[336]&m[683])|(m[98]&m[336]&m[683]))):InitCond[1146];
    m[428] = run?((((~m[99]&~m[352]&~m[684])|(m[99]&m[352]&~m[684]))&BiasedRNG[651])|(((m[99]&~m[352]&~m[684])|(~m[99]&m[352]&m[684]))&~BiasedRNG[651])|((~m[99]&~m[352]&m[684])|(m[99]&~m[352]&m[684])|(m[99]&m[352]&m[684]))):InitCond[1147];
    m[429] = run?((((~m[99]&~m[368]&~m[685])|(m[99]&m[368]&~m[685]))&BiasedRNG[652])|(((m[99]&~m[368]&~m[685])|(~m[99]&m[368]&m[685]))&~BiasedRNG[652])|((~m[99]&~m[368]&m[685])|(m[99]&~m[368]&m[685])|(m[99]&m[368]&m[685]))):InitCond[1148];
    m[430] = run?((((~m[99]&~m[384]&~m[686])|(m[99]&m[384]&~m[686]))&BiasedRNG[653])|(((m[99]&~m[384]&~m[686])|(~m[99]&m[384]&m[686]))&~BiasedRNG[653])|((~m[99]&~m[384]&m[686])|(m[99]&~m[384]&m[686])|(m[99]&m[384]&m[686]))):InitCond[1149];
    m[431] = run?((((~m[99]&~m[400]&~m[687])|(m[99]&m[400]&~m[687]))&BiasedRNG[654])|(((m[99]&~m[400]&~m[687])|(~m[99]&m[400]&m[687]))&~BiasedRNG[654])|((~m[99]&~m[400]&m[687])|(m[99]&~m[400]&m[687])|(m[99]&m[400]&m[687]))):InitCond[1150];
    m[432] = run?((((~m[100]&~m[161]&~m[688])|(m[100]&m[161]&~m[688]))&BiasedRNG[655])|(((m[100]&~m[161]&~m[688])|(~m[100]&m[161]&m[688]))&~BiasedRNG[655])|((~m[100]&~m[161]&m[688])|(m[100]&~m[161]&m[688])|(m[100]&m[161]&m[688]))):InitCond[1151];
    m[433] = run?((((~m[100]&~m[177]&~m[689])|(m[100]&m[177]&~m[689]))&BiasedRNG[656])|(((m[100]&~m[177]&~m[689])|(~m[100]&m[177]&m[689]))&~BiasedRNG[656])|((~m[100]&~m[177]&m[689])|(m[100]&~m[177]&m[689])|(m[100]&m[177]&m[689]))):InitCond[1152];
    m[434] = run?((((~m[100]&~m[193]&~m[690])|(m[100]&m[193]&~m[690]))&BiasedRNG[657])|(((m[100]&~m[193]&~m[690])|(~m[100]&m[193]&m[690]))&~BiasedRNG[657])|((~m[100]&~m[193]&m[690])|(m[100]&~m[193]&m[690])|(m[100]&m[193]&m[690]))):InitCond[1153];
    m[435] = run?((((~m[100]&~m[209]&~m[691])|(m[100]&m[209]&~m[691]))&BiasedRNG[658])|(((m[100]&~m[209]&~m[691])|(~m[100]&m[209]&m[691]))&~BiasedRNG[658])|((~m[100]&~m[209]&m[691])|(m[100]&~m[209]&m[691])|(m[100]&m[209]&m[691]))):InitCond[1154];
    m[436] = run?((((~m[101]&~m[225]&~m[692])|(m[101]&m[225]&~m[692]))&BiasedRNG[659])|(((m[101]&~m[225]&~m[692])|(~m[101]&m[225]&m[692]))&~BiasedRNG[659])|((~m[101]&~m[225]&m[692])|(m[101]&~m[225]&m[692])|(m[101]&m[225]&m[692]))):InitCond[1155];
    m[437] = run?((((~m[101]&~m[241]&~m[693])|(m[101]&m[241]&~m[693]))&BiasedRNG[660])|(((m[101]&~m[241]&~m[693])|(~m[101]&m[241]&m[693]))&~BiasedRNG[660])|((~m[101]&~m[241]&m[693])|(m[101]&~m[241]&m[693])|(m[101]&m[241]&m[693]))):InitCond[1156];
    m[438] = run?((((~m[101]&~m[257]&~m[694])|(m[101]&m[257]&~m[694]))&BiasedRNG[661])|(((m[101]&~m[257]&~m[694])|(~m[101]&m[257]&m[694]))&~BiasedRNG[661])|((~m[101]&~m[257]&m[694])|(m[101]&~m[257]&m[694])|(m[101]&m[257]&m[694]))):InitCond[1157];
    m[439] = run?((((~m[101]&~m[273]&~m[695])|(m[101]&m[273]&~m[695]))&BiasedRNG[662])|(((m[101]&~m[273]&~m[695])|(~m[101]&m[273]&m[695]))&~BiasedRNG[662])|((~m[101]&~m[273]&m[695])|(m[101]&~m[273]&m[695])|(m[101]&m[273]&m[695]))):InitCond[1158];
    m[440] = run?((((~m[102]&~m[289]&~m[696])|(m[102]&m[289]&~m[696]))&BiasedRNG[663])|(((m[102]&~m[289]&~m[696])|(~m[102]&m[289]&m[696]))&~BiasedRNG[663])|((~m[102]&~m[289]&m[696])|(m[102]&~m[289]&m[696])|(m[102]&m[289]&m[696]))):InitCond[1159];
    m[441] = run?((((~m[102]&~m[305]&~m[697])|(m[102]&m[305]&~m[697]))&BiasedRNG[664])|(((m[102]&~m[305]&~m[697])|(~m[102]&m[305]&m[697]))&~BiasedRNG[664])|((~m[102]&~m[305]&m[697])|(m[102]&~m[305]&m[697])|(m[102]&m[305]&m[697]))):InitCond[1160];
    m[442] = run?((((~m[102]&~m[321]&~m[698])|(m[102]&m[321]&~m[698]))&BiasedRNG[665])|(((m[102]&~m[321]&~m[698])|(~m[102]&m[321]&m[698]))&~BiasedRNG[665])|((~m[102]&~m[321]&m[698])|(m[102]&~m[321]&m[698])|(m[102]&m[321]&m[698]))):InitCond[1161];
    m[443] = run?((((~m[102]&~m[337]&~m[699])|(m[102]&m[337]&~m[699]))&BiasedRNG[666])|(((m[102]&~m[337]&~m[699])|(~m[102]&m[337]&m[699]))&~BiasedRNG[666])|((~m[102]&~m[337]&m[699])|(m[102]&~m[337]&m[699])|(m[102]&m[337]&m[699]))):InitCond[1162];
    m[444] = run?((((~m[103]&~m[353]&~m[700])|(m[103]&m[353]&~m[700]))&BiasedRNG[667])|(((m[103]&~m[353]&~m[700])|(~m[103]&m[353]&m[700]))&~BiasedRNG[667])|((~m[103]&~m[353]&m[700])|(m[103]&~m[353]&m[700])|(m[103]&m[353]&m[700]))):InitCond[1163];
    m[445] = run?((((~m[103]&~m[369]&~m[701])|(m[103]&m[369]&~m[701]))&BiasedRNG[668])|(((m[103]&~m[369]&~m[701])|(~m[103]&m[369]&m[701]))&~BiasedRNG[668])|((~m[103]&~m[369]&m[701])|(m[103]&~m[369]&m[701])|(m[103]&m[369]&m[701]))):InitCond[1164];
    m[446] = run?((((~m[103]&~m[385]&~m[702])|(m[103]&m[385]&~m[702]))&BiasedRNG[669])|(((m[103]&~m[385]&~m[702])|(~m[103]&m[385]&m[702]))&~BiasedRNG[669])|((~m[103]&~m[385]&m[702])|(m[103]&~m[385]&m[702])|(m[103]&m[385]&m[702]))):InitCond[1165];
    m[447] = run?((((~m[103]&~m[401]&~m[703])|(m[103]&m[401]&~m[703]))&BiasedRNG[670])|(((m[103]&~m[401]&~m[703])|(~m[103]&m[401]&m[703]))&~BiasedRNG[670])|((~m[103]&~m[401]&m[703])|(m[103]&~m[401]&m[703])|(m[103]&m[401]&m[703]))):InitCond[1166];
    m[448] = run?((((~m[104]&~m[162]&~m[704])|(m[104]&m[162]&~m[704]))&BiasedRNG[671])|(((m[104]&~m[162]&~m[704])|(~m[104]&m[162]&m[704]))&~BiasedRNG[671])|((~m[104]&~m[162]&m[704])|(m[104]&~m[162]&m[704])|(m[104]&m[162]&m[704]))):InitCond[1167];
    m[449] = run?((((~m[104]&~m[178]&~m[705])|(m[104]&m[178]&~m[705]))&BiasedRNG[672])|(((m[104]&~m[178]&~m[705])|(~m[104]&m[178]&m[705]))&~BiasedRNG[672])|((~m[104]&~m[178]&m[705])|(m[104]&~m[178]&m[705])|(m[104]&m[178]&m[705]))):InitCond[1168];
    m[450] = run?((((~m[104]&~m[194]&~m[706])|(m[104]&m[194]&~m[706]))&BiasedRNG[673])|(((m[104]&~m[194]&~m[706])|(~m[104]&m[194]&m[706]))&~BiasedRNG[673])|((~m[104]&~m[194]&m[706])|(m[104]&~m[194]&m[706])|(m[104]&m[194]&m[706]))):InitCond[1169];
    m[451] = run?((((~m[104]&~m[210]&~m[707])|(m[104]&m[210]&~m[707]))&BiasedRNG[674])|(((m[104]&~m[210]&~m[707])|(~m[104]&m[210]&m[707]))&~BiasedRNG[674])|((~m[104]&~m[210]&m[707])|(m[104]&~m[210]&m[707])|(m[104]&m[210]&m[707]))):InitCond[1170];
    m[452] = run?((((~m[105]&~m[226]&~m[708])|(m[105]&m[226]&~m[708]))&BiasedRNG[675])|(((m[105]&~m[226]&~m[708])|(~m[105]&m[226]&m[708]))&~BiasedRNG[675])|((~m[105]&~m[226]&m[708])|(m[105]&~m[226]&m[708])|(m[105]&m[226]&m[708]))):InitCond[1171];
    m[453] = run?((((~m[105]&~m[242]&~m[709])|(m[105]&m[242]&~m[709]))&BiasedRNG[676])|(((m[105]&~m[242]&~m[709])|(~m[105]&m[242]&m[709]))&~BiasedRNG[676])|((~m[105]&~m[242]&m[709])|(m[105]&~m[242]&m[709])|(m[105]&m[242]&m[709]))):InitCond[1172];
    m[454] = run?((((~m[105]&~m[258]&~m[710])|(m[105]&m[258]&~m[710]))&BiasedRNG[677])|(((m[105]&~m[258]&~m[710])|(~m[105]&m[258]&m[710]))&~BiasedRNG[677])|((~m[105]&~m[258]&m[710])|(m[105]&~m[258]&m[710])|(m[105]&m[258]&m[710]))):InitCond[1173];
    m[455] = run?((((~m[105]&~m[274]&~m[711])|(m[105]&m[274]&~m[711]))&BiasedRNG[678])|(((m[105]&~m[274]&~m[711])|(~m[105]&m[274]&m[711]))&~BiasedRNG[678])|((~m[105]&~m[274]&m[711])|(m[105]&~m[274]&m[711])|(m[105]&m[274]&m[711]))):InitCond[1174];
    m[456] = run?((((~m[106]&~m[290]&~m[712])|(m[106]&m[290]&~m[712]))&BiasedRNG[679])|(((m[106]&~m[290]&~m[712])|(~m[106]&m[290]&m[712]))&~BiasedRNG[679])|((~m[106]&~m[290]&m[712])|(m[106]&~m[290]&m[712])|(m[106]&m[290]&m[712]))):InitCond[1175];
    m[457] = run?((((~m[106]&~m[306]&~m[713])|(m[106]&m[306]&~m[713]))&BiasedRNG[680])|(((m[106]&~m[306]&~m[713])|(~m[106]&m[306]&m[713]))&~BiasedRNG[680])|((~m[106]&~m[306]&m[713])|(m[106]&~m[306]&m[713])|(m[106]&m[306]&m[713]))):InitCond[1176];
    m[458] = run?((((~m[106]&~m[322]&~m[714])|(m[106]&m[322]&~m[714]))&BiasedRNG[681])|(((m[106]&~m[322]&~m[714])|(~m[106]&m[322]&m[714]))&~BiasedRNG[681])|((~m[106]&~m[322]&m[714])|(m[106]&~m[322]&m[714])|(m[106]&m[322]&m[714]))):InitCond[1177];
    m[459] = run?((((~m[106]&~m[338]&~m[715])|(m[106]&m[338]&~m[715]))&BiasedRNG[682])|(((m[106]&~m[338]&~m[715])|(~m[106]&m[338]&m[715]))&~BiasedRNG[682])|((~m[106]&~m[338]&m[715])|(m[106]&~m[338]&m[715])|(m[106]&m[338]&m[715]))):InitCond[1178];
    m[460] = run?((((~m[107]&~m[354]&~m[716])|(m[107]&m[354]&~m[716]))&BiasedRNG[683])|(((m[107]&~m[354]&~m[716])|(~m[107]&m[354]&m[716]))&~BiasedRNG[683])|((~m[107]&~m[354]&m[716])|(m[107]&~m[354]&m[716])|(m[107]&m[354]&m[716]))):InitCond[1179];
    m[461] = run?((((~m[107]&~m[370]&~m[717])|(m[107]&m[370]&~m[717]))&BiasedRNG[684])|(((m[107]&~m[370]&~m[717])|(~m[107]&m[370]&m[717]))&~BiasedRNG[684])|((~m[107]&~m[370]&m[717])|(m[107]&~m[370]&m[717])|(m[107]&m[370]&m[717]))):InitCond[1180];
    m[462] = run?((((~m[107]&~m[386]&~m[718])|(m[107]&m[386]&~m[718]))&BiasedRNG[685])|(((m[107]&~m[386]&~m[718])|(~m[107]&m[386]&m[718]))&~BiasedRNG[685])|((~m[107]&~m[386]&m[718])|(m[107]&~m[386]&m[718])|(m[107]&m[386]&m[718]))):InitCond[1181];
    m[463] = run?((((~m[107]&~m[402]&~m[719])|(m[107]&m[402]&~m[719]))&BiasedRNG[686])|(((m[107]&~m[402]&~m[719])|(~m[107]&m[402]&m[719]))&~BiasedRNG[686])|((~m[107]&~m[402]&m[719])|(m[107]&~m[402]&m[719])|(m[107]&m[402]&m[719]))):InitCond[1182];
    m[464] = run?((((~m[108]&~m[163]&~m[720])|(m[108]&m[163]&~m[720]))&BiasedRNG[687])|(((m[108]&~m[163]&~m[720])|(~m[108]&m[163]&m[720]))&~BiasedRNG[687])|((~m[108]&~m[163]&m[720])|(m[108]&~m[163]&m[720])|(m[108]&m[163]&m[720]))):InitCond[1183];
    m[465] = run?((((~m[108]&~m[179]&~m[721])|(m[108]&m[179]&~m[721]))&BiasedRNG[688])|(((m[108]&~m[179]&~m[721])|(~m[108]&m[179]&m[721]))&~BiasedRNG[688])|((~m[108]&~m[179]&m[721])|(m[108]&~m[179]&m[721])|(m[108]&m[179]&m[721]))):InitCond[1184];
    m[466] = run?((((~m[108]&~m[195]&~m[722])|(m[108]&m[195]&~m[722]))&BiasedRNG[689])|(((m[108]&~m[195]&~m[722])|(~m[108]&m[195]&m[722]))&~BiasedRNG[689])|((~m[108]&~m[195]&m[722])|(m[108]&~m[195]&m[722])|(m[108]&m[195]&m[722]))):InitCond[1185];
    m[467] = run?((((~m[108]&~m[211]&~m[723])|(m[108]&m[211]&~m[723]))&BiasedRNG[690])|(((m[108]&~m[211]&~m[723])|(~m[108]&m[211]&m[723]))&~BiasedRNG[690])|((~m[108]&~m[211]&m[723])|(m[108]&~m[211]&m[723])|(m[108]&m[211]&m[723]))):InitCond[1186];
    m[468] = run?((((~m[109]&~m[227]&~m[724])|(m[109]&m[227]&~m[724]))&BiasedRNG[691])|(((m[109]&~m[227]&~m[724])|(~m[109]&m[227]&m[724]))&~BiasedRNG[691])|((~m[109]&~m[227]&m[724])|(m[109]&~m[227]&m[724])|(m[109]&m[227]&m[724]))):InitCond[1187];
    m[469] = run?((((~m[109]&~m[243]&~m[725])|(m[109]&m[243]&~m[725]))&BiasedRNG[692])|(((m[109]&~m[243]&~m[725])|(~m[109]&m[243]&m[725]))&~BiasedRNG[692])|((~m[109]&~m[243]&m[725])|(m[109]&~m[243]&m[725])|(m[109]&m[243]&m[725]))):InitCond[1188];
    m[470] = run?((((~m[109]&~m[259]&~m[726])|(m[109]&m[259]&~m[726]))&BiasedRNG[693])|(((m[109]&~m[259]&~m[726])|(~m[109]&m[259]&m[726]))&~BiasedRNG[693])|((~m[109]&~m[259]&m[726])|(m[109]&~m[259]&m[726])|(m[109]&m[259]&m[726]))):InitCond[1189];
    m[471] = run?((((~m[109]&~m[275]&~m[727])|(m[109]&m[275]&~m[727]))&BiasedRNG[694])|(((m[109]&~m[275]&~m[727])|(~m[109]&m[275]&m[727]))&~BiasedRNG[694])|((~m[109]&~m[275]&m[727])|(m[109]&~m[275]&m[727])|(m[109]&m[275]&m[727]))):InitCond[1190];
    m[472] = run?((((~m[110]&~m[291]&~m[728])|(m[110]&m[291]&~m[728]))&BiasedRNG[695])|(((m[110]&~m[291]&~m[728])|(~m[110]&m[291]&m[728]))&~BiasedRNG[695])|((~m[110]&~m[291]&m[728])|(m[110]&~m[291]&m[728])|(m[110]&m[291]&m[728]))):InitCond[1191];
    m[473] = run?((((~m[110]&~m[307]&~m[729])|(m[110]&m[307]&~m[729]))&BiasedRNG[696])|(((m[110]&~m[307]&~m[729])|(~m[110]&m[307]&m[729]))&~BiasedRNG[696])|((~m[110]&~m[307]&m[729])|(m[110]&~m[307]&m[729])|(m[110]&m[307]&m[729]))):InitCond[1192];
    m[474] = run?((((~m[110]&~m[323]&~m[730])|(m[110]&m[323]&~m[730]))&BiasedRNG[697])|(((m[110]&~m[323]&~m[730])|(~m[110]&m[323]&m[730]))&~BiasedRNG[697])|((~m[110]&~m[323]&m[730])|(m[110]&~m[323]&m[730])|(m[110]&m[323]&m[730]))):InitCond[1193];
    m[475] = run?((((~m[110]&~m[339]&~m[731])|(m[110]&m[339]&~m[731]))&BiasedRNG[698])|(((m[110]&~m[339]&~m[731])|(~m[110]&m[339]&m[731]))&~BiasedRNG[698])|((~m[110]&~m[339]&m[731])|(m[110]&~m[339]&m[731])|(m[110]&m[339]&m[731]))):InitCond[1194];
    m[476] = run?((((~m[111]&~m[355]&~m[732])|(m[111]&m[355]&~m[732]))&BiasedRNG[699])|(((m[111]&~m[355]&~m[732])|(~m[111]&m[355]&m[732]))&~BiasedRNG[699])|((~m[111]&~m[355]&m[732])|(m[111]&~m[355]&m[732])|(m[111]&m[355]&m[732]))):InitCond[1195];
    m[477] = run?((((~m[111]&~m[371]&~m[733])|(m[111]&m[371]&~m[733]))&BiasedRNG[700])|(((m[111]&~m[371]&~m[733])|(~m[111]&m[371]&m[733]))&~BiasedRNG[700])|((~m[111]&~m[371]&m[733])|(m[111]&~m[371]&m[733])|(m[111]&m[371]&m[733]))):InitCond[1196];
    m[478] = run?((((~m[111]&~m[387]&~m[734])|(m[111]&m[387]&~m[734]))&BiasedRNG[701])|(((m[111]&~m[387]&~m[734])|(~m[111]&m[387]&m[734]))&~BiasedRNG[701])|((~m[111]&~m[387]&m[734])|(m[111]&~m[387]&m[734])|(m[111]&m[387]&m[734]))):InitCond[1197];
    m[479] = run?((((~m[111]&~m[403]&~m[735])|(m[111]&m[403]&~m[735]))&BiasedRNG[702])|(((m[111]&~m[403]&~m[735])|(~m[111]&m[403]&m[735]))&~BiasedRNG[702])|((~m[111]&~m[403]&m[735])|(m[111]&~m[403]&m[735])|(m[111]&m[403]&m[735]))):InitCond[1198];
    m[480] = run?((((~m[112]&~m[164]&~m[736])|(m[112]&m[164]&~m[736]))&BiasedRNG[703])|(((m[112]&~m[164]&~m[736])|(~m[112]&m[164]&m[736]))&~BiasedRNG[703])|((~m[112]&~m[164]&m[736])|(m[112]&~m[164]&m[736])|(m[112]&m[164]&m[736]))):InitCond[1199];
    m[481] = run?((((~m[112]&~m[180]&~m[737])|(m[112]&m[180]&~m[737]))&BiasedRNG[704])|(((m[112]&~m[180]&~m[737])|(~m[112]&m[180]&m[737]))&~BiasedRNG[704])|((~m[112]&~m[180]&m[737])|(m[112]&~m[180]&m[737])|(m[112]&m[180]&m[737]))):InitCond[1200];
    m[482] = run?((((~m[112]&~m[196]&~m[738])|(m[112]&m[196]&~m[738]))&BiasedRNG[705])|(((m[112]&~m[196]&~m[738])|(~m[112]&m[196]&m[738]))&~BiasedRNG[705])|((~m[112]&~m[196]&m[738])|(m[112]&~m[196]&m[738])|(m[112]&m[196]&m[738]))):InitCond[1201];
    m[483] = run?((((~m[112]&~m[212]&~m[739])|(m[112]&m[212]&~m[739]))&BiasedRNG[706])|(((m[112]&~m[212]&~m[739])|(~m[112]&m[212]&m[739]))&~BiasedRNG[706])|((~m[112]&~m[212]&m[739])|(m[112]&~m[212]&m[739])|(m[112]&m[212]&m[739]))):InitCond[1202];
    m[484] = run?((((~m[113]&~m[228]&~m[740])|(m[113]&m[228]&~m[740]))&BiasedRNG[707])|(((m[113]&~m[228]&~m[740])|(~m[113]&m[228]&m[740]))&~BiasedRNG[707])|((~m[113]&~m[228]&m[740])|(m[113]&~m[228]&m[740])|(m[113]&m[228]&m[740]))):InitCond[1203];
    m[485] = run?((((~m[113]&~m[244]&~m[741])|(m[113]&m[244]&~m[741]))&BiasedRNG[708])|(((m[113]&~m[244]&~m[741])|(~m[113]&m[244]&m[741]))&~BiasedRNG[708])|((~m[113]&~m[244]&m[741])|(m[113]&~m[244]&m[741])|(m[113]&m[244]&m[741]))):InitCond[1204];
    m[486] = run?((((~m[113]&~m[260]&~m[742])|(m[113]&m[260]&~m[742]))&BiasedRNG[709])|(((m[113]&~m[260]&~m[742])|(~m[113]&m[260]&m[742]))&~BiasedRNG[709])|((~m[113]&~m[260]&m[742])|(m[113]&~m[260]&m[742])|(m[113]&m[260]&m[742]))):InitCond[1205];
    m[487] = run?((((~m[113]&~m[276]&~m[743])|(m[113]&m[276]&~m[743]))&BiasedRNG[710])|(((m[113]&~m[276]&~m[743])|(~m[113]&m[276]&m[743]))&~BiasedRNG[710])|((~m[113]&~m[276]&m[743])|(m[113]&~m[276]&m[743])|(m[113]&m[276]&m[743]))):InitCond[1206];
    m[488] = run?((((~m[114]&~m[292]&~m[744])|(m[114]&m[292]&~m[744]))&BiasedRNG[711])|(((m[114]&~m[292]&~m[744])|(~m[114]&m[292]&m[744]))&~BiasedRNG[711])|((~m[114]&~m[292]&m[744])|(m[114]&~m[292]&m[744])|(m[114]&m[292]&m[744]))):InitCond[1207];
    m[489] = run?((((~m[114]&~m[308]&~m[745])|(m[114]&m[308]&~m[745]))&BiasedRNG[712])|(((m[114]&~m[308]&~m[745])|(~m[114]&m[308]&m[745]))&~BiasedRNG[712])|((~m[114]&~m[308]&m[745])|(m[114]&~m[308]&m[745])|(m[114]&m[308]&m[745]))):InitCond[1208];
    m[490] = run?((((~m[114]&~m[324]&~m[746])|(m[114]&m[324]&~m[746]))&BiasedRNG[713])|(((m[114]&~m[324]&~m[746])|(~m[114]&m[324]&m[746]))&~BiasedRNG[713])|((~m[114]&~m[324]&m[746])|(m[114]&~m[324]&m[746])|(m[114]&m[324]&m[746]))):InitCond[1209];
    m[491] = run?((((~m[114]&~m[340]&~m[747])|(m[114]&m[340]&~m[747]))&BiasedRNG[714])|(((m[114]&~m[340]&~m[747])|(~m[114]&m[340]&m[747]))&~BiasedRNG[714])|((~m[114]&~m[340]&m[747])|(m[114]&~m[340]&m[747])|(m[114]&m[340]&m[747]))):InitCond[1210];
    m[492] = run?((((~m[115]&~m[356]&~m[748])|(m[115]&m[356]&~m[748]))&BiasedRNG[715])|(((m[115]&~m[356]&~m[748])|(~m[115]&m[356]&m[748]))&~BiasedRNG[715])|((~m[115]&~m[356]&m[748])|(m[115]&~m[356]&m[748])|(m[115]&m[356]&m[748]))):InitCond[1211];
    m[493] = run?((((~m[115]&~m[372]&~m[749])|(m[115]&m[372]&~m[749]))&BiasedRNG[716])|(((m[115]&~m[372]&~m[749])|(~m[115]&m[372]&m[749]))&~BiasedRNG[716])|((~m[115]&~m[372]&m[749])|(m[115]&~m[372]&m[749])|(m[115]&m[372]&m[749]))):InitCond[1212];
    m[494] = run?((((~m[115]&~m[388]&~m[750])|(m[115]&m[388]&~m[750]))&BiasedRNG[717])|(((m[115]&~m[388]&~m[750])|(~m[115]&m[388]&m[750]))&~BiasedRNG[717])|((~m[115]&~m[388]&m[750])|(m[115]&~m[388]&m[750])|(m[115]&m[388]&m[750]))):InitCond[1213];
    m[495] = run?((((~m[115]&~m[404]&~m[751])|(m[115]&m[404]&~m[751]))&BiasedRNG[718])|(((m[115]&~m[404]&~m[751])|(~m[115]&m[404]&m[751]))&~BiasedRNG[718])|((~m[115]&~m[404]&m[751])|(m[115]&~m[404]&m[751])|(m[115]&m[404]&m[751]))):InitCond[1214];
    m[496] = run?((((~m[116]&~m[165]&~m[752])|(m[116]&m[165]&~m[752]))&BiasedRNG[719])|(((m[116]&~m[165]&~m[752])|(~m[116]&m[165]&m[752]))&~BiasedRNG[719])|((~m[116]&~m[165]&m[752])|(m[116]&~m[165]&m[752])|(m[116]&m[165]&m[752]))):InitCond[1215];
    m[497] = run?((((~m[116]&~m[181]&~m[753])|(m[116]&m[181]&~m[753]))&BiasedRNG[720])|(((m[116]&~m[181]&~m[753])|(~m[116]&m[181]&m[753]))&~BiasedRNG[720])|((~m[116]&~m[181]&m[753])|(m[116]&~m[181]&m[753])|(m[116]&m[181]&m[753]))):InitCond[1216];
    m[498] = run?((((~m[116]&~m[197]&~m[754])|(m[116]&m[197]&~m[754]))&BiasedRNG[721])|(((m[116]&~m[197]&~m[754])|(~m[116]&m[197]&m[754]))&~BiasedRNG[721])|((~m[116]&~m[197]&m[754])|(m[116]&~m[197]&m[754])|(m[116]&m[197]&m[754]))):InitCond[1217];
    m[499] = run?((((~m[116]&~m[213]&~m[755])|(m[116]&m[213]&~m[755]))&BiasedRNG[722])|(((m[116]&~m[213]&~m[755])|(~m[116]&m[213]&m[755]))&~BiasedRNG[722])|((~m[116]&~m[213]&m[755])|(m[116]&~m[213]&m[755])|(m[116]&m[213]&m[755]))):InitCond[1218];
    m[500] = run?((((~m[117]&~m[229]&~m[756])|(m[117]&m[229]&~m[756]))&BiasedRNG[723])|(((m[117]&~m[229]&~m[756])|(~m[117]&m[229]&m[756]))&~BiasedRNG[723])|((~m[117]&~m[229]&m[756])|(m[117]&~m[229]&m[756])|(m[117]&m[229]&m[756]))):InitCond[1219];
    m[501] = run?((((~m[117]&~m[245]&~m[757])|(m[117]&m[245]&~m[757]))&BiasedRNG[724])|(((m[117]&~m[245]&~m[757])|(~m[117]&m[245]&m[757]))&~BiasedRNG[724])|((~m[117]&~m[245]&m[757])|(m[117]&~m[245]&m[757])|(m[117]&m[245]&m[757]))):InitCond[1220];
    m[502] = run?((((~m[117]&~m[261]&~m[758])|(m[117]&m[261]&~m[758]))&BiasedRNG[725])|(((m[117]&~m[261]&~m[758])|(~m[117]&m[261]&m[758]))&~BiasedRNG[725])|((~m[117]&~m[261]&m[758])|(m[117]&~m[261]&m[758])|(m[117]&m[261]&m[758]))):InitCond[1221];
    m[503] = run?((((~m[117]&~m[277]&~m[759])|(m[117]&m[277]&~m[759]))&BiasedRNG[726])|(((m[117]&~m[277]&~m[759])|(~m[117]&m[277]&m[759]))&~BiasedRNG[726])|((~m[117]&~m[277]&m[759])|(m[117]&~m[277]&m[759])|(m[117]&m[277]&m[759]))):InitCond[1222];
    m[504] = run?((((~m[118]&~m[293]&~m[760])|(m[118]&m[293]&~m[760]))&BiasedRNG[727])|(((m[118]&~m[293]&~m[760])|(~m[118]&m[293]&m[760]))&~BiasedRNG[727])|((~m[118]&~m[293]&m[760])|(m[118]&~m[293]&m[760])|(m[118]&m[293]&m[760]))):InitCond[1223];
    m[505] = run?((((~m[118]&~m[309]&~m[761])|(m[118]&m[309]&~m[761]))&BiasedRNG[728])|(((m[118]&~m[309]&~m[761])|(~m[118]&m[309]&m[761]))&~BiasedRNG[728])|((~m[118]&~m[309]&m[761])|(m[118]&~m[309]&m[761])|(m[118]&m[309]&m[761]))):InitCond[1224];
    m[506] = run?((((~m[118]&~m[325]&~m[762])|(m[118]&m[325]&~m[762]))&BiasedRNG[729])|(((m[118]&~m[325]&~m[762])|(~m[118]&m[325]&m[762]))&~BiasedRNG[729])|((~m[118]&~m[325]&m[762])|(m[118]&~m[325]&m[762])|(m[118]&m[325]&m[762]))):InitCond[1225];
    m[507] = run?((((~m[118]&~m[341]&~m[763])|(m[118]&m[341]&~m[763]))&BiasedRNG[730])|(((m[118]&~m[341]&~m[763])|(~m[118]&m[341]&m[763]))&~BiasedRNG[730])|((~m[118]&~m[341]&m[763])|(m[118]&~m[341]&m[763])|(m[118]&m[341]&m[763]))):InitCond[1226];
    m[508] = run?((((~m[119]&~m[357]&~m[764])|(m[119]&m[357]&~m[764]))&BiasedRNG[731])|(((m[119]&~m[357]&~m[764])|(~m[119]&m[357]&m[764]))&~BiasedRNG[731])|((~m[119]&~m[357]&m[764])|(m[119]&~m[357]&m[764])|(m[119]&m[357]&m[764]))):InitCond[1227];
    m[509] = run?((((~m[119]&~m[373]&~m[765])|(m[119]&m[373]&~m[765]))&BiasedRNG[732])|(((m[119]&~m[373]&~m[765])|(~m[119]&m[373]&m[765]))&~BiasedRNG[732])|((~m[119]&~m[373]&m[765])|(m[119]&~m[373]&m[765])|(m[119]&m[373]&m[765]))):InitCond[1228];
    m[510] = run?((((~m[119]&~m[389]&~m[766])|(m[119]&m[389]&~m[766]))&BiasedRNG[733])|(((m[119]&~m[389]&~m[766])|(~m[119]&m[389]&m[766]))&~BiasedRNG[733])|((~m[119]&~m[389]&m[766])|(m[119]&~m[389]&m[766])|(m[119]&m[389]&m[766]))):InitCond[1229];
    m[511] = run?((((~m[119]&~m[405]&~m[767])|(m[119]&m[405]&~m[767]))&BiasedRNG[734])|(((m[119]&~m[405]&~m[767])|(~m[119]&m[405]&m[767]))&~BiasedRNG[734])|((~m[119]&~m[405]&m[767])|(m[119]&~m[405]&m[767])|(m[119]&m[405]&m[767]))):InitCond[1230];
    m[512] = run?((((~m[120]&~m[166]&~m[768])|(m[120]&m[166]&~m[768]))&BiasedRNG[735])|(((m[120]&~m[166]&~m[768])|(~m[120]&m[166]&m[768]))&~BiasedRNG[735])|((~m[120]&~m[166]&m[768])|(m[120]&~m[166]&m[768])|(m[120]&m[166]&m[768]))):InitCond[1231];
    m[513] = run?((((~m[120]&~m[182]&~m[769])|(m[120]&m[182]&~m[769]))&BiasedRNG[736])|(((m[120]&~m[182]&~m[769])|(~m[120]&m[182]&m[769]))&~BiasedRNG[736])|((~m[120]&~m[182]&m[769])|(m[120]&~m[182]&m[769])|(m[120]&m[182]&m[769]))):InitCond[1232];
    m[514] = run?((((~m[120]&~m[198]&~m[770])|(m[120]&m[198]&~m[770]))&BiasedRNG[737])|(((m[120]&~m[198]&~m[770])|(~m[120]&m[198]&m[770]))&~BiasedRNG[737])|((~m[120]&~m[198]&m[770])|(m[120]&~m[198]&m[770])|(m[120]&m[198]&m[770]))):InitCond[1233];
    m[515] = run?((((~m[120]&~m[214]&~m[771])|(m[120]&m[214]&~m[771]))&BiasedRNG[738])|(((m[120]&~m[214]&~m[771])|(~m[120]&m[214]&m[771]))&~BiasedRNG[738])|((~m[120]&~m[214]&m[771])|(m[120]&~m[214]&m[771])|(m[120]&m[214]&m[771]))):InitCond[1234];
    m[516] = run?((((~m[121]&~m[230]&~m[772])|(m[121]&m[230]&~m[772]))&BiasedRNG[739])|(((m[121]&~m[230]&~m[772])|(~m[121]&m[230]&m[772]))&~BiasedRNG[739])|((~m[121]&~m[230]&m[772])|(m[121]&~m[230]&m[772])|(m[121]&m[230]&m[772]))):InitCond[1235];
    m[517] = run?((((~m[121]&~m[246]&~m[773])|(m[121]&m[246]&~m[773]))&BiasedRNG[740])|(((m[121]&~m[246]&~m[773])|(~m[121]&m[246]&m[773]))&~BiasedRNG[740])|((~m[121]&~m[246]&m[773])|(m[121]&~m[246]&m[773])|(m[121]&m[246]&m[773]))):InitCond[1236];
    m[518] = run?((((~m[121]&~m[262]&~m[774])|(m[121]&m[262]&~m[774]))&BiasedRNG[741])|(((m[121]&~m[262]&~m[774])|(~m[121]&m[262]&m[774]))&~BiasedRNG[741])|((~m[121]&~m[262]&m[774])|(m[121]&~m[262]&m[774])|(m[121]&m[262]&m[774]))):InitCond[1237];
    m[519] = run?((((~m[121]&~m[278]&~m[775])|(m[121]&m[278]&~m[775]))&BiasedRNG[742])|(((m[121]&~m[278]&~m[775])|(~m[121]&m[278]&m[775]))&~BiasedRNG[742])|((~m[121]&~m[278]&m[775])|(m[121]&~m[278]&m[775])|(m[121]&m[278]&m[775]))):InitCond[1238];
    m[520] = run?((((~m[122]&~m[294]&~m[776])|(m[122]&m[294]&~m[776]))&BiasedRNG[743])|(((m[122]&~m[294]&~m[776])|(~m[122]&m[294]&m[776]))&~BiasedRNG[743])|((~m[122]&~m[294]&m[776])|(m[122]&~m[294]&m[776])|(m[122]&m[294]&m[776]))):InitCond[1239];
    m[521] = run?((((~m[122]&~m[310]&~m[777])|(m[122]&m[310]&~m[777]))&BiasedRNG[744])|(((m[122]&~m[310]&~m[777])|(~m[122]&m[310]&m[777]))&~BiasedRNG[744])|((~m[122]&~m[310]&m[777])|(m[122]&~m[310]&m[777])|(m[122]&m[310]&m[777]))):InitCond[1240];
    m[522] = run?((((~m[122]&~m[326]&~m[778])|(m[122]&m[326]&~m[778]))&BiasedRNG[745])|(((m[122]&~m[326]&~m[778])|(~m[122]&m[326]&m[778]))&~BiasedRNG[745])|((~m[122]&~m[326]&m[778])|(m[122]&~m[326]&m[778])|(m[122]&m[326]&m[778]))):InitCond[1241];
    m[523] = run?((((~m[122]&~m[342]&~m[779])|(m[122]&m[342]&~m[779]))&BiasedRNG[746])|(((m[122]&~m[342]&~m[779])|(~m[122]&m[342]&m[779]))&~BiasedRNG[746])|((~m[122]&~m[342]&m[779])|(m[122]&~m[342]&m[779])|(m[122]&m[342]&m[779]))):InitCond[1242];
    m[524] = run?((((~m[123]&~m[358]&~m[780])|(m[123]&m[358]&~m[780]))&BiasedRNG[747])|(((m[123]&~m[358]&~m[780])|(~m[123]&m[358]&m[780]))&~BiasedRNG[747])|((~m[123]&~m[358]&m[780])|(m[123]&~m[358]&m[780])|(m[123]&m[358]&m[780]))):InitCond[1243];
    m[525] = run?((((~m[123]&~m[374]&~m[781])|(m[123]&m[374]&~m[781]))&BiasedRNG[748])|(((m[123]&~m[374]&~m[781])|(~m[123]&m[374]&m[781]))&~BiasedRNG[748])|((~m[123]&~m[374]&m[781])|(m[123]&~m[374]&m[781])|(m[123]&m[374]&m[781]))):InitCond[1244];
    m[526] = run?((((~m[123]&~m[390]&~m[782])|(m[123]&m[390]&~m[782]))&BiasedRNG[749])|(((m[123]&~m[390]&~m[782])|(~m[123]&m[390]&m[782]))&~BiasedRNG[749])|((~m[123]&~m[390]&m[782])|(m[123]&~m[390]&m[782])|(m[123]&m[390]&m[782]))):InitCond[1245];
    m[527] = run?((((~m[123]&~m[406]&~m[783])|(m[123]&m[406]&~m[783]))&BiasedRNG[750])|(((m[123]&~m[406]&~m[783])|(~m[123]&m[406]&m[783]))&~BiasedRNG[750])|((~m[123]&~m[406]&m[783])|(m[123]&~m[406]&m[783])|(m[123]&m[406]&m[783]))):InitCond[1246];
    m[528] = run?((((~m[124]&~m[167]&~m[784])|(m[124]&m[167]&~m[784]))&BiasedRNG[751])|(((m[124]&~m[167]&~m[784])|(~m[124]&m[167]&m[784]))&~BiasedRNG[751])|((~m[124]&~m[167]&m[784])|(m[124]&~m[167]&m[784])|(m[124]&m[167]&m[784]))):InitCond[1247];
    m[529] = run?((((~m[124]&~m[183]&~m[785])|(m[124]&m[183]&~m[785]))&BiasedRNG[752])|(((m[124]&~m[183]&~m[785])|(~m[124]&m[183]&m[785]))&~BiasedRNG[752])|((~m[124]&~m[183]&m[785])|(m[124]&~m[183]&m[785])|(m[124]&m[183]&m[785]))):InitCond[1248];
    m[530] = run?((((~m[124]&~m[199]&~m[786])|(m[124]&m[199]&~m[786]))&BiasedRNG[753])|(((m[124]&~m[199]&~m[786])|(~m[124]&m[199]&m[786]))&~BiasedRNG[753])|((~m[124]&~m[199]&m[786])|(m[124]&~m[199]&m[786])|(m[124]&m[199]&m[786]))):InitCond[1249];
    m[531] = run?((((~m[124]&~m[215]&~m[787])|(m[124]&m[215]&~m[787]))&BiasedRNG[754])|(((m[124]&~m[215]&~m[787])|(~m[124]&m[215]&m[787]))&~BiasedRNG[754])|((~m[124]&~m[215]&m[787])|(m[124]&~m[215]&m[787])|(m[124]&m[215]&m[787]))):InitCond[1250];
    m[532] = run?((((~m[125]&~m[231]&~m[788])|(m[125]&m[231]&~m[788]))&BiasedRNG[755])|(((m[125]&~m[231]&~m[788])|(~m[125]&m[231]&m[788]))&~BiasedRNG[755])|((~m[125]&~m[231]&m[788])|(m[125]&~m[231]&m[788])|(m[125]&m[231]&m[788]))):InitCond[1251];
    m[533] = run?((((~m[125]&~m[247]&~m[789])|(m[125]&m[247]&~m[789]))&BiasedRNG[756])|(((m[125]&~m[247]&~m[789])|(~m[125]&m[247]&m[789]))&~BiasedRNG[756])|((~m[125]&~m[247]&m[789])|(m[125]&~m[247]&m[789])|(m[125]&m[247]&m[789]))):InitCond[1252];
    m[534] = run?((((~m[125]&~m[263]&~m[790])|(m[125]&m[263]&~m[790]))&BiasedRNG[757])|(((m[125]&~m[263]&~m[790])|(~m[125]&m[263]&m[790]))&~BiasedRNG[757])|((~m[125]&~m[263]&m[790])|(m[125]&~m[263]&m[790])|(m[125]&m[263]&m[790]))):InitCond[1253];
    m[535] = run?((((~m[125]&~m[279]&~m[791])|(m[125]&m[279]&~m[791]))&BiasedRNG[758])|(((m[125]&~m[279]&~m[791])|(~m[125]&m[279]&m[791]))&~BiasedRNG[758])|((~m[125]&~m[279]&m[791])|(m[125]&~m[279]&m[791])|(m[125]&m[279]&m[791]))):InitCond[1254];
    m[536] = run?((((~m[126]&~m[295]&~m[792])|(m[126]&m[295]&~m[792]))&BiasedRNG[759])|(((m[126]&~m[295]&~m[792])|(~m[126]&m[295]&m[792]))&~BiasedRNG[759])|((~m[126]&~m[295]&m[792])|(m[126]&~m[295]&m[792])|(m[126]&m[295]&m[792]))):InitCond[1255];
    m[537] = run?((((~m[126]&~m[311]&~m[793])|(m[126]&m[311]&~m[793]))&BiasedRNG[760])|(((m[126]&~m[311]&~m[793])|(~m[126]&m[311]&m[793]))&~BiasedRNG[760])|((~m[126]&~m[311]&m[793])|(m[126]&~m[311]&m[793])|(m[126]&m[311]&m[793]))):InitCond[1256];
    m[538] = run?((((~m[126]&~m[327]&~m[794])|(m[126]&m[327]&~m[794]))&BiasedRNG[761])|(((m[126]&~m[327]&~m[794])|(~m[126]&m[327]&m[794]))&~BiasedRNG[761])|((~m[126]&~m[327]&m[794])|(m[126]&~m[327]&m[794])|(m[126]&m[327]&m[794]))):InitCond[1257];
    m[539] = run?((((~m[126]&~m[343]&~m[795])|(m[126]&m[343]&~m[795]))&BiasedRNG[762])|(((m[126]&~m[343]&~m[795])|(~m[126]&m[343]&m[795]))&~BiasedRNG[762])|((~m[126]&~m[343]&m[795])|(m[126]&~m[343]&m[795])|(m[126]&m[343]&m[795]))):InitCond[1258];
    m[540] = run?((((~m[127]&~m[359]&~m[796])|(m[127]&m[359]&~m[796]))&BiasedRNG[763])|(((m[127]&~m[359]&~m[796])|(~m[127]&m[359]&m[796]))&~BiasedRNG[763])|((~m[127]&~m[359]&m[796])|(m[127]&~m[359]&m[796])|(m[127]&m[359]&m[796]))):InitCond[1259];
    m[541] = run?((((~m[127]&~m[375]&~m[797])|(m[127]&m[375]&~m[797]))&BiasedRNG[764])|(((m[127]&~m[375]&~m[797])|(~m[127]&m[375]&m[797]))&~BiasedRNG[764])|((~m[127]&~m[375]&m[797])|(m[127]&~m[375]&m[797])|(m[127]&m[375]&m[797]))):InitCond[1260];
    m[542] = run?((((~m[127]&~m[391]&~m[798])|(m[127]&m[391]&~m[798]))&BiasedRNG[765])|(((m[127]&~m[391]&~m[798])|(~m[127]&m[391]&m[798]))&~BiasedRNG[765])|((~m[127]&~m[391]&m[798])|(m[127]&~m[391]&m[798])|(m[127]&m[391]&m[798]))):InitCond[1261];
    m[543] = run?((((~m[127]&~m[407]&~m[799])|(m[127]&m[407]&~m[799]))&BiasedRNG[766])|(((m[127]&~m[407]&~m[799])|(~m[127]&m[407]&m[799]))&~BiasedRNG[766])|((~m[127]&~m[407]&m[799])|(m[127]&~m[407]&m[799])|(m[127]&m[407]&m[799]))):InitCond[1262];
    m[544] = run?((((~m[128]&~m[168]&~m[800])|(m[128]&m[168]&~m[800]))&BiasedRNG[767])|(((m[128]&~m[168]&~m[800])|(~m[128]&m[168]&m[800]))&~BiasedRNG[767])|((~m[128]&~m[168]&m[800])|(m[128]&~m[168]&m[800])|(m[128]&m[168]&m[800]))):InitCond[1263];
    m[545] = run?((((~m[128]&~m[184]&~m[801])|(m[128]&m[184]&~m[801]))&BiasedRNG[768])|(((m[128]&~m[184]&~m[801])|(~m[128]&m[184]&m[801]))&~BiasedRNG[768])|((~m[128]&~m[184]&m[801])|(m[128]&~m[184]&m[801])|(m[128]&m[184]&m[801]))):InitCond[1264];
    m[546] = run?((((~m[128]&~m[200]&~m[802])|(m[128]&m[200]&~m[802]))&BiasedRNG[769])|(((m[128]&~m[200]&~m[802])|(~m[128]&m[200]&m[802]))&~BiasedRNG[769])|((~m[128]&~m[200]&m[802])|(m[128]&~m[200]&m[802])|(m[128]&m[200]&m[802]))):InitCond[1265];
    m[547] = run?((((~m[128]&~m[216]&~m[803])|(m[128]&m[216]&~m[803]))&BiasedRNG[770])|(((m[128]&~m[216]&~m[803])|(~m[128]&m[216]&m[803]))&~BiasedRNG[770])|((~m[128]&~m[216]&m[803])|(m[128]&~m[216]&m[803])|(m[128]&m[216]&m[803]))):InitCond[1266];
    m[548] = run?((((~m[129]&~m[232]&~m[804])|(m[129]&m[232]&~m[804]))&BiasedRNG[771])|(((m[129]&~m[232]&~m[804])|(~m[129]&m[232]&m[804]))&~BiasedRNG[771])|((~m[129]&~m[232]&m[804])|(m[129]&~m[232]&m[804])|(m[129]&m[232]&m[804]))):InitCond[1267];
    m[549] = run?((((~m[129]&~m[248]&~m[805])|(m[129]&m[248]&~m[805]))&BiasedRNG[772])|(((m[129]&~m[248]&~m[805])|(~m[129]&m[248]&m[805]))&~BiasedRNG[772])|((~m[129]&~m[248]&m[805])|(m[129]&~m[248]&m[805])|(m[129]&m[248]&m[805]))):InitCond[1268];
    m[550] = run?((((~m[129]&~m[264]&~m[806])|(m[129]&m[264]&~m[806]))&BiasedRNG[773])|(((m[129]&~m[264]&~m[806])|(~m[129]&m[264]&m[806]))&~BiasedRNG[773])|((~m[129]&~m[264]&m[806])|(m[129]&~m[264]&m[806])|(m[129]&m[264]&m[806]))):InitCond[1269];
    m[551] = run?((((~m[129]&~m[280]&~m[807])|(m[129]&m[280]&~m[807]))&BiasedRNG[774])|(((m[129]&~m[280]&~m[807])|(~m[129]&m[280]&m[807]))&~BiasedRNG[774])|((~m[129]&~m[280]&m[807])|(m[129]&~m[280]&m[807])|(m[129]&m[280]&m[807]))):InitCond[1270];
    m[552] = run?((((~m[130]&~m[296]&~m[808])|(m[130]&m[296]&~m[808]))&BiasedRNG[775])|(((m[130]&~m[296]&~m[808])|(~m[130]&m[296]&m[808]))&~BiasedRNG[775])|((~m[130]&~m[296]&m[808])|(m[130]&~m[296]&m[808])|(m[130]&m[296]&m[808]))):InitCond[1271];
    m[553] = run?((((~m[130]&~m[312]&~m[809])|(m[130]&m[312]&~m[809]))&BiasedRNG[776])|(((m[130]&~m[312]&~m[809])|(~m[130]&m[312]&m[809]))&~BiasedRNG[776])|((~m[130]&~m[312]&m[809])|(m[130]&~m[312]&m[809])|(m[130]&m[312]&m[809]))):InitCond[1272];
    m[554] = run?((((~m[130]&~m[328]&~m[810])|(m[130]&m[328]&~m[810]))&BiasedRNG[777])|(((m[130]&~m[328]&~m[810])|(~m[130]&m[328]&m[810]))&~BiasedRNG[777])|((~m[130]&~m[328]&m[810])|(m[130]&~m[328]&m[810])|(m[130]&m[328]&m[810]))):InitCond[1273];
    m[555] = run?((((~m[130]&~m[344]&~m[811])|(m[130]&m[344]&~m[811]))&BiasedRNG[778])|(((m[130]&~m[344]&~m[811])|(~m[130]&m[344]&m[811]))&~BiasedRNG[778])|((~m[130]&~m[344]&m[811])|(m[130]&~m[344]&m[811])|(m[130]&m[344]&m[811]))):InitCond[1274];
    m[556] = run?((((~m[131]&~m[360]&~m[812])|(m[131]&m[360]&~m[812]))&BiasedRNG[779])|(((m[131]&~m[360]&~m[812])|(~m[131]&m[360]&m[812]))&~BiasedRNG[779])|((~m[131]&~m[360]&m[812])|(m[131]&~m[360]&m[812])|(m[131]&m[360]&m[812]))):InitCond[1275];
    m[557] = run?((((~m[131]&~m[376]&~m[813])|(m[131]&m[376]&~m[813]))&BiasedRNG[780])|(((m[131]&~m[376]&~m[813])|(~m[131]&m[376]&m[813]))&~BiasedRNG[780])|((~m[131]&~m[376]&m[813])|(m[131]&~m[376]&m[813])|(m[131]&m[376]&m[813]))):InitCond[1276];
    m[558] = run?((((~m[131]&~m[392]&~m[814])|(m[131]&m[392]&~m[814]))&BiasedRNG[781])|(((m[131]&~m[392]&~m[814])|(~m[131]&m[392]&m[814]))&~BiasedRNG[781])|((~m[131]&~m[392]&m[814])|(m[131]&~m[392]&m[814])|(m[131]&m[392]&m[814]))):InitCond[1277];
    m[559] = run?((((~m[131]&~m[408]&~m[815])|(m[131]&m[408]&~m[815]))&BiasedRNG[782])|(((m[131]&~m[408]&~m[815])|(~m[131]&m[408]&m[815]))&~BiasedRNG[782])|((~m[131]&~m[408]&m[815])|(m[131]&~m[408]&m[815])|(m[131]&m[408]&m[815]))):InitCond[1278];
    m[560] = run?((((~m[132]&~m[169]&~m[816])|(m[132]&m[169]&~m[816]))&BiasedRNG[783])|(((m[132]&~m[169]&~m[816])|(~m[132]&m[169]&m[816]))&~BiasedRNG[783])|((~m[132]&~m[169]&m[816])|(m[132]&~m[169]&m[816])|(m[132]&m[169]&m[816]))):InitCond[1279];
    m[561] = run?((((~m[132]&~m[185]&~m[817])|(m[132]&m[185]&~m[817]))&BiasedRNG[784])|(((m[132]&~m[185]&~m[817])|(~m[132]&m[185]&m[817]))&~BiasedRNG[784])|((~m[132]&~m[185]&m[817])|(m[132]&~m[185]&m[817])|(m[132]&m[185]&m[817]))):InitCond[1280];
    m[562] = run?((((~m[132]&~m[201]&~m[818])|(m[132]&m[201]&~m[818]))&BiasedRNG[785])|(((m[132]&~m[201]&~m[818])|(~m[132]&m[201]&m[818]))&~BiasedRNG[785])|((~m[132]&~m[201]&m[818])|(m[132]&~m[201]&m[818])|(m[132]&m[201]&m[818]))):InitCond[1281];
    m[563] = run?((((~m[132]&~m[217]&~m[819])|(m[132]&m[217]&~m[819]))&BiasedRNG[786])|(((m[132]&~m[217]&~m[819])|(~m[132]&m[217]&m[819]))&~BiasedRNG[786])|((~m[132]&~m[217]&m[819])|(m[132]&~m[217]&m[819])|(m[132]&m[217]&m[819]))):InitCond[1282];
    m[564] = run?((((~m[133]&~m[233]&~m[820])|(m[133]&m[233]&~m[820]))&BiasedRNG[787])|(((m[133]&~m[233]&~m[820])|(~m[133]&m[233]&m[820]))&~BiasedRNG[787])|((~m[133]&~m[233]&m[820])|(m[133]&~m[233]&m[820])|(m[133]&m[233]&m[820]))):InitCond[1283];
    m[565] = run?((((~m[133]&~m[249]&~m[821])|(m[133]&m[249]&~m[821]))&BiasedRNG[788])|(((m[133]&~m[249]&~m[821])|(~m[133]&m[249]&m[821]))&~BiasedRNG[788])|((~m[133]&~m[249]&m[821])|(m[133]&~m[249]&m[821])|(m[133]&m[249]&m[821]))):InitCond[1284];
    m[566] = run?((((~m[133]&~m[265]&~m[822])|(m[133]&m[265]&~m[822]))&BiasedRNG[789])|(((m[133]&~m[265]&~m[822])|(~m[133]&m[265]&m[822]))&~BiasedRNG[789])|((~m[133]&~m[265]&m[822])|(m[133]&~m[265]&m[822])|(m[133]&m[265]&m[822]))):InitCond[1285];
    m[567] = run?((((~m[133]&~m[281]&~m[823])|(m[133]&m[281]&~m[823]))&BiasedRNG[790])|(((m[133]&~m[281]&~m[823])|(~m[133]&m[281]&m[823]))&~BiasedRNG[790])|((~m[133]&~m[281]&m[823])|(m[133]&~m[281]&m[823])|(m[133]&m[281]&m[823]))):InitCond[1286];
    m[568] = run?((((~m[134]&~m[297]&~m[824])|(m[134]&m[297]&~m[824]))&BiasedRNG[791])|(((m[134]&~m[297]&~m[824])|(~m[134]&m[297]&m[824]))&~BiasedRNG[791])|((~m[134]&~m[297]&m[824])|(m[134]&~m[297]&m[824])|(m[134]&m[297]&m[824]))):InitCond[1287];
    m[569] = run?((((~m[134]&~m[313]&~m[825])|(m[134]&m[313]&~m[825]))&BiasedRNG[792])|(((m[134]&~m[313]&~m[825])|(~m[134]&m[313]&m[825]))&~BiasedRNG[792])|((~m[134]&~m[313]&m[825])|(m[134]&~m[313]&m[825])|(m[134]&m[313]&m[825]))):InitCond[1288];
    m[570] = run?((((~m[134]&~m[329]&~m[826])|(m[134]&m[329]&~m[826]))&BiasedRNG[793])|(((m[134]&~m[329]&~m[826])|(~m[134]&m[329]&m[826]))&~BiasedRNG[793])|((~m[134]&~m[329]&m[826])|(m[134]&~m[329]&m[826])|(m[134]&m[329]&m[826]))):InitCond[1289];
    m[571] = run?((((~m[134]&~m[345]&~m[827])|(m[134]&m[345]&~m[827]))&BiasedRNG[794])|(((m[134]&~m[345]&~m[827])|(~m[134]&m[345]&m[827]))&~BiasedRNG[794])|((~m[134]&~m[345]&m[827])|(m[134]&~m[345]&m[827])|(m[134]&m[345]&m[827]))):InitCond[1290];
    m[572] = run?((((~m[135]&~m[361]&~m[828])|(m[135]&m[361]&~m[828]))&BiasedRNG[795])|(((m[135]&~m[361]&~m[828])|(~m[135]&m[361]&m[828]))&~BiasedRNG[795])|((~m[135]&~m[361]&m[828])|(m[135]&~m[361]&m[828])|(m[135]&m[361]&m[828]))):InitCond[1291];
    m[573] = run?((((~m[135]&~m[377]&~m[829])|(m[135]&m[377]&~m[829]))&BiasedRNG[796])|(((m[135]&~m[377]&~m[829])|(~m[135]&m[377]&m[829]))&~BiasedRNG[796])|((~m[135]&~m[377]&m[829])|(m[135]&~m[377]&m[829])|(m[135]&m[377]&m[829]))):InitCond[1292];
    m[574] = run?((((~m[135]&~m[393]&~m[830])|(m[135]&m[393]&~m[830]))&BiasedRNG[797])|(((m[135]&~m[393]&~m[830])|(~m[135]&m[393]&m[830]))&~BiasedRNG[797])|((~m[135]&~m[393]&m[830])|(m[135]&~m[393]&m[830])|(m[135]&m[393]&m[830]))):InitCond[1293];
    m[575] = run?((((~m[135]&~m[409]&~m[831])|(m[135]&m[409]&~m[831]))&BiasedRNG[798])|(((m[135]&~m[409]&~m[831])|(~m[135]&m[409]&m[831]))&~BiasedRNG[798])|((~m[135]&~m[409]&m[831])|(m[135]&~m[409]&m[831])|(m[135]&m[409]&m[831]))):InitCond[1294];
    m[576] = run?((((~m[136]&~m[170]&~m[832])|(m[136]&m[170]&~m[832]))&BiasedRNG[799])|(((m[136]&~m[170]&~m[832])|(~m[136]&m[170]&m[832]))&~BiasedRNG[799])|((~m[136]&~m[170]&m[832])|(m[136]&~m[170]&m[832])|(m[136]&m[170]&m[832]))):InitCond[1295];
    m[577] = run?((((~m[136]&~m[186]&~m[833])|(m[136]&m[186]&~m[833]))&BiasedRNG[800])|(((m[136]&~m[186]&~m[833])|(~m[136]&m[186]&m[833]))&~BiasedRNG[800])|((~m[136]&~m[186]&m[833])|(m[136]&~m[186]&m[833])|(m[136]&m[186]&m[833]))):InitCond[1296];
    m[578] = run?((((~m[136]&~m[202]&~m[834])|(m[136]&m[202]&~m[834]))&BiasedRNG[801])|(((m[136]&~m[202]&~m[834])|(~m[136]&m[202]&m[834]))&~BiasedRNG[801])|((~m[136]&~m[202]&m[834])|(m[136]&~m[202]&m[834])|(m[136]&m[202]&m[834]))):InitCond[1297];
    m[579] = run?((((~m[136]&~m[218]&~m[835])|(m[136]&m[218]&~m[835]))&BiasedRNG[802])|(((m[136]&~m[218]&~m[835])|(~m[136]&m[218]&m[835]))&~BiasedRNG[802])|((~m[136]&~m[218]&m[835])|(m[136]&~m[218]&m[835])|(m[136]&m[218]&m[835]))):InitCond[1298];
    m[580] = run?((((~m[137]&~m[234]&~m[836])|(m[137]&m[234]&~m[836]))&BiasedRNG[803])|(((m[137]&~m[234]&~m[836])|(~m[137]&m[234]&m[836]))&~BiasedRNG[803])|((~m[137]&~m[234]&m[836])|(m[137]&~m[234]&m[836])|(m[137]&m[234]&m[836]))):InitCond[1299];
    m[581] = run?((((~m[137]&~m[250]&~m[837])|(m[137]&m[250]&~m[837]))&BiasedRNG[804])|(((m[137]&~m[250]&~m[837])|(~m[137]&m[250]&m[837]))&~BiasedRNG[804])|((~m[137]&~m[250]&m[837])|(m[137]&~m[250]&m[837])|(m[137]&m[250]&m[837]))):InitCond[1300];
    m[582] = run?((((~m[137]&~m[266]&~m[838])|(m[137]&m[266]&~m[838]))&BiasedRNG[805])|(((m[137]&~m[266]&~m[838])|(~m[137]&m[266]&m[838]))&~BiasedRNG[805])|((~m[137]&~m[266]&m[838])|(m[137]&~m[266]&m[838])|(m[137]&m[266]&m[838]))):InitCond[1301];
    m[583] = run?((((~m[137]&~m[282]&~m[839])|(m[137]&m[282]&~m[839]))&BiasedRNG[806])|(((m[137]&~m[282]&~m[839])|(~m[137]&m[282]&m[839]))&~BiasedRNG[806])|((~m[137]&~m[282]&m[839])|(m[137]&~m[282]&m[839])|(m[137]&m[282]&m[839]))):InitCond[1302];
    m[584] = run?((((~m[138]&~m[298]&~m[840])|(m[138]&m[298]&~m[840]))&BiasedRNG[807])|(((m[138]&~m[298]&~m[840])|(~m[138]&m[298]&m[840]))&~BiasedRNG[807])|((~m[138]&~m[298]&m[840])|(m[138]&~m[298]&m[840])|(m[138]&m[298]&m[840]))):InitCond[1303];
    m[585] = run?((((~m[138]&~m[314]&~m[841])|(m[138]&m[314]&~m[841]))&BiasedRNG[808])|(((m[138]&~m[314]&~m[841])|(~m[138]&m[314]&m[841]))&~BiasedRNG[808])|((~m[138]&~m[314]&m[841])|(m[138]&~m[314]&m[841])|(m[138]&m[314]&m[841]))):InitCond[1304];
    m[586] = run?((((~m[138]&~m[330]&~m[842])|(m[138]&m[330]&~m[842]))&BiasedRNG[809])|(((m[138]&~m[330]&~m[842])|(~m[138]&m[330]&m[842]))&~BiasedRNG[809])|((~m[138]&~m[330]&m[842])|(m[138]&~m[330]&m[842])|(m[138]&m[330]&m[842]))):InitCond[1305];
    m[587] = run?((((~m[138]&~m[346]&~m[843])|(m[138]&m[346]&~m[843]))&BiasedRNG[810])|(((m[138]&~m[346]&~m[843])|(~m[138]&m[346]&m[843]))&~BiasedRNG[810])|((~m[138]&~m[346]&m[843])|(m[138]&~m[346]&m[843])|(m[138]&m[346]&m[843]))):InitCond[1306];
    m[588] = run?((((~m[139]&~m[362]&~m[844])|(m[139]&m[362]&~m[844]))&BiasedRNG[811])|(((m[139]&~m[362]&~m[844])|(~m[139]&m[362]&m[844]))&~BiasedRNG[811])|((~m[139]&~m[362]&m[844])|(m[139]&~m[362]&m[844])|(m[139]&m[362]&m[844]))):InitCond[1307];
    m[589] = run?((((~m[139]&~m[378]&~m[845])|(m[139]&m[378]&~m[845]))&BiasedRNG[812])|(((m[139]&~m[378]&~m[845])|(~m[139]&m[378]&m[845]))&~BiasedRNG[812])|((~m[139]&~m[378]&m[845])|(m[139]&~m[378]&m[845])|(m[139]&m[378]&m[845]))):InitCond[1308];
    m[590] = run?((((~m[139]&~m[394]&~m[846])|(m[139]&m[394]&~m[846]))&BiasedRNG[813])|(((m[139]&~m[394]&~m[846])|(~m[139]&m[394]&m[846]))&~BiasedRNG[813])|((~m[139]&~m[394]&m[846])|(m[139]&~m[394]&m[846])|(m[139]&m[394]&m[846]))):InitCond[1309];
    m[591] = run?((((~m[139]&~m[410]&~m[847])|(m[139]&m[410]&~m[847]))&BiasedRNG[814])|(((m[139]&~m[410]&~m[847])|(~m[139]&m[410]&m[847]))&~BiasedRNG[814])|((~m[139]&~m[410]&m[847])|(m[139]&~m[410]&m[847])|(m[139]&m[410]&m[847]))):InitCond[1310];
    m[592] = run?((((~m[140]&~m[171]&~m[848])|(m[140]&m[171]&~m[848]))&BiasedRNG[815])|(((m[140]&~m[171]&~m[848])|(~m[140]&m[171]&m[848]))&~BiasedRNG[815])|((~m[140]&~m[171]&m[848])|(m[140]&~m[171]&m[848])|(m[140]&m[171]&m[848]))):InitCond[1311];
    m[593] = run?((((~m[140]&~m[187]&~m[849])|(m[140]&m[187]&~m[849]))&BiasedRNG[816])|(((m[140]&~m[187]&~m[849])|(~m[140]&m[187]&m[849]))&~BiasedRNG[816])|((~m[140]&~m[187]&m[849])|(m[140]&~m[187]&m[849])|(m[140]&m[187]&m[849]))):InitCond[1312];
    m[594] = run?((((~m[140]&~m[203]&~m[850])|(m[140]&m[203]&~m[850]))&BiasedRNG[817])|(((m[140]&~m[203]&~m[850])|(~m[140]&m[203]&m[850]))&~BiasedRNG[817])|((~m[140]&~m[203]&m[850])|(m[140]&~m[203]&m[850])|(m[140]&m[203]&m[850]))):InitCond[1313];
    m[595] = run?((((~m[140]&~m[219]&~m[851])|(m[140]&m[219]&~m[851]))&BiasedRNG[818])|(((m[140]&~m[219]&~m[851])|(~m[140]&m[219]&m[851]))&~BiasedRNG[818])|((~m[140]&~m[219]&m[851])|(m[140]&~m[219]&m[851])|(m[140]&m[219]&m[851]))):InitCond[1314];
    m[596] = run?((((~m[141]&~m[235]&~m[852])|(m[141]&m[235]&~m[852]))&BiasedRNG[819])|(((m[141]&~m[235]&~m[852])|(~m[141]&m[235]&m[852]))&~BiasedRNG[819])|((~m[141]&~m[235]&m[852])|(m[141]&~m[235]&m[852])|(m[141]&m[235]&m[852]))):InitCond[1315];
    m[597] = run?((((~m[141]&~m[251]&~m[853])|(m[141]&m[251]&~m[853]))&BiasedRNG[820])|(((m[141]&~m[251]&~m[853])|(~m[141]&m[251]&m[853]))&~BiasedRNG[820])|((~m[141]&~m[251]&m[853])|(m[141]&~m[251]&m[853])|(m[141]&m[251]&m[853]))):InitCond[1316];
    m[598] = run?((((~m[141]&~m[267]&~m[854])|(m[141]&m[267]&~m[854]))&BiasedRNG[821])|(((m[141]&~m[267]&~m[854])|(~m[141]&m[267]&m[854]))&~BiasedRNG[821])|((~m[141]&~m[267]&m[854])|(m[141]&~m[267]&m[854])|(m[141]&m[267]&m[854]))):InitCond[1317];
    m[599] = run?((((~m[141]&~m[283]&~m[855])|(m[141]&m[283]&~m[855]))&BiasedRNG[822])|(((m[141]&~m[283]&~m[855])|(~m[141]&m[283]&m[855]))&~BiasedRNG[822])|((~m[141]&~m[283]&m[855])|(m[141]&~m[283]&m[855])|(m[141]&m[283]&m[855]))):InitCond[1318];
    m[600] = run?((((~m[142]&~m[299]&~m[856])|(m[142]&m[299]&~m[856]))&BiasedRNG[823])|(((m[142]&~m[299]&~m[856])|(~m[142]&m[299]&m[856]))&~BiasedRNG[823])|((~m[142]&~m[299]&m[856])|(m[142]&~m[299]&m[856])|(m[142]&m[299]&m[856]))):InitCond[1319];
    m[601] = run?((((~m[142]&~m[315]&~m[857])|(m[142]&m[315]&~m[857]))&BiasedRNG[824])|(((m[142]&~m[315]&~m[857])|(~m[142]&m[315]&m[857]))&~BiasedRNG[824])|((~m[142]&~m[315]&m[857])|(m[142]&~m[315]&m[857])|(m[142]&m[315]&m[857]))):InitCond[1320];
    m[602] = run?((((~m[142]&~m[331]&~m[858])|(m[142]&m[331]&~m[858]))&BiasedRNG[825])|(((m[142]&~m[331]&~m[858])|(~m[142]&m[331]&m[858]))&~BiasedRNG[825])|((~m[142]&~m[331]&m[858])|(m[142]&~m[331]&m[858])|(m[142]&m[331]&m[858]))):InitCond[1321];
    m[603] = run?((((~m[142]&~m[347]&~m[859])|(m[142]&m[347]&~m[859]))&BiasedRNG[826])|(((m[142]&~m[347]&~m[859])|(~m[142]&m[347]&m[859]))&~BiasedRNG[826])|((~m[142]&~m[347]&m[859])|(m[142]&~m[347]&m[859])|(m[142]&m[347]&m[859]))):InitCond[1322];
    m[604] = run?((((~m[143]&~m[363]&~m[860])|(m[143]&m[363]&~m[860]))&BiasedRNG[827])|(((m[143]&~m[363]&~m[860])|(~m[143]&m[363]&m[860]))&~BiasedRNG[827])|((~m[143]&~m[363]&m[860])|(m[143]&~m[363]&m[860])|(m[143]&m[363]&m[860]))):InitCond[1323];
    m[605] = run?((((~m[143]&~m[379]&~m[861])|(m[143]&m[379]&~m[861]))&BiasedRNG[828])|(((m[143]&~m[379]&~m[861])|(~m[143]&m[379]&m[861]))&~BiasedRNG[828])|((~m[143]&~m[379]&m[861])|(m[143]&~m[379]&m[861])|(m[143]&m[379]&m[861]))):InitCond[1324];
    m[606] = run?((((~m[143]&~m[395]&~m[862])|(m[143]&m[395]&~m[862]))&BiasedRNG[829])|(((m[143]&~m[395]&~m[862])|(~m[143]&m[395]&m[862]))&~BiasedRNG[829])|((~m[143]&~m[395]&m[862])|(m[143]&~m[395]&m[862])|(m[143]&m[395]&m[862]))):InitCond[1325];
    m[607] = run?((((~m[143]&~m[411]&~m[863])|(m[143]&m[411]&~m[863]))&BiasedRNG[830])|(((m[143]&~m[411]&~m[863])|(~m[143]&m[411]&m[863]))&~BiasedRNG[830])|((~m[143]&~m[411]&m[863])|(m[143]&~m[411]&m[863])|(m[143]&m[411]&m[863]))):InitCond[1326];
    m[608] = run?((((~m[144]&~m[172]&~m[864])|(m[144]&m[172]&~m[864]))&BiasedRNG[831])|(((m[144]&~m[172]&~m[864])|(~m[144]&m[172]&m[864]))&~BiasedRNG[831])|((~m[144]&~m[172]&m[864])|(m[144]&~m[172]&m[864])|(m[144]&m[172]&m[864]))):InitCond[1327];
    m[609] = run?((((~m[144]&~m[188]&~m[865])|(m[144]&m[188]&~m[865]))&BiasedRNG[832])|(((m[144]&~m[188]&~m[865])|(~m[144]&m[188]&m[865]))&~BiasedRNG[832])|((~m[144]&~m[188]&m[865])|(m[144]&~m[188]&m[865])|(m[144]&m[188]&m[865]))):InitCond[1328];
    m[610] = run?((((~m[144]&~m[204]&~m[866])|(m[144]&m[204]&~m[866]))&BiasedRNG[833])|(((m[144]&~m[204]&~m[866])|(~m[144]&m[204]&m[866]))&~BiasedRNG[833])|((~m[144]&~m[204]&m[866])|(m[144]&~m[204]&m[866])|(m[144]&m[204]&m[866]))):InitCond[1329];
    m[611] = run?((((~m[144]&~m[220]&~m[867])|(m[144]&m[220]&~m[867]))&BiasedRNG[834])|(((m[144]&~m[220]&~m[867])|(~m[144]&m[220]&m[867]))&~BiasedRNG[834])|((~m[144]&~m[220]&m[867])|(m[144]&~m[220]&m[867])|(m[144]&m[220]&m[867]))):InitCond[1330];
    m[612] = run?((((~m[145]&~m[236]&~m[868])|(m[145]&m[236]&~m[868]))&BiasedRNG[835])|(((m[145]&~m[236]&~m[868])|(~m[145]&m[236]&m[868]))&~BiasedRNG[835])|((~m[145]&~m[236]&m[868])|(m[145]&~m[236]&m[868])|(m[145]&m[236]&m[868]))):InitCond[1331];
    m[613] = run?((((~m[145]&~m[252]&~m[869])|(m[145]&m[252]&~m[869]))&BiasedRNG[836])|(((m[145]&~m[252]&~m[869])|(~m[145]&m[252]&m[869]))&~BiasedRNG[836])|((~m[145]&~m[252]&m[869])|(m[145]&~m[252]&m[869])|(m[145]&m[252]&m[869]))):InitCond[1332];
    m[614] = run?((((~m[145]&~m[268]&~m[870])|(m[145]&m[268]&~m[870]))&BiasedRNG[837])|(((m[145]&~m[268]&~m[870])|(~m[145]&m[268]&m[870]))&~BiasedRNG[837])|((~m[145]&~m[268]&m[870])|(m[145]&~m[268]&m[870])|(m[145]&m[268]&m[870]))):InitCond[1333];
    m[615] = run?((((~m[145]&~m[284]&~m[871])|(m[145]&m[284]&~m[871]))&BiasedRNG[838])|(((m[145]&~m[284]&~m[871])|(~m[145]&m[284]&m[871]))&~BiasedRNG[838])|((~m[145]&~m[284]&m[871])|(m[145]&~m[284]&m[871])|(m[145]&m[284]&m[871]))):InitCond[1334];
    m[616] = run?((((~m[146]&~m[300]&~m[872])|(m[146]&m[300]&~m[872]))&BiasedRNG[839])|(((m[146]&~m[300]&~m[872])|(~m[146]&m[300]&m[872]))&~BiasedRNG[839])|((~m[146]&~m[300]&m[872])|(m[146]&~m[300]&m[872])|(m[146]&m[300]&m[872]))):InitCond[1335];
    m[617] = run?((((~m[146]&~m[316]&~m[873])|(m[146]&m[316]&~m[873]))&BiasedRNG[840])|(((m[146]&~m[316]&~m[873])|(~m[146]&m[316]&m[873]))&~BiasedRNG[840])|((~m[146]&~m[316]&m[873])|(m[146]&~m[316]&m[873])|(m[146]&m[316]&m[873]))):InitCond[1336];
    m[618] = run?((((~m[146]&~m[332]&~m[874])|(m[146]&m[332]&~m[874]))&BiasedRNG[841])|(((m[146]&~m[332]&~m[874])|(~m[146]&m[332]&m[874]))&~BiasedRNG[841])|((~m[146]&~m[332]&m[874])|(m[146]&~m[332]&m[874])|(m[146]&m[332]&m[874]))):InitCond[1337];
    m[619] = run?((((~m[146]&~m[348]&~m[875])|(m[146]&m[348]&~m[875]))&BiasedRNG[842])|(((m[146]&~m[348]&~m[875])|(~m[146]&m[348]&m[875]))&~BiasedRNG[842])|((~m[146]&~m[348]&m[875])|(m[146]&~m[348]&m[875])|(m[146]&m[348]&m[875]))):InitCond[1338];
    m[620] = run?((((~m[147]&~m[364]&~m[876])|(m[147]&m[364]&~m[876]))&BiasedRNG[843])|(((m[147]&~m[364]&~m[876])|(~m[147]&m[364]&m[876]))&~BiasedRNG[843])|((~m[147]&~m[364]&m[876])|(m[147]&~m[364]&m[876])|(m[147]&m[364]&m[876]))):InitCond[1339];
    m[621] = run?((((~m[147]&~m[380]&~m[877])|(m[147]&m[380]&~m[877]))&BiasedRNG[844])|(((m[147]&~m[380]&~m[877])|(~m[147]&m[380]&m[877]))&~BiasedRNG[844])|((~m[147]&~m[380]&m[877])|(m[147]&~m[380]&m[877])|(m[147]&m[380]&m[877]))):InitCond[1340];
    m[622] = run?((((~m[147]&~m[396]&~m[878])|(m[147]&m[396]&~m[878]))&BiasedRNG[845])|(((m[147]&~m[396]&~m[878])|(~m[147]&m[396]&m[878]))&~BiasedRNG[845])|((~m[147]&~m[396]&m[878])|(m[147]&~m[396]&m[878])|(m[147]&m[396]&m[878]))):InitCond[1341];
    m[623] = run?((((~m[147]&~m[412]&~m[879])|(m[147]&m[412]&~m[879]))&BiasedRNG[846])|(((m[147]&~m[412]&~m[879])|(~m[147]&m[412]&m[879]))&~BiasedRNG[846])|((~m[147]&~m[412]&m[879])|(m[147]&~m[412]&m[879])|(m[147]&m[412]&m[879]))):InitCond[1342];
    m[624] = run?((((~m[148]&~m[173]&~m[880])|(m[148]&m[173]&~m[880]))&BiasedRNG[847])|(((m[148]&~m[173]&~m[880])|(~m[148]&m[173]&m[880]))&~BiasedRNG[847])|((~m[148]&~m[173]&m[880])|(m[148]&~m[173]&m[880])|(m[148]&m[173]&m[880]))):InitCond[1343];
    m[625] = run?((((~m[148]&~m[189]&~m[881])|(m[148]&m[189]&~m[881]))&BiasedRNG[848])|(((m[148]&~m[189]&~m[881])|(~m[148]&m[189]&m[881]))&~BiasedRNG[848])|((~m[148]&~m[189]&m[881])|(m[148]&~m[189]&m[881])|(m[148]&m[189]&m[881]))):InitCond[1344];
    m[626] = run?((((~m[148]&~m[205]&~m[882])|(m[148]&m[205]&~m[882]))&BiasedRNG[849])|(((m[148]&~m[205]&~m[882])|(~m[148]&m[205]&m[882]))&~BiasedRNG[849])|((~m[148]&~m[205]&m[882])|(m[148]&~m[205]&m[882])|(m[148]&m[205]&m[882]))):InitCond[1345];
    m[627] = run?((((~m[148]&~m[221]&~m[883])|(m[148]&m[221]&~m[883]))&BiasedRNG[850])|(((m[148]&~m[221]&~m[883])|(~m[148]&m[221]&m[883]))&~BiasedRNG[850])|((~m[148]&~m[221]&m[883])|(m[148]&~m[221]&m[883])|(m[148]&m[221]&m[883]))):InitCond[1346];
    m[628] = run?((((~m[149]&~m[237]&~m[884])|(m[149]&m[237]&~m[884]))&BiasedRNG[851])|(((m[149]&~m[237]&~m[884])|(~m[149]&m[237]&m[884]))&~BiasedRNG[851])|((~m[149]&~m[237]&m[884])|(m[149]&~m[237]&m[884])|(m[149]&m[237]&m[884]))):InitCond[1347];
    m[629] = run?((((~m[149]&~m[253]&~m[885])|(m[149]&m[253]&~m[885]))&BiasedRNG[852])|(((m[149]&~m[253]&~m[885])|(~m[149]&m[253]&m[885]))&~BiasedRNG[852])|((~m[149]&~m[253]&m[885])|(m[149]&~m[253]&m[885])|(m[149]&m[253]&m[885]))):InitCond[1348];
    m[630] = run?((((~m[149]&~m[269]&~m[886])|(m[149]&m[269]&~m[886]))&BiasedRNG[853])|(((m[149]&~m[269]&~m[886])|(~m[149]&m[269]&m[886]))&~BiasedRNG[853])|((~m[149]&~m[269]&m[886])|(m[149]&~m[269]&m[886])|(m[149]&m[269]&m[886]))):InitCond[1349];
    m[631] = run?((((~m[149]&~m[285]&~m[887])|(m[149]&m[285]&~m[887]))&BiasedRNG[854])|(((m[149]&~m[285]&~m[887])|(~m[149]&m[285]&m[887]))&~BiasedRNG[854])|((~m[149]&~m[285]&m[887])|(m[149]&~m[285]&m[887])|(m[149]&m[285]&m[887]))):InitCond[1350];
    m[632] = run?((((~m[150]&~m[301]&~m[888])|(m[150]&m[301]&~m[888]))&BiasedRNG[855])|(((m[150]&~m[301]&~m[888])|(~m[150]&m[301]&m[888]))&~BiasedRNG[855])|((~m[150]&~m[301]&m[888])|(m[150]&~m[301]&m[888])|(m[150]&m[301]&m[888]))):InitCond[1351];
    m[633] = run?((((~m[150]&~m[317]&~m[889])|(m[150]&m[317]&~m[889]))&BiasedRNG[856])|(((m[150]&~m[317]&~m[889])|(~m[150]&m[317]&m[889]))&~BiasedRNG[856])|((~m[150]&~m[317]&m[889])|(m[150]&~m[317]&m[889])|(m[150]&m[317]&m[889]))):InitCond[1352];
    m[634] = run?((((~m[150]&~m[333]&~m[890])|(m[150]&m[333]&~m[890]))&BiasedRNG[857])|(((m[150]&~m[333]&~m[890])|(~m[150]&m[333]&m[890]))&~BiasedRNG[857])|((~m[150]&~m[333]&m[890])|(m[150]&~m[333]&m[890])|(m[150]&m[333]&m[890]))):InitCond[1353];
    m[635] = run?((((~m[150]&~m[349]&~m[891])|(m[150]&m[349]&~m[891]))&BiasedRNG[858])|(((m[150]&~m[349]&~m[891])|(~m[150]&m[349]&m[891]))&~BiasedRNG[858])|((~m[150]&~m[349]&m[891])|(m[150]&~m[349]&m[891])|(m[150]&m[349]&m[891]))):InitCond[1354];
    m[636] = run?((((~m[151]&~m[365]&~m[892])|(m[151]&m[365]&~m[892]))&BiasedRNG[859])|(((m[151]&~m[365]&~m[892])|(~m[151]&m[365]&m[892]))&~BiasedRNG[859])|((~m[151]&~m[365]&m[892])|(m[151]&~m[365]&m[892])|(m[151]&m[365]&m[892]))):InitCond[1355];
    m[637] = run?((((~m[151]&~m[381]&~m[893])|(m[151]&m[381]&~m[893]))&BiasedRNG[860])|(((m[151]&~m[381]&~m[893])|(~m[151]&m[381]&m[893]))&~BiasedRNG[860])|((~m[151]&~m[381]&m[893])|(m[151]&~m[381]&m[893])|(m[151]&m[381]&m[893]))):InitCond[1356];
    m[638] = run?((((~m[151]&~m[397]&~m[894])|(m[151]&m[397]&~m[894]))&BiasedRNG[861])|(((m[151]&~m[397]&~m[894])|(~m[151]&m[397]&m[894]))&~BiasedRNG[861])|((~m[151]&~m[397]&m[894])|(m[151]&~m[397]&m[894])|(m[151]&m[397]&m[894]))):InitCond[1357];
    m[639] = run?((((~m[151]&~m[413]&~m[895])|(m[151]&m[413]&~m[895]))&BiasedRNG[862])|(((m[151]&~m[413]&~m[895])|(~m[151]&m[413]&m[895]))&~BiasedRNG[862])|((~m[151]&~m[413]&m[895])|(m[151]&~m[413]&m[895])|(m[151]&m[413]&m[895]))):InitCond[1358];
    m[640] = run?((((~m[152]&~m[174]&~m[896])|(m[152]&m[174]&~m[896]))&BiasedRNG[863])|(((m[152]&~m[174]&~m[896])|(~m[152]&m[174]&m[896]))&~BiasedRNG[863])|((~m[152]&~m[174]&m[896])|(m[152]&~m[174]&m[896])|(m[152]&m[174]&m[896]))):InitCond[1359];
    m[641] = run?((((~m[152]&~m[190]&~m[897])|(m[152]&m[190]&~m[897]))&BiasedRNG[864])|(((m[152]&~m[190]&~m[897])|(~m[152]&m[190]&m[897]))&~BiasedRNG[864])|((~m[152]&~m[190]&m[897])|(m[152]&~m[190]&m[897])|(m[152]&m[190]&m[897]))):InitCond[1360];
    m[642] = run?((((~m[152]&~m[206]&~m[898])|(m[152]&m[206]&~m[898]))&BiasedRNG[865])|(((m[152]&~m[206]&~m[898])|(~m[152]&m[206]&m[898]))&~BiasedRNG[865])|((~m[152]&~m[206]&m[898])|(m[152]&~m[206]&m[898])|(m[152]&m[206]&m[898]))):InitCond[1361];
    m[643] = run?((((~m[152]&~m[222]&~m[899])|(m[152]&m[222]&~m[899]))&BiasedRNG[866])|(((m[152]&~m[222]&~m[899])|(~m[152]&m[222]&m[899]))&~BiasedRNG[866])|((~m[152]&~m[222]&m[899])|(m[152]&~m[222]&m[899])|(m[152]&m[222]&m[899]))):InitCond[1362];
    m[644] = run?((((~m[153]&~m[238]&~m[900])|(m[153]&m[238]&~m[900]))&BiasedRNG[867])|(((m[153]&~m[238]&~m[900])|(~m[153]&m[238]&m[900]))&~BiasedRNG[867])|((~m[153]&~m[238]&m[900])|(m[153]&~m[238]&m[900])|(m[153]&m[238]&m[900]))):InitCond[1363];
    m[645] = run?((((~m[153]&~m[254]&~m[901])|(m[153]&m[254]&~m[901]))&BiasedRNG[868])|(((m[153]&~m[254]&~m[901])|(~m[153]&m[254]&m[901]))&~BiasedRNG[868])|((~m[153]&~m[254]&m[901])|(m[153]&~m[254]&m[901])|(m[153]&m[254]&m[901]))):InitCond[1364];
    m[646] = run?((((~m[153]&~m[270]&~m[902])|(m[153]&m[270]&~m[902]))&BiasedRNG[869])|(((m[153]&~m[270]&~m[902])|(~m[153]&m[270]&m[902]))&~BiasedRNG[869])|((~m[153]&~m[270]&m[902])|(m[153]&~m[270]&m[902])|(m[153]&m[270]&m[902]))):InitCond[1365];
    m[647] = run?((((~m[153]&~m[286]&~m[903])|(m[153]&m[286]&~m[903]))&BiasedRNG[870])|(((m[153]&~m[286]&~m[903])|(~m[153]&m[286]&m[903]))&~BiasedRNG[870])|((~m[153]&~m[286]&m[903])|(m[153]&~m[286]&m[903])|(m[153]&m[286]&m[903]))):InitCond[1366];
    m[648] = run?((((~m[154]&~m[302]&~m[904])|(m[154]&m[302]&~m[904]))&BiasedRNG[871])|(((m[154]&~m[302]&~m[904])|(~m[154]&m[302]&m[904]))&~BiasedRNG[871])|((~m[154]&~m[302]&m[904])|(m[154]&~m[302]&m[904])|(m[154]&m[302]&m[904]))):InitCond[1367];
    m[649] = run?((((~m[154]&~m[318]&~m[905])|(m[154]&m[318]&~m[905]))&BiasedRNG[872])|(((m[154]&~m[318]&~m[905])|(~m[154]&m[318]&m[905]))&~BiasedRNG[872])|((~m[154]&~m[318]&m[905])|(m[154]&~m[318]&m[905])|(m[154]&m[318]&m[905]))):InitCond[1368];
    m[650] = run?((((~m[154]&~m[334]&~m[906])|(m[154]&m[334]&~m[906]))&BiasedRNG[873])|(((m[154]&~m[334]&~m[906])|(~m[154]&m[334]&m[906]))&~BiasedRNG[873])|((~m[154]&~m[334]&m[906])|(m[154]&~m[334]&m[906])|(m[154]&m[334]&m[906]))):InitCond[1369];
    m[651] = run?((((~m[154]&~m[350]&~m[907])|(m[154]&m[350]&~m[907]))&BiasedRNG[874])|(((m[154]&~m[350]&~m[907])|(~m[154]&m[350]&m[907]))&~BiasedRNG[874])|((~m[154]&~m[350]&m[907])|(m[154]&~m[350]&m[907])|(m[154]&m[350]&m[907]))):InitCond[1370];
    m[652] = run?((((~m[155]&~m[366]&~m[908])|(m[155]&m[366]&~m[908]))&BiasedRNG[875])|(((m[155]&~m[366]&~m[908])|(~m[155]&m[366]&m[908]))&~BiasedRNG[875])|((~m[155]&~m[366]&m[908])|(m[155]&~m[366]&m[908])|(m[155]&m[366]&m[908]))):InitCond[1371];
    m[653] = run?((((~m[155]&~m[382]&~m[909])|(m[155]&m[382]&~m[909]))&BiasedRNG[876])|(((m[155]&~m[382]&~m[909])|(~m[155]&m[382]&m[909]))&~BiasedRNG[876])|((~m[155]&~m[382]&m[909])|(m[155]&~m[382]&m[909])|(m[155]&m[382]&m[909]))):InitCond[1372];
    m[654] = run?((((~m[155]&~m[398]&~m[910])|(m[155]&m[398]&~m[910]))&BiasedRNG[877])|(((m[155]&~m[398]&~m[910])|(~m[155]&m[398]&m[910]))&~BiasedRNG[877])|((~m[155]&~m[398]&m[910])|(m[155]&~m[398]&m[910])|(m[155]&m[398]&m[910]))):InitCond[1373];
    m[655] = run?((((~m[155]&~m[414]&~m[911])|(m[155]&m[414]&~m[911]))&BiasedRNG[878])|(((m[155]&~m[414]&~m[911])|(~m[155]&m[414]&m[911]))&~BiasedRNG[878])|((~m[155]&~m[414]&m[911])|(m[155]&~m[414]&m[911])|(m[155]&m[414]&m[911]))):InitCond[1374];
    m[656] = run?((((~m[156]&~m[175]&~m[912])|(m[156]&m[175]&~m[912]))&BiasedRNG[879])|(((m[156]&~m[175]&~m[912])|(~m[156]&m[175]&m[912]))&~BiasedRNG[879])|((~m[156]&~m[175]&m[912])|(m[156]&~m[175]&m[912])|(m[156]&m[175]&m[912]))):InitCond[1375];
    m[657] = run?((((~m[156]&~m[191]&~m[913])|(m[156]&m[191]&~m[913]))&BiasedRNG[880])|(((m[156]&~m[191]&~m[913])|(~m[156]&m[191]&m[913]))&~BiasedRNG[880])|((~m[156]&~m[191]&m[913])|(m[156]&~m[191]&m[913])|(m[156]&m[191]&m[913]))):InitCond[1376];
    m[658] = run?((((~m[156]&~m[207]&~m[914])|(m[156]&m[207]&~m[914]))&BiasedRNG[881])|(((m[156]&~m[207]&~m[914])|(~m[156]&m[207]&m[914]))&~BiasedRNG[881])|((~m[156]&~m[207]&m[914])|(m[156]&~m[207]&m[914])|(m[156]&m[207]&m[914]))):InitCond[1377];
    m[659] = run?((((~m[156]&~m[223]&~m[915])|(m[156]&m[223]&~m[915]))&BiasedRNG[882])|(((m[156]&~m[223]&~m[915])|(~m[156]&m[223]&m[915]))&~BiasedRNG[882])|((~m[156]&~m[223]&m[915])|(m[156]&~m[223]&m[915])|(m[156]&m[223]&m[915]))):InitCond[1378];
    m[660] = run?((((~m[157]&~m[239]&~m[916])|(m[157]&m[239]&~m[916]))&BiasedRNG[883])|(((m[157]&~m[239]&~m[916])|(~m[157]&m[239]&m[916]))&~BiasedRNG[883])|((~m[157]&~m[239]&m[916])|(m[157]&~m[239]&m[916])|(m[157]&m[239]&m[916]))):InitCond[1379];
    m[661] = run?((((~m[157]&~m[255]&~m[917])|(m[157]&m[255]&~m[917]))&BiasedRNG[884])|(((m[157]&~m[255]&~m[917])|(~m[157]&m[255]&m[917]))&~BiasedRNG[884])|((~m[157]&~m[255]&m[917])|(m[157]&~m[255]&m[917])|(m[157]&m[255]&m[917]))):InitCond[1380];
    m[662] = run?((((~m[157]&~m[271]&~m[918])|(m[157]&m[271]&~m[918]))&BiasedRNG[885])|(((m[157]&~m[271]&~m[918])|(~m[157]&m[271]&m[918]))&~BiasedRNG[885])|((~m[157]&~m[271]&m[918])|(m[157]&~m[271]&m[918])|(m[157]&m[271]&m[918]))):InitCond[1381];
    m[663] = run?((((~m[157]&~m[287]&~m[919])|(m[157]&m[287]&~m[919]))&BiasedRNG[886])|(((m[157]&~m[287]&~m[919])|(~m[157]&m[287]&m[919]))&~BiasedRNG[886])|((~m[157]&~m[287]&m[919])|(m[157]&~m[287]&m[919])|(m[157]&m[287]&m[919]))):InitCond[1382];
    m[664] = run?((((~m[158]&~m[303]&~m[920])|(m[158]&m[303]&~m[920]))&BiasedRNG[887])|(((m[158]&~m[303]&~m[920])|(~m[158]&m[303]&m[920]))&~BiasedRNG[887])|((~m[158]&~m[303]&m[920])|(m[158]&~m[303]&m[920])|(m[158]&m[303]&m[920]))):InitCond[1383];
    m[665] = run?((((~m[158]&~m[319]&~m[921])|(m[158]&m[319]&~m[921]))&BiasedRNG[888])|(((m[158]&~m[319]&~m[921])|(~m[158]&m[319]&m[921]))&~BiasedRNG[888])|((~m[158]&~m[319]&m[921])|(m[158]&~m[319]&m[921])|(m[158]&m[319]&m[921]))):InitCond[1384];
    m[666] = run?((((~m[158]&~m[335]&~m[922])|(m[158]&m[335]&~m[922]))&BiasedRNG[889])|(((m[158]&~m[335]&~m[922])|(~m[158]&m[335]&m[922]))&~BiasedRNG[889])|((~m[158]&~m[335]&m[922])|(m[158]&~m[335]&m[922])|(m[158]&m[335]&m[922]))):InitCond[1385];
    m[667] = run?((((~m[158]&~m[351]&~m[923])|(m[158]&m[351]&~m[923]))&BiasedRNG[890])|(((m[158]&~m[351]&~m[923])|(~m[158]&m[351]&m[923]))&~BiasedRNG[890])|((~m[158]&~m[351]&m[923])|(m[158]&~m[351]&m[923])|(m[158]&m[351]&m[923]))):InitCond[1386];
    m[668] = run?((((~m[159]&~m[367]&~m[924])|(m[159]&m[367]&~m[924]))&BiasedRNG[891])|(((m[159]&~m[367]&~m[924])|(~m[159]&m[367]&m[924]))&~BiasedRNG[891])|((~m[159]&~m[367]&m[924])|(m[159]&~m[367]&m[924])|(m[159]&m[367]&m[924]))):InitCond[1387];
    m[669] = run?((((~m[159]&~m[383]&~m[925])|(m[159]&m[383]&~m[925]))&BiasedRNG[892])|(((m[159]&~m[383]&~m[925])|(~m[159]&m[383]&m[925]))&~BiasedRNG[892])|((~m[159]&~m[383]&m[925])|(m[159]&~m[383]&m[925])|(m[159]&m[383]&m[925]))):InitCond[1388];
    m[670] = run?((((~m[159]&~m[399]&~m[926])|(m[159]&m[399]&~m[926]))&BiasedRNG[893])|(((m[159]&~m[399]&~m[926])|(~m[159]&m[399]&m[926]))&~BiasedRNG[893])|((~m[159]&~m[399]&m[926])|(m[159]&~m[399]&m[926])|(m[159]&m[399]&m[926]))):InitCond[1389];
    m[671] = run?((((~m[159]&~m[415]&~m[927])|(m[159]&m[415]&~m[927]))&BiasedRNG[894])|(((m[159]&~m[415]&~m[927])|(~m[159]&m[415]&m[927]))&~BiasedRNG[894])|((~m[159]&~m[415]&m[927])|(m[159]&~m[415]&m[927])|(m[159]&m[415]&m[927]))):InitCond[1390];
    m[929] = run?((((m[688]&~m[928]&~m[930]&~m[931]&~m[932])|(~m[688]&~m[928]&~m[930]&m[931]&~m[932])|(m[688]&m[928]&~m[930]&m[931]&~m[932])|(m[688]&~m[928]&m[930]&m[931]&~m[932])|(~m[688]&m[928]&~m[930]&~m[931]&m[932])|(~m[688]&~m[928]&m[930]&~m[931]&m[932])|(m[688]&m[928]&m[930]&~m[931]&m[932])|(~m[688]&m[928]&m[930]&m[931]&m[932]))&UnbiasedRNG[496])|((m[688]&~m[928]&~m[930]&m[931]&~m[932])|(~m[688]&~m[928]&~m[930]&~m[931]&m[932])|(m[688]&~m[928]&~m[930]&~m[931]&m[932])|(m[688]&m[928]&~m[930]&~m[931]&m[932])|(m[688]&~m[928]&m[930]&~m[931]&m[932])|(~m[688]&~m[928]&~m[930]&m[931]&m[932])|(m[688]&~m[928]&~m[930]&m[931]&m[932])|(~m[688]&m[928]&~m[930]&m[931]&m[932])|(m[688]&m[928]&~m[930]&m[931]&m[932])|(~m[688]&~m[928]&m[930]&m[931]&m[932])|(m[688]&~m[928]&m[930]&m[931]&m[932])|(m[688]&m[928]&m[930]&m[931]&m[932]))):InitCond[1391];
    m[934] = run?((((m[689]&~m[933]&~m[935]&~m[936]&~m[937])|(~m[689]&~m[933]&~m[935]&m[936]&~m[937])|(m[689]&m[933]&~m[935]&m[936]&~m[937])|(m[689]&~m[933]&m[935]&m[936]&~m[937])|(~m[689]&m[933]&~m[935]&~m[936]&m[937])|(~m[689]&~m[933]&m[935]&~m[936]&m[937])|(m[689]&m[933]&m[935]&~m[936]&m[937])|(~m[689]&m[933]&m[935]&m[936]&m[937]))&UnbiasedRNG[497])|((m[689]&~m[933]&~m[935]&m[936]&~m[937])|(~m[689]&~m[933]&~m[935]&~m[936]&m[937])|(m[689]&~m[933]&~m[935]&~m[936]&m[937])|(m[689]&m[933]&~m[935]&~m[936]&m[937])|(m[689]&~m[933]&m[935]&~m[936]&m[937])|(~m[689]&~m[933]&~m[935]&m[936]&m[937])|(m[689]&~m[933]&~m[935]&m[936]&m[937])|(~m[689]&m[933]&~m[935]&m[936]&m[937])|(m[689]&m[933]&~m[935]&m[936]&m[937])|(~m[689]&~m[933]&m[935]&m[936]&m[937])|(m[689]&~m[933]&m[935]&m[936]&m[937])|(m[689]&m[933]&m[935]&m[936]&m[937]))):InitCond[1392];
    m[939] = run?((((m[704]&~m[938]&~m[940]&~m[941]&~m[942])|(~m[704]&~m[938]&~m[940]&m[941]&~m[942])|(m[704]&m[938]&~m[940]&m[941]&~m[942])|(m[704]&~m[938]&m[940]&m[941]&~m[942])|(~m[704]&m[938]&~m[940]&~m[941]&m[942])|(~m[704]&~m[938]&m[940]&~m[941]&m[942])|(m[704]&m[938]&m[940]&~m[941]&m[942])|(~m[704]&m[938]&m[940]&m[941]&m[942]))&UnbiasedRNG[498])|((m[704]&~m[938]&~m[940]&m[941]&~m[942])|(~m[704]&~m[938]&~m[940]&~m[941]&m[942])|(m[704]&~m[938]&~m[940]&~m[941]&m[942])|(m[704]&m[938]&~m[940]&~m[941]&m[942])|(m[704]&~m[938]&m[940]&~m[941]&m[942])|(~m[704]&~m[938]&~m[940]&m[941]&m[942])|(m[704]&~m[938]&~m[940]&m[941]&m[942])|(~m[704]&m[938]&~m[940]&m[941]&m[942])|(m[704]&m[938]&~m[940]&m[941]&m[942])|(~m[704]&~m[938]&m[940]&m[941]&m[942])|(m[704]&~m[938]&m[940]&m[941]&m[942])|(m[704]&m[938]&m[940]&m[941]&m[942]))):InitCond[1393];
    m[944] = run?((((m[690]&~m[943]&~m[945]&~m[946]&~m[947])|(~m[690]&~m[943]&~m[945]&m[946]&~m[947])|(m[690]&m[943]&~m[945]&m[946]&~m[947])|(m[690]&~m[943]&m[945]&m[946]&~m[947])|(~m[690]&m[943]&~m[945]&~m[946]&m[947])|(~m[690]&~m[943]&m[945]&~m[946]&m[947])|(m[690]&m[943]&m[945]&~m[946]&m[947])|(~m[690]&m[943]&m[945]&m[946]&m[947]))&UnbiasedRNG[499])|((m[690]&~m[943]&~m[945]&m[946]&~m[947])|(~m[690]&~m[943]&~m[945]&~m[946]&m[947])|(m[690]&~m[943]&~m[945]&~m[946]&m[947])|(m[690]&m[943]&~m[945]&~m[946]&m[947])|(m[690]&~m[943]&m[945]&~m[946]&m[947])|(~m[690]&~m[943]&~m[945]&m[946]&m[947])|(m[690]&~m[943]&~m[945]&m[946]&m[947])|(~m[690]&m[943]&~m[945]&m[946]&m[947])|(m[690]&m[943]&~m[945]&m[946]&m[947])|(~m[690]&~m[943]&m[945]&m[946]&m[947])|(m[690]&~m[943]&m[945]&m[946]&m[947])|(m[690]&m[943]&m[945]&m[946]&m[947]))):InitCond[1394];
    m[949] = run?((((m[705]&~m[948]&~m[950]&~m[951]&~m[952])|(~m[705]&~m[948]&~m[950]&m[951]&~m[952])|(m[705]&m[948]&~m[950]&m[951]&~m[952])|(m[705]&~m[948]&m[950]&m[951]&~m[952])|(~m[705]&m[948]&~m[950]&~m[951]&m[952])|(~m[705]&~m[948]&m[950]&~m[951]&m[952])|(m[705]&m[948]&m[950]&~m[951]&m[952])|(~m[705]&m[948]&m[950]&m[951]&m[952]))&UnbiasedRNG[500])|((m[705]&~m[948]&~m[950]&m[951]&~m[952])|(~m[705]&~m[948]&~m[950]&~m[951]&m[952])|(m[705]&~m[948]&~m[950]&~m[951]&m[952])|(m[705]&m[948]&~m[950]&~m[951]&m[952])|(m[705]&~m[948]&m[950]&~m[951]&m[952])|(~m[705]&~m[948]&~m[950]&m[951]&m[952])|(m[705]&~m[948]&~m[950]&m[951]&m[952])|(~m[705]&m[948]&~m[950]&m[951]&m[952])|(m[705]&m[948]&~m[950]&m[951]&m[952])|(~m[705]&~m[948]&m[950]&m[951]&m[952])|(m[705]&~m[948]&m[950]&m[951]&m[952])|(m[705]&m[948]&m[950]&m[951]&m[952]))):InitCond[1395];
    m[954] = run?((((m[720]&~m[953]&~m[955]&~m[956]&~m[957])|(~m[720]&~m[953]&~m[955]&m[956]&~m[957])|(m[720]&m[953]&~m[955]&m[956]&~m[957])|(m[720]&~m[953]&m[955]&m[956]&~m[957])|(~m[720]&m[953]&~m[955]&~m[956]&m[957])|(~m[720]&~m[953]&m[955]&~m[956]&m[957])|(m[720]&m[953]&m[955]&~m[956]&m[957])|(~m[720]&m[953]&m[955]&m[956]&m[957]))&UnbiasedRNG[501])|((m[720]&~m[953]&~m[955]&m[956]&~m[957])|(~m[720]&~m[953]&~m[955]&~m[956]&m[957])|(m[720]&~m[953]&~m[955]&~m[956]&m[957])|(m[720]&m[953]&~m[955]&~m[956]&m[957])|(m[720]&~m[953]&m[955]&~m[956]&m[957])|(~m[720]&~m[953]&~m[955]&m[956]&m[957])|(m[720]&~m[953]&~m[955]&m[956]&m[957])|(~m[720]&m[953]&~m[955]&m[956]&m[957])|(m[720]&m[953]&~m[955]&m[956]&m[957])|(~m[720]&~m[953]&m[955]&m[956]&m[957])|(m[720]&~m[953]&m[955]&m[956]&m[957])|(m[720]&m[953]&m[955]&m[956]&m[957]))):InitCond[1396];
    m[959] = run?((((m[691]&~m[958]&~m[960]&~m[961]&~m[962])|(~m[691]&~m[958]&~m[960]&m[961]&~m[962])|(m[691]&m[958]&~m[960]&m[961]&~m[962])|(m[691]&~m[958]&m[960]&m[961]&~m[962])|(~m[691]&m[958]&~m[960]&~m[961]&m[962])|(~m[691]&~m[958]&m[960]&~m[961]&m[962])|(m[691]&m[958]&m[960]&~m[961]&m[962])|(~m[691]&m[958]&m[960]&m[961]&m[962]))&UnbiasedRNG[502])|((m[691]&~m[958]&~m[960]&m[961]&~m[962])|(~m[691]&~m[958]&~m[960]&~m[961]&m[962])|(m[691]&~m[958]&~m[960]&~m[961]&m[962])|(m[691]&m[958]&~m[960]&~m[961]&m[962])|(m[691]&~m[958]&m[960]&~m[961]&m[962])|(~m[691]&~m[958]&~m[960]&m[961]&m[962])|(m[691]&~m[958]&~m[960]&m[961]&m[962])|(~m[691]&m[958]&~m[960]&m[961]&m[962])|(m[691]&m[958]&~m[960]&m[961]&m[962])|(~m[691]&~m[958]&m[960]&m[961]&m[962])|(m[691]&~m[958]&m[960]&m[961]&m[962])|(m[691]&m[958]&m[960]&m[961]&m[962]))):InitCond[1397];
    m[964] = run?((((m[706]&~m[963]&~m[965]&~m[966]&~m[967])|(~m[706]&~m[963]&~m[965]&m[966]&~m[967])|(m[706]&m[963]&~m[965]&m[966]&~m[967])|(m[706]&~m[963]&m[965]&m[966]&~m[967])|(~m[706]&m[963]&~m[965]&~m[966]&m[967])|(~m[706]&~m[963]&m[965]&~m[966]&m[967])|(m[706]&m[963]&m[965]&~m[966]&m[967])|(~m[706]&m[963]&m[965]&m[966]&m[967]))&UnbiasedRNG[503])|((m[706]&~m[963]&~m[965]&m[966]&~m[967])|(~m[706]&~m[963]&~m[965]&~m[966]&m[967])|(m[706]&~m[963]&~m[965]&~m[966]&m[967])|(m[706]&m[963]&~m[965]&~m[966]&m[967])|(m[706]&~m[963]&m[965]&~m[966]&m[967])|(~m[706]&~m[963]&~m[965]&m[966]&m[967])|(m[706]&~m[963]&~m[965]&m[966]&m[967])|(~m[706]&m[963]&~m[965]&m[966]&m[967])|(m[706]&m[963]&~m[965]&m[966]&m[967])|(~m[706]&~m[963]&m[965]&m[966]&m[967])|(m[706]&~m[963]&m[965]&m[966]&m[967])|(m[706]&m[963]&m[965]&m[966]&m[967]))):InitCond[1398];
    m[969] = run?((((m[721]&~m[968]&~m[970]&~m[971]&~m[972])|(~m[721]&~m[968]&~m[970]&m[971]&~m[972])|(m[721]&m[968]&~m[970]&m[971]&~m[972])|(m[721]&~m[968]&m[970]&m[971]&~m[972])|(~m[721]&m[968]&~m[970]&~m[971]&m[972])|(~m[721]&~m[968]&m[970]&~m[971]&m[972])|(m[721]&m[968]&m[970]&~m[971]&m[972])|(~m[721]&m[968]&m[970]&m[971]&m[972]))&UnbiasedRNG[504])|((m[721]&~m[968]&~m[970]&m[971]&~m[972])|(~m[721]&~m[968]&~m[970]&~m[971]&m[972])|(m[721]&~m[968]&~m[970]&~m[971]&m[972])|(m[721]&m[968]&~m[970]&~m[971]&m[972])|(m[721]&~m[968]&m[970]&~m[971]&m[972])|(~m[721]&~m[968]&~m[970]&m[971]&m[972])|(m[721]&~m[968]&~m[970]&m[971]&m[972])|(~m[721]&m[968]&~m[970]&m[971]&m[972])|(m[721]&m[968]&~m[970]&m[971]&m[972])|(~m[721]&~m[968]&m[970]&m[971]&m[972])|(m[721]&~m[968]&m[970]&m[971]&m[972])|(m[721]&m[968]&m[970]&m[971]&m[972]))):InitCond[1399];
    m[974] = run?((((m[736]&~m[973]&~m[975]&~m[976]&~m[977])|(~m[736]&~m[973]&~m[975]&m[976]&~m[977])|(m[736]&m[973]&~m[975]&m[976]&~m[977])|(m[736]&~m[973]&m[975]&m[976]&~m[977])|(~m[736]&m[973]&~m[975]&~m[976]&m[977])|(~m[736]&~m[973]&m[975]&~m[976]&m[977])|(m[736]&m[973]&m[975]&~m[976]&m[977])|(~m[736]&m[973]&m[975]&m[976]&m[977]))&UnbiasedRNG[505])|((m[736]&~m[973]&~m[975]&m[976]&~m[977])|(~m[736]&~m[973]&~m[975]&~m[976]&m[977])|(m[736]&~m[973]&~m[975]&~m[976]&m[977])|(m[736]&m[973]&~m[975]&~m[976]&m[977])|(m[736]&~m[973]&m[975]&~m[976]&m[977])|(~m[736]&~m[973]&~m[975]&m[976]&m[977])|(m[736]&~m[973]&~m[975]&m[976]&m[977])|(~m[736]&m[973]&~m[975]&m[976]&m[977])|(m[736]&m[973]&~m[975]&m[976]&m[977])|(~m[736]&~m[973]&m[975]&m[976]&m[977])|(m[736]&~m[973]&m[975]&m[976]&m[977])|(m[736]&m[973]&m[975]&m[976]&m[977]))):InitCond[1400];
    m[979] = run?((((m[692]&~m[978]&~m[980]&~m[981]&~m[982])|(~m[692]&~m[978]&~m[980]&m[981]&~m[982])|(m[692]&m[978]&~m[980]&m[981]&~m[982])|(m[692]&~m[978]&m[980]&m[981]&~m[982])|(~m[692]&m[978]&~m[980]&~m[981]&m[982])|(~m[692]&~m[978]&m[980]&~m[981]&m[982])|(m[692]&m[978]&m[980]&~m[981]&m[982])|(~m[692]&m[978]&m[980]&m[981]&m[982]))&UnbiasedRNG[506])|((m[692]&~m[978]&~m[980]&m[981]&~m[982])|(~m[692]&~m[978]&~m[980]&~m[981]&m[982])|(m[692]&~m[978]&~m[980]&~m[981]&m[982])|(m[692]&m[978]&~m[980]&~m[981]&m[982])|(m[692]&~m[978]&m[980]&~m[981]&m[982])|(~m[692]&~m[978]&~m[980]&m[981]&m[982])|(m[692]&~m[978]&~m[980]&m[981]&m[982])|(~m[692]&m[978]&~m[980]&m[981]&m[982])|(m[692]&m[978]&~m[980]&m[981]&m[982])|(~m[692]&~m[978]&m[980]&m[981]&m[982])|(m[692]&~m[978]&m[980]&m[981]&m[982])|(m[692]&m[978]&m[980]&m[981]&m[982]))):InitCond[1401];
    m[984] = run?((((m[707]&~m[983]&~m[985]&~m[986]&~m[987])|(~m[707]&~m[983]&~m[985]&m[986]&~m[987])|(m[707]&m[983]&~m[985]&m[986]&~m[987])|(m[707]&~m[983]&m[985]&m[986]&~m[987])|(~m[707]&m[983]&~m[985]&~m[986]&m[987])|(~m[707]&~m[983]&m[985]&~m[986]&m[987])|(m[707]&m[983]&m[985]&~m[986]&m[987])|(~m[707]&m[983]&m[985]&m[986]&m[987]))&UnbiasedRNG[507])|((m[707]&~m[983]&~m[985]&m[986]&~m[987])|(~m[707]&~m[983]&~m[985]&~m[986]&m[987])|(m[707]&~m[983]&~m[985]&~m[986]&m[987])|(m[707]&m[983]&~m[985]&~m[986]&m[987])|(m[707]&~m[983]&m[985]&~m[986]&m[987])|(~m[707]&~m[983]&~m[985]&m[986]&m[987])|(m[707]&~m[983]&~m[985]&m[986]&m[987])|(~m[707]&m[983]&~m[985]&m[986]&m[987])|(m[707]&m[983]&~m[985]&m[986]&m[987])|(~m[707]&~m[983]&m[985]&m[986]&m[987])|(m[707]&~m[983]&m[985]&m[986]&m[987])|(m[707]&m[983]&m[985]&m[986]&m[987]))):InitCond[1402];
    m[989] = run?((((m[722]&~m[988]&~m[990]&~m[991]&~m[992])|(~m[722]&~m[988]&~m[990]&m[991]&~m[992])|(m[722]&m[988]&~m[990]&m[991]&~m[992])|(m[722]&~m[988]&m[990]&m[991]&~m[992])|(~m[722]&m[988]&~m[990]&~m[991]&m[992])|(~m[722]&~m[988]&m[990]&~m[991]&m[992])|(m[722]&m[988]&m[990]&~m[991]&m[992])|(~m[722]&m[988]&m[990]&m[991]&m[992]))&UnbiasedRNG[508])|((m[722]&~m[988]&~m[990]&m[991]&~m[992])|(~m[722]&~m[988]&~m[990]&~m[991]&m[992])|(m[722]&~m[988]&~m[990]&~m[991]&m[992])|(m[722]&m[988]&~m[990]&~m[991]&m[992])|(m[722]&~m[988]&m[990]&~m[991]&m[992])|(~m[722]&~m[988]&~m[990]&m[991]&m[992])|(m[722]&~m[988]&~m[990]&m[991]&m[992])|(~m[722]&m[988]&~m[990]&m[991]&m[992])|(m[722]&m[988]&~m[990]&m[991]&m[992])|(~m[722]&~m[988]&m[990]&m[991]&m[992])|(m[722]&~m[988]&m[990]&m[991]&m[992])|(m[722]&m[988]&m[990]&m[991]&m[992]))):InitCond[1403];
    m[994] = run?((((m[737]&~m[993]&~m[995]&~m[996]&~m[997])|(~m[737]&~m[993]&~m[995]&m[996]&~m[997])|(m[737]&m[993]&~m[995]&m[996]&~m[997])|(m[737]&~m[993]&m[995]&m[996]&~m[997])|(~m[737]&m[993]&~m[995]&~m[996]&m[997])|(~m[737]&~m[993]&m[995]&~m[996]&m[997])|(m[737]&m[993]&m[995]&~m[996]&m[997])|(~m[737]&m[993]&m[995]&m[996]&m[997]))&UnbiasedRNG[509])|((m[737]&~m[993]&~m[995]&m[996]&~m[997])|(~m[737]&~m[993]&~m[995]&~m[996]&m[997])|(m[737]&~m[993]&~m[995]&~m[996]&m[997])|(m[737]&m[993]&~m[995]&~m[996]&m[997])|(m[737]&~m[993]&m[995]&~m[996]&m[997])|(~m[737]&~m[993]&~m[995]&m[996]&m[997])|(m[737]&~m[993]&~m[995]&m[996]&m[997])|(~m[737]&m[993]&~m[995]&m[996]&m[997])|(m[737]&m[993]&~m[995]&m[996]&m[997])|(~m[737]&~m[993]&m[995]&m[996]&m[997])|(m[737]&~m[993]&m[995]&m[996]&m[997])|(m[737]&m[993]&m[995]&m[996]&m[997]))):InitCond[1404];
    m[999] = run?((((m[752]&~m[998]&~m[1000]&~m[1001]&~m[1002])|(~m[752]&~m[998]&~m[1000]&m[1001]&~m[1002])|(m[752]&m[998]&~m[1000]&m[1001]&~m[1002])|(m[752]&~m[998]&m[1000]&m[1001]&~m[1002])|(~m[752]&m[998]&~m[1000]&~m[1001]&m[1002])|(~m[752]&~m[998]&m[1000]&~m[1001]&m[1002])|(m[752]&m[998]&m[1000]&~m[1001]&m[1002])|(~m[752]&m[998]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[510])|((m[752]&~m[998]&~m[1000]&m[1001]&~m[1002])|(~m[752]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[752]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[752]&m[998]&~m[1000]&~m[1001]&m[1002])|(m[752]&~m[998]&m[1000]&~m[1001]&m[1002])|(~m[752]&~m[998]&~m[1000]&m[1001]&m[1002])|(m[752]&~m[998]&~m[1000]&m[1001]&m[1002])|(~m[752]&m[998]&~m[1000]&m[1001]&m[1002])|(m[752]&m[998]&~m[1000]&m[1001]&m[1002])|(~m[752]&~m[998]&m[1000]&m[1001]&m[1002])|(m[752]&~m[998]&m[1000]&m[1001]&m[1002])|(m[752]&m[998]&m[1000]&m[1001]&m[1002]))):InitCond[1405];
    m[1004] = run?((((m[693]&~m[1003]&~m[1005]&~m[1006]&~m[1007])|(~m[693]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(m[693]&m[1003]&~m[1005]&m[1006]&~m[1007])|(m[693]&~m[1003]&m[1005]&m[1006]&~m[1007])|(~m[693]&m[1003]&~m[1005]&~m[1006]&m[1007])|(~m[693]&~m[1003]&m[1005]&~m[1006]&m[1007])|(m[693]&m[1003]&m[1005]&~m[1006]&m[1007])|(~m[693]&m[1003]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[511])|((m[693]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(~m[693]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[693]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[693]&m[1003]&~m[1005]&~m[1006]&m[1007])|(m[693]&~m[1003]&m[1005]&~m[1006]&m[1007])|(~m[693]&~m[1003]&~m[1005]&m[1006]&m[1007])|(m[693]&~m[1003]&~m[1005]&m[1006]&m[1007])|(~m[693]&m[1003]&~m[1005]&m[1006]&m[1007])|(m[693]&m[1003]&~m[1005]&m[1006]&m[1007])|(~m[693]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[693]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[693]&m[1003]&m[1005]&m[1006]&m[1007]))):InitCond[1406];
    m[1009] = run?((((m[708]&~m[1008]&~m[1010]&~m[1011]&~m[1012])|(~m[708]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(m[708]&m[1008]&~m[1010]&m[1011]&~m[1012])|(m[708]&~m[1008]&m[1010]&m[1011]&~m[1012])|(~m[708]&m[1008]&~m[1010]&~m[1011]&m[1012])|(~m[708]&~m[1008]&m[1010]&~m[1011]&m[1012])|(m[708]&m[1008]&m[1010]&~m[1011]&m[1012])|(~m[708]&m[1008]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[512])|((m[708]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(~m[708]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[708]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[708]&m[1008]&~m[1010]&~m[1011]&m[1012])|(m[708]&~m[1008]&m[1010]&~m[1011]&m[1012])|(~m[708]&~m[1008]&~m[1010]&m[1011]&m[1012])|(m[708]&~m[1008]&~m[1010]&m[1011]&m[1012])|(~m[708]&m[1008]&~m[1010]&m[1011]&m[1012])|(m[708]&m[1008]&~m[1010]&m[1011]&m[1012])|(~m[708]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[708]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[708]&m[1008]&m[1010]&m[1011]&m[1012]))):InitCond[1407];
    m[1014] = run?((((m[723]&~m[1013]&~m[1015]&~m[1016]&~m[1017])|(~m[723]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(m[723]&m[1013]&~m[1015]&m[1016]&~m[1017])|(m[723]&~m[1013]&m[1015]&m[1016]&~m[1017])|(~m[723]&m[1013]&~m[1015]&~m[1016]&m[1017])|(~m[723]&~m[1013]&m[1015]&~m[1016]&m[1017])|(m[723]&m[1013]&m[1015]&~m[1016]&m[1017])|(~m[723]&m[1013]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[513])|((m[723]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(~m[723]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[723]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[723]&m[1013]&~m[1015]&~m[1016]&m[1017])|(m[723]&~m[1013]&m[1015]&~m[1016]&m[1017])|(~m[723]&~m[1013]&~m[1015]&m[1016]&m[1017])|(m[723]&~m[1013]&~m[1015]&m[1016]&m[1017])|(~m[723]&m[1013]&~m[1015]&m[1016]&m[1017])|(m[723]&m[1013]&~m[1015]&m[1016]&m[1017])|(~m[723]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[723]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[723]&m[1013]&m[1015]&m[1016]&m[1017]))):InitCond[1408];
    m[1019] = run?((((m[738]&~m[1018]&~m[1020]&~m[1021]&~m[1022])|(~m[738]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(m[738]&m[1018]&~m[1020]&m[1021]&~m[1022])|(m[738]&~m[1018]&m[1020]&m[1021]&~m[1022])|(~m[738]&m[1018]&~m[1020]&~m[1021]&m[1022])|(~m[738]&~m[1018]&m[1020]&~m[1021]&m[1022])|(m[738]&m[1018]&m[1020]&~m[1021]&m[1022])|(~m[738]&m[1018]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[514])|((m[738]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(~m[738]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[738]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[738]&m[1018]&~m[1020]&~m[1021]&m[1022])|(m[738]&~m[1018]&m[1020]&~m[1021]&m[1022])|(~m[738]&~m[1018]&~m[1020]&m[1021]&m[1022])|(m[738]&~m[1018]&~m[1020]&m[1021]&m[1022])|(~m[738]&m[1018]&~m[1020]&m[1021]&m[1022])|(m[738]&m[1018]&~m[1020]&m[1021]&m[1022])|(~m[738]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[738]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[738]&m[1018]&m[1020]&m[1021]&m[1022]))):InitCond[1409];
    m[1024] = run?((((m[753]&~m[1023]&~m[1025]&~m[1026]&~m[1027])|(~m[753]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(m[753]&m[1023]&~m[1025]&m[1026]&~m[1027])|(m[753]&~m[1023]&m[1025]&m[1026]&~m[1027])|(~m[753]&m[1023]&~m[1025]&~m[1026]&m[1027])|(~m[753]&~m[1023]&m[1025]&~m[1026]&m[1027])|(m[753]&m[1023]&m[1025]&~m[1026]&m[1027])|(~m[753]&m[1023]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[515])|((m[753]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(~m[753]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[753]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[753]&m[1023]&~m[1025]&~m[1026]&m[1027])|(m[753]&~m[1023]&m[1025]&~m[1026]&m[1027])|(~m[753]&~m[1023]&~m[1025]&m[1026]&m[1027])|(m[753]&~m[1023]&~m[1025]&m[1026]&m[1027])|(~m[753]&m[1023]&~m[1025]&m[1026]&m[1027])|(m[753]&m[1023]&~m[1025]&m[1026]&m[1027])|(~m[753]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[753]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[753]&m[1023]&m[1025]&m[1026]&m[1027]))):InitCond[1410];
    m[1029] = run?((((m[768]&~m[1028]&~m[1030]&~m[1031]&~m[1032])|(~m[768]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(m[768]&m[1028]&~m[1030]&m[1031]&~m[1032])|(m[768]&~m[1028]&m[1030]&m[1031]&~m[1032])|(~m[768]&m[1028]&~m[1030]&~m[1031]&m[1032])|(~m[768]&~m[1028]&m[1030]&~m[1031]&m[1032])|(m[768]&m[1028]&m[1030]&~m[1031]&m[1032])|(~m[768]&m[1028]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[516])|((m[768]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(~m[768]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[768]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[768]&m[1028]&~m[1030]&~m[1031]&m[1032])|(m[768]&~m[1028]&m[1030]&~m[1031]&m[1032])|(~m[768]&~m[1028]&~m[1030]&m[1031]&m[1032])|(m[768]&~m[1028]&~m[1030]&m[1031]&m[1032])|(~m[768]&m[1028]&~m[1030]&m[1031]&m[1032])|(m[768]&m[1028]&~m[1030]&m[1031]&m[1032])|(~m[768]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[768]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[768]&m[1028]&m[1030]&m[1031]&m[1032]))):InitCond[1411];
    m[1034] = run?((((m[694]&~m[1033]&~m[1035]&~m[1036]&~m[1037])|(~m[694]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(m[694]&m[1033]&~m[1035]&m[1036]&~m[1037])|(m[694]&~m[1033]&m[1035]&m[1036]&~m[1037])|(~m[694]&m[1033]&~m[1035]&~m[1036]&m[1037])|(~m[694]&~m[1033]&m[1035]&~m[1036]&m[1037])|(m[694]&m[1033]&m[1035]&~m[1036]&m[1037])|(~m[694]&m[1033]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[517])|((m[694]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(~m[694]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[694]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[694]&m[1033]&~m[1035]&~m[1036]&m[1037])|(m[694]&~m[1033]&m[1035]&~m[1036]&m[1037])|(~m[694]&~m[1033]&~m[1035]&m[1036]&m[1037])|(m[694]&~m[1033]&~m[1035]&m[1036]&m[1037])|(~m[694]&m[1033]&~m[1035]&m[1036]&m[1037])|(m[694]&m[1033]&~m[1035]&m[1036]&m[1037])|(~m[694]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[694]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[694]&m[1033]&m[1035]&m[1036]&m[1037]))):InitCond[1412];
    m[1039] = run?((((m[709]&~m[1038]&~m[1040]&~m[1041]&~m[1042])|(~m[709]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(m[709]&m[1038]&~m[1040]&m[1041]&~m[1042])|(m[709]&~m[1038]&m[1040]&m[1041]&~m[1042])|(~m[709]&m[1038]&~m[1040]&~m[1041]&m[1042])|(~m[709]&~m[1038]&m[1040]&~m[1041]&m[1042])|(m[709]&m[1038]&m[1040]&~m[1041]&m[1042])|(~m[709]&m[1038]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[518])|((m[709]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(~m[709]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[709]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[709]&m[1038]&~m[1040]&~m[1041]&m[1042])|(m[709]&~m[1038]&m[1040]&~m[1041]&m[1042])|(~m[709]&~m[1038]&~m[1040]&m[1041]&m[1042])|(m[709]&~m[1038]&~m[1040]&m[1041]&m[1042])|(~m[709]&m[1038]&~m[1040]&m[1041]&m[1042])|(m[709]&m[1038]&~m[1040]&m[1041]&m[1042])|(~m[709]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[709]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[709]&m[1038]&m[1040]&m[1041]&m[1042]))):InitCond[1413];
    m[1044] = run?((((m[724]&~m[1043]&~m[1045]&~m[1046]&~m[1047])|(~m[724]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(m[724]&m[1043]&~m[1045]&m[1046]&~m[1047])|(m[724]&~m[1043]&m[1045]&m[1046]&~m[1047])|(~m[724]&m[1043]&~m[1045]&~m[1046]&m[1047])|(~m[724]&~m[1043]&m[1045]&~m[1046]&m[1047])|(m[724]&m[1043]&m[1045]&~m[1046]&m[1047])|(~m[724]&m[1043]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[519])|((m[724]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(~m[724]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[724]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[724]&m[1043]&~m[1045]&~m[1046]&m[1047])|(m[724]&~m[1043]&m[1045]&~m[1046]&m[1047])|(~m[724]&~m[1043]&~m[1045]&m[1046]&m[1047])|(m[724]&~m[1043]&~m[1045]&m[1046]&m[1047])|(~m[724]&m[1043]&~m[1045]&m[1046]&m[1047])|(m[724]&m[1043]&~m[1045]&m[1046]&m[1047])|(~m[724]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[724]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[724]&m[1043]&m[1045]&m[1046]&m[1047]))):InitCond[1414];
    m[1049] = run?((((m[739]&~m[1048]&~m[1050]&~m[1051]&~m[1052])|(~m[739]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(m[739]&m[1048]&~m[1050]&m[1051]&~m[1052])|(m[739]&~m[1048]&m[1050]&m[1051]&~m[1052])|(~m[739]&m[1048]&~m[1050]&~m[1051]&m[1052])|(~m[739]&~m[1048]&m[1050]&~m[1051]&m[1052])|(m[739]&m[1048]&m[1050]&~m[1051]&m[1052])|(~m[739]&m[1048]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[520])|((m[739]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(~m[739]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[739]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[739]&m[1048]&~m[1050]&~m[1051]&m[1052])|(m[739]&~m[1048]&m[1050]&~m[1051]&m[1052])|(~m[739]&~m[1048]&~m[1050]&m[1051]&m[1052])|(m[739]&~m[1048]&~m[1050]&m[1051]&m[1052])|(~m[739]&m[1048]&~m[1050]&m[1051]&m[1052])|(m[739]&m[1048]&~m[1050]&m[1051]&m[1052])|(~m[739]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[739]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[739]&m[1048]&m[1050]&m[1051]&m[1052]))):InitCond[1415];
    m[1054] = run?((((m[754]&~m[1053]&~m[1055]&~m[1056]&~m[1057])|(~m[754]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(m[754]&m[1053]&~m[1055]&m[1056]&~m[1057])|(m[754]&~m[1053]&m[1055]&m[1056]&~m[1057])|(~m[754]&m[1053]&~m[1055]&~m[1056]&m[1057])|(~m[754]&~m[1053]&m[1055]&~m[1056]&m[1057])|(m[754]&m[1053]&m[1055]&~m[1056]&m[1057])|(~m[754]&m[1053]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[521])|((m[754]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(~m[754]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[754]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[754]&m[1053]&~m[1055]&~m[1056]&m[1057])|(m[754]&~m[1053]&m[1055]&~m[1056]&m[1057])|(~m[754]&~m[1053]&~m[1055]&m[1056]&m[1057])|(m[754]&~m[1053]&~m[1055]&m[1056]&m[1057])|(~m[754]&m[1053]&~m[1055]&m[1056]&m[1057])|(m[754]&m[1053]&~m[1055]&m[1056]&m[1057])|(~m[754]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[754]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[754]&m[1053]&m[1055]&m[1056]&m[1057]))):InitCond[1416];
    m[1059] = run?((((m[769]&~m[1058]&~m[1060]&~m[1061]&~m[1062])|(~m[769]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(m[769]&m[1058]&~m[1060]&m[1061]&~m[1062])|(m[769]&~m[1058]&m[1060]&m[1061]&~m[1062])|(~m[769]&m[1058]&~m[1060]&~m[1061]&m[1062])|(~m[769]&~m[1058]&m[1060]&~m[1061]&m[1062])|(m[769]&m[1058]&m[1060]&~m[1061]&m[1062])|(~m[769]&m[1058]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[522])|((m[769]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(~m[769]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[769]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[769]&m[1058]&~m[1060]&~m[1061]&m[1062])|(m[769]&~m[1058]&m[1060]&~m[1061]&m[1062])|(~m[769]&~m[1058]&~m[1060]&m[1061]&m[1062])|(m[769]&~m[1058]&~m[1060]&m[1061]&m[1062])|(~m[769]&m[1058]&~m[1060]&m[1061]&m[1062])|(m[769]&m[1058]&~m[1060]&m[1061]&m[1062])|(~m[769]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[769]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[769]&m[1058]&m[1060]&m[1061]&m[1062]))):InitCond[1417];
    m[1064] = run?((((m[784]&~m[1063]&~m[1065]&~m[1066]&~m[1067])|(~m[784]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(m[784]&m[1063]&~m[1065]&m[1066]&~m[1067])|(m[784]&~m[1063]&m[1065]&m[1066]&~m[1067])|(~m[784]&m[1063]&~m[1065]&~m[1066]&m[1067])|(~m[784]&~m[1063]&m[1065]&~m[1066]&m[1067])|(m[784]&m[1063]&m[1065]&~m[1066]&m[1067])|(~m[784]&m[1063]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[523])|((m[784]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(~m[784]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[784]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[784]&m[1063]&~m[1065]&~m[1066]&m[1067])|(m[784]&~m[1063]&m[1065]&~m[1066]&m[1067])|(~m[784]&~m[1063]&~m[1065]&m[1066]&m[1067])|(m[784]&~m[1063]&~m[1065]&m[1066]&m[1067])|(~m[784]&m[1063]&~m[1065]&m[1066]&m[1067])|(m[784]&m[1063]&~m[1065]&m[1066]&m[1067])|(~m[784]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[784]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[784]&m[1063]&m[1065]&m[1066]&m[1067]))):InitCond[1418];
    m[1069] = run?((((m[695]&~m[1068]&~m[1070]&~m[1071]&~m[1072])|(~m[695]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(m[695]&m[1068]&~m[1070]&m[1071]&~m[1072])|(m[695]&~m[1068]&m[1070]&m[1071]&~m[1072])|(~m[695]&m[1068]&~m[1070]&~m[1071]&m[1072])|(~m[695]&~m[1068]&m[1070]&~m[1071]&m[1072])|(m[695]&m[1068]&m[1070]&~m[1071]&m[1072])|(~m[695]&m[1068]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[524])|((m[695]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(~m[695]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[695]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[695]&m[1068]&~m[1070]&~m[1071]&m[1072])|(m[695]&~m[1068]&m[1070]&~m[1071]&m[1072])|(~m[695]&~m[1068]&~m[1070]&m[1071]&m[1072])|(m[695]&~m[1068]&~m[1070]&m[1071]&m[1072])|(~m[695]&m[1068]&~m[1070]&m[1071]&m[1072])|(m[695]&m[1068]&~m[1070]&m[1071]&m[1072])|(~m[695]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[695]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[695]&m[1068]&m[1070]&m[1071]&m[1072]))):InitCond[1419];
    m[1074] = run?((((m[710]&~m[1073]&~m[1075]&~m[1076]&~m[1077])|(~m[710]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(m[710]&m[1073]&~m[1075]&m[1076]&~m[1077])|(m[710]&~m[1073]&m[1075]&m[1076]&~m[1077])|(~m[710]&m[1073]&~m[1075]&~m[1076]&m[1077])|(~m[710]&~m[1073]&m[1075]&~m[1076]&m[1077])|(m[710]&m[1073]&m[1075]&~m[1076]&m[1077])|(~m[710]&m[1073]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[525])|((m[710]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(~m[710]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[710]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[710]&m[1073]&~m[1075]&~m[1076]&m[1077])|(m[710]&~m[1073]&m[1075]&~m[1076]&m[1077])|(~m[710]&~m[1073]&~m[1075]&m[1076]&m[1077])|(m[710]&~m[1073]&~m[1075]&m[1076]&m[1077])|(~m[710]&m[1073]&~m[1075]&m[1076]&m[1077])|(m[710]&m[1073]&~m[1075]&m[1076]&m[1077])|(~m[710]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[710]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[710]&m[1073]&m[1075]&m[1076]&m[1077]))):InitCond[1420];
    m[1079] = run?((((m[725]&~m[1078]&~m[1080]&~m[1081]&~m[1082])|(~m[725]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(m[725]&m[1078]&~m[1080]&m[1081]&~m[1082])|(m[725]&~m[1078]&m[1080]&m[1081]&~m[1082])|(~m[725]&m[1078]&~m[1080]&~m[1081]&m[1082])|(~m[725]&~m[1078]&m[1080]&~m[1081]&m[1082])|(m[725]&m[1078]&m[1080]&~m[1081]&m[1082])|(~m[725]&m[1078]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[526])|((m[725]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(~m[725]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[725]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[725]&m[1078]&~m[1080]&~m[1081]&m[1082])|(m[725]&~m[1078]&m[1080]&~m[1081]&m[1082])|(~m[725]&~m[1078]&~m[1080]&m[1081]&m[1082])|(m[725]&~m[1078]&~m[1080]&m[1081]&m[1082])|(~m[725]&m[1078]&~m[1080]&m[1081]&m[1082])|(m[725]&m[1078]&~m[1080]&m[1081]&m[1082])|(~m[725]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[725]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[725]&m[1078]&m[1080]&m[1081]&m[1082]))):InitCond[1421];
    m[1084] = run?((((m[740]&~m[1083]&~m[1085]&~m[1086]&~m[1087])|(~m[740]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(m[740]&m[1083]&~m[1085]&m[1086]&~m[1087])|(m[740]&~m[1083]&m[1085]&m[1086]&~m[1087])|(~m[740]&m[1083]&~m[1085]&~m[1086]&m[1087])|(~m[740]&~m[1083]&m[1085]&~m[1086]&m[1087])|(m[740]&m[1083]&m[1085]&~m[1086]&m[1087])|(~m[740]&m[1083]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[527])|((m[740]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(~m[740]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[740]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[740]&m[1083]&~m[1085]&~m[1086]&m[1087])|(m[740]&~m[1083]&m[1085]&~m[1086]&m[1087])|(~m[740]&~m[1083]&~m[1085]&m[1086]&m[1087])|(m[740]&~m[1083]&~m[1085]&m[1086]&m[1087])|(~m[740]&m[1083]&~m[1085]&m[1086]&m[1087])|(m[740]&m[1083]&~m[1085]&m[1086]&m[1087])|(~m[740]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[740]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[740]&m[1083]&m[1085]&m[1086]&m[1087]))):InitCond[1422];
    m[1089] = run?((((m[755]&~m[1088]&~m[1090]&~m[1091]&~m[1092])|(~m[755]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(m[755]&m[1088]&~m[1090]&m[1091]&~m[1092])|(m[755]&~m[1088]&m[1090]&m[1091]&~m[1092])|(~m[755]&m[1088]&~m[1090]&~m[1091]&m[1092])|(~m[755]&~m[1088]&m[1090]&~m[1091]&m[1092])|(m[755]&m[1088]&m[1090]&~m[1091]&m[1092])|(~m[755]&m[1088]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[528])|((m[755]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(~m[755]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[755]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[755]&m[1088]&~m[1090]&~m[1091]&m[1092])|(m[755]&~m[1088]&m[1090]&~m[1091]&m[1092])|(~m[755]&~m[1088]&~m[1090]&m[1091]&m[1092])|(m[755]&~m[1088]&~m[1090]&m[1091]&m[1092])|(~m[755]&m[1088]&~m[1090]&m[1091]&m[1092])|(m[755]&m[1088]&~m[1090]&m[1091]&m[1092])|(~m[755]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[755]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[755]&m[1088]&m[1090]&m[1091]&m[1092]))):InitCond[1423];
    m[1094] = run?((((m[770]&~m[1093]&~m[1095]&~m[1096]&~m[1097])|(~m[770]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(m[770]&m[1093]&~m[1095]&m[1096]&~m[1097])|(m[770]&~m[1093]&m[1095]&m[1096]&~m[1097])|(~m[770]&m[1093]&~m[1095]&~m[1096]&m[1097])|(~m[770]&~m[1093]&m[1095]&~m[1096]&m[1097])|(m[770]&m[1093]&m[1095]&~m[1096]&m[1097])|(~m[770]&m[1093]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[529])|((m[770]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(~m[770]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[770]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[770]&m[1093]&~m[1095]&~m[1096]&m[1097])|(m[770]&~m[1093]&m[1095]&~m[1096]&m[1097])|(~m[770]&~m[1093]&~m[1095]&m[1096]&m[1097])|(m[770]&~m[1093]&~m[1095]&m[1096]&m[1097])|(~m[770]&m[1093]&~m[1095]&m[1096]&m[1097])|(m[770]&m[1093]&~m[1095]&m[1096]&m[1097])|(~m[770]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[770]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[770]&m[1093]&m[1095]&m[1096]&m[1097]))):InitCond[1424];
    m[1099] = run?((((m[785]&~m[1098]&~m[1100]&~m[1101]&~m[1102])|(~m[785]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(m[785]&m[1098]&~m[1100]&m[1101]&~m[1102])|(m[785]&~m[1098]&m[1100]&m[1101]&~m[1102])|(~m[785]&m[1098]&~m[1100]&~m[1101]&m[1102])|(~m[785]&~m[1098]&m[1100]&~m[1101]&m[1102])|(m[785]&m[1098]&m[1100]&~m[1101]&m[1102])|(~m[785]&m[1098]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[530])|((m[785]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(~m[785]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[785]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[785]&m[1098]&~m[1100]&~m[1101]&m[1102])|(m[785]&~m[1098]&m[1100]&~m[1101]&m[1102])|(~m[785]&~m[1098]&~m[1100]&m[1101]&m[1102])|(m[785]&~m[1098]&~m[1100]&m[1101]&m[1102])|(~m[785]&m[1098]&~m[1100]&m[1101]&m[1102])|(m[785]&m[1098]&~m[1100]&m[1101]&m[1102])|(~m[785]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[785]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[785]&m[1098]&m[1100]&m[1101]&m[1102]))):InitCond[1425];
    m[1104] = run?((((m[800]&~m[1103]&~m[1105]&~m[1106]&~m[1107])|(~m[800]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(m[800]&m[1103]&~m[1105]&m[1106]&~m[1107])|(m[800]&~m[1103]&m[1105]&m[1106]&~m[1107])|(~m[800]&m[1103]&~m[1105]&~m[1106]&m[1107])|(~m[800]&~m[1103]&m[1105]&~m[1106]&m[1107])|(m[800]&m[1103]&m[1105]&~m[1106]&m[1107])|(~m[800]&m[1103]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[531])|((m[800]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(~m[800]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[800]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[800]&m[1103]&~m[1105]&~m[1106]&m[1107])|(m[800]&~m[1103]&m[1105]&~m[1106]&m[1107])|(~m[800]&~m[1103]&~m[1105]&m[1106]&m[1107])|(m[800]&~m[1103]&~m[1105]&m[1106]&m[1107])|(~m[800]&m[1103]&~m[1105]&m[1106]&m[1107])|(m[800]&m[1103]&~m[1105]&m[1106]&m[1107])|(~m[800]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[800]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[800]&m[1103]&m[1105]&m[1106]&m[1107]))):InitCond[1426];
    m[1109] = run?((((m[696]&~m[1108]&~m[1110]&~m[1111]&~m[1112])|(~m[696]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(m[696]&m[1108]&~m[1110]&m[1111]&~m[1112])|(m[696]&~m[1108]&m[1110]&m[1111]&~m[1112])|(~m[696]&m[1108]&~m[1110]&~m[1111]&m[1112])|(~m[696]&~m[1108]&m[1110]&~m[1111]&m[1112])|(m[696]&m[1108]&m[1110]&~m[1111]&m[1112])|(~m[696]&m[1108]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[532])|((m[696]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(~m[696]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[696]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[696]&m[1108]&~m[1110]&~m[1111]&m[1112])|(m[696]&~m[1108]&m[1110]&~m[1111]&m[1112])|(~m[696]&~m[1108]&~m[1110]&m[1111]&m[1112])|(m[696]&~m[1108]&~m[1110]&m[1111]&m[1112])|(~m[696]&m[1108]&~m[1110]&m[1111]&m[1112])|(m[696]&m[1108]&~m[1110]&m[1111]&m[1112])|(~m[696]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[696]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[696]&m[1108]&m[1110]&m[1111]&m[1112]))):InitCond[1427];
    m[1114] = run?((((m[711]&~m[1113]&~m[1115]&~m[1116]&~m[1117])|(~m[711]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(m[711]&m[1113]&~m[1115]&m[1116]&~m[1117])|(m[711]&~m[1113]&m[1115]&m[1116]&~m[1117])|(~m[711]&m[1113]&~m[1115]&~m[1116]&m[1117])|(~m[711]&~m[1113]&m[1115]&~m[1116]&m[1117])|(m[711]&m[1113]&m[1115]&~m[1116]&m[1117])|(~m[711]&m[1113]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[533])|((m[711]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(~m[711]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[711]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[711]&m[1113]&~m[1115]&~m[1116]&m[1117])|(m[711]&~m[1113]&m[1115]&~m[1116]&m[1117])|(~m[711]&~m[1113]&~m[1115]&m[1116]&m[1117])|(m[711]&~m[1113]&~m[1115]&m[1116]&m[1117])|(~m[711]&m[1113]&~m[1115]&m[1116]&m[1117])|(m[711]&m[1113]&~m[1115]&m[1116]&m[1117])|(~m[711]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[711]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[711]&m[1113]&m[1115]&m[1116]&m[1117]))):InitCond[1428];
    m[1119] = run?((((m[726]&~m[1118]&~m[1120]&~m[1121]&~m[1122])|(~m[726]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(m[726]&m[1118]&~m[1120]&m[1121]&~m[1122])|(m[726]&~m[1118]&m[1120]&m[1121]&~m[1122])|(~m[726]&m[1118]&~m[1120]&~m[1121]&m[1122])|(~m[726]&~m[1118]&m[1120]&~m[1121]&m[1122])|(m[726]&m[1118]&m[1120]&~m[1121]&m[1122])|(~m[726]&m[1118]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[534])|((m[726]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(~m[726]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[726]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[726]&m[1118]&~m[1120]&~m[1121]&m[1122])|(m[726]&~m[1118]&m[1120]&~m[1121]&m[1122])|(~m[726]&~m[1118]&~m[1120]&m[1121]&m[1122])|(m[726]&~m[1118]&~m[1120]&m[1121]&m[1122])|(~m[726]&m[1118]&~m[1120]&m[1121]&m[1122])|(m[726]&m[1118]&~m[1120]&m[1121]&m[1122])|(~m[726]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[726]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[726]&m[1118]&m[1120]&m[1121]&m[1122]))):InitCond[1429];
    m[1124] = run?((((m[741]&~m[1123]&~m[1125]&~m[1126]&~m[1127])|(~m[741]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(m[741]&m[1123]&~m[1125]&m[1126]&~m[1127])|(m[741]&~m[1123]&m[1125]&m[1126]&~m[1127])|(~m[741]&m[1123]&~m[1125]&~m[1126]&m[1127])|(~m[741]&~m[1123]&m[1125]&~m[1126]&m[1127])|(m[741]&m[1123]&m[1125]&~m[1126]&m[1127])|(~m[741]&m[1123]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[535])|((m[741]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(~m[741]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[741]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[741]&m[1123]&~m[1125]&~m[1126]&m[1127])|(m[741]&~m[1123]&m[1125]&~m[1126]&m[1127])|(~m[741]&~m[1123]&~m[1125]&m[1126]&m[1127])|(m[741]&~m[1123]&~m[1125]&m[1126]&m[1127])|(~m[741]&m[1123]&~m[1125]&m[1126]&m[1127])|(m[741]&m[1123]&~m[1125]&m[1126]&m[1127])|(~m[741]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[741]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[741]&m[1123]&m[1125]&m[1126]&m[1127]))):InitCond[1430];
    m[1129] = run?((((m[756]&~m[1128]&~m[1130]&~m[1131]&~m[1132])|(~m[756]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(m[756]&m[1128]&~m[1130]&m[1131]&~m[1132])|(m[756]&~m[1128]&m[1130]&m[1131]&~m[1132])|(~m[756]&m[1128]&~m[1130]&~m[1131]&m[1132])|(~m[756]&~m[1128]&m[1130]&~m[1131]&m[1132])|(m[756]&m[1128]&m[1130]&~m[1131]&m[1132])|(~m[756]&m[1128]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[536])|((m[756]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(~m[756]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[756]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[756]&m[1128]&~m[1130]&~m[1131]&m[1132])|(m[756]&~m[1128]&m[1130]&~m[1131]&m[1132])|(~m[756]&~m[1128]&~m[1130]&m[1131]&m[1132])|(m[756]&~m[1128]&~m[1130]&m[1131]&m[1132])|(~m[756]&m[1128]&~m[1130]&m[1131]&m[1132])|(m[756]&m[1128]&~m[1130]&m[1131]&m[1132])|(~m[756]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[756]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[756]&m[1128]&m[1130]&m[1131]&m[1132]))):InitCond[1431];
    m[1134] = run?((((m[771]&~m[1133]&~m[1135]&~m[1136]&~m[1137])|(~m[771]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(m[771]&m[1133]&~m[1135]&m[1136]&~m[1137])|(m[771]&~m[1133]&m[1135]&m[1136]&~m[1137])|(~m[771]&m[1133]&~m[1135]&~m[1136]&m[1137])|(~m[771]&~m[1133]&m[1135]&~m[1136]&m[1137])|(m[771]&m[1133]&m[1135]&~m[1136]&m[1137])|(~m[771]&m[1133]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[537])|((m[771]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(~m[771]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[771]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[771]&m[1133]&~m[1135]&~m[1136]&m[1137])|(m[771]&~m[1133]&m[1135]&~m[1136]&m[1137])|(~m[771]&~m[1133]&~m[1135]&m[1136]&m[1137])|(m[771]&~m[1133]&~m[1135]&m[1136]&m[1137])|(~m[771]&m[1133]&~m[1135]&m[1136]&m[1137])|(m[771]&m[1133]&~m[1135]&m[1136]&m[1137])|(~m[771]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[771]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[771]&m[1133]&m[1135]&m[1136]&m[1137]))):InitCond[1432];
    m[1139] = run?((((m[786]&~m[1138]&~m[1140]&~m[1141]&~m[1142])|(~m[786]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(m[786]&m[1138]&~m[1140]&m[1141]&~m[1142])|(m[786]&~m[1138]&m[1140]&m[1141]&~m[1142])|(~m[786]&m[1138]&~m[1140]&~m[1141]&m[1142])|(~m[786]&~m[1138]&m[1140]&~m[1141]&m[1142])|(m[786]&m[1138]&m[1140]&~m[1141]&m[1142])|(~m[786]&m[1138]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[538])|((m[786]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(~m[786]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[786]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[786]&m[1138]&~m[1140]&~m[1141]&m[1142])|(m[786]&~m[1138]&m[1140]&~m[1141]&m[1142])|(~m[786]&~m[1138]&~m[1140]&m[1141]&m[1142])|(m[786]&~m[1138]&~m[1140]&m[1141]&m[1142])|(~m[786]&m[1138]&~m[1140]&m[1141]&m[1142])|(m[786]&m[1138]&~m[1140]&m[1141]&m[1142])|(~m[786]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[786]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[786]&m[1138]&m[1140]&m[1141]&m[1142]))):InitCond[1433];
    m[1144] = run?((((m[801]&~m[1143]&~m[1145]&~m[1146]&~m[1147])|(~m[801]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(m[801]&m[1143]&~m[1145]&m[1146]&~m[1147])|(m[801]&~m[1143]&m[1145]&m[1146]&~m[1147])|(~m[801]&m[1143]&~m[1145]&~m[1146]&m[1147])|(~m[801]&~m[1143]&m[1145]&~m[1146]&m[1147])|(m[801]&m[1143]&m[1145]&~m[1146]&m[1147])|(~m[801]&m[1143]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[539])|((m[801]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(~m[801]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[801]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[801]&m[1143]&~m[1145]&~m[1146]&m[1147])|(m[801]&~m[1143]&m[1145]&~m[1146]&m[1147])|(~m[801]&~m[1143]&~m[1145]&m[1146]&m[1147])|(m[801]&~m[1143]&~m[1145]&m[1146]&m[1147])|(~m[801]&m[1143]&~m[1145]&m[1146]&m[1147])|(m[801]&m[1143]&~m[1145]&m[1146]&m[1147])|(~m[801]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[801]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[801]&m[1143]&m[1145]&m[1146]&m[1147]))):InitCond[1434];
    m[1149] = run?((((m[816]&~m[1148]&~m[1150]&~m[1151]&~m[1152])|(~m[816]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(m[816]&m[1148]&~m[1150]&m[1151]&~m[1152])|(m[816]&~m[1148]&m[1150]&m[1151]&~m[1152])|(~m[816]&m[1148]&~m[1150]&~m[1151]&m[1152])|(~m[816]&~m[1148]&m[1150]&~m[1151]&m[1152])|(m[816]&m[1148]&m[1150]&~m[1151]&m[1152])|(~m[816]&m[1148]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[540])|((m[816]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(~m[816]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[816]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[816]&m[1148]&~m[1150]&~m[1151]&m[1152])|(m[816]&~m[1148]&m[1150]&~m[1151]&m[1152])|(~m[816]&~m[1148]&~m[1150]&m[1151]&m[1152])|(m[816]&~m[1148]&~m[1150]&m[1151]&m[1152])|(~m[816]&m[1148]&~m[1150]&m[1151]&m[1152])|(m[816]&m[1148]&~m[1150]&m[1151]&m[1152])|(~m[816]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[816]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[816]&m[1148]&m[1150]&m[1151]&m[1152]))):InitCond[1435];
    m[1154] = run?((((m[697]&~m[1153]&~m[1155]&~m[1156]&~m[1157])|(~m[697]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(m[697]&m[1153]&~m[1155]&m[1156]&~m[1157])|(m[697]&~m[1153]&m[1155]&m[1156]&~m[1157])|(~m[697]&m[1153]&~m[1155]&~m[1156]&m[1157])|(~m[697]&~m[1153]&m[1155]&~m[1156]&m[1157])|(m[697]&m[1153]&m[1155]&~m[1156]&m[1157])|(~m[697]&m[1153]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[541])|((m[697]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(~m[697]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[697]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[697]&m[1153]&~m[1155]&~m[1156]&m[1157])|(m[697]&~m[1153]&m[1155]&~m[1156]&m[1157])|(~m[697]&~m[1153]&~m[1155]&m[1156]&m[1157])|(m[697]&~m[1153]&~m[1155]&m[1156]&m[1157])|(~m[697]&m[1153]&~m[1155]&m[1156]&m[1157])|(m[697]&m[1153]&~m[1155]&m[1156]&m[1157])|(~m[697]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[697]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[697]&m[1153]&m[1155]&m[1156]&m[1157]))):InitCond[1436];
    m[1159] = run?((((m[712]&~m[1158]&~m[1160]&~m[1161]&~m[1162])|(~m[712]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(m[712]&m[1158]&~m[1160]&m[1161]&~m[1162])|(m[712]&~m[1158]&m[1160]&m[1161]&~m[1162])|(~m[712]&m[1158]&~m[1160]&~m[1161]&m[1162])|(~m[712]&~m[1158]&m[1160]&~m[1161]&m[1162])|(m[712]&m[1158]&m[1160]&~m[1161]&m[1162])|(~m[712]&m[1158]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[542])|((m[712]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(~m[712]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[712]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[712]&m[1158]&~m[1160]&~m[1161]&m[1162])|(m[712]&~m[1158]&m[1160]&~m[1161]&m[1162])|(~m[712]&~m[1158]&~m[1160]&m[1161]&m[1162])|(m[712]&~m[1158]&~m[1160]&m[1161]&m[1162])|(~m[712]&m[1158]&~m[1160]&m[1161]&m[1162])|(m[712]&m[1158]&~m[1160]&m[1161]&m[1162])|(~m[712]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[712]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[712]&m[1158]&m[1160]&m[1161]&m[1162]))):InitCond[1437];
    m[1164] = run?((((m[727]&~m[1163]&~m[1165]&~m[1166]&~m[1167])|(~m[727]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(m[727]&m[1163]&~m[1165]&m[1166]&~m[1167])|(m[727]&~m[1163]&m[1165]&m[1166]&~m[1167])|(~m[727]&m[1163]&~m[1165]&~m[1166]&m[1167])|(~m[727]&~m[1163]&m[1165]&~m[1166]&m[1167])|(m[727]&m[1163]&m[1165]&~m[1166]&m[1167])|(~m[727]&m[1163]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[543])|((m[727]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(~m[727]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[727]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[727]&m[1163]&~m[1165]&~m[1166]&m[1167])|(m[727]&~m[1163]&m[1165]&~m[1166]&m[1167])|(~m[727]&~m[1163]&~m[1165]&m[1166]&m[1167])|(m[727]&~m[1163]&~m[1165]&m[1166]&m[1167])|(~m[727]&m[1163]&~m[1165]&m[1166]&m[1167])|(m[727]&m[1163]&~m[1165]&m[1166]&m[1167])|(~m[727]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[727]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[727]&m[1163]&m[1165]&m[1166]&m[1167]))):InitCond[1438];
    m[1169] = run?((((m[742]&~m[1168]&~m[1170]&~m[1171]&~m[1172])|(~m[742]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(m[742]&m[1168]&~m[1170]&m[1171]&~m[1172])|(m[742]&~m[1168]&m[1170]&m[1171]&~m[1172])|(~m[742]&m[1168]&~m[1170]&~m[1171]&m[1172])|(~m[742]&~m[1168]&m[1170]&~m[1171]&m[1172])|(m[742]&m[1168]&m[1170]&~m[1171]&m[1172])|(~m[742]&m[1168]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[544])|((m[742]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(~m[742]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[742]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[742]&m[1168]&~m[1170]&~m[1171]&m[1172])|(m[742]&~m[1168]&m[1170]&~m[1171]&m[1172])|(~m[742]&~m[1168]&~m[1170]&m[1171]&m[1172])|(m[742]&~m[1168]&~m[1170]&m[1171]&m[1172])|(~m[742]&m[1168]&~m[1170]&m[1171]&m[1172])|(m[742]&m[1168]&~m[1170]&m[1171]&m[1172])|(~m[742]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[742]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[742]&m[1168]&m[1170]&m[1171]&m[1172]))):InitCond[1439];
    m[1174] = run?((((m[757]&~m[1173]&~m[1175]&~m[1176]&~m[1177])|(~m[757]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(m[757]&m[1173]&~m[1175]&m[1176]&~m[1177])|(m[757]&~m[1173]&m[1175]&m[1176]&~m[1177])|(~m[757]&m[1173]&~m[1175]&~m[1176]&m[1177])|(~m[757]&~m[1173]&m[1175]&~m[1176]&m[1177])|(m[757]&m[1173]&m[1175]&~m[1176]&m[1177])|(~m[757]&m[1173]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[545])|((m[757]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(~m[757]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[757]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[757]&m[1173]&~m[1175]&~m[1176]&m[1177])|(m[757]&~m[1173]&m[1175]&~m[1176]&m[1177])|(~m[757]&~m[1173]&~m[1175]&m[1176]&m[1177])|(m[757]&~m[1173]&~m[1175]&m[1176]&m[1177])|(~m[757]&m[1173]&~m[1175]&m[1176]&m[1177])|(m[757]&m[1173]&~m[1175]&m[1176]&m[1177])|(~m[757]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[757]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[757]&m[1173]&m[1175]&m[1176]&m[1177]))):InitCond[1440];
    m[1179] = run?((((m[772]&~m[1178]&~m[1180]&~m[1181]&~m[1182])|(~m[772]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(m[772]&m[1178]&~m[1180]&m[1181]&~m[1182])|(m[772]&~m[1178]&m[1180]&m[1181]&~m[1182])|(~m[772]&m[1178]&~m[1180]&~m[1181]&m[1182])|(~m[772]&~m[1178]&m[1180]&~m[1181]&m[1182])|(m[772]&m[1178]&m[1180]&~m[1181]&m[1182])|(~m[772]&m[1178]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[546])|((m[772]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(~m[772]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[772]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[772]&m[1178]&~m[1180]&~m[1181]&m[1182])|(m[772]&~m[1178]&m[1180]&~m[1181]&m[1182])|(~m[772]&~m[1178]&~m[1180]&m[1181]&m[1182])|(m[772]&~m[1178]&~m[1180]&m[1181]&m[1182])|(~m[772]&m[1178]&~m[1180]&m[1181]&m[1182])|(m[772]&m[1178]&~m[1180]&m[1181]&m[1182])|(~m[772]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[772]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[772]&m[1178]&m[1180]&m[1181]&m[1182]))):InitCond[1441];
    m[1184] = run?((((m[787]&~m[1183]&~m[1185]&~m[1186]&~m[1187])|(~m[787]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(m[787]&m[1183]&~m[1185]&m[1186]&~m[1187])|(m[787]&~m[1183]&m[1185]&m[1186]&~m[1187])|(~m[787]&m[1183]&~m[1185]&~m[1186]&m[1187])|(~m[787]&~m[1183]&m[1185]&~m[1186]&m[1187])|(m[787]&m[1183]&m[1185]&~m[1186]&m[1187])|(~m[787]&m[1183]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[547])|((m[787]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(~m[787]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[787]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[787]&m[1183]&~m[1185]&~m[1186]&m[1187])|(m[787]&~m[1183]&m[1185]&~m[1186]&m[1187])|(~m[787]&~m[1183]&~m[1185]&m[1186]&m[1187])|(m[787]&~m[1183]&~m[1185]&m[1186]&m[1187])|(~m[787]&m[1183]&~m[1185]&m[1186]&m[1187])|(m[787]&m[1183]&~m[1185]&m[1186]&m[1187])|(~m[787]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[787]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[787]&m[1183]&m[1185]&m[1186]&m[1187]))):InitCond[1442];
    m[1189] = run?((((m[802]&~m[1188]&~m[1190]&~m[1191]&~m[1192])|(~m[802]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(m[802]&m[1188]&~m[1190]&m[1191]&~m[1192])|(m[802]&~m[1188]&m[1190]&m[1191]&~m[1192])|(~m[802]&m[1188]&~m[1190]&~m[1191]&m[1192])|(~m[802]&~m[1188]&m[1190]&~m[1191]&m[1192])|(m[802]&m[1188]&m[1190]&~m[1191]&m[1192])|(~m[802]&m[1188]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[548])|((m[802]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(~m[802]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[802]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[802]&m[1188]&~m[1190]&~m[1191]&m[1192])|(m[802]&~m[1188]&m[1190]&~m[1191]&m[1192])|(~m[802]&~m[1188]&~m[1190]&m[1191]&m[1192])|(m[802]&~m[1188]&~m[1190]&m[1191]&m[1192])|(~m[802]&m[1188]&~m[1190]&m[1191]&m[1192])|(m[802]&m[1188]&~m[1190]&m[1191]&m[1192])|(~m[802]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[802]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[802]&m[1188]&m[1190]&m[1191]&m[1192]))):InitCond[1443];
    m[1194] = run?((((m[817]&~m[1193]&~m[1195]&~m[1196]&~m[1197])|(~m[817]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(m[817]&m[1193]&~m[1195]&m[1196]&~m[1197])|(m[817]&~m[1193]&m[1195]&m[1196]&~m[1197])|(~m[817]&m[1193]&~m[1195]&~m[1196]&m[1197])|(~m[817]&~m[1193]&m[1195]&~m[1196]&m[1197])|(m[817]&m[1193]&m[1195]&~m[1196]&m[1197])|(~m[817]&m[1193]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[549])|((m[817]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(~m[817]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[817]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[817]&m[1193]&~m[1195]&~m[1196]&m[1197])|(m[817]&~m[1193]&m[1195]&~m[1196]&m[1197])|(~m[817]&~m[1193]&~m[1195]&m[1196]&m[1197])|(m[817]&~m[1193]&~m[1195]&m[1196]&m[1197])|(~m[817]&m[1193]&~m[1195]&m[1196]&m[1197])|(m[817]&m[1193]&~m[1195]&m[1196]&m[1197])|(~m[817]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[817]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[817]&m[1193]&m[1195]&m[1196]&m[1197]))):InitCond[1444];
    m[1199] = run?((((m[832]&~m[1198]&~m[1200]&~m[1201]&~m[1202])|(~m[832]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(m[832]&m[1198]&~m[1200]&m[1201]&~m[1202])|(m[832]&~m[1198]&m[1200]&m[1201]&~m[1202])|(~m[832]&m[1198]&~m[1200]&~m[1201]&m[1202])|(~m[832]&~m[1198]&m[1200]&~m[1201]&m[1202])|(m[832]&m[1198]&m[1200]&~m[1201]&m[1202])|(~m[832]&m[1198]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[550])|((m[832]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(~m[832]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[832]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[832]&m[1198]&~m[1200]&~m[1201]&m[1202])|(m[832]&~m[1198]&m[1200]&~m[1201]&m[1202])|(~m[832]&~m[1198]&~m[1200]&m[1201]&m[1202])|(m[832]&~m[1198]&~m[1200]&m[1201]&m[1202])|(~m[832]&m[1198]&~m[1200]&m[1201]&m[1202])|(m[832]&m[1198]&~m[1200]&m[1201]&m[1202])|(~m[832]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[832]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[832]&m[1198]&m[1200]&m[1201]&m[1202]))):InitCond[1445];
    m[1204] = run?((((m[698]&~m[1203]&~m[1205]&~m[1206]&~m[1207])|(~m[698]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(m[698]&m[1203]&~m[1205]&m[1206]&~m[1207])|(m[698]&~m[1203]&m[1205]&m[1206]&~m[1207])|(~m[698]&m[1203]&~m[1205]&~m[1206]&m[1207])|(~m[698]&~m[1203]&m[1205]&~m[1206]&m[1207])|(m[698]&m[1203]&m[1205]&~m[1206]&m[1207])|(~m[698]&m[1203]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[551])|((m[698]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(~m[698]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[698]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[698]&m[1203]&~m[1205]&~m[1206]&m[1207])|(m[698]&~m[1203]&m[1205]&~m[1206]&m[1207])|(~m[698]&~m[1203]&~m[1205]&m[1206]&m[1207])|(m[698]&~m[1203]&~m[1205]&m[1206]&m[1207])|(~m[698]&m[1203]&~m[1205]&m[1206]&m[1207])|(m[698]&m[1203]&~m[1205]&m[1206]&m[1207])|(~m[698]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[698]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[698]&m[1203]&m[1205]&m[1206]&m[1207]))):InitCond[1446];
    m[1209] = run?((((m[713]&~m[1208]&~m[1210]&~m[1211]&~m[1212])|(~m[713]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(m[713]&m[1208]&~m[1210]&m[1211]&~m[1212])|(m[713]&~m[1208]&m[1210]&m[1211]&~m[1212])|(~m[713]&m[1208]&~m[1210]&~m[1211]&m[1212])|(~m[713]&~m[1208]&m[1210]&~m[1211]&m[1212])|(m[713]&m[1208]&m[1210]&~m[1211]&m[1212])|(~m[713]&m[1208]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[552])|((m[713]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(~m[713]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[713]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[713]&m[1208]&~m[1210]&~m[1211]&m[1212])|(m[713]&~m[1208]&m[1210]&~m[1211]&m[1212])|(~m[713]&~m[1208]&~m[1210]&m[1211]&m[1212])|(m[713]&~m[1208]&~m[1210]&m[1211]&m[1212])|(~m[713]&m[1208]&~m[1210]&m[1211]&m[1212])|(m[713]&m[1208]&~m[1210]&m[1211]&m[1212])|(~m[713]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[713]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[713]&m[1208]&m[1210]&m[1211]&m[1212]))):InitCond[1447];
    m[1214] = run?((((m[728]&~m[1213]&~m[1215]&~m[1216]&~m[1217])|(~m[728]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(m[728]&m[1213]&~m[1215]&m[1216]&~m[1217])|(m[728]&~m[1213]&m[1215]&m[1216]&~m[1217])|(~m[728]&m[1213]&~m[1215]&~m[1216]&m[1217])|(~m[728]&~m[1213]&m[1215]&~m[1216]&m[1217])|(m[728]&m[1213]&m[1215]&~m[1216]&m[1217])|(~m[728]&m[1213]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[553])|((m[728]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(~m[728]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[728]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[728]&m[1213]&~m[1215]&~m[1216]&m[1217])|(m[728]&~m[1213]&m[1215]&~m[1216]&m[1217])|(~m[728]&~m[1213]&~m[1215]&m[1216]&m[1217])|(m[728]&~m[1213]&~m[1215]&m[1216]&m[1217])|(~m[728]&m[1213]&~m[1215]&m[1216]&m[1217])|(m[728]&m[1213]&~m[1215]&m[1216]&m[1217])|(~m[728]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[728]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[728]&m[1213]&m[1215]&m[1216]&m[1217]))):InitCond[1448];
    m[1219] = run?((((m[743]&~m[1218]&~m[1220]&~m[1221]&~m[1222])|(~m[743]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(m[743]&m[1218]&~m[1220]&m[1221]&~m[1222])|(m[743]&~m[1218]&m[1220]&m[1221]&~m[1222])|(~m[743]&m[1218]&~m[1220]&~m[1221]&m[1222])|(~m[743]&~m[1218]&m[1220]&~m[1221]&m[1222])|(m[743]&m[1218]&m[1220]&~m[1221]&m[1222])|(~m[743]&m[1218]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[554])|((m[743]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(~m[743]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[743]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[743]&m[1218]&~m[1220]&~m[1221]&m[1222])|(m[743]&~m[1218]&m[1220]&~m[1221]&m[1222])|(~m[743]&~m[1218]&~m[1220]&m[1221]&m[1222])|(m[743]&~m[1218]&~m[1220]&m[1221]&m[1222])|(~m[743]&m[1218]&~m[1220]&m[1221]&m[1222])|(m[743]&m[1218]&~m[1220]&m[1221]&m[1222])|(~m[743]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[743]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[743]&m[1218]&m[1220]&m[1221]&m[1222]))):InitCond[1449];
    m[1224] = run?((((m[758]&~m[1223]&~m[1225]&~m[1226]&~m[1227])|(~m[758]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(m[758]&m[1223]&~m[1225]&m[1226]&~m[1227])|(m[758]&~m[1223]&m[1225]&m[1226]&~m[1227])|(~m[758]&m[1223]&~m[1225]&~m[1226]&m[1227])|(~m[758]&~m[1223]&m[1225]&~m[1226]&m[1227])|(m[758]&m[1223]&m[1225]&~m[1226]&m[1227])|(~m[758]&m[1223]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[555])|((m[758]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(~m[758]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[758]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[758]&m[1223]&~m[1225]&~m[1226]&m[1227])|(m[758]&~m[1223]&m[1225]&~m[1226]&m[1227])|(~m[758]&~m[1223]&~m[1225]&m[1226]&m[1227])|(m[758]&~m[1223]&~m[1225]&m[1226]&m[1227])|(~m[758]&m[1223]&~m[1225]&m[1226]&m[1227])|(m[758]&m[1223]&~m[1225]&m[1226]&m[1227])|(~m[758]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[758]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[758]&m[1223]&m[1225]&m[1226]&m[1227]))):InitCond[1450];
    m[1229] = run?((((m[773]&~m[1228]&~m[1230]&~m[1231]&~m[1232])|(~m[773]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(m[773]&m[1228]&~m[1230]&m[1231]&~m[1232])|(m[773]&~m[1228]&m[1230]&m[1231]&~m[1232])|(~m[773]&m[1228]&~m[1230]&~m[1231]&m[1232])|(~m[773]&~m[1228]&m[1230]&~m[1231]&m[1232])|(m[773]&m[1228]&m[1230]&~m[1231]&m[1232])|(~m[773]&m[1228]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[556])|((m[773]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(~m[773]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[773]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[773]&m[1228]&~m[1230]&~m[1231]&m[1232])|(m[773]&~m[1228]&m[1230]&~m[1231]&m[1232])|(~m[773]&~m[1228]&~m[1230]&m[1231]&m[1232])|(m[773]&~m[1228]&~m[1230]&m[1231]&m[1232])|(~m[773]&m[1228]&~m[1230]&m[1231]&m[1232])|(m[773]&m[1228]&~m[1230]&m[1231]&m[1232])|(~m[773]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[773]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[773]&m[1228]&m[1230]&m[1231]&m[1232]))):InitCond[1451];
    m[1234] = run?((((m[788]&~m[1233]&~m[1235]&~m[1236]&~m[1237])|(~m[788]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(m[788]&m[1233]&~m[1235]&m[1236]&~m[1237])|(m[788]&~m[1233]&m[1235]&m[1236]&~m[1237])|(~m[788]&m[1233]&~m[1235]&~m[1236]&m[1237])|(~m[788]&~m[1233]&m[1235]&~m[1236]&m[1237])|(m[788]&m[1233]&m[1235]&~m[1236]&m[1237])|(~m[788]&m[1233]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[557])|((m[788]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(~m[788]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[788]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[788]&m[1233]&~m[1235]&~m[1236]&m[1237])|(m[788]&~m[1233]&m[1235]&~m[1236]&m[1237])|(~m[788]&~m[1233]&~m[1235]&m[1236]&m[1237])|(m[788]&~m[1233]&~m[1235]&m[1236]&m[1237])|(~m[788]&m[1233]&~m[1235]&m[1236]&m[1237])|(m[788]&m[1233]&~m[1235]&m[1236]&m[1237])|(~m[788]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[788]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[788]&m[1233]&m[1235]&m[1236]&m[1237]))):InitCond[1452];
    m[1239] = run?((((m[803]&~m[1238]&~m[1240]&~m[1241]&~m[1242])|(~m[803]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(m[803]&m[1238]&~m[1240]&m[1241]&~m[1242])|(m[803]&~m[1238]&m[1240]&m[1241]&~m[1242])|(~m[803]&m[1238]&~m[1240]&~m[1241]&m[1242])|(~m[803]&~m[1238]&m[1240]&~m[1241]&m[1242])|(m[803]&m[1238]&m[1240]&~m[1241]&m[1242])|(~m[803]&m[1238]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[558])|((m[803]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(~m[803]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[803]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[803]&m[1238]&~m[1240]&~m[1241]&m[1242])|(m[803]&~m[1238]&m[1240]&~m[1241]&m[1242])|(~m[803]&~m[1238]&~m[1240]&m[1241]&m[1242])|(m[803]&~m[1238]&~m[1240]&m[1241]&m[1242])|(~m[803]&m[1238]&~m[1240]&m[1241]&m[1242])|(m[803]&m[1238]&~m[1240]&m[1241]&m[1242])|(~m[803]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[803]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[803]&m[1238]&m[1240]&m[1241]&m[1242]))):InitCond[1453];
    m[1244] = run?((((m[818]&~m[1243]&~m[1245]&~m[1246]&~m[1247])|(~m[818]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(m[818]&m[1243]&~m[1245]&m[1246]&~m[1247])|(m[818]&~m[1243]&m[1245]&m[1246]&~m[1247])|(~m[818]&m[1243]&~m[1245]&~m[1246]&m[1247])|(~m[818]&~m[1243]&m[1245]&~m[1246]&m[1247])|(m[818]&m[1243]&m[1245]&~m[1246]&m[1247])|(~m[818]&m[1243]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[559])|((m[818]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(~m[818]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[818]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[818]&m[1243]&~m[1245]&~m[1246]&m[1247])|(m[818]&~m[1243]&m[1245]&~m[1246]&m[1247])|(~m[818]&~m[1243]&~m[1245]&m[1246]&m[1247])|(m[818]&~m[1243]&~m[1245]&m[1246]&m[1247])|(~m[818]&m[1243]&~m[1245]&m[1246]&m[1247])|(m[818]&m[1243]&~m[1245]&m[1246]&m[1247])|(~m[818]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[818]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[818]&m[1243]&m[1245]&m[1246]&m[1247]))):InitCond[1454];
    m[1249] = run?((((m[833]&~m[1248]&~m[1250]&~m[1251]&~m[1252])|(~m[833]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(m[833]&m[1248]&~m[1250]&m[1251]&~m[1252])|(m[833]&~m[1248]&m[1250]&m[1251]&~m[1252])|(~m[833]&m[1248]&~m[1250]&~m[1251]&m[1252])|(~m[833]&~m[1248]&m[1250]&~m[1251]&m[1252])|(m[833]&m[1248]&m[1250]&~m[1251]&m[1252])|(~m[833]&m[1248]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[560])|((m[833]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(~m[833]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[833]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[833]&m[1248]&~m[1250]&~m[1251]&m[1252])|(m[833]&~m[1248]&m[1250]&~m[1251]&m[1252])|(~m[833]&~m[1248]&~m[1250]&m[1251]&m[1252])|(m[833]&~m[1248]&~m[1250]&m[1251]&m[1252])|(~m[833]&m[1248]&~m[1250]&m[1251]&m[1252])|(m[833]&m[1248]&~m[1250]&m[1251]&m[1252])|(~m[833]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[833]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[833]&m[1248]&m[1250]&m[1251]&m[1252]))):InitCond[1455];
    m[1254] = run?((((m[848]&~m[1253]&~m[1255]&~m[1256]&~m[1257])|(~m[848]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(m[848]&m[1253]&~m[1255]&m[1256]&~m[1257])|(m[848]&~m[1253]&m[1255]&m[1256]&~m[1257])|(~m[848]&m[1253]&~m[1255]&~m[1256]&m[1257])|(~m[848]&~m[1253]&m[1255]&~m[1256]&m[1257])|(m[848]&m[1253]&m[1255]&~m[1256]&m[1257])|(~m[848]&m[1253]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[561])|((m[848]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(~m[848]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[848]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[848]&m[1253]&~m[1255]&~m[1256]&m[1257])|(m[848]&~m[1253]&m[1255]&~m[1256]&m[1257])|(~m[848]&~m[1253]&~m[1255]&m[1256]&m[1257])|(m[848]&~m[1253]&~m[1255]&m[1256]&m[1257])|(~m[848]&m[1253]&~m[1255]&m[1256]&m[1257])|(m[848]&m[1253]&~m[1255]&m[1256]&m[1257])|(~m[848]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[848]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[848]&m[1253]&m[1255]&m[1256]&m[1257]))):InitCond[1456];
    m[1259] = run?((((m[699]&~m[1258]&~m[1260]&~m[1261]&~m[1262])|(~m[699]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(m[699]&m[1258]&~m[1260]&m[1261]&~m[1262])|(m[699]&~m[1258]&m[1260]&m[1261]&~m[1262])|(~m[699]&m[1258]&~m[1260]&~m[1261]&m[1262])|(~m[699]&~m[1258]&m[1260]&~m[1261]&m[1262])|(m[699]&m[1258]&m[1260]&~m[1261]&m[1262])|(~m[699]&m[1258]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[562])|((m[699]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(~m[699]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[699]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[699]&m[1258]&~m[1260]&~m[1261]&m[1262])|(m[699]&~m[1258]&m[1260]&~m[1261]&m[1262])|(~m[699]&~m[1258]&~m[1260]&m[1261]&m[1262])|(m[699]&~m[1258]&~m[1260]&m[1261]&m[1262])|(~m[699]&m[1258]&~m[1260]&m[1261]&m[1262])|(m[699]&m[1258]&~m[1260]&m[1261]&m[1262])|(~m[699]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[699]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[699]&m[1258]&m[1260]&m[1261]&m[1262]))):InitCond[1457];
    m[1264] = run?((((m[714]&~m[1263]&~m[1265]&~m[1266]&~m[1267])|(~m[714]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(m[714]&m[1263]&~m[1265]&m[1266]&~m[1267])|(m[714]&~m[1263]&m[1265]&m[1266]&~m[1267])|(~m[714]&m[1263]&~m[1265]&~m[1266]&m[1267])|(~m[714]&~m[1263]&m[1265]&~m[1266]&m[1267])|(m[714]&m[1263]&m[1265]&~m[1266]&m[1267])|(~m[714]&m[1263]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[563])|((m[714]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(~m[714]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[714]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[714]&m[1263]&~m[1265]&~m[1266]&m[1267])|(m[714]&~m[1263]&m[1265]&~m[1266]&m[1267])|(~m[714]&~m[1263]&~m[1265]&m[1266]&m[1267])|(m[714]&~m[1263]&~m[1265]&m[1266]&m[1267])|(~m[714]&m[1263]&~m[1265]&m[1266]&m[1267])|(m[714]&m[1263]&~m[1265]&m[1266]&m[1267])|(~m[714]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[714]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[714]&m[1263]&m[1265]&m[1266]&m[1267]))):InitCond[1458];
    m[1269] = run?((((m[729]&~m[1268]&~m[1270]&~m[1271]&~m[1272])|(~m[729]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(m[729]&m[1268]&~m[1270]&m[1271]&~m[1272])|(m[729]&~m[1268]&m[1270]&m[1271]&~m[1272])|(~m[729]&m[1268]&~m[1270]&~m[1271]&m[1272])|(~m[729]&~m[1268]&m[1270]&~m[1271]&m[1272])|(m[729]&m[1268]&m[1270]&~m[1271]&m[1272])|(~m[729]&m[1268]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[564])|((m[729]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(~m[729]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[729]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[729]&m[1268]&~m[1270]&~m[1271]&m[1272])|(m[729]&~m[1268]&m[1270]&~m[1271]&m[1272])|(~m[729]&~m[1268]&~m[1270]&m[1271]&m[1272])|(m[729]&~m[1268]&~m[1270]&m[1271]&m[1272])|(~m[729]&m[1268]&~m[1270]&m[1271]&m[1272])|(m[729]&m[1268]&~m[1270]&m[1271]&m[1272])|(~m[729]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[729]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[729]&m[1268]&m[1270]&m[1271]&m[1272]))):InitCond[1459];
    m[1274] = run?((((m[744]&~m[1273]&~m[1275]&~m[1276]&~m[1277])|(~m[744]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(m[744]&m[1273]&~m[1275]&m[1276]&~m[1277])|(m[744]&~m[1273]&m[1275]&m[1276]&~m[1277])|(~m[744]&m[1273]&~m[1275]&~m[1276]&m[1277])|(~m[744]&~m[1273]&m[1275]&~m[1276]&m[1277])|(m[744]&m[1273]&m[1275]&~m[1276]&m[1277])|(~m[744]&m[1273]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[565])|((m[744]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(~m[744]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[744]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[744]&m[1273]&~m[1275]&~m[1276]&m[1277])|(m[744]&~m[1273]&m[1275]&~m[1276]&m[1277])|(~m[744]&~m[1273]&~m[1275]&m[1276]&m[1277])|(m[744]&~m[1273]&~m[1275]&m[1276]&m[1277])|(~m[744]&m[1273]&~m[1275]&m[1276]&m[1277])|(m[744]&m[1273]&~m[1275]&m[1276]&m[1277])|(~m[744]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[744]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[744]&m[1273]&m[1275]&m[1276]&m[1277]))):InitCond[1460];
    m[1279] = run?((((m[759]&~m[1278]&~m[1280]&~m[1281]&~m[1282])|(~m[759]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(m[759]&m[1278]&~m[1280]&m[1281]&~m[1282])|(m[759]&~m[1278]&m[1280]&m[1281]&~m[1282])|(~m[759]&m[1278]&~m[1280]&~m[1281]&m[1282])|(~m[759]&~m[1278]&m[1280]&~m[1281]&m[1282])|(m[759]&m[1278]&m[1280]&~m[1281]&m[1282])|(~m[759]&m[1278]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[566])|((m[759]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(~m[759]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[759]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[759]&m[1278]&~m[1280]&~m[1281]&m[1282])|(m[759]&~m[1278]&m[1280]&~m[1281]&m[1282])|(~m[759]&~m[1278]&~m[1280]&m[1281]&m[1282])|(m[759]&~m[1278]&~m[1280]&m[1281]&m[1282])|(~m[759]&m[1278]&~m[1280]&m[1281]&m[1282])|(m[759]&m[1278]&~m[1280]&m[1281]&m[1282])|(~m[759]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[759]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[759]&m[1278]&m[1280]&m[1281]&m[1282]))):InitCond[1461];
    m[1284] = run?((((m[774]&~m[1283]&~m[1285]&~m[1286]&~m[1287])|(~m[774]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(m[774]&m[1283]&~m[1285]&m[1286]&~m[1287])|(m[774]&~m[1283]&m[1285]&m[1286]&~m[1287])|(~m[774]&m[1283]&~m[1285]&~m[1286]&m[1287])|(~m[774]&~m[1283]&m[1285]&~m[1286]&m[1287])|(m[774]&m[1283]&m[1285]&~m[1286]&m[1287])|(~m[774]&m[1283]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[567])|((m[774]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(~m[774]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[774]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[774]&m[1283]&~m[1285]&~m[1286]&m[1287])|(m[774]&~m[1283]&m[1285]&~m[1286]&m[1287])|(~m[774]&~m[1283]&~m[1285]&m[1286]&m[1287])|(m[774]&~m[1283]&~m[1285]&m[1286]&m[1287])|(~m[774]&m[1283]&~m[1285]&m[1286]&m[1287])|(m[774]&m[1283]&~m[1285]&m[1286]&m[1287])|(~m[774]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[774]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[774]&m[1283]&m[1285]&m[1286]&m[1287]))):InitCond[1462];
    m[1289] = run?((((m[789]&~m[1288]&~m[1290]&~m[1291]&~m[1292])|(~m[789]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(m[789]&m[1288]&~m[1290]&m[1291]&~m[1292])|(m[789]&~m[1288]&m[1290]&m[1291]&~m[1292])|(~m[789]&m[1288]&~m[1290]&~m[1291]&m[1292])|(~m[789]&~m[1288]&m[1290]&~m[1291]&m[1292])|(m[789]&m[1288]&m[1290]&~m[1291]&m[1292])|(~m[789]&m[1288]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[568])|((m[789]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(~m[789]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[789]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[789]&m[1288]&~m[1290]&~m[1291]&m[1292])|(m[789]&~m[1288]&m[1290]&~m[1291]&m[1292])|(~m[789]&~m[1288]&~m[1290]&m[1291]&m[1292])|(m[789]&~m[1288]&~m[1290]&m[1291]&m[1292])|(~m[789]&m[1288]&~m[1290]&m[1291]&m[1292])|(m[789]&m[1288]&~m[1290]&m[1291]&m[1292])|(~m[789]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[789]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[789]&m[1288]&m[1290]&m[1291]&m[1292]))):InitCond[1463];
    m[1294] = run?((((m[804]&~m[1293]&~m[1295]&~m[1296]&~m[1297])|(~m[804]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(m[804]&m[1293]&~m[1295]&m[1296]&~m[1297])|(m[804]&~m[1293]&m[1295]&m[1296]&~m[1297])|(~m[804]&m[1293]&~m[1295]&~m[1296]&m[1297])|(~m[804]&~m[1293]&m[1295]&~m[1296]&m[1297])|(m[804]&m[1293]&m[1295]&~m[1296]&m[1297])|(~m[804]&m[1293]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[569])|((m[804]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(~m[804]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[804]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[804]&m[1293]&~m[1295]&~m[1296]&m[1297])|(m[804]&~m[1293]&m[1295]&~m[1296]&m[1297])|(~m[804]&~m[1293]&~m[1295]&m[1296]&m[1297])|(m[804]&~m[1293]&~m[1295]&m[1296]&m[1297])|(~m[804]&m[1293]&~m[1295]&m[1296]&m[1297])|(m[804]&m[1293]&~m[1295]&m[1296]&m[1297])|(~m[804]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[804]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[804]&m[1293]&m[1295]&m[1296]&m[1297]))):InitCond[1464];
    m[1299] = run?((((m[819]&~m[1298]&~m[1300]&~m[1301]&~m[1302])|(~m[819]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(m[819]&m[1298]&~m[1300]&m[1301]&~m[1302])|(m[819]&~m[1298]&m[1300]&m[1301]&~m[1302])|(~m[819]&m[1298]&~m[1300]&~m[1301]&m[1302])|(~m[819]&~m[1298]&m[1300]&~m[1301]&m[1302])|(m[819]&m[1298]&m[1300]&~m[1301]&m[1302])|(~m[819]&m[1298]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[570])|((m[819]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(~m[819]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[819]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[819]&m[1298]&~m[1300]&~m[1301]&m[1302])|(m[819]&~m[1298]&m[1300]&~m[1301]&m[1302])|(~m[819]&~m[1298]&~m[1300]&m[1301]&m[1302])|(m[819]&~m[1298]&~m[1300]&m[1301]&m[1302])|(~m[819]&m[1298]&~m[1300]&m[1301]&m[1302])|(m[819]&m[1298]&~m[1300]&m[1301]&m[1302])|(~m[819]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[819]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[819]&m[1298]&m[1300]&m[1301]&m[1302]))):InitCond[1465];
    m[1304] = run?((((m[834]&~m[1303]&~m[1305]&~m[1306]&~m[1307])|(~m[834]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(m[834]&m[1303]&~m[1305]&m[1306]&~m[1307])|(m[834]&~m[1303]&m[1305]&m[1306]&~m[1307])|(~m[834]&m[1303]&~m[1305]&~m[1306]&m[1307])|(~m[834]&~m[1303]&m[1305]&~m[1306]&m[1307])|(m[834]&m[1303]&m[1305]&~m[1306]&m[1307])|(~m[834]&m[1303]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[571])|((m[834]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(~m[834]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[834]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[834]&m[1303]&~m[1305]&~m[1306]&m[1307])|(m[834]&~m[1303]&m[1305]&~m[1306]&m[1307])|(~m[834]&~m[1303]&~m[1305]&m[1306]&m[1307])|(m[834]&~m[1303]&~m[1305]&m[1306]&m[1307])|(~m[834]&m[1303]&~m[1305]&m[1306]&m[1307])|(m[834]&m[1303]&~m[1305]&m[1306]&m[1307])|(~m[834]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[834]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[834]&m[1303]&m[1305]&m[1306]&m[1307]))):InitCond[1466];
    m[1309] = run?((((m[849]&~m[1308]&~m[1310]&~m[1311]&~m[1312])|(~m[849]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(m[849]&m[1308]&~m[1310]&m[1311]&~m[1312])|(m[849]&~m[1308]&m[1310]&m[1311]&~m[1312])|(~m[849]&m[1308]&~m[1310]&~m[1311]&m[1312])|(~m[849]&~m[1308]&m[1310]&~m[1311]&m[1312])|(m[849]&m[1308]&m[1310]&~m[1311]&m[1312])|(~m[849]&m[1308]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[572])|((m[849]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(~m[849]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[849]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[849]&m[1308]&~m[1310]&~m[1311]&m[1312])|(m[849]&~m[1308]&m[1310]&~m[1311]&m[1312])|(~m[849]&~m[1308]&~m[1310]&m[1311]&m[1312])|(m[849]&~m[1308]&~m[1310]&m[1311]&m[1312])|(~m[849]&m[1308]&~m[1310]&m[1311]&m[1312])|(m[849]&m[1308]&~m[1310]&m[1311]&m[1312])|(~m[849]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[849]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[849]&m[1308]&m[1310]&m[1311]&m[1312]))):InitCond[1467];
    m[1314] = run?((((m[864]&~m[1313]&~m[1315]&~m[1316]&~m[1317])|(~m[864]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(m[864]&m[1313]&~m[1315]&m[1316]&~m[1317])|(m[864]&~m[1313]&m[1315]&m[1316]&~m[1317])|(~m[864]&m[1313]&~m[1315]&~m[1316]&m[1317])|(~m[864]&~m[1313]&m[1315]&~m[1316]&m[1317])|(m[864]&m[1313]&m[1315]&~m[1316]&m[1317])|(~m[864]&m[1313]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[573])|((m[864]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(~m[864]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[864]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[864]&m[1313]&~m[1315]&~m[1316]&m[1317])|(m[864]&~m[1313]&m[1315]&~m[1316]&m[1317])|(~m[864]&~m[1313]&~m[1315]&m[1316]&m[1317])|(m[864]&~m[1313]&~m[1315]&m[1316]&m[1317])|(~m[864]&m[1313]&~m[1315]&m[1316]&m[1317])|(m[864]&m[1313]&~m[1315]&m[1316]&m[1317])|(~m[864]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[864]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[864]&m[1313]&m[1315]&m[1316]&m[1317]))):InitCond[1468];
    m[1319] = run?((((m[700]&~m[1318]&~m[1320]&~m[1321]&~m[1322])|(~m[700]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(m[700]&m[1318]&~m[1320]&m[1321]&~m[1322])|(m[700]&~m[1318]&m[1320]&m[1321]&~m[1322])|(~m[700]&m[1318]&~m[1320]&~m[1321]&m[1322])|(~m[700]&~m[1318]&m[1320]&~m[1321]&m[1322])|(m[700]&m[1318]&m[1320]&~m[1321]&m[1322])|(~m[700]&m[1318]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[574])|((m[700]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(~m[700]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[700]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[700]&m[1318]&~m[1320]&~m[1321]&m[1322])|(m[700]&~m[1318]&m[1320]&~m[1321]&m[1322])|(~m[700]&~m[1318]&~m[1320]&m[1321]&m[1322])|(m[700]&~m[1318]&~m[1320]&m[1321]&m[1322])|(~m[700]&m[1318]&~m[1320]&m[1321]&m[1322])|(m[700]&m[1318]&~m[1320]&m[1321]&m[1322])|(~m[700]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[700]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[700]&m[1318]&m[1320]&m[1321]&m[1322]))):InitCond[1469];
    m[1324] = run?((((m[715]&~m[1323]&~m[1325]&~m[1326]&~m[1327])|(~m[715]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(m[715]&m[1323]&~m[1325]&m[1326]&~m[1327])|(m[715]&~m[1323]&m[1325]&m[1326]&~m[1327])|(~m[715]&m[1323]&~m[1325]&~m[1326]&m[1327])|(~m[715]&~m[1323]&m[1325]&~m[1326]&m[1327])|(m[715]&m[1323]&m[1325]&~m[1326]&m[1327])|(~m[715]&m[1323]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[575])|((m[715]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(~m[715]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[715]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[715]&m[1323]&~m[1325]&~m[1326]&m[1327])|(m[715]&~m[1323]&m[1325]&~m[1326]&m[1327])|(~m[715]&~m[1323]&~m[1325]&m[1326]&m[1327])|(m[715]&~m[1323]&~m[1325]&m[1326]&m[1327])|(~m[715]&m[1323]&~m[1325]&m[1326]&m[1327])|(m[715]&m[1323]&~m[1325]&m[1326]&m[1327])|(~m[715]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[715]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[715]&m[1323]&m[1325]&m[1326]&m[1327]))):InitCond[1470];
    m[1329] = run?((((m[730]&~m[1328]&~m[1330]&~m[1331]&~m[1332])|(~m[730]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(m[730]&m[1328]&~m[1330]&m[1331]&~m[1332])|(m[730]&~m[1328]&m[1330]&m[1331]&~m[1332])|(~m[730]&m[1328]&~m[1330]&~m[1331]&m[1332])|(~m[730]&~m[1328]&m[1330]&~m[1331]&m[1332])|(m[730]&m[1328]&m[1330]&~m[1331]&m[1332])|(~m[730]&m[1328]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[576])|((m[730]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(~m[730]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[730]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[730]&m[1328]&~m[1330]&~m[1331]&m[1332])|(m[730]&~m[1328]&m[1330]&~m[1331]&m[1332])|(~m[730]&~m[1328]&~m[1330]&m[1331]&m[1332])|(m[730]&~m[1328]&~m[1330]&m[1331]&m[1332])|(~m[730]&m[1328]&~m[1330]&m[1331]&m[1332])|(m[730]&m[1328]&~m[1330]&m[1331]&m[1332])|(~m[730]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[730]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[730]&m[1328]&m[1330]&m[1331]&m[1332]))):InitCond[1471];
    m[1334] = run?((((m[745]&~m[1333]&~m[1335]&~m[1336]&~m[1337])|(~m[745]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(m[745]&m[1333]&~m[1335]&m[1336]&~m[1337])|(m[745]&~m[1333]&m[1335]&m[1336]&~m[1337])|(~m[745]&m[1333]&~m[1335]&~m[1336]&m[1337])|(~m[745]&~m[1333]&m[1335]&~m[1336]&m[1337])|(m[745]&m[1333]&m[1335]&~m[1336]&m[1337])|(~m[745]&m[1333]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[577])|((m[745]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(~m[745]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[745]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[745]&m[1333]&~m[1335]&~m[1336]&m[1337])|(m[745]&~m[1333]&m[1335]&~m[1336]&m[1337])|(~m[745]&~m[1333]&~m[1335]&m[1336]&m[1337])|(m[745]&~m[1333]&~m[1335]&m[1336]&m[1337])|(~m[745]&m[1333]&~m[1335]&m[1336]&m[1337])|(m[745]&m[1333]&~m[1335]&m[1336]&m[1337])|(~m[745]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[745]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[745]&m[1333]&m[1335]&m[1336]&m[1337]))):InitCond[1472];
    m[1339] = run?((((m[760]&~m[1338]&~m[1340]&~m[1341]&~m[1342])|(~m[760]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(m[760]&m[1338]&~m[1340]&m[1341]&~m[1342])|(m[760]&~m[1338]&m[1340]&m[1341]&~m[1342])|(~m[760]&m[1338]&~m[1340]&~m[1341]&m[1342])|(~m[760]&~m[1338]&m[1340]&~m[1341]&m[1342])|(m[760]&m[1338]&m[1340]&~m[1341]&m[1342])|(~m[760]&m[1338]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[578])|((m[760]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(~m[760]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[760]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[760]&m[1338]&~m[1340]&~m[1341]&m[1342])|(m[760]&~m[1338]&m[1340]&~m[1341]&m[1342])|(~m[760]&~m[1338]&~m[1340]&m[1341]&m[1342])|(m[760]&~m[1338]&~m[1340]&m[1341]&m[1342])|(~m[760]&m[1338]&~m[1340]&m[1341]&m[1342])|(m[760]&m[1338]&~m[1340]&m[1341]&m[1342])|(~m[760]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[760]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[760]&m[1338]&m[1340]&m[1341]&m[1342]))):InitCond[1473];
    m[1344] = run?((((m[775]&~m[1343]&~m[1345]&~m[1346]&~m[1347])|(~m[775]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(m[775]&m[1343]&~m[1345]&m[1346]&~m[1347])|(m[775]&~m[1343]&m[1345]&m[1346]&~m[1347])|(~m[775]&m[1343]&~m[1345]&~m[1346]&m[1347])|(~m[775]&~m[1343]&m[1345]&~m[1346]&m[1347])|(m[775]&m[1343]&m[1345]&~m[1346]&m[1347])|(~m[775]&m[1343]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[579])|((m[775]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(~m[775]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[775]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[775]&m[1343]&~m[1345]&~m[1346]&m[1347])|(m[775]&~m[1343]&m[1345]&~m[1346]&m[1347])|(~m[775]&~m[1343]&~m[1345]&m[1346]&m[1347])|(m[775]&~m[1343]&~m[1345]&m[1346]&m[1347])|(~m[775]&m[1343]&~m[1345]&m[1346]&m[1347])|(m[775]&m[1343]&~m[1345]&m[1346]&m[1347])|(~m[775]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[775]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[775]&m[1343]&m[1345]&m[1346]&m[1347]))):InitCond[1474];
    m[1349] = run?((((m[790]&~m[1348]&~m[1350]&~m[1351]&~m[1352])|(~m[790]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(m[790]&m[1348]&~m[1350]&m[1351]&~m[1352])|(m[790]&~m[1348]&m[1350]&m[1351]&~m[1352])|(~m[790]&m[1348]&~m[1350]&~m[1351]&m[1352])|(~m[790]&~m[1348]&m[1350]&~m[1351]&m[1352])|(m[790]&m[1348]&m[1350]&~m[1351]&m[1352])|(~m[790]&m[1348]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[580])|((m[790]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(~m[790]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[790]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[790]&m[1348]&~m[1350]&~m[1351]&m[1352])|(m[790]&~m[1348]&m[1350]&~m[1351]&m[1352])|(~m[790]&~m[1348]&~m[1350]&m[1351]&m[1352])|(m[790]&~m[1348]&~m[1350]&m[1351]&m[1352])|(~m[790]&m[1348]&~m[1350]&m[1351]&m[1352])|(m[790]&m[1348]&~m[1350]&m[1351]&m[1352])|(~m[790]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[790]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[790]&m[1348]&m[1350]&m[1351]&m[1352]))):InitCond[1475];
    m[1354] = run?((((m[805]&~m[1353]&~m[1355]&~m[1356]&~m[1357])|(~m[805]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(m[805]&m[1353]&~m[1355]&m[1356]&~m[1357])|(m[805]&~m[1353]&m[1355]&m[1356]&~m[1357])|(~m[805]&m[1353]&~m[1355]&~m[1356]&m[1357])|(~m[805]&~m[1353]&m[1355]&~m[1356]&m[1357])|(m[805]&m[1353]&m[1355]&~m[1356]&m[1357])|(~m[805]&m[1353]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[581])|((m[805]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(~m[805]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[805]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[805]&m[1353]&~m[1355]&~m[1356]&m[1357])|(m[805]&~m[1353]&m[1355]&~m[1356]&m[1357])|(~m[805]&~m[1353]&~m[1355]&m[1356]&m[1357])|(m[805]&~m[1353]&~m[1355]&m[1356]&m[1357])|(~m[805]&m[1353]&~m[1355]&m[1356]&m[1357])|(m[805]&m[1353]&~m[1355]&m[1356]&m[1357])|(~m[805]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[805]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[805]&m[1353]&m[1355]&m[1356]&m[1357]))):InitCond[1476];
    m[1359] = run?((((m[820]&~m[1358]&~m[1360]&~m[1361]&~m[1362])|(~m[820]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(m[820]&m[1358]&~m[1360]&m[1361]&~m[1362])|(m[820]&~m[1358]&m[1360]&m[1361]&~m[1362])|(~m[820]&m[1358]&~m[1360]&~m[1361]&m[1362])|(~m[820]&~m[1358]&m[1360]&~m[1361]&m[1362])|(m[820]&m[1358]&m[1360]&~m[1361]&m[1362])|(~m[820]&m[1358]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[582])|((m[820]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(~m[820]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[820]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[820]&m[1358]&~m[1360]&~m[1361]&m[1362])|(m[820]&~m[1358]&m[1360]&~m[1361]&m[1362])|(~m[820]&~m[1358]&~m[1360]&m[1361]&m[1362])|(m[820]&~m[1358]&~m[1360]&m[1361]&m[1362])|(~m[820]&m[1358]&~m[1360]&m[1361]&m[1362])|(m[820]&m[1358]&~m[1360]&m[1361]&m[1362])|(~m[820]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[820]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[820]&m[1358]&m[1360]&m[1361]&m[1362]))):InitCond[1477];
    m[1364] = run?((((m[835]&~m[1363]&~m[1365]&~m[1366]&~m[1367])|(~m[835]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(m[835]&m[1363]&~m[1365]&m[1366]&~m[1367])|(m[835]&~m[1363]&m[1365]&m[1366]&~m[1367])|(~m[835]&m[1363]&~m[1365]&~m[1366]&m[1367])|(~m[835]&~m[1363]&m[1365]&~m[1366]&m[1367])|(m[835]&m[1363]&m[1365]&~m[1366]&m[1367])|(~m[835]&m[1363]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[583])|((m[835]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(~m[835]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[835]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[835]&m[1363]&~m[1365]&~m[1366]&m[1367])|(m[835]&~m[1363]&m[1365]&~m[1366]&m[1367])|(~m[835]&~m[1363]&~m[1365]&m[1366]&m[1367])|(m[835]&~m[1363]&~m[1365]&m[1366]&m[1367])|(~m[835]&m[1363]&~m[1365]&m[1366]&m[1367])|(m[835]&m[1363]&~m[1365]&m[1366]&m[1367])|(~m[835]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[835]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[835]&m[1363]&m[1365]&m[1366]&m[1367]))):InitCond[1478];
    m[1369] = run?((((m[850]&~m[1368]&~m[1370]&~m[1371]&~m[1372])|(~m[850]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(m[850]&m[1368]&~m[1370]&m[1371]&~m[1372])|(m[850]&~m[1368]&m[1370]&m[1371]&~m[1372])|(~m[850]&m[1368]&~m[1370]&~m[1371]&m[1372])|(~m[850]&~m[1368]&m[1370]&~m[1371]&m[1372])|(m[850]&m[1368]&m[1370]&~m[1371]&m[1372])|(~m[850]&m[1368]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[584])|((m[850]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(~m[850]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[850]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[850]&m[1368]&~m[1370]&~m[1371]&m[1372])|(m[850]&~m[1368]&m[1370]&~m[1371]&m[1372])|(~m[850]&~m[1368]&~m[1370]&m[1371]&m[1372])|(m[850]&~m[1368]&~m[1370]&m[1371]&m[1372])|(~m[850]&m[1368]&~m[1370]&m[1371]&m[1372])|(m[850]&m[1368]&~m[1370]&m[1371]&m[1372])|(~m[850]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[850]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[850]&m[1368]&m[1370]&m[1371]&m[1372]))):InitCond[1479];
    m[1374] = run?((((m[865]&~m[1373]&~m[1375]&~m[1376]&~m[1377])|(~m[865]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(m[865]&m[1373]&~m[1375]&m[1376]&~m[1377])|(m[865]&~m[1373]&m[1375]&m[1376]&~m[1377])|(~m[865]&m[1373]&~m[1375]&~m[1376]&m[1377])|(~m[865]&~m[1373]&m[1375]&~m[1376]&m[1377])|(m[865]&m[1373]&m[1375]&~m[1376]&m[1377])|(~m[865]&m[1373]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[585])|((m[865]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(~m[865]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[865]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[865]&m[1373]&~m[1375]&~m[1376]&m[1377])|(m[865]&~m[1373]&m[1375]&~m[1376]&m[1377])|(~m[865]&~m[1373]&~m[1375]&m[1376]&m[1377])|(m[865]&~m[1373]&~m[1375]&m[1376]&m[1377])|(~m[865]&m[1373]&~m[1375]&m[1376]&m[1377])|(m[865]&m[1373]&~m[1375]&m[1376]&m[1377])|(~m[865]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[865]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[865]&m[1373]&m[1375]&m[1376]&m[1377]))):InitCond[1480];
    m[1379] = run?((((m[880]&~m[1378]&~m[1380]&~m[1381]&~m[1382])|(~m[880]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(m[880]&m[1378]&~m[1380]&m[1381]&~m[1382])|(m[880]&~m[1378]&m[1380]&m[1381]&~m[1382])|(~m[880]&m[1378]&~m[1380]&~m[1381]&m[1382])|(~m[880]&~m[1378]&m[1380]&~m[1381]&m[1382])|(m[880]&m[1378]&m[1380]&~m[1381]&m[1382])|(~m[880]&m[1378]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[586])|((m[880]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(~m[880]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[880]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[880]&m[1378]&~m[1380]&~m[1381]&m[1382])|(m[880]&~m[1378]&m[1380]&~m[1381]&m[1382])|(~m[880]&~m[1378]&~m[1380]&m[1381]&m[1382])|(m[880]&~m[1378]&~m[1380]&m[1381]&m[1382])|(~m[880]&m[1378]&~m[1380]&m[1381]&m[1382])|(m[880]&m[1378]&~m[1380]&m[1381]&m[1382])|(~m[880]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[880]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[880]&m[1378]&m[1380]&m[1381]&m[1382]))):InitCond[1481];
    m[1384] = run?((((m[701]&~m[1383]&~m[1385]&~m[1386]&~m[1387])|(~m[701]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(m[701]&m[1383]&~m[1385]&m[1386]&~m[1387])|(m[701]&~m[1383]&m[1385]&m[1386]&~m[1387])|(~m[701]&m[1383]&~m[1385]&~m[1386]&m[1387])|(~m[701]&~m[1383]&m[1385]&~m[1386]&m[1387])|(m[701]&m[1383]&m[1385]&~m[1386]&m[1387])|(~m[701]&m[1383]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[587])|((m[701]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(~m[701]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[701]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[701]&m[1383]&~m[1385]&~m[1386]&m[1387])|(m[701]&~m[1383]&m[1385]&~m[1386]&m[1387])|(~m[701]&~m[1383]&~m[1385]&m[1386]&m[1387])|(m[701]&~m[1383]&~m[1385]&m[1386]&m[1387])|(~m[701]&m[1383]&~m[1385]&m[1386]&m[1387])|(m[701]&m[1383]&~m[1385]&m[1386]&m[1387])|(~m[701]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[701]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[701]&m[1383]&m[1385]&m[1386]&m[1387]))):InitCond[1482];
    m[1389] = run?((((m[716]&~m[1388]&~m[1390]&~m[1391]&~m[1392])|(~m[716]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(m[716]&m[1388]&~m[1390]&m[1391]&~m[1392])|(m[716]&~m[1388]&m[1390]&m[1391]&~m[1392])|(~m[716]&m[1388]&~m[1390]&~m[1391]&m[1392])|(~m[716]&~m[1388]&m[1390]&~m[1391]&m[1392])|(m[716]&m[1388]&m[1390]&~m[1391]&m[1392])|(~m[716]&m[1388]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[588])|((m[716]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(~m[716]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[716]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[716]&m[1388]&~m[1390]&~m[1391]&m[1392])|(m[716]&~m[1388]&m[1390]&~m[1391]&m[1392])|(~m[716]&~m[1388]&~m[1390]&m[1391]&m[1392])|(m[716]&~m[1388]&~m[1390]&m[1391]&m[1392])|(~m[716]&m[1388]&~m[1390]&m[1391]&m[1392])|(m[716]&m[1388]&~m[1390]&m[1391]&m[1392])|(~m[716]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[716]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[716]&m[1388]&m[1390]&m[1391]&m[1392]))):InitCond[1483];
    m[1394] = run?((((m[731]&~m[1393]&~m[1395]&~m[1396]&~m[1397])|(~m[731]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(m[731]&m[1393]&~m[1395]&m[1396]&~m[1397])|(m[731]&~m[1393]&m[1395]&m[1396]&~m[1397])|(~m[731]&m[1393]&~m[1395]&~m[1396]&m[1397])|(~m[731]&~m[1393]&m[1395]&~m[1396]&m[1397])|(m[731]&m[1393]&m[1395]&~m[1396]&m[1397])|(~m[731]&m[1393]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[589])|((m[731]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(~m[731]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[731]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[731]&m[1393]&~m[1395]&~m[1396]&m[1397])|(m[731]&~m[1393]&m[1395]&~m[1396]&m[1397])|(~m[731]&~m[1393]&~m[1395]&m[1396]&m[1397])|(m[731]&~m[1393]&~m[1395]&m[1396]&m[1397])|(~m[731]&m[1393]&~m[1395]&m[1396]&m[1397])|(m[731]&m[1393]&~m[1395]&m[1396]&m[1397])|(~m[731]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[731]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[731]&m[1393]&m[1395]&m[1396]&m[1397]))):InitCond[1484];
    m[1399] = run?((((m[746]&~m[1398]&~m[1400]&~m[1401]&~m[1402])|(~m[746]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(m[746]&m[1398]&~m[1400]&m[1401]&~m[1402])|(m[746]&~m[1398]&m[1400]&m[1401]&~m[1402])|(~m[746]&m[1398]&~m[1400]&~m[1401]&m[1402])|(~m[746]&~m[1398]&m[1400]&~m[1401]&m[1402])|(m[746]&m[1398]&m[1400]&~m[1401]&m[1402])|(~m[746]&m[1398]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[590])|((m[746]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(~m[746]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[746]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[746]&m[1398]&~m[1400]&~m[1401]&m[1402])|(m[746]&~m[1398]&m[1400]&~m[1401]&m[1402])|(~m[746]&~m[1398]&~m[1400]&m[1401]&m[1402])|(m[746]&~m[1398]&~m[1400]&m[1401]&m[1402])|(~m[746]&m[1398]&~m[1400]&m[1401]&m[1402])|(m[746]&m[1398]&~m[1400]&m[1401]&m[1402])|(~m[746]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[746]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[746]&m[1398]&m[1400]&m[1401]&m[1402]))):InitCond[1485];
    m[1404] = run?((((m[761]&~m[1403]&~m[1405]&~m[1406]&~m[1407])|(~m[761]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(m[761]&m[1403]&~m[1405]&m[1406]&~m[1407])|(m[761]&~m[1403]&m[1405]&m[1406]&~m[1407])|(~m[761]&m[1403]&~m[1405]&~m[1406]&m[1407])|(~m[761]&~m[1403]&m[1405]&~m[1406]&m[1407])|(m[761]&m[1403]&m[1405]&~m[1406]&m[1407])|(~m[761]&m[1403]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[591])|((m[761]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(~m[761]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[761]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[761]&m[1403]&~m[1405]&~m[1406]&m[1407])|(m[761]&~m[1403]&m[1405]&~m[1406]&m[1407])|(~m[761]&~m[1403]&~m[1405]&m[1406]&m[1407])|(m[761]&~m[1403]&~m[1405]&m[1406]&m[1407])|(~m[761]&m[1403]&~m[1405]&m[1406]&m[1407])|(m[761]&m[1403]&~m[1405]&m[1406]&m[1407])|(~m[761]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[761]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[761]&m[1403]&m[1405]&m[1406]&m[1407]))):InitCond[1486];
    m[1409] = run?((((m[776]&~m[1408]&~m[1410]&~m[1411]&~m[1412])|(~m[776]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(m[776]&m[1408]&~m[1410]&m[1411]&~m[1412])|(m[776]&~m[1408]&m[1410]&m[1411]&~m[1412])|(~m[776]&m[1408]&~m[1410]&~m[1411]&m[1412])|(~m[776]&~m[1408]&m[1410]&~m[1411]&m[1412])|(m[776]&m[1408]&m[1410]&~m[1411]&m[1412])|(~m[776]&m[1408]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[592])|((m[776]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(~m[776]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[776]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[776]&m[1408]&~m[1410]&~m[1411]&m[1412])|(m[776]&~m[1408]&m[1410]&~m[1411]&m[1412])|(~m[776]&~m[1408]&~m[1410]&m[1411]&m[1412])|(m[776]&~m[1408]&~m[1410]&m[1411]&m[1412])|(~m[776]&m[1408]&~m[1410]&m[1411]&m[1412])|(m[776]&m[1408]&~m[1410]&m[1411]&m[1412])|(~m[776]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[776]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[776]&m[1408]&m[1410]&m[1411]&m[1412]))):InitCond[1487];
    m[1414] = run?((((m[791]&~m[1413]&~m[1415]&~m[1416]&~m[1417])|(~m[791]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(m[791]&m[1413]&~m[1415]&m[1416]&~m[1417])|(m[791]&~m[1413]&m[1415]&m[1416]&~m[1417])|(~m[791]&m[1413]&~m[1415]&~m[1416]&m[1417])|(~m[791]&~m[1413]&m[1415]&~m[1416]&m[1417])|(m[791]&m[1413]&m[1415]&~m[1416]&m[1417])|(~m[791]&m[1413]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[593])|((m[791]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(~m[791]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[791]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[791]&m[1413]&~m[1415]&~m[1416]&m[1417])|(m[791]&~m[1413]&m[1415]&~m[1416]&m[1417])|(~m[791]&~m[1413]&~m[1415]&m[1416]&m[1417])|(m[791]&~m[1413]&~m[1415]&m[1416]&m[1417])|(~m[791]&m[1413]&~m[1415]&m[1416]&m[1417])|(m[791]&m[1413]&~m[1415]&m[1416]&m[1417])|(~m[791]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[791]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[791]&m[1413]&m[1415]&m[1416]&m[1417]))):InitCond[1488];
    m[1419] = run?((((m[806]&~m[1418]&~m[1420]&~m[1421]&~m[1422])|(~m[806]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(m[806]&m[1418]&~m[1420]&m[1421]&~m[1422])|(m[806]&~m[1418]&m[1420]&m[1421]&~m[1422])|(~m[806]&m[1418]&~m[1420]&~m[1421]&m[1422])|(~m[806]&~m[1418]&m[1420]&~m[1421]&m[1422])|(m[806]&m[1418]&m[1420]&~m[1421]&m[1422])|(~m[806]&m[1418]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[594])|((m[806]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(~m[806]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[806]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[806]&m[1418]&~m[1420]&~m[1421]&m[1422])|(m[806]&~m[1418]&m[1420]&~m[1421]&m[1422])|(~m[806]&~m[1418]&~m[1420]&m[1421]&m[1422])|(m[806]&~m[1418]&~m[1420]&m[1421]&m[1422])|(~m[806]&m[1418]&~m[1420]&m[1421]&m[1422])|(m[806]&m[1418]&~m[1420]&m[1421]&m[1422])|(~m[806]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[806]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[806]&m[1418]&m[1420]&m[1421]&m[1422]))):InitCond[1489];
    m[1424] = run?((((m[821]&~m[1423]&~m[1425]&~m[1426]&~m[1427])|(~m[821]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(m[821]&m[1423]&~m[1425]&m[1426]&~m[1427])|(m[821]&~m[1423]&m[1425]&m[1426]&~m[1427])|(~m[821]&m[1423]&~m[1425]&~m[1426]&m[1427])|(~m[821]&~m[1423]&m[1425]&~m[1426]&m[1427])|(m[821]&m[1423]&m[1425]&~m[1426]&m[1427])|(~m[821]&m[1423]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[595])|((m[821]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(~m[821]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[821]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[821]&m[1423]&~m[1425]&~m[1426]&m[1427])|(m[821]&~m[1423]&m[1425]&~m[1426]&m[1427])|(~m[821]&~m[1423]&~m[1425]&m[1426]&m[1427])|(m[821]&~m[1423]&~m[1425]&m[1426]&m[1427])|(~m[821]&m[1423]&~m[1425]&m[1426]&m[1427])|(m[821]&m[1423]&~m[1425]&m[1426]&m[1427])|(~m[821]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[821]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[821]&m[1423]&m[1425]&m[1426]&m[1427]))):InitCond[1490];
    m[1429] = run?((((m[836]&~m[1428]&~m[1430]&~m[1431]&~m[1432])|(~m[836]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(m[836]&m[1428]&~m[1430]&m[1431]&~m[1432])|(m[836]&~m[1428]&m[1430]&m[1431]&~m[1432])|(~m[836]&m[1428]&~m[1430]&~m[1431]&m[1432])|(~m[836]&~m[1428]&m[1430]&~m[1431]&m[1432])|(m[836]&m[1428]&m[1430]&~m[1431]&m[1432])|(~m[836]&m[1428]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[596])|((m[836]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(~m[836]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[836]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[836]&m[1428]&~m[1430]&~m[1431]&m[1432])|(m[836]&~m[1428]&m[1430]&~m[1431]&m[1432])|(~m[836]&~m[1428]&~m[1430]&m[1431]&m[1432])|(m[836]&~m[1428]&~m[1430]&m[1431]&m[1432])|(~m[836]&m[1428]&~m[1430]&m[1431]&m[1432])|(m[836]&m[1428]&~m[1430]&m[1431]&m[1432])|(~m[836]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[836]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[836]&m[1428]&m[1430]&m[1431]&m[1432]))):InitCond[1491];
    m[1434] = run?((((m[851]&~m[1433]&~m[1435]&~m[1436]&~m[1437])|(~m[851]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(m[851]&m[1433]&~m[1435]&m[1436]&~m[1437])|(m[851]&~m[1433]&m[1435]&m[1436]&~m[1437])|(~m[851]&m[1433]&~m[1435]&~m[1436]&m[1437])|(~m[851]&~m[1433]&m[1435]&~m[1436]&m[1437])|(m[851]&m[1433]&m[1435]&~m[1436]&m[1437])|(~m[851]&m[1433]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[597])|((m[851]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(~m[851]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[851]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[851]&m[1433]&~m[1435]&~m[1436]&m[1437])|(m[851]&~m[1433]&m[1435]&~m[1436]&m[1437])|(~m[851]&~m[1433]&~m[1435]&m[1436]&m[1437])|(m[851]&~m[1433]&~m[1435]&m[1436]&m[1437])|(~m[851]&m[1433]&~m[1435]&m[1436]&m[1437])|(m[851]&m[1433]&~m[1435]&m[1436]&m[1437])|(~m[851]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[851]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[851]&m[1433]&m[1435]&m[1436]&m[1437]))):InitCond[1492];
    m[1439] = run?((((m[866]&~m[1438]&~m[1440]&~m[1441]&~m[1442])|(~m[866]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(m[866]&m[1438]&~m[1440]&m[1441]&~m[1442])|(m[866]&~m[1438]&m[1440]&m[1441]&~m[1442])|(~m[866]&m[1438]&~m[1440]&~m[1441]&m[1442])|(~m[866]&~m[1438]&m[1440]&~m[1441]&m[1442])|(m[866]&m[1438]&m[1440]&~m[1441]&m[1442])|(~m[866]&m[1438]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[598])|((m[866]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(~m[866]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[866]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[866]&m[1438]&~m[1440]&~m[1441]&m[1442])|(m[866]&~m[1438]&m[1440]&~m[1441]&m[1442])|(~m[866]&~m[1438]&~m[1440]&m[1441]&m[1442])|(m[866]&~m[1438]&~m[1440]&m[1441]&m[1442])|(~m[866]&m[1438]&~m[1440]&m[1441]&m[1442])|(m[866]&m[1438]&~m[1440]&m[1441]&m[1442])|(~m[866]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[866]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[866]&m[1438]&m[1440]&m[1441]&m[1442]))):InitCond[1493];
    m[1444] = run?((((m[881]&~m[1443]&~m[1445]&~m[1446]&~m[1447])|(~m[881]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(m[881]&m[1443]&~m[1445]&m[1446]&~m[1447])|(m[881]&~m[1443]&m[1445]&m[1446]&~m[1447])|(~m[881]&m[1443]&~m[1445]&~m[1446]&m[1447])|(~m[881]&~m[1443]&m[1445]&~m[1446]&m[1447])|(m[881]&m[1443]&m[1445]&~m[1446]&m[1447])|(~m[881]&m[1443]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[599])|((m[881]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(~m[881]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[881]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[881]&m[1443]&~m[1445]&~m[1446]&m[1447])|(m[881]&~m[1443]&m[1445]&~m[1446]&m[1447])|(~m[881]&~m[1443]&~m[1445]&m[1446]&m[1447])|(m[881]&~m[1443]&~m[1445]&m[1446]&m[1447])|(~m[881]&m[1443]&~m[1445]&m[1446]&m[1447])|(m[881]&m[1443]&~m[1445]&m[1446]&m[1447])|(~m[881]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[881]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[881]&m[1443]&m[1445]&m[1446]&m[1447]))):InitCond[1494];
    m[1449] = run?((((m[896]&~m[1448]&~m[1450]&~m[1451]&~m[1452])|(~m[896]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(m[896]&m[1448]&~m[1450]&m[1451]&~m[1452])|(m[896]&~m[1448]&m[1450]&m[1451]&~m[1452])|(~m[896]&m[1448]&~m[1450]&~m[1451]&m[1452])|(~m[896]&~m[1448]&m[1450]&~m[1451]&m[1452])|(m[896]&m[1448]&m[1450]&~m[1451]&m[1452])|(~m[896]&m[1448]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[600])|((m[896]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(~m[896]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[896]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[896]&m[1448]&~m[1450]&~m[1451]&m[1452])|(m[896]&~m[1448]&m[1450]&~m[1451]&m[1452])|(~m[896]&~m[1448]&~m[1450]&m[1451]&m[1452])|(m[896]&~m[1448]&~m[1450]&m[1451]&m[1452])|(~m[896]&m[1448]&~m[1450]&m[1451]&m[1452])|(m[896]&m[1448]&~m[1450]&m[1451]&m[1452])|(~m[896]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[896]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[896]&m[1448]&m[1450]&m[1451]&m[1452]))):InitCond[1495];
    m[1454] = run?((((m[702]&~m[1453]&~m[1455]&~m[1456]&~m[1457])|(~m[702]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(m[702]&m[1453]&~m[1455]&m[1456]&~m[1457])|(m[702]&~m[1453]&m[1455]&m[1456]&~m[1457])|(~m[702]&m[1453]&~m[1455]&~m[1456]&m[1457])|(~m[702]&~m[1453]&m[1455]&~m[1456]&m[1457])|(m[702]&m[1453]&m[1455]&~m[1456]&m[1457])|(~m[702]&m[1453]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[601])|((m[702]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(~m[702]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[702]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[702]&m[1453]&~m[1455]&~m[1456]&m[1457])|(m[702]&~m[1453]&m[1455]&~m[1456]&m[1457])|(~m[702]&~m[1453]&~m[1455]&m[1456]&m[1457])|(m[702]&~m[1453]&~m[1455]&m[1456]&m[1457])|(~m[702]&m[1453]&~m[1455]&m[1456]&m[1457])|(m[702]&m[1453]&~m[1455]&m[1456]&m[1457])|(~m[702]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[702]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[702]&m[1453]&m[1455]&m[1456]&m[1457]))):InitCond[1496];
    m[1459] = run?((((m[717]&~m[1458]&~m[1460]&~m[1461]&~m[1462])|(~m[717]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(m[717]&m[1458]&~m[1460]&m[1461]&~m[1462])|(m[717]&~m[1458]&m[1460]&m[1461]&~m[1462])|(~m[717]&m[1458]&~m[1460]&~m[1461]&m[1462])|(~m[717]&~m[1458]&m[1460]&~m[1461]&m[1462])|(m[717]&m[1458]&m[1460]&~m[1461]&m[1462])|(~m[717]&m[1458]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[602])|((m[717]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(~m[717]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[717]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[717]&m[1458]&~m[1460]&~m[1461]&m[1462])|(m[717]&~m[1458]&m[1460]&~m[1461]&m[1462])|(~m[717]&~m[1458]&~m[1460]&m[1461]&m[1462])|(m[717]&~m[1458]&~m[1460]&m[1461]&m[1462])|(~m[717]&m[1458]&~m[1460]&m[1461]&m[1462])|(m[717]&m[1458]&~m[1460]&m[1461]&m[1462])|(~m[717]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[717]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[717]&m[1458]&m[1460]&m[1461]&m[1462]))):InitCond[1497];
    m[1464] = run?((((m[732]&~m[1463]&~m[1465]&~m[1466]&~m[1467])|(~m[732]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(m[732]&m[1463]&~m[1465]&m[1466]&~m[1467])|(m[732]&~m[1463]&m[1465]&m[1466]&~m[1467])|(~m[732]&m[1463]&~m[1465]&~m[1466]&m[1467])|(~m[732]&~m[1463]&m[1465]&~m[1466]&m[1467])|(m[732]&m[1463]&m[1465]&~m[1466]&m[1467])|(~m[732]&m[1463]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[603])|((m[732]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(~m[732]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[732]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[732]&m[1463]&~m[1465]&~m[1466]&m[1467])|(m[732]&~m[1463]&m[1465]&~m[1466]&m[1467])|(~m[732]&~m[1463]&~m[1465]&m[1466]&m[1467])|(m[732]&~m[1463]&~m[1465]&m[1466]&m[1467])|(~m[732]&m[1463]&~m[1465]&m[1466]&m[1467])|(m[732]&m[1463]&~m[1465]&m[1466]&m[1467])|(~m[732]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[732]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[732]&m[1463]&m[1465]&m[1466]&m[1467]))):InitCond[1498];
    m[1469] = run?((((m[747]&~m[1468]&~m[1470]&~m[1471]&~m[1472])|(~m[747]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(m[747]&m[1468]&~m[1470]&m[1471]&~m[1472])|(m[747]&~m[1468]&m[1470]&m[1471]&~m[1472])|(~m[747]&m[1468]&~m[1470]&~m[1471]&m[1472])|(~m[747]&~m[1468]&m[1470]&~m[1471]&m[1472])|(m[747]&m[1468]&m[1470]&~m[1471]&m[1472])|(~m[747]&m[1468]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[604])|((m[747]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(~m[747]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[747]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[747]&m[1468]&~m[1470]&~m[1471]&m[1472])|(m[747]&~m[1468]&m[1470]&~m[1471]&m[1472])|(~m[747]&~m[1468]&~m[1470]&m[1471]&m[1472])|(m[747]&~m[1468]&~m[1470]&m[1471]&m[1472])|(~m[747]&m[1468]&~m[1470]&m[1471]&m[1472])|(m[747]&m[1468]&~m[1470]&m[1471]&m[1472])|(~m[747]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[747]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[747]&m[1468]&m[1470]&m[1471]&m[1472]))):InitCond[1499];
    m[1474] = run?((((m[762]&~m[1473]&~m[1475]&~m[1476]&~m[1477])|(~m[762]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(m[762]&m[1473]&~m[1475]&m[1476]&~m[1477])|(m[762]&~m[1473]&m[1475]&m[1476]&~m[1477])|(~m[762]&m[1473]&~m[1475]&~m[1476]&m[1477])|(~m[762]&~m[1473]&m[1475]&~m[1476]&m[1477])|(m[762]&m[1473]&m[1475]&~m[1476]&m[1477])|(~m[762]&m[1473]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[605])|((m[762]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(~m[762]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[762]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[762]&m[1473]&~m[1475]&~m[1476]&m[1477])|(m[762]&~m[1473]&m[1475]&~m[1476]&m[1477])|(~m[762]&~m[1473]&~m[1475]&m[1476]&m[1477])|(m[762]&~m[1473]&~m[1475]&m[1476]&m[1477])|(~m[762]&m[1473]&~m[1475]&m[1476]&m[1477])|(m[762]&m[1473]&~m[1475]&m[1476]&m[1477])|(~m[762]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[762]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[762]&m[1473]&m[1475]&m[1476]&m[1477]))):InitCond[1500];
    m[1479] = run?((((m[777]&~m[1478]&~m[1480]&~m[1481]&~m[1482])|(~m[777]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(m[777]&m[1478]&~m[1480]&m[1481]&~m[1482])|(m[777]&~m[1478]&m[1480]&m[1481]&~m[1482])|(~m[777]&m[1478]&~m[1480]&~m[1481]&m[1482])|(~m[777]&~m[1478]&m[1480]&~m[1481]&m[1482])|(m[777]&m[1478]&m[1480]&~m[1481]&m[1482])|(~m[777]&m[1478]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[606])|((m[777]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(~m[777]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[777]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[777]&m[1478]&~m[1480]&~m[1481]&m[1482])|(m[777]&~m[1478]&m[1480]&~m[1481]&m[1482])|(~m[777]&~m[1478]&~m[1480]&m[1481]&m[1482])|(m[777]&~m[1478]&~m[1480]&m[1481]&m[1482])|(~m[777]&m[1478]&~m[1480]&m[1481]&m[1482])|(m[777]&m[1478]&~m[1480]&m[1481]&m[1482])|(~m[777]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[777]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[777]&m[1478]&m[1480]&m[1481]&m[1482]))):InitCond[1501];
    m[1484] = run?((((m[792]&~m[1483]&~m[1485]&~m[1486]&~m[1487])|(~m[792]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(m[792]&m[1483]&~m[1485]&m[1486]&~m[1487])|(m[792]&~m[1483]&m[1485]&m[1486]&~m[1487])|(~m[792]&m[1483]&~m[1485]&~m[1486]&m[1487])|(~m[792]&~m[1483]&m[1485]&~m[1486]&m[1487])|(m[792]&m[1483]&m[1485]&~m[1486]&m[1487])|(~m[792]&m[1483]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[607])|((m[792]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(~m[792]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[792]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[792]&m[1483]&~m[1485]&~m[1486]&m[1487])|(m[792]&~m[1483]&m[1485]&~m[1486]&m[1487])|(~m[792]&~m[1483]&~m[1485]&m[1486]&m[1487])|(m[792]&~m[1483]&~m[1485]&m[1486]&m[1487])|(~m[792]&m[1483]&~m[1485]&m[1486]&m[1487])|(m[792]&m[1483]&~m[1485]&m[1486]&m[1487])|(~m[792]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[792]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[792]&m[1483]&m[1485]&m[1486]&m[1487]))):InitCond[1502];
    m[1489] = run?((((m[807]&~m[1488]&~m[1490]&~m[1491]&~m[1492])|(~m[807]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(m[807]&m[1488]&~m[1490]&m[1491]&~m[1492])|(m[807]&~m[1488]&m[1490]&m[1491]&~m[1492])|(~m[807]&m[1488]&~m[1490]&~m[1491]&m[1492])|(~m[807]&~m[1488]&m[1490]&~m[1491]&m[1492])|(m[807]&m[1488]&m[1490]&~m[1491]&m[1492])|(~m[807]&m[1488]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[608])|((m[807]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(~m[807]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[807]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[807]&m[1488]&~m[1490]&~m[1491]&m[1492])|(m[807]&~m[1488]&m[1490]&~m[1491]&m[1492])|(~m[807]&~m[1488]&~m[1490]&m[1491]&m[1492])|(m[807]&~m[1488]&~m[1490]&m[1491]&m[1492])|(~m[807]&m[1488]&~m[1490]&m[1491]&m[1492])|(m[807]&m[1488]&~m[1490]&m[1491]&m[1492])|(~m[807]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[807]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[807]&m[1488]&m[1490]&m[1491]&m[1492]))):InitCond[1503];
    m[1494] = run?((((m[822]&~m[1493]&~m[1495]&~m[1496]&~m[1497])|(~m[822]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(m[822]&m[1493]&~m[1495]&m[1496]&~m[1497])|(m[822]&~m[1493]&m[1495]&m[1496]&~m[1497])|(~m[822]&m[1493]&~m[1495]&~m[1496]&m[1497])|(~m[822]&~m[1493]&m[1495]&~m[1496]&m[1497])|(m[822]&m[1493]&m[1495]&~m[1496]&m[1497])|(~m[822]&m[1493]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[609])|((m[822]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(~m[822]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[822]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[822]&m[1493]&~m[1495]&~m[1496]&m[1497])|(m[822]&~m[1493]&m[1495]&~m[1496]&m[1497])|(~m[822]&~m[1493]&~m[1495]&m[1496]&m[1497])|(m[822]&~m[1493]&~m[1495]&m[1496]&m[1497])|(~m[822]&m[1493]&~m[1495]&m[1496]&m[1497])|(m[822]&m[1493]&~m[1495]&m[1496]&m[1497])|(~m[822]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[822]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[822]&m[1493]&m[1495]&m[1496]&m[1497]))):InitCond[1504];
    m[1499] = run?((((m[837]&~m[1498]&~m[1500]&~m[1501]&~m[1502])|(~m[837]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(m[837]&m[1498]&~m[1500]&m[1501]&~m[1502])|(m[837]&~m[1498]&m[1500]&m[1501]&~m[1502])|(~m[837]&m[1498]&~m[1500]&~m[1501]&m[1502])|(~m[837]&~m[1498]&m[1500]&~m[1501]&m[1502])|(m[837]&m[1498]&m[1500]&~m[1501]&m[1502])|(~m[837]&m[1498]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[610])|((m[837]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(~m[837]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[837]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[837]&m[1498]&~m[1500]&~m[1501]&m[1502])|(m[837]&~m[1498]&m[1500]&~m[1501]&m[1502])|(~m[837]&~m[1498]&~m[1500]&m[1501]&m[1502])|(m[837]&~m[1498]&~m[1500]&m[1501]&m[1502])|(~m[837]&m[1498]&~m[1500]&m[1501]&m[1502])|(m[837]&m[1498]&~m[1500]&m[1501]&m[1502])|(~m[837]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[837]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[837]&m[1498]&m[1500]&m[1501]&m[1502]))):InitCond[1505];
    m[1504] = run?((((m[852]&~m[1503]&~m[1505]&~m[1506]&~m[1507])|(~m[852]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(m[852]&m[1503]&~m[1505]&m[1506]&~m[1507])|(m[852]&~m[1503]&m[1505]&m[1506]&~m[1507])|(~m[852]&m[1503]&~m[1505]&~m[1506]&m[1507])|(~m[852]&~m[1503]&m[1505]&~m[1506]&m[1507])|(m[852]&m[1503]&m[1505]&~m[1506]&m[1507])|(~m[852]&m[1503]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[611])|((m[852]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(~m[852]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[852]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[852]&m[1503]&~m[1505]&~m[1506]&m[1507])|(m[852]&~m[1503]&m[1505]&~m[1506]&m[1507])|(~m[852]&~m[1503]&~m[1505]&m[1506]&m[1507])|(m[852]&~m[1503]&~m[1505]&m[1506]&m[1507])|(~m[852]&m[1503]&~m[1505]&m[1506]&m[1507])|(m[852]&m[1503]&~m[1505]&m[1506]&m[1507])|(~m[852]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[852]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[852]&m[1503]&m[1505]&m[1506]&m[1507]))):InitCond[1506];
    m[1509] = run?((((m[867]&~m[1508]&~m[1510]&~m[1511]&~m[1512])|(~m[867]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(m[867]&m[1508]&~m[1510]&m[1511]&~m[1512])|(m[867]&~m[1508]&m[1510]&m[1511]&~m[1512])|(~m[867]&m[1508]&~m[1510]&~m[1511]&m[1512])|(~m[867]&~m[1508]&m[1510]&~m[1511]&m[1512])|(m[867]&m[1508]&m[1510]&~m[1511]&m[1512])|(~m[867]&m[1508]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[612])|((m[867]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(~m[867]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[867]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[867]&m[1508]&~m[1510]&~m[1511]&m[1512])|(m[867]&~m[1508]&m[1510]&~m[1511]&m[1512])|(~m[867]&~m[1508]&~m[1510]&m[1511]&m[1512])|(m[867]&~m[1508]&~m[1510]&m[1511]&m[1512])|(~m[867]&m[1508]&~m[1510]&m[1511]&m[1512])|(m[867]&m[1508]&~m[1510]&m[1511]&m[1512])|(~m[867]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[867]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[867]&m[1508]&m[1510]&m[1511]&m[1512]))):InitCond[1507];
    m[1514] = run?((((m[882]&~m[1513]&~m[1515]&~m[1516]&~m[1517])|(~m[882]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(m[882]&m[1513]&~m[1515]&m[1516]&~m[1517])|(m[882]&~m[1513]&m[1515]&m[1516]&~m[1517])|(~m[882]&m[1513]&~m[1515]&~m[1516]&m[1517])|(~m[882]&~m[1513]&m[1515]&~m[1516]&m[1517])|(m[882]&m[1513]&m[1515]&~m[1516]&m[1517])|(~m[882]&m[1513]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[613])|((m[882]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(~m[882]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[882]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[882]&m[1513]&~m[1515]&~m[1516]&m[1517])|(m[882]&~m[1513]&m[1515]&~m[1516]&m[1517])|(~m[882]&~m[1513]&~m[1515]&m[1516]&m[1517])|(m[882]&~m[1513]&~m[1515]&m[1516]&m[1517])|(~m[882]&m[1513]&~m[1515]&m[1516]&m[1517])|(m[882]&m[1513]&~m[1515]&m[1516]&m[1517])|(~m[882]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[882]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[882]&m[1513]&m[1515]&m[1516]&m[1517]))):InitCond[1508];
    m[1519] = run?((((m[897]&~m[1518]&~m[1520]&~m[1521]&~m[1522])|(~m[897]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(m[897]&m[1518]&~m[1520]&m[1521]&~m[1522])|(m[897]&~m[1518]&m[1520]&m[1521]&~m[1522])|(~m[897]&m[1518]&~m[1520]&~m[1521]&m[1522])|(~m[897]&~m[1518]&m[1520]&~m[1521]&m[1522])|(m[897]&m[1518]&m[1520]&~m[1521]&m[1522])|(~m[897]&m[1518]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[614])|((m[897]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(~m[897]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[897]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[897]&m[1518]&~m[1520]&~m[1521]&m[1522])|(m[897]&~m[1518]&m[1520]&~m[1521]&m[1522])|(~m[897]&~m[1518]&~m[1520]&m[1521]&m[1522])|(m[897]&~m[1518]&~m[1520]&m[1521]&m[1522])|(~m[897]&m[1518]&~m[1520]&m[1521]&m[1522])|(m[897]&m[1518]&~m[1520]&m[1521]&m[1522])|(~m[897]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[897]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[897]&m[1518]&m[1520]&m[1521]&m[1522]))):InitCond[1509];
    m[1524] = run?((((m[912]&~m[1523]&~m[1525]&~m[1526]&~m[1527])|(~m[912]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(m[912]&m[1523]&~m[1525]&m[1526]&~m[1527])|(m[912]&~m[1523]&m[1525]&m[1526]&~m[1527])|(~m[912]&m[1523]&~m[1525]&~m[1526]&m[1527])|(~m[912]&~m[1523]&m[1525]&~m[1526]&m[1527])|(m[912]&m[1523]&m[1525]&~m[1526]&m[1527])|(~m[912]&m[1523]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[615])|((m[912]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(~m[912]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[912]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[912]&m[1523]&~m[1525]&~m[1526]&m[1527])|(m[912]&~m[1523]&m[1525]&~m[1526]&m[1527])|(~m[912]&~m[1523]&~m[1525]&m[1526]&m[1527])|(m[912]&~m[1523]&~m[1525]&m[1526]&m[1527])|(~m[912]&m[1523]&~m[1525]&m[1526]&m[1527])|(m[912]&m[1523]&~m[1525]&m[1526]&m[1527])|(~m[912]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[912]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[912]&m[1523]&m[1525]&m[1526]&m[1527]))):InitCond[1510];
    m[1529] = run?((((m[703]&~m[1528]&~m[1530]&~m[1531]&~m[1532])|(~m[703]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(m[703]&m[1528]&~m[1530]&m[1531]&~m[1532])|(m[703]&~m[1528]&m[1530]&m[1531]&~m[1532])|(~m[703]&m[1528]&~m[1530]&~m[1531]&m[1532])|(~m[703]&~m[1528]&m[1530]&~m[1531]&m[1532])|(m[703]&m[1528]&m[1530]&~m[1531]&m[1532])|(~m[703]&m[1528]&m[1530]&m[1531]&m[1532]))&UnbiasedRNG[616])|((m[703]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(~m[703]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[703]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[703]&m[1528]&~m[1530]&~m[1531]&m[1532])|(m[703]&~m[1528]&m[1530]&~m[1531]&m[1532])|(~m[703]&~m[1528]&~m[1530]&m[1531]&m[1532])|(m[703]&~m[1528]&~m[1530]&m[1531]&m[1532])|(~m[703]&m[1528]&~m[1530]&m[1531]&m[1532])|(m[703]&m[1528]&~m[1530]&m[1531]&m[1532])|(~m[703]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[703]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[703]&m[1528]&m[1530]&m[1531]&m[1532]))):InitCond[1511];
    m[1534] = run?((((m[718]&~m[1533]&~m[1535]&~m[1536]&~m[1537])|(~m[718]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(m[718]&m[1533]&~m[1535]&m[1536]&~m[1537])|(m[718]&~m[1533]&m[1535]&m[1536]&~m[1537])|(~m[718]&m[1533]&~m[1535]&~m[1536]&m[1537])|(~m[718]&~m[1533]&m[1535]&~m[1536]&m[1537])|(m[718]&m[1533]&m[1535]&~m[1536]&m[1537])|(~m[718]&m[1533]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[617])|((m[718]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(~m[718]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[718]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[718]&m[1533]&~m[1535]&~m[1536]&m[1537])|(m[718]&~m[1533]&m[1535]&~m[1536]&m[1537])|(~m[718]&~m[1533]&~m[1535]&m[1536]&m[1537])|(m[718]&~m[1533]&~m[1535]&m[1536]&m[1537])|(~m[718]&m[1533]&~m[1535]&m[1536]&m[1537])|(m[718]&m[1533]&~m[1535]&m[1536]&m[1537])|(~m[718]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[718]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[718]&m[1533]&m[1535]&m[1536]&m[1537]))):InitCond[1512];
    m[1539] = run?((((m[733]&~m[1538]&~m[1540]&~m[1541]&~m[1542])|(~m[733]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(m[733]&m[1538]&~m[1540]&m[1541]&~m[1542])|(m[733]&~m[1538]&m[1540]&m[1541]&~m[1542])|(~m[733]&m[1538]&~m[1540]&~m[1541]&m[1542])|(~m[733]&~m[1538]&m[1540]&~m[1541]&m[1542])|(m[733]&m[1538]&m[1540]&~m[1541]&m[1542])|(~m[733]&m[1538]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[618])|((m[733]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(~m[733]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[733]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[733]&m[1538]&~m[1540]&~m[1541]&m[1542])|(m[733]&~m[1538]&m[1540]&~m[1541]&m[1542])|(~m[733]&~m[1538]&~m[1540]&m[1541]&m[1542])|(m[733]&~m[1538]&~m[1540]&m[1541]&m[1542])|(~m[733]&m[1538]&~m[1540]&m[1541]&m[1542])|(m[733]&m[1538]&~m[1540]&m[1541]&m[1542])|(~m[733]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[733]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[733]&m[1538]&m[1540]&m[1541]&m[1542]))):InitCond[1513];
    m[1544] = run?((((m[748]&~m[1543]&~m[1545]&~m[1546]&~m[1547])|(~m[748]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(m[748]&m[1543]&~m[1545]&m[1546]&~m[1547])|(m[748]&~m[1543]&m[1545]&m[1546]&~m[1547])|(~m[748]&m[1543]&~m[1545]&~m[1546]&m[1547])|(~m[748]&~m[1543]&m[1545]&~m[1546]&m[1547])|(m[748]&m[1543]&m[1545]&~m[1546]&m[1547])|(~m[748]&m[1543]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[619])|((m[748]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(~m[748]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[748]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[748]&m[1543]&~m[1545]&~m[1546]&m[1547])|(m[748]&~m[1543]&m[1545]&~m[1546]&m[1547])|(~m[748]&~m[1543]&~m[1545]&m[1546]&m[1547])|(m[748]&~m[1543]&~m[1545]&m[1546]&m[1547])|(~m[748]&m[1543]&~m[1545]&m[1546]&m[1547])|(m[748]&m[1543]&~m[1545]&m[1546]&m[1547])|(~m[748]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[748]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[748]&m[1543]&m[1545]&m[1546]&m[1547]))):InitCond[1514];
    m[1549] = run?((((m[763]&~m[1548]&~m[1550]&~m[1551]&~m[1552])|(~m[763]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(m[763]&m[1548]&~m[1550]&m[1551]&~m[1552])|(m[763]&~m[1548]&m[1550]&m[1551]&~m[1552])|(~m[763]&m[1548]&~m[1550]&~m[1551]&m[1552])|(~m[763]&~m[1548]&m[1550]&~m[1551]&m[1552])|(m[763]&m[1548]&m[1550]&~m[1551]&m[1552])|(~m[763]&m[1548]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[620])|((m[763]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(~m[763]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[763]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[763]&m[1548]&~m[1550]&~m[1551]&m[1552])|(m[763]&~m[1548]&m[1550]&~m[1551]&m[1552])|(~m[763]&~m[1548]&~m[1550]&m[1551]&m[1552])|(m[763]&~m[1548]&~m[1550]&m[1551]&m[1552])|(~m[763]&m[1548]&~m[1550]&m[1551]&m[1552])|(m[763]&m[1548]&~m[1550]&m[1551]&m[1552])|(~m[763]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[763]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[763]&m[1548]&m[1550]&m[1551]&m[1552]))):InitCond[1515];
    m[1554] = run?((((m[778]&~m[1553]&~m[1555]&~m[1556]&~m[1557])|(~m[778]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(m[778]&m[1553]&~m[1555]&m[1556]&~m[1557])|(m[778]&~m[1553]&m[1555]&m[1556]&~m[1557])|(~m[778]&m[1553]&~m[1555]&~m[1556]&m[1557])|(~m[778]&~m[1553]&m[1555]&~m[1556]&m[1557])|(m[778]&m[1553]&m[1555]&~m[1556]&m[1557])|(~m[778]&m[1553]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[621])|((m[778]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(~m[778]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[778]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[778]&m[1553]&~m[1555]&~m[1556]&m[1557])|(m[778]&~m[1553]&m[1555]&~m[1556]&m[1557])|(~m[778]&~m[1553]&~m[1555]&m[1556]&m[1557])|(m[778]&~m[1553]&~m[1555]&m[1556]&m[1557])|(~m[778]&m[1553]&~m[1555]&m[1556]&m[1557])|(m[778]&m[1553]&~m[1555]&m[1556]&m[1557])|(~m[778]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[778]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[778]&m[1553]&m[1555]&m[1556]&m[1557]))):InitCond[1516];
    m[1559] = run?((((m[793]&~m[1558]&~m[1560]&~m[1561]&~m[1562])|(~m[793]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(m[793]&m[1558]&~m[1560]&m[1561]&~m[1562])|(m[793]&~m[1558]&m[1560]&m[1561]&~m[1562])|(~m[793]&m[1558]&~m[1560]&~m[1561]&m[1562])|(~m[793]&~m[1558]&m[1560]&~m[1561]&m[1562])|(m[793]&m[1558]&m[1560]&~m[1561]&m[1562])|(~m[793]&m[1558]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[622])|((m[793]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(~m[793]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[793]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[793]&m[1558]&~m[1560]&~m[1561]&m[1562])|(m[793]&~m[1558]&m[1560]&~m[1561]&m[1562])|(~m[793]&~m[1558]&~m[1560]&m[1561]&m[1562])|(m[793]&~m[1558]&~m[1560]&m[1561]&m[1562])|(~m[793]&m[1558]&~m[1560]&m[1561]&m[1562])|(m[793]&m[1558]&~m[1560]&m[1561]&m[1562])|(~m[793]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[793]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[793]&m[1558]&m[1560]&m[1561]&m[1562]))):InitCond[1517];
    m[1564] = run?((((m[808]&~m[1563]&~m[1565]&~m[1566]&~m[1567])|(~m[808]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(m[808]&m[1563]&~m[1565]&m[1566]&~m[1567])|(m[808]&~m[1563]&m[1565]&m[1566]&~m[1567])|(~m[808]&m[1563]&~m[1565]&~m[1566]&m[1567])|(~m[808]&~m[1563]&m[1565]&~m[1566]&m[1567])|(m[808]&m[1563]&m[1565]&~m[1566]&m[1567])|(~m[808]&m[1563]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[623])|((m[808]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(~m[808]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[808]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[808]&m[1563]&~m[1565]&~m[1566]&m[1567])|(m[808]&~m[1563]&m[1565]&~m[1566]&m[1567])|(~m[808]&~m[1563]&~m[1565]&m[1566]&m[1567])|(m[808]&~m[1563]&~m[1565]&m[1566]&m[1567])|(~m[808]&m[1563]&~m[1565]&m[1566]&m[1567])|(m[808]&m[1563]&~m[1565]&m[1566]&m[1567])|(~m[808]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[808]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[808]&m[1563]&m[1565]&m[1566]&m[1567]))):InitCond[1518];
    m[1569] = run?((((m[823]&~m[1568]&~m[1570]&~m[1571]&~m[1572])|(~m[823]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(m[823]&m[1568]&~m[1570]&m[1571]&~m[1572])|(m[823]&~m[1568]&m[1570]&m[1571]&~m[1572])|(~m[823]&m[1568]&~m[1570]&~m[1571]&m[1572])|(~m[823]&~m[1568]&m[1570]&~m[1571]&m[1572])|(m[823]&m[1568]&m[1570]&~m[1571]&m[1572])|(~m[823]&m[1568]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[624])|((m[823]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(~m[823]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[823]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[823]&m[1568]&~m[1570]&~m[1571]&m[1572])|(m[823]&~m[1568]&m[1570]&~m[1571]&m[1572])|(~m[823]&~m[1568]&~m[1570]&m[1571]&m[1572])|(m[823]&~m[1568]&~m[1570]&m[1571]&m[1572])|(~m[823]&m[1568]&~m[1570]&m[1571]&m[1572])|(m[823]&m[1568]&~m[1570]&m[1571]&m[1572])|(~m[823]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[823]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[823]&m[1568]&m[1570]&m[1571]&m[1572]))):InitCond[1519];
    m[1574] = run?((((m[838]&~m[1573]&~m[1575]&~m[1576]&~m[1577])|(~m[838]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(m[838]&m[1573]&~m[1575]&m[1576]&~m[1577])|(m[838]&~m[1573]&m[1575]&m[1576]&~m[1577])|(~m[838]&m[1573]&~m[1575]&~m[1576]&m[1577])|(~m[838]&~m[1573]&m[1575]&~m[1576]&m[1577])|(m[838]&m[1573]&m[1575]&~m[1576]&m[1577])|(~m[838]&m[1573]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[625])|((m[838]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(~m[838]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[838]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[838]&m[1573]&~m[1575]&~m[1576]&m[1577])|(m[838]&~m[1573]&m[1575]&~m[1576]&m[1577])|(~m[838]&~m[1573]&~m[1575]&m[1576]&m[1577])|(m[838]&~m[1573]&~m[1575]&m[1576]&m[1577])|(~m[838]&m[1573]&~m[1575]&m[1576]&m[1577])|(m[838]&m[1573]&~m[1575]&m[1576]&m[1577])|(~m[838]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[838]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[838]&m[1573]&m[1575]&m[1576]&m[1577]))):InitCond[1520];
    m[1579] = run?((((m[853]&~m[1578]&~m[1580]&~m[1581]&~m[1582])|(~m[853]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(m[853]&m[1578]&~m[1580]&m[1581]&~m[1582])|(m[853]&~m[1578]&m[1580]&m[1581]&~m[1582])|(~m[853]&m[1578]&~m[1580]&~m[1581]&m[1582])|(~m[853]&~m[1578]&m[1580]&~m[1581]&m[1582])|(m[853]&m[1578]&m[1580]&~m[1581]&m[1582])|(~m[853]&m[1578]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[626])|((m[853]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(~m[853]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[853]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[853]&m[1578]&~m[1580]&~m[1581]&m[1582])|(m[853]&~m[1578]&m[1580]&~m[1581]&m[1582])|(~m[853]&~m[1578]&~m[1580]&m[1581]&m[1582])|(m[853]&~m[1578]&~m[1580]&m[1581]&m[1582])|(~m[853]&m[1578]&~m[1580]&m[1581]&m[1582])|(m[853]&m[1578]&~m[1580]&m[1581]&m[1582])|(~m[853]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[853]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[853]&m[1578]&m[1580]&m[1581]&m[1582]))):InitCond[1521];
    m[1584] = run?((((m[868]&~m[1583]&~m[1585]&~m[1586]&~m[1587])|(~m[868]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(m[868]&m[1583]&~m[1585]&m[1586]&~m[1587])|(m[868]&~m[1583]&m[1585]&m[1586]&~m[1587])|(~m[868]&m[1583]&~m[1585]&~m[1586]&m[1587])|(~m[868]&~m[1583]&m[1585]&~m[1586]&m[1587])|(m[868]&m[1583]&m[1585]&~m[1586]&m[1587])|(~m[868]&m[1583]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[627])|((m[868]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(~m[868]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[868]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[868]&m[1583]&~m[1585]&~m[1586]&m[1587])|(m[868]&~m[1583]&m[1585]&~m[1586]&m[1587])|(~m[868]&~m[1583]&~m[1585]&m[1586]&m[1587])|(m[868]&~m[1583]&~m[1585]&m[1586]&m[1587])|(~m[868]&m[1583]&~m[1585]&m[1586]&m[1587])|(m[868]&m[1583]&~m[1585]&m[1586]&m[1587])|(~m[868]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[868]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[868]&m[1583]&m[1585]&m[1586]&m[1587]))):InitCond[1522];
    m[1589] = run?((((m[883]&~m[1588]&~m[1590]&~m[1591]&~m[1592])|(~m[883]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(m[883]&m[1588]&~m[1590]&m[1591]&~m[1592])|(m[883]&~m[1588]&m[1590]&m[1591]&~m[1592])|(~m[883]&m[1588]&~m[1590]&~m[1591]&m[1592])|(~m[883]&~m[1588]&m[1590]&~m[1591]&m[1592])|(m[883]&m[1588]&m[1590]&~m[1591]&m[1592])|(~m[883]&m[1588]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[628])|((m[883]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(~m[883]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[883]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[883]&m[1588]&~m[1590]&~m[1591]&m[1592])|(m[883]&~m[1588]&m[1590]&~m[1591]&m[1592])|(~m[883]&~m[1588]&~m[1590]&m[1591]&m[1592])|(m[883]&~m[1588]&~m[1590]&m[1591]&m[1592])|(~m[883]&m[1588]&~m[1590]&m[1591]&m[1592])|(m[883]&m[1588]&~m[1590]&m[1591]&m[1592])|(~m[883]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[883]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[883]&m[1588]&m[1590]&m[1591]&m[1592]))):InitCond[1523];
    m[1594] = run?((((m[898]&~m[1593]&~m[1595]&~m[1596]&~m[1597])|(~m[898]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(m[898]&m[1593]&~m[1595]&m[1596]&~m[1597])|(m[898]&~m[1593]&m[1595]&m[1596]&~m[1597])|(~m[898]&m[1593]&~m[1595]&~m[1596]&m[1597])|(~m[898]&~m[1593]&m[1595]&~m[1596]&m[1597])|(m[898]&m[1593]&m[1595]&~m[1596]&m[1597])|(~m[898]&m[1593]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[629])|((m[898]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(~m[898]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[898]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[898]&m[1593]&~m[1595]&~m[1596]&m[1597])|(m[898]&~m[1593]&m[1595]&~m[1596]&m[1597])|(~m[898]&~m[1593]&~m[1595]&m[1596]&m[1597])|(m[898]&~m[1593]&~m[1595]&m[1596]&m[1597])|(~m[898]&m[1593]&~m[1595]&m[1596]&m[1597])|(m[898]&m[1593]&~m[1595]&m[1596]&m[1597])|(~m[898]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[898]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[898]&m[1593]&m[1595]&m[1596]&m[1597]))):InitCond[1524];
    m[1599] = run?((((m[913]&~m[1598]&~m[1600]&~m[1601]&~m[1602])|(~m[913]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(m[913]&m[1598]&~m[1600]&m[1601]&~m[1602])|(m[913]&~m[1598]&m[1600]&m[1601]&~m[1602])|(~m[913]&m[1598]&~m[1600]&~m[1601]&m[1602])|(~m[913]&~m[1598]&m[1600]&~m[1601]&m[1602])|(m[913]&m[1598]&m[1600]&~m[1601]&m[1602])|(~m[913]&m[1598]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[630])|((m[913]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(~m[913]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[913]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[913]&m[1598]&~m[1600]&~m[1601]&m[1602])|(m[913]&~m[1598]&m[1600]&~m[1601]&m[1602])|(~m[913]&~m[1598]&~m[1600]&m[1601]&m[1602])|(m[913]&~m[1598]&~m[1600]&m[1601]&m[1602])|(~m[913]&m[1598]&~m[1600]&m[1601]&m[1602])|(m[913]&m[1598]&~m[1600]&m[1601]&m[1602])|(~m[913]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[913]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[913]&m[1598]&m[1600]&m[1601]&m[1602]))):InitCond[1525];
    m[1604] = run?((((m[719]&~m[1603]&~m[1605]&~m[1606]&~m[1607])|(~m[719]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(m[719]&m[1603]&~m[1605]&m[1606]&~m[1607])|(m[719]&~m[1603]&m[1605]&m[1606]&~m[1607])|(~m[719]&m[1603]&~m[1605]&~m[1606]&m[1607])|(~m[719]&~m[1603]&m[1605]&~m[1606]&m[1607])|(m[719]&m[1603]&m[1605]&~m[1606]&m[1607])|(~m[719]&m[1603]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[631])|((m[719]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(~m[719]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[719]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[719]&m[1603]&~m[1605]&~m[1606]&m[1607])|(m[719]&~m[1603]&m[1605]&~m[1606]&m[1607])|(~m[719]&~m[1603]&~m[1605]&m[1606]&m[1607])|(m[719]&~m[1603]&~m[1605]&m[1606]&m[1607])|(~m[719]&m[1603]&~m[1605]&m[1606]&m[1607])|(m[719]&m[1603]&~m[1605]&m[1606]&m[1607])|(~m[719]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[719]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[719]&m[1603]&m[1605]&m[1606]&m[1607]))):InitCond[1526];
    m[1609] = run?((((m[734]&~m[1608]&~m[1610]&~m[1611]&~m[1612])|(~m[734]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(m[734]&m[1608]&~m[1610]&m[1611]&~m[1612])|(m[734]&~m[1608]&m[1610]&m[1611]&~m[1612])|(~m[734]&m[1608]&~m[1610]&~m[1611]&m[1612])|(~m[734]&~m[1608]&m[1610]&~m[1611]&m[1612])|(m[734]&m[1608]&m[1610]&~m[1611]&m[1612])|(~m[734]&m[1608]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[632])|((m[734]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(~m[734]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[734]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[734]&m[1608]&~m[1610]&~m[1611]&m[1612])|(m[734]&~m[1608]&m[1610]&~m[1611]&m[1612])|(~m[734]&~m[1608]&~m[1610]&m[1611]&m[1612])|(m[734]&~m[1608]&~m[1610]&m[1611]&m[1612])|(~m[734]&m[1608]&~m[1610]&m[1611]&m[1612])|(m[734]&m[1608]&~m[1610]&m[1611]&m[1612])|(~m[734]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[734]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[734]&m[1608]&m[1610]&m[1611]&m[1612]))):InitCond[1527];
    m[1614] = run?((((m[749]&~m[1613]&~m[1615]&~m[1616]&~m[1617])|(~m[749]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(m[749]&m[1613]&~m[1615]&m[1616]&~m[1617])|(m[749]&~m[1613]&m[1615]&m[1616]&~m[1617])|(~m[749]&m[1613]&~m[1615]&~m[1616]&m[1617])|(~m[749]&~m[1613]&m[1615]&~m[1616]&m[1617])|(m[749]&m[1613]&m[1615]&~m[1616]&m[1617])|(~m[749]&m[1613]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[633])|((m[749]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(~m[749]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[749]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[749]&m[1613]&~m[1615]&~m[1616]&m[1617])|(m[749]&~m[1613]&m[1615]&~m[1616]&m[1617])|(~m[749]&~m[1613]&~m[1615]&m[1616]&m[1617])|(m[749]&~m[1613]&~m[1615]&m[1616]&m[1617])|(~m[749]&m[1613]&~m[1615]&m[1616]&m[1617])|(m[749]&m[1613]&~m[1615]&m[1616]&m[1617])|(~m[749]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[749]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[749]&m[1613]&m[1615]&m[1616]&m[1617]))):InitCond[1528];
    m[1619] = run?((((m[764]&~m[1618]&~m[1620]&~m[1621]&~m[1622])|(~m[764]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(m[764]&m[1618]&~m[1620]&m[1621]&~m[1622])|(m[764]&~m[1618]&m[1620]&m[1621]&~m[1622])|(~m[764]&m[1618]&~m[1620]&~m[1621]&m[1622])|(~m[764]&~m[1618]&m[1620]&~m[1621]&m[1622])|(m[764]&m[1618]&m[1620]&~m[1621]&m[1622])|(~m[764]&m[1618]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[634])|((m[764]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(~m[764]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[764]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[764]&m[1618]&~m[1620]&~m[1621]&m[1622])|(m[764]&~m[1618]&m[1620]&~m[1621]&m[1622])|(~m[764]&~m[1618]&~m[1620]&m[1621]&m[1622])|(m[764]&~m[1618]&~m[1620]&m[1621]&m[1622])|(~m[764]&m[1618]&~m[1620]&m[1621]&m[1622])|(m[764]&m[1618]&~m[1620]&m[1621]&m[1622])|(~m[764]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[764]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[764]&m[1618]&m[1620]&m[1621]&m[1622]))):InitCond[1529];
    m[1624] = run?((((m[779]&~m[1623]&~m[1625]&~m[1626]&~m[1627])|(~m[779]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(m[779]&m[1623]&~m[1625]&m[1626]&~m[1627])|(m[779]&~m[1623]&m[1625]&m[1626]&~m[1627])|(~m[779]&m[1623]&~m[1625]&~m[1626]&m[1627])|(~m[779]&~m[1623]&m[1625]&~m[1626]&m[1627])|(m[779]&m[1623]&m[1625]&~m[1626]&m[1627])|(~m[779]&m[1623]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[635])|((m[779]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(~m[779]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[779]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[779]&m[1623]&~m[1625]&~m[1626]&m[1627])|(m[779]&~m[1623]&m[1625]&~m[1626]&m[1627])|(~m[779]&~m[1623]&~m[1625]&m[1626]&m[1627])|(m[779]&~m[1623]&~m[1625]&m[1626]&m[1627])|(~m[779]&m[1623]&~m[1625]&m[1626]&m[1627])|(m[779]&m[1623]&~m[1625]&m[1626]&m[1627])|(~m[779]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[779]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[779]&m[1623]&m[1625]&m[1626]&m[1627]))):InitCond[1530];
    m[1629] = run?((((m[794]&~m[1628]&~m[1630]&~m[1631]&~m[1632])|(~m[794]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(m[794]&m[1628]&~m[1630]&m[1631]&~m[1632])|(m[794]&~m[1628]&m[1630]&m[1631]&~m[1632])|(~m[794]&m[1628]&~m[1630]&~m[1631]&m[1632])|(~m[794]&~m[1628]&m[1630]&~m[1631]&m[1632])|(m[794]&m[1628]&m[1630]&~m[1631]&m[1632])|(~m[794]&m[1628]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[636])|((m[794]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(~m[794]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[794]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[794]&m[1628]&~m[1630]&~m[1631]&m[1632])|(m[794]&~m[1628]&m[1630]&~m[1631]&m[1632])|(~m[794]&~m[1628]&~m[1630]&m[1631]&m[1632])|(m[794]&~m[1628]&~m[1630]&m[1631]&m[1632])|(~m[794]&m[1628]&~m[1630]&m[1631]&m[1632])|(m[794]&m[1628]&~m[1630]&m[1631]&m[1632])|(~m[794]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[794]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[794]&m[1628]&m[1630]&m[1631]&m[1632]))):InitCond[1531];
    m[1634] = run?((((m[809]&~m[1633]&~m[1635]&~m[1636]&~m[1637])|(~m[809]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(m[809]&m[1633]&~m[1635]&m[1636]&~m[1637])|(m[809]&~m[1633]&m[1635]&m[1636]&~m[1637])|(~m[809]&m[1633]&~m[1635]&~m[1636]&m[1637])|(~m[809]&~m[1633]&m[1635]&~m[1636]&m[1637])|(m[809]&m[1633]&m[1635]&~m[1636]&m[1637])|(~m[809]&m[1633]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[637])|((m[809]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(~m[809]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[809]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[809]&m[1633]&~m[1635]&~m[1636]&m[1637])|(m[809]&~m[1633]&m[1635]&~m[1636]&m[1637])|(~m[809]&~m[1633]&~m[1635]&m[1636]&m[1637])|(m[809]&~m[1633]&~m[1635]&m[1636]&m[1637])|(~m[809]&m[1633]&~m[1635]&m[1636]&m[1637])|(m[809]&m[1633]&~m[1635]&m[1636]&m[1637])|(~m[809]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[809]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[809]&m[1633]&m[1635]&m[1636]&m[1637]))):InitCond[1532];
    m[1639] = run?((((m[824]&~m[1638]&~m[1640]&~m[1641]&~m[1642])|(~m[824]&~m[1638]&~m[1640]&m[1641]&~m[1642])|(m[824]&m[1638]&~m[1640]&m[1641]&~m[1642])|(m[824]&~m[1638]&m[1640]&m[1641]&~m[1642])|(~m[824]&m[1638]&~m[1640]&~m[1641]&m[1642])|(~m[824]&~m[1638]&m[1640]&~m[1641]&m[1642])|(m[824]&m[1638]&m[1640]&~m[1641]&m[1642])|(~m[824]&m[1638]&m[1640]&m[1641]&m[1642]))&UnbiasedRNG[638])|((m[824]&~m[1638]&~m[1640]&m[1641]&~m[1642])|(~m[824]&~m[1638]&~m[1640]&~m[1641]&m[1642])|(m[824]&~m[1638]&~m[1640]&~m[1641]&m[1642])|(m[824]&m[1638]&~m[1640]&~m[1641]&m[1642])|(m[824]&~m[1638]&m[1640]&~m[1641]&m[1642])|(~m[824]&~m[1638]&~m[1640]&m[1641]&m[1642])|(m[824]&~m[1638]&~m[1640]&m[1641]&m[1642])|(~m[824]&m[1638]&~m[1640]&m[1641]&m[1642])|(m[824]&m[1638]&~m[1640]&m[1641]&m[1642])|(~m[824]&~m[1638]&m[1640]&m[1641]&m[1642])|(m[824]&~m[1638]&m[1640]&m[1641]&m[1642])|(m[824]&m[1638]&m[1640]&m[1641]&m[1642]))):InitCond[1533];
    m[1644] = run?((((m[839]&~m[1643]&~m[1645]&~m[1646]&~m[1647])|(~m[839]&~m[1643]&~m[1645]&m[1646]&~m[1647])|(m[839]&m[1643]&~m[1645]&m[1646]&~m[1647])|(m[839]&~m[1643]&m[1645]&m[1646]&~m[1647])|(~m[839]&m[1643]&~m[1645]&~m[1646]&m[1647])|(~m[839]&~m[1643]&m[1645]&~m[1646]&m[1647])|(m[839]&m[1643]&m[1645]&~m[1646]&m[1647])|(~m[839]&m[1643]&m[1645]&m[1646]&m[1647]))&UnbiasedRNG[639])|((m[839]&~m[1643]&~m[1645]&m[1646]&~m[1647])|(~m[839]&~m[1643]&~m[1645]&~m[1646]&m[1647])|(m[839]&~m[1643]&~m[1645]&~m[1646]&m[1647])|(m[839]&m[1643]&~m[1645]&~m[1646]&m[1647])|(m[839]&~m[1643]&m[1645]&~m[1646]&m[1647])|(~m[839]&~m[1643]&~m[1645]&m[1646]&m[1647])|(m[839]&~m[1643]&~m[1645]&m[1646]&m[1647])|(~m[839]&m[1643]&~m[1645]&m[1646]&m[1647])|(m[839]&m[1643]&~m[1645]&m[1646]&m[1647])|(~m[839]&~m[1643]&m[1645]&m[1646]&m[1647])|(m[839]&~m[1643]&m[1645]&m[1646]&m[1647])|(m[839]&m[1643]&m[1645]&m[1646]&m[1647]))):InitCond[1534];
    m[1649] = run?((((m[854]&~m[1648]&~m[1650]&~m[1651]&~m[1652])|(~m[854]&~m[1648]&~m[1650]&m[1651]&~m[1652])|(m[854]&m[1648]&~m[1650]&m[1651]&~m[1652])|(m[854]&~m[1648]&m[1650]&m[1651]&~m[1652])|(~m[854]&m[1648]&~m[1650]&~m[1651]&m[1652])|(~m[854]&~m[1648]&m[1650]&~m[1651]&m[1652])|(m[854]&m[1648]&m[1650]&~m[1651]&m[1652])|(~m[854]&m[1648]&m[1650]&m[1651]&m[1652]))&UnbiasedRNG[640])|((m[854]&~m[1648]&~m[1650]&m[1651]&~m[1652])|(~m[854]&~m[1648]&~m[1650]&~m[1651]&m[1652])|(m[854]&~m[1648]&~m[1650]&~m[1651]&m[1652])|(m[854]&m[1648]&~m[1650]&~m[1651]&m[1652])|(m[854]&~m[1648]&m[1650]&~m[1651]&m[1652])|(~m[854]&~m[1648]&~m[1650]&m[1651]&m[1652])|(m[854]&~m[1648]&~m[1650]&m[1651]&m[1652])|(~m[854]&m[1648]&~m[1650]&m[1651]&m[1652])|(m[854]&m[1648]&~m[1650]&m[1651]&m[1652])|(~m[854]&~m[1648]&m[1650]&m[1651]&m[1652])|(m[854]&~m[1648]&m[1650]&m[1651]&m[1652])|(m[854]&m[1648]&m[1650]&m[1651]&m[1652]))):InitCond[1535];
    m[1654] = run?((((m[869]&~m[1653]&~m[1655]&~m[1656]&~m[1657])|(~m[869]&~m[1653]&~m[1655]&m[1656]&~m[1657])|(m[869]&m[1653]&~m[1655]&m[1656]&~m[1657])|(m[869]&~m[1653]&m[1655]&m[1656]&~m[1657])|(~m[869]&m[1653]&~m[1655]&~m[1656]&m[1657])|(~m[869]&~m[1653]&m[1655]&~m[1656]&m[1657])|(m[869]&m[1653]&m[1655]&~m[1656]&m[1657])|(~m[869]&m[1653]&m[1655]&m[1656]&m[1657]))&UnbiasedRNG[641])|((m[869]&~m[1653]&~m[1655]&m[1656]&~m[1657])|(~m[869]&~m[1653]&~m[1655]&~m[1656]&m[1657])|(m[869]&~m[1653]&~m[1655]&~m[1656]&m[1657])|(m[869]&m[1653]&~m[1655]&~m[1656]&m[1657])|(m[869]&~m[1653]&m[1655]&~m[1656]&m[1657])|(~m[869]&~m[1653]&~m[1655]&m[1656]&m[1657])|(m[869]&~m[1653]&~m[1655]&m[1656]&m[1657])|(~m[869]&m[1653]&~m[1655]&m[1656]&m[1657])|(m[869]&m[1653]&~m[1655]&m[1656]&m[1657])|(~m[869]&~m[1653]&m[1655]&m[1656]&m[1657])|(m[869]&~m[1653]&m[1655]&m[1656]&m[1657])|(m[869]&m[1653]&m[1655]&m[1656]&m[1657]))):InitCond[1536];
    m[1659] = run?((((m[884]&~m[1658]&~m[1660]&~m[1661]&~m[1662])|(~m[884]&~m[1658]&~m[1660]&m[1661]&~m[1662])|(m[884]&m[1658]&~m[1660]&m[1661]&~m[1662])|(m[884]&~m[1658]&m[1660]&m[1661]&~m[1662])|(~m[884]&m[1658]&~m[1660]&~m[1661]&m[1662])|(~m[884]&~m[1658]&m[1660]&~m[1661]&m[1662])|(m[884]&m[1658]&m[1660]&~m[1661]&m[1662])|(~m[884]&m[1658]&m[1660]&m[1661]&m[1662]))&UnbiasedRNG[642])|((m[884]&~m[1658]&~m[1660]&m[1661]&~m[1662])|(~m[884]&~m[1658]&~m[1660]&~m[1661]&m[1662])|(m[884]&~m[1658]&~m[1660]&~m[1661]&m[1662])|(m[884]&m[1658]&~m[1660]&~m[1661]&m[1662])|(m[884]&~m[1658]&m[1660]&~m[1661]&m[1662])|(~m[884]&~m[1658]&~m[1660]&m[1661]&m[1662])|(m[884]&~m[1658]&~m[1660]&m[1661]&m[1662])|(~m[884]&m[1658]&~m[1660]&m[1661]&m[1662])|(m[884]&m[1658]&~m[1660]&m[1661]&m[1662])|(~m[884]&~m[1658]&m[1660]&m[1661]&m[1662])|(m[884]&~m[1658]&m[1660]&m[1661]&m[1662])|(m[884]&m[1658]&m[1660]&m[1661]&m[1662]))):InitCond[1537];
    m[1664] = run?((((m[899]&~m[1663]&~m[1665]&~m[1666]&~m[1667])|(~m[899]&~m[1663]&~m[1665]&m[1666]&~m[1667])|(m[899]&m[1663]&~m[1665]&m[1666]&~m[1667])|(m[899]&~m[1663]&m[1665]&m[1666]&~m[1667])|(~m[899]&m[1663]&~m[1665]&~m[1666]&m[1667])|(~m[899]&~m[1663]&m[1665]&~m[1666]&m[1667])|(m[899]&m[1663]&m[1665]&~m[1666]&m[1667])|(~m[899]&m[1663]&m[1665]&m[1666]&m[1667]))&UnbiasedRNG[643])|((m[899]&~m[1663]&~m[1665]&m[1666]&~m[1667])|(~m[899]&~m[1663]&~m[1665]&~m[1666]&m[1667])|(m[899]&~m[1663]&~m[1665]&~m[1666]&m[1667])|(m[899]&m[1663]&~m[1665]&~m[1666]&m[1667])|(m[899]&~m[1663]&m[1665]&~m[1666]&m[1667])|(~m[899]&~m[1663]&~m[1665]&m[1666]&m[1667])|(m[899]&~m[1663]&~m[1665]&m[1666]&m[1667])|(~m[899]&m[1663]&~m[1665]&m[1666]&m[1667])|(m[899]&m[1663]&~m[1665]&m[1666]&m[1667])|(~m[899]&~m[1663]&m[1665]&m[1666]&m[1667])|(m[899]&~m[1663]&m[1665]&m[1666]&m[1667])|(m[899]&m[1663]&m[1665]&m[1666]&m[1667]))):InitCond[1538];
    m[1669] = run?((((m[914]&~m[1668]&~m[1670]&~m[1671]&~m[1672])|(~m[914]&~m[1668]&~m[1670]&m[1671]&~m[1672])|(m[914]&m[1668]&~m[1670]&m[1671]&~m[1672])|(m[914]&~m[1668]&m[1670]&m[1671]&~m[1672])|(~m[914]&m[1668]&~m[1670]&~m[1671]&m[1672])|(~m[914]&~m[1668]&m[1670]&~m[1671]&m[1672])|(m[914]&m[1668]&m[1670]&~m[1671]&m[1672])|(~m[914]&m[1668]&m[1670]&m[1671]&m[1672]))&UnbiasedRNG[644])|((m[914]&~m[1668]&~m[1670]&m[1671]&~m[1672])|(~m[914]&~m[1668]&~m[1670]&~m[1671]&m[1672])|(m[914]&~m[1668]&~m[1670]&~m[1671]&m[1672])|(m[914]&m[1668]&~m[1670]&~m[1671]&m[1672])|(m[914]&~m[1668]&m[1670]&~m[1671]&m[1672])|(~m[914]&~m[1668]&~m[1670]&m[1671]&m[1672])|(m[914]&~m[1668]&~m[1670]&m[1671]&m[1672])|(~m[914]&m[1668]&~m[1670]&m[1671]&m[1672])|(m[914]&m[1668]&~m[1670]&m[1671]&m[1672])|(~m[914]&~m[1668]&m[1670]&m[1671]&m[1672])|(m[914]&~m[1668]&m[1670]&m[1671]&m[1672])|(m[914]&m[1668]&m[1670]&m[1671]&m[1672]))):InitCond[1539];
    m[1674] = run?((((m[735]&~m[1673]&~m[1675]&~m[1676]&~m[1677])|(~m[735]&~m[1673]&~m[1675]&m[1676]&~m[1677])|(m[735]&m[1673]&~m[1675]&m[1676]&~m[1677])|(m[735]&~m[1673]&m[1675]&m[1676]&~m[1677])|(~m[735]&m[1673]&~m[1675]&~m[1676]&m[1677])|(~m[735]&~m[1673]&m[1675]&~m[1676]&m[1677])|(m[735]&m[1673]&m[1675]&~m[1676]&m[1677])|(~m[735]&m[1673]&m[1675]&m[1676]&m[1677]))&UnbiasedRNG[645])|((m[735]&~m[1673]&~m[1675]&m[1676]&~m[1677])|(~m[735]&~m[1673]&~m[1675]&~m[1676]&m[1677])|(m[735]&~m[1673]&~m[1675]&~m[1676]&m[1677])|(m[735]&m[1673]&~m[1675]&~m[1676]&m[1677])|(m[735]&~m[1673]&m[1675]&~m[1676]&m[1677])|(~m[735]&~m[1673]&~m[1675]&m[1676]&m[1677])|(m[735]&~m[1673]&~m[1675]&m[1676]&m[1677])|(~m[735]&m[1673]&~m[1675]&m[1676]&m[1677])|(m[735]&m[1673]&~m[1675]&m[1676]&m[1677])|(~m[735]&~m[1673]&m[1675]&m[1676]&m[1677])|(m[735]&~m[1673]&m[1675]&m[1676]&m[1677])|(m[735]&m[1673]&m[1675]&m[1676]&m[1677]))):InitCond[1540];
    m[1679] = run?((((m[750]&~m[1678]&~m[1680]&~m[1681]&~m[1682])|(~m[750]&~m[1678]&~m[1680]&m[1681]&~m[1682])|(m[750]&m[1678]&~m[1680]&m[1681]&~m[1682])|(m[750]&~m[1678]&m[1680]&m[1681]&~m[1682])|(~m[750]&m[1678]&~m[1680]&~m[1681]&m[1682])|(~m[750]&~m[1678]&m[1680]&~m[1681]&m[1682])|(m[750]&m[1678]&m[1680]&~m[1681]&m[1682])|(~m[750]&m[1678]&m[1680]&m[1681]&m[1682]))&UnbiasedRNG[646])|((m[750]&~m[1678]&~m[1680]&m[1681]&~m[1682])|(~m[750]&~m[1678]&~m[1680]&~m[1681]&m[1682])|(m[750]&~m[1678]&~m[1680]&~m[1681]&m[1682])|(m[750]&m[1678]&~m[1680]&~m[1681]&m[1682])|(m[750]&~m[1678]&m[1680]&~m[1681]&m[1682])|(~m[750]&~m[1678]&~m[1680]&m[1681]&m[1682])|(m[750]&~m[1678]&~m[1680]&m[1681]&m[1682])|(~m[750]&m[1678]&~m[1680]&m[1681]&m[1682])|(m[750]&m[1678]&~m[1680]&m[1681]&m[1682])|(~m[750]&~m[1678]&m[1680]&m[1681]&m[1682])|(m[750]&~m[1678]&m[1680]&m[1681]&m[1682])|(m[750]&m[1678]&m[1680]&m[1681]&m[1682]))):InitCond[1541];
    m[1684] = run?((((m[765]&~m[1683]&~m[1685]&~m[1686]&~m[1687])|(~m[765]&~m[1683]&~m[1685]&m[1686]&~m[1687])|(m[765]&m[1683]&~m[1685]&m[1686]&~m[1687])|(m[765]&~m[1683]&m[1685]&m[1686]&~m[1687])|(~m[765]&m[1683]&~m[1685]&~m[1686]&m[1687])|(~m[765]&~m[1683]&m[1685]&~m[1686]&m[1687])|(m[765]&m[1683]&m[1685]&~m[1686]&m[1687])|(~m[765]&m[1683]&m[1685]&m[1686]&m[1687]))&UnbiasedRNG[647])|((m[765]&~m[1683]&~m[1685]&m[1686]&~m[1687])|(~m[765]&~m[1683]&~m[1685]&~m[1686]&m[1687])|(m[765]&~m[1683]&~m[1685]&~m[1686]&m[1687])|(m[765]&m[1683]&~m[1685]&~m[1686]&m[1687])|(m[765]&~m[1683]&m[1685]&~m[1686]&m[1687])|(~m[765]&~m[1683]&~m[1685]&m[1686]&m[1687])|(m[765]&~m[1683]&~m[1685]&m[1686]&m[1687])|(~m[765]&m[1683]&~m[1685]&m[1686]&m[1687])|(m[765]&m[1683]&~m[1685]&m[1686]&m[1687])|(~m[765]&~m[1683]&m[1685]&m[1686]&m[1687])|(m[765]&~m[1683]&m[1685]&m[1686]&m[1687])|(m[765]&m[1683]&m[1685]&m[1686]&m[1687]))):InitCond[1542];
    m[1689] = run?((((m[780]&~m[1688]&~m[1690]&~m[1691]&~m[1692])|(~m[780]&~m[1688]&~m[1690]&m[1691]&~m[1692])|(m[780]&m[1688]&~m[1690]&m[1691]&~m[1692])|(m[780]&~m[1688]&m[1690]&m[1691]&~m[1692])|(~m[780]&m[1688]&~m[1690]&~m[1691]&m[1692])|(~m[780]&~m[1688]&m[1690]&~m[1691]&m[1692])|(m[780]&m[1688]&m[1690]&~m[1691]&m[1692])|(~m[780]&m[1688]&m[1690]&m[1691]&m[1692]))&UnbiasedRNG[648])|((m[780]&~m[1688]&~m[1690]&m[1691]&~m[1692])|(~m[780]&~m[1688]&~m[1690]&~m[1691]&m[1692])|(m[780]&~m[1688]&~m[1690]&~m[1691]&m[1692])|(m[780]&m[1688]&~m[1690]&~m[1691]&m[1692])|(m[780]&~m[1688]&m[1690]&~m[1691]&m[1692])|(~m[780]&~m[1688]&~m[1690]&m[1691]&m[1692])|(m[780]&~m[1688]&~m[1690]&m[1691]&m[1692])|(~m[780]&m[1688]&~m[1690]&m[1691]&m[1692])|(m[780]&m[1688]&~m[1690]&m[1691]&m[1692])|(~m[780]&~m[1688]&m[1690]&m[1691]&m[1692])|(m[780]&~m[1688]&m[1690]&m[1691]&m[1692])|(m[780]&m[1688]&m[1690]&m[1691]&m[1692]))):InitCond[1543];
    m[1694] = run?((((m[795]&~m[1693]&~m[1695]&~m[1696]&~m[1697])|(~m[795]&~m[1693]&~m[1695]&m[1696]&~m[1697])|(m[795]&m[1693]&~m[1695]&m[1696]&~m[1697])|(m[795]&~m[1693]&m[1695]&m[1696]&~m[1697])|(~m[795]&m[1693]&~m[1695]&~m[1696]&m[1697])|(~m[795]&~m[1693]&m[1695]&~m[1696]&m[1697])|(m[795]&m[1693]&m[1695]&~m[1696]&m[1697])|(~m[795]&m[1693]&m[1695]&m[1696]&m[1697]))&UnbiasedRNG[649])|((m[795]&~m[1693]&~m[1695]&m[1696]&~m[1697])|(~m[795]&~m[1693]&~m[1695]&~m[1696]&m[1697])|(m[795]&~m[1693]&~m[1695]&~m[1696]&m[1697])|(m[795]&m[1693]&~m[1695]&~m[1696]&m[1697])|(m[795]&~m[1693]&m[1695]&~m[1696]&m[1697])|(~m[795]&~m[1693]&~m[1695]&m[1696]&m[1697])|(m[795]&~m[1693]&~m[1695]&m[1696]&m[1697])|(~m[795]&m[1693]&~m[1695]&m[1696]&m[1697])|(m[795]&m[1693]&~m[1695]&m[1696]&m[1697])|(~m[795]&~m[1693]&m[1695]&m[1696]&m[1697])|(m[795]&~m[1693]&m[1695]&m[1696]&m[1697])|(m[795]&m[1693]&m[1695]&m[1696]&m[1697]))):InitCond[1544];
    m[1699] = run?((((m[810]&~m[1698]&~m[1700]&~m[1701]&~m[1702])|(~m[810]&~m[1698]&~m[1700]&m[1701]&~m[1702])|(m[810]&m[1698]&~m[1700]&m[1701]&~m[1702])|(m[810]&~m[1698]&m[1700]&m[1701]&~m[1702])|(~m[810]&m[1698]&~m[1700]&~m[1701]&m[1702])|(~m[810]&~m[1698]&m[1700]&~m[1701]&m[1702])|(m[810]&m[1698]&m[1700]&~m[1701]&m[1702])|(~m[810]&m[1698]&m[1700]&m[1701]&m[1702]))&UnbiasedRNG[650])|((m[810]&~m[1698]&~m[1700]&m[1701]&~m[1702])|(~m[810]&~m[1698]&~m[1700]&~m[1701]&m[1702])|(m[810]&~m[1698]&~m[1700]&~m[1701]&m[1702])|(m[810]&m[1698]&~m[1700]&~m[1701]&m[1702])|(m[810]&~m[1698]&m[1700]&~m[1701]&m[1702])|(~m[810]&~m[1698]&~m[1700]&m[1701]&m[1702])|(m[810]&~m[1698]&~m[1700]&m[1701]&m[1702])|(~m[810]&m[1698]&~m[1700]&m[1701]&m[1702])|(m[810]&m[1698]&~m[1700]&m[1701]&m[1702])|(~m[810]&~m[1698]&m[1700]&m[1701]&m[1702])|(m[810]&~m[1698]&m[1700]&m[1701]&m[1702])|(m[810]&m[1698]&m[1700]&m[1701]&m[1702]))):InitCond[1545];
    m[1704] = run?((((m[825]&~m[1703]&~m[1705]&~m[1706]&~m[1707])|(~m[825]&~m[1703]&~m[1705]&m[1706]&~m[1707])|(m[825]&m[1703]&~m[1705]&m[1706]&~m[1707])|(m[825]&~m[1703]&m[1705]&m[1706]&~m[1707])|(~m[825]&m[1703]&~m[1705]&~m[1706]&m[1707])|(~m[825]&~m[1703]&m[1705]&~m[1706]&m[1707])|(m[825]&m[1703]&m[1705]&~m[1706]&m[1707])|(~m[825]&m[1703]&m[1705]&m[1706]&m[1707]))&UnbiasedRNG[651])|((m[825]&~m[1703]&~m[1705]&m[1706]&~m[1707])|(~m[825]&~m[1703]&~m[1705]&~m[1706]&m[1707])|(m[825]&~m[1703]&~m[1705]&~m[1706]&m[1707])|(m[825]&m[1703]&~m[1705]&~m[1706]&m[1707])|(m[825]&~m[1703]&m[1705]&~m[1706]&m[1707])|(~m[825]&~m[1703]&~m[1705]&m[1706]&m[1707])|(m[825]&~m[1703]&~m[1705]&m[1706]&m[1707])|(~m[825]&m[1703]&~m[1705]&m[1706]&m[1707])|(m[825]&m[1703]&~m[1705]&m[1706]&m[1707])|(~m[825]&~m[1703]&m[1705]&m[1706]&m[1707])|(m[825]&~m[1703]&m[1705]&m[1706]&m[1707])|(m[825]&m[1703]&m[1705]&m[1706]&m[1707]))):InitCond[1546];
    m[1709] = run?((((m[840]&~m[1708]&~m[1710]&~m[1711]&~m[1712])|(~m[840]&~m[1708]&~m[1710]&m[1711]&~m[1712])|(m[840]&m[1708]&~m[1710]&m[1711]&~m[1712])|(m[840]&~m[1708]&m[1710]&m[1711]&~m[1712])|(~m[840]&m[1708]&~m[1710]&~m[1711]&m[1712])|(~m[840]&~m[1708]&m[1710]&~m[1711]&m[1712])|(m[840]&m[1708]&m[1710]&~m[1711]&m[1712])|(~m[840]&m[1708]&m[1710]&m[1711]&m[1712]))&UnbiasedRNG[652])|((m[840]&~m[1708]&~m[1710]&m[1711]&~m[1712])|(~m[840]&~m[1708]&~m[1710]&~m[1711]&m[1712])|(m[840]&~m[1708]&~m[1710]&~m[1711]&m[1712])|(m[840]&m[1708]&~m[1710]&~m[1711]&m[1712])|(m[840]&~m[1708]&m[1710]&~m[1711]&m[1712])|(~m[840]&~m[1708]&~m[1710]&m[1711]&m[1712])|(m[840]&~m[1708]&~m[1710]&m[1711]&m[1712])|(~m[840]&m[1708]&~m[1710]&m[1711]&m[1712])|(m[840]&m[1708]&~m[1710]&m[1711]&m[1712])|(~m[840]&~m[1708]&m[1710]&m[1711]&m[1712])|(m[840]&~m[1708]&m[1710]&m[1711]&m[1712])|(m[840]&m[1708]&m[1710]&m[1711]&m[1712]))):InitCond[1547];
    m[1714] = run?((((m[855]&~m[1713]&~m[1715]&~m[1716]&~m[1717])|(~m[855]&~m[1713]&~m[1715]&m[1716]&~m[1717])|(m[855]&m[1713]&~m[1715]&m[1716]&~m[1717])|(m[855]&~m[1713]&m[1715]&m[1716]&~m[1717])|(~m[855]&m[1713]&~m[1715]&~m[1716]&m[1717])|(~m[855]&~m[1713]&m[1715]&~m[1716]&m[1717])|(m[855]&m[1713]&m[1715]&~m[1716]&m[1717])|(~m[855]&m[1713]&m[1715]&m[1716]&m[1717]))&UnbiasedRNG[653])|((m[855]&~m[1713]&~m[1715]&m[1716]&~m[1717])|(~m[855]&~m[1713]&~m[1715]&~m[1716]&m[1717])|(m[855]&~m[1713]&~m[1715]&~m[1716]&m[1717])|(m[855]&m[1713]&~m[1715]&~m[1716]&m[1717])|(m[855]&~m[1713]&m[1715]&~m[1716]&m[1717])|(~m[855]&~m[1713]&~m[1715]&m[1716]&m[1717])|(m[855]&~m[1713]&~m[1715]&m[1716]&m[1717])|(~m[855]&m[1713]&~m[1715]&m[1716]&m[1717])|(m[855]&m[1713]&~m[1715]&m[1716]&m[1717])|(~m[855]&~m[1713]&m[1715]&m[1716]&m[1717])|(m[855]&~m[1713]&m[1715]&m[1716]&m[1717])|(m[855]&m[1713]&m[1715]&m[1716]&m[1717]))):InitCond[1548];
    m[1719] = run?((((m[870]&~m[1718]&~m[1720]&~m[1721]&~m[1722])|(~m[870]&~m[1718]&~m[1720]&m[1721]&~m[1722])|(m[870]&m[1718]&~m[1720]&m[1721]&~m[1722])|(m[870]&~m[1718]&m[1720]&m[1721]&~m[1722])|(~m[870]&m[1718]&~m[1720]&~m[1721]&m[1722])|(~m[870]&~m[1718]&m[1720]&~m[1721]&m[1722])|(m[870]&m[1718]&m[1720]&~m[1721]&m[1722])|(~m[870]&m[1718]&m[1720]&m[1721]&m[1722]))&UnbiasedRNG[654])|((m[870]&~m[1718]&~m[1720]&m[1721]&~m[1722])|(~m[870]&~m[1718]&~m[1720]&~m[1721]&m[1722])|(m[870]&~m[1718]&~m[1720]&~m[1721]&m[1722])|(m[870]&m[1718]&~m[1720]&~m[1721]&m[1722])|(m[870]&~m[1718]&m[1720]&~m[1721]&m[1722])|(~m[870]&~m[1718]&~m[1720]&m[1721]&m[1722])|(m[870]&~m[1718]&~m[1720]&m[1721]&m[1722])|(~m[870]&m[1718]&~m[1720]&m[1721]&m[1722])|(m[870]&m[1718]&~m[1720]&m[1721]&m[1722])|(~m[870]&~m[1718]&m[1720]&m[1721]&m[1722])|(m[870]&~m[1718]&m[1720]&m[1721]&m[1722])|(m[870]&m[1718]&m[1720]&m[1721]&m[1722]))):InitCond[1549];
    m[1724] = run?((((m[885]&~m[1723]&~m[1725]&~m[1726]&~m[1727])|(~m[885]&~m[1723]&~m[1725]&m[1726]&~m[1727])|(m[885]&m[1723]&~m[1725]&m[1726]&~m[1727])|(m[885]&~m[1723]&m[1725]&m[1726]&~m[1727])|(~m[885]&m[1723]&~m[1725]&~m[1726]&m[1727])|(~m[885]&~m[1723]&m[1725]&~m[1726]&m[1727])|(m[885]&m[1723]&m[1725]&~m[1726]&m[1727])|(~m[885]&m[1723]&m[1725]&m[1726]&m[1727]))&UnbiasedRNG[655])|((m[885]&~m[1723]&~m[1725]&m[1726]&~m[1727])|(~m[885]&~m[1723]&~m[1725]&~m[1726]&m[1727])|(m[885]&~m[1723]&~m[1725]&~m[1726]&m[1727])|(m[885]&m[1723]&~m[1725]&~m[1726]&m[1727])|(m[885]&~m[1723]&m[1725]&~m[1726]&m[1727])|(~m[885]&~m[1723]&~m[1725]&m[1726]&m[1727])|(m[885]&~m[1723]&~m[1725]&m[1726]&m[1727])|(~m[885]&m[1723]&~m[1725]&m[1726]&m[1727])|(m[885]&m[1723]&~m[1725]&m[1726]&m[1727])|(~m[885]&~m[1723]&m[1725]&m[1726]&m[1727])|(m[885]&~m[1723]&m[1725]&m[1726]&m[1727])|(m[885]&m[1723]&m[1725]&m[1726]&m[1727]))):InitCond[1550];
    m[1729] = run?((((m[900]&~m[1728]&~m[1730]&~m[1731]&~m[1732])|(~m[900]&~m[1728]&~m[1730]&m[1731]&~m[1732])|(m[900]&m[1728]&~m[1730]&m[1731]&~m[1732])|(m[900]&~m[1728]&m[1730]&m[1731]&~m[1732])|(~m[900]&m[1728]&~m[1730]&~m[1731]&m[1732])|(~m[900]&~m[1728]&m[1730]&~m[1731]&m[1732])|(m[900]&m[1728]&m[1730]&~m[1731]&m[1732])|(~m[900]&m[1728]&m[1730]&m[1731]&m[1732]))&UnbiasedRNG[656])|((m[900]&~m[1728]&~m[1730]&m[1731]&~m[1732])|(~m[900]&~m[1728]&~m[1730]&~m[1731]&m[1732])|(m[900]&~m[1728]&~m[1730]&~m[1731]&m[1732])|(m[900]&m[1728]&~m[1730]&~m[1731]&m[1732])|(m[900]&~m[1728]&m[1730]&~m[1731]&m[1732])|(~m[900]&~m[1728]&~m[1730]&m[1731]&m[1732])|(m[900]&~m[1728]&~m[1730]&m[1731]&m[1732])|(~m[900]&m[1728]&~m[1730]&m[1731]&m[1732])|(m[900]&m[1728]&~m[1730]&m[1731]&m[1732])|(~m[900]&~m[1728]&m[1730]&m[1731]&m[1732])|(m[900]&~m[1728]&m[1730]&m[1731]&m[1732])|(m[900]&m[1728]&m[1730]&m[1731]&m[1732]))):InitCond[1551];
    m[1734] = run?((((m[915]&~m[1733]&~m[1735]&~m[1736]&~m[1737])|(~m[915]&~m[1733]&~m[1735]&m[1736]&~m[1737])|(m[915]&m[1733]&~m[1735]&m[1736]&~m[1737])|(m[915]&~m[1733]&m[1735]&m[1736]&~m[1737])|(~m[915]&m[1733]&~m[1735]&~m[1736]&m[1737])|(~m[915]&~m[1733]&m[1735]&~m[1736]&m[1737])|(m[915]&m[1733]&m[1735]&~m[1736]&m[1737])|(~m[915]&m[1733]&m[1735]&m[1736]&m[1737]))&UnbiasedRNG[657])|((m[915]&~m[1733]&~m[1735]&m[1736]&~m[1737])|(~m[915]&~m[1733]&~m[1735]&~m[1736]&m[1737])|(m[915]&~m[1733]&~m[1735]&~m[1736]&m[1737])|(m[915]&m[1733]&~m[1735]&~m[1736]&m[1737])|(m[915]&~m[1733]&m[1735]&~m[1736]&m[1737])|(~m[915]&~m[1733]&~m[1735]&m[1736]&m[1737])|(m[915]&~m[1733]&~m[1735]&m[1736]&m[1737])|(~m[915]&m[1733]&~m[1735]&m[1736]&m[1737])|(m[915]&m[1733]&~m[1735]&m[1736]&m[1737])|(~m[915]&~m[1733]&m[1735]&m[1736]&m[1737])|(m[915]&~m[1733]&m[1735]&m[1736]&m[1737])|(m[915]&m[1733]&m[1735]&m[1736]&m[1737]))):InitCond[1552];
    m[1739] = run?((((m[751]&~m[1738]&~m[1740]&~m[1741]&~m[1742])|(~m[751]&~m[1738]&~m[1740]&m[1741]&~m[1742])|(m[751]&m[1738]&~m[1740]&m[1741]&~m[1742])|(m[751]&~m[1738]&m[1740]&m[1741]&~m[1742])|(~m[751]&m[1738]&~m[1740]&~m[1741]&m[1742])|(~m[751]&~m[1738]&m[1740]&~m[1741]&m[1742])|(m[751]&m[1738]&m[1740]&~m[1741]&m[1742])|(~m[751]&m[1738]&m[1740]&m[1741]&m[1742]))&UnbiasedRNG[658])|((m[751]&~m[1738]&~m[1740]&m[1741]&~m[1742])|(~m[751]&~m[1738]&~m[1740]&~m[1741]&m[1742])|(m[751]&~m[1738]&~m[1740]&~m[1741]&m[1742])|(m[751]&m[1738]&~m[1740]&~m[1741]&m[1742])|(m[751]&~m[1738]&m[1740]&~m[1741]&m[1742])|(~m[751]&~m[1738]&~m[1740]&m[1741]&m[1742])|(m[751]&~m[1738]&~m[1740]&m[1741]&m[1742])|(~m[751]&m[1738]&~m[1740]&m[1741]&m[1742])|(m[751]&m[1738]&~m[1740]&m[1741]&m[1742])|(~m[751]&~m[1738]&m[1740]&m[1741]&m[1742])|(m[751]&~m[1738]&m[1740]&m[1741]&m[1742])|(m[751]&m[1738]&m[1740]&m[1741]&m[1742]))):InitCond[1553];
    m[1744] = run?((((m[766]&~m[1743]&~m[1745]&~m[1746]&~m[1747])|(~m[766]&~m[1743]&~m[1745]&m[1746]&~m[1747])|(m[766]&m[1743]&~m[1745]&m[1746]&~m[1747])|(m[766]&~m[1743]&m[1745]&m[1746]&~m[1747])|(~m[766]&m[1743]&~m[1745]&~m[1746]&m[1747])|(~m[766]&~m[1743]&m[1745]&~m[1746]&m[1747])|(m[766]&m[1743]&m[1745]&~m[1746]&m[1747])|(~m[766]&m[1743]&m[1745]&m[1746]&m[1747]))&UnbiasedRNG[659])|((m[766]&~m[1743]&~m[1745]&m[1746]&~m[1747])|(~m[766]&~m[1743]&~m[1745]&~m[1746]&m[1747])|(m[766]&~m[1743]&~m[1745]&~m[1746]&m[1747])|(m[766]&m[1743]&~m[1745]&~m[1746]&m[1747])|(m[766]&~m[1743]&m[1745]&~m[1746]&m[1747])|(~m[766]&~m[1743]&~m[1745]&m[1746]&m[1747])|(m[766]&~m[1743]&~m[1745]&m[1746]&m[1747])|(~m[766]&m[1743]&~m[1745]&m[1746]&m[1747])|(m[766]&m[1743]&~m[1745]&m[1746]&m[1747])|(~m[766]&~m[1743]&m[1745]&m[1746]&m[1747])|(m[766]&~m[1743]&m[1745]&m[1746]&m[1747])|(m[766]&m[1743]&m[1745]&m[1746]&m[1747]))):InitCond[1554];
    m[1749] = run?((((m[781]&~m[1748]&~m[1750]&~m[1751]&~m[1752])|(~m[781]&~m[1748]&~m[1750]&m[1751]&~m[1752])|(m[781]&m[1748]&~m[1750]&m[1751]&~m[1752])|(m[781]&~m[1748]&m[1750]&m[1751]&~m[1752])|(~m[781]&m[1748]&~m[1750]&~m[1751]&m[1752])|(~m[781]&~m[1748]&m[1750]&~m[1751]&m[1752])|(m[781]&m[1748]&m[1750]&~m[1751]&m[1752])|(~m[781]&m[1748]&m[1750]&m[1751]&m[1752]))&UnbiasedRNG[660])|((m[781]&~m[1748]&~m[1750]&m[1751]&~m[1752])|(~m[781]&~m[1748]&~m[1750]&~m[1751]&m[1752])|(m[781]&~m[1748]&~m[1750]&~m[1751]&m[1752])|(m[781]&m[1748]&~m[1750]&~m[1751]&m[1752])|(m[781]&~m[1748]&m[1750]&~m[1751]&m[1752])|(~m[781]&~m[1748]&~m[1750]&m[1751]&m[1752])|(m[781]&~m[1748]&~m[1750]&m[1751]&m[1752])|(~m[781]&m[1748]&~m[1750]&m[1751]&m[1752])|(m[781]&m[1748]&~m[1750]&m[1751]&m[1752])|(~m[781]&~m[1748]&m[1750]&m[1751]&m[1752])|(m[781]&~m[1748]&m[1750]&m[1751]&m[1752])|(m[781]&m[1748]&m[1750]&m[1751]&m[1752]))):InitCond[1555];
    m[1754] = run?((((m[796]&~m[1753]&~m[1755]&~m[1756]&~m[1757])|(~m[796]&~m[1753]&~m[1755]&m[1756]&~m[1757])|(m[796]&m[1753]&~m[1755]&m[1756]&~m[1757])|(m[796]&~m[1753]&m[1755]&m[1756]&~m[1757])|(~m[796]&m[1753]&~m[1755]&~m[1756]&m[1757])|(~m[796]&~m[1753]&m[1755]&~m[1756]&m[1757])|(m[796]&m[1753]&m[1755]&~m[1756]&m[1757])|(~m[796]&m[1753]&m[1755]&m[1756]&m[1757]))&UnbiasedRNG[661])|((m[796]&~m[1753]&~m[1755]&m[1756]&~m[1757])|(~m[796]&~m[1753]&~m[1755]&~m[1756]&m[1757])|(m[796]&~m[1753]&~m[1755]&~m[1756]&m[1757])|(m[796]&m[1753]&~m[1755]&~m[1756]&m[1757])|(m[796]&~m[1753]&m[1755]&~m[1756]&m[1757])|(~m[796]&~m[1753]&~m[1755]&m[1756]&m[1757])|(m[796]&~m[1753]&~m[1755]&m[1756]&m[1757])|(~m[796]&m[1753]&~m[1755]&m[1756]&m[1757])|(m[796]&m[1753]&~m[1755]&m[1756]&m[1757])|(~m[796]&~m[1753]&m[1755]&m[1756]&m[1757])|(m[796]&~m[1753]&m[1755]&m[1756]&m[1757])|(m[796]&m[1753]&m[1755]&m[1756]&m[1757]))):InitCond[1556];
    m[1759] = run?((((m[811]&~m[1758]&~m[1760]&~m[1761]&~m[1762])|(~m[811]&~m[1758]&~m[1760]&m[1761]&~m[1762])|(m[811]&m[1758]&~m[1760]&m[1761]&~m[1762])|(m[811]&~m[1758]&m[1760]&m[1761]&~m[1762])|(~m[811]&m[1758]&~m[1760]&~m[1761]&m[1762])|(~m[811]&~m[1758]&m[1760]&~m[1761]&m[1762])|(m[811]&m[1758]&m[1760]&~m[1761]&m[1762])|(~m[811]&m[1758]&m[1760]&m[1761]&m[1762]))&UnbiasedRNG[662])|((m[811]&~m[1758]&~m[1760]&m[1761]&~m[1762])|(~m[811]&~m[1758]&~m[1760]&~m[1761]&m[1762])|(m[811]&~m[1758]&~m[1760]&~m[1761]&m[1762])|(m[811]&m[1758]&~m[1760]&~m[1761]&m[1762])|(m[811]&~m[1758]&m[1760]&~m[1761]&m[1762])|(~m[811]&~m[1758]&~m[1760]&m[1761]&m[1762])|(m[811]&~m[1758]&~m[1760]&m[1761]&m[1762])|(~m[811]&m[1758]&~m[1760]&m[1761]&m[1762])|(m[811]&m[1758]&~m[1760]&m[1761]&m[1762])|(~m[811]&~m[1758]&m[1760]&m[1761]&m[1762])|(m[811]&~m[1758]&m[1760]&m[1761]&m[1762])|(m[811]&m[1758]&m[1760]&m[1761]&m[1762]))):InitCond[1557];
    m[1764] = run?((((m[826]&~m[1763]&~m[1765]&~m[1766]&~m[1767])|(~m[826]&~m[1763]&~m[1765]&m[1766]&~m[1767])|(m[826]&m[1763]&~m[1765]&m[1766]&~m[1767])|(m[826]&~m[1763]&m[1765]&m[1766]&~m[1767])|(~m[826]&m[1763]&~m[1765]&~m[1766]&m[1767])|(~m[826]&~m[1763]&m[1765]&~m[1766]&m[1767])|(m[826]&m[1763]&m[1765]&~m[1766]&m[1767])|(~m[826]&m[1763]&m[1765]&m[1766]&m[1767]))&UnbiasedRNG[663])|((m[826]&~m[1763]&~m[1765]&m[1766]&~m[1767])|(~m[826]&~m[1763]&~m[1765]&~m[1766]&m[1767])|(m[826]&~m[1763]&~m[1765]&~m[1766]&m[1767])|(m[826]&m[1763]&~m[1765]&~m[1766]&m[1767])|(m[826]&~m[1763]&m[1765]&~m[1766]&m[1767])|(~m[826]&~m[1763]&~m[1765]&m[1766]&m[1767])|(m[826]&~m[1763]&~m[1765]&m[1766]&m[1767])|(~m[826]&m[1763]&~m[1765]&m[1766]&m[1767])|(m[826]&m[1763]&~m[1765]&m[1766]&m[1767])|(~m[826]&~m[1763]&m[1765]&m[1766]&m[1767])|(m[826]&~m[1763]&m[1765]&m[1766]&m[1767])|(m[826]&m[1763]&m[1765]&m[1766]&m[1767]))):InitCond[1558];
    m[1769] = run?((((m[841]&~m[1768]&~m[1770]&~m[1771]&~m[1772])|(~m[841]&~m[1768]&~m[1770]&m[1771]&~m[1772])|(m[841]&m[1768]&~m[1770]&m[1771]&~m[1772])|(m[841]&~m[1768]&m[1770]&m[1771]&~m[1772])|(~m[841]&m[1768]&~m[1770]&~m[1771]&m[1772])|(~m[841]&~m[1768]&m[1770]&~m[1771]&m[1772])|(m[841]&m[1768]&m[1770]&~m[1771]&m[1772])|(~m[841]&m[1768]&m[1770]&m[1771]&m[1772]))&UnbiasedRNG[664])|((m[841]&~m[1768]&~m[1770]&m[1771]&~m[1772])|(~m[841]&~m[1768]&~m[1770]&~m[1771]&m[1772])|(m[841]&~m[1768]&~m[1770]&~m[1771]&m[1772])|(m[841]&m[1768]&~m[1770]&~m[1771]&m[1772])|(m[841]&~m[1768]&m[1770]&~m[1771]&m[1772])|(~m[841]&~m[1768]&~m[1770]&m[1771]&m[1772])|(m[841]&~m[1768]&~m[1770]&m[1771]&m[1772])|(~m[841]&m[1768]&~m[1770]&m[1771]&m[1772])|(m[841]&m[1768]&~m[1770]&m[1771]&m[1772])|(~m[841]&~m[1768]&m[1770]&m[1771]&m[1772])|(m[841]&~m[1768]&m[1770]&m[1771]&m[1772])|(m[841]&m[1768]&m[1770]&m[1771]&m[1772]))):InitCond[1559];
    m[1774] = run?((((m[856]&~m[1773]&~m[1775]&~m[1776]&~m[1777])|(~m[856]&~m[1773]&~m[1775]&m[1776]&~m[1777])|(m[856]&m[1773]&~m[1775]&m[1776]&~m[1777])|(m[856]&~m[1773]&m[1775]&m[1776]&~m[1777])|(~m[856]&m[1773]&~m[1775]&~m[1776]&m[1777])|(~m[856]&~m[1773]&m[1775]&~m[1776]&m[1777])|(m[856]&m[1773]&m[1775]&~m[1776]&m[1777])|(~m[856]&m[1773]&m[1775]&m[1776]&m[1777]))&UnbiasedRNG[665])|((m[856]&~m[1773]&~m[1775]&m[1776]&~m[1777])|(~m[856]&~m[1773]&~m[1775]&~m[1776]&m[1777])|(m[856]&~m[1773]&~m[1775]&~m[1776]&m[1777])|(m[856]&m[1773]&~m[1775]&~m[1776]&m[1777])|(m[856]&~m[1773]&m[1775]&~m[1776]&m[1777])|(~m[856]&~m[1773]&~m[1775]&m[1776]&m[1777])|(m[856]&~m[1773]&~m[1775]&m[1776]&m[1777])|(~m[856]&m[1773]&~m[1775]&m[1776]&m[1777])|(m[856]&m[1773]&~m[1775]&m[1776]&m[1777])|(~m[856]&~m[1773]&m[1775]&m[1776]&m[1777])|(m[856]&~m[1773]&m[1775]&m[1776]&m[1777])|(m[856]&m[1773]&m[1775]&m[1776]&m[1777]))):InitCond[1560];
    m[1779] = run?((((m[871]&~m[1778]&~m[1780]&~m[1781]&~m[1782])|(~m[871]&~m[1778]&~m[1780]&m[1781]&~m[1782])|(m[871]&m[1778]&~m[1780]&m[1781]&~m[1782])|(m[871]&~m[1778]&m[1780]&m[1781]&~m[1782])|(~m[871]&m[1778]&~m[1780]&~m[1781]&m[1782])|(~m[871]&~m[1778]&m[1780]&~m[1781]&m[1782])|(m[871]&m[1778]&m[1780]&~m[1781]&m[1782])|(~m[871]&m[1778]&m[1780]&m[1781]&m[1782]))&UnbiasedRNG[666])|((m[871]&~m[1778]&~m[1780]&m[1781]&~m[1782])|(~m[871]&~m[1778]&~m[1780]&~m[1781]&m[1782])|(m[871]&~m[1778]&~m[1780]&~m[1781]&m[1782])|(m[871]&m[1778]&~m[1780]&~m[1781]&m[1782])|(m[871]&~m[1778]&m[1780]&~m[1781]&m[1782])|(~m[871]&~m[1778]&~m[1780]&m[1781]&m[1782])|(m[871]&~m[1778]&~m[1780]&m[1781]&m[1782])|(~m[871]&m[1778]&~m[1780]&m[1781]&m[1782])|(m[871]&m[1778]&~m[1780]&m[1781]&m[1782])|(~m[871]&~m[1778]&m[1780]&m[1781]&m[1782])|(m[871]&~m[1778]&m[1780]&m[1781]&m[1782])|(m[871]&m[1778]&m[1780]&m[1781]&m[1782]))):InitCond[1561];
    m[1784] = run?((((m[886]&~m[1783]&~m[1785]&~m[1786]&~m[1787])|(~m[886]&~m[1783]&~m[1785]&m[1786]&~m[1787])|(m[886]&m[1783]&~m[1785]&m[1786]&~m[1787])|(m[886]&~m[1783]&m[1785]&m[1786]&~m[1787])|(~m[886]&m[1783]&~m[1785]&~m[1786]&m[1787])|(~m[886]&~m[1783]&m[1785]&~m[1786]&m[1787])|(m[886]&m[1783]&m[1785]&~m[1786]&m[1787])|(~m[886]&m[1783]&m[1785]&m[1786]&m[1787]))&UnbiasedRNG[667])|((m[886]&~m[1783]&~m[1785]&m[1786]&~m[1787])|(~m[886]&~m[1783]&~m[1785]&~m[1786]&m[1787])|(m[886]&~m[1783]&~m[1785]&~m[1786]&m[1787])|(m[886]&m[1783]&~m[1785]&~m[1786]&m[1787])|(m[886]&~m[1783]&m[1785]&~m[1786]&m[1787])|(~m[886]&~m[1783]&~m[1785]&m[1786]&m[1787])|(m[886]&~m[1783]&~m[1785]&m[1786]&m[1787])|(~m[886]&m[1783]&~m[1785]&m[1786]&m[1787])|(m[886]&m[1783]&~m[1785]&m[1786]&m[1787])|(~m[886]&~m[1783]&m[1785]&m[1786]&m[1787])|(m[886]&~m[1783]&m[1785]&m[1786]&m[1787])|(m[886]&m[1783]&m[1785]&m[1786]&m[1787]))):InitCond[1562];
    m[1789] = run?((((m[901]&~m[1788]&~m[1790]&~m[1791]&~m[1792])|(~m[901]&~m[1788]&~m[1790]&m[1791]&~m[1792])|(m[901]&m[1788]&~m[1790]&m[1791]&~m[1792])|(m[901]&~m[1788]&m[1790]&m[1791]&~m[1792])|(~m[901]&m[1788]&~m[1790]&~m[1791]&m[1792])|(~m[901]&~m[1788]&m[1790]&~m[1791]&m[1792])|(m[901]&m[1788]&m[1790]&~m[1791]&m[1792])|(~m[901]&m[1788]&m[1790]&m[1791]&m[1792]))&UnbiasedRNG[668])|((m[901]&~m[1788]&~m[1790]&m[1791]&~m[1792])|(~m[901]&~m[1788]&~m[1790]&~m[1791]&m[1792])|(m[901]&~m[1788]&~m[1790]&~m[1791]&m[1792])|(m[901]&m[1788]&~m[1790]&~m[1791]&m[1792])|(m[901]&~m[1788]&m[1790]&~m[1791]&m[1792])|(~m[901]&~m[1788]&~m[1790]&m[1791]&m[1792])|(m[901]&~m[1788]&~m[1790]&m[1791]&m[1792])|(~m[901]&m[1788]&~m[1790]&m[1791]&m[1792])|(m[901]&m[1788]&~m[1790]&m[1791]&m[1792])|(~m[901]&~m[1788]&m[1790]&m[1791]&m[1792])|(m[901]&~m[1788]&m[1790]&m[1791]&m[1792])|(m[901]&m[1788]&m[1790]&m[1791]&m[1792]))):InitCond[1563];
    m[1794] = run?((((m[916]&~m[1793]&~m[1795]&~m[1796]&~m[1797])|(~m[916]&~m[1793]&~m[1795]&m[1796]&~m[1797])|(m[916]&m[1793]&~m[1795]&m[1796]&~m[1797])|(m[916]&~m[1793]&m[1795]&m[1796]&~m[1797])|(~m[916]&m[1793]&~m[1795]&~m[1796]&m[1797])|(~m[916]&~m[1793]&m[1795]&~m[1796]&m[1797])|(m[916]&m[1793]&m[1795]&~m[1796]&m[1797])|(~m[916]&m[1793]&m[1795]&m[1796]&m[1797]))&UnbiasedRNG[669])|((m[916]&~m[1793]&~m[1795]&m[1796]&~m[1797])|(~m[916]&~m[1793]&~m[1795]&~m[1796]&m[1797])|(m[916]&~m[1793]&~m[1795]&~m[1796]&m[1797])|(m[916]&m[1793]&~m[1795]&~m[1796]&m[1797])|(m[916]&~m[1793]&m[1795]&~m[1796]&m[1797])|(~m[916]&~m[1793]&~m[1795]&m[1796]&m[1797])|(m[916]&~m[1793]&~m[1795]&m[1796]&m[1797])|(~m[916]&m[1793]&~m[1795]&m[1796]&m[1797])|(m[916]&m[1793]&~m[1795]&m[1796]&m[1797])|(~m[916]&~m[1793]&m[1795]&m[1796]&m[1797])|(m[916]&~m[1793]&m[1795]&m[1796]&m[1797])|(m[916]&m[1793]&m[1795]&m[1796]&m[1797]))):InitCond[1564];
    m[1799] = run?((((m[767]&~m[1798]&~m[1800]&~m[1801]&~m[1802])|(~m[767]&~m[1798]&~m[1800]&m[1801]&~m[1802])|(m[767]&m[1798]&~m[1800]&m[1801]&~m[1802])|(m[767]&~m[1798]&m[1800]&m[1801]&~m[1802])|(~m[767]&m[1798]&~m[1800]&~m[1801]&m[1802])|(~m[767]&~m[1798]&m[1800]&~m[1801]&m[1802])|(m[767]&m[1798]&m[1800]&~m[1801]&m[1802])|(~m[767]&m[1798]&m[1800]&m[1801]&m[1802]))&UnbiasedRNG[670])|((m[767]&~m[1798]&~m[1800]&m[1801]&~m[1802])|(~m[767]&~m[1798]&~m[1800]&~m[1801]&m[1802])|(m[767]&~m[1798]&~m[1800]&~m[1801]&m[1802])|(m[767]&m[1798]&~m[1800]&~m[1801]&m[1802])|(m[767]&~m[1798]&m[1800]&~m[1801]&m[1802])|(~m[767]&~m[1798]&~m[1800]&m[1801]&m[1802])|(m[767]&~m[1798]&~m[1800]&m[1801]&m[1802])|(~m[767]&m[1798]&~m[1800]&m[1801]&m[1802])|(m[767]&m[1798]&~m[1800]&m[1801]&m[1802])|(~m[767]&~m[1798]&m[1800]&m[1801]&m[1802])|(m[767]&~m[1798]&m[1800]&m[1801]&m[1802])|(m[767]&m[1798]&m[1800]&m[1801]&m[1802]))):InitCond[1565];
    m[1804] = run?((((m[782]&~m[1803]&~m[1805]&~m[1806]&~m[1807])|(~m[782]&~m[1803]&~m[1805]&m[1806]&~m[1807])|(m[782]&m[1803]&~m[1805]&m[1806]&~m[1807])|(m[782]&~m[1803]&m[1805]&m[1806]&~m[1807])|(~m[782]&m[1803]&~m[1805]&~m[1806]&m[1807])|(~m[782]&~m[1803]&m[1805]&~m[1806]&m[1807])|(m[782]&m[1803]&m[1805]&~m[1806]&m[1807])|(~m[782]&m[1803]&m[1805]&m[1806]&m[1807]))&UnbiasedRNG[671])|((m[782]&~m[1803]&~m[1805]&m[1806]&~m[1807])|(~m[782]&~m[1803]&~m[1805]&~m[1806]&m[1807])|(m[782]&~m[1803]&~m[1805]&~m[1806]&m[1807])|(m[782]&m[1803]&~m[1805]&~m[1806]&m[1807])|(m[782]&~m[1803]&m[1805]&~m[1806]&m[1807])|(~m[782]&~m[1803]&~m[1805]&m[1806]&m[1807])|(m[782]&~m[1803]&~m[1805]&m[1806]&m[1807])|(~m[782]&m[1803]&~m[1805]&m[1806]&m[1807])|(m[782]&m[1803]&~m[1805]&m[1806]&m[1807])|(~m[782]&~m[1803]&m[1805]&m[1806]&m[1807])|(m[782]&~m[1803]&m[1805]&m[1806]&m[1807])|(m[782]&m[1803]&m[1805]&m[1806]&m[1807]))):InitCond[1566];
    m[1809] = run?((((m[797]&~m[1808]&~m[1810]&~m[1811]&~m[1812])|(~m[797]&~m[1808]&~m[1810]&m[1811]&~m[1812])|(m[797]&m[1808]&~m[1810]&m[1811]&~m[1812])|(m[797]&~m[1808]&m[1810]&m[1811]&~m[1812])|(~m[797]&m[1808]&~m[1810]&~m[1811]&m[1812])|(~m[797]&~m[1808]&m[1810]&~m[1811]&m[1812])|(m[797]&m[1808]&m[1810]&~m[1811]&m[1812])|(~m[797]&m[1808]&m[1810]&m[1811]&m[1812]))&UnbiasedRNG[672])|((m[797]&~m[1808]&~m[1810]&m[1811]&~m[1812])|(~m[797]&~m[1808]&~m[1810]&~m[1811]&m[1812])|(m[797]&~m[1808]&~m[1810]&~m[1811]&m[1812])|(m[797]&m[1808]&~m[1810]&~m[1811]&m[1812])|(m[797]&~m[1808]&m[1810]&~m[1811]&m[1812])|(~m[797]&~m[1808]&~m[1810]&m[1811]&m[1812])|(m[797]&~m[1808]&~m[1810]&m[1811]&m[1812])|(~m[797]&m[1808]&~m[1810]&m[1811]&m[1812])|(m[797]&m[1808]&~m[1810]&m[1811]&m[1812])|(~m[797]&~m[1808]&m[1810]&m[1811]&m[1812])|(m[797]&~m[1808]&m[1810]&m[1811]&m[1812])|(m[797]&m[1808]&m[1810]&m[1811]&m[1812]))):InitCond[1567];
    m[1814] = run?((((m[812]&~m[1813]&~m[1815]&~m[1816]&~m[1817])|(~m[812]&~m[1813]&~m[1815]&m[1816]&~m[1817])|(m[812]&m[1813]&~m[1815]&m[1816]&~m[1817])|(m[812]&~m[1813]&m[1815]&m[1816]&~m[1817])|(~m[812]&m[1813]&~m[1815]&~m[1816]&m[1817])|(~m[812]&~m[1813]&m[1815]&~m[1816]&m[1817])|(m[812]&m[1813]&m[1815]&~m[1816]&m[1817])|(~m[812]&m[1813]&m[1815]&m[1816]&m[1817]))&UnbiasedRNG[673])|((m[812]&~m[1813]&~m[1815]&m[1816]&~m[1817])|(~m[812]&~m[1813]&~m[1815]&~m[1816]&m[1817])|(m[812]&~m[1813]&~m[1815]&~m[1816]&m[1817])|(m[812]&m[1813]&~m[1815]&~m[1816]&m[1817])|(m[812]&~m[1813]&m[1815]&~m[1816]&m[1817])|(~m[812]&~m[1813]&~m[1815]&m[1816]&m[1817])|(m[812]&~m[1813]&~m[1815]&m[1816]&m[1817])|(~m[812]&m[1813]&~m[1815]&m[1816]&m[1817])|(m[812]&m[1813]&~m[1815]&m[1816]&m[1817])|(~m[812]&~m[1813]&m[1815]&m[1816]&m[1817])|(m[812]&~m[1813]&m[1815]&m[1816]&m[1817])|(m[812]&m[1813]&m[1815]&m[1816]&m[1817]))):InitCond[1568];
    m[1819] = run?((((m[827]&~m[1818]&~m[1820]&~m[1821]&~m[1822])|(~m[827]&~m[1818]&~m[1820]&m[1821]&~m[1822])|(m[827]&m[1818]&~m[1820]&m[1821]&~m[1822])|(m[827]&~m[1818]&m[1820]&m[1821]&~m[1822])|(~m[827]&m[1818]&~m[1820]&~m[1821]&m[1822])|(~m[827]&~m[1818]&m[1820]&~m[1821]&m[1822])|(m[827]&m[1818]&m[1820]&~m[1821]&m[1822])|(~m[827]&m[1818]&m[1820]&m[1821]&m[1822]))&UnbiasedRNG[674])|((m[827]&~m[1818]&~m[1820]&m[1821]&~m[1822])|(~m[827]&~m[1818]&~m[1820]&~m[1821]&m[1822])|(m[827]&~m[1818]&~m[1820]&~m[1821]&m[1822])|(m[827]&m[1818]&~m[1820]&~m[1821]&m[1822])|(m[827]&~m[1818]&m[1820]&~m[1821]&m[1822])|(~m[827]&~m[1818]&~m[1820]&m[1821]&m[1822])|(m[827]&~m[1818]&~m[1820]&m[1821]&m[1822])|(~m[827]&m[1818]&~m[1820]&m[1821]&m[1822])|(m[827]&m[1818]&~m[1820]&m[1821]&m[1822])|(~m[827]&~m[1818]&m[1820]&m[1821]&m[1822])|(m[827]&~m[1818]&m[1820]&m[1821]&m[1822])|(m[827]&m[1818]&m[1820]&m[1821]&m[1822]))):InitCond[1569];
    m[1824] = run?((((m[842]&~m[1823]&~m[1825]&~m[1826]&~m[1827])|(~m[842]&~m[1823]&~m[1825]&m[1826]&~m[1827])|(m[842]&m[1823]&~m[1825]&m[1826]&~m[1827])|(m[842]&~m[1823]&m[1825]&m[1826]&~m[1827])|(~m[842]&m[1823]&~m[1825]&~m[1826]&m[1827])|(~m[842]&~m[1823]&m[1825]&~m[1826]&m[1827])|(m[842]&m[1823]&m[1825]&~m[1826]&m[1827])|(~m[842]&m[1823]&m[1825]&m[1826]&m[1827]))&UnbiasedRNG[675])|((m[842]&~m[1823]&~m[1825]&m[1826]&~m[1827])|(~m[842]&~m[1823]&~m[1825]&~m[1826]&m[1827])|(m[842]&~m[1823]&~m[1825]&~m[1826]&m[1827])|(m[842]&m[1823]&~m[1825]&~m[1826]&m[1827])|(m[842]&~m[1823]&m[1825]&~m[1826]&m[1827])|(~m[842]&~m[1823]&~m[1825]&m[1826]&m[1827])|(m[842]&~m[1823]&~m[1825]&m[1826]&m[1827])|(~m[842]&m[1823]&~m[1825]&m[1826]&m[1827])|(m[842]&m[1823]&~m[1825]&m[1826]&m[1827])|(~m[842]&~m[1823]&m[1825]&m[1826]&m[1827])|(m[842]&~m[1823]&m[1825]&m[1826]&m[1827])|(m[842]&m[1823]&m[1825]&m[1826]&m[1827]))):InitCond[1570];
    m[1829] = run?((((m[857]&~m[1828]&~m[1830]&~m[1831]&~m[1832])|(~m[857]&~m[1828]&~m[1830]&m[1831]&~m[1832])|(m[857]&m[1828]&~m[1830]&m[1831]&~m[1832])|(m[857]&~m[1828]&m[1830]&m[1831]&~m[1832])|(~m[857]&m[1828]&~m[1830]&~m[1831]&m[1832])|(~m[857]&~m[1828]&m[1830]&~m[1831]&m[1832])|(m[857]&m[1828]&m[1830]&~m[1831]&m[1832])|(~m[857]&m[1828]&m[1830]&m[1831]&m[1832]))&UnbiasedRNG[676])|((m[857]&~m[1828]&~m[1830]&m[1831]&~m[1832])|(~m[857]&~m[1828]&~m[1830]&~m[1831]&m[1832])|(m[857]&~m[1828]&~m[1830]&~m[1831]&m[1832])|(m[857]&m[1828]&~m[1830]&~m[1831]&m[1832])|(m[857]&~m[1828]&m[1830]&~m[1831]&m[1832])|(~m[857]&~m[1828]&~m[1830]&m[1831]&m[1832])|(m[857]&~m[1828]&~m[1830]&m[1831]&m[1832])|(~m[857]&m[1828]&~m[1830]&m[1831]&m[1832])|(m[857]&m[1828]&~m[1830]&m[1831]&m[1832])|(~m[857]&~m[1828]&m[1830]&m[1831]&m[1832])|(m[857]&~m[1828]&m[1830]&m[1831]&m[1832])|(m[857]&m[1828]&m[1830]&m[1831]&m[1832]))):InitCond[1571];
    m[1834] = run?((((m[872]&~m[1833]&~m[1835]&~m[1836]&~m[1837])|(~m[872]&~m[1833]&~m[1835]&m[1836]&~m[1837])|(m[872]&m[1833]&~m[1835]&m[1836]&~m[1837])|(m[872]&~m[1833]&m[1835]&m[1836]&~m[1837])|(~m[872]&m[1833]&~m[1835]&~m[1836]&m[1837])|(~m[872]&~m[1833]&m[1835]&~m[1836]&m[1837])|(m[872]&m[1833]&m[1835]&~m[1836]&m[1837])|(~m[872]&m[1833]&m[1835]&m[1836]&m[1837]))&UnbiasedRNG[677])|((m[872]&~m[1833]&~m[1835]&m[1836]&~m[1837])|(~m[872]&~m[1833]&~m[1835]&~m[1836]&m[1837])|(m[872]&~m[1833]&~m[1835]&~m[1836]&m[1837])|(m[872]&m[1833]&~m[1835]&~m[1836]&m[1837])|(m[872]&~m[1833]&m[1835]&~m[1836]&m[1837])|(~m[872]&~m[1833]&~m[1835]&m[1836]&m[1837])|(m[872]&~m[1833]&~m[1835]&m[1836]&m[1837])|(~m[872]&m[1833]&~m[1835]&m[1836]&m[1837])|(m[872]&m[1833]&~m[1835]&m[1836]&m[1837])|(~m[872]&~m[1833]&m[1835]&m[1836]&m[1837])|(m[872]&~m[1833]&m[1835]&m[1836]&m[1837])|(m[872]&m[1833]&m[1835]&m[1836]&m[1837]))):InitCond[1572];
    m[1839] = run?((((m[887]&~m[1838]&~m[1840]&~m[1841]&~m[1842])|(~m[887]&~m[1838]&~m[1840]&m[1841]&~m[1842])|(m[887]&m[1838]&~m[1840]&m[1841]&~m[1842])|(m[887]&~m[1838]&m[1840]&m[1841]&~m[1842])|(~m[887]&m[1838]&~m[1840]&~m[1841]&m[1842])|(~m[887]&~m[1838]&m[1840]&~m[1841]&m[1842])|(m[887]&m[1838]&m[1840]&~m[1841]&m[1842])|(~m[887]&m[1838]&m[1840]&m[1841]&m[1842]))&UnbiasedRNG[678])|((m[887]&~m[1838]&~m[1840]&m[1841]&~m[1842])|(~m[887]&~m[1838]&~m[1840]&~m[1841]&m[1842])|(m[887]&~m[1838]&~m[1840]&~m[1841]&m[1842])|(m[887]&m[1838]&~m[1840]&~m[1841]&m[1842])|(m[887]&~m[1838]&m[1840]&~m[1841]&m[1842])|(~m[887]&~m[1838]&~m[1840]&m[1841]&m[1842])|(m[887]&~m[1838]&~m[1840]&m[1841]&m[1842])|(~m[887]&m[1838]&~m[1840]&m[1841]&m[1842])|(m[887]&m[1838]&~m[1840]&m[1841]&m[1842])|(~m[887]&~m[1838]&m[1840]&m[1841]&m[1842])|(m[887]&~m[1838]&m[1840]&m[1841]&m[1842])|(m[887]&m[1838]&m[1840]&m[1841]&m[1842]))):InitCond[1573];
    m[1844] = run?((((m[902]&~m[1843]&~m[1845]&~m[1846]&~m[1847])|(~m[902]&~m[1843]&~m[1845]&m[1846]&~m[1847])|(m[902]&m[1843]&~m[1845]&m[1846]&~m[1847])|(m[902]&~m[1843]&m[1845]&m[1846]&~m[1847])|(~m[902]&m[1843]&~m[1845]&~m[1846]&m[1847])|(~m[902]&~m[1843]&m[1845]&~m[1846]&m[1847])|(m[902]&m[1843]&m[1845]&~m[1846]&m[1847])|(~m[902]&m[1843]&m[1845]&m[1846]&m[1847]))&UnbiasedRNG[679])|((m[902]&~m[1843]&~m[1845]&m[1846]&~m[1847])|(~m[902]&~m[1843]&~m[1845]&~m[1846]&m[1847])|(m[902]&~m[1843]&~m[1845]&~m[1846]&m[1847])|(m[902]&m[1843]&~m[1845]&~m[1846]&m[1847])|(m[902]&~m[1843]&m[1845]&~m[1846]&m[1847])|(~m[902]&~m[1843]&~m[1845]&m[1846]&m[1847])|(m[902]&~m[1843]&~m[1845]&m[1846]&m[1847])|(~m[902]&m[1843]&~m[1845]&m[1846]&m[1847])|(m[902]&m[1843]&~m[1845]&m[1846]&m[1847])|(~m[902]&~m[1843]&m[1845]&m[1846]&m[1847])|(m[902]&~m[1843]&m[1845]&m[1846]&m[1847])|(m[902]&m[1843]&m[1845]&m[1846]&m[1847]))):InitCond[1574];
    m[1849] = run?((((m[917]&~m[1848]&~m[1850]&~m[1851]&~m[1852])|(~m[917]&~m[1848]&~m[1850]&m[1851]&~m[1852])|(m[917]&m[1848]&~m[1850]&m[1851]&~m[1852])|(m[917]&~m[1848]&m[1850]&m[1851]&~m[1852])|(~m[917]&m[1848]&~m[1850]&~m[1851]&m[1852])|(~m[917]&~m[1848]&m[1850]&~m[1851]&m[1852])|(m[917]&m[1848]&m[1850]&~m[1851]&m[1852])|(~m[917]&m[1848]&m[1850]&m[1851]&m[1852]))&UnbiasedRNG[680])|((m[917]&~m[1848]&~m[1850]&m[1851]&~m[1852])|(~m[917]&~m[1848]&~m[1850]&~m[1851]&m[1852])|(m[917]&~m[1848]&~m[1850]&~m[1851]&m[1852])|(m[917]&m[1848]&~m[1850]&~m[1851]&m[1852])|(m[917]&~m[1848]&m[1850]&~m[1851]&m[1852])|(~m[917]&~m[1848]&~m[1850]&m[1851]&m[1852])|(m[917]&~m[1848]&~m[1850]&m[1851]&m[1852])|(~m[917]&m[1848]&~m[1850]&m[1851]&m[1852])|(m[917]&m[1848]&~m[1850]&m[1851]&m[1852])|(~m[917]&~m[1848]&m[1850]&m[1851]&m[1852])|(m[917]&~m[1848]&m[1850]&m[1851]&m[1852])|(m[917]&m[1848]&m[1850]&m[1851]&m[1852]))):InitCond[1575];
    m[1854] = run?((((m[783]&~m[1853]&~m[1855]&~m[1856]&~m[1857])|(~m[783]&~m[1853]&~m[1855]&m[1856]&~m[1857])|(m[783]&m[1853]&~m[1855]&m[1856]&~m[1857])|(m[783]&~m[1853]&m[1855]&m[1856]&~m[1857])|(~m[783]&m[1853]&~m[1855]&~m[1856]&m[1857])|(~m[783]&~m[1853]&m[1855]&~m[1856]&m[1857])|(m[783]&m[1853]&m[1855]&~m[1856]&m[1857])|(~m[783]&m[1853]&m[1855]&m[1856]&m[1857]))&UnbiasedRNG[681])|((m[783]&~m[1853]&~m[1855]&m[1856]&~m[1857])|(~m[783]&~m[1853]&~m[1855]&~m[1856]&m[1857])|(m[783]&~m[1853]&~m[1855]&~m[1856]&m[1857])|(m[783]&m[1853]&~m[1855]&~m[1856]&m[1857])|(m[783]&~m[1853]&m[1855]&~m[1856]&m[1857])|(~m[783]&~m[1853]&~m[1855]&m[1856]&m[1857])|(m[783]&~m[1853]&~m[1855]&m[1856]&m[1857])|(~m[783]&m[1853]&~m[1855]&m[1856]&m[1857])|(m[783]&m[1853]&~m[1855]&m[1856]&m[1857])|(~m[783]&~m[1853]&m[1855]&m[1856]&m[1857])|(m[783]&~m[1853]&m[1855]&m[1856]&m[1857])|(m[783]&m[1853]&m[1855]&m[1856]&m[1857]))):InitCond[1576];
    m[1859] = run?((((m[798]&~m[1858]&~m[1860]&~m[1861]&~m[1862])|(~m[798]&~m[1858]&~m[1860]&m[1861]&~m[1862])|(m[798]&m[1858]&~m[1860]&m[1861]&~m[1862])|(m[798]&~m[1858]&m[1860]&m[1861]&~m[1862])|(~m[798]&m[1858]&~m[1860]&~m[1861]&m[1862])|(~m[798]&~m[1858]&m[1860]&~m[1861]&m[1862])|(m[798]&m[1858]&m[1860]&~m[1861]&m[1862])|(~m[798]&m[1858]&m[1860]&m[1861]&m[1862]))&UnbiasedRNG[682])|((m[798]&~m[1858]&~m[1860]&m[1861]&~m[1862])|(~m[798]&~m[1858]&~m[1860]&~m[1861]&m[1862])|(m[798]&~m[1858]&~m[1860]&~m[1861]&m[1862])|(m[798]&m[1858]&~m[1860]&~m[1861]&m[1862])|(m[798]&~m[1858]&m[1860]&~m[1861]&m[1862])|(~m[798]&~m[1858]&~m[1860]&m[1861]&m[1862])|(m[798]&~m[1858]&~m[1860]&m[1861]&m[1862])|(~m[798]&m[1858]&~m[1860]&m[1861]&m[1862])|(m[798]&m[1858]&~m[1860]&m[1861]&m[1862])|(~m[798]&~m[1858]&m[1860]&m[1861]&m[1862])|(m[798]&~m[1858]&m[1860]&m[1861]&m[1862])|(m[798]&m[1858]&m[1860]&m[1861]&m[1862]))):InitCond[1577];
    m[1864] = run?((((m[813]&~m[1863]&~m[1865]&~m[1866]&~m[1867])|(~m[813]&~m[1863]&~m[1865]&m[1866]&~m[1867])|(m[813]&m[1863]&~m[1865]&m[1866]&~m[1867])|(m[813]&~m[1863]&m[1865]&m[1866]&~m[1867])|(~m[813]&m[1863]&~m[1865]&~m[1866]&m[1867])|(~m[813]&~m[1863]&m[1865]&~m[1866]&m[1867])|(m[813]&m[1863]&m[1865]&~m[1866]&m[1867])|(~m[813]&m[1863]&m[1865]&m[1866]&m[1867]))&UnbiasedRNG[683])|((m[813]&~m[1863]&~m[1865]&m[1866]&~m[1867])|(~m[813]&~m[1863]&~m[1865]&~m[1866]&m[1867])|(m[813]&~m[1863]&~m[1865]&~m[1866]&m[1867])|(m[813]&m[1863]&~m[1865]&~m[1866]&m[1867])|(m[813]&~m[1863]&m[1865]&~m[1866]&m[1867])|(~m[813]&~m[1863]&~m[1865]&m[1866]&m[1867])|(m[813]&~m[1863]&~m[1865]&m[1866]&m[1867])|(~m[813]&m[1863]&~m[1865]&m[1866]&m[1867])|(m[813]&m[1863]&~m[1865]&m[1866]&m[1867])|(~m[813]&~m[1863]&m[1865]&m[1866]&m[1867])|(m[813]&~m[1863]&m[1865]&m[1866]&m[1867])|(m[813]&m[1863]&m[1865]&m[1866]&m[1867]))):InitCond[1578];
    m[1869] = run?((((m[828]&~m[1868]&~m[1870]&~m[1871]&~m[1872])|(~m[828]&~m[1868]&~m[1870]&m[1871]&~m[1872])|(m[828]&m[1868]&~m[1870]&m[1871]&~m[1872])|(m[828]&~m[1868]&m[1870]&m[1871]&~m[1872])|(~m[828]&m[1868]&~m[1870]&~m[1871]&m[1872])|(~m[828]&~m[1868]&m[1870]&~m[1871]&m[1872])|(m[828]&m[1868]&m[1870]&~m[1871]&m[1872])|(~m[828]&m[1868]&m[1870]&m[1871]&m[1872]))&UnbiasedRNG[684])|((m[828]&~m[1868]&~m[1870]&m[1871]&~m[1872])|(~m[828]&~m[1868]&~m[1870]&~m[1871]&m[1872])|(m[828]&~m[1868]&~m[1870]&~m[1871]&m[1872])|(m[828]&m[1868]&~m[1870]&~m[1871]&m[1872])|(m[828]&~m[1868]&m[1870]&~m[1871]&m[1872])|(~m[828]&~m[1868]&~m[1870]&m[1871]&m[1872])|(m[828]&~m[1868]&~m[1870]&m[1871]&m[1872])|(~m[828]&m[1868]&~m[1870]&m[1871]&m[1872])|(m[828]&m[1868]&~m[1870]&m[1871]&m[1872])|(~m[828]&~m[1868]&m[1870]&m[1871]&m[1872])|(m[828]&~m[1868]&m[1870]&m[1871]&m[1872])|(m[828]&m[1868]&m[1870]&m[1871]&m[1872]))):InitCond[1579];
    m[1874] = run?((((m[843]&~m[1873]&~m[1875]&~m[1876]&~m[1877])|(~m[843]&~m[1873]&~m[1875]&m[1876]&~m[1877])|(m[843]&m[1873]&~m[1875]&m[1876]&~m[1877])|(m[843]&~m[1873]&m[1875]&m[1876]&~m[1877])|(~m[843]&m[1873]&~m[1875]&~m[1876]&m[1877])|(~m[843]&~m[1873]&m[1875]&~m[1876]&m[1877])|(m[843]&m[1873]&m[1875]&~m[1876]&m[1877])|(~m[843]&m[1873]&m[1875]&m[1876]&m[1877]))&UnbiasedRNG[685])|((m[843]&~m[1873]&~m[1875]&m[1876]&~m[1877])|(~m[843]&~m[1873]&~m[1875]&~m[1876]&m[1877])|(m[843]&~m[1873]&~m[1875]&~m[1876]&m[1877])|(m[843]&m[1873]&~m[1875]&~m[1876]&m[1877])|(m[843]&~m[1873]&m[1875]&~m[1876]&m[1877])|(~m[843]&~m[1873]&~m[1875]&m[1876]&m[1877])|(m[843]&~m[1873]&~m[1875]&m[1876]&m[1877])|(~m[843]&m[1873]&~m[1875]&m[1876]&m[1877])|(m[843]&m[1873]&~m[1875]&m[1876]&m[1877])|(~m[843]&~m[1873]&m[1875]&m[1876]&m[1877])|(m[843]&~m[1873]&m[1875]&m[1876]&m[1877])|(m[843]&m[1873]&m[1875]&m[1876]&m[1877]))):InitCond[1580];
    m[1879] = run?((((m[858]&~m[1878]&~m[1880]&~m[1881]&~m[1882])|(~m[858]&~m[1878]&~m[1880]&m[1881]&~m[1882])|(m[858]&m[1878]&~m[1880]&m[1881]&~m[1882])|(m[858]&~m[1878]&m[1880]&m[1881]&~m[1882])|(~m[858]&m[1878]&~m[1880]&~m[1881]&m[1882])|(~m[858]&~m[1878]&m[1880]&~m[1881]&m[1882])|(m[858]&m[1878]&m[1880]&~m[1881]&m[1882])|(~m[858]&m[1878]&m[1880]&m[1881]&m[1882]))&UnbiasedRNG[686])|((m[858]&~m[1878]&~m[1880]&m[1881]&~m[1882])|(~m[858]&~m[1878]&~m[1880]&~m[1881]&m[1882])|(m[858]&~m[1878]&~m[1880]&~m[1881]&m[1882])|(m[858]&m[1878]&~m[1880]&~m[1881]&m[1882])|(m[858]&~m[1878]&m[1880]&~m[1881]&m[1882])|(~m[858]&~m[1878]&~m[1880]&m[1881]&m[1882])|(m[858]&~m[1878]&~m[1880]&m[1881]&m[1882])|(~m[858]&m[1878]&~m[1880]&m[1881]&m[1882])|(m[858]&m[1878]&~m[1880]&m[1881]&m[1882])|(~m[858]&~m[1878]&m[1880]&m[1881]&m[1882])|(m[858]&~m[1878]&m[1880]&m[1881]&m[1882])|(m[858]&m[1878]&m[1880]&m[1881]&m[1882]))):InitCond[1581];
    m[1884] = run?((((m[873]&~m[1883]&~m[1885]&~m[1886]&~m[1887])|(~m[873]&~m[1883]&~m[1885]&m[1886]&~m[1887])|(m[873]&m[1883]&~m[1885]&m[1886]&~m[1887])|(m[873]&~m[1883]&m[1885]&m[1886]&~m[1887])|(~m[873]&m[1883]&~m[1885]&~m[1886]&m[1887])|(~m[873]&~m[1883]&m[1885]&~m[1886]&m[1887])|(m[873]&m[1883]&m[1885]&~m[1886]&m[1887])|(~m[873]&m[1883]&m[1885]&m[1886]&m[1887]))&UnbiasedRNG[687])|((m[873]&~m[1883]&~m[1885]&m[1886]&~m[1887])|(~m[873]&~m[1883]&~m[1885]&~m[1886]&m[1887])|(m[873]&~m[1883]&~m[1885]&~m[1886]&m[1887])|(m[873]&m[1883]&~m[1885]&~m[1886]&m[1887])|(m[873]&~m[1883]&m[1885]&~m[1886]&m[1887])|(~m[873]&~m[1883]&~m[1885]&m[1886]&m[1887])|(m[873]&~m[1883]&~m[1885]&m[1886]&m[1887])|(~m[873]&m[1883]&~m[1885]&m[1886]&m[1887])|(m[873]&m[1883]&~m[1885]&m[1886]&m[1887])|(~m[873]&~m[1883]&m[1885]&m[1886]&m[1887])|(m[873]&~m[1883]&m[1885]&m[1886]&m[1887])|(m[873]&m[1883]&m[1885]&m[1886]&m[1887]))):InitCond[1582];
    m[1889] = run?((((m[888]&~m[1888]&~m[1890]&~m[1891]&~m[1892])|(~m[888]&~m[1888]&~m[1890]&m[1891]&~m[1892])|(m[888]&m[1888]&~m[1890]&m[1891]&~m[1892])|(m[888]&~m[1888]&m[1890]&m[1891]&~m[1892])|(~m[888]&m[1888]&~m[1890]&~m[1891]&m[1892])|(~m[888]&~m[1888]&m[1890]&~m[1891]&m[1892])|(m[888]&m[1888]&m[1890]&~m[1891]&m[1892])|(~m[888]&m[1888]&m[1890]&m[1891]&m[1892]))&UnbiasedRNG[688])|((m[888]&~m[1888]&~m[1890]&m[1891]&~m[1892])|(~m[888]&~m[1888]&~m[1890]&~m[1891]&m[1892])|(m[888]&~m[1888]&~m[1890]&~m[1891]&m[1892])|(m[888]&m[1888]&~m[1890]&~m[1891]&m[1892])|(m[888]&~m[1888]&m[1890]&~m[1891]&m[1892])|(~m[888]&~m[1888]&~m[1890]&m[1891]&m[1892])|(m[888]&~m[1888]&~m[1890]&m[1891]&m[1892])|(~m[888]&m[1888]&~m[1890]&m[1891]&m[1892])|(m[888]&m[1888]&~m[1890]&m[1891]&m[1892])|(~m[888]&~m[1888]&m[1890]&m[1891]&m[1892])|(m[888]&~m[1888]&m[1890]&m[1891]&m[1892])|(m[888]&m[1888]&m[1890]&m[1891]&m[1892]))):InitCond[1583];
    m[1894] = run?((((m[903]&~m[1893]&~m[1895]&~m[1896]&~m[1897])|(~m[903]&~m[1893]&~m[1895]&m[1896]&~m[1897])|(m[903]&m[1893]&~m[1895]&m[1896]&~m[1897])|(m[903]&~m[1893]&m[1895]&m[1896]&~m[1897])|(~m[903]&m[1893]&~m[1895]&~m[1896]&m[1897])|(~m[903]&~m[1893]&m[1895]&~m[1896]&m[1897])|(m[903]&m[1893]&m[1895]&~m[1896]&m[1897])|(~m[903]&m[1893]&m[1895]&m[1896]&m[1897]))&UnbiasedRNG[689])|((m[903]&~m[1893]&~m[1895]&m[1896]&~m[1897])|(~m[903]&~m[1893]&~m[1895]&~m[1896]&m[1897])|(m[903]&~m[1893]&~m[1895]&~m[1896]&m[1897])|(m[903]&m[1893]&~m[1895]&~m[1896]&m[1897])|(m[903]&~m[1893]&m[1895]&~m[1896]&m[1897])|(~m[903]&~m[1893]&~m[1895]&m[1896]&m[1897])|(m[903]&~m[1893]&~m[1895]&m[1896]&m[1897])|(~m[903]&m[1893]&~m[1895]&m[1896]&m[1897])|(m[903]&m[1893]&~m[1895]&m[1896]&m[1897])|(~m[903]&~m[1893]&m[1895]&m[1896]&m[1897])|(m[903]&~m[1893]&m[1895]&m[1896]&m[1897])|(m[903]&m[1893]&m[1895]&m[1896]&m[1897]))):InitCond[1584];
    m[1899] = run?((((m[918]&~m[1898]&~m[1900]&~m[1901]&~m[1902])|(~m[918]&~m[1898]&~m[1900]&m[1901]&~m[1902])|(m[918]&m[1898]&~m[1900]&m[1901]&~m[1902])|(m[918]&~m[1898]&m[1900]&m[1901]&~m[1902])|(~m[918]&m[1898]&~m[1900]&~m[1901]&m[1902])|(~m[918]&~m[1898]&m[1900]&~m[1901]&m[1902])|(m[918]&m[1898]&m[1900]&~m[1901]&m[1902])|(~m[918]&m[1898]&m[1900]&m[1901]&m[1902]))&UnbiasedRNG[690])|((m[918]&~m[1898]&~m[1900]&m[1901]&~m[1902])|(~m[918]&~m[1898]&~m[1900]&~m[1901]&m[1902])|(m[918]&~m[1898]&~m[1900]&~m[1901]&m[1902])|(m[918]&m[1898]&~m[1900]&~m[1901]&m[1902])|(m[918]&~m[1898]&m[1900]&~m[1901]&m[1902])|(~m[918]&~m[1898]&~m[1900]&m[1901]&m[1902])|(m[918]&~m[1898]&~m[1900]&m[1901]&m[1902])|(~m[918]&m[1898]&~m[1900]&m[1901]&m[1902])|(m[918]&m[1898]&~m[1900]&m[1901]&m[1902])|(~m[918]&~m[1898]&m[1900]&m[1901]&m[1902])|(m[918]&~m[1898]&m[1900]&m[1901]&m[1902])|(m[918]&m[1898]&m[1900]&m[1901]&m[1902]))):InitCond[1585];
    m[1904] = run?((((m[799]&~m[1903]&~m[1905]&~m[1906]&~m[1907])|(~m[799]&~m[1903]&~m[1905]&m[1906]&~m[1907])|(m[799]&m[1903]&~m[1905]&m[1906]&~m[1907])|(m[799]&~m[1903]&m[1905]&m[1906]&~m[1907])|(~m[799]&m[1903]&~m[1905]&~m[1906]&m[1907])|(~m[799]&~m[1903]&m[1905]&~m[1906]&m[1907])|(m[799]&m[1903]&m[1905]&~m[1906]&m[1907])|(~m[799]&m[1903]&m[1905]&m[1906]&m[1907]))&UnbiasedRNG[691])|((m[799]&~m[1903]&~m[1905]&m[1906]&~m[1907])|(~m[799]&~m[1903]&~m[1905]&~m[1906]&m[1907])|(m[799]&~m[1903]&~m[1905]&~m[1906]&m[1907])|(m[799]&m[1903]&~m[1905]&~m[1906]&m[1907])|(m[799]&~m[1903]&m[1905]&~m[1906]&m[1907])|(~m[799]&~m[1903]&~m[1905]&m[1906]&m[1907])|(m[799]&~m[1903]&~m[1905]&m[1906]&m[1907])|(~m[799]&m[1903]&~m[1905]&m[1906]&m[1907])|(m[799]&m[1903]&~m[1905]&m[1906]&m[1907])|(~m[799]&~m[1903]&m[1905]&m[1906]&m[1907])|(m[799]&~m[1903]&m[1905]&m[1906]&m[1907])|(m[799]&m[1903]&m[1905]&m[1906]&m[1907]))):InitCond[1586];
    m[1909] = run?((((m[814]&~m[1908]&~m[1910]&~m[1911]&~m[1912])|(~m[814]&~m[1908]&~m[1910]&m[1911]&~m[1912])|(m[814]&m[1908]&~m[1910]&m[1911]&~m[1912])|(m[814]&~m[1908]&m[1910]&m[1911]&~m[1912])|(~m[814]&m[1908]&~m[1910]&~m[1911]&m[1912])|(~m[814]&~m[1908]&m[1910]&~m[1911]&m[1912])|(m[814]&m[1908]&m[1910]&~m[1911]&m[1912])|(~m[814]&m[1908]&m[1910]&m[1911]&m[1912]))&UnbiasedRNG[692])|((m[814]&~m[1908]&~m[1910]&m[1911]&~m[1912])|(~m[814]&~m[1908]&~m[1910]&~m[1911]&m[1912])|(m[814]&~m[1908]&~m[1910]&~m[1911]&m[1912])|(m[814]&m[1908]&~m[1910]&~m[1911]&m[1912])|(m[814]&~m[1908]&m[1910]&~m[1911]&m[1912])|(~m[814]&~m[1908]&~m[1910]&m[1911]&m[1912])|(m[814]&~m[1908]&~m[1910]&m[1911]&m[1912])|(~m[814]&m[1908]&~m[1910]&m[1911]&m[1912])|(m[814]&m[1908]&~m[1910]&m[1911]&m[1912])|(~m[814]&~m[1908]&m[1910]&m[1911]&m[1912])|(m[814]&~m[1908]&m[1910]&m[1911]&m[1912])|(m[814]&m[1908]&m[1910]&m[1911]&m[1912]))):InitCond[1587];
    m[1914] = run?((((m[829]&~m[1913]&~m[1915]&~m[1916]&~m[1917])|(~m[829]&~m[1913]&~m[1915]&m[1916]&~m[1917])|(m[829]&m[1913]&~m[1915]&m[1916]&~m[1917])|(m[829]&~m[1913]&m[1915]&m[1916]&~m[1917])|(~m[829]&m[1913]&~m[1915]&~m[1916]&m[1917])|(~m[829]&~m[1913]&m[1915]&~m[1916]&m[1917])|(m[829]&m[1913]&m[1915]&~m[1916]&m[1917])|(~m[829]&m[1913]&m[1915]&m[1916]&m[1917]))&UnbiasedRNG[693])|((m[829]&~m[1913]&~m[1915]&m[1916]&~m[1917])|(~m[829]&~m[1913]&~m[1915]&~m[1916]&m[1917])|(m[829]&~m[1913]&~m[1915]&~m[1916]&m[1917])|(m[829]&m[1913]&~m[1915]&~m[1916]&m[1917])|(m[829]&~m[1913]&m[1915]&~m[1916]&m[1917])|(~m[829]&~m[1913]&~m[1915]&m[1916]&m[1917])|(m[829]&~m[1913]&~m[1915]&m[1916]&m[1917])|(~m[829]&m[1913]&~m[1915]&m[1916]&m[1917])|(m[829]&m[1913]&~m[1915]&m[1916]&m[1917])|(~m[829]&~m[1913]&m[1915]&m[1916]&m[1917])|(m[829]&~m[1913]&m[1915]&m[1916]&m[1917])|(m[829]&m[1913]&m[1915]&m[1916]&m[1917]))):InitCond[1588];
    m[1919] = run?((((m[844]&~m[1918]&~m[1920]&~m[1921]&~m[1922])|(~m[844]&~m[1918]&~m[1920]&m[1921]&~m[1922])|(m[844]&m[1918]&~m[1920]&m[1921]&~m[1922])|(m[844]&~m[1918]&m[1920]&m[1921]&~m[1922])|(~m[844]&m[1918]&~m[1920]&~m[1921]&m[1922])|(~m[844]&~m[1918]&m[1920]&~m[1921]&m[1922])|(m[844]&m[1918]&m[1920]&~m[1921]&m[1922])|(~m[844]&m[1918]&m[1920]&m[1921]&m[1922]))&UnbiasedRNG[694])|((m[844]&~m[1918]&~m[1920]&m[1921]&~m[1922])|(~m[844]&~m[1918]&~m[1920]&~m[1921]&m[1922])|(m[844]&~m[1918]&~m[1920]&~m[1921]&m[1922])|(m[844]&m[1918]&~m[1920]&~m[1921]&m[1922])|(m[844]&~m[1918]&m[1920]&~m[1921]&m[1922])|(~m[844]&~m[1918]&~m[1920]&m[1921]&m[1922])|(m[844]&~m[1918]&~m[1920]&m[1921]&m[1922])|(~m[844]&m[1918]&~m[1920]&m[1921]&m[1922])|(m[844]&m[1918]&~m[1920]&m[1921]&m[1922])|(~m[844]&~m[1918]&m[1920]&m[1921]&m[1922])|(m[844]&~m[1918]&m[1920]&m[1921]&m[1922])|(m[844]&m[1918]&m[1920]&m[1921]&m[1922]))):InitCond[1589];
    m[1924] = run?((((m[859]&~m[1923]&~m[1925]&~m[1926]&~m[1927])|(~m[859]&~m[1923]&~m[1925]&m[1926]&~m[1927])|(m[859]&m[1923]&~m[1925]&m[1926]&~m[1927])|(m[859]&~m[1923]&m[1925]&m[1926]&~m[1927])|(~m[859]&m[1923]&~m[1925]&~m[1926]&m[1927])|(~m[859]&~m[1923]&m[1925]&~m[1926]&m[1927])|(m[859]&m[1923]&m[1925]&~m[1926]&m[1927])|(~m[859]&m[1923]&m[1925]&m[1926]&m[1927]))&UnbiasedRNG[695])|((m[859]&~m[1923]&~m[1925]&m[1926]&~m[1927])|(~m[859]&~m[1923]&~m[1925]&~m[1926]&m[1927])|(m[859]&~m[1923]&~m[1925]&~m[1926]&m[1927])|(m[859]&m[1923]&~m[1925]&~m[1926]&m[1927])|(m[859]&~m[1923]&m[1925]&~m[1926]&m[1927])|(~m[859]&~m[1923]&~m[1925]&m[1926]&m[1927])|(m[859]&~m[1923]&~m[1925]&m[1926]&m[1927])|(~m[859]&m[1923]&~m[1925]&m[1926]&m[1927])|(m[859]&m[1923]&~m[1925]&m[1926]&m[1927])|(~m[859]&~m[1923]&m[1925]&m[1926]&m[1927])|(m[859]&~m[1923]&m[1925]&m[1926]&m[1927])|(m[859]&m[1923]&m[1925]&m[1926]&m[1927]))):InitCond[1590];
    m[1929] = run?((((m[874]&~m[1928]&~m[1930]&~m[1931]&~m[1932])|(~m[874]&~m[1928]&~m[1930]&m[1931]&~m[1932])|(m[874]&m[1928]&~m[1930]&m[1931]&~m[1932])|(m[874]&~m[1928]&m[1930]&m[1931]&~m[1932])|(~m[874]&m[1928]&~m[1930]&~m[1931]&m[1932])|(~m[874]&~m[1928]&m[1930]&~m[1931]&m[1932])|(m[874]&m[1928]&m[1930]&~m[1931]&m[1932])|(~m[874]&m[1928]&m[1930]&m[1931]&m[1932]))&UnbiasedRNG[696])|((m[874]&~m[1928]&~m[1930]&m[1931]&~m[1932])|(~m[874]&~m[1928]&~m[1930]&~m[1931]&m[1932])|(m[874]&~m[1928]&~m[1930]&~m[1931]&m[1932])|(m[874]&m[1928]&~m[1930]&~m[1931]&m[1932])|(m[874]&~m[1928]&m[1930]&~m[1931]&m[1932])|(~m[874]&~m[1928]&~m[1930]&m[1931]&m[1932])|(m[874]&~m[1928]&~m[1930]&m[1931]&m[1932])|(~m[874]&m[1928]&~m[1930]&m[1931]&m[1932])|(m[874]&m[1928]&~m[1930]&m[1931]&m[1932])|(~m[874]&~m[1928]&m[1930]&m[1931]&m[1932])|(m[874]&~m[1928]&m[1930]&m[1931]&m[1932])|(m[874]&m[1928]&m[1930]&m[1931]&m[1932]))):InitCond[1591];
    m[1934] = run?((((m[889]&~m[1933]&~m[1935]&~m[1936]&~m[1937])|(~m[889]&~m[1933]&~m[1935]&m[1936]&~m[1937])|(m[889]&m[1933]&~m[1935]&m[1936]&~m[1937])|(m[889]&~m[1933]&m[1935]&m[1936]&~m[1937])|(~m[889]&m[1933]&~m[1935]&~m[1936]&m[1937])|(~m[889]&~m[1933]&m[1935]&~m[1936]&m[1937])|(m[889]&m[1933]&m[1935]&~m[1936]&m[1937])|(~m[889]&m[1933]&m[1935]&m[1936]&m[1937]))&UnbiasedRNG[697])|((m[889]&~m[1933]&~m[1935]&m[1936]&~m[1937])|(~m[889]&~m[1933]&~m[1935]&~m[1936]&m[1937])|(m[889]&~m[1933]&~m[1935]&~m[1936]&m[1937])|(m[889]&m[1933]&~m[1935]&~m[1936]&m[1937])|(m[889]&~m[1933]&m[1935]&~m[1936]&m[1937])|(~m[889]&~m[1933]&~m[1935]&m[1936]&m[1937])|(m[889]&~m[1933]&~m[1935]&m[1936]&m[1937])|(~m[889]&m[1933]&~m[1935]&m[1936]&m[1937])|(m[889]&m[1933]&~m[1935]&m[1936]&m[1937])|(~m[889]&~m[1933]&m[1935]&m[1936]&m[1937])|(m[889]&~m[1933]&m[1935]&m[1936]&m[1937])|(m[889]&m[1933]&m[1935]&m[1936]&m[1937]))):InitCond[1592];
    m[1939] = run?((((m[904]&~m[1938]&~m[1940]&~m[1941]&~m[1942])|(~m[904]&~m[1938]&~m[1940]&m[1941]&~m[1942])|(m[904]&m[1938]&~m[1940]&m[1941]&~m[1942])|(m[904]&~m[1938]&m[1940]&m[1941]&~m[1942])|(~m[904]&m[1938]&~m[1940]&~m[1941]&m[1942])|(~m[904]&~m[1938]&m[1940]&~m[1941]&m[1942])|(m[904]&m[1938]&m[1940]&~m[1941]&m[1942])|(~m[904]&m[1938]&m[1940]&m[1941]&m[1942]))&UnbiasedRNG[698])|((m[904]&~m[1938]&~m[1940]&m[1941]&~m[1942])|(~m[904]&~m[1938]&~m[1940]&~m[1941]&m[1942])|(m[904]&~m[1938]&~m[1940]&~m[1941]&m[1942])|(m[904]&m[1938]&~m[1940]&~m[1941]&m[1942])|(m[904]&~m[1938]&m[1940]&~m[1941]&m[1942])|(~m[904]&~m[1938]&~m[1940]&m[1941]&m[1942])|(m[904]&~m[1938]&~m[1940]&m[1941]&m[1942])|(~m[904]&m[1938]&~m[1940]&m[1941]&m[1942])|(m[904]&m[1938]&~m[1940]&m[1941]&m[1942])|(~m[904]&~m[1938]&m[1940]&m[1941]&m[1942])|(m[904]&~m[1938]&m[1940]&m[1941]&m[1942])|(m[904]&m[1938]&m[1940]&m[1941]&m[1942]))):InitCond[1593];
    m[1944] = run?((((m[919]&~m[1943]&~m[1945]&~m[1946]&~m[1947])|(~m[919]&~m[1943]&~m[1945]&m[1946]&~m[1947])|(m[919]&m[1943]&~m[1945]&m[1946]&~m[1947])|(m[919]&~m[1943]&m[1945]&m[1946]&~m[1947])|(~m[919]&m[1943]&~m[1945]&~m[1946]&m[1947])|(~m[919]&~m[1943]&m[1945]&~m[1946]&m[1947])|(m[919]&m[1943]&m[1945]&~m[1946]&m[1947])|(~m[919]&m[1943]&m[1945]&m[1946]&m[1947]))&UnbiasedRNG[699])|((m[919]&~m[1943]&~m[1945]&m[1946]&~m[1947])|(~m[919]&~m[1943]&~m[1945]&~m[1946]&m[1947])|(m[919]&~m[1943]&~m[1945]&~m[1946]&m[1947])|(m[919]&m[1943]&~m[1945]&~m[1946]&m[1947])|(m[919]&~m[1943]&m[1945]&~m[1946]&m[1947])|(~m[919]&~m[1943]&~m[1945]&m[1946]&m[1947])|(m[919]&~m[1943]&~m[1945]&m[1946]&m[1947])|(~m[919]&m[1943]&~m[1945]&m[1946]&m[1947])|(m[919]&m[1943]&~m[1945]&m[1946]&m[1947])|(~m[919]&~m[1943]&m[1945]&m[1946]&m[1947])|(m[919]&~m[1943]&m[1945]&m[1946]&m[1947])|(m[919]&m[1943]&m[1945]&m[1946]&m[1947]))):InitCond[1594];
    m[1949] = run?((((m[815]&~m[1948]&~m[1950]&~m[1951]&~m[1952])|(~m[815]&~m[1948]&~m[1950]&m[1951]&~m[1952])|(m[815]&m[1948]&~m[1950]&m[1951]&~m[1952])|(m[815]&~m[1948]&m[1950]&m[1951]&~m[1952])|(~m[815]&m[1948]&~m[1950]&~m[1951]&m[1952])|(~m[815]&~m[1948]&m[1950]&~m[1951]&m[1952])|(m[815]&m[1948]&m[1950]&~m[1951]&m[1952])|(~m[815]&m[1948]&m[1950]&m[1951]&m[1952]))&UnbiasedRNG[700])|((m[815]&~m[1948]&~m[1950]&m[1951]&~m[1952])|(~m[815]&~m[1948]&~m[1950]&~m[1951]&m[1952])|(m[815]&~m[1948]&~m[1950]&~m[1951]&m[1952])|(m[815]&m[1948]&~m[1950]&~m[1951]&m[1952])|(m[815]&~m[1948]&m[1950]&~m[1951]&m[1952])|(~m[815]&~m[1948]&~m[1950]&m[1951]&m[1952])|(m[815]&~m[1948]&~m[1950]&m[1951]&m[1952])|(~m[815]&m[1948]&~m[1950]&m[1951]&m[1952])|(m[815]&m[1948]&~m[1950]&m[1951]&m[1952])|(~m[815]&~m[1948]&m[1950]&m[1951]&m[1952])|(m[815]&~m[1948]&m[1950]&m[1951]&m[1952])|(m[815]&m[1948]&m[1950]&m[1951]&m[1952]))):InitCond[1595];
    m[1954] = run?((((m[830]&~m[1953]&~m[1955]&~m[1956]&~m[1957])|(~m[830]&~m[1953]&~m[1955]&m[1956]&~m[1957])|(m[830]&m[1953]&~m[1955]&m[1956]&~m[1957])|(m[830]&~m[1953]&m[1955]&m[1956]&~m[1957])|(~m[830]&m[1953]&~m[1955]&~m[1956]&m[1957])|(~m[830]&~m[1953]&m[1955]&~m[1956]&m[1957])|(m[830]&m[1953]&m[1955]&~m[1956]&m[1957])|(~m[830]&m[1953]&m[1955]&m[1956]&m[1957]))&UnbiasedRNG[701])|((m[830]&~m[1953]&~m[1955]&m[1956]&~m[1957])|(~m[830]&~m[1953]&~m[1955]&~m[1956]&m[1957])|(m[830]&~m[1953]&~m[1955]&~m[1956]&m[1957])|(m[830]&m[1953]&~m[1955]&~m[1956]&m[1957])|(m[830]&~m[1953]&m[1955]&~m[1956]&m[1957])|(~m[830]&~m[1953]&~m[1955]&m[1956]&m[1957])|(m[830]&~m[1953]&~m[1955]&m[1956]&m[1957])|(~m[830]&m[1953]&~m[1955]&m[1956]&m[1957])|(m[830]&m[1953]&~m[1955]&m[1956]&m[1957])|(~m[830]&~m[1953]&m[1955]&m[1956]&m[1957])|(m[830]&~m[1953]&m[1955]&m[1956]&m[1957])|(m[830]&m[1953]&m[1955]&m[1956]&m[1957]))):InitCond[1596];
    m[1959] = run?((((m[845]&~m[1958]&~m[1960]&~m[1961]&~m[1962])|(~m[845]&~m[1958]&~m[1960]&m[1961]&~m[1962])|(m[845]&m[1958]&~m[1960]&m[1961]&~m[1962])|(m[845]&~m[1958]&m[1960]&m[1961]&~m[1962])|(~m[845]&m[1958]&~m[1960]&~m[1961]&m[1962])|(~m[845]&~m[1958]&m[1960]&~m[1961]&m[1962])|(m[845]&m[1958]&m[1960]&~m[1961]&m[1962])|(~m[845]&m[1958]&m[1960]&m[1961]&m[1962]))&UnbiasedRNG[702])|((m[845]&~m[1958]&~m[1960]&m[1961]&~m[1962])|(~m[845]&~m[1958]&~m[1960]&~m[1961]&m[1962])|(m[845]&~m[1958]&~m[1960]&~m[1961]&m[1962])|(m[845]&m[1958]&~m[1960]&~m[1961]&m[1962])|(m[845]&~m[1958]&m[1960]&~m[1961]&m[1962])|(~m[845]&~m[1958]&~m[1960]&m[1961]&m[1962])|(m[845]&~m[1958]&~m[1960]&m[1961]&m[1962])|(~m[845]&m[1958]&~m[1960]&m[1961]&m[1962])|(m[845]&m[1958]&~m[1960]&m[1961]&m[1962])|(~m[845]&~m[1958]&m[1960]&m[1961]&m[1962])|(m[845]&~m[1958]&m[1960]&m[1961]&m[1962])|(m[845]&m[1958]&m[1960]&m[1961]&m[1962]))):InitCond[1597];
    m[1964] = run?((((m[860]&~m[1963]&~m[1965]&~m[1966]&~m[1967])|(~m[860]&~m[1963]&~m[1965]&m[1966]&~m[1967])|(m[860]&m[1963]&~m[1965]&m[1966]&~m[1967])|(m[860]&~m[1963]&m[1965]&m[1966]&~m[1967])|(~m[860]&m[1963]&~m[1965]&~m[1966]&m[1967])|(~m[860]&~m[1963]&m[1965]&~m[1966]&m[1967])|(m[860]&m[1963]&m[1965]&~m[1966]&m[1967])|(~m[860]&m[1963]&m[1965]&m[1966]&m[1967]))&UnbiasedRNG[703])|((m[860]&~m[1963]&~m[1965]&m[1966]&~m[1967])|(~m[860]&~m[1963]&~m[1965]&~m[1966]&m[1967])|(m[860]&~m[1963]&~m[1965]&~m[1966]&m[1967])|(m[860]&m[1963]&~m[1965]&~m[1966]&m[1967])|(m[860]&~m[1963]&m[1965]&~m[1966]&m[1967])|(~m[860]&~m[1963]&~m[1965]&m[1966]&m[1967])|(m[860]&~m[1963]&~m[1965]&m[1966]&m[1967])|(~m[860]&m[1963]&~m[1965]&m[1966]&m[1967])|(m[860]&m[1963]&~m[1965]&m[1966]&m[1967])|(~m[860]&~m[1963]&m[1965]&m[1966]&m[1967])|(m[860]&~m[1963]&m[1965]&m[1966]&m[1967])|(m[860]&m[1963]&m[1965]&m[1966]&m[1967]))):InitCond[1598];
    m[1969] = run?((((m[875]&~m[1968]&~m[1970]&~m[1971]&~m[1972])|(~m[875]&~m[1968]&~m[1970]&m[1971]&~m[1972])|(m[875]&m[1968]&~m[1970]&m[1971]&~m[1972])|(m[875]&~m[1968]&m[1970]&m[1971]&~m[1972])|(~m[875]&m[1968]&~m[1970]&~m[1971]&m[1972])|(~m[875]&~m[1968]&m[1970]&~m[1971]&m[1972])|(m[875]&m[1968]&m[1970]&~m[1971]&m[1972])|(~m[875]&m[1968]&m[1970]&m[1971]&m[1972]))&UnbiasedRNG[704])|((m[875]&~m[1968]&~m[1970]&m[1971]&~m[1972])|(~m[875]&~m[1968]&~m[1970]&~m[1971]&m[1972])|(m[875]&~m[1968]&~m[1970]&~m[1971]&m[1972])|(m[875]&m[1968]&~m[1970]&~m[1971]&m[1972])|(m[875]&~m[1968]&m[1970]&~m[1971]&m[1972])|(~m[875]&~m[1968]&~m[1970]&m[1971]&m[1972])|(m[875]&~m[1968]&~m[1970]&m[1971]&m[1972])|(~m[875]&m[1968]&~m[1970]&m[1971]&m[1972])|(m[875]&m[1968]&~m[1970]&m[1971]&m[1972])|(~m[875]&~m[1968]&m[1970]&m[1971]&m[1972])|(m[875]&~m[1968]&m[1970]&m[1971]&m[1972])|(m[875]&m[1968]&m[1970]&m[1971]&m[1972]))):InitCond[1599];
    m[1974] = run?((((m[890]&~m[1973]&~m[1975]&~m[1976]&~m[1977])|(~m[890]&~m[1973]&~m[1975]&m[1976]&~m[1977])|(m[890]&m[1973]&~m[1975]&m[1976]&~m[1977])|(m[890]&~m[1973]&m[1975]&m[1976]&~m[1977])|(~m[890]&m[1973]&~m[1975]&~m[1976]&m[1977])|(~m[890]&~m[1973]&m[1975]&~m[1976]&m[1977])|(m[890]&m[1973]&m[1975]&~m[1976]&m[1977])|(~m[890]&m[1973]&m[1975]&m[1976]&m[1977]))&UnbiasedRNG[705])|((m[890]&~m[1973]&~m[1975]&m[1976]&~m[1977])|(~m[890]&~m[1973]&~m[1975]&~m[1976]&m[1977])|(m[890]&~m[1973]&~m[1975]&~m[1976]&m[1977])|(m[890]&m[1973]&~m[1975]&~m[1976]&m[1977])|(m[890]&~m[1973]&m[1975]&~m[1976]&m[1977])|(~m[890]&~m[1973]&~m[1975]&m[1976]&m[1977])|(m[890]&~m[1973]&~m[1975]&m[1976]&m[1977])|(~m[890]&m[1973]&~m[1975]&m[1976]&m[1977])|(m[890]&m[1973]&~m[1975]&m[1976]&m[1977])|(~m[890]&~m[1973]&m[1975]&m[1976]&m[1977])|(m[890]&~m[1973]&m[1975]&m[1976]&m[1977])|(m[890]&m[1973]&m[1975]&m[1976]&m[1977]))):InitCond[1600];
    m[1979] = run?((((m[905]&~m[1978]&~m[1980]&~m[1981]&~m[1982])|(~m[905]&~m[1978]&~m[1980]&m[1981]&~m[1982])|(m[905]&m[1978]&~m[1980]&m[1981]&~m[1982])|(m[905]&~m[1978]&m[1980]&m[1981]&~m[1982])|(~m[905]&m[1978]&~m[1980]&~m[1981]&m[1982])|(~m[905]&~m[1978]&m[1980]&~m[1981]&m[1982])|(m[905]&m[1978]&m[1980]&~m[1981]&m[1982])|(~m[905]&m[1978]&m[1980]&m[1981]&m[1982]))&UnbiasedRNG[706])|((m[905]&~m[1978]&~m[1980]&m[1981]&~m[1982])|(~m[905]&~m[1978]&~m[1980]&~m[1981]&m[1982])|(m[905]&~m[1978]&~m[1980]&~m[1981]&m[1982])|(m[905]&m[1978]&~m[1980]&~m[1981]&m[1982])|(m[905]&~m[1978]&m[1980]&~m[1981]&m[1982])|(~m[905]&~m[1978]&~m[1980]&m[1981]&m[1982])|(m[905]&~m[1978]&~m[1980]&m[1981]&m[1982])|(~m[905]&m[1978]&~m[1980]&m[1981]&m[1982])|(m[905]&m[1978]&~m[1980]&m[1981]&m[1982])|(~m[905]&~m[1978]&m[1980]&m[1981]&m[1982])|(m[905]&~m[1978]&m[1980]&m[1981]&m[1982])|(m[905]&m[1978]&m[1980]&m[1981]&m[1982]))):InitCond[1601];
    m[1984] = run?((((m[920]&~m[1983]&~m[1985]&~m[1986]&~m[1987])|(~m[920]&~m[1983]&~m[1985]&m[1986]&~m[1987])|(m[920]&m[1983]&~m[1985]&m[1986]&~m[1987])|(m[920]&~m[1983]&m[1985]&m[1986]&~m[1987])|(~m[920]&m[1983]&~m[1985]&~m[1986]&m[1987])|(~m[920]&~m[1983]&m[1985]&~m[1986]&m[1987])|(m[920]&m[1983]&m[1985]&~m[1986]&m[1987])|(~m[920]&m[1983]&m[1985]&m[1986]&m[1987]))&UnbiasedRNG[707])|((m[920]&~m[1983]&~m[1985]&m[1986]&~m[1987])|(~m[920]&~m[1983]&~m[1985]&~m[1986]&m[1987])|(m[920]&~m[1983]&~m[1985]&~m[1986]&m[1987])|(m[920]&m[1983]&~m[1985]&~m[1986]&m[1987])|(m[920]&~m[1983]&m[1985]&~m[1986]&m[1987])|(~m[920]&~m[1983]&~m[1985]&m[1986]&m[1987])|(m[920]&~m[1983]&~m[1985]&m[1986]&m[1987])|(~m[920]&m[1983]&~m[1985]&m[1986]&m[1987])|(m[920]&m[1983]&~m[1985]&m[1986]&m[1987])|(~m[920]&~m[1983]&m[1985]&m[1986]&m[1987])|(m[920]&~m[1983]&m[1985]&m[1986]&m[1987])|(m[920]&m[1983]&m[1985]&m[1986]&m[1987]))):InitCond[1602];
    m[1989] = run?((((m[831]&~m[1988]&~m[1990]&~m[1991]&~m[1992])|(~m[831]&~m[1988]&~m[1990]&m[1991]&~m[1992])|(m[831]&m[1988]&~m[1990]&m[1991]&~m[1992])|(m[831]&~m[1988]&m[1990]&m[1991]&~m[1992])|(~m[831]&m[1988]&~m[1990]&~m[1991]&m[1992])|(~m[831]&~m[1988]&m[1990]&~m[1991]&m[1992])|(m[831]&m[1988]&m[1990]&~m[1991]&m[1992])|(~m[831]&m[1988]&m[1990]&m[1991]&m[1992]))&UnbiasedRNG[708])|((m[831]&~m[1988]&~m[1990]&m[1991]&~m[1992])|(~m[831]&~m[1988]&~m[1990]&~m[1991]&m[1992])|(m[831]&~m[1988]&~m[1990]&~m[1991]&m[1992])|(m[831]&m[1988]&~m[1990]&~m[1991]&m[1992])|(m[831]&~m[1988]&m[1990]&~m[1991]&m[1992])|(~m[831]&~m[1988]&~m[1990]&m[1991]&m[1992])|(m[831]&~m[1988]&~m[1990]&m[1991]&m[1992])|(~m[831]&m[1988]&~m[1990]&m[1991]&m[1992])|(m[831]&m[1988]&~m[1990]&m[1991]&m[1992])|(~m[831]&~m[1988]&m[1990]&m[1991]&m[1992])|(m[831]&~m[1988]&m[1990]&m[1991]&m[1992])|(m[831]&m[1988]&m[1990]&m[1991]&m[1992]))):InitCond[1603];
    m[1994] = run?((((m[846]&~m[1993]&~m[1995]&~m[1996]&~m[1997])|(~m[846]&~m[1993]&~m[1995]&m[1996]&~m[1997])|(m[846]&m[1993]&~m[1995]&m[1996]&~m[1997])|(m[846]&~m[1993]&m[1995]&m[1996]&~m[1997])|(~m[846]&m[1993]&~m[1995]&~m[1996]&m[1997])|(~m[846]&~m[1993]&m[1995]&~m[1996]&m[1997])|(m[846]&m[1993]&m[1995]&~m[1996]&m[1997])|(~m[846]&m[1993]&m[1995]&m[1996]&m[1997]))&UnbiasedRNG[709])|((m[846]&~m[1993]&~m[1995]&m[1996]&~m[1997])|(~m[846]&~m[1993]&~m[1995]&~m[1996]&m[1997])|(m[846]&~m[1993]&~m[1995]&~m[1996]&m[1997])|(m[846]&m[1993]&~m[1995]&~m[1996]&m[1997])|(m[846]&~m[1993]&m[1995]&~m[1996]&m[1997])|(~m[846]&~m[1993]&~m[1995]&m[1996]&m[1997])|(m[846]&~m[1993]&~m[1995]&m[1996]&m[1997])|(~m[846]&m[1993]&~m[1995]&m[1996]&m[1997])|(m[846]&m[1993]&~m[1995]&m[1996]&m[1997])|(~m[846]&~m[1993]&m[1995]&m[1996]&m[1997])|(m[846]&~m[1993]&m[1995]&m[1996]&m[1997])|(m[846]&m[1993]&m[1995]&m[1996]&m[1997]))):InitCond[1604];
    m[1999] = run?((((m[861]&~m[1998]&~m[2000]&~m[2001]&~m[2002])|(~m[861]&~m[1998]&~m[2000]&m[2001]&~m[2002])|(m[861]&m[1998]&~m[2000]&m[2001]&~m[2002])|(m[861]&~m[1998]&m[2000]&m[2001]&~m[2002])|(~m[861]&m[1998]&~m[2000]&~m[2001]&m[2002])|(~m[861]&~m[1998]&m[2000]&~m[2001]&m[2002])|(m[861]&m[1998]&m[2000]&~m[2001]&m[2002])|(~m[861]&m[1998]&m[2000]&m[2001]&m[2002]))&UnbiasedRNG[710])|((m[861]&~m[1998]&~m[2000]&m[2001]&~m[2002])|(~m[861]&~m[1998]&~m[2000]&~m[2001]&m[2002])|(m[861]&~m[1998]&~m[2000]&~m[2001]&m[2002])|(m[861]&m[1998]&~m[2000]&~m[2001]&m[2002])|(m[861]&~m[1998]&m[2000]&~m[2001]&m[2002])|(~m[861]&~m[1998]&~m[2000]&m[2001]&m[2002])|(m[861]&~m[1998]&~m[2000]&m[2001]&m[2002])|(~m[861]&m[1998]&~m[2000]&m[2001]&m[2002])|(m[861]&m[1998]&~m[2000]&m[2001]&m[2002])|(~m[861]&~m[1998]&m[2000]&m[2001]&m[2002])|(m[861]&~m[1998]&m[2000]&m[2001]&m[2002])|(m[861]&m[1998]&m[2000]&m[2001]&m[2002]))):InitCond[1605];
    m[2004] = run?((((m[876]&~m[2003]&~m[2005]&~m[2006]&~m[2007])|(~m[876]&~m[2003]&~m[2005]&m[2006]&~m[2007])|(m[876]&m[2003]&~m[2005]&m[2006]&~m[2007])|(m[876]&~m[2003]&m[2005]&m[2006]&~m[2007])|(~m[876]&m[2003]&~m[2005]&~m[2006]&m[2007])|(~m[876]&~m[2003]&m[2005]&~m[2006]&m[2007])|(m[876]&m[2003]&m[2005]&~m[2006]&m[2007])|(~m[876]&m[2003]&m[2005]&m[2006]&m[2007]))&UnbiasedRNG[711])|((m[876]&~m[2003]&~m[2005]&m[2006]&~m[2007])|(~m[876]&~m[2003]&~m[2005]&~m[2006]&m[2007])|(m[876]&~m[2003]&~m[2005]&~m[2006]&m[2007])|(m[876]&m[2003]&~m[2005]&~m[2006]&m[2007])|(m[876]&~m[2003]&m[2005]&~m[2006]&m[2007])|(~m[876]&~m[2003]&~m[2005]&m[2006]&m[2007])|(m[876]&~m[2003]&~m[2005]&m[2006]&m[2007])|(~m[876]&m[2003]&~m[2005]&m[2006]&m[2007])|(m[876]&m[2003]&~m[2005]&m[2006]&m[2007])|(~m[876]&~m[2003]&m[2005]&m[2006]&m[2007])|(m[876]&~m[2003]&m[2005]&m[2006]&m[2007])|(m[876]&m[2003]&m[2005]&m[2006]&m[2007]))):InitCond[1606];
    m[2009] = run?((((m[891]&~m[2008]&~m[2010]&~m[2011]&~m[2012])|(~m[891]&~m[2008]&~m[2010]&m[2011]&~m[2012])|(m[891]&m[2008]&~m[2010]&m[2011]&~m[2012])|(m[891]&~m[2008]&m[2010]&m[2011]&~m[2012])|(~m[891]&m[2008]&~m[2010]&~m[2011]&m[2012])|(~m[891]&~m[2008]&m[2010]&~m[2011]&m[2012])|(m[891]&m[2008]&m[2010]&~m[2011]&m[2012])|(~m[891]&m[2008]&m[2010]&m[2011]&m[2012]))&UnbiasedRNG[712])|((m[891]&~m[2008]&~m[2010]&m[2011]&~m[2012])|(~m[891]&~m[2008]&~m[2010]&~m[2011]&m[2012])|(m[891]&~m[2008]&~m[2010]&~m[2011]&m[2012])|(m[891]&m[2008]&~m[2010]&~m[2011]&m[2012])|(m[891]&~m[2008]&m[2010]&~m[2011]&m[2012])|(~m[891]&~m[2008]&~m[2010]&m[2011]&m[2012])|(m[891]&~m[2008]&~m[2010]&m[2011]&m[2012])|(~m[891]&m[2008]&~m[2010]&m[2011]&m[2012])|(m[891]&m[2008]&~m[2010]&m[2011]&m[2012])|(~m[891]&~m[2008]&m[2010]&m[2011]&m[2012])|(m[891]&~m[2008]&m[2010]&m[2011]&m[2012])|(m[891]&m[2008]&m[2010]&m[2011]&m[2012]))):InitCond[1607];
    m[2014] = run?((((m[906]&~m[2013]&~m[2015]&~m[2016]&~m[2017])|(~m[906]&~m[2013]&~m[2015]&m[2016]&~m[2017])|(m[906]&m[2013]&~m[2015]&m[2016]&~m[2017])|(m[906]&~m[2013]&m[2015]&m[2016]&~m[2017])|(~m[906]&m[2013]&~m[2015]&~m[2016]&m[2017])|(~m[906]&~m[2013]&m[2015]&~m[2016]&m[2017])|(m[906]&m[2013]&m[2015]&~m[2016]&m[2017])|(~m[906]&m[2013]&m[2015]&m[2016]&m[2017]))&UnbiasedRNG[713])|((m[906]&~m[2013]&~m[2015]&m[2016]&~m[2017])|(~m[906]&~m[2013]&~m[2015]&~m[2016]&m[2017])|(m[906]&~m[2013]&~m[2015]&~m[2016]&m[2017])|(m[906]&m[2013]&~m[2015]&~m[2016]&m[2017])|(m[906]&~m[2013]&m[2015]&~m[2016]&m[2017])|(~m[906]&~m[2013]&~m[2015]&m[2016]&m[2017])|(m[906]&~m[2013]&~m[2015]&m[2016]&m[2017])|(~m[906]&m[2013]&~m[2015]&m[2016]&m[2017])|(m[906]&m[2013]&~m[2015]&m[2016]&m[2017])|(~m[906]&~m[2013]&m[2015]&m[2016]&m[2017])|(m[906]&~m[2013]&m[2015]&m[2016]&m[2017])|(m[906]&m[2013]&m[2015]&m[2016]&m[2017]))):InitCond[1608];
    m[2019] = run?((((m[921]&~m[2018]&~m[2020]&~m[2021]&~m[2022])|(~m[921]&~m[2018]&~m[2020]&m[2021]&~m[2022])|(m[921]&m[2018]&~m[2020]&m[2021]&~m[2022])|(m[921]&~m[2018]&m[2020]&m[2021]&~m[2022])|(~m[921]&m[2018]&~m[2020]&~m[2021]&m[2022])|(~m[921]&~m[2018]&m[2020]&~m[2021]&m[2022])|(m[921]&m[2018]&m[2020]&~m[2021]&m[2022])|(~m[921]&m[2018]&m[2020]&m[2021]&m[2022]))&UnbiasedRNG[714])|((m[921]&~m[2018]&~m[2020]&m[2021]&~m[2022])|(~m[921]&~m[2018]&~m[2020]&~m[2021]&m[2022])|(m[921]&~m[2018]&~m[2020]&~m[2021]&m[2022])|(m[921]&m[2018]&~m[2020]&~m[2021]&m[2022])|(m[921]&~m[2018]&m[2020]&~m[2021]&m[2022])|(~m[921]&~m[2018]&~m[2020]&m[2021]&m[2022])|(m[921]&~m[2018]&~m[2020]&m[2021]&m[2022])|(~m[921]&m[2018]&~m[2020]&m[2021]&m[2022])|(m[921]&m[2018]&~m[2020]&m[2021]&m[2022])|(~m[921]&~m[2018]&m[2020]&m[2021]&m[2022])|(m[921]&~m[2018]&m[2020]&m[2021]&m[2022])|(m[921]&m[2018]&m[2020]&m[2021]&m[2022]))):InitCond[1609];
    m[2024] = run?((((m[847]&~m[2023]&~m[2025]&~m[2026]&~m[2027])|(~m[847]&~m[2023]&~m[2025]&m[2026]&~m[2027])|(m[847]&m[2023]&~m[2025]&m[2026]&~m[2027])|(m[847]&~m[2023]&m[2025]&m[2026]&~m[2027])|(~m[847]&m[2023]&~m[2025]&~m[2026]&m[2027])|(~m[847]&~m[2023]&m[2025]&~m[2026]&m[2027])|(m[847]&m[2023]&m[2025]&~m[2026]&m[2027])|(~m[847]&m[2023]&m[2025]&m[2026]&m[2027]))&UnbiasedRNG[715])|((m[847]&~m[2023]&~m[2025]&m[2026]&~m[2027])|(~m[847]&~m[2023]&~m[2025]&~m[2026]&m[2027])|(m[847]&~m[2023]&~m[2025]&~m[2026]&m[2027])|(m[847]&m[2023]&~m[2025]&~m[2026]&m[2027])|(m[847]&~m[2023]&m[2025]&~m[2026]&m[2027])|(~m[847]&~m[2023]&~m[2025]&m[2026]&m[2027])|(m[847]&~m[2023]&~m[2025]&m[2026]&m[2027])|(~m[847]&m[2023]&~m[2025]&m[2026]&m[2027])|(m[847]&m[2023]&~m[2025]&m[2026]&m[2027])|(~m[847]&~m[2023]&m[2025]&m[2026]&m[2027])|(m[847]&~m[2023]&m[2025]&m[2026]&m[2027])|(m[847]&m[2023]&m[2025]&m[2026]&m[2027]))):InitCond[1610];
    m[2029] = run?((((m[862]&~m[2028]&~m[2030]&~m[2031]&~m[2032])|(~m[862]&~m[2028]&~m[2030]&m[2031]&~m[2032])|(m[862]&m[2028]&~m[2030]&m[2031]&~m[2032])|(m[862]&~m[2028]&m[2030]&m[2031]&~m[2032])|(~m[862]&m[2028]&~m[2030]&~m[2031]&m[2032])|(~m[862]&~m[2028]&m[2030]&~m[2031]&m[2032])|(m[862]&m[2028]&m[2030]&~m[2031]&m[2032])|(~m[862]&m[2028]&m[2030]&m[2031]&m[2032]))&UnbiasedRNG[716])|((m[862]&~m[2028]&~m[2030]&m[2031]&~m[2032])|(~m[862]&~m[2028]&~m[2030]&~m[2031]&m[2032])|(m[862]&~m[2028]&~m[2030]&~m[2031]&m[2032])|(m[862]&m[2028]&~m[2030]&~m[2031]&m[2032])|(m[862]&~m[2028]&m[2030]&~m[2031]&m[2032])|(~m[862]&~m[2028]&~m[2030]&m[2031]&m[2032])|(m[862]&~m[2028]&~m[2030]&m[2031]&m[2032])|(~m[862]&m[2028]&~m[2030]&m[2031]&m[2032])|(m[862]&m[2028]&~m[2030]&m[2031]&m[2032])|(~m[862]&~m[2028]&m[2030]&m[2031]&m[2032])|(m[862]&~m[2028]&m[2030]&m[2031]&m[2032])|(m[862]&m[2028]&m[2030]&m[2031]&m[2032]))):InitCond[1611];
    m[2034] = run?((((m[877]&~m[2033]&~m[2035]&~m[2036]&~m[2037])|(~m[877]&~m[2033]&~m[2035]&m[2036]&~m[2037])|(m[877]&m[2033]&~m[2035]&m[2036]&~m[2037])|(m[877]&~m[2033]&m[2035]&m[2036]&~m[2037])|(~m[877]&m[2033]&~m[2035]&~m[2036]&m[2037])|(~m[877]&~m[2033]&m[2035]&~m[2036]&m[2037])|(m[877]&m[2033]&m[2035]&~m[2036]&m[2037])|(~m[877]&m[2033]&m[2035]&m[2036]&m[2037]))&UnbiasedRNG[717])|((m[877]&~m[2033]&~m[2035]&m[2036]&~m[2037])|(~m[877]&~m[2033]&~m[2035]&~m[2036]&m[2037])|(m[877]&~m[2033]&~m[2035]&~m[2036]&m[2037])|(m[877]&m[2033]&~m[2035]&~m[2036]&m[2037])|(m[877]&~m[2033]&m[2035]&~m[2036]&m[2037])|(~m[877]&~m[2033]&~m[2035]&m[2036]&m[2037])|(m[877]&~m[2033]&~m[2035]&m[2036]&m[2037])|(~m[877]&m[2033]&~m[2035]&m[2036]&m[2037])|(m[877]&m[2033]&~m[2035]&m[2036]&m[2037])|(~m[877]&~m[2033]&m[2035]&m[2036]&m[2037])|(m[877]&~m[2033]&m[2035]&m[2036]&m[2037])|(m[877]&m[2033]&m[2035]&m[2036]&m[2037]))):InitCond[1612];
    m[2039] = run?((((m[892]&~m[2038]&~m[2040]&~m[2041]&~m[2042])|(~m[892]&~m[2038]&~m[2040]&m[2041]&~m[2042])|(m[892]&m[2038]&~m[2040]&m[2041]&~m[2042])|(m[892]&~m[2038]&m[2040]&m[2041]&~m[2042])|(~m[892]&m[2038]&~m[2040]&~m[2041]&m[2042])|(~m[892]&~m[2038]&m[2040]&~m[2041]&m[2042])|(m[892]&m[2038]&m[2040]&~m[2041]&m[2042])|(~m[892]&m[2038]&m[2040]&m[2041]&m[2042]))&UnbiasedRNG[718])|((m[892]&~m[2038]&~m[2040]&m[2041]&~m[2042])|(~m[892]&~m[2038]&~m[2040]&~m[2041]&m[2042])|(m[892]&~m[2038]&~m[2040]&~m[2041]&m[2042])|(m[892]&m[2038]&~m[2040]&~m[2041]&m[2042])|(m[892]&~m[2038]&m[2040]&~m[2041]&m[2042])|(~m[892]&~m[2038]&~m[2040]&m[2041]&m[2042])|(m[892]&~m[2038]&~m[2040]&m[2041]&m[2042])|(~m[892]&m[2038]&~m[2040]&m[2041]&m[2042])|(m[892]&m[2038]&~m[2040]&m[2041]&m[2042])|(~m[892]&~m[2038]&m[2040]&m[2041]&m[2042])|(m[892]&~m[2038]&m[2040]&m[2041]&m[2042])|(m[892]&m[2038]&m[2040]&m[2041]&m[2042]))):InitCond[1613];
    m[2044] = run?((((m[907]&~m[2043]&~m[2045]&~m[2046]&~m[2047])|(~m[907]&~m[2043]&~m[2045]&m[2046]&~m[2047])|(m[907]&m[2043]&~m[2045]&m[2046]&~m[2047])|(m[907]&~m[2043]&m[2045]&m[2046]&~m[2047])|(~m[907]&m[2043]&~m[2045]&~m[2046]&m[2047])|(~m[907]&~m[2043]&m[2045]&~m[2046]&m[2047])|(m[907]&m[2043]&m[2045]&~m[2046]&m[2047])|(~m[907]&m[2043]&m[2045]&m[2046]&m[2047]))&UnbiasedRNG[719])|((m[907]&~m[2043]&~m[2045]&m[2046]&~m[2047])|(~m[907]&~m[2043]&~m[2045]&~m[2046]&m[2047])|(m[907]&~m[2043]&~m[2045]&~m[2046]&m[2047])|(m[907]&m[2043]&~m[2045]&~m[2046]&m[2047])|(m[907]&~m[2043]&m[2045]&~m[2046]&m[2047])|(~m[907]&~m[2043]&~m[2045]&m[2046]&m[2047])|(m[907]&~m[2043]&~m[2045]&m[2046]&m[2047])|(~m[907]&m[2043]&~m[2045]&m[2046]&m[2047])|(m[907]&m[2043]&~m[2045]&m[2046]&m[2047])|(~m[907]&~m[2043]&m[2045]&m[2046]&m[2047])|(m[907]&~m[2043]&m[2045]&m[2046]&m[2047])|(m[907]&m[2043]&m[2045]&m[2046]&m[2047]))):InitCond[1614];
    m[2049] = run?((((m[922]&~m[2048]&~m[2050]&~m[2051]&~m[2052])|(~m[922]&~m[2048]&~m[2050]&m[2051]&~m[2052])|(m[922]&m[2048]&~m[2050]&m[2051]&~m[2052])|(m[922]&~m[2048]&m[2050]&m[2051]&~m[2052])|(~m[922]&m[2048]&~m[2050]&~m[2051]&m[2052])|(~m[922]&~m[2048]&m[2050]&~m[2051]&m[2052])|(m[922]&m[2048]&m[2050]&~m[2051]&m[2052])|(~m[922]&m[2048]&m[2050]&m[2051]&m[2052]))&UnbiasedRNG[720])|((m[922]&~m[2048]&~m[2050]&m[2051]&~m[2052])|(~m[922]&~m[2048]&~m[2050]&~m[2051]&m[2052])|(m[922]&~m[2048]&~m[2050]&~m[2051]&m[2052])|(m[922]&m[2048]&~m[2050]&~m[2051]&m[2052])|(m[922]&~m[2048]&m[2050]&~m[2051]&m[2052])|(~m[922]&~m[2048]&~m[2050]&m[2051]&m[2052])|(m[922]&~m[2048]&~m[2050]&m[2051]&m[2052])|(~m[922]&m[2048]&~m[2050]&m[2051]&m[2052])|(m[922]&m[2048]&~m[2050]&m[2051]&m[2052])|(~m[922]&~m[2048]&m[2050]&m[2051]&m[2052])|(m[922]&~m[2048]&m[2050]&m[2051]&m[2052])|(m[922]&m[2048]&m[2050]&m[2051]&m[2052]))):InitCond[1615];
    m[2054] = run?((((m[863]&~m[2053]&~m[2055]&~m[2056]&~m[2057])|(~m[863]&~m[2053]&~m[2055]&m[2056]&~m[2057])|(m[863]&m[2053]&~m[2055]&m[2056]&~m[2057])|(m[863]&~m[2053]&m[2055]&m[2056]&~m[2057])|(~m[863]&m[2053]&~m[2055]&~m[2056]&m[2057])|(~m[863]&~m[2053]&m[2055]&~m[2056]&m[2057])|(m[863]&m[2053]&m[2055]&~m[2056]&m[2057])|(~m[863]&m[2053]&m[2055]&m[2056]&m[2057]))&UnbiasedRNG[721])|((m[863]&~m[2053]&~m[2055]&m[2056]&~m[2057])|(~m[863]&~m[2053]&~m[2055]&~m[2056]&m[2057])|(m[863]&~m[2053]&~m[2055]&~m[2056]&m[2057])|(m[863]&m[2053]&~m[2055]&~m[2056]&m[2057])|(m[863]&~m[2053]&m[2055]&~m[2056]&m[2057])|(~m[863]&~m[2053]&~m[2055]&m[2056]&m[2057])|(m[863]&~m[2053]&~m[2055]&m[2056]&m[2057])|(~m[863]&m[2053]&~m[2055]&m[2056]&m[2057])|(m[863]&m[2053]&~m[2055]&m[2056]&m[2057])|(~m[863]&~m[2053]&m[2055]&m[2056]&m[2057])|(m[863]&~m[2053]&m[2055]&m[2056]&m[2057])|(m[863]&m[2053]&m[2055]&m[2056]&m[2057]))):InitCond[1616];
    m[2059] = run?((((m[878]&~m[2058]&~m[2060]&~m[2061]&~m[2062])|(~m[878]&~m[2058]&~m[2060]&m[2061]&~m[2062])|(m[878]&m[2058]&~m[2060]&m[2061]&~m[2062])|(m[878]&~m[2058]&m[2060]&m[2061]&~m[2062])|(~m[878]&m[2058]&~m[2060]&~m[2061]&m[2062])|(~m[878]&~m[2058]&m[2060]&~m[2061]&m[2062])|(m[878]&m[2058]&m[2060]&~m[2061]&m[2062])|(~m[878]&m[2058]&m[2060]&m[2061]&m[2062]))&UnbiasedRNG[722])|((m[878]&~m[2058]&~m[2060]&m[2061]&~m[2062])|(~m[878]&~m[2058]&~m[2060]&~m[2061]&m[2062])|(m[878]&~m[2058]&~m[2060]&~m[2061]&m[2062])|(m[878]&m[2058]&~m[2060]&~m[2061]&m[2062])|(m[878]&~m[2058]&m[2060]&~m[2061]&m[2062])|(~m[878]&~m[2058]&~m[2060]&m[2061]&m[2062])|(m[878]&~m[2058]&~m[2060]&m[2061]&m[2062])|(~m[878]&m[2058]&~m[2060]&m[2061]&m[2062])|(m[878]&m[2058]&~m[2060]&m[2061]&m[2062])|(~m[878]&~m[2058]&m[2060]&m[2061]&m[2062])|(m[878]&~m[2058]&m[2060]&m[2061]&m[2062])|(m[878]&m[2058]&m[2060]&m[2061]&m[2062]))):InitCond[1617];
    m[2064] = run?((((m[893]&~m[2063]&~m[2065]&~m[2066]&~m[2067])|(~m[893]&~m[2063]&~m[2065]&m[2066]&~m[2067])|(m[893]&m[2063]&~m[2065]&m[2066]&~m[2067])|(m[893]&~m[2063]&m[2065]&m[2066]&~m[2067])|(~m[893]&m[2063]&~m[2065]&~m[2066]&m[2067])|(~m[893]&~m[2063]&m[2065]&~m[2066]&m[2067])|(m[893]&m[2063]&m[2065]&~m[2066]&m[2067])|(~m[893]&m[2063]&m[2065]&m[2066]&m[2067]))&UnbiasedRNG[723])|((m[893]&~m[2063]&~m[2065]&m[2066]&~m[2067])|(~m[893]&~m[2063]&~m[2065]&~m[2066]&m[2067])|(m[893]&~m[2063]&~m[2065]&~m[2066]&m[2067])|(m[893]&m[2063]&~m[2065]&~m[2066]&m[2067])|(m[893]&~m[2063]&m[2065]&~m[2066]&m[2067])|(~m[893]&~m[2063]&~m[2065]&m[2066]&m[2067])|(m[893]&~m[2063]&~m[2065]&m[2066]&m[2067])|(~m[893]&m[2063]&~m[2065]&m[2066]&m[2067])|(m[893]&m[2063]&~m[2065]&m[2066]&m[2067])|(~m[893]&~m[2063]&m[2065]&m[2066]&m[2067])|(m[893]&~m[2063]&m[2065]&m[2066]&m[2067])|(m[893]&m[2063]&m[2065]&m[2066]&m[2067]))):InitCond[1618];
    m[2069] = run?((((m[908]&~m[2068]&~m[2070]&~m[2071]&~m[2072])|(~m[908]&~m[2068]&~m[2070]&m[2071]&~m[2072])|(m[908]&m[2068]&~m[2070]&m[2071]&~m[2072])|(m[908]&~m[2068]&m[2070]&m[2071]&~m[2072])|(~m[908]&m[2068]&~m[2070]&~m[2071]&m[2072])|(~m[908]&~m[2068]&m[2070]&~m[2071]&m[2072])|(m[908]&m[2068]&m[2070]&~m[2071]&m[2072])|(~m[908]&m[2068]&m[2070]&m[2071]&m[2072]))&UnbiasedRNG[724])|((m[908]&~m[2068]&~m[2070]&m[2071]&~m[2072])|(~m[908]&~m[2068]&~m[2070]&~m[2071]&m[2072])|(m[908]&~m[2068]&~m[2070]&~m[2071]&m[2072])|(m[908]&m[2068]&~m[2070]&~m[2071]&m[2072])|(m[908]&~m[2068]&m[2070]&~m[2071]&m[2072])|(~m[908]&~m[2068]&~m[2070]&m[2071]&m[2072])|(m[908]&~m[2068]&~m[2070]&m[2071]&m[2072])|(~m[908]&m[2068]&~m[2070]&m[2071]&m[2072])|(m[908]&m[2068]&~m[2070]&m[2071]&m[2072])|(~m[908]&~m[2068]&m[2070]&m[2071]&m[2072])|(m[908]&~m[2068]&m[2070]&m[2071]&m[2072])|(m[908]&m[2068]&m[2070]&m[2071]&m[2072]))):InitCond[1619];
    m[2074] = run?((((m[923]&~m[2073]&~m[2075]&~m[2076]&~m[2077])|(~m[923]&~m[2073]&~m[2075]&m[2076]&~m[2077])|(m[923]&m[2073]&~m[2075]&m[2076]&~m[2077])|(m[923]&~m[2073]&m[2075]&m[2076]&~m[2077])|(~m[923]&m[2073]&~m[2075]&~m[2076]&m[2077])|(~m[923]&~m[2073]&m[2075]&~m[2076]&m[2077])|(m[923]&m[2073]&m[2075]&~m[2076]&m[2077])|(~m[923]&m[2073]&m[2075]&m[2076]&m[2077]))&UnbiasedRNG[725])|((m[923]&~m[2073]&~m[2075]&m[2076]&~m[2077])|(~m[923]&~m[2073]&~m[2075]&~m[2076]&m[2077])|(m[923]&~m[2073]&~m[2075]&~m[2076]&m[2077])|(m[923]&m[2073]&~m[2075]&~m[2076]&m[2077])|(m[923]&~m[2073]&m[2075]&~m[2076]&m[2077])|(~m[923]&~m[2073]&~m[2075]&m[2076]&m[2077])|(m[923]&~m[2073]&~m[2075]&m[2076]&m[2077])|(~m[923]&m[2073]&~m[2075]&m[2076]&m[2077])|(m[923]&m[2073]&~m[2075]&m[2076]&m[2077])|(~m[923]&~m[2073]&m[2075]&m[2076]&m[2077])|(m[923]&~m[2073]&m[2075]&m[2076]&m[2077])|(m[923]&m[2073]&m[2075]&m[2076]&m[2077]))):InitCond[1620];
    m[2079] = run?((((m[879]&~m[2078]&~m[2080]&~m[2081]&~m[2082])|(~m[879]&~m[2078]&~m[2080]&m[2081]&~m[2082])|(m[879]&m[2078]&~m[2080]&m[2081]&~m[2082])|(m[879]&~m[2078]&m[2080]&m[2081]&~m[2082])|(~m[879]&m[2078]&~m[2080]&~m[2081]&m[2082])|(~m[879]&~m[2078]&m[2080]&~m[2081]&m[2082])|(m[879]&m[2078]&m[2080]&~m[2081]&m[2082])|(~m[879]&m[2078]&m[2080]&m[2081]&m[2082]))&UnbiasedRNG[726])|((m[879]&~m[2078]&~m[2080]&m[2081]&~m[2082])|(~m[879]&~m[2078]&~m[2080]&~m[2081]&m[2082])|(m[879]&~m[2078]&~m[2080]&~m[2081]&m[2082])|(m[879]&m[2078]&~m[2080]&~m[2081]&m[2082])|(m[879]&~m[2078]&m[2080]&~m[2081]&m[2082])|(~m[879]&~m[2078]&~m[2080]&m[2081]&m[2082])|(m[879]&~m[2078]&~m[2080]&m[2081]&m[2082])|(~m[879]&m[2078]&~m[2080]&m[2081]&m[2082])|(m[879]&m[2078]&~m[2080]&m[2081]&m[2082])|(~m[879]&~m[2078]&m[2080]&m[2081]&m[2082])|(m[879]&~m[2078]&m[2080]&m[2081]&m[2082])|(m[879]&m[2078]&m[2080]&m[2081]&m[2082]))):InitCond[1621];
    m[2084] = run?((((m[894]&~m[2083]&~m[2085]&~m[2086]&~m[2087])|(~m[894]&~m[2083]&~m[2085]&m[2086]&~m[2087])|(m[894]&m[2083]&~m[2085]&m[2086]&~m[2087])|(m[894]&~m[2083]&m[2085]&m[2086]&~m[2087])|(~m[894]&m[2083]&~m[2085]&~m[2086]&m[2087])|(~m[894]&~m[2083]&m[2085]&~m[2086]&m[2087])|(m[894]&m[2083]&m[2085]&~m[2086]&m[2087])|(~m[894]&m[2083]&m[2085]&m[2086]&m[2087]))&UnbiasedRNG[727])|((m[894]&~m[2083]&~m[2085]&m[2086]&~m[2087])|(~m[894]&~m[2083]&~m[2085]&~m[2086]&m[2087])|(m[894]&~m[2083]&~m[2085]&~m[2086]&m[2087])|(m[894]&m[2083]&~m[2085]&~m[2086]&m[2087])|(m[894]&~m[2083]&m[2085]&~m[2086]&m[2087])|(~m[894]&~m[2083]&~m[2085]&m[2086]&m[2087])|(m[894]&~m[2083]&~m[2085]&m[2086]&m[2087])|(~m[894]&m[2083]&~m[2085]&m[2086]&m[2087])|(m[894]&m[2083]&~m[2085]&m[2086]&m[2087])|(~m[894]&~m[2083]&m[2085]&m[2086]&m[2087])|(m[894]&~m[2083]&m[2085]&m[2086]&m[2087])|(m[894]&m[2083]&m[2085]&m[2086]&m[2087]))):InitCond[1622];
    m[2089] = run?((((m[909]&~m[2088]&~m[2090]&~m[2091]&~m[2092])|(~m[909]&~m[2088]&~m[2090]&m[2091]&~m[2092])|(m[909]&m[2088]&~m[2090]&m[2091]&~m[2092])|(m[909]&~m[2088]&m[2090]&m[2091]&~m[2092])|(~m[909]&m[2088]&~m[2090]&~m[2091]&m[2092])|(~m[909]&~m[2088]&m[2090]&~m[2091]&m[2092])|(m[909]&m[2088]&m[2090]&~m[2091]&m[2092])|(~m[909]&m[2088]&m[2090]&m[2091]&m[2092]))&UnbiasedRNG[728])|((m[909]&~m[2088]&~m[2090]&m[2091]&~m[2092])|(~m[909]&~m[2088]&~m[2090]&~m[2091]&m[2092])|(m[909]&~m[2088]&~m[2090]&~m[2091]&m[2092])|(m[909]&m[2088]&~m[2090]&~m[2091]&m[2092])|(m[909]&~m[2088]&m[2090]&~m[2091]&m[2092])|(~m[909]&~m[2088]&~m[2090]&m[2091]&m[2092])|(m[909]&~m[2088]&~m[2090]&m[2091]&m[2092])|(~m[909]&m[2088]&~m[2090]&m[2091]&m[2092])|(m[909]&m[2088]&~m[2090]&m[2091]&m[2092])|(~m[909]&~m[2088]&m[2090]&m[2091]&m[2092])|(m[909]&~m[2088]&m[2090]&m[2091]&m[2092])|(m[909]&m[2088]&m[2090]&m[2091]&m[2092]))):InitCond[1623];
    m[2094] = run?((((m[924]&~m[2093]&~m[2095]&~m[2096]&~m[2097])|(~m[924]&~m[2093]&~m[2095]&m[2096]&~m[2097])|(m[924]&m[2093]&~m[2095]&m[2096]&~m[2097])|(m[924]&~m[2093]&m[2095]&m[2096]&~m[2097])|(~m[924]&m[2093]&~m[2095]&~m[2096]&m[2097])|(~m[924]&~m[2093]&m[2095]&~m[2096]&m[2097])|(m[924]&m[2093]&m[2095]&~m[2096]&m[2097])|(~m[924]&m[2093]&m[2095]&m[2096]&m[2097]))&UnbiasedRNG[729])|((m[924]&~m[2093]&~m[2095]&m[2096]&~m[2097])|(~m[924]&~m[2093]&~m[2095]&~m[2096]&m[2097])|(m[924]&~m[2093]&~m[2095]&~m[2096]&m[2097])|(m[924]&m[2093]&~m[2095]&~m[2096]&m[2097])|(m[924]&~m[2093]&m[2095]&~m[2096]&m[2097])|(~m[924]&~m[2093]&~m[2095]&m[2096]&m[2097])|(m[924]&~m[2093]&~m[2095]&m[2096]&m[2097])|(~m[924]&m[2093]&~m[2095]&m[2096]&m[2097])|(m[924]&m[2093]&~m[2095]&m[2096]&m[2097])|(~m[924]&~m[2093]&m[2095]&m[2096]&m[2097])|(m[924]&~m[2093]&m[2095]&m[2096]&m[2097])|(m[924]&m[2093]&m[2095]&m[2096]&m[2097]))):InitCond[1624];
    m[2099] = run?((((m[895]&~m[2098]&~m[2100]&~m[2101]&~m[2102])|(~m[895]&~m[2098]&~m[2100]&m[2101]&~m[2102])|(m[895]&m[2098]&~m[2100]&m[2101]&~m[2102])|(m[895]&~m[2098]&m[2100]&m[2101]&~m[2102])|(~m[895]&m[2098]&~m[2100]&~m[2101]&m[2102])|(~m[895]&~m[2098]&m[2100]&~m[2101]&m[2102])|(m[895]&m[2098]&m[2100]&~m[2101]&m[2102])|(~m[895]&m[2098]&m[2100]&m[2101]&m[2102]))&UnbiasedRNG[730])|((m[895]&~m[2098]&~m[2100]&m[2101]&~m[2102])|(~m[895]&~m[2098]&~m[2100]&~m[2101]&m[2102])|(m[895]&~m[2098]&~m[2100]&~m[2101]&m[2102])|(m[895]&m[2098]&~m[2100]&~m[2101]&m[2102])|(m[895]&~m[2098]&m[2100]&~m[2101]&m[2102])|(~m[895]&~m[2098]&~m[2100]&m[2101]&m[2102])|(m[895]&~m[2098]&~m[2100]&m[2101]&m[2102])|(~m[895]&m[2098]&~m[2100]&m[2101]&m[2102])|(m[895]&m[2098]&~m[2100]&m[2101]&m[2102])|(~m[895]&~m[2098]&m[2100]&m[2101]&m[2102])|(m[895]&~m[2098]&m[2100]&m[2101]&m[2102])|(m[895]&m[2098]&m[2100]&m[2101]&m[2102]))):InitCond[1625];
    m[2104] = run?((((m[910]&~m[2103]&~m[2105]&~m[2106]&~m[2107])|(~m[910]&~m[2103]&~m[2105]&m[2106]&~m[2107])|(m[910]&m[2103]&~m[2105]&m[2106]&~m[2107])|(m[910]&~m[2103]&m[2105]&m[2106]&~m[2107])|(~m[910]&m[2103]&~m[2105]&~m[2106]&m[2107])|(~m[910]&~m[2103]&m[2105]&~m[2106]&m[2107])|(m[910]&m[2103]&m[2105]&~m[2106]&m[2107])|(~m[910]&m[2103]&m[2105]&m[2106]&m[2107]))&UnbiasedRNG[731])|((m[910]&~m[2103]&~m[2105]&m[2106]&~m[2107])|(~m[910]&~m[2103]&~m[2105]&~m[2106]&m[2107])|(m[910]&~m[2103]&~m[2105]&~m[2106]&m[2107])|(m[910]&m[2103]&~m[2105]&~m[2106]&m[2107])|(m[910]&~m[2103]&m[2105]&~m[2106]&m[2107])|(~m[910]&~m[2103]&~m[2105]&m[2106]&m[2107])|(m[910]&~m[2103]&~m[2105]&m[2106]&m[2107])|(~m[910]&m[2103]&~m[2105]&m[2106]&m[2107])|(m[910]&m[2103]&~m[2105]&m[2106]&m[2107])|(~m[910]&~m[2103]&m[2105]&m[2106]&m[2107])|(m[910]&~m[2103]&m[2105]&m[2106]&m[2107])|(m[910]&m[2103]&m[2105]&m[2106]&m[2107]))):InitCond[1626];
    m[2109] = run?((((m[925]&~m[2108]&~m[2110]&~m[2111]&~m[2112])|(~m[925]&~m[2108]&~m[2110]&m[2111]&~m[2112])|(m[925]&m[2108]&~m[2110]&m[2111]&~m[2112])|(m[925]&~m[2108]&m[2110]&m[2111]&~m[2112])|(~m[925]&m[2108]&~m[2110]&~m[2111]&m[2112])|(~m[925]&~m[2108]&m[2110]&~m[2111]&m[2112])|(m[925]&m[2108]&m[2110]&~m[2111]&m[2112])|(~m[925]&m[2108]&m[2110]&m[2111]&m[2112]))&UnbiasedRNG[732])|((m[925]&~m[2108]&~m[2110]&m[2111]&~m[2112])|(~m[925]&~m[2108]&~m[2110]&~m[2111]&m[2112])|(m[925]&~m[2108]&~m[2110]&~m[2111]&m[2112])|(m[925]&m[2108]&~m[2110]&~m[2111]&m[2112])|(m[925]&~m[2108]&m[2110]&~m[2111]&m[2112])|(~m[925]&~m[2108]&~m[2110]&m[2111]&m[2112])|(m[925]&~m[2108]&~m[2110]&m[2111]&m[2112])|(~m[925]&m[2108]&~m[2110]&m[2111]&m[2112])|(m[925]&m[2108]&~m[2110]&m[2111]&m[2112])|(~m[925]&~m[2108]&m[2110]&m[2111]&m[2112])|(m[925]&~m[2108]&m[2110]&m[2111]&m[2112])|(m[925]&m[2108]&m[2110]&m[2111]&m[2112]))):InitCond[1627];
    m[2114] = run?((((m[911]&~m[2113]&~m[2115]&~m[2116]&~m[2117])|(~m[911]&~m[2113]&~m[2115]&m[2116]&~m[2117])|(m[911]&m[2113]&~m[2115]&m[2116]&~m[2117])|(m[911]&~m[2113]&m[2115]&m[2116]&~m[2117])|(~m[911]&m[2113]&~m[2115]&~m[2116]&m[2117])|(~m[911]&~m[2113]&m[2115]&~m[2116]&m[2117])|(m[911]&m[2113]&m[2115]&~m[2116]&m[2117])|(~m[911]&m[2113]&m[2115]&m[2116]&m[2117]))&UnbiasedRNG[733])|((m[911]&~m[2113]&~m[2115]&m[2116]&~m[2117])|(~m[911]&~m[2113]&~m[2115]&~m[2116]&m[2117])|(m[911]&~m[2113]&~m[2115]&~m[2116]&m[2117])|(m[911]&m[2113]&~m[2115]&~m[2116]&m[2117])|(m[911]&~m[2113]&m[2115]&~m[2116]&m[2117])|(~m[911]&~m[2113]&~m[2115]&m[2116]&m[2117])|(m[911]&~m[2113]&~m[2115]&m[2116]&m[2117])|(~m[911]&m[2113]&~m[2115]&m[2116]&m[2117])|(m[911]&m[2113]&~m[2115]&m[2116]&m[2117])|(~m[911]&~m[2113]&m[2115]&m[2116]&m[2117])|(m[911]&~m[2113]&m[2115]&m[2116]&m[2117])|(m[911]&m[2113]&m[2115]&m[2116]&m[2117]))):InitCond[1628];
    m[2119] = run?((((m[926]&~m[2118]&~m[2120]&~m[2121]&~m[2122])|(~m[926]&~m[2118]&~m[2120]&m[2121]&~m[2122])|(m[926]&m[2118]&~m[2120]&m[2121]&~m[2122])|(m[926]&~m[2118]&m[2120]&m[2121]&~m[2122])|(~m[926]&m[2118]&~m[2120]&~m[2121]&m[2122])|(~m[926]&~m[2118]&m[2120]&~m[2121]&m[2122])|(m[926]&m[2118]&m[2120]&~m[2121]&m[2122])|(~m[926]&m[2118]&m[2120]&m[2121]&m[2122]))&UnbiasedRNG[734])|((m[926]&~m[2118]&~m[2120]&m[2121]&~m[2122])|(~m[926]&~m[2118]&~m[2120]&~m[2121]&m[2122])|(m[926]&~m[2118]&~m[2120]&~m[2121]&m[2122])|(m[926]&m[2118]&~m[2120]&~m[2121]&m[2122])|(m[926]&~m[2118]&m[2120]&~m[2121]&m[2122])|(~m[926]&~m[2118]&~m[2120]&m[2121]&m[2122])|(m[926]&~m[2118]&~m[2120]&m[2121]&m[2122])|(~m[926]&m[2118]&~m[2120]&m[2121]&m[2122])|(m[926]&m[2118]&~m[2120]&m[2121]&m[2122])|(~m[926]&~m[2118]&m[2120]&m[2121]&m[2122])|(m[926]&~m[2118]&m[2120]&m[2121]&m[2122])|(m[926]&m[2118]&m[2120]&m[2121]&m[2122]))):InitCond[1629];
    m[2124] = run?((((m[927]&~m[2123]&~m[2125]&~m[2126]&~m[2127])|(~m[927]&~m[2123]&~m[2125]&m[2126]&~m[2127])|(m[927]&m[2123]&~m[2125]&m[2126]&~m[2127])|(m[927]&~m[2123]&m[2125]&m[2126]&~m[2127])|(~m[927]&m[2123]&~m[2125]&~m[2126]&m[2127])|(~m[927]&~m[2123]&m[2125]&~m[2126]&m[2127])|(m[927]&m[2123]&m[2125]&~m[2126]&m[2127])|(~m[927]&m[2123]&m[2125]&m[2126]&m[2127]))&UnbiasedRNG[735])|((m[927]&~m[2123]&~m[2125]&m[2126]&~m[2127])|(~m[927]&~m[2123]&~m[2125]&~m[2126]&m[2127])|(m[927]&~m[2123]&~m[2125]&~m[2126]&m[2127])|(m[927]&m[2123]&~m[2125]&~m[2126]&m[2127])|(m[927]&~m[2123]&m[2125]&~m[2126]&m[2127])|(~m[927]&~m[2123]&~m[2125]&m[2126]&m[2127])|(m[927]&~m[2123]&~m[2125]&m[2126]&m[2127])|(~m[927]&m[2123]&~m[2125]&m[2126]&m[2127])|(m[927]&m[2123]&~m[2125]&m[2126]&m[2127])|(~m[927]&~m[2123]&m[2125]&m[2126]&m[2127])|(m[927]&~m[2123]&m[2125]&m[2126]&m[2127])|(m[927]&m[2123]&m[2125]&m[2126]&m[2127]))):InitCond[1630];
end

always @(posedge color3_clk) begin
    m[936] = run?((((m[933]&~m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&~m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&m[937]&~m[938])|(~m[933]&~m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&m[937]&m[938])|(m[933]&~m[934]&m[935]&m[937]&m[938])|(~m[933]&m[934]&m[935]&m[937]&m[938]))&UnbiasedRNG[736])|((m[933]&m[934]&~m[935]&~m[937]&~m[938])|(m[933]&~m[934]&m[935]&~m[937]&~m[938])|(~m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&~m[934]&~m[935]&~m[937]&m[938])|(~m[933]&m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&~m[937]&m[938])|(~m[933]&~m[934]&m[935]&~m[937]&m[938])|(m[933]&~m[934]&m[935]&~m[937]&m[938])|(~m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&m[937]&m[938]))):InitCond[1631];
    m[946] = run?((((m[943]&~m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&~m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&m[947]&~m[948])|(~m[943]&~m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&m[947]&m[948])|(m[943]&~m[944]&m[945]&m[947]&m[948])|(~m[943]&m[944]&m[945]&m[947]&m[948]))&UnbiasedRNG[737])|((m[943]&m[944]&~m[945]&~m[947]&~m[948])|(m[943]&~m[944]&m[945]&~m[947]&~m[948])|(~m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&~m[944]&~m[945]&~m[947]&m[948])|(~m[943]&m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&~m[947]&m[948])|(~m[943]&~m[944]&m[945]&~m[947]&m[948])|(m[943]&~m[944]&m[945]&~m[947]&m[948])|(~m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&m[947]&m[948]))):InitCond[1632];
    m[951] = run?((((m[948]&~m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&~m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&m[952]&~m[953])|(~m[948]&~m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&m[952]&m[953])|(m[948]&~m[949]&m[950]&m[952]&m[953])|(~m[948]&m[949]&m[950]&m[952]&m[953]))&UnbiasedRNG[738])|((m[948]&m[949]&~m[950]&~m[952]&~m[953])|(m[948]&~m[949]&m[950]&~m[952]&~m[953])|(~m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&~m[949]&~m[950]&~m[952]&m[953])|(~m[948]&m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&~m[952]&m[953])|(~m[948]&~m[949]&m[950]&~m[952]&m[953])|(m[948]&~m[949]&m[950]&~m[952]&m[953])|(~m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&m[952]&m[953]))):InitCond[1633];
    m[961] = run?((((m[958]&~m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&~m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&m[962]&~m[963])|(~m[958]&~m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&m[962]&m[963])|(m[958]&~m[959]&m[960]&m[962]&m[963])|(~m[958]&m[959]&m[960]&m[962]&m[963]))&UnbiasedRNG[739])|((m[958]&m[959]&~m[960]&~m[962]&~m[963])|(m[958]&~m[959]&m[960]&~m[962]&~m[963])|(~m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&~m[959]&~m[960]&~m[962]&m[963])|(~m[958]&m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&~m[962]&m[963])|(~m[958]&~m[959]&m[960]&~m[962]&m[963])|(m[958]&~m[959]&m[960]&~m[962]&m[963])|(~m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&m[962]&m[963]))):InitCond[1634];
    m[966] = run?((((m[963]&~m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&~m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&m[967]&~m[968])|(~m[963]&~m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&m[967]&m[968])|(m[963]&~m[964]&m[965]&m[967]&m[968])|(~m[963]&m[964]&m[965]&m[967]&m[968]))&UnbiasedRNG[740])|((m[963]&m[964]&~m[965]&~m[967]&~m[968])|(m[963]&~m[964]&m[965]&~m[967]&~m[968])|(~m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&~m[964]&~m[965]&~m[967]&m[968])|(~m[963]&m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&~m[967]&m[968])|(~m[963]&~m[964]&m[965]&~m[967]&m[968])|(m[963]&~m[964]&m[965]&~m[967]&m[968])|(~m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&m[967]&m[968]))):InitCond[1635];
    m[971] = run?((((m[968]&~m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&~m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&m[972]&~m[973])|(~m[968]&~m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&m[972]&m[973])|(m[968]&~m[969]&m[970]&m[972]&m[973])|(~m[968]&m[969]&m[970]&m[972]&m[973]))&UnbiasedRNG[741])|((m[968]&m[969]&~m[970]&~m[972]&~m[973])|(m[968]&~m[969]&m[970]&~m[972]&~m[973])|(~m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&~m[969]&~m[970]&~m[972]&m[973])|(~m[968]&m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&~m[972]&m[973])|(~m[968]&~m[969]&m[970]&~m[972]&m[973])|(m[968]&~m[969]&m[970]&~m[972]&m[973])|(~m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&m[972]&m[973]))):InitCond[1636];
    m[981] = run?((((m[978]&~m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&~m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&m[982]&~m[983])|(~m[978]&~m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&m[982]&m[983])|(m[978]&~m[979]&m[980]&m[982]&m[983])|(~m[978]&m[979]&m[980]&m[982]&m[983]))&UnbiasedRNG[742])|((m[978]&m[979]&~m[980]&~m[982]&~m[983])|(m[978]&~m[979]&m[980]&~m[982]&~m[983])|(~m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&~m[979]&~m[980]&~m[982]&m[983])|(~m[978]&m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&~m[982]&m[983])|(~m[978]&~m[979]&m[980]&~m[982]&m[983])|(m[978]&~m[979]&m[980]&~m[982]&m[983])|(~m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&m[982]&m[983]))):InitCond[1637];
    m[986] = run?((((m[983]&~m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&~m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&m[987]&~m[988])|(~m[983]&~m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&m[987]&m[988])|(m[983]&~m[984]&m[985]&m[987]&m[988])|(~m[983]&m[984]&m[985]&m[987]&m[988]))&UnbiasedRNG[743])|((m[983]&m[984]&~m[985]&~m[987]&~m[988])|(m[983]&~m[984]&m[985]&~m[987]&~m[988])|(~m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&~m[984]&~m[985]&~m[987]&m[988])|(~m[983]&m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&~m[987]&m[988])|(~m[983]&~m[984]&m[985]&~m[987]&m[988])|(m[983]&~m[984]&m[985]&~m[987]&m[988])|(~m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&m[987]&m[988]))):InitCond[1638];
    m[991] = run?((((m[988]&~m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&~m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&m[992]&~m[993])|(~m[988]&~m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&m[992]&m[993])|(m[988]&~m[989]&m[990]&m[992]&m[993])|(~m[988]&m[989]&m[990]&m[992]&m[993]))&UnbiasedRNG[744])|((m[988]&m[989]&~m[990]&~m[992]&~m[993])|(m[988]&~m[989]&m[990]&~m[992]&~m[993])|(~m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&~m[989]&~m[990]&~m[992]&m[993])|(~m[988]&m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&~m[992]&m[993])|(~m[988]&~m[989]&m[990]&~m[992]&m[993])|(m[988]&~m[989]&m[990]&~m[992]&m[993])|(~m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&m[992]&m[993]))):InitCond[1639];
    m[996] = run?((((m[993]&~m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&~m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&m[997]&~m[998])|(~m[993]&~m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&m[997]&m[998])|(m[993]&~m[994]&m[995]&m[997]&m[998])|(~m[993]&m[994]&m[995]&m[997]&m[998]))&UnbiasedRNG[745])|((m[993]&m[994]&~m[995]&~m[997]&~m[998])|(m[993]&~m[994]&m[995]&~m[997]&~m[998])|(~m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&~m[994]&~m[995]&~m[997]&m[998])|(~m[993]&m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&~m[997]&m[998])|(~m[993]&~m[994]&m[995]&~m[997]&m[998])|(m[993]&~m[994]&m[995]&~m[997]&m[998])|(~m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&m[997]&m[998]))):InitCond[1640];
    m[1006] = run?((((m[1003]&~m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&~m[1008])|(~m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&m[1007]&m[1008]))&UnbiasedRNG[746])|((m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&m[1008]))):InitCond[1641];
    m[1011] = run?((((m[1008]&~m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&~m[1013])|(~m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))&UnbiasedRNG[747])|((m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))):InitCond[1642];
    m[1016] = run?((((m[1013]&~m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&~m[1018])|(~m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))&UnbiasedRNG[748])|((m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))):InitCond[1643];
    m[1021] = run?((((m[1018]&~m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&~m[1023])|(~m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))&UnbiasedRNG[749])|((m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))):InitCond[1644];
    m[1026] = run?((((m[1023]&~m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&~m[1028])|(~m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))&UnbiasedRNG[750])|((m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))):InitCond[1645];
    m[1036] = run?((((m[1033]&~m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&~m[1038])|(~m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))&UnbiasedRNG[751])|((m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))):InitCond[1646];
    m[1041] = run?((((m[1038]&~m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&~m[1043])|(~m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))&UnbiasedRNG[752])|((m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))):InitCond[1647];
    m[1046] = run?((((m[1043]&~m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&~m[1048])|(~m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&m[1047]&m[1048]))&UnbiasedRNG[753])|((m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&m[1048]))):InitCond[1648];
    m[1051] = run?((((m[1048]&~m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&~m[1053])|(~m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))&UnbiasedRNG[754])|((m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))):InitCond[1649];
    m[1056] = run?((((m[1053]&~m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&~m[1058])|(~m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&m[1057]&m[1058]))&UnbiasedRNG[755])|((m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&m[1058]))):InitCond[1650];
    m[1061] = run?((((m[1058]&~m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&~m[1063])|(~m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))&UnbiasedRNG[756])|((m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))):InitCond[1651];
    m[1071] = run?((((m[1068]&~m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&~m[1073])|(~m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))&UnbiasedRNG[757])|((m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))):InitCond[1652];
    m[1076] = run?((((m[1073]&~m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&~m[1078])|(~m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))&UnbiasedRNG[758])|((m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))):InitCond[1653];
    m[1081] = run?((((m[1078]&~m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&~m[1083])|(~m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&m[1082]&m[1083]))&UnbiasedRNG[759])|((m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&m[1083]))):InitCond[1654];
    m[1086] = run?((((m[1083]&~m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&~m[1088])|(~m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))&UnbiasedRNG[760])|((m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))):InitCond[1655];
    m[1091] = run?((((m[1088]&~m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&~m[1093])|(~m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))&UnbiasedRNG[761])|((m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))):InitCond[1656];
    m[1096] = run?((((m[1093]&~m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&~m[1098])|(~m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))&UnbiasedRNG[762])|((m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))):InitCond[1657];
    m[1101] = run?((((m[1098]&~m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&~m[1103])|(~m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))&UnbiasedRNG[763])|((m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))):InitCond[1658];
    m[1111] = run?((((m[1108]&~m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&~m[1113])|(~m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&m[1112]&m[1113]))&UnbiasedRNG[764])|((m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&m[1113]))):InitCond[1659];
    m[1116] = run?((((m[1113]&~m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&~m[1118])|(~m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&m[1117]&m[1118]))&UnbiasedRNG[765])|((m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&m[1118]))):InitCond[1660];
    m[1121] = run?((((m[1118]&~m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&~m[1123])|(~m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))&UnbiasedRNG[766])|((m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))):InitCond[1661];
    m[1126] = run?((((m[1123]&~m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&~m[1128])|(~m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))&UnbiasedRNG[767])|((m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))):InitCond[1662];
    m[1131] = run?((((m[1128]&~m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&~m[1133])|(~m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))&UnbiasedRNG[768])|((m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))):InitCond[1663];
    m[1136] = run?((((m[1133]&~m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&~m[1138])|(~m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&m[1137]&m[1138]))&UnbiasedRNG[769])|((m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&m[1138]))):InitCond[1664];
    m[1141] = run?((((m[1138]&~m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&~m[1143])|(~m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))&UnbiasedRNG[770])|((m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))):InitCond[1665];
    m[1146] = run?((((m[1143]&~m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&~m[1148])|(~m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))&UnbiasedRNG[771])|((m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))):InitCond[1666];
    m[1156] = run?((((m[1153]&~m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&~m[1158])|(~m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&m[1157]&m[1158]))&UnbiasedRNG[772])|((m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&m[1158]))):InitCond[1667];
    m[1161] = run?((((m[1158]&~m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&~m[1163])|(~m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))&UnbiasedRNG[773])|((m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))):InitCond[1668];
    m[1166] = run?((((m[1163]&~m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&~m[1168])|(~m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))&UnbiasedRNG[774])|((m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))):InitCond[1669];
    m[1171] = run?((((m[1168]&~m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&~m[1173])|(~m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&m[1172]&m[1173]))&UnbiasedRNG[775])|((m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&m[1173]))):InitCond[1670];
    m[1176] = run?((((m[1173]&~m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&~m[1178])|(~m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))&UnbiasedRNG[776])|((m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))):InitCond[1671];
    m[1181] = run?((((m[1178]&~m[1179]&~m[1180]&~m[1182]&~m[1183])|(~m[1178]&m[1179]&~m[1180]&~m[1182]&~m[1183])|(~m[1178]&~m[1179]&m[1180]&~m[1182]&~m[1183])|(m[1178]&m[1179]&m[1180]&m[1182]&~m[1183])|(~m[1178]&~m[1179]&~m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&~m[1180]&m[1182]&m[1183])|(m[1178]&~m[1179]&m[1180]&m[1182]&m[1183])|(~m[1178]&m[1179]&m[1180]&m[1182]&m[1183]))&UnbiasedRNG[777])|((m[1178]&m[1179]&~m[1180]&~m[1182]&~m[1183])|(m[1178]&~m[1179]&m[1180]&~m[1182]&~m[1183])|(~m[1178]&m[1179]&m[1180]&~m[1182]&~m[1183])|(m[1178]&m[1179]&m[1180]&~m[1182]&~m[1183])|(m[1178]&~m[1179]&~m[1180]&~m[1182]&m[1183])|(~m[1178]&m[1179]&~m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&~m[1180]&~m[1182]&m[1183])|(~m[1178]&~m[1179]&m[1180]&~m[1182]&m[1183])|(m[1178]&~m[1179]&m[1180]&~m[1182]&m[1183])|(~m[1178]&m[1179]&m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&m[1180]&~m[1182]&m[1183])|(m[1178]&m[1179]&m[1180]&m[1182]&m[1183]))):InitCond[1672];
    m[1186] = run?((((m[1183]&~m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&~m[1188])|(~m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&m[1187]&m[1188]))&UnbiasedRNG[778])|((m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&m[1188]))):InitCond[1673];
    m[1191] = run?((((m[1188]&~m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&~m[1193])|(~m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&m[1192]&m[1193]))&UnbiasedRNG[779])|((m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&m[1193]))):InitCond[1674];
    m[1196] = run?((((m[1193]&~m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&~m[1198])|(~m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&m[1197]&m[1198]))&UnbiasedRNG[780])|((m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&m[1198]))):InitCond[1675];
    m[1206] = run?((((m[1203]&~m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&~m[1208])|(~m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&m[1207]&m[1208]))&UnbiasedRNG[781])|((m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&m[1208]))):InitCond[1676];
    m[1211] = run?((((m[1208]&~m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&~m[1213])|(~m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&m[1212]&m[1213]))&UnbiasedRNG[782])|((m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&m[1213]))):InitCond[1677];
    m[1216] = run?((((m[1213]&~m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&~m[1218])|(~m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&m[1217]&m[1218]))&UnbiasedRNG[783])|((m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&m[1218]))):InitCond[1678];
    m[1221] = run?((((m[1218]&~m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&~m[1223])|(~m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&m[1222]&m[1223]))&UnbiasedRNG[784])|((m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&m[1223]))):InitCond[1679];
    m[1226] = run?((((m[1223]&~m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&~m[1228])|(~m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&m[1227]&m[1228]))&UnbiasedRNG[785])|((m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&m[1228]))):InitCond[1680];
    m[1231] = run?((((m[1228]&~m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&~m[1233])|(~m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&m[1232]&m[1233]))&UnbiasedRNG[786])|((m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&m[1233]))):InitCond[1681];
    m[1236] = run?((((m[1233]&~m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&~m[1238])|(~m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&m[1237]&m[1238]))&UnbiasedRNG[787])|((m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&m[1238]))):InitCond[1682];
    m[1241] = run?((((m[1238]&~m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&~m[1243])|(~m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&m[1242]&m[1243]))&UnbiasedRNG[788])|((m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&m[1243]))):InitCond[1683];
    m[1246] = run?((((m[1243]&~m[1244]&~m[1245]&~m[1247]&~m[1248])|(~m[1243]&m[1244]&~m[1245]&~m[1247]&~m[1248])|(~m[1243]&~m[1244]&m[1245]&~m[1247]&~m[1248])|(m[1243]&m[1244]&m[1245]&m[1247]&~m[1248])|(~m[1243]&~m[1244]&~m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&~m[1245]&m[1247]&m[1248])|(m[1243]&~m[1244]&m[1245]&m[1247]&m[1248])|(~m[1243]&m[1244]&m[1245]&m[1247]&m[1248]))&UnbiasedRNG[789])|((m[1243]&m[1244]&~m[1245]&~m[1247]&~m[1248])|(m[1243]&~m[1244]&m[1245]&~m[1247]&~m[1248])|(~m[1243]&m[1244]&m[1245]&~m[1247]&~m[1248])|(m[1243]&m[1244]&m[1245]&~m[1247]&~m[1248])|(m[1243]&~m[1244]&~m[1245]&~m[1247]&m[1248])|(~m[1243]&m[1244]&~m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&~m[1245]&~m[1247]&m[1248])|(~m[1243]&~m[1244]&m[1245]&~m[1247]&m[1248])|(m[1243]&~m[1244]&m[1245]&~m[1247]&m[1248])|(~m[1243]&m[1244]&m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&m[1245]&~m[1247]&m[1248])|(m[1243]&m[1244]&m[1245]&m[1247]&m[1248]))):InitCond[1684];
    m[1251] = run?((((m[1248]&~m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&~m[1253])|(~m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&m[1252]&m[1253]))&UnbiasedRNG[790])|((m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&m[1253]))):InitCond[1685];
    m[1261] = run?((((m[1258]&~m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&~m[1263])|(~m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&m[1262]&m[1263]))&UnbiasedRNG[791])|((m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&m[1263]))):InitCond[1686];
    m[1266] = run?((((m[1263]&~m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&~m[1268])|(~m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&m[1267]&m[1268]))&UnbiasedRNG[792])|((m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&m[1268]))):InitCond[1687];
    m[1271] = run?((((m[1268]&~m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&~m[1273])|(~m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&m[1272]&m[1273]))&UnbiasedRNG[793])|((m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&m[1273]))):InitCond[1688];
    m[1276] = run?((((m[1273]&~m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&~m[1278])|(~m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&m[1277]&m[1278]))&UnbiasedRNG[794])|((m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&m[1278]))):InitCond[1689];
    m[1281] = run?((((m[1278]&~m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&~m[1283])|(~m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&m[1282]&m[1283]))&UnbiasedRNG[795])|((m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&m[1283]))):InitCond[1690];
    m[1286] = run?((((m[1283]&~m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&~m[1288])|(~m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&m[1287]&m[1288]))&UnbiasedRNG[796])|((m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&m[1288]))):InitCond[1691];
    m[1291] = run?((((m[1288]&~m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&~m[1293])|(~m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&m[1292]&m[1293]))&UnbiasedRNG[797])|((m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&m[1293]))):InitCond[1692];
    m[1296] = run?((((m[1293]&~m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&~m[1298])|(~m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&m[1297]&m[1298]))&UnbiasedRNG[798])|((m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&m[1298]))):InitCond[1693];
    m[1301] = run?((((m[1298]&~m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&~m[1303])|(~m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&m[1302]&m[1303]))&UnbiasedRNG[799])|((m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&m[1303]))):InitCond[1694];
    m[1306] = run?((((m[1303]&~m[1304]&~m[1305]&~m[1307]&~m[1308])|(~m[1303]&m[1304]&~m[1305]&~m[1307]&~m[1308])|(~m[1303]&~m[1304]&m[1305]&~m[1307]&~m[1308])|(m[1303]&m[1304]&m[1305]&m[1307]&~m[1308])|(~m[1303]&~m[1304]&~m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&~m[1305]&m[1307]&m[1308])|(m[1303]&~m[1304]&m[1305]&m[1307]&m[1308])|(~m[1303]&m[1304]&m[1305]&m[1307]&m[1308]))&UnbiasedRNG[800])|((m[1303]&m[1304]&~m[1305]&~m[1307]&~m[1308])|(m[1303]&~m[1304]&m[1305]&~m[1307]&~m[1308])|(~m[1303]&m[1304]&m[1305]&~m[1307]&~m[1308])|(m[1303]&m[1304]&m[1305]&~m[1307]&~m[1308])|(m[1303]&~m[1304]&~m[1305]&~m[1307]&m[1308])|(~m[1303]&m[1304]&~m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&~m[1305]&~m[1307]&m[1308])|(~m[1303]&~m[1304]&m[1305]&~m[1307]&m[1308])|(m[1303]&~m[1304]&m[1305]&~m[1307]&m[1308])|(~m[1303]&m[1304]&m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&m[1305]&~m[1307]&m[1308])|(m[1303]&m[1304]&m[1305]&m[1307]&m[1308]))):InitCond[1695];
    m[1311] = run?((((m[1308]&~m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&~m[1313])|(~m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&m[1312]&m[1313]))&UnbiasedRNG[801])|((m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&m[1313]))):InitCond[1696];
    m[1321] = run?((((m[1318]&~m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&~m[1323])|(~m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&m[1322]&m[1323]))&UnbiasedRNG[802])|((m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&m[1323]))):InitCond[1697];
    m[1326] = run?((((m[1323]&~m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&~m[1328])|(~m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&m[1327]&m[1328]))&UnbiasedRNG[803])|((m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&m[1328]))):InitCond[1698];
    m[1331] = run?((((m[1328]&~m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&~m[1333])|(~m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&m[1332]&m[1333]))&UnbiasedRNG[804])|((m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&m[1333]))):InitCond[1699];
    m[1336] = run?((((m[1333]&~m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&~m[1338])|(~m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&m[1337]&m[1338]))&UnbiasedRNG[805])|((m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&m[1338]))):InitCond[1700];
    m[1341] = run?((((m[1338]&~m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&~m[1343])|(~m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&m[1342]&m[1343]))&UnbiasedRNG[806])|((m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&m[1343]))):InitCond[1701];
    m[1346] = run?((((m[1343]&~m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&~m[1348])|(~m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&m[1347]&m[1348]))&UnbiasedRNG[807])|((m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&m[1348]))):InitCond[1702];
    m[1351] = run?((((m[1348]&~m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&~m[1353])|(~m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&m[1352]&m[1353]))&UnbiasedRNG[808])|((m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&m[1353]))):InitCond[1703];
    m[1356] = run?((((m[1353]&~m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&~m[1358])|(~m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&m[1357]&m[1358]))&UnbiasedRNG[809])|((m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&m[1358]))):InitCond[1704];
    m[1361] = run?((((m[1358]&~m[1359]&~m[1360]&~m[1362]&~m[1363])|(~m[1358]&m[1359]&~m[1360]&~m[1362]&~m[1363])|(~m[1358]&~m[1359]&m[1360]&~m[1362]&~m[1363])|(m[1358]&m[1359]&m[1360]&m[1362]&~m[1363])|(~m[1358]&~m[1359]&~m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&~m[1360]&m[1362]&m[1363])|(m[1358]&~m[1359]&m[1360]&m[1362]&m[1363])|(~m[1358]&m[1359]&m[1360]&m[1362]&m[1363]))&UnbiasedRNG[810])|((m[1358]&m[1359]&~m[1360]&~m[1362]&~m[1363])|(m[1358]&~m[1359]&m[1360]&~m[1362]&~m[1363])|(~m[1358]&m[1359]&m[1360]&~m[1362]&~m[1363])|(m[1358]&m[1359]&m[1360]&~m[1362]&~m[1363])|(m[1358]&~m[1359]&~m[1360]&~m[1362]&m[1363])|(~m[1358]&m[1359]&~m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&~m[1360]&~m[1362]&m[1363])|(~m[1358]&~m[1359]&m[1360]&~m[1362]&m[1363])|(m[1358]&~m[1359]&m[1360]&~m[1362]&m[1363])|(~m[1358]&m[1359]&m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&m[1360]&~m[1362]&m[1363])|(m[1358]&m[1359]&m[1360]&m[1362]&m[1363]))):InitCond[1705];
    m[1366] = run?((((m[1363]&~m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&~m[1368])|(~m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&m[1367]&m[1368]))&UnbiasedRNG[811])|((m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&m[1368]))):InitCond[1706];
    m[1371] = run?((((m[1368]&~m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&~m[1373])|(~m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&m[1372]&m[1373]))&UnbiasedRNG[812])|((m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&m[1373]))):InitCond[1707];
    m[1376] = run?((((m[1373]&~m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&~m[1378])|(~m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&m[1377]&m[1378]))&UnbiasedRNG[813])|((m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&m[1378]))):InitCond[1708];
    m[1386] = run?((((m[1383]&~m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&~m[1388])|(~m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&m[1387]&m[1388]))&UnbiasedRNG[814])|((m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&m[1388]))):InitCond[1709];
    m[1391] = run?((((m[1388]&~m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&~m[1393])|(~m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&m[1392]&m[1393]))&UnbiasedRNG[815])|((m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&m[1393]))):InitCond[1710];
    m[1396] = run?((((m[1393]&~m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&~m[1398])|(~m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&m[1397]&m[1398]))&UnbiasedRNG[816])|((m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&m[1398]))):InitCond[1711];
    m[1401] = run?((((m[1398]&~m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&~m[1403])|(~m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&m[1402]&m[1403]))&UnbiasedRNG[817])|((m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&m[1403]))):InitCond[1712];
    m[1406] = run?((((m[1403]&~m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&~m[1408])|(~m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&m[1407]&m[1408]))&UnbiasedRNG[818])|((m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&m[1408]))):InitCond[1713];
    m[1411] = run?((((m[1408]&~m[1409]&~m[1410]&~m[1412]&~m[1413])|(~m[1408]&m[1409]&~m[1410]&~m[1412]&~m[1413])|(~m[1408]&~m[1409]&m[1410]&~m[1412]&~m[1413])|(m[1408]&m[1409]&m[1410]&m[1412]&~m[1413])|(~m[1408]&~m[1409]&~m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&~m[1410]&m[1412]&m[1413])|(m[1408]&~m[1409]&m[1410]&m[1412]&m[1413])|(~m[1408]&m[1409]&m[1410]&m[1412]&m[1413]))&UnbiasedRNG[819])|((m[1408]&m[1409]&~m[1410]&~m[1412]&~m[1413])|(m[1408]&~m[1409]&m[1410]&~m[1412]&~m[1413])|(~m[1408]&m[1409]&m[1410]&~m[1412]&~m[1413])|(m[1408]&m[1409]&m[1410]&~m[1412]&~m[1413])|(m[1408]&~m[1409]&~m[1410]&~m[1412]&m[1413])|(~m[1408]&m[1409]&~m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&~m[1410]&~m[1412]&m[1413])|(~m[1408]&~m[1409]&m[1410]&~m[1412]&m[1413])|(m[1408]&~m[1409]&m[1410]&~m[1412]&m[1413])|(~m[1408]&m[1409]&m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&m[1410]&~m[1412]&m[1413])|(m[1408]&m[1409]&m[1410]&m[1412]&m[1413]))):InitCond[1714];
    m[1416] = run?((((m[1413]&~m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&~m[1418])|(~m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&m[1417]&m[1418]))&UnbiasedRNG[820])|((m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&m[1418]))):InitCond[1715];
    m[1421] = run?((((m[1418]&~m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&~m[1423])|(~m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&m[1422]&m[1423]))&UnbiasedRNG[821])|((m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&m[1423]))):InitCond[1716];
    m[1426] = run?((((m[1423]&~m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&~m[1428])|(~m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&m[1427]&m[1428]))&UnbiasedRNG[822])|((m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&m[1428]))):InitCond[1717];
    m[1431] = run?((((m[1428]&~m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&~m[1433])|(~m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&m[1432]&m[1433]))&UnbiasedRNG[823])|((m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&m[1433]))):InitCond[1718];
    m[1436] = run?((((m[1433]&~m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&~m[1438])|(~m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&m[1437]&m[1438]))&UnbiasedRNG[824])|((m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&m[1438]))):InitCond[1719];
    m[1441] = run?((((m[1438]&~m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&~m[1443])|(~m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&m[1442]&m[1443]))&UnbiasedRNG[825])|((m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&m[1443]))):InitCond[1720];
    m[1446] = run?((((m[1443]&~m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&~m[1448])|(~m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&m[1447]&m[1448]))&UnbiasedRNG[826])|((m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&m[1448]))):InitCond[1721];
    m[1456] = run?((((m[1453]&~m[1454]&~m[1455]&~m[1457]&~m[1458])|(~m[1453]&m[1454]&~m[1455]&~m[1457]&~m[1458])|(~m[1453]&~m[1454]&m[1455]&~m[1457]&~m[1458])|(m[1453]&m[1454]&m[1455]&m[1457]&~m[1458])|(~m[1453]&~m[1454]&~m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&~m[1455]&m[1457]&m[1458])|(m[1453]&~m[1454]&m[1455]&m[1457]&m[1458])|(~m[1453]&m[1454]&m[1455]&m[1457]&m[1458]))&UnbiasedRNG[827])|((m[1453]&m[1454]&~m[1455]&~m[1457]&~m[1458])|(m[1453]&~m[1454]&m[1455]&~m[1457]&~m[1458])|(~m[1453]&m[1454]&m[1455]&~m[1457]&~m[1458])|(m[1453]&m[1454]&m[1455]&~m[1457]&~m[1458])|(m[1453]&~m[1454]&~m[1455]&~m[1457]&m[1458])|(~m[1453]&m[1454]&~m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&~m[1455]&~m[1457]&m[1458])|(~m[1453]&~m[1454]&m[1455]&~m[1457]&m[1458])|(m[1453]&~m[1454]&m[1455]&~m[1457]&m[1458])|(~m[1453]&m[1454]&m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&m[1455]&~m[1457]&m[1458])|(m[1453]&m[1454]&m[1455]&m[1457]&m[1458]))):InitCond[1722];
    m[1461] = run?((((m[1458]&~m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&~m[1463])|(~m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&m[1462]&m[1463]))&UnbiasedRNG[828])|((m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&m[1463]))):InitCond[1723];
    m[1466] = run?((((m[1463]&~m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&~m[1468])|(~m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&m[1467]&m[1468]))&UnbiasedRNG[829])|((m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&m[1468]))):InitCond[1724];
    m[1471] = run?((((m[1468]&~m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&~m[1473])|(~m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&m[1472]&m[1473]))&UnbiasedRNG[830])|((m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&m[1473]))):InitCond[1725];
    m[1476] = run?((((m[1473]&~m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&~m[1478])|(~m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&m[1477]&m[1478]))&UnbiasedRNG[831])|((m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&m[1478]))):InitCond[1726];
    m[1481] = run?((((m[1478]&~m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&~m[1483])|(~m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&m[1482]&m[1483]))&UnbiasedRNG[832])|((m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&m[1483]))):InitCond[1727];
    m[1486] = run?((((m[1483]&~m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&~m[1488])|(~m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&m[1487]&m[1488]))&UnbiasedRNG[833])|((m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&m[1488]))):InitCond[1728];
    m[1491] = run?((((m[1488]&~m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&~m[1493])|(~m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&m[1492]&m[1493]))&UnbiasedRNG[834])|((m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&m[1493]))):InitCond[1729];
    m[1496] = run?((((m[1493]&~m[1494]&~m[1495]&~m[1497]&~m[1498])|(~m[1493]&m[1494]&~m[1495]&~m[1497]&~m[1498])|(~m[1493]&~m[1494]&m[1495]&~m[1497]&~m[1498])|(m[1493]&m[1494]&m[1495]&m[1497]&~m[1498])|(~m[1493]&~m[1494]&~m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&~m[1495]&m[1497]&m[1498])|(m[1493]&~m[1494]&m[1495]&m[1497]&m[1498])|(~m[1493]&m[1494]&m[1495]&m[1497]&m[1498]))&UnbiasedRNG[835])|((m[1493]&m[1494]&~m[1495]&~m[1497]&~m[1498])|(m[1493]&~m[1494]&m[1495]&~m[1497]&~m[1498])|(~m[1493]&m[1494]&m[1495]&~m[1497]&~m[1498])|(m[1493]&m[1494]&m[1495]&~m[1497]&~m[1498])|(m[1493]&~m[1494]&~m[1495]&~m[1497]&m[1498])|(~m[1493]&m[1494]&~m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&~m[1495]&~m[1497]&m[1498])|(~m[1493]&~m[1494]&m[1495]&~m[1497]&m[1498])|(m[1493]&~m[1494]&m[1495]&~m[1497]&m[1498])|(~m[1493]&m[1494]&m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&m[1495]&~m[1497]&m[1498])|(m[1493]&m[1494]&m[1495]&m[1497]&m[1498]))):InitCond[1730];
    m[1501] = run?((((m[1498]&~m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&~m[1503])|(~m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&m[1502]&m[1503]))&UnbiasedRNG[836])|((m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&m[1503]))):InitCond[1731];
    m[1506] = run?((((m[1503]&~m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&~m[1508])|(~m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&m[1507]&m[1508]))&UnbiasedRNG[837])|((m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&m[1508]))):InitCond[1732];
    m[1511] = run?((((m[1508]&~m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&~m[1513])|(~m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&m[1512]&m[1513]))&UnbiasedRNG[838])|((m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&m[1513]))):InitCond[1733];
    m[1516] = run?((((m[1513]&~m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&~m[1518])|(~m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&m[1517]&m[1518]))&UnbiasedRNG[839])|((m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&m[1518]))):InitCond[1734];
    m[1521] = run?((((m[1518]&~m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&~m[1523])|(~m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&m[1522]&m[1523]))&UnbiasedRNG[840])|((m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&m[1523]))):InitCond[1735];
    m[1531] = run?((((m[1528]&~m[1529]&~m[1530]&~m[1532]&~m[1533])|(~m[1528]&m[1529]&~m[1530]&~m[1532]&~m[1533])|(~m[1528]&~m[1529]&m[1530]&~m[1532]&~m[1533])|(m[1528]&m[1529]&m[1530]&m[1532]&~m[1533])|(~m[1528]&~m[1529]&~m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&~m[1530]&m[1532]&m[1533])|(m[1528]&~m[1529]&m[1530]&m[1532]&m[1533])|(~m[1528]&m[1529]&m[1530]&m[1532]&m[1533]))&UnbiasedRNG[841])|((m[1528]&m[1529]&~m[1530]&~m[1532]&~m[1533])|(m[1528]&~m[1529]&m[1530]&~m[1532]&~m[1533])|(~m[1528]&m[1529]&m[1530]&~m[1532]&~m[1533])|(m[1528]&m[1529]&m[1530]&~m[1532]&~m[1533])|(m[1528]&~m[1529]&~m[1530]&~m[1532]&m[1533])|(~m[1528]&m[1529]&~m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&~m[1530]&~m[1532]&m[1533])|(~m[1528]&~m[1529]&m[1530]&~m[1532]&m[1533])|(m[1528]&~m[1529]&m[1530]&~m[1532]&m[1533])|(~m[1528]&m[1529]&m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&m[1530]&~m[1532]&m[1533])|(m[1528]&m[1529]&m[1530]&m[1532]&m[1533]))):InitCond[1736];
    m[1536] = run?((((m[1533]&~m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&~m[1538])|(~m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&m[1537]&m[1538]))&UnbiasedRNG[842])|((m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&m[1538]))):InitCond[1737];
    m[1541] = run?((((m[1538]&~m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&~m[1543])|(~m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&m[1542]&m[1543]))&UnbiasedRNG[843])|((m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&m[1543]))):InitCond[1738];
    m[1546] = run?((((m[1543]&~m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&~m[1548])|(~m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&m[1547]&m[1548]))&UnbiasedRNG[844])|((m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&m[1548]))):InitCond[1739];
    m[1551] = run?((((m[1548]&~m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&~m[1553])|(~m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&m[1552]&m[1553]))&UnbiasedRNG[845])|((m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&m[1553]))):InitCond[1740];
    m[1556] = run?((((m[1553]&~m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&~m[1558])|(~m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&m[1557]&m[1558]))&UnbiasedRNG[846])|((m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&m[1558]))):InitCond[1741];
    m[1561] = run?((((m[1558]&~m[1559]&~m[1560]&~m[1562]&~m[1563])|(~m[1558]&m[1559]&~m[1560]&~m[1562]&~m[1563])|(~m[1558]&~m[1559]&m[1560]&~m[1562]&~m[1563])|(m[1558]&m[1559]&m[1560]&m[1562]&~m[1563])|(~m[1558]&~m[1559]&~m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&~m[1560]&m[1562]&m[1563])|(m[1558]&~m[1559]&m[1560]&m[1562]&m[1563])|(~m[1558]&m[1559]&m[1560]&m[1562]&m[1563]))&UnbiasedRNG[847])|((m[1558]&m[1559]&~m[1560]&~m[1562]&~m[1563])|(m[1558]&~m[1559]&m[1560]&~m[1562]&~m[1563])|(~m[1558]&m[1559]&m[1560]&~m[1562]&~m[1563])|(m[1558]&m[1559]&m[1560]&~m[1562]&~m[1563])|(m[1558]&~m[1559]&~m[1560]&~m[1562]&m[1563])|(~m[1558]&m[1559]&~m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&~m[1560]&~m[1562]&m[1563])|(~m[1558]&~m[1559]&m[1560]&~m[1562]&m[1563])|(m[1558]&~m[1559]&m[1560]&~m[1562]&m[1563])|(~m[1558]&m[1559]&m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&m[1560]&~m[1562]&m[1563])|(m[1558]&m[1559]&m[1560]&m[1562]&m[1563]))):InitCond[1742];
    m[1566] = run?((((m[1563]&~m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&~m[1568])|(~m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&m[1567]&m[1568]))&UnbiasedRNG[848])|((m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&m[1568]))):InitCond[1743];
    m[1571] = run?((((m[1568]&~m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&~m[1573])|(~m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&m[1572]&m[1573]))&UnbiasedRNG[849])|((m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&m[1573]))):InitCond[1744];
    m[1576] = run?((((m[1573]&~m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&~m[1578])|(~m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&m[1577]&m[1578]))&UnbiasedRNG[850])|((m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&m[1578]))):InitCond[1745];
    m[1581] = run?((((m[1578]&~m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&~m[1583])|(~m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&m[1582]&m[1583]))&UnbiasedRNG[851])|((m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&m[1583]))):InitCond[1746];
    m[1586] = run?((((m[1583]&~m[1584]&~m[1585]&~m[1587]&~m[1588])|(~m[1583]&m[1584]&~m[1585]&~m[1587]&~m[1588])|(~m[1583]&~m[1584]&m[1585]&~m[1587]&~m[1588])|(m[1583]&m[1584]&m[1585]&m[1587]&~m[1588])|(~m[1583]&~m[1584]&~m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&~m[1585]&m[1587]&m[1588])|(m[1583]&~m[1584]&m[1585]&m[1587]&m[1588])|(~m[1583]&m[1584]&m[1585]&m[1587]&m[1588]))&UnbiasedRNG[852])|((m[1583]&m[1584]&~m[1585]&~m[1587]&~m[1588])|(m[1583]&~m[1584]&m[1585]&~m[1587]&~m[1588])|(~m[1583]&m[1584]&m[1585]&~m[1587]&~m[1588])|(m[1583]&m[1584]&m[1585]&~m[1587]&~m[1588])|(m[1583]&~m[1584]&~m[1585]&~m[1587]&m[1588])|(~m[1583]&m[1584]&~m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&~m[1585]&~m[1587]&m[1588])|(~m[1583]&~m[1584]&m[1585]&~m[1587]&m[1588])|(m[1583]&~m[1584]&m[1585]&~m[1587]&m[1588])|(~m[1583]&m[1584]&m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&m[1585]&~m[1587]&m[1588])|(m[1583]&m[1584]&m[1585]&m[1587]&m[1588]))):InitCond[1747];
    m[1591] = run?((((m[1588]&~m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&~m[1593])|(~m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&m[1592]&m[1593]))&UnbiasedRNG[853])|((m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&m[1593]))):InitCond[1748];
    m[1596] = run?((((m[1593]&~m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&~m[1598])|(~m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&m[1597]&m[1598]))&UnbiasedRNG[854])|((m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&m[1598]))):InitCond[1749];
    m[1606] = run?((((m[1603]&~m[1604]&~m[1605]&~m[1607]&~m[1608])|(~m[1603]&m[1604]&~m[1605]&~m[1607]&~m[1608])|(~m[1603]&~m[1604]&m[1605]&~m[1607]&~m[1608])|(m[1603]&m[1604]&m[1605]&m[1607]&~m[1608])|(~m[1603]&~m[1604]&~m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&~m[1605]&m[1607]&m[1608])|(m[1603]&~m[1604]&m[1605]&m[1607]&m[1608])|(~m[1603]&m[1604]&m[1605]&m[1607]&m[1608]))&UnbiasedRNG[855])|((m[1603]&m[1604]&~m[1605]&~m[1607]&~m[1608])|(m[1603]&~m[1604]&m[1605]&~m[1607]&~m[1608])|(~m[1603]&m[1604]&m[1605]&~m[1607]&~m[1608])|(m[1603]&m[1604]&m[1605]&~m[1607]&~m[1608])|(m[1603]&~m[1604]&~m[1605]&~m[1607]&m[1608])|(~m[1603]&m[1604]&~m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&~m[1605]&~m[1607]&m[1608])|(~m[1603]&~m[1604]&m[1605]&~m[1607]&m[1608])|(m[1603]&~m[1604]&m[1605]&~m[1607]&m[1608])|(~m[1603]&m[1604]&m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&m[1605]&~m[1607]&m[1608])|(m[1603]&m[1604]&m[1605]&m[1607]&m[1608]))):InitCond[1750];
    m[1611] = run?((((m[1608]&~m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&~m[1613])|(~m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&m[1612]&m[1613]))&UnbiasedRNG[856])|((m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&m[1613]))):InitCond[1751];
    m[1616] = run?((((m[1613]&~m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&~m[1618])|(~m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&m[1617]&m[1618]))&UnbiasedRNG[857])|((m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&m[1618]))):InitCond[1752];
    m[1621] = run?((((m[1618]&~m[1619]&~m[1620]&~m[1622]&~m[1623])|(~m[1618]&m[1619]&~m[1620]&~m[1622]&~m[1623])|(~m[1618]&~m[1619]&m[1620]&~m[1622]&~m[1623])|(m[1618]&m[1619]&m[1620]&m[1622]&~m[1623])|(~m[1618]&~m[1619]&~m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&~m[1620]&m[1622]&m[1623])|(m[1618]&~m[1619]&m[1620]&m[1622]&m[1623])|(~m[1618]&m[1619]&m[1620]&m[1622]&m[1623]))&UnbiasedRNG[858])|((m[1618]&m[1619]&~m[1620]&~m[1622]&~m[1623])|(m[1618]&~m[1619]&m[1620]&~m[1622]&~m[1623])|(~m[1618]&m[1619]&m[1620]&~m[1622]&~m[1623])|(m[1618]&m[1619]&m[1620]&~m[1622]&~m[1623])|(m[1618]&~m[1619]&~m[1620]&~m[1622]&m[1623])|(~m[1618]&m[1619]&~m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&~m[1620]&~m[1622]&m[1623])|(~m[1618]&~m[1619]&m[1620]&~m[1622]&m[1623])|(m[1618]&~m[1619]&m[1620]&~m[1622]&m[1623])|(~m[1618]&m[1619]&m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&m[1620]&~m[1622]&m[1623])|(m[1618]&m[1619]&m[1620]&m[1622]&m[1623]))):InitCond[1753];
    m[1626] = run?((((m[1623]&~m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&~m[1628])|(~m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&m[1627]&m[1628]))&UnbiasedRNG[859])|((m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&m[1628]))):InitCond[1754];
    m[1631] = run?((((m[1628]&~m[1629]&~m[1630]&~m[1632]&~m[1633])|(~m[1628]&m[1629]&~m[1630]&~m[1632]&~m[1633])|(~m[1628]&~m[1629]&m[1630]&~m[1632]&~m[1633])|(m[1628]&m[1629]&m[1630]&m[1632]&~m[1633])|(~m[1628]&~m[1629]&~m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&~m[1630]&m[1632]&m[1633])|(m[1628]&~m[1629]&m[1630]&m[1632]&m[1633])|(~m[1628]&m[1629]&m[1630]&m[1632]&m[1633]))&UnbiasedRNG[860])|((m[1628]&m[1629]&~m[1630]&~m[1632]&~m[1633])|(m[1628]&~m[1629]&m[1630]&~m[1632]&~m[1633])|(~m[1628]&m[1629]&m[1630]&~m[1632]&~m[1633])|(m[1628]&m[1629]&m[1630]&~m[1632]&~m[1633])|(m[1628]&~m[1629]&~m[1630]&~m[1632]&m[1633])|(~m[1628]&m[1629]&~m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&~m[1630]&~m[1632]&m[1633])|(~m[1628]&~m[1629]&m[1630]&~m[1632]&m[1633])|(m[1628]&~m[1629]&m[1630]&~m[1632]&m[1633])|(~m[1628]&m[1629]&m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&m[1630]&~m[1632]&m[1633])|(m[1628]&m[1629]&m[1630]&m[1632]&m[1633]))):InitCond[1755];
    m[1636] = run?((((m[1633]&~m[1634]&~m[1635]&~m[1637]&~m[1638])|(~m[1633]&m[1634]&~m[1635]&~m[1637]&~m[1638])|(~m[1633]&~m[1634]&m[1635]&~m[1637]&~m[1638])|(m[1633]&m[1634]&m[1635]&m[1637]&~m[1638])|(~m[1633]&~m[1634]&~m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&~m[1635]&m[1637]&m[1638])|(m[1633]&~m[1634]&m[1635]&m[1637]&m[1638])|(~m[1633]&m[1634]&m[1635]&m[1637]&m[1638]))&UnbiasedRNG[861])|((m[1633]&m[1634]&~m[1635]&~m[1637]&~m[1638])|(m[1633]&~m[1634]&m[1635]&~m[1637]&~m[1638])|(~m[1633]&m[1634]&m[1635]&~m[1637]&~m[1638])|(m[1633]&m[1634]&m[1635]&~m[1637]&~m[1638])|(m[1633]&~m[1634]&~m[1635]&~m[1637]&m[1638])|(~m[1633]&m[1634]&~m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&~m[1635]&~m[1637]&m[1638])|(~m[1633]&~m[1634]&m[1635]&~m[1637]&m[1638])|(m[1633]&~m[1634]&m[1635]&~m[1637]&m[1638])|(~m[1633]&m[1634]&m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&m[1635]&~m[1637]&m[1638])|(m[1633]&m[1634]&m[1635]&m[1637]&m[1638]))):InitCond[1756];
    m[1641] = run?((((m[1638]&~m[1639]&~m[1640]&~m[1642]&~m[1643])|(~m[1638]&m[1639]&~m[1640]&~m[1642]&~m[1643])|(~m[1638]&~m[1639]&m[1640]&~m[1642]&~m[1643])|(m[1638]&m[1639]&m[1640]&m[1642]&~m[1643])|(~m[1638]&~m[1639]&~m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&~m[1640]&m[1642]&m[1643])|(m[1638]&~m[1639]&m[1640]&m[1642]&m[1643])|(~m[1638]&m[1639]&m[1640]&m[1642]&m[1643]))&UnbiasedRNG[862])|((m[1638]&m[1639]&~m[1640]&~m[1642]&~m[1643])|(m[1638]&~m[1639]&m[1640]&~m[1642]&~m[1643])|(~m[1638]&m[1639]&m[1640]&~m[1642]&~m[1643])|(m[1638]&m[1639]&m[1640]&~m[1642]&~m[1643])|(m[1638]&~m[1639]&~m[1640]&~m[1642]&m[1643])|(~m[1638]&m[1639]&~m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&~m[1640]&~m[1642]&m[1643])|(~m[1638]&~m[1639]&m[1640]&~m[1642]&m[1643])|(m[1638]&~m[1639]&m[1640]&~m[1642]&m[1643])|(~m[1638]&m[1639]&m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&m[1640]&~m[1642]&m[1643])|(m[1638]&m[1639]&m[1640]&m[1642]&m[1643]))):InitCond[1757];
    m[1646] = run?((((m[1643]&~m[1644]&~m[1645]&~m[1647]&~m[1648])|(~m[1643]&m[1644]&~m[1645]&~m[1647]&~m[1648])|(~m[1643]&~m[1644]&m[1645]&~m[1647]&~m[1648])|(m[1643]&m[1644]&m[1645]&m[1647]&~m[1648])|(~m[1643]&~m[1644]&~m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&~m[1645]&m[1647]&m[1648])|(m[1643]&~m[1644]&m[1645]&m[1647]&m[1648])|(~m[1643]&m[1644]&m[1645]&m[1647]&m[1648]))&UnbiasedRNG[863])|((m[1643]&m[1644]&~m[1645]&~m[1647]&~m[1648])|(m[1643]&~m[1644]&m[1645]&~m[1647]&~m[1648])|(~m[1643]&m[1644]&m[1645]&~m[1647]&~m[1648])|(m[1643]&m[1644]&m[1645]&~m[1647]&~m[1648])|(m[1643]&~m[1644]&~m[1645]&~m[1647]&m[1648])|(~m[1643]&m[1644]&~m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&~m[1645]&~m[1647]&m[1648])|(~m[1643]&~m[1644]&m[1645]&~m[1647]&m[1648])|(m[1643]&~m[1644]&m[1645]&~m[1647]&m[1648])|(~m[1643]&m[1644]&m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&m[1645]&~m[1647]&m[1648])|(m[1643]&m[1644]&m[1645]&m[1647]&m[1648]))):InitCond[1758];
    m[1651] = run?((((m[1648]&~m[1649]&~m[1650]&~m[1652]&~m[1653])|(~m[1648]&m[1649]&~m[1650]&~m[1652]&~m[1653])|(~m[1648]&~m[1649]&m[1650]&~m[1652]&~m[1653])|(m[1648]&m[1649]&m[1650]&m[1652]&~m[1653])|(~m[1648]&~m[1649]&~m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&~m[1650]&m[1652]&m[1653])|(m[1648]&~m[1649]&m[1650]&m[1652]&m[1653])|(~m[1648]&m[1649]&m[1650]&m[1652]&m[1653]))&UnbiasedRNG[864])|((m[1648]&m[1649]&~m[1650]&~m[1652]&~m[1653])|(m[1648]&~m[1649]&m[1650]&~m[1652]&~m[1653])|(~m[1648]&m[1649]&m[1650]&~m[1652]&~m[1653])|(m[1648]&m[1649]&m[1650]&~m[1652]&~m[1653])|(m[1648]&~m[1649]&~m[1650]&~m[1652]&m[1653])|(~m[1648]&m[1649]&~m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&~m[1650]&~m[1652]&m[1653])|(~m[1648]&~m[1649]&m[1650]&~m[1652]&m[1653])|(m[1648]&~m[1649]&m[1650]&~m[1652]&m[1653])|(~m[1648]&m[1649]&m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&m[1650]&~m[1652]&m[1653])|(m[1648]&m[1649]&m[1650]&m[1652]&m[1653]))):InitCond[1759];
    m[1656] = run?((((m[1653]&~m[1654]&~m[1655]&~m[1657]&~m[1658])|(~m[1653]&m[1654]&~m[1655]&~m[1657]&~m[1658])|(~m[1653]&~m[1654]&m[1655]&~m[1657]&~m[1658])|(m[1653]&m[1654]&m[1655]&m[1657]&~m[1658])|(~m[1653]&~m[1654]&~m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&~m[1655]&m[1657]&m[1658])|(m[1653]&~m[1654]&m[1655]&m[1657]&m[1658])|(~m[1653]&m[1654]&m[1655]&m[1657]&m[1658]))&UnbiasedRNG[865])|((m[1653]&m[1654]&~m[1655]&~m[1657]&~m[1658])|(m[1653]&~m[1654]&m[1655]&~m[1657]&~m[1658])|(~m[1653]&m[1654]&m[1655]&~m[1657]&~m[1658])|(m[1653]&m[1654]&m[1655]&~m[1657]&~m[1658])|(m[1653]&~m[1654]&~m[1655]&~m[1657]&m[1658])|(~m[1653]&m[1654]&~m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&~m[1655]&~m[1657]&m[1658])|(~m[1653]&~m[1654]&m[1655]&~m[1657]&m[1658])|(m[1653]&~m[1654]&m[1655]&~m[1657]&m[1658])|(~m[1653]&m[1654]&m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&m[1655]&~m[1657]&m[1658])|(m[1653]&m[1654]&m[1655]&m[1657]&m[1658]))):InitCond[1760];
    m[1661] = run?((((m[1658]&~m[1659]&~m[1660]&~m[1662]&~m[1663])|(~m[1658]&m[1659]&~m[1660]&~m[1662]&~m[1663])|(~m[1658]&~m[1659]&m[1660]&~m[1662]&~m[1663])|(m[1658]&m[1659]&m[1660]&m[1662]&~m[1663])|(~m[1658]&~m[1659]&~m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&~m[1660]&m[1662]&m[1663])|(m[1658]&~m[1659]&m[1660]&m[1662]&m[1663])|(~m[1658]&m[1659]&m[1660]&m[1662]&m[1663]))&UnbiasedRNG[866])|((m[1658]&m[1659]&~m[1660]&~m[1662]&~m[1663])|(m[1658]&~m[1659]&m[1660]&~m[1662]&~m[1663])|(~m[1658]&m[1659]&m[1660]&~m[1662]&~m[1663])|(m[1658]&m[1659]&m[1660]&~m[1662]&~m[1663])|(m[1658]&~m[1659]&~m[1660]&~m[1662]&m[1663])|(~m[1658]&m[1659]&~m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&~m[1660]&~m[1662]&m[1663])|(~m[1658]&~m[1659]&m[1660]&~m[1662]&m[1663])|(m[1658]&~m[1659]&m[1660]&~m[1662]&m[1663])|(~m[1658]&m[1659]&m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&m[1660]&~m[1662]&m[1663])|(m[1658]&m[1659]&m[1660]&m[1662]&m[1663]))):InitCond[1761];
    m[1666] = run?((((m[1663]&~m[1664]&~m[1665]&~m[1667]&~m[1668])|(~m[1663]&m[1664]&~m[1665]&~m[1667]&~m[1668])|(~m[1663]&~m[1664]&m[1665]&~m[1667]&~m[1668])|(m[1663]&m[1664]&m[1665]&m[1667]&~m[1668])|(~m[1663]&~m[1664]&~m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&~m[1665]&m[1667]&m[1668])|(m[1663]&~m[1664]&m[1665]&m[1667]&m[1668])|(~m[1663]&m[1664]&m[1665]&m[1667]&m[1668]))&UnbiasedRNG[867])|((m[1663]&m[1664]&~m[1665]&~m[1667]&~m[1668])|(m[1663]&~m[1664]&m[1665]&~m[1667]&~m[1668])|(~m[1663]&m[1664]&m[1665]&~m[1667]&~m[1668])|(m[1663]&m[1664]&m[1665]&~m[1667]&~m[1668])|(m[1663]&~m[1664]&~m[1665]&~m[1667]&m[1668])|(~m[1663]&m[1664]&~m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&~m[1665]&~m[1667]&m[1668])|(~m[1663]&~m[1664]&m[1665]&~m[1667]&m[1668])|(m[1663]&~m[1664]&m[1665]&~m[1667]&m[1668])|(~m[1663]&m[1664]&m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&m[1665]&~m[1667]&m[1668])|(m[1663]&m[1664]&m[1665]&m[1667]&m[1668]))):InitCond[1762];
    m[1676] = run?((((m[1673]&~m[1674]&~m[1675]&~m[1677]&~m[1678])|(~m[1673]&m[1674]&~m[1675]&~m[1677]&~m[1678])|(~m[1673]&~m[1674]&m[1675]&~m[1677]&~m[1678])|(m[1673]&m[1674]&m[1675]&m[1677]&~m[1678])|(~m[1673]&~m[1674]&~m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&~m[1675]&m[1677]&m[1678])|(m[1673]&~m[1674]&m[1675]&m[1677]&m[1678])|(~m[1673]&m[1674]&m[1675]&m[1677]&m[1678]))&UnbiasedRNG[868])|((m[1673]&m[1674]&~m[1675]&~m[1677]&~m[1678])|(m[1673]&~m[1674]&m[1675]&~m[1677]&~m[1678])|(~m[1673]&m[1674]&m[1675]&~m[1677]&~m[1678])|(m[1673]&m[1674]&m[1675]&~m[1677]&~m[1678])|(m[1673]&~m[1674]&~m[1675]&~m[1677]&m[1678])|(~m[1673]&m[1674]&~m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&~m[1675]&~m[1677]&m[1678])|(~m[1673]&~m[1674]&m[1675]&~m[1677]&m[1678])|(m[1673]&~m[1674]&m[1675]&~m[1677]&m[1678])|(~m[1673]&m[1674]&m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&m[1675]&~m[1677]&m[1678])|(m[1673]&m[1674]&m[1675]&m[1677]&m[1678]))):InitCond[1763];
    m[1681] = run?((((m[1678]&~m[1679]&~m[1680]&~m[1682]&~m[1683])|(~m[1678]&m[1679]&~m[1680]&~m[1682]&~m[1683])|(~m[1678]&~m[1679]&m[1680]&~m[1682]&~m[1683])|(m[1678]&m[1679]&m[1680]&m[1682]&~m[1683])|(~m[1678]&~m[1679]&~m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&~m[1680]&m[1682]&m[1683])|(m[1678]&~m[1679]&m[1680]&m[1682]&m[1683])|(~m[1678]&m[1679]&m[1680]&m[1682]&m[1683]))&UnbiasedRNG[869])|((m[1678]&m[1679]&~m[1680]&~m[1682]&~m[1683])|(m[1678]&~m[1679]&m[1680]&~m[1682]&~m[1683])|(~m[1678]&m[1679]&m[1680]&~m[1682]&~m[1683])|(m[1678]&m[1679]&m[1680]&~m[1682]&~m[1683])|(m[1678]&~m[1679]&~m[1680]&~m[1682]&m[1683])|(~m[1678]&m[1679]&~m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&~m[1680]&~m[1682]&m[1683])|(~m[1678]&~m[1679]&m[1680]&~m[1682]&m[1683])|(m[1678]&~m[1679]&m[1680]&~m[1682]&m[1683])|(~m[1678]&m[1679]&m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&m[1680]&~m[1682]&m[1683])|(m[1678]&m[1679]&m[1680]&m[1682]&m[1683]))):InitCond[1764];
    m[1686] = run?((((m[1683]&~m[1684]&~m[1685]&~m[1687]&~m[1688])|(~m[1683]&m[1684]&~m[1685]&~m[1687]&~m[1688])|(~m[1683]&~m[1684]&m[1685]&~m[1687]&~m[1688])|(m[1683]&m[1684]&m[1685]&m[1687]&~m[1688])|(~m[1683]&~m[1684]&~m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&~m[1685]&m[1687]&m[1688])|(m[1683]&~m[1684]&m[1685]&m[1687]&m[1688])|(~m[1683]&m[1684]&m[1685]&m[1687]&m[1688]))&UnbiasedRNG[870])|((m[1683]&m[1684]&~m[1685]&~m[1687]&~m[1688])|(m[1683]&~m[1684]&m[1685]&~m[1687]&~m[1688])|(~m[1683]&m[1684]&m[1685]&~m[1687]&~m[1688])|(m[1683]&m[1684]&m[1685]&~m[1687]&~m[1688])|(m[1683]&~m[1684]&~m[1685]&~m[1687]&m[1688])|(~m[1683]&m[1684]&~m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&~m[1685]&~m[1687]&m[1688])|(~m[1683]&~m[1684]&m[1685]&~m[1687]&m[1688])|(m[1683]&~m[1684]&m[1685]&~m[1687]&m[1688])|(~m[1683]&m[1684]&m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&m[1685]&~m[1687]&m[1688])|(m[1683]&m[1684]&m[1685]&m[1687]&m[1688]))):InitCond[1765];
    m[1691] = run?((((m[1688]&~m[1689]&~m[1690]&~m[1692]&~m[1693])|(~m[1688]&m[1689]&~m[1690]&~m[1692]&~m[1693])|(~m[1688]&~m[1689]&m[1690]&~m[1692]&~m[1693])|(m[1688]&m[1689]&m[1690]&m[1692]&~m[1693])|(~m[1688]&~m[1689]&~m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&~m[1690]&m[1692]&m[1693])|(m[1688]&~m[1689]&m[1690]&m[1692]&m[1693])|(~m[1688]&m[1689]&m[1690]&m[1692]&m[1693]))&UnbiasedRNG[871])|((m[1688]&m[1689]&~m[1690]&~m[1692]&~m[1693])|(m[1688]&~m[1689]&m[1690]&~m[1692]&~m[1693])|(~m[1688]&m[1689]&m[1690]&~m[1692]&~m[1693])|(m[1688]&m[1689]&m[1690]&~m[1692]&~m[1693])|(m[1688]&~m[1689]&~m[1690]&~m[1692]&m[1693])|(~m[1688]&m[1689]&~m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&~m[1690]&~m[1692]&m[1693])|(~m[1688]&~m[1689]&m[1690]&~m[1692]&m[1693])|(m[1688]&~m[1689]&m[1690]&~m[1692]&m[1693])|(~m[1688]&m[1689]&m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&m[1690]&~m[1692]&m[1693])|(m[1688]&m[1689]&m[1690]&m[1692]&m[1693]))):InitCond[1766];
    m[1696] = run?((((m[1693]&~m[1694]&~m[1695]&~m[1697]&~m[1698])|(~m[1693]&m[1694]&~m[1695]&~m[1697]&~m[1698])|(~m[1693]&~m[1694]&m[1695]&~m[1697]&~m[1698])|(m[1693]&m[1694]&m[1695]&m[1697]&~m[1698])|(~m[1693]&~m[1694]&~m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&~m[1695]&m[1697]&m[1698])|(m[1693]&~m[1694]&m[1695]&m[1697]&m[1698])|(~m[1693]&m[1694]&m[1695]&m[1697]&m[1698]))&UnbiasedRNG[872])|((m[1693]&m[1694]&~m[1695]&~m[1697]&~m[1698])|(m[1693]&~m[1694]&m[1695]&~m[1697]&~m[1698])|(~m[1693]&m[1694]&m[1695]&~m[1697]&~m[1698])|(m[1693]&m[1694]&m[1695]&~m[1697]&~m[1698])|(m[1693]&~m[1694]&~m[1695]&~m[1697]&m[1698])|(~m[1693]&m[1694]&~m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&~m[1695]&~m[1697]&m[1698])|(~m[1693]&~m[1694]&m[1695]&~m[1697]&m[1698])|(m[1693]&~m[1694]&m[1695]&~m[1697]&m[1698])|(~m[1693]&m[1694]&m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&m[1695]&~m[1697]&m[1698])|(m[1693]&m[1694]&m[1695]&m[1697]&m[1698]))):InitCond[1767];
    m[1701] = run?((((m[1698]&~m[1699]&~m[1700]&~m[1702]&~m[1703])|(~m[1698]&m[1699]&~m[1700]&~m[1702]&~m[1703])|(~m[1698]&~m[1699]&m[1700]&~m[1702]&~m[1703])|(m[1698]&m[1699]&m[1700]&m[1702]&~m[1703])|(~m[1698]&~m[1699]&~m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&~m[1700]&m[1702]&m[1703])|(m[1698]&~m[1699]&m[1700]&m[1702]&m[1703])|(~m[1698]&m[1699]&m[1700]&m[1702]&m[1703]))&UnbiasedRNG[873])|((m[1698]&m[1699]&~m[1700]&~m[1702]&~m[1703])|(m[1698]&~m[1699]&m[1700]&~m[1702]&~m[1703])|(~m[1698]&m[1699]&m[1700]&~m[1702]&~m[1703])|(m[1698]&m[1699]&m[1700]&~m[1702]&~m[1703])|(m[1698]&~m[1699]&~m[1700]&~m[1702]&m[1703])|(~m[1698]&m[1699]&~m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&~m[1700]&~m[1702]&m[1703])|(~m[1698]&~m[1699]&m[1700]&~m[1702]&m[1703])|(m[1698]&~m[1699]&m[1700]&~m[1702]&m[1703])|(~m[1698]&m[1699]&m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&m[1700]&~m[1702]&m[1703])|(m[1698]&m[1699]&m[1700]&m[1702]&m[1703]))):InitCond[1768];
    m[1706] = run?((((m[1703]&~m[1704]&~m[1705]&~m[1707]&~m[1708])|(~m[1703]&m[1704]&~m[1705]&~m[1707]&~m[1708])|(~m[1703]&~m[1704]&m[1705]&~m[1707]&~m[1708])|(m[1703]&m[1704]&m[1705]&m[1707]&~m[1708])|(~m[1703]&~m[1704]&~m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&~m[1705]&m[1707]&m[1708])|(m[1703]&~m[1704]&m[1705]&m[1707]&m[1708])|(~m[1703]&m[1704]&m[1705]&m[1707]&m[1708]))&UnbiasedRNG[874])|((m[1703]&m[1704]&~m[1705]&~m[1707]&~m[1708])|(m[1703]&~m[1704]&m[1705]&~m[1707]&~m[1708])|(~m[1703]&m[1704]&m[1705]&~m[1707]&~m[1708])|(m[1703]&m[1704]&m[1705]&~m[1707]&~m[1708])|(m[1703]&~m[1704]&~m[1705]&~m[1707]&m[1708])|(~m[1703]&m[1704]&~m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&~m[1705]&~m[1707]&m[1708])|(~m[1703]&~m[1704]&m[1705]&~m[1707]&m[1708])|(m[1703]&~m[1704]&m[1705]&~m[1707]&m[1708])|(~m[1703]&m[1704]&m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&m[1705]&~m[1707]&m[1708])|(m[1703]&m[1704]&m[1705]&m[1707]&m[1708]))):InitCond[1769];
    m[1711] = run?((((m[1708]&~m[1709]&~m[1710]&~m[1712]&~m[1713])|(~m[1708]&m[1709]&~m[1710]&~m[1712]&~m[1713])|(~m[1708]&~m[1709]&m[1710]&~m[1712]&~m[1713])|(m[1708]&m[1709]&m[1710]&m[1712]&~m[1713])|(~m[1708]&~m[1709]&~m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&~m[1710]&m[1712]&m[1713])|(m[1708]&~m[1709]&m[1710]&m[1712]&m[1713])|(~m[1708]&m[1709]&m[1710]&m[1712]&m[1713]))&UnbiasedRNG[875])|((m[1708]&m[1709]&~m[1710]&~m[1712]&~m[1713])|(m[1708]&~m[1709]&m[1710]&~m[1712]&~m[1713])|(~m[1708]&m[1709]&m[1710]&~m[1712]&~m[1713])|(m[1708]&m[1709]&m[1710]&~m[1712]&~m[1713])|(m[1708]&~m[1709]&~m[1710]&~m[1712]&m[1713])|(~m[1708]&m[1709]&~m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&~m[1710]&~m[1712]&m[1713])|(~m[1708]&~m[1709]&m[1710]&~m[1712]&m[1713])|(m[1708]&~m[1709]&m[1710]&~m[1712]&m[1713])|(~m[1708]&m[1709]&m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&m[1710]&~m[1712]&m[1713])|(m[1708]&m[1709]&m[1710]&m[1712]&m[1713]))):InitCond[1770];
    m[1716] = run?((((m[1713]&~m[1714]&~m[1715]&~m[1717]&~m[1718])|(~m[1713]&m[1714]&~m[1715]&~m[1717]&~m[1718])|(~m[1713]&~m[1714]&m[1715]&~m[1717]&~m[1718])|(m[1713]&m[1714]&m[1715]&m[1717]&~m[1718])|(~m[1713]&~m[1714]&~m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&~m[1715]&m[1717]&m[1718])|(m[1713]&~m[1714]&m[1715]&m[1717]&m[1718])|(~m[1713]&m[1714]&m[1715]&m[1717]&m[1718]))&UnbiasedRNG[876])|((m[1713]&m[1714]&~m[1715]&~m[1717]&~m[1718])|(m[1713]&~m[1714]&m[1715]&~m[1717]&~m[1718])|(~m[1713]&m[1714]&m[1715]&~m[1717]&~m[1718])|(m[1713]&m[1714]&m[1715]&~m[1717]&~m[1718])|(m[1713]&~m[1714]&~m[1715]&~m[1717]&m[1718])|(~m[1713]&m[1714]&~m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&~m[1715]&~m[1717]&m[1718])|(~m[1713]&~m[1714]&m[1715]&~m[1717]&m[1718])|(m[1713]&~m[1714]&m[1715]&~m[1717]&m[1718])|(~m[1713]&m[1714]&m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&m[1715]&~m[1717]&m[1718])|(m[1713]&m[1714]&m[1715]&m[1717]&m[1718]))):InitCond[1771];
    m[1721] = run?((((m[1718]&~m[1719]&~m[1720]&~m[1722]&~m[1723])|(~m[1718]&m[1719]&~m[1720]&~m[1722]&~m[1723])|(~m[1718]&~m[1719]&m[1720]&~m[1722]&~m[1723])|(m[1718]&m[1719]&m[1720]&m[1722]&~m[1723])|(~m[1718]&~m[1719]&~m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&~m[1720]&m[1722]&m[1723])|(m[1718]&~m[1719]&m[1720]&m[1722]&m[1723])|(~m[1718]&m[1719]&m[1720]&m[1722]&m[1723]))&UnbiasedRNG[877])|((m[1718]&m[1719]&~m[1720]&~m[1722]&~m[1723])|(m[1718]&~m[1719]&m[1720]&~m[1722]&~m[1723])|(~m[1718]&m[1719]&m[1720]&~m[1722]&~m[1723])|(m[1718]&m[1719]&m[1720]&~m[1722]&~m[1723])|(m[1718]&~m[1719]&~m[1720]&~m[1722]&m[1723])|(~m[1718]&m[1719]&~m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&~m[1720]&~m[1722]&m[1723])|(~m[1718]&~m[1719]&m[1720]&~m[1722]&m[1723])|(m[1718]&~m[1719]&m[1720]&~m[1722]&m[1723])|(~m[1718]&m[1719]&m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&m[1720]&~m[1722]&m[1723])|(m[1718]&m[1719]&m[1720]&m[1722]&m[1723]))):InitCond[1772];
    m[1726] = run?((((m[1723]&~m[1724]&~m[1725]&~m[1727]&~m[1728])|(~m[1723]&m[1724]&~m[1725]&~m[1727]&~m[1728])|(~m[1723]&~m[1724]&m[1725]&~m[1727]&~m[1728])|(m[1723]&m[1724]&m[1725]&m[1727]&~m[1728])|(~m[1723]&~m[1724]&~m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&~m[1725]&m[1727]&m[1728])|(m[1723]&~m[1724]&m[1725]&m[1727]&m[1728])|(~m[1723]&m[1724]&m[1725]&m[1727]&m[1728]))&UnbiasedRNG[878])|((m[1723]&m[1724]&~m[1725]&~m[1727]&~m[1728])|(m[1723]&~m[1724]&m[1725]&~m[1727]&~m[1728])|(~m[1723]&m[1724]&m[1725]&~m[1727]&~m[1728])|(m[1723]&m[1724]&m[1725]&~m[1727]&~m[1728])|(m[1723]&~m[1724]&~m[1725]&~m[1727]&m[1728])|(~m[1723]&m[1724]&~m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&~m[1725]&~m[1727]&m[1728])|(~m[1723]&~m[1724]&m[1725]&~m[1727]&m[1728])|(m[1723]&~m[1724]&m[1725]&~m[1727]&m[1728])|(~m[1723]&m[1724]&m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&m[1725]&~m[1727]&m[1728])|(m[1723]&m[1724]&m[1725]&m[1727]&m[1728]))):InitCond[1773];
    m[1731] = run?((((m[1728]&~m[1729]&~m[1730]&~m[1732]&~m[1733])|(~m[1728]&m[1729]&~m[1730]&~m[1732]&~m[1733])|(~m[1728]&~m[1729]&m[1730]&~m[1732]&~m[1733])|(m[1728]&m[1729]&m[1730]&m[1732]&~m[1733])|(~m[1728]&~m[1729]&~m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&~m[1730]&m[1732]&m[1733])|(m[1728]&~m[1729]&m[1730]&m[1732]&m[1733])|(~m[1728]&m[1729]&m[1730]&m[1732]&m[1733]))&UnbiasedRNG[879])|((m[1728]&m[1729]&~m[1730]&~m[1732]&~m[1733])|(m[1728]&~m[1729]&m[1730]&~m[1732]&~m[1733])|(~m[1728]&m[1729]&m[1730]&~m[1732]&~m[1733])|(m[1728]&m[1729]&m[1730]&~m[1732]&~m[1733])|(m[1728]&~m[1729]&~m[1730]&~m[1732]&m[1733])|(~m[1728]&m[1729]&~m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&~m[1730]&~m[1732]&m[1733])|(~m[1728]&~m[1729]&m[1730]&~m[1732]&m[1733])|(m[1728]&~m[1729]&m[1730]&~m[1732]&m[1733])|(~m[1728]&m[1729]&m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&m[1730]&~m[1732]&m[1733])|(m[1728]&m[1729]&m[1730]&m[1732]&m[1733]))):InitCond[1774];
    m[1741] = run?((((m[1738]&~m[1739]&~m[1740]&~m[1742]&~m[1743])|(~m[1738]&m[1739]&~m[1740]&~m[1742]&~m[1743])|(~m[1738]&~m[1739]&m[1740]&~m[1742]&~m[1743])|(m[1738]&m[1739]&m[1740]&m[1742]&~m[1743])|(~m[1738]&~m[1739]&~m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&~m[1740]&m[1742]&m[1743])|(m[1738]&~m[1739]&m[1740]&m[1742]&m[1743])|(~m[1738]&m[1739]&m[1740]&m[1742]&m[1743]))&UnbiasedRNG[880])|((m[1738]&m[1739]&~m[1740]&~m[1742]&~m[1743])|(m[1738]&~m[1739]&m[1740]&~m[1742]&~m[1743])|(~m[1738]&m[1739]&m[1740]&~m[1742]&~m[1743])|(m[1738]&m[1739]&m[1740]&~m[1742]&~m[1743])|(m[1738]&~m[1739]&~m[1740]&~m[1742]&m[1743])|(~m[1738]&m[1739]&~m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&~m[1740]&~m[1742]&m[1743])|(~m[1738]&~m[1739]&m[1740]&~m[1742]&m[1743])|(m[1738]&~m[1739]&m[1740]&~m[1742]&m[1743])|(~m[1738]&m[1739]&m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&m[1740]&~m[1742]&m[1743])|(m[1738]&m[1739]&m[1740]&m[1742]&m[1743]))):InitCond[1775];
    m[1746] = run?((((m[1743]&~m[1744]&~m[1745]&~m[1747]&~m[1748])|(~m[1743]&m[1744]&~m[1745]&~m[1747]&~m[1748])|(~m[1743]&~m[1744]&m[1745]&~m[1747]&~m[1748])|(m[1743]&m[1744]&m[1745]&m[1747]&~m[1748])|(~m[1743]&~m[1744]&~m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&~m[1745]&m[1747]&m[1748])|(m[1743]&~m[1744]&m[1745]&m[1747]&m[1748])|(~m[1743]&m[1744]&m[1745]&m[1747]&m[1748]))&UnbiasedRNG[881])|((m[1743]&m[1744]&~m[1745]&~m[1747]&~m[1748])|(m[1743]&~m[1744]&m[1745]&~m[1747]&~m[1748])|(~m[1743]&m[1744]&m[1745]&~m[1747]&~m[1748])|(m[1743]&m[1744]&m[1745]&~m[1747]&~m[1748])|(m[1743]&~m[1744]&~m[1745]&~m[1747]&m[1748])|(~m[1743]&m[1744]&~m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&~m[1745]&~m[1747]&m[1748])|(~m[1743]&~m[1744]&m[1745]&~m[1747]&m[1748])|(m[1743]&~m[1744]&m[1745]&~m[1747]&m[1748])|(~m[1743]&m[1744]&m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&m[1745]&~m[1747]&m[1748])|(m[1743]&m[1744]&m[1745]&m[1747]&m[1748]))):InitCond[1776];
    m[1751] = run?((((m[1748]&~m[1749]&~m[1750]&~m[1752]&~m[1753])|(~m[1748]&m[1749]&~m[1750]&~m[1752]&~m[1753])|(~m[1748]&~m[1749]&m[1750]&~m[1752]&~m[1753])|(m[1748]&m[1749]&m[1750]&m[1752]&~m[1753])|(~m[1748]&~m[1749]&~m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&~m[1750]&m[1752]&m[1753])|(m[1748]&~m[1749]&m[1750]&m[1752]&m[1753])|(~m[1748]&m[1749]&m[1750]&m[1752]&m[1753]))&UnbiasedRNG[882])|((m[1748]&m[1749]&~m[1750]&~m[1752]&~m[1753])|(m[1748]&~m[1749]&m[1750]&~m[1752]&~m[1753])|(~m[1748]&m[1749]&m[1750]&~m[1752]&~m[1753])|(m[1748]&m[1749]&m[1750]&~m[1752]&~m[1753])|(m[1748]&~m[1749]&~m[1750]&~m[1752]&m[1753])|(~m[1748]&m[1749]&~m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&~m[1750]&~m[1752]&m[1753])|(~m[1748]&~m[1749]&m[1750]&~m[1752]&m[1753])|(m[1748]&~m[1749]&m[1750]&~m[1752]&m[1753])|(~m[1748]&m[1749]&m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&m[1750]&~m[1752]&m[1753])|(m[1748]&m[1749]&m[1750]&m[1752]&m[1753]))):InitCond[1777];
    m[1756] = run?((((m[1753]&~m[1754]&~m[1755]&~m[1757]&~m[1758])|(~m[1753]&m[1754]&~m[1755]&~m[1757]&~m[1758])|(~m[1753]&~m[1754]&m[1755]&~m[1757]&~m[1758])|(m[1753]&m[1754]&m[1755]&m[1757]&~m[1758])|(~m[1753]&~m[1754]&~m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&~m[1755]&m[1757]&m[1758])|(m[1753]&~m[1754]&m[1755]&m[1757]&m[1758])|(~m[1753]&m[1754]&m[1755]&m[1757]&m[1758]))&UnbiasedRNG[883])|((m[1753]&m[1754]&~m[1755]&~m[1757]&~m[1758])|(m[1753]&~m[1754]&m[1755]&~m[1757]&~m[1758])|(~m[1753]&m[1754]&m[1755]&~m[1757]&~m[1758])|(m[1753]&m[1754]&m[1755]&~m[1757]&~m[1758])|(m[1753]&~m[1754]&~m[1755]&~m[1757]&m[1758])|(~m[1753]&m[1754]&~m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&~m[1755]&~m[1757]&m[1758])|(~m[1753]&~m[1754]&m[1755]&~m[1757]&m[1758])|(m[1753]&~m[1754]&m[1755]&~m[1757]&m[1758])|(~m[1753]&m[1754]&m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&m[1755]&~m[1757]&m[1758])|(m[1753]&m[1754]&m[1755]&m[1757]&m[1758]))):InitCond[1778];
    m[1761] = run?((((m[1758]&~m[1759]&~m[1760]&~m[1762]&~m[1763])|(~m[1758]&m[1759]&~m[1760]&~m[1762]&~m[1763])|(~m[1758]&~m[1759]&m[1760]&~m[1762]&~m[1763])|(m[1758]&m[1759]&m[1760]&m[1762]&~m[1763])|(~m[1758]&~m[1759]&~m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&~m[1760]&m[1762]&m[1763])|(m[1758]&~m[1759]&m[1760]&m[1762]&m[1763])|(~m[1758]&m[1759]&m[1760]&m[1762]&m[1763]))&UnbiasedRNG[884])|((m[1758]&m[1759]&~m[1760]&~m[1762]&~m[1763])|(m[1758]&~m[1759]&m[1760]&~m[1762]&~m[1763])|(~m[1758]&m[1759]&m[1760]&~m[1762]&~m[1763])|(m[1758]&m[1759]&m[1760]&~m[1762]&~m[1763])|(m[1758]&~m[1759]&~m[1760]&~m[1762]&m[1763])|(~m[1758]&m[1759]&~m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&~m[1760]&~m[1762]&m[1763])|(~m[1758]&~m[1759]&m[1760]&~m[1762]&m[1763])|(m[1758]&~m[1759]&m[1760]&~m[1762]&m[1763])|(~m[1758]&m[1759]&m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&m[1760]&~m[1762]&m[1763])|(m[1758]&m[1759]&m[1760]&m[1762]&m[1763]))):InitCond[1779];
    m[1766] = run?((((m[1763]&~m[1764]&~m[1765]&~m[1767]&~m[1768])|(~m[1763]&m[1764]&~m[1765]&~m[1767]&~m[1768])|(~m[1763]&~m[1764]&m[1765]&~m[1767]&~m[1768])|(m[1763]&m[1764]&m[1765]&m[1767]&~m[1768])|(~m[1763]&~m[1764]&~m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&~m[1765]&m[1767]&m[1768])|(m[1763]&~m[1764]&m[1765]&m[1767]&m[1768])|(~m[1763]&m[1764]&m[1765]&m[1767]&m[1768]))&UnbiasedRNG[885])|((m[1763]&m[1764]&~m[1765]&~m[1767]&~m[1768])|(m[1763]&~m[1764]&m[1765]&~m[1767]&~m[1768])|(~m[1763]&m[1764]&m[1765]&~m[1767]&~m[1768])|(m[1763]&m[1764]&m[1765]&~m[1767]&~m[1768])|(m[1763]&~m[1764]&~m[1765]&~m[1767]&m[1768])|(~m[1763]&m[1764]&~m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&~m[1765]&~m[1767]&m[1768])|(~m[1763]&~m[1764]&m[1765]&~m[1767]&m[1768])|(m[1763]&~m[1764]&m[1765]&~m[1767]&m[1768])|(~m[1763]&m[1764]&m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&m[1765]&~m[1767]&m[1768])|(m[1763]&m[1764]&m[1765]&m[1767]&m[1768]))):InitCond[1780];
    m[1771] = run?((((m[1768]&~m[1769]&~m[1770]&~m[1772]&~m[1773])|(~m[1768]&m[1769]&~m[1770]&~m[1772]&~m[1773])|(~m[1768]&~m[1769]&m[1770]&~m[1772]&~m[1773])|(m[1768]&m[1769]&m[1770]&m[1772]&~m[1773])|(~m[1768]&~m[1769]&~m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&~m[1770]&m[1772]&m[1773])|(m[1768]&~m[1769]&m[1770]&m[1772]&m[1773])|(~m[1768]&m[1769]&m[1770]&m[1772]&m[1773]))&UnbiasedRNG[886])|((m[1768]&m[1769]&~m[1770]&~m[1772]&~m[1773])|(m[1768]&~m[1769]&m[1770]&~m[1772]&~m[1773])|(~m[1768]&m[1769]&m[1770]&~m[1772]&~m[1773])|(m[1768]&m[1769]&m[1770]&~m[1772]&~m[1773])|(m[1768]&~m[1769]&~m[1770]&~m[1772]&m[1773])|(~m[1768]&m[1769]&~m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&~m[1770]&~m[1772]&m[1773])|(~m[1768]&~m[1769]&m[1770]&~m[1772]&m[1773])|(m[1768]&~m[1769]&m[1770]&~m[1772]&m[1773])|(~m[1768]&m[1769]&m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&m[1770]&~m[1772]&m[1773])|(m[1768]&m[1769]&m[1770]&m[1772]&m[1773]))):InitCond[1781];
    m[1776] = run?((((m[1773]&~m[1774]&~m[1775]&~m[1777]&~m[1778])|(~m[1773]&m[1774]&~m[1775]&~m[1777]&~m[1778])|(~m[1773]&~m[1774]&m[1775]&~m[1777]&~m[1778])|(m[1773]&m[1774]&m[1775]&m[1777]&~m[1778])|(~m[1773]&~m[1774]&~m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&~m[1775]&m[1777]&m[1778])|(m[1773]&~m[1774]&m[1775]&m[1777]&m[1778])|(~m[1773]&m[1774]&m[1775]&m[1777]&m[1778]))&UnbiasedRNG[887])|((m[1773]&m[1774]&~m[1775]&~m[1777]&~m[1778])|(m[1773]&~m[1774]&m[1775]&~m[1777]&~m[1778])|(~m[1773]&m[1774]&m[1775]&~m[1777]&~m[1778])|(m[1773]&m[1774]&m[1775]&~m[1777]&~m[1778])|(m[1773]&~m[1774]&~m[1775]&~m[1777]&m[1778])|(~m[1773]&m[1774]&~m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&~m[1775]&~m[1777]&m[1778])|(~m[1773]&~m[1774]&m[1775]&~m[1777]&m[1778])|(m[1773]&~m[1774]&m[1775]&~m[1777]&m[1778])|(~m[1773]&m[1774]&m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&m[1775]&~m[1777]&m[1778])|(m[1773]&m[1774]&m[1775]&m[1777]&m[1778]))):InitCond[1782];
    m[1781] = run?((((m[1778]&~m[1779]&~m[1780]&~m[1782]&~m[1783])|(~m[1778]&m[1779]&~m[1780]&~m[1782]&~m[1783])|(~m[1778]&~m[1779]&m[1780]&~m[1782]&~m[1783])|(m[1778]&m[1779]&m[1780]&m[1782]&~m[1783])|(~m[1778]&~m[1779]&~m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&~m[1780]&m[1782]&m[1783])|(m[1778]&~m[1779]&m[1780]&m[1782]&m[1783])|(~m[1778]&m[1779]&m[1780]&m[1782]&m[1783]))&UnbiasedRNG[888])|((m[1778]&m[1779]&~m[1780]&~m[1782]&~m[1783])|(m[1778]&~m[1779]&m[1780]&~m[1782]&~m[1783])|(~m[1778]&m[1779]&m[1780]&~m[1782]&~m[1783])|(m[1778]&m[1779]&m[1780]&~m[1782]&~m[1783])|(m[1778]&~m[1779]&~m[1780]&~m[1782]&m[1783])|(~m[1778]&m[1779]&~m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&~m[1780]&~m[1782]&m[1783])|(~m[1778]&~m[1779]&m[1780]&~m[1782]&m[1783])|(m[1778]&~m[1779]&m[1780]&~m[1782]&m[1783])|(~m[1778]&m[1779]&m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&m[1780]&~m[1782]&m[1783])|(m[1778]&m[1779]&m[1780]&m[1782]&m[1783]))):InitCond[1783];
    m[1786] = run?((((m[1783]&~m[1784]&~m[1785]&~m[1787]&~m[1788])|(~m[1783]&m[1784]&~m[1785]&~m[1787]&~m[1788])|(~m[1783]&~m[1784]&m[1785]&~m[1787]&~m[1788])|(m[1783]&m[1784]&m[1785]&m[1787]&~m[1788])|(~m[1783]&~m[1784]&~m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&~m[1785]&m[1787]&m[1788])|(m[1783]&~m[1784]&m[1785]&m[1787]&m[1788])|(~m[1783]&m[1784]&m[1785]&m[1787]&m[1788]))&UnbiasedRNG[889])|((m[1783]&m[1784]&~m[1785]&~m[1787]&~m[1788])|(m[1783]&~m[1784]&m[1785]&~m[1787]&~m[1788])|(~m[1783]&m[1784]&m[1785]&~m[1787]&~m[1788])|(m[1783]&m[1784]&m[1785]&~m[1787]&~m[1788])|(m[1783]&~m[1784]&~m[1785]&~m[1787]&m[1788])|(~m[1783]&m[1784]&~m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&~m[1785]&~m[1787]&m[1788])|(~m[1783]&~m[1784]&m[1785]&~m[1787]&m[1788])|(m[1783]&~m[1784]&m[1785]&~m[1787]&m[1788])|(~m[1783]&m[1784]&m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&m[1785]&~m[1787]&m[1788])|(m[1783]&m[1784]&m[1785]&m[1787]&m[1788]))):InitCond[1784];
    m[1791] = run?((((m[1788]&~m[1789]&~m[1790]&~m[1792]&~m[1793])|(~m[1788]&m[1789]&~m[1790]&~m[1792]&~m[1793])|(~m[1788]&~m[1789]&m[1790]&~m[1792]&~m[1793])|(m[1788]&m[1789]&m[1790]&m[1792]&~m[1793])|(~m[1788]&~m[1789]&~m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&~m[1790]&m[1792]&m[1793])|(m[1788]&~m[1789]&m[1790]&m[1792]&m[1793])|(~m[1788]&m[1789]&m[1790]&m[1792]&m[1793]))&UnbiasedRNG[890])|((m[1788]&m[1789]&~m[1790]&~m[1792]&~m[1793])|(m[1788]&~m[1789]&m[1790]&~m[1792]&~m[1793])|(~m[1788]&m[1789]&m[1790]&~m[1792]&~m[1793])|(m[1788]&m[1789]&m[1790]&~m[1792]&~m[1793])|(m[1788]&~m[1789]&~m[1790]&~m[1792]&m[1793])|(~m[1788]&m[1789]&~m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&~m[1790]&~m[1792]&m[1793])|(~m[1788]&~m[1789]&m[1790]&~m[1792]&m[1793])|(m[1788]&~m[1789]&m[1790]&~m[1792]&m[1793])|(~m[1788]&m[1789]&m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&m[1790]&~m[1792]&m[1793])|(m[1788]&m[1789]&m[1790]&m[1792]&m[1793]))):InitCond[1785];
    m[1801] = run?((((m[1798]&~m[1799]&~m[1800]&~m[1802]&~m[1803])|(~m[1798]&m[1799]&~m[1800]&~m[1802]&~m[1803])|(~m[1798]&~m[1799]&m[1800]&~m[1802]&~m[1803])|(m[1798]&m[1799]&m[1800]&m[1802]&~m[1803])|(~m[1798]&~m[1799]&~m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&~m[1800]&m[1802]&m[1803])|(m[1798]&~m[1799]&m[1800]&m[1802]&m[1803])|(~m[1798]&m[1799]&m[1800]&m[1802]&m[1803]))&UnbiasedRNG[891])|((m[1798]&m[1799]&~m[1800]&~m[1802]&~m[1803])|(m[1798]&~m[1799]&m[1800]&~m[1802]&~m[1803])|(~m[1798]&m[1799]&m[1800]&~m[1802]&~m[1803])|(m[1798]&m[1799]&m[1800]&~m[1802]&~m[1803])|(m[1798]&~m[1799]&~m[1800]&~m[1802]&m[1803])|(~m[1798]&m[1799]&~m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&~m[1800]&~m[1802]&m[1803])|(~m[1798]&~m[1799]&m[1800]&~m[1802]&m[1803])|(m[1798]&~m[1799]&m[1800]&~m[1802]&m[1803])|(~m[1798]&m[1799]&m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&m[1800]&~m[1802]&m[1803])|(m[1798]&m[1799]&m[1800]&m[1802]&m[1803]))):InitCond[1786];
    m[1806] = run?((((m[1803]&~m[1804]&~m[1805]&~m[1807]&~m[1808])|(~m[1803]&m[1804]&~m[1805]&~m[1807]&~m[1808])|(~m[1803]&~m[1804]&m[1805]&~m[1807]&~m[1808])|(m[1803]&m[1804]&m[1805]&m[1807]&~m[1808])|(~m[1803]&~m[1804]&~m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&~m[1805]&m[1807]&m[1808])|(m[1803]&~m[1804]&m[1805]&m[1807]&m[1808])|(~m[1803]&m[1804]&m[1805]&m[1807]&m[1808]))&UnbiasedRNG[892])|((m[1803]&m[1804]&~m[1805]&~m[1807]&~m[1808])|(m[1803]&~m[1804]&m[1805]&~m[1807]&~m[1808])|(~m[1803]&m[1804]&m[1805]&~m[1807]&~m[1808])|(m[1803]&m[1804]&m[1805]&~m[1807]&~m[1808])|(m[1803]&~m[1804]&~m[1805]&~m[1807]&m[1808])|(~m[1803]&m[1804]&~m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&~m[1805]&~m[1807]&m[1808])|(~m[1803]&~m[1804]&m[1805]&~m[1807]&m[1808])|(m[1803]&~m[1804]&m[1805]&~m[1807]&m[1808])|(~m[1803]&m[1804]&m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&m[1805]&~m[1807]&m[1808])|(m[1803]&m[1804]&m[1805]&m[1807]&m[1808]))):InitCond[1787];
    m[1811] = run?((((m[1808]&~m[1809]&~m[1810]&~m[1812]&~m[1813])|(~m[1808]&m[1809]&~m[1810]&~m[1812]&~m[1813])|(~m[1808]&~m[1809]&m[1810]&~m[1812]&~m[1813])|(m[1808]&m[1809]&m[1810]&m[1812]&~m[1813])|(~m[1808]&~m[1809]&~m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&~m[1810]&m[1812]&m[1813])|(m[1808]&~m[1809]&m[1810]&m[1812]&m[1813])|(~m[1808]&m[1809]&m[1810]&m[1812]&m[1813]))&UnbiasedRNG[893])|((m[1808]&m[1809]&~m[1810]&~m[1812]&~m[1813])|(m[1808]&~m[1809]&m[1810]&~m[1812]&~m[1813])|(~m[1808]&m[1809]&m[1810]&~m[1812]&~m[1813])|(m[1808]&m[1809]&m[1810]&~m[1812]&~m[1813])|(m[1808]&~m[1809]&~m[1810]&~m[1812]&m[1813])|(~m[1808]&m[1809]&~m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&~m[1810]&~m[1812]&m[1813])|(~m[1808]&~m[1809]&m[1810]&~m[1812]&m[1813])|(m[1808]&~m[1809]&m[1810]&~m[1812]&m[1813])|(~m[1808]&m[1809]&m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&m[1810]&~m[1812]&m[1813])|(m[1808]&m[1809]&m[1810]&m[1812]&m[1813]))):InitCond[1788];
    m[1816] = run?((((m[1813]&~m[1814]&~m[1815]&~m[1817]&~m[1818])|(~m[1813]&m[1814]&~m[1815]&~m[1817]&~m[1818])|(~m[1813]&~m[1814]&m[1815]&~m[1817]&~m[1818])|(m[1813]&m[1814]&m[1815]&m[1817]&~m[1818])|(~m[1813]&~m[1814]&~m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&~m[1815]&m[1817]&m[1818])|(m[1813]&~m[1814]&m[1815]&m[1817]&m[1818])|(~m[1813]&m[1814]&m[1815]&m[1817]&m[1818]))&UnbiasedRNG[894])|((m[1813]&m[1814]&~m[1815]&~m[1817]&~m[1818])|(m[1813]&~m[1814]&m[1815]&~m[1817]&~m[1818])|(~m[1813]&m[1814]&m[1815]&~m[1817]&~m[1818])|(m[1813]&m[1814]&m[1815]&~m[1817]&~m[1818])|(m[1813]&~m[1814]&~m[1815]&~m[1817]&m[1818])|(~m[1813]&m[1814]&~m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&~m[1815]&~m[1817]&m[1818])|(~m[1813]&~m[1814]&m[1815]&~m[1817]&m[1818])|(m[1813]&~m[1814]&m[1815]&~m[1817]&m[1818])|(~m[1813]&m[1814]&m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&m[1815]&~m[1817]&m[1818])|(m[1813]&m[1814]&m[1815]&m[1817]&m[1818]))):InitCond[1789];
    m[1821] = run?((((m[1818]&~m[1819]&~m[1820]&~m[1822]&~m[1823])|(~m[1818]&m[1819]&~m[1820]&~m[1822]&~m[1823])|(~m[1818]&~m[1819]&m[1820]&~m[1822]&~m[1823])|(m[1818]&m[1819]&m[1820]&m[1822]&~m[1823])|(~m[1818]&~m[1819]&~m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&~m[1820]&m[1822]&m[1823])|(m[1818]&~m[1819]&m[1820]&m[1822]&m[1823])|(~m[1818]&m[1819]&m[1820]&m[1822]&m[1823]))&UnbiasedRNG[895])|((m[1818]&m[1819]&~m[1820]&~m[1822]&~m[1823])|(m[1818]&~m[1819]&m[1820]&~m[1822]&~m[1823])|(~m[1818]&m[1819]&m[1820]&~m[1822]&~m[1823])|(m[1818]&m[1819]&m[1820]&~m[1822]&~m[1823])|(m[1818]&~m[1819]&~m[1820]&~m[1822]&m[1823])|(~m[1818]&m[1819]&~m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&~m[1820]&~m[1822]&m[1823])|(~m[1818]&~m[1819]&m[1820]&~m[1822]&m[1823])|(m[1818]&~m[1819]&m[1820]&~m[1822]&m[1823])|(~m[1818]&m[1819]&m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&m[1820]&~m[1822]&m[1823])|(m[1818]&m[1819]&m[1820]&m[1822]&m[1823]))):InitCond[1790];
    m[1826] = run?((((m[1823]&~m[1824]&~m[1825]&~m[1827]&~m[1828])|(~m[1823]&m[1824]&~m[1825]&~m[1827]&~m[1828])|(~m[1823]&~m[1824]&m[1825]&~m[1827]&~m[1828])|(m[1823]&m[1824]&m[1825]&m[1827]&~m[1828])|(~m[1823]&~m[1824]&~m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&~m[1825]&m[1827]&m[1828])|(m[1823]&~m[1824]&m[1825]&m[1827]&m[1828])|(~m[1823]&m[1824]&m[1825]&m[1827]&m[1828]))&UnbiasedRNG[896])|((m[1823]&m[1824]&~m[1825]&~m[1827]&~m[1828])|(m[1823]&~m[1824]&m[1825]&~m[1827]&~m[1828])|(~m[1823]&m[1824]&m[1825]&~m[1827]&~m[1828])|(m[1823]&m[1824]&m[1825]&~m[1827]&~m[1828])|(m[1823]&~m[1824]&~m[1825]&~m[1827]&m[1828])|(~m[1823]&m[1824]&~m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&~m[1825]&~m[1827]&m[1828])|(~m[1823]&~m[1824]&m[1825]&~m[1827]&m[1828])|(m[1823]&~m[1824]&m[1825]&~m[1827]&m[1828])|(~m[1823]&m[1824]&m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&m[1825]&~m[1827]&m[1828])|(m[1823]&m[1824]&m[1825]&m[1827]&m[1828]))):InitCond[1791];
    m[1831] = run?((((m[1828]&~m[1829]&~m[1830]&~m[1832]&~m[1833])|(~m[1828]&m[1829]&~m[1830]&~m[1832]&~m[1833])|(~m[1828]&~m[1829]&m[1830]&~m[1832]&~m[1833])|(m[1828]&m[1829]&m[1830]&m[1832]&~m[1833])|(~m[1828]&~m[1829]&~m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&~m[1830]&m[1832]&m[1833])|(m[1828]&~m[1829]&m[1830]&m[1832]&m[1833])|(~m[1828]&m[1829]&m[1830]&m[1832]&m[1833]))&UnbiasedRNG[897])|((m[1828]&m[1829]&~m[1830]&~m[1832]&~m[1833])|(m[1828]&~m[1829]&m[1830]&~m[1832]&~m[1833])|(~m[1828]&m[1829]&m[1830]&~m[1832]&~m[1833])|(m[1828]&m[1829]&m[1830]&~m[1832]&~m[1833])|(m[1828]&~m[1829]&~m[1830]&~m[1832]&m[1833])|(~m[1828]&m[1829]&~m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&~m[1830]&~m[1832]&m[1833])|(~m[1828]&~m[1829]&m[1830]&~m[1832]&m[1833])|(m[1828]&~m[1829]&m[1830]&~m[1832]&m[1833])|(~m[1828]&m[1829]&m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&m[1830]&~m[1832]&m[1833])|(m[1828]&m[1829]&m[1830]&m[1832]&m[1833]))):InitCond[1792];
    m[1836] = run?((((m[1833]&~m[1834]&~m[1835]&~m[1837]&~m[1838])|(~m[1833]&m[1834]&~m[1835]&~m[1837]&~m[1838])|(~m[1833]&~m[1834]&m[1835]&~m[1837]&~m[1838])|(m[1833]&m[1834]&m[1835]&m[1837]&~m[1838])|(~m[1833]&~m[1834]&~m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&~m[1835]&m[1837]&m[1838])|(m[1833]&~m[1834]&m[1835]&m[1837]&m[1838])|(~m[1833]&m[1834]&m[1835]&m[1837]&m[1838]))&UnbiasedRNG[898])|((m[1833]&m[1834]&~m[1835]&~m[1837]&~m[1838])|(m[1833]&~m[1834]&m[1835]&~m[1837]&~m[1838])|(~m[1833]&m[1834]&m[1835]&~m[1837]&~m[1838])|(m[1833]&m[1834]&m[1835]&~m[1837]&~m[1838])|(m[1833]&~m[1834]&~m[1835]&~m[1837]&m[1838])|(~m[1833]&m[1834]&~m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&~m[1835]&~m[1837]&m[1838])|(~m[1833]&~m[1834]&m[1835]&~m[1837]&m[1838])|(m[1833]&~m[1834]&m[1835]&~m[1837]&m[1838])|(~m[1833]&m[1834]&m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&m[1835]&~m[1837]&m[1838])|(m[1833]&m[1834]&m[1835]&m[1837]&m[1838]))):InitCond[1793];
    m[1841] = run?((((m[1838]&~m[1839]&~m[1840]&~m[1842]&~m[1843])|(~m[1838]&m[1839]&~m[1840]&~m[1842]&~m[1843])|(~m[1838]&~m[1839]&m[1840]&~m[1842]&~m[1843])|(m[1838]&m[1839]&m[1840]&m[1842]&~m[1843])|(~m[1838]&~m[1839]&~m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&~m[1840]&m[1842]&m[1843])|(m[1838]&~m[1839]&m[1840]&m[1842]&m[1843])|(~m[1838]&m[1839]&m[1840]&m[1842]&m[1843]))&UnbiasedRNG[899])|((m[1838]&m[1839]&~m[1840]&~m[1842]&~m[1843])|(m[1838]&~m[1839]&m[1840]&~m[1842]&~m[1843])|(~m[1838]&m[1839]&m[1840]&~m[1842]&~m[1843])|(m[1838]&m[1839]&m[1840]&~m[1842]&~m[1843])|(m[1838]&~m[1839]&~m[1840]&~m[1842]&m[1843])|(~m[1838]&m[1839]&~m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&~m[1840]&~m[1842]&m[1843])|(~m[1838]&~m[1839]&m[1840]&~m[1842]&m[1843])|(m[1838]&~m[1839]&m[1840]&~m[1842]&m[1843])|(~m[1838]&m[1839]&m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&m[1840]&~m[1842]&m[1843])|(m[1838]&m[1839]&m[1840]&m[1842]&m[1843]))):InitCond[1794];
    m[1846] = run?((((m[1843]&~m[1844]&~m[1845]&~m[1847]&~m[1848])|(~m[1843]&m[1844]&~m[1845]&~m[1847]&~m[1848])|(~m[1843]&~m[1844]&m[1845]&~m[1847]&~m[1848])|(m[1843]&m[1844]&m[1845]&m[1847]&~m[1848])|(~m[1843]&~m[1844]&~m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&~m[1845]&m[1847]&m[1848])|(m[1843]&~m[1844]&m[1845]&m[1847]&m[1848])|(~m[1843]&m[1844]&m[1845]&m[1847]&m[1848]))&UnbiasedRNG[900])|((m[1843]&m[1844]&~m[1845]&~m[1847]&~m[1848])|(m[1843]&~m[1844]&m[1845]&~m[1847]&~m[1848])|(~m[1843]&m[1844]&m[1845]&~m[1847]&~m[1848])|(m[1843]&m[1844]&m[1845]&~m[1847]&~m[1848])|(m[1843]&~m[1844]&~m[1845]&~m[1847]&m[1848])|(~m[1843]&m[1844]&~m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&~m[1845]&~m[1847]&m[1848])|(~m[1843]&~m[1844]&m[1845]&~m[1847]&m[1848])|(m[1843]&~m[1844]&m[1845]&~m[1847]&m[1848])|(~m[1843]&m[1844]&m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&m[1845]&~m[1847]&m[1848])|(m[1843]&m[1844]&m[1845]&m[1847]&m[1848]))):InitCond[1795];
    m[1856] = run?((((m[1853]&~m[1854]&~m[1855]&~m[1857]&~m[1858])|(~m[1853]&m[1854]&~m[1855]&~m[1857]&~m[1858])|(~m[1853]&~m[1854]&m[1855]&~m[1857]&~m[1858])|(m[1853]&m[1854]&m[1855]&m[1857]&~m[1858])|(~m[1853]&~m[1854]&~m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&~m[1855]&m[1857]&m[1858])|(m[1853]&~m[1854]&m[1855]&m[1857]&m[1858])|(~m[1853]&m[1854]&m[1855]&m[1857]&m[1858]))&UnbiasedRNG[901])|((m[1853]&m[1854]&~m[1855]&~m[1857]&~m[1858])|(m[1853]&~m[1854]&m[1855]&~m[1857]&~m[1858])|(~m[1853]&m[1854]&m[1855]&~m[1857]&~m[1858])|(m[1853]&m[1854]&m[1855]&~m[1857]&~m[1858])|(m[1853]&~m[1854]&~m[1855]&~m[1857]&m[1858])|(~m[1853]&m[1854]&~m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&~m[1855]&~m[1857]&m[1858])|(~m[1853]&~m[1854]&m[1855]&~m[1857]&m[1858])|(m[1853]&~m[1854]&m[1855]&~m[1857]&m[1858])|(~m[1853]&m[1854]&m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&m[1855]&~m[1857]&m[1858])|(m[1853]&m[1854]&m[1855]&m[1857]&m[1858]))):InitCond[1796];
    m[1861] = run?((((m[1858]&~m[1859]&~m[1860]&~m[1862]&~m[1863])|(~m[1858]&m[1859]&~m[1860]&~m[1862]&~m[1863])|(~m[1858]&~m[1859]&m[1860]&~m[1862]&~m[1863])|(m[1858]&m[1859]&m[1860]&m[1862]&~m[1863])|(~m[1858]&~m[1859]&~m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&~m[1860]&m[1862]&m[1863])|(m[1858]&~m[1859]&m[1860]&m[1862]&m[1863])|(~m[1858]&m[1859]&m[1860]&m[1862]&m[1863]))&UnbiasedRNG[902])|((m[1858]&m[1859]&~m[1860]&~m[1862]&~m[1863])|(m[1858]&~m[1859]&m[1860]&~m[1862]&~m[1863])|(~m[1858]&m[1859]&m[1860]&~m[1862]&~m[1863])|(m[1858]&m[1859]&m[1860]&~m[1862]&~m[1863])|(m[1858]&~m[1859]&~m[1860]&~m[1862]&m[1863])|(~m[1858]&m[1859]&~m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&~m[1860]&~m[1862]&m[1863])|(~m[1858]&~m[1859]&m[1860]&~m[1862]&m[1863])|(m[1858]&~m[1859]&m[1860]&~m[1862]&m[1863])|(~m[1858]&m[1859]&m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&m[1860]&~m[1862]&m[1863])|(m[1858]&m[1859]&m[1860]&m[1862]&m[1863]))):InitCond[1797];
    m[1866] = run?((((m[1863]&~m[1864]&~m[1865]&~m[1867]&~m[1868])|(~m[1863]&m[1864]&~m[1865]&~m[1867]&~m[1868])|(~m[1863]&~m[1864]&m[1865]&~m[1867]&~m[1868])|(m[1863]&m[1864]&m[1865]&m[1867]&~m[1868])|(~m[1863]&~m[1864]&~m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&~m[1865]&m[1867]&m[1868])|(m[1863]&~m[1864]&m[1865]&m[1867]&m[1868])|(~m[1863]&m[1864]&m[1865]&m[1867]&m[1868]))&UnbiasedRNG[903])|((m[1863]&m[1864]&~m[1865]&~m[1867]&~m[1868])|(m[1863]&~m[1864]&m[1865]&~m[1867]&~m[1868])|(~m[1863]&m[1864]&m[1865]&~m[1867]&~m[1868])|(m[1863]&m[1864]&m[1865]&~m[1867]&~m[1868])|(m[1863]&~m[1864]&~m[1865]&~m[1867]&m[1868])|(~m[1863]&m[1864]&~m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&~m[1865]&~m[1867]&m[1868])|(~m[1863]&~m[1864]&m[1865]&~m[1867]&m[1868])|(m[1863]&~m[1864]&m[1865]&~m[1867]&m[1868])|(~m[1863]&m[1864]&m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&m[1865]&~m[1867]&m[1868])|(m[1863]&m[1864]&m[1865]&m[1867]&m[1868]))):InitCond[1798];
    m[1871] = run?((((m[1868]&~m[1869]&~m[1870]&~m[1872]&~m[1873])|(~m[1868]&m[1869]&~m[1870]&~m[1872]&~m[1873])|(~m[1868]&~m[1869]&m[1870]&~m[1872]&~m[1873])|(m[1868]&m[1869]&m[1870]&m[1872]&~m[1873])|(~m[1868]&~m[1869]&~m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&~m[1870]&m[1872]&m[1873])|(m[1868]&~m[1869]&m[1870]&m[1872]&m[1873])|(~m[1868]&m[1869]&m[1870]&m[1872]&m[1873]))&UnbiasedRNG[904])|((m[1868]&m[1869]&~m[1870]&~m[1872]&~m[1873])|(m[1868]&~m[1869]&m[1870]&~m[1872]&~m[1873])|(~m[1868]&m[1869]&m[1870]&~m[1872]&~m[1873])|(m[1868]&m[1869]&m[1870]&~m[1872]&~m[1873])|(m[1868]&~m[1869]&~m[1870]&~m[1872]&m[1873])|(~m[1868]&m[1869]&~m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&~m[1870]&~m[1872]&m[1873])|(~m[1868]&~m[1869]&m[1870]&~m[1872]&m[1873])|(m[1868]&~m[1869]&m[1870]&~m[1872]&m[1873])|(~m[1868]&m[1869]&m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&m[1870]&~m[1872]&m[1873])|(m[1868]&m[1869]&m[1870]&m[1872]&m[1873]))):InitCond[1799];
    m[1876] = run?((((m[1873]&~m[1874]&~m[1875]&~m[1877]&~m[1878])|(~m[1873]&m[1874]&~m[1875]&~m[1877]&~m[1878])|(~m[1873]&~m[1874]&m[1875]&~m[1877]&~m[1878])|(m[1873]&m[1874]&m[1875]&m[1877]&~m[1878])|(~m[1873]&~m[1874]&~m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&~m[1875]&m[1877]&m[1878])|(m[1873]&~m[1874]&m[1875]&m[1877]&m[1878])|(~m[1873]&m[1874]&m[1875]&m[1877]&m[1878]))&UnbiasedRNG[905])|((m[1873]&m[1874]&~m[1875]&~m[1877]&~m[1878])|(m[1873]&~m[1874]&m[1875]&~m[1877]&~m[1878])|(~m[1873]&m[1874]&m[1875]&~m[1877]&~m[1878])|(m[1873]&m[1874]&m[1875]&~m[1877]&~m[1878])|(m[1873]&~m[1874]&~m[1875]&~m[1877]&m[1878])|(~m[1873]&m[1874]&~m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&~m[1875]&~m[1877]&m[1878])|(~m[1873]&~m[1874]&m[1875]&~m[1877]&m[1878])|(m[1873]&~m[1874]&m[1875]&~m[1877]&m[1878])|(~m[1873]&m[1874]&m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&m[1875]&~m[1877]&m[1878])|(m[1873]&m[1874]&m[1875]&m[1877]&m[1878]))):InitCond[1800];
    m[1881] = run?((((m[1878]&~m[1879]&~m[1880]&~m[1882]&~m[1883])|(~m[1878]&m[1879]&~m[1880]&~m[1882]&~m[1883])|(~m[1878]&~m[1879]&m[1880]&~m[1882]&~m[1883])|(m[1878]&m[1879]&m[1880]&m[1882]&~m[1883])|(~m[1878]&~m[1879]&~m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&~m[1880]&m[1882]&m[1883])|(m[1878]&~m[1879]&m[1880]&m[1882]&m[1883])|(~m[1878]&m[1879]&m[1880]&m[1882]&m[1883]))&UnbiasedRNG[906])|((m[1878]&m[1879]&~m[1880]&~m[1882]&~m[1883])|(m[1878]&~m[1879]&m[1880]&~m[1882]&~m[1883])|(~m[1878]&m[1879]&m[1880]&~m[1882]&~m[1883])|(m[1878]&m[1879]&m[1880]&~m[1882]&~m[1883])|(m[1878]&~m[1879]&~m[1880]&~m[1882]&m[1883])|(~m[1878]&m[1879]&~m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&~m[1880]&~m[1882]&m[1883])|(~m[1878]&~m[1879]&m[1880]&~m[1882]&m[1883])|(m[1878]&~m[1879]&m[1880]&~m[1882]&m[1883])|(~m[1878]&m[1879]&m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&m[1880]&~m[1882]&m[1883])|(m[1878]&m[1879]&m[1880]&m[1882]&m[1883]))):InitCond[1801];
    m[1886] = run?((((m[1883]&~m[1884]&~m[1885]&~m[1887]&~m[1888])|(~m[1883]&m[1884]&~m[1885]&~m[1887]&~m[1888])|(~m[1883]&~m[1884]&m[1885]&~m[1887]&~m[1888])|(m[1883]&m[1884]&m[1885]&m[1887]&~m[1888])|(~m[1883]&~m[1884]&~m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&~m[1885]&m[1887]&m[1888])|(m[1883]&~m[1884]&m[1885]&m[1887]&m[1888])|(~m[1883]&m[1884]&m[1885]&m[1887]&m[1888]))&UnbiasedRNG[907])|((m[1883]&m[1884]&~m[1885]&~m[1887]&~m[1888])|(m[1883]&~m[1884]&m[1885]&~m[1887]&~m[1888])|(~m[1883]&m[1884]&m[1885]&~m[1887]&~m[1888])|(m[1883]&m[1884]&m[1885]&~m[1887]&~m[1888])|(m[1883]&~m[1884]&~m[1885]&~m[1887]&m[1888])|(~m[1883]&m[1884]&~m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&~m[1885]&~m[1887]&m[1888])|(~m[1883]&~m[1884]&m[1885]&~m[1887]&m[1888])|(m[1883]&~m[1884]&m[1885]&~m[1887]&m[1888])|(~m[1883]&m[1884]&m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&m[1885]&~m[1887]&m[1888])|(m[1883]&m[1884]&m[1885]&m[1887]&m[1888]))):InitCond[1802];
    m[1891] = run?((((m[1888]&~m[1889]&~m[1890]&~m[1892]&~m[1893])|(~m[1888]&m[1889]&~m[1890]&~m[1892]&~m[1893])|(~m[1888]&~m[1889]&m[1890]&~m[1892]&~m[1893])|(m[1888]&m[1889]&m[1890]&m[1892]&~m[1893])|(~m[1888]&~m[1889]&~m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&~m[1890]&m[1892]&m[1893])|(m[1888]&~m[1889]&m[1890]&m[1892]&m[1893])|(~m[1888]&m[1889]&m[1890]&m[1892]&m[1893]))&UnbiasedRNG[908])|((m[1888]&m[1889]&~m[1890]&~m[1892]&~m[1893])|(m[1888]&~m[1889]&m[1890]&~m[1892]&~m[1893])|(~m[1888]&m[1889]&m[1890]&~m[1892]&~m[1893])|(m[1888]&m[1889]&m[1890]&~m[1892]&~m[1893])|(m[1888]&~m[1889]&~m[1890]&~m[1892]&m[1893])|(~m[1888]&m[1889]&~m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&~m[1890]&~m[1892]&m[1893])|(~m[1888]&~m[1889]&m[1890]&~m[1892]&m[1893])|(m[1888]&~m[1889]&m[1890]&~m[1892]&m[1893])|(~m[1888]&m[1889]&m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&m[1890]&~m[1892]&m[1893])|(m[1888]&m[1889]&m[1890]&m[1892]&m[1893]))):InitCond[1803];
    m[1896] = run?((((m[1893]&~m[1894]&~m[1895]&~m[1897]&~m[1898])|(~m[1893]&m[1894]&~m[1895]&~m[1897]&~m[1898])|(~m[1893]&~m[1894]&m[1895]&~m[1897]&~m[1898])|(m[1893]&m[1894]&m[1895]&m[1897]&~m[1898])|(~m[1893]&~m[1894]&~m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&~m[1895]&m[1897]&m[1898])|(m[1893]&~m[1894]&m[1895]&m[1897]&m[1898])|(~m[1893]&m[1894]&m[1895]&m[1897]&m[1898]))&UnbiasedRNG[909])|((m[1893]&m[1894]&~m[1895]&~m[1897]&~m[1898])|(m[1893]&~m[1894]&m[1895]&~m[1897]&~m[1898])|(~m[1893]&m[1894]&m[1895]&~m[1897]&~m[1898])|(m[1893]&m[1894]&m[1895]&~m[1897]&~m[1898])|(m[1893]&~m[1894]&~m[1895]&~m[1897]&m[1898])|(~m[1893]&m[1894]&~m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&~m[1895]&~m[1897]&m[1898])|(~m[1893]&~m[1894]&m[1895]&~m[1897]&m[1898])|(m[1893]&~m[1894]&m[1895]&~m[1897]&m[1898])|(~m[1893]&m[1894]&m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&m[1895]&~m[1897]&m[1898])|(m[1893]&m[1894]&m[1895]&m[1897]&m[1898]))):InitCond[1804];
    m[1906] = run?((((m[1903]&~m[1904]&~m[1905]&~m[1907]&~m[1908])|(~m[1903]&m[1904]&~m[1905]&~m[1907]&~m[1908])|(~m[1903]&~m[1904]&m[1905]&~m[1907]&~m[1908])|(m[1903]&m[1904]&m[1905]&m[1907]&~m[1908])|(~m[1903]&~m[1904]&~m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&~m[1905]&m[1907]&m[1908])|(m[1903]&~m[1904]&m[1905]&m[1907]&m[1908])|(~m[1903]&m[1904]&m[1905]&m[1907]&m[1908]))&UnbiasedRNG[910])|((m[1903]&m[1904]&~m[1905]&~m[1907]&~m[1908])|(m[1903]&~m[1904]&m[1905]&~m[1907]&~m[1908])|(~m[1903]&m[1904]&m[1905]&~m[1907]&~m[1908])|(m[1903]&m[1904]&m[1905]&~m[1907]&~m[1908])|(m[1903]&~m[1904]&~m[1905]&~m[1907]&m[1908])|(~m[1903]&m[1904]&~m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&~m[1905]&~m[1907]&m[1908])|(~m[1903]&~m[1904]&m[1905]&~m[1907]&m[1908])|(m[1903]&~m[1904]&m[1905]&~m[1907]&m[1908])|(~m[1903]&m[1904]&m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&m[1905]&~m[1907]&m[1908])|(m[1903]&m[1904]&m[1905]&m[1907]&m[1908]))):InitCond[1805];
    m[1911] = run?((((m[1908]&~m[1909]&~m[1910]&~m[1912]&~m[1913])|(~m[1908]&m[1909]&~m[1910]&~m[1912]&~m[1913])|(~m[1908]&~m[1909]&m[1910]&~m[1912]&~m[1913])|(m[1908]&m[1909]&m[1910]&m[1912]&~m[1913])|(~m[1908]&~m[1909]&~m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&~m[1910]&m[1912]&m[1913])|(m[1908]&~m[1909]&m[1910]&m[1912]&m[1913])|(~m[1908]&m[1909]&m[1910]&m[1912]&m[1913]))&UnbiasedRNG[911])|((m[1908]&m[1909]&~m[1910]&~m[1912]&~m[1913])|(m[1908]&~m[1909]&m[1910]&~m[1912]&~m[1913])|(~m[1908]&m[1909]&m[1910]&~m[1912]&~m[1913])|(m[1908]&m[1909]&m[1910]&~m[1912]&~m[1913])|(m[1908]&~m[1909]&~m[1910]&~m[1912]&m[1913])|(~m[1908]&m[1909]&~m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&~m[1910]&~m[1912]&m[1913])|(~m[1908]&~m[1909]&m[1910]&~m[1912]&m[1913])|(m[1908]&~m[1909]&m[1910]&~m[1912]&m[1913])|(~m[1908]&m[1909]&m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&m[1910]&~m[1912]&m[1913])|(m[1908]&m[1909]&m[1910]&m[1912]&m[1913]))):InitCond[1806];
    m[1916] = run?((((m[1913]&~m[1914]&~m[1915]&~m[1917]&~m[1918])|(~m[1913]&m[1914]&~m[1915]&~m[1917]&~m[1918])|(~m[1913]&~m[1914]&m[1915]&~m[1917]&~m[1918])|(m[1913]&m[1914]&m[1915]&m[1917]&~m[1918])|(~m[1913]&~m[1914]&~m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&~m[1915]&m[1917]&m[1918])|(m[1913]&~m[1914]&m[1915]&m[1917]&m[1918])|(~m[1913]&m[1914]&m[1915]&m[1917]&m[1918]))&UnbiasedRNG[912])|((m[1913]&m[1914]&~m[1915]&~m[1917]&~m[1918])|(m[1913]&~m[1914]&m[1915]&~m[1917]&~m[1918])|(~m[1913]&m[1914]&m[1915]&~m[1917]&~m[1918])|(m[1913]&m[1914]&m[1915]&~m[1917]&~m[1918])|(m[1913]&~m[1914]&~m[1915]&~m[1917]&m[1918])|(~m[1913]&m[1914]&~m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&~m[1915]&~m[1917]&m[1918])|(~m[1913]&~m[1914]&m[1915]&~m[1917]&m[1918])|(m[1913]&~m[1914]&m[1915]&~m[1917]&m[1918])|(~m[1913]&m[1914]&m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&m[1915]&~m[1917]&m[1918])|(m[1913]&m[1914]&m[1915]&m[1917]&m[1918]))):InitCond[1807];
    m[1921] = run?((((m[1918]&~m[1919]&~m[1920]&~m[1922]&~m[1923])|(~m[1918]&m[1919]&~m[1920]&~m[1922]&~m[1923])|(~m[1918]&~m[1919]&m[1920]&~m[1922]&~m[1923])|(m[1918]&m[1919]&m[1920]&m[1922]&~m[1923])|(~m[1918]&~m[1919]&~m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&~m[1920]&m[1922]&m[1923])|(m[1918]&~m[1919]&m[1920]&m[1922]&m[1923])|(~m[1918]&m[1919]&m[1920]&m[1922]&m[1923]))&UnbiasedRNG[913])|((m[1918]&m[1919]&~m[1920]&~m[1922]&~m[1923])|(m[1918]&~m[1919]&m[1920]&~m[1922]&~m[1923])|(~m[1918]&m[1919]&m[1920]&~m[1922]&~m[1923])|(m[1918]&m[1919]&m[1920]&~m[1922]&~m[1923])|(m[1918]&~m[1919]&~m[1920]&~m[1922]&m[1923])|(~m[1918]&m[1919]&~m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&~m[1920]&~m[1922]&m[1923])|(~m[1918]&~m[1919]&m[1920]&~m[1922]&m[1923])|(m[1918]&~m[1919]&m[1920]&~m[1922]&m[1923])|(~m[1918]&m[1919]&m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&m[1920]&~m[1922]&m[1923])|(m[1918]&m[1919]&m[1920]&m[1922]&m[1923]))):InitCond[1808];
    m[1926] = run?((((m[1923]&~m[1924]&~m[1925]&~m[1927]&~m[1928])|(~m[1923]&m[1924]&~m[1925]&~m[1927]&~m[1928])|(~m[1923]&~m[1924]&m[1925]&~m[1927]&~m[1928])|(m[1923]&m[1924]&m[1925]&m[1927]&~m[1928])|(~m[1923]&~m[1924]&~m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&~m[1925]&m[1927]&m[1928])|(m[1923]&~m[1924]&m[1925]&m[1927]&m[1928])|(~m[1923]&m[1924]&m[1925]&m[1927]&m[1928]))&UnbiasedRNG[914])|((m[1923]&m[1924]&~m[1925]&~m[1927]&~m[1928])|(m[1923]&~m[1924]&m[1925]&~m[1927]&~m[1928])|(~m[1923]&m[1924]&m[1925]&~m[1927]&~m[1928])|(m[1923]&m[1924]&m[1925]&~m[1927]&~m[1928])|(m[1923]&~m[1924]&~m[1925]&~m[1927]&m[1928])|(~m[1923]&m[1924]&~m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&~m[1925]&~m[1927]&m[1928])|(~m[1923]&~m[1924]&m[1925]&~m[1927]&m[1928])|(m[1923]&~m[1924]&m[1925]&~m[1927]&m[1928])|(~m[1923]&m[1924]&m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&m[1925]&~m[1927]&m[1928])|(m[1923]&m[1924]&m[1925]&m[1927]&m[1928]))):InitCond[1809];
    m[1931] = run?((((m[1928]&~m[1929]&~m[1930]&~m[1932]&~m[1933])|(~m[1928]&m[1929]&~m[1930]&~m[1932]&~m[1933])|(~m[1928]&~m[1929]&m[1930]&~m[1932]&~m[1933])|(m[1928]&m[1929]&m[1930]&m[1932]&~m[1933])|(~m[1928]&~m[1929]&~m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&~m[1930]&m[1932]&m[1933])|(m[1928]&~m[1929]&m[1930]&m[1932]&m[1933])|(~m[1928]&m[1929]&m[1930]&m[1932]&m[1933]))&UnbiasedRNG[915])|((m[1928]&m[1929]&~m[1930]&~m[1932]&~m[1933])|(m[1928]&~m[1929]&m[1930]&~m[1932]&~m[1933])|(~m[1928]&m[1929]&m[1930]&~m[1932]&~m[1933])|(m[1928]&m[1929]&m[1930]&~m[1932]&~m[1933])|(m[1928]&~m[1929]&~m[1930]&~m[1932]&m[1933])|(~m[1928]&m[1929]&~m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&~m[1930]&~m[1932]&m[1933])|(~m[1928]&~m[1929]&m[1930]&~m[1932]&m[1933])|(m[1928]&~m[1929]&m[1930]&~m[1932]&m[1933])|(~m[1928]&m[1929]&m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&m[1930]&~m[1932]&m[1933])|(m[1928]&m[1929]&m[1930]&m[1932]&m[1933]))):InitCond[1810];
    m[1936] = run?((((m[1933]&~m[1934]&~m[1935]&~m[1937]&~m[1938])|(~m[1933]&m[1934]&~m[1935]&~m[1937]&~m[1938])|(~m[1933]&~m[1934]&m[1935]&~m[1937]&~m[1938])|(m[1933]&m[1934]&m[1935]&m[1937]&~m[1938])|(~m[1933]&~m[1934]&~m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&~m[1935]&m[1937]&m[1938])|(m[1933]&~m[1934]&m[1935]&m[1937]&m[1938])|(~m[1933]&m[1934]&m[1935]&m[1937]&m[1938]))&UnbiasedRNG[916])|((m[1933]&m[1934]&~m[1935]&~m[1937]&~m[1938])|(m[1933]&~m[1934]&m[1935]&~m[1937]&~m[1938])|(~m[1933]&m[1934]&m[1935]&~m[1937]&~m[1938])|(m[1933]&m[1934]&m[1935]&~m[1937]&~m[1938])|(m[1933]&~m[1934]&~m[1935]&~m[1937]&m[1938])|(~m[1933]&m[1934]&~m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&~m[1935]&~m[1937]&m[1938])|(~m[1933]&~m[1934]&m[1935]&~m[1937]&m[1938])|(m[1933]&~m[1934]&m[1935]&~m[1937]&m[1938])|(~m[1933]&m[1934]&m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&m[1935]&~m[1937]&m[1938])|(m[1933]&m[1934]&m[1935]&m[1937]&m[1938]))):InitCond[1811];
    m[1941] = run?((((m[1938]&~m[1939]&~m[1940]&~m[1942]&~m[1943])|(~m[1938]&m[1939]&~m[1940]&~m[1942]&~m[1943])|(~m[1938]&~m[1939]&m[1940]&~m[1942]&~m[1943])|(m[1938]&m[1939]&m[1940]&m[1942]&~m[1943])|(~m[1938]&~m[1939]&~m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&~m[1940]&m[1942]&m[1943])|(m[1938]&~m[1939]&m[1940]&m[1942]&m[1943])|(~m[1938]&m[1939]&m[1940]&m[1942]&m[1943]))&UnbiasedRNG[917])|((m[1938]&m[1939]&~m[1940]&~m[1942]&~m[1943])|(m[1938]&~m[1939]&m[1940]&~m[1942]&~m[1943])|(~m[1938]&m[1939]&m[1940]&~m[1942]&~m[1943])|(m[1938]&m[1939]&m[1940]&~m[1942]&~m[1943])|(m[1938]&~m[1939]&~m[1940]&~m[1942]&m[1943])|(~m[1938]&m[1939]&~m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&~m[1940]&~m[1942]&m[1943])|(~m[1938]&~m[1939]&m[1940]&~m[1942]&m[1943])|(m[1938]&~m[1939]&m[1940]&~m[1942]&m[1943])|(~m[1938]&m[1939]&m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&m[1940]&~m[1942]&m[1943])|(m[1938]&m[1939]&m[1940]&m[1942]&m[1943]))):InitCond[1812];
    m[1951] = run?((((m[1948]&~m[1949]&~m[1950]&~m[1952]&~m[1953])|(~m[1948]&m[1949]&~m[1950]&~m[1952]&~m[1953])|(~m[1948]&~m[1949]&m[1950]&~m[1952]&~m[1953])|(m[1948]&m[1949]&m[1950]&m[1952]&~m[1953])|(~m[1948]&~m[1949]&~m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&~m[1950]&m[1952]&m[1953])|(m[1948]&~m[1949]&m[1950]&m[1952]&m[1953])|(~m[1948]&m[1949]&m[1950]&m[1952]&m[1953]))&UnbiasedRNG[918])|((m[1948]&m[1949]&~m[1950]&~m[1952]&~m[1953])|(m[1948]&~m[1949]&m[1950]&~m[1952]&~m[1953])|(~m[1948]&m[1949]&m[1950]&~m[1952]&~m[1953])|(m[1948]&m[1949]&m[1950]&~m[1952]&~m[1953])|(m[1948]&~m[1949]&~m[1950]&~m[1952]&m[1953])|(~m[1948]&m[1949]&~m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&~m[1950]&~m[1952]&m[1953])|(~m[1948]&~m[1949]&m[1950]&~m[1952]&m[1953])|(m[1948]&~m[1949]&m[1950]&~m[1952]&m[1953])|(~m[1948]&m[1949]&m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&m[1950]&~m[1952]&m[1953])|(m[1948]&m[1949]&m[1950]&m[1952]&m[1953]))):InitCond[1813];
    m[1956] = run?((((m[1953]&~m[1954]&~m[1955]&~m[1957]&~m[1958])|(~m[1953]&m[1954]&~m[1955]&~m[1957]&~m[1958])|(~m[1953]&~m[1954]&m[1955]&~m[1957]&~m[1958])|(m[1953]&m[1954]&m[1955]&m[1957]&~m[1958])|(~m[1953]&~m[1954]&~m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&~m[1955]&m[1957]&m[1958])|(m[1953]&~m[1954]&m[1955]&m[1957]&m[1958])|(~m[1953]&m[1954]&m[1955]&m[1957]&m[1958]))&UnbiasedRNG[919])|((m[1953]&m[1954]&~m[1955]&~m[1957]&~m[1958])|(m[1953]&~m[1954]&m[1955]&~m[1957]&~m[1958])|(~m[1953]&m[1954]&m[1955]&~m[1957]&~m[1958])|(m[1953]&m[1954]&m[1955]&~m[1957]&~m[1958])|(m[1953]&~m[1954]&~m[1955]&~m[1957]&m[1958])|(~m[1953]&m[1954]&~m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&~m[1955]&~m[1957]&m[1958])|(~m[1953]&~m[1954]&m[1955]&~m[1957]&m[1958])|(m[1953]&~m[1954]&m[1955]&~m[1957]&m[1958])|(~m[1953]&m[1954]&m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&m[1955]&~m[1957]&m[1958])|(m[1953]&m[1954]&m[1955]&m[1957]&m[1958]))):InitCond[1814];
    m[1961] = run?((((m[1958]&~m[1959]&~m[1960]&~m[1962]&~m[1963])|(~m[1958]&m[1959]&~m[1960]&~m[1962]&~m[1963])|(~m[1958]&~m[1959]&m[1960]&~m[1962]&~m[1963])|(m[1958]&m[1959]&m[1960]&m[1962]&~m[1963])|(~m[1958]&~m[1959]&~m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&~m[1960]&m[1962]&m[1963])|(m[1958]&~m[1959]&m[1960]&m[1962]&m[1963])|(~m[1958]&m[1959]&m[1960]&m[1962]&m[1963]))&UnbiasedRNG[920])|((m[1958]&m[1959]&~m[1960]&~m[1962]&~m[1963])|(m[1958]&~m[1959]&m[1960]&~m[1962]&~m[1963])|(~m[1958]&m[1959]&m[1960]&~m[1962]&~m[1963])|(m[1958]&m[1959]&m[1960]&~m[1962]&~m[1963])|(m[1958]&~m[1959]&~m[1960]&~m[1962]&m[1963])|(~m[1958]&m[1959]&~m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&~m[1960]&~m[1962]&m[1963])|(~m[1958]&~m[1959]&m[1960]&~m[1962]&m[1963])|(m[1958]&~m[1959]&m[1960]&~m[1962]&m[1963])|(~m[1958]&m[1959]&m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&m[1960]&~m[1962]&m[1963])|(m[1958]&m[1959]&m[1960]&m[1962]&m[1963]))):InitCond[1815];
    m[1966] = run?((((m[1963]&~m[1964]&~m[1965]&~m[1967]&~m[1968])|(~m[1963]&m[1964]&~m[1965]&~m[1967]&~m[1968])|(~m[1963]&~m[1964]&m[1965]&~m[1967]&~m[1968])|(m[1963]&m[1964]&m[1965]&m[1967]&~m[1968])|(~m[1963]&~m[1964]&~m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&~m[1965]&m[1967]&m[1968])|(m[1963]&~m[1964]&m[1965]&m[1967]&m[1968])|(~m[1963]&m[1964]&m[1965]&m[1967]&m[1968]))&UnbiasedRNG[921])|((m[1963]&m[1964]&~m[1965]&~m[1967]&~m[1968])|(m[1963]&~m[1964]&m[1965]&~m[1967]&~m[1968])|(~m[1963]&m[1964]&m[1965]&~m[1967]&~m[1968])|(m[1963]&m[1964]&m[1965]&~m[1967]&~m[1968])|(m[1963]&~m[1964]&~m[1965]&~m[1967]&m[1968])|(~m[1963]&m[1964]&~m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&~m[1965]&~m[1967]&m[1968])|(~m[1963]&~m[1964]&m[1965]&~m[1967]&m[1968])|(m[1963]&~m[1964]&m[1965]&~m[1967]&m[1968])|(~m[1963]&m[1964]&m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&m[1965]&~m[1967]&m[1968])|(m[1963]&m[1964]&m[1965]&m[1967]&m[1968]))):InitCond[1816];
    m[1971] = run?((((m[1968]&~m[1969]&~m[1970]&~m[1972]&~m[1973])|(~m[1968]&m[1969]&~m[1970]&~m[1972]&~m[1973])|(~m[1968]&~m[1969]&m[1970]&~m[1972]&~m[1973])|(m[1968]&m[1969]&m[1970]&m[1972]&~m[1973])|(~m[1968]&~m[1969]&~m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&~m[1970]&m[1972]&m[1973])|(m[1968]&~m[1969]&m[1970]&m[1972]&m[1973])|(~m[1968]&m[1969]&m[1970]&m[1972]&m[1973]))&UnbiasedRNG[922])|((m[1968]&m[1969]&~m[1970]&~m[1972]&~m[1973])|(m[1968]&~m[1969]&m[1970]&~m[1972]&~m[1973])|(~m[1968]&m[1969]&m[1970]&~m[1972]&~m[1973])|(m[1968]&m[1969]&m[1970]&~m[1972]&~m[1973])|(m[1968]&~m[1969]&~m[1970]&~m[1972]&m[1973])|(~m[1968]&m[1969]&~m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&~m[1970]&~m[1972]&m[1973])|(~m[1968]&~m[1969]&m[1970]&~m[1972]&m[1973])|(m[1968]&~m[1969]&m[1970]&~m[1972]&m[1973])|(~m[1968]&m[1969]&m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&m[1970]&~m[1972]&m[1973])|(m[1968]&m[1969]&m[1970]&m[1972]&m[1973]))):InitCond[1817];
    m[1976] = run?((((m[1973]&~m[1974]&~m[1975]&~m[1977]&~m[1978])|(~m[1973]&m[1974]&~m[1975]&~m[1977]&~m[1978])|(~m[1973]&~m[1974]&m[1975]&~m[1977]&~m[1978])|(m[1973]&m[1974]&m[1975]&m[1977]&~m[1978])|(~m[1973]&~m[1974]&~m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&~m[1975]&m[1977]&m[1978])|(m[1973]&~m[1974]&m[1975]&m[1977]&m[1978])|(~m[1973]&m[1974]&m[1975]&m[1977]&m[1978]))&UnbiasedRNG[923])|((m[1973]&m[1974]&~m[1975]&~m[1977]&~m[1978])|(m[1973]&~m[1974]&m[1975]&~m[1977]&~m[1978])|(~m[1973]&m[1974]&m[1975]&~m[1977]&~m[1978])|(m[1973]&m[1974]&m[1975]&~m[1977]&~m[1978])|(m[1973]&~m[1974]&~m[1975]&~m[1977]&m[1978])|(~m[1973]&m[1974]&~m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&~m[1975]&~m[1977]&m[1978])|(~m[1973]&~m[1974]&m[1975]&~m[1977]&m[1978])|(m[1973]&~m[1974]&m[1975]&~m[1977]&m[1978])|(~m[1973]&m[1974]&m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&m[1975]&~m[1977]&m[1978])|(m[1973]&m[1974]&m[1975]&m[1977]&m[1978]))):InitCond[1818];
    m[1981] = run?((((m[1978]&~m[1979]&~m[1980]&~m[1982]&~m[1983])|(~m[1978]&m[1979]&~m[1980]&~m[1982]&~m[1983])|(~m[1978]&~m[1979]&m[1980]&~m[1982]&~m[1983])|(m[1978]&m[1979]&m[1980]&m[1982]&~m[1983])|(~m[1978]&~m[1979]&~m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&~m[1980]&m[1982]&m[1983])|(m[1978]&~m[1979]&m[1980]&m[1982]&m[1983])|(~m[1978]&m[1979]&m[1980]&m[1982]&m[1983]))&UnbiasedRNG[924])|((m[1978]&m[1979]&~m[1980]&~m[1982]&~m[1983])|(m[1978]&~m[1979]&m[1980]&~m[1982]&~m[1983])|(~m[1978]&m[1979]&m[1980]&~m[1982]&~m[1983])|(m[1978]&m[1979]&m[1980]&~m[1982]&~m[1983])|(m[1978]&~m[1979]&~m[1980]&~m[1982]&m[1983])|(~m[1978]&m[1979]&~m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&~m[1980]&~m[1982]&m[1983])|(~m[1978]&~m[1979]&m[1980]&~m[1982]&m[1983])|(m[1978]&~m[1979]&m[1980]&~m[1982]&m[1983])|(~m[1978]&m[1979]&m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&m[1980]&~m[1982]&m[1983])|(m[1978]&m[1979]&m[1980]&m[1982]&m[1983]))):InitCond[1819];
    m[1991] = run?((((m[1988]&~m[1989]&~m[1990]&~m[1992]&~m[1993])|(~m[1988]&m[1989]&~m[1990]&~m[1992]&~m[1993])|(~m[1988]&~m[1989]&m[1990]&~m[1992]&~m[1993])|(m[1988]&m[1989]&m[1990]&m[1992]&~m[1993])|(~m[1988]&~m[1989]&~m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&~m[1990]&m[1992]&m[1993])|(m[1988]&~m[1989]&m[1990]&m[1992]&m[1993])|(~m[1988]&m[1989]&m[1990]&m[1992]&m[1993]))&UnbiasedRNG[925])|((m[1988]&m[1989]&~m[1990]&~m[1992]&~m[1993])|(m[1988]&~m[1989]&m[1990]&~m[1992]&~m[1993])|(~m[1988]&m[1989]&m[1990]&~m[1992]&~m[1993])|(m[1988]&m[1989]&m[1990]&~m[1992]&~m[1993])|(m[1988]&~m[1989]&~m[1990]&~m[1992]&m[1993])|(~m[1988]&m[1989]&~m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&~m[1990]&~m[1992]&m[1993])|(~m[1988]&~m[1989]&m[1990]&~m[1992]&m[1993])|(m[1988]&~m[1989]&m[1990]&~m[1992]&m[1993])|(~m[1988]&m[1989]&m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&m[1990]&~m[1992]&m[1993])|(m[1988]&m[1989]&m[1990]&m[1992]&m[1993]))):InitCond[1820];
    m[1996] = run?((((m[1993]&~m[1994]&~m[1995]&~m[1997]&~m[1998])|(~m[1993]&m[1994]&~m[1995]&~m[1997]&~m[1998])|(~m[1993]&~m[1994]&m[1995]&~m[1997]&~m[1998])|(m[1993]&m[1994]&m[1995]&m[1997]&~m[1998])|(~m[1993]&~m[1994]&~m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&~m[1995]&m[1997]&m[1998])|(m[1993]&~m[1994]&m[1995]&m[1997]&m[1998])|(~m[1993]&m[1994]&m[1995]&m[1997]&m[1998]))&UnbiasedRNG[926])|((m[1993]&m[1994]&~m[1995]&~m[1997]&~m[1998])|(m[1993]&~m[1994]&m[1995]&~m[1997]&~m[1998])|(~m[1993]&m[1994]&m[1995]&~m[1997]&~m[1998])|(m[1993]&m[1994]&m[1995]&~m[1997]&~m[1998])|(m[1993]&~m[1994]&~m[1995]&~m[1997]&m[1998])|(~m[1993]&m[1994]&~m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&~m[1995]&~m[1997]&m[1998])|(~m[1993]&~m[1994]&m[1995]&~m[1997]&m[1998])|(m[1993]&~m[1994]&m[1995]&~m[1997]&m[1998])|(~m[1993]&m[1994]&m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&m[1995]&~m[1997]&m[1998])|(m[1993]&m[1994]&m[1995]&m[1997]&m[1998]))):InitCond[1821];
    m[2001] = run?((((m[1998]&~m[1999]&~m[2000]&~m[2002]&~m[2003])|(~m[1998]&m[1999]&~m[2000]&~m[2002]&~m[2003])|(~m[1998]&~m[1999]&m[2000]&~m[2002]&~m[2003])|(m[1998]&m[1999]&m[2000]&m[2002]&~m[2003])|(~m[1998]&~m[1999]&~m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&~m[2000]&m[2002]&m[2003])|(m[1998]&~m[1999]&m[2000]&m[2002]&m[2003])|(~m[1998]&m[1999]&m[2000]&m[2002]&m[2003]))&UnbiasedRNG[927])|((m[1998]&m[1999]&~m[2000]&~m[2002]&~m[2003])|(m[1998]&~m[1999]&m[2000]&~m[2002]&~m[2003])|(~m[1998]&m[1999]&m[2000]&~m[2002]&~m[2003])|(m[1998]&m[1999]&m[2000]&~m[2002]&~m[2003])|(m[1998]&~m[1999]&~m[2000]&~m[2002]&m[2003])|(~m[1998]&m[1999]&~m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&~m[2000]&~m[2002]&m[2003])|(~m[1998]&~m[1999]&m[2000]&~m[2002]&m[2003])|(m[1998]&~m[1999]&m[2000]&~m[2002]&m[2003])|(~m[1998]&m[1999]&m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&m[2000]&~m[2002]&m[2003])|(m[1998]&m[1999]&m[2000]&m[2002]&m[2003]))):InitCond[1822];
    m[2006] = run?((((m[2003]&~m[2004]&~m[2005]&~m[2007]&~m[2008])|(~m[2003]&m[2004]&~m[2005]&~m[2007]&~m[2008])|(~m[2003]&~m[2004]&m[2005]&~m[2007]&~m[2008])|(m[2003]&m[2004]&m[2005]&m[2007]&~m[2008])|(~m[2003]&~m[2004]&~m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&~m[2005]&m[2007]&m[2008])|(m[2003]&~m[2004]&m[2005]&m[2007]&m[2008])|(~m[2003]&m[2004]&m[2005]&m[2007]&m[2008]))&UnbiasedRNG[928])|((m[2003]&m[2004]&~m[2005]&~m[2007]&~m[2008])|(m[2003]&~m[2004]&m[2005]&~m[2007]&~m[2008])|(~m[2003]&m[2004]&m[2005]&~m[2007]&~m[2008])|(m[2003]&m[2004]&m[2005]&~m[2007]&~m[2008])|(m[2003]&~m[2004]&~m[2005]&~m[2007]&m[2008])|(~m[2003]&m[2004]&~m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&~m[2005]&~m[2007]&m[2008])|(~m[2003]&~m[2004]&m[2005]&~m[2007]&m[2008])|(m[2003]&~m[2004]&m[2005]&~m[2007]&m[2008])|(~m[2003]&m[2004]&m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&m[2005]&~m[2007]&m[2008])|(m[2003]&m[2004]&m[2005]&m[2007]&m[2008]))):InitCond[1823];
    m[2011] = run?((((m[2008]&~m[2009]&~m[2010]&~m[2012]&~m[2013])|(~m[2008]&m[2009]&~m[2010]&~m[2012]&~m[2013])|(~m[2008]&~m[2009]&m[2010]&~m[2012]&~m[2013])|(m[2008]&m[2009]&m[2010]&m[2012]&~m[2013])|(~m[2008]&~m[2009]&~m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&~m[2010]&m[2012]&m[2013])|(m[2008]&~m[2009]&m[2010]&m[2012]&m[2013])|(~m[2008]&m[2009]&m[2010]&m[2012]&m[2013]))&UnbiasedRNG[929])|((m[2008]&m[2009]&~m[2010]&~m[2012]&~m[2013])|(m[2008]&~m[2009]&m[2010]&~m[2012]&~m[2013])|(~m[2008]&m[2009]&m[2010]&~m[2012]&~m[2013])|(m[2008]&m[2009]&m[2010]&~m[2012]&~m[2013])|(m[2008]&~m[2009]&~m[2010]&~m[2012]&m[2013])|(~m[2008]&m[2009]&~m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&~m[2010]&~m[2012]&m[2013])|(~m[2008]&~m[2009]&m[2010]&~m[2012]&m[2013])|(m[2008]&~m[2009]&m[2010]&~m[2012]&m[2013])|(~m[2008]&m[2009]&m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&m[2010]&~m[2012]&m[2013])|(m[2008]&m[2009]&m[2010]&m[2012]&m[2013]))):InitCond[1824];
    m[2016] = run?((((m[2013]&~m[2014]&~m[2015]&~m[2017]&~m[2018])|(~m[2013]&m[2014]&~m[2015]&~m[2017]&~m[2018])|(~m[2013]&~m[2014]&m[2015]&~m[2017]&~m[2018])|(m[2013]&m[2014]&m[2015]&m[2017]&~m[2018])|(~m[2013]&~m[2014]&~m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&~m[2015]&m[2017]&m[2018])|(m[2013]&~m[2014]&m[2015]&m[2017]&m[2018])|(~m[2013]&m[2014]&m[2015]&m[2017]&m[2018]))&UnbiasedRNG[930])|((m[2013]&m[2014]&~m[2015]&~m[2017]&~m[2018])|(m[2013]&~m[2014]&m[2015]&~m[2017]&~m[2018])|(~m[2013]&m[2014]&m[2015]&~m[2017]&~m[2018])|(m[2013]&m[2014]&m[2015]&~m[2017]&~m[2018])|(m[2013]&~m[2014]&~m[2015]&~m[2017]&m[2018])|(~m[2013]&m[2014]&~m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&~m[2015]&~m[2017]&m[2018])|(~m[2013]&~m[2014]&m[2015]&~m[2017]&m[2018])|(m[2013]&~m[2014]&m[2015]&~m[2017]&m[2018])|(~m[2013]&m[2014]&m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&m[2015]&~m[2017]&m[2018])|(m[2013]&m[2014]&m[2015]&m[2017]&m[2018]))):InitCond[1825];
    m[2026] = run?((((m[2023]&~m[2024]&~m[2025]&~m[2027]&~m[2028])|(~m[2023]&m[2024]&~m[2025]&~m[2027]&~m[2028])|(~m[2023]&~m[2024]&m[2025]&~m[2027]&~m[2028])|(m[2023]&m[2024]&m[2025]&m[2027]&~m[2028])|(~m[2023]&~m[2024]&~m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&~m[2025]&m[2027]&m[2028])|(m[2023]&~m[2024]&m[2025]&m[2027]&m[2028])|(~m[2023]&m[2024]&m[2025]&m[2027]&m[2028]))&UnbiasedRNG[931])|((m[2023]&m[2024]&~m[2025]&~m[2027]&~m[2028])|(m[2023]&~m[2024]&m[2025]&~m[2027]&~m[2028])|(~m[2023]&m[2024]&m[2025]&~m[2027]&~m[2028])|(m[2023]&m[2024]&m[2025]&~m[2027]&~m[2028])|(m[2023]&~m[2024]&~m[2025]&~m[2027]&m[2028])|(~m[2023]&m[2024]&~m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&~m[2025]&~m[2027]&m[2028])|(~m[2023]&~m[2024]&m[2025]&~m[2027]&m[2028])|(m[2023]&~m[2024]&m[2025]&~m[2027]&m[2028])|(~m[2023]&m[2024]&m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&m[2025]&~m[2027]&m[2028])|(m[2023]&m[2024]&m[2025]&m[2027]&m[2028]))):InitCond[1826];
    m[2031] = run?((((m[2028]&~m[2029]&~m[2030]&~m[2032]&~m[2033])|(~m[2028]&m[2029]&~m[2030]&~m[2032]&~m[2033])|(~m[2028]&~m[2029]&m[2030]&~m[2032]&~m[2033])|(m[2028]&m[2029]&m[2030]&m[2032]&~m[2033])|(~m[2028]&~m[2029]&~m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&~m[2030]&m[2032]&m[2033])|(m[2028]&~m[2029]&m[2030]&m[2032]&m[2033])|(~m[2028]&m[2029]&m[2030]&m[2032]&m[2033]))&UnbiasedRNG[932])|((m[2028]&m[2029]&~m[2030]&~m[2032]&~m[2033])|(m[2028]&~m[2029]&m[2030]&~m[2032]&~m[2033])|(~m[2028]&m[2029]&m[2030]&~m[2032]&~m[2033])|(m[2028]&m[2029]&m[2030]&~m[2032]&~m[2033])|(m[2028]&~m[2029]&~m[2030]&~m[2032]&m[2033])|(~m[2028]&m[2029]&~m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&~m[2030]&~m[2032]&m[2033])|(~m[2028]&~m[2029]&m[2030]&~m[2032]&m[2033])|(m[2028]&~m[2029]&m[2030]&~m[2032]&m[2033])|(~m[2028]&m[2029]&m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&m[2030]&~m[2032]&m[2033])|(m[2028]&m[2029]&m[2030]&m[2032]&m[2033]))):InitCond[1827];
    m[2036] = run?((((m[2033]&~m[2034]&~m[2035]&~m[2037]&~m[2038])|(~m[2033]&m[2034]&~m[2035]&~m[2037]&~m[2038])|(~m[2033]&~m[2034]&m[2035]&~m[2037]&~m[2038])|(m[2033]&m[2034]&m[2035]&m[2037]&~m[2038])|(~m[2033]&~m[2034]&~m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&~m[2035]&m[2037]&m[2038])|(m[2033]&~m[2034]&m[2035]&m[2037]&m[2038])|(~m[2033]&m[2034]&m[2035]&m[2037]&m[2038]))&UnbiasedRNG[933])|((m[2033]&m[2034]&~m[2035]&~m[2037]&~m[2038])|(m[2033]&~m[2034]&m[2035]&~m[2037]&~m[2038])|(~m[2033]&m[2034]&m[2035]&~m[2037]&~m[2038])|(m[2033]&m[2034]&m[2035]&~m[2037]&~m[2038])|(m[2033]&~m[2034]&~m[2035]&~m[2037]&m[2038])|(~m[2033]&m[2034]&~m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&~m[2035]&~m[2037]&m[2038])|(~m[2033]&~m[2034]&m[2035]&~m[2037]&m[2038])|(m[2033]&~m[2034]&m[2035]&~m[2037]&m[2038])|(~m[2033]&m[2034]&m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&m[2035]&~m[2037]&m[2038])|(m[2033]&m[2034]&m[2035]&m[2037]&m[2038]))):InitCond[1828];
    m[2041] = run?((((m[2038]&~m[2039]&~m[2040]&~m[2042]&~m[2043])|(~m[2038]&m[2039]&~m[2040]&~m[2042]&~m[2043])|(~m[2038]&~m[2039]&m[2040]&~m[2042]&~m[2043])|(m[2038]&m[2039]&m[2040]&m[2042]&~m[2043])|(~m[2038]&~m[2039]&~m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&~m[2040]&m[2042]&m[2043])|(m[2038]&~m[2039]&m[2040]&m[2042]&m[2043])|(~m[2038]&m[2039]&m[2040]&m[2042]&m[2043]))&UnbiasedRNG[934])|((m[2038]&m[2039]&~m[2040]&~m[2042]&~m[2043])|(m[2038]&~m[2039]&m[2040]&~m[2042]&~m[2043])|(~m[2038]&m[2039]&m[2040]&~m[2042]&~m[2043])|(m[2038]&m[2039]&m[2040]&~m[2042]&~m[2043])|(m[2038]&~m[2039]&~m[2040]&~m[2042]&m[2043])|(~m[2038]&m[2039]&~m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&~m[2040]&~m[2042]&m[2043])|(~m[2038]&~m[2039]&m[2040]&~m[2042]&m[2043])|(m[2038]&~m[2039]&m[2040]&~m[2042]&m[2043])|(~m[2038]&m[2039]&m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&m[2040]&~m[2042]&m[2043])|(m[2038]&m[2039]&m[2040]&m[2042]&m[2043]))):InitCond[1829];
    m[2046] = run?((((m[2043]&~m[2044]&~m[2045]&~m[2047]&~m[2048])|(~m[2043]&m[2044]&~m[2045]&~m[2047]&~m[2048])|(~m[2043]&~m[2044]&m[2045]&~m[2047]&~m[2048])|(m[2043]&m[2044]&m[2045]&m[2047]&~m[2048])|(~m[2043]&~m[2044]&~m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&~m[2045]&m[2047]&m[2048])|(m[2043]&~m[2044]&m[2045]&m[2047]&m[2048])|(~m[2043]&m[2044]&m[2045]&m[2047]&m[2048]))&UnbiasedRNG[935])|((m[2043]&m[2044]&~m[2045]&~m[2047]&~m[2048])|(m[2043]&~m[2044]&m[2045]&~m[2047]&~m[2048])|(~m[2043]&m[2044]&m[2045]&~m[2047]&~m[2048])|(m[2043]&m[2044]&m[2045]&~m[2047]&~m[2048])|(m[2043]&~m[2044]&~m[2045]&~m[2047]&m[2048])|(~m[2043]&m[2044]&~m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&~m[2045]&~m[2047]&m[2048])|(~m[2043]&~m[2044]&m[2045]&~m[2047]&m[2048])|(m[2043]&~m[2044]&m[2045]&~m[2047]&m[2048])|(~m[2043]&m[2044]&m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&m[2045]&~m[2047]&m[2048])|(m[2043]&m[2044]&m[2045]&m[2047]&m[2048]))):InitCond[1830];
    m[2056] = run?((((m[2053]&~m[2054]&~m[2055]&~m[2057]&~m[2058])|(~m[2053]&m[2054]&~m[2055]&~m[2057]&~m[2058])|(~m[2053]&~m[2054]&m[2055]&~m[2057]&~m[2058])|(m[2053]&m[2054]&m[2055]&m[2057]&~m[2058])|(~m[2053]&~m[2054]&~m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&~m[2055]&m[2057]&m[2058])|(m[2053]&~m[2054]&m[2055]&m[2057]&m[2058])|(~m[2053]&m[2054]&m[2055]&m[2057]&m[2058]))&UnbiasedRNG[936])|((m[2053]&m[2054]&~m[2055]&~m[2057]&~m[2058])|(m[2053]&~m[2054]&m[2055]&~m[2057]&~m[2058])|(~m[2053]&m[2054]&m[2055]&~m[2057]&~m[2058])|(m[2053]&m[2054]&m[2055]&~m[2057]&~m[2058])|(m[2053]&~m[2054]&~m[2055]&~m[2057]&m[2058])|(~m[2053]&m[2054]&~m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&~m[2055]&~m[2057]&m[2058])|(~m[2053]&~m[2054]&m[2055]&~m[2057]&m[2058])|(m[2053]&~m[2054]&m[2055]&~m[2057]&m[2058])|(~m[2053]&m[2054]&m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&m[2055]&~m[2057]&m[2058])|(m[2053]&m[2054]&m[2055]&m[2057]&m[2058]))):InitCond[1831];
    m[2061] = run?((((m[2058]&~m[2059]&~m[2060]&~m[2062]&~m[2063])|(~m[2058]&m[2059]&~m[2060]&~m[2062]&~m[2063])|(~m[2058]&~m[2059]&m[2060]&~m[2062]&~m[2063])|(m[2058]&m[2059]&m[2060]&m[2062]&~m[2063])|(~m[2058]&~m[2059]&~m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&~m[2060]&m[2062]&m[2063])|(m[2058]&~m[2059]&m[2060]&m[2062]&m[2063])|(~m[2058]&m[2059]&m[2060]&m[2062]&m[2063]))&UnbiasedRNG[937])|((m[2058]&m[2059]&~m[2060]&~m[2062]&~m[2063])|(m[2058]&~m[2059]&m[2060]&~m[2062]&~m[2063])|(~m[2058]&m[2059]&m[2060]&~m[2062]&~m[2063])|(m[2058]&m[2059]&m[2060]&~m[2062]&~m[2063])|(m[2058]&~m[2059]&~m[2060]&~m[2062]&m[2063])|(~m[2058]&m[2059]&~m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&~m[2060]&~m[2062]&m[2063])|(~m[2058]&~m[2059]&m[2060]&~m[2062]&m[2063])|(m[2058]&~m[2059]&m[2060]&~m[2062]&m[2063])|(~m[2058]&m[2059]&m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&m[2060]&~m[2062]&m[2063])|(m[2058]&m[2059]&m[2060]&m[2062]&m[2063]))):InitCond[1832];
    m[2066] = run?((((m[2063]&~m[2064]&~m[2065]&~m[2067]&~m[2068])|(~m[2063]&m[2064]&~m[2065]&~m[2067]&~m[2068])|(~m[2063]&~m[2064]&m[2065]&~m[2067]&~m[2068])|(m[2063]&m[2064]&m[2065]&m[2067]&~m[2068])|(~m[2063]&~m[2064]&~m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&~m[2065]&m[2067]&m[2068])|(m[2063]&~m[2064]&m[2065]&m[2067]&m[2068])|(~m[2063]&m[2064]&m[2065]&m[2067]&m[2068]))&UnbiasedRNG[938])|((m[2063]&m[2064]&~m[2065]&~m[2067]&~m[2068])|(m[2063]&~m[2064]&m[2065]&~m[2067]&~m[2068])|(~m[2063]&m[2064]&m[2065]&~m[2067]&~m[2068])|(m[2063]&m[2064]&m[2065]&~m[2067]&~m[2068])|(m[2063]&~m[2064]&~m[2065]&~m[2067]&m[2068])|(~m[2063]&m[2064]&~m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&~m[2065]&~m[2067]&m[2068])|(~m[2063]&~m[2064]&m[2065]&~m[2067]&m[2068])|(m[2063]&~m[2064]&m[2065]&~m[2067]&m[2068])|(~m[2063]&m[2064]&m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&m[2065]&~m[2067]&m[2068])|(m[2063]&m[2064]&m[2065]&m[2067]&m[2068]))):InitCond[1833];
    m[2071] = run?((((m[2068]&~m[2069]&~m[2070]&~m[2072]&~m[2073])|(~m[2068]&m[2069]&~m[2070]&~m[2072]&~m[2073])|(~m[2068]&~m[2069]&m[2070]&~m[2072]&~m[2073])|(m[2068]&m[2069]&m[2070]&m[2072]&~m[2073])|(~m[2068]&~m[2069]&~m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&~m[2070]&m[2072]&m[2073])|(m[2068]&~m[2069]&m[2070]&m[2072]&m[2073])|(~m[2068]&m[2069]&m[2070]&m[2072]&m[2073]))&UnbiasedRNG[939])|((m[2068]&m[2069]&~m[2070]&~m[2072]&~m[2073])|(m[2068]&~m[2069]&m[2070]&~m[2072]&~m[2073])|(~m[2068]&m[2069]&m[2070]&~m[2072]&~m[2073])|(m[2068]&m[2069]&m[2070]&~m[2072]&~m[2073])|(m[2068]&~m[2069]&~m[2070]&~m[2072]&m[2073])|(~m[2068]&m[2069]&~m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&~m[2070]&~m[2072]&m[2073])|(~m[2068]&~m[2069]&m[2070]&~m[2072]&m[2073])|(m[2068]&~m[2069]&m[2070]&~m[2072]&m[2073])|(~m[2068]&m[2069]&m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&m[2070]&~m[2072]&m[2073])|(m[2068]&m[2069]&m[2070]&m[2072]&m[2073]))):InitCond[1834];
    m[2081] = run?((((m[2078]&~m[2079]&~m[2080]&~m[2082]&~m[2083])|(~m[2078]&m[2079]&~m[2080]&~m[2082]&~m[2083])|(~m[2078]&~m[2079]&m[2080]&~m[2082]&~m[2083])|(m[2078]&m[2079]&m[2080]&m[2082]&~m[2083])|(~m[2078]&~m[2079]&~m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&~m[2080]&m[2082]&m[2083])|(m[2078]&~m[2079]&m[2080]&m[2082]&m[2083])|(~m[2078]&m[2079]&m[2080]&m[2082]&m[2083]))&UnbiasedRNG[940])|((m[2078]&m[2079]&~m[2080]&~m[2082]&~m[2083])|(m[2078]&~m[2079]&m[2080]&~m[2082]&~m[2083])|(~m[2078]&m[2079]&m[2080]&~m[2082]&~m[2083])|(m[2078]&m[2079]&m[2080]&~m[2082]&~m[2083])|(m[2078]&~m[2079]&~m[2080]&~m[2082]&m[2083])|(~m[2078]&m[2079]&~m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&~m[2080]&~m[2082]&m[2083])|(~m[2078]&~m[2079]&m[2080]&~m[2082]&m[2083])|(m[2078]&~m[2079]&m[2080]&~m[2082]&m[2083])|(~m[2078]&m[2079]&m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&m[2080]&~m[2082]&m[2083])|(m[2078]&m[2079]&m[2080]&m[2082]&m[2083]))):InitCond[1835];
    m[2086] = run?((((m[2083]&~m[2084]&~m[2085]&~m[2087]&~m[2088])|(~m[2083]&m[2084]&~m[2085]&~m[2087]&~m[2088])|(~m[2083]&~m[2084]&m[2085]&~m[2087]&~m[2088])|(m[2083]&m[2084]&m[2085]&m[2087]&~m[2088])|(~m[2083]&~m[2084]&~m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&~m[2085]&m[2087]&m[2088])|(m[2083]&~m[2084]&m[2085]&m[2087]&m[2088])|(~m[2083]&m[2084]&m[2085]&m[2087]&m[2088]))&UnbiasedRNG[941])|((m[2083]&m[2084]&~m[2085]&~m[2087]&~m[2088])|(m[2083]&~m[2084]&m[2085]&~m[2087]&~m[2088])|(~m[2083]&m[2084]&m[2085]&~m[2087]&~m[2088])|(m[2083]&m[2084]&m[2085]&~m[2087]&~m[2088])|(m[2083]&~m[2084]&~m[2085]&~m[2087]&m[2088])|(~m[2083]&m[2084]&~m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&~m[2085]&~m[2087]&m[2088])|(~m[2083]&~m[2084]&m[2085]&~m[2087]&m[2088])|(m[2083]&~m[2084]&m[2085]&~m[2087]&m[2088])|(~m[2083]&m[2084]&m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&m[2085]&~m[2087]&m[2088])|(m[2083]&m[2084]&m[2085]&m[2087]&m[2088]))):InitCond[1836];
    m[2091] = run?((((m[2088]&~m[2089]&~m[2090]&~m[2092]&~m[2093])|(~m[2088]&m[2089]&~m[2090]&~m[2092]&~m[2093])|(~m[2088]&~m[2089]&m[2090]&~m[2092]&~m[2093])|(m[2088]&m[2089]&m[2090]&m[2092]&~m[2093])|(~m[2088]&~m[2089]&~m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&~m[2090]&m[2092]&m[2093])|(m[2088]&~m[2089]&m[2090]&m[2092]&m[2093])|(~m[2088]&m[2089]&m[2090]&m[2092]&m[2093]))&UnbiasedRNG[942])|((m[2088]&m[2089]&~m[2090]&~m[2092]&~m[2093])|(m[2088]&~m[2089]&m[2090]&~m[2092]&~m[2093])|(~m[2088]&m[2089]&m[2090]&~m[2092]&~m[2093])|(m[2088]&m[2089]&m[2090]&~m[2092]&~m[2093])|(m[2088]&~m[2089]&~m[2090]&~m[2092]&m[2093])|(~m[2088]&m[2089]&~m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&~m[2090]&~m[2092]&m[2093])|(~m[2088]&~m[2089]&m[2090]&~m[2092]&m[2093])|(m[2088]&~m[2089]&m[2090]&~m[2092]&m[2093])|(~m[2088]&m[2089]&m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&m[2090]&~m[2092]&m[2093])|(m[2088]&m[2089]&m[2090]&m[2092]&m[2093]))):InitCond[1837];
    m[2101] = run?((((m[2098]&~m[2099]&~m[2100]&~m[2102]&~m[2103])|(~m[2098]&m[2099]&~m[2100]&~m[2102]&~m[2103])|(~m[2098]&~m[2099]&m[2100]&~m[2102]&~m[2103])|(m[2098]&m[2099]&m[2100]&m[2102]&~m[2103])|(~m[2098]&~m[2099]&~m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&~m[2100]&m[2102]&m[2103])|(m[2098]&~m[2099]&m[2100]&m[2102]&m[2103])|(~m[2098]&m[2099]&m[2100]&m[2102]&m[2103]))&UnbiasedRNG[943])|((m[2098]&m[2099]&~m[2100]&~m[2102]&~m[2103])|(m[2098]&~m[2099]&m[2100]&~m[2102]&~m[2103])|(~m[2098]&m[2099]&m[2100]&~m[2102]&~m[2103])|(m[2098]&m[2099]&m[2100]&~m[2102]&~m[2103])|(m[2098]&~m[2099]&~m[2100]&~m[2102]&m[2103])|(~m[2098]&m[2099]&~m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&~m[2100]&~m[2102]&m[2103])|(~m[2098]&~m[2099]&m[2100]&~m[2102]&m[2103])|(m[2098]&~m[2099]&m[2100]&~m[2102]&m[2103])|(~m[2098]&m[2099]&m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&m[2100]&~m[2102]&m[2103])|(m[2098]&m[2099]&m[2100]&m[2102]&m[2103]))):InitCond[1838];
    m[2106] = run?((((m[2103]&~m[2104]&~m[2105]&~m[2107]&~m[2108])|(~m[2103]&m[2104]&~m[2105]&~m[2107]&~m[2108])|(~m[2103]&~m[2104]&m[2105]&~m[2107]&~m[2108])|(m[2103]&m[2104]&m[2105]&m[2107]&~m[2108])|(~m[2103]&~m[2104]&~m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&~m[2105]&m[2107]&m[2108])|(m[2103]&~m[2104]&m[2105]&m[2107]&m[2108])|(~m[2103]&m[2104]&m[2105]&m[2107]&m[2108]))&UnbiasedRNG[944])|((m[2103]&m[2104]&~m[2105]&~m[2107]&~m[2108])|(m[2103]&~m[2104]&m[2105]&~m[2107]&~m[2108])|(~m[2103]&m[2104]&m[2105]&~m[2107]&~m[2108])|(m[2103]&m[2104]&m[2105]&~m[2107]&~m[2108])|(m[2103]&~m[2104]&~m[2105]&~m[2107]&m[2108])|(~m[2103]&m[2104]&~m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&~m[2105]&~m[2107]&m[2108])|(~m[2103]&~m[2104]&m[2105]&~m[2107]&m[2108])|(m[2103]&~m[2104]&m[2105]&~m[2107]&m[2108])|(~m[2103]&m[2104]&m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&m[2105]&~m[2107]&m[2108])|(m[2103]&m[2104]&m[2105]&m[2107]&m[2108]))):InitCond[1839];
    m[2116] = run?((((m[2113]&~m[2114]&~m[2115]&~m[2117]&~m[2118])|(~m[2113]&m[2114]&~m[2115]&~m[2117]&~m[2118])|(~m[2113]&~m[2114]&m[2115]&~m[2117]&~m[2118])|(m[2113]&m[2114]&m[2115]&m[2117]&~m[2118])|(~m[2113]&~m[2114]&~m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&~m[2115]&m[2117]&m[2118])|(m[2113]&~m[2114]&m[2115]&m[2117]&m[2118])|(~m[2113]&m[2114]&m[2115]&m[2117]&m[2118]))&UnbiasedRNG[945])|((m[2113]&m[2114]&~m[2115]&~m[2117]&~m[2118])|(m[2113]&~m[2114]&m[2115]&~m[2117]&~m[2118])|(~m[2113]&m[2114]&m[2115]&~m[2117]&~m[2118])|(m[2113]&m[2114]&m[2115]&~m[2117]&~m[2118])|(m[2113]&~m[2114]&~m[2115]&~m[2117]&m[2118])|(~m[2113]&m[2114]&~m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&~m[2115]&~m[2117]&m[2118])|(~m[2113]&~m[2114]&m[2115]&~m[2117]&m[2118])|(m[2113]&~m[2114]&m[2115]&~m[2117]&m[2118])|(~m[2113]&m[2114]&m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&m[2115]&~m[2117]&m[2118])|(m[2113]&m[2114]&m[2115]&m[2117]&m[2118]))):InitCond[1840];
end

always @(posedge color4_clk) begin
    m[932] = run?((((m[928]&~m[929]&~m[930]&~m[931]&~m[935])|(~m[928]&m[929]&~m[930]&~m[931]&~m[935])|(~m[928]&~m[929]&m[930]&~m[931]&~m[935])|(m[928]&m[929]&~m[930]&m[931]&~m[935])|(m[928]&~m[929]&m[930]&m[931]&~m[935])|(~m[928]&m[929]&m[930]&m[931]&~m[935]))&BiasedRNG[895])|(((m[928]&~m[929]&~m[930]&~m[931]&m[935])|(~m[928]&m[929]&~m[930]&~m[931]&m[935])|(~m[928]&~m[929]&m[930]&~m[931]&m[935])|(m[928]&m[929]&~m[930]&m[931]&m[935])|(m[928]&~m[929]&m[930]&m[931]&m[935])|(~m[928]&m[929]&m[930]&m[931]&m[935]))&~BiasedRNG[895])|((m[928]&m[929]&~m[930]&~m[931]&~m[935])|(m[928]&~m[929]&m[930]&~m[931]&~m[935])|(~m[928]&m[929]&m[930]&~m[931]&~m[935])|(m[928]&m[929]&m[930]&~m[931]&~m[935])|(m[928]&m[929]&m[930]&m[931]&~m[935])|(m[928]&m[929]&~m[930]&~m[931]&m[935])|(m[928]&~m[929]&m[930]&~m[931]&m[935])|(~m[928]&m[929]&m[930]&~m[931]&m[935])|(m[928]&m[929]&m[930]&~m[931]&m[935])|(m[928]&m[929]&m[930]&m[931]&m[935]))):InitCond[1841];
    m[937] = run?((((m[933]&~m[934]&~m[935]&~m[936]&~m[945])|(~m[933]&m[934]&~m[935]&~m[936]&~m[945])|(~m[933]&~m[934]&m[935]&~m[936]&~m[945])|(m[933]&m[934]&~m[935]&m[936]&~m[945])|(m[933]&~m[934]&m[935]&m[936]&~m[945])|(~m[933]&m[934]&m[935]&m[936]&~m[945]))&BiasedRNG[896])|(((m[933]&~m[934]&~m[935]&~m[936]&m[945])|(~m[933]&m[934]&~m[935]&~m[936]&m[945])|(~m[933]&~m[934]&m[935]&~m[936]&m[945])|(m[933]&m[934]&~m[935]&m[936]&m[945])|(m[933]&~m[934]&m[935]&m[936]&m[945])|(~m[933]&m[934]&m[935]&m[936]&m[945]))&~BiasedRNG[896])|((m[933]&m[934]&~m[935]&~m[936]&~m[945])|(m[933]&~m[934]&m[935]&~m[936]&~m[945])|(~m[933]&m[934]&m[935]&~m[936]&~m[945])|(m[933]&m[934]&m[935]&~m[936]&~m[945])|(m[933]&m[934]&m[935]&m[936]&~m[945])|(m[933]&m[934]&~m[935]&~m[936]&m[945])|(m[933]&~m[934]&m[935]&~m[936]&m[945])|(~m[933]&m[934]&m[935]&~m[936]&m[945])|(m[933]&m[934]&m[935]&~m[936]&m[945])|(m[933]&m[934]&m[935]&m[936]&m[945]))):InitCond[1842];
    m[942] = run?((((m[938]&~m[939]&~m[940]&~m[941]&~m[950])|(~m[938]&m[939]&~m[940]&~m[941]&~m[950])|(~m[938]&~m[939]&m[940]&~m[941]&~m[950])|(m[938]&m[939]&~m[940]&m[941]&~m[950])|(m[938]&~m[939]&m[940]&m[941]&~m[950])|(~m[938]&m[939]&m[940]&m[941]&~m[950]))&BiasedRNG[897])|(((m[938]&~m[939]&~m[940]&~m[941]&m[950])|(~m[938]&m[939]&~m[940]&~m[941]&m[950])|(~m[938]&~m[939]&m[940]&~m[941]&m[950])|(m[938]&m[939]&~m[940]&m[941]&m[950])|(m[938]&~m[939]&m[940]&m[941]&m[950])|(~m[938]&m[939]&m[940]&m[941]&m[950]))&~BiasedRNG[897])|((m[938]&m[939]&~m[940]&~m[941]&~m[950])|(m[938]&~m[939]&m[940]&~m[941]&~m[950])|(~m[938]&m[939]&m[940]&~m[941]&~m[950])|(m[938]&m[939]&m[940]&~m[941]&~m[950])|(m[938]&m[939]&m[940]&m[941]&~m[950])|(m[938]&m[939]&~m[940]&~m[941]&m[950])|(m[938]&~m[939]&m[940]&~m[941]&m[950])|(~m[938]&m[939]&m[940]&~m[941]&m[950])|(m[938]&m[939]&m[940]&~m[941]&m[950])|(m[938]&m[939]&m[940]&m[941]&m[950]))):InitCond[1843];
    m[947] = run?((((m[943]&~m[944]&~m[945]&~m[946]&~m[960])|(~m[943]&m[944]&~m[945]&~m[946]&~m[960])|(~m[943]&~m[944]&m[945]&~m[946]&~m[960])|(m[943]&m[944]&~m[945]&m[946]&~m[960])|(m[943]&~m[944]&m[945]&m[946]&~m[960])|(~m[943]&m[944]&m[945]&m[946]&~m[960]))&BiasedRNG[898])|(((m[943]&~m[944]&~m[945]&~m[946]&m[960])|(~m[943]&m[944]&~m[945]&~m[946]&m[960])|(~m[943]&~m[944]&m[945]&~m[946]&m[960])|(m[943]&m[944]&~m[945]&m[946]&m[960])|(m[943]&~m[944]&m[945]&m[946]&m[960])|(~m[943]&m[944]&m[945]&m[946]&m[960]))&~BiasedRNG[898])|((m[943]&m[944]&~m[945]&~m[946]&~m[960])|(m[943]&~m[944]&m[945]&~m[946]&~m[960])|(~m[943]&m[944]&m[945]&~m[946]&~m[960])|(m[943]&m[944]&m[945]&~m[946]&~m[960])|(m[943]&m[944]&m[945]&m[946]&~m[960])|(m[943]&m[944]&~m[945]&~m[946]&m[960])|(m[943]&~m[944]&m[945]&~m[946]&m[960])|(~m[943]&m[944]&m[945]&~m[946]&m[960])|(m[943]&m[944]&m[945]&~m[946]&m[960])|(m[943]&m[944]&m[945]&m[946]&m[960]))):InitCond[1844];
    m[952] = run?((((m[948]&~m[949]&~m[950]&~m[951]&~m[965])|(~m[948]&m[949]&~m[950]&~m[951]&~m[965])|(~m[948]&~m[949]&m[950]&~m[951]&~m[965])|(m[948]&m[949]&~m[950]&m[951]&~m[965])|(m[948]&~m[949]&m[950]&m[951]&~m[965])|(~m[948]&m[949]&m[950]&m[951]&~m[965]))&BiasedRNG[899])|(((m[948]&~m[949]&~m[950]&~m[951]&m[965])|(~m[948]&m[949]&~m[950]&~m[951]&m[965])|(~m[948]&~m[949]&m[950]&~m[951]&m[965])|(m[948]&m[949]&~m[950]&m[951]&m[965])|(m[948]&~m[949]&m[950]&m[951]&m[965])|(~m[948]&m[949]&m[950]&m[951]&m[965]))&~BiasedRNG[899])|((m[948]&m[949]&~m[950]&~m[951]&~m[965])|(m[948]&~m[949]&m[950]&~m[951]&~m[965])|(~m[948]&m[949]&m[950]&~m[951]&~m[965])|(m[948]&m[949]&m[950]&~m[951]&~m[965])|(m[948]&m[949]&m[950]&m[951]&~m[965])|(m[948]&m[949]&~m[950]&~m[951]&m[965])|(m[948]&~m[949]&m[950]&~m[951]&m[965])|(~m[948]&m[949]&m[950]&~m[951]&m[965])|(m[948]&m[949]&m[950]&~m[951]&m[965])|(m[948]&m[949]&m[950]&m[951]&m[965]))):InitCond[1845];
    m[957] = run?((((m[953]&~m[954]&~m[955]&~m[956]&~m[970])|(~m[953]&m[954]&~m[955]&~m[956]&~m[970])|(~m[953]&~m[954]&m[955]&~m[956]&~m[970])|(m[953]&m[954]&~m[955]&m[956]&~m[970])|(m[953]&~m[954]&m[955]&m[956]&~m[970])|(~m[953]&m[954]&m[955]&m[956]&~m[970]))&BiasedRNG[900])|(((m[953]&~m[954]&~m[955]&~m[956]&m[970])|(~m[953]&m[954]&~m[955]&~m[956]&m[970])|(~m[953]&~m[954]&m[955]&~m[956]&m[970])|(m[953]&m[954]&~m[955]&m[956]&m[970])|(m[953]&~m[954]&m[955]&m[956]&m[970])|(~m[953]&m[954]&m[955]&m[956]&m[970]))&~BiasedRNG[900])|((m[953]&m[954]&~m[955]&~m[956]&~m[970])|(m[953]&~m[954]&m[955]&~m[956]&~m[970])|(~m[953]&m[954]&m[955]&~m[956]&~m[970])|(m[953]&m[954]&m[955]&~m[956]&~m[970])|(m[953]&m[954]&m[955]&m[956]&~m[970])|(m[953]&m[954]&~m[955]&~m[956]&m[970])|(m[953]&~m[954]&m[955]&~m[956]&m[970])|(~m[953]&m[954]&m[955]&~m[956]&m[970])|(m[953]&m[954]&m[955]&~m[956]&m[970])|(m[953]&m[954]&m[955]&m[956]&m[970]))):InitCond[1846];
    m[962] = run?((((m[958]&~m[959]&~m[960]&~m[961]&~m[980])|(~m[958]&m[959]&~m[960]&~m[961]&~m[980])|(~m[958]&~m[959]&m[960]&~m[961]&~m[980])|(m[958]&m[959]&~m[960]&m[961]&~m[980])|(m[958]&~m[959]&m[960]&m[961]&~m[980])|(~m[958]&m[959]&m[960]&m[961]&~m[980]))&BiasedRNG[901])|(((m[958]&~m[959]&~m[960]&~m[961]&m[980])|(~m[958]&m[959]&~m[960]&~m[961]&m[980])|(~m[958]&~m[959]&m[960]&~m[961]&m[980])|(m[958]&m[959]&~m[960]&m[961]&m[980])|(m[958]&~m[959]&m[960]&m[961]&m[980])|(~m[958]&m[959]&m[960]&m[961]&m[980]))&~BiasedRNG[901])|((m[958]&m[959]&~m[960]&~m[961]&~m[980])|(m[958]&~m[959]&m[960]&~m[961]&~m[980])|(~m[958]&m[959]&m[960]&~m[961]&~m[980])|(m[958]&m[959]&m[960]&~m[961]&~m[980])|(m[958]&m[959]&m[960]&m[961]&~m[980])|(m[958]&m[959]&~m[960]&~m[961]&m[980])|(m[958]&~m[959]&m[960]&~m[961]&m[980])|(~m[958]&m[959]&m[960]&~m[961]&m[980])|(m[958]&m[959]&m[960]&~m[961]&m[980])|(m[958]&m[959]&m[960]&m[961]&m[980]))):InitCond[1847];
    m[967] = run?((((m[963]&~m[964]&~m[965]&~m[966]&~m[985])|(~m[963]&m[964]&~m[965]&~m[966]&~m[985])|(~m[963]&~m[964]&m[965]&~m[966]&~m[985])|(m[963]&m[964]&~m[965]&m[966]&~m[985])|(m[963]&~m[964]&m[965]&m[966]&~m[985])|(~m[963]&m[964]&m[965]&m[966]&~m[985]))&BiasedRNG[902])|(((m[963]&~m[964]&~m[965]&~m[966]&m[985])|(~m[963]&m[964]&~m[965]&~m[966]&m[985])|(~m[963]&~m[964]&m[965]&~m[966]&m[985])|(m[963]&m[964]&~m[965]&m[966]&m[985])|(m[963]&~m[964]&m[965]&m[966]&m[985])|(~m[963]&m[964]&m[965]&m[966]&m[985]))&~BiasedRNG[902])|((m[963]&m[964]&~m[965]&~m[966]&~m[985])|(m[963]&~m[964]&m[965]&~m[966]&~m[985])|(~m[963]&m[964]&m[965]&~m[966]&~m[985])|(m[963]&m[964]&m[965]&~m[966]&~m[985])|(m[963]&m[964]&m[965]&m[966]&~m[985])|(m[963]&m[964]&~m[965]&~m[966]&m[985])|(m[963]&~m[964]&m[965]&~m[966]&m[985])|(~m[963]&m[964]&m[965]&~m[966]&m[985])|(m[963]&m[964]&m[965]&~m[966]&m[985])|(m[963]&m[964]&m[965]&m[966]&m[985]))):InitCond[1848];
    m[972] = run?((((m[968]&~m[969]&~m[970]&~m[971]&~m[990])|(~m[968]&m[969]&~m[970]&~m[971]&~m[990])|(~m[968]&~m[969]&m[970]&~m[971]&~m[990])|(m[968]&m[969]&~m[970]&m[971]&~m[990])|(m[968]&~m[969]&m[970]&m[971]&~m[990])|(~m[968]&m[969]&m[970]&m[971]&~m[990]))&BiasedRNG[903])|(((m[968]&~m[969]&~m[970]&~m[971]&m[990])|(~m[968]&m[969]&~m[970]&~m[971]&m[990])|(~m[968]&~m[969]&m[970]&~m[971]&m[990])|(m[968]&m[969]&~m[970]&m[971]&m[990])|(m[968]&~m[969]&m[970]&m[971]&m[990])|(~m[968]&m[969]&m[970]&m[971]&m[990]))&~BiasedRNG[903])|((m[968]&m[969]&~m[970]&~m[971]&~m[990])|(m[968]&~m[969]&m[970]&~m[971]&~m[990])|(~m[968]&m[969]&m[970]&~m[971]&~m[990])|(m[968]&m[969]&m[970]&~m[971]&~m[990])|(m[968]&m[969]&m[970]&m[971]&~m[990])|(m[968]&m[969]&~m[970]&~m[971]&m[990])|(m[968]&~m[969]&m[970]&~m[971]&m[990])|(~m[968]&m[969]&m[970]&~m[971]&m[990])|(m[968]&m[969]&m[970]&~m[971]&m[990])|(m[968]&m[969]&m[970]&m[971]&m[990]))):InitCond[1849];
    m[977] = run?((((m[973]&~m[974]&~m[975]&~m[976]&~m[995])|(~m[973]&m[974]&~m[975]&~m[976]&~m[995])|(~m[973]&~m[974]&m[975]&~m[976]&~m[995])|(m[973]&m[974]&~m[975]&m[976]&~m[995])|(m[973]&~m[974]&m[975]&m[976]&~m[995])|(~m[973]&m[974]&m[975]&m[976]&~m[995]))&BiasedRNG[904])|(((m[973]&~m[974]&~m[975]&~m[976]&m[995])|(~m[973]&m[974]&~m[975]&~m[976]&m[995])|(~m[973]&~m[974]&m[975]&~m[976]&m[995])|(m[973]&m[974]&~m[975]&m[976]&m[995])|(m[973]&~m[974]&m[975]&m[976]&m[995])|(~m[973]&m[974]&m[975]&m[976]&m[995]))&~BiasedRNG[904])|((m[973]&m[974]&~m[975]&~m[976]&~m[995])|(m[973]&~m[974]&m[975]&~m[976]&~m[995])|(~m[973]&m[974]&m[975]&~m[976]&~m[995])|(m[973]&m[974]&m[975]&~m[976]&~m[995])|(m[973]&m[974]&m[975]&m[976]&~m[995])|(m[973]&m[974]&~m[975]&~m[976]&m[995])|(m[973]&~m[974]&m[975]&~m[976]&m[995])|(~m[973]&m[974]&m[975]&~m[976]&m[995])|(m[973]&m[974]&m[975]&~m[976]&m[995])|(m[973]&m[974]&m[975]&m[976]&m[995]))):InitCond[1850];
    m[982] = run?((((m[978]&~m[979]&~m[980]&~m[981]&~m[1005])|(~m[978]&m[979]&~m[980]&~m[981]&~m[1005])|(~m[978]&~m[979]&m[980]&~m[981]&~m[1005])|(m[978]&m[979]&~m[980]&m[981]&~m[1005])|(m[978]&~m[979]&m[980]&m[981]&~m[1005])|(~m[978]&m[979]&m[980]&m[981]&~m[1005]))&BiasedRNG[905])|(((m[978]&~m[979]&~m[980]&~m[981]&m[1005])|(~m[978]&m[979]&~m[980]&~m[981]&m[1005])|(~m[978]&~m[979]&m[980]&~m[981]&m[1005])|(m[978]&m[979]&~m[980]&m[981]&m[1005])|(m[978]&~m[979]&m[980]&m[981]&m[1005])|(~m[978]&m[979]&m[980]&m[981]&m[1005]))&~BiasedRNG[905])|((m[978]&m[979]&~m[980]&~m[981]&~m[1005])|(m[978]&~m[979]&m[980]&~m[981]&~m[1005])|(~m[978]&m[979]&m[980]&~m[981]&~m[1005])|(m[978]&m[979]&m[980]&~m[981]&~m[1005])|(m[978]&m[979]&m[980]&m[981]&~m[1005])|(m[978]&m[979]&~m[980]&~m[981]&m[1005])|(m[978]&~m[979]&m[980]&~m[981]&m[1005])|(~m[978]&m[979]&m[980]&~m[981]&m[1005])|(m[978]&m[979]&m[980]&~m[981]&m[1005])|(m[978]&m[979]&m[980]&m[981]&m[1005]))):InitCond[1851];
    m[987] = run?((((m[983]&~m[984]&~m[985]&~m[986]&~m[1010])|(~m[983]&m[984]&~m[985]&~m[986]&~m[1010])|(~m[983]&~m[984]&m[985]&~m[986]&~m[1010])|(m[983]&m[984]&~m[985]&m[986]&~m[1010])|(m[983]&~m[984]&m[985]&m[986]&~m[1010])|(~m[983]&m[984]&m[985]&m[986]&~m[1010]))&BiasedRNG[906])|(((m[983]&~m[984]&~m[985]&~m[986]&m[1010])|(~m[983]&m[984]&~m[985]&~m[986]&m[1010])|(~m[983]&~m[984]&m[985]&~m[986]&m[1010])|(m[983]&m[984]&~m[985]&m[986]&m[1010])|(m[983]&~m[984]&m[985]&m[986]&m[1010])|(~m[983]&m[984]&m[985]&m[986]&m[1010]))&~BiasedRNG[906])|((m[983]&m[984]&~m[985]&~m[986]&~m[1010])|(m[983]&~m[984]&m[985]&~m[986]&~m[1010])|(~m[983]&m[984]&m[985]&~m[986]&~m[1010])|(m[983]&m[984]&m[985]&~m[986]&~m[1010])|(m[983]&m[984]&m[985]&m[986]&~m[1010])|(m[983]&m[984]&~m[985]&~m[986]&m[1010])|(m[983]&~m[984]&m[985]&~m[986]&m[1010])|(~m[983]&m[984]&m[985]&~m[986]&m[1010])|(m[983]&m[984]&m[985]&~m[986]&m[1010])|(m[983]&m[984]&m[985]&m[986]&m[1010]))):InitCond[1852];
    m[992] = run?((((m[988]&~m[989]&~m[990]&~m[991]&~m[1015])|(~m[988]&m[989]&~m[990]&~m[991]&~m[1015])|(~m[988]&~m[989]&m[990]&~m[991]&~m[1015])|(m[988]&m[989]&~m[990]&m[991]&~m[1015])|(m[988]&~m[989]&m[990]&m[991]&~m[1015])|(~m[988]&m[989]&m[990]&m[991]&~m[1015]))&BiasedRNG[907])|(((m[988]&~m[989]&~m[990]&~m[991]&m[1015])|(~m[988]&m[989]&~m[990]&~m[991]&m[1015])|(~m[988]&~m[989]&m[990]&~m[991]&m[1015])|(m[988]&m[989]&~m[990]&m[991]&m[1015])|(m[988]&~m[989]&m[990]&m[991]&m[1015])|(~m[988]&m[989]&m[990]&m[991]&m[1015]))&~BiasedRNG[907])|((m[988]&m[989]&~m[990]&~m[991]&~m[1015])|(m[988]&~m[989]&m[990]&~m[991]&~m[1015])|(~m[988]&m[989]&m[990]&~m[991]&~m[1015])|(m[988]&m[989]&m[990]&~m[991]&~m[1015])|(m[988]&m[989]&m[990]&m[991]&~m[1015])|(m[988]&m[989]&~m[990]&~m[991]&m[1015])|(m[988]&~m[989]&m[990]&~m[991]&m[1015])|(~m[988]&m[989]&m[990]&~m[991]&m[1015])|(m[988]&m[989]&m[990]&~m[991]&m[1015])|(m[988]&m[989]&m[990]&m[991]&m[1015]))):InitCond[1853];
    m[997] = run?((((m[993]&~m[994]&~m[995]&~m[996]&~m[1020])|(~m[993]&m[994]&~m[995]&~m[996]&~m[1020])|(~m[993]&~m[994]&m[995]&~m[996]&~m[1020])|(m[993]&m[994]&~m[995]&m[996]&~m[1020])|(m[993]&~m[994]&m[995]&m[996]&~m[1020])|(~m[993]&m[994]&m[995]&m[996]&~m[1020]))&BiasedRNG[908])|(((m[993]&~m[994]&~m[995]&~m[996]&m[1020])|(~m[993]&m[994]&~m[995]&~m[996]&m[1020])|(~m[993]&~m[994]&m[995]&~m[996]&m[1020])|(m[993]&m[994]&~m[995]&m[996]&m[1020])|(m[993]&~m[994]&m[995]&m[996]&m[1020])|(~m[993]&m[994]&m[995]&m[996]&m[1020]))&~BiasedRNG[908])|((m[993]&m[994]&~m[995]&~m[996]&~m[1020])|(m[993]&~m[994]&m[995]&~m[996]&~m[1020])|(~m[993]&m[994]&m[995]&~m[996]&~m[1020])|(m[993]&m[994]&m[995]&~m[996]&~m[1020])|(m[993]&m[994]&m[995]&m[996]&~m[1020])|(m[993]&m[994]&~m[995]&~m[996]&m[1020])|(m[993]&~m[994]&m[995]&~m[996]&m[1020])|(~m[993]&m[994]&m[995]&~m[996]&m[1020])|(m[993]&m[994]&m[995]&~m[996]&m[1020])|(m[993]&m[994]&m[995]&m[996]&m[1020]))):InitCond[1854];
    m[1002] = run?((((m[998]&~m[999]&~m[1000]&~m[1001]&~m[1025])|(~m[998]&m[999]&~m[1000]&~m[1001]&~m[1025])|(~m[998]&~m[999]&m[1000]&~m[1001]&~m[1025])|(m[998]&m[999]&~m[1000]&m[1001]&~m[1025])|(m[998]&~m[999]&m[1000]&m[1001]&~m[1025])|(~m[998]&m[999]&m[1000]&m[1001]&~m[1025]))&BiasedRNG[909])|(((m[998]&~m[999]&~m[1000]&~m[1001]&m[1025])|(~m[998]&m[999]&~m[1000]&~m[1001]&m[1025])|(~m[998]&~m[999]&m[1000]&~m[1001]&m[1025])|(m[998]&m[999]&~m[1000]&m[1001]&m[1025])|(m[998]&~m[999]&m[1000]&m[1001]&m[1025])|(~m[998]&m[999]&m[1000]&m[1001]&m[1025]))&~BiasedRNG[909])|((m[998]&m[999]&~m[1000]&~m[1001]&~m[1025])|(m[998]&~m[999]&m[1000]&~m[1001]&~m[1025])|(~m[998]&m[999]&m[1000]&~m[1001]&~m[1025])|(m[998]&m[999]&m[1000]&~m[1001]&~m[1025])|(m[998]&m[999]&m[1000]&m[1001]&~m[1025])|(m[998]&m[999]&~m[1000]&~m[1001]&m[1025])|(m[998]&~m[999]&m[1000]&~m[1001]&m[1025])|(~m[998]&m[999]&m[1000]&~m[1001]&m[1025])|(m[998]&m[999]&m[1000]&~m[1001]&m[1025])|(m[998]&m[999]&m[1000]&m[1001]&m[1025]))):InitCond[1855];
    m[1007] = run?((((m[1003]&~m[1004]&~m[1005]&~m[1006]&~m[1035])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1035])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1035])|(m[1003]&m[1004]&~m[1005]&m[1006]&~m[1035])|(m[1003]&~m[1004]&m[1005]&m[1006]&~m[1035])|(~m[1003]&m[1004]&m[1005]&m[1006]&~m[1035]))&BiasedRNG[910])|(((m[1003]&~m[1004]&~m[1005]&~m[1006]&m[1035])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&m[1035])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&m[1035])|(m[1003]&m[1004]&~m[1005]&m[1006]&m[1035])|(m[1003]&~m[1004]&m[1005]&m[1006]&m[1035])|(~m[1003]&m[1004]&m[1005]&m[1006]&m[1035]))&~BiasedRNG[910])|((m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1035])|(m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1035])|(~m[1003]&m[1004]&m[1005]&~m[1006]&~m[1035])|(m[1003]&m[1004]&m[1005]&~m[1006]&~m[1035])|(m[1003]&m[1004]&m[1005]&m[1006]&~m[1035])|(m[1003]&m[1004]&~m[1005]&~m[1006]&m[1035])|(m[1003]&~m[1004]&m[1005]&~m[1006]&m[1035])|(~m[1003]&m[1004]&m[1005]&~m[1006]&m[1035])|(m[1003]&m[1004]&m[1005]&~m[1006]&m[1035])|(m[1003]&m[1004]&m[1005]&m[1006]&m[1035]))):InitCond[1856];
    m[1012] = run?((((m[1008]&~m[1009]&~m[1010]&~m[1011]&~m[1040])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1040])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1040])|(m[1008]&m[1009]&~m[1010]&m[1011]&~m[1040])|(m[1008]&~m[1009]&m[1010]&m[1011]&~m[1040])|(~m[1008]&m[1009]&m[1010]&m[1011]&~m[1040]))&BiasedRNG[911])|(((m[1008]&~m[1009]&~m[1010]&~m[1011]&m[1040])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&m[1040])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&m[1040])|(m[1008]&m[1009]&~m[1010]&m[1011]&m[1040])|(m[1008]&~m[1009]&m[1010]&m[1011]&m[1040])|(~m[1008]&m[1009]&m[1010]&m[1011]&m[1040]))&~BiasedRNG[911])|((m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1040])|(m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1040])|(~m[1008]&m[1009]&m[1010]&~m[1011]&~m[1040])|(m[1008]&m[1009]&m[1010]&~m[1011]&~m[1040])|(m[1008]&m[1009]&m[1010]&m[1011]&~m[1040])|(m[1008]&m[1009]&~m[1010]&~m[1011]&m[1040])|(m[1008]&~m[1009]&m[1010]&~m[1011]&m[1040])|(~m[1008]&m[1009]&m[1010]&~m[1011]&m[1040])|(m[1008]&m[1009]&m[1010]&~m[1011]&m[1040])|(m[1008]&m[1009]&m[1010]&m[1011]&m[1040]))):InitCond[1857];
    m[1017] = run?((((m[1013]&~m[1014]&~m[1015]&~m[1016]&~m[1045])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1045])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1045])|(m[1013]&m[1014]&~m[1015]&m[1016]&~m[1045])|(m[1013]&~m[1014]&m[1015]&m[1016]&~m[1045])|(~m[1013]&m[1014]&m[1015]&m[1016]&~m[1045]))&BiasedRNG[912])|(((m[1013]&~m[1014]&~m[1015]&~m[1016]&m[1045])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&m[1045])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&m[1045])|(m[1013]&m[1014]&~m[1015]&m[1016]&m[1045])|(m[1013]&~m[1014]&m[1015]&m[1016]&m[1045])|(~m[1013]&m[1014]&m[1015]&m[1016]&m[1045]))&~BiasedRNG[912])|((m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1045])|(m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1045])|(~m[1013]&m[1014]&m[1015]&~m[1016]&~m[1045])|(m[1013]&m[1014]&m[1015]&~m[1016]&~m[1045])|(m[1013]&m[1014]&m[1015]&m[1016]&~m[1045])|(m[1013]&m[1014]&~m[1015]&~m[1016]&m[1045])|(m[1013]&~m[1014]&m[1015]&~m[1016]&m[1045])|(~m[1013]&m[1014]&m[1015]&~m[1016]&m[1045])|(m[1013]&m[1014]&m[1015]&~m[1016]&m[1045])|(m[1013]&m[1014]&m[1015]&m[1016]&m[1045]))):InitCond[1858];
    m[1022] = run?((((m[1018]&~m[1019]&~m[1020]&~m[1021]&~m[1050])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1050])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1050])|(m[1018]&m[1019]&~m[1020]&m[1021]&~m[1050])|(m[1018]&~m[1019]&m[1020]&m[1021]&~m[1050])|(~m[1018]&m[1019]&m[1020]&m[1021]&~m[1050]))&BiasedRNG[913])|(((m[1018]&~m[1019]&~m[1020]&~m[1021]&m[1050])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&m[1050])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&m[1050])|(m[1018]&m[1019]&~m[1020]&m[1021]&m[1050])|(m[1018]&~m[1019]&m[1020]&m[1021]&m[1050])|(~m[1018]&m[1019]&m[1020]&m[1021]&m[1050]))&~BiasedRNG[913])|((m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1050])|(m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1050])|(~m[1018]&m[1019]&m[1020]&~m[1021]&~m[1050])|(m[1018]&m[1019]&m[1020]&~m[1021]&~m[1050])|(m[1018]&m[1019]&m[1020]&m[1021]&~m[1050])|(m[1018]&m[1019]&~m[1020]&~m[1021]&m[1050])|(m[1018]&~m[1019]&m[1020]&~m[1021]&m[1050])|(~m[1018]&m[1019]&m[1020]&~m[1021]&m[1050])|(m[1018]&m[1019]&m[1020]&~m[1021]&m[1050])|(m[1018]&m[1019]&m[1020]&m[1021]&m[1050]))):InitCond[1859];
    m[1027] = run?((((m[1023]&~m[1024]&~m[1025]&~m[1026]&~m[1055])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1055])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1055])|(m[1023]&m[1024]&~m[1025]&m[1026]&~m[1055])|(m[1023]&~m[1024]&m[1025]&m[1026]&~m[1055])|(~m[1023]&m[1024]&m[1025]&m[1026]&~m[1055]))&BiasedRNG[914])|(((m[1023]&~m[1024]&~m[1025]&~m[1026]&m[1055])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&m[1055])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&m[1055])|(m[1023]&m[1024]&~m[1025]&m[1026]&m[1055])|(m[1023]&~m[1024]&m[1025]&m[1026]&m[1055])|(~m[1023]&m[1024]&m[1025]&m[1026]&m[1055]))&~BiasedRNG[914])|((m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1055])|(m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1055])|(~m[1023]&m[1024]&m[1025]&~m[1026]&~m[1055])|(m[1023]&m[1024]&m[1025]&~m[1026]&~m[1055])|(m[1023]&m[1024]&m[1025]&m[1026]&~m[1055])|(m[1023]&m[1024]&~m[1025]&~m[1026]&m[1055])|(m[1023]&~m[1024]&m[1025]&~m[1026]&m[1055])|(~m[1023]&m[1024]&m[1025]&~m[1026]&m[1055])|(m[1023]&m[1024]&m[1025]&~m[1026]&m[1055])|(m[1023]&m[1024]&m[1025]&m[1026]&m[1055]))):InitCond[1860];
    m[1032] = run?((((m[1028]&~m[1029]&~m[1030]&~m[1031]&~m[1060])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1060])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1060])|(m[1028]&m[1029]&~m[1030]&m[1031]&~m[1060])|(m[1028]&~m[1029]&m[1030]&m[1031]&~m[1060])|(~m[1028]&m[1029]&m[1030]&m[1031]&~m[1060]))&BiasedRNG[915])|(((m[1028]&~m[1029]&~m[1030]&~m[1031]&m[1060])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&m[1060])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&m[1060])|(m[1028]&m[1029]&~m[1030]&m[1031]&m[1060])|(m[1028]&~m[1029]&m[1030]&m[1031]&m[1060])|(~m[1028]&m[1029]&m[1030]&m[1031]&m[1060]))&~BiasedRNG[915])|((m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1060])|(m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1060])|(~m[1028]&m[1029]&m[1030]&~m[1031]&~m[1060])|(m[1028]&m[1029]&m[1030]&~m[1031]&~m[1060])|(m[1028]&m[1029]&m[1030]&m[1031]&~m[1060])|(m[1028]&m[1029]&~m[1030]&~m[1031]&m[1060])|(m[1028]&~m[1029]&m[1030]&~m[1031]&m[1060])|(~m[1028]&m[1029]&m[1030]&~m[1031]&m[1060])|(m[1028]&m[1029]&m[1030]&~m[1031]&m[1060])|(m[1028]&m[1029]&m[1030]&m[1031]&m[1060]))):InitCond[1861];
    m[1037] = run?((((m[1033]&~m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&~m[1070]))&BiasedRNG[916])|(((m[1033]&~m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&m[1070]))&~BiasedRNG[916])|((m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&m[1070]))):InitCond[1862];
    m[1042] = run?((((m[1038]&~m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&~m[1075]))&BiasedRNG[917])|(((m[1038]&~m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&m[1075]))&~BiasedRNG[917])|((m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&m[1075]))):InitCond[1863];
    m[1047] = run?((((m[1043]&~m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&~m[1080]))&BiasedRNG[918])|(((m[1043]&~m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&m[1080]))&~BiasedRNG[918])|((m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&m[1080]))):InitCond[1864];
    m[1052] = run?((((m[1048]&~m[1049]&~m[1050]&~m[1051]&~m[1085])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1085])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1085])|(m[1048]&m[1049]&~m[1050]&m[1051]&~m[1085])|(m[1048]&~m[1049]&m[1050]&m[1051]&~m[1085])|(~m[1048]&m[1049]&m[1050]&m[1051]&~m[1085]))&BiasedRNG[919])|(((m[1048]&~m[1049]&~m[1050]&~m[1051]&m[1085])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&m[1085])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&m[1085])|(m[1048]&m[1049]&~m[1050]&m[1051]&m[1085])|(m[1048]&~m[1049]&m[1050]&m[1051]&m[1085])|(~m[1048]&m[1049]&m[1050]&m[1051]&m[1085]))&~BiasedRNG[919])|((m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1085])|(m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1085])|(~m[1048]&m[1049]&m[1050]&~m[1051]&~m[1085])|(m[1048]&m[1049]&m[1050]&~m[1051]&~m[1085])|(m[1048]&m[1049]&m[1050]&m[1051]&~m[1085])|(m[1048]&m[1049]&~m[1050]&~m[1051]&m[1085])|(m[1048]&~m[1049]&m[1050]&~m[1051]&m[1085])|(~m[1048]&m[1049]&m[1050]&~m[1051]&m[1085])|(m[1048]&m[1049]&m[1050]&~m[1051]&m[1085])|(m[1048]&m[1049]&m[1050]&m[1051]&m[1085]))):InitCond[1865];
    m[1057] = run?((((m[1053]&~m[1054]&~m[1055]&~m[1056]&~m[1090])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1090])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1090])|(m[1053]&m[1054]&~m[1055]&m[1056]&~m[1090])|(m[1053]&~m[1054]&m[1055]&m[1056]&~m[1090])|(~m[1053]&m[1054]&m[1055]&m[1056]&~m[1090]))&BiasedRNG[920])|(((m[1053]&~m[1054]&~m[1055]&~m[1056]&m[1090])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&m[1090])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&m[1090])|(m[1053]&m[1054]&~m[1055]&m[1056]&m[1090])|(m[1053]&~m[1054]&m[1055]&m[1056]&m[1090])|(~m[1053]&m[1054]&m[1055]&m[1056]&m[1090]))&~BiasedRNG[920])|((m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1090])|(m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1090])|(~m[1053]&m[1054]&m[1055]&~m[1056]&~m[1090])|(m[1053]&m[1054]&m[1055]&~m[1056]&~m[1090])|(m[1053]&m[1054]&m[1055]&m[1056]&~m[1090])|(m[1053]&m[1054]&~m[1055]&~m[1056]&m[1090])|(m[1053]&~m[1054]&m[1055]&~m[1056]&m[1090])|(~m[1053]&m[1054]&m[1055]&~m[1056]&m[1090])|(m[1053]&m[1054]&m[1055]&~m[1056]&m[1090])|(m[1053]&m[1054]&m[1055]&m[1056]&m[1090]))):InitCond[1866];
    m[1062] = run?((((m[1058]&~m[1059]&~m[1060]&~m[1061]&~m[1095])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1095])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1095])|(m[1058]&m[1059]&~m[1060]&m[1061]&~m[1095])|(m[1058]&~m[1059]&m[1060]&m[1061]&~m[1095])|(~m[1058]&m[1059]&m[1060]&m[1061]&~m[1095]))&BiasedRNG[921])|(((m[1058]&~m[1059]&~m[1060]&~m[1061]&m[1095])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&m[1095])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&m[1095])|(m[1058]&m[1059]&~m[1060]&m[1061]&m[1095])|(m[1058]&~m[1059]&m[1060]&m[1061]&m[1095])|(~m[1058]&m[1059]&m[1060]&m[1061]&m[1095]))&~BiasedRNG[921])|((m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1095])|(m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1095])|(~m[1058]&m[1059]&m[1060]&~m[1061]&~m[1095])|(m[1058]&m[1059]&m[1060]&~m[1061]&~m[1095])|(m[1058]&m[1059]&m[1060]&m[1061]&~m[1095])|(m[1058]&m[1059]&~m[1060]&~m[1061]&m[1095])|(m[1058]&~m[1059]&m[1060]&~m[1061]&m[1095])|(~m[1058]&m[1059]&m[1060]&~m[1061]&m[1095])|(m[1058]&m[1059]&m[1060]&~m[1061]&m[1095])|(m[1058]&m[1059]&m[1060]&m[1061]&m[1095]))):InitCond[1867];
    m[1067] = run?((((m[1063]&~m[1064]&~m[1065]&~m[1066]&~m[1100])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1100])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1100])|(m[1063]&m[1064]&~m[1065]&m[1066]&~m[1100])|(m[1063]&~m[1064]&m[1065]&m[1066]&~m[1100])|(~m[1063]&m[1064]&m[1065]&m[1066]&~m[1100]))&BiasedRNG[922])|(((m[1063]&~m[1064]&~m[1065]&~m[1066]&m[1100])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&m[1100])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&m[1100])|(m[1063]&m[1064]&~m[1065]&m[1066]&m[1100])|(m[1063]&~m[1064]&m[1065]&m[1066]&m[1100])|(~m[1063]&m[1064]&m[1065]&m[1066]&m[1100]))&~BiasedRNG[922])|((m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1100])|(m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1100])|(~m[1063]&m[1064]&m[1065]&~m[1066]&~m[1100])|(m[1063]&m[1064]&m[1065]&~m[1066]&~m[1100])|(m[1063]&m[1064]&m[1065]&m[1066]&~m[1100])|(m[1063]&m[1064]&~m[1065]&~m[1066]&m[1100])|(m[1063]&~m[1064]&m[1065]&~m[1066]&m[1100])|(~m[1063]&m[1064]&m[1065]&~m[1066]&m[1100])|(m[1063]&m[1064]&m[1065]&~m[1066]&m[1100])|(m[1063]&m[1064]&m[1065]&m[1066]&m[1100]))):InitCond[1868];
    m[1072] = run?((((m[1068]&~m[1069]&~m[1070]&~m[1071]&~m[1110])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1110])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1110])|(m[1068]&m[1069]&~m[1070]&m[1071]&~m[1110])|(m[1068]&~m[1069]&m[1070]&m[1071]&~m[1110])|(~m[1068]&m[1069]&m[1070]&m[1071]&~m[1110]))&BiasedRNG[923])|(((m[1068]&~m[1069]&~m[1070]&~m[1071]&m[1110])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&m[1110])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&m[1110])|(m[1068]&m[1069]&~m[1070]&m[1071]&m[1110])|(m[1068]&~m[1069]&m[1070]&m[1071]&m[1110])|(~m[1068]&m[1069]&m[1070]&m[1071]&m[1110]))&~BiasedRNG[923])|((m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1110])|(m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1110])|(~m[1068]&m[1069]&m[1070]&~m[1071]&~m[1110])|(m[1068]&m[1069]&m[1070]&~m[1071]&~m[1110])|(m[1068]&m[1069]&m[1070]&m[1071]&~m[1110])|(m[1068]&m[1069]&~m[1070]&~m[1071]&m[1110])|(m[1068]&~m[1069]&m[1070]&~m[1071]&m[1110])|(~m[1068]&m[1069]&m[1070]&~m[1071]&m[1110])|(m[1068]&m[1069]&m[1070]&~m[1071]&m[1110])|(m[1068]&m[1069]&m[1070]&m[1071]&m[1110]))):InitCond[1869];
    m[1077] = run?((((m[1073]&~m[1074]&~m[1075]&~m[1076]&~m[1115])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1115])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1115])|(m[1073]&m[1074]&~m[1075]&m[1076]&~m[1115])|(m[1073]&~m[1074]&m[1075]&m[1076]&~m[1115])|(~m[1073]&m[1074]&m[1075]&m[1076]&~m[1115]))&BiasedRNG[924])|(((m[1073]&~m[1074]&~m[1075]&~m[1076]&m[1115])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&m[1115])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&m[1115])|(m[1073]&m[1074]&~m[1075]&m[1076]&m[1115])|(m[1073]&~m[1074]&m[1075]&m[1076]&m[1115])|(~m[1073]&m[1074]&m[1075]&m[1076]&m[1115]))&~BiasedRNG[924])|((m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1115])|(m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1115])|(~m[1073]&m[1074]&m[1075]&~m[1076]&~m[1115])|(m[1073]&m[1074]&m[1075]&~m[1076]&~m[1115])|(m[1073]&m[1074]&m[1075]&m[1076]&~m[1115])|(m[1073]&m[1074]&~m[1075]&~m[1076]&m[1115])|(m[1073]&~m[1074]&m[1075]&~m[1076]&m[1115])|(~m[1073]&m[1074]&m[1075]&~m[1076]&m[1115])|(m[1073]&m[1074]&m[1075]&~m[1076]&m[1115])|(m[1073]&m[1074]&m[1075]&m[1076]&m[1115]))):InitCond[1870];
    m[1082] = run?((((m[1078]&~m[1079]&~m[1080]&~m[1081]&~m[1120])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1120])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1120])|(m[1078]&m[1079]&~m[1080]&m[1081]&~m[1120])|(m[1078]&~m[1079]&m[1080]&m[1081]&~m[1120])|(~m[1078]&m[1079]&m[1080]&m[1081]&~m[1120]))&BiasedRNG[925])|(((m[1078]&~m[1079]&~m[1080]&~m[1081]&m[1120])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&m[1120])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&m[1120])|(m[1078]&m[1079]&~m[1080]&m[1081]&m[1120])|(m[1078]&~m[1079]&m[1080]&m[1081]&m[1120])|(~m[1078]&m[1079]&m[1080]&m[1081]&m[1120]))&~BiasedRNG[925])|((m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1120])|(m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1120])|(~m[1078]&m[1079]&m[1080]&~m[1081]&~m[1120])|(m[1078]&m[1079]&m[1080]&~m[1081]&~m[1120])|(m[1078]&m[1079]&m[1080]&m[1081]&~m[1120])|(m[1078]&m[1079]&~m[1080]&~m[1081]&m[1120])|(m[1078]&~m[1079]&m[1080]&~m[1081]&m[1120])|(~m[1078]&m[1079]&m[1080]&~m[1081]&m[1120])|(m[1078]&m[1079]&m[1080]&~m[1081]&m[1120])|(m[1078]&m[1079]&m[1080]&m[1081]&m[1120]))):InitCond[1871];
    m[1087] = run?((((m[1083]&~m[1084]&~m[1085]&~m[1086]&~m[1125])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1125])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1125])|(m[1083]&m[1084]&~m[1085]&m[1086]&~m[1125])|(m[1083]&~m[1084]&m[1085]&m[1086]&~m[1125])|(~m[1083]&m[1084]&m[1085]&m[1086]&~m[1125]))&BiasedRNG[926])|(((m[1083]&~m[1084]&~m[1085]&~m[1086]&m[1125])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&m[1125])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&m[1125])|(m[1083]&m[1084]&~m[1085]&m[1086]&m[1125])|(m[1083]&~m[1084]&m[1085]&m[1086]&m[1125])|(~m[1083]&m[1084]&m[1085]&m[1086]&m[1125]))&~BiasedRNG[926])|((m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1125])|(m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1125])|(~m[1083]&m[1084]&m[1085]&~m[1086]&~m[1125])|(m[1083]&m[1084]&m[1085]&~m[1086]&~m[1125])|(m[1083]&m[1084]&m[1085]&m[1086]&~m[1125])|(m[1083]&m[1084]&~m[1085]&~m[1086]&m[1125])|(m[1083]&~m[1084]&m[1085]&~m[1086]&m[1125])|(~m[1083]&m[1084]&m[1085]&~m[1086]&m[1125])|(m[1083]&m[1084]&m[1085]&~m[1086]&m[1125])|(m[1083]&m[1084]&m[1085]&m[1086]&m[1125]))):InitCond[1872];
    m[1092] = run?((((m[1088]&~m[1089]&~m[1090]&~m[1091]&~m[1130])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1130])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1130])|(m[1088]&m[1089]&~m[1090]&m[1091]&~m[1130])|(m[1088]&~m[1089]&m[1090]&m[1091]&~m[1130])|(~m[1088]&m[1089]&m[1090]&m[1091]&~m[1130]))&BiasedRNG[927])|(((m[1088]&~m[1089]&~m[1090]&~m[1091]&m[1130])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&m[1130])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&m[1130])|(m[1088]&m[1089]&~m[1090]&m[1091]&m[1130])|(m[1088]&~m[1089]&m[1090]&m[1091]&m[1130])|(~m[1088]&m[1089]&m[1090]&m[1091]&m[1130]))&~BiasedRNG[927])|((m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1130])|(m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1130])|(~m[1088]&m[1089]&m[1090]&~m[1091]&~m[1130])|(m[1088]&m[1089]&m[1090]&~m[1091]&~m[1130])|(m[1088]&m[1089]&m[1090]&m[1091]&~m[1130])|(m[1088]&m[1089]&~m[1090]&~m[1091]&m[1130])|(m[1088]&~m[1089]&m[1090]&~m[1091]&m[1130])|(~m[1088]&m[1089]&m[1090]&~m[1091]&m[1130])|(m[1088]&m[1089]&m[1090]&~m[1091]&m[1130])|(m[1088]&m[1089]&m[1090]&m[1091]&m[1130]))):InitCond[1873];
    m[1097] = run?((((m[1093]&~m[1094]&~m[1095]&~m[1096]&~m[1135])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1135])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1135])|(m[1093]&m[1094]&~m[1095]&m[1096]&~m[1135])|(m[1093]&~m[1094]&m[1095]&m[1096]&~m[1135])|(~m[1093]&m[1094]&m[1095]&m[1096]&~m[1135]))&BiasedRNG[928])|(((m[1093]&~m[1094]&~m[1095]&~m[1096]&m[1135])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&m[1135])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&m[1135])|(m[1093]&m[1094]&~m[1095]&m[1096]&m[1135])|(m[1093]&~m[1094]&m[1095]&m[1096]&m[1135])|(~m[1093]&m[1094]&m[1095]&m[1096]&m[1135]))&~BiasedRNG[928])|((m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1135])|(m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1135])|(~m[1093]&m[1094]&m[1095]&~m[1096]&~m[1135])|(m[1093]&m[1094]&m[1095]&~m[1096]&~m[1135])|(m[1093]&m[1094]&m[1095]&m[1096]&~m[1135])|(m[1093]&m[1094]&~m[1095]&~m[1096]&m[1135])|(m[1093]&~m[1094]&m[1095]&~m[1096]&m[1135])|(~m[1093]&m[1094]&m[1095]&~m[1096]&m[1135])|(m[1093]&m[1094]&m[1095]&~m[1096]&m[1135])|(m[1093]&m[1094]&m[1095]&m[1096]&m[1135]))):InitCond[1874];
    m[1102] = run?((((m[1098]&~m[1099]&~m[1100]&~m[1101]&~m[1140])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1140])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1140])|(m[1098]&m[1099]&~m[1100]&m[1101]&~m[1140])|(m[1098]&~m[1099]&m[1100]&m[1101]&~m[1140])|(~m[1098]&m[1099]&m[1100]&m[1101]&~m[1140]))&BiasedRNG[929])|(((m[1098]&~m[1099]&~m[1100]&~m[1101]&m[1140])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&m[1140])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&m[1140])|(m[1098]&m[1099]&~m[1100]&m[1101]&m[1140])|(m[1098]&~m[1099]&m[1100]&m[1101]&m[1140])|(~m[1098]&m[1099]&m[1100]&m[1101]&m[1140]))&~BiasedRNG[929])|((m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1140])|(m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1140])|(~m[1098]&m[1099]&m[1100]&~m[1101]&~m[1140])|(m[1098]&m[1099]&m[1100]&~m[1101]&~m[1140])|(m[1098]&m[1099]&m[1100]&m[1101]&~m[1140])|(m[1098]&m[1099]&~m[1100]&~m[1101]&m[1140])|(m[1098]&~m[1099]&m[1100]&~m[1101]&m[1140])|(~m[1098]&m[1099]&m[1100]&~m[1101]&m[1140])|(m[1098]&m[1099]&m[1100]&~m[1101]&m[1140])|(m[1098]&m[1099]&m[1100]&m[1101]&m[1140]))):InitCond[1875];
    m[1107] = run?((((m[1103]&~m[1104]&~m[1105]&~m[1106]&~m[1145])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1145])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1145])|(m[1103]&m[1104]&~m[1105]&m[1106]&~m[1145])|(m[1103]&~m[1104]&m[1105]&m[1106]&~m[1145])|(~m[1103]&m[1104]&m[1105]&m[1106]&~m[1145]))&BiasedRNG[930])|(((m[1103]&~m[1104]&~m[1105]&~m[1106]&m[1145])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&m[1145])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&m[1145])|(m[1103]&m[1104]&~m[1105]&m[1106]&m[1145])|(m[1103]&~m[1104]&m[1105]&m[1106]&m[1145])|(~m[1103]&m[1104]&m[1105]&m[1106]&m[1145]))&~BiasedRNG[930])|((m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1145])|(m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1145])|(~m[1103]&m[1104]&m[1105]&~m[1106]&~m[1145])|(m[1103]&m[1104]&m[1105]&~m[1106]&~m[1145])|(m[1103]&m[1104]&m[1105]&m[1106]&~m[1145])|(m[1103]&m[1104]&~m[1105]&~m[1106]&m[1145])|(m[1103]&~m[1104]&m[1105]&~m[1106]&m[1145])|(~m[1103]&m[1104]&m[1105]&~m[1106]&m[1145])|(m[1103]&m[1104]&m[1105]&~m[1106]&m[1145])|(m[1103]&m[1104]&m[1105]&m[1106]&m[1145]))):InitCond[1876];
    m[1112] = run?((((m[1108]&~m[1109]&~m[1110]&~m[1111]&~m[1155])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1155])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1155])|(m[1108]&m[1109]&~m[1110]&m[1111]&~m[1155])|(m[1108]&~m[1109]&m[1110]&m[1111]&~m[1155])|(~m[1108]&m[1109]&m[1110]&m[1111]&~m[1155]))&BiasedRNG[931])|(((m[1108]&~m[1109]&~m[1110]&~m[1111]&m[1155])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&m[1155])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&m[1155])|(m[1108]&m[1109]&~m[1110]&m[1111]&m[1155])|(m[1108]&~m[1109]&m[1110]&m[1111]&m[1155])|(~m[1108]&m[1109]&m[1110]&m[1111]&m[1155]))&~BiasedRNG[931])|((m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1155])|(m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1155])|(~m[1108]&m[1109]&m[1110]&~m[1111]&~m[1155])|(m[1108]&m[1109]&m[1110]&~m[1111]&~m[1155])|(m[1108]&m[1109]&m[1110]&m[1111]&~m[1155])|(m[1108]&m[1109]&~m[1110]&~m[1111]&m[1155])|(m[1108]&~m[1109]&m[1110]&~m[1111]&m[1155])|(~m[1108]&m[1109]&m[1110]&~m[1111]&m[1155])|(m[1108]&m[1109]&m[1110]&~m[1111]&m[1155])|(m[1108]&m[1109]&m[1110]&m[1111]&m[1155]))):InitCond[1877];
    m[1117] = run?((((m[1113]&~m[1114]&~m[1115]&~m[1116]&~m[1160])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1160])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1160])|(m[1113]&m[1114]&~m[1115]&m[1116]&~m[1160])|(m[1113]&~m[1114]&m[1115]&m[1116]&~m[1160])|(~m[1113]&m[1114]&m[1115]&m[1116]&~m[1160]))&BiasedRNG[932])|(((m[1113]&~m[1114]&~m[1115]&~m[1116]&m[1160])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&m[1160])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&m[1160])|(m[1113]&m[1114]&~m[1115]&m[1116]&m[1160])|(m[1113]&~m[1114]&m[1115]&m[1116]&m[1160])|(~m[1113]&m[1114]&m[1115]&m[1116]&m[1160]))&~BiasedRNG[932])|((m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1160])|(m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1160])|(~m[1113]&m[1114]&m[1115]&~m[1116]&~m[1160])|(m[1113]&m[1114]&m[1115]&~m[1116]&~m[1160])|(m[1113]&m[1114]&m[1115]&m[1116]&~m[1160])|(m[1113]&m[1114]&~m[1115]&~m[1116]&m[1160])|(m[1113]&~m[1114]&m[1115]&~m[1116]&m[1160])|(~m[1113]&m[1114]&m[1115]&~m[1116]&m[1160])|(m[1113]&m[1114]&m[1115]&~m[1116]&m[1160])|(m[1113]&m[1114]&m[1115]&m[1116]&m[1160]))):InitCond[1878];
    m[1122] = run?((((m[1118]&~m[1119]&~m[1120]&~m[1121]&~m[1165])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1165])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1165])|(m[1118]&m[1119]&~m[1120]&m[1121]&~m[1165])|(m[1118]&~m[1119]&m[1120]&m[1121]&~m[1165])|(~m[1118]&m[1119]&m[1120]&m[1121]&~m[1165]))&BiasedRNG[933])|(((m[1118]&~m[1119]&~m[1120]&~m[1121]&m[1165])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&m[1165])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&m[1165])|(m[1118]&m[1119]&~m[1120]&m[1121]&m[1165])|(m[1118]&~m[1119]&m[1120]&m[1121]&m[1165])|(~m[1118]&m[1119]&m[1120]&m[1121]&m[1165]))&~BiasedRNG[933])|((m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1165])|(m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1165])|(~m[1118]&m[1119]&m[1120]&~m[1121]&~m[1165])|(m[1118]&m[1119]&m[1120]&~m[1121]&~m[1165])|(m[1118]&m[1119]&m[1120]&m[1121]&~m[1165])|(m[1118]&m[1119]&~m[1120]&~m[1121]&m[1165])|(m[1118]&~m[1119]&m[1120]&~m[1121]&m[1165])|(~m[1118]&m[1119]&m[1120]&~m[1121]&m[1165])|(m[1118]&m[1119]&m[1120]&~m[1121]&m[1165])|(m[1118]&m[1119]&m[1120]&m[1121]&m[1165]))):InitCond[1879];
    m[1127] = run?((((m[1123]&~m[1124]&~m[1125]&~m[1126]&~m[1170])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1170])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1170])|(m[1123]&m[1124]&~m[1125]&m[1126]&~m[1170])|(m[1123]&~m[1124]&m[1125]&m[1126]&~m[1170])|(~m[1123]&m[1124]&m[1125]&m[1126]&~m[1170]))&BiasedRNG[934])|(((m[1123]&~m[1124]&~m[1125]&~m[1126]&m[1170])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&m[1170])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&m[1170])|(m[1123]&m[1124]&~m[1125]&m[1126]&m[1170])|(m[1123]&~m[1124]&m[1125]&m[1126]&m[1170])|(~m[1123]&m[1124]&m[1125]&m[1126]&m[1170]))&~BiasedRNG[934])|((m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1170])|(m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1170])|(~m[1123]&m[1124]&m[1125]&~m[1126]&~m[1170])|(m[1123]&m[1124]&m[1125]&~m[1126]&~m[1170])|(m[1123]&m[1124]&m[1125]&m[1126]&~m[1170])|(m[1123]&m[1124]&~m[1125]&~m[1126]&m[1170])|(m[1123]&~m[1124]&m[1125]&~m[1126]&m[1170])|(~m[1123]&m[1124]&m[1125]&~m[1126]&m[1170])|(m[1123]&m[1124]&m[1125]&~m[1126]&m[1170])|(m[1123]&m[1124]&m[1125]&m[1126]&m[1170]))):InitCond[1880];
    m[1132] = run?((((m[1128]&~m[1129]&~m[1130]&~m[1131]&~m[1175])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1175])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1175])|(m[1128]&m[1129]&~m[1130]&m[1131]&~m[1175])|(m[1128]&~m[1129]&m[1130]&m[1131]&~m[1175])|(~m[1128]&m[1129]&m[1130]&m[1131]&~m[1175]))&BiasedRNG[935])|(((m[1128]&~m[1129]&~m[1130]&~m[1131]&m[1175])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&m[1175])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&m[1175])|(m[1128]&m[1129]&~m[1130]&m[1131]&m[1175])|(m[1128]&~m[1129]&m[1130]&m[1131]&m[1175])|(~m[1128]&m[1129]&m[1130]&m[1131]&m[1175]))&~BiasedRNG[935])|((m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1175])|(m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1175])|(~m[1128]&m[1129]&m[1130]&~m[1131]&~m[1175])|(m[1128]&m[1129]&m[1130]&~m[1131]&~m[1175])|(m[1128]&m[1129]&m[1130]&m[1131]&~m[1175])|(m[1128]&m[1129]&~m[1130]&~m[1131]&m[1175])|(m[1128]&~m[1129]&m[1130]&~m[1131]&m[1175])|(~m[1128]&m[1129]&m[1130]&~m[1131]&m[1175])|(m[1128]&m[1129]&m[1130]&~m[1131]&m[1175])|(m[1128]&m[1129]&m[1130]&m[1131]&m[1175]))):InitCond[1881];
    m[1137] = run?((((m[1133]&~m[1134]&~m[1135]&~m[1136]&~m[1180])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1180])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1180])|(m[1133]&m[1134]&~m[1135]&m[1136]&~m[1180])|(m[1133]&~m[1134]&m[1135]&m[1136]&~m[1180])|(~m[1133]&m[1134]&m[1135]&m[1136]&~m[1180]))&BiasedRNG[936])|(((m[1133]&~m[1134]&~m[1135]&~m[1136]&m[1180])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&m[1180])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&m[1180])|(m[1133]&m[1134]&~m[1135]&m[1136]&m[1180])|(m[1133]&~m[1134]&m[1135]&m[1136]&m[1180])|(~m[1133]&m[1134]&m[1135]&m[1136]&m[1180]))&~BiasedRNG[936])|((m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1180])|(m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1180])|(~m[1133]&m[1134]&m[1135]&~m[1136]&~m[1180])|(m[1133]&m[1134]&m[1135]&~m[1136]&~m[1180])|(m[1133]&m[1134]&m[1135]&m[1136]&~m[1180])|(m[1133]&m[1134]&~m[1135]&~m[1136]&m[1180])|(m[1133]&~m[1134]&m[1135]&~m[1136]&m[1180])|(~m[1133]&m[1134]&m[1135]&~m[1136]&m[1180])|(m[1133]&m[1134]&m[1135]&~m[1136]&m[1180])|(m[1133]&m[1134]&m[1135]&m[1136]&m[1180]))):InitCond[1882];
    m[1142] = run?((((m[1138]&~m[1139]&~m[1140]&~m[1141]&~m[1185])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1185])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1185])|(m[1138]&m[1139]&~m[1140]&m[1141]&~m[1185])|(m[1138]&~m[1139]&m[1140]&m[1141]&~m[1185])|(~m[1138]&m[1139]&m[1140]&m[1141]&~m[1185]))&BiasedRNG[937])|(((m[1138]&~m[1139]&~m[1140]&~m[1141]&m[1185])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&m[1185])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&m[1185])|(m[1138]&m[1139]&~m[1140]&m[1141]&m[1185])|(m[1138]&~m[1139]&m[1140]&m[1141]&m[1185])|(~m[1138]&m[1139]&m[1140]&m[1141]&m[1185]))&~BiasedRNG[937])|((m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1185])|(m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1185])|(~m[1138]&m[1139]&m[1140]&~m[1141]&~m[1185])|(m[1138]&m[1139]&m[1140]&~m[1141]&~m[1185])|(m[1138]&m[1139]&m[1140]&m[1141]&~m[1185])|(m[1138]&m[1139]&~m[1140]&~m[1141]&m[1185])|(m[1138]&~m[1139]&m[1140]&~m[1141]&m[1185])|(~m[1138]&m[1139]&m[1140]&~m[1141]&m[1185])|(m[1138]&m[1139]&m[1140]&~m[1141]&m[1185])|(m[1138]&m[1139]&m[1140]&m[1141]&m[1185]))):InitCond[1883];
    m[1147] = run?((((m[1143]&~m[1144]&~m[1145]&~m[1146]&~m[1190])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1190])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1190])|(m[1143]&m[1144]&~m[1145]&m[1146]&~m[1190])|(m[1143]&~m[1144]&m[1145]&m[1146]&~m[1190])|(~m[1143]&m[1144]&m[1145]&m[1146]&~m[1190]))&BiasedRNG[938])|(((m[1143]&~m[1144]&~m[1145]&~m[1146]&m[1190])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&m[1190])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&m[1190])|(m[1143]&m[1144]&~m[1145]&m[1146]&m[1190])|(m[1143]&~m[1144]&m[1145]&m[1146]&m[1190])|(~m[1143]&m[1144]&m[1145]&m[1146]&m[1190]))&~BiasedRNG[938])|((m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1190])|(m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1190])|(~m[1143]&m[1144]&m[1145]&~m[1146]&~m[1190])|(m[1143]&m[1144]&m[1145]&~m[1146]&~m[1190])|(m[1143]&m[1144]&m[1145]&m[1146]&~m[1190])|(m[1143]&m[1144]&~m[1145]&~m[1146]&m[1190])|(m[1143]&~m[1144]&m[1145]&~m[1146]&m[1190])|(~m[1143]&m[1144]&m[1145]&~m[1146]&m[1190])|(m[1143]&m[1144]&m[1145]&~m[1146]&m[1190])|(m[1143]&m[1144]&m[1145]&m[1146]&m[1190]))):InitCond[1884];
    m[1152] = run?((((m[1148]&~m[1149]&~m[1150]&~m[1151]&~m[1195])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1195])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1195])|(m[1148]&m[1149]&~m[1150]&m[1151]&~m[1195])|(m[1148]&~m[1149]&m[1150]&m[1151]&~m[1195])|(~m[1148]&m[1149]&m[1150]&m[1151]&~m[1195]))&BiasedRNG[939])|(((m[1148]&~m[1149]&~m[1150]&~m[1151]&m[1195])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&m[1195])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&m[1195])|(m[1148]&m[1149]&~m[1150]&m[1151]&m[1195])|(m[1148]&~m[1149]&m[1150]&m[1151]&m[1195])|(~m[1148]&m[1149]&m[1150]&m[1151]&m[1195]))&~BiasedRNG[939])|((m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1195])|(m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1195])|(~m[1148]&m[1149]&m[1150]&~m[1151]&~m[1195])|(m[1148]&m[1149]&m[1150]&~m[1151]&~m[1195])|(m[1148]&m[1149]&m[1150]&m[1151]&~m[1195])|(m[1148]&m[1149]&~m[1150]&~m[1151]&m[1195])|(m[1148]&~m[1149]&m[1150]&~m[1151]&m[1195])|(~m[1148]&m[1149]&m[1150]&~m[1151]&m[1195])|(m[1148]&m[1149]&m[1150]&~m[1151]&m[1195])|(m[1148]&m[1149]&m[1150]&m[1151]&m[1195]))):InitCond[1885];
    m[1157] = run?((((m[1153]&~m[1154]&~m[1155]&~m[1156]&~m[1205])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1205])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1205])|(m[1153]&m[1154]&~m[1155]&m[1156]&~m[1205])|(m[1153]&~m[1154]&m[1155]&m[1156]&~m[1205])|(~m[1153]&m[1154]&m[1155]&m[1156]&~m[1205]))&BiasedRNG[940])|(((m[1153]&~m[1154]&~m[1155]&~m[1156]&m[1205])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&m[1205])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&m[1205])|(m[1153]&m[1154]&~m[1155]&m[1156]&m[1205])|(m[1153]&~m[1154]&m[1155]&m[1156]&m[1205])|(~m[1153]&m[1154]&m[1155]&m[1156]&m[1205]))&~BiasedRNG[940])|((m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1205])|(m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1205])|(~m[1153]&m[1154]&m[1155]&~m[1156]&~m[1205])|(m[1153]&m[1154]&m[1155]&~m[1156]&~m[1205])|(m[1153]&m[1154]&m[1155]&m[1156]&~m[1205])|(m[1153]&m[1154]&~m[1155]&~m[1156]&m[1205])|(m[1153]&~m[1154]&m[1155]&~m[1156]&m[1205])|(~m[1153]&m[1154]&m[1155]&~m[1156]&m[1205])|(m[1153]&m[1154]&m[1155]&~m[1156]&m[1205])|(m[1153]&m[1154]&m[1155]&m[1156]&m[1205]))):InitCond[1886];
    m[1162] = run?((((m[1158]&~m[1159]&~m[1160]&~m[1161]&~m[1210])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1210])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1210])|(m[1158]&m[1159]&~m[1160]&m[1161]&~m[1210])|(m[1158]&~m[1159]&m[1160]&m[1161]&~m[1210])|(~m[1158]&m[1159]&m[1160]&m[1161]&~m[1210]))&BiasedRNG[941])|(((m[1158]&~m[1159]&~m[1160]&~m[1161]&m[1210])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&m[1210])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&m[1210])|(m[1158]&m[1159]&~m[1160]&m[1161]&m[1210])|(m[1158]&~m[1159]&m[1160]&m[1161]&m[1210])|(~m[1158]&m[1159]&m[1160]&m[1161]&m[1210]))&~BiasedRNG[941])|((m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1210])|(m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1210])|(~m[1158]&m[1159]&m[1160]&~m[1161]&~m[1210])|(m[1158]&m[1159]&m[1160]&~m[1161]&~m[1210])|(m[1158]&m[1159]&m[1160]&m[1161]&~m[1210])|(m[1158]&m[1159]&~m[1160]&~m[1161]&m[1210])|(m[1158]&~m[1159]&m[1160]&~m[1161]&m[1210])|(~m[1158]&m[1159]&m[1160]&~m[1161]&m[1210])|(m[1158]&m[1159]&m[1160]&~m[1161]&m[1210])|(m[1158]&m[1159]&m[1160]&m[1161]&m[1210]))):InitCond[1887];
    m[1167] = run?((((m[1163]&~m[1164]&~m[1165]&~m[1166]&~m[1215])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1215])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1215])|(m[1163]&m[1164]&~m[1165]&m[1166]&~m[1215])|(m[1163]&~m[1164]&m[1165]&m[1166]&~m[1215])|(~m[1163]&m[1164]&m[1165]&m[1166]&~m[1215]))&BiasedRNG[942])|(((m[1163]&~m[1164]&~m[1165]&~m[1166]&m[1215])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&m[1215])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&m[1215])|(m[1163]&m[1164]&~m[1165]&m[1166]&m[1215])|(m[1163]&~m[1164]&m[1165]&m[1166]&m[1215])|(~m[1163]&m[1164]&m[1165]&m[1166]&m[1215]))&~BiasedRNG[942])|((m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1215])|(m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1215])|(~m[1163]&m[1164]&m[1165]&~m[1166]&~m[1215])|(m[1163]&m[1164]&m[1165]&~m[1166]&~m[1215])|(m[1163]&m[1164]&m[1165]&m[1166]&~m[1215])|(m[1163]&m[1164]&~m[1165]&~m[1166]&m[1215])|(m[1163]&~m[1164]&m[1165]&~m[1166]&m[1215])|(~m[1163]&m[1164]&m[1165]&~m[1166]&m[1215])|(m[1163]&m[1164]&m[1165]&~m[1166]&m[1215])|(m[1163]&m[1164]&m[1165]&m[1166]&m[1215]))):InitCond[1888];
    m[1172] = run?((((m[1168]&~m[1169]&~m[1170]&~m[1171]&~m[1220])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1220])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1220])|(m[1168]&m[1169]&~m[1170]&m[1171]&~m[1220])|(m[1168]&~m[1169]&m[1170]&m[1171]&~m[1220])|(~m[1168]&m[1169]&m[1170]&m[1171]&~m[1220]))&BiasedRNG[943])|(((m[1168]&~m[1169]&~m[1170]&~m[1171]&m[1220])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&m[1220])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&m[1220])|(m[1168]&m[1169]&~m[1170]&m[1171]&m[1220])|(m[1168]&~m[1169]&m[1170]&m[1171]&m[1220])|(~m[1168]&m[1169]&m[1170]&m[1171]&m[1220]))&~BiasedRNG[943])|((m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1220])|(m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1220])|(~m[1168]&m[1169]&m[1170]&~m[1171]&~m[1220])|(m[1168]&m[1169]&m[1170]&~m[1171]&~m[1220])|(m[1168]&m[1169]&m[1170]&m[1171]&~m[1220])|(m[1168]&m[1169]&~m[1170]&~m[1171]&m[1220])|(m[1168]&~m[1169]&m[1170]&~m[1171]&m[1220])|(~m[1168]&m[1169]&m[1170]&~m[1171]&m[1220])|(m[1168]&m[1169]&m[1170]&~m[1171]&m[1220])|(m[1168]&m[1169]&m[1170]&m[1171]&m[1220]))):InitCond[1889];
    m[1177] = run?((((m[1173]&~m[1174]&~m[1175]&~m[1176]&~m[1225])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1225])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1225])|(m[1173]&m[1174]&~m[1175]&m[1176]&~m[1225])|(m[1173]&~m[1174]&m[1175]&m[1176]&~m[1225])|(~m[1173]&m[1174]&m[1175]&m[1176]&~m[1225]))&BiasedRNG[944])|(((m[1173]&~m[1174]&~m[1175]&~m[1176]&m[1225])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&m[1225])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&m[1225])|(m[1173]&m[1174]&~m[1175]&m[1176]&m[1225])|(m[1173]&~m[1174]&m[1175]&m[1176]&m[1225])|(~m[1173]&m[1174]&m[1175]&m[1176]&m[1225]))&~BiasedRNG[944])|((m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1225])|(m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1225])|(~m[1173]&m[1174]&m[1175]&~m[1176]&~m[1225])|(m[1173]&m[1174]&m[1175]&~m[1176]&~m[1225])|(m[1173]&m[1174]&m[1175]&m[1176]&~m[1225])|(m[1173]&m[1174]&~m[1175]&~m[1176]&m[1225])|(m[1173]&~m[1174]&m[1175]&~m[1176]&m[1225])|(~m[1173]&m[1174]&m[1175]&~m[1176]&m[1225])|(m[1173]&m[1174]&m[1175]&~m[1176]&m[1225])|(m[1173]&m[1174]&m[1175]&m[1176]&m[1225]))):InitCond[1890];
    m[1182] = run?((((m[1178]&~m[1179]&~m[1180]&~m[1181]&~m[1230])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1230])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1230])|(m[1178]&m[1179]&~m[1180]&m[1181]&~m[1230])|(m[1178]&~m[1179]&m[1180]&m[1181]&~m[1230])|(~m[1178]&m[1179]&m[1180]&m[1181]&~m[1230]))&BiasedRNG[945])|(((m[1178]&~m[1179]&~m[1180]&~m[1181]&m[1230])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&m[1230])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&m[1230])|(m[1178]&m[1179]&~m[1180]&m[1181]&m[1230])|(m[1178]&~m[1179]&m[1180]&m[1181]&m[1230])|(~m[1178]&m[1179]&m[1180]&m[1181]&m[1230]))&~BiasedRNG[945])|((m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1230])|(m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1230])|(~m[1178]&m[1179]&m[1180]&~m[1181]&~m[1230])|(m[1178]&m[1179]&m[1180]&~m[1181]&~m[1230])|(m[1178]&m[1179]&m[1180]&m[1181]&~m[1230])|(m[1178]&m[1179]&~m[1180]&~m[1181]&m[1230])|(m[1178]&~m[1179]&m[1180]&~m[1181]&m[1230])|(~m[1178]&m[1179]&m[1180]&~m[1181]&m[1230])|(m[1178]&m[1179]&m[1180]&~m[1181]&m[1230])|(m[1178]&m[1179]&m[1180]&m[1181]&m[1230]))):InitCond[1891];
    m[1187] = run?((((m[1183]&~m[1184]&~m[1185]&~m[1186]&~m[1235])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1235])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1235])|(m[1183]&m[1184]&~m[1185]&m[1186]&~m[1235])|(m[1183]&~m[1184]&m[1185]&m[1186]&~m[1235])|(~m[1183]&m[1184]&m[1185]&m[1186]&~m[1235]))&BiasedRNG[946])|(((m[1183]&~m[1184]&~m[1185]&~m[1186]&m[1235])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&m[1235])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&m[1235])|(m[1183]&m[1184]&~m[1185]&m[1186]&m[1235])|(m[1183]&~m[1184]&m[1185]&m[1186]&m[1235])|(~m[1183]&m[1184]&m[1185]&m[1186]&m[1235]))&~BiasedRNG[946])|((m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1235])|(m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1235])|(~m[1183]&m[1184]&m[1185]&~m[1186]&~m[1235])|(m[1183]&m[1184]&m[1185]&~m[1186]&~m[1235])|(m[1183]&m[1184]&m[1185]&m[1186]&~m[1235])|(m[1183]&m[1184]&~m[1185]&~m[1186]&m[1235])|(m[1183]&~m[1184]&m[1185]&~m[1186]&m[1235])|(~m[1183]&m[1184]&m[1185]&~m[1186]&m[1235])|(m[1183]&m[1184]&m[1185]&~m[1186]&m[1235])|(m[1183]&m[1184]&m[1185]&m[1186]&m[1235]))):InitCond[1892];
    m[1192] = run?((((m[1188]&~m[1189]&~m[1190]&~m[1191]&~m[1240])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1240])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1240])|(m[1188]&m[1189]&~m[1190]&m[1191]&~m[1240])|(m[1188]&~m[1189]&m[1190]&m[1191]&~m[1240])|(~m[1188]&m[1189]&m[1190]&m[1191]&~m[1240]))&BiasedRNG[947])|(((m[1188]&~m[1189]&~m[1190]&~m[1191]&m[1240])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&m[1240])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&m[1240])|(m[1188]&m[1189]&~m[1190]&m[1191]&m[1240])|(m[1188]&~m[1189]&m[1190]&m[1191]&m[1240])|(~m[1188]&m[1189]&m[1190]&m[1191]&m[1240]))&~BiasedRNG[947])|((m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1240])|(m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1240])|(~m[1188]&m[1189]&m[1190]&~m[1191]&~m[1240])|(m[1188]&m[1189]&m[1190]&~m[1191]&~m[1240])|(m[1188]&m[1189]&m[1190]&m[1191]&~m[1240])|(m[1188]&m[1189]&~m[1190]&~m[1191]&m[1240])|(m[1188]&~m[1189]&m[1190]&~m[1191]&m[1240])|(~m[1188]&m[1189]&m[1190]&~m[1191]&m[1240])|(m[1188]&m[1189]&m[1190]&~m[1191]&m[1240])|(m[1188]&m[1189]&m[1190]&m[1191]&m[1240]))):InitCond[1893];
    m[1197] = run?((((m[1193]&~m[1194]&~m[1195]&~m[1196]&~m[1245])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1245])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1245])|(m[1193]&m[1194]&~m[1195]&m[1196]&~m[1245])|(m[1193]&~m[1194]&m[1195]&m[1196]&~m[1245])|(~m[1193]&m[1194]&m[1195]&m[1196]&~m[1245]))&BiasedRNG[948])|(((m[1193]&~m[1194]&~m[1195]&~m[1196]&m[1245])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&m[1245])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&m[1245])|(m[1193]&m[1194]&~m[1195]&m[1196]&m[1245])|(m[1193]&~m[1194]&m[1195]&m[1196]&m[1245])|(~m[1193]&m[1194]&m[1195]&m[1196]&m[1245]))&~BiasedRNG[948])|((m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1245])|(m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1245])|(~m[1193]&m[1194]&m[1195]&~m[1196]&~m[1245])|(m[1193]&m[1194]&m[1195]&~m[1196]&~m[1245])|(m[1193]&m[1194]&m[1195]&m[1196]&~m[1245])|(m[1193]&m[1194]&~m[1195]&~m[1196]&m[1245])|(m[1193]&~m[1194]&m[1195]&~m[1196]&m[1245])|(~m[1193]&m[1194]&m[1195]&~m[1196]&m[1245])|(m[1193]&m[1194]&m[1195]&~m[1196]&m[1245])|(m[1193]&m[1194]&m[1195]&m[1196]&m[1245]))):InitCond[1894];
    m[1202] = run?((((m[1198]&~m[1199]&~m[1200]&~m[1201]&~m[1250])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1250])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1250])|(m[1198]&m[1199]&~m[1200]&m[1201]&~m[1250])|(m[1198]&~m[1199]&m[1200]&m[1201]&~m[1250])|(~m[1198]&m[1199]&m[1200]&m[1201]&~m[1250]))&BiasedRNG[949])|(((m[1198]&~m[1199]&~m[1200]&~m[1201]&m[1250])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&m[1250])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&m[1250])|(m[1198]&m[1199]&~m[1200]&m[1201]&m[1250])|(m[1198]&~m[1199]&m[1200]&m[1201]&m[1250])|(~m[1198]&m[1199]&m[1200]&m[1201]&m[1250]))&~BiasedRNG[949])|((m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1250])|(m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1250])|(~m[1198]&m[1199]&m[1200]&~m[1201]&~m[1250])|(m[1198]&m[1199]&m[1200]&~m[1201]&~m[1250])|(m[1198]&m[1199]&m[1200]&m[1201]&~m[1250])|(m[1198]&m[1199]&~m[1200]&~m[1201]&m[1250])|(m[1198]&~m[1199]&m[1200]&~m[1201]&m[1250])|(~m[1198]&m[1199]&m[1200]&~m[1201]&m[1250])|(m[1198]&m[1199]&m[1200]&~m[1201]&m[1250])|(m[1198]&m[1199]&m[1200]&m[1201]&m[1250]))):InitCond[1895];
    m[1207] = run?((((m[1203]&~m[1204]&~m[1205]&~m[1206]&~m[1260])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1260])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1260])|(m[1203]&m[1204]&~m[1205]&m[1206]&~m[1260])|(m[1203]&~m[1204]&m[1205]&m[1206]&~m[1260])|(~m[1203]&m[1204]&m[1205]&m[1206]&~m[1260]))&BiasedRNG[950])|(((m[1203]&~m[1204]&~m[1205]&~m[1206]&m[1260])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&m[1260])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&m[1260])|(m[1203]&m[1204]&~m[1205]&m[1206]&m[1260])|(m[1203]&~m[1204]&m[1205]&m[1206]&m[1260])|(~m[1203]&m[1204]&m[1205]&m[1206]&m[1260]))&~BiasedRNG[950])|((m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1260])|(m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1260])|(~m[1203]&m[1204]&m[1205]&~m[1206]&~m[1260])|(m[1203]&m[1204]&m[1205]&~m[1206]&~m[1260])|(m[1203]&m[1204]&m[1205]&m[1206]&~m[1260])|(m[1203]&m[1204]&~m[1205]&~m[1206]&m[1260])|(m[1203]&~m[1204]&m[1205]&~m[1206]&m[1260])|(~m[1203]&m[1204]&m[1205]&~m[1206]&m[1260])|(m[1203]&m[1204]&m[1205]&~m[1206]&m[1260])|(m[1203]&m[1204]&m[1205]&m[1206]&m[1260]))):InitCond[1896];
    m[1212] = run?((((m[1208]&~m[1209]&~m[1210]&~m[1211]&~m[1265])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1265])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1265])|(m[1208]&m[1209]&~m[1210]&m[1211]&~m[1265])|(m[1208]&~m[1209]&m[1210]&m[1211]&~m[1265])|(~m[1208]&m[1209]&m[1210]&m[1211]&~m[1265]))&BiasedRNG[951])|(((m[1208]&~m[1209]&~m[1210]&~m[1211]&m[1265])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&m[1265])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&m[1265])|(m[1208]&m[1209]&~m[1210]&m[1211]&m[1265])|(m[1208]&~m[1209]&m[1210]&m[1211]&m[1265])|(~m[1208]&m[1209]&m[1210]&m[1211]&m[1265]))&~BiasedRNG[951])|((m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1265])|(m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1265])|(~m[1208]&m[1209]&m[1210]&~m[1211]&~m[1265])|(m[1208]&m[1209]&m[1210]&~m[1211]&~m[1265])|(m[1208]&m[1209]&m[1210]&m[1211]&~m[1265])|(m[1208]&m[1209]&~m[1210]&~m[1211]&m[1265])|(m[1208]&~m[1209]&m[1210]&~m[1211]&m[1265])|(~m[1208]&m[1209]&m[1210]&~m[1211]&m[1265])|(m[1208]&m[1209]&m[1210]&~m[1211]&m[1265])|(m[1208]&m[1209]&m[1210]&m[1211]&m[1265]))):InitCond[1897];
    m[1217] = run?((((m[1213]&~m[1214]&~m[1215]&~m[1216]&~m[1270])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1270])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1270])|(m[1213]&m[1214]&~m[1215]&m[1216]&~m[1270])|(m[1213]&~m[1214]&m[1215]&m[1216]&~m[1270])|(~m[1213]&m[1214]&m[1215]&m[1216]&~m[1270]))&BiasedRNG[952])|(((m[1213]&~m[1214]&~m[1215]&~m[1216]&m[1270])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&m[1270])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&m[1270])|(m[1213]&m[1214]&~m[1215]&m[1216]&m[1270])|(m[1213]&~m[1214]&m[1215]&m[1216]&m[1270])|(~m[1213]&m[1214]&m[1215]&m[1216]&m[1270]))&~BiasedRNG[952])|((m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1270])|(m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1270])|(~m[1213]&m[1214]&m[1215]&~m[1216]&~m[1270])|(m[1213]&m[1214]&m[1215]&~m[1216]&~m[1270])|(m[1213]&m[1214]&m[1215]&m[1216]&~m[1270])|(m[1213]&m[1214]&~m[1215]&~m[1216]&m[1270])|(m[1213]&~m[1214]&m[1215]&~m[1216]&m[1270])|(~m[1213]&m[1214]&m[1215]&~m[1216]&m[1270])|(m[1213]&m[1214]&m[1215]&~m[1216]&m[1270])|(m[1213]&m[1214]&m[1215]&m[1216]&m[1270]))):InitCond[1898];
    m[1222] = run?((((m[1218]&~m[1219]&~m[1220]&~m[1221]&~m[1275])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1275])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1275])|(m[1218]&m[1219]&~m[1220]&m[1221]&~m[1275])|(m[1218]&~m[1219]&m[1220]&m[1221]&~m[1275])|(~m[1218]&m[1219]&m[1220]&m[1221]&~m[1275]))&BiasedRNG[953])|(((m[1218]&~m[1219]&~m[1220]&~m[1221]&m[1275])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&m[1275])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&m[1275])|(m[1218]&m[1219]&~m[1220]&m[1221]&m[1275])|(m[1218]&~m[1219]&m[1220]&m[1221]&m[1275])|(~m[1218]&m[1219]&m[1220]&m[1221]&m[1275]))&~BiasedRNG[953])|((m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1275])|(m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1275])|(~m[1218]&m[1219]&m[1220]&~m[1221]&~m[1275])|(m[1218]&m[1219]&m[1220]&~m[1221]&~m[1275])|(m[1218]&m[1219]&m[1220]&m[1221]&~m[1275])|(m[1218]&m[1219]&~m[1220]&~m[1221]&m[1275])|(m[1218]&~m[1219]&m[1220]&~m[1221]&m[1275])|(~m[1218]&m[1219]&m[1220]&~m[1221]&m[1275])|(m[1218]&m[1219]&m[1220]&~m[1221]&m[1275])|(m[1218]&m[1219]&m[1220]&m[1221]&m[1275]))):InitCond[1899];
    m[1227] = run?((((m[1223]&~m[1224]&~m[1225]&~m[1226]&~m[1280])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1280])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1280])|(m[1223]&m[1224]&~m[1225]&m[1226]&~m[1280])|(m[1223]&~m[1224]&m[1225]&m[1226]&~m[1280])|(~m[1223]&m[1224]&m[1225]&m[1226]&~m[1280]))&BiasedRNG[954])|(((m[1223]&~m[1224]&~m[1225]&~m[1226]&m[1280])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&m[1280])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&m[1280])|(m[1223]&m[1224]&~m[1225]&m[1226]&m[1280])|(m[1223]&~m[1224]&m[1225]&m[1226]&m[1280])|(~m[1223]&m[1224]&m[1225]&m[1226]&m[1280]))&~BiasedRNG[954])|((m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1280])|(m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1280])|(~m[1223]&m[1224]&m[1225]&~m[1226]&~m[1280])|(m[1223]&m[1224]&m[1225]&~m[1226]&~m[1280])|(m[1223]&m[1224]&m[1225]&m[1226]&~m[1280])|(m[1223]&m[1224]&~m[1225]&~m[1226]&m[1280])|(m[1223]&~m[1224]&m[1225]&~m[1226]&m[1280])|(~m[1223]&m[1224]&m[1225]&~m[1226]&m[1280])|(m[1223]&m[1224]&m[1225]&~m[1226]&m[1280])|(m[1223]&m[1224]&m[1225]&m[1226]&m[1280]))):InitCond[1900];
    m[1232] = run?((((m[1228]&~m[1229]&~m[1230]&~m[1231]&~m[1285])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1285])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1285])|(m[1228]&m[1229]&~m[1230]&m[1231]&~m[1285])|(m[1228]&~m[1229]&m[1230]&m[1231]&~m[1285])|(~m[1228]&m[1229]&m[1230]&m[1231]&~m[1285]))&BiasedRNG[955])|(((m[1228]&~m[1229]&~m[1230]&~m[1231]&m[1285])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&m[1285])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&m[1285])|(m[1228]&m[1229]&~m[1230]&m[1231]&m[1285])|(m[1228]&~m[1229]&m[1230]&m[1231]&m[1285])|(~m[1228]&m[1229]&m[1230]&m[1231]&m[1285]))&~BiasedRNG[955])|((m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1285])|(m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1285])|(~m[1228]&m[1229]&m[1230]&~m[1231]&~m[1285])|(m[1228]&m[1229]&m[1230]&~m[1231]&~m[1285])|(m[1228]&m[1229]&m[1230]&m[1231]&~m[1285])|(m[1228]&m[1229]&~m[1230]&~m[1231]&m[1285])|(m[1228]&~m[1229]&m[1230]&~m[1231]&m[1285])|(~m[1228]&m[1229]&m[1230]&~m[1231]&m[1285])|(m[1228]&m[1229]&m[1230]&~m[1231]&m[1285])|(m[1228]&m[1229]&m[1230]&m[1231]&m[1285]))):InitCond[1901];
    m[1237] = run?((((m[1233]&~m[1234]&~m[1235]&~m[1236]&~m[1290])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1290])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1290])|(m[1233]&m[1234]&~m[1235]&m[1236]&~m[1290])|(m[1233]&~m[1234]&m[1235]&m[1236]&~m[1290])|(~m[1233]&m[1234]&m[1235]&m[1236]&~m[1290]))&BiasedRNG[956])|(((m[1233]&~m[1234]&~m[1235]&~m[1236]&m[1290])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&m[1290])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&m[1290])|(m[1233]&m[1234]&~m[1235]&m[1236]&m[1290])|(m[1233]&~m[1234]&m[1235]&m[1236]&m[1290])|(~m[1233]&m[1234]&m[1235]&m[1236]&m[1290]))&~BiasedRNG[956])|((m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1290])|(m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1290])|(~m[1233]&m[1234]&m[1235]&~m[1236]&~m[1290])|(m[1233]&m[1234]&m[1235]&~m[1236]&~m[1290])|(m[1233]&m[1234]&m[1235]&m[1236]&~m[1290])|(m[1233]&m[1234]&~m[1235]&~m[1236]&m[1290])|(m[1233]&~m[1234]&m[1235]&~m[1236]&m[1290])|(~m[1233]&m[1234]&m[1235]&~m[1236]&m[1290])|(m[1233]&m[1234]&m[1235]&~m[1236]&m[1290])|(m[1233]&m[1234]&m[1235]&m[1236]&m[1290]))):InitCond[1902];
    m[1242] = run?((((m[1238]&~m[1239]&~m[1240]&~m[1241]&~m[1295])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1295])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1295])|(m[1238]&m[1239]&~m[1240]&m[1241]&~m[1295])|(m[1238]&~m[1239]&m[1240]&m[1241]&~m[1295])|(~m[1238]&m[1239]&m[1240]&m[1241]&~m[1295]))&BiasedRNG[957])|(((m[1238]&~m[1239]&~m[1240]&~m[1241]&m[1295])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&m[1295])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&m[1295])|(m[1238]&m[1239]&~m[1240]&m[1241]&m[1295])|(m[1238]&~m[1239]&m[1240]&m[1241]&m[1295])|(~m[1238]&m[1239]&m[1240]&m[1241]&m[1295]))&~BiasedRNG[957])|((m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1295])|(m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1295])|(~m[1238]&m[1239]&m[1240]&~m[1241]&~m[1295])|(m[1238]&m[1239]&m[1240]&~m[1241]&~m[1295])|(m[1238]&m[1239]&m[1240]&m[1241]&~m[1295])|(m[1238]&m[1239]&~m[1240]&~m[1241]&m[1295])|(m[1238]&~m[1239]&m[1240]&~m[1241]&m[1295])|(~m[1238]&m[1239]&m[1240]&~m[1241]&m[1295])|(m[1238]&m[1239]&m[1240]&~m[1241]&m[1295])|(m[1238]&m[1239]&m[1240]&m[1241]&m[1295]))):InitCond[1903];
    m[1247] = run?((((m[1243]&~m[1244]&~m[1245]&~m[1246]&~m[1300])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1300])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1300])|(m[1243]&m[1244]&~m[1245]&m[1246]&~m[1300])|(m[1243]&~m[1244]&m[1245]&m[1246]&~m[1300])|(~m[1243]&m[1244]&m[1245]&m[1246]&~m[1300]))&BiasedRNG[958])|(((m[1243]&~m[1244]&~m[1245]&~m[1246]&m[1300])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&m[1300])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&m[1300])|(m[1243]&m[1244]&~m[1245]&m[1246]&m[1300])|(m[1243]&~m[1244]&m[1245]&m[1246]&m[1300])|(~m[1243]&m[1244]&m[1245]&m[1246]&m[1300]))&~BiasedRNG[958])|((m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1300])|(m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1300])|(~m[1243]&m[1244]&m[1245]&~m[1246]&~m[1300])|(m[1243]&m[1244]&m[1245]&~m[1246]&~m[1300])|(m[1243]&m[1244]&m[1245]&m[1246]&~m[1300])|(m[1243]&m[1244]&~m[1245]&~m[1246]&m[1300])|(m[1243]&~m[1244]&m[1245]&~m[1246]&m[1300])|(~m[1243]&m[1244]&m[1245]&~m[1246]&m[1300])|(m[1243]&m[1244]&m[1245]&~m[1246]&m[1300])|(m[1243]&m[1244]&m[1245]&m[1246]&m[1300]))):InitCond[1904];
    m[1252] = run?((((m[1248]&~m[1249]&~m[1250]&~m[1251]&~m[1305])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1305])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1305])|(m[1248]&m[1249]&~m[1250]&m[1251]&~m[1305])|(m[1248]&~m[1249]&m[1250]&m[1251]&~m[1305])|(~m[1248]&m[1249]&m[1250]&m[1251]&~m[1305]))&BiasedRNG[959])|(((m[1248]&~m[1249]&~m[1250]&~m[1251]&m[1305])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&m[1305])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&m[1305])|(m[1248]&m[1249]&~m[1250]&m[1251]&m[1305])|(m[1248]&~m[1249]&m[1250]&m[1251]&m[1305])|(~m[1248]&m[1249]&m[1250]&m[1251]&m[1305]))&~BiasedRNG[959])|((m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1305])|(m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1305])|(~m[1248]&m[1249]&m[1250]&~m[1251]&~m[1305])|(m[1248]&m[1249]&m[1250]&~m[1251]&~m[1305])|(m[1248]&m[1249]&m[1250]&m[1251]&~m[1305])|(m[1248]&m[1249]&~m[1250]&~m[1251]&m[1305])|(m[1248]&~m[1249]&m[1250]&~m[1251]&m[1305])|(~m[1248]&m[1249]&m[1250]&~m[1251]&m[1305])|(m[1248]&m[1249]&m[1250]&~m[1251]&m[1305])|(m[1248]&m[1249]&m[1250]&m[1251]&m[1305]))):InitCond[1905];
    m[1257] = run?((((m[1253]&~m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&~m[1310]))&BiasedRNG[960])|(((m[1253]&~m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&m[1310]))&~BiasedRNG[960])|((m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&m[1310]))):InitCond[1906];
    m[1262] = run?((((m[1258]&~m[1259]&~m[1260]&~m[1261]&~m[1320])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1320])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1320])|(m[1258]&m[1259]&~m[1260]&m[1261]&~m[1320])|(m[1258]&~m[1259]&m[1260]&m[1261]&~m[1320])|(~m[1258]&m[1259]&m[1260]&m[1261]&~m[1320]))&BiasedRNG[961])|(((m[1258]&~m[1259]&~m[1260]&~m[1261]&m[1320])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&m[1320])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&m[1320])|(m[1258]&m[1259]&~m[1260]&m[1261]&m[1320])|(m[1258]&~m[1259]&m[1260]&m[1261]&m[1320])|(~m[1258]&m[1259]&m[1260]&m[1261]&m[1320]))&~BiasedRNG[961])|((m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1320])|(m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1320])|(~m[1258]&m[1259]&m[1260]&~m[1261]&~m[1320])|(m[1258]&m[1259]&m[1260]&~m[1261]&~m[1320])|(m[1258]&m[1259]&m[1260]&m[1261]&~m[1320])|(m[1258]&m[1259]&~m[1260]&~m[1261]&m[1320])|(m[1258]&~m[1259]&m[1260]&~m[1261]&m[1320])|(~m[1258]&m[1259]&m[1260]&~m[1261]&m[1320])|(m[1258]&m[1259]&m[1260]&~m[1261]&m[1320])|(m[1258]&m[1259]&m[1260]&m[1261]&m[1320]))):InitCond[1907];
    m[1267] = run?((((m[1263]&~m[1264]&~m[1265]&~m[1266]&~m[1325])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1325])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1325])|(m[1263]&m[1264]&~m[1265]&m[1266]&~m[1325])|(m[1263]&~m[1264]&m[1265]&m[1266]&~m[1325])|(~m[1263]&m[1264]&m[1265]&m[1266]&~m[1325]))&BiasedRNG[962])|(((m[1263]&~m[1264]&~m[1265]&~m[1266]&m[1325])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&m[1325])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&m[1325])|(m[1263]&m[1264]&~m[1265]&m[1266]&m[1325])|(m[1263]&~m[1264]&m[1265]&m[1266]&m[1325])|(~m[1263]&m[1264]&m[1265]&m[1266]&m[1325]))&~BiasedRNG[962])|((m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1325])|(m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1325])|(~m[1263]&m[1264]&m[1265]&~m[1266]&~m[1325])|(m[1263]&m[1264]&m[1265]&~m[1266]&~m[1325])|(m[1263]&m[1264]&m[1265]&m[1266]&~m[1325])|(m[1263]&m[1264]&~m[1265]&~m[1266]&m[1325])|(m[1263]&~m[1264]&m[1265]&~m[1266]&m[1325])|(~m[1263]&m[1264]&m[1265]&~m[1266]&m[1325])|(m[1263]&m[1264]&m[1265]&~m[1266]&m[1325])|(m[1263]&m[1264]&m[1265]&m[1266]&m[1325]))):InitCond[1908];
    m[1272] = run?((((m[1268]&~m[1269]&~m[1270]&~m[1271]&~m[1330])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1330])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1330])|(m[1268]&m[1269]&~m[1270]&m[1271]&~m[1330])|(m[1268]&~m[1269]&m[1270]&m[1271]&~m[1330])|(~m[1268]&m[1269]&m[1270]&m[1271]&~m[1330]))&BiasedRNG[963])|(((m[1268]&~m[1269]&~m[1270]&~m[1271]&m[1330])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&m[1330])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&m[1330])|(m[1268]&m[1269]&~m[1270]&m[1271]&m[1330])|(m[1268]&~m[1269]&m[1270]&m[1271]&m[1330])|(~m[1268]&m[1269]&m[1270]&m[1271]&m[1330]))&~BiasedRNG[963])|((m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1330])|(m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1330])|(~m[1268]&m[1269]&m[1270]&~m[1271]&~m[1330])|(m[1268]&m[1269]&m[1270]&~m[1271]&~m[1330])|(m[1268]&m[1269]&m[1270]&m[1271]&~m[1330])|(m[1268]&m[1269]&~m[1270]&~m[1271]&m[1330])|(m[1268]&~m[1269]&m[1270]&~m[1271]&m[1330])|(~m[1268]&m[1269]&m[1270]&~m[1271]&m[1330])|(m[1268]&m[1269]&m[1270]&~m[1271]&m[1330])|(m[1268]&m[1269]&m[1270]&m[1271]&m[1330]))):InitCond[1909];
    m[1277] = run?((((m[1273]&~m[1274]&~m[1275]&~m[1276]&~m[1335])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1335])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1335])|(m[1273]&m[1274]&~m[1275]&m[1276]&~m[1335])|(m[1273]&~m[1274]&m[1275]&m[1276]&~m[1335])|(~m[1273]&m[1274]&m[1275]&m[1276]&~m[1335]))&BiasedRNG[964])|(((m[1273]&~m[1274]&~m[1275]&~m[1276]&m[1335])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&m[1335])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&m[1335])|(m[1273]&m[1274]&~m[1275]&m[1276]&m[1335])|(m[1273]&~m[1274]&m[1275]&m[1276]&m[1335])|(~m[1273]&m[1274]&m[1275]&m[1276]&m[1335]))&~BiasedRNG[964])|((m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1335])|(m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1335])|(~m[1273]&m[1274]&m[1275]&~m[1276]&~m[1335])|(m[1273]&m[1274]&m[1275]&~m[1276]&~m[1335])|(m[1273]&m[1274]&m[1275]&m[1276]&~m[1335])|(m[1273]&m[1274]&~m[1275]&~m[1276]&m[1335])|(m[1273]&~m[1274]&m[1275]&~m[1276]&m[1335])|(~m[1273]&m[1274]&m[1275]&~m[1276]&m[1335])|(m[1273]&m[1274]&m[1275]&~m[1276]&m[1335])|(m[1273]&m[1274]&m[1275]&m[1276]&m[1335]))):InitCond[1910];
    m[1282] = run?((((m[1278]&~m[1279]&~m[1280]&~m[1281]&~m[1340])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1340])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1340])|(m[1278]&m[1279]&~m[1280]&m[1281]&~m[1340])|(m[1278]&~m[1279]&m[1280]&m[1281]&~m[1340])|(~m[1278]&m[1279]&m[1280]&m[1281]&~m[1340]))&BiasedRNG[965])|(((m[1278]&~m[1279]&~m[1280]&~m[1281]&m[1340])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&m[1340])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&m[1340])|(m[1278]&m[1279]&~m[1280]&m[1281]&m[1340])|(m[1278]&~m[1279]&m[1280]&m[1281]&m[1340])|(~m[1278]&m[1279]&m[1280]&m[1281]&m[1340]))&~BiasedRNG[965])|((m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1340])|(m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1340])|(~m[1278]&m[1279]&m[1280]&~m[1281]&~m[1340])|(m[1278]&m[1279]&m[1280]&~m[1281]&~m[1340])|(m[1278]&m[1279]&m[1280]&m[1281]&~m[1340])|(m[1278]&m[1279]&~m[1280]&~m[1281]&m[1340])|(m[1278]&~m[1279]&m[1280]&~m[1281]&m[1340])|(~m[1278]&m[1279]&m[1280]&~m[1281]&m[1340])|(m[1278]&m[1279]&m[1280]&~m[1281]&m[1340])|(m[1278]&m[1279]&m[1280]&m[1281]&m[1340]))):InitCond[1911];
    m[1287] = run?((((m[1283]&~m[1284]&~m[1285]&~m[1286]&~m[1345])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1345])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1345])|(m[1283]&m[1284]&~m[1285]&m[1286]&~m[1345])|(m[1283]&~m[1284]&m[1285]&m[1286]&~m[1345])|(~m[1283]&m[1284]&m[1285]&m[1286]&~m[1345]))&BiasedRNG[966])|(((m[1283]&~m[1284]&~m[1285]&~m[1286]&m[1345])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&m[1345])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&m[1345])|(m[1283]&m[1284]&~m[1285]&m[1286]&m[1345])|(m[1283]&~m[1284]&m[1285]&m[1286]&m[1345])|(~m[1283]&m[1284]&m[1285]&m[1286]&m[1345]))&~BiasedRNG[966])|((m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1345])|(m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1345])|(~m[1283]&m[1284]&m[1285]&~m[1286]&~m[1345])|(m[1283]&m[1284]&m[1285]&~m[1286]&~m[1345])|(m[1283]&m[1284]&m[1285]&m[1286]&~m[1345])|(m[1283]&m[1284]&~m[1285]&~m[1286]&m[1345])|(m[1283]&~m[1284]&m[1285]&~m[1286]&m[1345])|(~m[1283]&m[1284]&m[1285]&~m[1286]&m[1345])|(m[1283]&m[1284]&m[1285]&~m[1286]&m[1345])|(m[1283]&m[1284]&m[1285]&m[1286]&m[1345]))):InitCond[1912];
    m[1292] = run?((((m[1288]&~m[1289]&~m[1290]&~m[1291]&~m[1350])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1350])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1350])|(m[1288]&m[1289]&~m[1290]&m[1291]&~m[1350])|(m[1288]&~m[1289]&m[1290]&m[1291]&~m[1350])|(~m[1288]&m[1289]&m[1290]&m[1291]&~m[1350]))&BiasedRNG[967])|(((m[1288]&~m[1289]&~m[1290]&~m[1291]&m[1350])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&m[1350])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&m[1350])|(m[1288]&m[1289]&~m[1290]&m[1291]&m[1350])|(m[1288]&~m[1289]&m[1290]&m[1291]&m[1350])|(~m[1288]&m[1289]&m[1290]&m[1291]&m[1350]))&~BiasedRNG[967])|((m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1350])|(m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1350])|(~m[1288]&m[1289]&m[1290]&~m[1291]&~m[1350])|(m[1288]&m[1289]&m[1290]&~m[1291]&~m[1350])|(m[1288]&m[1289]&m[1290]&m[1291]&~m[1350])|(m[1288]&m[1289]&~m[1290]&~m[1291]&m[1350])|(m[1288]&~m[1289]&m[1290]&~m[1291]&m[1350])|(~m[1288]&m[1289]&m[1290]&~m[1291]&m[1350])|(m[1288]&m[1289]&m[1290]&~m[1291]&m[1350])|(m[1288]&m[1289]&m[1290]&m[1291]&m[1350]))):InitCond[1913];
    m[1297] = run?((((m[1293]&~m[1294]&~m[1295]&~m[1296]&~m[1355])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1355])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1355])|(m[1293]&m[1294]&~m[1295]&m[1296]&~m[1355])|(m[1293]&~m[1294]&m[1295]&m[1296]&~m[1355])|(~m[1293]&m[1294]&m[1295]&m[1296]&~m[1355]))&BiasedRNG[968])|(((m[1293]&~m[1294]&~m[1295]&~m[1296]&m[1355])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&m[1355])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&m[1355])|(m[1293]&m[1294]&~m[1295]&m[1296]&m[1355])|(m[1293]&~m[1294]&m[1295]&m[1296]&m[1355])|(~m[1293]&m[1294]&m[1295]&m[1296]&m[1355]))&~BiasedRNG[968])|((m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1355])|(m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1355])|(~m[1293]&m[1294]&m[1295]&~m[1296]&~m[1355])|(m[1293]&m[1294]&m[1295]&~m[1296]&~m[1355])|(m[1293]&m[1294]&m[1295]&m[1296]&~m[1355])|(m[1293]&m[1294]&~m[1295]&~m[1296]&m[1355])|(m[1293]&~m[1294]&m[1295]&~m[1296]&m[1355])|(~m[1293]&m[1294]&m[1295]&~m[1296]&m[1355])|(m[1293]&m[1294]&m[1295]&~m[1296]&m[1355])|(m[1293]&m[1294]&m[1295]&m[1296]&m[1355]))):InitCond[1914];
    m[1302] = run?((((m[1298]&~m[1299]&~m[1300]&~m[1301]&~m[1360])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1360])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1360])|(m[1298]&m[1299]&~m[1300]&m[1301]&~m[1360])|(m[1298]&~m[1299]&m[1300]&m[1301]&~m[1360])|(~m[1298]&m[1299]&m[1300]&m[1301]&~m[1360]))&BiasedRNG[969])|(((m[1298]&~m[1299]&~m[1300]&~m[1301]&m[1360])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&m[1360])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&m[1360])|(m[1298]&m[1299]&~m[1300]&m[1301]&m[1360])|(m[1298]&~m[1299]&m[1300]&m[1301]&m[1360])|(~m[1298]&m[1299]&m[1300]&m[1301]&m[1360]))&~BiasedRNG[969])|((m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1360])|(m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1360])|(~m[1298]&m[1299]&m[1300]&~m[1301]&~m[1360])|(m[1298]&m[1299]&m[1300]&~m[1301]&~m[1360])|(m[1298]&m[1299]&m[1300]&m[1301]&~m[1360])|(m[1298]&m[1299]&~m[1300]&~m[1301]&m[1360])|(m[1298]&~m[1299]&m[1300]&~m[1301]&m[1360])|(~m[1298]&m[1299]&m[1300]&~m[1301]&m[1360])|(m[1298]&m[1299]&m[1300]&~m[1301]&m[1360])|(m[1298]&m[1299]&m[1300]&m[1301]&m[1360]))):InitCond[1915];
    m[1307] = run?((((m[1303]&~m[1304]&~m[1305]&~m[1306]&~m[1365])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1365])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1365])|(m[1303]&m[1304]&~m[1305]&m[1306]&~m[1365])|(m[1303]&~m[1304]&m[1305]&m[1306]&~m[1365])|(~m[1303]&m[1304]&m[1305]&m[1306]&~m[1365]))&BiasedRNG[970])|(((m[1303]&~m[1304]&~m[1305]&~m[1306]&m[1365])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&m[1365])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&m[1365])|(m[1303]&m[1304]&~m[1305]&m[1306]&m[1365])|(m[1303]&~m[1304]&m[1305]&m[1306]&m[1365])|(~m[1303]&m[1304]&m[1305]&m[1306]&m[1365]))&~BiasedRNG[970])|((m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1365])|(m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1365])|(~m[1303]&m[1304]&m[1305]&~m[1306]&~m[1365])|(m[1303]&m[1304]&m[1305]&~m[1306]&~m[1365])|(m[1303]&m[1304]&m[1305]&m[1306]&~m[1365])|(m[1303]&m[1304]&~m[1305]&~m[1306]&m[1365])|(m[1303]&~m[1304]&m[1305]&~m[1306]&m[1365])|(~m[1303]&m[1304]&m[1305]&~m[1306]&m[1365])|(m[1303]&m[1304]&m[1305]&~m[1306]&m[1365])|(m[1303]&m[1304]&m[1305]&m[1306]&m[1365]))):InitCond[1916];
    m[1312] = run?((((m[1308]&~m[1309]&~m[1310]&~m[1311]&~m[1370])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1370])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1370])|(m[1308]&m[1309]&~m[1310]&m[1311]&~m[1370])|(m[1308]&~m[1309]&m[1310]&m[1311]&~m[1370])|(~m[1308]&m[1309]&m[1310]&m[1311]&~m[1370]))&BiasedRNG[971])|(((m[1308]&~m[1309]&~m[1310]&~m[1311]&m[1370])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&m[1370])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&m[1370])|(m[1308]&m[1309]&~m[1310]&m[1311]&m[1370])|(m[1308]&~m[1309]&m[1310]&m[1311]&m[1370])|(~m[1308]&m[1309]&m[1310]&m[1311]&m[1370]))&~BiasedRNG[971])|((m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1370])|(m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1370])|(~m[1308]&m[1309]&m[1310]&~m[1311]&~m[1370])|(m[1308]&m[1309]&m[1310]&~m[1311]&~m[1370])|(m[1308]&m[1309]&m[1310]&m[1311]&~m[1370])|(m[1308]&m[1309]&~m[1310]&~m[1311]&m[1370])|(m[1308]&~m[1309]&m[1310]&~m[1311]&m[1370])|(~m[1308]&m[1309]&m[1310]&~m[1311]&m[1370])|(m[1308]&m[1309]&m[1310]&~m[1311]&m[1370])|(m[1308]&m[1309]&m[1310]&m[1311]&m[1370]))):InitCond[1917];
    m[1317] = run?((((m[1313]&~m[1314]&~m[1315]&~m[1316]&~m[1375])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1375])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1375])|(m[1313]&m[1314]&~m[1315]&m[1316]&~m[1375])|(m[1313]&~m[1314]&m[1315]&m[1316]&~m[1375])|(~m[1313]&m[1314]&m[1315]&m[1316]&~m[1375]))&BiasedRNG[972])|(((m[1313]&~m[1314]&~m[1315]&~m[1316]&m[1375])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&m[1375])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&m[1375])|(m[1313]&m[1314]&~m[1315]&m[1316]&m[1375])|(m[1313]&~m[1314]&m[1315]&m[1316]&m[1375])|(~m[1313]&m[1314]&m[1315]&m[1316]&m[1375]))&~BiasedRNG[972])|((m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1375])|(m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1375])|(~m[1313]&m[1314]&m[1315]&~m[1316]&~m[1375])|(m[1313]&m[1314]&m[1315]&~m[1316]&~m[1375])|(m[1313]&m[1314]&m[1315]&m[1316]&~m[1375])|(m[1313]&m[1314]&~m[1315]&~m[1316]&m[1375])|(m[1313]&~m[1314]&m[1315]&~m[1316]&m[1375])|(~m[1313]&m[1314]&m[1315]&~m[1316]&m[1375])|(m[1313]&m[1314]&m[1315]&~m[1316]&m[1375])|(m[1313]&m[1314]&m[1315]&m[1316]&m[1375]))):InitCond[1918];
    m[1322] = run?((((m[1318]&~m[1319]&~m[1320]&~m[1321]&~m[1385])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1385])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1385])|(m[1318]&m[1319]&~m[1320]&m[1321]&~m[1385])|(m[1318]&~m[1319]&m[1320]&m[1321]&~m[1385])|(~m[1318]&m[1319]&m[1320]&m[1321]&~m[1385]))&BiasedRNG[973])|(((m[1318]&~m[1319]&~m[1320]&~m[1321]&m[1385])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&m[1385])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&m[1385])|(m[1318]&m[1319]&~m[1320]&m[1321]&m[1385])|(m[1318]&~m[1319]&m[1320]&m[1321]&m[1385])|(~m[1318]&m[1319]&m[1320]&m[1321]&m[1385]))&~BiasedRNG[973])|((m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1385])|(m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1385])|(~m[1318]&m[1319]&m[1320]&~m[1321]&~m[1385])|(m[1318]&m[1319]&m[1320]&~m[1321]&~m[1385])|(m[1318]&m[1319]&m[1320]&m[1321]&~m[1385])|(m[1318]&m[1319]&~m[1320]&~m[1321]&m[1385])|(m[1318]&~m[1319]&m[1320]&~m[1321]&m[1385])|(~m[1318]&m[1319]&m[1320]&~m[1321]&m[1385])|(m[1318]&m[1319]&m[1320]&~m[1321]&m[1385])|(m[1318]&m[1319]&m[1320]&m[1321]&m[1385]))):InitCond[1919];
    m[1327] = run?((((m[1323]&~m[1324]&~m[1325]&~m[1326]&~m[1390])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1390])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1390])|(m[1323]&m[1324]&~m[1325]&m[1326]&~m[1390])|(m[1323]&~m[1324]&m[1325]&m[1326]&~m[1390])|(~m[1323]&m[1324]&m[1325]&m[1326]&~m[1390]))&BiasedRNG[974])|(((m[1323]&~m[1324]&~m[1325]&~m[1326]&m[1390])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&m[1390])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&m[1390])|(m[1323]&m[1324]&~m[1325]&m[1326]&m[1390])|(m[1323]&~m[1324]&m[1325]&m[1326]&m[1390])|(~m[1323]&m[1324]&m[1325]&m[1326]&m[1390]))&~BiasedRNG[974])|((m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1390])|(m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1390])|(~m[1323]&m[1324]&m[1325]&~m[1326]&~m[1390])|(m[1323]&m[1324]&m[1325]&~m[1326]&~m[1390])|(m[1323]&m[1324]&m[1325]&m[1326]&~m[1390])|(m[1323]&m[1324]&~m[1325]&~m[1326]&m[1390])|(m[1323]&~m[1324]&m[1325]&~m[1326]&m[1390])|(~m[1323]&m[1324]&m[1325]&~m[1326]&m[1390])|(m[1323]&m[1324]&m[1325]&~m[1326]&m[1390])|(m[1323]&m[1324]&m[1325]&m[1326]&m[1390]))):InitCond[1920];
    m[1332] = run?((((m[1328]&~m[1329]&~m[1330]&~m[1331]&~m[1395])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1395])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1395])|(m[1328]&m[1329]&~m[1330]&m[1331]&~m[1395])|(m[1328]&~m[1329]&m[1330]&m[1331]&~m[1395])|(~m[1328]&m[1329]&m[1330]&m[1331]&~m[1395]))&BiasedRNG[975])|(((m[1328]&~m[1329]&~m[1330]&~m[1331]&m[1395])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&m[1395])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&m[1395])|(m[1328]&m[1329]&~m[1330]&m[1331]&m[1395])|(m[1328]&~m[1329]&m[1330]&m[1331]&m[1395])|(~m[1328]&m[1329]&m[1330]&m[1331]&m[1395]))&~BiasedRNG[975])|((m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1395])|(m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1395])|(~m[1328]&m[1329]&m[1330]&~m[1331]&~m[1395])|(m[1328]&m[1329]&m[1330]&~m[1331]&~m[1395])|(m[1328]&m[1329]&m[1330]&m[1331]&~m[1395])|(m[1328]&m[1329]&~m[1330]&~m[1331]&m[1395])|(m[1328]&~m[1329]&m[1330]&~m[1331]&m[1395])|(~m[1328]&m[1329]&m[1330]&~m[1331]&m[1395])|(m[1328]&m[1329]&m[1330]&~m[1331]&m[1395])|(m[1328]&m[1329]&m[1330]&m[1331]&m[1395]))):InitCond[1921];
    m[1337] = run?((((m[1333]&~m[1334]&~m[1335]&~m[1336]&~m[1400])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1400])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1400])|(m[1333]&m[1334]&~m[1335]&m[1336]&~m[1400])|(m[1333]&~m[1334]&m[1335]&m[1336]&~m[1400])|(~m[1333]&m[1334]&m[1335]&m[1336]&~m[1400]))&BiasedRNG[976])|(((m[1333]&~m[1334]&~m[1335]&~m[1336]&m[1400])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&m[1400])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&m[1400])|(m[1333]&m[1334]&~m[1335]&m[1336]&m[1400])|(m[1333]&~m[1334]&m[1335]&m[1336]&m[1400])|(~m[1333]&m[1334]&m[1335]&m[1336]&m[1400]))&~BiasedRNG[976])|((m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1400])|(m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1400])|(~m[1333]&m[1334]&m[1335]&~m[1336]&~m[1400])|(m[1333]&m[1334]&m[1335]&~m[1336]&~m[1400])|(m[1333]&m[1334]&m[1335]&m[1336]&~m[1400])|(m[1333]&m[1334]&~m[1335]&~m[1336]&m[1400])|(m[1333]&~m[1334]&m[1335]&~m[1336]&m[1400])|(~m[1333]&m[1334]&m[1335]&~m[1336]&m[1400])|(m[1333]&m[1334]&m[1335]&~m[1336]&m[1400])|(m[1333]&m[1334]&m[1335]&m[1336]&m[1400]))):InitCond[1922];
    m[1342] = run?((((m[1338]&~m[1339]&~m[1340]&~m[1341]&~m[1405])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1405])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1405])|(m[1338]&m[1339]&~m[1340]&m[1341]&~m[1405])|(m[1338]&~m[1339]&m[1340]&m[1341]&~m[1405])|(~m[1338]&m[1339]&m[1340]&m[1341]&~m[1405]))&BiasedRNG[977])|(((m[1338]&~m[1339]&~m[1340]&~m[1341]&m[1405])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&m[1405])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&m[1405])|(m[1338]&m[1339]&~m[1340]&m[1341]&m[1405])|(m[1338]&~m[1339]&m[1340]&m[1341]&m[1405])|(~m[1338]&m[1339]&m[1340]&m[1341]&m[1405]))&~BiasedRNG[977])|((m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1405])|(m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1405])|(~m[1338]&m[1339]&m[1340]&~m[1341]&~m[1405])|(m[1338]&m[1339]&m[1340]&~m[1341]&~m[1405])|(m[1338]&m[1339]&m[1340]&m[1341]&~m[1405])|(m[1338]&m[1339]&~m[1340]&~m[1341]&m[1405])|(m[1338]&~m[1339]&m[1340]&~m[1341]&m[1405])|(~m[1338]&m[1339]&m[1340]&~m[1341]&m[1405])|(m[1338]&m[1339]&m[1340]&~m[1341]&m[1405])|(m[1338]&m[1339]&m[1340]&m[1341]&m[1405]))):InitCond[1923];
    m[1347] = run?((((m[1343]&~m[1344]&~m[1345]&~m[1346]&~m[1410])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1410])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1410])|(m[1343]&m[1344]&~m[1345]&m[1346]&~m[1410])|(m[1343]&~m[1344]&m[1345]&m[1346]&~m[1410])|(~m[1343]&m[1344]&m[1345]&m[1346]&~m[1410]))&BiasedRNG[978])|(((m[1343]&~m[1344]&~m[1345]&~m[1346]&m[1410])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&m[1410])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&m[1410])|(m[1343]&m[1344]&~m[1345]&m[1346]&m[1410])|(m[1343]&~m[1344]&m[1345]&m[1346]&m[1410])|(~m[1343]&m[1344]&m[1345]&m[1346]&m[1410]))&~BiasedRNG[978])|((m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1410])|(m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1410])|(~m[1343]&m[1344]&m[1345]&~m[1346]&~m[1410])|(m[1343]&m[1344]&m[1345]&~m[1346]&~m[1410])|(m[1343]&m[1344]&m[1345]&m[1346]&~m[1410])|(m[1343]&m[1344]&~m[1345]&~m[1346]&m[1410])|(m[1343]&~m[1344]&m[1345]&~m[1346]&m[1410])|(~m[1343]&m[1344]&m[1345]&~m[1346]&m[1410])|(m[1343]&m[1344]&m[1345]&~m[1346]&m[1410])|(m[1343]&m[1344]&m[1345]&m[1346]&m[1410]))):InitCond[1924];
    m[1352] = run?((((m[1348]&~m[1349]&~m[1350]&~m[1351]&~m[1415])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1415])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1415])|(m[1348]&m[1349]&~m[1350]&m[1351]&~m[1415])|(m[1348]&~m[1349]&m[1350]&m[1351]&~m[1415])|(~m[1348]&m[1349]&m[1350]&m[1351]&~m[1415]))&BiasedRNG[979])|(((m[1348]&~m[1349]&~m[1350]&~m[1351]&m[1415])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&m[1415])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&m[1415])|(m[1348]&m[1349]&~m[1350]&m[1351]&m[1415])|(m[1348]&~m[1349]&m[1350]&m[1351]&m[1415])|(~m[1348]&m[1349]&m[1350]&m[1351]&m[1415]))&~BiasedRNG[979])|((m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1415])|(m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1415])|(~m[1348]&m[1349]&m[1350]&~m[1351]&~m[1415])|(m[1348]&m[1349]&m[1350]&~m[1351]&~m[1415])|(m[1348]&m[1349]&m[1350]&m[1351]&~m[1415])|(m[1348]&m[1349]&~m[1350]&~m[1351]&m[1415])|(m[1348]&~m[1349]&m[1350]&~m[1351]&m[1415])|(~m[1348]&m[1349]&m[1350]&~m[1351]&m[1415])|(m[1348]&m[1349]&m[1350]&~m[1351]&m[1415])|(m[1348]&m[1349]&m[1350]&m[1351]&m[1415]))):InitCond[1925];
    m[1357] = run?((((m[1353]&~m[1354]&~m[1355]&~m[1356]&~m[1420])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1420])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1420])|(m[1353]&m[1354]&~m[1355]&m[1356]&~m[1420])|(m[1353]&~m[1354]&m[1355]&m[1356]&~m[1420])|(~m[1353]&m[1354]&m[1355]&m[1356]&~m[1420]))&BiasedRNG[980])|(((m[1353]&~m[1354]&~m[1355]&~m[1356]&m[1420])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&m[1420])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&m[1420])|(m[1353]&m[1354]&~m[1355]&m[1356]&m[1420])|(m[1353]&~m[1354]&m[1355]&m[1356]&m[1420])|(~m[1353]&m[1354]&m[1355]&m[1356]&m[1420]))&~BiasedRNG[980])|((m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1420])|(m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1420])|(~m[1353]&m[1354]&m[1355]&~m[1356]&~m[1420])|(m[1353]&m[1354]&m[1355]&~m[1356]&~m[1420])|(m[1353]&m[1354]&m[1355]&m[1356]&~m[1420])|(m[1353]&m[1354]&~m[1355]&~m[1356]&m[1420])|(m[1353]&~m[1354]&m[1355]&~m[1356]&m[1420])|(~m[1353]&m[1354]&m[1355]&~m[1356]&m[1420])|(m[1353]&m[1354]&m[1355]&~m[1356]&m[1420])|(m[1353]&m[1354]&m[1355]&m[1356]&m[1420]))):InitCond[1926];
    m[1362] = run?((((m[1358]&~m[1359]&~m[1360]&~m[1361]&~m[1425])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1425])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1425])|(m[1358]&m[1359]&~m[1360]&m[1361]&~m[1425])|(m[1358]&~m[1359]&m[1360]&m[1361]&~m[1425])|(~m[1358]&m[1359]&m[1360]&m[1361]&~m[1425]))&BiasedRNG[981])|(((m[1358]&~m[1359]&~m[1360]&~m[1361]&m[1425])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&m[1425])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&m[1425])|(m[1358]&m[1359]&~m[1360]&m[1361]&m[1425])|(m[1358]&~m[1359]&m[1360]&m[1361]&m[1425])|(~m[1358]&m[1359]&m[1360]&m[1361]&m[1425]))&~BiasedRNG[981])|((m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1425])|(m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1425])|(~m[1358]&m[1359]&m[1360]&~m[1361]&~m[1425])|(m[1358]&m[1359]&m[1360]&~m[1361]&~m[1425])|(m[1358]&m[1359]&m[1360]&m[1361]&~m[1425])|(m[1358]&m[1359]&~m[1360]&~m[1361]&m[1425])|(m[1358]&~m[1359]&m[1360]&~m[1361]&m[1425])|(~m[1358]&m[1359]&m[1360]&~m[1361]&m[1425])|(m[1358]&m[1359]&m[1360]&~m[1361]&m[1425])|(m[1358]&m[1359]&m[1360]&m[1361]&m[1425]))):InitCond[1927];
    m[1367] = run?((((m[1363]&~m[1364]&~m[1365]&~m[1366]&~m[1430])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1430])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1430])|(m[1363]&m[1364]&~m[1365]&m[1366]&~m[1430])|(m[1363]&~m[1364]&m[1365]&m[1366]&~m[1430])|(~m[1363]&m[1364]&m[1365]&m[1366]&~m[1430]))&BiasedRNG[982])|(((m[1363]&~m[1364]&~m[1365]&~m[1366]&m[1430])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&m[1430])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&m[1430])|(m[1363]&m[1364]&~m[1365]&m[1366]&m[1430])|(m[1363]&~m[1364]&m[1365]&m[1366]&m[1430])|(~m[1363]&m[1364]&m[1365]&m[1366]&m[1430]))&~BiasedRNG[982])|((m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1430])|(m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1430])|(~m[1363]&m[1364]&m[1365]&~m[1366]&~m[1430])|(m[1363]&m[1364]&m[1365]&~m[1366]&~m[1430])|(m[1363]&m[1364]&m[1365]&m[1366]&~m[1430])|(m[1363]&m[1364]&~m[1365]&~m[1366]&m[1430])|(m[1363]&~m[1364]&m[1365]&~m[1366]&m[1430])|(~m[1363]&m[1364]&m[1365]&~m[1366]&m[1430])|(m[1363]&m[1364]&m[1365]&~m[1366]&m[1430])|(m[1363]&m[1364]&m[1365]&m[1366]&m[1430]))):InitCond[1928];
    m[1372] = run?((((m[1368]&~m[1369]&~m[1370]&~m[1371]&~m[1435])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1435])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1435])|(m[1368]&m[1369]&~m[1370]&m[1371]&~m[1435])|(m[1368]&~m[1369]&m[1370]&m[1371]&~m[1435])|(~m[1368]&m[1369]&m[1370]&m[1371]&~m[1435]))&BiasedRNG[983])|(((m[1368]&~m[1369]&~m[1370]&~m[1371]&m[1435])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&m[1435])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&m[1435])|(m[1368]&m[1369]&~m[1370]&m[1371]&m[1435])|(m[1368]&~m[1369]&m[1370]&m[1371]&m[1435])|(~m[1368]&m[1369]&m[1370]&m[1371]&m[1435]))&~BiasedRNG[983])|((m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1435])|(m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1435])|(~m[1368]&m[1369]&m[1370]&~m[1371]&~m[1435])|(m[1368]&m[1369]&m[1370]&~m[1371]&~m[1435])|(m[1368]&m[1369]&m[1370]&m[1371]&~m[1435])|(m[1368]&m[1369]&~m[1370]&~m[1371]&m[1435])|(m[1368]&~m[1369]&m[1370]&~m[1371]&m[1435])|(~m[1368]&m[1369]&m[1370]&~m[1371]&m[1435])|(m[1368]&m[1369]&m[1370]&~m[1371]&m[1435])|(m[1368]&m[1369]&m[1370]&m[1371]&m[1435]))):InitCond[1929];
    m[1377] = run?((((m[1373]&~m[1374]&~m[1375]&~m[1376]&~m[1440])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1440])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1440])|(m[1373]&m[1374]&~m[1375]&m[1376]&~m[1440])|(m[1373]&~m[1374]&m[1375]&m[1376]&~m[1440])|(~m[1373]&m[1374]&m[1375]&m[1376]&~m[1440]))&BiasedRNG[984])|(((m[1373]&~m[1374]&~m[1375]&~m[1376]&m[1440])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&m[1440])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&m[1440])|(m[1373]&m[1374]&~m[1375]&m[1376]&m[1440])|(m[1373]&~m[1374]&m[1375]&m[1376]&m[1440])|(~m[1373]&m[1374]&m[1375]&m[1376]&m[1440]))&~BiasedRNG[984])|((m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1440])|(m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1440])|(~m[1373]&m[1374]&m[1375]&~m[1376]&~m[1440])|(m[1373]&m[1374]&m[1375]&~m[1376]&~m[1440])|(m[1373]&m[1374]&m[1375]&m[1376]&~m[1440])|(m[1373]&m[1374]&~m[1375]&~m[1376]&m[1440])|(m[1373]&~m[1374]&m[1375]&~m[1376]&m[1440])|(~m[1373]&m[1374]&m[1375]&~m[1376]&m[1440])|(m[1373]&m[1374]&m[1375]&~m[1376]&m[1440])|(m[1373]&m[1374]&m[1375]&m[1376]&m[1440]))):InitCond[1930];
    m[1382] = run?((((m[1378]&~m[1379]&~m[1380]&~m[1381]&~m[1445])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1445])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1445])|(m[1378]&m[1379]&~m[1380]&m[1381]&~m[1445])|(m[1378]&~m[1379]&m[1380]&m[1381]&~m[1445])|(~m[1378]&m[1379]&m[1380]&m[1381]&~m[1445]))&BiasedRNG[985])|(((m[1378]&~m[1379]&~m[1380]&~m[1381]&m[1445])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&m[1445])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&m[1445])|(m[1378]&m[1379]&~m[1380]&m[1381]&m[1445])|(m[1378]&~m[1379]&m[1380]&m[1381]&m[1445])|(~m[1378]&m[1379]&m[1380]&m[1381]&m[1445]))&~BiasedRNG[985])|((m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1445])|(m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1445])|(~m[1378]&m[1379]&m[1380]&~m[1381]&~m[1445])|(m[1378]&m[1379]&m[1380]&~m[1381]&~m[1445])|(m[1378]&m[1379]&m[1380]&m[1381]&~m[1445])|(m[1378]&m[1379]&~m[1380]&~m[1381]&m[1445])|(m[1378]&~m[1379]&m[1380]&~m[1381]&m[1445])|(~m[1378]&m[1379]&m[1380]&~m[1381]&m[1445])|(m[1378]&m[1379]&m[1380]&~m[1381]&m[1445])|(m[1378]&m[1379]&m[1380]&m[1381]&m[1445]))):InitCond[1931];
    m[1387] = run?((((m[1383]&~m[1384]&~m[1385]&~m[1386]&~m[1455])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1455])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1455])|(m[1383]&m[1384]&~m[1385]&m[1386]&~m[1455])|(m[1383]&~m[1384]&m[1385]&m[1386]&~m[1455])|(~m[1383]&m[1384]&m[1385]&m[1386]&~m[1455]))&BiasedRNG[986])|(((m[1383]&~m[1384]&~m[1385]&~m[1386]&m[1455])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&m[1455])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&m[1455])|(m[1383]&m[1384]&~m[1385]&m[1386]&m[1455])|(m[1383]&~m[1384]&m[1385]&m[1386]&m[1455])|(~m[1383]&m[1384]&m[1385]&m[1386]&m[1455]))&~BiasedRNG[986])|((m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1455])|(m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1455])|(~m[1383]&m[1384]&m[1385]&~m[1386]&~m[1455])|(m[1383]&m[1384]&m[1385]&~m[1386]&~m[1455])|(m[1383]&m[1384]&m[1385]&m[1386]&~m[1455])|(m[1383]&m[1384]&~m[1385]&~m[1386]&m[1455])|(m[1383]&~m[1384]&m[1385]&~m[1386]&m[1455])|(~m[1383]&m[1384]&m[1385]&~m[1386]&m[1455])|(m[1383]&m[1384]&m[1385]&~m[1386]&m[1455])|(m[1383]&m[1384]&m[1385]&m[1386]&m[1455]))):InitCond[1932];
    m[1392] = run?((((m[1388]&~m[1389]&~m[1390]&~m[1391]&~m[1460])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1460])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1460])|(m[1388]&m[1389]&~m[1390]&m[1391]&~m[1460])|(m[1388]&~m[1389]&m[1390]&m[1391]&~m[1460])|(~m[1388]&m[1389]&m[1390]&m[1391]&~m[1460]))&BiasedRNG[987])|(((m[1388]&~m[1389]&~m[1390]&~m[1391]&m[1460])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&m[1460])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&m[1460])|(m[1388]&m[1389]&~m[1390]&m[1391]&m[1460])|(m[1388]&~m[1389]&m[1390]&m[1391]&m[1460])|(~m[1388]&m[1389]&m[1390]&m[1391]&m[1460]))&~BiasedRNG[987])|((m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1460])|(m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1460])|(~m[1388]&m[1389]&m[1390]&~m[1391]&~m[1460])|(m[1388]&m[1389]&m[1390]&~m[1391]&~m[1460])|(m[1388]&m[1389]&m[1390]&m[1391]&~m[1460])|(m[1388]&m[1389]&~m[1390]&~m[1391]&m[1460])|(m[1388]&~m[1389]&m[1390]&~m[1391]&m[1460])|(~m[1388]&m[1389]&m[1390]&~m[1391]&m[1460])|(m[1388]&m[1389]&m[1390]&~m[1391]&m[1460])|(m[1388]&m[1389]&m[1390]&m[1391]&m[1460]))):InitCond[1933];
    m[1397] = run?((((m[1393]&~m[1394]&~m[1395]&~m[1396]&~m[1465])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1465])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1465])|(m[1393]&m[1394]&~m[1395]&m[1396]&~m[1465])|(m[1393]&~m[1394]&m[1395]&m[1396]&~m[1465])|(~m[1393]&m[1394]&m[1395]&m[1396]&~m[1465]))&BiasedRNG[988])|(((m[1393]&~m[1394]&~m[1395]&~m[1396]&m[1465])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&m[1465])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&m[1465])|(m[1393]&m[1394]&~m[1395]&m[1396]&m[1465])|(m[1393]&~m[1394]&m[1395]&m[1396]&m[1465])|(~m[1393]&m[1394]&m[1395]&m[1396]&m[1465]))&~BiasedRNG[988])|((m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1465])|(m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1465])|(~m[1393]&m[1394]&m[1395]&~m[1396]&~m[1465])|(m[1393]&m[1394]&m[1395]&~m[1396]&~m[1465])|(m[1393]&m[1394]&m[1395]&m[1396]&~m[1465])|(m[1393]&m[1394]&~m[1395]&~m[1396]&m[1465])|(m[1393]&~m[1394]&m[1395]&~m[1396]&m[1465])|(~m[1393]&m[1394]&m[1395]&~m[1396]&m[1465])|(m[1393]&m[1394]&m[1395]&~m[1396]&m[1465])|(m[1393]&m[1394]&m[1395]&m[1396]&m[1465]))):InitCond[1934];
    m[1402] = run?((((m[1398]&~m[1399]&~m[1400]&~m[1401]&~m[1470])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1470])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1470])|(m[1398]&m[1399]&~m[1400]&m[1401]&~m[1470])|(m[1398]&~m[1399]&m[1400]&m[1401]&~m[1470])|(~m[1398]&m[1399]&m[1400]&m[1401]&~m[1470]))&BiasedRNG[989])|(((m[1398]&~m[1399]&~m[1400]&~m[1401]&m[1470])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&m[1470])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&m[1470])|(m[1398]&m[1399]&~m[1400]&m[1401]&m[1470])|(m[1398]&~m[1399]&m[1400]&m[1401]&m[1470])|(~m[1398]&m[1399]&m[1400]&m[1401]&m[1470]))&~BiasedRNG[989])|((m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1470])|(m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1470])|(~m[1398]&m[1399]&m[1400]&~m[1401]&~m[1470])|(m[1398]&m[1399]&m[1400]&~m[1401]&~m[1470])|(m[1398]&m[1399]&m[1400]&m[1401]&~m[1470])|(m[1398]&m[1399]&~m[1400]&~m[1401]&m[1470])|(m[1398]&~m[1399]&m[1400]&~m[1401]&m[1470])|(~m[1398]&m[1399]&m[1400]&~m[1401]&m[1470])|(m[1398]&m[1399]&m[1400]&~m[1401]&m[1470])|(m[1398]&m[1399]&m[1400]&m[1401]&m[1470]))):InitCond[1935];
    m[1407] = run?((((m[1403]&~m[1404]&~m[1405]&~m[1406]&~m[1475])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1475])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1475])|(m[1403]&m[1404]&~m[1405]&m[1406]&~m[1475])|(m[1403]&~m[1404]&m[1405]&m[1406]&~m[1475])|(~m[1403]&m[1404]&m[1405]&m[1406]&~m[1475]))&BiasedRNG[990])|(((m[1403]&~m[1404]&~m[1405]&~m[1406]&m[1475])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&m[1475])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&m[1475])|(m[1403]&m[1404]&~m[1405]&m[1406]&m[1475])|(m[1403]&~m[1404]&m[1405]&m[1406]&m[1475])|(~m[1403]&m[1404]&m[1405]&m[1406]&m[1475]))&~BiasedRNG[990])|((m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1475])|(m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1475])|(~m[1403]&m[1404]&m[1405]&~m[1406]&~m[1475])|(m[1403]&m[1404]&m[1405]&~m[1406]&~m[1475])|(m[1403]&m[1404]&m[1405]&m[1406]&~m[1475])|(m[1403]&m[1404]&~m[1405]&~m[1406]&m[1475])|(m[1403]&~m[1404]&m[1405]&~m[1406]&m[1475])|(~m[1403]&m[1404]&m[1405]&~m[1406]&m[1475])|(m[1403]&m[1404]&m[1405]&~m[1406]&m[1475])|(m[1403]&m[1404]&m[1405]&m[1406]&m[1475]))):InitCond[1936];
    m[1412] = run?((((m[1408]&~m[1409]&~m[1410]&~m[1411]&~m[1480])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1480])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1480])|(m[1408]&m[1409]&~m[1410]&m[1411]&~m[1480])|(m[1408]&~m[1409]&m[1410]&m[1411]&~m[1480])|(~m[1408]&m[1409]&m[1410]&m[1411]&~m[1480]))&BiasedRNG[991])|(((m[1408]&~m[1409]&~m[1410]&~m[1411]&m[1480])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&m[1480])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&m[1480])|(m[1408]&m[1409]&~m[1410]&m[1411]&m[1480])|(m[1408]&~m[1409]&m[1410]&m[1411]&m[1480])|(~m[1408]&m[1409]&m[1410]&m[1411]&m[1480]))&~BiasedRNG[991])|((m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1480])|(m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1480])|(~m[1408]&m[1409]&m[1410]&~m[1411]&~m[1480])|(m[1408]&m[1409]&m[1410]&~m[1411]&~m[1480])|(m[1408]&m[1409]&m[1410]&m[1411]&~m[1480])|(m[1408]&m[1409]&~m[1410]&~m[1411]&m[1480])|(m[1408]&~m[1409]&m[1410]&~m[1411]&m[1480])|(~m[1408]&m[1409]&m[1410]&~m[1411]&m[1480])|(m[1408]&m[1409]&m[1410]&~m[1411]&m[1480])|(m[1408]&m[1409]&m[1410]&m[1411]&m[1480]))):InitCond[1937];
    m[1417] = run?((((m[1413]&~m[1414]&~m[1415]&~m[1416]&~m[1485])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1485])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1485])|(m[1413]&m[1414]&~m[1415]&m[1416]&~m[1485])|(m[1413]&~m[1414]&m[1415]&m[1416]&~m[1485])|(~m[1413]&m[1414]&m[1415]&m[1416]&~m[1485]))&BiasedRNG[992])|(((m[1413]&~m[1414]&~m[1415]&~m[1416]&m[1485])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&m[1485])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&m[1485])|(m[1413]&m[1414]&~m[1415]&m[1416]&m[1485])|(m[1413]&~m[1414]&m[1415]&m[1416]&m[1485])|(~m[1413]&m[1414]&m[1415]&m[1416]&m[1485]))&~BiasedRNG[992])|((m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1485])|(m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1485])|(~m[1413]&m[1414]&m[1415]&~m[1416]&~m[1485])|(m[1413]&m[1414]&m[1415]&~m[1416]&~m[1485])|(m[1413]&m[1414]&m[1415]&m[1416]&~m[1485])|(m[1413]&m[1414]&~m[1415]&~m[1416]&m[1485])|(m[1413]&~m[1414]&m[1415]&~m[1416]&m[1485])|(~m[1413]&m[1414]&m[1415]&~m[1416]&m[1485])|(m[1413]&m[1414]&m[1415]&~m[1416]&m[1485])|(m[1413]&m[1414]&m[1415]&m[1416]&m[1485]))):InitCond[1938];
    m[1422] = run?((((m[1418]&~m[1419]&~m[1420]&~m[1421]&~m[1490])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1490])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1490])|(m[1418]&m[1419]&~m[1420]&m[1421]&~m[1490])|(m[1418]&~m[1419]&m[1420]&m[1421]&~m[1490])|(~m[1418]&m[1419]&m[1420]&m[1421]&~m[1490]))&BiasedRNG[993])|(((m[1418]&~m[1419]&~m[1420]&~m[1421]&m[1490])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&m[1490])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&m[1490])|(m[1418]&m[1419]&~m[1420]&m[1421]&m[1490])|(m[1418]&~m[1419]&m[1420]&m[1421]&m[1490])|(~m[1418]&m[1419]&m[1420]&m[1421]&m[1490]))&~BiasedRNG[993])|((m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1490])|(m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1490])|(~m[1418]&m[1419]&m[1420]&~m[1421]&~m[1490])|(m[1418]&m[1419]&m[1420]&~m[1421]&~m[1490])|(m[1418]&m[1419]&m[1420]&m[1421]&~m[1490])|(m[1418]&m[1419]&~m[1420]&~m[1421]&m[1490])|(m[1418]&~m[1419]&m[1420]&~m[1421]&m[1490])|(~m[1418]&m[1419]&m[1420]&~m[1421]&m[1490])|(m[1418]&m[1419]&m[1420]&~m[1421]&m[1490])|(m[1418]&m[1419]&m[1420]&m[1421]&m[1490]))):InitCond[1939];
    m[1427] = run?((((m[1423]&~m[1424]&~m[1425]&~m[1426]&~m[1495])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1495])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1495])|(m[1423]&m[1424]&~m[1425]&m[1426]&~m[1495])|(m[1423]&~m[1424]&m[1425]&m[1426]&~m[1495])|(~m[1423]&m[1424]&m[1425]&m[1426]&~m[1495]))&BiasedRNG[994])|(((m[1423]&~m[1424]&~m[1425]&~m[1426]&m[1495])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&m[1495])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&m[1495])|(m[1423]&m[1424]&~m[1425]&m[1426]&m[1495])|(m[1423]&~m[1424]&m[1425]&m[1426]&m[1495])|(~m[1423]&m[1424]&m[1425]&m[1426]&m[1495]))&~BiasedRNG[994])|((m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1495])|(m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1495])|(~m[1423]&m[1424]&m[1425]&~m[1426]&~m[1495])|(m[1423]&m[1424]&m[1425]&~m[1426]&~m[1495])|(m[1423]&m[1424]&m[1425]&m[1426]&~m[1495])|(m[1423]&m[1424]&~m[1425]&~m[1426]&m[1495])|(m[1423]&~m[1424]&m[1425]&~m[1426]&m[1495])|(~m[1423]&m[1424]&m[1425]&~m[1426]&m[1495])|(m[1423]&m[1424]&m[1425]&~m[1426]&m[1495])|(m[1423]&m[1424]&m[1425]&m[1426]&m[1495]))):InitCond[1940];
    m[1432] = run?((((m[1428]&~m[1429]&~m[1430]&~m[1431]&~m[1500])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1500])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1500])|(m[1428]&m[1429]&~m[1430]&m[1431]&~m[1500])|(m[1428]&~m[1429]&m[1430]&m[1431]&~m[1500])|(~m[1428]&m[1429]&m[1430]&m[1431]&~m[1500]))&BiasedRNG[995])|(((m[1428]&~m[1429]&~m[1430]&~m[1431]&m[1500])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&m[1500])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&m[1500])|(m[1428]&m[1429]&~m[1430]&m[1431]&m[1500])|(m[1428]&~m[1429]&m[1430]&m[1431]&m[1500])|(~m[1428]&m[1429]&m[1430]&m[1431]&m[1500]))&~BiasedRNG[995])|((m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1500])|(m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1500])|(~m[1428]&m[1429]&m[1430]&~m[1431]&~m[1500])|(m[1428]&m[1429]&m[1430]&~m[1431]&~m[1500])|(m[1428]&m[1429]&m[1430]&m[1431]&~m[1500])|(m[1428]&m[1429]&~m[1430]&~m[1431]&m[1500])|(m[1428]&~m[1429]&m[1430]&~m[1431]&m[1500])|(~m[1428]&m[1429]&m[1430]&~m[1431]&m[1500])|(m[1428]&m[1429]&m[1430]&~m[1431]&m[1500])|(m[1428]&m[1429]&m[1430]&m[1431]&m[1500]))):InitCond[1941];
    m[1437] = run?((((m[1433]&~m[1434]&~m[1435]&~m[1436]&~m[1505])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1505])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1505])|(m[1433]&m[1434]&~m[1435]&m[1436]&~m[1505])|(m[1433]&~m[1434]&m[1435]&m[1436]&~m[1505])|(~m[1433]&m[1434]&m[1435]&m[1436]&~m[1505]))&BiasedRNG[996])|(((m[1433]&~m[1434]&~m[1435]&~m[1436]&m[1505])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&m[1505])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&m[1505])|(m[1433]&m[1434]&~m[1435]&m[1436]&m[1505])|(m[1433]&~m[1434]&m[1435]&m[1436]&m[1505])|(~m[1433]&m[1434]&m[1435]&m[1436]&m[1505]))&~BiasedRNG[996])|((m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1505])|(m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1505])|(~m[1433]&m[1434]&m[1435]&~m[1436]&~m[1505])|(m[1433]&m[1434]&m[1435]&~m[1436]&~m[1505])|(m[1433]&m[1434]&m[1435]&m[1436]&~m[1505])|(m[1433]&m[1434]&~m[1435]&~m[1436]&m[1505])|(m[1433]&~m[1434]&m[1435]&~m[1436]&m[1505])|(~m[1433]&m[1434]&m[1435]&~m[1436]&m[1505])|(m[1433]&m[1434]&m[1435]&~m[1436]&m[1505])|(m[1433]&m[1434]&m[1435]&m[1436]&m[1505]))):InitCond[1942];
    m[1442] = run?((((m[1438]&~m[1439]&~m[1440]&~m[1441]&~m[1510])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1510])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1510])|(m[1438]&m[1439]&~m[1440]&m[1441]&~m[1510])|(m[1438]&~m[1439]&m[1440]&m[1441]&~m[1510])|(~m[1438]&m[1439]&m[1440]&m[1441]&~m[1510]))&BiasedRNG[997])|(((m[1438]&~m[1439]&~m[1440]&~m[1441]&m[1510])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&m[1510])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&m[1510])|(m[1438]&m[1439]&~m[1440]&m[1441]&m[1510])|(m[1438]&~m[1439]&m[1440]&m[1441]&m[1510])|(~m[1438]&m[1439]&m[1440]&m[1441]&m[1510]))&~BiasedRNG[997])|((m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1510])|(m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1510])|(~m[1438]&m[1439]&m[1440]&~m[1441]&~m[1510])|(m[1438]&m[1439]&m[1440]&~m[1441]&~m[1510])|(m[1438]&m[1439]&m[1440]&m[1441]&~m[1510])|(m[1438]&m[1439]&~m[1440]&~m[1441]&m[1510])|(m[1438]&~m[1439]&m[1440]&~m[1441]&m[1510])|(~m[1438]&m[1439]&m[1440]&~m[1441]&m[1510])|(m[1438]&m[1439]&m[1440]&~m[1441]&m[1510])|(m[1438]&m[1439]&m[1440]&m[1441]&m[1510]))):InitCond[1943];
    m[1447] = run?((((m[1443]&~m[1444]&~m[1445]&~m[1446]&~m[1515])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1515])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1515])|(m[1443]&m[1444]&~m[1445]&m[1446]&~m[1515])|(m[1443]&~m[1444]&m[1445]&m[1446]&~m[1515])|(~m[1443]&m[1444]&m[1445]&m[1446]&~m[1515]))&BiasedRNG[998])|(((m[1443]&~m[1444]&~m[1445]&~m[1446]&m[1515])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&m[1515])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&m[1515])|(m[1443]&m[1444]&~m[1445]&m[1446]&m[1515])|(m[1443]&~m[1444]&m[1445]&m[1446]&m[1515])|(~m[1443]&m[1444]&m[1445]&m[1446]&m[1515]))&~BiasedRNG[998])|((m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1515])|(m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1515])|(~m[1443]&m[1444]&m[1445]&~m[1446]&~m[1515])|(m[1443]&m[1444]&m[1445]&~m[1446]&~m[1515])|(m[1443]&m[1444]&m[1445]&m[1446]&~m[1515])|(m[1443]&m[1444]&~m[1445]&~m[1446]&m[1515])|(m[1443]&~m[1444]&m[1445]&~m[1446]&m[1515])|(~m[1443]&m[1444]&m[1445]&~m[1446]&m[1515])|(m[1443]&m[1444]&m[1445]&~m[1446]&m[1515])|(m[1443]&m[1444]&m[1445]&m[1446]&m[1515]))):InitCond[1944];
    m[1452] = run?((((m[1448]&~m[1449]&~m[1450]&~m[1451]&~m[1520])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1520])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1520])|(m[1448]&m[1449]&~m[1450]&m[1451]&~m[1520])|(m[1448]&~m[1449]&m[1450]&m[1451]&~m[1520])|(~m[1448]&m[1449]&m[1450]&m[1451]&~m[1520]))&BiasedRNG[999])|(((m[1448]&~m[1449]&~m[1450]&~m[1451]&m[1520])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&m[1520])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&m[1520])|(m[1448]&m[1449]&~m[1450]&m[1451]&m[1520])|(m[1448]&~m[1449]&m[1450]&m[1451]&m[1520])|(~m[1448]&m[1449]&m[1450]&m[1451]&m[1520]))&~BiasedRNG[999])|((m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1520])|(m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1520])|(~m[1448]&m[1449]&m[1450]&~m[1451]&~m[1520])|(m[1448]&m[1449]&m[1450]&~m[1451]&~m[1520])|(m[1448]&m[1449]&m[1450]&m[1451]&~m[1520])|(m[1448]&m[1449]&~m[1450]&~m[1451]&m[1520])|(m[1448]&~m[1449]&m[1450]&~m[1451]&m[1520])|(~m[1448]&m[1449]&m[1450]&~m[1451]&m[1520])|(m[1448]&m[1449]&m[1450]&~m[1451]&m[1520])|(m[1448]&m[1449]&m[1450]&m[1451]&m[1520]))):InitCond[1945];
    m[1457] = run?((((m[1453]&~m[1454]&~m[1455]&~m[1456]&~m[1530])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1530])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1530])|(m[1453]&m[1454]&~m[1455]&m[1456]&~m[1530])|(m[1453]&~m[1454]&m[1455]&m[1456]&~m[1530])|(~m[1453]&m[1454]&m[1455]&m[1456]&~m[1530]))&BiasedRNG[1000])|(((m[1453]&~m[1454]&~m[1455]&~m[1456]&m[1530])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&m[1530])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&m[1530])|(m[1453]&m[1454]&~m[1455]&m[1456]&m[1530])|(m[1453]&~m[1454]&m[1455]&m[1456]&m[1530])|(~m[1453]&m[1454]&m[1455]&m[1456]&m[1530]))&~BiasedRNG[1000])|((m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1530])|(m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1530])|(~m[1453]&m[1454]&m[1455]&~m[1456]&~m[1530])|(m[1453]&m[1454]&m[1455]&~m[1456]&~m[1530])|(m[1453]&m[1454]&m[1455]&m[1456]&~m[1530])|(m[1453]&m[1454]&~m[1455]&~m[1456]&m[1530])|(m[1453]&~m[1454]&m[1455]&~m[1456]&m[1530])|(~m[1453]&m[1454]&m[1455]&~m[1456]&m[1530])|(m[1453]&m[1454]&m[1455]&~m[1456]&m[1530])|(m[1453]&m[1454]&m[1455]&m[1456]&m[1530]))):InitCond[1946];
    m[1462] = run?((((m[1458]&~m[1459]&~m[1460]&~m[1461]&~m[1535])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1535])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1535])|(m[1458]&m[1459]&~m[1460]&m[1461]&~m[1535])|(m[1458]&~m[1459]&m[1460]&m[1461]&~m[1535])|(~m[1458]&m[1459]&m[1460]&m[1461]&~m[1535]))&BiasedRNG[1001])|(((m[1458]&~m[1459]&~m[1460]&~m[1461]&m[1535])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&m[1535])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&m[1535])|(m[1458]&m[1459]&~m[1460]&m[1461]&m[1535])|(m[1458]&~m[1459]&m[1460]&m[1461]&m[1535])|(~m[1458]&m[1459]&m[1460]&m[1461]&m[1535]))&~BiasedRNG[1001])|((m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1535])|(m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1535])|(~m[1458]&m[1459]&m[1460]&~m[1461]&~m[1535])|(m[1458]&m[1459]&m[1460]&~m[1461]&~m[1535])|(m[1458]&m[1459]&m[1460]&m[1461]&~m[1535])|(m[1458]&m[1459]&~m[1460]&~m[1461]&m[1535])|(m[1458]&~m[1459]&m[1460]&~m[1461]&m[1535])|(~m[1458]&m[1459]&m[1460]&~m[1461]&m[1535])|(m[1458]&m[1459]&m[1460]&~m[1461]&m[1535])|(m[1458]&m[1459]&m[1460]&m[1461]&m[1535]))):InitCond[1947];
    m[1467] = run?((((m[1463]&~m[1464]&~m[1465]&~m[1466]&~m[1540])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1540])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1540])|(m[1463]&m[1464]&~m[1465]&m[1466]&~m[1540])|(m[1463]&~m[1464]&m[1465]&m[1466]&~m[1540])|(~m[1463]&m[1464]&m[1465]&m[1466]&~m[1540]))&BiasedRNG[1002])|(((m[1463]&~m[1464]&~m[1465]&~m[1466]&m[1540])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&m[1540])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&m[1540])|(m[1463]&m[1464]&~m[1465]&m[1466]&m[1540])|(m[1463]&~m[1464]&m[1465]&m[1466]&m[1540])|(~m[1463]&m[1464]&m[1465]&m[1466]&m[1540]))&~BiasedRNG[1002])|((m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1540])|(m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1540])|(~m[1463]&m[1464]&m[1465]&~m[1466]&~m[1540])|(m[1463]&m[1464]&m[1465]&~m[1466]&~m[1540])|(m[1463]&m[1464]&m[1465]&m[1466]&~m[1540])|(m[1463]&m[1464]&~m[1465]&~m[1466]&m[1540])|(m[1463]&~m[1464]&m[1465]&~m[1466]&m[1540])|(~m[1463]&m[1464]&m[1465]&~m[1466]&m[1540])|(m[1463]&m[1464]&m[1465]&~m[1466]&m[1540])|(m[1463]&m[1464]&m[1465]&m[1466]&m[1540]))):InitCond[1948];
    m[1472] = run?((((m[1468]&~m[1469]&~m[1470]&~m[1471]&~m[1545])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1545])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1545])|(m[1468]&m[1469]&~m[1470]&m[1471]&~m[1545])|(m[1468]&~m[1469]&m[1470]&m[1471]&~m[1545])|(~m[1468]&m[1469]&m[1470]&m[1471]&~m[1545]))&BiasedRNG[1003])|(((m[1468]&~m[1469]&~m[1470]&~m[1471]&m[1545])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&m[1545])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&m[1545])|(m[1468]&m[1469]&~m[1470]&m[1471]&m[1545])|(m[1468]&~m[1469]&m[1470]&m[1471]&m[1545])|(~m[1468]&m[1469]&m[1470]&m[1471]&m[1545]))&~BiasedRNG[1003])|((m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1545])|(m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1545])|(~m[1468]&m[1469]&m[1470]&~m[1471]&~m[1545])|(m[1468]&m[1469]&m[1470]&~m[1471]&~m[1545])|(m[1468]&m[1469]&m[1470]&m[1471]&~m[1545])|(m[1468]&m[1469]&~m[1470]&~m[1471]&m[1545])|(m[1468]&~m[1469]&m[1470]&~m[1471]&m[1545])|(~m[1468]&m[1469]&m[1470]&~m[1471]&m[1545])|(m[1468]&m[1469]&m[1470]&~m[1471]&m[1545])|(m[1468]&m[1469]&m[1470]&m[1471]&m[1545]))):InitCond[1949];
    m[1477] = run?((((m[1473]&~m[1474]&~m[1475]&~m[1476]&~m[1550])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1550])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1550])|(m[1473]&m[1474]&~m[1475]&m[1476]&~m[1550])|(m[1473]&~m[1474]&m[1475]&m[1476]&~m[1550])|(~m[1473]&m[1474]&m[1475]&m[1476]&~m[1550]))&BiasedRNG[1004])|(((m[1473]&~m[1474]&~m[1475]&~m[1476]&m[1550])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&m[1550])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&m[1550])|(m[1473]&m[1474]&~m[1475]&m[1476]&m[1550])|(m[1473]&~m[1474]&m[1475]&m[1476]&m[1550])|(~m[1473]&m[1474]&m[1475]&m[1476]&m[1550]))&~BiasedRNG[1004])|((m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1550])|(m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1550])|(~m[1473]&m[1474]&m[1475]&~m[1476]&~m[1550])|(m[1473]&m[1474]&m[1475]&~m[1476]&~m[1550])|(m[1473]&m[1474]&m[1475]&m[1476]&~m[1550])|(m[1473]&m[1474]&~m[1475]&~m[1476]&m[1550])|(m[1473]&~m[1474]&m[1475]&~m[1476]&m[1550])|(~m[1473]&m[1474]&m[1475]&~m[1476]&m[1550])|(m[1473]&m[1474]&m[1475]&~m[1476]&m[1550])|(m[1473]&m[1474]&m[1475]&m[1476]&m[1550]))):InitCond[1950];
    m[1482] = run?((((m[1478]&~m[1479]&~m[1480]&~m[1481]&~m[1555])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1555])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1555])|(m[1478]&m[1479]&~m[1480]&m[1481]&~m[1555])|(m[1478]&~m[1479]&m[1480]&m[1481]&~m[1555])|(~m[1478]&m[1479]&m[1480]&m[1481]&~m[1555]))&BiasedRNG[1005])|(((m[1478]&~m[1479]&~m[1480]&~m[1481]&m[1555])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&m[1555])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&m[1555])|(m[1478]&m[1479]&~m[1480]&m[1481]&m[1555])|(m[1478]&~m[1479]&m[1480]&m[1481]&m[1555])|(~m[1478]&m[1479]&m[1480]&m[1481]&m[1555]))&~BiasedRNG[1005])|((m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1555])|(m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1555])|(~m[1478]&m[1479]&m[1480]&~m[1481]&~m[1555])|(m[1478]&m[1479]&m[1480]&~m[1481]&~m[1555])|(m[1478]&m[1479]&m[1480]&m[1481]&~m[1555])|(m[1478]&m[1479]&~m[1480]&~m[1481]&m[1555])|(m[1478]&~m[1479]&m[1480]&~m[1481]&m[1555])|(~m[1478]&m[1479]&m[1480]&~m[1481]&m[1555])|(m[1478]&m[1479]&m[1480]&~m[1481]&m[1555])|(m[1478]&m[1479]&m[1480]&m[1481]&m[1555]))):InitCond[1951];
    m[1487] = run?((((m[1483]&~m[1484]&~m[1485]&~m[1486]&~m[1560])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1560])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1560])|(m[1483]&m[1484]&~m[1485]&m[1486]&~m[1560])|(m[1483]&~m[1484]&m[1485]&m[1486]&~m[1560])|(~m[1483]&m[1484]&m[1485]&m[1486]&~m[1560]))&BiasedRNG[1006])|(((m[1483]&~m[1484]&~m[1485]&~m[1486]&m[1560])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&m[1560])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&m[1560])|(m[1483]&m[1484]&~m[1485]&m[1486]&m[1560])|(m[1483]&~m[1484]&m[1485]&m[1486]&m[1560])|(~m[1483]&m[1484]&m[1485]&m[1486]&m[1560]))&~BiasedRNG[1006])|((m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1560])|(m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1560])|(~m[1483]&m[1484]&m[1485]&~m[1486]&~m[1560])|(m[1483]&m[1484]&m[1485]&~m[1486]&~m[1560])|(m[1483]&m[1484]&m[1485]&m[1486]&~m[1560])|(m[1483]&m[1484]&~m[1485]&~m[1486]&m[1560])|(m[1483]&~m[1484]&m[1485]&~m[1486]&m[1560])|(~m[1483]&m[1484]&m[1485]&~m[1486]&m[1560])|(m[1483]&m[1484]&m[1485]&~m[1486]&m[1560])|(m[1483]&m[1484]&m[1485]&m[1486]&m[1560]))):InitCond[1952];
    m[1492] = run?((((m[1488]&~m[1489]&~m[1490]&~m[1491]&~m[1565])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1565])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1565])|(m[1488]&m[1489]&~m[1490]&m[1491]&~m[1565])|(m[1488]&~m[1489]&m[1490]&m[1491]&~m[1565])|(~m[1488]&m[1489]&m[1490]&m[1491]&~m[1565]))&BiasedRNG[1007])|(((m[1488]&~m[1489]&~m[1490]&~m[1491]&m[1565])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&m[1565])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&m[1565])|(m[1488]&m[1489]&~m[1490]&m[1491]&m[1565])|(m[1488]&~m[1489]&m[1490]&m[1491]&m[1565])|(~m[1488]&m[1489]&m[1490]&m[1491]&m[1565]))&~BiasedRNG[1007])|((m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1565])|(m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1565])|(~m[1488]&m[1489]&m[1490]&~m[1491]&~m[1565])|(m[1488]&m[1489]&m[1490]&~m[1491]&~m[1565])|(m[1488]&m[1489]&m[1490]&m[1491]&~m[1565])|(m[1488]&m[1489]&~m[1490]&~m[1491]&m[1565])|(m[1488]&~m[1489]&m[1490]&~m[1491]&m[1565])|(~m[1488]&m[1489]&m[1490]&~m[1491]&m[1565])|(m[1488]&m[1489]&m[1490]&~m[1491]&m[1565])|(m[1488]&m[1489]&m[1490]&m[1491]&m[1565]))):InitCond[1953];
    m[1497] = run?((((m[1493]&~m[1494]&~m[1495]&~m[1496]&~m[1570])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1570])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1570])|(m[1493]&m[1494]&~m[1495]&m[1496]&~m[1570])|(m[1493]&~m[1494]&m[1495]&m[1496]&~m[1570])|(~m[1493]&m[1494]&m[1495]&m[1496]&~m[1570]))&BiasedRNG[1008])|(((m[1493]&~m[1494]&~m[1495]&~m[1496]&m[1570])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&m[1570])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&m[1570])|(m[1493]&m[1494]&~m[1495]&m[1496]&m[1570])|(m[1493]&~m[1494]&m[1495]&m[1496]&m[1570])|(~m[1493]&m[1494]&m[1495]&m[1496]&m[1570]))&~BiasedRNG[1008])|((m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1570])|(m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1570])|(~m[1493]&m[1494]&m[1495]&~m[1496]&~m[1570])|(m[1493]&m[1494]&m[1495]&~m[1496]&~m[1570])|(m[1493]&m[1494]&m[1495]&m[1496]&~m[1570])|(m[1493]&m[1494]&~m[1495]&~m[1496]&m[1570])|(m[1493]&~m[1494]&m[1495]&~m[1496]&m[1570])|(~m[1493]&m[1494]&m[1495]&~m[1496]&m[1570])|(m[1493]&m[1494]&m[1495]&~m[1496]&m[1570])|(m[1493]&m[1494]&m[1495]&m[1496]&m[1570]))):InitCond[1954];
    m[1502] = run?((((m[1498]&~m[1499]&~m[1500]&~m[1501]&~m[1575])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1575])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1575])|(m[1498]&m[1499]&~m[1500]&m[1501]&~m[1575])|(m[1498]&~m[1499]&m[1500]&m[1501]&~m[1575])|(~m[1498]&m[1499]&m[1500]&m[1501]&~m[1575]))&BiasedRNG[1009])|(((m[1498]&~m[1499]&~m[1500]&~m[1501]&m[1575])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&m[1575])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&m[1575])|(m[1498]&m[1499]&~m[1500]&m[1501]&m[1575])|(m[1498]&~m[1499]&m[1500]&m[1501]&m[1575])|(~m[1498]&m[1499]&m[1500]&m[1501]&m[1575]))&~BiasedRNG[1009])|((m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1575])|(m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1575])|(~m[1498]&m[1499]&m[1500]&~m[1501]&~m[1575])|(m[1498]&m[1499]&m[1500]&~m[1501]&~m[1575])|(m[1498]&m[1499]&m[1500]&m[1501]&~m[1575])|(m[1498]&m[1499]&~m[1500]&~m[1501]&m[1575])|(m[1498]&~m[1499]&m[1500]&~m[1501]&m[1575])|(~m[1498]&m[1499]&m[1500]&~m[1501]&m[1575])|(m[1498]&m[1499]&m[1500]&~m[1501]&m[1575])|(m[1498]&m[1499]&m[1500]&m[1501]&m[1575]))):InitCond[1955];
    m[1507] = run?((((m[1503]&~m[1504]&~m[1505]&~m[1506]&~m[1580])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1580])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1580])|(m[1503]&m[1504]&~m[1505]&m[1506]&~m[1580])|(m[1503]&~m[1504]&m[1505]&m[1506]&~m[1580])|(~m[1503]&m[1504]&m[1505]&m[1506]&~m[1580]))&BiasedRNG[1010])|(((m[1503]&~m[1504]&~m[1505]&~m[1506]&m[1580])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&m[1580])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&m[1580])|(m[1503]&m[1504]&~m[1505]&m[1506]&m[1580])|(m[1503]&~m[1504]&m[1505]&m[1506]&m[1580])|(~m[1503]&m[1504]&m[1505]&m[1506]&m[1580]))&~BiasedRNG[1010])|((m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1580])|(m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1580])|(~m[1503]&m[1504]&m[1505]&~m[1506]&~m[1580])|(m[1503]&m[1504]&m[1505]&~m[1506]&~m[1580])|(m[1503]&m[1504]&m[1505]&m[1506]&~m[1580])|(m[1503]&m[1504]&~m[1505]&~m[1506]&m[1580])|(m[1503]&~m[1504]&m[1505]&~m[1506]&m[1580])|(~m[1503]&m[1504]&m[1505]&~m[1506]&m[1580])|(m[1503]&m[1504]&m[1505]&~m[1506]&m[1580])|(m[1503]&m[1504]&m[1505]&m[1506]&m[1580]))):InitCond[1956];
    m[1512] = run?((((m[1508]&~m[1509]&~m[1510]&~m[1511]&~m[1585])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1585])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1585])|(m[1508]&m[1509]&~m[1510]&m[1511]&~m[1585])|(m[1508]&~m[1509]&m[1510]&m[1511]&~m[1585])|(~m[1508]&m[1509]&m[1510]&m[1511]&~m[1585]))&BiasedRNG[1011])|(((m[1508]&~m[1509]&~m[1510]&~m[1511]&m[1585])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&m[1585])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&m[1585])|(m[1508]&m[1509]&~m[1510]&m[1511]&m[1585])|(m[1508]&~m[1509]&m[1510]&m[1511]&m[1585])|(~m[1508]&m[1509]&m[1510]&m[1511]&m[1585]))&~BiasedRNG[1011])|((m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1585])|(m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1585])|(~m[1508]&m[1509]&m[1510]&~m[1511]&~m[1585])|(m[1508]&m[1509]&m[1510]&~m[1511]&~m[1585])|(m[1508]&m[1509]&m[1510]&m[1511]&~m[1585])|(m[1508]&m[1509]&~m[1510]&~m[1511]&m[1585])|(m[1508]&~m[1509]&m[1510]&~m[1511]&m[1585])|(~m[1508]&m[1509]&m[1510]&~m[1511]&m[1585])|(m[1508]&m[1509]&m[1510]&~m[1511]&m[1585])|(m[1508]&m[1509]&m[1510]&m[1511]&m[1585]))):InitCond[1957];
    m[1517] = run?((((m[1513]&~m[1514]&~m[1515]&~m[1516]&~m[1590])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1590])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1590])|(m[1513]&m[1514]&~m[1515]&m[1516]&~m[1590])|(m[1513]&~m[1514]&m[1515]&m[1516]&~m[1590])|(~m[1513]&m[1514]&m[1515]&m[1516]&~m[1590]))&BiasedRNG[1012])|(((m[1513]&~m[1514]&~m[1515]&~m[1516]&m[1590])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&m[1590])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&m[1590])|(m[1513]&m[1514]&~m[1515]&m[1516]&m[1590])|(m[1513]&~m[1514]&m[1515]&m[1516]&m[1590])|(~m[1513]&m[1514]&m[1515]&m[1516]&m[1590]))&~BiasedRNG[1012])|((m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1590])|(m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1590])|(~m[1513]&m[1514]&m[1515]&~m[1516]&~m[1590])|(m[1513]&m[1514]&m[1515]&~m[1516]&~m[1590])|(m[1513]&m[1514]&m[1515]&m[1516]&~m[1590])|(m[1513]&m[1514]&~m[1515]&~m[1516]&m[1590])|(m[1513]&~m[1514]&m[1515]&~m[1516]&m[1590])|(~m[1513]&m[1514]&m[1515]&~m[1516]&m[1590])|(m[1513]&m[1514]&m[1515]&~m[1516]&m[1590])|(m[1513]&m[1514]&m[1515]&m[1516]&m[1590]))):InitCond[1958];
    m[1522] = run?((((m[1518]&~m[1519]&~m[1520]&~m[1521]&~m[1595])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1595])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1595])|(m[1518]&m[1519]&~m[1520]&m[1521]&~m[1595])|(m[1518]&~m[1519]&m[1520]&m[1521]&~m[1595])|(~m[1518]&m[1519]&m[1520]&m[1521]&~m[1595]))&BiasedRNG[1013])|(((m[1518]&~m[1519]&~m[1520]&~m[1521]&m[1595])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&m[1595])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&m[1595])|(m[1518]&m[1519]&~m[1520]&m[1521]&m[1595])|(m[1518]&~m[1519]&m[1520]&m[1521]&m[1595])|(~m[1518]&m[1519]&m[1520]&m[1521]&m[1595]))&~BiasedRNG[1013])|((m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1595])|(m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1595])|(~m[1518]&m[1519]&m[1520]&~m[1521]&~m[1595])|(m[1518]&m[1519]&m[1520]&~m[1521]&~m[1595])|(m[1518]&m[1519]&m[1520]&m[1521]&~m[1595])|(m[1518]&m[1519]&~m[1520]&~m[1521]&m[1595])|(m[1518]&~m[1519]&m[1520]&~m[1521]&m[1595])|(~m[1518]&m[1519]&m[1520]&~m[1521]&m[1595])|(m[1518]&m[1519]&m[1520]&~m[1521]&m[1595])|(m[1518]&m[1519]&m[1520]&m[1521]&m[1595]))):InitCond[1959];
    m[1527] = run?((((m[1523]&~m[1524]&~m[1525]&~m[1526]&~m[1600])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1600])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1600])|(m[1523]&m[1524]&~m[1525]&m[1526]&~m[1600])|(m[1523]&~m[1524]&m[1525]&m[1526]&~m[1600])|(~m[1523]&m[1524]&m[1525]&m[1526]&~m[1600]))&BiasedRNG[1014])|(((m[1523]&~m[1524]&~m[1525]&~m[1526]&m[1600])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&m[1600])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&m[1600])|(m[1523]&m[1524]&~m[1525]&m[1526]&m[1600])|(m[1523]&~m[1524]&m[1525]&m[1526]&m[1600])|(~m[1523]&m[1524]&m[1525]&m[1526]&m[1600]))&~BiasedRNG[1014])|((m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1600])|(m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1600])|(~m[1523]&m[1524]&m[1525]&~m[1526]&~m[1600])|(m[1523]&m[1524]&m[1525]&~m[1526]&~m[1600])|(m[1523]&m[1524]&m[1525]&m[1526]&~m[1600])|(m[1523]&m[1524]&~m[1525]&~m[1526]&m[1600])|(m[1523]&~m[1524]&m[1525]&~m[1526]&m[1600])|(~m[1523]&m[1524]&m[1525]&~m[1526]&m[1600])|(m[1523]&m[1524]&m[1525]&~m[1526]&m[1600])|(m[1523]&m[1524]&m[1525]&m[1526]&m[1600]))):InitCond[1960];
    m[1532] = run?((((m[1528]&~m[1529]&~m[1530]&~m[1531]&~m[1603])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1603])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1603])|(m[1528]&m[1529]&~m[1530]&m[1531]&~m[1603])|(m[1528]&~m[1529]&m[1530]&m[1531]&~m[1603])|(~m[1528]&m[1529]&m[1530]&m[1531]&~m[1603]))&BiasedRNG[1015])|(((m[1528]&~m[1529]&~m[1530]&~m[1531]&m[1603])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&m[1603])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&m[1603])|(m[1528]&m[1529]&~m[1530]&m[1531]&m[1603])|(m[1528]&~m[1529]&m[1530]&m[1531]&m[1603])|(~m[1528]&m[1529]&m[1530]&m[1531]&m[1603]))&~BiasedRNG[1015])|((m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1603])|(m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1603])|(~m[1528]&m[1529]&m[1530]&~m[1531]&~m[1603])|(m[1528]&m[1529]&m[1530]&~m[1531]&~m[1603])|(m[1528]&m[1529]&m[1530]&m[1531]&~m[1603])|(m[1528]&m[1529]&~m[1530]&~m[1531]&m[1603])|(m[1528]&~m[1529]&m[1530]&~m[1531]&m[1603])|(~m[1528]&m[1529]&m[1530]&~m[1531]&m[1603])|(m[1528]&m[1529]&m[1530]&~m[1531]&m[1603])|(m[1528]&m[1529]&m[1530]&m[1531]&m[1603]))):InitCond[1961];
    m[1537] = run?((((m[1533]&~m[1534]&~m[1535]&~m[1536]&~m[1605])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1605])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1605])|(m[1533]&m[1534]&~m[1535]&m[1536]&~m[1605])|(m[1533]&~m[1534]&m[1535]&m[1536]&~m[1605])|(~m[1533]&m[1534]&m[1535]&m[1536]&~m[1605]))&BiasedRNG[1016])|(((m[1533]&~m[1534]&~m[1535]&~m[1536]&m[1605])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&m[1605])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&m[1605])|(m[1533]&m[1534]&~m[1535]&m[1536]&m[1605])|(m[1533]&~m[1534]&m[1535]&m[1536]&m[1605])|(~m[1533]&m[1534]&m[1535]&m[1536]&m[1605]))&~BiasedRNG[1016])|((m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1605])|(m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1605])|(~m[1533]&m[1534]&m[1535]&~m[1536]&~m[1605])|(m[1533]&m[1534]&m[1535]&~m[1536]&~m[1605])|(m[1533]&m[1534]&m[1535]&m[1536]&~m[1605])|(m[1533]&m[1534]&~m[1535]&~m[1536]&m[1605])|(m[1533]&~m[1534]&m[1535]&~m[1536]&m[1605])|(~m[1533]&m[1534]&m[1535]&~m[1536]&m[1605])|(m[1533]&m[1534]&m[1535]&~m[1536]&m[1605])|(m[1533]&m[1534]&m[1535]&m[1536]&m[1605]))):InitCond[1962];
    m[1542] = run?((((m[1538]&~m[1539]&~m[1540]&~m[1541]&~m[1610])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1610])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1610])|(m[1538]&m[1539]&~m[1540]&m[1541]&~m[1610])|(m[1538]&~m[1539]&m[1540]&m[1541]&~m[1610])|(~m[1538]&m[1539]&m[1540]&m[1541]&~m[1610]))&BiasedRNG[1017])|(((m[1538]&~m[1539]&~m[1540]&~m[1541]&m[1610])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&m[1610])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&m[1610])|(m[1538]&m[1539]&~m[1540]&m[1541]&m[1610])|(m[1538]&~m[1539]&m[1540]&m[1541]&m[1610])|(~m[1538]&m[1539]&m[1540]&m[1541]&m[1610]))&~BiasedRNG[1017])|((m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1610])|(m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1610])|(~m[1538]&m[1539]&m[1540]&~m[1541]&~m[1610])|(m[1538]&m[1539]&m[1540]&~m[1541]&~m[1610])|(m[1538]&m[1539]&m[1540]&m[1541]&~m[1610])|(m[1538]&m[1539]&~m[1540]&~m[1541]&m[1610])|(m[1538]&~m[1539]&m[1540]&~m[1541]&m[1610])|(~m[1538]&m[1539]&m[1540]&~m[1541]&m[1610])|(m[1538]&m[1539]&m[1540]&~m[1541]&m[1610])|(m[1538]&m[1539]&m[1540]&m[1541]&m[1610]))):InitCond[1963];
    m[1547] = run?((((m[1543]&~m[1544]&~m[1545]&~m[1546]&~m[1615])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1615])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1615])|(m[1543]&m[1544]&~m[1545]&m[1546]&~m[1615])|(m[1543]&~m[1544]&m[1545]&m[1546]&~m[1615])|(~m[1543]&m[1544]&m[1545]&m[1546]&~m[1615]))&BiasedRNG[1018])|(((m[1543]&~m[1544]&~m[1545]&~m[1546]&m[1615])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&m[1615])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&m[1615])|(m[1543]&m[1544]&~m[1545]&m[1546]&m[1615])|(m[1543]&~m[1544]&m[1545]&m[1546]&m[1615])|(~m[1543]&m[1544]&m[1545]&m[1546]&m[1615]))&~BiasedRNG[1018])|((m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1615])|(m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1615])|(~m[1543]&m[1544]&m[1545]&~m[1546]&~m[1615])|(m[1543]&m[1544]&m[1545]&~m[1546]&~m[1615])|(m[1543]&m[1544]&m[1545]&m[1546]&~m[1615])|(m[1543]&m[1544]&~m[1545]&~m[1546]&m[1615])|(m[1543]&~m[1544]&m[1545]&~m[1546]&m[1615])|(~m[1543]&m[1544]&m[1545]&~m[1546]&m[1615])|(m[1543]&m[1544]&m[1545]&~m[1546]&m[1615])|(m[1543]&m[1544]&m[1545]&m[1546]&m[1615]))):InitCond[1964];
    m[1552] = run?((((m[1548]&~m[1549]&~m[1550]&~m[1551]&~m[1620])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1620])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1620])|(m[1548]&m[1549]&~m[1550]&m[1551]&~m[1620])|(m[1548]&~m[1549]&m[1550]&m[1551]&~m[1620])|(~m[1548]&m[1549]&m[1550]&m[1551]&~m[1620]))&BiasedRNG[1019])|(((m[1548]&~m[1549]&~m[1550]&~m[1551]&m[1620])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&m[1620])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&m[1620])|(m[1548]&m[1549]&~m[1550]&m[1551]&m[1620])|(m[1548]&~m[1549]&m[1550]&m[1551]&m[1620])|(~m[1548]&m[1549]&m[1550]&m[1551]&m[1620]))&~BiasedRNG[1019])|((m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1620])|(m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1620])|(~m[1548]&m[1549]&m[1550]&~m[1551]&~m[1620])|(m[1548]&m[1549]&m[1550]&~m[1551]&~m[1620])|(m[1548]&m[1549]&m[1550]&m[1551]&~m[1620])|(m[1548]&m[1549]&~m[1550]&~m[1551]&m[1620])|(m[1548]&~m[1549]&m[1550]&~m[1551]&m[1620])|(~m[1548]&m[1549]&m[1550]&~m[1551]&m[1620])|(m[1548]&m[1549]&m[1550]&~m[1551]&m[1620])|(m[1548]&m[1549]&m[1550]&m[1551]&m[1620]))):InitCond[1965];
    m[1557] = run?((((m[1553]&~m[1554]&~m[1555]&~m[1556]&~m[1625])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1625])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1625])|(m[1553]&m[1554]&~m[1555]&m[1556]&~m[1625])|(m[1553]&~m[1554]&m[1555]&m[1556]&~m[1625])|(~m[1553]&m[1554]&m[1555]&m[1556]&~m[1625]))&BiasedRNG[1020])|(((m[1553]&~m[1554]&~m[1555]&~m[1556]&m[1625])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&m[1625])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&m[1625])|(m[1553]&m[1554]&~m[1555]&m[1556]&m[1625])|(m[1553]&~m[1554]&m[1555]&m[1556]&m[1625])|(~m[1553]&m[1554]&m[1555]&m[1556]&m[1625]))&~BiasedRNG[1020])|((m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1625])|(m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1625])|(~m[1553]&m[1554]&m[1555]&~m[1556]&~m[1625])|(m[1553]&m[1554]&m[1555]&~m[1556]&~m[1625])|(m[1553]&m[1554]&m[1555]&m[1556]&~m[1625])|(m[1553]&m[1554]&~m[1555]&~m[1556]&m[1625])|(m[1553]&~m[1554]&m[1555]&~m[1556]&m[1625])|(~m[1553]&m[1554]&m[1555]&~m[1556]&m[1625])|(m[1553]&m[1554]&m[1555]&~m[1556]&m[1625])|(m[1553]&m[1554]&m[1555]&m[1556]&m[1625]))):InitCond[1966];
    m[1562] = run?((((m[1558]&~m[1559]&~m[1560]&~m[1561]&~m[1630])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1630])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1630])|(m[1558]&m[1559]&~m[1560]&m[1561]&~m[1630])|(m[1558]&~m[1559]&m[1560]&m[1561]&~m[1630])|(~m[1558]&m[1559]&m[1560]&m[1561]&~m[1630]))&BiasedRNG[1021])|(((m[1558]&~m[1559]&~m[1560]&~m[1561]&m[1630])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&m[1630])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&m[1630])|(m[1558]&m[1559]&~m[1560]&m[1561]&m[1630])|(m[1558]&~m[1559]&m[1560]&m[1561]&m[1630])|(~m[1558]&m[1559]&m[1560]&m[1561]&m[1630]))&~BiasedRNG[1021])|((m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1630])|(m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1630])|(~m[1558]&m[1559]&m[1560]&~m[1561]&~m[1630])|(m[1558]&m[1559]&m[1560]&~m[1561]&~m[1630])|(m[1558]&m[1559]&m[1560]&m[1561]&~m[1630])|(m[1558]&m[1559]&~m[1560]&~m[1561]&m[1630])|(m[1558]&~m[1559]&m[1560]&~m[1561]&m[1630])|(~m[1558]&m[1559]&m[1560]&~m[1561]&m[1630])|(m[1558]&m[1559]&m[1560]&~m[1561]&m[1630])|(m[1558]&m[1559]&m[1560]&m[1561]&m[1630]))):InitCond[1967];
    m[1567] = run?((((m[1563]&~m[1564]&~m[1565]&~m[1566]&~m[1635])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1635])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1635])|(m[1563]&m[1564]&~m[1565]&m[1566]&~m[1635])|(m[1563]&~m[1564]&m[1565]&m[1566]&~m[1635])|(~m[1563]&m[1564]&m[1565]&m[1566]&~m[1635]))&BiasedRNG[1022])|(((m[1563]&~m[1564]&~m[1565]&~m[1566]&m[1635])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&m[1635])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&m[1635])|(m[1563]&m[1564]&~m[1565]&m[1566]&m[1635])|(m[1563]&~m[1564]&m[1565]&m[1566]&m[1635])|(~m[1563]&m[1564]&m[1565]&m[1566]&m[1635]))&~BiasedRNG[1022])|((m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1635])|(m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1635])|(~m[1563]&m[1564]&m[1565]&~m[1566]&~m[1635])|(m[1563]&m[1564]&m[1565]&~m[1566]&~m[1635])|(m[1563]&m[1564]&m[1565]&m[1566]&~m[1635])|(m[1563]&m[1564]&~m[1565]&~m[1566]&m[1635])|(m[1563]&~m[1564]&m[1565]&~m[1566]&m[1635])|(~m[1563]&m[1564]&m[1565]&~m[1566]&m[1635])|(m[1563]&m[1564]&m[1565]&~m[1566]&m[1635])|(m[1563]&m[1564]&m[1565]&m[1566]&m[1635]))):InitCond[1968];
    m[1572] = run?((((m[1568]&~m[1569]&~m[1570]&~m[1571]&~m[1640])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1640])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1640])|(m[1568]&m[1569]&~m[1570]&m[1571]&~m[1640])|(m[1568]&~m[1569]&m[1570]&m[1571]&~m[1640])|(~m[1568]&m[1569]&m[1570]&m[1571]&~m[1640]))&BiasedRNG[1023])|(((m[1568]&~m[1569]&~m[1570]&~m[1571]&m[1640])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&m[1640])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&m[1640])|(m[1568]&m[1569]&~m[1570]&m[1571]&m[1640])|(m[1568]&~m[1569]&m[1570]&m[1571]&m[1640])|(~m[1568]&m[1569]&m[1570]&m[1571]&m[1640]))&~BiasedRNG[1023])|((m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1640])|(m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1640])|(~m[1568]&m[1569]&m[1570]&~m[1571]&~m[1640])|(m[1568]&m[1569]&m[1570]&~m[1571]&~m[1640])|(m[1568]&m[1569]&m[1570]&m[1571]&~m[1640])|(m[1568]&m[1569]&~m[1570]&~m[1571]&m[1640])|(m[1568]&~m[1569]&m[1570]&~m[1571]&m[1640])|(~m[1568]&m[1569]&m[1570]&~m[1571]&m[1640])|(m[1568]&m[1569]&m[1570]&~m[1571]&m[1640])|(m[1568]&m[1569]&m[1570]&m[1571]&m[1640]))):InitCond[1969];
    m[1577] = run?((((m[1573]&~m[1574]&~m[1575]&~m[1576]&~m[1645])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1645])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1645])|(m[1573]&m[1574]&~m[1575]&m[1576]&~m[1645])|(m[1573]&~m[1574]&m[1575]&m[1576]&~m[1645])|(~m[1573]&m[1574]&m[1575]&m[1576]&~m[1645]))&BiasedRNG[1024])|(((m[1573]&~m[1574]&~m[1575]&~m[1576]&m[1645])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&m[1645])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&m[1645])|(m[1573]&m[1574]&~m[1575]&m[1576]&m[1645])|(m[1573]&~m[1574]&m[1575]&m[1576]&m[1645])|(~m[1573]&m[1574]&m[1575]&m[1576]&m[1645]))&~BiasedRNG[1024])|((m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1645])|(m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1645])|(~m[1573]&m[1574]&m[1575]&~m[1576]&~m[1645])|(m[1573]&m[1574]&m[1575]&~m[1576]&~m[1645])|(m[1573]&m[1574]&m[1575]&m[1576]&~m[1645])|(m[1573]&m[1574]&~m[1575]&~m[1576]&m[1645])|(m[1573]&~m[1574]&m[1575]&~m[1576]&m[1645])|(~m[1573]&m[1574]&m[1575]&~m[1576]&m[1645])|(m[1573]&m[1574]&m[1575]&~m[1576]&m[1645])|(m[1573]&m[1574]&m[1575]&m[1576]&m[1645]))):InitCond[1970];
    m[1582] = run?((((m[1578]&~m[1579]&~m[1580]&~m[1581]&~m[1650])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1650])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1650])|(m[1578]&m[1579]&~m[1580]&m[1581]&~m[1650])|(m[1578]&~m[1579]&m[1580]&m[1581]&~m[1650])|(~m[1578]&m[1579]&m[1580]&m[1581]&~m[1650]))&BiasedRNG[1025])|(((m[1578]&~m[1579]&~m[1580]&~m[1581]&m[1650])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&m[1650])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&m[1650])|(m[1578]&m[1579]&~m[1580]&m[1581]&m[1650])|(m[1578]&~m[1579]&m[1580]&m[1581]&m[1650])|(~m[1578]&m[1579]&m[1580]&m[1581]&m[1650]))&~BiasedRNG[1025])|((m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1650])|(m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1650])|(~m[1578]&m[1579]&m[1580]&~m[1581]&~m[1650])|(m[1578]&m[1579]&m[1580]&~m[1581]&~m[1650])|(m[1578]&m[1579]&m[1580]&m[1581]&~m[1650])|(m[1578]&m[1579]&~m[1580]&~m[1581]&m[1650])|(m[1578]&~m[1579]&m[1580]&~m[1581]&m[1650])|(~m[1578]&m[1579]&m[1580]&~m[1581]&m[1650])|(m[1578]&m[1579]&m[1580]&~m[1581]&m[1650])|(m[1578]&m[1579]&m[1580]&m[1581]&m[1650]))):InitCond[1971];
    m[1587] = run?((((m[1583]&~m[1584]&~m[1585]&~m[1586]&~m[1655])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1655])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1655])|(m[1583]&m[1584]&~m[1585]&m[1586]&~m[1655])|(m[1583]&~m[1584]&m[1585]&m[1586]&~m[1655])|(~m[1583]&m[1584]&m[1585]&m[1586]&~m[1655]))&BiasedRNG[1026])|(((m[1583]&~m[1584]&~m[1585]&~m[1586]&m[1655])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&m[1655])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&m[1655])|(m[1583]&m[1584]&~m[1585]&m[1586]&m[1655])|(m[1583]&~m[1584]&m[1585]&m[1586]&m[1655])|(~m[1583]&m[1584]&m[1585]&m[1586]&m[1655]))&~BiasedRNG[1026])|((m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1655])|(m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1655])|(~m[1583]&m[1584]&m[1585]&~m[1586]&~m[1655])|(m[1583]&m[1584]&m[1585]&~m[1586]&~m[1655])|(m[1583]&m[1584]&m[1585]&m[1586]&~m[1655])|(m[1583]&m[1584]&~m[1585]&~m[1586]&m[1655])|(m[1583]&~m[1584]&m[1585]&~m[1586]&m[1655])|(~m[1583]&m[1584]&m[1585]&~m[1586]&m[1655])|(m[1583]&m[1584]&m[1585]&~m[1586]&m[1655])|(m[1583]&m[1584]&m[1585]&m[1586]&m[1655]))):InitCond[1972];
    m[1592] = run?((((m[1588]&~m[1589]&~m[1590]&~m[1591]&~m[1660])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1660])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1660])|(m[1588]&m[1589]&~m[1590]&m[1591]&~m[1660])|(m[1588]&~m[1589]&m[1590]&m[1591]&~m[1660])|(~m[1588]&m[1589]&m[1590]&m[1591]&~m[1660]))&BiasedRNG[1027])|(((m[1588]&~m[1589]&~m[1590]&~m[1591]&m[1660])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&m[1660])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&m[1660])|(m[1588]&m[1589]&~m[1590]&m[1591]&m[1660])|(m[1588]&~m[1589]&m[1590]&m[1591]&m[1660])|(~m[1588]&m[1589]&m[1590]&m[1591]&m[1660]))&~BiasedRNG[1027])|((m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1660])|(m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1660])|(~m[1588]&m[1589]&m[1590]&~m[1591]&~m[1660])|(m[1588]&m[1589]&m[1590]&~m[1591]&~m[1660])|(m[1588]&m[1589]&m[1590]&m[1591]&~m[1660])|(m[1588]&m[1589]&~m[1590]&~m[1591]&m[1660])|(m[1588]&~m[1589]&m[1590]&~m[1591]&m[1660])|(~m[1588]&m[1589]&m[1590]&~m[1591]&m[1660])|(m[1588]&m[1589]&m[1590]&~m[1591]&m[1660])|(m[1588]&m[1589]&m[1590]&m[1591]&m[1660]))):InitCond[1973];
    m[1597] = run?((((m[1593]&~m[1594]&~m[1595]&~m[1596]&~m[1665])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1665])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1665])|(m[1593]&m[1594]&~m[1595]&m[1596]&~m[1665])|(m[1593]&~m[1594]&m[1595]&m[1596]&~m[1665])|(~m[1593]&m[1594]&m[1595]&m[1596]&~m[1665]))&BiasedRNG[1028])|(((m[1593]&~m[1594]&~m[1595]&~m[1596]&m[1665])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&m[1665])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&m[1665])|(m[1593]&m[1594]&~m[1595]&m[1596]&m[1665])|(m[1593]&~m[1594]&m[1595]&m[1596]&m[1665])|(~m[1593]&m[1594]&m[1595]&m[1596]&m[1665]))&~BiasedRNG[1028])|((m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1665])|(m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1665])|(~m[1593]&m[1594]&m[1595]&~m[1596]&~m[1665])|(m[1593]&m[1594]&m[1595]&~m[1596]&~m[1665])|(m[1593]&m[1594]&m[1595]&m[1596]&~m[1665])|(m[1593]&m[1594]&~m[1595]&~m[1596]&m[1665])|(m[1593]&~m[1594]&m[1595]&~m[1596]&m[1665])|(~m[1593]&m[1594]&m[1595]&~m[1596]&m[1665])|(m[1593]&m[1594]&m[1595]&~m[1596]&m[1665])|(m[1593]&m[1594]&m[1595]&m[1596]&m[1665]))):InitCond[1974];
    m[1602] = run?((((m[1598]&~m[1599]&~m[1600]&~m[1601]&~m[1670])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1670])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1670])|(m[1598]&m[1599]&~m[1600]&m[1601]&~m[1670])|(m[1598]&~m[1599]&m[1600]&m[1601]&~m[1670])|(~m[1598]&m[1599]&m[1600]&m[1601]&~m[1670]))&BiasedRNG[1029])|(((m[1598]&~m[1599]&~m[1600]&~m[1601]&m[1670])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&m[1670])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&m[1670])|(m[1598]&m[1599]&~m[1600]&m[1601]&m[1670])|(m[1598]&~m[1599]&m[1600]&m[1601]&m[1670])|(~m[1598]&m[1599]&m[1600]&m[1601]&m[1670]))&~BiasedRNG[1029])|((m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1670])|(m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1670])|(~m[1598]&m[1599]&m[1600]&~m[1601]&~m[1670])|(m[1598]&m[1599]&m[1600]&~m[1601]&~m[1670])|(m[1598]&m[1599]&m[1600]&m[1601]&~m[1670])|(m[1598]&m[1599]&~m[1600]&~m[1601]&m[1670])|(m[1598]&~m[1599]&m[1600]&~m[1601]&m[1670])|(~m[1598]&m[1599]&m[1600]&~m[1601]&m[1670])|(m[1598]&m[1599]&m[1600]&~m[1601]&m[1670])|(m[1598]&m[1599]&m[1600]&m[1601]&m[1670]))):InitCond[1975];
    m[1607] = run?((((m[1603]&~m[1604]&~m[1605]&~m[1606]&~m[1673])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1673])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1673])|(m[1603]&m[1604]&~m[1605]&m[1606]&~m[1673])|(m[1603]&~m[1604]&m[1605]&m[1606]&~m[1673])|(~m[1603]&m[1604]&m[1605]&m[1606]&~m[1673]))&BiasedRNG[1030])|(((m[1603]&~m[1604]&~m[1605]&~m[1606]&m[1673])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&m[1673])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&m[1673])|(m[1603]&m[1604]&~m[1605]&m[1606]&m[1673])|(m[1603]&~m[1604]&m[1605]&m[1606]&m[1673])|(~m[1603]&m[1604]&m[1605]&m[1606]&m[1673]))&~BiasedRNG[1030])|((m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1673])|(m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1673])|(~m[1603]&m[1604]&m[1605]&~m[1606]&~m[1673])|(m[1603]&m[1604]&m[1605]&~m[1606]&~m[1673])|(m[1603]&m[1604]&m[1605]&m[1606]&~m[1673])|(m[1603]&m[1604]&~m[1605]&~m[1606]&m[1673])|(m[1603]&~m[1604]&m[1605]&~m[1606]&m[1673])|(~m[1603]&m[1604]&m[1605]&~m[1606]&m[1673])|(m[1603]&m[1604]&m[1605]&~m[1606]&m[1673])|(m[1603]&m[1604]&m[1605]&m[1606]&m[1673]))):InitCond[1976];
    m[1612] = run?((((m[1608]&~m[1609]&~m[1610]&~m[1611]&~m[1675])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1675])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1675])|(m[1608]&m[1609]&~m[1610]&m[1611]&~m[1675])|(m[1608]&~m[1609]&m[1610]&m[1611]&~m[1675])|(~m[1608]&m[1609]&m[1610]&m[1611]&~m[1675]))&BiasedRNG[1031])|(((m[1608]&~m[1609]&~m[1610]&~m[1611]&m[1675])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&m[1675])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&m[1675])|(m[1608]&m[1609]&~m[1610]&m[1611]&m[1675])|(m[1608]&~m[1609]&m[1610]&m[1611]&m[1675])|(~m[1608]&m[1609]&m[1610]&m[1611]&m[1675]))&~BiasedRNG[1031])|((m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1675])|(m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1675])|(~m[1608]&m[1609]&m[1610]&~m[1611]&~m[1675])|(m[1608]&m[1609]&m[1610]&~m[1611]&~m[1675])|(m[1608]&m[1609]&m[1610]&m[1611]&~m[1675])|(m[1608]&m[1609]&~m[1610]&~m[1611]&m[1675])|(m[1608]&~m[1609]&m[1610]&~m[1611]&m[1675])|(~m[1608]&m[1609]&m[1610]&~m[1611]&m[1675])|(m[1608]&m[1609]&m[1610]&~m[1611]&m[1675])|(m[1608]&m[1609]&m[1610]&m[1611]&m[1675]))):InitCond[1977];
    m[1617] = run?((((m[1613]&~m[1614]&~m[1615]&~m[1616]&~m[1680])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1680])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1680])|(m[1613]&m[1614]&~m[1615]&m[1616]&~m[1680])|(m[1613]&~m[1614]&m[1615]&m[1616]&~m[1680])|(~m[1613]&m[1614]&m[1615]&m[1616]&~m[1680]))&BiasedRNG[1032])|(((m[1613]&~m[1614]&~m[1615]&~m[1616]&m[1680])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&m[1680])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&m[1680])|(m[1613]&m[1614]&~m[1615]&m[1616]&m[1680])|(m[1613]&~m[1614]&m[1615]&m[1616]&m[1680])|(~m[1613]&m[1614]&m[1615]&m[1616]&m[1680]))&~BiasedRNG[1032])|((m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1680])|(m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1680])|(~m[1613]&m[1614]&m[1615]&~m[1616]&~m[1680])|(m[1613]&m[1614]&m[1615]&~m[1616]&~m[1680])|(m[1613]&m[1614]&m[1615]&m[1616]&~m[1680])|(m[1613]&m[1614]&~m[1615]&~m[1616]&m[1680])|(m[1613]&~m[1614]&m[1615]&~m[1616]&m[1680])|(~m[1613]&m[1614]&m[1615]&~m[1616]&m[1680])|(m[1613]&m[1614]&m[1615]&~m[1616]&m[1680])|(m[1613]&m[1614]&m[1615]&m[1616]&m[1680]))):InitCond[1978];
    m[1622] = run?((((m[1618]&~m[1619]&~m[1620]&~m[1621]&~m[1685])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1685])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1685])|(m[1618]&m[1619]&~m[1620]&m[1621]&~m[1685])|(m[1618]&~m[1619]&m[1620]&m[1621]&~m[1685])|(~m[1618]&m[1619]&m[1620]&m[1621]&~m[1685]))&BiasedRNG[1033])|(((m[1618]&~m[1619]&~m[1620]&~m[1621]&m[1685])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&m[1685])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&m[1685])|(m[1618]&m[1619]&~m[1620]&m[1621]&m[1685])|(m[1618]&~m[1619]&m[1620]&m[1621]&m[1685])|(~m[1618]&m[1619]&m[1620]&m[1621]&m[1685]))&~BiasedRNG[1033])|((m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1685])|(m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1685])|(~m[1618]&m[1619]&m[1620]&~m[1621]&~m[1685])|(m[1618]&m[1619]&m[1620]&~m[1621]&~m[1685])|(m[1618]&m[1619]&m[1620]&m[1621]&~m[1685])|(m[1618]&m[1619]&~m[1620]&~m[1621]&m[1685])|(m[1618]&~m[1619]&m[1620]&~m[1621]&m[1685])|(~m[1618]&m[1619]&m[1620]&~m[1621]&m[1685])|(m[1618]&m[1619]&m[1620]&~m[1621]&m[1685])|(m[1618]&m[1619]&m[1620]&m[1621]&m[1685]))):InitCond[1979];
    m[1627] = run?((((m[1623]&~m[1624]&~m[1625]&~m[1626]&~m[1690])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1690])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1690])|(m[1623]&m[1624]&~m[1625]&m[1626]&~m[1690])|(m[1623]&~m[1624]&m[1625]&m[1626]&~m[1690])|(~m[1623]&m[1624]&m[1625]&m[1626]&~m[1690]))&BiasedRNG[1034])|(((m[1623]&~m[1624]&~m[1625]&~m[1626]&m[1690])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&m[1690])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&m[1690])|(m[1623]&m[1624]&~m[1625]&m[1626]&m[1690])|(m[1623]&~m[1624]&m[1625]&m[1626]&m[1690])|(~m[1623]&m[1624]&m[1625]&m[1626]&m[1690]))&~BiasedRNG[1034])|((m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1690])|(m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1690])|(~m[1623]&m[1624]&m[1625]&~m[1626]&~m[1690])|(m[1623]&m[1624]&m[1625]&~m[1626]&~m[1690])|(m[1623]&m[1624]&m[1625]&m[1626]&~m[1690])|(m[1623]&m[1624]&~m[1625]&~m[1626]&m[1690])|(m[1623]&~m[1624]&m[1625]&~m[1626]&m[1690])|(~m[1623]&m[1624]&m[1625]&~m[1626]&m[1690])|(m[1623]&m[1624]&m[1625]&~m[1626]&m[1690])|(m[1623]&m[1624]&m[1625]&m[1626]&m[1690]))):InitCond[1980];
    m[1632] = run?((((m[1628]&~m[1629]&~m[1630]&~m[1631]&~m[1695])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1695])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1695])|(m[1628]&m[1629]&~m[1630]&m[1631]&~m[1695])|(m[1628]&~m[1629]&m[1630]&m[1631]&~m[1695])|(~m[1628]&m[1629]&m[1630]&m[1631]&~m[1695]))&BiasedRNG[1035])|(((m[1628]&~m[1629]&~m[1630]&~m[1631]&m[1695])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&m[1695])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&m[1695])|(m[1628]&m[1629]&~m[1630]&m[1631]&m[1695])|(m[1628]&~m[1629]&m[1630]&m[1631]&m[1695])|(~m[1628]&m[1629]&m[1630]&m[1631]&m[1695]))&~BiasedRNG[1035])|((m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1695])|(m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1695])|(~m[1628]&m[1629]&m[1630]&~m[1631]&~m[1695])|(m[1628]&m[1629]&m[1630]&~m[1631]&~m[1695])|(m[1628]&m[1629]&m[1630]&m[1631]&~m[1695])|(m[1628]&m[1629]&~m[1630]&~m[1631]&m[1695])|(m[1628]&~m[1629]&m[1630]&~m[1631]&m[1695])|(~m[1628]&m[1629]&m[1630]&~m[1631]&m[1695])|(m[1628]&m[1629]&m[1630]&~m[1631]&m[1695])|(m[1628]&m[1629]&m[1630]&m[1631]&m[1695]))):InitCond[1981];
    m[1637] = run?((((m[1633]&~m[1634]&~m[1635]&~m[1636]&~m[1700])|(~m[1633]&m[1634]&~m[1635]&~m[1636]&~m[1700])|(~m[1633]&~m[1634]&m[1635]&~m[1636]&~m[1700])|(m[1633]&m[1634]&~m[1635]&m[1636]&~m[1700])|(m[1633]&~m[1634]&m[1635]&m[1636]&~m[1700])|(~m[1633]&m[1634]&m[1635]&m[1636]&~m[1700]))&BiasedRNG[1036])|(((m[1633]&~m[1634]&~m[1635]&~m[1636]&m[1700])|(~m[1633]&m[1634]&~m[1635]&~m[1636]&m[1700])|(~m[1633]&~m[1634]&m[1635]&~m[1636]&m[1700])|(m[1633]&m[1634]&~m[1635]&m[1636]&m[1700])|(m[1633]&~m[1634]&m[1635]&m[1636]&m[1700])|(~m[1633]&m[1634]&m[1635]&m[1636]&m[1700]))&~BiasedRNG[1036])|((m[1633]&m[1634]&~m[1635]&~m[1636]&~m[1700])|(m[1633]&~m[1634]&m[1635]&~m[1636]&~m[1700])|(~m[1633]&m[1634]&m[1635]&~m[1636]&~m[1700])|(m[1633]&m[1634]&m[1635]&~m[1636]&~m[1700])|(m[1633]&m[1634]&m[1635]&m[1636]&~m[1700])|(m[1633]&m[1634]&~m[1635]&~m[1636]&m[1700])|(m[1633]&~m[1634]&m[1635]&~m[1636]&m[1700])|(~m[1633]&m[1634]&m[1635]&~m[1636]&m[1700])|(m[1633]&m[1634]&m[1635]&~m[1636]&m[1700])|(m[1633]&m[1634]&m[1635]&m[1636]&m[1700]))):InitCond[1982];
    m[1642] = run?((((m[1638]&~m[1639]&~m[1640]&~m[1641]&~m[1705])|(~m[1638]&m[1639]&~m[1640]&~m[1641]&~m[1705])|(~m[1638]&~m[1639]&m[1640]&~m[1641]&~m[1705])|(m[1638]&m[1639]&~m[1640]&m[1641]&~m[1705])|(m[1638]&~m[1639]&m[1640]&m[1641]&~m[1705])|(~m[1638]&m[1639]&m[1640]&m[1641]&~m[1705]))&BiasedRNG[1037])|(((m[1638]&~m[1639]&~m[1640]&~m[1641]&m[1705])|(~m[1638]&m[1639]&~m[1640]&~m[1641]&m[1705])|(~m[1638]&~m[1639]&m[1640]&~m[1641]&m[1705])|(m[1638]&m[1639]&~m[1640]&m[1641]&m[1705])|(m[1638]&~m[1639]&m[1640]&m[1641]&m[1705])|(~m[1638]&m[1639]&m[1640]&m[1641]&m[1705]))&~BiasedRNG[1037])|((m[1638]&m[1639]&~m[1640]&~m[1641]&~m[1705])|(m[1638]&~m[1639]&m[1640]&~m[1641]&~m[1705])|(~m[1638]&m[1639]&m[1640]&~m[1641]&~m[1705])|(m[1638]&m[1639]&m[1640]&~m[1641]&~m[1705])|(m[1638]&m[1639]&m[1640]&m[1641]&~m[1705])|(m[1638]&m[1639]&~m[1640]&~m[1641]&m[1705])|(m[1638]&~m[1639]&m[1640]&~m[1641]&m[1705])|(~m[1638]&m[1639]&m[1640]&~m[1641]&m[1705])|(m[1638]&m[1639]&m[1640]&~m[1641]&m[1705])|(m[1638]&m[1639]&m[1640]&m[1641]&m[1705]))):InitCond[1983];
    m[1647] = run?((((m[1643]&~m[1644]&~m[1645]&~m[1646]&~m[1710])|(~m[1643]&m[1644]&~m[1645]&~m[1646]&~m[1710])|(~m[1643]&~m[1644]&m[1645]&~m[1646]&~m[1710])|(m[1643]&m[1644]&~m[1645]&m[1646]&~m[1710])|(m[1643]&~m[1644]&m[1645]&m[1646]&~m[1710])|(~m[1643]&m[1644]&m[1645]&m[1646]&~m[1710]))&BiasedRNG[1038])|(((m[1643]&~m[1644]&~m[1645]&~m[1646]&m[1710])|(~m[1643]&m[1644]&~m[1645]&~m[1646]&m[1710])|(~m[1643]&~m[1644]&m[1645]&~m[1646]&m[1710])|(m[1643]&m[1644]&~m[1645]&m[1646]&m[1710])|(m[1643]&~m[1644]&m[1645]&m[1646]&m[1710])|(~m[1643]&m[1644]&m[1645]&m[1646]&m[1710]))&~BiasedRNG[1038])|((m[1643]&m[1644]&~m[1645]&~m[1646]&~m[1710])|(m[1643]&~m[1644]&m[1645]&~m[1646]&~m[1710])|(~m[1643]&m[1644]&m[1645]&~m[1646]&~m[1710])|(m[1643]&m[1644]&m[1645]&~m[1646]&~m[1710])|(m[1643]&m[1644]&m[1645]&m[1646]&~m[1710])|(m[1643]&m[1644]&~m[1645]&~m[1646]&m[1710])|(m[1643]&~m[1644]&m[1645]&~m[1646]&m[1710])|(~m[1643]&m[1644]&m[1645]&~m[1646]&m[1710])|(m[1643]&m[1644]&m[1645]&~m[1646]&m[1710])|(m[1643]&m[1644]&m[1645]&m[1646]&m[1710]))):InitCond[1984];
    m[1652] = run?((((m[1648]&~m[1649]&~m[1650]&~m[1651]&~m[1715])|(~m[1648]&m[1649]&~m[1650]&~m[1651]&~m[1715])|(~m[1648]&~m[1649]&m[1650]&~m[1651]&~m[1715])|(m[1648]&m[1649]&~m[1650]&m[1651]&~m[1715])|(m[1648]&~m[1649]&m[1650]&m[1651]&~m[1715])|(~m[1648]&m[1649]&m[1650]&m[1651]&~m[1715]))&BiasedRNG[1039])|(((m[1648]&~m[1649]&~m[1650]&~m[1651]&m[1715])|(~m[1648]&m[1649]&~m[1650]&~m[1651]&m[1715])|(~m[1648]&~m[1649]&m[1650]&~m[1651]&m[1715])|(m[1648]&m[1649]&~m[1650]&m[1651]&m[1715])|(m[1648]&~m[1649]&m[1650]&m[1651]&m[1715])|(~m[1648]&m[1649]&m[1650]&m[1651]&m[1715]))&~BiasedRNG[1039])|((m[1648]&m[1649]&~m[1650]&~m[1651]&~m[1715])|(m[1648]&~m[1649]&m[1650]&~m[1651]&~m[1715])|(~m[1648]&m[1649]&m[1650]&~m[1651]&~m[1715])|(m[1648]&m[1649]&m[1650]&~m[1651]&~m[1715])|(m[1648]&m[1649]&m[1650]&m[1651]&~m[1715])|(m[1648]&m[1649]&~m[1650]&~m[1651]&m[1715])|(m[1648]&~m[1649]&m[1650]&~m[1651]&m[1715])|(~m[1648]&m[1649]&m[1650]&~m[1651]&m[1715])|(m[1648]&m[1649]&m[1650]&~m[1651]&m[1715])|(m[1648]&m[1649]&m[1650]&m[1651]&m[1715]))):InitCond[1985];
    m[1657] = run?((((m[1653]&~m[1654]&~m[1655]&~m[1656]&~m[1720])|(~m[1653]&m[1654]&~m[1655]&~m[1656]&~m[1720])|(~m[1653]&~m[1654]&m[1655]&~m[1656]&~m[1720])|(m[1653]&m[1654]&~m[1655]&m[1656]&~m[1720])|(m[1653]&~m[1654]&m[1655]&m[1656]&~m[1720])|(~m[1653]&m[1654]&m[1655]&m[1656]&~m[1720]))&BiasedRNG[1040])|(((m[1653]&~m[1654]&~m[1655]&~m[1656]&m[1720])|(~m[1653]&m[1654]&~m[1655]&~m[1656]&m[1720])|(~m[1653]&~m[1654]&m[1655]&~m[1656]&m[1720])|(m[1653]&m[1654]&~m[1655]&m[1656]&m[1720])|(m[1653]&~m[1654]&m[1655]&m[1656]&m[1720])|(~m[1653]&m[1654]&m[1655]&m[1656]&m[1720]))&~BiasedRNG[1040])|((m[1653]&m[1654]&~m[1655]&~m[1656]&~m[1720])|(m[1653]&~m[1654]&m[1655]&~m[1656]&~m[1720])|(~m[1653]&m[1654]&m[1655]&~m[1656]&~m[1720])|(m[1653]&m[1654]&m[1655]&~m[1656]&~m[1720])|(m[1653]&m[1654]&m[1655]&m[1656]&~m[1720])|(m[1653]&m[1654]&~m[1655]&~m[1656]&m[1720])|(m[1653]&~m[1654]&m[1655]&~m[1656]&m[1720])|(~m[1653]&m[1654]&m[1655]&~m[1656]&m[1720])|(m[1653]&m[1654]&m[1655]&~m[1656]&m[1720])|(m[1653]&m[1654]&m[1655]&m[1656]&m[1720]))):InitCond[1986];
    m[1662] = run?((((m[1658]&~m[1659]&~m[1660]&~m[1661]&~m[1725])|(~m[1658]&m[1659]&~m[1660]&~m[1661]&~m[1725])|(~m[1658]&~m[1659]&m[1660]&~m[1661]&~m[1725])|(m[1658]&m[1659]&~m[1660]&m[1661]&~m[1725])|(m[1658]&~m[1659]&m[1660]&m[1661]&~m[1725])|(~m[1658]&m[1659]&m[1660]&m[1661]&~m[1725]))&BiasedRNG[1041])|(((m[1658]&~m[1659]&~m[1660]&~m[1661]&m[1725])|(~m[1658]&m[1659]&~m[1660]&~m[1661]&m[1725])|(~m[1658]&~m[1659]&m[1660]&~m[1661]&m[1725])|(m[1658]&m[1659]&~m[1660]&m[1661]&m[1725])|(m[1658]&~m[1659]&m[1660]&m[1661]&m[1725])|(~m[1658]&m[1659]&m[1660]&m[1661]&m[1725]))&~BiasedRNG[1041])|((m[1658]&m[1659]&~m[1660]&~m[1661]&~m[1725])|(m[1658]&~m[1659]&m[1660]&~m[1661]&~m[1725])|(~m[1658]&m[1659]&m[1660]&~m[1661]&~m[1725])|(m[1658]&m[1659]&m[1660]&~m[1661]&~m[1725])|(m[1658]&m[1659]&m[1660]&m[1661]&~m[1725])|(m[1658]&m[1659]&~m[1660]&~m[1661]&m[1725])|(m[1658]&~m[1659]&m[1660]&~m[1661]&m[1725])|(~m[1658]&m[1659]&m[1660]&~m[1661]&m[1725])|(m[1658]&m[1659]&m[1660]&~m[1661]&m[1725])|(m[1658]&m[1659]&m[1660]&m[1661]&m[1725]))):InitCond[1987];
    m[1667] = run?((((m[1663]&~m[1664]&~m[1665]&~m[1666]&~m[1730])|(~m[1663]&m[1664]&~m[1665]&~m[1666]&~m[1730])|(~m[1663]&~m[1664]&m[1665]&~m[1666]&~m[1730])|(m[1663]&m[1664]&~m[1665]&m[1666]&~m[1730])|(m[1663]&~m[1664]&m[1665]&m[1666]&~m[1730])|(~m[1663]&m[1664]&m[1665]&m[1666]&~m[1730]))&BiasedRNG[1042])|(((m[1663]&~m[1664]&~m[1665]&~m[1666]&m[1730])|(~m[1663]&m[1664]&~m[1665]&~m[1666]&m[1730])|(~m[1663]&~m[1664]&m[1665]&~m[1666]&m[1730])|(m[1663]&m[1664]&~m[1665]&m[1666]&m[1730])|(m[1663]&~m[1664]&m[1665]&m[1666]&m[1730])|(~m[1663]&m[1664]&m[1665]&m[1666]&m[1730]))&~BiasedRNG[1042])|((m[1663]&m[1664]&~m[1665]&~m[1666]&~m[1730])|(m[1663]&~m[1664]&m[1665]&~m[1666]&~m[1730])|(~m[1663]&m[1664]&m[1665]&~m[1666]&~m[1730])|(m[1663]&m[1664]&m[1665]&~m[1666]&~m[1730])|(m[1663]&m[1664]&m[1665]&m[1666]&~m[1730])|(m[1663]&m[1664]&~m[1665]&~m[1666]&m[1730])|(m[1663]&~m[1664]&m[1665]&~m[1666]&m[1730])|(~m[1663]&m[1664]&m[1665]&~m[1666]&m[1730])|(m[1663]&m[1664]&m[1665]&~m[1666]&m[1730])|(m[1663]&m[1664]&m[1665]&m[1666]&m[1730]))):InitCond[1988];
    m[1672] = run?((((m[1668]&~m[1669]&~m[1670]&~m[1671]&~m[1735])|(~m[1668]&m[1669]&~m[1670]&~m[1671]&~m[1735])|(~m[1668]&~m[1669]&m[1670]&~m[1671]&~m[1735])|(m[1668]&m[1669]&~m[1670]&m[1671]&~m[1735])|(m[1668]&~m[1669]&m[1670]&m[1671]&~m[1735])|(~m[1668]&m[1669]&m[1670]&m[1671]&~m[1735]))&BiasedRNG[1043])|(((m[1668]&~m[1669]&~m[1670]&~m[1671]&m[1735])|(~m[1668]&m[1669]&~m[1670]&~m[1671]&m[1735])|(~m[1668]&~m[1669]&m[1670]&~m[1671]&m[1735])|(m[1668]&m[1669]&~m[1670]&m[1671]&m[1735])|(m[1668]&~m[1669]&m[1670]&m[1671]&m[1735])|(~m[1668]&m[1669]&m[1670]&m[1671]&m[1735]))&~BiasedRNG[1043])|((m[1668]&m[1669]&~m[1670]&~m[1671]&~m[1735])|(m[1668]&~m[1669]&m[1670]&~m[1671]&~m[1735])|(~m[1668]&m[1669]&m[1670]&~m[1671]&~m[1735])|(m[1668]&m[1669]&m[1670]&~m[1671]&~m[1735])|(m[1668]&m[1669]&m[1670]&m[1671]&~m[1735])|(m[1668]&m[1669]&~m[1670]&~m[1671]&m[1735])|(m[1668]&~m[1669]&m[1670]&~m[1671]&m[1735])|(~m[1668]&m[1669]&m[1670]&~m[1671]&m[1735])|(m[1668]&m[1669]&m[1670]&~m[1671]&m[1735])|(m[1668]&m[1669]&m[1670]&m[1671]&m[1735]))):InitCond[1989];
    m[1677] = run?((((m[1673]&~m[1674]&~m[1675]&~m[1676]&~m[1738])|(~m[1673]&m[1674]&~m[1675]&~m[1676]&~m[1738])|(~m[1673]&~m[1674]&m[1675]&~m[1676]&~m[1738])|(m[1673]&m[1674]&~m[1675]&m[1676]&~m[1738])|(m[1673]&~m[1674]&m[1675]&m[1676]&~m[1738])|(~m[1673]&m[1674]&m[1675]&m[1676]&~m[1738]))&BiasedRNG[1044])|(((m[1673]&~m[1674]&~m[1675]&~m[1676]&m[1738])|(~m[1673]&m[1674]&~m[1675]&~m[1676]&m[1738])|(~m[1673]&~m[1674]&m[1675]&~m[1676]&m[1738])|(m[1673]&m[1674]&~m[1675]&m[1676]&m[1738])|(m[1673]&~m[1674]&m[1675]&m[1676]&m[1738])|(~m[1673]&m[1674]&m[1675]&m[1676]&m[1738]))&~BiasedRNG[1044])|((m[1673]&m[1674]&~m[1675]&~m[1676]&~m[1738])|(m[1673]&~m[1674]&m[1675]&~m[1676]&~m[1738])|(~m[1673]&m[1674]&m[1675]&~m[1676]&~m[1738])|(m[1673]&m[1674]&m[1675]&~m[1676]&~m[1738])|(m[1673]&m[1674]&m[1675]&m[1676]&~m[1738])|(m[1673]&m[1674]&~m[1675]&~m[1676]&m[1738])|(m[1673]&~m[1674]&m[1675]&~m[1676]&m[1738])|(~m[1673]&m[1674]&m[1675]&~m[1676]&m[1738])|(m[1673]&m[1674]&m[1675]&~m[1676]&m[1738])|(m[1673]&m[1674]&m[1675]&m[1676]&m[1738]))):InitCond[1990];
    m[1682] = run?((((m[1678]&~m[1679]&~m[1680]&~m[1681]&~m[1740])|(~m[1678]&m[1679]&~m[1680]&~m[1681]&~m[1740])|(~m[1678]&~m[1679]&m[1680]&~m[1681]&~m[1740])|(m[1678]&m[1679]&~m[1680]&m[1681]&~m[1740])|(m[1678]&~m[1679]&m[1680]&m[1681]&~m[1740])|(~m[1678]&m[1679]&m[1680]&m[1681]&~m[1740]))&BiasedRNG[1045])|(((m[1678]&~m[1679]&~m[1680]&~m[1681]&m[1740])|(~m[1678]&m[1679]&~m[1680]&~m[1681]&m[1740])|(~m[1678]&~m[1679]&m[1680]&~m[1681]&m[1740])|(m[1678]&m[1679]&~m[1680]&m[1681]&m[1740])|(m[1678]&~m[1679]&m[1680]&m[1681]&m[1740])|(~m[1678]&m[1679]&m[1680]&m[1681]&m[1740]))&~BiasedRNG[1045])|((m[1678]&m[1679]&~m[1680]&~m[1681]&~m[1740])|(m[1678]&~m[1679]&m[1680]&~m[1681]&~m[1740])|(~m[1678]&m[1679]&m[1680]&~m[1681]&~m[1740])|(m[1678]&m[1679]&m[1680]&~m[1681]&~m[1740])|(m[1678]&m[1679]&m[1680]&m[1681]&~m[1740])|(m[1678]&m[1679]&~m[1680]&~m[1681]&m[1740])|(m[1678]&~m[1679]&m[1680]&~m[1681]&m[1740])|(~m[1678]&m[1679]&m[1680]&~m[1681]&m[1740])|(m[1678]&m[1679]&m[1680]&~m[1681]&m[1740])|(m[1678]&m[1679]&m[1680]&m[1681]&m[1740]))):InitCond[1991];
    m[1687] = run?((((m[1683]&~m[1684]&~m[1685]&~m[1686]&~m[1745])|(~m[1683]&m[1684]&~m[1685]&~m[1686]&~m[1745])|(~m[1683]&~m[1684]&m[1685]&~m[1686]&~m[1745])|(m[1683]&m[1684]&~m[1685]&m[1686]&~m[1745])|(m[1683]&~m[1684]&m[1685]&m[1686]&~m[1745])|(~m[1683]&m[1684]&m[1685]&m[1686]&~m[1745]))&BiasedRNG[1046])|(((m[1683]&~m[1684]&~m[1685]&~m[1686]&m[1745])|(~m[1683]&m[1684]&~m[1685]&~m[1686]&m[1745])|(~m[1683]&~m[1684]&m[1685]&~m[1686]&m[1745])|(m[1683]&m[1684]&~m[1685]&m[1686]&m[1745])|(m[1683]&~m[1684]&m[1685]&m[1686]&m[1745])|(~m[1683]&m[1684]&m[1685]&m[1686]&m[1745]))&~BiasedRNG[1046])|((m[1683]&m[1684]&~m[1685]&~m[1686]&~m[1745])|(m[1683]&~m[1684]&m[1685]&~m[1686]&~m[1745])|(~m[1683]&m[1684]&m[1685]&~m[1686]&~m[1745])|(m[1683]&m[1684]&m[1685]&~m[1686]&~m[1745])|(m[1683]&m[1684]&m[1685]&m[1686]&~m[1745])|(m[1683]&m[1684]&~m[1685]&~m[1686]&m[1745])|(m[1683]&~m[1684]&m[1685]&~m[1686]&m[1745])|(~m[1683]&m[1684]&m[1685]&~m[1686]&m[1745])|(m[1683]&m[1684]&m[1685]&~m[1686]&m[1745])|(m[1683]&m[1684]&m[1685]&m[1686]&m[1745]))):InitCond[1992];
    m[1692] = run?((((m[1688]&~m[1689]&~m[1690]&~m[1691]&~m[1750])|(~m[1688]&m[1689]&~m[1690]&~m[1691]&~m[1750])|(~m[1688]&~m[1689]&m[1690]&~m[1691]&~m[1750])|(m[1688]&m[1689]&~m[1690]&m[1691]&~m[1750])|(m[1688]&~m[1689]&m[1690]&m[1691]&~m[1750])|(~m[1688]&m[1689]&m[1690]&m[1691]&~m[1750]))&BiasedRNG[1047])|(((m[1688]&~m[1689]&~m[1690]&~m[1691]&m[1750])|(~m[1688]&m[1689]&~m[1690]&~m[1691]&m[1750])|(~m[1688]&~m[1689]&m[1690]&~m[1691]&m[1750])|(m[1688]&m[1689]&~m[1690]&m[1691]&m[1750])|(m[1688]&~m[1689]&m[1690]&m[1691]&m[1750])|(~m[1688]&m[1689]&m[1690]&m[1691]&m[1750]))&~BiasedRNG[1047])|((m[1688]&m[1689]&~m[1690]&~m[1691]&~m[1750])|(m[1688]&~m[1689]&m[1690]&~m[1691]&~m[1750])|(~m[1688]&m[1689]&m[1690]&~m[1691]&~m[1750])|(m[1688]&m[1689]&m[1690]&~m[1691]&~m[1750])|(m[1688]&m[1689]&m[1690]&m[1691]&~m[1750])|(m[1688]&m[1689]&~m[1690]&~m[1691]&m[1750])|(m[1688]&~m[1689]&m[1690]&~m[1691]&m[1750])|(~m[1688]&m[1689]&m[1690]&~m[1691]&m[1750])|(m[1688]&m[1689]&m[1690]&~m[1691]&m[1750])|(m[1688]&m[1689]&m[1690]&m[1691]&m[1750]))):InitCond[1993];
    m[1697] = run?((((m[1693]&~m[1694]&~m[1695]&~m[1696]&~m[1755])|(~m[1693]&m[1694]&~m[1695]&~m[1696]&~m[1755])|(~m[1693]&~m[1694]&m[1695]&~m[1696]&~m[1755])|(m[1693]&m[1694]&~m[1695]&m[1696]&~m[1755])|(m[1693]&~m[1694]&m[1695]&m[1696]&~m[1755])|(~m[1693]&m[1694]&m[1695]&m[1696]&~m[1755]))&BiasedRNG[1048])|(((m[1693]&~m[1694]&~m[1695]&~m[1696]&m[1755])|(~m[1693]&m[1694]&~m[1695]&~m[1696]&m[1755])|(~m[1693]&~m[1694]&m[1695]&~m[1696]&m[1755])|(m[1693]&m[1694]&~m[1695]&m[1696]&m[1755])|(m[1693]&~m[1694]&m[1695]&m[1696]&m[1755])|(~m[1693]&m[1694]&m[1695]&m[1696]&m[1755]))&~BiasedRNG[1048])|((m[1693]&m[1694]&~m[1695]&~m[1696]&~m[1755])|(m[1693]&~m[1694]&m[1695]&~m[1696]&~m[1755])|(~m[1693]&m[1694]&m[1695]&~m[1696]&~m[1755])|(m[1693]&m[1694]&m[1695]&~m[1696]&~m[1755])|(m[1693]&m[1694]&m[1695]&m[1696]&~m[1755])|(m[1693]&m[1694]&~m[1695]&~m[1696]&m[1755])|(m[1693]&~m[1694]&m[1695]&~m[1696]&m[1755])|(~m[1693]&m[1694]&m[1695]&~m[1696]&m[1755])|(m[1693]&m[1694]&m[1695]&~m[1696]&m[1755])|(m[1693]&m[1694]&m[1695]&m[1696]&m[1755]))):InitCond[1994];
    m[1702] = run?((((m[1698]&~m[1699]&~m[1700]&~m[1701]&~m[1760])|(~m[1698]&m[1699]&~m[1700]&~m[1701]&~m[1760])|(~m[1698]&~m[1699]&m[1700]&~m[1701]&~m[1760])|(m[1698]&m[1699]&~m[1700]&m[1701]&~m[1760])|(m[1698]&~m[1699]&m[1700]&m[1701]&~m[1760])|(~m[1698]&m[1699]&m[1700]&m[1701]&~m[1760]))&BiasedRNG[1049])|(((m[1698]&~m[1699]&~m[1700]&~m[1701]&m[1760])|(~m[1698]&m[1699]&~m[1700]&~m[1701]&m[1760])|(~m[1698]&~m[1699]&m[1700]&~m[1701]&m[1760])|(m[1698]&m[1699]&~m[1700]&m[1701]&m[1760])|(m[1698]&~m[1699]&m[1700]&m[1701]&m[1760])|(~m[1698]&m[1699]&m[1700]&m[1701]&m[1760]))&~BiasedRNG[1049])|((m[1698]&m[1699]&~m[1700]&~m[1701]&~m[1760])|(m[1698]&~m[1699]&m[1700]&~m[1701]&~m[1760])|(~m[1698]&m[1699]&m[1700]&~m[1701]&~m[1760])|(m[1698]&m[1699]&m[1700]&~m[1701]&~m[1760])|(m[1698]&m[1699]&m[1700]&m[1701]&~m[1760])|(m[1698]&m[1699]&~m[1700]&~m[1701]&m[1760])|(m[1698]&~m[1699]&m[1700]&~m[1701]&m[1760])|(~m[1698]&m[1699]&m[1700]&~m[1701]&m[1760])|(m[1698]&m[1699]&m[1700]&~m[1701]&m[1760])|(m[1698]&m[1699]&m[1700]&m[1701]&m[1760]))):InitCond[1995];
    m[1707] = run?((((m[1703]&~m[1704]&~m[1705]&~m[1706]&~m[1765])|(~m[1703]&m[1704]&~m[1705]&~m[1706]&~m[1765])|(~m[1703]&~m[1704]&m[1705]&~m[1706]&~m[1765])|(m[1703]&m[1704]&~m[1705]&m[1706]&~m[1765])|(m[1703]&~m[1704]&m[1705]&m[1706]&~m[1765])|(~m[1703]&m[1704]&m[1705]&m[1706]&~m[1765]))&BiasedRNG[1050])|(((m[1703]&~m[1704]&~m[1705]&~m[1706]&m[1765])|(~m[1703]&m[1704]&~m[1705]&~m[1706]&m[1765])|(~m[1703]&~m[1704]&m[1705]&~m[1706]&m[1765])|(m[1703]&m[1704]&~m[1705]&m[1706]&m[1765])|(m[1703]&~m[1704]&m[1705]&m[1706]&m[1765])|(~m[1703]&m[1704]&m[1705]&m[1706]&m[1765]))&~BiasedRNG[1050])|((m[1703]&m[1704]&~m[1705]&~m[1706]&~m[1765])|(m[1703]&~m[1704]&m[1705]&~m[1706]&~m[1765])|(~m[1703]&m[1704]&m[1705]&~m[1706]&~m[1765])|(m[1703]&m[1704]&m[1705]&~m[1706]&~m[1765])|(m[1703]&m[1704]&m[1705]&m[1706]&~m[1765])|(m[1703]&m[1704]&~m[1705]&~m[1706]&m[1765])|(m[1703]&~m[1704]&m[1705]&~m[1706]&m[1765])|(~m[1703]&m[1704]&m[1705]&~m[1706]&m[1765])|(m[1703]&m[1704]&m[1705]&~m[1706]&m[1765])|(m[1703]&m[1704]&m[1705]&m[1706]&m[1765]))):InitCond[1996];
    m[1712] = run?((((m[1708]&~m[1709]&~m[1710]&~m[1711]&~m[1770])|(~m[1708]&m[1709]&~m[1710]&~m[1711]&~m[1770])|(~m[1708]&~m[1709]&m[1710]&~m[1711]&~m[1770])|(m[1708]&m[1709]&~m[1710]&m[1711]&~m[1770])|(m[1708]&~m[1709]&m[1710]&m[1711]&~m[1770])|(~m[1708]&m[1709]&m[1710]&m[1711]&~m[1770]))&BiasedRNG[1051])|(((m[1708]&~m[1709]&~m[1710]&~m[1711]&m[1770])|(~m[1708]&m[1709]&~m[1710]&~m[1711]&m[1770])|(~m[1708]&~m[1709]&m[1710]&~m[1711]&m[1770])|(m[1708]&m[1709]&~m[1710]&m[1711]&m[1770])|(m[1708]&~m[1709]&m[1710]&m[1711]&m[1770])|(~m[1708]&m[1709]&m[1710]&m[1711]&m[1770]))&~BiasedRNG[1051])|((m[1708]&m[1709]&~m[1710]&~m[1711]&~m[1770])|(m[1708]&~m[1709]&m[1710]&~m[1711]&~m[1770])|(~m[1708]&m[1709]&m[1710]&~m[1711]&~m[1770])|(m[1708]&m[1709]&m[1710]&~m[1711]&~m[1770])|(m[1708]&m[1709]&m[1710]&m[1711]&~m[1770])|(m[1708]&m[1709]&~m[1710]&~m[1711]&m[1770])|(m[1708]&~m[1709]&m[1710]&~m[1711]&m[1770])|(~m[1708]&m[1709]&m[1710]&~m[1711]&m[1770])|(m[1708]&m[1709]&m[1710]&~m[1711]&m[1770])|(m[1708]&m[1709]&m[1710]&m[1711]&m[1770]))):InitCond[1997];
    m[1717] = run?((((m[1713]&~m[1714]&~m[1715]&~m[1716]&~m[1775])|(~m[1713]&m[1714]&~m[1715]&~m[1716]&~m[1775])|(~m[1713]&~m[1714]&m[1715]&~m[1716]&~m[1775])|(m[1713]&m[1714]&~m[1715]&m[1716]&~m[1775])|(m[1713]&~m[1714]&m[1715]&m[1716]&~m[1775])|(~m[1713]&m[1714]&m[1715]&m[1716]&~m[1775]))&BiasedRNG[1052])|(((m[1713]&~m[1714]&~m[1715]&~m[1716]&m[1775])|(~m[1713]&m[1714]&~m[1715]&~m[1716]&m[1775])|(~m[1713]&~m[1714]&m[1715]&~m[1716]&m[1775])|(m[1713]&m[1714]&~m[1715]&m[1716]&m[1775])|(m[1713]&~m[1714]&m[1715]&m[1716]&m[1775])|(~m[1713]&m[1714]&m[1715]&m[1716]&m[1775]))&~BiasedRNG[1052])|((m[1713]&m[1714]&~m[1715]&~m[1716]&~m[1775])|(m[1713]&~m[1714]&m[1715]&~m[1716]&~m[1775])|(~m[1713]&m[1714]&m[1715]&~m[1716]&~m[1775])|(m[1713]&m[1714]&m[1715]&~m[1716]&~m[1775])|(m[1713]&m[1714]&m[1715]&m[1716]&~m[1775])|(m[1713]&m[1714]&~m[1715]&~m[1716]&m[1775])|(m[1713]&~m[1714]&m[1715]&~m[1716]&m[1775])|(~m[1713]&m[1714]&m[1715]&~m[1716]&m[1775])|(m[1713]&m[1714]&m[1715]&~m[1716]&m[1775])|(m[1713]&m[1714]&m[1715]&m[1716]&m[1775]))):InitCond[1998];
    m[1722] = run?((((m[1718]&~m[1719]&~m[1720]&~m[1721]&~m[1780])|(~m[1718]&m[1719]&~m[1720]&~m[1721]&~m[1780])|(~m[1718]&~m[1719]&m[1720]&~m[1721]&~m[1780])|(m[1718]&m[1719]&~m[1720]&m[1721]&~m[1780])|(m[1718]&~m[1719]&m[1720]&m[1721]&~m[1780])|(~m[1718]&m[1719]&m[1720]&m[1721]&~m[1780]))&BiasedRNG[1053])|(((m[1718]&~m[1719]&~m[1720]&~m[1721]&m[1780])|(~m[1718]&m[1719]&~m[1720]&~m[1721]&m[1780])|(~m[1718]&~m[1719]&m[1720]&~m[1721]&m[1780])|(m[1718]&m[1719]&~m[1720]&m[1721]&m[1780])|(m[1718]&~m[1719]&m[1720]&m[1721]&m[1780])|(~m[1718]&m[1719]&m[1720]&m[1721]&m[1780]))&~BiasedRNG[1053])|((m[1718]&m[1719]&~m[1720]&~m[1721]&~m[1780])|(m[1718]&~m[1719]&m[1720]&~m[1721]&~m[1780])|(~m[1718]&m[1719]&m[1720]&~m[1721]&~m[1780])|(m[1718]&m[1719]&m[1720]&~m[1721]&~m[1780])|(m[1718]&m[1719]&m[1720]&m[1721]&~m[1780])|(m[1718]&m[1719]&~m[1720]&~m[1721]&m[1780])|(m[1718]&~m[1719]&m[1720]&~m[1721]&m[1780])|(~m[1718]&m[1719]&m[1720]&~m[1721]&m[1780])|(m[1718]&m[1719]&m[1720]&~m[1721]&m[1780])|(m[1718]&m[1719]&m[1720]&m[1721]&m[1780]))):InitCond[1999];
    m[1727] = run?((((m[1723]&~m[1724]&~m[1725]&~m[1726]&~m[1785])|(~m[1723]&m[1724]&~m[1725]&~m[1726]&~m[1785])|(~m[1723]&~m[1724]&m[1725]&~m[1726]&~m[1785])|(m[1723]&m[1724]&~m[1725]&m[1726]&~m[1785])|(m[1723]&~m[1724]&m[1725]&m[1726]&~m[1785])|(~m[1723]&m[1724]&m[1725]&m[1726]&~m[1785]))&BiasedRNG[1054])|(((m[1723]&~m[1724]&~m[1725]&~m[1726]&m[1785])|(~m[1723]&m[1724]&~m[1725]&~m[1726]&m[1785])|(~m[1723]&~m[1724]&m[1725]&~m[1726]&m[1785])|(m[1723]&m[1724]&~m[1725]&m[1726]&m[1785])|(m[1723]&~m[1724]&m[1725]&m[1726]&m[1785])|(~m[1723]&m[1724]&m[1725]&m[1726]&m[1785]))&~BiasedRNG[1054])|((m[1723]&m[1724]&~m[1725]&~m[1726]&~m[1785])|(m[1723]&~m[1724]&m[1725]&~m[1726]&~m[1785])|(~m[1723]&m[1724]&m[1725]&~m[1726]&~m[1785])|(m[1723]&m[1724]&m[1725]&~m[1726]&~m[1785])|(m[1723]&m[1724]&m[1725]&m[1726]&~m[1785])|(m[1723]&m[1724]&~m[1725]&~m[1726]&m[1785])|(m[1723]&~m[1724]&m[1725]&~m[1726]&m[1785])|(~m[1723]&m[1724]&m[1725]&~m[1726]&m[1785])|(m[1723]&m[1724]&m[1725]&~m[1726]&m[1785])|(m[1723]&m[1724]&m[1725]&m[1726]&m[1785]))):InitCond[2000];
    m[1732] = run?((((m[1728]&~m[1729]&~m[1730]&~m[1731]&~m[1790])|(~m[1728]&m[1729]&~m[1730]&~m[1731]&~m[1790])|(~m[1728]&~m[1729]&m[1730]&~m[1731]&~m[1790])|(m[1728]&m[1729]&~m[1730]&m[1731]&~m[1790])|(m[1728]&~m[1729]&m[1730]&m[1731]&~m[1790])|(~m[1728]&m[1729]&m[1730]&m[1731]&~m[1790]))&BiasedRNG[1055])|(((m[1728]&~m[1729]&~m[1730]&~m[1731]&m[1790])|(~m[1728]&m[1729]&~m[1730]&~m[1731]&m[1790])|(~m[1728]&~m[1729]&m[1730]&~m[1731]&m[1790])|(m[1728]&m[1729]&~m[1730]&m[1731]&m[1790])|(m[1728]&~m[1729]&m[1730]&m[1731]&m[1790])|(~m[1728]&m[1729]&m[1730]&m[1731]&m[1790]))&~BiasedRNG[1055])|((m[1728]&m[1729]&~m[1730]&~m[1731]&~m[1790])|(m[1728]&~m[1729]&m[1730]&~m[1731]&~m[1790])|(~m[1728]&m[1729]&m[1730]&~m[1731]&~m[1790])|(m[1728]&m[1729]&m[1730]&~m[1731]&~m[1790])|(m[1728]&m[1729]&m[1730]&m[1731]&~m[1790])|(m[1728]&m[1729]&~m[1730]&~m[1731]&m[1790])|(m[1728]&~m[1729]&m[1730]&~m[1731]&m[1790])|(~m[1728]&m[1729]&m[1730]&~m[1731]&m[1790])|(m[1728]&m[1729]&m[1730]&~m[1731]&m[1790])|(m[1728]&m[1729]&m[1730]&m[1731]&m[1790]))):InitCond[2001];
    m[1737] = run?((((m[1733]&~m[1734]&~m[1735]&~m[1736]&~m[1795])|(~m[1733]&m[1734]&~m[1735]&~m[1736]&~m[1795])|(~m[1733]&~m[1734]&m[1735]&~m[1736]&~m[1795])|(m[1733]&m[1734]&~m[1735]&m[1736]&~m[1795])|(m[1733]&~m[1734]&m[1735]&m[1736]&~m[1795])|(~m[1733]&m[1734]&m[1735]&m[1736]&~m[1795]))&BiasedRNG[1056])|(((m[1733]&~m[1734]&~m[1735]&~m[1736]&m[1795])|(~m[1733]&m[1734]&~m[1735]&~m[1736]&m[1795])|(~m[1733]&~m[1734]&m[1735]&~m[1736]&m[1795])|(m[1733]&m[1734]&~m[1735]&m[1736]&m[1795])|(m[1733]&~m[1734]&m[1735]&m[1736]&m[1795])|(~m[1733]&m[1734]&m[1735]&m[1736]&m[1795]))&~BiasedRNG[1056])|((m[1733]&m[1734]&~m[1735]&~m[1736]&~m[1795])|(m[1733]&~m[1734]&m[1735]&~m[1736]&~m[1795])|(~m[1733]&m[1734]&m[1735]&~m[1736]&~m[1795])|(m[1733]&m[1734]&m[1735]&~m[1736]&~m[1795])|(m[1733]&m[1734]&m[1735]&m[1736]&~m[1795])|(m[1733]&m[1734]&~m[1735]&~m[1736]&m[1795])|(m[1733]&~m[1734]&m[1735]&~m[1736]&m[1795])|(~m[1733]&m[1734]&m[1735]&~m[1736]&m[1795])|(m[1733]&m[1734]&m[1735]&~m[1736]&m[1795])|(m[1733]&m[1734]&m[1735]&m[1736]&m[1795]))):InitCond[2002];
    m[1742] = run?((((m[1738]&~m[1739]&~m[1740]&~m[1741]&~m[1798])|(~m[1738]&m[1739]&~m[1740]&~m[1741]&~m[1798])|(~m[1738]&~m[1739]&m[1740]&~m[1741]&~m[1798])|(m[1738]&m[1739]&~m[1740]&m[1741]&~m[1798])|(m[1738]&~m[1739]&m[1740]&m[1741]&~m[1798])|(~m[1738]&m[1739]&m[1740]&m[1741]&~m[1798]))&BiasedRNG[1057])|(((m[1738]&~m[1739]&~m[1740]&~m[1741]&m[1798])|(~m[1738]&m[1739]&~m[1740]&~m[1741]&m[1798])|(~m[1738]&~m[1739]&m[1740]&~m[1741]&m[1798])|(m[1738]&m[1739]&~m[1740]&m[1741]&m[1798])|(m[1738]&~m[1739]&m[1740]&m[1741]&m[1798])|(~m[1738]&m[1739]&m[1740]&m[1741]&m[1798]))&~BiasedRNG[1057])|((m[1738]&m[1739]&~m[1740]&~m[1741]&~m[1798])|(m[1738]&~m[1739]&m[1740]&~m[1741]&~m[1798])|(~m[1738]&m[1739]&m[1740]&~m[1741]&~m[1798])|(m[1738]&m[1739]&m[1740]&~m[1741]&~m[1798])|(m[1738]&m[1739]&m[1740]&m[1741]&~m[1798])|(m[1738]&m[1739]&~m[1740]&~m[1741]&m[1798])|(m[1738]&~m[1739]&m[1740]&~m[1741]&m[1798])|(~m[1738]&m[1739]&m[1740]&~m[1741]&m[1798])|(m[1738]&m[1739]&m[1740]&~m[1741]&m[1798])|(m[1738]&m[1739]&m[1740]&m[1741]&m[1798]))):InitCond[2003];
    m[1747] = run?((((m[1743]&~m[1744]&~m[1745]&~m[1746]&~m[1800])|(~m[1743]&m[1744]&~m[1745]&~m[1746]&~m[1800])|(~m[1743]&~m[1744]&m[1745]&~m[1746]&~m[1800])|(m[1743]&m[1744]&~m[1745]&m[1746]&~m[1800])|(m[1743]&~m[1744]&m[1745]&m[1746]&~m[1800])|(~m[1743]&m[1744]&m[1745]&m[1746]&~m[1800]))&BiasedRNG[1058])|(((m[1743]&~m[1744]&~m[1745]&~m[1746]&m[1800])|(~m[1743]&m[1744]&~m[1745]&~m[1746]&m[1800])|(~m[1743]&~m[1744]&m[1745]&~m[1746]&m[1800])|(m[1743]&m[1744]&~m[1745]&m[1746]&m[1800])|(m[1743]&~m[1744]&m[1745]&m[1746]&m[1800])|(~m[1743]&m[1744]&m[1745]&m[1746]&m[1800]))&~BiasedRNG[1058])|((m[1743]&m[1744]&~m[1745]&~m[1746]&~m[1800])|(m[1743]&~m[1744]&m[1745]&~m[1746]&~m[1800])|(~m[1743]&m[1744]&m[1745]&~m[1746]&~m[1800])|(m[1743]&m[1744]&m[1745]&~m[1746]&~m[1800])|(m[1743]&m[1744]&m[1745]&m[1746]&~m[1800])|(m[1743]&m[1744]&~m[1745]&~m[1746]&m[1800])|(m[1743]&~m[1744]&m[1745]&~m[1746]&m[1800])|(~m[1743]&m[1744]&m[1745]&~m[1746]&m[1800])|(m[1743]&m[1744]&m[1745]&~m[1746]&m[1800])|(m[1743]&m[1744]&m[1745]&m[1746]&m[1800]))):InitCond[2004];
    m[1752] = run?((((m[1748]&~m[1749]&~m[1750]&~m[1751]&~m[1805])|(~m[1748]&m[1749]&~m[1750]&~m[1751]&~m[1805])|(~m[1748]&~m[1749]&m[1750]&~m[1751]&~m[1805])|(m[1748]&m[1749]&~m[1750]&m[1751]&~m[1805])|(m[1748]&~m[1749]&m[1750]&m[1751]&~m[1805])|(~m[1748]&m[1749]&m[1750]&m[1751]&~m[1805]))&BiasedRNG[1059])|(((m[1748]&~m[1749]&~m[1750]&~m[1751]&m[1805])|(~m[1748]&m[1749]&~m[1750]&~m[1751]&m[1805])|(~m[1748]&~m[1749]&m[1750]&~m[1751]&m[1805])|(m[1748]&m[1749]&~m[1750]&m[1751]&m[1805])|(m[1748]&~m[1749]&m[1750]&m[1751]&m[1805])|(~m[1748]&m[1749]&m[1750]&m[1751]&m[1805]))&~BiasedRNG[1059])|((m[1748]&m[1749]&~m[1750]&~m[1751]&~m[1805])|(m[1748]&~m[1749]&m[1750]&~m[1751]&~m[1805])|(~m[1748]&m[1749]&m[1750]&~m[1751]&~m[1805])|(m[1748]&m[1749]&m[1750]&~m[1751]&~m[1805])|(m[1748]&m[1749]&m[1750]&m[1751]&~m[1805])|(m[1748]&m[1749]&~m[1750]&~m[1751]&m[1805])|(m[1748]&~m[1749]&m[1750]&~m[1751]&m[1805])|(~m[1748]&m[1749]&m[1750]&~m[1751]&m[1805])|(m[1748]&m[1749]&m[1750]&~m[1751]&m[1805])|(m[1748]&m[1749]&m[1750]&m[1751]&m[1805]))):InitCond[2005];
    m[1757] = run?((((m[1753]&~m[1754]&~m[1755]&~m[1756]&~m[1810])|(~m[1753]&m[1754]&~m[1755]&~m[1756]&~m[1810])|(~m[1753]&~m[1754]&m[1755]&~m[1756]&~m[1810])|(m[1753]&m[1754]&~m[1755]&m[1756]&~m[1810])|(m[1753]&~m[1754]&m[1755]&m[1756]&~m[1810])|(~m[1753]&m[1754]&m[1755]&m[1756]&~m[1810]))&BiasedRNG[1060])|(((m[1753]&~m[1754]&~m[1755]&~m[1756]&m[1810])|(~m[1753]&m[1754]&~m[1755]&~m[1756]&m[1810])|(~m[1753]&~m[1754]&m[1755]&~m[1756]&m[1810])|(m[1753]&m[1754]&~m[1755]&m[1756]&m[1810])|(m[1753]&~m[1754]&m[1755]&m[1756]&m[1810])|(~m[1753]&m[1754]&m[1755]&m[1756]&m[1810]))&~BiasedRNG[1060])|((m[1753]&m[1754]&~m[1755]&~m[1756]&~m[1810])|(m[1753]&~m[1754]&m[1755]&~m[1756]&~m[1810])|(~m[1753]&m[1754]&m[1755]&~m[1756]&~m[1810])|(m[1753]&m[1754]&m[1755]&~m[1756]&~m[1810])|(m[1753]&m[1754]&m[1755]&m[1756]&~m[1810])|(m[1753]&m[1754]&~m[1755]&~m[1756]&m[1810])|(m[1753]&~m[1754]&m[1755]&~m[1756]&m[1810])|(~m[1753]&m[1754]&m[1755]&~m[1756]&m[1810])|(m[1753]&m[1754]&m[1755]&~m[1756]&m[1810])|(m[1753]&m[1754]&m[1755]&m[1756]&m[1810]))):InitCond[2006];
    m[1762] = run?((((m[1758]&~m[1759]&~m[1760]&~m[1761]&~m[1815])|(~m[1758]&m[1759]&~m[1760]&~m[1761]&~m[1815])|(~m[1758]&~m[1759]&m[1760]&~m[1761]&~m[1815])|(m[1758]&m[1759]&~m[1760]&m[1761]&~m[1815])|(m[1758]&~m[1759]&m[1760]&m[1761]&~m[1815])|(~m[1758]&m[1759]&m[1760]&m[1761]&~m[1815]))&BiasedRNG[1061])|(((m[1758]&~m[1759]&~m[1760]&~m[1761]&m[1815])|(~m[1758]&m[1759]&~m[1760]&~m[1761]&m[1815])|(~m[1758]&~m[1759]&m[1760]&~m[1761]&m[1815])|(m[1758]&m[1759]&~m[1760]&m[1761]&m[1815])|(m[1758]&~m[1759]&m[1760]&m[1761]&m[1815])|(~m[1758]&m[1759]&m[1760]&m[1761]&m[1815]))&~BiasedRNG[1061])|((m[1758]&m[1759]&~m[1760]&~m[1761]&~m[1815])|(m[1758]&~m[1759]&m[1760]&~m[1761]&~m[1815])|(~m[1758]&m[1759]&m[1760]&~m[1761]&~m[1815])|(m[1758]&m[1759]&m[1760]&~m[1761]&~m[1815])|(m[1758]&m[1759]&m[1760]&m[1761]&~m[1815])|(m[1758]&m[1759]&~m[1760]&~m[1761]&m[1815])|(m[1758]&~m[1759]&m[1760]&~m[1761]&m[1815])|(~m[1758]&m[1759]&m[1760]&~m[1761]&m[1815])|(m[1758]&m[1759]&m[1760]&~m[1761]&m[1815])|(m[1758]&m[1759]&m[1760]&m[1761]&m[1815]))):InitCond[2007];
    m[1767] = run?((((m[1763]&~m[1764]&~m[1765]&~m[1766]&~m[1820])|(~m[1763]&m[1764]&~m[1765]&~m[1766]&~m[1820])|(~m[1763]&~m[1764]&m[1765]&~m[1766]&~m[1820])|(m[1763]&m[1764]&~m[1765]&m[1766]&~m[1820])|(m[1763]&~m[1764]&m[1765]&m[1766]&~m[1820])|(~m[1763]&m[1764]&m[1765]&m[1766]&~m[1820]))&BiasedRNG[1062])|(((m[1763]&~m[1764]&~m[1765]&~m[1766]&m[1820])|(~m[1763]&m[1764]&~m[1765]&~m[1766]&m[1820])|(~m[1763]&~m[1764]&m[1765]&~m[1766]&m[1820])|(m[1763]&m[1764]&~m[1765]&m[1766]&m[1820])|(m[1763]&~m[1764]&m[1765]&m[1766]&m[1820])|(~m[1763]&m[1764]&m[1765]&m[1766]&m[1820]))&~BiasedRNG[1062])|((m[1763]&m[1764]&~m[1765]&~m[1766]&~m[1820])|(m[1763]&~m[1764]&m[1765]&~m[1766]&~m[1820])|(~m[1763]&m[1764]&m[1765]&~m[1766]&~m[1820])|(m[1763]&m[1764]&m[1765]&~m[1766]&~m[1820])|(m[1763]&m[1764]&m[1765]&m[1766]&~m[1820])|(m[1763]&m[1764]&~m[1765]&~m[1766]&m[1820])|(m[1763]&~m[1764]&m[1765]&~m[1766]&m[1820])|(~m[1763]&m[1764]&m[1765]&~m[1766]&m[1820])|(m[1763]&m[1764]&m[1765]&~m[1766]&m[1820])|(m[1763]&m[1764]&m[1765]&m[1766]&m[1820]))):InitCond[2008];
    m[1772] = run?((((m[1768]&~m[1769]&~m[1770]&~m[1771]&~m[1825])|(~m[1768]&m[1769]&~m[1770]&~m[1771]&~m[1825])|(~m[1768]&~m[1769]&m[1770]&~m[1771]&~m[1825])|(m[1768]&m[1769]&~m[1770]&m[1771]&~m[1825])|(m[1768]&~m[1769]&m[1770]&m[1771]&~m[1825])|(~m[1768]&m[1769]&m[1770]&m[1771]&~m[1825]))&BiasedRNG[1063])|(((m[1768]&~m[1769]&~m[1770]&~m[1771]&m[1825])|(~m[1768]&m[1769]&~m[1770]&~m[1771]&m[1825])|(~m[1768]&~m[1769]&m[1770]&~m[1771]&m[1825])|(m[1768]&m[1769]&~m[1770]&m[1771]&m[1825])|(m[1768]&~m[1769]&m[1770]&m[1771]&m[1825])|(~m[1768]&m[1769]&m[1770]&m[1771]&m[1825]))&~BiasedRNG[1063])|((m[1768]&m[1769]&~m[1770]&~m[1771]&~m[1825])|(m[1768]&~m[1769]&m[1770]&~m[1771]&~m[1825])|(~m[1768]&m[1769]&m[1770]&~m[1771]&~m[1825])|(m[1768]&m[1769]&m[1770]&~m[1771]&~m[1825])|(m[1768]&m[1769]&m[1770]&m[1771]&~m[1825])|(m[1768]&m[1769]&~m[1770]&~m[1771]&m[1825])|(m[1768]&~m[1769]&m[1770]&~m[1771]&m[1825])|(~m[1768]&m[1769]&m[1770]&~m[1771]&m[1825])|(m[1768]&m[1769]&m[1770]&~m[1771]&m[1825])|(m[1768]&m[1769]&m[1770]&m[1771]&m[1825]))):InitCond[2009];
    m[1777] = run?((((m[1773]&~m[1774]&~m[1775]&~m[1776]&~m[1830])|(~m[1773]&m[1774]&~m[1775]&~m[1776]&~m[1830])|(~m[1773]&~m[1774]&m[1775]&~m[1776]&~m[1830])|(m[1773]&m[1774]&~m[1775]&m[1776]&~m[1830])|(m[1773]&~m[1774]&m[1775]&m[1776]&~m[1830])|(~m[1773]&m[1774]&m[1775]&m[1776]&~m[1830]))&BiasedRNG[1064])|(((m[1773]&~m[1774]&~m[1775]&~m[1776]&m[1830])|(~m[1773]&m[1774]&~m[1775]&~m[1776]&m[1830])|(~m[1773]&~m[1774]&m[1775]&~m[1776]&m[1830])|(m[1773]&m[1774]&~m[1775]&m[1776]&m[1830])|(m[1773]&~m[1774]&m[1775]&m[1776]&m[1830])|(~m[1773]&m[1774]&m[1775]&m[1776]&m[1830]))&~BiasedRNG[1064])|((m[1773]&m[1774]&~m[1775]&~m[1776]&~m[1830])|(m[1773]&~m[1774]&m[1775]&~m[1776]&~m[1830])|(~m[1773]&m[1774]&m[1775]&~m[1776]&~m[1830])|(m[1773]&m[1774]&m[1775]&~m[1776]&~m[1830])|(m[1773]&m[1774]&m[1775]&m[1776]&~m[1830])|(m[1773]&m[1774]&~m[1775]&~m[1776]&m[1830])|(m[1773]&~m[1774]&m[1775]&~m[1776]&m[1830])|(~m[1773]&m[1774]&m[1775]&~m[1776]&m[1830])|(m[1773]&m[1774]&m[1775]&~m[1776]&m[1830])|(m[1773]&m[1774]&m[1775]&m[1776]&m[1830]))):InitCond[2010];
    m[1782] = run?((((m[1778]&~m[1779]&~m[1780]&~m[1781]&~m[1835])|(~m[1778]&m[1779]&~m[1780]&~m[1781]&~m[1835])|(~m[1778]&~m[1779]&m[1780]&~m[1781]&~m[1835])|(m[1778]&m[1779]&~m[1780]&m[1781]&~m[1835])|(m[1778]&~m[1779]&m[1780]&m[1781]&~m[1835])|(~m[1778]&m[1779]&m[1780]&m[1781]&~m[1835]))&BiasedRNG[1065])|(((m[1778]&~m[1779]&~m[1780]&~m[1781]&m[1835])|(~m[1778]&m[1779]&~m[1780]&~m[1781]&m[1835])|(~m[1778]&~m[1779]&m[1780]&~m[1781]&m[1835])|(m[1778]&m[1779]&~m[1780]&m[1781]&m[1835])|(m[1778]&~m[1779]&m[1780]&m[1781]&m[1835])|(~m[1778]&m[1779]&m[1780]&m[1781]&m[1835]))&~BiasedRNG[1065])|((m[1778]&m[1779]&~m[1780]&~m[1781]&~m[1835])|(m[1778]&~m[1779]&m[1780]&~m[1781]&~m[1835])|(~m[1778]&m[1779]&m[1780]&~m[1781]&~m[1835])|(m[1778]&m[1779]&m[1780]&~m[1781]&~m[1835])|(m[1778]&m[1779]&m[1780]&m[1781]&~m[1835])|(m[1778]&m[1779]&~m[1780]&~m[1781]&m[1835])|(m[1778]&~m[1779]&m[1780]&~m[1781]&m[1835])|(~m[1778]&m[1779]&m[1780]&~m[1781]&m[1835])|(m[1778]&m[1779]&m[1780]&~m[1781]&m[1835])|(m[1778]&m[1779]&m[1780]&m[1781]&m[1835]))):InitCond[2011];
    m[1787] = run?((((m[1783]&~m[1784]&~m[1785]&~m[1786]&~m[1840])|(~m[1783]&m[1784]&~m[1785]&~m[1786]&~m[1840])|(~m[1783]&~m[1784]&m[1785]&~m[1786]&~m[1840])|(m[1783]&m[1784]&~m[1785]&m[1786]&~m[1840])|(m[1783]&~m[1784]&m[1785]&m[1786]&~m[1840])|(~m[1783]&m[1784]&m[1785]&m[1786]&~m[1840]))&BiasedRNG[1066])|(((m[1783]&~m[1784]&~m[1785]&~m[1786]&m[1840])|(~m[1783]&m[1784]&~m[1785]&~m[1786]&m[1840])|(~m[1783]&~m[1784]&m[1785]&~m[1786]&m[1840])|(m[1783]&m[1784]&~m[1785]&m[1786]&m[1840])|(m[1783]&~m[1784]&m[1785]&m[1786]&m[1840])|(~m[1783]&m[1784]&m[1785]&m[1786]&m[1840]))&~BiasedRNG[1066])|((m[1783]&m[1784]&~m[1785]&~m[1786]&~m[1840])|(m[1783]&~m[1784]&m[1785]&~m[1786]&~m[1840])|(~m[1783]&m[1784]&m[1785]&~m[1786]&~m[1840])|(m[1783]&m[1784]&m[1785]&~m[1786]&~m[1840])|(m[1783]&m[1784]&m[1785]&m[1786]&~m[1840])|(m[1783]&m[1784]&~m[1785]&~m[1786]&m[1840])|(m[1783]&~m[1784]&m[1785]&~m[1786]&m[1840])|(~m[1783]&m[1784]&m[1785]&~m[1786]&m[1840])|(m[1783]&m[1784]&m[1785]&~m[1786]&m[1840])|(m[1783]&m[1784]&m[1785]&m[1786]&m[1840]))):InitCond[2012];
    m[1792] = run?((((m[1788]&~m[1789]&~m[1790]&~m[1791]&~m[1845])|(~m[1788]&m[1789]&~m[1790]&~m[1791]&~m[1845])|(~m[1788]&~m[1789]&m[1790]&~m[1791]&~m[1845])|(m[1788]&m[1789]&~m[1790]&m[1791]&~m[1845])|(m[1788]&~m[1789]&m[1790]&m[1791]&~m[1845])|(~m[1788]&m[1789]&m[1790]&m[1791]&~m[1845]))&BiasedRNG[1067])|(((m[1788]&~m[1789]&~m[1790]&~m[1791]&m[1845])|(~m[1788]&m[1789]&~m[1790]&~m[1791]&m[1845])|(~m[1788]&~m[1789]&m[1790]&~m[1791]&m[1845])|(m[1788]&m[1789]&~m[1790]&m[1791]&m[1845])|(m[1788]&~m[1789]&m[1790]&m[1791]&m[1845])|(~m[1788]&m[1789]&m[1790]&m[1791]&m[1845]))&~BiasedRNG[1067])|((m[1788]&m[1789]&~m[1790]&~m[1791]&~m[1845])|(m[1788]&~m[1789]&m[1790]&~m[1791]&~m[1845])|(~m[1788]&m[1789]&m[1790]&~m[1791]&~m[1845])|(m[1788]&m[1789]&m[1790]&~m[1791]&~m[1845])|(m[1788]&m[1789]&m[1790]&m[1791]&~m[1845])|(m[1788]&m[1789]&~m[1790]&~m[1791]&m[1845])|(m[1788]&~m[1789]&m[1790]&~m[1791]&m[1845])|(~m[1788]&m[1789]&m[1790]&~m[1791]&m[1845])|(m[1788]&m[1789]&m[1790]&~m[1791]&m[1845])|(m[1788]&m[1789]&m[1790]&m[1791]&m[1845]))):InitCond[2013];
    m[1797] = run?((((m[1793]&~m[1794]&~m[1795]&~m[1796]&~m[1850])|(~m[1793]&m[1794]&~m[1795]&~m[1796]&~m[1850])|(~m[1793]&~m[1794]&m[1795]&~m[1796]&~m[1850])|(m[1793]&m[1794]&~m[1795]&m[1796]&~m[1850])|(m[1793]&~m[1794]&m[1795]&m[1796]&~m[1850])|(~m[1793]&m[1794]&m[1795]&m[1796]&~m[1850]))&BiasedRNG[1068])|(((m[1793]&~m[1794]&~m[1795]&~m[1796]&m[1850])|(~m[1793]&m[1794]&~m[1795]&~m[1796]&m[1850])|(~m[1793]&~m[1794]&m[1795]&~m[1796]&m[1850])|(m[1793]&m[1794]&~m[1795]&m[1796]&m[1850])|(m[1793]&~m[1794]&m[1795]&m[1796]&m[1850])|(~m[1793]&m[1794]&m[1795]&m[1796]&m[1850]))&~BiasedRNG[1068])|((m[1793]&m[1794]&~m[1795]&~m[1796]&~m[1850])|(m[1793]&~m[1794]&m[1795]&~m[1796]&~m[1850])|(~m[1793]&m[1794]&m[1795]&~m[1796]&~m[1850])|(m[1793]&m[1794]&m[1795]&~m[1796]&~m[1850])|(m[1793]&m[1794]&m[1795]&m[1796]&~m[1850])|(m[1793]&m[1794]&~m[1795]&~m[1796]&m[1850])|(m[1793]&~m[1794]&m[1795]&~m[1796]&m[1850])|(~m[1793]&m[1794]&m[1795]&~m[1796]&m[1850])|(m[1793]&m[1794]&m[1795]&~m[1796]&m[1850])|(m[1793]&m[1794]&m[1795]&m[1796]&m[1850]))):InitCond[2014];
    m[1802] = run?((((m[1798]&~m[1799]&~m[1800]&~m[1801]&~m[1853])|(~m[1798]&m[1799]&~m[1800]&~m[1801]&~m[1853])|(~m[1798]&~m[1799]&m[1800]&~m[1801]&~m[1853])|(m[1798]&m[1799]&~m[1800]&m[1801]&~m[1853])|(m[1798]&~m[1799]&m[1800]&m[1801]&~m[1853])|(~m[1798]&m[1799]&m[1800]&m[1801]&~m[1853]))&BiasedRNG[1069])|(((m[1798]&~m[1799]&~m[1800]&~m[1801]&m[1853])|(~m[1798]&m[1799]&~m[1800]&~m[1801]&m[1853])|(~m[1798]&~m[1799]&m[1800]&~m[1801]&m[1853])|(m[1798]&m[1799]&~m[1800]&m[1801]&m[1853])|(m[1798]&~m[1799]&m[1800]&m[1801]&m[1853])|(~m[1798]&m[1799]&m[1800]&m[1801]&m[1853]))&~BiasedRNG[1069])|((m[1798]&m[1799]&~m[1800]&~m[1801]&~m[1853])|(m[1798]&~m[1799]&m[1800]&~m[1801]&~m[1853])|(~m[1798]&m[1799]&m[1800]&~m[1801]&~m[1853])|(m[1798]&m[1799]&m[1800]&~m[1801]&~m[1853])|(m[1798]&m[1799]&m[1800]&m[1801]&~m[1853])|(m[1798]&m[1799]&~m[1800]&~m[1801]&m[1853])|(m[1798]&~m[1799]&m[1800]&~m[1801]&m[1853])|(~m[1798]&m[1799]&m[1800]&~m[1801]&m[1853])|(m[1798]&m[1799]&m[1800]&~m[1801]&m[1853])|(m[1798]&m[1799]&m[1800]&m[1801]&m[1853]))):InitCond[2015];
    m[1807] = run?((((m[1803]&~m[1804]&~m[1805]&~m[1806]&~m[1855])|(~m[1803]&m[1804]&~m[1805]&~m[1806]&~m[1855])|(~m[1803]&~m[1804]&m[1805]&~m[1806]&~m[1855])|(m[1803]&m[1804]&~m[1805]&m[1806]&~m[1855])|(m[1803]&~m[1804]&m[1805]&m[1806]&~m[1855])|(~m[1803]&m[1804]&m[1805]&m[1806]&~m[1855]))&BiasedRNG[1070])|(((m[1803]&~m[1804]&~m[1805]&~m[1806]&m[1855])|(~m[1803]&m[1804]&~m[1805]&~m[1806]&m[1855])|(~m[1803]&~m[1804]&m[1805]&~m[1806]&m[1855])|(m[1803]&m[1804]&~m[1805]&m[1806]&m[1855])|(m[1803]&~m[1804]&m[1805]&m[1806]&m[1855])|(~m[1803]&m[1804]&m[1805]&m[1806]&m[1855]))&~BiasedRNG[1070])|((m[1803]&m[1804]&~m[1805]&~m[1806]&~m[1855])|(m[1803]&~m[1804]&m[1805]&~m[1806]&~m[1855])|(~m[1803]&m[1804]&m[1805]&~m[1806]&~m[1855])|(m[1803]&m[1804]&m[1805]&~m[1806]&~m[1855])|(m[1803]&m[1804]&m[1805]&m[1806]&~m[1855])|(m[1803]&m[1804]&~m[1805]&~m[1806]&m[1855])|(m[1803]&~m[1804]&m[1805]&~m[1806]&m[1855])|(~m[1803]&m[1804]&m[1805]&~m[1806]&m[1855])|(m[1803]&m[1804]&m[1805]&~m[1806]&m[1855])|(m[1803]&m[1804]&m[1805]&m[1806]&m[1855]))):InitCond[2016];
    m[1812] = run?((((m[1808]&~m[1809]&~m[1810]&~m[1811]&~m[1860])|(~m[1808]&m[1809]&~m[1810]&~m[1811]&~m[1860])|(~m[1808]&~m[1809]&m[1810]&~m[1811]&~m[1860])|(m[1808]&m[1809]&~m[1810]&m[1811]&~m[1860])|(m[1808]&~m[1809]&m[1810]&m[1811]&~m[1860])|(~m[1808]&m[1809]&m[1810]&m[1811]&~m[1860]))&BiasedRNG[1071])|(((m[1808]&~m[1809]&~m[1810]&~m[1811]&m[1860])|(~m[1808]&m[1809]&~m[1810]&~m[1811]&m[1860])|(~m[1808]&~m[1809]&m[1810]&~m[1811]&m[1860])|(m[1808]&m[1809]&~m[1810]&m[1811]&m[1860])|(m[1808]&~m[1809]&m[1810]&m[1811]&m[1860])|(~m[1808]&m[1809]&m[1810]&m[1811]&m[1860]))&~BiasedRNG[1071])|((m[1808]&m[1809]&~m[1810]&~m[1811]&~m[1860])|(m[1808]&~m[1809]&m[1810]&~m[1811]&~m[1860])|(~m[1808]&m[1809]&m[1810]&~m[1811]&~m[1860])|(m[1808]&m[1809]&m[1810]&~m[1811]&~m[1860])|(m[1808]&m[1809]&m[1810]&m[1811]&~m[1860])|(m[1808]&m[1809]&~m[1810]&~m[1811]&m[1860])|(m[1808]&~m[1809]&m[1810]&~m[1811]&m[1860])|(~m[1808]&m[1809]&m[1810]&~m[1811]&m[1860])|(m[1808]&m[1809]&m[1810]&~m[1811]&m[1860])|(m[1808]&m[1809]&m[1810]&m[1811]&m[1860]))):InitCond[2017];
    m[1817] = run?((((m[1813]&~m[1814]&~m[1815]&~m[1816]&~m[1865])|(~m[1813]&m[1814]&~m[1815]&~m[1816]&~m[1865])|(~m[1813]&~m[1814]&m[1815]&~m[1816]&~m[1865])|(m[1813]&m[1814]&~m[1815]&m[1816]&~m[1865])|(m[1813]&~m[1814]&m[1815]&m[1816]&~m[1865])|(~m[1813]&m[1814]&m[1815]&m[1816]&~m[1865]))&BiasedRNG[1072])|(((m[1813]&~m[1814]&~m[1815]&~m[1816]&m[1865])|(~m[1813]&m[1814]&~m[1815]&~m[1816]&m[1865])|(~m[1813]&~m[1814]&m[1815]&~m[1816]&m[1865])|(m[1813]&m[1814]&~m[1815]&m[1816]&m[1865])|(m[1813]&~m[1814]&m[1815]&m[1816]&m[1865])|(~m[1813]&m[1814]&m[1815]&m[1816]&m[1865]))&~BiasedRNG[1072])|((m[1813]&m[1814]&~m[1815]&~m[1816]&~m[1865])|(m[1813]&~m[1814]&m[1815]&~m[1816]&~m[1865])|(~m[1813]&m[1814]&m[1815]&~m[1816]&~m[1865])|(m[1813]&m[1814]&m[1815]&~m[1816]&~m[1865])|(m[1813]&m[1814]&m[1815]&m[1816]&~m[1865])|(m[1813]&m[1814]&~m[1815]&~m[1816]&m[1865])|(m[1813]&~m[1814]&m[1815]&~m[1816]&m[1865])|(~m[1813]&m[1814]&m[1815]&~m[1816]&m[1865])|(m[1813]&m[1814]&m[1815]&~m[1816]&m[1865])|(m[1813]&m[1814]&m[1815]&m[1816]&m[1865]))):InitCond[2018];
    m[1822] = run?((((m[1818]&~m[1819]&~m[1820]&~m[1821]&~m[1870])|(~m[1818]&m[1819]&~m[1820]&~m[1821]&~m[1870])|(~m[1818]&~m[1819]&m[1820]&~m[1821]&~m[1870])|(m[1818]&m[1819]&~m[1820]&m[1821]&~m[1870])|(m[1818]&~m[1819]&m[1820]&m[1821]&~m[1870])|(~m[1818]&m[1819]&m[1820]&m[1821]&~m[1870]))&BiasedRNG[1073])|(((m[1818]&~m[1819]&~m[1820]&~m[1821]&m[1870])|(~m[1818]&m[1819]&~m[1820]&~m[1821]&m[1870])|(~m[1818]&~m[1819]&m[1820]&~m[1821]&m[1870])|(m[1818]&m[1819]&~m[1820]&m[1821]&m[1870])|(m[1818]&~m[1819]&m[1820]&m[1821]&m[1870])|(~m[1818]&m[1819]&m[1820]&m[1821]&m[1870]))&~BiasedRNG[1073])|((m[1818]&m[1819]&~m[1820]&~m[1821]&~m[1870])|(m[1818]&~m[1819]&m[1820]&~m[1821]&~m[1870])|(~m[1818]&m[1819]&m[1820]&~m[1821]&~m[1870])|(m[1818]&m[1819]&m[1820]&~m[1821]&~m[1870])|(m[1818]&m[1819]&m[1820]&m[1821]&~m[1870])|(m[1818]&m[1819]&~m[1820]&~m[1821]&m[1870])|(m[1818]&~m[1819]&m[1820]&~m[1821]&m[1870])|(~m[1818]&m[1819]&m[1820]&~m[1821]&m[1870])|(m[1818]&m[1819]&m[1820]&~m[1821]&m[1870])|(m[1818]&m[1819]&m[1820]&m[1821]&m[1870]))):InitCond[2019];
    m[1827] = run?((((m[1823]&~m[1824]&~m[1825]&~m[1826]&~m[1875])|(~m[1823]&m[1824]&~m[1825]&~m[1826]&~m[1875])|(~m[1823]&~m[1824]&m[1825]&~m[1826]&~m[1875])|(m[1823]&m[1824]&~m[1825]&m[1826]&~m[1875])|(m[1823]&~m[1824]&m[1825]&m[1826]&~m[1875])|(~m[1823]&m[1824]&m[1825]&m[1826]&~m[1875]))&BiasedRNG[1074])|(((m[1823]&~m[1824]&~m[1825]&~m[1826]&m[1875])|(~m[1823]&m[1824]&~m[1825]&~m[1826]&m[1875])|(~m[1823]&~m[1824]&m[1825]&~m[1826]&m[1875])|(m[1823]&m[1824]&~m[1825]&m[1826]&m[1875])|(m[1823]&~m[1824]&m[1825]&m[1826]&m[1875])|(~m[1823]&m[1824]&m[1825]&m[1826]&m[1875]))&~BiasedRNG[1074])|((m[1823]&m[1824]&~m[1825]&~m[1826]&~m[1875])|(m[1823]&~m[1824]&m[1825]&~m[1826]&~m[1875])|(~m[1823]&m[1824]&m[1825]&~m[1826]&~m[1875])|(m[1823]&m[1824]&m[1825]&~m[1826]&~m[1875])|(m[1823]&m[1824]&m[1825]&m[1826]&~m[1875])|(m[1823]&m[1824]&~m[1825]&~m[1826]&m[1875])|(m[1823]&~m[1824]&m[1825]&~m[1826]&m[1875])|(~m[1823]&m[1824]&m[1825]&~m[1826]&m[1875])|(m[1823]&m[1824]&m[1825]&~m[1826]&m[1875])|(m[1823]&m[1824]&m[1825]&m[1826]&m[1875]))):InitCond[2020];
    m[1832] = run?((((m[1828]&~m[1829]&~m[1830]&~m[1831]&~m[1880])|(~m[1828]&m[1829]&~m[1830]&~m[1831]&~m[1880])|(~m[1828]&~m[1829]&m[1830]&~m[1831]&~m[1880])|(m[1828]&m[1829]&~m[1830]&m[1831]&~m[1880])|(m[1828]&~m[1829]&m[1830]&m[1831]&~m[1880])|(~m[1828]&m[1829]&m[1830]&m[1831]&~m[1880]))&BiasedRNG[1075])|(((m[1828]&~m[1829]&~m[1830]&~m[1831]&m[1880])|(~m[1828]&m[1829]&~m[1830]&~m[1831]&m[1880])|(~m[1828]&~m[1829]&m[1830]&~m[1831]&m[1880])|(m[1828]&m[1829]&~m[1830]&m[1831]&m[1880])|(m[1828]&~m[1829]&m[1830]&m[1831]&m[1880])|(~m[1828]&m[1829]&m[1830]&m[1831]&m[1880]))&~BiasedRNG[1075])|((m[1828]&m[1829]&~m[1830]&~m[1831]&~m[1880])|(m[1828]&~m[1829]&m[1830]&~m[1831]&~m[1880])|(~m[1828]&m[1829]&m[1830]&~m[1831]&~m[1880])|(m[1828]&m[1829]&m[1830]&~m[1831]&~m[1880])|(m[1828]&m[1829]&m[1830]&m[1831]&~m[1880])|(m[1828]&m[1829]&~m[1830]&~m[1831]&m[1880])|(m[1828]&~m[1829]&m[1830]&~m[1831]&m[1880])|(~m[1828]&m[1829]&m[1830]&~m[1831]&m[1880])|(m[1828]&m[1829]&m[1830]&~m[1831]&m[1880])|(m[1828]&m[1829]&m[1830]&m[1831]&m[1880]))):InitCond[2021];
    m[1837] = run?((((m[1833]&~m[1834]&~m[1835]&~m[1836]&~m[1885])|(~m[1833]&m[1834]&~m[1835]&~m[1836]&~m[1885])|(~m[1833]&~m[1834]&m[1835]&~m[1836]&~m[1885])|(m[1833]&m[1834]&~m[1835]&m[1836]&~m[1885])|(m[1833]&~m[1834]&m[1835]&m[1836]&~m[1885])|(~m[1833]&m[1834]&m[1835]&m[1836]&~m[1885]))&BiasedRNG[1076])|(((m[1833]&~m[1834]&~m[1835]&~m[1836]&m[1885])|(~m[1833]&m[1834]&~m[1835]&~m[1836]&m[1885])|(~m[1833]&~m[1834]&m[1835]&~m[1836]&m[1885])|(m[1833]&m[1834]&~m[1835]&m[1836]&m[1885])|(m[1833]&~m[1834]&m[1835]&m[1836]&m[1885])|(~m[1833]&m[1834]&m[1835]&m[1836]&m[1885]))&~BiasedRNG[1076])|((m[1833]&m[1834]&~m[1835]&~m[1836]&~m[1885])|(m[1833]&~m[1834]&m[1835]&~m[1836]&~m[1885])|(~m[1833]&m[1834]&m[1835]&~m[1836]&~m[1885])|(m[1833]&m[1834]&m[1835]&~m[1836]&~m[1885])|(m[1833]&m[1834]&m[1835]&m[1836]&~m[1885])|(m[1833]&m[1834]&~m[1835]&~m[1836]&m[1885])|(m[1833]&~m[1834]&m[1835]&~m[1836]&m[1885])|(~m[1833]&m[1834]&m[1835]&~m[1836]&m[1885])|(m[1833]&m[1834]&m[1835]&~m[1836]&m[1885])|(m[1833]&m[1834]&m[1835]&m[1836]&m[1885]))):InitCond[2022];
    m[1842] = run?((((m[1838]&~m[1839]&~m[1840]&~m[1841]&~m[1890])|(~m[1838]&m[1839]&~m[1840]&~m[1841]&~m[1890])|(~m[1838]&~m[1839]&m[1840]&~m[1841]&~m[1890])|(m[1838]&m[1839]&~m[1840]&m[1841]&~m[1890])|(m[1838]&~m[1839]&m[1840]&m[1841]&~m[1890])|(~m[1838]&m[1839]&m[1840]&m[1841]&~m[1890]))&BiasedRNG[1077])|(((m[1838]&~m[1839]&~m[1840]&~m[1841]&m[1890])|(~m[1838]&m[1839]&~m[1840]&~m[1841]&m[1890])|(~m[1838]&~m[1839]&m[1840]&~m[1841]&m[1890])|(m[1838]&m[1839]&~m[1840]&m[1841]&m[1890])|(m[1838]&~m[1839]&m[1840]&m[1841]&m[1890])|(~m[1838]&m[1839]&m[1840]&m[1841]&m[1890]))&~BiasedRNG[1077])|((m[1838]&m[1839]&~m[1840]&~m[1841]&~m[1890])|(m[1838]&~m[1839]&m[1840]&~m[1841]&~m[1890])|(~m[1838]&m[1839]&m[1840]&~m[1841]&~m[1890])|(m[1838]&m[1839]&m[1840]&~m[1841]&~m[1890])|(m[1838]&m[1839]&m[1840]&m[1841]&~m[1890])|(m[1838]&m[1839]&~m[1840]&~m[1841]&m[1890])|(m[1838]&~m[1839]&m[1840]&~m[1841]&m[1890])|(~m[1838]&m[1839]&m[1840]&~m[1841]&m[1890])|(m[1838]&m[1839]&m[1840]&~m[1841]&m[1890])|(m[1838]&m[1839]&m[1840]&m[1841]&m[1890]))):InitCond[2023];
    m[1847] = run?((((m[1843]&~m[1844]&~m[1845]&~m[1846]&~m[1895])|(~m[1843]&m[1844]&~m[1845]&~m[1846]&~m[1895])|(~m[1843]&~m[1844]&m[1845]&~m[1846]&~m[1895])|(m[1843]&m[1844]&~m[1845]&m[1846]&~m[1895])|(m[1843]&~m[1844]&m[1845]&m[1846]&~m[1895])|(~m[1843]&m[1844]&m[1845]&m[1846]&~m[1895]))&BiasedRNG[1078])|(((m[1843]&~m[1844]&~m[1845]&~m[1846]&m[1895])|(~m[1843]&m[1844]&~m[1845]&~m[1846]&m[1895])|(~m[1843]&~m[1844]&m[1845]&~m[1846]&m[1895])|(m[1843]&m[1844]&~m[1845]&m[1846]&m[1895])|(m[1843]&~m[1844]&m[1845]&m[1846]&m[1895])|(~m[1843]&m[1844]&m[1845]&m[1846]&m[1895]))&~BiasedRNG[1078])|((m[1843]&m[1844]&~m[1845]&~m[1846]&~m[1895])|(m[1843]&~m[1844]&m[1845]&~m[1846]&~m[1895])|(~m[1843]&m[1844]&m[1845]&~m[1846]&~m[1895])|(m[1843]&m[1844]&m[1845]&~m[1846]&~m[1895])|(m[1843]&m[1844]&m[1845]&m[1846]&~m[1895])|(m[1843]&m[1844]&~m[1845]&~m[1846]&m[1895])|(m[1843]&~m[1844]&m[1845]&~m[1846]&m[1895])|(~m[1843]&m[1844]&m[1845]&~m[1846]&m[1895])|(m[1843]&m[1844]&m[1845]&~m[1846]&m[1895])|(m[1843]&m[1844]&m[1845]&m[1846]&m[1895]))):InitCond[2024];
    m[1852] = run?((((m[1848]&~m[1849]&~m[1850]&~m[1851]&~m[1900])|(~m[1848]&m[1849]&~m[1850]&~m[1851]&~m[1900])|(~m[1848]&~m[1849]&m[1850]&~m[1851]&~m[1900])|(m[1848]&m[1849]&~m[1850]&m[1851]&~m[1900])|(m[1848]&~m[1849]&m[1850]&m[1851]&~m[1900])|(~m[1848]&m[1849]&m[1850]&m[1851]&~m[1900]))&BiasedRNG[1079])|(((m[1848]&~m[1849]&~m[1850]&~m[1851]&m[1900])|(~m[1848]&m[1849]&~m[1850]&~m[1851]&m[1900])|(~m[1848]&~m[1849]&m[1850]&~m[1851]&m[1900])|(m[1848]&m[1849]&~m[1850]&m[1851]&m[1900])|(m[1848]&~m[1849]&m[1850]&m[1851]&m[1900])|(~m[1848]&m[1849]&m[1850]&m[1851]&m[1900]))&~BiasedRNG[1079])|((m[1848]&m[1849]&~m[1850]&~m[1851]&~m[1900])|(m[1848]&~m[1849]&m[1850]&~m[1851]&~m[1900])|(~m[1848]&m[1849]&m[1850]&~m[1851]&~m[1900])|(m[1848]&m[1849]&m[1850]&~m[1851]&~m[1900])|(m[1848]&m[1849]&m[1850]&m[1851]&~m[1900])|(m[1848]&m[1849]&~m[1850]&~m[1851]&m[1900])|(m[1848]&~m[1849]&m[1850]&~m[1851]&m[1900])|(~m[1848]&m[1849]&m[1850]&~m[1851]&m[1900])|(m[1848]&m[1849]&m[1850]&~m[1851]&m[1900])|(m[1848]&m[1849]&m[1850]&m[1851]&m[1900]))):InitCond[2025];
    m[1857] = run?((((m[1853]&~m[1854]&~m[1855]&~m[1856]&~m[1903])|(~m[1853]&m[1854]&~m[1855]&~m[1856]&~m[1903])|(~m[1853]&~m[1854]&m[1855]&~m[1856]&~m[1903])|(m[1853]&m[1854]&~m[1855]&m[1856]&~m[1903])|(m[1853]&~m[1854]&m[1855]&m[1856]&~m[1903])|(~m[1853]&m[1854]&m[1855]&m[1856]&~m[1903]))&BiasedRNG[1080])|(((m[1853]&~m[1854]&~m[1855]&~m[1856]&m[1903])|(~m[1853]&m[1854]&~m[1855]&~m[1856]&m[1903])|(~m[1853]&~m[1854]&m[1855]&~m[1856]&m[1903])|(m[1853]&m[1854]&~m[1855]&m[1856]&m[1903])|(m[1853]&~m[1854]&m[1855]&m[1856]&m[1903])|(~m[1853]&m[1854]&m[1855]&m[1856]&m[1903]))&~BiasedRNG[1080])|((m[1853]&m[1854]&~m[1855]&~m[1856]&~m[1903])|(m[1853]&~m[1854]&m[1855]&~m[1856]&~m[1903])|(~m[1853]&m[1854]&m[1855]&~m[1856]&~m[1903])|(m[1853]&m[1854]&m[1855]&~m[1856]&~m[1903])|(m[1853]&m[1854]&m[1855]&m[1856]&~m[1903])|(m[1853]&m[1854]&~m[1855]&~m[1856]&m[1903])|(m[1853]&~m[1854]&m[1855]&~m[1856]&m[1903])|(~m[1853]&m[1854]&m[1855]&~m[1856]&m[1903])|(m[1853]&m[1854]&m[1855]&~m[1856]&m[1903])|(m[1853]&m[1854]&m[1855]&m[1856]&m[1903]))):InitCond[2026];
    m[1862] = run?((((m[1858]&~m[1859]&~m[1860]&~m[1861]&~m[1905])|(~m[1858]&m[1859]&~m[1860]&~m[1861]&~m[1905])|(~m[1858]&~m[1859]&m[1860]&~m[1861]&~m[1905])|(m[1858]&m[1859]&~m[1860]&m[1861]&~m[1905])|(m[1858]&~m[1859]&m[1860]&m[1861]&~m[1905])|(~m[1858]&m[1859]&m[1860]&m[1861]&~m[1905]))&BiasedRNG[1081])|(((m[1858]&~m[1859]&~m[1860]&~m[1861]&m[1905])|(~m[1858]&m[1859]&~m[1860]&~m[1861]&m[1905])|(~m[1858]&~m[1859]&m[1860]&~m[1861]&m[1905])|(m[1858]&m[1859]&~m[1860]&m[1861]&m[1905])|(m[1858]&~m[1859]&m[1860]&m[1861]&m[1905])|(~m[1858]&m[1859]&m[1860]&m[1861]&m[1905]))&~BiasedRNG[1081])|((m[1858]&m[1859]&~m[1860]&~m[1861]&~m[1905])|(m[1858]&~m[1859]&m[1860]&~m[1861]&~m[1905])|(~m[1858]&m[1859]&m[1860]&~m[1861]&~m[1905])|(m[1858]&m[1859]&m[1860]&~m[1861]&~m[1905])|(m[1858]&m[1859]&m[1860]&m[1861]&~m[1905])|(m[1858]&m[1859]&~m[1860]&~m[1861]&m[1905])|(m[1858]&~m[1859]&m[1860]&~m[1861]&m[1905])|(~m[1858]&m[1859]&m[1860]&~m[1861]&m[1905])|(m[1858]&m[1859]&m[1860]&~m[1861]&m[1905])|(m[1858]&m[1859]&m[1860]&m[1861]&m[1905]))):InitCond[2027];
    m[1867] = run?((((m[1863]&~m[1864]&~m[1865]&~m[1866]&~m[1910])|(~m[1863]&m[1864]&~m[1865]&~m[1866]&~m[1910])|(~m[1863]&~m[1864]&m[1865]&~m[1866]&~m[1910])|(m[1863]&m[1864]&~m[1865]&m[1866]&~m[1910])|(m[1863]&~m[1864]&m[1865]&m[1866]&~m[1910])|(~m[1863]&m[1864]&m[1865]&m[1866]&~m[1910]))&BiasedRNG[1082])|(((m[1863]&~m[1864]&~m[1865]&~m[1866]&m[1910])|(~m[1863]&m[1864]&~m[1865]&~m[1866]&m[1910])|(~m[1863]&~m[1864]&m[1865]&~m[1866]&m[1910])|(m[1863]&m[1864]&~m[1865]&m[1866]&m[1910])|(m[1863]&~m[1864]&m[1865]&m[1866]&m[1910])|(~m[1863]&m[1864]&m[1865]&m[1866]&m[1910]))&~BiasedRNG[1082])|((m[1863]&m[1864]&~m[1865]&~m[1866]&~m[1910])|(m[1863]&~m[1864]&m[1865]&~m[1866]&~m[1910])|(~m[1863]&m[1864]&m[1865]&~m[1866]&~m[1910])|(m[1863]&m[1864]&m[1865]&~m[1866]&~m[1910])|(m[1863]&m[1864]&m[1865]&m[1866]&~m[1910])|(m[1863]&m[1864]&~m[1865]&~m[1866]&m[1910])|(m[1863]&~m[1864]&m[1865]&~m[1866]&m[1910])|(~m[1863]&m[1864]&m[1865]&~m[1866]&m[1910])|(m[1863]&m[1864]&m[1865]&~m[1866]&m[1910])|(m[1863]&m[1864]&m[1865]&m[1866]&m[1910]))):InitCond[2028];
    m[1872] = run?((((m[1868]&~m[1869]&~m[1870]&~m[1871]&~m[1915])|(~m[1868]&m[1869]&~m[1870]&~m[1871]&~m[1915])|(~m[1868]&~m[1869]&m[1870]&~m[1871]&~m[1915])|(m[1868]&m[1869]&~m[1870]&m[1871]&~m[1915])|(m[1868]&~m[1869]&m[1870]&m[1871]&~m[1915])|(~m[1868]&m[1869]&m[1870]&m[1871]&~m[1915]))&BiasedRNG[1083])|(((m[1868]&~m[1869]&~m[1870]&~m[1871]&m[1915])|(~m[1868]&m[1869]&~m[1870]&~m[1871]&m[1915])|(~m[1868]&~m[1869]&m[1870]&~m[1871]&m[1915])|(m[1868]&m[1869]&~m[1870]&m[1871]&m[1915])|(m[1868]&~m[1869]&m[1870]&m[1871]&m[1915])|(~m[1868]&m[1869]&m[1870]&m[1871]&m[1915]))&~BiasedRNG[1083])|((m[1868]&m[1869]&~m[1870]&~m[1871]&~m[1915])|(m[1868]&~m[1869]&m[1870]&~m[1871]&~m[1915])|(~m[1868]&m[1869]&m[1870]&~m[1871]&~m[1915])|(m[1868]&m[1869]&m[1870]&~m[1871]&~m[1915])|(m[1868]&m[1869]&m[1870]&m[1871]&~m[1915])|(m[1868]&m[1869]&~m[1870]&~m[1871]&m[1915])|(m[1868]&~m[1869]&m[1870]&~m[1871]&m[1915])|(~m[1868]&m[1869]&m[1870]&~m[1871]&m[1915])|(m[1868]&m[1869]&m[1870]&~m[1871]&m[1915])|(m[1868]&m[1869]&m[1870]&m[1871]&m[1915]))):InitCond[2029];
    m[1877] = run?((((m[1873]&~m[1874]&~m[1875]&~m[1876]&~m[1920])|(~m[1873]&m[1874]&~m[1875]&~m[1876]&~m[1920])|(~m[1873]&~m[1874]&m[1875]&~m[1876]&~m[1920])|(m[1873]&m[1874]&~m[1875]&m[1876]&~m[1920])|(m[1873]&~m[1874]&m[1875]&m[1876]&~m[1920])|(~m[1873]&m[1874]&m[1875]&m[1876]&~m[1920]))&BiasedRNG[1084])|(((m[1873]&~m[1874]&~m[1875]&~m[1876]&m[1920])|(~m[1873]&m[1874]&~m[1875]&~m[1876]&m[1920])|(~m[1873]&~m[1874]&m[1875]&~m[1876]&m[1920])|(m[1873]&m[1874]&~m[1875]&m[1876]&m[1920])|(m[1873]&~m[1874]&m[1875]&m[1876]&m[1920])|(~m[1873]&m[1874]&m[1875]&m[1876]&m[1920]))&~BiasedRNG[1084])|((m[1873]&m[1874]&~m[1875]&~m[1876]&~m[1920])|(m[1873]&~m[1874]&m[1875]&~m[1876]&~m[1920])|(~m[1873]&m[1874]&m[1875]&~m[1876]&~m[1920])|(m[1873]&m[1874]&m[1875]&~m[1876]&~m[1920])|(m[1873]&m[1874]&m[1875]&m[1876]&~m[1920])|(m[1873]&m[1874]&~m[1875]&~m[1876]&m[1920])|(m[1873]&~m[1874]&m[1875]&~m[1876]&m[1920])|(~m[1873]&m[1874]&m[1875]&~m[1876]&m[1920])|(m[1873]&m[1874]&m[1875]&~m[1876]&m[1920])|(m[1873]&m[1874]&m[1875]&m[1876]&m[1920]))):InitCond[2030];
    m[1882] = run?((((m[1878]&~m[1879]&~m[1880]&~m[1881]&~m[1925])|(~m[1878]&m[1879]&~m[1880]&~m[1881]&~m[1925])|(~m[1878]&~m[1879]&m[1880]&~m[1881]&~m[1925])|(m[1878]&m[1879]&~m[1880]&m[1881]&~m[1925])|(m[1878]&~m[1879]&m[1880]&m[1881]&~m[1925])|(~m[1878]&m[1879]&m[1880]&m[1881]&~m[1925]))&BiasedRNG[1085])|(((m[1878]&~m[1879]&~m[1880]&~m[1881]&m[1925])|(~m[1878]&m[1879]&~m[1880]&~m[1881]&m[1925])|(~m[1878]&~m[1879]&m[1880]&~m[1881]&m[1925])|(m[1878]&m[1879]&~m[1880]&m[1881]&m[1925])|(m[1878]&~m[1879]&m[1880]&m[1881]&m[1925])|(~m[1878]&m[1879]&m[1880]&m[1881]&m[1925]))&~BiasedRNG[1085])|((m[1878]&m[1879]&~m[1880]&~m[1881]&~m[1925])|(m[1878]&~m[1879]&m[1880]&~m[1881]&~m[1925])|(~m[1878]&m[1879]&m[1880]&~m[1881]&~m[1925])|(m[1878]&m[1879]&m[1880]&~m[1881]&~m[1925])|(m[1878]&m[1879]&m[1880]&m[1881]&~m[1925])|(m[1878]&m[1879]&~m[1880]&~m[1881]&m[1925])|(m[1878]&~m[1879]&m[1880]&~m[1881]&m[1925])|(~m[1878]&m[1879]&m[1880]&~m[1881]&m[1925])|(m[1878]&m[1879]&m[1880]&~m[1881]&m[1925])|(m[1878]&m[1879]&m[1880]&m[1881]&m[1925]))):InitCond[2031];
    m[1887] = run?((((m[1883]&~m[1884]&~m[1885]&~m[1886]&~m[1930])|(~m[1883]&m[1884]&~m[1885]&~m[1886]&~m[1930])|(~m[1883]&~m[1884]&m[1885]&~m[1886]&~m[1930])|(m[1883]&m[1884]&~m[1885]&m[1886]&~m[1930])|(m[1883]&~m[1884]&m[1885]&m[1886]&~m[1930])|(~m[1883]&m[1884]&m[1885]&m[1886]&~m[1930]))&BiasedRNG[1086])|(((m[1883]&~m[1884]&~m[1885]&~m[1886]&m[1930])|(~m[1883]&m[1884]&~m[1885]&~m[1886]&m[1930])|(~m[1883]&~m[1884]&m[1885]&~m[1886]&m[1930])|(m[1883]&m[1884]&~m[1885]&m[1886]&m[1930])|(m[1883]&~m[1884]&m[1885]&m[1886]&m[1930])|(~m[1883]&m[1884]&m[1885]&m[1886]&m[1930]))&~BiasedRNG[1086])|((m[1883]&m[1884]&~m[1885]&~m[1886]&~m[1930])|(m[1883]&~m[1884]&m[1885]&~m[1886]&~m[1930])|(~m[1883]&m[1884]&m[1885]&~m[1886]&~m[1930])|(m[1883]&m[1884]&m[1885]&~m[1886]&~m[1930])|(m[1883]&m[1884]&m[1885]&m[1886]&~m[1930])|(m[1883]&m[1884]&~m[1885]&~m[1886]&m[1930])|(m[1883]&~m[1884]&m[1885]&~m[1886]&m[1930])|(~m[1883]&m[1884]&m[1885]&~m[1886]&m[1930])|(m[1883]&m[1884]&m[1885]&~m[1886]&m[1930])|(m[1883]&m[1884]&m[1885]&m[1886]&m[1930]))):InitCond[2032];
    m[1892] = run?((((m[1888]&~m[1889]&~m[1890]&~m[1891]&~m[1935])|(~m[1888]&m[1889]&~m[1890]&~m[1891]&~m[1935])|(~m[1888]&~m[1889]&m[1890]&~m[1891]&~m[1935])|(m[1888]&m[1889]&~m[1890]&m[1891]&~m[1935])|(m[1888]&~m[1889]&m[1890]&m[1891]&~m[1935])|(~m[1888]&m[1889]&m[1890]&m[1891]&~m[1935]))&BiasedRNG[1087])|(((m[1888]&~m[1889]&~m[1890]&~m[1891]&m[1935])|(~m[1888]&m[1889]&~m[1890]&~m[1891]&m[1935])|(~m[1888]&~m[1889]&m[1890]&~m[1891]&m[1935])|(m[1888]&m[1889]&~m[1890]&m[1891]&m[1935])|(m[1888]&~m[1889]&m[1890]&m[1891]&m[1935])|(~m[1888]&m[1889]&m[1890]&m[1891]&m[1935]))&~BiasedRNG[1087])|((m[1888]&m[1889]&~m[1890]&~m[1891]&~m[1935])|(m[1888]&~m[1889]&m[1890]&~m[1891]&~m[1935])|(~m[1888]&m[1889]&m[1890]&~m[1891]&~m[1935])|(m[1888]&m[1889]&m[1890]&~m[1891]&~m[1935])|(m[1888]&m[1889]&m[1890]&m[1891]&~m[1935])|(m[1888]&m[1889]&~m[1890]&~m[1891]&m[1935])|(m[1888]&~m[1889]&m[1890]&~m[1891]&m[1935])|(~m[1888]&m[1889]&m[1890]&~m[1891]&m[1935])|(m[1888]&m[1889]&m[1890]&~m[1891]&m[1935])|(m[1888]&m[1889]&m[1890]&m[1891]&m[1935]))):InitCond[2033];
    m[1897] = run?((((m[1893]&~m[1894]&~m[1895]&~m[1896]&~m[1940])|(~m[1893]&m[1894]&~m[1895]&~m[1896]&~m[1940])|(~m[1893]&~m[1894]&m[1895]&~m[1896]&~m[1940])|(m[1893]&m[1894]&~m[1895]&m[1896]&~m[1940])|(m[1893]&~m[1894]&m[1895]&m[1896]&~m[1940])|(~m[1893]&m[1894]&m[1895]&m[1896]&~m[1940]))&BiasedRNG[1088])|(((m[1893]&~m[1894]&~m[1895]&~m[1896]&m[1940])|(~m[1893]&m[1894]&~m[1895]&~m[1896]&m[1940])|(~m[1893]&~m[1894]&m[1895]&~m[1896]&m[1940])|(m[1893]&m[1894]&~m[1895]&m[1896]&m[1940])|(m[1893]&~m[1894]&m[1895]&m[1896]&m[1940])|(~m[1893]&m[1894]&m[1895]&m[1896]&m[1940]))&~BiasedRNG[1088])|((m[1893]&m[1894]&~m[1895]&~m[1896]&~m[1940])|(m[1893]&~m[1894]&m[1895]&~m[1896]&~m[1940])|(~m[1893]&m[1894]&m[1895]&~m[1896]&~m[1940])|(m[1893]&m[1894]&m[1895]&~m[1896]&~m[1940])|(m[1893]&m[1894]&m[1895]&m[1896]&~m[1940])|(m[1893]&m[1894]&~m[1895]&~m[1896]&m[1940])|(m[1893]&~m[1894]&m[1895]&~m[1896]&m[1940])|(~m[1893]&m[1894]&m[1895]&~m[1896]&m[1940])|(m[1893]&m[1894]&m[1895]&~m[1896]&m[1940])|(m[1893]&m[1894]&m[1895]&m[1896]&m[1940]))):InitCond[2034];
    m[1902] = run?((((m[1898]&~m[1899]&~m[1900]&~m[1901]&~m[1945])|(~m[1898]&m[1899]&~m[1900]&~m[1901]&~m[1945])|(~m[1898]&~m[1899]&m[1900]&~m[1901]&~m[1945])|(m[1898]&m[1899]&~m[1900]&m[1901]&~m[1945])|(m[1898]&~m[1899]&m[1900]&m[1901]&~m[1945])|(~m[1898]&m[1899]&m[1900]&m[1901]&~m[1945]))&BiasedRNG[1089])|(((m[1898]&~m[1899]&~m[1900]&~m[1901]&m[1945])|(~m[1898]&m[1899]&~m[1900]&~m[1901]&m[1945])|(~m[1898]&~m[1899]&m[1900]&~m[1901]&m[1945])|(m[1898]&m[1899]&~m[1900]&m[1901]&m[1945])|(m[1898]&~m[1899]&m[1900]&m[1901]&m[1945])|(~m[1898]&m[1899]&m[1900]&m[1901]&m[1945]))&~BiasedRNG[1089])|((m[1898]&m[1899]&~m[1900]&~m[1901]&~m[1945])|(m[1898]&~m[1899]&m[1900]&~m[1901]&~m[1945])|(~m[1898]&m[1899]&m[1900]&~m[1901]&~m[1945])|(m[1898]&m[1899]&m[1900]&~m[1901]&~m[1945])|(m[1898]&m[1899]&m[1900]&m[1901]&~m[1945])|(m[1898]&m[1899]&~m[1900]&~m[1901]&m[1945])|(m[1898]&~m[1899]&m[1900]&~m[1901]&m[1945])|(~m[1898]&m[1899]&m[1900]&~m[1901]&m[1945])|(m[1898]&m[1899]&m[1900]&~m[1901]&m[1945])|(m[1898]&m[1899]&m[1900]&m[1901]&m[1945]))):InitCond[2035];
    m[1907] = run?((((m[1903]&~m[1904]&~m[1905]&~m[1906]&~m[1948])|(~m[1903]&m[1904]&~m[1905]&~m[1906]&~m[1948])|(~m[1903]&~m[1904]&m[1905]&~m[1906]&~m[1948])|(m[1903]&m[1904]&~m[1905]&m[1906]&~m[1948])|(m[1903]&~m[1904]&m[1905]&m[1906]&~m[1948])|(~m[1903]&m[1904]&m[1905]&m[1906]&~m[1948]))&BiasedRNG[1090])|(((m[1903]&~m[1904]&~m[1905]&~m[1906]&m[1948])|(~m[1903]&m[1904]&~m[1905]&~m[1906]&m[1948])|(~m[1903]&~m[1904]&m[1905]&~m[1906]&m[1948])|(m[1903]&m[1904]&~m[1905]&m[1906]&m[1948])|(m[1903]&~m[1904]&m[1905]&m[1906]&m[1948])|(~m[1903]&m[1904]&m[1905]&m[1906]&m[1948]))&~BiasedRNG[1090])|((m[1903]&m[1904]&~m[1905]&~m[1906]&~m[1948])|(m[1903]&~m[1904]&m[1905]&~m[1906]&~m[1948])|(~m[1903]&m[1904]&m[1905]&~m[1906]&~m[1948])|(m[1903]&m[1904]&m[1905]&~m[1906]&~m[1948])|(m[1903]&m[1904]&m[1905]&m[1906]&~m[1948])|(m[1903]&m[1904]&~m[1905]&~m[1906]&m[1948])|(m[1903]&~m[1904]&m[1905]&~m[1906]&m[1948])|(~m[1903]&m[1904]&m[1905]&~m[1906]&m[1948])|(m[1903]&m[1904]&m[1905]&~m[1906]&m[1948])|(m[1903]&m[1904]&m[1905]&m[1906]&m[1948]))):InitCond[2036];
    m[1912] = run?((((m[1908]&~m[1909]&~m[1910]&~m[1911]&~m[1950])|(~m[1908]&m[1909]&~m[1910]&~m[1911]&~m[1950])|(~m[1908]&~m[1909]&m[1910]&~m[1911]&~m[1950])|(m[1908]&m[1909]&~m[1910]&m[1911]&~m[1950])|(m[1908]&~m[1909]&m[1910]&m[1911]&~m[1950])|(~m[1908]&m[1909]&m[1910]&m[1911]&~m[1950]))&BiasedRNG[1091])|(((m[1908]&~m[1909]&~m[1910]&~m[1911]&m[1950])|(~m[1908]&m[1909]&~m[1910]&~m[1911]&m[1950])|(~m[1908]&~m[1909]&m[1910]&~m[1911]&m[1950])|(m[1908]&m[1909]&~m[1910]&m[1911]&m[1950])|(m[1908]&~m[1909]&m[1910]&m[1911]&m[1950])|(~m[1908]&m[1909]&m[1910]&m[1911]&m[1950]))&~BiasedRNG[1091])|((m[1908]&m[1909]&~m[1910]&~m[1911]&~m[1950])|(m[1908]&~m[1909]&m[1910]&~m[1911]&~m[1950])|(~m[1908]&m[1909]&m[1910]&~m[1911]&~m[1950])|(m[1908]&m[1909]&m[1910]&~m[1911]&~m[1950])|(m[1908]&m[1909]&m[1910]&m[1911]&~m[1950])|(m[1908]&m[1909]&~m[1910]&~m[1911]&m[1950])|(m[1908]&~m[1909]&m[1910]&~m[1911]&m[1950])|(~m[1908]&m[1909]&m[1910]&~m[1911]&m[1950])|(m[1908]&m[1909]&m[1910]&~m[1911]&m[1950])|(m[1908]&m[1909]&m[1910]&m[1911]&m[1950]))):InitCond[2037];
    m[1917] = run?((((m[1913]&~m[1914]&~m[1915]&~m[1916]&~m[1955])|(~m[1913]&m[1914]&~m[1915]&~m[1916]&~m[1955])|(~m[1913]&~m[1914]&m[1915]&~m[1916]&~m[1955])|(m[1913]&m[1914]&~m[1915]&m[1916]&~m[1955])|(m[1913]&~m[1914]&m[1915]&m[1916]&~m[1955])|(~m[1913]&m[1914]&m[1915]&m[1916]&~m[1955]))&BiasedRNG[1092])|(((m[1913]&~m[1914]&~m[1915]&~m[1916]&m[1955])|(~m[1913]&m[1914]&~m[1915]&~m[1916]&m[1955])|(~m[1913]&~m[1914]&m[1915]&~m[1916]&m[1955])|(m[1913]&m[1914]&~m[1915]&m[1916]&m[1955])|(m[1913]&~m[1914]&m[1915]&m[1916]&m[1955])|(~m[1913]&m[1914]&m[1915]&m[1916]&m[1955]))&~BiasedRNG[1092])|((m[1913]&m[1914]&~m[1915]&~m[1916]&~m[1955])|(m[1913]&~m[1914]&m[1915]&~m[1916]&~m[1955])|(~m[1913]&m[1914]&m[1915]&~m[1916]&~m[1955])|(m[1913]&m[1914]&m[1915]&~m[1916]&~m[1955])|(m[1913]&m[1914]&m[1915]&m[1916]&~m[1955])|(m[1913]&m[1914]&~m[1915]&~m[1916]&m[1955])|(m[1913]&~m[1914]&m[1915]&~m[1916]&m[1955])|(~m[1913]&m[1914]&m[1915]&~m[1916]&m[1955])|(m[1913]&m[1914]&m[1915]&~m[1916]&m[1955])|(m[1913]&m[1914]&m[1915]&m[1916]&m[1955]))):InitCond[2038];
    m[1922] = run?((((m[1918]&~m[1919]&~m[1920]&~m[1921]&~m[1960])|(~m[1918]&m[1919]&~m[1920]&~m[1921]&~m[1960])|(~m[1918]&~m[1919]&m[1920]&~m[1921]&~m[1960])|(m[1918]&m[1919]&~m[1920]&m[1921]&~m[1960])|(m[1918]&~m[1919]&m[1920]&m[1921]&~m[1960])|(~m[1918]&m[1919]&m[1920]&m[1921]&~m[1960]))&BiasedRNG[1093])|(((m[1918]&~m[1919]&~m[1920]&~m[1921]&m[1960])|(~m[1918]&m[1919]&~m[1920]&~m[1921]&m[1960])|(~m[1918]&~m[1919]&m[1920]&~m[1921]&m[1960])|(m[1918]&m[1919]&~m[1920]&m[1921]&m[1960])|(m[1918]&~m[1919]&m[1920]&m[1921]&m[1960])|(~m[1918]&m[1919]&m[1920]&m[1921]&m[1960]))&~BiasedRNG[1093])|((m[1918]&m[1919]&~m[1920]&~m[1921]&~m[1960])|(m[1918]&~m[1919]&m[1920]&~m[1921]&~m[1960])|(~m[1918]&m[1919]&m[1920]&~m[1921]&~m[1960])|(m[1918]&m[1919]&m[1920]&~m[1921]&~m[1960])|(m[1918]&m[1919]&m[1920]&m[1921]&~m[1960])|(m[1918]&m[1919]&~m[1920]&~m[1921]&m[1960])|(m[1918]&~m[1919]&m[1920]&~m[1921]&m[1960])|(~m[1918]&m[1919]&m[1920]&~m[1921]&m[1960])|(m[1918]&m[1919]&m[1920]&~m[1921]&m[1960])|(m[1918]&m[1919]&m[1920]&m[1921]&m[1960]))):InitCond[2039];
    m[1927] = run?((((m[1923]&~m[1924]&~m[1925]&~m[1926]&~m[1965])|(~m[1923]&m[1924]&~m[1925]&~m[1926]&~m[1965])|(~m[1923]&~m[1924]&m[1925]&~m[1926]&~m[1965])|(m[1923]&m[1924]&~m[1925]&m[1926]&~m[1965])|(m[1923]&~m[1924]&m[1925]&m[1926]&~m[1965])|(~m[1923]&m[1924]&m[1925]&m[1926]&~m[1965]))&BiasedRNG[1094])|(((m[1923]&~m[1924]&~m[1925]&~m[1926]&m[1965])|(~m[1923]&m[1924]&~m[1925]&~m[1926]&m[1965])|(~m[1923]&~m[1924]&m[1925]&~m[1926]&m[1965])|(m[1923]&m[1924]&~m[1925]&m[1926]&m[1965])|(m[1923]&~m[1924]&m[1925]&m[1926]&m[1965])|(~m[1923]&m[1924]&m[1925]&m[1926]&m[1965]))&~BiasedRNG[1094])|((m[1923]&m[1924]&~m[1925]&~m[1926]&~m[1965])|(m[1923]&~m[1924]&m[1925]&~m[1926]&~m[1965])|(~m[1923]&m[1924]&m[1925]&~m[1926]&~m[1965])|(m[1923]&m[1924]&m[1925]&~m[1926]&~m[1965])|(m[1923]&m[1924]&m[1925]&m[1926]&~m[1965])|(m[1923]&m[1924]&~m[1925]&~m[1926]&m[1965])|(m[1923]&~m[1924]&m[1925]&~m[1926]&m[1965])|(~m[1923]&m[1924]&m[1925]&~m[1926]&m[1965])|(m[1923]&m[1924]&m[1925]&~m[1926]&m[1965])|(m[1923]&m[1924]&m[1925]&m[1926]&m[1965]))):InitCond[2040];
    m[1932] = run?((((m[1928]&~m[1929]&~m[1930]&~m[1931]&~m[1970])|(~m[1928]&m[1929]&~m[1930]&~m[1931]&~m[1970])|(~m[1928]&~m[1929]&m[1930]&~m[1931]&~m[1970])|(m[1928]&m[1929]&~m[1930]&m[1931]&~m[1970])|(m[1928]&~m[1929]&m[1930]&m[1931]&~m[1970])|(~m[1928]&m[1929]&m[1930]&m[1931]&~m[1970]))&BiasedRNG[1095])|(((m[1928]&~m[1929]&~m[1930]&~m[1931]&m[1970])|(~m[1928]&m[1929]&~m[1930]&~m[1931]&m[1970])|(~m[1928]&~m[1929]&m[1930]&~m[1931]&m[1970])|(m[1928]&m[1929]&~m[1930]&m[1931]&m[1970])|(m[1928]&~m[1929]&m[1930]&m[1931]&m[1970])|(~m[1928]&m[1929]&m[1930]&m[1931]&m[1970]))&~BiasedRNG[1095])|((m[1928]&m[1929]&~m[1930]&~m[1931]&~m[1970])|(m[1928]&~m[1929]&m[1930]&~m[1931]&~m[1970])|(~m[1928]&m[1929]&m[1930]&~m[1931]&~m[1970])|(m[1928]&m[1929]&m[1930]&~m[1931]&~m[1970])|(m[1928]&m[1929]&m[1930]&m[1931]&~m[1970])|(m[1928]&m[1929]&~m[1930]&~m[1931]&m[1970])|(m[1928]&~m[1929]&m[1930]&~m[1931]&m[1970])|(~m[1928]&m[1929]&m[1930]&~m[1931]&m[1970])|(m[1928]&m[1929]&m[1930]&~m[1931]&m[1970])|(m[1928]&m[1929]&m[1930]&m[1931]&m[1970]))):InitCond[2041];
    m[1937] = run?((((m[1933]&~m[1934]&~m[1935]&~m[1936]&~m[1975])|(~m[1933]&m[1934]&~m[1935]&~m[1936]&~m[1975])|(~m[1933]&~m[1934]&m[1935]&~m[1936]&~m[1975])|(m[1933]&m[1934]&~m[1935]&m[1936]&~m[1975])|(m[1933]&~m[1934]&m[1935]&m[1936]&~m[1975])|(~m[1933]&m[1934]&m[1935]&m[1936]&~m[1975]))&BiasedRNG[1096])|(((m[1933]&~m[1934]&~m[1935]&~m[1936]&m[1975])|(~m[1933]&m[1934]&~m[1935]&~m[1936]&m[1975])|(~m[1933]&~m[1934]&m[1935]&~m[1936]&m[1975])|(m[1933]&m[1934]&~m[1935]&m[1936]&m[1975])|(m[1933]&~m[1934]&m[1935]&m[1936]&m[1975])|(~m[1933]&m[1934]&m[1935]&m[1936]&m[1975]))&~BiasedRNG[1096])|((m[1933]&m[1934]&~m[1935]&~m[1936]&~m[1975])|(m[1933]&~m[1934]&m[1935]&~m[1936]&~m[1975])|(~m[1933]&m[1934]&m[1935]&~m[1936]&~m[1975])|(m[1933]&m[1934]&m[1935]&~m[1936]&~m[1975])|(m[1933]&m[1934]&m[1935]&m[1936]&~m[1975])|(m[1933]&m[1934]&~m[1935]&~m[1936]&m[1975])|(m[1933]&~m[1934]&m[1935]&~m[1936]&m[1975])|(~m[1933]&m[1934]&m[1935]&~m[1936]&m[1975])|(m[1933]&m[1934]&m[1935]&~m[1936]&m[1975])|(m[1933]&m[1934]&m[1935]&m[1936]&m[1975]))):InitCond[2042];
    m[1942] = run?((((m[1938]&~m[1939]&~m[1940]&~m[1941]&~m[1980])|(~m[1938]&m[1939]&~m[1940]&~m[1941]&~m[1980])|(~m[1938]&~m[1939]&m[1940]&~m[1941]&~m[1980])|(m[1938]&m[1939]&~m[1940]&m[1941]&~m[1980])|(m[1938]&~m[1939]&m[1940]&m[1941]&~m[1980])|(~m[1938]&m[1939]&m[1940]&m[1941]&~m[1980]))&BiasedRNG[1097])|(((m[1938]&~m[1939]&~m[1940]&~m[1941]&m[1980])|(~m[1938]&m[1939]&~m[1940]&~m[1941]&m[1980])|(~m[1938]&~m[1939]&m[1940]&~m[1941]&m[1980])|(m[1938]&m[1939]&~m[1940]&m[1941]&m[1980])|(m[1938]&~m[1939]&m[1940]&m[1941]&m[1980])|(~m[1938]&m[1939]&m[1940]&m[1941]&m[1980]))&~BiasedRNG[1097])|((m[1938]&m[1939]&~m[1940]&~m[1941]&~m[1980])|(m[1938]&~m[1939]&m[1940]&~m[1941]&~m[1980])|(~m[1938]&m[1939]&m[1940]&~m[1941]&~m[1980])|(m[1938]&m[1939]&m[1940]&~m[1941]&~m[1980])|(m[1938]&m[1939]&m[1940]&m[1941]&~m[1980])|(m[1938]&m[1939]&~m[1940]&~m[1941]&m[1980])|(m[1938]&~m[1939]&m[1940]&~m[1941]&m[1980])|(~m[1938]&m[1939]&m[1940]&~m[1941]&m[1980])|(m[1938]&m[1939]&m[1940]&~m[1941]&m[1980])|(m[1938]&m[1939]&m[1940]&m[1941]&m[1980]))):InitCond[2043];
    m[1947] = run?((((m[1943]&~m[1944]&~m[1945]&~m[1946]&~m[1985])|(~m[1943]&m[1944]&~m[1945]&~m[1946]&~m[1985])|(~m[1943]&~m[1944]&m[1945]&~m[1946]&~m[1985])|(m[1943]&m[1944]&~m[1945]&m[1946]&~m[1985])|(m[1943]&~m[1944]&m[1945]&m[1946]&~m[1985])|(~m[1943]&m[1944]&m[1945]&m[1946]&~m[1985]))&BiasedRNG[1098])|(((m[1943]&~m[1944]&~m[1945]&~m[1946]&m[1985])|(~m[1943]&m[1944]&~m[1945]&~m[1946]&m[1985])|(~m[1943]&~m[1944]&m[1945]&~m[1946]&m[1985])|(m[1943]&m[1944]&~m[1945]&m[1946]&m[1985])|(m[1943]&~m[1944]&m[1945]&m[1946]&m[1985])|(~m[1943]&m[1944]&m[1945]&m[1946]&m[1985]))&~BiasedRNG[1098])|((m[1943]&m[1944]&~m[1945]&~m[1946]&~m[1985])|(m[1943]&~m[1944]&m[1945]&~m[1946]&~m[1985])|(~m[1943]&m[1944]&m[1945]&~m[1946]&~m[1985])|(m[1943]&m[1944]&m[1945]&~m[1946]&~m[1985])|(m[1943]&m[1944]&m[1945]&m[1946]&~m[1985])|(m[1943]&m[1944]&~m[1945]&~m[1946]&m[1985])|(m[1943]&~m[1944]&m[1945]&~m[1946]&m[1985])|(~m[1943]&m[1944]&m[1945]&~m[1946]&m[1985])|(m[1943]&m[1944]&m[1945]&~m[1946]&m[1985])|(m[1943]&m[1944]&m[1945]&m[1946]&m[1985]))):InitCond[2044];
    m[1952] = run?((((m[1948]&~m[1949]&~m[1950]&~m[1951]&~m[1988])|(~m[1948]&m[1949]&~m[1950]&~m[1951]&~m[1988])|(~m[1948]&~m[1949]&m[1950]&~m[1951]&~m[1988])|(m[1948]&m[1949]&~m[1950]&m[1951]&~m[1988])|(m[1948]&~m[1949]&m[1950]&m[1951]&~m[1988])|(~m[1948]&m[1949]&m[1950]&m[1951]&~m[1988]))&BiasedRNG[1099])|(((m[1948]&~m[1949]&~m[1950]&~m[1951]&m[1988])|(~m[1948]&m[1949]&~m[1950]&~m[1951]&m[1988])|(~m[1948]&~m[1949]&m[1950]&~m[1951]&m[1988])|(m[1948]&m[1949]&~m[1950]&m[1951]&m[1988])|(m[1948]&~m[1949]&m[1950]&m[1951]&m[1988])|(~m[1948]&m[1949]&m[1950]&m[1951]&m[1988]))&~BiasedRNG[1099])|((m[1948]&m[1949]&~m[1950]&~m[1951]&~m[1988])|(m[1948]&~m[1949]&m[1950]&~m[1951]&~m[1988])|(~m[1948]&m[1949]&m[1950]&~m[1951]&~m[1988])|(m[1948]&m[1949]&m[1950]&~m[1951]&~m[1988])|(m[1948]&m[1949]&m[1950]&m[1951]&~m[1988])|(m[1948]&m[1949]&~m[1950]&~m[1951]&m[1988])|(m[1948]&~m[1949]&m[1950]&~m[1951]&m[1988])|(~m[1948]&m[1949]&m[1950]&~m[1951]&m[1988])|(m[1948]&m[1949]&m[1950]&~m[1951]&m[1988])|(m[1948]&m[1949]&m[1950]&m[1951]&m[1988]))):InitCond[2045];
    m[1957] = run?((((m[1953]&~m[1954]&~m[1955]&~m[1956]&~m[1990])|(~m[1953]&m[1954]&~m[1955]&~m[1956]&~m[1990])|(~m[1953]&~m[1954]&m[1955]&~m[1956]&~m[1990])|(m[1953]&m[1954]&~m[1955]&m[1956]&~m[1990])|(m[1953]&~m[1954]&m[1955]&m[1956]&~m[1990])|(~m[1953]&m[1954]&m[1955]&m[1956]&~m[1990]))&BiasedRNG[1100])|(((m[1953]&~m[1954]&~m[1955]&~m[1956]&m[1990])|(~m[1953]&m[1954]&~m[1955]&~m[1956]&m[1990])|(~m[1953]&~m[1954]&m[1955]&~m[1956]&m[1990])|(m[1953]&m[1954]&~m[1955]&m[1956]&m[1990])|(m[1953]&~m[1954]&m[1955]&m[1956]&m[1990])|(~m[1953]&m[1954]&m[1955]&m[1956]&m[1990]))&~BiasedRNG[1100])|((m[1953]&m[1954]&~m[1955]&~m[1956]&~m[1990])|(m[1953]&~m[1954]&m[1955]&~m[1956]&~m[1990])|(~m[1953]&m[1954]&m[1955]&~m[1956]&~m[1990])|(m[1953]&m[1954]&m[1955]&~m[1956]&~m[1990])|(m[1953]&m[1954]&m[1955]&m[1956]&~m[1990])|(m[1953]&m[1954]&~m[1955]&~m[1956]&m[1990])|(m[1953]&~m[1954]&m[1955]&~m[1956]&m[1990])|(~m[1953]&m[1954]&m[1955]&~m[1956]&m[1990])|(m[1953]&m[1954]&m[1955]&~m[1956]&m[1990])|(m[1953]&m[1954]&m[1955]&m[1956]&m[1990]))):InitCond[2046];
    m[1962] = run?((((m[1958]&~m[1959]&~m[1960]&~m[1961]&~m[1995])|(~m[1958]&m[1959]&~m[1960]&~m[1961]&~m[1995])|(~m[1958]&~m[1959]&m[1960]&~m[1961]&~m[1995])|(m[1958]&m[1959]&~m[1960]&m[1961]&~m[1995])|(m[1958]&~m[1959]&m[1960]&m[1961]&~m[1995])|(~m[1958]&m[1959]&m[1960]&m[1961]&~m[1995]))&BiasedRNG[1101])|(((m[1958]&~m[1959]&~m[1960]&~m[1961]&m[1995])|(~m[1958]&m[1959]&~m[1960]&~m[1961]&m[1995])|(~m[1958]&~m[1959]&m[1960]&~m[1961]&m[1995])|(m[1958]&m[1959]&~m[1960]&m[1961]&m[1995])|(m[1958]&~m[1959]&m[1960]&m[1961]&m[1995])|(~m[1958]&m[1959]&m[1960]&m[1961]&m[1995]))&~BiasedRNG[1101])|((m[1958]&m[1959]&~m[1960]&~m[1961]&~m[1995])|(m[1958]&~m[1959]&m[1960]&~m[1961]&~m[1995])|(~m[1958]&m[1959]&m[1960]&~m[1961]&~m[1995])|(m[1958]&m[1959]&m[1960]&~m[1961]&~m[1995])|(m[1958]&m[1959]&m[1960]&m[1961]&~m[1995])|(m[1958]&m[1959]&~m[1960]&~m[1961]&m[1995])|(m[1958]&~m[1959]&m[1960]&~m[1961]&m[1995])|(~m[1958]&m[1959]&m[1960]&~m[1961]&m[1995])|(m[1958]&m[1959]&m[1960]&~m[1961]&m[1995])|(m[1958]&m[1959]&m[1960]&m[1961]&m[1995]))):InitCond[2047];
    m[1967] = run?((((m[1963]&~m[1964]&~m[1965]&~m[1966]&~m[2000])|(~m[1963]&m[1964]&~m[1965]&~m[1966]&~m[2000])|(~m[1963]&~m[1964]&m[1965]&~m[1966]&~m[2000])|(m[1963]&m[1964]&~m[1965]&m[1966]&~m[2000])|(m[1963]&~m[1964]&m[1965]&m[1966]&~m[2000])|(~m[1963]&m[1964]&m[1965]&m[1966]&~m[2000]))&BiasedRNG[1102])|(((m[1963]&~m[1964]&~m[1965]&~m[1966]&m[2000])|(~m[1963]&m[1964]&~m[1965]&~m[1966]&m[2000])|(~m[1963]&~m[1964]&m[1965]&~m[1966]&m[2000])|(m[1963]&m[1964]&~m[1965]&m[1966]&m[2000])|(m[1963]&~m[1964]&m[1965]&m[1966]&m[2000])|(~m[1963]&m[1964]&m[1965]&m[1966]&m[2000]))&~BiasedRNG[1102])|((m[1963]&m[1964]&~m[1965]&~m[1966]&~m[2000])|(m[1963]&~m[1964]&m[1965]&~m[1966]&~m[2000])|(~m[1963]&m[1964]&m[1965]&~m[1966]&~m[2000])|(m[1963]&m[1964]&m[1965]&~m[1966]&~m[2000])|(m[1963]&m[1964]&m[1965]&m[1966]&~m[2000])|(m[1963]&m[1964]&~m[1965]&~m[1966]&m[2000])|(m[1963]&~m[1964]&m[1965]&~m[1966]&m[2000])|(~m[1963]&m[1964]&m[1965]&~m[1966]&m[2000])|(m[1963]&m[1964]&m[1965]&~m[1966]&m[2000])|(m[1963]&m[1964]&m[1965]&m[1966]&m[2000]))):InitCond[2048];
    m[1972] = run?((((m[1968]&~m[1969]&~m[1970]&~m[1971]&~m[2005])|(~m[1968]&m[1969]&~m[1970]&~m[1971]&~m[2005])|(~m[1968]&~m[1969]&m[1970]&~m[1971]&~m[2005])|(m[1968]&m[1969]&~m[1970]&m[1971]&~m[2005])|(m[1968]&~m[1969]&m[1970]&m[1971]&~m[2005])|(~m[1968]&m[1969]&m[1970]&m[1971]&~m[2005]))&BiasedRNG[1103])|(((m[1968]&~m[1969]&~m[1970]&~m[1971]&m[2005])|(~m[1968]&m[1969]&~m[1970]&~m[1971]&m[2005])|(~m[1968]&~m[1969]&m[1970]&~m[1971]&m[2005])|(m[1968]&m[1969]&~m[1970]&m[1971]&m[2005])|(m[1968]&~m[1969]&m[1970]&m[1971]&m[2005])|(~m[1968]&m[1969]&m[1970]&m[1971]&m[2005]))&~BiasedRNG[1103])|((m[1968]&m[1969]&~m[1970]&~m[1971]&~m[2005])|(m[1968]&~m[1969]&m[1970]&~m[1971]&~m[2005])|(~m[1968]&m[1969]&m[1970]&~m[1971]&~m[2005])|(m[1968]&m[1969]&m[1970]&~m[1971]&~m[2005])|(m[1968]&m[1969]&m[1970]&m[1971]&~m[2005])|(m[1968]&m[1969]&~m[1970]&~m[1971]&m[2005])|(m[1968]&~m[1969]&m[1970]&~m[1971]&m[2005])|(~m[1968]&m[1969]&m[1970]&~m[1971]&m[2005])|(m[1968]&m[1969]&m[1970]&~m[1971]&m[2005])|(m[1968]&m[1969]&m[1970]&m[1971]&m[2005]))):InitCond[2049];
    m[1977] = run?((((m[1973]&~m[1974]&~m[1975]&~m[1976]&~m[2010])|(~m[1973]&m[1974]&~m[1975]&~m[1976]&~m[2010])|(~m[1973]&~m[1974]&m[1975]&~m[1976]&~m[2010])|(m[1973]&m[1974]&~m[1975]&m[1976]&~m[2010])|(m[1973]&~m[1974]&m[1975]&m[1976]&~m[2010])|(~m[1973]&m[1974]&m[1975]&m[1976]&~m[2010]))&BiasedRNG[1104])|(((m[1973]&~m[1974]&~m[1975]&~m[1976]&m[2010])|(~m[1973]&m[1974]&~m[1975]&~m[1976]&m[2010])|(~m[1973]&~m[1974]&m[1975]&~m[1976]&m[2010])|(m[1973]&m[1974]&~m[1975]&m[1976]&m[2010])|(m[1973]&~m[1974]&m[1975]&m[1976]&m[2010])|(~m[1973]&m[1974]&m[1975]&m[1976]&m[2010]))&~BiasedRNG[1104])|((m[1973]&m[1974]&~m[1975]&~m[1976]&~m[2010])|(m[1973]&~m[1974]&m[1975]&~m[1976]&~m[2010])|(~m[1973]&m[1974]&m[1975]&~m[1976]&~m[2010])|(m[1973]&m[1974]&m[1975]&~m[1976]&~m[2010])|(m[1973]&m[1974]&m[1975]&m[1976]&~m[2010])|(m[1973]&m[1974]&~m[1975]&~m[1976]&m[2010])|(m[1973]&~m[1974]&m[1975]&~m[1976]&m[2010])|(~m[1973]&m[1974]&m[1975]&~m[1976]&m[2010])|(m[1973]&m[1974]&m[1975]&~m[1976]&m[2010])|(m[1973]&m[1974]&m[1975]&m[1976]&m[2010]))):InitCond[2050];
    m[1982] = run?((((m[1978]&~m[1979]&~m[1980]&~m[1981]&~m[2015])|(~m[1978]&m[1979]&~m[1980]&~m[1981]&~m[2015])|(~m[1978]&~m[1979]&m[1980]&~m[1981]&~m[2015])|(m[1978]&m[1979]&~m[1980]&m[1981]&~m[2015])|(m[1978]&~m[1979]&m[1980]&m[1981]&~m[2015])|(~m[1978]&m[1979]&m[1980]&m[1981]&~m[2015]))&BiasedRNG[1105])|(((m[1978]&~m[1979]&~m[1980]&~m[1981]&m[2015])|(~m[1978]&m[1979]&~m[1980]&~m[1981]&m[2015])|(~m[1978]&~m[1979]&m[1980]&~m[1981]&m[2015])|(m[1978]&m[1979]&~m[1980]&m[1981]&m[2015])|(m[1978]&~m[1979]&m[1980]&m[1981]&m[2015])|(~m[1978]&m[1979]&m[1980]&m[1981]&m[2015]))&~BiasedRNG[1105])|((m[1978]&m[1979]&~m[1980]&~m[1981]&~m[2015])|(m[1978]&~m[1979]&m[1980]&~m[1981]&~m[2015])|(~m[1978]&m[1979]&m[1980]&~m[1981]&~m[2015])|(m[1978]&m[1979]&m[1980]&~m[1981]&~m[2015])|(m[1978]&m[1979]&m[1980]&m[1981]&~m[2015])|(m[1978]&m[1979]&~m[1980]&~m[1981]&m[2015])|(m[1978]&~m[1979]&m[1980]&~m[1981]&m[2015])|(~m[1978]&m[1979]&m[1980]&~m[1981]&m[2015])|(m[1978]&m[1979]&m[1980]&~m[1981]&m[2015])|(m[1978]&m[1979]&m[1980]&m[1981]&m[2015]))):InitCond[2051];
    m[1987] = run?((((m[1983]&~m[1984]&~m[1985]&~m[1986]&~m[2020])|(~m[1983]&m[1984]&~m[1985]&~m[1986]&~m[2020])|(~m[1983]&~m[1984]&m[1985]&~m[1986]&~m[2020])|(m[1983]&m[1984]&~m[1985]&m[1986]&~m[2020])|(m[1983]&~m[1984]&m[1985]&m[1986]&~m[2020])|(~m[1983]&m[1984]&m[1985]&m[1986]&~m[2020]))&BiasedRNG[1106])|(((m[1983]&~m[1984]&~m[1985]&~m[1986]&m[2020])|(~m[1983]&m[1984]&~m[1985]&~m[1986]&m[2020])|(~m[1983]&~m[1984]&m[1985]&~m[1986]&m[2020])|(m[1983]&m[1984]&~m[1985]&m[1986]&m[2020])|(m[1983]&~m[1984]&m[1985]&m[1986]&m[2020])|(~m[1983]&m[1984]&m[1985]&m[1986]&m[2020]))&~BiasedRNG[1106])|((m[1983]&m[1984]&~m[1985]&~m[1986]&~m[2020])|(m[1983]&~m[1984]&m[1985]&~m[1986]&~m[2020])|(~m[1983]&m[1984]&m[1985]&~m[1986]&~m[2020])|(m[1983]&m[1984]&m[1985]&~m[1986]&~m[2020])|(m[1983]&m[1984]&m[1985]&m[1986]&~m[2020])|(m[1983]&m[1984]&~m[1985]&~m[1986]&m[2020])|(m[1983]&~m[1984]&m[1985]&~m[1986]&m[2020])|(~m[1983]&m[1984]&m[1985]&~m[1986]&m[2020])|(m[1983]&m[1984]&m[1985]&~m[1986]&m[2020])|(m[1983]&m[1984]&m[1985]&m[1986]&m[2020]))):InitCond[2052];
    m[1992] = run?((((m[1988]&~m[1989]&~m[1990]&~m[1991]&~m[2023])|(~m[1988]&m[1989]&~m[1990]&~m[1991]&~m[2023])|(~m[1988]&~m[1989]&m[1990]&~m[1991]&~m[2023])|(m[1988]&m[1989]&~m[1990]&m[1991]&~m[2023])|(m[1988]&~m[1989]&m[1990]&m[1991]&~m[2023])|(~m[1988]&m[1989]&m[1990]&m[1991]&~m[2023]))&BiasedRNG[1107])|(((m[1988]&~m[1989]&~m[1990]&~m[1991]&m[2023])|(~m[1988]&m[1989]&~m[1990]&~m[1991]&m[2023])|(~m[1988]&~m[1989]&m[1990]&~m[1991]&m[2023])|(m[1988]&m[1989]&~m[1990]&m[1991]&m[2023])|(m[1988]&~m[1989]&m[1990]&m[1991]&m[2023])|(~m[1988]&m[1989]&m[1990]&m[1991]&m[2023]))&~BiasedRNG[1107])|((m[1988]&m[1989]&~m[1990]&~m[1991]&~m[2023])|(m[1988]&~m[1989]&m[1990]&~m[1991]&~m[2023])|(~m[1988]&m[1989]&m[1990]&~m[1991]&~m[2023])|(m[1988]&m[1989]&m[1990]&~m[1991]&~m[2023])|(m[1988]&m[1989]&m[1990]&m[1991]&~m[2023])|(m[1988]&m[1989]&~m[1990]&~m[1991]&m[2023])|(m[1988]&~m[1989]&m[1990]&~m[1991]&m[2023])|(~m[1988]&m[1989]&m[1990]&~m[1991]&m[2023])|(m[1988]&m[1989]&m[1990]&~m[1991]&m[2023])|(m[1988]&m[1989]&m[1990]&m[1991]&m[2023]))):InitCond[2053];
    m[1997] = run?((((m[1993]&~m[1994]&~m[1995]&~m[1996]&~m[2025])|(~m[1993]&m[1994]&~m[1995]&~m[1996]&~m[2025])|(~m[1993]&~m[1994]&m[1995]&~m[1996]&~m[2025])|(m[1993]&m[1994]&~m[1995]&m[1996]&~m[2025])|(m[1993]&~m[1994]&m[1995]&m[1996]&~m[2025])|(~m[1993]&m[1994]&m[1995]&m[1996]&~m[2025]))&BiasedRNG[1108])|(((m[1993]&~m[1994]&~m[1995]&~m[1996]&m[2025])|(~m[1993]&m[1994]&~m[1995]&~m[1996]&m[2025])|(~m[1993]&~m[1994]&m[1995]&~m[1996]&m[2025])|(m[1993]&m[1994]&~m[1995]&m[1996]&m[2025])|(m[1993]&~m[1994]&m[1995]&m[1996]&m[2025])|(~m[1993]&m[1994]&m[1995]&m[1996]&m[2025]))&~BiasedRNG[1108])|((m[1993]&m[1994]&~m[1995]&~m[1996]&~m[2025])|(m[1993]&~m[1994]&m[1995]&~m[1996]&~m[2025])|(~m[1993]&m[1994]&m[1995]&~m[1996]&~m[2025])|(m[1993]&m[1994]&m[1995]&~m[1996]&~m[2025])|(m[1993]&m[1994]&m[1995]&m[1996]&~m[2025])|(m[1993]&m[1994]&~m[1995]&~m[1996]&m[2025])|(m[1993]&~m[1994]&m[1995]&~m[1996]&m[2025])|(~m[1993]&m[1994]&m[1995]&~m[1996]&m[2025])|(m[1993]&m[1994]&m[1995]&~m[1996]&m[2025])|(m[1993]&m[1994]&m[1995]&m[1996]&m[2025]))):InitCond[2054];
    m[2002] = run?((((m[1998]&~m[1999]&~m[2000]&~m[2001]&~m[2030])|(~m[1998]&m[1999]&~m[2000]&~m[2001]&~m[2030])|(~m[1998]&~m[1999]&m[2000]&~m[2001]&~m[2030])|(m[1998]&m[1999]&~m[2000]&m[2001]&~m[2030])|(m[1998]&~m[1999]&m[2000]&m[2001]&~m[2030])|(~m[1998]&m[1999]&m[2000]&m[2001]&~m[2030]))&BiasedRNG[1109])|(((m[1998]&~m[1999]&~m[2000]&~m[2001]&m[2030])|(~m[1998]&m[1999]&~m[2000]&~m[2001]&m[2030])|(~m[1998]&~m[1999]&m[2000]&~m[2001]&m[2030])|(m[1998]&m[1999]&~m[2000]&m[2001]&m[2030])|(m[1998]&~m[1999]&m[2000]&m[2001]&m[2030])|(~m[1998]&m[1999]&m[2000]&m[2001]&m[2030]))&~BiasedRNG[1109])|((m[1998]&m[1999]&~m[2000]&~m[2001]&~m[2030])|(m[1998]&~m[1999]&m[2000]&~m[2001]&~m[2030])|(~m[1998]&m[1999]&m[2000]&~m[2001]&~m[2030])|(m[1998]&m[1999]&m[2000]&~m[2001]&~m[2030])|(m[1998]&m[1999]&m[2000]&m[2001]&~m[2030])|(m[1998]&m[1999]&~m[2000]&~m[2001]&m[2030])|(m[1998]&~m[1999]&m[2000]&~m[2001]&m[2030])|(~m[1998]&m[1999]&m[2000]&~m[2001]&m[2030])|(m[1998]&m[1999]&m[2000]&~m[2001]&m[2030])|(m[1998]&m[1999]&m[2000]&m[2001]&m[2030]))):InitCond[2055];
    m[2007] = run?((((m[2003]&~m[2004]&~m[2005]&~m[2006]&~m[2035])|(~m[2003]&m[2004]&~m[2005]&~m[2006]&~m[2035])|(~m[2003]&~m[2004]&m[2005]&~m[2006]&~m[2035])|(m[2003]&m[2004]&~m[2005]&m[2006]&~m[2035])|(m[2003]&~m[2004]&m[2005]&m[2006]&~m[2035])|(~m[2003]&m[2004]&m[2005]&m[2006]&~m[2035]))&BiasedRNG[1110])|(((m[2003]&~m[2004]&~m[2005]&~m[2006]&m[2035])|(~m[2003]&m[2004]&~m[2005]&~m[2006]&m[2035])|(~m[2003]&~m[2004]&m[2005]&~m[2006]&m[2035])|(m[2003]&m[2004]&~m[2005]&m[2006]&m[2035])|(m[2003]&~m[2004]&m[2005]&m[2006]&m[2035])|(~m[2003]&m[2004]&m[2005]&m[2006]&m[2035]))&~BiasedRNG[1110])|((m[2003]&m[2004]&~m[2005]&~m[2006]&~m[2035])|(m[2003]&~m[2004]&m[2005]&~m[2006]&~m[2035])|(~m[2003]&m[2004]&m[2005]&~m[2006]&~m[2035])|(m[2003]&m[2004]&m[2005]&~m[2006]&~m[2035])|(m[2003]&m[2004]&m[2005]&m[2006]&~m[2035])|(m[2003]&m[2004]&~m[2005]&~m[2006]&m[2035])|(m[2003]&~m[2004]&m[2005]&~m[2006]&m[2035])|(~m[2003]&m[2004]&m[2005]&~m[2006]&m[2035])|(m[2003]&m[2004]&m[2005]&~m[2006]&m[2035])|(m[2003]&m[2004]&m[2005]&m[2006]&m[2035]))):InitCond[2056];
    m[2012] = run?((((m[2008]&~m[2009]&~m[2010]&~m[2011]&~m[2040])|(~m[2008]&m[2009]&~m[2010]&~m[2011]&~m[2040])|(~m[2008]&~m[2009]&m[2010]&~m[2011]&~m[2040])|(m[2008]&m[2009]&~m[2010]&m[2011]&~m[2040])|(m[2008]&~m[2009]&m[2010]&m[2011]&~m[2040])|(~m[2008]&m[2009]&m[2010]&m[2011]&~m[2040]))&BiasedRNG[1111])|(((m[2008]&~m[2009]&~m[2010]&~m[2011]&m[2040])|(~m[2008]&m[2009]&~m[2010]&~m[2011]&m[2040])|(~m[2008]&~m[2009]&m[2010]&~m[2011]&m[2040])|(m[2008]&m[2009]&~m[2010]&m[2011]&m[2040])|(m[2008]&~m[2009]&m[2010]&m[2011]&m[2040])|(~m[2008]&m[2009]&m[2010]&m[2011]&m[2040]))&~BiasedRNG[1111])|((m[2008]&m[2009]&~m[2010]&~m[2011]&~m[2040])|(m[2008]&~m[2009]&m[2010]&~m[2011]&~m[2040])|(~m[2008]&m[2009]&m[2010]&~m[2011]&~m[2040])|(m[2008]&m[2009]&m[2010]&~m[2011]&~m[2040])|(m[2008]&m[2009]&m[2010]&m[2011]&~m[2040])|(m[2008]&m[2009]&~m[2010]&~m[2011]&m[2040])|(m[2008]&~m[2009]&m[2010]&~m[2011]&m[2040])|(~m[2008]&m[2009]&m[2010]&~m[2011]&m[2040])|(m[2008]&m[2009]&m[2010]&~m[2011]&m[2040])|(m[2008]&m[2009]&m[2010]&m[2011]&m[2040]))):InitCond[2057];
    m[2017] = run?((((m[2013]&~m[2014]&~m[2015]&~m[2016]&~m[2045])|(~m[2013]&m[2014]&~m[2015]&~m[2016]&~m[2045])|(~m[2013]&~m[2014]&m[2015]&~m[2016]&~m[2045])|(m[2013]&m[2014]&~m[2015]&m[2016]&~m[2045])|(m[2013]&~m[2014]&m[2015]&m[2016]&~m[2045])|(~m[2013]&m[2014]&m[2015]&m[2016]&~m[2045]))&BiasedRNG[1112])|(((m[2013]&~m[2014]&~m[2015]&~m[2016]&m[2045])|(~m[2013]&m[2014]&~m[2015]&~m[2016]&m[2045])|(~m[2013]&~m[2014]&m[2015]&~m[2016]&m[2045])|(m[2013]&m[2014]&~m[2015]&m[2016]&m[2045])|(m[2013]&~m[2014]&m[2015]&m[2016]&m[2045])|(~m[2013]&m[2014]&m[2015]&m[2016]&m[2045]))&~BiasedRNG[1112])|((m[2013]&m[2014]&~m[2015]&~m[2016]&~m[2045])|(m[2013]&~m[2014]&m[2015]&~m[2016]&~m[2045])|(~m[2013]&m[2014]&m[2015]&~m[2016]&~m[2045])|(m[2013]&m[2014]&m[2015]&~m[2016]&~m[2045])|(m[2013]&m[2014]&m[2015]&m[2016]&~m[2045])|(m[2013]&m[2014]&~m[2015]&~m[2016]&m[2045])|(m[2013]&~m[2014]&m[2015]&~m[2016]&m[2045])|(~m[2013]&m[2014]&m[2015]&~m[2016]&m[2045])|(m[2013]&m[2014]&m[2015]&~m[2016]&m[2045])|(m[2013]&m[2014]&m[2015]&m[2016]&m[2045]))):InitCond[2058];
    m[2022] = run?((((m[2018]&~m[2019]&~m[2020]&~m[2021]&~m[2050])|(~m[2018]&m[2019]&~m[2020]&~m[2021]&~m[2050])|(~m[2018]&~m[2019]&m[2020]&~m[2021]&~m[2050])|(m[2018]&m[2019]&~m[2020]&m[2021]&~m[2050])|(m[2018]&~m[2019]&m[2020]&m[2021]&~m[2050])|(~m[2018]&m[2019]&m[2020]&m[2021]&~m[2050]))&BiasedRNG[1113])|(((m[2018]&~m[2019]&~m[2020]&~m[2021]&m[2050])|(~m[2018]&m[2019]&~m[2020]&~m[2021]&m[2050])|(~m[2018]&~m[2019]&m[2020]&~m[2021]&m[2050])|(m[2018]&m[2019]&~m[2020]&m[2021]&m[2050])|(m[2018]&~m[2019]&m[2020]&m[2021]&m[2050])|(~m[2018]&m[2019]&m[2020]&m[2021]&m[2050]))&~BiasedRNG[1113])|((m[2018]&m[2019]&~m[2020]&~m[2021]&~m[2050])|(m[2018]&~m[2019]&m[2020]&~m[2021]&~m[2050])|(~m[2018]&m[2019]&m[2020]&~m[2021]&~m[2050])|(m[2018]&m[2019]&m[2020]&~m[2021]&~m[2050])|(m[2018]&m[2019]&m[2020]&m[2021]&~m[2050])|(m[2018]&m[2019]&~m[2020]&~m[2021]&m[2050])|(m[2018]&~m[2019]&m[2020]&~m[2021]&m[2050])|(~m[2018]&m[2019]&m[2020]&~m[2021]&m[2050])|(m[2018]&m[2019]&m[2020]&~m[2021]&m[2050])|(m[2018]&m[2019]&m[2020]&m[2021]&m[2050]))):InitCond[2059];
    m[2027] = run?((((m[2023]&~m[2024]&~m[2025]&~m[2026]&~m[2053])|(~m[2023]&m[2024]&~m[2025]&~m[2026]&~m[2053])|(~m[2023]&~m[2024]&m[2025]&~m[2026]&~m[2053])|(m[2023]&m[2024]&~m[2025]&m[2026]&~m[2053])|(m[2023]&~m[2024]&m[2025]&m[2026]&~m[2053])|(~m[2023]&m[2024]&m[2025]&m[2026]&~m[2053]))&BiasedRNG[1114])|(((m[2023]&~m[2024]&~m[2025]&~m[2026]&m[2053])|(~m[2023]&m[2024]&~m[2025]&~m[2026]&m[2053])|(~m[2023]&~m[2024]&m[2025]&~m[2026]&m[2053])|(m[2023]&m[2024]&~m[2025]&m[2026]&m[2053])|(m[2023]&~m[2024]&m[2025]&m[2026]&m[2053])|(~m[2023]&m[2024]&m[2025]&m[2026]&m[2053]))&~BiasedRNG[1114])|((m[2023]&m[2024]&~m[2025]&~m[2026]&~m[2053])|(m[2023]&~m[2024]&m[2025]&~m[2026]&~m[2053])|(~m[2023]&m[2024]&m[2025]&~m[2026]&~m[2053])|(m[2023]&m[2024]&m[2025]&~m[2026]&~m[2053])|(m[2023]&m[2024]&m[2025]&m[2026]&~m[2053])|(m[2023]&m[2024]&~m[2025]&~m[2026]&m[2053])|(m[2023]&~m[2024]&m[2025]&~m[2026]&m[2053])|(~m[2023]&m[2024]&m[2025]&~m[2026]&m[2053])|(m[2023]&m[2024]&m[2025]&~m[2026]&m[2053])|(m[2023]&m[2024]&m[2025]&m[2026]&m[2053]))):InitCond[2060];
    m[2032] = run?((((m[2028]&~m[2029]&~m[2030]&~m[2031]&~m[2055])|(~m[2028]&m[2029]&~m[2030]&~m[2031]&~m[2055])|(~m[2028]&~m[2029]&m[2030]&~m[2031]&~m[2055])|(m[2028]&m[2029]&~m[2030]&m[2031]&~m[2055])|(m[2028]&~m[2029]&m[2030]&m[2031]&~m[2055])|(~m[2028]&m[2029]&m[2030]&m[2031]&~m[2055]))&BiasedRNG[1115])|(((m[2028]&~m[2029]&~m[2030]&~m[2031]&m[2055])|(~m[2028]&m[2029]&~m[2030]&~m[2031]&m[2055])|(~m[2028]&~m[2029]&m[2030]&~m[2031]&m[2055])|(m[2028]&m[2029]&~m[2030]&m[2031]&m[2055])|(m[2028]&~m[2029]&m[2030]&m[2031]&m[2055])|(~m[2028]&m[2029]&m[2030]&m[2031]&m[2055]))&~BiasedRNG[1115])|((m[2028]&m[2029]&~m[2030]&~m[2031]&~m[2055])|(m[2028]&~m[2029]&m[2030]&~m[2031]&~m[2055])|(~m[2028]&m[2029]&m[2030]&~m[2031]&~m[2055])|(m[2028]&m[2029]&m[2030]&~m[2031]&~m[2055])|(m[2028]&m[2029]&m[2030]&m[2031]&~m[2055])|(m[2028]&m[2029]&~m[2030]&~m[2031]&m[2055])|(m[2028]&~m[2029]&m[2030]&~m[2031]&m[2055])|(~m[2028]&m[2029]&m[2030]&~m[2031]&m[2055])|(m[2028]&m[2029]&m[2030]&~m[2031]&m[2055])|(m[2028]&m[2029]&m[2030]&m[2031]&m[2055]))):InitCond[2061];
    m[2037] = run?((((m[2033]&~m[2034]&~m[2035]&~m[2036]&~m[2060])|(~m[2033]&m[2034]&~m[2035]&~m[2036]&~m[2060])|(~m[2033]&~m[2034]&m[2035]&~m[2036]&~m[2060])|(m[2033]&m[2034]&~m[2035]&m[2036]&~m[2060])|(m[2033]&~m[2034]&m[2035]&m[2036]&~m[2060])|(~m[2033]&m[2034]&m[2035]&m[2036]&~m[2060]))&BiasedRNG[1116])|(((m[2033]&~m[2034]&~m[2035]&~m[2036]&m[2060])|(~m[2033]&m[2034]&~m[2035]&~m[2036]&m[2060])|(~m[2033]&~m[2034]&m[2035]&~m[2036]&m[2060])|(m[2033]&m[2034]&~m[2035]&m[2036]&m[2060])|(m[2033]&~m[2034]&m[2035]&m[2036]&m[2060])|(~m[2033]&m[2034]&m[2035]&m[2036]&m[2060]))&~BiasedRNG[1116])|((m[2033]&m[2034]&~m[2035]&~m[2036]&~m[2060])|(m[2033]&~m[2034]&m[2035]&~m[2036]&~m[2060])|(~m[2033]&m[2034]&m[2035]&~m[2036]&~m[2060])|(m[2033]&m[2034]&m[2035]&~m[2036]&~m[2060])|(m[2033]&m[2034]&m[2035]&m[2036]&~m[2060])|(m[2033]&m[2034]&~m[2035]&~m[2036]&m[2060])|(m[2033]&~m[2034]&m[2035]&~m[2036]&m[2060])|(~m[2033]&m[2034]&m[2035]&~m[2036]&m[2060])|(m[2033]&m[2034]&m[2035]&~m[2036]&m[2060])|(m[2033]&m[2034]&m[2035]&m[2036]&m[2060]))):InitCond[2062];
    m[2042] = run?((((m[2038]&~m[2039]&~m[2040]&~m[2041]&~m[2065])|(~m[2038]&m[2039]&~m[2040]&~m[2041]&~m[2065])|(~m[2038]&~m[2039]&m[2040]&~m[2041]&~m[2065])|(m[2038]&m[2039]&~m[2040]&m[2041]&~m[2065])|(m[2038]&~m[2039]&m[2040]&m[2041]&~m[2065])|(~m[2038]&m[2039]&m[2040]&m[2041]&~m[2065]))&BiasedRNG[1117])|(((m[2038]&~m[2039]&~m[2040]&~m[2041]&m[2065])|(~m[2038]&m[2039]&~m[2040]&~m[2041]&m[2065])|(~m[2038]&~m[2039]&m[2040]&~m[2041]&m[2065])|(m[2038]&m[2039]&~m[2040]&m[2041]&m[2065])|(m[2038]&~m[2039]&m[2040]&m[2041]&m[2065])|(~m[2038]&m[2039]&m[2040]&m[2041]&m[2065]))&~BiasedRNG[1117])|((m[2038]&m[2039]&~m[2040]&~m[2041]&~m[2065])|(m[2038]&~m[2039]&m[2040]&~m[2041]&~m[2065])|(~m[2038]&m[2039]&m[2040]&~m[2041]&~m[2065])|(m[2038]&m[2039]&m[2040]&~m[2041]&~m[2065])|(m[2038]&m[2039]&m[2040]&m[2041]&~m[2065])|(m[2038]&m[2039]&~m[2040]&~m[2041]&m[2065])|(m[2038]&~m[2039]&m[2040]&~m[2041]&m[2065])|(~m[2038]&m[2039]&m[2040]&~m[2041]&m[2065])|(m[2038]&m[2039]&m[2040]&~m[2041]&m[2065])|(m[2038]&m[2039]&m[2040]&m[2041]&m[2065]))):InitCond[2063];
    m[2047] = run?((((m[2043]&~m[2044]&~m[2045]&~m[2046]&~m[2070])|(~m[2043]&m[2044]&~m[2045]&~m[2046]&~m[2070])|(~m[2043]&~m[2044]&m[2045]&~m[2046]&~m[2070])|(m[2043]&m[2044]&~m[2045]&m[2046]&~m[2070])|(m[2043]&~m[2044]&m[2045]&m[2046]&~m[2070])|(~m[2043]&m[2044]&m[2045]&m[2046]&~m[2070]))&BiasedRNG[1118])|(((m[2043]&~m[2044]&~m[2045]&~m[2046]&m[2070])|(~m[2043]&m[2044]&~m[2045]&~m[2046]&m[2070])|(~m[2043]&~m[2044]&m[2045]&~m[2046]&m[2070])|(m[2043]&m[2044]&~m[2045]&m[2046]&m[2070])|(m[2043]&~m[2044]&m[2045]&m[2046]&m[2070])|(~m[2043]&m[2044]&m[2045]&m[2046]&m[2070]))&~BiasedRNG[1118])|((m[2043]&m[2044]&~m[2045]&~m[2046]&~m[2070])|(m[2043]&~m[2044]&m[2045]&~m[2046]&~m[2070])|(~m[2043]&m[2044]&m[2045]&~m[2046]&~m[2070])|(m[2043]&m[2044]&m[2045]&~m[2046]&~m[2070])|(m[2043]&m[2044]&m[2045]&m[2046]&~m[2070])|(m[2043]&m[2044]&~m[2045]&~m[2046]&m[2070])|(m[2043]&~m[2044]&m[2045]&~m[2046]&m[2070])|(~m[2043]&m[2044]&m[2045]&~m[2046]&m[2070])|(m[2043]&m[2044]&m[2045]&~m[2046]&m[2070])|(m[2043]&m[2044]&m[2045]&m[2046]&m[2070]))):InitCond[2064];
    m[2052] = run?((((m[2048]&~m[2049]&~m[2050]&~m[2051]&~m[2075])|(~m[2048]&m[2049]&~m[2050]&~m[2051]&~m[2075])|(~m[2048]&~m[2049]&m[2050]&~m[2051]&~m[2075])|(m[2048]&m[2049]&~m[2050]&m[2051]&~m[2075])|(m[2048]&~m[2049]&m[2050]&m[2051]&~m[2075])|(~m[2048]&m[2049]&m[2050]&m[2051]&~m[2075]))&BiasedRNG[1119])|(((m[2048]&~m[2049]&~m[2050]&~m[2051]&m[2075])|(~m[2048]&m[2049]&~m[2050]&~m[2051]&m[2075])|(~m[2048]&~m[2049]&m[2050]&~m[2051]&m[2075])|(m[2048]&m[2049]&~m[2050]&m[2051]&m[2075])|(m[2048]&~m[2049]&m[2050]&m[2051]&m[2075])|(~m[2048]&m[2049]&m[2050]&m[2051]&m[2075]))&~BiasedRNG[1119])|((m[2048]&m[2049]&~m[2050]&~m[2051]&~m[2075])|(m[2048]&~m[2049]&m[2050]&~m[2051]&~m[2075])|(~m[2048]&m[2049]&m[2050]&~m[2051]&~m[2075])|(m[2048]&m[2049]&m[2050]&~m[2051]&~m[2075])|(m[2048]&m[2049]&m[2050]&m[2051]&~m[2075])|(m[2048]&m[2049]&~m[2050]&~m[2051]&m[2075])|(m[2048]&~m[2049]&m[2050]&~m[2051]&m[2075])|(~m[2048]&m[2049]&m[2050]&~m[2051]&m[2075])|(m[2048]&m[2049]&m[2050]&~m[2051]&m[2075])|(m[2048]&m[2049]&m[2050]&m[2051]&m[2075]))):InitCond[2065];
    m[2057] = run?((((m[2053]&~m[2054]&~m[2055]&~m[2056]&~m[2078])|(~m[2053]&m[2054]&~m[2055]&~m[2056]&~m[2078])|(~m[2053]&~m[2054]&m[2055]&~m[2056]&~m[2078])|(m[2053]&m[2054]&~m[2055]&m[2056]&~m[2078])|(m[2053]&~m[2054]&m[2055]&m[2056]&~m[2078])|(~m[2053]&m[2054]&m[2055]&m[2056]&~m[2078]))&BiasedRNG[1120])|(((m[2053]&~m[2054]&~m[2055]&~m[2056]&m[2078])|(~m[2053]&m[2054]&~m[2055]&~m[2056]&m[2078])|(~m[2053]&~m[2054]&m[2055]&~m[2056]&m[2078])|(m[2053]&m[2054]&~m[2055]&m[2056]&m[2078])|(m[2053]&~m[2054]&m[2055]&m[2056]&m[2078])|(~m[2053]&m[2054]&m[2055]&m[2056]&m[2078]))&~BiasedRNG[1120])|((m[2053]&m[2054]&~m[2055]&~m[2056]&~m[2078])|(m[2053]&~m[2054]&m[2055]&~m[2056]&~m[2078])|(~m[2053]&m[2054]&m[2055]&~m[2056]&~m[2078])|(m[2053]&m[2054]&m[2055]&~m[2056]&~m[2078])|(m[2053]&m[2054]&m[2055]&m[2056]&~m[2078])|(m[2053]&m[2054]&~m[2055]&~m[2056]&m[2078])|(m[2053]&~m[2054]&m[2055]&~m[2056]&m[2078])|(~m[2053]&m[2054]&m[2055]&~m[2056]&m[2078])|(m[2053]&m[2054]&m[2055]&~m[2056]&m[2078])|(m[2053]&m[2054]&m[2055]&m[2056]&m[2078]))):InitCond[2066];
    m[2062] = run?((((m[2058]&~m[2059]&~m[2060]&~m[2061]&~m[2080])|(~m[2058]&m[2059]&~m[2060]&~m[2061]&~m[2080])|(~m[2058]&~m[2059]&m[2060]&~m[2061]&~m[2080])|(m[2058]&m[2059]&~m[2060]&m[2061]&~m[2080])|(m[2058]&~m[2059]&m[2060]&m[2061]&~m[2080])|(~m[2058]&m[2059]&m[2060]&m[2061]&~m[2080]))&BiasedRNG[1121])|(((m[2058]&~m[2059]&~m[2060]&~m[2061]&m[2080])|(~m[2058]&m[2059]&~m[2060]&~m[2061]&m[2080])|(~m[2058]&~m[2059]&m[2060]&~m[2061]&m[2080])|(m[2058]&m[2059]&~m[2060]&m[2061]&m[2080])|(m[2058]&~m[2059]&m[2060]&m[2061]&m[2080])|(~m[2058]&m[2059]&m[2060]&m[2061]&m[2080]))&~BiasedRNG[1121])|((m[2058]&m[2059]&~m[2060]&~m[2061]&~m[2080])|(m[2058]&~m[2059]&m[2060]&~m[2061]&~m[2080])|(~m[2058]&m[2059]&m[2060]&~m[2061]&~m[2080])|(m[2058]&m[2059]&m[2060]&~m[2061]&~m[2080])|(m[2058]&m[2059]&m[2060]&m[2061]&~m[2080])|(m[2058]&m[2059]&~m[2060]&~m[2061]&m[2080])|(m[2058]&~m[2059]&m[2060]&~m[2061]&m[2080])|(~m[2058]&m[2059]&m[2060]&~m[2061]&m[2080])|(m[2058]&m[2059]&m[2060]&~m[2061]&m[2080])|(m[2058]&m[2059]&m[2060]&m[2061]&m[2080]))):InitCond[2067];
    m[2067] = run?((((m[2063]&~m[2064]&~m[2065]&~m[2066]&~m[2085])|(~m[2063]&m[2064]&~m[2065]&~m[2066]&~m[2085])|(~m[2063]&~m[2064]&m[2065]&~m[2066]&~m[2085])|(m[2063]&m[2064]&~m[2065]&m[2066]&~m[2085])|(m[2063]&~m[2064]&m[2065]&m[2066]&~m[2085])|(~m[2063]&m[2064]&m[2065]&m[2066]&~m[2085]))&BiasedRNG[1122])|(((m[2063]&~m[2064]&~m[2065]&~m[2066]&m[2085])|(~m[2063]&m[2064]&~m[2065]&~m[2066]&m[2085])|(~m[2063]&~m[2064]&m[2065]&~m[2066]&m[2085])|(m[2063]&m[2064]&~m[2065]&m[2066]&m[2085])|(m[2063]&~m[2064]&m[2065]&m[2066]&m[2085])|(~m[2063]&m[2064]&m[2065]&m[2066]&m[2085]))&~BiasedRNG[1122])|((m[2063]&m[2064]&~m[2065]&~m[2066]&~m[2085])|(m[2063]&~m[2064]&m[2065]&~m[2066]&~m[2085])|(~m[2063]&m[2064]&m[2065]&~m[2066]&~m[2085])|(m[2063]&m[2064]&m[2065]&~m[2066]&~m[2085])|(m[2063]&m[2064]&m[2065]&m[2066]&~m[2085])|(m[2063]&m[2064]&~m[2065]&~m[2066]&m[2085])|(m[2063]&~m[2064]&m[2065]&~m[2066]&m[2085])|(~m[2063]&m[2064]&m[2065]&~m[2066]&m[2085])|(m[2063]&m[2064]&m[2065]&~m[2066]&m[2085])|(m[2063]&m[2064]&m[2065]&m[2066]&m[2085]))):InitCond[2068];
    m[2072] = run?((((m[2068]&~m[2069]&~m[2070]&~m[2071]&~m[2090])|(~m[2068]&m[2069]&~m[2070]&~m[2071]&~m[2090])|(~m[2068]&~m[2069]&m[2070]&~m[2071]&~m[2090])|(m[2068]&m[2069]&~m[2070]&m[2071]&~m[2090])|(m[2068]&~m[2069]&m[2070]&m[2071]&~m[2090])|(~m[2068]&m[2069]&m[2070]&m[2071]&~m[2090]))&BiasedRNG[1123])|(((m[2068]&~m[2069]&~m[2070]&~m[2071]&m[2090])|(~m[2068]&m[2069]&~m[2070]&~m[2071]&m[2090])|(~m[2068]&~m[2069]&m[2070]&~m[2071]&m[2090])|(m[2068]&m[2069]&~m[2070]&m[2071]&m[2090])|(m[2068]&~m[2069]&m[2070]&m[2071]&m[2090])|(~m[2068]&m[2069]&m[2070]&m[2071]&m[2090]))&~BiasedRNG[1123])|((m[2068]&m[2069]&~m[2070]&~m[2071]&~m[2090])|(m[2068]&~m[2069]&m[2070]&~m[2071]&~m[2090])|(~m[2068]&m[2069]&m[2070]&~m[2071]&~m[2090])|(m[2068]&m[2069]&m[2070]&~m[2071]&~m[2090])|(m[2068]&m[2069]&m[2070]&m[2071]&~m[2090])|(m[2068]&m[2069]&~m[2070]&~m[2071]&m[2090])|(m[2068]&~m[2069]&m[2070]&~m[2071]&m[2090])|(~m[2068]&m[2069]&m[2070]&~m[2071]&m[2090])|(m[2068]&m[2069]&m[2070]&~m[2071]&m[2090])|(m[2068]&m[2069]&m[2070]&m[2071]&m[2090]))):InitCond[2069];
    m[2077] = run?((((m[2073]&~m[2074]&~m[2075]&~m[2076]&~m[2095])|(~m[2073]&m[2074]&~m[2075]&~m[2076]&~m[2095])|(~m[2073]&~m[2074]&m[2075]&~m[2076]&~m[2095])|(m[2073]&m[2074]&~m[2075]&m[2076]&~m[2095])|(m[2073]&~m[2074]&m[2075]&m[2076]&~m[2095])|(~m[2073]&m[2074]&m[2075]&m[2076]&~m[2095]))&BiasedRNG[1124])|(((m[2073]&~m[2074]&~m[2075]&~m[2076]&m[2095])|(~m[2073]&m[2074]&~m[2075]&~m[2076]&m[2095])|(~m[2073]&~m[2074]&m[2075]&~m[2076]&m[2095])|(m[2073]&m[2074]&~m[2075]&m[2076]&m[2095])|(m[2073]&~m[2074]&m[2075]&m[2076]&m[2095])|(~m[2073]&m[2074]&m[2075]&m[2076]&m[2095]))&~BiasedRNG[1124])|((m[2073]&m[2074]&~m[2075]&~m[2076]&~m[2095])|(m[2073]&~m[2074]&m[2075]&~m[2076]&~m[2095])|(~m[2073]&m[2074]&m[2075]&~m[2076]&~m[2095])|(m[2073]&m[2074]&m[2075]&~m[2076]&~m[2095])|(m[2073]&m[2074]&m[2075]&m[2076]&~m[2095])|(m[2073]&m[2074]&~m[2075]&~m[2076]&m[2095])|(m[2073]&~m[2074]&m[2075]&~m[2076]&m[2095])|(~m[2073]&m[2074]&m[2075]&~m[2076]&m[2095])|(m[2073]&m[2074]&m[2075]&~m[2076]&m[2095])|(m[2073]&m[2074]&m[2075]&m[2076]&m[2095]))):InitCond[2070];
    m[2082] = run?((((m[2078]&~m[2079]&~m[2080]&~m[2081]&~m[2098])|(~m[2078]&m[2079]&~m[2080]&~m[2081]&~m[2098])|(~m[2078]&~m[2079]&m[2080]&~m[2081]&~m[2098])|(m[2078]&m[2079]&~m[2080]&m[2081]&~m[2098])|(m[2078]&~m[2079]&m[2080]&m[2081]&~m[2098])|(~m[2078]&m[2079]&m[2080]&m[2081]&~m[2098]))&BiasedRNG[1125])|(((m[2078]&~m[2079]&~m[2080]&~m[2081]&m[2098])|(~m[2078]&m[2079]&~m[2080]&~m[2081]&m[2098])|(~m[2078]&~m[2079]&m[2080]&~m[2081]&m[2098])|(m[2078]&m[2079]&~m[2080]&m[2081]&m[2098])|(m[2078]&~m[2079]&m[2080]&m[2081]&m[2098])|(~m[2078]&m[2079]&m[2080]&m[2081]&m[2098]))&~BiasedRNG[1125])|((m[2078]&m[2079]&~m[2080]&~m[2081]&~m[2098])|(m[2078]&~m[2079]&m[2080]&~m[2081]&~m[2098])|(~m[2078]&m[2079]&m[2080]&~m[2081]&~m[2098])|(m[2078]&m[2079]&m[2080]&~m[2081]&~m[2098])|(m[2078]&m[2079]&m[2080]&m[2081]&~m[2098])|(m[2078]&m[2079]&~m[2080]&~m[2081]&m[2098])|(m[2078]&~m[2079]&m[2080]&~m[2081]&m[2098])|(~m[2078]&m[2079]&m[2080]&~m[2081]&m[2098])|(m[2078]&m[2079]&m[2080]&~m[2081]&m[2098])|(m[2078]&m[2079]&m[2080]&m[2081]&m[2098]))):InitCond[2071];
    m[2087] = run?((((m[2083]&~m[2084]&~m[2085]&~m[2086]&~m[2100])|(~m[2083]&m[2084]&~m[2085]&~m[2086]&~m[2100])|(~m[2083]&~m[2084]&m[2085]&~m[2086]&~m[2100])|(m[2083]&m[2084]&~m[2085]&m[2086]&~m[2100])|(m[2083]&~m[2084]&m[2085]&m[2086]&~m[2100])|(~m[2083]&m[2084]&m[2085]&m[2086]&~m[2100]))&BiasedRNG[1126])|(((m[2083]&~m[2084]&~m[2085]&~m[2086]&m[2100])|(~m[2083]&m[2084]&~m[2085]&~m[2086]&m[2100])|(~m[2083]&~m[2084]&m[2085]&~m[2086]&m[2100])|(m[2083]&m[2084]&~m[2085]&m[2086]&m[2100])|(m[2083]&~m[2084]&m[2085]&m[2086]&m[2100])|(~m[2083]&m[2084]&m[2085]&m[2086]&m[2100]))&~BiasedRNG[1126])|((m[2083]&m[2084]&~m[2085]&~m[2086]&~m[2100])|(m[2083]&~m[2084]&m[2085]&~m[2086]&~m[2100])|(~m[2083]&m[2084]&m[2085]&~m[2086]&~m[2100])|(m[2083]&m[2084]&m[2085]&~m[2086]&~m[2100])|(m[2083]&m[2084]&m[2085]&m[2086]&~m[2100])|(m[2083]&m[2084]&~m[2085]&~m[2086]&m[2100])|(m[2083]&~m[2084]&m[2085]&~m[2086]&m[2100])|(~m[2083]&m[2084]&m[2085]&~m[2086]&m[2100])|(m[2083]&m[2084]&m[2085]&~m[2086]&m[2100])|(m[2083]&m[2084]&m[2085]&m[2086]&m[2100]))):InitCond[2072];
    m[2092] = run?((((m[2088]&~m[2089]&~m[2090]&~m[2091]&~m[2105])|(~m[2088]&m[2089]&~m[2090]&~m[2091]&~m[2105])|(~m[2088]&~m[2089]&m[2090]&~m[2091]&~m[2105])|(m[2088]&m[2089]&~m[2090]&m[2091]&~m[2105])|(m[2088]&~m[2089]&m[2090]&m[2091]&~m[2105])|(~m[2088]&m[2089]&m[2090]&m[2091]&~m[2105]))&BiasedRNG[1127])|(((m[2088]&~m[2089]&~m[2090]&~m[2091]&m[2105])|(~m[2088]&m[2089]&~m[2090]&~m[2091]&m[2105])|(~m[2088]&~m[2089]&m[2090]&~m[2091]&m[2105])|(m[2088]&m[2089]&~m[2090]&m[2091]&m[2105])|(m[2088]&~m[2089]&m[2090]&m[2091]&m[2105])|(~m[2088]&m[2089]&m[2090]&m[2091]&m[2105]))&~BiasedRNG[1127])|((m[2088]&m[2089]&~m[2090]&~m[2091]&~m[2105])|(m[2088]&~m[2089]&m[2090]&~m[2091]&~m[2105])|(~m[2088]&m[2089]&m[2090]&~m[2091]&~m[2105])|(m[2088]&m[2089]&m[2090]&~m[2091]&~m[2105])|(m[2088]&m[2089]&m[2090]&m[2091]&~m[2105])|(m[2088]&m[2089]&~m[2090]&~m[2091]&m[2105])|(m[2088]&~m[2089]&m[2090]&~m[2091]&m[2105])|(~m[2088]&m[2089]&m[2090]&~m[2091]&m[2105])|(m[2088]&m[2089]&m[2090]&~m[2091]&m[2105])|(m[2088]&m[2089]&m[2090]&m[2091]&m[2105]))):InitCond[2073];
    m[2097] = run?((((m[2093]&~m[2094]&~m[2095]&~m[2096]&~m[2110])|(~m[2093]&m[2094]&~m[2095]&~m[2096]&~m[2110])|(~m[2093]&~m[2094]&m[2095]&~m[2096]&~m[2110])|(m[2093]&m[2094]&~m[2095]&m[2096]&~m[2110])|(m[2093]&~m[2094]&m[2095]&m[2096]&~m[2110])|(~m[2093]&m[2094]&m[2095]&m[2096]&~m[2110]))&BiasedRNG[1128])|(((m[2093]&~m[2094]&~m[2095]&~m[2096]&m[2110])|(~m[2093]&m[2094]&~m[2095]&~m[2096]&m[2110])|(~m[2093]&~m[2094]&m[2095]&~m[2096]&m[2110])|(m[2093]&m[2094]&~m[2095]&m[2096]&m[2110])|(m[2093]&~m[2094]&m[2095]&m[2096]&m[2110])|(~m[2093]&m[2094]&m[2095]&m[2096]&m[2110]))&~BiasedRNG[1128])|((m[2093]&m[2094]&~m[2095]&~m[2096]&~m[2110])|(m[2093]&~m[2094]&m[2095]&~m[2096]&~m[2110])|(~m[2093]&m[2094]&m[2095]&~m[2096]&~m[2110])|(m[2093]&m[2094]&m[2095]&~m[2096]&~m[2110])|(m[2093]&m[2094]&m[2095]&m[2096]&~m[2110])|(m[2093]&m[2094]&~m[2095]&~m[2096]&m[2110])|(m[2093]&~m[2094]&m[2095]&~m[2096]&m[2110])|(~m[2093]&m[2094]&m[2095]&~m[2096]&m[2110])|(m[2093]&m[2094]&m[2095]&~m[2096]&m[2110])|(m[2093]&m[2094]&m[2095]&m[2096]&m[2110]))):InitCond[2074];
    m[2102] = run?((((m[2098]&~m[2099]&~m[2100]&~m[2101]&~m[2113])|(~m[2098]&m[2099]&~m[2100]&~m[2101]&~m[2113])|(~m[2098]&~m[2099]&m[2100]&~m[2101]&~m[2113])|(m[2098]&m[2099]&~m[2100]&m[2101]&~m[2113])|(m[2098]&~m[2099]&m[2100]&m[2101]&~m[2113])|(~m[2098]&m[2099]&m[2100]&m[2101]&~m[2113]))&BiasedRNG[1129])|(((m[2098]&~m[2099]&~m[2100]&~m[2101]&m[2113])|(~m[2098]&m[2099]&~m[2100]&~m[2101]&m[2113])|(~m[2098]&~m[2099]&m[2100]&~m[2101]&m[2113])|(m[2098]&m[2099]&~m[2100]&m[2101]&m[2113])|(m[2098]&~m[2099]&m[2100]&m[2101]&m[2113])|(~m[2098]&m[2099]&m[2100]&m[2101]&m[2113]))&~BiasedRNG[1129])|((m[2098]&m[2099]&~m[2100]&~m[2101]&~m[2113])|(m[2098]&~m[2099]&m[2100]&~m[2101]&~m[2113])|(~m[2098]&m[2099]&m[2100]&~m[2101]&~m[2113])|(m[2098]&m[2099]&m[2100]&~m[2101]&~m[2113])|(m[2098]&m[2099]&m[2100]&m[2101]&~m[2113])|(m[2098]&m[2099]&~m[2100]&~m[2101]&m[2113])|(m[2098]&~m[2099]&m[2100]&~m[2101]&m[2113])|(~m[2098]&m[2099]&m[2100]&~m[2101]&m[2113])|(m[2098]&m[2099]&m[2100]&~m[2101]&m[2113])|(m[2098]&m[2099]&m[2100]&m[2101]&m[2113]))):InitCond[2075];
    m[2107] = run?((((m[2103]&~m[2104]&~m[2105]&~m[2106]&~m[2115])|(~m[2103]&m[2104]&~m[2105]&~m[2106]&~m[2115])|(~m[2103]&~m[2104]&m[2105]&~m[2106]&~m[2115])|(m[2103]&m[2104]&~m[2105]&m[2106]&~m[2115])|(m[2103]&~m[2104]&m[2105]&m[2106]&~m[2115])|(~m[2103]&m[2104]&m[2105]&m[2106]&~m[2115]))&BiasedRNG[1130])|(((m[2103]&~m[2104]&~m[2105]&~m[2106]&m[2115])|(~m[2103]&m[2104]&~m[2105]&~m[2106]&m[2115])|(~m[2103]&~m[2104]&m[2105]&~m[2106]&m[2115])|(m[2103]&m[2104]&~m[2105]&m[2106]&m[2115])|(m[2103]&~m[2104]&m[2105]&m[2106]&m[2115])|(~m[2103]&m[2104]&m[2105]&m[2106]&m[2115]))&~BiasedRNG[1130])|((m[2103]&m[2104]&~m[2105]&~m[2106]&~m[2115])|(m[2103]&~m[2104]&m[2105]&~m[2106]&~m[2115])|(~m[2103]&m[2104]&m[2105]&~m[2106]&~m[2115])|(m[2103]&m[2104]&m[2105]&~m[2106]&~m[2115])|(m[2103]&m[2104]&m[2105]&m[2106]&~m[2115])|(m[2103]&m[2104]&~m[2105]&~m[2106]&m[2115])|(m[2103]&~m[2104]&m[2105]&~m[2106]&m[2115])|(~m[2103]&m[2104]&m[2105]&~m[2106]&m[2115])|(m[2103]&m[2104]&m[2105]&~m[2106]&m[2115])|(m[2103]&m[2104]&m[2105]&m[2106]&m[2115]))):InitCond[2076];
    m[2112] = run?((((m[2108]&~m[2109]&~m[2110]&~m[2111]&~m[2120])|(~m[2108]&m[2109]&~m[2110]&~m[2111]&~m[2120])|(~m[2108]&~m[2109]&m[2110]&~m[2111]&~m[2120])|(m[2108]&m[2109]&~m[2110]&m[2111]&~m[2120])|(m[2108]&~m[2109]&m[2110]&m[2111]&~m[2120])|(~m[2108]&m[2109]&m[2110]&m[2111]&~m[2120]))&BiasedRNG[1131])|(((m[2108]&~m[2109]&~m[2110]&~m[2111]&m[2120])|(~m[2108]&m[2109]&~m[2110]&~m[2111]&m[2120])|(~m[2108]&~m[2109]&m[2110]&~m[2111]&m[2120])|(m[2108]&m[2109]&~m[2110]&m[2111]&m[2120])|(m[2108]&~m[2109]&m[2110]&m[2111]&m[2120])|(~m[2108]&m[2109]&m[2110]&m[2111]&m[2120]))&~BiasedRNG[1131])|((m[2108]&m[2109]&~m[2110]&~m[2111]&~m[2120])|(m[2108]&~m[2109]&m[2110]&~m[2111]&~m[2120])|(~m[2108]&m[2109]&m[2110]&~m[2111]&~m[2120])|(m[2108]&m[2109]&m[2110]&~m[2111]&~m[2120])|(m[2108]&m[2109]&m[2110]&m[2111]&~m[2120])|(m[2108]&m[2109]&~m[2110]&~m[2111]&m[2120])|(m[2108]&~m[2109]&m[2110]&~m[2111]&m[2120])|(~m[2108]&m[2109]&m[2110]&~m[2111]&m[2120])|(m[2108]&m[2109]&m[2110]&~m[2111]&m[2120])|(m[2108]&m[2109]&m[2110]&m[2111]&m[2120]))):InitCond[2077];
    m[2117] = run?((((m[2113]&~m[2114]&~m[2115]&~m[2116]&~m[2123])|(~m[2113]&m[2114]&~m[2115]&~m[2116]&~m[2123])|(~m[2113]&~m[2114]&m[2115]&~m[2116]&~m[2123])|(m[2113]&m[2114]&~m[2115]&m[2116]&~m[2123])|(m[2113]&~m[2114]&m[2115]&m[2116]&~m[2123])|(~m[2113]&m[2114]&m[2115]&m[2116]&~m[2123]))&BiasedRNG[1132])|(((m[2113]&~m[2114]&~m[2115]&~m[2116]&m[2123])|(~m[2113]&m[2114]&~m[2115]&~m[2116]&m[2123])|(~m[2113]&~m[2114]&m[2115]&~m[2116]&m[2123])|(m[2113]&m[2114]&~m[2115]&m[2116]&m[2123])|(m[2113]&~m[2114]&m[2115]&m[2116]&m[2123])|(~m[2113]&m[2114]&m[2115]&m[2116]&m[2123]))&~BiasedRNG[1132])|((m[2113]&m[2114]&~m[2115]&~m[2116]&~m[2123])|(m[2113]&~m[2114]&m[2115]&~m[2116]&~m[2123])|(~m[2113]&m[2114]&m[2115]&~m[2116]&~m[2123])|(m[2113]&m[2114]&m[2115]&~m[2116]&~m[2123])|(m[2113]&m[2114]&m[2115]&m[2116]&~m[2123])|(m[2113]&m[2114]&~m[2115]&~m[2116]&m[2123])|(m[2113]&~m[2114]&m[2115]&~m[2116]&m[2123])|(~m[2113]&m[2114]&m[2115]&~m[2116]&m[2123])|(m[2113]&m[2114]&m[2115]&~m[2116]&m[2123])|(m[2113]&m[2114]&m[2115]&m[2116]&m[2123]))):InitCond[2078];
    m[2122] = run?((((m[2118]&~m[2119]&~m[2120]&~m[2121]&~m[2125])|(~m[2118]&m[2119]&~m[2120]&~m[2121]&~m[2125])|(~m[2118]&~m[2119]&m[2120]&~m[2121]&~m[2125])|(m[2118]&m[2119]&~m[2120]&m[2121]&~m[2125])|(m[2118]&~m[2119]&m[2120]&m[2121]&~m[2125])|(~m[2118]&m[2119]&m[2120]&m[2121]&~m[2125]))&BiasedRNG[1133])|(((m[2118]&~m[2119]&~m[2120]&~m[2121]&m[2125])|(~m[2118]&m[2119]&~m[2120]&~m[2121]&m[2125])|(~m[2118]&~m[2119]&m[2120]&~m[2121]&m[2125])|(m[2118]&m[2119]&~m[2120]&m[2121]&m[2125])|(m[2118]&~m[2119]&m[2120]&m[2121]&m[2125])|(~m[2118]&m[2119]&m[2120]&m[2121]&m[2125]))&~BiasedRNG[1133])|((m[2118]&m[2119]&~m[2120]&~m[2121]&~m[2125])|(m[2118]&~m[2119]&m[2120]&~m[2121]&~m[2125])|(~m[2118]&m[2119]&m[2120]&~m[2121]&~m[2125])|(m[2118]&m[2119]&m[2120]&~m[2121]&~m[2125])|(m[2118]&m[2119]&m[2120]&m[2121]&~m[2125])|(m[2118]&m[2119]&~m[2120]&~m[2121]&m[2125])|(m[2118]&~m[2119]&m[2120]&~m[2121]&m[2125])|(~m[2118]&m[2119]&m[2120]&~m[2121]&m[2125])|(m[2118]&m[2119]&m[2120]&~m[2121]&m[2125])|(m[2118]&m[2119]&m[2120]&m[2121]&m[2125]))):InitCond[2079];
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[1312]&LFSRcolor0[817]&LFSRcolor0[884]&LFSRcolor0[555]);
    BiasedRNG[1] = (LFSRcolor0[1094]&LFSRcolor0[146]&LFSRcolor0[1104]&LFSRcolor0[453]);
    BiasedRNG[2] = (LFSRcolor0[995]&LFSRcolor0[584]&LFSRcolor0[105]&LFSRcolor0[1168]);
    BiasedRNG[3] = (LFSRcolor0[971]&LFSRcolor0[353]&LFSRcolor0[990]&LFSRcolor0[688]);
    BiasedRNG[4] = (LFSRcolor0[102]&LFSRcolor0[934]&LFSRcolor0[790]&LFSRcolor0[897]);
    BiasedRNG[5] = (LFSRcolor0[1192]&LFSRcolor0[756]&LFSRcolor0[499]&LFSRcolor0[282]);
    BiasedRNG[6] = (LFSRcolor0[415]&LFSRcolor0[94]&LFSRcolor0[550]&LFSRcolor0[459]);
    BiasedRNG[7] = (LFSRcolor0[137]&LFSRcolor0[476]&LFSRcolor0[518]&LFSRcolor0[967]);
    BiasedRNG[8] = (LFSRcolor0[761]&LFSRcolor0[770]&LFSRcolor0[565]&LFSRcolor0[1193]);
    BiasedRNG[9] = (LFSRcolor0[948]&LFSRcolor0[525]&LFSRcolor0[197]&LFSRcolor0[607]);
    BiasedRNG[10] = (LFSRcolor0[95]&LFSRcolor0[408]&LFSRcolor0[717]&LFSRcolor0[332]);
    BiasedRNG[11] = (LFSRcolor0[177]&LFSRcolor0[952]&LFSRcolor0[987]&LFSRcolor0[778]);
    BiasedRNG[12] = (LFSRcolor0[41]&LFSRcolor0[920]&LFSRcolor0[936]&LFSRcolor0[113]);
    BiasedRNG[13] = (LFSRcolor0[1170]&LFSRcolor0[372]&LFSRcolor0[483]&LFSRcolor0[1133]);
    BiasedRNG[14] = (LFSRcolor0[25]&LFSRcolor0[479]&LFSRcolor0[201]&LFSRcolor0[1138]);
    BiasedRNG[15] = (LFSRcolor0[517]&LFSRcolor0[676]&LFSRcolor0[766]&LFSRcolor0[579]);
    BiasedRNG[16] = (LFSRcolor0[705]&LFSRcolor0[1061]&LFSRcolor0[190]&LFSRcolor0[1247]);
    BiasedRNG[17] = (LFSRcolor0[460]&LFSRcolor0[585]&LFSRcolor0[1290]&LFSRcolor0[1221]);
    BiasedRNG[18] = (LFSRcolor0[1049]&LFSRcolor0[1174]&LFSRcolor0[154]&LFSRcolor0[1008]);
    BiasedRNG[19] = (LFSRcolor0[194]&LFSRcolor0[17]&LFSRcolor0[998]&LFSRcolor0[1158]);
    BiasedRNG[20] = (LFSRcolor0[131]&LFSRcolor0[1275]&LFSRcolor0[1019]&LFSRcolor0[260]);
    BiasedRNG[21] = (LFSRcolor0[819]&LFSRcolor0[1035]&LFSRcolor0[1281]&LFSRcolor0[816]);
    BiasedRNG[22] = (LFSRcolor0[70]&LFSRcolor0[624]&LFSRcolor0[1197]&LFSRcolor0[242]);
    BiasedRNG[23] = (LFSRcolor0[93]&LFSRcolor0[88]&LFSRcolor0[600]&LFSRcolor0[123]);
    BiasedRNG[24] = (LFSRcolor0[931]&LFSRcolor0[1141]&LFSRcolor0[845]&LFSRcolor0[589]);
    BiasedRNG[25] = (LFSRcolor0[49]&LFSRcolor0[856]&LFSRcolor0[500]&LFSRcolor0[143]);
    BiasedRNG[26] = (LFSRcolor0[619]&LFSRcolor0[874]&LFSRcolor0[445]&LFSRcolor0[1128]);
    BiasedRNG[27] = (LFSRcolor0[1022]&LFSRcolor0[1236]&LFSRcolor0[329]&LFSRcolor0[323]);
    BiasedRNG[28] = (LFSRcolor0[250]&LFSRcolor0[150]&LFSRcolor0[366]&LFSRcolor0[905]);
    BiasedRNG[29] = (LFSRcolor0[863]&LFSRcolor0[1200]&LFSRcolor0[321]&LFSRcolor0[29]);
    BiasedRNG[30] = (LFSRcolor0[679]&LFSRcolor0[1320]&LFSRcolor0[792]&LFSRcolor0[84]);
    BiasedRNG[31] = (LFSRcolor0[208]&LFSRcolor0[338]&LFSRcolor0[660]&LFSRcolor0[846]);
    BiasedRNG[32] = (LFSRcolor0[294]&LFSRcolor0[765]&LFSRcolor0[0]&LFSRcolor0[340]);
    BiasedRNG[33] = (LFSRcolor0[295]&LFSRcolor0[433]&LFSRcolor0[657]&LFSRcolor0[1028]);
    BiasedRNG[34] = (LFSRcolor0[414]&LFSRcolor0[992]&LFSRcolor0[1187]&LFSRcolor0[754]);
    BiasedRNG[35] = (LFSRcolor0[215]&LFSRcolor0[156]&LFSRcolor0[1217]&LFSRcolor0[1242]);
    BiasedRNG[36] = (LFSRcolor0[159]&LFSRcolor0[1273]&LFSRcolor0[121]&LFSRcolor0[1212]);
    BiasedRNG[37] = (LFSRcolor0[1060]&LFSRcolor0[248]&LFSRcolor0[434]&LFSRcolor0[956]);
    BiasedRNG[38] = (LFSRcolor0[597]&LFSRcolor0[777]&LFSRcolor0[348]&LFSRcolor0[354]);
    BiasedRNG[39] = (LFSRcolor0[397]&LFSRcolor0[1089]&LFSRcolor0[165]&LFSRcolor0[596]);
    BiasedRNG[40] = (LFSRcolor0[975]&LFSRcolor0[1253]&LFSRcolor0[728]&LFSRcolor0[945]);
    BiasedRNG[41] = (LFSRcolor0[768]&LFSRcolor0[279]&LFSRcolor0[539]&LFSRcolor0[1189]);
    BiasedRNG[42] = (LFSRcolor0[245]&LFSRcolor0[652]&LFSRcolor0[1093]&LFSRcolor0[36]);
    BiasedRNG[43] = (LFSRcolor0[485]&LFSRcolor0[1153]&LFSRcolor0[877]&LFSRcolor0[663]);
    BiasedRNG[44] = (LFSRcolor0[955]&LFSRcolor0[511]&LFSRcolor0[1124]&LFSRcolor0[388]);
    BiasedRNG[45] = (LFSRcolor0[82]&LFSRcolor0[1159]&LFSRcolor0[136]&LFSRcolor0[832]);
    BiasedRNG[46] = (LFSRcolor0[502]&LFSRcolor0[664]&LFSRcolor0[733]&LFSRcolor0[200]);
    BiasedRNG[47] = (LFSRcolor0[708]&LFSRcolor0[148]&LFSRcolor0[1001]&LFSRcolor0[1092]);
    BiasedRNG[48] = (LFSRcolor0[457]&LFSRcolor0[1263]&LFSRcolor0[1127]&LFSRcolor0[801]);
    BiasedRNG[49] = (LFSRcolor0[814]&LFSRcolor0[784]&LFSRcolor0[595]&LFSRcolor0[75]);
    BiasedRNG[50] = (LFSRcolor0[382]&LFSRcolor0[526]&LFSRcolor0[166]&LFSRcolor0[394]);
    BiasedRNG[51] = (LFSRcolor0[763]&LFSRcolor0[196]&LFSRcolor0[737]&LFSRcolor0[883]);
    BiasedRNG[52] = (LFSRcolor0[358]&LFSRcolor0[1286]&LFSRcolor0[1121]&LFSRcolor0[1292]);
    BiasedRNG[53] = (LFSRcolor0[1239]&LFSRcolor0[224]&LFSRcolor0[376]&LFSRcolor0[642]);
    BiasedRNG[54] = (LFSRcolor0[773]&LFSRcolor0[537]&LFSRcolor0[1002]&LFSRcolor0[629]);
    BiasedRNG[55] = (LFSRcolor0[669]&LFSRcolor0[848]&LFSRcolor0[783]&LFSRcolor0[942]);
    BiasedRNG[56] = (LFSRcolor0[346]&LFSRcolor0[780]&LFSRcolor0[573]&LFSRcolor0[1143]);
    BiasedRNG[57] = (LFSRcolor0[843]&LFSRcolor0[741]&LFSRcolor0[1]&LFSRcolor0[370]);
    BiasedRNG[58] = (LFSRcolor0[1333]&LFSRcolor0[745]&LFSRcolor0[900]&LFSRcolor0[1037]);
    BiasedRNG[59] = (LFSRcolor0[1126]&LFSRcolor0[544]&LFSRcolor0[842]&LFSRcolor0[724]);
    BiasedRNG[60] = (LFSRcolor0[574]&LFSRcolor0[949]&LFSRcolor0[1216]&LFSRcolor0[730]);
    BiasedRNG[61] = (LFSRcolor0[450]&LFSRcolor0[130]&LFSRcolor0[899]&LFSRcolor0[230]);
    BiasedRNG[62] = (LFSRcolor0[1299]&LFSRcolor0[1006]&LFSRcolor0[379]&LFSRcolor0[1183]);
    BiasedRNG[63] = (LFSRcolor0[7]&LFSRcolor0[925]&LFSRcolor0[923]&LFSRcolor0[490]);
    BiasedRNG[64] = (LFSRcolor0[692]&LFSRcolor0[261]&LFSRcolor0[515]&LFSRcolor0[505]);
    BiasedRNG[65] = (LFSRcolor0[1070]&LFSRcolor0[641]&LFSRcolor0[61]&LFSRcolor0[1240]);
    BiasedRNG[66] = (LFSRcolor0[129]&LFSRcolor0[960]&LFSRcolor0[72]&LFSRcolor0[638]);
    BiasedRNG[67] = (LFSRcolor0[97]&LFSRcolor0[1155]&LFSRcolor0[1063]&LFSRcolor0[1079]);
    BiasedRNG[68] = (LFSRcolor0[1098]&LFSRcolor0[1171]&LFSRcolor0[1199]&LFSRcolor0[994]);
    BiasedRNG[69] = (LFSRcolor0[586]&LFSRcolor0[1026]&LFSRcolor0[1258]&LFSRcolor0[240]);
    BiasedRNG[70] = (LFSRcolor0[1140]&LFSRcolor0[873]&LFSRcolor0[513]&LFSRcolor0[540]);
    BiasedRNG[71] = (LFSRcolor0[1235]&LFSRcolor0[1250]&LFSRcolor0[1167]&LFSRcolor0[176]);
    BiasedRNG[72] = (LFSRcolor0[1271]&LFSRcolor0[714]&LFSRcolor0[1194]&LFSRcolor0[301]);
    BiasedRNG[73] = (LFSRcolor0[673]&LFSRcolor0[946]&LFSRcolor0[1027]&LFSRcolor0[860]);
    BiasedRNG[74] = (LFSRcolor0[55]&LFSRcolor0[1324]&LFSRcolor0[1261]&LFSRcolor0[1228]);
    BiasedRNG[75] = (LFSRcolor0[1066]&LFSRcolor0[1234]&LFSRcolor0[147]&LFSRcolor0[769]);
    BiasedRNG[76] = (LFSRcolor0[81]&LFSRcolor0[371]&LFSRcolor0[625]&LFSRcolor0[569]);
    BiasedRNG[77] = (LFSRcolor0[443]&LFSRcolor0[1000]&LFSRcolor0[1316]&LFSRcolor0[1114]);
    BiasedRNG[78] = (LFSRcolor0[411]&LFSRcolor0[344]&LFSRcolor0[861]&LFSRcolor0[719]);
    BiasedRNG[79] = (LFSRcolor0[1005]&LFSRcolor0[1254]&LFSRcolor0[670]&LFSRcolor0[299]);
    BiasedRNG[80] = (LFSRcolor0[1314]&LFSRcolor0[480]&LFSRcolor0[913]&LFSRcolor0[825]);
    BiasedRNG[81] = (LFSRcolor0[690]&LFSRcolor0[1137]&LFSRcolor0[12]&LFSRcolor0[1057]);
    BiasedRNG[82] = (LFSRcolor0[1191]&LFSRcolor0[606]&LFSRcolor0[300]&LFSRcolor0[138]);
    BiasedRNG[83] = (LFSRcolor0[941]&LFSRcolor0[319]&LFSRcolor0[1132]&LFSRcolor0[864]);
    BiasedRNG[84] = (LFSRcolor0[599]&LFSRcolor0[1303]&LFSRcolor0[189]&LFSRcolor0[1190]);
    BiasedRNG[85] = (LFSRcolor0[922]&LFSRcolor0[986]&LFSRcolor0[594]&LFSRcolor0[616]);
    BiasedRNG[86] = (LFSRcolor0[895]&LFSRcolor0[976]&LFSRcolor0[465]&LFSRcolor0[988]);
    BiasedRNG[87] = (LFSRcolor0[222]&LFSRcolor0[824]&LFSRcolor0[646]&LFSRcolor0[424]);
    BiasedRNG[88] = (LFSRcolor0[109]&LFSRcolor0[1294]&LFSRcolor0[760]&LFSRcolor0[439]);
    BiasedRNG[89] = (LFSRcolor0[605]&LFSRcolor0[903]&LFSRcolor0[1210]&LFSRcolor0[545]);
    BiasedRNG[90] = (LFSRcolor0[1246]&LFSRcolor0[609]&LFSRcolor0[648]&LFSRcolor0[283]);
    BiasedRNG[91] = (LFSRcolor0[964]&LFSRcolor0[1306]&LFSRcolor0[1220]&LFSRcolor0[810]);
    BiasedRNG[92] = (LFSRcolor0[682]&LFSRcolor0[1195]&LFSRcolor0[336]&LFSRcolor0[375]);
    BiasedRNG[93] = (LFSRcolor0[644]&LFSRcolor0[892]&LFSRcolor0[51]&LFSRcolor0[806]);
    BiasedRNG[94] = (LFSRcolor0[116]&LFSRcolor0[1023]&LFSRcolor0[822]&LFSRcolor0[588]);
    BiasedRNG[95] = (LFSRcolor0[716]&LFSRcolor0[455]&LFSRcolor0[420]&LFSRcolor0[398]);
    BiasedRNG[96] = (LFSRcolor0[314]&LFSRcolor0[689]&LFSRcolor0[1052]&LFSRcolor0[772]);
    BiasedRNG[97] = (LFSRcolor0[1186]&LFSRcolor0[331]&LFSRcolor0[651]&LFSRcolor0[39]);
    BiasedRNG[98] = (LFSRcolor0[885]&LFSRcolor0[111]&LFSRcolor0[1219]&LFSRcolor0[878]);
    BiasedRNG[99] = (LFSRcolor0[1188]&LFSRcolor0[1321]&LFSRcolor0[441]&LFSRcolor0[229]);
    BiasedRNG[100] = (LFSRcolor0[590]&LFSRcolor0[277]&LFSRcolor0[970]&LFSRcolor0[151]);
    BiasedRNG[101] = (LFSRcolor0[1102]&LFSRcolor0[426]&LFSRcolor0[1178]&LFSRcolor0[27]);
    BiasedRNG[102] = (LFSRcolor0[127]&LFSRcolor0[775]&LFSRcolor0[254]&LFSRcolor0[118]);
    BiasedRNG[103] = (LFSRcolor0[78]&LFSRcolor0[125]&LFSRcolor0[738]&LFSRcolor0[418]);
    BiasedRNG[104] = (LFSRcolor0[495]&LFSRcolor0[1135]&LFSRcolor0[767]&LFSRcolor0[636]);
    BiasedRNG[105] = (LFSRcolor0[1149]&LFSRcolor0[407]&LFSRcolor0[867]&LFSRcolor0[328]);
    BiasedRNG[106] = (LFSRcolor0[1116]&LFSRcolor0[626]&LFSRcolor0[850]&LFSRcolor0[727]);
    BiasedRNG[107] = (LFSRcolor0[437]&LFSRcolor0[937]&LFSRcolor0[1122]&LFSRcolor0[467]);
    BiasedRNG[108] = (LFSRcolor0[725]&LFSRcolor0[306]&LFSRcolor0[1293]&LFSRcolor0[493]);
    BiasedRNG[109] = (LFSRcolor0[310]&LFSRcolor0[364]&LFSRcolor0[278]&LFSRcolor0[195]);
    BiasedRNG[110] = (LFSRcolor0[1095]&LFSRcolor0[811]&LFSRcolor0[34]&LFSRcolor0[706]);
    BiasedRNG[111] = (LFSRcolor0[1179]&LFSRcolor0[1125]&LFSRcolor0[1308]&LFSRcolor0[1296]);
    BiasedRNG[112] = (LFSRcolor0[360]&LFSRcolor0[417]&LFSRcolor0[563]&LFSRcolor0[210]);
    BiasedRNG[113] = (LFSRcolor0[28]&LFSRcolor0[576]&LFSRcolor0[1145]&LFSRcolor0[172]);
    BiasedRNG[114] = (LFSRcolor0[225]&LFSRcolor0[915]&LFSRcolor0[337]&LFSRcolor0[813]);
    BiasedRNG[115] = (LFSRcolor0[735]&LFSRcolor0[1310]&LFSRcolor0[1329]&LFSRcolor0[841]);
    BiasedRNG[116] = (LFSRcolor0[838]&LFSRcolor0[898]&LFSRcolor0[630]&LFSRcolor0[536]);
    BiasedRNG[117] = (LFSRcolor0[577]&LFSRcolor0[1325]&LFSRcolor0[582]&LFSRcolor0[933]);
    BiasedRNG[118] = (LFSRcolor0[9]&LFSRcolor0[423]&LFSRcolor0[313]&LFSRcolor0[674]);
    BiasedRNG[119] = (LFSRcolor0[1184]&LFSRcolor0[1043]&LFSRcolor0[381]&LFSRcolor0[162]);
    BiasedRNG[120] = (LFSRcolor0[184]&LFSRcolor0[270]&LFSRcolor0[1161]&LFSRcolor0[972]);
    BiasedRNG[121] = (LFSRcolor0[788]&LFSRcolor0[1050]&LFSRcolor0[671]&LFSRcolor0[698]);
    BiasedRNG[122] = (LFSRcolor0[1185]&LFSRcolor0[155]&LFSRcolor0[1332]&LFSRcolor0[509]);
    BiasedRNG[123] = (LFSRcolor0[1058]&LFSRcolor0[100]&LFSRcolor0[870]&LFSRcolor0[1154]);
    BiasedRNG[124] = (LFSRcolor0[86]&LFSRcolor0[681]&LFSRcolor0[290]&LFSRcolor0[1091]);
    BiasedRNG[125] = (LFSRcolor0[157]&LFSRcolor0[1039]&LFSRcolor0[1289]&LFSRcolor0[474]);
    BiasedRNG[126] = (LFSRcolor0[206]&LFSRcolor0[977]&LFSRcolor0[1172]&LFSRcolor0[531]);
    BiasedRNG[127] = (LFSRcolor0[950]&LFSRcolor0[896]&LFSRcolor0[98]&LFSRcolor0[752]);
    BiasedRNG[128] = (LFSRcolor0[293]&LFSRcolor0[454]&LFSRcolor0[558]&LFSRcolor0[298]);
    BiasedRNG[129] = (LFSRcolor0[74]&LFSRcolor0[1209]&LFSRcolor0[377]&LFSRcolor0[1330]);
    BiasedRNG[130] = (LFSRcolor0[1107]&LFSRcolor0[880]&LFSRcolor0[68]&LFSRcolor0[982]);
    BiasedRNG[131] = (LFSRcolor0[209]&LFSRcolor0[117]&LFSRcolor0[1272]&LFSRcolor0[902]);
    BiasedRNG[132] = (LFSRcolor0[581]&LFSRcolor0[1208]&LFSRcolor0[753]&LFSRcolor0[567]);
    BiasedRNG[133] = (LFSRcolor0[732]&LFSRcolor0[48]&LFSRcolor0[268]&LFSRcolor0[410]);
    BiasedRNG[134] = (LFSRcolor0[330]&LFSRcolor0[851]&LFSRcolor0[687]&LFSRcolor0[830]);
    BiasedRNG[135] = (LFSRcolor0[887]&LFSRcolor0[1004]&LFSRcolor0[736]&LFSRcolor0[359]);
    BiasedRNG[136] = (LFSRcolor0[703]&LFSRcolor0[186]&LFSRcolor0[622]&LFSRcolor0[1232]);
    BiasedRNG[137] = (LFSRcolor0[959]&LFSRcolor0[436]&LFSRcolor0[1142]&LFSRcolor0[541]);
    BiasedRNG[138] = (LFSRcolor0[999]&LFSRcolor0[1120]&LFSRcolor0[1169]&LFSRcolor0[939]);
    BiasedRNG[139] = (LFSRcolor0[1072]&LFSRcolor0[1304]&LFSRcolor0[1031]&LFSRcolor0[809]);
    BiasedRNG[140] = (LFSRcolor0[869]&LFSRcolor0[747]&LFSRcolor0[1313]&LFSRcolor0[1003]);
    BiasedRNG[141] = (LFSRcolor0[702]&LFSRcolor0[362]&LFSRcolor0[965]&LFSRcolor0[428]);
    BiasedRNG[142] = (LFSRcolor0[2]&LFSRcolor0[711]&LFSRcolor0[1311]&LFSRcolor0[1211]);
    BiasedRNG[143] = (LFSRcolor0[315]&LFSRcolor0[935]&LFSRcolor0[8]&LFSRcolor0[1030]);
    BiasedRNG[144] = (LFSRcolor0[1139]&LFSRcolor0[365]&LFSRcolor0[1119]&LFSRcolor0[233]);
    BiasedRNG[145] = (LFSRcolor0[289]&LFSRcolor0[859]&LFSRcolor0[1032]&LFSRcolor0[559]);
    BiasedRNG[146] = (LFSRcolor0[794]&LFSRcolor0[991]&LFSRcolor0[1156]&LFSRcolor0[409]);
    BiasedRNG[147] = (LFSRcolor0[175]&LFSRcolor0[774]&LFSRcolor0[789]&LFSRcolor0[307]);
    BiasedRNG[148] = (LFSRcolor0[980]&LFSRcolor0[378]&LFSRcolor0[911]&LFSRcolor0[334]);
    BiasedRNG[149] = (LFSRcolor0[968]&LFSRcolor0[665]&LFSRcolor0[628]&LFSRcolor0[1229]);
    BiasedRNG[150] = (LFSRcolor0[5]&LFSRcolor0[89]&LFSRcolor0[60]&LFSRcolor0[1231]);
    BiasedRNG[151] = (LFSRcolor0[380]&LFSRcolor0[1280]&LFSRcolor0[471]&LFSRcolor0[546]);
    BiasedRNG[152] = (LFSRcolor0[1270]&LFSRcolor0[65]&LFSRcolor0[56]&LFSRcolor0[345]);
    BiasedRNG[153] = (LFSRcolor0[693]&LFSRcolor0[570]&LFSRcolor0[390]&LFSRcolor0[996]);
    BiasedRNG[154] = (LFSRcolor0[341]&LFSRcolor0[369]&LFSRcolor0[1260]&LFSRcolor0[361]);
    BiasedRNG[155] = (LFSRcolor0[83]&LFSRcolor0[342]&LFSRcolor0[530]&LFSRcolor0[239]);
    BiasedRNG[156] = (LFSRcolor0[335]&LFSRcolor0[1097]&LFSRcolor0[1157]&LFSRcolor0[1252]);
    BiasedRNG[157] = (LFSRcolor0[1078]&LFSRcolor0[385]&LFSRcolor0[291]&LFSRcolor0[1257]);
    BiasedRNG[158] = (LFSRcolor0[1251]&LFSRcolor0[153]&LFSRcolor0[272]&LFSRcolor0[984]);
    BiasedRNG[159] = (LFSRcolor0[221]&LFSRcolor0[472]&LFSRcolor0[661]&LFSRcolor0[1298]);
    BiasedRNG[160] = (LFSRcolor0[691]&LFSRcolor0[1196]&LFSRcolor0[758]&LFSRcolor0[14]);
    BiasedRNG[161] = (LFSRcolor0[1020]&LFSRcolor0[894]&LFSRcolor0[442]&LFSRcolor0[562]);
    BiasedRNG[162] = (LFSRcolor0[183]&LFSRcolor0[312]&LFSRcolor0[1068]&LFSRcolor0[80]);
    BiasedRNG[163] = (LFSRcolor0[1059]&LFSRcolor0[35]&LFSRcolor0[42]&LFSRcolor0[496]);
    BiasedRNG[164] = (LFSRcolor0[875]&LFSRcolor0[267]&LFSRcolor0[909]&LFSRcolor0[1284]);
    BiasedRNG[165] = (LFSRcolor0[820]&LFSRcolor0[1108]&LFSRcolor0[750]&LFSRcolor0[721]);
    BiasedRNG[166] = (LFSRcolor0[1248]&LFSRcolor0[553]&LFSRcolor0[797]&LFSRcolor0[1036]);
    BiasedRNG[167] = (LFSRcolor0[1160]&LFSRcolor0[1276]&LFSRcolor0[11]&LFSRcolor0[401]);
    BiasedRNG[168] = (LFSRcolor0[343]&LFSRcolor0[857]&LFSRcolor0[1326]&LFSRcolor0[486]);
    BiasedRNG[169] = (LFSRcolor0[1164]&LFSRcolor0[551]&LFSRcolor0[617]&LFSRcolor0[508]);
    BiasedRNG[170] = (LFSRcolor0[468]&LFSRcolor0[1123]&LFSRcolor0[168]&LFSRcolor0[557]);
    BiasedRNG[171] = (LFSRcolor0[449]&LFSRcolor0[640]&LFSRcolor0[1328]&LFSRcolor0[163]);
    BiasedRNG[172] = (LFSRcolor0[320]&LFSRcolor0[1082]&LFSRcolor0[649]&LFSRcolor0[548]);
    BiasedRNG[173] = (LFSRcolor0[566]&LFSRcolor0[680]&LFSRcolor0[1131]&LFSRcolor0[466]);
    BiasedRNG[174] = (LFSRcolor0[1064]&LFSRcolor0[771]&LFSRcolor0[107]&LFSRcolor0[1130]);
    BiasedRNG[175] = (LFSRcolor0[170]&LFSRcolor0[43]&LFSRcolor0[512]&LFSRcolor0[477]);
    BiasedRNG[176] = (LFSRcolor0[182]&LFSRcolor0[879]&LFSRcolor0[1025]&LFSRcolor0[203]);
    BiasedRNG[177] = (LFSRcolor0[1077]&LFSRcolor0[918]&LFSRcolor0[1051]&LFSRcolor0[1071]);
    BiasedRNG[178] = (LFSRcolor0[64]&LFSRcolor0[85]&LFSRcolor0[288]&LFSRcolor0[799]);
    BiasedRNG[179] = (LFSRcolor0[1282]&LFSRcolor0[1148]&LFSRcolor0[256]&LFSRcolor0[140]);
    BiasedRNG[180] = (LFSRcolor0[405]&LFSRcolor0[458]&LFSRcolor0[389]&LFSRcolor0[795]);
    BiasedRNG[181] = (LFSRcolor0[473]&LFSRcolor0[492]&LFSRcolor0[1083]&LFSRcolor0[1309]);
    BiasedRNG[182] = (LFSRcolor0[347]&LFSRcolor0[908]&LFSRcolor0[249]&LFSRcolor0[452]);
    BiasedRNG[183] = (LFSRcolor0[185]&LFSRcolor0[917]&LFSRcolor0[124]&LFSRcolor0[658]);
    BiasedRNG[184] = (LFSRcolor0[962]&LFSRcolor0[826]&LFSRcolor0[919]&LFSRcolor0[470]);
    BiasedRNG[185] = (LFSRcolor0[269]&LFSRcolor0[1021]&LFSRcolor0[818]&LFSRcolor0[700]);
    BiasedRNG[186] = (LFSRcolor0[858]&LFSRcolor0[79]&LFSRcolor0[710]&LFSRcolor0[621]);
    BiasedRNG[187] = (LFSRcolor0[759]&LFSRcolor0[601]&LFSRcolor0[906]&LFSRcolor0[1053]);
    BiasedRNG[188] = (LFSRcolor0[273]&LFSRcolor0[252]&LFSRcolor0[1065]&LFSRcolor0[808]);
    BiasedRNG[189] = (LFSRcolor0[1056]&LFSRcolor0[675]&LFSRcolor0[19]&LFSRcolor0[174]);
    BiasedRNG[190] = (LFSRcolor0[1241]&LFSRcolor0[253]&LFSRcolor0[391]&LFSRcolor0[464]);
    BiasedRNG[191] = (LFSRcolor0[1129]&LFSRcolor0[357]&LFSRcolor0[264]&LFSRcolor0[444]);
    BiasedRNG[192] = (LFSRcolor0[339]&LFSRcolor0[45]&LFSRcolor0[866]&LFSRcolor0[961]);
    BiasedRNG[193] = (LFSRcolor0[974]&LFSRcolor0[614]&LFSRcolor0[1177]&LFSRcolor0[1226]);
    BiasedRNG[194] = (LFSRcolor0[115]&LFSRcolor0[623]&LFSRcolor0[271]&LFSRcolor0[1233]);
    BiasedRNG[195] = (LFSRcolor0[187]&LFSRcolor0[938]&LFSRcolor0[779]&LFSRcolor0[33]);
    BiasedRNG[196] = (LFSRcolor0[198]&LFSRcolor0[787]&LFSRcolor0[1113]&LFSRcolor0[729]);
    BiasedRNG[197] = (LFSRcolor0[20]&LFSRcolor0[1225]&LFSRcolor0[891]&LFSRcolor0[528]);
    BiasedRNG[198] = (LFSRcolor0[287]&LFSRcolor0[1150]&LFSRcolor0[516]&LFSRcolor0[828]);
    BiasedRNG[199] = (LFSRcolor0[603]&LFSRcolor0[191]&LFSRcolor0[620]&LFSRcolor0[461]);
    BiasedRNG[200] = (LFSRcolor0[1096]&LFSRcolor0[355]&LFSRcolor0[23]&LFSRcolor0[363]);
    BiasedRNG[201] = (LFSRcolor0[1323]&LFSRcolor0[1046]&LFSRcolor0[1105]&LFSRcolor0[507]);
    BiasedRNG[202] = (LFSRcolor0[399]&LFSRcolor0[1012]&LFSRcolor0[549]&LFSRcolor0[1283]);
    BiasedRNG[203] = (LFSRcolor0[1266]&LFSRcolor0[1207]&LFSRcolor0[764]&LFSRcolor0[608]);
    BiasedRNG[204] = (LFSRcolor0[1227]&LFSRcolor0[104]&LFSRcolor0[234]&LFSRcolor0[114]);
    BiasedRNG[205] = (LFSRcolor0[52]&LFSRcolor0[90]&LFSRcolor0[92]&LFSRcolor0[501]);
    BiasedRNG[206] = (LFSRcolor0[1264]&LFSRcolor0[571]&LFSRcolor0[927]&LFSRcolor0[1014]);
    BiasedRNG[207] = (LFSRcolor0[1112]&LFSRcolor0[232]&LFSRcolor0[853]&LFSRcolor0[47]);
    BiasedRNG[208] = (LFSRcolor0[1045]&LFSRcolor0[69]&LFSRcolor0[1106]&LFSRcolor0[40]);
    BiasedRNG[209] = (LFSRcolor0[62]&LFSRcolor0[659]&LFSRcolor0[227]&LFSRcolor0[1165]);
    BiasedRNG[210] = (LFSRcolor0[743]&LFSRcolor0[1327]&LFSRcolor0[805]&LFSRcolor0[67]);
    BiasedRNG[211] = (LFSRcolor0[255]&LFSRcolor0[205]&LFSRcolor0[456]&LFSRcolor0[101]);
    BiasedRNG[212] = (LFSRcolor0[1218]&LFSRcolor0[1297]&LFSRcolor0[506]&LFSRcolor0[726]);
    BiasedRNG[213] = (LFSRcolor0[367]&LFSRcolor0[755]&LFSRcolor0[568]&LFSRcolor0[132]);
    BiasedRNG[214] = (LFSRcolor0[178]&LFSRcolor0[1080]&LFSRcolor0[776]&LFSRcolor0[1010]);
    BiasedRNG[215] = (LFSRcolor0[932]&LFSRcolor0[647]&LFSRcolor0[929]&LFSRcolor0[161]);
    BiasedRNG[216] = (LFSRcolor0[823]&LFSRcolor0[1146]&LFSRcolor0[807]&LFSRcolor0[793]);
    BiasedRNG[217] = (LFSRcolor0[547]&LFSRcolor0[1182]&LFSRcolor0[685]&LFSRcolor0[575]);
    BiasedRNG[218] = (LFSRcolor0[1322]&LFSRcolor0[488]&LFSRcolor0[108]&LFSRcolor0[1084]);
    BiasedRNG[219] = (LFSRcolor0[804]&LFSRcolor0[219]&LFSRcolor0[834]&LFSRcolor0[1267]);
    BiasedRNG[220] = (LFSRcolor0[169]&LFSRcolor0[697]&LFSRcolor0[901]&LFSRcolor0[214]);
    BiasedRNG[221] = (LFSRcolor0[653]&LFSRcolor0[1269]&LFSRcolor0[1110]&LFSRcolor0[266]);
    BiasedRNG[222] = (LFSRcolor0[749]&LFSRcolor0[538]&LFSRcolor0[1166]&LFSRcolor0[618]);
    BiasedRNG[223] = (LFSRcolor0[1085]&LFSRcolor0[997]&LFSRcolor0[1024]&LFSRcolor0[610]);
    BiasedRNG[224] = (LFSRcolor0[1249]&LFSRcolor0[871]&LFSRcolor0[4]&LFSRcolor0[1147]);
    BiasedRNG[225] = (LFSRcolor0[1244]&LFSRcolor0[134]&LFSRcolor0[973]&LFSRcolor0[734]);
    BiasedRNG[226] = (LFSRcolor0[1224]&LFSRcolor0[882]&LFSRcolor0[683]&LFSRcolor0[297]);
    BiasedRNG[227] = (LFSRcolor0[709]&LFSRcolor0[236]&LFSRcolor0[827]&LFSRcolor0[218]);
    BiasedRNG[228] = (LFSRcolor0[13]&LFSRcolor0[611]&LFSRcolor0[228]&LFSRcolor0[31]);
    BiasedRNG[229] = (LFSRcolor0[757]&LFSRcolor0[482]&LFSRcolor0[519]&LFSRcolor0[1118]);
    BiasedRNG[230] = (LFSRcolor0[333]&LFSRcolor0[149]&LFSRcolor0[662]&LFSRcolor0[383]);
    BiasedRNG[231] = (LFSRcolor0[1088]&LFSRcolor0[1291]&LFSRcolor0[462]&LFSRcolor0[835]);
    BiasedRNG[232] = (LFSRcolor0[316]&LFSRcolor0[139]&LFSRcolor0[1062]&LFSRcolor0[435]);
    BiasedRNG[233] = (LFSRcolor0[751]&LFSRcolor0[821]&LFSRcolor0[504]&LFSRcolor0[914]);
    BiasedRNG[234] = (LFSRcolor0[57]&LFSRcolor0[179]&LFSRcolor0[231]&LFSRcolor0[71]);
    BiasedRNG[235] = (LFSRcolor0[812]&LFSRcolor0[6]&LFSRcolor0[966]&LFSRcolor0[593]);
    BiasedRNG[236] = (LFSRcolor0[1301]&LFSRcolor0[650]&LFSRcolor0[26]&LFSRcolor0[746]);
    BiasedRNG[237] = (LFSRcolor0[978]&LFSRcolor0[484]&LFSRcolor0[1201]&LFSRcolor0[940]);
    BiasedRNG[238] = (LFSRcolor0[1331]&LFSRcolor0[930]&LFSRcolor0[1237]&LFSRcolor0[50]);
    BiasedRNG[239] = (LFSRcolor0[837]&LFSRcolor0[326]&LFSRcolor0[304]&LFSRcolor0[489]);
    BiasedRNG[240] = (LFSRcolor0[368]&LFSRcolor0[322]&LFSRcolor0[1245]&LFSRcolor0[235]);
    BiasedRNG[241] = (LFSRcolor0[989]&LFSRcolor0[16]&LFSRcolor0[46]&LFSRcolor0[943]);
    BiasedRNG[242] = (LFSRcolor0[286]&LFSRcolor0[969]&LFSRcolor0[1111]&LFSRcolor0[96]);
    BiasedRNG[243] = (LFSRcolor0[947]&LFSRcolor0[387]&LFSRcolor0[1205]&LFSRcolor0[678]);
    BiasedRNG[244] = (LFSRcolor0[246]&LFSRcolor0[928]&LFSRcolor0[422]&LFSRcolor0[440]);
    BiasedRNG[245] = (LFSRcolor0[193]&LFSRcolor0[303]&LFSRcolor0[1034]&LFSRcolor0[704]);
    BiasedRNG[246] = (LFSRcolor0[1214]&LFSRcolor0[855]&LFSRcolor0[637]&LFSRcolor0[167]);
    BiasedRNG[247] = (LFSRcolor0[32]&LFSRcolor0[144]&LFSRcolor0[317]&LFSRcolor0[522]);
    BiasedRNG[248] = (LFSRcolor0[572]&LFSRcolor0[723]&LFSRcolor0[633]&LFSRcolor0[276]);
    BiasedRNG[249] = (LFSRcolor0[192]&LFSRcolor0[592]&LFSRcolor0[829]&LFSRcolor0[634]);
    BiasedRNG[250] = (LFSRcolor0[904]&LFSRcolor0[1277]&LFSRcolor0[392]&LFSRcolor0[1075]);
    BiasedRNG[251] = (LFSRcolor0[416]&LFSRcolor0[655]&LFSRcolor0[1319]&LFSRcolor0[1100]);
    BiasedRNG[252] = (LFSRcolor0[400]&LFSRcolor0[889]&LFSRcolor0[1033]&LFSRcolor0[404]);
    BiasedRNG[253] = (LFSRcolor0[1076]&LFSRcolor0[510]&LFSRcolor0[839]&LFSRcolor0[106]);
    BiasedRNG[254] = (LFSRcolor0[325]&LFSRcolor0[1101]&LFSRcolor0[204]&LFSRcolor0[503]);
    BiasedRNG[255] = (LFSRcolor0[910]&LFSRcolor0[280]&LFSRcolor0[142]&LFSRcolor0[373]);
    UnbiasedRNG[0] = LFSRcolor0[907];
    UnbiasedRNG[1] = LFSRcolor0[1115];
    UnbiasedRNG[2] = LFSRcolor0[854];
    UnbiasedRNG[3] = LFSRcolor0[598];
    UnbiasedRNG[4] = LFSRcolor0[762];
    UnbiasedRNG[5] = LFSRcolor0[419];
    UnbiasedRNG[6] = LFSRcolor0[1203];
    UnbiasedRNG[7] = LFSRcolor0[430];
    UnbiasedRNG[8] = LFSRcolor0[311];
    UnbiasedRNG[9] = LFSRcolor0[1213];
    UnbiasedRNG[10] = LFSRcolor0[63];
    UnbiasedRNG[11] = LFSRcolor0[99];
    UnbiasedRNG[12] = LFSRcolor0[604];
    UnbiasedRNG[13] = LFSRcolor0[521];
    UnbiasedRNG[14] = LFSRcolor0[1007];
    UnbiasedRNG[15] = LFSRcolor0[552];
    UnbiasedRNG[16] = LFSRcolor0[207];
    UnbiasedRNG[17] = LFSRcolor0[446];
    UnbiasedRNG[18] = LFSRcolor0[349];
    UnbiasedRNG[19] = LFSRcolor0[448];
    UnbiasedRNG[20] = LFSRcolor0[1202];
    UnbiasedRNG[21] = LFSRcolor0[713];
    UnbiasedRNG[22] = LFSRcolor0[958];
    UnbiasedRNG[23] = LFSRcolor0[308];
    UnbiasedRNG[24] = LFSRcolor0[1230];
    UnbiasedRNG[25] = LFSRcolor0[535];
    UnbiasedRNG[26] = LFSRcolor0[715];
    UnbiasedRNG[27] = LFSRcolor0[145];
    UnbiasedRNG[28] = LFSRcolor0[785];
    UnbiasedRNG[29] = LFSRcolor0[529];
    UnbiasedRNG[30] = LFSRcolor0[791];
    UnbiasedRNG[31] = LFSRcolor0[1074];
    UnbiasedRNG[32] = LFSRcolor0[1016];
    UnbiasedRNG[33] = LFSRcolor0[37];
    UnbiasedRNG[34] = LFSRcolor0[265];
    UnbiasedRNG[35] = LFSRcolor0[1215];
    UnbiasedRNG[36] = LFSRcolor0[396];
    UnbiasedRNG[37] = LFSRcolor0[110];
    UnbiasedRNG[38] = LFSRcolor0[15];
    UnbiasedRNG[39] = LFSRcolor0[247];
    UnbiasedRNG[40] = LFSRcolor0[1318];
    UnbiasedRNG[41] = LFSRcolor0[872];
    UnbiasedRNG[42] = LFSRcolor0[1223];
    UnbiasedRNG[43] = LFSRcolor0[583];
    UnbiasedRNG[44] = LFSRcolor0[412];
    UnbiasedRNG[45] = LFSRcolor0[1259];
    UnbiasedRNG[46] = LFSRcolor0[916];
    UnbiasedRNG[47] = LFSRcolor0[523];
    UnbiasedRNG[48] = LFSRcolor0[119];
    UnbiasedRNG[49] = LFSRcolor0[742];
    UnbiasedRNG[50] = LFSRcolor0[251];
    UnbiasedRNG[51] = LFSRcolor0[1018];
    UnbiasedRNG[52] = LFSRcolor0[395];
    UnbiasedRNG[53] = LFSRcolor0[1086];
    UnbiasedRNG[54] = LFSRcolor0[798];
    UnbiasedRNG[55] = LFSRcolor0[954];
    UnbiasedRNG[56] = LFSRcolor0[656];
    UnbiasedRNG[57] = LFSRcolor0[425];
    UnbiasedRNG[58] = LFSRcolor0[1238];
    UnbiasedRNG[59] = LFSRcolor0[87];
    UnbiasedRNG[60] = LFSRcolor0[556];
    UnbiasedRNG[61] = LFSRcolor0[1144];
    UnbiasedRNG[62] = LFSRcolor0[38];
    UnbiasedRNG[63] = LFSRcolor0[285];
    UnbiasedRNG[64] = LFSRcolor0[212];
    UnbiasedRNG[65] = LFSRcolor0[30];
    UnbiasedRNG[66] = LFSRcolor0[1044];
    UnbiasedRNG[67] = LFSRcolor0[612];
    UnbiasedRNG[68] = LFSRcolor0[639];
    UnbiasedRNG[69] = LFSRcolor0[542];
    UnbiasedRNG[70] = LFSRcolor0[22];
    UnbiasedRNG[71] = LFSRcolor0[886];
    UnbiasedRNG[72] = LFSRcolor0[481];
    UnbiasedRNG[73] = LFSRcolor0[199];
    UnbiasedRNG[74] = LFSRcolor0[1262];
    UnbiasedRNG[75] = LFSRcolor0[351];
    UnbiasedRNG[76] = LFSRcolor0[386];
    UnbiasedRNG[77] = LFSRcolor0[578];
    UnbiasedRNG[78] = LFSRcolor0[21];
    UnbiasedRNG[79] = LFSRcolor0[91];
    UnbiasedRNG[80] = LFSRcolor0[1206];
    UnbiasedRNG[81] = LFSRcolor0[438];
    UnbiasedRNG[82] = LFSRcolor0[1222];
    UnbiasedRNG[83] = LFSRcolor0[1295];
    UnbiasedRNG[84] = LFSRcolor0[847];
    UnbiasedRNG[85] = LFSRcolor0[1285];
    UnbiasedRNG[86] = LFSRcolor0[1315];
    UnbiasedRNG[87] = LFSRcolor0[1279];
    UnbiasedRNG[88] = LFSRcolor0[327];
    UnbiasedRNG[89] = LFSRcolor0[296];
    UnbiasedRNG[90] = LFSRcolor0[1163];
    UnbiasedRNG[91] = LFSRcolor0[491];
    UnbiasedRNG[92] = LFSRcolor0[957];
    UnbiasedRNG[93] = LFSRcolor0[318];
    UnbiasedRNG[94] = LFSRcolor0[1274];
    UnbiasedRNG[95] = LFSRcolor0[171];
    UnbiasedRNG[96] = LFSRcolor0[1204];
    UnbiasedRNG[97] = LFSRcolor0[120];
    UnbiasedRNG[98] = LFSRcolor0[494];
    UnbiasedRNG[99] = LFSRcolor0[202];
    UnbiasedRNG[100] = LFSRcolor0[66];
    UnbiasedRNG[101] = LFSRcolor0[893];
    UnbiasedRNG[102] = LFSRcolor0[1243];
    UnbiasedRNG[103] = LFSRcolor0[217];
    UnbiasedRNG[104] = LFSRcolor0[1067];
    UnbiasedRNG[105] = LFSRcolor0[1152];
    UnbiasedRNG[106] = LFSRcolor0[921];
    UnbiasedRNG[107] = LFSRcolor0[554];
    UnbiasedRNG[108] = LFSRcolor0[1017];
    UnbiasedRNG[109] = LFSRcolor0[284];
    UnbiasedRNG[110] = LFSRcolor0[1307];
    UnbiasedRNG[111] = LFSRcolor0[1081];
    UnbiasedRNG[112] = LFSRcolor0[1011];
    UnbiasedRNG[113] = LFSRcolor0[1136];
    UnbiasedRNG[114] = LFSRcolor0[831];
    UnbiasedRNG[115] = LFSRcolor0[815];
    UnbiasedRNG[116] = LFSRcolor0[173];
    UnbiasedRNG[117] = LFSRcolor0[112];
    UnbiasedRNG[118] = LFSRcolor0[613];
    UnbiasedRNG[119] = LFSRcolor0[384];
    UnbiasedRNG[120] = LFSRcolor0[1173];
    UnbiasedRNG[121] = LFSRcolor0[258];
    UnbiasedRNG[122] = LFSRcolor0[865];
    UnbiasedRNG[123] = LFSRcolor0[10];
    UnbiasedRNG[124] = LFSRcolor0[76];
    UnbiasedRNG[125] = LFSRcolor0[356];
    UnbiasedRNG[126] = LFSRcolor0[686];
    UnbiasedRNG[127] = LFSRcolor0[77];
    UnbiasedRNG[128] = LFSRcolor0[985];
    UnbiasedRNG[129] = LFSRcolor0[1013];
    UnbiasedRNG[130] = LFSRcolor0[238];
    UnbiasedRNG[131] = LFSRcolor0[1288];
    UnbiasedRNG[132] = LFSRcolor0[836];
    UnbiasedRNG[133] = LFSRcolor0[53];
    UnbiasedRNG[134] = LFSRcolor0[677];
    UnbiasedRNG[135] = LFSRcolor0[667];
    UnbiasedRNG[136] = LFSRcolor0[631];
    UnbiasedRNG[137] = LFSRcolor0[262];
    UnbiasedRNG[138] = LFSRcolor0[292];
    UnbiasedRNG[139] = LFSRcolor0[1054];
    UnbiasedRNG[140] = LFSRcolor0[654];
    UnbiasedRNG[141] = LFSRcolor0[1117];
    UnbiasedRNG[142] = LFSRcolor0[722];
    UnbiasedRNG[143] = LFSRcolor0[406];
    UnbiasedRNG[144] = LFSRcolor0[431];
    UnbiasedRNG[145] = LFSRcolor0[220];
    UnbiasedRNG[146] = LFSRcolor0[24];
    UnbiasedRNG[147] = LFSRcolor0[469];
    UnbiasedRNG[148] = LFSRcolor0[862];
    UnbiasedRNG[149] = LFSRcolor0[263];
    UnbiasedRNG[150] = LFSRcolor0[696];
    UnbiasedRNG[151] = LFSRcolor0[243];
    UnbiasedRNG[152] = LFSRcolor0[59];
    UnbiasedRNG[153] = LFSRcolor0[699];
    UnbiasedRNG[154] = LFSRcolor0[564];
    UnbiasedRNG[155] = LFSRcolor0[740];
    UnbiasedRNG[156] = LFSRcolor0[447];
    UnbiasedRNG[157] = LFSRcolor0[1181];
    UnbiasedRNG[158] = LFSRcolor0[237];
    UnbiasedRNG[159] = LFSRcolor0[520];
    UnbiasedRNG[160] = LFSRcolor0[122];
    UnbiasedRNG[161] = LFSRcolor0[1134];
    UnbiasedRNG[162] = LFSRcolor0[852];
    UnbiasedRNG[163] = LFSRcolor0[152];
    UnbiasedRNG[164] = LFSRcolor0[731];
    UnbiasedRNG[165] = LFSRcolor0[514];
    UnbiasedRNG[166] = LFSRcolor0[707];
    UnbiasedRNG[167] = LFSRcolor0[560];
    UnbiasedRNG[168] = LFSRcolor0[800];
    UnbiasedRNG[169] = LFSRcolor0[712];
    UnbiasedRNG[170] = LFSRcolor0[213];
    UnbiasedRNG[171] = LFSRcolor0[1268];
    UnbiasedRNG[172] = LFSRcolor0[1255];
    UnbiasedRNG[173] = LFSRcolor0[158];
    UnbiasedRNG[174] = LFSRcolor0[403];
    UnbiasedRNG[175] = LFSRcolor0[802];
    UnbiasedRNG[176] = LFSRcolor0[188];
    UnbiasedRNG[177] = LFSRcolor0[627];
    UnbiasedRNG[178] = LFSRcolor0[128];
    UnbiasedRNG[179] = LFSRcolor0[54];
    UnbiasedRNG[180] = LFSRcolor0[890];
    UnbiasedRNG[181] = LFSRcolor0[944];
    UnbiasedRNG[182] = LFSRcolor0[635];
    UnbiasedRNG[183] = LFSRcolor0[402];
    UnbiasedRNG[184] = LFSRcolor0[1256];
    UnbiasedRNG[185] = LFSRcolor0[413];
    UnbiasedRNG[186] = LFSRcolor0[632];
    UnbiasedRNG[187] = LFSRcolor0[309];
    UnbiasedRNG[188] = LFSRcolor0[1038];
    UnbiasedRNG[189] = LFSRcolor0[1048];
    UnbiasedRNG[190] = LFSRcolor0[981];
    UnbiasedRNG[191] = LFSRcolor0[1109];
    UnbiasedRNG[192] = LFSRcolor0[350];
    UnbiasedRNG[193] = LFSRcolor0[543];
    UnbiasedRNG[194] = LFSRcolor0[781];
    UnbiasedRNG[195] = LFSRcolor0[1302];
    UnbiasedRNG[196] = LFSRcolor0[672];
    UnbiasedRNG[197] = LFSRcolor0[1087];
    UnbiasedRNG[198] = LFSRcolor0[963];
    UnbiasedRNG[199] = LFSRcolor0[888];
    UnbiasedRNG[200] = LFSRcolor0[739];
    UnbiasedRNG[201] = LFSRcolor0[881];
    UnbiasedRNG[202] = LFSRcolor0[302];
    UnbiasedRNG[203] = LFSRcolor0[744];
    UnbiasedRNG[204] = LFSRcolor0[701];
    UnbiasedRNG[205] = LFSRcolor0[979];
    UnbiasedRNG[206] = LFSRcolor0[1029];
    UnbiasedRNG[207] = LFSRcolor0[953];
    UnbiasedRNG[208] = LFSRcolor0[281];
    UnbiasedRNG[209] = LFSRcolor0[587];
    UnbiasedRNG[210] = LFSRcolor0[451];
    UnbiasedRNG[211] = LFSRcolor0[849];
    UnbiasedRNG[212] = LFSRcolor0[324];
    UnbiasedRNG[213] = LFSRcolor0[216];
    UnbiasedRNG[214] = LFSRcolor0[666];
    UnbiasedRNG[215] = LFSRcolor0[180];
    UnbiasedRNG[216] = LFSRcolor0[844];
    UnbiasedRNG[217] = LFSRcolor0[44];
    UnbiasedRNG[218] = LFSRcolor0[1278];
    UnbiasedRNG[219] = LFSRcolor0[374];
    UnbiasedRNG[220] = LFSRcolor0[58];
    UnbiasedRNG[221] = LFSRcolor0[244];
    UnbiasedRNG[222] = LFSRcolor0[1090];
    UnbiasedRNG[223] = LFSRcolor0[748];
    UnbiasedRNG[224] = LFSRcolor0[718];
    UnbiasedRNG[225] = LFSRcolor0[580];
    UnbiasedRNG[226] = LFSRcolor0[103];
    UnbiasedRNG[227] = LFSRcolor0[645];
    UnbiasedRNG[228] = LFSRcolor0[840];
    UnbiasedRNG[229] = LFSRcolor0[668];
    UnbiasedRNG[230] = LFSRcolor0[720];
    UnbiasedRNG[231] = LFSRcolor0[1175];
    UnbiasedRNG[232] = LFSRcolor0[796];
    UnbiasedRNG[233] = LFSRcolor0[912];
    UnbiasedRNG[234] = LFSRcolor0[1047];
    UnbiasedRNG[235] = LFSRcolor0[876];
    UnbiasedRNG[236] = LFSRcolor0[1176];
    UnbiasedRNG[237] = LFSRcolor0[1069];
    UnbiasedRNG[238] = LFSRcolor0[695];
    UnbiasedRNG[239] = LFSRcolor0[1151];
    UnbiasedRNG[240] = LFSRcolor0[427];
    UnbiasedRNG[241] = LFSRcolor0[164];
    UnbiasedRNG[242] = LFSRcolor0[786];
    UnbiasedRNG[243] = LFSRcolor0[259];
    UnbiasedRNG[244] = LFSRcolor0[1009];
    UnbiasedRNG[245] = LFSRcolor0[983];
    UnbiasedRNG[246] = LFSRcolor0[181];
    UnbiasedRNG[247] = LFSRcolor0[924];
    UnbiasedRNG[248] = LFSRcolor0[951];
    UnbiasedRNG[249] = LFSRcolor0[429];
    UnbiasedRNG[250] = LFSRcolor0[305];
    UnbiasedRNG[251] = LFSRcolor0[803];
    UnbiasedRNG[252] = LFSRcolor0[993];
    UnbiasedRNG[253] = LFSRcolor0[524];
    UnbiasedRNG[254] = LFSRcolor0[223];
    UnbiasedRNG[255] = LFSRcolor0[393];
    UnbiasedRNG[256] = LFSRcolor0[141];
    UnbiasedRNG[257] = LFSRcolor0[211];
    UnbiasedRNG[258] = LFSRcolor0[478];
    UnbiasedRNG[259] = LFSRcolor0[241];
    UnbiasedRNG[260] = LFSRcolor0[602];
    UnbiasedRNG[261] = LFSRcolor0[257];
    UnbiasedRNG[262] = LFSRcolor0[1198];
    UnbiasedRNG[263] = LFSRcolor0[533];
    UnbiasedRNG[264] = LFSRcolor0[487];
    UnbiasedRNG[265] = LFSRcolor0[274];
    UnbiasedRNG[266] = LFSRcolor0[126];
    UnbiasedRNG[267] = LFSRcolor0[1055];
    UnbiasedRNG[268] = LFSRcolor0[926];
    UnbiasedRNG[269] = LFSRcolor0[643];
    UnbiasedRNG[270] = LFSRcolor0[1317];
end

always @(posedge color0_clk) begin
    BiasedRNG[256] = (LFSRcolor1[1048]&LFSRcolor1[677]&LFSRcolor1[1280]&LFSRcolor1[398]);
    BiasedRNG[257] = (LFSRcolor1[299]&LFSRcolor1[1351]&LFSRcolor1[1755]&LFSRcolor1[672]);
    BiasedRNG[258] = (LFSRcolor1[1634]&LFSRcolor1[573]&LFSRcolor1[278]&LFSRcolor1[208]);
    BiasedRNG[259] = (LFSRcolor1[1501]&LFSRcolor1[501]&LFSRcolor1[785]&LFSRcolor1[1193]);
    BiasedRNG[260] = (LFSRcolor1[796]&LFSRcolor1[1598]&LFSRcolor1[1445]&LFSRcolor1[1083]);
    BiasedRNG[261] = (LFSRcolor1[273]&LFSRcolor1[1288]&LFSRcolor1[1019]&LFSRcolor1[1683]);
    BiasedRNG[262] = (LFSRcolor1[229]&LFSRcolor1[160]&LFSRcolor1[1769]&LFSRcolor1[1188]);
    BiasedRNG[263] = (LFSRcolor1[1054]&LFSRcolor1[456]&LFSRcolor1[690]&LFSRcolor1[238]);
    BiasedRNG[264] = (LFSRcolor1[641]&LFSRcolor1[246]&LFSRcolor1[786]&LFSRcolor1[1085]);
    BiasedRNG[265] = (LFSRcolor1[4]&LFSRcolor1[1091]&LFSRcolor1[1562]&LFSRcolor1[696]);
    BiasedRNG[266] = (LFSRcolor1[523]&LFSRcolor1[1706]&LFSRcolor1[1664]&LFSRcolor1[461]);
    BiasedRNG[267] = (LFSRcolor1[470]&LFSRcolor1[50]&LFSRcolor1[992]&LFSRcolor1[59]);
    BiasedRNG[268] = (LFSRcolor1[1062]&LFSRcolor1[874]&LFSRcolor1[106]&LFSRcolor1[729]);
    BiasedRNG[269] = (LFSRcolor1[1382]&LFSRcolor1[1028]&LFSRcolor1[1530]&LFSRcolor1[536]);
    BiasedRNG[270] = (LFSRcolor1[1785]&LFSRcolor1[198]&LFSRcolor1[436]&LFSRcolor1[636]);
    BiasedRNG[271] = (LFSRcolor1[1184]&LFSRcolor1[773]&LFSRcolor1[1169]&LFSRcolor1[1330]);
    BiasedRNG[272] = (LFSRcolor1[1248]&LFSRcolor1[621]&LFSRcolor1[1380]&LFSRcolor1[853]);
    BiasedRNG[273] = (LFSRcolor1[1496]&LFSRcolor1[1057]&LFSRcolor1[430]&LFSRcolor1[814]);
    BiasedRNG[274] = (LFSRcolor1[1182]&LFSRcolor1[1262]&LFSRcolor1[224]&LFSRcolor1[1637]);
    BiasedRNG[275] = (LFSRcolor1[910]&LFSRcolor1[311]&LFSRcolor1[1052]&LFSRcolor1[364]);
    BiasedRNG[276] = (LFSRcolor1[421]&LFSRcolor1[680]&LFSRcolor1[1369]&LFSRcolor1[93]);
    BiasedRNG[277] = (LFSRcolor1[1521]&LFSRcolor1[1323]&LFSRcolor1[1488]&LFSRcolor1[597]);
    BiasedRNG[278] = (LFSRcolor1[85]&LFSRcolor1[728]&LFSRcolor1[1286]&LFSRcolor1[906]);
    BiasedRNG[279] = (LFSRcolor1[528]&LFSRcolor1[262]&LFSRcolor1[359]&LFSRcolor1[1651]);
    BiasedRNG[280] = (LFSRcolor1[345]&LFSRcolor1[979]&LFSRcolor1[542]&LFSRcolor1[617]);
    BiasedRNG[281] = (LFSRcolor1[165]&LFSRcolor1[1660]&LFSRcolor1[1309]&LFSRcolor1[587]);
    BiasedRNG[282] = (LFSRcolor1[998]&LFSRcolor1[74]&LFSRcolor1[404]&LFSRcolor1[584]);
    BiasedRNG[283] = (LFSRcolor1[1332]&LFSRcolor1[288]&LFSRcolor1[1700]&LFSRcolor1[768]);
    BiasedRNG[284] = (LFSRcolor1[904]&LFSRcolor1[1114]&LFSRcolor1[1538]&LFSRcolor1[1476]);
    BiasedRNG[285] = (LFSRcolor1[1224]&LFSRcolor1[261]&LFSRcolor1[691]&LFSRcolor1[350]);
    BiasedRNG[286] = (LFSRcolor1[1561]&LFSRcolor1[757]&LFSRcolor1[154]&LFSRcolor1[1559]);
    BiasedRNG[287] = (LFSRcolor1[1069]&LFSRcolor1[294]&LFSRcolor1[1344]&LFSRcolor1[651]);
    BiasedRNG[288] = (LFSRcolor1[283]&LFSRcolor1[632]&LFSRcolor1[511]&LFSRcolor1[504]);
    BiasedRNG[289] = (LFSRcolor1[1168]&LFSRcolor1[806]&LFSRcolor1[158]&LFSRcolor1[1543]);
    BiasedRNG[290] = (LFSRcolor1[20]&LFSRcolor1[570]&LFSRcolor1[891]&LFSRcolor1[1347]);
    BiasedRNG[291] = (LFSRcolor1[450]&LFSRcolor1[847]&LFSRcolor1[790]&LFSRcolor1[42]);
    BiasedRNG[292] = (LFSRcolor1[991]&LFSRcolor1[118]&LFSRcolor1[424]&LFSRcolor1[1267]);
    BiasedRNG[293] = (LFSRcolor1[1076]&LFSRcolor1[1061]&LFSRcolor1[811]&LFSRcolor1[1682]);
    BiasedRNG[294] = (LFSRcolor1[656]&LFSRcolor1[1746]&LFSRcolor1[1459]&LFSRcolor1[655]);
    BiasedRNG[295] = (LFSRcolor1[1460]&LFSRcolor1[1038]&LFSRcolor1[1234]&LFSRcolor1[639]);
    BiasedRNG[296] = (LFSRcolor1[1597]&LFSRcolor1[661]&LFSRcolor1[589]&LFSRcolor1[1339]);
    BiasedRNG[297] = (LFSRcolor1[1241]&LFSRcolor1[1120]&LFSRcolor1[342]&LFSRcolor1[480]);
    BiasedRNG[298] = (LFSRcolor1[371]&LFSRcolor1[1620]&LFSRcolor1[315]&LFSRcolor1[627]);
    BiasedRNG[299] = (LFSRcolor1[1606]&LFSRcolor1[494]&LFSRcolor1[391]&LFSRcolor1[380]);
    BiasedRNG[300] = (LFSRcolor1[1283]&LFSRcolor1[1163]&LFSRcolor1[778]&LFSRcolor1[509]);
    BiasedRNG[301] = (LFSRcolor1[1406]&LFSRcolor1[755]&LFSRcolor1[1509]&LFSRcolor1[1695]);
    BiasedRNG[302] = (LFSRcolor1[1750]&LFSRcolor1[604]&LFSRcolor1[1471]&LFSRcolor1[1304]);
    BiasedRNG[303] = (LFSRcolor1[1552]&LFSRcolor1[351]&LFSRcolor1[1222]&LFSRcolor1[1490]);
    BiasedRNG[304] = (LFSRcolor1[647]&LFSRcolor1[190]&LFSRcolor1[113]&LFSRcolor1[1692]);
    BiasedRNG[305] = (LFSRcolor1[683]&LFSRcolor1[775]&LFSRcolor1[750]&LFSRcolor1[1625]);
    BiasedRNG[306] = (LFSRcolor1[1440]&LFSRcolor1[1602]&LFSRcolor1[507]&LFSRcolor1[823]);
    BiasedRNG[307] = (LFSRcolor1[1110]&LFSRcolor1[183]&LFSRcolor1[754]&LFSRcolor1[1191]);
    BiasedRNG[308] = (LFSRcolor1[601]&LFSRcolor1[867]&LFSRcolor1[1481]&LFSRcolor1[1420]);
    BiasedRNG[309] = (LFSRcolor1[694]&LFSRcolor1[574]&LFSRcolor1[1009]&LFSRcolor1[78]);
    BiasedRNG[310] = (LFSRcolor1[277]&LFSRcolor1[389]&LFSRcolor1[433]&LFSRcolor1[1467]);
    BiasedRNG[311] = (LFSRcolor1[1022]&LFSRcolor1[684]&LFSRcolor1[1721]&LFSRcolor1[196]);
    BiasedRNG[312] = (LFSRcolor1[1043]&LFSRcolor1[581]&LFSRcolor1[782]&LFSRcolor1[1164]);
    BiasedRNG[313] = (LFSRcolor1[833]&LFSRcolor1[1671]&LFSRcolor1[1599]&LFSRcolor1[894]);
    BiasedRNG[314] = (LFSRcolor1[1282]&LFSRcolor1[1278]&LFSRcolor1[1544]&LFSRcolor1[187]);
    BiasedRNG[315] = (LFSRcolor1[1665]&LFSRcolor1[1541]&LFSRcolor1[537]&LFSRcolor1[1722]);
    BiasedRNG[316] = (LFSRcolor1[486]&LFSRcolor1[312]&LFSRcolor1[538]&LFSRcolor1[900]);
    BiasedRNG[317] = (LFSRcolor1[825]&LFSRcolor1[459]&LFSRcolor1[925]&LFSRcolor1[1029]);
    BiasedRNG[318] = (LFSRcolor1[1174]&LFSRcolor1[919]&LFSRcolor1[993]&LFSRcolor1[241]);
    BiasedRNG[319] = (LFSRcolor1[1197]&LFSRcolor1[413]&LFSRcolor1[170]&LFSRcolor1[640]);
    BiasedRNG[320] = (LFSRcolor1[868]&LFSRcolor1[446]&LFSRcolor1[1461]&LFSRcolor1[422]);
    BiasedRNG[321] = (LFSRcolor1[397]&LFSRcolor1[929]&LFSRcolor1[1423]&LFSRcolor1[846]);
    BiasedRNG[322] = (LFSRcolor1[1441]&LFSRcolor1[1242]&LFSRcolor1[1446]&LFSRcolor1[356]);
    BiasedRNG[323] = (LFSRcolor1[1387]&LFSRcolor1[1104]&LFSRcolor1[378]&LFSRcolor1[736]);
    BiasedRNG[324] = (LFSRcolor1[1698]&LFSRcolor1[265]&LFSRcolor1[855]&LFSRcolor1[94]);
    BiasedRNG[325] = (LFSRcolor1[733]&LFSRcolor1[68]&LFSRcolor1[225]&LFSRcolor1[1108]);
    BiasedRNG[326] = (LFSRcolor1[1112]&LFSRcolor1[1724]&LFSRcolor1[1495]&LFSRcolor1[415]);
    BiasedRNG[327] = (LFSRcolor1[1199]&LFSRcolor1[172]&LFSRcolor1[1153]&LFSRcolor1[1428]);
    BiasedRNG[328] = (LFSRcolor1[1152]&LFSRcolor1[401]&LFSRcolor1[291]&LFSRcolor1[447]);
    BiasedRNG[329] = (LFSRcolor1[107]&LFSRcolor1[1058]&LFSRcolor1[321]&LFSRcolor1[65]);
    BiasedRNG[330] = (LFSRcolor1[1659]&LFSRcolor1[1626]&LFSRcolor1[988]&LFSRcolor1[1210]);
    BiasedRNG[331] = (LFSRcolor1[805]&LFSRcolor1[1192]&LFSRcolor1[1247]&LFSRcolor1[517]);
    BiasedRNG[332] = (LFSRcolor1[396]&LFSRcolor1[88]&LFSRcolor1[1713]&LFSRcolor1[1765]);
    BiasedRNG[333] = (LFSRcolor1[1514]&LFSRcolor1[917]&LFSRcolor1[1001]&LFSRcolor1[1055]);
    BiasedRNG[334] = (LFSRcolor1[652]&LFSRcolor1[791]&LFSRcolor1[1591]&LFSRcolor1[281]);
    BiasedRNG[335] = (LFSRcolor1[1277]&LFSRcolor1[409]&LFSRcolor1[1573]&LFSRcolor1[1741]);
    BiasedRNG[336] = (LFSRcolor1[1523]&LFSRcolor1[673]&LFSRcolor1[1293]&LFSRcolor1[594]);
    BiasedRNG[337] = (LFSRcolor1[477]&LFSRcolor1[1528]&LFSRcolor1[1498]&LFSRcolor1[551]);
    BiasedRNG[338] = (LFSRcolor1[1452]&LFSRcolor1[173]&LFSRcolor1[1784]&LFSRcolor1[1274]);
    BiasedRNG[339] = (LFSRcolor1[1074]&LFSRcolor1[1125]&LFSRcolor1[475]&LFSRcolor1[333]);
    BiasedRNG[340] = (LFSRcolor1[465]&LFSRcolor1[1263]&LFSRcolor1[616]&LFSRcolor1[1571]);
    BiasedRNG[341] = (LFSRcolor1[449]&LFSRcolor1[698]&LFSRcolor1[727]&LFSRcolor1[860]);
    BiasedRNG[342] = (LFSRcolor1[298]&LFSRcolor1[526]&LFSRcolor1[822]&LFSRcolor1[590]);
    BiasedRNG[343] = (LFSRcolor1[452]&LFSRcolor1[1143]&LFSRcolor1[1711]&LFSRcolor1[362]);
    BiasedRNG[344] = (LFSRcolor1[127]&LFSRcolor1[1179]&LFSRcolor1[268]&LFSRcolor1[1566]);
    BiasedRNG[345] = (LFSRcolor1[361]&LFSRcolor1[1699]&LFSRcolor1[1186]&LFSRcolor1[1313]);
    BiasedRNG[346] = (LFSRcolor1[1362]&LFSRcolor1[886]&LFSRcolor1[210]&LFSRcolor1[957]);
    BiasedRNG[347] = (LFSRcolor1[188]&LFSRcolor1[821]&LFSRcolor1[105]&LFSRcolor1[1401]);
    BiasedRNG[348] = (LFSRcolor1[1284]&LFSRcolor1[1118]&LFSRcolor1[890]&LFSRcolor1[560]);
    BiasedRNG[349] = (LFSRcolor1[1775]&LFSRcolor1[379]&LFSRcolor1[175]&LFSRcolor1[1653]);
    BiasedRNG[350] = (LFSRcolor1[1424]&LFSRcolor1[1772]&LFSRcolor1[1458]&LFSRcolor1[923]);
    BiasedRNG[351] = (LFSRcolor1[664]&LFSRcolor1[568]&LFSRcolor1[1209]&LFSRcolor1[1427]);
    BiasedRNG[352] = (LFSRcolor1[1738]&LFSRcolor1[146]&LFSRcolor1[1616]&LFSRcolor1[1771]);
    BiasedRNG[353] = (LFSRcolor1[603]&LFSRcolor1[799]&LFSRcolor1[1223]&LFSRcolor1[1133]);
    BiasedRNG[354] = (LFSRcolor1[1124]&LFSRcolor1[1726]&LFSRcolor1[302]&LFSRcolor1[1273]);
    BiasedRNG[355] = (LFSRcolor1[1582]&LFSRcolor1[1506]&LFSRcolor1[235]&LFSRcolor1[203]);
    BiasedRNG[356] = (LFSRcolor1[687]&LFSRcolor1[1455]&LFSRcolor1[567]&LFSRcolor1[13]);
    BiasedRNG[357] = (LFSRcolor1[1053]&LFSRcolor1[242]&LFSRcolor1[1770]&LFSRcolor1[1757]);
    BiasedRNG[358] = (LFSRcolor1[1610]&LFSRcolor1[615]&LFSRcolor1[676]&LFSRcolor1[1397]);
    BiasedRNG[359] = (LFSRcolor1[301]&LFSRcolor1[431]&LFSRcolor1[387]&LFSRcolor1[240]);
    BiasedRNG[360] = (LFSRcolor1[56]&LFSRcolor1[488]&LFSRcolor1[592]&LFSRcolor1[1676]);
    BiasedRNG[361] = (LFSRcolor1[827]&LFSRcolor1[1754]&LFSRcolor1[1556]&LFSRcolor1[329]);
    BiasedRNG[362] = (LFSRcolor1[583]&LFSRcolor1[503]&LFSRcolor1[1486]&LFSRcolor1[186]);
    BiasedRNG[363] = (LFSRcolor1[275]&LFSRcolor1[1730]&LFSRcolor1[844]&LFSRcolor1[1758]);
    BiasedRNG[364] = (LFSRcolor1[879]&LFSRcolor1[1296]&LFSRcolor1[716]&LFSRcolor1[1714]);
    BiasedRNG[365] = (LFSRcolor1[1639]&LFSRcolor1[1231]&LFSRcolor1[487]&LFSRcolor1[711]);
    BiasedRNG[366] = (LFSRcolor1[539]&LFSRcolor1[1520]&LFSRcolor1[1047]&LFSRcolor1[1761]);
    BiasedRNG[367] = (LFSRcolor1[1244]&LFSRcolor1[1733]&LFSRcolor1[1281]&LFSRcolor1[180]);
    BiasedRNG[368] = (LFSRcolor1[982]&LFSRcolor1[646]&LFSRcolor1[1492]&LFSRcolor1[1448]);
    BiasedRNG[369] = (LFSRcolor1[1400]&LFSRcolor1[21]&LFSRcolor1[1583]&LFSRcolor1[1405]);
    BiasedRNG[370] = (LFSRcolor1[963]&LFSRcolor1[323]&LFSRcolor1[1728]&LFSRcolor1[18]);
    BiasedRNG[371] = (LFSRcolor1[1742]&LFSRcolor1[1317]&LFSRcolor1[213]&LFSRcolor1[739]);
    BiasedRNG[372] = (LFSRcolor1[370]&LFSRcolor1[1553]&LFSRcolor1[922]&LFSRcolor1[1259]);
    BiasedRNG[373] = (LFSRcolor1[1450]&LFSRcolor1[1203]&LFSRcolor1[706]&LFSRcolor1[1516]);
    BiasedRNG[374] = (LFSRcolor1[608]&LFSRcolor1[337]&LFSRcolor1[1513]&LFSRcolor1[1403]);
    BiasedRNG[375] = (LFSRcolor1[330]&LFSRcolor1[168]&LFSRcolor1[482]&LFSRcolor1[514]);
    BiasedRNG[376] = (LFSRcolor1[865]&LFSRcolor1[1285]&LFSRcolor1[132]&LFSRcolor1[474]);
    BiasedRNG[377] = (LFSRcolor1[193]&LFSRcolor1[1404]&LFSRcolor1[521]&LFSRcolor1[961]);
    BiasedRNG[378] = (LFSRcolor1[230]&LFSRcolor1[1790]&LFSRcolor1[1236]&LFSRcolor1[519]);
    BiasedRNG[379] = (LFSRcolor1[284]&LFSRcolor1[912]&LFSRcolor1[1150]&LFSRcolor1[1010]);
    BiasedRNG[380] = (LFSRcolor1[1654]&LFSRcolor1[1144]&LFSRcolor1[496]&LFSRcolor1[1198]);
    BiasedRNG[381] = (LFSRcolor1[215]&LFSRcolor1[1276]&LFSRcolor1[777]&LFSRcolor1[610]);
    BiasedRNG[382] = (LFSRcolor1[958]&LFSRcolor1[204]&LFSRcolor1[1791]&LFSRcolor1[625]);
    BiasedRNG[383] = (LFSRcolor1[293]&LFSRcolor1[1580]&LFSRcolor1[141]&LFSRcolor1[1574]);
    BiasedRNG[384] = (LFSRcolor1[338]&LFSRcolor1[1645]&LFSRcolor1[829]&LFSRcolor1[510]);
    BiasedRNG[385] = (LFSRcolor1[1256]&LFSRcolor1[869]&LFSRcolor1[481]&LFSRcolor1[1303]);
    BiasedRNG[386] = (LFSRcolor1[374]&LFSRcolor1[9]&LFSRcolor1[1158]&LFSRcolor1[1723]);
    BiasedRNG[387] = (LFSRcolor1[492]&LFSRcolor1[1740]&LFSRcolor1[942]&LFSRcolor1[873]);
    BiasedRNG[388] = (LFSRcolor1[1097]&LFSRcolor1[55]&LFSRcolor1[92]&LFSRcolor1[662]);
    BiasedRNG[389] = (LFSRcolor1[956]&LFSRcolor1[1385]&LFSRcolor1[813]&LFSRcolor1[1178]);
    BiasedRNG[390] = (LFSRcolor1[1527]&LFSRcolor1[1340]&LFSRcolor1[1099]&LFSRcolor1[289]);
    BiasedRNG[391] = (LFSRcolor1[1375]&LFSRcolor1[740]&LFSRcolor1[419]&LFSRcolor1[642]);
    BiasedRNG[392] = (LFSRcolor1[572]&LFSRcolor1[845]&LFSRcolor1[1250]&LFSRcolor1[1046]);
    BiasedRNG[393] = (LFSRcolor1[780]&LFSRcolor1[606]&LFSRcolor1[1066]&LFSRcolor1[882]);
    BiasedRNG[394] = (LFSRcolor1[667]&LFSRcolor1[975]&LFSRcolor1[971]&LFSRcolor1[1454]);
    BiasedRNG[395] = (LFSRcolor1[1697]&LFSRcolor1[1589]&LFSRcolor1[1564]&LFSRcolor1[1220]);
    BiasedRNG[396] = (LFSRcolor1[1594]&LFSRcolor1[157]&LFSRcolor1[1111]&LFSRcolor1[820]);
    BiasedRNG[397] = (LFSRcolor1[162]&LFSRcolor1[233]&LFSRcolor1[1491]&LFSRcolor1[239]);
    BiasedRNG[398] = (LFSRcolor1[1675]&LFSRcolor1[471]&LFSRcolor1[803]&LFSRcolor1[1008]);
    BiasedRNG[399] = (LFSRcolor1[544]&LFSRcolor1[264]&LFSRcolor1[668]&LFSRcolor1[741]);
    BiasedRNG[400] = (LFSRcolor1[148]&LFSRcolor1[654]&LFSRcolor1[279]&LFSRcolor1[735]);
    BiasedRNG[401] = (LFSRcolor1[100]&LFSRcolor1[947]&LFSRcolor1[365]&LFSRcolor1[1018]);
    BiasedRNG[402] = (LFSRcolor1[1684]&LFSRcolor1[1253]&LFSRcolor1[566]&LFSRcolor1[300]);
    BiasedRNG[403] = (LFSRcolor1[1079]&LFSRcolor1[1050]&LFSRcolor1[1444]&LFSRcolor1[1792]);
    BiasedRNG[404] = (LFSRcolor1[1302]&LFSRcolor1[732]&LFSRcolor1[527]&LFSRcolor1[776]);
    BiasedRNG[405] = (LFSRcolor1[967]&LFSRcolor1[1127]&LFSRcolor1[506]&LFSRcolor1[562]);
    BiasedRNG[406] = (LFSRcolor1[864]&LFSRcolor1[1702]&LFSRcolor1[1640]&LFSRcolor1[1147]);
    BiasedRNG[407] = (LFSRcolor1[1202]&LFSRcolor1[326]&LFSRcolor1[637]&LFSRcolor1[395]);
    BiasedRNG[408] = (LFSRcolor1[1389]&LFSRcolor1[1013]&LFSRcolor1[1685]&LFSRcolor1[473]);
    BiasedRNG[409] = (LFSRcolor1[792]&LFSRcolor1[466]&LFSRcolor1[334]&LFSRcolor1[1297]);
    BiasedRNG[410] = (LFSRcolor1[838]&LFSRcolor1[1151]&LFSRcolor1[1525]&LFSRcolor1[400]);
    BiasedRNG[411] = (LFSRcolor1[256]&LFSRcolor1[842]&LFSRcolor1[455]&LFSRcolor1[1672]);
    BiasedRNG[412] = (LFSRcolor1[1005]&LFSRcolor1[439]&LFSRcolor1[1155]&LFSRcolor1[1100]);
    BiasedRNG[413] = (LFSRcolor1[406]&LFSRcolor1[403]&LFSRcolor1[1352]&LFSRcolor1[850]);
    BiasedRNG[414] = (LFSRcolor1[1609]&LFSRcolor1[1252]&LFSRcolor1[1305]&LFSRcolor1[1381]);
    BiasedRNG[415] = (LFSRcolor1[658]&LFSRcolor1[1355]&LFSRcolor1[1260]&LFSRcolor1[1780]);
    BiasedRNG[416] = (LFSRcolor1[940]&LFSRcolor1[102]&LFSRcolor1[631]&LFSRcolor1[1107]);
    BiasedRNG[417] = (LFSRcolor1[73]&LFSRcolor1[1629]&LFSRcolor1[1652]&LFSRcolor1[650]);
    BiasedRNG[418] = (LFSRcolor1[1668]&LFSRcolor1[1534]&LFSRcolor1[211]&LFSRcolor1[1181]);
    BiasedRNG[419] = (LFSRcolor1[1628]&LFSRcolor1[714]&LFSRcolor1[81]&LFSRcolor1[804]);
    BiasedRNG[420] = (LFSRcolor1[497]&LFSRcolor1[1663]&LFSRcolor1[819]&LFSRcolor1[1307]);
    BiasedRNG[421] = (LFSRcolor1[1216]&LFSRcolor1[810]&LFSRcolor1[1291]&LFSRcolor1[1033]);
    BiasedRNG[422] = (LFSRcolor1[98]&LFSRcolor1[1542]&LFSRcolor1[1679]&LFSRcolor1[255]);
    BiasedRNG[423] = (LFSRcolor1[788]&LFSRcolor1[237]&LFSRcolor1[1778]&LFSRcolor1[888]);
    BiasedRNG[424] = (LFSRcolor1[410]&LFSRcolor1[1195]&LFSRcolor1[1557]&LFSRcolor1[795]);
    BiasedRNG[425] = (LFSRcolor1[1311]&LFSRcolor1[1732]&LFSRcolor1[898]&LFSRcolor1[5]);
    BiasedRNG[426] = (LFSRcolor1[575]&LFSRcolor1[31]&LFSRcolor1[1425]&LFSRcolor1[1254]);
    BiasedRNG[427] = (LFSRcolor1[828]&LFSRcolor1[1788]&LFSRcolor1[505]&LFSRcolor1[765]);
    BiasedRNG[428] = (LFSRcolor1[686]&LFSRcolor1[1226]&LFSRcolor1[1270]&LFSRcolor1[1690]);
    BiasedRNG[429] = (LFSRcolor1[1088]&LFSRcolor1[166]&LFSRcolor1[989]&LFSRcolor1[1632]);
    BiasedRNG[430] = (LFSRcolor1[19]&LFSRcolor1[1023]&LFSRcolor1[34]&LFSRcolor1[336]);
    BiasedRNG[431] = (LFSRcolor1[1363]&LFSRcolor1[1457]&LFSRcolor1[981]&LFSRcolor1[1656]);
    BiasedRNG[432] = (LFSRcolor1[1658]&LFSRcolor1[248]&LFSRcolor1[761]&LFSRcolor1[685]);
    BiasedRNG[433] = (LFSRcolor1[1781]&LFSRcolor1[1185]&LFSRcolor1[174]&LFSRcolor1[263]);
    BiasedRNG[434] = (LFSRcolor1[1753]&LFSRcolor1[36]&LFSRcolor1[937]&LFSRcolor1[783]);
    BiasedRNG[435] = (LFSRcolor1[1670]&LFSRcolor1[1157]&LFSRcolor1[427]&LFSRcolor1[665]);
    BiasedRNG[436] = (LFSRcolor1[223]&LFSRcolor1[554]&LFSRcolor1[1774]&LFSRcolor1[1014]);
    BiasedRNG[437] = (LFSRcolor1[1434]&LFSRcolor1[1529]&LFSRcolor1[987]&LFSRcolor1[1535]);
    BiasedRNG[438] = (LFSRcolor1[1171]&LFSRcolor1[354]&LFSRcolor1[156]&LFSRcolor1[1522]);
    BiasedRNG[439] = (LFSRcolor1[306]&LFSRcolor1[495]&LFSRcolor1[270]&LFSRcolor1[969]);
    BiasedRNG[440] = (LFSRcolor1[124]&LFSRcolor1[644]&LFSRcolor1[458]&LFSRcolor1[897]);
    BiasedRNG[441] = (LFSRcolor1[307]&LFSRcolor1[525]&LFSRcolor1[1419]&LFSRcolor1[131]);
    BiasedRNG[442] = (LFSRcolor1[1624]&LFSRcolor1[493]&LFSRcolor1[390]&LFSRcolor1[144]);
    BiasedRNG[443] = (LFSRcolor1[1443]&LFSRcolor1[340]&LFSRcolor1[214]&LFSRcolor1[1357]);
    BiasedRNG[444] = (LFSRcolor1[876]&LFSRcolor1[1229]&LFSRcolor1[695]&LFSRcolor1[564]);
    BiasedRNG[445] = (LFSRcolor1[1265]&LFSRcolor1[1167]&LFSRcolor1[70]&LFSRcolor1[1484]);
    BiasedRNG[446] = (LFSRcolor1[1575]&LFSRcolor1[547]&LFSRcolor1[1130]&LFSRcolor1[508]);
    BiasedRNG[447] = (LFSRcolor1[76]&LFSRcolor1[22]&LFSRcolor1[1678]&LFSRcolor1[7]);
    BiasedRNG[448] = (LFSRcolor1[258]&LFSRcolor1[414]&LFSRcolor1[434]&LFSRcolor1[161]);
    BiasedRNG[449] = (LFSRcolor1[1207]&LFSRcolor1[1334]&LFSRcolor1[80]&LFSRcolor1[1708]);
    BiasedRNG[450] = (LFSRcolor1[600]&LFSRcolor1[1370]&LFSRcolor1[290]&LFSRcolor1[902]);
    BiasedRNG[451] = (LFSRcolor1[938]&LFSRcolor1[1408]&LFSRcolor1[1603]&LFSRcolor1[1601]);
    BiasedRNG[452] = (LFSRcolor1[1719]&LFSRcolor1[69]&LFSRcolor1[82]&LFSRcolor1[558]);
    BiasedRNG[453] = (LFSRcolor1[1123]&LFSRcolor1[123]&LFSRcolor1[1479]&LFSRcolor1[1103]);
    BiasedRNG[454] = (LFSRcolor1[1237]&LFSRcolor1[797]&LFSRcolor1[620]&LFSRcolor1[1696]);
    BiasedRNG[455] = (LFSRcolor1[478]&LFSRcolor1[366]&LFSRcolor1[1243]&LFSRcolor1[14]);
    BiasedRNG[456] = (LFSRcolor1[27]&LFSRcolor1[502]&LFSRcolor1[1051]&LFSRcolor1[479]);
    BiasedRNG[457] = (LFSRcolor1[420]&LFSRcolor1[793]&LFSRcolor1[816]&LFSRcolor1[1249]);
    BiasedRNG[458] = (LFSRcolor1[416]&LFSRcolor1[725]&LFSRcolor1[1453]&LFSRcolor1[95]);
    BiasedRNG[459] = (LFSRcolor1[79]&LFSRcolor1[1470]&LFSRcolor1[1673]&LFSRcolor1[199]);
    BiasedRNG[460] = (LFSRcolor1[1680]&LFSRcolor1[1140]&LFSRcolor1[83]&LFSRcolor1[1737]);
    BiasedRNG[461] = (LFSRcolor1[1377]&LFSRcolor1[71]&LFSRcolor1[1605]&LFSRcolor1[946]);
    BiasedRNG[462] = (LFSRcolor1[1314]&LFSRcolor1[1578]&LFSRcolor1[341]&LFSRcolor1[1190]);
    BiasedRNG[463] = (LFSRcolor1[460]&LFSRcolor1[442]&LFSRcolor1[405]&LFSRcolor1[1301]);
    BiasedRNG[464] = (LFSRcolor1[1655]&LFSRcolor1[895]&LFSRcolor1[423]&LFSRcolor1[1555]);
    BiasedRNG[465] = (LFSRcolor1[1392]&LFSRcolor1[1608]&LFSRcolor1[1217]&LFSRcolor1[1462]);
    BiasedRNG[466] = (LFSRcolor1[375]&LFSRcolor1[1275]&LFSRcolor1[1762]&LFSRcolor1[349]);
    BiasedRNG[467] = (LFSRcolor1[1494]&LFSRcolor1[355]&LFSRcolor1[638]&LFSRcolor1[1617]);
    BiasedRNG[468] = (LFSRcolor1[1517]&LFSRcolor1[1084]&LFSRcolor1[1098]&LFSRcolor1[1271]);
    BiasedRNG[469] = (LFSRcolor1[1393]&LFSRcolor1[1004]&LFSRcolor1[292]&LFSRcolor1[363]);
    BiasedRNG[470] = (LFSRcolor1[1507]&LFSRcolor1[140]&LFSRcolor1[1438]&LFSRcolor1[1464]);
    BiasedRNG[471] = (LFSRcolor1[901]&LFSRcolor1[875]&LFSRcolor1[759]&LFSRcolor1[1101]);
    BiasedRNG[472] = (LFSRcolor1[936]&LFSRcolor1[109]&LFSRcolor1[1748]&LFSRcolor1[195]);
    BiasedRNG[473] = (LFSRcolor1[457]&LFSRcolor1[159]&LFSRcolor1[871]&LFSRcolor1[1593]);
    BiasedRNG[474] = (LFSRcolor1[220]&LFSRcolor1[701]&LFSRcolor1[878]&LFSRcolor1[1166]);
    BiasedRNG[475] = (LFSRcolor1[682]&LFSRcolor1[1327]&LFSRcolor1[201]&LFSRcolor1[353]);
    BiasedRNG[476] = (LFSRcolor1[1218]&LFSRcolor1[854]&LFSRcolor1[674]&LFSRcolor1[185]);
    BiasedRNG[477] = (LFSRcolor1[16]&LFSRcolor1[1568]&LFSRcolor1[1550]&LFSRcolor1[1213]);
    BiasedRNG[478] = (LFSRcolor1[1482]&LFSRcolor1[206]&LFSRcolor1[57]&LFSRcolor1[1077]);
    BiasedRNG[479] = (LFSRcolor1[1487]&LFSRcolor1[742]&LFSRcolor1[310]&LFSRcolor1[1430]);
    BiasedRNG[480] = (LFSRcolor1[522]&LFSRcolor1[950]&LFSRcolor1[216]&LFSRcolor1[563]);
    BiasedRNG[481] = (LFSRcolor1[115]&LFSRcolor1[812]&LFSRcolor1[12]&LFSRcolor1[815]);
    BiasedRNG[482] = (LFSRcolor1[1709]&LFSRcolor1[1070]&LFSRcolor1[1094]&LFSRcolor1[1090]);
    BiasedRNG[483] = (LFSRcolor1[1080]&LFSRcolor1[934]&LFSRcolor1[1376]&LFSRcolor1[29]);
    BiasedRNG[484] = (LFSRcolor1[862]&LFSRcolor1[908]&LFSRcolor1[303]&LFSRcolor1[1451]);
    BiasedRNG[485] = (LFSRcolor1[51]&LFSRcolor1[970]&LFSRcolor1[1636]&LFSRcolor1[15]);
    BiasedRNG[486] = (LFSRcolor1[181]&LFSRcolor1[712]&LFSRcolor1[531]&LFSRcolor1[756]);
    BiasedRNG[487] = (LFSRcolor1[1402]&LFSRcolor1[976]&LFSRcolor1[763]&LFSRcolor1[1214]);
    BiasedRNG[488] = (LFSRcolor1[1786]&LFSRcolor1[296]&LFSRcolor1[626]&LFSRcolor1[393]);
    BiasedRNG[489] = (LFSRcolor1[1413]&LFSRcolor1[914]&LFSRcolor1[679]&LFSRcolor1[1312]);
    BiasedRNG[490] = (LFSRcolor1[1793]&LFSRcolor1[121]&LFSRcolor1[1136]&LFSRcolor1[319]);
    BiasedRNG[491] = (LFSRcolor1[624]&LFSRcolor1[357]&LFSRcolor1[1519]&LFSRcolor1[807]);
    BiasedRNG[492] = (LFSRcolor1[718]&LFSRcolor1[128]&LFSRcolor1[535]&LFSRcolor1[1264]);
    BiasedRNG[493] = (LFSRcolor1[1060]&LFSRcolor1[697]&LFSRcolor1[669]&LFSRcolor1[444]);
    BiasedRNG[494] = (LFSRcolor1[1546]&LFSRcolor1[1745]&LFSRcolor1[46]&LFSRcolor1[630]);
    BiasedRNG[495] = (LFSRcolor1[476]&LFSRcolor1[1777]&LFSRcolor1[1417]&LFSRcolor1[1040]);
    BiasedRNG[496] = (LFSRcolor1[1142]&LFSRcolor1[746]&LFSRcolor1[1439]&LFSRcolor1[1649]);
    BiasedRNG[497] = (LFSRcolor1[675]&LFSRcolor1[885]&LFSRcolor1[72]&LFSRcolor1[145]);
    BiasedRNG[498] = (LFSRcolor1[689]&LFSRcolor1[1082]&LFSRcolor1[45]&LFSRcolor1[1731]);
    BiasedRNG[499] = (LFSRcolor1[1162]&LFSRcolor1[150]&LFSRcolor1[1502]&LFSRcolor1[599]);
    BiasedRNG[500] = (LFSRcolor1[1701]&LFSRcolor1[653]&LFSRcolor1[693]&LFSRcolor1[41]);
    BiasedRNG[501] = (LFSRcolor1[1266]&LFSRcolor1[1346]&LFSRcolor1[468]&LFSRcolor1[830]);
    BiasedRNG[502] = (LFSRcolor1[324]&LFSRcolor1[1141]&LFSRcolor1[1328]&LFSRcolor1[108]);
    BiasedRNG[503] = (LFSRcolor1[25]&LFSRcolor1[962]&LFSRcolor1[723]&LFSRcolor1[1586]);
    BiasedRNG[504] = (LFSRcolor1[751]&LFSRcolor1[1478]&LFSRcolor1[179]&LFSRcolor1[1073]);
    BiasedRNG[505] = (LFSRcolor1[1364]&LFSRcolor1[1474]&LFSRcolor1[184]&LFSRcolor1[305]);
    BiasedRNG[506] = (LFSRcolor1[951]&LFSRcolor1[818]&LFSRcolor1[1418]&LFSRcolor1[125]);
    BiasedRNG[507] = (LFSRcolor1[817]&LFSRcolor1[1691]&LFSRcolor1[1246]&LFSRcolor1[231]);
    BiasedRNG[508] = (LFSRcolor1[276]&LFSRcolor1[1409]&LFSRcolor1[1044]&LFSRcolor1[1315]);
    BiasedRNG[509] = (LFSRcolor1[1768]&LFSRcolor1[1547]&LFSRcolor1[1384]&LFSRcolor1[28]);
    BiasedRNG[510] = (LFSRcolor1[1576]&LFSRcolor1[565]&LFSRcolor1[1065]&LFSRcolor1[995]);
    BiasedRNG[511] = (LFSRcolor1[429]&LFSRcolor1[1725]&LFSRcolor1[1093]&LFSRcolor1[1071]);
    BiasedRNG[512] = (LFSRcolor1[1134]&LFSRcolor1[1595]&LFSRcolor1[1776]&LFSRcolor1[1623]);
    BiasedRNG[513] = (LFSRcolor1[927]&LFSRcolor1[205]&LFSRcolor1[1592]&LFSRcolor1[454]);
    BiasedRNG[514] = (LFSRcolor1[848]&LFSRcolor1[724]&LFSRcolor1[217]&LFSRcolor1[119]);
    BiasedRNG[515] = (LFSRcolor1[1704]&LFSRcolor1[111]&LFSRcolor1[163]&LFSRcolor1[1326]);
    BiasedRNG[516] = (LFSRcolor1[135]&LFSRcolor1[1666]&LFSRcolor1[130]&LFSRcolor1[48]);
    BiasedRNG[517] = (LFSRcolor1[808]&LFSRcolor1[1643]&LFSRcolor1[126]&LFSRcolor1[703]);
    BiasedRNG[518] = (LFSRcolor1[999]&LFSRcolor1[1611]&LFSRcolor1[634]&LFSRcolor1[1383]);
    BiasedRNG[519] = (LFSRcolor1[985]&LFSRcolor1[760]&LFSRcolor1[43]&LFSRcolor1[1356]);
    BiasedRNG[520] = (LFSRcolor1[44]&LFSRcolor1[1485]&LFSRcolor1[1365]&LFSRcolor1[924]);
    BiasedRNG[521] = (LFSRcolor1[1548]&LFSRcolor1[832]&LFSRcolor1[1015]&LFSRcolor1[1705]);
    BiasedRNG[522] = (LFSRcolor1[1113]&LFSRcolor1[1426]&LFSRcolor1[699]&LFSRcolor1[670]);
    BiasedRNG[523] = (LFSRcolor1[464]&LFSRcolor1[809]&LFSRcolor1[933]&LFSRcolor1[1343]);
    BiasedRNG[524] = (LFSRcolor1[253]&LFSRcolor1[1333]&LFSRcolor1[1407]&LFSRcolor1[984]);
    BiasedRNG[525] = (LFSRcolor1[1261]&LFSRcolor1[1642]&LFSRcolor1[1394]&LFSRcolor1[591]);
    BiasedRNG[526] = (LFSRcolor1[96]&LFSRcolor1[194]&LFSRcolor1[53]&LFSRcolor1[1075]);
    BiasedRNG[527] = (LFSRcolor1[1515]&LFSRcolor1[671]&LFSRcolor1[960]&LFSRcolor1[1059]);
    BiasedRNG[528] = (LFSRcolor1[861]&LFSRcolor1[543]&LFSRcolor1[192]&LFSRcolor1[1729]);
    BiasedRNG[529] = (LFSRcolor1[200]&LFSRcolor1[779]&LFSRcolor1[1067]&LFSRcolor1[1206]);
    BiasedRNG[530] = (LFSRcolor1[1225]&LFSRcolor1[1]&LFSRcolor1[533]&LFSRcolor1[66]);
    BiasedRNG[531] = (LFSRcolor1[997]&LFSRcolor1[764]&LFSRcolor1[86]&LFSRcolor1[1787]);
    BiasedRNG[532] = (LFSRcolor1[1739]&LFSRcolor1[1449]&LFSRcolor1[1122]&LFSRcolor1[588]);
    BiasedRNG[533] = (LFSRcolor1[841]&LFSRcolor1[541]&LFSRcolor1[1289]&LFSRcolor1[708]);
    BiasedRNG[534] = (LFSRcolor1[1138]&LFSRcolor1[114]&LFSRcolor1[498]&LFSRcolor1[789]);
    BiasedRNG[535] = (LFSRcolor1[251]&LFSRcolor1[1034]&LFSRcolor1[612]&LFSRcolor1[1681]);
    BiasedRNG[536] = (LFSRcolor1[207]&LFSRcolor1[1360]&LFSRcolor1[707]&LFSRcolor1[1290]);
    BiasedRNG[537] = (LFSRcolor1[1504]&LFSRcolor1[483]&LFSRcolor1[138]&LFSRcolor1[836]);
    BiasedRNG[538] = (LFSRcolor1[1587]&LFSRcolor1[1779]&LFSRcolor1[308]&LFSRcolor1[889]);
    BiasedRNG[539] = (LFSRcolor1[1627]&LFSRcolor1[1359]&LFSRcolor1[602]&LFSRcolor1[189]);
    BiasedRNG[540] = (LFSRcolor1[771]&LFSRcolor1[1176]&LFSRcolor1[1024]&LFSRcolor1[1358]);
    BiasedRNG[541] = (LFSRcolor1[1433]&LFSRcolor1[129]&LFSRcolor1[139]&LFSRcolor1[182]);
    BiasedRNG[542] = (LFSRcolor1[32]&LFSRcolor1[1087]&LFSRcolor1[112]&LFSRcolor1[1512]);
    BiasedRNG[543] = (LFSRcolor1[609]&LFSRcolor1[1751]&LFSRcolor1[943]&LFSRcolor1[1016]);
    BiasedRNG[544] = (LFSRcolor1[35]&LFSRcolor1[1532]&LFSRcolor1[663]&LFSRcolor1[1341]);
    BiasedRNG[545] = (LFSRcolor1[994]&LFSRcolor1[499]&LFSRcolor1[411]&LFSRcolor1[1577]);
    BiasedRNG[546] = (LFSRcolor1[1508]&LFSRcolor1[717]&LFSRcolor1[347]&LFSRcolor1[866]);
    BiasedRNG[547] = (LFSRcolor1[843]&LFSRcolor1[660]&LFSRcolor1[64]&LFSRcolor1[197]);
    BiasedRNG[548] = (LFSRcolor1[1579]&LFSRcolor1[332]&LFSRcolor1[1388]&LFSRcolor1[408]);
    BiasedRNG[549] = (LFSRcolor1[1378]&LFSRcolor1[425]&LFSRcolor1[623]&LFSRcolor1[167]);
    BiasedRNG[550] = (LFSRcolor1[611]&LFSRcolor1[681]&LFSRcolor1[1089]&LFSRcolor1[965]);
    BiasedRNG[551] = (LFSRcolor1[1279]&LFSRcolor1[1316]&LFSRcolor1[954]&LFSRcolor1[392]);
    BiasedRNG[552] = (LFSRcolor1[1221]&LFSRcolor1[688]&LFSRcolor1[1227]&LFSRcolor1[155]);
    BiasedRNG[553] = (LFSRcolor1[297]&LFSRcolor1[142]&LFSRcolor1[441]&LFSRcolor1[935]);
    BiasedRNG[554] = (LFSRcolor1[1161]&LFSRcolor1[1391]&LFSRcolor1[835]&LFSRcolor1[151]);
    BiasedRNG[555] = (LFSRcolor1[593]&LFSRcolor1[1002]&LFSRcolor1[881]&LFSRcolor1[372]);
    BiasedRNG[556] = (LFSRcolor1[1475]&LFSRcolor1[840]&LFSRcolor1[218]&LFSRcolor1[1641]);
    BiasedRNG[557] = (LFSRcolor1[1092]&LFSRcolor1[62]&LFSRcolor1[1483]&LFSRcolor1[1773]);
    BiasedRNG[558] = (LFSRcolor1[955]&LFSRcolor1[752]&LFSRcolor1[1416]&LFSRcolor1[939]);
    BiasedRNG[559] = (LFSRcolor1[1148]&LFSRcolor1[1635]&LFSRcolor1[77]&LFSRcolor1[1614]);
    BiasedRNG[560] = (LFSRcolor1[628]&LFSRcolor1[1049]&LFSRcolor1[1064]&LFSRcolor1[932]);
    BiasedRNG[561] = (LFSRcolor1[870]&LFSRcolor1[1379]&LFSRcolor1[1563]&LFSRcolor1[1096]);
    BiasedRNG[562] = (LFSRcolor1[1390]&LFSRcolor1[1612]&LFSRcolor1[318]&LFSRcolor1[1109]);
    BiasedRNG[563] = (LFSRcolor1[1036]&LFSRcolor1[47]&LFSRcolor1[1415]&LFSRcolor1[1622]);
    BiasedRNG[564] = (LFSRcolor1[120]&LFSRcolor1[343]&LFSRcolor1[1063]&LFSRcolor1[1505]);
    BiasedRNG[565] = (LFSRcolor1[916]&LFSRcolor1[872]&LFSRcolor1[438]&LFSRcolor1[1117]);
    BiasedRNG[566] = (LFSRcolor1[1646]&LFSRcolor1[1412]&LFSRcolor1[339]&LFSRcolor1[743]);
    BiasedRNG[567] = (LFSRcolor1[1056]&LFSRcolor1[726]&LFSRcolor1[445]&LFSRcolor1[1354]);
    BiasedRNG[568] = (LFSRcolor1[1533]&LFSRcolor1[1027]&LFSRcolor1[1102]&LFSRcolor1[952]);
    BiasedRNG[569] = (LFSRcolor1[1121]&LFSRcolor1[1473]&LFSRcolor1[271]&LFSRcolor1[383]);
    BiasedRNG[570] = (LFSRcolor1[346]&LFSRcolor1[1238]&LFSRcolor1[1716]&LFSRcolor1[147]);
    BiasedRNG[571] = (LFSRcolor1[884]&LFSRcolor1[973]&LFSRcolor1[974]&LFSRcolor1[287]);
    BiasedRNG[572] = (LFSRcolor1[734]&LFSRcolor1[1715]&LFSRcolor1[585]&LFSRcolor1[101]);
    BiasedRNG[573] = (LFSRcolor1[1693]&LFSRcolor1[1421]&LFSRcolor1[1287]&LFSRcolor1[1782]);
    BiasedRNG[574] = (LFSRcolor1[1510]&LFSRcolor1[1456]&LFSRcolor1[54]&LFSRcolor1[1319]);
    BiasedRNG[575] = (LFSRcolor1[905]&LFSRcolor1[918]&LFSRcolor1[1030]&LFSRcolor1[1688]);
    BiasedRNG[576] = (LFSRcolor1[1095]&LFSRcolor1[949]&LFSRcolor1[529]&LFSRcolor1[1647]);
    BiasedRNG[577] = (LFSRcolor1[8]&LFSRcolor1[1045]&LFSRcolor1[177]&LFSRcolor1[103]);
    BiasedRNG[578] = (LFSRcolor1[1531]&LFSRcolor1[1736]&LFSRcolor1[191]&LFSRcolor1[1031]);
    BiasedRNG[579] = (LFSRcolor1[1350]&LFSRcolor1[709]&LFSRcolor1[692]&LFSRcolor1[972]);
    BiasedRNG[580] = (LFSRcolor1[1560]&LFSRcolor1[512]&LFSRcolor1[266]&LFSRcolor1[931]);
    BiasedRNG[581] = (LFSRcolor1[1661]&LFSRcolor1[1156]&LFSRcolor1[605]&LFSRcolor1[1630]);
    BiasedRNG[582] = (LFSRcolor1[63]&LFSRcolor1[1257]&LFSRcolor1[99]&LFSRcolor1[831]);
    BiasedRNG[583] = (LFSRcolor1[896]&LFSRcolor1[657]&LFSRcolor1[1437]&LFSRcolor1[49]);
    BiasedRNG[584] = (LFSRcolor1[1549]&LFSRcolor1[1763]&LFSRcolor1[178]&LFSRcolor1[67]);
    BiasedRNG[585] = (LFSRcolor1[91]&LFSRcolor1[983]&LFSRcolor1[39]&LFSRcolor1[1230]);
    BiasedRNG[586] = (LFSRcolor1[426]&LFSRcolor1[877]&LFSRcolor1[3]&LFSRcolor1[1756]);
    BiasedRNG[587] = (LFSRcolor1[1017]&LFSRcolor1[1233]&LFSRcolor1[580]&LFSRcolor1[309]);
    BiasedRNG[588] = (LFSRcolor1[462]&LFSRcolor1[317]&LFSRcolor1[328]&LFSRcolor1[834]);
    BiasedRNG[589] = (LFSRcolor1[1137]&LFSRcolor1[313]&LFSRcolor1[252]&LFSRcolor1[267]);
    BiasedRNG[590] = (LFSRcolor1[578]&LFSRcolor1[1020]&LFSRcolor1[758]&LFSRcolor1[1743]);
    BiasedRNG[591] = (LFSRcolor1[883]&LFSRcolor1[327]&LFSRcolor1[388]&LFSRcolor1[596]);
    BiasedRNG[592] = (LFSRcolor1[622]&LFSRcolor1[659]&LFSRcolor1[122]&LFSRcolor1[491]);
    BiasedRNG[593] = (LFSRcolor1[1300]&LFSRcolor1[1524]&LFSRcolor1[1135]&LFSRcolor1[635]);
    BiasedRNG[594] = (LFSRcolor1[1411]&LFSRcolor1[1613]&LFSRcolor1[2]&LFSRcolor1[17]);
    BiasedRNG[595] = (LFSRcolor1[1650]&LFSRcolor1[801]&LFSRcolor1[1146]&LFSRcolor1[137]);
    BiasedRNG[596] = (LFSRcolor1[1442]&LFSRcolor1[1235]&LFSRcolor1[280]&LFSRcolor1[133]);
    BiasedRNG[597] = (LFSRcolor1[1194]&LFSRcolor1[6]&LFSRcolor1[472]&LFSRcolor1[1707]);
    BiasedRNG[598] = (LFSRcolor1[232]&LFSRcolor1[1749]&LFSRcolor1[209]&LFSRcolor1[90]);
    BiasedRNG[599] = (LFSRcolor1[1766]&LFSRcolor1[1011]&LFSRcolor1[545]&LFSRcolor1[515]);
    BiasedRNG[600] = (LFSRcolor1[376]&LFSRcolor1[1689]&LFSRcolor1[1255]&LFSRcolor1[1489]);
    BiasedRNG[601] = (LFSRcolor1[37]&LFSRcolor1[247]&LFSRcolor1[1588]&LFSRcolor1[75]);
    BiasedRNG[602] = (LFSRcolor1[1299]&LFSRcolor1[1345]&LFSRcolor1[1183]&LFSRcolor1[490]);
    BiasedRNG[603] = (LFSRcolor1[1126]&LFSRcolor1[550]&LFSRcolor1[1211]&LFSRcolor1[1615]);
    BiasedRNG[604] = (LFSRcolor1[944]&LFSRcolor1[1041]&LFSRcolor1[1078]&LFSRcolor1[959]);
    BiasedRNG[605] = (LFSRcolor1[451]&LFSRcolor1[1175]&LFSRcolor1[721]&LFSRcolor1[953]);
    BiasedRNG[606] = (LFSRcolor1[1325]&LFSRcolor1[556]&LFSRcolor1[532]&LFSRcolor1[61]);
    BiasedRNG[607] = (LFSRcolor1[176]&LFSRcolor1[629]&LFSRcolor1[715]&LFSRcolor1[1349]);
    BiasedRNG[608] = (LFSRcolor1[1129]&LFSRcolor1[1747]&LFSRcolor1[453]&LFSRcolor1[222]);
    BiasedRNG[609] = (LFSRcolor1[402]&LFSRcolor1[282]&LFSRcolor1[1035]&LFSRcolor1[762]);
    BiasedRNG[610] = (LFSRcolor1[87]&LFSRcolor1[704]&LFSRcolor1[1145]&LFSRcolor1[1395]);
    BiasedRNG[611] = (LFSRcolor1[1294]&LFSRcolor1[1324]&LFSRcolor1[557]&LFSRcolor1[1477]);
    BiasedRNG[612] = (LFSRcolor1[134]&LFSRcolor1[548]&LFSRcolor1[1429]&LFSRcolor1[1187]);
    BiasedRNG[613] = (LFSRcolor1[1177]&LFSRcolor1[559]&LFSRcolor1[1604]&LFSRcolor1[325]);
    BiasedRNG[614] = (LFSRcolor1[1321]&LFSRcolor1[1386]&LFSRcolor1[966]&LFSRcolor1[720]);
    BiasedRNG[615] = (LFSRcolor1[858]&LFSRcolor1[666]&LFSRcolor1[1596]&LFSRcolor1[913]);
    BiasedRNG[616] = (LFSRcolor1[619]&LFSRcolor1[171]&LFSRcolor1[443]&LFSRcolor1[555]);
    BiasedRNG[617] = (LFSRcolor1[784]&LFSRcolor1[1196]&LFSRcolor1[513]&LFSRcolor1[1585]);
    BiasedRNG[618] = (LFSRcolor1[254]&LFSRcolor1[772]&LFSRcolor1[986]&LFSRcolor1[770]);
    BiasedRNG[619] = (LFSRcolor1[1320]&LFSRcolor1[990]&LFSRcolor1[1106]&LFSRcolor1[1007]);
    BiasedRNG[620] = (LFSRcolor1[702]&LFSRcolor1[1764]&LFSRcolor1[377]&LFSRcolor1[463]);
    BiasedRNG[621] = (LFSRcolor1[643]&LFSRcolor1[534]&LFSRcolor1[1584]&LFSRcolor1[1338]);
    BiasedRNG[622] = (LFSRcolor1[802]&LFSRcolor1[399]&LFSRcolor1[1212]&LFSRcolor1[1115]);
    BiasedRNG[623] = (LFSRcolor1[1735]&LFSRcolor1[23]&LFSRcolor1[1694]&LFSRcolor1[518]);
    BiasedRNG[624] = (LFSRcolor1[1638]&LFSRcolor1[921]&LFSRcolor1[1463]&LFSRcolor1[920]);
    BiasedRNG[625] = (LFSRcolor1[1292]&LFSRcolor1[1322]&LFSRcolor1[417]&LFSRcolor1[335]);
    BiasedRNG[626] = (LFSRcolor1[500]&LFSRcolor1[1600]&LFSRcolor1[899]&LFSRcolor1[1567]);
    BiasedRNG[627] = (LFSRcolor1[295]&LFSRcolor1[1337]&LFSRcolor1[358]&LFSRcolor1[1662]);
    BiasedRNG[628] = (LFSRcolor1[826]&LFSRcolor1[569]&LFSRcolor1[1180]&LFSRcolor1[169]);
    BiasedRNG[629] = (LFSRcolor1[1173]&LFSRcolor1[234]&LFSRcolor1[1251]&LFSRcolor1[1310]);
    BiasedRNG[630] = (LFSRcolor1[1215]&LFSRcolor1[348]&LFSRcolor1[1619]&LFSRcolor1[0]);
    BiasedRNG[631] = (LFSRcolor1[945]&LFSRcolor1[713]&LFSRcolor1[10]&LFSRcolor1[1500]);
    BiasedRNG[632] = (LFSRcolor1[705]&LFSRcolor1[440]&LFSRcolor1[228]&LFSRcolor1[1565]);
    BiasedRNG[633] = (LFSRcolor1[38]&LFSRcolor1[227]&LFSRcolor1[435]&LFSRcolor1[1239]);
    BiasedRNG[634] = (LFSRcolor1[26]&LFSRcolor1[1687]&LFSRcolor1[30]&LFSRcolor1[618]);
    BiasedRNG[635] = (LFSRcolor1[530]&LFSRcolor1[1298]&LFSRcolor1[903]&LFSRcolor1[1431]);
    BiasedRNG[636] = (LFSRcolor1[1674]&LFSRcolor1[1131]&LFSRcolor1[1268]&LFSRcolor1[1306]);
    BiasedRNG[637] = (LFSRcolor1[1371]&LFSRcolor1[579]&LFSRcolor1[373]&LFSRcolor1[116]);
    BiasedRNG[638] = (LFSRcolor1[485]&LFSRcolor1[1657]&LFSRcolor1[1308]&LFSRcolor1[1410]);
    UnbiasedRNG[271] = LFSRcolor1[586];
    UnbiasedRNG[272] = LFSRcolor1[744];
    UnbiasedRNG[273] = LFSRcolor1[1336];
    UnbiasedRNG[274] = LFSRcolor1[1537];
    UnbiasedRNG[275] = LFSRcolor1[582];
    UnbiasedRNG[276] = LFSRcolor1[202];
    UnbiasedRNG[277] = LFSRcolor1[553];
    UnbiasedRNG[278] = LFSRcolor1[1703];
    UnbiasedRNG[279] = LFSRcolor1[722];
    UnbiasedRNG[280] = LFSRcolor1[700];
    UnbiasedRNG[281] = LFSRcolor1[1200];
    UnbiasedRNG[282] = LFSRcolor1[607];
    UnbiasedRNG[283] = LFSRcolor1[260];
    UnbiasedRNG[284] = LFSRcolor1[1435];
    UnbiasedRNG[285] = LFSRcolor1[304];
    UnbiasedRNG[286] = LFSRcolor1[930];
    UnbiasedRNG[287] = LFSRcolor1[893];
    UnbiasedRNG[288] = LFSRcolor1[737];
    UnbiasedRNG[289] = LFSRcolor1[1367];
    UnbiasedRNG[290] = LFSRcolor1[285];
    UnbiasedRNG[291] = LFSRcolor1[219];
    UnbiasedRNG[292] = LFSRcolor1[1789];
    UnbiasedRNG[293] = LFSRcolor1[432];
    UnbiasedRNG[294] = LFSRcolor1[412];
    UnbiasedRNG[295] = LFSRcolor1[1000];
    UnbiasedRNG[296] = LFSRcolor1[1759];
    UnbiasedRNG[297] = LFSRcolor1[546];
    UnbiasedRNG[298] = LFSRcolor1[552];
    UnbiasedRNG[299] = LFSRcolor1[244];
    UnbiasedRNG[300] = LFSRcolor1[418];
    UnbiasedRNG[301] = LFSRcolor1[1710];
    UnbiasedRNG[302] = LFSRcolor1[331];
    UnbiasedRNG[303] = LFSRcolor1[1466];
    UnbiasedRNG[304] = LFSRcolor1[322];
    UnbiasedRNG[305] = LFSRcolor1[117];
    UnbiasedRNG[306] = LFSRcolor1[257];
    UnbiasedRNG[307] = LFSRcolor1[648];
    UnbiasedRNG[308] = LFSRcolor1[852];
    UnbiasedRNG[309] = LFSRcolor1[1422];
    UnbiasedRNG[310] = LFSRcolor1[104];
    UnbiasedRNG[311] = LFSRcolor1[1712];
    UnbiasedRNG[312] = LFSRcolor1[1398];
    UnbiasedRNG[313] = LFSRcolor1[226];
    UnbiasedRNG[314] = LFSRcolor1[1373];
    UnbiasedRNG[315] = LFSRcolor1[369];
    UnbiasedRNG[316] = LFSRcolor1[250];
    UnbiasedRNG[317] = LFSRcolor1[1558];
    UnbiasedRNG[318] = LFSRcolor1[1436];
    UnbiasedRNG[319] = LFSRcolor1[1744];
    UnbiasedRNG[320] = LFSRcolor1[1469];
    UnbiasedRNG[321] = LFSRcolor1[980];
    UnbiasedRNG[322] = LFSRcolor1[915];
    UnbiasedRNG[323] = LFSRcolor1[1480];
    UnbiasedRNG[324] = LFSRcolor1[892];
    UnbiasedRNG[325] = LFSRcolor1[1204];
    UnbiasedRNG[326] = LFSRcolor1[221];
    UnbiasedRNG[327] = LFSRcolor1[1631];
    UnbiasedRNG[328] = LFSRcolor1[385];
    UnbiasedRNG[329] = LFSRcolor1[1734];
    UnbiasedRNG[330] = LFSRcolor1[1518];
    UnbiasedRNG[331] = LFSRcolor1[911];
    UnbiasedRNG[332] = LFSRcolor1[1342];
    UnbiasedRNG[333] = LFSRcolor1[1677];
    UnbiasedRNG[334] = LFSRcolor1[1170];
    UnbiasedRNG[335] = LFSRcolor1[1590];
    UnbiasedRNG[336] = LFSRcolor1[1669];
    UnbiasedRNG[337] = LFSRcolor1[1039];
    UnbiasedRNG[338] = LFSRcolor1[1572];
    UnbiasedRNG[339] = LFSRcolor1[837];
    UnbiasedRNG[340] = LFSRcolor1[1245];
    UnbiasedRNG[341] = LFSRcolor1[407];
    UnbiasedRNG[342] = LFSRcolor1[1012];
    UnbiasedRNG[343] = LFSRcolor1[386];
    UnbiasedRNG[344] = LFSRcolor1[1767];
    UnbiasedRNG[345] = LFSRcolor1[1240];
    UnbiasedRNG[346] = LFSRcolor1[968];
    UnbiasedRNG[347] = LFSRcolor1[839];
    UnbiasedRNG[348] = LFSRcolor1[212];
    UnbiasedRNG[349] = LFSRcolor1[24];
    UnbiasedRNG[350] = LFSRcolor1[1348];
    UnbiasedRNG[351] = LFSRcolor1[428];
    UnbiasedRNG[352] = LFSRcolor1[1545];
    UnbiasedRNG[353] = LFSRcolor1[1539];
    UnbiasedRNG[354] = LFSRcolor1[1159];
    UnbiasedRNG[355] = LFSRcolor1[1648];
    UnbiasedRNG[356] = LFSRcolor1[33];
    UnbiasedRNG[357] = LFSRcolor1[352];
    UnbiasedRNG[358] = LFSRcolor1[1718];
    UnbiasedRNG[359] = LFSRcolor1[747];
    UnbiasedRNG[360] = LFSRcolor1[738];
    UnbiasedRNG[361] = LFSRcolor1[448];
    UnbiasedRNG[362] = LFSRcolor1[540];
    UnbiasedRNG[363] = LFSRcolor1[1353];
    UnbiasedRNG[364] = LFSRcolor1[1329];
    UnbiasedRNG[365] = LFSRcolor1[136];
    UnbiasedRNG[366] = LFSRcolor1[1368];
    UnbiasedRNG[367] = LFSRcolor1[571];
    UnbiasedRNG[368] = LFSRcolor1[1201];
    UnbiasedRNG[369] = LFSRcolor1[320];
    UnbiasedRNG[370] = LFSRcolor1[794];
    UnbiasedRNG[371] = LFSRcolor1[1068];
    UnbiasedRNG[372] = LFSRcolor1[316];
    UnbiasedRNG[373] = LFSRcolor1[1228];
    UnbiasedRNG[374] = LFSRcolor1[384];
    UnbiasedRNG[375] = LFSRcolor1[849];
    UnbiasedRNG[376] = LFSRcolor1[856];
    UnbiasedRNG[377] = LFSRcolor1[1717];
    UnbiasedRNG[378] = LFSRcolor1[1633];
    UnbiasedRNG[379] = LFSRcolor1[948];
    UnbiasedRNG[380] = LFSRcolor1[1621];
    UnbiasedRNG[381] = LFSRcolor1[977];
    UnbiasedRNG[382] = LFSRcolor1[245];
    UnbiasedRNG[383] = LFSRcolor1[1511];
    UnbiasedRNG[384] = LFSRcolor1[1132];
    UnbiasedRNG[385] = LFSRcolor1[243];
    UnbiasedRNG[386] = LFSRcolor1[769];
    UnbiasedRNG[387] = LFSRcolor1[520];
    UnbiasedRNG[388] = LFSRcolor1[767];
    UnbiasedRNG[389] = LFSRcolor1[748];
    UnbiasedRNG[390] = LFSRcolor1[1331];
    UnbiasedRNG[391] = LFSRcolor1[89];
    UnbiasedRNG[392] = LFSRcolor1[1232];
    UnbiasedRNG[393] = LFSRcolor1[1208];
    UnbiasedRNG[394] = LFSRcolor1[367];
    UnbiasedRNG[395] = LFSRcolor1[1116];
    UnbiasedRNG[396] = LFSRcolor1[1540];
    UnbiasedRNG[397] = LFSRcolor1[1006];
    UnbiasedRNG[398] = LFSRcolor1[851];
    UnbiasedRNG[399] = LFSRcolor1[381];
    UnbiasedRNG[400] = LFSRcolor1[753];
    UnbiasedRNG[401] = LFSRcolor1[1554];
    UnbiasedRNG[402] = LFSRcolor1[1042];
    UnbiasedRNG[403] = LFSRcolor1[97];
    UnbiasedRNG[404] = LFSRcolor1[344];
    UnbiasedRNG[405] = LFSRcolor1[1526];
    UnbiasedRNG[406] = LFSRcolor1[731];
    UnbiasedRNG[407] = LFSRcolor1[1269];
    UnbiasedRNG[408] = LFSRcolor1[1783];
    UnbiasedRNG[409] = LFSRcolor1[1026];
    UnbiasedRNG[410] = LFSRcolor1[1644];
    UnbiasedRNG[411] = LFSRcolor1[1686];
    UnbiasedRNG[412] = LFSRcolor1[1037];
    UnbiasedRNG[413] = LFSRcolor1[1154];
    UnbiasedRNG[414] = LFSRcolor1[1667];
    UnbiasedRNG[415] = LFSRcolor1[516];
    UnbiasedRNG[416] = LFSRcolor1[1205];
    UnbiasedRNG[417] = LFSRcolor1[749];
    UnbiasedRNG[418] = LFSRcolor1[719];
    UnbiasedRNG[419] = LFSRcolor1[382];
    UnbiasedRNG[420] = LFSRcolor1[549];
    UnbiasedRNG[421] = LFSRcolor1[645];
    UnbiasedRNG[422] = LFSRcolor1[1752];
    UnbiasedRNG[423] = LFSRcolor1[978];
    UnbiasedRNG[424] = LFSRcolor1[60];
    UnbiasedRNG[425] = LFSRcolor1[1072];
    UnbiasedRNG[426] = LFSRcolor1[857];
    UnbiasedRNG[427] = LFSRcolor1[1366];
    UnbiasedRNG[428] = LFSRcolor1[1189];
    UnbiasedRNG[429] = LFSRcolor1[863];
    UnbiasedRNG[430] = LFSRcolor1[110];
    UnbiasedRNG[431] = LFSRcolor1[1318];
    UnbiasedRNG[432] = LFSRcolor1[926];
    UnbiasedRNG[433] = LFSRcolor1[1607];
    UnbiasedRNG[434] = LFSRcolor1[595];
    UnbiasedRNG[435] = LFSRcolor1[152];
    UnbiasedRNG[436] = LFSRcolor1[1372];
    UnbiasedRNG[437] = LFSRcolor1[887];
    UnbiasedRNG[438] = LFSRcolor1[1295];
    UnbiasedRNG[439] = LFSRcolor1[314];
    UnbiasedRNG[440] = LFSRcolor1[1086];
    UnbiasedRNG[441] = LFSRcolor1[941];
    UnbiasedRNG[442] = LFSRcolor1[614];
    UnbiasedRNG[443] = LFSRcolor1[766];
    UnbiasedRNG[444] = LFSRcolor1[1472];
    UnbiasedRNG[445] = LFSRcolor1[269];
    UnbiasedRNG[446] = LFSRcolor1[1432];
    UnbiasedRNG[447] = LFSRcolor1[11];
    UnbiasedRNG[448] = LFSRcolor1[1618];
    UnbiasedRNG[449] = LFSRcolor1[781];
    UnbiasedRNG[450] = LFSRcolor1[598];
    UnbiasedRNG[451] = LFSRcolor1[286];
    UnbiasedRNG[452] = LFSRcolor1[1581];
    UnbiasedRNG[453] = LFSRcolor1[880];
    UnbiasedRNG[454] = LFSRcolor1[1172];
    UnbiasedRNG[455] = LFSRcolor1[649];
    UnbiasedRNG[456] = LFSRcolor1[1335];
    UnbiasedRNG[457] = LFSRcolor1[996];
    UnbiasedRNG[458] = LFSRcolor1[1503];
    UnbiasedRNG[459] = LFSRcolor1[964];
    UnbiasedRNG[460] = LFSRcolor1[1569];
    UnbiasedRNG[461] = LFSRcolor1[368];
    UnbiasedRNG[462] = LFSRcolor1[1165];
    UnbiasedRNG[463] = LFSRcolor1[1536];
    UnbiasedRNG[464] = LFSRcolor1[143];
    UnbiasedRNG[465] = LFSRcolor1[745];
    UnbiasedRNG[466] = LFSRcolor1[524];
    UnbiasedRNG[467] = LFSRcolor1[800];
    UnbiasedRNG[468] = LFSRcolor1[249];
    UnbiasedRNG[469] = LFSRcolor1[561];
    UnbiasedRNG[470] = LFSRcolor1[259];
    UnbiasedRNG[471] = LFSRcolor1[1258];
    UnbiasedRNG[472] = LFSRcolor1[274];
    UnbiasedRNG[473] = LFSRcolor1[52];
    UnbiasedRNG[474] = LFSRcolor1[1465];
    UnbiasedRNG[475] = LFSRcolor1[613];
    UnbiasedRNG[476] = LFSRcolor1[1760];
    UnbiasedRNG[477] = LFSRcolor1[1499];
    UnbiasedRNG[478] = LFSRcolor1[1105];
    UnbiasedRNG[479] = LFSRcolor1[149];
    UnbiasedRNG[480] = LFSRcolor1[467];
    UnbiasedRNG[481] = LFSRcolor1[1374];
    UnbiasedRNG[482] = LFSRcolor1[1003];
    UnbiasedRNG[483] = LFSRcolor1[394];
    UnbiasedRNG[484] = LFSRcolor1[774];
    UnbiasedRNG[485] = LFSRcolor1[1021];
    UnbiasedRNG[486] = LFSRcolor1[678];
    UnbiasedRNG[487] = LFSRcolor1[272];
    UnbiasedRNG[488] = LFSRcolor1[824];
    UnbiasedRNG[489] = LFSRcolor1[469];
    UnbiasedRNG[490] = LFSRcolor1[577];
    UnbiasedRNG[491] = LFSRcolor1[1119];
    UnbiasedRNG[492] = LFSRcolor1[1497];
    UnbiasedRNG[493] = LFSRcolor1[1396];
    UnbiasedRNG[494] = LFSRcolor1[1447];
    UnbiasedRNG[495] = LFSRcolor1[730];
end

always @(posedge color1_clk) begin
    BiasedRNG[639] = (LFSRcolor2[1175]&LFSRcolor2[1110]&LFSRcolor2[627]&LFSRcolor2[833]);
    BiasedRNG[640] = (LFSRcolor2[197]&LFSRcolor2[805]&LFSRcolor2[385]&LFSRcolor2[1250]);
    BiasedRNG[641] = (LFSRcolor2[354]&LFSRcolor2[50]&LFSRcolor2[167]&LFSRcolor2[911]);
    BiasedRNG[642] = (LFSRcolor2[411]&LFSRcolor2[1132]&LFSRcolor2[362]&LFSRcolor2[307]);
    BiasedRNG[643] = (LFSRcolor2[449]&LFSRcolor2[583]&LFSRcolor2[782]&LFSRcolor2[978]);
    BiasedRNG[644] = (LFSRcolor2[318]&LFSRcolor2[301]&LFSRcolor2[421]&LFSRcolor2[161]);
    BiasedRNG[645] = (LFSRcolor2[1249]&LFSRcolor2[539]&LFSRcolor2[586]&LFSRcolor2[595]);
    BiasedRNG[646] = (LFSRcolor2[210]&LFSRcolor2[1059]&LFSRcolor2[728]&LFSRcolor2[196]);
    BiasedRNG[647] = (LFSRcolor2[156]&LFSRcolor2[419]&LFSRcolor2[729]&LFSRcolor2[1042]);
    BiasedRNG[648] = (LFSRcolor2[64]&LFSRcolor2[256]&LFSRcolor2[683]&LFSRcolor2[479]);
    BiasedRNG[649] = (LFSRcolor2[828]&LFSRcolor2[1053]&LFSRcolor2[46]&LFSRcolor2[959]);
    BiasedRNG[650] = (LFSRcolor2[15]&LFSRcolor2[731]&LFSRcolor2[206]&LFSRcolor2[192]);
    BiasedRNG[651] = (LFSRcolor2[618]&LFSRcolor2[773]&LFSRcolor2[1035]&LFSRcolor2[893]);
    BiasedRNG[652] = (LFSRcolor2[662]&LFSRcolor2[455]&LFSRcolor2[43]&LFSRcolor2[151]);
    BiasedRNG[653] = (LFSRcolor2[1199]&LFSRcolor2[1234]&LFSRcolor2[358]&LFSRcolor2[425]);
    BiasedRNG[654] = (LFSRcolor2[520]&LFSRcolor2[483]&LFSRcolor2[100]&LFSRcolor2[1099]);
    BiasedRNG[655] = (LFSRcolor2[562]&LFSRcolor2[293]&LFSRcolor2[235]&LFSRcolor2[656]);
    BiasedRNG[656] = (LFSRcolor2[839]&LFSRcolor2[604]&LFSRcolor2[84]&LFSRcolor2[56]);
    BiasedRNG[657] = (LFSRcolor2[277]&LFSRcolor2[970]&LFSRcolor2[719]&LFSRcolor2[1131]);
    BiasedRNG[658] = (LFSRcolor2[767]&LFSRcolor2[780]&LFSRcolor2[446]&LFSRcolor2[1260]);
    BiasedRNG[659] = (LFSRcolor2[681]&LFSRcolor2[493]&LFSRcolor2[1101]&LFSRcolor2[1102]);
    BiasedRNG[660] = (LFSRcolor2[749]&LFSRcolor2[874]&LFSRcolor2[311]&LFSRcolor2[772]);
    BiasedRNG[661] = (LFSRcolor2[159]&LFSRcolor2[1082]&LFSRcolor2[559]&LFSRcolor2[689]);
    BiasedRNG[662] = (LFSRcolor2[120]&LFSRcolor2[879]&LFSRcolor2[185]&LFSRcolor2[1067]);
    BiasedRNG[663] = (LFSRcolor2[32]&LFSRcolor2[848]&LFSRcolor2[612]&LFSRcolor2[245]);
    BiasedRNG[664] = (LFSRcolor2[330]&LFSRcolor2[867]&LFSRcolor2[889]&LFSRcolor2[510]);
    BiasedRNG[665] = (LFSRcolor2[1213]&LFSRcolor2[601]&LFSRcolor2[300]&LFSRcolor2[506]);
    BiasedRNG[666] = (LFSRcolor2[613]&LFSRcolor2[608]&LFSRcolor2[1052]&LFSRcolor2[57]);
    BiasedRNG[667] = (LFSRcolor2[1159]&LFSRcolor2[993]&LFSRcolor2[1272]&LFSRcolor2[1214]);
    BiasedRNG[668] = (LFSRcolor2[966]&LFSRcolor2[1275]&LFSRcolor2[576]&LFSRcolor2[588]);
    BiasedRNG[669] = (LFSRcolor2[1073]&LFSRcolor2[1142]&LFSRcolor2[958]&LFSRcolor2[1271]);
    BiasedRNG[670] = (LFSRcolor2[814]&LFSRcolor2[1242]&LFSRcolor2[883]&LFSRcolor2[896]);
    BiasedRNG[671] = (LFSRcolor2[325]&LFSRcolor2[1243]&LFSRcolor2[1174]&LFSRcolor2[974]);
    BiasedRNG[672] = (LFSRcolor2[873]&LFSRcolor2[438]&LFSRcolor2[653]&LFSRcolor2[254]);
    BiasedRNG[673] = (LFSRcolor2[442]&LFSRcolor2[427]&LFSRcolor2[226]&LFSRcolor2[503]);
    BiasedRNG[674] = (LFSRcolor2[1138]&LFSRcolor2[452]&LFSRcolor2[847]&LFSRcolor2[1049]);
    BiasedRNG[675] = (LFSRcolor2[363]&LFSRcolor2[1098]&LFSRcolor2[834]&LFSRcolor2[775]);
    BiasedRNG[676] = (LFSRcolor2[920]&LFSRcolor2[276]&LFSRcolor2[851]&LFSRcolor2[1133]);
    BiasedRNG[677] = (LFSRcolor2[759]&LFSRcolor2[285]&LFSRcolor2[956]&LFSRcolor2[10]);
    BiasedRNG[678] = (LFSRcolor2[1125]&LFSRcolor2[263]&LFSRcolor2[85]&LFSRcolor2[81]);
    BiasedRNG[679] = (LFSRcolor2[718]&LFSRcolor2[399]&LFSRcolor2[1165]&LFSRcolor2[30]);
    BiasedRNG[680] = (LFSRcolor2[1156]&LFSRcolor2[371]&LFSRcolor2[615]&LFSRcolor2[1072]);
    BiasedRNG[681] = (LFSRcolor2[690]&LFSRcolor2[467]&LFSRcolor2[141]&LFSRcolor2[323]);
    BiasedRNG[682] = (LFSRcolor2[1149]&LFSRcolor2[1157]&LFSRcolor2[435]&LFSRcolor2[216]);
    BiasedRNG[683] = (LFSRcolor2[727]&LFSRcolor2[591]&LFSRcolor2[529]&LFSRcolor2[526]);
    BiasedRNG[684] = (LFSRcolor2[175]&LFSRcolor2[725]&LFSRcolor2[995]&LFSRcolor2[496]);
    BiasedRNG[685] = (LFSRcolor2[969]&LFSRcolor2[1160]&LFSRcolor2[976]&LFSRcolor2[297]);
    BiasedRNG[686] = (LFSRcolor2[1254]&LFSRcolor2[800]&LFSRcolor2[132]&LFSRcolor2[204]);
    BiasedRNG[687] = (LFSRcolor2[439]&LFSRcolor2[762]&LFSRcolor2[1038]&LFSRcolor2[855]);
    BiasedRNG[688] = (LFSRcolor2[716]&LFSRcolor2[1218]&LFSRcolor2[31]&LFSRcolor2[74]);
    BiasedRNG[689] = (LFSRcolor2[941]&LFSRcolor2[985]&LFSRcolor2[696]&LFSRcolor2[975]);
    BiasedRNG[690] = (LFSRcolor2[447]&LFSRcolor2[157]&LFSRcolor2[625]&LFSRcolor2[545]);
    BiasedRNG[691] = (LFSRcolor2[1189]&LFSRcolor2[269]&LFSRcolor2[426]&LFSRcolor2[791]);
    BiasedRNG[692] = (LFSRcolor2[471]&LFSRcolor2[1029]&LFSRcolor2[919]&LFSRcolor2[594]);
    BiasedRNG[693] = (LFSRcolor2[1139]&LFSRcolor2[304]&LFSRcolor2[650]&LFSRcolor2[553]);
    BiasedRNG[694] = (LFSRcolor2[955]&LFSRcolor2[459]&LFSRcolor2[55]&LFSRcolor2[367]);
    BiasedRNG[695] = (LFSRcolor2[628]&LFSRcolor2[39]&LFSRcolor2[774]&LFSRcolor2[133]);
    BiasedRNG[696] = (LFSRcolor2[864]&LFSRcolor2[850]&LFSRcolor2[95]&LFSRcolor2[1155]);
    BiasedRNG[697] = (LFSRcolor2[918]&LFSRcolor2[785]&LFSRcolor2[434]&LFSRcolor2[1060]);
    BiasedRNG[698] = (LFSRcolor2[870]&LFSRcolor2[581]&LFSRcolor2[306]&LFSRcolor2[1066]);
    BiasedRNG[699] = (LFSRcolor2[756]&LFSRcolor2[199]&LFSRcolor2[1032]&LFSRcolor2[887]);
    BiasedRNG[700] = (LFSRcolor2[417]&LFSRcolor2[1203]&LFSRcolor2[209]&LFSRcolor2[266]);
    BiasedRNG[701] = (LFSRcolor2[1144]&LFSRcolor2[212]&LFSRcolor2[538]&LFSRcolor2[303]);
    BiasedRNG[702] = (LFSRcolor2[465]&LFSRcolor2[1166]&LFSRcolor2[954]&LFSRcolor2[910]);
    BiasedRNG[703] = (LFSRcolor2[28]&LFSRcolor2[368]&LFSRcolor2[645]&LFSRcolor2[784]);
    BiasedRNG[704] = (LFSRcolor2[657]&LFSRcolor2[579]&LFSRcolor2[220]&LFSRcolor2[965]);
    BiasedRNG[705] = (LFSRcolor2[374]&LFSRcolor2[207]&LFSRcolor2[807]&LFSRcolor2[20]);
    BiasedRNG[706] = (LFSRcolor2[332]&LFSRcolor2[977]&LFSRcolor2[1173]&LFSRcolor2[160]);
    BiasedRNG[707] = (LFSRcolor2[355]&LFSRcolor2[981]&LFSRcolor2[68]&LFSRcolor2[692]);
    BiasedRNG[708] = (LFSRcolor2[989]&LFSRcolor2[183]&LFSRcolor2[1248]&LFSRcolor2[1253]);
    BiasedRNG[709] = (LFSRcolor2[916]&LFSRcolor2[1143]&LFSRcolor2[428]&LFSRcolor2[139]);
    BiasedRNG[710] = (LFSRcolor2[1216]&LFSRcolor2[992]&LFSRcolor2[1020]&LFSRcolor2[166]);
    BiasedRNG[711] = (LFSRcolor2[878]&LFSRcolor2[1071]&LFSRcolor2[1235]&LFSRcolor2[131]);
    BiasedRNG[712] = (LFSRcolor2[97]&LFSRcolor2[513]&LFSRcolor2[1074]&LFSRcolor2[1113]);
    BiasedRNG[713] = (LFSRcolor2[240]&LFSRcolor2[638]&LFSRcolor2[616]&LFSRcolor2[248]);
    BiasedRNG[714] = (LFSRcolor2[934]&LFSRcolor2[302]&LFSRcolor2[611]&LFSRcolor2[605]);
    BiasedRNG[715] = (LFSRcolor2[478]&LFSRcolor2[331]&LFSRcolor2[580]&LFSRcolor2[232]);
    BiasedRNG[716] = (LFSRcolor2[988]&LFSRcolor2[633]&LFSRcolor2[474]&LFSRcolor2[24]);
    BiasedRNG[717] = (LFSRcolor2[624]&LFSRcolor2[554]&LFSRcolor2[821]&LFSRcolor2[685]);
    BiasedRNG[718] = (LFSRcolor2[723]&LFSRcolor2[1036]&LFSRcolor2[922]&LFSRcolor2[700]);
    BiasedRNG[719] = (LFSRcolor2[983]&LFSRcolor2[812]&LFSRcolor2[825]&LFSRcolor2[602]);
    BiasedRNG[720] = (LFSRcolor2[518]&LFSRcolor2[877]&LFSRcolor2[83]&LFSRcolor2[1280]);
    BiasedRNG[721] = (LFSRcolor2[1107]&LFSRcolor2[103]&LFSRcolor2[708]&LFSRcolor2[1024]);
    BiasedRNG[722] = (LFSRcolor2[392]&LFSRcolor2[322]&LFSRcolor2[171]&LFSRcolor2[957]);
    BiasedRNG[723] = (LFSRcolor2[1191]&LFSRcolor2[40]&LFSRcolor2[463]&LFSRcolor2[675]);
    BiasedRNG[724] = (LFSRcolor2[908]&LFSRcolor2[8]&LFSRcolor2[1092]&LFSRcolor2[69]);
    BiasedRNG[725] = (LFSRcolor2[1037]&LFSRcolor2[1122]&LFSRcolor2[566]&LFSRcolor2[714]);
    BiasedRNG[726] = (LFSRcolor2[54]&LFSRcolor2[1120]&LFSRcolor2[316]&LFSRcolor2[203]);
    BiasedRNG[727] = (LFSRcolor2[664]&LFSRcolor2[128]&LFSRcolor2[1180]&LFSRcolor2[164]);
    BiasedRNG[728] = (LFSRcolor2[414]&LFSRcolor2[257]&LFSRcolor2[511]&LFSRcolor2[1231]);
    BiasedRNG[729] = (LFSRcolor2[1169]&LFSRcolor2[1207]&LFSRcolor2[211]&LFSRcolor2[963]);
    BiasedRNG[730] = (LFSRcolor2[1255]&LFSRcolor2[231]&LFSRcolor2[949]&LFSRcolor2[72]);
    BiasedRNG[731] = (LFSRcolor2[541]&LFSRcolor2[505]&LFSRcolor2[241]&LFSRcolor2[748]);
    BiasedRNG[732] = (LFSRcolor2[516]&LFSRcolor2[17]&LFSRcolor2[461]&LFSRcolor2[1278]);
    BiasedRNG[733] = (LFSRcolor2[726]&LFSRcolor2[1028]&LFSRcolor2[906]&LFSRcolor2[381]);
    BiasedRNG[734] = (LFSRcolor2[1018]&LFSRcolor2[366]&LFSRcolor2[1274]&LFSRcolor2[398]);
    BiasedRNG[735] = (LFSRcolor2[663]&LFSRcolor2[676]&LFSRcolor2[1094]&LFSRcolor2[945]);
    BiasedRNG[736] = (LFSRcolor2[1246]&LFSRcolor2[630]&LFSRcolor2[309]&LFSRcolor2[312]);
    BiasedRNG[737] = (LFSRcolor2[942]&LFSRcolor2[1033]&LFSRcolor2[1109]&LFSRcolor2[902]);
    BiasedRNG[738] = (LFSRcolor2[482]&LFSRcolor2[1261]&LFSRcolor2[107]&LFSRcolor2[557]);
    BiasedRNG[739] = (LFSRcolor2[1006]&LFSRcolor2[946]&LFSRcolor2[710]&LFSRcolor2[243]);
    BiasedRNG[740] = (LFSRcolor2[512]&LFSRcolor2[349]&LFSRcolor2[578]&LFSRcolor2[432]);
    BiasedRNG[741] = (LFSRcolor2[1239]&LFSRcolor2[213]&LFSRcolor2[409]&LFSRcolor2[750]);
    BiasedRNG[742] = (LFSRcolor2[693]&LFSRcolor2[904]&LFSRcolor2[1123]&LFSRcolor2[238]);
    BiasedRNG[743] = (LFSRcolor2[440]&LFSRcolor2[950]&LFSRcolor2[666]&LFSRcolor2[1140]);
    BiasedRNG[744] = (LFSRcolor2[181]&LFSRcolor2[990]&LFSRcolor2[1075]&LFSRcolor2[561]);
    BiasedRNG[745] = (LFSRcolor2[1034]&LFSRcolor2[777]&LFSRcolor2[261]&LFSRcolor2[781]);
    BiasedRNG[746] = (LFSRcolor2[619]&LFSRcolor2[629]&LFSRcolor2[912]&LFSRcolor2[565]);
    BiasedRNG[747] = (LFSRcolor2[917]&LFSRcolor2[191]&LFSRcolor2[822]&LFSRcolor2[960]);
    BiasedRNG[748] = (LFSRcolor2[694]&LFSRcolor2[907]&LFSRcolor2[356]&LFSRcolor2[1056]);
    BiasedRNG[749] = (LFSRcolor2[1198]&LFSRcolor2[999]&LFSRcolor2[1057]&LFSRcolor2[44]);
    BiasedRNG[750] = (LFSRcolor2[386]&LFSRcolor2[485]&LFSRcolor2[458]&LFSRcolor2[473]);
    BiasedRNG[751] = (LFSRcolor2[445]&LFSRcolor2[1116]&LFSRcolor2[674]&LFSRcolor2[658]);
    BiasedRNG[752] = (LFSRcolor2[888]&LFSRcolor2[603]&LFSRcolor2[222]&LFSRcolor2[1091]);
    BiasedRNG[753] = (LFSRcolor2[1114]&LFSRcolor2[1043]&LFSRcolor2[375]&LFSRcolor2[393]);
    BiasedRNG[754] = (LFSRcolor2[838]&LFSRcolor2[4]&LFSRcolor2[486]&LFSRcolor2[1085]);
    BiasedRNG[755] = (LFSRcolor2[1217]&LFSRcolor2[536]&LFSRcolor2[378]&LFSRcolor2[1244]);
    BiasedRNG[756] = (LFSRcolor2[1230]&LFSRcolor2[333]&LFSRcolor2[670]&LFSRcolor2[407]);
    BiasedRNG[757] = (LFSRcolor2[1023]&LFSRcolor2[1130]&LFSRcolor2[687]&LFSRcolor2[188]);
    BiasedRNG[758] = (LFSRcolor2[1093]&LFSRcolor2[34]&LFSRcolor2[1224]&LFSRcolor2[424]);
    BiasedRNG[759] = (LFSRcolor2[453]&LFSRcolor2[768]&LFSRcolor2[487]&LFSRcolor2[475]);
    BiasedRNG[760] = (LFSRcolor2[412]&LFSRcolor2[765]&LFSRcolor2[163]&LFSRcolor2[1177]);
    BiasedRNG[761] = (LFSRcolor2[678]&LFSRcolor2[1025]&LFSRcolor2[1058]&LFSRcolor2[1245]);
    BiasedRNG[762] = (LFSRcolor2[1204]&LFSRcolor2[1237]&LFSRcolor2[94]&LFSRcolor2[75]);
    BiasedRNG[763] = (LFSRcolor2[802]&LFSRcolor2[489]&LFSRcolor2[430]&LFSRcolor2[18]);
    BiasedRNG[764] = (LFSRcolor2[270]&LFSRcolor2[158]&LFSRcolor2[469]&LFSRcolor2[326]);
    BiasedRNG[765] = (LFSRcolor2[149]&LFSRcolor2[590]&LFSRcolor2[609]&LFSRcolor2[353]);
    BiasedRNG[766] = (LFSRcolor2[147]&LFSRcolor2[679]&LFSRcolor2[972]&LFSRcolor2[868]);
    BiasedRNG[767] = (LFSRcolor2[413]&LFSRcolor2[672]&LFSRcolor2[940]&LFSRcolor2[875]);
    BiasedRNG[768] = (LFSRcolor2[1076]&LFSRcolor2[1027]&LFSRcolor2[1196]&LFSRcolor2[707]);
    BiasedRNG[769] = (LFSRcolor2[1048]&LFSRcolor2[234]&LFSRcolor2[262]&LFSRcolor2[253]);
    BiasedRNG[770] = (LFSRcolor2[6]&LFSRcolor2[876]&LFSRcolor2[556]&LFSRcolor2[964]);
    BiasedRNG[771] = (LFSRcolor2[218]&LFSRcolor2[1087]&LFSRcolor2[314]&LFSRcolor2[1268]);
    BiasedRNG[772] = (LFSRcolor2[109]&LFSRcolor2[1229]&LFSRcolor2[587]&LFSRcolor2[1262]);
    BiasedRNG[773] = (LFSRcolor2[1287]&LFSRcolor2[1267]&LFSRcolor2[747]&LFSRcolor2[620]);
    BiasedRNG[774] = (LFSRcolor2[639]&LFSRcolor2[494]&LFSRcolor2[1005]&LFSRcolor2[490]);
    BiasedRNG[775] = (LFSRcolor2[1031]&LFSRcolor2[859]&LFSRcolor2[315]&LFSRcolor2[1004]);
    BiasedRNG[776] = (LFSRcolor2[324]&LFSRcolor2[384]&LFSRcolor2[1070]&LFSRcolor2[610]);
    BiasedRNG[777] = (LFSRcolor2[264]&LFSRcolor2[251]&LFSRcolor2[2]&LFSRcolor2[382]);
    BiasedRNG[778] = (LFSRcolor2[239]&LFSRcolor2[845]&LFSRcolor2[110]&LFSRcolor2[67]);
    BiasedRNG[779] = (LFSRcolor2[933]&LFSRcolor2[659]&LFSRcolor2[655]&LFSRcolor2[1182]);
    BiasedRNG[780] = (LFSRcolor2[810]&LFSRcolor2[668]&LFSRcolor2[346]&LFSRcolor2[36]);
    BiasedRNG[781] = (LFSRcolor2[745]&LFSRcolor2[1021]&LFSRcolor2[201]&LFSRcolor2[574]);
    BiasedRNG[782] = (LFSRcolor2[287]&LFSRcolor2[737]&LFSRcolor2[905]&LFSRcolor2[236]);
    BiasedRNG[783] = (LFSRcolor2[186]&LFSRcolor2[1201]&LFSRcolor2[947]&LFSRcolor2[636]);
    BiasedRNG[784] = (LFSRcolor2[600]&LFSRcolor2[1014]&LFSRcolor2[152]&LFSRcolor2[524]);
    BiasedRNG[785] = (LFSRcolor2[189]&LFSRcolor2[892]&LFSRcolor2[472]&LFSRcolor2[273]);
    BiasedRNG[786] = (LFSRcolor2[373]&LFSRcolor2[401]&LFSRcolor2[1178]&LFSRcolor2[460]);
    BiasedRNG[787] = (LFSRcolor2[813]&LFSRcolor2[7]&LFSRcolor2[1270]&LFSRcolor2[746]);
    BiasedRNG[788] = (LFSRcolor2[1247]&LFSRcolor2[1127]&LFSRcolor2[347]&LFSRcolor2[779]);
    BiasedRNG[789] = (LFSRcolor2[1062]&LFSRcolor2[1000]&LFSRcolor2[134]&LFSRcolor2[415]);
    BiasedRNG[790] = (LFSRcolor2[684]&LFSRcolor2[14]&LFSRcolor2[1016]&LFSRcolor2[555]);
    BiasedRNG[791] = (LFSRcolor2[11]&LFSRcolor2[359]&LFSRcolor2[1045]&LFSRcolor2[820]);
    BiasedRNG[792] = (LFSRcolor2[247]&LFSRcolor2[70]&LFSRcolor2[626]&LFSRcolor2[89]);
    BiasedRNG[793] = (LFSRcolor2[860]&LFSRcolor2[1212]&LFSRcolor2[734]&LFSRcolor2[643]);
    BiasedRNG[794] = (LFSRcolor2[351]&LFSRcolor2[1170]&LFSRcolor2[1022]&LFSRcolor2[1080]);
    BiasedRNG[795] = (LFSRcolor2[1054]&LFSRcolor2[205]&LFSRcolor2[935]&LFSRcolor2[1118]);
    BiasedRNG[796] = (LFSRcolor2[1001]&LFSRcolor2[766]&LFSRcolor2[631]&LFSRcolor2[344]);
    BiasedRNG[797] = (LFSRcolor2[289]&LFSRcolor2[715]&LFSRcolor2[436]&LFSRcolor2[923]);
    BiasedRNG[798] = (LFSRcolor2[114]&LFSRcolor2[1010]&LFSRcolor2[1226]&LFSRcolor2[1129]);
    BiasedRNG[799] = (LFSRcolor2[170]&LFSRcolor2[504]&LFSRcolor2[65]&LFSRcolor2[388]);
    BiasedRNG[800] = (LFSRcolor2[1269]&LFSRcolor2[63]&LFSRcolor2[376]&LFSRcolor2[104]);
    BiasedRNG[801] = (LFSRcolor2[948]&LFSRcolor2[1104]&LFSRcolor2[927]&LFSRcolor2[682]);
    BiasedRNG[802] = (LFSRcolor2[431]&LFSRcolor2[836]&LFSRcolor2[35]&LFSRcolor2[319]);
    BiasedRNG[803] = (LFSRcolor2[732]&LFSRcolor2[1068]&LFSRcolor2[930]&LFSRcolor2[1220]);
    BiasedRNG[804] = (LFSRcolor2[703]&LFSRcolor2[1179]&LFSRcolor2[770]&LFSRcolor2[394]);
    BiasedRNG[805] = (LFSRcolor2[327]&LFSRcolor2[408]&LFSRcolor2[1090]&LFSRcolor2[743]);
    BiasedRNG[806] = (LFSRcolor2[533]&LFSRcolor2[404]&LFSRcolor2[1282]&LFSRcolor2[909]);
    BiasedRNG[807] = (LFSRcolor2[162]&LFSRcolor2[597]&LFSRcolor2[647]&LFSRcolor2[1009]);
    BiasedRNG[808] = (LFSRcolor2[369]&LFSRcolor2[361]&LFSRcolor2[507]&LFSRcolor2[313]);
    BiasedRNG[809] = (LFSRcolor2[991]&LFSRcolor2[937]&LFSRcolor2[924]&LFSRcolor2[865]);
    BiasedRNG[810] = (LFSRcolor2[429]&LFSRcolor2[1097]&LFSRcolor2[763]&LFSRcolor2[570]);
    BiasedRNG[811] = (LFSRcolor2[758]&LFSRcolor2[819]&LFSRcolor2[798]&LFSRcolor2[736]);
    BiasedRNG[812] = (LFSRcolor2[1095]&LFSRcolor2[644]&LFSRcolor2[811]&LFSRcolor2[788]);
    BiasedRNG[813] = (LFSRcolor2[418]&LFSRcolor2[1188]&LFSRcolor2[1017]&LFSRcolor2[560]);
    BiasedRNG[814] = (LFSRcolor2[502]&LFSRcolor2[1086]&LFSRcolor2[783]&LFSRcolor2[722]);
    BiasedRNG[815] = (LFSRcolor2[654]&LFSRcolor2[195]&LFSRcolor2[126]&LFSRcolor2[115]);
    BiasedRNG[816] = (LFSRcolor2[1121]&LFSRcolor2[577]&LFSRcolor2[21]&LFSRcolor2[1257]);
    BiasedRNG[817] = (LFSRcolor2[1141]&LFSRcolor2[1084]&LFSRcolor2[568]&LFSRcolor2[898]);
    BiasedRNG[818] = (LFSRcolor2[290]&LFSRcolor2[477]&LFSRcolor2[897]&LFSRcolor2[66]);
    BiasedRNG[819] = (LFSRcolor2[457]&LFSRcolor2[793]&LFSRcolor2[340]&LFSRcolor2[416]);
    BiasedRNG[820] = (LFSRcolor2[1222]&LFSRcolor2[823]&LFSRcolor2[441]&LFSRcolor2[336]);
    BiasedRNG[821] = (LFSRcolor2[771]&LFSRcolor2[444]&LFSRcolor2[776]&LFSRcolor2[379]);
    BiasedRNG[822] = (LFSRcolor2[58]&LFSRcolor2[174]&LFSRcolor2[968]&LFSRcolor2[829]);
    BiasedRNG[823] = (LFSRcolor2[334]&LFSRcolor2[422]&LFSRcolor2[830]&LFSRcolor2[1153]);
    BiasedRNG[824] = (LFSRcolor2[899]&LFSRcolor2[172]&LFSRcolor2[468]&LFSRcolor2[1200]);
    BiasedRNG[825] = (LFSRcolor2[614]&LFSRcolor2[1251]&LFSRcolor2[741]&LFSRcolor2[1167]);
    BiasedRNG[826] = (LFSRcolor2[1223]&LFSRcolor2[721]&LFSRcolor2[1]&LFSRcolor2[547]);
    BiasedRNG[827] = (LFSRcolor2[826]&LFSRcolor2[343]&LFSRcolor2[671]&LFSRcolor2[1111]);
    BiasedRNG[828] = (LFSRcolor2[395]&LFSRcolor2[106]&LFSRcolor2[136]&LFSRcolor2[928]);
    BiasedRNG[829] = (LFSRcolor2[1003]&LFSRcolor2[320]&LFSRcolor2[789]&LFSRcolor2[1100]);
    BiasedRNG[830] = (LFSRcolor2[522]&LFSRcolor2[962]&LFSRcolor2[660]&LFSRcolor2[1026]);
    BiasedRNG[831] = (LFSRcolor2[1146]&LFSRcolor2[317]&LFSRcolor2[1194]&LFSRcolor2[1186]);
    BiasedRNG[832] = (LFSRcolor2[1013]&LFSRcolor2[786]&LFSRcolor2[1208]&LFSRcolor2[1030]);
    BiasedRNG[833] = (LFSRcolor2[295]&LFSRcolor2[842]&LFSRcolor2[515]&LFSRcolor2[1206]);
    BiasedRNG[834] = (LFSRcolor2[462]&LFSRcolor2[1050]&LFSRcolor2[79]&LFSRcolor2[1233]);
    BiasedRNG[835] = (LFSRcolor2[352]&LFSRcolor2[1063]&LFSRcolor2[667]&LFSRcolor2[755]);
    BiasedRNG[836] = (LFSRcolor2[971]&LFSRcolor2[481]&LFSRcolor2[19]&LFSRcolor2[60]);
    BiasedRNG[837] = (LFSRcolor2[90]&LFSRcolor2[701]&LFSRcolor2[1215]&LFSRcolor2[0]);
    BiasedRNG[838] = (LFSRcolor2[886]&LFSRcolor2[1281]&LFSRcolor2[348]&LFSRcolor2[1081]);
    BiasedRNG[839] = (LFSRcolor2[61]&LFSRcolor2[357]&LFSRcolor2[816]&LFSRcolor2[544]);
    BiasedRNG[840] = (LFSRcolor2[832]&LFSRcolor2[537]&LFSRcolor2[987]&LFSRcolor2[984]);
    BiasedRNG[841] = (LFSRcolor2[73]&LFSRcolor2[1041]&LFSRcolor2[1211]&LFSRcolor2[1105]);
    BiasedRNG[842] = (LFSRcolor2[1176]&LFSRcolor2[148]&LFSRcolor2[1044]&LFSRcolor2[871]);
    BiasedRNG[843] = (LFSRcolor2[1154]&LFSRcolor2[882]&LFSRcolor2[282]&LFSRcolor2[299]);
    BiasedRNG[844] = (LFSRcolor2[420]&LFSRcolor2[53]&LFSRcolor2[1047]&LFSRcolor2[751]);
    BiasedRNG[845] = (LFSRcolor2[952]&LFSRcolor2[853]&LFSRcolor2[492]&LFSRcolor2[584]);
    BiasedRNG[846] = (LFSRcolor2[593]&LFSRcolor2[1252]&LFSRcolor2[221]&LFSRcolor2[178]);
    BiasedRNG[847] = (LFSRcolor2[380]&LFSRcolor2[450]&LFSRcolor2[1115]&LFSRcolor2[996]);
    BiasedRNG[848] = (LFSRcolor2[951]&LFSRcolor2[841]&LFSRcolor2[1256]&LFSRcolor2[792]);
    BiasedRNG[849] = (LFSRcolor2[495]&LFSRcolor2[530]&LFSRcolor2[501]&LFSRcolor2[824]);
    BiasedRNG[850] = (LFSRcolor2[1106]&LFSRcolor2[852]&LFSRcolor2[866]&LFSRcolor2[16]);
    BiasedRNG[851] = (LFSRcolor2[1210]&LFSRcolor2[497]&LFSRcolor2[686]&LFSRcolor2[464]);
    BiasedRNG[852] = (LFSRcolor2[1163]&LFSRcolor2[854]&LFSRcolor2[194]&LFSRcolor2[1164]);
    BiasedRNG[853] = (LFSRcolor2[1236]&LFSRcolor2[127]&LFSRcolor2[476]&LFSRcolor2[370]);
    BiasedRNG[854] = (LFSRcolor2[939]&LFSRcolor2[112]&LFSRcolor2[321]&LFSRcolor2[641]);
    BiasedRNG[855] = (LFSRcolor2[831]&LFSRcolor2[153]&LFSRcolor2[155]&LFSRcolor2[1285]);
    BiasedRNG[856] = (LFSRcolor2[1039]&LFSRcolor2[177]&LFSRcolor2[778]&LFSRcolor2[764]);
    BiasedRNG[857] = (LFSRcolor2[931]&LFSRcolor2[227]&LFSRcolor2[673]&LFSRcolor2[1145]);
    BiasedRNG[858] = (LFSRcolor2[699]&LFSRcolor2[272]&LFSRcolor2[96]&LFSRcolor2[499]);
    BiasedRNG[859] = (LFSRcolor2[665]&LFSRcolor2[863]&LFSRcolor2[200]&LFSRcolor2[1069]);
    BiasedRNG[860] = (LFSRcolor2[278]&LFSRcolor2[423]&LFSRcolor2[154]&LFSRcolor2[329]);
    BiasedRNG[861] = (LFSRcolor2[596]&LFSRcolor2[338]&LFSRcolor2[190]&LFSRcolor2[396]);
    BiasedRNG[862] = (LFSRcolor2[47]&LFSRcolor2[1061]&LFSRcolor2[1168]&LFSRcolor2[551]);
    BiasedRNG[863] = (LFSRcolor2[124]&LFSRcolor2[1064]&LFSRcolor2[997]&LFSRcolor2[144]);
    BiasedRNG[864] = (LFSRcolor2[291]&LFSRcolor2[246]&LFSRcolor2[125]&LFSRcolor2[350]);
    BiasedRNG[865] = (LFSRcolor2[697]&LFSRcolor2[730]&LFSRcolor2[550]&LFSRcolor2[669]);
    BiasedRNG[866] = (LFSRcolor2[733]&LFSRcolor2[1172]&LFSRcolor2[795]&LFSRcolor2[540]);
    BiasedRNG[867] = (LFSRcolor2[288]&LFSRcolor2[130]&LFSRcolor2[484]&LFSRcolor2[224]);
    BiasedRNG[868] = (LFSRcolor2[1008]&LFSRcolor2[827]&LFSRcolor2[915]&LFSRcolor2[525]);
    BiasedRNG[869] = (LFSRcolor2[635]&LFSRcolor2[488]&LFSRcolor2[849]&LFSRcolor2[1117]);
    BiasedRNG[870] = (LFSRcolor2[558]&LFSRcolor2[895]&LFSRcolor2[249]&LFSRcolor2[244]);
    BiasedRNG[871] = (LFSRcolor2[335]&LFSRcolor2[345]&LFSRcolor2[622]&LFSRcolor2[546]);
    BiasedRNG[872] = (LFSRcolor2[648]&LFSRcolor2[1148]&LFSRcolor2[1161]&LFSRcolor2[869]);
    BiasedRNG[873] = (LFSRcolor2[268]&LFSRcolor2[1279]&LFSRcolor2[514]&LFSRcolor2[979]);
    BiasedRNG[874] = (LFSRcolor2[914]&LFSRcolor2[283]&LFSRcolor2[5]&LFSRcolor2[1202]);
    BiasedRNG[875] = (LFSRcolor2[738]&LFSRcolor2[573]&LFSRcolor2[808]&LFSRcolor2[129]);
    BiasedRNG[876] = (LFSRcolor2[1283]&LFSRcolor2[572]&LFSRcolor2[651]&LFSRcolor2[448]);
    BiasedRNG[877] = (LFSRcolor2[23]&LFSRcolor2[582]&LFSRcolor2[880]&LFSRcolor2[640]);
    BiasedRNG[878] = (LFSRcolor2[229]&LFSRcolor2[389]&LFSRcolor2[861]&LFSRcolor2[1011]);
    BiasedRNG[879] = (LFSRcolor2[9]&LFSRcolor2[623]&LFSRcolor2[102]&LFSRcolor2[1162]);
    BiasedRNG[880] = (LFSRcolor2[534]&LFSRcolor2[279]&LFSRcolor2[77]&LFSRcolor2[1135]);
    BiasedRNG[881] = (LFSRcolor2[1183]&LFSRcolor2[99]&LFSRcolor2[1103]&LFSRcolor2[900]);
    BiasedRNG[882] = (LFSRcolor2[739]&LFSRcolor2[184]&LFSRcolor2[599]&LFSRcolor2[936]);
    BiasedRNG[883] = (LFSRcolor2[403]&LFSRcolor2[563]&LFSRcolor2[400]&LFSRcolor2[138]);
    BiasedRNG[884] = (LFSRcolor2[122]&LFSRcolor2[1171]&LFSRcolor2[521]&LFSRcolor2[140]);
    BiasedRNG[885] = (LFSRcolor2[1228]&LFSRcolor2[1152]&LFSRcolor2[410]&LFSRcolor2[585]);
    BiasedRNG[886] = (LFSRcolor2[118]&LFSRcolor2[642]&LFSRcolor2[41]&LFSRcolor2[365]);
    BiasedRNG[887] = (LFSRcolor2[1181]&LFSRcolor2[480]&LFSRcolor2[310]&LFSRcolor2[858]);
    BiasedRNG[888] = (LFSRcolor2[713]&LFSRcolor2[119]&LFSRcolor2[891]&LFSRcolor2[101]);
    BiasedRNG[889] = (LFSRcolor2[52]&LFSRcolor2[255]&LFSRcolor2[757]&LFSRcolor2[535]);
    BiasedRNG[890] = (LFSRcolor2[1128]&LFSRcolor2[1137]&LFSRcolor2[498]&LFSRcolor2[451]);
    BiasedRNG[891] = (LFSRcolor2[637]&LFSRcolor2[88]&LFSRcolor2[1089]&LFSRcolor2[994]);
    BiasedRNG[892] = (LFSRcolor2[146]&LFSRcolor2[443]&LFSRcolor2[598]&LFSRcolor2[1259]);
    BiasedRNG[893] = (LFSRcolor2[840]&LFSRcolor2[769]&LFSRcolor2[857]&LFSRcolor2[187]);
    BiasedRNG[894] = (LFSRcolor2[284]&LFSRcolor2[49]&LFSRcolor2[1209]&LFSRcolor2[214]);
    UnbiasedRNG[496] = LFSRcolor2[796];
    UnbiasedRNG[497] = LFSRcolor2[105];
    UnbiasedRNG[498] = LFSRcolor2[402];
    UnbiasedRNG[499] = LFSRcolor2[815];
    UnbiasedRNG[500] = LFSRcolor2[986];
    UnbiasedRNG[501] = LFSRcolor2[1264];
    UnbiasedRNG[502] = LFSRcolor2[702];
    UnbiasedRNG[503] = LFSRcolor2[1265];
    UnbiasedRNG[504] = LFSRcolor2[274];
    UnbiasedRNG[505] = LFSRcolor2[1088];
    UnbiasedRNG[506] = LFSRcolor2[980];
    UnbiasedRNG[507] = LFSRcolor2[862];
    UnbiasedRNG[508] = LFSRcolor2[169];
    UnbiasedRNG[509] = LFSRcolor2[1258];
    UnbiasedRNG[510] = LFSRcolor2[500];
    UnbiasedRNG[511] = LFSRcolor2[71];
    UnbiasedRNG[512] = LFSRcolor2[142];
    UnbiasedRNG[513] = LFSRcolor2[250];
    UnbiasedRNG[514] = LFSRcolor2[27];
    UnbiasedRNG[515] = LFSRcolor2[135];
    UnbiasedRNG[516] = LFSRcolor2[837];
    UnbiasedRNG[517] = LFSRcolor2[760];
    UnbiasedRNG[518] = LFSRcolor2[173];
    UnbiasedRNG[519] = LFSRcolor2[387];
    UnbiasedRNG[520] = LFSRcolor2[884];
    UnbiasedRNG[521] = LFSRcolor2[617];
    UnbiasedRNG[522] = LFSRcolor2[37];
    UnbiasedRNG[523] = LFSRcolor2[42];
    UnbiasedRNG[524] = LFSRcolor2[292];
    UnbiasedRNG[525] = LFSRcolor2[29];
    UnbiasedRNG[526] = LFSRcolor2[117];
    UnbiasedRNG[527] = LFSRcolor2[564];
    UnbiasedRNG[528] = LFSRcolor2[1079];
    UnbiasedRNG[529] = LFSRcolor2[143];
    UnbiasedRNG[530] = LFSRcolor2[397];
    UnbiasedRNG[531] = LFSRcolor2[267];
    UnbiasedRNG[532] = LFSRcolor2[1078];
    UnbiasedRNG[533] = LFSRcolor2[804];
    UnbiasedRNG[534] = LFSRcolor2[1266];
    UnbiasedRNG[535] = LFSRcolor2[176];
    UnbiasedRNG[536] = LFSRcolor2[92];
    UnbiasedRNG[537] = LFSRcolor2[225];
    UnbiasedRNG[538] = LFSRcolor2[406];
    UnbiasedRNG[539] = LFSRcolor2[549];
    UnbiasedRNG[540] = LFSRcolor2[59];
    UnbiasedRNG[541] = LFSRcolor2[182];
    UnbiasedRNG[542] = LFSRcolor2[111];
    UnbiasedRNG[543] = LFSRcolor2[592];
    UnbiasedRNG[544] = LFSRcolor2[1108];
    UnbiasedRNG[545] = LFSRcolor2[519];
    UnbiasedRNG[546] = LFSRcolor2[1119];
    UnbiasedRNG[547] = LFSRcolor2[527];
    UnbiasedRNG[548] = LFSRcolor2[1046];
    UnbiasedRNG[549] = LFSRcolor2[569];
    UnbiasedRNG[550] = LFSRcolor2[1112];
    UnbiasedRNG[551] = LFSRcolor2[48];
    UnbiasedRNG[552] = LFSRcolor2[794];
    UnbiasedRNG[553] = LFSRcolor2[790];
    UnbiasedRNG[554] = LFSRcolor2[856];
    UnbiasedRNG[555] = LFSRcolor2[711];
    UnbiasedRNG[556] = LFSRcolor2[228];
    UnbiasedRNG[557] = LFSRcolor2[219];
    UnbiasedRNG[558] = LFSRcolor2[1192];
    UnbiasedRNG[559] = LFSRcolor2[1096];
    UnbiasedRNG[560] = LFSRcolor2[724];
    UnbiasedRNG[561] = LFSRcolor2[1015];
    UnbiasedRNG[562] = LFSRcolor2[607];
    UnbiasedRNG[563] = LFSRcolor2[294];
    UnbiasedRNG[564] = LFSRcolor2[22];
    UnbiasedRNG[565] = LFSRcolor2[818];
    UnbiasedRNG[566] = LFSRcolor2[677];
    UnbiasedRNG[567] = LFSRcolor2[217];
    UnbiasedRNG[568] = LFSRcolor2[801];
    UnbiasedRNG[569] = LFSRcolor2[938];
    UnbiasedRNG[570] = LFSRcolor2[13];
    UnbiasedRNG[571] = LFSRcolor2[1219];
    UnbiasedRNG[572] = LFSRcolor2[339];
    UnbiasedRNG[573] = LFSRcolor2[913];
    UnbiasedRNG[574] = LFSRcolor2[634];
    UnbiasedRNG[575] = LFSRcolor2[265];
    UnbiasedRNG[576] = LFSRcolor2[606];
    UnbiasedRNG[577] = LFSRcolor2[973];
    UnbiasedRNG[578] = LFSRcolor2[87];
    UnbiasedRNG[579] = LFSRcolor2[967];
    UnbiasedRNG[580] = LFSRcolor2[93];
    UnbiasedRNG[581] = LFSRcolor2[337];
    UnbiasedRNG[582] = LFSRcolor2[744];
    UnbiasedRNG[583] = LFSRcolor2[296];
    UnbiasedRNG[584] = LFSRcolor2[391];
    UnbiasedRNG[585] = LFSRcolor2[1195];
    UnbiasedRNG[586] = LFSRcolor2[1197];
    UnbiasedRNG[587] = LFSRcolor2[286];
    UnbiasedRNG[588] = LFSRcolor2[237];
    UnbiasedRNG[589] = LFSRcolor2[1240];
    UnbiasedRNG[590] = LFSRcolor2[25];
    UnbiasedRNG[591] = LFSRcolor2[230];
    UnbiasedRNG[592] = LFSRcolor2[1051];
    UnbiasedRNG[593] = LFSRcolor2[341];
    UnbiasedRNG[594] = LFSRcolor2[437];
    UnbiasedRNG[595] = LFSRcolor2[1284];
    UnbiasedRNG[596] = LFSRcolor2[740];
    UnbiasedRNG[597] = LFSRcolor2[1134];
    UnbiasedRNG[598] = LFSRcolor2[1263];
    UnbiasedRNG[599] = LFSRcolor2[717];
    UnbiasedRNG[600] = LFSRcolor2[706];
    UnbiasedRNG[601] = LFSRcolor2[1184];
    UnbiasedRNG[602] = LFSRcolor2[1286];
    UnbiasedRNG[603] = LFSRcolor2[589];
    UnbiasedRNG[604] = LFSRcolor2[1065];
    UnbiasedRNG[605] = LFSRcolor2[405];
    UnbiasedRNG[606] = LFSRcolor2[86];
    UnbiasedRNG[607] = LFSRcolor2[1277];
    UnbiasedRNG[608] = LFSRcolor2[929];
    UnbiasedRNG[609] = LFSRcolor2[890];
    UnbiasedRNG[610] = LFSRcolor2[1124];
    UnbiasedRNG[611] = LFSRcolor2[932];
    UnbiasedRNG[612] = LFSRcolor2[646];
    UnbiasedRNG[613] = LFSRcolor2[252];
    UnbiasedRNG[614] = LFSRcolor2[652];
    UnbiasedRNG[615] = LFSRcolor2[305];
    UnbiasedRNG[616] = LFSRcolor2[180];
    UnbiasedRNG[617] = LFSRcolor2[12];
    UnbiasedRNG[618] = LFSRcolor2[925];
    UnbiasedRNG[619] = LFSRcolor2[62];
    UnbiasedRNG[620] = LFSRcolor2[179];
    UnbiasedRNG[621] = LFSRcolor2[844];
    UnbiasedRNG[622] = LFSRcolor2[691];
    UnbiasedRNG[623] = LFSRcolor2[1007];
    UnbiasedRNG[624] = LFSRcolor2[835];
    UnbiasedRNG[625] = LFSRcolor2[943];
    UnbiasedRNG[626] = LFSRcolor2[82];
    UnbiasedRNG[627] = LFSRcolor2[698];
    UnbiasedRNG[628] = LFSRcolor2[470];
    UnbiasedRNG[629] = LFSRcolor2[799];
    UnbiasedRNG[630] = LFSRcolor2[621];
    UnbiasedRNG[631] = LFSRcolor2[275];
    UnbiasedRNG[632] = LFSRcolor2[1273];
    UnbiasedRNG[633] = LFSRcolor2[1040];
    UnbiasedRNG[634] = LFSRcolor2[926];
    UnbiasedRNG[635] = LFSRcolor2[998];
    UnbiasedRNG[636] = LFSRcolor2[150];
    UnbiasedRNG[637] = LFSRcolor2[695];
    UnbiasedRNG[638] = LFSRcolor2[364];
    UnbiasedRNG[639] = LFSRcolor2[233];
    UnbiasedRNG[640] = LFSRcolor2[208];
    UnbiasedRNG[641] = LFSRcolor2[752];
    UnbiasedRNG[642] = LFSRcolor2[1083];
    UnbiasedRNG[643] = LFSRcolor2[342];
    UnbiasedRNG[644] = LFSRcolor2[1019];
    UnbiasedRNG[645] = LFSRcolor2[720];
    UnbiasedRNG[646] = LFSRcolor2[215];
    UnbiasedRNG[647] = LFSRcolor2[548];
    UnbiasedRNG[648] = LFSRcolor2[532];
    UnbiasedRNG[649] = LFSRcolor2[901];
    UnbiasedRNG[650] = LFSRcolor2[38];
    UnbiasedRNG[651] = LFSRcolor2[632];
    UnbiasedRNG[652] = LFSRcolor2[761];
    UnbiasedRNG[653] = LFSRcolor2[308];
    UnbiasedRNG[654] = LFSRcolor2[903];
    UnbiasedRNG[655] = LFSRcolor2[116];
    UnbiasedRNG[656] = LFSRcolor2[567];
    UnbiasedRNG[657] = LFSRcolor2[523];
    UnbiasedRNG[658] = LFSRcolor2[797];
    UnbiasedRNG[659] = LFSRcolor2[280];
    UnbiasedRNG[660] = LFSRcolor2[1190];
    UnbiasedRNG[661] = LFSRcolor2[298];
    UnbiasedRNG[662] = LFSRcolor2[1002];
    UnbiasedRNG[663] = LFSRcolor2[1012];
    UnbiasedRNG[664] = LFSRcolor2[78];
    UnbiasedRNG[665] = LFSRcolor2[753];
    UnbiasedRNG[666] = LFSRcolor2[704];
    UnbiasedRNG[667] = LFSRcolor2[872];
    UnbiasedRNG[668] = LFSRcolor2[885];
    UnbiasedRNG[669] = LFSRcolor2[552];
    UnbiasedRNG[670] = LFSRcolor2[1147];
    UnbiasedRNG[671] = LFSRcolor2[98];
    UnbiasedRNG[672] = LFSRcolor2[1158];
    UnbiasedRNG[673] = LFSRcolor2[108];
    UnbiasedRNG[674] = LFSRcolor2[649];
    UnbiasedRNG[675] = LFSRcolor2[1227];
    UnbiasedRNG[676] = LFSRcolor2[1276];
    UnbiasedRNG[677] = LFSRcolor2[113];
    UnbiasedRNG[678] = LFSRcolor2[260];
    UnbiasedRNG[679] = LFSRcolor2[508];
    UnbiasedRNG[680] = LFSRcolor2[360];
    UnbiasedRNG[681] = LFSRcolor2[91];
    UnbiasedRNG[682] = LFSRcolor2[1238];
    UnbiasedRNG[683] = LFSRcolor2[517];
    UnbiasedRNG[684] = LFSRcolor2[1232];
    UnbiasedRNG[685] = LFSRcolor2[271];
    UnbiasedRNG[686] = LFSRcolor2[982];
    UnbiasedRNG[687] = LFSRcolor2[168];
    UnbiasedRNG[688] = LFSRcolor2[571];
    UnbiasedRNG[689] = LFSRcolor2[705];
    UnbiasedRNG[690] = LFSRcolor2[491];
    UnbiasedRNG[691] = LFSRcolor2[193];
    UnbiasedRNG[692] = LFSRcolor2[787];
    UnbiasedRNG[693] = LFSRcolor2[1150];
    UnbiasedRNG[694] = LFSRcolor2[45];
    UnbiasedRNG[695] = LFSRcolor2[377];
    UnbiasedRNG[696] = LFSRcolor2[921];
    UnbiasedRNG[697] = LFSRcolor2[454];
    UnbiasedRNG[698] = LFSRcolor2[328];
    UnbiasedRNG[699] = LFSRcolor2[121];
    UnbiasedRNG[700] = LFSRcolor2[817];
    UnbiasedRNG[701] = LFSRcolor2[1205];
    UnbiasedRNG[702] = LFSRcolor2[1151];
    UnbiasedRNG[703] = LFSRcolor2[843];
    UnbiasedRNG[704] = LFSRcolor2[1055];
    UnbiasedRNG[705] = LFSRcolor2[258];
    UnbiasedRNG[706] = LFSRcolor2[543];
    UnbiasedRNG[707] = LFSRcolor2[846];
    UnbiasedRNG[708] = LFSRcolor2[894];
    UnbiasedRNG[709] = LFSRcolor2[709];
    UnbiasedRNG[710] = LFSRcolor2[165];
    UnbiasedRNG[711] = LFSRcolor2[383];
    UnbiasedRNG[712] = LFSRcolor2[528];
    UnbiasedRNG[713] = LFSRcolor2[223];
    UnbiasedRNG[714] = LFSRcolor2[80];
    UnbiasedRNG[715] = LFSRcolor2[202];
    UnbiasedRNG[716] = LFSRcolor2[661];
    UnbiasedRNG[717] = LFSRcolor2[688];
    UnbiasedRNG[718] = LFSRcolor2[754];
    UnbiasedRNG[719] = LFSRcolor2[531];
    UnbiasedRNG[720] = LFSRcolor2[3];
    UnbiasedRNG[721] = LFSRcolor2[76];
    UnbiasedRNG[722] = LFSRcolor2[433];
    UnbiasedRNG[723] = LFSRcolor2[1221];
    UnbiasedRNG[724] = LFSRcolor2[198];
    UnbiasedRNG[725] = LFSRcolor2[145];
    UnbiasedRNG[726] = LFSRcolor2[1136];
    UnbiasedRNG[727] = LFSRcolor2[881];
    UnbiasedRNG[728] = LFSRcolor2[123];
    UnbiasedRNG[729] = LFSRcolor2[51];
    UnbiasedRNG[730] = LFSRcolor2[953];
    UnbiasedRNG[731] = LFSRcolor2[1126];
    UnbiasedRNG[732] = LFSRcolor2[259];
    UnbiasedRNG[733] = LFSRcolor2[712];
    UnbiasedRNG[734] = LFSRcolor2[806];
    UnbiasedRNG[735] = LFSRcolor2[466];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[736] = LFSRcolor3[46];
    UnbiasedRNG[737] = LFSRcolor3[195];
    UnbiasedRNG[738] = LFSRcolor3[86];
    UnbiasedRNG[739] = LFSRcolor3[24];
    UnbiasedRNG[740] = LFSRcolor3[19];
    UnbiasedRNG[741] = LFSRcolor3[5];
    UnbiasedRNG[742] = LFSRcolor3[39];
    UnbiasedRNG[743] = LFSRcolor3[107];
    UnbiasedRNG[744] = LFSRcolor3[104];
    UnbiasedRNG[745] = LFSRcolor3[84];
    UnbiasedRNG[746] = LFSRcolor3[186];
    UnbiasedRNG[747] = LFSRcolor3[70];
    UnbiasedRNG[748] = LFSRcolor3[220];
    UnbiasedRNG[749] = LFSRcolor3[37];
    UnbiasedRNG[750] = LFSRcolor3[58];
    UnbiasedRNG[751] = LFSRcolor3[26];
    UnbiasedRNG[752] = LFSRcolor3[181];
    UnbiasedRNG[753] = LFSRcolor3[217];
    UnbiasedRNG[754] = LFSRcolor3[187];
    UnbiasedRNG[755] = LFSRcolor3[203];
    UnbiasedRNG[756] = LFSRcolor3[214];
    UnbiasedRNG[757] = LFSRcolor3[216];
    UnbiasedRNG[758] = LFSRcolor3[172];
    UnbiasedRNG[759] = LFSRcolor3[158];
    UnbiasedRNG[760] = LFSRcolor3[171];
    UnbiasedRNG[761] = LFSRcolor3[1];
    UnbiasedRNG[762] = LFSRcolor3[153];
    UnbiasedRNG[763] = LFSRcolor3[89];
    UnbiasedRNG[764] = LFSRcolor3[174];
    UnbiasedRNG[765] = LFSRcolor3[112];
    UnbiasedRNG[766] = LFSRcolor3[2];
    UnbiasedRNG[767] = LFSRcolor3[177];
    UnbiasedRNG[768] = LFSRcolor3[140];
    UnbiasedRNG[769] = LFSRcolor3[152];
    UnbiasedRNG[770] = LFSRcolor3[10];
    UnbiasedRNG[771] = LFSRcolor3[98];
    UnbiasedRNG[772] = LFSRcolor3[115];
    UnbiasedRNG[773] = LFSRcolor3[80];
    UnbiasedRNG[774] = LFSRcolor3[78];
    UnbiasedRNG[775] = LFSRcolor3[179];
    UnbiasedRNG[776] = LFSRcolor3[71];
    UnbiasedRNG[777] = LFSRcolor3[51];
    UnbiasedRNG[778] = LFSRcolor3[62];
    UnbiasedRNG[779] = LFSRcolor3[116];
    UnbiasedRNG[780] = LFSRcolor3[8];
    UnbiasedRNG[781] = LFSRcolor3[36];
    UnbiasedRNG[782] = LFSRcolor3[28];
    UnbiasedRNG[783] = LFSRcolor3[184];
    UnbiasedRNG[784] = LFSRcolor3[47];
    UnbiasedRNG[785] = LFSRcolor3[126];
    UnbiasedRNG[786] = LFSRcolor3[161];
    UnbiasedRNG[787] = LFSRcolor3[27];
    UnbiasedRNG[788] = LFSRcolor3[200];
    UnbiasedRNG[789] = LFSRcolor3[97];
    UnbiasedRNG[790] = LFSRcolor3[149];
    UnbiasedRNG[791] = LFSRcolor3[48];
    UnbiasedRNG[792] = LFSRcolor3[207];
    UnbiasedRNG[793] = LFSRcolor3[148];
    UnbiasedRNG[794] = LFSRcolor3[64];
    UnbiasedRNG[795] = LFSRcolor3[227];
    UnbiasedRNG[796] = LFSRcolor3[137];
    UnbiasedRNG[797] = LFSRcolor3[210];
    UnbiasedRNG[798] = LFSRcolor3[23];
    UnbiasedRNG[799] = LFSRcolor3[75];
    UnbiasedRNG[800] = LFSRcolor3[4];
    UnbiasedRNG[801] = LFSRcolor3[132];
    UnbiasedRNG[802] = LFSRcolor3[156];
    UnbiasedRNG[803] = LFSRcolor3[69];
    UnbiasedRNG[804] = LFSRcolor3[73];
    UnbiasedRNG[805] = LFSRcolor3[81];
    UnbiasedRNG[806] = LFSRcolor3[52];
    UnbiasedRNG[807] = LFSRcolor3[213];
    UnbiasedRNG[808] = LFSRcolor3[111];
    UnbiasedRNG[809] = LFSRcolor3[99];
    UnbiasedRNG[810] = LFSRcolor3[65];
    UnbiasedRNG[811] = LFSRcolor3[165];
    UnbiasedRNG[812] = LFSRcolor3[68];
    UnbiasedRNG[813] = LFSRcolor3[20];
    UnbiasedRNG[814] = LFSRcolor3[185];
    UnbiasedRNG[815] = LFSRcolor3[163];
    UnbiasedRNG[816] = LFSRcolor3[110];
    UnbiasedRNG[817] = LFSRcolor3[169];
    UnbiasedRNG[818] = LFSRcolor3[125];
    UnbiasedRNG[819] = LFSRcolor3[94];
    UnbiasedRNG[820] = LFSRcolor3[168];
    UnbiasedRNG[821] = LFSRcolor3[67];
    UnbiasedRNG[822] = LFSRcolor3[175];
    UnbiasedRNG[823] = LFSRcolor3[82];
    UnbiasedRNG[824] = LFSRcolor3[121];
    UnbiasedRNG[825] = LFSRcolor3[204];
    UnbiasedRNG[826] = LFSRcolor3[190];
    UnbiasedRNG[827] = LFSRcolor3[120];
    UnbiasedRNG[828] = LFSRcolor3[167];
    UnbiasedRNG[829] = LFSRcolor3[42];
    UnbiasedRNG[830] = LFSRcolor3[154];
    UnbiasedRNG[831] = LFSRcolor3[95];
    UnbiasedRNG[832] = LFSRcolor3[142];
    UnbiasedRNG[833] = LFSRcolor3[219];
    UnbiasedRNG[834] = LFSRcolor3[201];
    UnbiasedRNG[835] = LFSRcolor3[32];
    UnbiasedRNG[836] = LFSRcolor3[87];
    UnbiasedRNG[837] = LFSRcolor3[21];
    UnbiasedRNG[838] = LFSRcolor3[41];
    UnbiasedRNG[839] = LFSRcolor3[193];
    UnbiasedRNG[840] = LFSRcolor3[109];
    UnbiasedRNG[841] = LFSRcolor3[133];
    UnbiasedRNG[842] = LFSRcolor3[85];
    UnbiasedRNG[843] = LFSRcolor3[22];
    UnbiasedRNG[844] = LFSRcolor3[128];
    UnbiasedRNG[845] = LFSRcolor3[117];
    UnbiasedRNG[846] = LFSRcolor3[212];
    UnbiasedRNG[847] = LFSRcolor3[194];
    UnbiasedRNG[848] = LFSRcolor3[206];
    UnbiasedRNG[849] = LFSRcolor3[40];
    UnbiasedRNG[850] = LFSRcolor3[29];
    UnbiasedRNG[851] = LFSRcolor3[218];
    UnbiasedRNG[852] = LFSRcolor3[76];
    UnbiasedRNG[853] = LFSRcolor3[77];
    UnbiasedRNG[854] = LFSRcolor3[45];
    UnbiasedRNG[855] = LFSRcolor3[54];
    UnbiasedRNG[856] = LFSRcolor3[50];
    UnbiasedRNG[857] = LFSRcolor3[113];
    UnbiasedRNG[858] = LFSRcolor3[30];
    UnbiasedRNG[859] = LFSRcolor3[160];
    UnbiasedRNG[860] = LFSRcolor3[182];
    UnbiasedRNG[861] = LFSRcolor3[103];
    UnbiasedRNG[862] = LFSRcolor3[145];
    UnbiasedRNG[863] = LFSRcolor3[224];
    UnbiasedRNG[864] = LFSRcolor3[12];
    UnbiasedRNG[865] = LFSRcolor3[53];
    UnbiasedRNG[866] = LFSRcolor3[198];
    UnbiasedRNG[867] = LFSRcolor3[100];
    UnbiasedRNG[868] = LFSRcolor3[176];
    UnbiasedRNG[869] = LFSRcolor3[101];
    UnbiasedRNG[870] = LFSRcolor3[93];
    UnbiasedRNG[871] = LFSRcolor3[211];
    UnbiasedRNG[872] = LFSRcolor3[199];
    UnbiasedRNG[873] = LFSRcolor3[197];
    UnbiasedRNG[874] = LFSRcolor3[61];
    UnbiasedRNG[875] = LFSRcolor3[222];
    UnbiasedRNG[876] = LFSRcolor3[88];
    UnbiasedRNG[877] = LFSRcolor3[134];
    UnbiasedRNG[878] = LFSRcolor3[178];
    UnbiasedRNG[879] = LFSRcolor3[25];
    UnbiasedRNG[880] = LFSRcolor3[13];
    UnbiasedRNG[881] = LFSRcolor3[221];
    UnbiasedRNG[882] = LFSRcolor3[74];
    UnbiasedRNG[883] = LFSRcolor3[146];
    UnbiasedRNG[884] = LFSRcolor3[18];
    UnbiasedRNG[885] = LFSRcolor3[202];
    UnbiasedRNG[886] = LFSRcolor3[124];
    UnbiasedRNG[887] = LFSRcolor3[43];
    UnbiasedRNG[888] = LFSRcolor3[229];
    UnbiasedRNG[889] = LFSRcolor3[90];
    UnbiasedRNG[890] = LFSRcolor3[139];
    UnbiasedRNG[891] = LFSRcolor3[226];
    UnbiasedRNG[892] = LFSRcolor3[180];
    UnbiasedRNG[893] = LFSRcolor3[144];
    UnbiasedRNG[894] = LFSRcolor3[114];
    UnbiasedRNG[895] = LFSRcolor3[59];
    UnbiasedRNG[896] = LFSRcolor3[155];
    UnbiasedRNG[897] = LFSRcolor3[72];
    UnbiasedRNG[898] = LFSRcolor3[17];
    UnbiasedRNG[899] = LFSRcolor3[16];
    UnbiasedRNG[900] = LFSRcolor3[122];
    UnbiasedRNG[901] = LFSRcolor3[79];
    UnbiasedRNG[902] = LFSRcolor3[130];
    UnbiasedRNG[903] = LFSRcolor3[129];
    UnbiasedRNG[904] = LFSRcolor3[189];
    UnbiasedRNG[905] = LFSRcolor3[205];
    UnbiasedRNG[906] = LFSRcolor3[188];
    UnbiasedRNG[907] = LFSRcolor3[66];
    UnbiasedRNG[908] = LFSRcolor3[208];
    UnbiasedRNG[909] = LFSRcolor3[143];
    UnbiasedRNG[910] = LFSRcolor3[166];
    UnbiasedRNG[911] = LFSRcolor3[192];
    UnbiasedRNG[912] = LFSRcolor3[63];
    UnbiasedRNG[913] = LFSRcolor3[157];
    UnbiasedRNG[914] = LFSRcolor3[151];
    UnbiasedRNG[915] = LFSRcolor3[56];
    UnbiasedRNG[916] = LFSRcolor3[196];
    UnbiasedRNG[917] = LFSRcolor3[14];
    UnbiasedRNG[918] = LFSRcolor3[173];
    UnbiasedRNG[919] = LFSRcolor3[147];
    UnbiasedRNG[920] = LFSRcolor3[209];
    UnbiasedRNG[921] = LFSRcolor3[33];
    UnbiasedRNG[922] = LFSRcolor3[7];
    UnbiasedRNG[923] = LFSRcolor3[60];
    UnbiasedRNG[924] = LFSRcolor3[123];
    UnbiasedRNG[925] = LFSRcolor3[31];
    UnbiasedRNG[926] = LFSRcolor3[9];
    UnbiasedRNG[927] = LFSRcolor3[150];
    UnbiasedRNG[928] = LFSRcolor3[106];
    UnbiasedRNG[929] = LFSRcolor3[0];
    UnbiasedRNG[930] = LFSRcolor3[11];
    UnbiasedRNG[931] = LFSRcolor3[102];
    UnbiasedRNG[932] = LFSRcolor3[228];
    UnbiasedRNG[933] = LFSRcolor3[223];
    UnbiasedRNG[934] = LFSRcolor3[138];
    UnbiasedRNG[935] = LFSRcolor3[92];
    UnbiasedRNG[936] = LFSRcolor3[108];
    UnbiasedRNG[937] = LFSRcolor3[135];
    UnbiasedRNG[938] = LFSRcolor3[118];
    UnbiasedRNG[939] = LFSRcolor3[91];
    UnbiasedRNG[940] = LFSRcolor3[83];
    UnbiasedRNG[941] = LFSRcolor3[15];
    UnbiasedRNG[942] = LFSRcolor3[127];
    UnbiasedRNG[943] = LFSRcolor3[183];
    UnbiasedRNG[944] = LFSRcolor3[55];
    UnbiasedRNG[945] = LFSRcolor3[57];
end

always @(posedge color3_clk) begin
    BiasedRNG[895] = (LFSRcolor4[777]&LFSRcolor4[891]&LFSRcolor4[151]&LFSRcolor4[863]);
    BiasedRNG[896] = (LFSRcolor4[451]&LFSRcolor4[763]&LFSRcolor4[622]&LFSRcolor4[686]);
    BiasedRNG[897] = (LFSRcolor4[39]&LFSRcolor4[66]&LFSRcolor4[603]&LFSRcolor4[546]);
    BiasedRNG[898] = (LFSRcolor4[859]&LFSRcolor4[676]&LFSRcolor4[926]&LFSRcolor4[215]);
    BiasedRNG[899] = (LFSRcolor4[209]&LFSRcolor4[761]&LFSRcolor4[821]&LFSRcolor4[797]);
    BiasedRNG[900] = (LFSRcolor4[724]&LFSRcolor4[35]&LFSRcolor4[135]&LFSRcolor4[943]);
    BiasedRNG[901] = (LFSRcolor4[652]&LFSRcolor4[198]&LFSRcolor4[455]&LFSRcolor4[359]);
    BiasedRNG[902] = (LFSRcolor4[261]&LFSRcolor4[816]&LFSRcolor4[239]&LFSRcolor4[281]);
    BiasedRNG[903] = (LFSRcolor4[568]&LFSRcolor4[313]&LFSRcolor4[872]&LFSRcolor4[138]);
    BiasedRNG[904] = (LFSRcolor4[785]&LFSRcolor4[256]&LFSRcolor4[612]&LFSRcolor4[526]);
    BiasedRNG[905] = (LFSRcolor4[255]&LFSRcolor4[807]&LFSRcolor4[611]&LFSRcolor4[132]);
    BiasedRNG[906] = (LFSRcolor4[440]&LFSRcolor4[49]&LFSRcolor4[391]&LFSRcolor4[702]);
    BiasedRNG[907] = (LFSRcolor4[713]&LFSRcolor4[541]&LFSRcolor4[375]&LFSRcolor4[202]);
    BiasedRNG[908] = (LFSRcolor4[108]&LFSRcolor4[574]&LFSRcolor4[457]&LFSRcolor4[908]);
    BiasedRNG[909] = (LFSRcolor4[741]&LFSRcolor4[715]&LFSRcolor4[836]&LFSRcolor4[540]);
    BiasedRNG[910] = (LFSRcolor4[576]&LFSRcolor4[409]&LFSRcolor4[382]&LFSRcolor4[760]);
    BiasedRNG[911] = (LFSRcolor4[271]&LFSRcolor4[607]&LFSRcolor4[698]&LFSRcolor4[648]);
    BiasedRNG[912] = (LFSRcolor4[111]&LFSRcolor4[792]&LFSRcolor4[819]&LFSRcolor4[822]);
    BiasedRNG[913] = (LFSRcolor4[303]&LFSRcolor4[827]&LFSRcolor4[98]&LFSRcolor4[858]);
    BiasedRNG[914] = (LFSRcolor4[380]&LFSRcolor4[466]&LFSRcolor4[245]&LFSRcolor4[894]);
    BiasedRNG[915] = (LFSRcolor4[877]&LFSRcolor4[678]&LFSRcolor4[22]&LFSRcolor4[498]);
    BiasedRNG[916] = (LFSRcolor4[532]&LFSRcolor4[887]&LFSRcolor4[448]&LFSRcolor4[627]);
    BiasedRNG[917] = (LFSRcolor4[572]&LFSRcolor4[589]&LFSRcolor4[264]&LFSRcolor4[673]);
    BiasedRNG[918] = (LFSRcolor4[250]&LFSRcolor4[731]&LFSRcolor4[125]&LFSRcolor4[77]);
    BiasedRNG[919] = (LFSRcolor4[205]&LFSRcolor4[25]&LFSRcolor4[240]&LFSRcolor4[140]);
    BiasedRNG[920] = (LFSRcolor4[505]&LFSRcolor4[55]&LFSRcolor4[742]&LFSRcolor4[6]);
    BiasedRNG[921] = (LFSRcolor4[835]&LFSRcolor4[578]&LFSRcolor4[89]&LFSRcolor4[306]);
    BiasedRNG[922] = (LFSRcolor4[591]&LFSRcolor4[844]&LFSRcolor4[638]&LFSRcolor4[867]);
    BiasedRNG[923] = (LFSRcolor4[280]&LFSRcolor4[60]&LFSRcolor4[637]&LFSRcolor4[459]);
    BiasedRNG[924] = (LFSRcolor4[865]&LFSRcolor4[107]&LFSRcolor4[404]&LFSRcolor4[928]);
    BiasedRNG[925] = (LFSRcolor4[482]&LFSRcolor4[486]&LFSRcolor4[598]&LFSRcolor4[879]);
    BiasedRNG[926] = (LFSRcolor4[524]&LFSRcolor4[600]&LFSRcolor4[137]&LFSRcolor4[300]);
    BiasedRNG[927] = (LFSRcolor4[10]&LFSRcolor4[178]&LFSRcolor4[421]&LFSRcolor4[784]);
    BiasedRNG[928] = (LFSRcolor4[8]&LFSRcolor4[463]&LFSRcolor4[387]&LFSRcolor4[737]);
    BiasedRNG[929] = (LFSRcolor4[90]&LFSRcolor4[259]&LFSRcolor4[664]&LFSRcolor4[383]);
    BiasedRNG[930] = (LFSRcolor4[224]&LFSRcolor4[18]&LFSRcolor4[438]&LFSRcolor4[295]);
    BiasedRNG[931] = (LFSRcolor4[292]&LFSRcolor4[927]&LFSRcolor4[272]&LFSRcolor4[832]);
    BiasedRNG[932] = (LFSRcolor4[919]&LFSRcolor4[144]&LFSRcolor4[754]&LFSRcolor4[308]);
    BiasedRNG[933] = (LFSRcolor4[839]&LFSRcolor4[374]&LFSRcolor4[284]&LFSRcolor4[503]);
    BiasedRNG[934] = (LFSRcolor4[901]&LFSRcolor4[62]&LFSRcolor4[458]&LFSRcolor4[182]);
    BiasedRNG[935] = (LFSRcolor4[762]&LFSRcolor4[353]&LFSRcolor4[251]&LFSRcolor4[393]);
    BiasedRNG[936] = (LFSRcolor4[207]&LFSRcolor4[615]&LFSRcolor4[142]&LFSRcolor4[770]);
    BiasedRNG[937] = (LFSRcolor4[947]&LFSRcolor4[34]&LFSRcolor4[502]&LFSRcolor4[536]);
    BiasedRNG[938] = (LFSRcolor4[512]&LFSRcolor4[586]&LFSRcolor4[806]&LFSRcolor4[917]);
    BiasedRNG[939] = (LFSRcolor4[848]&LFSRcolor4[156]&LFSRcolor4[845]&LFSRcolor4[340]);
    BiasedRNG[940] = (LFSRcolor4[361]&LFSRcolor4[525]&LFSRcolor4[67]&LFSRcolor4[236]);
    BiasedRNG[941] = (LFSRcolor4[543]&LFSRcolor4[320]&LFSRcolor4[783]&LFSRcolor4[475]);
    BiasedRNG[942] = (LFSRcolor4[467]&LFSRcolor4[247]&LFSRcolor4[237]&LFSRcolor4[685]);
    BiasedRNG[943] = (LFSRcolor4[561]&LFSRcolor4[623]&LFSRcolor4[874]&LFSRcolor4[902]);
    BiasedRNG[944] = (LFSRcolor4[403]&LFSRcolor4[496]&LFSRcolor4[213]&LFSRcolor4[59]);
    BiasedRNG[945] = (LFSRcolor4[95]&LFSRcolor4[921]&LFSRcolor4[871]&LFSRcolor4[483]);
    BiasedRNG[946] = (LFSRcolor4[857]&LFSRcolor4[775]&LFSRcolor4[700]&LFSRcolor4[217]);
    BiasedRNG[947] = (LFSRcolor4[220]&LFSRcolor4[799]&LFSRcolor4[196]&LFSRcolor4[100]);
    BiasedRNG[948] = (LFSRcolor4[704]&LFSRcolor4[314]&LFSRcolor4[804]&LFSRcolor4[558]);
    BiasedRNG[949] = (LFSRcolor4[932]&LFSRcolor4[109]&LFSRcolor4[516]&LFSRcolor4[515]);
    BiasedRNG[950] = (LFSRcolor4[534]&LFSRcolor4[682]&LFSRcolor4[618]&LFSRcolor4[273]);
    BiasedRNG[951] = (LFSRcolor4[155]&LFSRcolor4[439]&LFSRcolor4[697]&LFSRcolor4[658]);
    BiasedRNG[952] = (LFSRcolor4[955]&LFSRcolor4[692]&LFSRcolor4[771]&LFSRcolor4[379]);
    BiasedRNG[953] = (LFSRcolor4[657]&LFSRcolor4[352]&LFSRcolor4[789]&LFSRcolor4[290]);
    BiasedRNG[954] = (LFSRcolor4[630]&LFSRcolor4[212]&LFSRcolor4[252]&LFSRcolor4[766]);
    BiasedRNG[955] = (LFSRcolor4[841]&LFSRcolor4[934]&LFSRcolor4[720]&LFSRcolor4[276]);
    BiasedRNG[956] = (LFSRcolor4[473]&LFSRcolor4[84]&LFSRcolor4[206]&LFSRcolor4[581]);
    BiasedRNG[957] = (LFSRcolor4[339]&LFSRcolor4[895]&LFSRcolor4[952]&LFSRcolor4[399]);
    BiasedRNG[958] = (LFSRcolor4[930]&LFSRcolor4[559]&LFSRcolor4[412]&LFSRcolor4[656]);
    BiasedRNG[959] = (LFSRcolor4[794]&LFSRcolor4[531]&LFSRcolor4[868]&LFSRcolor4[74]);
    BiasedRNG[960] = (LFSRcolor4[809]&LFSRcolor4[661]&LFSRcolor4[873]&LFSRcolor4[402]);
    BiasedRNG[961] = (LFSRcolor4[378]&LFSRcolor4[398]&LFSRcolor4[925]&LFSRcolor4[755]);
    BiasedRNG[962] = (LFSRcolor4[406]&LFSRcolor4[668]&LFSRcolor4[106]&LFSRcolor4[756]);
    BiasedRNG[963] = (LFSRcolor4[291]&LFSRcolor4[386]&LFSRcolor4[265]&LFSRcolor4[604]);
    BiasedRNG[964] = (LFSRcolor4[343]&LFSRcolor4[850]&LFSRcolor4[726]&LFSRcolor4[548]);
    BiasedRNG[965] = (LFSRcolor4[26]&LFSRcolor4[218]&LFSRcolor4[170]&LFSRcolor4[547]);
    BiasedRNG[966] = (LFSRcolor4[727]&LFSRcolor4[86]&LFSRcolor4[800]&LFSRcolor4[563]);
    BiasedRNG[967] = (LFSRcolor4[157]&LFSRcolor4[187]&LFSRcolor4[164]&LFSRcolor4[1]);
    BiasedRNG[968] = (LFSRcolor4[434]&LFSRcolor4[776]&LFSRcolor4[730]&LFSRcolor4[945]);
    BiasedRNG[969] = (LFSRcolor4[659]&LFSRcolor4[556]&LFSRcolor4[179]&LFSRcolor4[282]);
    BiasedRNG[970] = (LFSRcolor4[93]&LFSRcolor4[58]&LFSRcolor4[263]&LFSRcolor4[900]);
    BiasedRNG[971] = (LFSRcolor4[30]&LFSRcolor4[485]&LFSRcolor4[75]&LFSRcolor4[780]);
    BiasedRNG[972] = (LFSRcolor4[560]&LFSRcolor4[192]&LFSRcolor4[76]&LFSRcolor4[21]);
    BiasedRNG[973] = (LFSRcolor4[266]&LFSRcolor4[162]&LFSRcolor4[687]&LFSRcolor4[233]);
    BiasedRNG[974] = (LFSRcolor4[99]&LFSRcolor4[294]&LFSRcolor4[829]&LFSRcolor4[96]);
    BiasedRNG[975] = (LFSRcolor4[430]&LFSRcolor4[453]&LFSRcolor4[298]&LFSRcolor4[511]);
    BiasedRNG[976] = (LFSRcolor4[176]&LFSRcolor4[920]&LFSRcolor4[337]&LFSRcolor4[166]);
    BiasedRNG[977] = (LFSRcolor4[751]&LFSRcolor4[562]&LFSRcolor4[768]&LFSRcolor4[585]);
    BiasedRNG[978] = (LFSRcolor4[624]&LFSRcolor4[653]&LFSRcolor4[45]&LFSRcolor4[332]);
    BiasedRNG[979] = (LFSRcolor4[92]&LFSRcolor4[960]&LFSRcolor4[414]&LFSRcolor4[573]);
    BiasedRNG[980] = (LFSRcolor4[454]&LFSRcolor4[721]&LFSRcolor4[331]&LFSRcolor4[283]);
    BiasedRNG[981] = (LFSRcolor4[47]&LFSRcolor4[51]&LFSRcolor4[165]&LFSRcolor4[348]);
    BiasedRNG[982] = (LFSRcolor4[14]&LFSRcolor4[351]&LFSRcolor4[5]&LFSRcolor4[241]);
    BiasedRNG[983] = (LFSRcolor4[429]&LFSRcolor4[257]&LFSRcolor4[452]&LFSRcolor4[167]);
    BiasedRNG[984] = (LFSRcolor4[954]&LFSRcolor4[708]&LFSRcolor4[326]&LFSRcolor4[961]);
    BiasedRNG[985] = (LFSRcolor4[666]&LFSRcolor4[234]&LFSRcolor4[826]&LFSRcolor4[823]);
    BiasedRNG[986] = (LFSRcolor4[669]&LFSRcolor4[680]&LFSRcolor4[905]&LFSRcolor4[684]);
    BiasedRNG[987] = (LFSRcolor4[544]&LFSRcolor4[449]&LFSRcolor4[53]&LFSRcolor4[501]);
    BiasedRNG[988] = (LFSRcolor4[87]&LFSRcolor4[805]&LFSRcolor4[173]&LFSRcolor4[376]);
    BiasedRNG[989] = (LFSRcolor4[513]&LFSRcolor4[175]&LFSRcolor4[594]&LFSRcolor4[147]);
    BiasedRNG[990] = (LFSRcolor4[3]&LFSRcolor4[275]&LFSRcolor4[91]&LFSRcolor4[958]);
    BiasedRNG[991] = (LFSRcolor4[83]&LFSRcolor4[959]&LFSRcolor4[221]&LFSRcolor4[450]);
    BiasedRNG[992] = (LFSRcolor4[679]&LFSRcolor4[104]&LFSRcolor4[420]&LFSRcolor4[788]);
    BiasedRNG[993] = (LFSRcolor4[145]&LFSRcolor4[222]&LFSRcolor4[688]&LFSRcolor4[631]);
    BiasedRNG[994] = (LFSRcolor4[843]&LFSRcolor4[601]&LFSRcolor4[929]&LFSRcolor4[4]);
    BiasedRNG[995] = (LFSRcolor4[81]&LFSRcolor4[113]&LFSRcolor4[923]&LFSRcolor4[181]);
    BiasedRNG[996] = (LFSRcolor4[767]&LFSRcolor4[293]&LFSRcolor4[133]&LFSRcolor4[646]);
    BiasedRNG[997] = (LFSRcolor4[941]&LFSRcolor4[599]&LFSRcolor4[408]&LFSRcolor4[335]);
    BiasedRNG[998] = (LFSRcolor4[748]&LFSRcolor4[169]&LFSRcolor4[535]&LFSRcolor4[707]);
    BiasedRNG[999] = (LFSRcolor4[9]&LFSRcolor4[861]&LFSRcolor4[738]&LFSRcolor4[232]);
    BiasedRNG[1000] = (LFSRcolor4[595]&LFSRcolor4[518]&LFSRcolor4[23]&LFSRcolor4[411]);
    BiasedRNG[1001] = (LFSRcolor4[20]&LFSRcolor4[831]&LFSRcolor4[711]&LFSRcolor4[349]);
    BiasedRNG[1002] = (LFSRcolor4[191]&LFSRcolor4[72]&LFSRcolor4[719]&LFSRcolor4[931]);
    BiasedRNG[1003] = (LFSRcolor4[898]&LFSRcolor4[476]&LFSRcolor4[946]&LFSRcolor4[287]);
    BiasedRNG[1004] = (LFSRcolor4[225]&LFSRcolor4[253]&LFSRcolor4[61]&LFSRcolor4[285]);
    BiasedRNG[1005] = (LFSRcolor4[577]&LFSRcolor4[171]&LFSRcolor4[878]&LFSRcolor4[712]);
    BiasedRNG[1006] = (LFSRcolor4[608]&LFSRcolor4[640]&LFSRcolor4[949]&LFSRcolor4[937]);
    BiasedRNG[1007] = (LFSRcolor4[19]&LFSRcolor4[787]&LFSRcolor4[956]&LFSRcolor4[413]);
    BiasedRNG[1008] = (LFSRcolor4[838]&LFSRcolor4[64]&LFSRcolor4[551]&LFSRcolor4[345]);
    BiasedRNG[1009] = (LFSRcolor4[765]&LFSRcolor4[350]&LFSRcolor4[200]&LFSRcolor4[365]);
    BiasedRNG[1010] = (LFSRcolor4[675]&LFSRcolor4[862]&LFSRcolor4[88]&LFSRcolor4[670]);
    BiasedRNG[1011] = (LFSRcolor4[249]&LFSRcolor4[325]&LFSRcolor4[694]&LFSRcolor4[395]);
    BiasedRNG[1012] = (LFSRcolor4[231]&LFSRcolor4[567]&LFSRcolor4[299]&LFSRcolor4[469]);
    BiasedRNG[1013] = (LFSRcolor4[914]&LFSRcolor4[663]&LFSRcolor4[758]&LFSRcolor4[401]);
    BiasedRNG[1014] = (LFSRcolor4[210]&LFSRcolor4[681]&LFSRcolor4[305]&LFSRcolor4[79]);
    BiasedRNG[1015] = (LFSRcolor4[590]&LFSRcolor4[153]&LFSRcolor4[899]&LFSRcolor4[286]);
    BiasedRNG[1016] = (LFSRcolor4[443]&LFSRcolor4[609]&LFSRcolor4[159]&LFSRcolor4[364]);
    BiasedRNG[1017] = (LFSRcolor4[17]&LFSRcolor4[509]&LFSRcolor4[654]&LFSRcolor4[46]);
    BiasedRNG[1018] = (LFSRcolor4[860]&LFSRcolor4[696]&LFSRcolor4[433]&LFSRcolor4[129]);
    BiasedRNG[1019] = (LFSRcolor4[368]&LFSRcolor4[722]&LFSRcolor4[655]&LFSRcolor4[371]);
    BiasedRNG[1020] = (LFSRcolor4[82]&LFSRcolor4[651]&LFSRcolor4[366]&LFSRcolor4[397]);
    BiasedRNG[1021] = (LFSRcolor4[367]&LFSRcolor4[297]&LFSRcolor4[520]&LFSRcolor4[321]);
    BiasedRNG[1022] = (LFSRcolor4[143]&LFSRcolor4[703]&LFSRcolor4[842]&LFSRcolor4[174]);
    BiasedRNG[1023] = (LFSRcolor4[405]&LFSRcolor4[953]&LFSRcolor4[818]&LFSRcolor4[533]);
    BiasedRNG[1024] = (LFSRcolor4[415]&LFSRcolor4[246]&LFSRcolor4[880]&LFSRcolor4[922]);
    BiasedRNG[1025] = (LFSRcolor4[110]&LFSRcolor4[16]&LFSRcolor4[270]&LFSRcolor4[596]);
    BiasedRNG[1026] = (LFSRcolor4[723]&LFSRcolor4[614]&LFSRcolor4[665]&LFSRcolor4[128]);
    BiasedRNG[1027] = (LFSRcolor4[833]&LFSRcolor4[360]&LFSRcolor4[309]&LFSRcolor4[370]);
    BiasedRNG[1028] = (LFSRcolor4[32]&LFSRcolor4[38]&LFSRcolor4[791]&LFSRcolor4[565]);
    BiasedRNG[1029] = (LFSRcolor4[334]&LFSRcolor4[813]&LFSRcolor4[936]&LFSRcolor4[517]);
    BiasedRNG[1030] = (LFSRcolor4[571]&LFSRcolor4[820]&LFSRcolor4[744]&LFSRcolor4[499]);
    BiasedRNG[1031] = (LFSRcolor4[570]&LFSRcolor4[223]&LFSRcolor4[588]&LFSRcolor4[781]);
    BiasedRNG[1032] = (LFSRcolor4[444]&LFSRcolor4[418]&LFSRcolor4[136]&LFSRcolor4[619]);
    BiasedRNG[1033] = (LFSRcolor4[341]&LFSRcolor4[769]&LFSRcolor4[706]&LFSRcolor4[602]);
    BiasedRNG[1034] = (LFSRcolor4[671]&LFSRcolor4[146]&LFSRcolor4[477]&LFSRcolor4[492]);
    BiasedRNG[1035] = (LFSRcolor4[950]&LFSRcolor4[94]&LFSRcolor4[392]&LFSRcolor4[114]);
    BiasedRNG[1036] = (LFSRcolor4[825]&LFSRcolor4[417]&LFSRcolor4[267]&LFSRcolor4[582]);
    BiasedRNG[1037] = (LFSRcolor4[795]&LFSRcolor4[484]&LFSRcolor4[388]&LFSRcolor4[728]);
    BiasedRNG[1038] = (LFSRcolor4[903]&LFSRcolor4[667]&LFSRcolor4[248]&LFSRcolor4[884]);
    BiasedRNG[1039] = (LFSRcolor4[310]&LFSRcolor4[390]&LFSRcolor4[85]&LFSRcolor4[881]);
    BiasedRNG[1040] = (LFSRcolor4[828]&LFSRcolor4[461]&LFSRcolor4[752]&LFSRcolor4[316]);
    BiasedRNG[1041] = (LFSRcolor4[36]&LFSRcolor4[662]&LFSRcolor4[793]&LFSRcolor4[268]);
    BiasedRNG[1042] = (LFSRcolor4[538]&LFSRcolor4[944]&LFSRcolor4[628]&LFSRcolor4[564]);
    BiasedRNG[1043] = (LFSRcolor4[824]&LFSRcolor4[228]&LFSRcolor4[42]&LFSRcolor4[396]);
    BiasedRNG[1044] = (LFSRcolor4[897]&LFSRcolor4[13]&LFSRcolor4[190]&LFSRcolor4[203]);
    BiasedRNG[1045] = (LFSRcolor4[242]&LFSRcolor4[633]&LFSRcolor4[52]&LFSRcolor4[480]);
    BiasedRNG[1046] = (LFSRcolor4[889]&LFSRcolor4[933]&LFSRcolor4[759]&LFSRcolor4[834]);
    BiasedRNG[1047] = (LFSRcolor4[119]&LFSRcolor4[199]&LFSRcolor4[435]&LFSRcolor4[864]);
    BiasedRNG[1048] = (LFSRcolor4[606]&LFSRcolor4[195]&LFSRcolor4[909]&LFSRcolor4[948]);
    BiasedRNG[1049] = (LFSRcolor4[425]&LFSRcolor4[229]&LFSRcolor4[918]&LFSRcolor4[416]);
    BiasedRNG[1050] = (LFSRcolor4[753]&LFSRcolor4[172]&LFSRcolor4[437]&LFSRcolor4[70]);
    BiasedRNG[1051] = (LFSRcolor4[322]&LFSRcolor4[189]&LFSRcolor4[629]&LFSRcolor4[892]);
    BiasedRNG[1052] = (LFSRcolor4[885]&LFSRcolor4[238]&LFSRcolor4[693]&LFSRcolor4[219]);
    BiasedRNG[1053] = (LFSRcolor4[134]&LFSRcolor4[796]&LFSRcolor4[964]&LFSRcolor4[916]);
    BiasedRNG[1054] = (LFSRcolor4[122]&LFSRcolor4[307]&LFSRcolor4[63]&LFSRcolor4[890]);
    BiasedRNG[1055] = (LFSRcolor4[866]&LFSRcolor4[910]&LFSRcolor4[886]&LFSRcolor4[734]);
    BiasedRNG[1056] = (LFSRcolor4[319]&LFSRcolor4[186]&LFSRcolor4[846]&LFSRcolor4[288]);
    BiasedRNG[1057] = (LFSRcolor4[141]&LFSRcolor4[185]&LFSRcolor4[139]&LFSRcolor4[621]);
    BiasedRNG[1058] = (LFSRcolor4[56]&LFSRcolor4[725]&LFSRcolor4[354]&LFSRcolor4[150]);
    BiasedRNG[1059] = (LFSRcolor4[495]&LFSRcolor4[460]&LFSRcolor4[344]&LFSRcolor4[216]);
    BiasedRNG[1060] = (LFSRcolor4[705]&LFSRcolor4[747]&LFSRcolor4[552]&LFSRcolor4[346]);
    BiasedRNG[1061] = (LFSRcolor4[647]&LFSRcolor4[940]&LFSRcolor4[68]&LFSRcolor4[852]);
    BiasedRNG[1062] = (LFSRcolor4[695]&LFSRcolor4[514]&LFSRcolor4[31]&LFSRcolor4[962]);
    BiasedRNG[1063] = (LFSRcolor4[851]&LFSRcolor4[424]&LFSRcolor4[7]&LFSRcolor4[124]);
    BiasedRNG[1064] = (LFSRcolor4[342]&LFSRcolor4[904]&LFSRcolor4[338]&LFSRcolor4[530]);
    BiasedRNG[1065] = (LFSRcolor4[394]&LFSRcolor4[152]&LFSRcolor4[774]&LFSRcolor4[462]);
    BiasedRNG[1066] = (LFSRcolor4[269]&LFSRcolor4[330]&LFSRcolor4[154]&LFSRcolor4[357]);
    BiasedRNG[1067] = (LFSRcolor4[131]&LFSRcolor4[812]&LFSRcolor4[553]&LFSRcolor4[71]);
    BiasedRNG[1068] = (LFSRcolor4[2]&LFSRcolor4[876]&LFSRcolor4[54]&LFSRcolor4[80]);
    BiasedRNG[1069] = (LFSRcolor4[888]&LFSRcolor4[732]&LFSRcolor4[523]&LFSRcolor4[0]);
    BiasedRNG[1070] = (LFSRcolor4[24]&LFSRcolor4[951]&LFSRcolor4[432]&LFSRcolor4[112]);
    BiasedRNG[1071] = (LFSRcolor4[121]&LFSRcolor4[363]&LFSRcolor4[105]&LFSRcolor4[407]);
    BiasedRNG[1072] = (LFSRcolor4[915]&LFSRcolor4[468]&LFSRcolor4[935]&LFSRcolor4[481]);
    BiasedRNG[1073] = (LFSRcolor4[302]&LFSRcolor4[634]&LFSRcolor4[235]&LFSRcolor4[500]);
    BiasedRNG[1074] = (LFSRcolor4[494]&LFSRcolor4[537]&LFSRcolor4[912]&LFSRcolor4[279]);
    BiasedRNG[1075] = (LFSRcolor4[464]&LFSRcolor4[750]&LFSRcolor4[478]&LFSRcolor4[592]);
    BiasedRNG[1076] = (LFSRcolor4[377]&LFSRcolor4[815]&LFSRcolor4[50]&LFSRcolor4[130]);
    BiasedRNG[1077] = (LFSRcolor4[635]&LFSRcolor4[431]&LFSRcolor4[605]&LFSRcolor4[569]);
    BiasedRNG[1078] = (LFSRcolor4[384]&LFSRcolor4[158]&LFSRcolor4[616]&LFSRcolor4[782]);
    BiasedRNG[1079] = (LFSRcolor4[854]&LFSRcolor4[183]&LFSRcolor4[736]&LFSRcolor4[214]);
    BiasedRNG[1080] = (LFSRcolor4[650]&LFSRcolor4[798]&LFSRcolor4[893]&LFSRcolor4[436]);
    BiasedRNG[1081] = (LFSRcolor4[710]&LFSRcolor4[906]&LFSRcolor4[230]&LFSRcolor4[278]);
    BiasedRNG[1082] = (LFSRcolor4[625]&LFSRcolor4[372]&LFSRcolor4[48]&LFSRcolor4[479]);
    BiasedRNG[1083] = (LFSRcolor4[474]&LFSRcolor4[942]&LFSRcolor4[506]&LFSRcolor4[817]);
    BiasedRNG[1084] = (LFSRcolor4[510]&LFSRcolor4[938]&LFSRcolor4[690]&LFSRcolor4[549]);
    BiasedRNG[1085] = (LFSRcolor4[689]&LFSRcolor4[57]&LFSRcolor4[579]&LFSRcolor4[78]);
    BiasedRNG[1086] = (LFSRcolor4[632]&LFSRcolor4[400]&LFSRcolor4[691]&LFSRcolor4[593]);
    BiasedRNG[1087] = (LFSRcolor4[126]&LFSRcolor4[853]&LFSRcolor4[856]&LFSRcolor4[963]);
    BiasedRNG[1088] = (LFSRcolor4[410]&LFSRcolor4[490]&LFSRcolor4[701]&LFSRcolor4[69]);
    BiasedRNG[1089] = (LFSRcolor4[566]&LFSRcolor4[957]&LFSRcolor4[422]&LFSRcolor4[802]);
    BiasedRNG[1090] = (LFSRcolor4[441]&LFSRcolor4[123]&LFSRcolor4[296]&LFSRcolor4[116]);
    BiasedRNG[1091] = (LFSRcolor4[674]&LFSRcolor4[317]&LFSRcolor4[587]&LFSRcolor4[896]);
    BiasedRNG[1092] = (LFSRcolor4[227]&LFSRcolor4[118]&LFSRcolor4[743]&LFSRcolor4[550]);
    BiasedRNG[1093] = (LFSRcolor4[254]&LFSRcolor4[472]&LFSRcolor4[177]&LFSRcolor4[323]);
    BiasedRNG[1094] = (LFSRcolor4[749]&LFSRcolor4[65]&LFSRcolor4[336]&LFSRcolor4[115]);
    BiasedRNG[1095] = (LFSRcolor4[790]&LFSRcolor4[641]&LFSRcolor4[939]&LFSRcolor4[869]);
    BiasedRNG[1096] = (LFSRcolor4[324]&LFSRcolor4[913]&LFSRcolor4[735]&LFSRcolor4[44]);
    BiasedRNG[1097] = (LFSRcolor4[672]&LFSRcolor4[645]&LFSRcolor4[636]&LFSRcolor4[764]);
    BiasedRNG[1098] = (LFSRcolor4[643]&LFSRcolor4[649]&LFSRcolor4[327]&LFSRcolor4[369]);
    BiasedRNG[1099] = (LFSRcolor4[883]&LFSRcolor4[584]&LFSRcolor4[882]&LFSRcolor4[274]);
    BiasedRNG[1100] = (LFSRcolor4[729]&LFSRcolor4[642]&LFSRcolor4[847]&LFSRcolor4[801]);
    BiasedRNG[1101] = (LFSRcolor4[814]&LFSRcolor4[965]&LFSRcolor4[493]&LFSRcolor4[620]);
    BiasedRNG[1102] = (LFSRcolor4[120]&LFSRcolor4[127]&LFSRcolor4[180]&LFSRcolor4[786]);
    BiasedRNG[1103] = (LFSRcolor4[426]&LFSRcolor4[557]&LFSRcolor4[677]&LFSRcolor4[508]);
    BiasedRNG[1104] = (LFSRcolor4[389]&LFSRcolor4[37]&LFSRcolor4[193]&LFSRcolor4[362]);
    BiasedRNG[1105] = (LFSRcolor4[745]&LFSRcolor4[117]&LFSRcolor4[924]&LFSRcolor4[356]);
    BiasedRNG[1106] = (LFSRcolor4[580]&LFSRcolor4[746]&LFSRcolor4[11]&LFSRcolor4[315]);
    BiasedRNG[1107] = (LFSRcolor4[311]&LFSRcolor4[521]&LFSRcolor4[197]&LFSRcolor4[529]);
    BiasedRNG[1108] = (LFSRcolor4[575]&LFSRcolor4[810]&LFSRcolor4[381]&LFSRcolor4[739]);
    BiasedRNG[1109] = (LFSRcolor4[149]&LFSRcolor4[304]&LFSRcolor4[446]&LFSRcolor4[639]);
    BiasedRNG[1110] = (LFSRcolor4[610]&LFSRcolor4[73]&LFSRcolor4[442]&LFSRcolor4[840]);
    BiasedRNG[1111] = (LFSRcolor4[329]&LFSRcolor4[683]&LFSRcolor4[803]&LFSRcolor4[188]);
    BiasedRNG[1112] = (LFSRcolor4[773]&LFSRcolor4[161]&LFSRcolor4[102]&LFSRcolor4[427]);
    BiasedRNG[1113] = (LFSRcolor4[260]&LFSRcolor4[28]&LFSRcolor4[148]&LFSRcolor4[29]);
    BiasedRNG[1114] = (LFSRcolor4[97]&LFSRcolor4[201]&LFSRcolor4[757]&LFSRcolor4[644]);
    BiasedRNG[1115] = (LFSRcolor4[911]&LFSRcolor4[733]&LFSRcolor4[507]&LFSRcolor4[226]);
    BiasedRNG[1116] = (LFSRcolor4[542]&LFSRcolor4[204]&LFSRcolor4[489]&LFSRcolor4[358]);
    BiasedRNG[1117] = (LFSRcolor4[907]&LFSRcolor4[312]&LFSRcolor4[849]&LFSRcolor4[522]);
    BiasedRNG[1118] = (LFSRcolor4[772]&LFSRcolor4[244]&LFSRcolor4[43]&LFSRcolor4[373]);
    BiasedRNG[1119] = (LFSRcolor4[545]&LFSRcolor4[385]&LFSRcolor4[447]&LFSRcolor4[718]);
    BiasedRNG[1120] = (LFSRcolor4[613]&LFSRcolor4[470]&LFSRcolor4[243]&LFSRcolor4[504]);
    BiasedRNG[1121] = (LFSRcolor4[528]&LFSRcolor4[33]&LFSRcolor4[837]&LFSRcolor4[740]);
    BiasedRNG[1122] = (LFSRcolor4[258]&LFSRcolor4[445]&LFSRcolor4[194]&LFSRcolor4[41]);
    BiasedRNG[1123] = (LFSRcolor4[870]&LFSRcolor4[716]&LFSRcolor4[717]&LFSRcolor4[660]);
    BiasedRNG[1124] = (LFSRcolor4[301]&LFSRcolor4[699]&LFSRcolor4[168]&LFSRcolor4[208]);
    BiasedRNG[1125] = (LFSRcolor4[779]&LFSRcolor4[328]&LFSRcolor4[40]&LFSRcolor4[830]);
    BiasedRNG[1126] = (LFSRcolor4[465]&LFSRcolor4[626]&LFSRcolor4[15]&LFSRcolor4[778]);
    BiasedRNG[1127] = (LFSRcolor4[318]&LFSRcolor4[347]&LFSRcolor4[277]&LFSRcolor4[160]);
    BiasedRNG[1128] = (LFSRcolor4[554]&LFSRcolor4[419]&LFSRcolor4[497]&LFSRcolor4[617]);
    BiasedRNG[1129] = (LFSRcolor4[163]&LFSRcolor4[519]&LFSRcolor4[355]&LFSRcolor4[428]);
    BiasedRNG[1130] = (LFSRcolor4[12]&LFSRcolor4[487]&LFSRcolor4[101]&LFSRcolor4[289]);
    BiasedRNG[1131] = (LFSRcolor4[423]&LFSRcolor4[555]&LFSRcolor4[488]&LFSRcolor4[103]);
    BiasedRNG[1132] = (LFSRcolor4[333]&LFSRcolor4[811]&LFSRcolor4[539]&LFSRcolor4[456]);
    BiasedRNG[1133] = (LFSRcolor4[211]&LFSRcolor4[855]&LFSRcolor4[471]&LFSRcolor4[709]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

//Generate the ILA for data collection:
ila_0 ILAinst(.clk(sample_clk),.probe0(run),.probe1(solution_flag),.probe2(failure),.probe3(counter[37:0]));

//Instantiate VIO:
vio_0 VIOinst (.clk(sample_clk),.probe_out0(reset),.probe_out1(solution_set[31:0]));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule