//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [23:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [827:0] LFSRcolor0;
wire [1011:0] LFSRcolor1;
wire [735:0] LFSRcolor2;
wire [137:0] LFSRcolor3;
wire [551:0] LFSRcolor4;
reg [657:0] BiasedRNG;       //For I=+/-1 cases
reg [493:0] UnbiasedRNG;   //For I=0 cases
reg [0:1187] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[384] = 1'b1;
initial m[531] = 1'b0;
initial m[541] = 1'b1;
initial m[556] = 1'b1;
initial m[576] = 1'b1;
initial m[601] = 1'b1;
initial m[631] = 1'b1;
initial m[666] = 1'b1;
initial m[706] = 1'b0;
initial m[751] = 1'b1;
initial m[801] = 1'b0;
initial m[856] = 1'b0;
initial m[911] = 1'b0;
initial m[961] = 1'b1;
initial m[1006] = 1'b0;
initial m[1046] = 1'b0;
initial m[1081] = 1'b0;
initial m[1111] = 1'b0;
initial m[1136] = 1'b1;
initial m[1156] = 1'b1;
initial m[1171] = 1'b1;
initial m[1181] = 1'b1;
initial m[1186] = 1'b1;
initial m[1187] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[530] = 1'b0;
initial m[540] = 1'b0;
initial m[555] = 1'b0;
initial m[575] = 1'b0;
initial m[600] = 1'b0;
initial m[630] = 1'b0;
initial m[665] = 1'b0;
initial m[705] = 1'b0;
initial m[750] = 1'b0;
initial m[800] = 1'b0;
initial m[855] = 1'b0;
initial m[858] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR0_11(.LFSRregister(LFSRcolor0[551:506]),.clk(sample_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR0_12(.LFSRregister(LFSRcolor0[597:552]),.clk(sample_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR0_13(.LFSRregister(LFSRcolor0[643:598]),.clk(sample_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR0_14(.LFSRregister(LFSRcolor0[689:644]),.clk(sample_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR0_15(.LFSRregister(LFSRcolor0[735:690]),.clk(sample_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR0_16(.LFSRregister(LFSRcolor0[781:736]),.clk(sample_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR0_17(.LFSRregister(LFSRcolor0[827:782]),.clk(sample_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR1_15(.LFSRregister(LFSRcolor1[735:690]),.clk(color0_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR1_16(.LFSRregister(LFSRcolor1[781:736]),.clk(color0_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR1_17(.LFSRregister(LFSRcolor1[827:782]),.clk(color0_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR1_18(.LFSRregister(LFSRcolor1[873:828]),.clk(color0_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR1_19(.LFSRregister(LFSRcolor1[919:874]),.clk(color0_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR1_20(.LFSRregister(LFSRcolor1[965:920]),.clk(color0_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR1_21(.LFSRregister(LFSRcolor1[1011:966]),.clk(color0_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b0011001000010001001111001110101111011111000110)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b0101000110100000010101001000010000101101100110)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b1110011010010011001010111010100101111111100000)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b1001111000010100100001100010110000001111101011)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b0011101001111100110111000000010000101100111110)) LFSR2_11(.LFSRregister(LFSRcolor2[551:506]),.clk(color1_clk));
lfsr #(.seed(46'b1010111010001100001100010110010011100100101100)) LFSR2_12(.LFSRregister(LFSRcolor2[597:552]),.clk(color1_clk));
lfsr #(.seed(46'b1101010000110001000001011010110100010000110101)) LFSR2_13(.LFSRregister(LFSRcolor2[643:598]),.clk(color1_clk));
lfsr #(.seed(46'b0111111000001001010001100011001110110101101001)) LFSR2_14(.LFSRregister(LFSRcolor2[689:644]),.clk(color1_clk));
lfsr #(.seed(46'b0111011110101100100001111000001001111001010010)) LFSR2_15(.LFSRregister(LFSRcolor2[735:690]),.clk(color1_clk));
lfsr #(.seed(46'b0110010001011011111100000000110011011110000100)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b1100101101001001110010011101110000001110111111)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b1110010100000011100111110011000001001000000101)) LFSR3_2(.LFSRregister(LFSRcolor3[137:92]),.clk(color2_clk));
lfsr #(.seed(46'b1100111110111110000101110101010111111010101000)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1101101000110111001110111111011011100011111101)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1011100111101011110000001101111100001111100011)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b1000011101010100110111010000000111000111010111)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b0011001001101100101110110001011100100100110000)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b0011110010011101000111111110100110110100101000)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b1100000100011100010111001011000000101100110100)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b1001101001101101001001111001110100110001100010)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));
lfsr #(.seed(46'b1000000000001101011011010100000001101001001111)) LFSR4_8(.LFSRregister(LFSRcolor4[413:368]),.clk(color3_clk));
lfsr #(.seed(46'b1000011000100000010011100100110100001010000001)) LFSR4_9(.LFSRregister(LFSRcolor4[459:414]),.clk(color3_clk));
lfsr #(.seed(46'b0101000011110010010110011011111101010101011010)) LFSR4_10(.LFSRregister(LFSRcolor4[505:460]),.clk(color3_clk));
lfsr #(.seed(46'b0011111001110010110000110100101000000000100010)) LFSR4_11(.LFSRregister(LFSRcolor4[551:506]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 0;
initial m[1] = 0;
initial m[2] = 1;
initial m[3] = 1;
initial m[4] = 1;
initial m[5] = 0;
initial m[6] = 1;
initial m[7] = 0;
initial m[8] = 0;
initial m[9] = 1;
initial m[10] = 1;
initial m[11] = 1;
initial m[12] = 0;
initial m[13] = 1;
initial m[14] = 0;
initial m[15] = 0;
initial m[16] = 1;
initial m[17] = 0;
initial m[18] = 1;
initial m[19] = 1;
initial m[20] = 0;
initial m[21] = 1;
initial m[22] = 1;
initial m[23] = 1;
initial m[24] = 1;
initial m[25] = 1;
initial m[26] = 0;
initial m[27] = 0;
initial m[28] = 1;
initial m[29] = 0;
initial m[30] = 1;
initial m[31] = 0;
initial m[32] = 1;
initial m[33] = 0;
initial m[34] = 1;
initial m[35] = 0;
initial m[36] = 1;
initial m[37] = 1;
initial m[38] = 0;
initial m[39] = 0;
initial m[40] = 1;
initial m[41] = 1;
initial m[42] = 0;
initial m[43] = 0;
initial m[44] = 0;
initial m[45] = 0;
initial m[46] = 1;
initial m[47] = 1;
initial m[48] = 0;
initial m[49] = 0;
initial m[50] = 1;
initial m[51] = 1;
initial m[52] = 1;
initial m[53] = 1;
initial m[54] = 0;
initial m[55] = 0;
initial m[56] = 0;
initial m[57] = 0;
initial m[58] = 1;
initial m[59] = 1;
initial m[60] = 1;
initial m[61] = 1;
initial m[62] = 0;
initial m[63] = 1;
initial m[64] = 0;
initial m[65] = 1;
initial m[66] = 1;
initial m[67] = 1;
initial m[68] = 0;
initial m[69] = 1;
initial m[70] = 1;
initial m[71] = 1;
initial m[72] = 0;
initial m[73] = 0;
initial m[74] = 0;
initial m[75] = 1;
initial m[76] = 1;
initial m[77] = 1;
initial m[78] = 1;
initial m[79] = 0;
initial m[80] = 0;
initial m[81] = 0;
initial m[82] = 1;
initial m[83] = 0;
initial m[84] = 1;
initial m[85] = 0;
initial m[86] = 1;
initial m[87] = 1;
initial m[88] = 0;
initial m[89] = 0;
initial m[90] = 1;
initial m[91] = 1;
initial m[92] = 0;
initial m[93] = 1;
initial m[94] = 0;
initial m[95] = 1;
initial m[96] = 1;
initial m[97] = 0;
initial m[98] = 1;
initial m[99] = 1;
initial m[100] = 1;
initial m[101] = 1;
initial m[102] = 1;
initial m[103] = 1;
initial m[104] = 1;
initial m[105] = 0;
initial m[106] = 0;
initial m[107] = 0;
initial m[108] = 1;
initial m[109] = 0;
initial m[110] = 1;
initial m[111] = 1;
initial m[112] = 1;
initial m[113] = 1;
initial m[114] = 1;
initial m[115] = 0;
initial m[116] = 1;
initial m[117] = 0;
initial m[118] = 1;
initial m[119] = 0;
initial m[120] = 1;
initial m[121] = 1;
initial m[122] = 1;
initial m[123] = 1;
initial m[124] = 0;
initial m[125] = 1;
initial m[126] = 1;
initial m[127] = 0;
initial m[128] = 0;
initial m[129] = 0;
initial m[130] = 1;
initial m[131] = 1;
initial m[132] = 1;
initial m[133] = 1;
initial m[134] = 0;
initial m[135] = 0;
initial m[136] = 1;
initial m[137] = 1;
initial m[138] = 1;
initial m[139] = 1;
initial m[140] = 0;
initial m[141] = 0;
initial m[142] = 1;
initial m[143] = 0;
initial m[144] = 1;
initial m[145] = 1;
initial m[146] = 0;
initial m[147] = 1;
initial m[148] = 1;
initial m[149] = 0;
initial m[150] = 1;
initial m[151] = 1;
initial m[152] = 1;
initial m[153] = 1;
initial m[154] = 1;
initial m[155] = 0;
initial m[156] = 0;
initial m[157] = 1;
initial m[158] = 0;
initial m[159] = 0;
initial m[160] = 1;
initial m[161] = 1;
initial m[162] = 1;
initial m[163] = 0;
initial m[164] = 1;
initial m[165] = 1;
initial m[166] = 1;
initial m[167] = 1;
initial m[168] = 0;
initial m[169] = 1;
initial m[170] = 1;
initial m[171] = 1;
initial m[172] = 0;
initial m[173] = 1;
initial m[174] = 0;
initial m[175] = 0;
initial m[176] = 1;
initial m[177] = 0;
initial m[178] = 1;
initial m[179] = 0;
initial m[180] = 0;
initial m[181] = 1;
initial m[182] = 0;
initial m[183] = 0;
initial m[184] = 0;
initial m[185] = 1;
initial m[186] = 1;
initial m[187] = 0;
initial m[188] = 0;
initial m[189] = 0;
initial m[190] = 1;
initial m[191] = 1;
initial m[192] = 1;
initial m[193] = 0;
initial m[194] = 0;
initial m[195] = 1;
initial m[196] = 0;
initial m[197] = 0;
initial m[198] = 1;
initial m[199] = 1;
initial m[200] = 0;
initial m[201] = 1;
initial m[202] = 0;
initial m[203] = 1;
initial m[204] = 0;
initial m[205] = 0;
initial m[206] = 1;
initial m[207] = 0;
initial m[208] = 1;
initial m[209] = 0;
initial m[210] = 1;
initial m[211] = 0;
initial m[212] = 0;
initial m[213] = 1;
initial m[214] = 0;
initial m[215] = 0;
initial m[216] = 1;
initial m[217] = 0;
initial m[218] = 1;
initial m[219] = 0;
initial m[220] = 0;
initial m[221] = 1;
initial m[222] = 0;
initial m[223] = 0;
initial m[224] = 0;
initial m[225] = 1;
initial m[226] = 1;
initial m[227] = 0;
initial m[228] = 0;
initial m[229] = 0;
initial m[230] = 0;
initial m[231] = 0;
initial m[232] = 1;
initial m[233] = 0;
initial m[234] = 1;
initial m[235] = 0;
initial m[236] = 1;
initial m[237] = 1;
initial m[238] = 1;
initial m[239] = 1;
initial m[240] = 1;
initial m[241] = 0;
initial m[242] = 1;
initial m[243] = 0;
initial m[244] = 1;
initial m[245] = 1;
initial m[246] = 0;
initial m[247] = 0;
initial m[248] = 1;
initial m[249] = 1;
initial m[250] = 1;
initial m[251] = 0;
initial m[252] = 1;
initial m[253] = 0;
initial m[254] = 0;
initial m[255] = 0;
initial m[256] = 0;
initial m[257] = 1;
initial m[258] = 1;
initial m[259] = 1;
initial m[260] = 0;
initial m[261] = 0;
initial m[262] = 1;
initial m[263] = 1;
initial m[264] = 0;
initial m[265] = 0;
initial m[266] = 0;
initial m[267] = 1;
initial m[268] = 0;
initial m[269] = 0;
initial m[270] = 0;
initial m[271] = 0;
initial m[272] = 1;
initial m[273] = 0;
initial m[274] = 0;
initial m[275] = 1;
initial m[276] = 0;
initial m[277] = 1;
initial m[278] = 0;
initial m[279] = 0;
initial m[280] = 1;
initial m[281] = 1;
initial m[282] = 0;
initial m[283] = 1;
initial m[284] = 0;
initial m[285] = 0;
initial m[286] = 1;
initial m[287] = 0;
initial m[288] = 1;
initial m[289] = 0;
initial m[290] = 0;
initial m[291] = 0;
initial m[292] = 1;
initial m[293] = 1;
initial m[294] = 0;
initial m[295] = 0;
initial m[296] = 0;
initial m[297] = 1;
initial m[298] = 0;
initial m[299] = 0;
initial m[300] = 0;
initial m[301] = 1;
initial m[302] = 1;
initial m[303] = 0;
initial m[304] = 1;
initial m[305] = 0;
initial m[306] = 1;
initial m[307] = 0;
initial m[308] = 1;
initial m[309] = 0;
initial m[310] = 0;
initial m[311] = 0;
initial m[312] = 1;
initial m[313] = 1;
initial m[314] = 1;
initial m[315] = 0;
initial m[316] = 1;
initial m[317] = 0;
initial m[318] = 0;
initial m[319] = 1;
initial m[320] = 0;
initial m[321] = 1;
initial m[322] = 1;
initial m[323] = 1;
initial m[324] = 1;
initial m[325] = 1;
initial m[326] = 0;
initial m[327] = 1;
initial m[328] = 0;
initial m[329] = 0;
initial m[330] = 1;
initial m[331] = 1;
initial m[332] = 0;
initial m[333] = 1;
initial m[334] = 0;
initial m[335] = 0;
initial m[336] = 0;
initial m[337] = 1;
initial m[338] = 0;
initial m[339] = 1;
initial m[340] = 1;
initial m[341] = 1;
initial m[342] = 1;
initial m[343] = 1;
initial m[344] = 1;
initial m[345] = 1;
initial m[346] = 0;
initial m[347] = 0;
initial m[348] = 1;
initial m[349] = 1;
initial m[350] = 0;
initial m[351] = 1;
initial m[352] = 1;
initial m[353] = 1;
initial m[354] = 1;
initial m[355] = 1;
initial m[356] = 0;
initial m[357] = 1;
initial m[358] = 1;
initial m[359] = 1;
initial m[360] = 1;
initial m[361] = 1;
initial m[362] = 0;
initial m[363] = 1;
initial m[364] = 1;
initial m[365] = 0;
initial m[366] = 1;
initial m[367] = 0;
initial m[368] = 0;
initial m[369] = 0;
initial m[370] = 1;
initial m[371] = 1;
initial m[372] = 0;
initial m[373] = 0;
initial m[374] = 0;
initial m[375] = 0;
initial m[376] = 1;
initial m[377] = 0;
initial m[378] = 0;
initial m[379] = 0;
initial m[380] = 1;
initial m[381] = 1;
initial m[382] = 0;
initial m[383] = 1;
initial m[385] = 0;
initial m[386] = 1;
initial m[387] = 1;
initial m[388] = 1;
initial m[389] = 0;
initial m[390] = 0;
initial m[391] = 1;
initial m[392] = 0;
initial m[393] = 1;
initial m[394] = 0;
initial m[395] = 1;
initial m[396] = 1;
initial m[397] = 1;
initial m[398] = 1;
initial m[399] = 1;
initial m[400] = 1;
initial m[401] = 0;
initial m[402] = 1;
initial m[403] = 0;
initial m[404] = 1;
initial m[405] = 0;
initial m[406] = 0;
initial m[407] = 0;
initial m[408] = 1;
initial m[409] = 0;
initial m[410] = 1;
initial m[411] = 0;
initial m[412] = 1;
initial m[413] = 1;
initial m[414] = 1;
initial m[415] = 0;
initial m[416] = 0;
initial m[417] = 1;
initial m[418] = 1;
initial m[419] = 0;
initial m[420] = 1;
initial m[421] = 0;
initial m[422] = 0;
initial m[423] = 1;
initial m[424] = 1;
initial m[425] = 0;
initial m[426] = 1;
initial m[427] = 1;
initial m[428] = 0;
initial m[429] = 0;
initial m[430] = 0;
initial m[431] = 1;
initial m[432] = 0;
initial m[433] = 0;
initial m[434] = 1;
initial m[435] = 1;
initial m[436] = 1;
initial m[437] = 0;
initial m[438] = 1;
initial m[439] = 1;
initial m[440] = 1;
initial m[441] = 0;
initial m[442] = 0;
initial m[443] = 0;
initial m[444] = 1;
initial m[445] = 0;
initial m[446] = 0;
initial m[447] = 0;
initial m[448] = 0;
initial m[449] = 0;
initial m[450] = 0;
initial m[451] = 1;
initial m[452] = 1;
initial m[453] = 1;
initial m[454] = 0;
initial m[455] = 0;
initial m[456] = 0;
initial m[457] = 1;
initial m[458] = 1;
initial m[459] = 1;
initial m[460] = 0;
initial m[461] = 0;
initial m[462] = 0;
initial m[463] = 1;
initial m[464] = 0;
initial m[465] = 1;
initial m[466] = 1;
initial m[467] = 0;
initial m[468] = 0;
initial m[469] = 0;
initial m[470] = 0;
initial m[471] = 0;
initial m[472] = 1;
initial m[473] = 1;
initial m[474] = 1;
initial m[475] = 1;
initial m[476] = 1;
initial m[477] = 1;
initial m[478] = 1;
initial m[479] = 1;
initial m[480] = 1;
initial m[481] = 1;
initial m[482] = 1;
initial m[483] = 1;
initial m[484] = 0;
initial m[485] = 1;
initial m[486] = 0;
initial m[487] = 0;
initial m[488] = 0;
initial m[489] = 1;
initial m[490] = 1;
initial m[491] = 1;
initial m[492] = 1;
initial m[493] = 0;
initial m[494] = 1;
initial m[495] = 1;
initial m[496] = 1;
initial m[497] = 1;
initial m[498] = 1;
initial m[499] = 0;
initial m[500] = 0;
initial m[501] = 1;
initial m[502] = 0;
initial m[503] = 1;
initial m[504] = 0;
initial m[505] = 0;
initial m[506] = 0;
initial m[507] = 1;
initial m[508] = 1;
initial m[509] = 1;
initial m[510] = 0;
initial m[511] = 0;
initial m[512] = 0;
initial m[513] = 0;
initial m[514] = 1;
initial m[515] = 1;
initial m[516] = 0;
initial m[517] = 0;
initial m[518] = 1;
initial m[519] = 0;
initial m[520] = 0;
initial m[521] = 1;
initial m[522] = 0;
initial m[523] = 1;
initial m[524] = 0;
initial m[525] = 0;
initial m[526] = 1;
initial m[527] = 1;
initial m[528] = 0;
initial m[529] = 0;
initial m[532] = 0;
initial m[533] = 0;
initial m[534] = 1;
initial m[535] = 1;
initial m[536] = 0;
initial m[537] = 0;
initial m[538] = 1;
initial m[539] = 0;
initial m[542] = 0;
initial m[543] = 0;
initial m[544] = 0;
initial m[545] = 0;
initial m[546] = 1;
initial m[547] = 1;
initial m[548] = 1;
initial m[549] = 1;
initial m[550] = 1;
initial m[551] = 1;
initial m[552] = 0;
initial m[553] = 0;
initial m[554] = 1;
initial m[557] = 1;
initial m[558] = 0;
initial m[559] = 0;
initial m[560] = 0;
initial m[561] = 1;
initial m[562] = 1;
initial m[563] = 1;
initial m[564] = 0;
initial m[565] = 1;
initial m[566] = 1;
initial m[567] = 0;
initial m[568] = 0;
initial m[569] = 0;
initial m[570] = 1;
initial m[571] = 0;
initial m[572] = 0;
initial m[573] = 1;
initial m[574] = 0;
initial m[577] = 1;
initial m[578] = 1;
initial m[579] = 1;
initial m[580] = 1;
initial m[581] = 1;
initial m[582] = 0;
initial m[583] = 0;
initial m[584] = 0;
initial m[585] = 0;
initial m[586] = 1;
initial m[587] = 0;
initial m[588] = 0;
initial m[589] = 0;
initial m[590] = 0;
initial m[591] = 1;
initial m[592] = 0;
initial m[593] = 1;
initial m[594] = 1;
initial m[595] = 0;
initial m[596] = 0;
initial m[597] = 0;
initial m[598] = 1;
initial m[599] = 1;
initial m[602] = 0;
initial m[603] = 0;
initial m[604] = 0;
initial m[605] = 1;
initial m[606] = 1;
initial m[607] = 0;
initial m[608] = 1;
initial m[609] = 0;
initial m[610] = 0;
initial m[611] = 1;
initial m[612] = 0;
initial m[613] = 0;
initial m[614] = 0;
initial m[615] = 1;
initial m[616] = 0;
initial m[617] = 1;
initial m[618] = 0;
initial m[619] = 1;
initial m[620] = 1;
initial m[621] = 1;
initial m[622] = 0;
initial m[623] = 0;
initial m[624] = 1;
initial m[625] = 0;
initial m[626] = 0;
initial m[627] = 0;
initial m[628] = 0;
initial m[629] = 1;
initial m[632] = 1;
initial m[633] = 1;
initial m[634] = 1;
initial m[635] = 0;
initial m[636] = 1;
initial m[637] = 1;
initial m[638] = 0;
initial m[639] = 1;
initial m[640] = 1;
initial m[641] = 0;
initial m[642] = 1;
initial m[643] = 1;
initial m[644] = 0;
initial m[645] = 1;
initial m[646] = 0;
initial m[647] = 0;
initial m[648] = 0;
initial m[649] = 0;
initial m[650] = 1;
initial m[651] = 0;
initial m[652] = 0;
initial m[653] = 1;
initial m[654] = 0;
initial m[655] = 1;
initial m[656] = 1;
initial m[657] = 1;
initial m[658] = 0;
initial m[659] = 1;
initial m[660] = 0;
initial m[661] = 1;
initial m[662] = 1;
initial m[663] = 1;
initial m[664] = 1;
initial m[667] = 1;
initial m[668] = 0;
initial m[669] = 0;
initial m[670] = 1;
initial m[671] = 0;
initial m[672] = 1;
initial m[673] = 0;
initial m[674] = 0;
initial m[675] = 1;
initial m[676] = 0;
initial m[677] = 0;
initial m[678] = 0;
initial m[679] = 0;
initial m[680] = 0;
initial m[681] = 1;
initial m[682] = 0;
initial m[683] = 0;
initial m[684] = 1;
initial m[685] = 1;
initial m[686] = 1;
initial m[687] = 1;
initial m[688] = 1;
initial m[689] = 1;
initial m[690] = 1;
initial m[691] = 1;
initial m[692] = 1;
initial m[693] = 1;
initial m[694] = 0;
initial m[695] = 1;
initial m[696] = 0;
initial m[697] = 1;
initial m[698] = 0;
initial m[699] = 1;
initial m[700] = 0;
initial m[701] = 1;
initial m[702] = 0;
initial m[703] = 1;
initial m[704] = 1;
initial m[707] = 0;
initial m[708] = 0;
initial m[709] = 0;
initial m[710] = 0;
initial m[711] = 0;
initial m[712] = 0;
initial m[713] = 1;
initial m[714] = 1;
initial m[715] = 0;
initial m[716] = 1;
initial m[717] = 0;
initial m[718] = 1;
initial m[719] = 0;
initial m[720] = 0;
initial m[721] = 1;
initial m[722] = 0;
initial m[723] = 1;
initial m[724] = 0;
initial m[725] = 1;
initial m[726] = 1;
initial m[727] = 1;
initial m[728] = 0;
initial m[729] = 0;
initial m[730] = 1;
initial m[731] = 0;
initial m[732] = 0;
initial m[733] = 0;
initial m[734] = 0;
initial m[735] = 0;
initial m[736] = 0;
initial m[737] = 1;
initial m[738] = 1;
initial m[739] = 1;
initial m[740] = 0;
initial m[741] = 1;
initial m[742] = 1;
initial m[743] = 1;
initial m[744] = 1;
initial m[745] = 0;
initial m[746] = 0;
initial m[747] = 0;
initial m[748] = 0;
initial m[749] = 0;
initial m[752] = 0;
initial m[753] = 0;
initial m[754] = 0;
initial m[755] = 0;
initial m[756] = 0;
initial m[757] = 0;
initial m[758] = 1;
initial m[759] = 1;
initial m[760] = 0;
initial m[761] = 1;
initial m[762] = 0;
initial m[763] = 1;
initial m[764] = 1;
initial m[765] = 1;
initial m[766] = 1;
initial m[767] = 0;
initial m[768] = 0;
initial m[769] = 0;
initial m[770] = 1;
initial m[771] = 1;
initial m[772] = 0;
initial m[773] = 1;
initial m[774] = 0;
initial m[775] = 0;
initial m[776] = 1;
initial m[777] = 1;
initial m[778] = 0;
initial m[779] = 1;
initial m[780] = 0;
initial m[781] = 0;
initial m[782] = 1;
initial m[783] = 1;
initial m[784] = 1;
initial m[785] = 1;
initial m[786] = 1;
initial m[787] = 1;
initial m[788] = 1;
initial m[789] = 0;
initial m[790] = 1;
initial m[791] = 1;
initial m[792] = 1;
initial m[793] = 0;
initial m[794] = 1;
initial m[795] = 0;
initial m[796] = 0;
initial m[797] = 1;
initial m[798] = 0;
initial m[799] = 1;
initial m[802] = 0;
initial m[803] = 1;
initial m[804] = 0;
initial m[805] = 1;
initial m[806] = 0;
initial m[807] = 1;
initial m[808] = 1;
initial m[809] = 1;
initial m[810] = 0;
initial m[811] = 1;
initial m[812] = 0;
initial m[813] = 0;
initial m[814] = 1;
initial m[815] = 1;
initial m[816] = 0;
initial m[817] = 1;
initial m[818] = 0;
initial m[819] = 1;
initial m[820] = 0;
initial m[821] = 1;
initial m[822] = 0;
initial m[823] = 0;
initial m[824] = 0;
initial m[825] = 1;
initial m[826] = 1;
initial m[827] = 1;
initial m[828] = 0;
initial m[829] = 1;
initial m[830] = 0;
initial m[831] = 0;
initial m[832] = 0;
initial m[833] = 1;
initial m[834] = 0;
initial m[835] = 0;
initial m[836] = 0;
initial m[837] = 0;
initial m[838] = 1;
initial m[839] = 0;
initial m[840] = 0;
initial m[841] = 1;
initial m[842] = 1;
initial m[843] = 1;
initial m[844] = 1;
initial m[845] = 0;
initial m[846] = 1;
initial m[847] = 1;
initial m[848] = 1;
initial m[849] = 0;
initial m[850] = 0;
initial m[851] = 0;
initial m[852] = 1;
initial m[853] = 1;
initial m[854] = 0;
initial m[857] = 0;
initial m[859] = 1;
initial m[860] = 0;
initial m[861] = 1;
initial m[862] = 1;
initial m[863] = 1;
initial m[864] = 1;
initial m[865] = 1;
initial m[866] = 1;
initial m[867] = 0;
initial m[868] = 1;
initial m[869] = 0;
initial m[870] = 1;
initial m[871] = 0;
initial m[872] = 1;
initial m[873] = 0;
initial m[874] = 1;
initial m[875] = 1;
initial m[876] = 1;
initial m[877] = 1;
initial m[878] = 1;
initial m[879] = 1;
initial m[880] = 1;
initial m[881] = 0;
initial m[882] = 0;
initial m[883] = 1;
initial m[884] = 0;
initial m[885] = 1;
initial m[886] = 1;
initial m[887] = 1;
initial m[888] = 1;
initial m[889] = 0;
initial m[890] = 0;
initial m[891] = 0;
initial m[892] = 0;
initial m[893] = 0;
initial m[894] = 0;
initial m[895] = 0;
initial m[896] = 1;
initial m[897] = 1;
initial m[898] = 1;
initial m[899] = 1;
initial m[900] = 1;
initial m[901] = 0;
initial m[902] = 1;
initial m[903] = 1;
initial m[904] = 0;
initial m[905] = 0;
initial m[906] = 1;
initial m[907] = 1;
initial m[908] = 1;
initial m[909] = 0;
initial m[910] = 1;
initial m[912] = 1;
initial m[913] = 1;
initial m[914] = 1;
initial m[915] = 1;
initial m[916] = 0;
initial m[917] = 0;
initial m[918] = 0;
initial m[919] = 0;
initial m[920] = 0;
initial m[921] = 0;
initial m[922] = 0;
initial m[923] = 1;
initial m[924] = 0;
initial m[925] = 1;
initial m[926] = 1;
initial m[927] = 1;
initial m[928] = 0;
initial m[929] = 0;
initial m[930] = 0;
initial m[931] = 1;
initial m[932] = 1;
initial m[933] = 0;
initial m[934] = 1;
initial m[935] = 0;
initial m[936] = 0;
initial m[937] = 1;
initial m[938] = 0;
initial m[939] = 1;
initial m[940] = 0;
initial m[941] = 0;
initial m[942] = 1;
initial m[943] = 0;
initial m[944] = 1;
initial m[945] = 1;
initial m[946] = 1;
initial m[947] = 1;
initial m[948] = 0;
initial m[949] = 1;
initial m[950] = 0;
initial m[951] = 1;
initial m[952] = 0;
initial m[953] = 1;
initial m[954] = 1;
initial m[955] = 0;
initial m[956] = 1;
initial m[957] = 1;
initial m[958] = 0;
initial m[959] = 1;
initial m[960] = 0;
initial m[962] = 1;
initial m[963] = 0;
initial m[964] = 1;
initial m[965] = 0;
initial m[966] = 1;
initial m[967] = 1;
initial m[968] = 0;
initial m[969] = 0;
initial m[970] = 1;
initial m[971] = 1;
initial m[972] = 1;
initial m[973] = 0;
initial m[974] = 1;
initial m[975] = 1;
initial m[976] = 0;
initial m[977] = 1;
initial m[978] = 1;
initial m[979] = 0;
initial m[980] = 1;
initial m[981] = 0;
initial m[982] = 0;
initial m[983] = 1;
initial m[984] = 0;
initial m[985] = 0;
initial m[986] = 1;
initial m[987] = 1;
initial m[988] = 0;
initial m[989] = 1;
initial m[990] = 1;
initial m[991] = 0;
initial m[992] = 0;
initial m[993] = 0;
initial m[994] = 1;
initial m[995] = 1;
initial m[996] = 1;
initial m[997] = 1;
initial m[998] = 1;
initial m[999] = 1;
initial m[1000] = 1;
initial m[1001] = 1;
initial m[1002] = 1;
initial m[1003] = 0;
initial m[1004] = 0;
initial m[1005] = 0;
initial m[1007] = 0;
initial m[1008] = 0;
initial m[1009] = 0;
initial m[1010] = 0;
initial m[1011] = 0;
initial m[1012] = 0;
initial m[1013] = 0;
initial m[1014] = 0;
initial m[1015] = 0;
initial m[1016] = 1;
initial m[1017] = 1;
initial m[1018] = 1;
initial m[1019] = 0;
initial m[1020] = 1;
initial m[1021] = 0;
initial m[1022] = 0;
initial m[1023] = 1;
initial m[1024] = 0;
initial m[1025] = 0;
initial m[1026] = 0;
initial m[1027] = 1;
initial m[1028] = 0;
initial m[1029] = 1;
initial m[1030] = 1;
initial m[1031] = 1;
initial m[1032] = 0;
initial m[1033] = 1;
initial m[1034] = 1;
initial m[1035] = 1;
initial m[1036] = 0;
initial m[1037] = 1;
initial m[1038] = 1;
initial m[1039] = 0;
initial m[1040] = 1;
initial m[1041] = 1;
initial m[1042] = 1;
initial m[1043] = 1;
initial m[1044] = 1;
initial m[1045] = 1;
initial m[1047] = 1;
initial m[1048] = 1;
initial m[1049] = 1;
initial m[1050] = 0;
initial m[1051] = 0;
initial m[1052] = 0;
initial m[1053] = 0;
initial m[1054] = 0;
initial m[1055] = 0;
initial m[1056] = 0;
initial m[1057] = 0;
initial m[1058] = 1;
initial m[1059] = 0;
initial m[1060] = 1;
initial m[1061] = 0;
initial m[1062] = 1;
initial m[1063] = 0;
initial m[1064] = 0;
initial m[1065] = 1;
initial m[1066] = 0;
initial m[1067] = 1;
initial m[1068] = 1;
initial m[1069] = 0;
initial m[1070] = 0;
initial m[1071] = 1;
initial m[1072] = 1;
initial m[1073] = 1;
initial m[1074] = 0;
initial m[1075] = 0;
initial m[1076] = 0;
initial m[1077] = 0;
initial m[1078] = 0;
initial m[1079] = 0;
initial m[1080] = 0;
initial m[1082] = 1;
initial m[1083] = 0;
initial m[1084] = 1;
initial m[1085] = 1;
initial m[1086] = 1;
initial m[1087] = 0;
initial m[1088] = 0;
initial m[1089] = 1;
initial m[1090] = 0;
initial m[1091] = 1;
initial m[1092] = 1;
initial m[1093] = 1;
initial m[1094] = 0;
initial m[1095] = 0;
initial m[1096] = 0;
initial m[1097] = 1;
initial m[1098] = 1;
initial m[1099] = 0;
initial m[1100] = 0;
initial m[1101] = 1;
initial m[1102] = 0;
initial m[1103] = 0;
initial m[1104] = 0;
initial m[1105] = 0;
initial m[1106] = 0;
initial m[1107] = 0;
initial m[1108] = 0;
initial m[1109] = 1;
initial m[1110] = 1;
initial m[1112] = 0;
initial m[1113] = 1;
initial m[1114] = 0;
initial m[1115] = 0;
initial m[1116] = 0;
initial m[1117] = 1;
initial m[1118] = 1;
initial m[1119] = 0;
initial m[1120] = 1;
initial m[1121] = 1;
initial m[1122] = 0;
initial m[1123] = 0;
initial m[1124] = 1;
initial m[1125] = 1;
initial m[1126] = 0;
initial m[1127] = 1;
initial m[1128] = 0;
initial m[1129] = 0;
initial m[1130] = 0;
initial m[1131] = 0;
initial m[1132] = 0;
initial m[1133] = 0;
initial m[1134] = 1;
initial m[1135] = 1;
initial m[1137] = 0;
initial m[1138] = 1;
initial m[1139] = 1;
initial m[1140] = 0;
initial m[1141] = 1;
initial m[1142] = 0;
initial m[1143] = 1;
initial m[1144] = 1;
initial m[1145] = 0;
initial m[1146] = 0;
initial m[1147] = 0;
initial m[1148] = 1;
initial m[1149] = 1;
initial m[1150] = 0;
initial m[1151] = 1;
initial m[1152] = 1;
initial m[1153] = 1;
initial m[1154] = 1;
initial m[1155] = 0;
initial m[1157] = 0;
initial m[1158] = 1;
initial m[1159] = 0;
initial m[1160] = 1;
initial m[1161] = 0;
initial m[1162] = 0;
initial m[1163] = 1;
initial m[1164] = 1;
initial m[1165] = 0;
initial m[1166] = 0;
initial m[1167] = 0;
initial m[1168] = 1;
initial m[1169] = 1;
initial m[1170] = 0;
initial m[1172] = 1;
initial m[1173] = 0;
initial m[1174] = 1;
initial m[1175] = 0;
initial m[1176] = 0;
initial m[1177] = 1;
initial m[1178] = 1;
initial m[1179] = 1;
initial m[1180] = 0;
initial m[1182] = 0;
initial m[1183] = 1;
initial m[1184] = 1;
initial m[1185] = 1;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[11],m[10],m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[23],m[22],m[21],m[20],m[19],m[18],m[17],m[16],m[15],m[14],m[13],m[12]};
end

always @(negedge sample_clk) begin
    if (solution == 24'b111111000010001011111101)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[24]&~m[25]&~m[26])|(~m[24]&m[25]&~m[26])|(~m[24]&~m[25]&m[26]))&BiasedRNG[0])|(((m[24]&m[25]&~m[26])|(m[24]&~m[25]&m[26])|(~m[24]&m[25]&m[26]))&~BiasedRNG[0])|((m[24]&m[25]&m[26]));
    m[1] = (((m[27]&~m[28]&~m[29])|(~m[27]&m[28]&~m[29])|(~m[27]&~m[28]&m[29]))&BiasedRNG[1])|(((m[27]&m[28]&~m[29])|(m[27]&~m[28]&m[29])|(~m[27]&m[28]&m[29]))&~BiasedRNG[1])|((m[27]&m[28]&m[29]));
    m[2] = (((m[30]&~m[31]&~m[32])|(~m[30]&m[31]&~m[32])|(~m[30]&~m[31]&m[32]))&BiasedRNG[2])|(((m[30]&m[31]&~m[32])|(m[30]&~m[31]&m[32])|(~m[30]&m[31]&m[32]))&~BiasedRNG[2])|((m[30]&m[31]&m[32]));
    m[3] = (((m[33]&~m[34]&~m[35])|(~m[33]&m[34]&~m[35])|(~m[33]&~m[34]&m[35]))&BiasedRNG[3])|(((m[33]&m[34]&~m[35])|(m[33]&~m[34]&m[35])|(~m[33]&m[34]&m[35]))&~BiasedRNG[3])|((m[33]&m[34]&m[35]));
    m[4] = (((m[36]&~m[37]&~m[38])|(~m[36]&m[37]&~m[38])|(~m[36]&~m[37]&m[38]))&BiasedRNG[4])|(((m[36]&m[37]&~m[38])|(m[36]&~m[37]&m[38])|(~m[36]&m[37]&m[38]))&~BiasedRNG[4])|((m[36]&m[37]&m[38]));
    m[5] = (((m[39]&~m[40]&~m[41])|(~m[39]&m[40]&~m[41])|(~m[39]&~m[40]&m[41]))&BiasedRNG[5])|(((m[39]&m[40]&~m[41])|(m[39]&~m[40]&m[41])|(~m[39]&m[40]&m[41]))&~BiasedRNG[5])|((m[39]&m[40]&m[41]));
    m[6] = (((m[42]&~m[43]&~m[44])|(~m[42]&m[43]&~m[44])|(~m[42]&~m[43]&m[44]))&BiasedRNG[6])|(((m[42]&m[43]&~m[44])|(m[42]&~m[43]&m[44])|(~m[42]&m[43]&m[44]))&~BiasedRNG[6])|((m[42]&m[43]&m[44]));
    m[7] = (((m[45]&~m[46]&~m[47])|(~m[45]&m[46]&~m[47])|(~m[45]&~m[46]&m[47]))&BiasedRNG[7])|(((m[45]&m[46]&~m[47])|(m[45]&~m[46]&m[47])|(~m[45]&m[46]&m[47]))&~BiasedRNG[7])|((m[45]&m[46]&m[47]));
    m[8] = (((m[48]&~m[49]&~m[50])|(~m[48]&m[49]&~m[50])|(~m[48]&~m[49]&m[50]))&BiasedRNG[8])|(((m[48]&m[49]&~m[50])|(m[48]&~m[49]&m[50])|(~m[48]&m[49]&m[50]))&~BiasedRNG[8])|((m[48]&m[49]&m[50]));
    m[9] = (((m[51]&~m[52]&~m[53])|(~m[51]&m[52]&~m[53])|(~m[51]&~m[52]&m[53]))&BiasedRNG[9])|(((m[51]&m[52]&~m[53])|(m[51]&~m[52]&m[53])|(~m[51]&m[52]&m[53]))&~BiasedRNG[9])|((m[51]&m[52]&m[53]));
    m[10] = (((m[54]&~m[55]&~m[56])|(~m[54]&m[55]&~m[56])|(~m[54]&~m[55]&m[56]))&BiasedRNG[10])|(((m[54]&m[55]&~m[56])|(m[54]&~m[55]&m[56])|(~m[54]&m[55]&m[56]))&~BiasedRNG[10])|((m[54]&m[55]&m[56]));
    m[11] = (((m[57]&~m[58]&~m[59])|(~m[57]&m[58]&~m[59])|(~m[57]&~m[58]&m[59]))&BiasedRNG[11])|(((m[57]&m[58]&~m[59])|(m[57]&~m[58]&m[59])|(~m[57]&m[58]&m[59]))&~BiasedRNG[11])|((m[57]&m[58]&m[59]));
    m[12] = (((m[60]&~m[61]&~m[62])|(~m[60]&m[61]&~m[62])|(~m[60]&~m[61]&m[62]))&BiasedRNG[12])|(((m[60]&m[61]&~m[62])|(m[60]&~m[61]&m[62])|(~m[60]&m[61]&m[62]))&~BiasedRNG[12])|((m[60]&m[61]&m[62]));
    m[13] = (((m[63]&~m[64]&~m[65])|(~m[63]&m[64]&~m[65])|(~m[63]&~m[64]&m[65]))&BiasedRNG[13])|(((m[63]&m[64]&~m[65])|(m[63]&~m[64]&m[65])|(~m[63]&m[64]&m[65]))&~BiasedRNG[13])|((m[63]&m[64]&m[65]));
    m[14] = (((m[66]&~m[67]&~m[68])|(~m[66]&m[67]&~m[68])|(~m[66]&~m[67]&m[68]))&BiasedRNG[14])|(((m[66]&m[67]&~m[68])|(m[66]&~m[67]&m[68])|(~m[66]&m[67]&m[68]))&~BiasedRNG[14])|((m[66]&m[67]&m[68]));
    m[15] = (((m[69]&~m[70]&~m[71])|(~m[69]&m[70]&~m[71])|(~m[69]&~m[70]&m[71]))&BiasedRNG[15])|(((m[69]&m[70]&~m[71])|(m[69]&~m[70]&m[71])|(~m[69]&m[70]&m[71]))&~BiasedRNG[15])|((m[69]&m[70]&m[71]));
    m[16] = (((m[72]&~m[73]&~m[74])|(~m[72]&m[73]&~m[74])|(~m[72]&~m[73]&m[74]))&BiasedRNG[16])|(((m[72]&m[73]&~m[74])|(m[72]&~m[73]&m[74])|(~m[72]&m[73]&m[74]))&~BiasedRNG[16])|((m[72]&m[73]&m[74]));
    m[17] = (((m[75]&~m[76]&~m[77])|(~m[75]&m[76]&~m[77])|(~m[75]&~m[76]&m[77]))&BiasedRNG[17])|(((m[75]&m[76]&~m[77])|(m[75]&~m[76]&m[77])|(~m[75]&m[76]&m[77]))&~BiasedRNG[17])|((m[75]&m[76]&m[77]));
    m[18] = (((m[78]&~m[79]&~m[80])|(~m[78]&m[79]&~m[80])|(~m[78]&~m[79]&m[80]))&BiasedRNG[18])|(((m[78]&m[79]&~m[80])|(m[78]&~m[79]&m[80])|(~m[78]&m[79]&m[80]))&~BiasedRNG[18])|((m[78]&m[79]&m[80]));
    m[19] = (((m[81]&~m[82]&~m[83])|(~m[81]&m[82]&~m[83])|(~m[81]&~m[82]&m[83]))&BiasedRNG[19])|(((m[81]&m[82]&~m[83])|(m[81]&~m[82]&m[83])|(~m[81]&m[82]&m[83]))&~BiasedRNG[19])|((m[81]&m[82]&m[83]));
    m[20] = (((m[84]&~m[85]&~m[86])|(~m[84]&m[85]&~m[86])|(~m[84]&~m[85]&m[86]))&BiasedRNG[20])|(((m[84]&m[85]&~m[86])|(m[84]&~m[85]&m[86])|(~m[84]&m[85]&m[86]))&~BiasedRNG[20])|((m[84]&m[85]&m[86]));
    m[21] = (((m[87]&~m[88]&~m[89])|(~m[87]&m[88]&~m[89])|(~m[87]&~m[88]&m[89]))&BiasedRNG[21])|(((m[87]&m[88]&~m[89])|(m[87]&~m[88]&m[89])|(~m[87]&m[88]&m[89]))&~BiasedRNG[21])|((m[87]&m[88]&m[89]));
    m[22] = (((m[90]&~m[91]&~m[92])|(~m[90]&m[91]&~m[92])|(~m[90]&~m[91]&m[92]))&BiasedRNG[22])|(((m[90]&m[91]&~m[92])|(m[90]&~m[91]&m[92])|(~m[90]&m[91]&m[92]))&~BiasedRNG[22])|((m[90]&m[91]&m[92]));
    m[23] = (((m[93]&~m[94]&~m[95])|(~m[93]&m[94]&~m[95])|(~m[93]&~m[94]&m[95]))&BiasedRNG[23])|(((m[93]&m[94]&~m[95])|(m[93]&~m[94]&m[95])|(~m[93]&m[94]&m[95]))&~BiasedRNG[23])|((m[93]&m[94]&m[95]));
    m[96] = (((~m[24]&~m[240]&~m[384])|(m[24]&m[240]&~m[384]))&BiasedRNG[24])|(((m[24]&~m[240]&~m[384])|(~m[24]&m[240]&m[384]))&~BiasedRNG[24])|((~m[24]&~m[240]&m[384])|(m[24]&~m[240]&m[384])|(m[24]&m[240]&m[384]));
    m[97] = (((~m[24]&~m[252]&~m[396])|(m[24]&m[252]&~m[396]))&BiasedRNG[25])|(((m[24]&~m[252]&~m[396])|(~m[24]&m[252]&m[396]))&~BiasedRNG[25])|((~m[24]&~m[252]&m[396])|(m[24]&~m[252]&m[396])|(m[24]&m[252]&m[396]));
    m[98] = (((~m[24]&~m[264]&~m[408])|(m[24]&m[264]&~m[408]))&BiasedRNG[26])|(((m[24]&~m[264]&~m[408])|(~m[24]&m[264]&m[408]))&~BiasedRNG[26])|((~m[24]&~m[264]&m[408])|(m[24]&~m[264]&m[408])|(m[24]&m[264]&m[408]));
    m[99] = (((~m[24]&~m[276]&~m[420])|(m[24]&m[276]&~m[420]))&BiasedRNG[27])|(((m[24]&~m[276]&~m[420])|(~m[24]&m[276]&m[420]))&~BiasedRNG[27])|((~m[24]&~m[276]&m[420])|(m[24]&~m[276]&m[420])|(m[24]&m[276]&m[420]));
    m[100] = (((~m[25]&~m[288]&~m[432])|(m[25]&m[288]&~m[432]))&BiasedRNG[28])|(((m[25]&~m[288]&~m[432])|(~m[25]&m[288]&m[432]))&~BiasedRNG[28])|((~m[25]&~m[288]&m[432])|(m[25]&~m[288]&m[432])|(m[25]&m[288]&m[432]));
    m[101] = (((~m[25]&~m[300]&~m[444])|(m[25]&m[300]&~m[444]))&BiasedRNG[29])|(((m[25]&~m[300]&~m[444])|(~m[25]&m[300]&m[444]))&~BiasedRNG[29])|((~m[25]&~m[300]&m[444])|(m[25]&~m[300]&m[444])|(m[25]&m[300]&m[444]));
    m[102] = (((~m[25]&~m[312]&~m[456])|(m[25]&m[312]&~m[456]))&BiasedRNG[30])|(((m[25]&~m[312]&~m[456])|(~m[25]&m[312]&m[456]))&~BiasedRNG[30])|((~m[25]&~m[312]&m[456])|(m[25]&~m[312]&m[456])|(m[25]&m[312]&m[456]));
    m[103] = (((~m[25]&~m[324]&~m[468])|(m[25]&m[324]&~m[468]))&BiasedRNG[31])|(((m[25]&~m[324]&~m[468])|(~m[25]&m[324]&m[468]))&~BiasedRNG[31])|((~m[25]&~m[324]&m[468])|(m[25]&~m[324]&m[468])|(m[25]&m[324]&m[468]));
    m[104] = (((~m[26]&~m[336]&~m[480])|(m[26]&m[336]&~m[480]))&BiasedRNG[32])|(((m[26]&~m[336]&~m[480])|(~m[26]&m[336]&m[480]))&~BiasedRNG[32])|((~m[26]&~m[336]&m[480])|(m[26]&~m[336]&m[480])|(m[26]&m[336]&m[480]));
    m[105] = (((~m[26]&~m[348]&~m[492])|(m[26]&m[348]&~m[492]))&BiasedRNG[33])|(((m[26]&~m[348]&~m[492])|(~m[26]&m[348]&m[492]))&~BiasedRNG[33])|((~m[26]&~m[348]&m[492])|(m[26]&~m[348]&m[492])|(m[26]&m[348]&m[492]));
    m[106] = (((~m[26]&~m[360]&~m[504])|(m[26]&m[360]&~m[504]))&BiasedRNG[34])|(((m[26]&~m[360]&~m[504])|(~m[26]&m[360]&m[504]))&~BiasedRNG[34])|((~m[26]&~m[360]&m[504])|(m[26]&~m[360]&m[504])|(m[26]&m[360]&m[504]));
    m[107] = (((~m[26]&~m[372]&~m[516])|(m[26]&m[372]&~m[516]))&BiasedRNG[35])|(((m[26]&~m[372]&~m[516])|(~m[26]&m[372]&m[516]))&~BiasedRNG[35])|((~m[26]&~m[372]&m[516])|(m[26]&~m[372]&m[516])|(m[26]&m[372]&m[516]));
    m[108] = (((~m[27]&~m[241]&~m[385])|(m[27]&m[241]&~m[385]))&BiasedRNG[36])|(((m[27]&~m[241]&~m[385])|(~m[27]&m[241]&m[385]))&~BiasedRNG[36])|((~m[27]&~m[241]&m[385])|(m[27]&~m[241]&m[385])|(m[27]&m[241]&m[385]));
    m[109] = (((~m[27]&~m[253]&~m[397])|(m[27]&m[253]&~m[397]))&BiasedRNG[37])|(((m[27]&~m[253]&~m[397])|(~m[27]&m[253]&m[397]))&~BiasedRNG[37])|((~m[27]&~m[253]&m[397])|(m[27]&~m[253]&m[397])|(m[27]&m[253]&m[397]));
    m[110] = (((~m[27]&~m[265]&~m[409])|(m[27]&m[265]&~m[409]))&BiasedRNG[38])|(((m[27]&~m[265]&~m[409])|(~m[27]&m[265]&m[409]))&~BiasedRNG[38])|((~m[27]&~m[265]&m[409])|(m[27]&~m[265]&m[409])|(m[27]&m[265]&m[409]));
    m[111] = (((~m[27]&~m[277]&~m[421])|(m[27]&m[277]&~m[421]))&BiasedRNG[39])|(((m[27]&~m[277]&~m[421])|(~m[27]&m[277]&m[421]))&~BiasedRNG[39])|((~m[27]&~m[277]&m[421])|(m[27]&~m[277]&m[421])|(m[27]&m[277]&m[421]));
    m[112] = (((~m[28]&~m[289]&~m[433])|(m[28]&m[289]&~m[433]))&BiasedRNG[40])|(((m[28]&~m[289]&~m[433])|(~m[28]&m[289]&m[433]))&~BiasedRNG[40])|((~m[28]&~m[289]&m[433])|(m[28]&~m[289]&m[433])|(m[28]&m[289]&m[433]));
    m[113] = (((~m[28]&~m[301]&~m[445])|(m[28]&m[301]&~m[445]))&BiasedRNG[41])|(((m[28]&~m[301]&~m[445])|(~m[28]&m[301]&m[445]))&~BiasedRNG[41])|((~m[28]&~m[301]&m[445])|(m[28]&~m[301]&m[445])|(m[28]&m[301]&m[445]));
    m[114] = (((~m[28]&~m[313]&~m[457])|(m[28]&m[313]&~m[457]))&BiasedRNG[42])|(((m[28]&~m[313]&~m[457])|(~m[28]&m[313]&m[457]))&~BiasedRNG[42])|((~m[28]&~m[313]&m[457])|(m[28]&~m[313]&m[457])|(m[28]&m[313]&m[457]));
    m[115] = (((~m[28]&~m[325]&~m[469])|(m[28]&m[325]&~m[469]))&BiasedRNG[43])|(((m[28]&~m[325]&~m[469])|(~m[28]&m[325]&m[469]))&~BiasedRNG[43])|((~m[28]&~m[325]&m[469])|(m[28]&~m[325]&m[469])|(m[28]&m[325]&m[469]));
    m[116] = (((~m[29]&~m[337]&~m[481])|(m[29]&m[337]&~m[481]))&BiasedRNG[44])|(((m[29]&~m[337]&~m[481])|(~m[29]&m[337]&m[481]))&~BiasedRNG[44])|((~m[29]&~m[337]&m[481])|(m[29]&~m[337]&m[481])|(m[29]&m[337]&m[481]));
    m[117] = (((~m[29]&~m[349]&~m[493])|(m[29]&m[349]&~m[493]))&BiasedRNG[45])|(((m[29]&~m[349]&~m[493])|(~m[29]&m[349]&m[493]))&~BiasedRNG[45])|((~m[29]&~m[349]&m[493])|(m[29]&~m[349]&m[493])|(m[29]&m[349]&m[493]));
    m[118] = (((~m[29]&~m[361]&~m[505])|(m[29]&m[361]&~m[505]))&BiasedRNG[46])|(((m[29]&~m[361]&~m[505])|(~m[29]&m[361]&m[505]))&~BiasedRNG[46])|((~m[29]&~m[361]&m[505])|(m[29]&~m[361]&m[505])|(m[29]&m[361]&m[505]));
    m[119] = (((~m[29]&~m[373]&~m[517])|(m[29]&m[373]&~m[517]))&BiasedRNG[47])|(((m[29]&~m[373]&~m[517])|(~m[29]&m[373]&m[517]))&~BiasedRNG[47])|((~m[29]&~m[373]&m[517])|(m[29]&~m[373]&m[517])|(m[29]&m[373]&m[517]));
    m[120] = (((~m[30]&~m[242]&~m[386])|(m[30]&m[242]&~m[386]))&BiasedRNG[48])|(((m[30]&~m[242]&~m[386])|(~m[30]&m[242]&m[386]))&~BiasedRNG[48])|((~m[30]&~m[242]&m[386])|(m[30]&~m[242]&m[386])|(m[30]&m[242]&m[386]));
    m[121] = (((~m[30]&~m[254]&~m[398])|(m[30]&m[254]&~m[398]))&BiasedRNG[49])|(((m[30]&~m[254]&~m[398])|(~m[30]&m[254]&m[398]))&~BiasedRNG[49])|((~m[30]&~m[254]&m[398])|(m[30]&~m[254]&m[398])|(m[30]&m[254]&m[398]));
    m[122] = (((~m[30]&~m[266]&~m[410])|(m[30]&m[266]&~m[410]))&BiasedRNG[50])|(((m[30]&~m[266]&~m[410])|(~m[30]&m[266]&m[410]))&~BiasedRNG[50])|((~m[30]&~m[266]&m[410])|(m[30]&~m[266]&m[410])|(m[30]&m[266]&m[410]));
    m[123] = (((~m[30]&~m[278]&~m[422])|(m[30]&m[278]&~m[422]))&BiasedRNG[51])|(((m[30]&~m[278]&~m[422])|(~m[30]&m[278]&m[422]))&~BiasedRNG[51])|((~m[30]&~m[278]&m[422])|(m[30]&~m[278]&m[422])|(m[30]&m[278]&m[422]));
    m[124] = (((~m[31]&~m[290]&~m[434])|(m[31]&m[290]&~m[434]))&BiasedRNG[52])|(((m[31]&~m[290]&~m[434])|(~m[31]&m[290]&m[434]))&~BiasedRNG[52])|((~m[31]&~m[290]&m[434])|(m[31]&~m[290]&m[434])|(m[31]&m[290]&m[434]));
    m[125] = (((~m[31]&~m[302]&~m[446])|(m[31]&m[302]&~m[446]))&BiasedRNG[53])|(((m[31]&~m[302]&~m[446])|(~m[31]&m[302]&m[446]))&~BiasedRNG[53])|((~m[31]&~m[302]&m[446])|(m[31]&~m[302]&m[446])|(m[31]&m[302]&m[446]));
    m[126] = (((~m[31]&~m[314]&~m[458])|(m[31]&m[314]&~m[458]))&BiasedRNG[54])|(((m[31]&~m[314]&~m[458])|(~m[31]&m[314]&m[458]))&~BiasedRNG[54])|((~m[31]&~m[314]&m[458])|(m[31]&~m[314]&m[458])|(m[31]&m[314]&m[458]));
    m[127] = (((~m[31]&~m[326]&~m[470])|(m[31]&m[326]&~m[470]))&BiasedRNG[55])|(((m[31]&~m[326]&~m[470])|(~m[31]&m[326]&m[470]))&~BiasedRNG[55])|((~m[31]&~m[326]&m[470])|(m[31]&~m[326]&m[470])|(m[31]&m[326]&m[470]));
    m[128] = (((~m[32]&~m[338]&~m[482])|(m[32]&m[338]&~m[482]))&BiasedRNG[56])|(((m[32]&~m[338]&~m[482])|(~m[32]&m[338]&m[482]))&~BiasedRNG[56])|((~m[32]&~m[338]&m[482])|(m[32]&~m[338]&m[482])|(m[32]&m[338]&m[482]));
    m[129] = (((~m[32]&~m[350]&~m[494])|(m[32]&m[350]&~m[494]))&BiasedRNG[57])|(((m[32]&~m[350]&~m[494])|(~m[32]&m[350]&m[494]))&~BiasedRNG[57])|((~m[32]&~m[350]&m[494])|(m[32]&~m[350]&m[494])|(m[32]&m[350]&m[494]));
    m[130] = (((~m[32]&~m[362]&~m[506])|(m[32]&m[362]&~m[506]))&BiasedRNG[58])|(((m[32]&~m[362]&~m[506])|(~m[32]&m[362]&m[506]))&~BiasedRNG[58])|((~m[32]&~m[362]&m[506])|(m[32]&~m[362]&m[506])|(m[32]&m[362]&m[506]));
    m[131] = (((~m[32]&~m[374]&~m[518])|(m[32]&m[374]&~m[518]))&BiasedRNG[59])|(((m[32]&~m[374]&~m[518])|(~m[32]&m[374]&m[518]))&~BiasedRNG[59])|((~m[32]&~m[374]&m[518])|(m[32]&~m[374]&m[518])|(m[32]&m[374]&m[518]));
    m[132] = (((~m[33]&~m[243]&~m[387])|(m[33]&m[243]&~m[387]))&BiasedRNG[60])|(((m[33]&~m[243]&~m[387])|(~m[33]&m[243]&m[387]))&~BiasedRNG[60])|((~m[33]&~m[243]&m[387])|(m[33]&~m[243]&m[387])|(m[33]&m[243]&m[387]));
    m[133] = (((~m[33]&~m[255]&~m[399])|(m[33]&m[255]&~m[399]))&BiasedRNG[61])|(((m[33]&~m[255]&~m[399])|(~m[33]&m[255]&m[399]))&~BiasedRNG[61])|((~m[33]&~m[255]&m[399])|(m[33]&~m[255]&m[399])|(m[33]&m[255]&m[399]));
    m[134] = (((~m[33]&~m[267]&~m[411])|(m[33]&m[267]&~m[411]))&BiasedRNG[62])|(((m[33]&~m[267]&~m[411])|(~m[33]&m[267]&m[411]))&~BiasedRNG[62])|((~m[33]&~m[267]&m[411])|(m[33]&~m[267]&m[411])|(m[33]&m[267]&m[411]));
    m[135] = (((~m[33]&~m[279]&~m[423])|(m[33]&m[279]&~m[423]))&BiasedRNG[63])|(((m[33]&~m[279]&~m[423])|(~m[33]&m[279]&m[423]))&~BiasedRNG[63])|((~m[33]&~m[279]&m[423])|(m[33]&~m[279]&m[423])|(m[33]&m[279]&m[423]));
    m[136] = (((~m[34]&~m[291]&~m[435])|(m[34]&m[291]&~m[435]))&BiasedRNG[64])|(((m[34]&~m[291]&~m[435])|(~m[34]&m[291]&m[435]))&~BiasedRNG[64])|((~m[34]&~m[291]&m[435])|(m[34]&~m[291]&m[435])|(m[34]&m[291]&m[435]));
    m[137] = (((~m[34]&~m[303]&~m[447])|(m[34]&m[303]&~m[447]))&BiasedRNG[65])|(((m[34]&~m[303]&~m[447])|(~m[34]&m[303]&m[447]))&~BiasedRNG[65])|((~m[34]&~m[303]&m[447])|(m[34]&~m[303]&m[447])|(m[34]&m[303]&m[447]));
    m[138] = (((~m[34]&~m[315]&~m[459])|(m[34]&m[315]&~m[459]))&BiasedRNG[66])|(((m[34]&~m[315]&~m[459])|(~m[34]&m[315]&m[459]))&~BiasedRNG[66])|((~m[34]&~m[315]&m[459])|(m[34]&~m[315]&m[459])|(m[34]&m[315]&m[459]));
    m[139] = (((~m[34]&~m[327]&~m[471])|(m[34]&m[327]&~m[471]))&BiasedRNG[67])|(((m[34]&~m[327]&~m[471])|(~m[34]&m[327]&m[471]))&~BiasedRNG[67])|((~m[34]&~m[327]&m[471])|(m[34]&~m[327]&m[471])|(m[34]&m[327]&m[471]));
    m[140] = (((~m[35]&~m[339]&~m[483])|(m[35]&m[339]&~m[483]))&BiasedRNG[68])|(((m[35]&~m[339]&~m[483])|(~m[35]&m[339]&m[483]))&~BiasedRNG[68])|((~m[35]&~m[339]&m[483])|(m[35]&~m[339]&m[483])|(m[35]&m[339]&m[483]));
    m[141] = (((~m[35]&~m[351]&~m[495])|(m[35]&m[351]&~m[495]))&BiasedRNG[69])|(((m[35]&~m[351]&~m[495])|(~m[35]&m[351]&m[495]))&~BiasedRNG[69])|((~m[35]&~m[351]&m[495])|(m[35]&~m[351]&m[495])|(m[35]&m[351]&m[495]));
    m[142] = (((~m[35]&~m[363]&~m[507])|(m[35]&m[363]&~m[507]))&BiasedRNG[70])|(((m[35]&~m[363]&~m[507])|(~m[35]&m[363]&m[507]))&~BiasedRNG[70])|((~m[35]&~m[363]&m[507])|(m[35]&~m[363]&m[507])|(m[35]&m[363]&m[507]));
    m[143] = (((~m[35]&~m[375]&~m[519])|(m[35]&m[375]&~m[519]))&BiasedRNG[71])|(((m[35]&~m[375]&~m[519])|(~m[35]&m[375]&m[519]))&~BiasedRNG[71])|((~m[35]&~m[375]&m[519])|(m[35]&~m[375]&m[519])|(m[35]&m[375]&m[519]));
    m[144] = (((~m[36]&~m[244]&~m[388])|(m[36]&m[244]&~m[388]))&BiasedRNG[72])|(((m[36]&~m[244]&~m[388])|(~m[36]&m[244]&m[388]))&~BiasedRNG[72])|((~m[36]&~m[244]&m[388])|(m[36]&~m[244]&m[388])|(m[36]&m[244]&m[388]));
    m[145] = (((~m[36]&~m[256]&~m[400])|(m[36]&m[256]&~m[400]))&BiasedRNG[73])|(((m[36]&~m[256]&~m[400])|(~m[36]&m[256]&m[400]))&~BiasedRNG[73])|((~m[36]&~m[256]&m[400])|(m[36]&~m[256]&m[400])|(m[36]&m[256]&m[400]));
    m[146] = (((~m[36]&~m[268]&~m[412])|(m[36]&m[268]&~m[412]))&BiasedRNG[74])|(((m[36]&~m[268]&~m[412])|(~m[36]&m[268]&m[412]))&~BiasedRNG[74])|((~m[36]&~m[268]&m[412])|(m[36]&~m[268]&m[412])|(m[36]&m[268]&m[412]));
    m[147] = (((~m[36]&~m[280]&~m[424])|(m[36]&m[280]&~m[424]))&BiasedRNG[75])|(((m[36]&~m[280]&~m[424])|(~m[36]&m[280]&m[424]))&~BiasedRNG[75])|((~m[36]&~m[280]&m[424])|(m[36]&~m[280]&m[424])|(m[36]&m[280]&m[424]));
    m[148] = (((~m[37]&~m[292]&~m[436])|(m[37]&m[292]&~m[436]))&BiasedRNG[76])|(((m[37]&~m[292]&~m[436])|(~m[37]&m[292]&m[436]))&~BiasedRNG[76])|((~m[37]&~m[292]&m[436])|(m[37]&~m[292]&m[436])|(m[37]&m[292]&m[436]));
    m[149] = (((~m[37]&~m[304]&~m[448])|(m[37]&m[304]&~m[448]))&BiasedRNG[77])|(((m[37]&~m[304]&~m[448])|(~m[37]&m[304]&m[448]))&~BiasedRNG[77])|((~m[37]&~m[304]&m[448])|(m[37]&~m[304]&m[448])|(m[37]&m[304]&m[448]));
    m[150] = (((~m[37]&~m[316]&~m[460])|(m[37]&m[316]&~m[460]))&BiasedRNG[78])|(((m[37]&~m[316]&~m[460])|(~m[37]&m[316]&m[460]))&~BiasedRNG[78])|((~m[37]&~m[316]&m[460])|(m[37]&~m[316]&m[460])|(m[37]&m[316]&m[460]));
    m[151] = (((~m[37]&~m[328]&~m[472])|(m[37]&m[328]&~m[472]))&BiasedRNG[79])|(((m[37]&~m[328]&~m[472])|(~m[37]&m[328]&m[472]))&~BiasedRNG[79])|((~m[37]&~m[328]&m[472])|(m[37]&~m[328]&m[472])|(m[37]&m[328]&m[472]));
    m[152] = (((~m[38]&~m[340]&~m[484])|(m[38]&m[340]&~m[484]))&BiasedRNG[80])|(((m[38]&~m[340]&~m[484])|(~m[38]&m[340]&m[484]))&~BiasedRNG[80])|((~m[38]&~m[340]&m[484])|(m[38]&~m[340]&m[484])|(m[38]&m[340]&m[484]));
    m[153] = (((~m[38]&~m[352]&~m[496])|(m[38]&m[352]&~m[496]))&BiasedRNG[81])|(((m[38]&~m[352]&~m[496])|(~m[38]&m[352]&m[496]))&~BiasedRNG[81])|((~m[38]&~m[352]&m[496])|(m[38]&~m[352]&m[496])|(m[38]&m[352]&m[496]));
    m[154] = (((~m[38]&~m[364]&~m[508])|(m[38]&m[364]&~m[508]))&BiasedRNG[82])|(((m[38]&~m[364]&~m[508])|(~m[38]&m[364]&m[508]))&~BiasedRNG[82])|((~m[38]&~m[364]&m[508])|(m[38]&~m[364]&m[508])|(m[38]&m[364]&m[508]));
    m[155] = (((~m[38]&~m[376]&~m[520])|(m[38]&m[376]&~m[520]))&BiasedRNG[83])|(((m[38]&~m[376]&~m[520])|(~m[38]&m[376]&m[520]))&~BiasedRNG[83])|((~m[38]&~m[376]&m[520])|(m[38]&~m[376]&m[520])|(m[38]&m[376]&m[520]));
    m[156] = (((~m[39]&~m[245]&~m[389])|(m[39]&m[245]&~m[389]))&BiasedRNG[84])|(((m[39]&~m[245]&~m[389])|(~m[39]&m[245]&m[389]))&~BiasedRNG[84])|((~m[39]&~m[245]&m[389])|(m[39]&~m[245]&m[389])|(m[39]&m[245]&m[389]));
    m[157] = (((~m[39]&~m[257]&~m[401])|(m[39]&m[257]&~m[401]))&BiasedRNG[85])|(((m[39]&~m[257]&~m[401])|(~m[39]&m[257]&m[401]))&~BiasedRNG[85])|((~m[39]&~m[257]&m[401])|(m[39]&~m[257]&m[401])|(m[39]&m[257]&m[401]));
    m[158] = (((~m[39]&~m[269]&~m[413])|(m[39]&m[269]&~m[413]))&BiasedRNG[86])|(((m[39]&~m[269]&~m[413])|(~m[39]&m[269]&m[413]))&~BiasedRNG[86])|((~m[39]&~m[269]&m[413])|(m[39]&~m[269]&m[413])|(m[39]&m[269]&m[413]));
    m[159] = (((~m[39]&~m[281]&~m[425])|(m[39]&m[281]&~m[425]))&BiasedRNG[87])|(((m[39]&~m[281]&~m[425])|(~m[39]&m[281]&m[425]))&~BiasedRNG[87])|((~m[39]&~m[281]&m[425])|(m[39]&~m[281]&m[425])|(m[39]&m[281]&m[425]));
    m[160] = (((~m[40]&~m[293]&~m[437])|(m[40]&m[293]&~m[437]))&BiasedRNG[88])|(((m[40]&~m[293]&~m[437])|(~m[40]&m[293]&m[437]))&~BiasedRNG[88])|((~m[40]&~m[293]&m[437])|(m[40]&~m[293]&m[437])|(m[40]&m[293]&m[437]));
    m[161] = (((~m[40]&~m[305]&~m[449])|(m[40]&m[305]&~m[449]))&BiasedRNG[89])|(((m[40]&~m[305]&~m[449])|(~m[40]&m[305]&m[449]))&~BiasedRNG[89])|((~m[40]&~m[305]&m[449])|(m[40]&~m[305]&m[449])|(m[40]&m[305]&m[449]));
    m[162] = (((~m[40]&~m[317]&~m[461])|(m[40]&m[317]&~m[461]))&BiasedRNG[90])|(((m[40]&~m[317]&~m[461])|(~m[40]&m[317]&m[461]))&~BiasedRNG[90])|((~m[40]&~m[317]&m[461])|(m[40]&~m[317]&m[461])|(m[40]&m[317]&m[461]));
    m[163] = (((~m[40]&~m[329]&~m[473])|(m[40]&m[329]&~m[473]))&BiasedRNG[91])|(((m[40]&~m[329]&~m[473])|(~m[40]&m[329]&m[473]))&~BiasedRNG[91])|((~m[40]&~m[329]&m[473])|(m[40]&~m[329]&m[473])|(m[40]&m[329]&m[473]));
    m[164] = (((~m[41]&~m[341]&~m[485])|(m[41]&m[341]&~m[485]))&BiasedRNG[92])|(((m[41]&~m[341]&~m[485])|(~m[41]&m[341]&m[485]))&~BiasedRNG[92])|((~m[41]&~m[341]&m[485])|(m[41]&~m[341]&m[485])|(m[41]&m[341]&m[485]));
    m[165] = (((~m[41]&~m[353]&~m[497])|(m[41]&m[353]&~m[497]))&BiasedRNG[93])|(((m[41]&~m[353]&~m[497])|(~m[41]&m[353]&m[497]))&~BiasedRNG[93])|((~m[41]&~m[353]&m[497])|(m[41]&~m[353]&m[497])|(m[41]&m[353]&m[497]));
    m[166] = (((~m[41]&~m[365]&~m[509])|(m[41]&m[365]&~m[509]))&BiasedRNG[94])|(((m[41]&~m[365]&~m[509])|(~m[41]&m[365]&m[509]))&~BiasedRNG[94])|((~m[41]&~m[365]&m[509])|(m[41]&~m[365]&m[509])|(m[41]&m[365]&m[509]));
    m[167] = (((~m[41]&~m[377]&~m[521])|(m[41]&m[377]&~m[521]))&BiasedRNG[95])|(((m[41]&~m[377]&~m[521])|(~m[41]&m[377]&m[521]))&~BiasedRNG[95])|((~m[41]&~m[377]&m[521])|(m[41]&~m[377]&m[521])|(m[41]&m[377]&m[521]));
    m[168] = (((~m[42]&~m[246]&~m[390])|(m[42]&m[246]&~m[390]))&BiasedRNG[96])|(((m[42]&~m[246]&~m[390])|(~m[42]&m[246]&m[390]))&~BiasedRNG[96])|((~m[42]&~m[246]&m[390])|(m[42]&~m[246]&m[390])|(m[42]&m[246]&m[390]));
    m[169] = (((~m[42]&~m[258]&~m[402])|(m[42]&m[258]&~m[402]))&BiasedRNG[97])|(((m[42]&~m[258]&~m[402])|(~m[42]&m[258]&m[402]))&~BiasedRNG[97])|((~m[42]&~m[258]&m[402])|(m[42]&~m[258]&m[402])|(m[42]&m[258]&m[402]));
    m[170] = (((~m[42]&~m[270]&~m[414])|(m[42]&m[270]&~m[414]))&BiasedRNG[98])|(((m[42]&~m[270]&~m[414])|(~m[42]&m[270]&m[414]))&~BiasedRNG[98])|((~m[42]&~m[270]&m[414])|(m[42]&~m[270]&m[414])|(m[42]&m[270]&m[414]));
    m[171] = (((~m[42]&~m[282]&~m[426])|(m[42]&m[282]&~m[426]))&BiasedRNG[99])|(((m[42]&~m[282]&~m[426])|(~m[42]&m[282]&m[426]))&~BiasedRNG[99])|((~m[42]&~m[282]&m[426])|(m[42]&~m[282]&m[426])|(m[42]&m[282]&m[426]));
    m[172] = (((~m[43]&~m[294]&~m[438])|(m[43]&m[294]&~m[438]))&BiasedRNG[100])|(((m[43]&~m[294]&~m[438])|(~m[43]&m[294]&m[438]))&~BiasedRNG[100])|((~m[43]&~m[294]&m[438])|(m[43]&~m[294]&m[438])|(m[43]&m[294]&m[438]));
    m[173] = (((~m[43]&~m[306]&~m[450])|(m[43]&m[306]&~m[450]))&BiasedRNG[101])|(((m[43]&~m[306]&~m[450])|(~m[43]&m[306]&m[450]))&~BiasedRNG[101])|((~m[43]&~m[306]&m[450])|(m[43]&~m[306]&m[450])|(m[43]&m[306]&m[450]));
    m[174] = (((~m[43]&~m[318]&~m[462])|(m[43]&m[318]&~m[462]))&BiasedRNG[102])|(((m[43]&~m[318]&~m[462])|(~m[43]&m[318]&m[462]))&~BiasedRNG[102])|((~m[43]&~m[318]&m[462])|(m[43]&~m[318]&m[462])|(m[43]&m[318]&m[462]));
    m[175] = (((~m[43]&~m[330]&~m[474])|(m[43]&m[330]&~m[474]))&BiasedRNG[103])|(((m[43]&~m[330]&~m[474])|(~m[43]&m[330]&m[474]))&~BiasedRNG[103])|((~m[43]&~m[330]&m[474])|(m[43]&~m[330]&m[474])|(m[43]&m[330]&m[474]));
    m[176] = (((~m[44]&~m[342]&~m[486])|(m[44]&m[342]&~m[486]))&BiasedRNG[104])|(((m[44]&~m[342]&~m[486])|(~m[44]&m[342]&m[486]))&~BiasedRNG[104])|((~m[44]&~m[342]&m[486])|(m[44]&~m[342]&m[486])|(m[44]&m[342]&m[486]));
    m[177] = (((~m[44]&~m[354]&~m[498])|(m[44]&m[354]&~m[498]))&BiasedRNG[105])|(((m[44]&~m[354]&~m[498])|(~m[44]&m[354]&m[498]))&~BiasedRNG[105])|((~m[44]&~m[354]&m[498])|(m[44]&~m[354]&m[498])|(m[44]&m[354]&m[498]));
    m[178] = (((~m[44]&~m[366]&~m[510])|(m[44]&m[366]&~m[510]))&BiasedRNG[106])|(((m[44]&~m[366]&~m[510])|(~m[44]&m[366]&m[510]))&~BiasedRNG[106])|((~m[44]&~m[366]&m[510])|(m[44]&~m[366]&m[510])|(m[44]&m[366]&m[510]));
    m[179] = (((~m[44]&~m[378]&~m[522])|(m[44]&m[378]&~m[522]))&BiasedRNG[107])|(((m[44]&~m[378]&~m[522])|(~m[44]&m[378]&m[522]))&~BiasedRNG[107])|((~m[44]&~m[378]&m[522])|(m[44]&~m[378]&m[522])|(m[44]&m[378]&m[522]));
    m[180] = (((~m[45]&~m[247]&~m[391])|(m[45]&m[247]&~m[391]))&BiasedRNG[108])|(((m[45]&~m[247]&~m[391])|(~m[45]&m[247]&m[391]))&~BiasedRNG[108])|((~m[45]&~m[247]&m[391])|(m[45]&~m[247]&m[391])|(m[45]&m[247]&m[391]));
    m[181] = (((~m[45]&~m[259]&~m[403])|(m[45]&m[259]&~m[403]))&BiasedRNG[109])|(((m[45]&~m[259]&~m[403])|(~m[45]&m[259]&m[403]))&~BiasedRNG[109])|((~m[45]&~m[259]&m[403])|(m[45]&~m[259]&m[403])|(m[45]&m[259]&m[403]));
    m[182] = (((~m[45]&~m[271]&~m[415])|(m[45]&m[271]&~m[415]))&BiasedRNG[110])|(((m[45]&~m[271]&~m[415])|(~m[45]&m[271]&m[415]))&~BiasedRNG[110])|((~m[45]&~m[271]&m[415])|(m[45]&~m[271]&m[415])|(m[45]&m[271]&m[415]));
    m[183] = (((~m[45]&~m[283]&~m[427])|(m[45]&m[283]&~m[427]))&BiasedRNG[111])|(((m[45]&~m[283]&~m[427])|(~m[45]&m[283]&m[427]))&~BiasedRNG[111])|((~m[45]&~m[283]&m[427])|(m[45]&~m[283]&m[427])|(m[45]&m[283]&m[427]));
    m[184] = (((~m[46]&~m[295]&~m[439])|(m[46]&m[295]&~m[439]))&BiasedRNG[112])|(((m[46]&~m[295]&~m[439])|(~m[46]&m[295]&m[439]))&~BiasedRNG[112])|((~m[46]&~m[295]&m[439])|(m[46]&~m[295]&m[439])|(m[46]&m[295]&m[439]));
    m[185] = (((~m[46]&~m[307]&~m[451])|(m[46]&m[307]&~m[451]))&BiasedRNG[113])|(((m[46]&~m[307]&~m[451])|(~m[46]&m[307]&m[451]))&~BiasedRNG[113])|((~m[46]&~m[307]&m[451])|(m[46]&~m[307]&m[451])|(m[46]&m[307]&m[451]));
    m[186] = (((~m[46]&~m[319]&~m[463])|(m[46]&m[319]&~m[463]))&BiasedRNG[114])|(((m[46]&~m[319]&~m[463])|(~m[46]&m[319]&m[463]))&~BiasedRNG[114])|((~m[46]&~m[319]&m[463])|(m[46]&~m[319]&m[463])|(m[46]&m[319]&m[463]));
    m[187] = (((~m[46]&~m[331]&~m[475])|(m[46]&m[331]&~m[475]))&BiasedRNG[115])|(((m[46]&~m[331]&~m[475])|(~m[46]&m[331]&m[475]))&~BiasedRNG[115])|((~m[46]&~m[331]&m[475])|(m[46]&~m[331]&m[475])|(m[46]&m[331]&m[475]));
    m[188] = (((~m[47]&~m[343]&~m[487])|(m[47]&m[343]&~m[487]))&BiasedRNG[116])|(((m[47]&~m[343]&~m[487])|(~m[47]&m[343]&m[487]))&~BiasedRNG[116])|((~m[47]&~m[343]&m[487])|(m[47]&~m[343]&m[487])|(m[47]&m[343]&m[487]));
    m[189] = (((~m[47]&~m[355]&~m[499])|(m[47]&m[355]&~m[499]))&BiasedRNG[117])|(((m[47]&~m[355]&~m[499])|(~m[47]&m[355]&m[499]))&~BiasedRNG[117])|((~m[47]&~m[355]&m[499])|(m[47]&~m[355]&m[499])|(m[47]&m[355]&m[499]));
    m[190] = (((~m[47]&~m[367]&~m[511])|(m[47]&m[367]&~m[511]))&BiasedRNG[118])|(((m[47]&~m[367]&~m[511])|(~m[47]&m[367]&m[511]))&~BiasedRNG[118])|((~m[47]&~m[367]&m[511])|(m[47]&~m[367]&m[511])|(m[47]&m[367]&m[511]));
    m[191] = (((~m[47]&~m[379]&~m[523])|(m[47]&m[379]&~m[523]))&BiasedRNG[119])|(((m[47]&~m[379]&~m[523])|(~m[47]&m[379]&m[523]))&~BiasedRNG[119])|((~m[47]&~m[379]&m[523])|(m[47]&~m[379]&m[523])|(m[47]&m[379]&m[523]));
    m[192] = (((~m[48]&~m[248]&~m[392])|(m[48]&m[248]&~m[392]))&BiasedRNG[120])|(((m[48]&~m[248]&~m[392])|(~m[48]&m[248]&m[392]))&~BiasedRNG[120])|((~m[48]&~m[248]&m[392])|(m[48]&~m[248]&m[392])|(m[48]&m[248]&m[392]));
    m[193] = (((~m[48]&~m[260]&~m[404])|(m[48]&m[260]&~m[404]))&BiasedRNG[121])|(((m[48]&~m[260]&~m[404])|(~m[48]&m[260]&m[404]))&~BiasedRNG[121])|((~m[48]&~m[260]&m[404])|(m[48]&~m[260]&m[404])|(m[48]&m[260]&m[404]));
    m[194] = (((~m[48]&~m[272]&~m[416])|(m[48]&m[272]&~m[416]))&BiasedRNG[122])|(((m[48]&~m[272]&~m[416])|(~m[48]&m[272]&m[416]))&~BiasedRNG[122])|((~m[48]&~m[272]&m[416])|(m[48]&~m[272]&m[416])|(m[48]&m[272]&m[416]));
    m[195] = (((~m[48]&~m[284]&~m[428])|(m[48]&m[284]&~m[428]))&BiasedRNG[123])|(((m[48]&~m[284]&~m[428])|(~m[48]&m[284]&m[428]))&~BiasedRNG[123])|((~m[48]&~m[284]&m[428])|(m[48]&~m[284]&m[428])|(m[48]&m[284]&m[428]));
    m[196] = (((~m[49]&~m[296]&~m[440])|(m[49]&m[296]&~m[440]))&BiasedRNG[124])|(((m[49]&~m[296]&~m[440])|(~m[49]&m[296]&m[440]))&~BiasedRNG[124])|((~m[49]&~m[296]&m[440])|(m[49]&~m[296]&m[440])|(m[49]&m[296]&m[440]));
    m[197] = (((~m[49]&~m[308]&~m[452])|(m[49]&m[308]&~m[452]))&BiasedRNG[125])|(((m[49]&~m[308]&~m[452])|(~m[49]&m[308]&m[452]))&~BiasedRNG[125])|((~m[49]&~m[308]&m[452])|(m[49]&~m[308]&m[452])|(m[49]&m[308]&m[452]));
    m[198] = (((~m[49]&~m[320]&~m[464])|(m[49]&m[320]&~m[464]))&BiasedRNG[126])|(((m[49]&~m[320]&~m[464])|(~m[49]&m[320]&m[464]))&~BiasedRNG[126])|((~m[49]&~m[320]&m[464])|(m[49]&~m[320]&m[464])|(m[49]&m[320]&m[464]));
    m[199] = (((~m[49]&~m[332]&~m[476])|(m[49]&m[332]&~m[476]))&BiasedRNG[127])|(((m[49]&~m[332]&~m[476])|(~m[49]&m[332]&m[476]))&~BiasedRNG[127])|((~m[49]&~m[332]&m[476])|(m[49]&~m[332]&m[476])|(m[49]&m[332]&m[476]));
    m[200] = (((~m[50]&~m[344]&~m[488])|(m[50]&m[344]&~m[488]))&BiasedRNG[128])|(((m[50]&~m[344]&~m[488])|(~m[50]&m[344]&m[488]))&~BiasedRNG[128])|((~m[50]&~m[344]&m[488])|(m[50]&~m[344]&m[488])|(m[50]&m[344]&m[488]));
    m[201] = (((~m[50]&~m[356]&~m[500])|(m[50]&m[356]&~m[500]))&BiasedRNG[129])|(((m[50]&~m[356]&~m[500])|(~m[50]&m[356]&m[500]))&~BiasedRNG[129])|((~m[50]&~m[356]&m[500])|(m[50]&~m[356]&m[500])|(m[50]&m[356]&m[500]));
    m[202] = (((~m[50]&~m[368]&~m[512])|(m[50]&m[368]&~m[512]))&BiasedRNG[130])|(((m[50]&~m[368]&~m[512])|(~m[50]&m[368]&m[512]))&~BiasedRNG[130])|((~m[50]&~m[368]&m[512])|(m[50]&~m[368]&m[512])|(m[50]&m[368]&m[512]));
    m[203] = (((~m[50]&~m[380]&~m[524])|(m[50]&m[380]&~m[524]))&BiasedRNG[131])|(((m[50]&~m[380]&~m[524])|(~m[50]&m[380]&m[524]))&~BiasedRNG[131])|((~m[50]&~m[380]&m[524])|(m[50]&~m[380]&m[524])|(m[50]&m[380]&m[524]));
    m[204] = (((~m[51]&~m[249]&~m[393])|(m[51]&m[249]&~m[393]))&BiasedRNG[132])|(((m[51]&~m[249]&~m[393])|(~m[51]&m[249]&m[393]))&~BiasedRNG[132])|((~m[51]&~m[249]&m[393])|(m[51]&~m[249]&m[393])|(m[51]&m[249]&m[393]));
    m[205] = (((~m[51]&~m[261]&~m[405])|(m[51]&m[261]&~m[405]))&BiasedRNG[133])|(((m[51]&~m[261]&~m[405])|(~m[51]&m[261]&m[405]))&~BiasedRNG[133])|((~m[51]&~m[261]&m[405])|(m[51]&~m[261]&m[405])|(m[51]&m[261]&m[405]));
    m[206] = (((~m[51]&~m[273]&~m[417])|(m[51]&m[273]&~m[417]))&BiasedRNG[134])|(((m[51]&~m[273]&~m[417])|(~m[51]&m[273]&m[417]))&~BiasedRNG[134])|((~m[51]&~m[273]&m[417])|(m[51]&~m[273]&m[417])|(m[51]&m[273]&m[417]));
    m[207] = (((~m[51]&~m[285]&~m[429])|(m[51]&m[285]&~m[429]))&BiasedRNG[135])|(((m[51]&~m[285]&~m[429])|(~m[51]&m[285]&m[429]))&~BiasedRNG[135])|((~m[51]&~m[285]&m[429])|(m[51]&~m[285]&m[429])|(m[51]&m[285]&m[429]));
    m[208] = (((~m[52]&~m[297]&~m[441])|(m[52]&m[297]&~m[441]))&BiasedRNG[136])|(((m[52]&~m[297]&~m[441])|(~m[52]&m[297]&m[441]))&~BiasedRNG[136])|((~m[52]&~m[297]&m[441])|(m[52]&~m[297]&m[441])|(m[52]&m[297]&m[441]));
    m[209] = (((~m[52]&~m[309]&~m[453])|(m[52]&m[309]&~m[453]))&BiasedRNG[137])|(((m[52]&~m[309]&~m[453])|(~m[52]&m[309]&m[453]))&~BiasedRNG[137])|((~m[52]&~m[309]&m[453])|(m[52]&~m[309]&m[453])|(m[52]&m[309]&m[453]));
    m[210] = (((~m[52]&~m[321]&~m[465])|(m[52]&m[321]&~m[465]))&BiasedRNG[138])|(((m[52]&~m[321]&~m[465])|(~m[52]&m[321]&m[465]))&~BiasedRNG[138])|((~m[52]&~m[321]&m[465])|(m[52]&~m[321]&m[465])|(m[52]&m[321]&m[465]));
    m[211] = (((~m[52]&~m[333]&~m[477])|(m[52]&m[333]&~m[477]))&BiasedRNG[139])|(((m[52]&~m[333]&~m[477])|(~m[52]&m[333]&m[477]))&~BiasedRNG[139])|((~m[52]&~m[333]&m[477])|(m[52]&~m[333]&m[477])|(m[52]&m[333]&m[477]));
    m[212] = (((~m[53]&~m[345]&~m[489])|(m[53]&m[345]&~m[489]))&BiasedRNG[140])|(((m[53]&~m[345]&~m[489])|(~m[53]&m[345]&m[489]))&~BiasedRNG[140])|((~m[53]&~m[345]&m[489])|(m[53]&~m[345]&m[489])|(m[53]&m[345]&m[489]));
    m[213] = (((~m[53]&~m[357]&~m[501])|(m[53]&m[357]&~m[501]))&BiasedRNG[141])|(((m[53]&~m[357]&~m[501])|(~m[53]&m[357]&m[501]))&~BiasedRNG[141])|((~m[53]&~m[357]&m[501])|(m[53]&~m[357]&m[501])|(m[53]&m[357]&m[501]));
    m[214] = (((~m[53]&~m[369]&~m[513])|(m[53]&m[369]&~m[513]))&BiasedRNG[142])|(((m[53]&~m[369]&~m[513])|(~m[53]&m[369]&m[513]))&~BiasedRNG[142])|((~m[53]&~m[369]&m[513])|(m[53]&~m[369]&m[513])|(m[53]&m[369]&m[513]));
    m[215] = (((~m[53]&~m[381]&~m[525])|(m[53]&m[381]&~m[525]))&BiasedRNG[143])|(((m[53]&~m[381]&~m[525])|(~m[53]&m[381]&m[525]))&~BiasedRNG[143])|((~m[53]&~m[381]&m[525])|(m[53]&~m[381]&m[525])|(m[53]&m[381]&m[525]));
    m[216] = (((~m[54]&~m[250]&~m[394])|(m[54]&m[250]&~m[394]))&BiasedRNG[144])|(((m[54]&~m[250]&~m[394])|(~m[54]&m[250]&m[394]))&~BiasedRNG[144])|((~m[54]&~m[250]&m[394])|(m[54]&~m[250]&m[394])|(m[54]&m[250]&m[394]));
    m[217] = (((~m[54]&~m[262]&~m[406])|(m[54]&m[262]&~m[406]))&BiasedRNG[145])|(((m[54]&~m[262]&~m[406])|(~m[54]&m[262]&m[406]))&~BiasedRNG[145])|((~m[54]&~m[262]&m[406])|(m[54]&~m[262]&m[406])|(m[54]&m[262]&m[406]));
    m[218] = (((~m[54]&~m[274]&~m[418])|(m[54]&m[274]&~m[418]))&BiasedRNG[146])|(((m[54]&~m[274]&~m[418])|(~m[54]&m[274]&m[418]))&~BiasedRNG[146])|((~m[54]&~m[274]&m[418])|(m[54]&~m[274]&m[418])|(m[54]&m[274]&m[418]));
    m[219] = (((~m[54]&~m[286]&~m[430])|(m[54]&m[286]&~m[430]))&BiasedRNG[147])|(((m[54]&~m[286]&~m[430])|(~m[54]&m[286]&m[430]))&~BiasedRNG[147])|((~m[54]&~m[286]&m[430])|(m[54]&~m[286]&m[430])|(m[54]&m[286]&m[430]));
    m[220] = (((~m[55]&~m[298]&~m[442])|(m[55]&m[298]&~m[442]))&BiasedRNG[148])|(((m[55]&~m[298]&~m[442])|(~m[55]&m[298]&m[442]))&~BiasedRNG[148])|((~m[55]&~m[298]&m[442])|(m[55]&~m[298]&m[442])|(m[55]&m[298]&m[442]));
    m[221] = (((~m[55]&~m[310]&~m[454])|(m[55]&m[310]&~m[454]))&BiasedRNG[149])|(((m[55]&~m[310]&~m[454])|(~m[55]&m[310]&m[454]))&~BiasedRNG[149])|((~m[55]&~m[310]&m[454])|(m[55]&~m[310]&m[454])|(m[55]&m[310]&m[454]));
    m[222] = (((~m[55]&~m[322]&~m[466])|(m[55]&m[322]&~m[466]))&BiasedRNG[150])|(((m[55]&~m[322]&~m[466])|(~m[55]&m[322]&m[466]))&~BiasedRNG[150])|((~m[55]&~m[322]&m[466])|(m[55]&~m[322]&m[466])|(m[55]&m[322]&m[466]));
    m[223] = (((~m[55]&~m[334]&~m[478])|(m[55]&m[334]&~m[478]))&BiasedRNG[151])|(((m[55]&~m[334]&~m[478])|(~m[55]&m[334]&m[478]))&~BiasedRNG[151])|((~m[55]&~m[334]&m[478])|(m[55]&~m[334]&m[478])|(m[55]&m[334]&m[478]));
    m[224] = (((~m[56]&~m[346]&~m[490])|(m[56]&m[346]&~m[490]))&BiasedRNG[152])|(((m[56]&~m[346]&~m[490])|(~m[56]&m[346]&m[490]))&~BiasedRNG[152])|((~m[56]&~m[346]&m[490])|(m[56]&~m[346]&m[490])|(m[56]&m[346]&m[490]));
    m[225] = (((~m[56]&~m[358]&~m[502])|(m[56]&m[358]&~m[502]))&BiasedRNG[153])|(((m[56]&~m[358]&~m[502])|(~m[56]&m[358]&m[502]))&~BiasedRNG[153])|((~m[56]&~m[358]&m[502])|(m[56]&~m[358]&m[502])|(m[56]&m[358]&m[502]));
    m[226] = (((~m[56]&~m[370]&~m[514])|(m[56]&m[370]&~m[514]))&BiasedRNG[154])|(((m[56]&~m[370]&~m[514])|(~m[56]&m[370]&m[514]))&~BiasedRNG[154])|((~m[56]&~m[370]&m[514])|(m[56]&~m[370]&m[514])|(m[56]&m[370]&m[514]));
    m[227] = (((~m[56]&~m[382]&~m[526])|(m[56]&m[382]&~m[526]))&BiasedRNG[155])|(((m[56]&~m[382]&~m[526])|(~m[56]&m[382]&m[526]))&~BiasedRNG[155])|((~m[56]&~m[382]&m[526])|(m[56]&~m[382]&m[526])|(m[56]&m[382]&m[526]));
    m[228] = (((~m[57]&~m[251]&~m[395])|(m[57]&m[251]&~m[395]))&BiasedRNG[156])|(((m[57]&~m[251]&~m[395])|(~m[57]&m[251]&m[395]))&~BiasedRNG[156])|((~m[57]&~m[251]&m[395])|(m[57]&~m[251]&m[395])|(m[57]&m[251]&m[395]));
    m[229] = (((~m[57]&~m[263]&~m[407])|(m[57]&m[263]&~m[407]))&BiasedRNG[157])|(((m[57]&~m[263]&~m[407])|(~m[57]&m[263]&m[407]))&~BiasedRNG[157])|((~m[57]&~m[263]&m[407])|(m[57]&~m[263]&m[407])|(m[57]&m[263]&m[407]));
    m[230] = (((~m[57]&~m[275]&~m[419])|(m[57]&m[275]&~m[419]))&BiasedRNG[158])|(((m[57]&~m[275]&~m[419])|(~m[57]&m[275]&m[419]))&~BiasedRNG[158])|((~m[57]&~m[275]&m[419])|(m[57]&~m[275]&m[419])|(m[57]&m[275]&m[419]));
    m[231] = (((~m[57]&~m[287]&~m[431])|(m[57]&m[287]&~m[431]))&BiasedRNG[159])|(((m[57]&~m[287]&~m[431])|(~m[57]&m[287]&m[431]))&~BiasedRNG[159])|((~m[57]&~m[287]&m[431])|(m[57]&~m[287]&m[431])|(m[57]&m[287]&m[431]));
    m[232] = (((~m[58]&~m[299]&~m[443])|(m[58]&m[299]&~m[443]))&BiasedRNG[160])|(((m[58]&~m[299]&~m[443])|(~m[58]&m[299]&m[443]))&~BiasedRNG[160])|((~m[58]&~m[299]&m[443])|(m[58]&~m[299]&m[443])|(m[58]&m[299]&m[443]));
    m[233] = (((~m[58]&~m[311]&~m[455])|(m[58]&m[311]&~m[455]))&BiasedRNG[161])|(((m[58]&~m[311]&~m[455])|(~m[58]&m[311]&m[455]))&~BiasedRNG[161])|((~m[58]&~m[311]&m[455])|(m[58]&~m[311]&m[455])|(m[58]&m[311]&m[455]));
    m[234] = (((~m[58]&~m[323]&~m[467])|(m[58]&m[323]&~m[467]))&BiasedRNG[162])|(((m[58]&~m[323]&~m[467])|(~m[58]&m[323]&m[467]))&~BiasedRNG[162])|((~m[58]&~m[323]&m[467])|(m[58]&~m[323]&m[467])|(m[58]&m[323]&m[467]));
    m[235] = (((~m[58]&~m[335]&~m[479])|(m[58]&m[335]&~m[479]))&BiasedRNG[163])|(((m[58]&~m[335]&~m[479])|(~m[58]&m[335]&m[479]))&~BiasedRNG[163])|((~m[58]&~m[335]&m[479])|(m[58]&~m[335]&m[479])|(m[58]&m[335]&m[479]));
    m[236] = (((~m[59]&~m[347]&~m[491])|(m[59]&m[347]&~m[491]))&BiasedRNG[164])|(((m[59]&~m[347]&~m[491])|(~m[59]&m[347]&m[491]))&~BiasedRNG[164])|((~m[59]&~m[347]&m[491])|(m[59]&~m[347]&m[491])|(m[59]&m[347]&m[491]));
    m[237] = (((~m[59]&~m[359]&~m[503])|(m[59]&m[359]&~m[503]))&BiasedRNG[165])|(((m[59]&~m[359]&~m[503])|(~m[59]&m[359]&m[503]))&~BiasedRNG[165])|((~m[59]&~m[359]&m[503])|(m[59]&~m[359]&m[503])|(m[59]&m[359]&m[503]));
    m[238] = (((~m[59]&~m[371]&~m[515])|(m[59]&m[371]&~m[515]))&BiasedRNG[166])|(((m[59]&~m[371]&~m[515])|(~m[59]&m[371]&m[515]))&~BiasedRNG[166])|((~m[59]&~m[371]&m[515])|(m[59]&~m[371]&m[515])|(m[59]&m[371]&m[515]));
    m[239] = (((~m[59]&~m[383]&~m[527])|(m[59]&m[383]&~m[527]))&BiasedRNG[167])|(((m[59]&~m[383]&~m[527])|(~m[59]&m[383]&m[527]))&~BiasedRNG[167])|((~m[59]&~m[383]&m[527])|(m[59]&~m[383]&m[527])|(m[59]&m[383]&m[527]));
    m[528] = (((m[385]&~m[529]&~m[530]&~m[531]&~m[532])|(~m[385]&~m[529]&~m[530]&m[531]&~m[532])|(m[385]&m[529]&~m[530]&m[531]&~m[532])|(m[385]&~m[529]&m[530]&m[531]&~m[532])|(~m[385]&m[529]&~m[530]&~m[531]&m[532])|(~m[385]&~m[529]&m[530]&~m[531]&m[532])|(m[385]&m[529]&m[530]&~m[531]&m[532])|(~m[385]&m[529]&m[530]&m[531]&m[532]))&UnbiasedRNG[0])|((m[385]&~m[529]&~m[530]&m[531]&~m[532])|(~m[385]&~m[529]&~m[530]&~m[531]&m[532])|(m[385]&~m[529]&~m[530]&~m[531]&m[532])|(m[385]&m[529]&~m[530]&~m[531]&m[532])|(m[385]&~m[529]&m[530]&~m[531]&m[532])|(~m[385]&~m[529]&~m[530]&m[531]&m[532])|(m[385]&~m[529]&~m[530]&m[531]&m[532])|(~m[385]&m[529]&~m[530]&m[531]&m[532])|(m[385]&m[529]&~m[530]&m[531]&m[532])|(~m[385]&~m[529]&m[530]&m[531]&m[532])|(m[385]&~m[529]&m[530]&m[531]&m[532])|(m[385]&m[529]&m[530]&m[531]&m[532]));
    m[533] = (((m[386]&~m[534]&~m[535]&~m[536]&~m[537])|(~m[386]&~m[534]&~m[535]&m[536]&~m[537])|(m[386]&m[534]&~m[535]&m[536]&~m[537])|(m[386]&~m[534]&m[535]&m[536]&~m[537])|(~m[386]&m[534]&~m[535]&~m[536]&m[537])|(~m[386]&~m[534]&m[535]&~m[536]&m[537])|(m[386]&m[534]&m[535]&~m[536]&m[537])|(~m[386]&m[534]&m[535]&m[536]&m[537]))&UnbiasedRNG[1])|((m[386]&~m[534]&~m[535]&m[536]&~m[537])|(~m[386]&~m[534]&~m[535]&~m[536]&m[537])|(m[386]&~m[534]&~m[535]&~m[536]&m[537])|(m[386]&m[534]&~m[535]&~m[536]&m[537])|(m[386]&~m[534]&m[535]&~m[536]&m[537])|(~m[386]&~m[534]&~m[535]&m[536]&m[537])|(m[386]&~m[534]&~m[535]&m[536]&m[537])|(~m[386]&m[534]&~m[535]&m[536]&m[537])|(m[386]&m[534]&~m[535]&m[536]&m[537])|(~m[386]&~m[534]&m[535]&m[536]&m[537])|(m[386]&~m[534]&m[535]&m[536]&m[537])|(m[386]&m[534]&m[535]&m[536]&m[537]));
    m[538] = (((m[536]&~m[539]&~m[540]&~m[541]&~m[542])|(~m[536]&~m[539]&~m[540]&m[541]&~m[542])|(m[536]&m[539]&~m[540]&m[541]&~m[542])|(m[536]&~m[539]&m[540]&m[541]&~m[542])|(~m[536]&m[539]&~m[540]&~m[541]&m[542])|(~m[536]&~m[539]&m[540]&~m[541]&m[542])|(m[536]&m[539]&m[540]&~m[541]&m[542])|(~m[536]&m[539]&m[540]&m[541]&m[542]))&UnbiasedRNG[2])|((m[536]&~m[539]&~m[540]&m[541]&~m[542])|(~m[536]&~m[539]&~m[540]&~m[541]&m[542])|(m[536]&~m[539]&~m[540]&~m[541]&m[542])|(m[536]&m[539]&~m[540]&~m[541]&m[542])|(m[536]&~m[539]&m[540]&~m[541]&m[542])|(~m[536]&~m[539]&~m[540]&m[541]&m[542])|(m[536]&~m[539]&~m[540]&m[541]&m[542])|(~m[536]&m[539]&~m[540]&m[541]&m[542])|(m[536]&m[539]&~m[540]&m[541]&m[542])|(~m[536]&~m[539]&m[540]&m[541]&m[542])|(m[536]&~m[539]&m[540]&m[541]&m[542])|(m[536]&m[539]&m[540]&m[541]&m[542]));
    m[543] = (((m[387]&~m[544]&~m[545]&~m[546]&~m[547])|(~m[387]&~m[544]&~m[545]&m[546]&~m[547])|(m[387]&m[544]&~m[545]&m[546]&~m[547])|(m[387]&~m[544]&m[545]&m[546]&~m[547])|(~m[387]&m[544]&~m[545]&~m[546]&m[547])|(~m[387]&~m[544]&m[545]&~m[546]&m[547])|(m[387]&m[544]&m[545]&~m[546]&m[547])|(~m[387]&m[544]&m[545]&m[546]&m[547]))&UnbiasedRNG[3])|((m[387]&~m[544]&~m[545]&m[546]&~m[547])|(~m[387]&~m[544]&~m[545]&~m[546]&m[547])|(m[387]&~m[544]&~m[545]&~m[546]&m[547])|(m[387]&m[544]&~m[545]&~m[546]&m[547])|(m[387]&~m[544]&m[545]&~m[546]&m[547])|(~m[387]&~m[544]&~m[545]&m[546]&m[547])|(m[387]&~m[544]&~m[545]&m[546]&m[547])|(~m[387]&m[544]&~m[545]&m[546]&m[547])|(m[387]&m[544]&~m[545]&m[546]&m[547])|(~m[387]&~m[544]&m[545]&m[546]&m[547])|(m[387]&~m[544]&m[545]&m[546]&m[547])|(m[387]&m[544]&m[545]&m[546]&m[547]));
    m[548] = (((m[546]&~m[549]&~m[550]&~m[551]&~m[552])|(~m[546]&~m[549]&~m[550]&m[551]&~m[552])|(m[546]&m[549]&~m[550]&m[551]&~m[552])|(m[546]&~m[549]&m[550]&m[551]&~m[552])|(~m[546]&m[549]&~m[550]&~m[551]&m[552])|(~m[546]&~m[549]&m[550]&~m[551]&m[552])|(m[546]&m[549]&m[550]&~m[551]&m[552])|(~m[546]&m[549]&m[550]&m[551]&m[552]))&UnbiasedRNG[4])|((m[546]&~m[549]&~m[550]&m[551]&~m[552])|(~m[546]&~m[549]&~m[550]&~m[551]&m[552])|(m[546]&~m[549]&~m[550]&~m[551]&m[552])|(m[546]&m[549]&~m[550]&~m[551]&m[552])|(m[546]&~m[549]&m[550]&~m[551]&m[552])|(~m[546]&~m[549]&~m[550]&m[551]&m[552])|(m[546]&~m[549]&~m[550]&m[551]&m[552])|(~m[546]&m[549]&~m[550]&m[551]&m[552])|(m[546]&m[549]&~m[550]&m[551]&m[552])|(~m[546]&~m[549]&m[550]&m[551]&m[552])|(m[546]&~m[549]&m[550]&m[551]&m[552])|(m[546]&m[549]&m[550]&m[551]&m[552]));
    m[553] = (((m[551]&~m[554]&~m[555]&~m[556]&~m[557])|(~m[551]&~m[554]&~m[555]&m[556]&~m[557])|(m[551]&m[554]&~m[555]&m[556]&~m[557])|(m[551]&~m[554]&m[555]&m[556]&~m[557])|(~m[551]&m[554]&~m[555]&~m[556]&m[557])|(~m[551]&~m[554]&m[555]&~m[556]&m[557])|(m[551]&m[554]&m[555]&~m[556]&m[557])|(~m[551]&m[554]&m[555]&m[556]&m[557]))&UnbiasedRNG[5])|((m[551]&~m[554]&~m[555]&m[556]&~m[557])|(~m[551]&~m[554]&~m[555]&~m[556]&m[557])|(m[551]&~m[554]&~m[555]&~m[556]&m[557])|(m[551]&m[554]&~m[555]&~m[556]&m[557])|(m[551]&~m[554]&m[555]&~m[556]&m[557])|(~m[551]&~m[554]&~m[555]&m[556]&m[557])|(m[551]&~m[554]&~m[555]&m[556]&m[557])|(~m[551]&m[554]&~m[555]&m[556]&m[557])|(m[551]&m[554]&~m[555]&m[556]&m[557])|(~m[551]&~m[554]&m[555]&m[556]&m[557])|(m[551]&~m[554]&m[555]&m[556]&m[557])|(m[551]&m[554]&m[555]&m[556]&m[557]));
    m[558] = (((m[388]&~m[559]&~m[560]&~m[561]&~m[562])|(~m[388]&~m[559]&~m[560]&m[561]&~m[562])|(m[388]&m[559]&~m[560]&m[561]&~m[562])|(m[388]&~m[559]&m[560]&m[561]&~m[562])|(~m[388]&m[559]&~m[560]&~m[561]&m[562])|(~m[388]&~m[559]&m[560]&~m[561]&m[562])|(m[388]&m[559]&m[560]&~m[561]&m[562])|(~m[388]&m[559]&m[560]&m[561]&m[562]))&UnbiasedRNG[6])|((m[388]&~m[559]&~m[560]&m[561]&~m[562])|(~m[388]&~m[559]&~m[560]&~m[561]&m[562])|(m[388]&~m[559]&~m[560]&~m[561]&m[562])|(m[388]&m[559]&~m[560]&~m[561]&m[562])|(m[388]&~m[559]&m[560]&~m[561]&m[562])|(~m[388]&~m[559]&~m[560]&m[561]&m[562])|(m[388]&~m[559]&~m[560]&m[561]&m[562])|(~m[388]&m[559]&~m[560]&m[561]&m[562])|(m[388]&m[559]&~m[560]&m[561]&m[562])|(~m[388]&~m[559]&m[560]&m[561]&m[562])|(m[388]&~m[559]&m[560]&m[561]&m[562])|(m[388]&m[559]&m[560]&m[561]&m[562]));
    m[563] = (((m[561]&~m[564]&~m[565]&~m[566]&~m[567])|(~m[561]&~m[564]&~m[565]&m[566]&~m[567])|(m[561]&m[564]&~m[565]&m[566]&~m[567])|(m[561]&~m[564]&m[565]&m[566]&~m[567])|(~m[561]&m[564]&~m[565]&~m[566]&m[567])|(~m[561]&~m[564]&m[565]&~m[566]&m[567])|(m[561]&m[564]&m[565]&~m[566]&m[567])|(~m[561]&m[564]&m[565]&m[566]&m[567]))&UnbiasedRNG[7])|((m[561]&~m[564]&~m[565]&m[566]&~m[567])|(~m[561]&~m[564]&~m[565]&~m[566]&m[567])|(m[561]&~m[564]&~m[565]&~m[566]&m[567])|(m[561]&m[564]&~m[565]&~m[566]&m[567])|(m[561]&~m[564]&m[565]&~m[566]&m[567])|(~m[561]&~m[564]&~m[565]&m[566]&m[567])|(m[561]&~m[564]&~m[565]&m[566]&m[567])|(~m[561]&m[564]&~m[565]&m[566]&m[567])|(m[561]&m[564]&~m[565]&m[566]&m[567])|(~m[561]&~m[564]&m[565]&m[566]&m[567])|(m[561]&~m[564]&m[565]&m[566]&m[567])|(m[561]&m[564]&m[565]&m[566]&m[567]));
    m[568] = (((m[566]&~m[569]&~m[570]&~m[571]&~m[572])|(~m[566]&~m[569]&~m[570]&m[571]&~m[572])|(m[566]&m[569]&~m[570]&m[571]&~m[572])|(m[566]&~m[569]&m[570]&m[571]&~m[572])|(~m[566]&m[569]&~m[570]&~m[571]&m[572])|(~m[566]&~m[569]&m[570]&~m[571]&m[572])|(m[566]&m[569]&m[570]&~m[571]&m[572])|(~m[566]&m[569]&m[570]&m[571]&m[572]))&UnbiasedRNG[8])|((m[566]&~m[569]&~m[570]&m[571]&~m[572])|(~m[566]&~m[569]&~m[570]&~m[571]&m[572])|(m[566]&~m[569]&~m[570]&~m[571]&m[572])|(m[566]&m[569]&~m[570]&~m[571]&m[572])|(m[566]&~m[569]&m[570]&~m[571]&m[572])|(~m[566]&~m[569]&~m[570]&m[571]&m[572])|(m[566]&~m[569]&~m[570]&m[571]&m[572])|(~m[566]&m[569]&~m[570]&m[571]&m[572])|(m[566]&m[569]&~m[570]&m[571]&m[572])|(~m[566]&~m[569]&m[570]&m[571]&m[572])|(m[566]&~m[569]&m[570]&m[571]&m[572])|(m[566]&m[569]&m[570]&m[571]&m[572]));
    m[573] = (((m[571]&~m[574]&~m[575]&~m[576]&~m[577])|(~m[571]&~m[574]&~m[575]&m[576]&~m[577])|(m[571]&m[574]&~m[575]&m[576]&~m[577])|(m[571]&~m[574]&m[575]&m[576]&~m[577])|(~m[571]&m[574]&~m[575]&~m[576]&m[577])|(~m[571]&~m[574]&m[575]&~m[576]&m[577])|(m[571]&m[574]&m[575]&~m[576]&m[577])|(~m[571]&m[574]&m[575]&m[576]&m[577]))&UnbiasedRNG[9])|((m[571]&~m[574]&~m[575]&m[576]&~m[577])|(~m[571]&~m[574]&~m[575]&~m[576]&m[577])|(m[571]&~m[574]&~m[575]&~m[576]&m[577])|(m[571]&m[574]&~m[575]&~m[576]&m[577])|(m[571]&~m[574]&m[575]&~m[576]&m[577])|(~m[571]&~m[574]&~m[575]&m[576]&m[577])|(m[571]&~m[574]&~m[575]&m[576]&m[577])|(~m[571]&m[574]&~m[575]&m[576]&m[577])|(m[571]&m[574]&~m[575]&m[576]&m[577])|(~m[571]&~m[574]&m[575]&m[576]&m[577])|(m[571]&~m[574]&m[575]&m[576]&m[577])|(m[571]&m[574]&m[575]&m[576]&m[577]));
    m[578] = (((m[389]&~m[579]&~m[580]&~m[581]&~m[582])|(~m[389]&~m[579]&~m[580]&m[581]&~m[582])|(m[389]&m[579]&~m[580]&m[581]&~m[582])|(m[389]&~m[579]&m[580]&m[581]&~m[582])|(~m[389]&m[579]&~m[580]&~m[581]&m[582])|(~m[389]&~m[579]&m[580]&~m[581]&m[582])|(m[389]&m[579]&m[580]&~m[581]&m[582])|(~m[389]&m[579]&m[580]&m[581]&m[582]))&UnbiasedRNG[10])|((m[389]&~m[579]&~m[580]&m[581]&~m[582])|(~m[389]&~m[579]&~m[580]&~m[581]&m[582])|(m[389]&~m[579]&~m[580]&~m[581]&m[582])|(m[389]&m[579]&~m[580]&~m[581]&m[582])|(m[389]&~m[579]&m[580]&~m[581]&m[582])|(~m[389]&~m[579]&~m[580]&m[581]&m[582])|(m[389]&~m[579]&~m[580]&m[581]&m[582])|(~m[389]&m[579]&~m[580]&m[581]&m[582])|(m[389]&m[579]&~m[580]&m[581]&m[582])|(~m[389]&~m[579]&m[580]&m[581]&m[582])|(m[389]&~m[579]&m[580]&m[581]&m[582])|(m[389]&m[579]&m[580]&m[581]&m[582]));
    m[583] = (((m[581]&~m[584]&~m[585]&~m[586]&~m[587])|(~m[581]&~m[584]&~m[585]&m[586]&~m[587])|(m[581]&m[584]&~m[585]&m[586]&~m[587])|(m[581]&~m[584]&m[585]&m[586]&~m[587])|(~m[581]&m[584]&~m[585]&~m[586]&m[587])|(~m[581]&~m[584]&m[585]&~m[586]&m[587])|(m[581]&m[584]&m[585]&~m[586]&m[587])|(~m[581]&m[584]&m[585]&m[586]&m[587]))&UnbiasedRNG[11])|((m[581]&~m[584]&~m[585]&m[586]&~m[587])|(~m[581]&~m[584]&~m[585]&~m[586]&m[587])|(m[581]&~m[584]&~m[585]&~m[586]&m[587])|(m[581]&m[584]&~m[585]&~m[586]&m[587])|(m[581]&~m[584]&m[585]&~m[586]&m[587])|(~m[581]&~m[584]&~m[585]&m[586]&m[587])|(m[581]&~m[584]&~m[585]&m[586]&m[587])|(~m[581]&m[584]&~m[585]&m[586]&m[587])|(m[581]&m[584]&~m[585]&m[586]&m[587])|(~m[581]&~m[584]&m[585]&m[586]&m[587])|(m[581]&~m[584]&m[585]&m[586]&m[587])|(m[581]&m[584]&m[585]&m[586]&m[587]));
    m[588] = (((m[586]&~m[589]&~m[590]&~m[591]&~m[592])|(~m[586]&~m[589]&~m[590]&m[591]&~m[592])|(m[586]&m[589]&~m[590]&m[591]&~m[592])|(m[586]&~m[589]&m[590]&m[591]&~m[592])|(~m[586]&m[589]&~m[590]&~m[591]&m[592])|(~m[586]&~m[589]&m[590]&~m[591]&m[592])|(m[586]&m[589]&m[590]&~m[591]&m[592])|(~m[586]&m[589]&m[590]&m[591]&m[592]))&UnbiasedRNG[12])|((m[586]&~m[589]&~m[590]&m[591]&~m[592])|(~m[586]&~m[589]&~m[590]&~m[591]&m[592])|(m[586]&~m[589]&~m[590]&~m[591]&m[592])|(m[586]&m[589]&~m[590]&~m[591]&m[592])|(m[586]&~m[589]&m[590]&~m[591]&m[592])|(~m[586]&~m[589]&~m[590]&m[591]&m[592])|(m[586]&~m[589]&~m[590]&m[591]&m[592])|(~m[586]&m[589]&~m[590]&m[591]&m[592])|(m[586]&m[589]&~m[590]&m[591]&m[592])|(~m[586]&~m[589]&m[590]&m[591]&m[592])|(m[586]&~m[589]&m[590]&m[591]&m[592])|(m[586]&m[589]&m[590]&m[591]&m[592]));
    m[593] = (((m[591]&~m[594]&~m[595]&~m[596]&~m[597])|(~m[591]&~m[594]&~m[595]&m[596]&~m[597])|(m[591]&m[594]&~m[595]&m[596]&~m[597])|(m[591]&~m[594]&m[595]&m[596]&~m[597])|(~m[591]&m[594]&~m[595]&~m[596]&m[597])|(~m[591]&~m[594]&m[595]&~m[596]&m[597])|(m[591]&m[594]&m[595]&~m[596]&m[597])|(~m[591]&m[594]&m[595]&m[596]&m[597]))&UnbiasedRNG[13])|((m[591]&~m[594]&~m[595]&m[596]&~m[597])|(~m[591]&~m[594]&~m[595]&~m[596]&m[597])|(m[591]&~m[594]&~m[595]&~m[596]&m[597])|(m[591]&m[594]&~m[595]&~m[596]&m[597])|(m[591]&~m[594]&m[595]&~m[596]&m[597])|(~m[591]&~m[594]&~m[595]&m[596]&m[597])|(m[591]&~m[594]&~m[595]&m[596]&m[597])|(~m[591]&m[594]&~m[595]&m[596]&m[597])|(m[591]&m[594]&~m[595]&m[596]&m[597])|(~m[591]&~m[594]&m[595]&m[596]&m[597])|(m[591]&~m[594]&m[595]&m[596]&m[597])|(m[591]&m[594]&m[595]&m[596]&m[597]));
    m[598] = (((m[596]&~m[599]&~m[600]&~m[601]&~m[602])|(~m[596]&~m[599]&~m[600]&m[601]&~m[602])|(m[596]&m[599]&~m[600]&m[601]&~m[602])|(m[596]&~m[599]&m[600]&m[601]&~m[602])|(~m[596]&m[599]&~m[600]&~m[601]&m[602])|(~m[596]&~m[599]&m[600]&~m[601]&m[602])|(m[596]&m[599]&m[600]&~m[601]&m[602])|(~m[596]&m[599]&m[600]&m[601]&m[602]))&UnbiasedRNG[14])|((m[596]&~m[599]&~m[600]&m[601]&~m[602])|(~m[596]&~m[599]&~m[600]&~m[601]&m[602])|(m[596]&~m[599]&~m[600]&~m[601]&m[602])|(m[596]&m[599]&~m[600]&~m[601]&m[602])|(m[596]&~m[599]&m[600]&~m[601]&m[602])|(~m[596]&~m[599]&~m[600]&m[601]&m[602])|(m[596]&~m[599]&~m[600]&m[601]&m[602])|(~m[596]&m[599]&~m[600]&m[601]&m[602])|(m[596]&m[599]&~m[600]&m[601]&m[602])|(~m[596]&~m[599]&m[600]&m[601]&m[602])|(m[596]&~m[599]&m[600]&m[601]&m[602])|(m[596]&m[599]&m[600]&m[601]&m[602]));
    m[603] = (((m[390]&~m[604]&~m[605]&~m[606]&~m[607])|(~m[390]&~m[604]&~m[605]&m[606]&~m[607])|(m[390]&m[604]&~m[605]&m[606]&~m[607])|(m[390]&~m[604]&m[605]&m[606]&~m[607])|(~m[390]&m[604]&~m[605]&~m[606]&m[607])|(~m[390]&~m[604]&m[605]&~m[606]&m[607])|(m[390]&m[604]&m[605]&~m[606]&m[607])|(~m[390]&m[604]&m[605]&m[606]&m[607]))&UnbiasedRNG[15])|((m[390]&~m[604]&~m[605]&m[606]&~m[607])|(~m[390]&~m[604]&~m[605]&~m[606]&m[607])|(m[390]&~m[604]&~m[605]&~m[606]&m[607])|(m[390]&m[604]&~m[605]&~m[606]&m[607])|(m[390]&~m[604]&m[605]&~m[606]&m[607])|(~m[390]&~m[604]&~m[605]&m[606]&m[607])|(m[390]&~m[604]&~m[605]&m[606]&m[607])|(~m[390]&m[604]&~m[605]&m[606]&m[607])|(m[390]&m[604]&~m[605]&m[606]&m[607])|(~m[390]&~m[604]&m[605]&m[606]&m[607])|(m[390]&~m[604]&m[605]&m[606]&m[607])|(m[390]&m[604]&m[605]&m[606]&m[607]));
    m[608] = (((m[606]&~m[609]&~m[610]&~m[611]&~m[612])|(~m[606]&~m[609]&~m[610]&m[611]&~m[612])|(m[606]&m[609]&~m[610]&m[611]&~m[612])|(m[606]&~m[609]&m[610]&m[611]&~m[612])|(~m[606]&m[609]&~m[610]&~m[611]&m[612])|(~m[606]&~m[609]&m[610]&~m[611]&m[612])|(m[606]&m[609]&m[610]&~m[611]&m[612])|(~m[606]&m[609]&m[610]&m[611]&m[612]))&UnbiasedRNG[16])|((m[606]&~m[609]&~m[610]&m[611]&~m[612])|(~m[606]&~m[609]&~m[610]&~m[611]&m[612])|(m[606]&~m[609]&~m[610]&~m[611]&m[612])|(m[606]&m[609]&~m[610]&~m[611]&m[612])|(m[606]&~m[609]&m[610]&~m[611]&m[612])|(~m[606]&~m[609]&~m[610]&m[611]&m[612])|(m[606]&~m[609]&~m[610]&m[611]&m[612])|(~m[606]&m[609]&~m[610]&m[611]&m[612])|(m[606]&m[609]&~m[610]&m[611]&m[612])|(~m[606]&~m[609]&m[610]&m[611]&m[612])|(m[606]&~m[609]&m[610]&m[611]&m[612])|(m[606]&m[609]&m[610]&m[611]&m[612]));
    m[613] = (((m[611]&~m[614]&~m[615]&~m[616]&~m[617])|(~m[611]&~m[614]&~m[615]&m[616]&~m[617])|(m[611]&m[614]&~m[615]&m[616]&~m[617])|(m[611]&~m[614]&m[615]&m[616]&~m[617])|(~m[611]&m[614]&~m[615]&~m[616]&m[617])|(~m[611]&~m[614]&m[615]&~m[616]&m[617])|(m[611]&m[614]&m[615]&~m[616]&m[617])|(~m[611]&m[614]&m[615]&m[616]&m[617]))&UnbiasedRNG[17])|((m[611]&~m[614]&~m[615]&m[616]&~m[617])|(~m[611]&~m[614]&~m[615]&~m[616]&m[617])|(m[611]&~m[614]&~m[615]&~m[616]&m[617])|(m[611]&m[614]&~m[615]&~m[616]&m[617])|(m[611]&~m[614]&m[615]&~m[616]&m[617])|(~m[611]&~m[614]&~m[615]&m[616]&m[617])|(m[611]&~m[614]&~m[615]&m[616]&m[617])|(~m[611]&m[614]&~m[615]&m[616]&m[617])|(m[611]&m[614]&~m[615]&m[616]&m[617])|(~m[611]&~m[614]&m[615]&m[616]&m[617])|(m[611]&~m[614]&m[615]&m[616]&m[617])|(m[611]&m[614]&m[615]&m[616]&m[617]));
    m[618] = (((m[616]&~m[619]&~m[620]&~m[621]&~m[622])|(~m[616]&~m[619]&~m[620]&m[621]&~m[622])|(m[616]&m[619]&~m[620]&m[621]&~m[622])|(m[616]&~m[619]&m[620]&m[621]&~m[622])|(~m[616]&m[619]&~m[620]&~m[621]&m[622])|(~m[616]&~m[619]&m[620]&~m[621]&m[622])|(m[616]&m[619]&m[620]&~m[621]&m[622])|(~m[616]&m[619]&m[620]&m[621]&m[622]))&UnbiasedRNG[18])|((m[616]&~m[619]&~m[620]&m[621]&~m[622])|(~m[616]&~m[619]&~m[620]&~m[621]&m[622])|(m[616]&~m[619]&~m[620]&~m[621]&m[622])|(m[616]&m[619]&~m[620]&~m[621]&m[622])|(m[616]&~m[619]&m[620]&~m[621]&m[622])|(~m[616]&~m[619]&~m[620]&m[621]&m[622])|(m[616]&~m[619]&~m[620]&m[621]&m[622])|(~m[616]&m[619]&~m[620]&m[621]&m[622])|(m[616]&m[619]&~m[620]&m[621]&m[622])|(~m[616]&~m[619]&m[620]&m[621]&m[622])|(m[616]&~m[619]&m[620]&m[621]&m[622])|(m[616]&m[619]&m[620]&m[621]&m[622]));
    m[623] = (((m[621]&~m[624]&~m[625]&~m[626]&~m[627])|(~m[621]&~m[624]&~m[625]&m[626]&~m[627])|(m[621]&m[624]&~m[625]&m[626]&~m[627])|(m[621]&~m[624]&m[625]&m[626]&~m[627])|(~m[621]&m[624]&~m[625]&~m[626]&m[627])|(~m[621]&~m[624]&m[625]&~m[626]&m[627])|(m[621]&m[624]&m[625]&~m[626]&m[627])|(~m[621]&m[624]&m[625]&m[626]&m[627]))&UnbiasedRNG[19])|((m[621]&~m[624]&~m[625]&m[626]&~m[627])|(~m[621]&~m[624]&~m[625]&~m[626]&m[627])|(m[621]&~m[624]&~m[625]&~m[626]&m[627])|(m[621]&m[624]&~m[625]&~m[626]&m[627])|(m[621]&~m[624]&m[625]&~m[626]&m[627])|(~m[621]&~m[624]&~m[625]&m[626]&m[627])|(m[621]&~m[624]&~m[625]&m[626]&m[627])|(~m[621]&m[624]&~m[625]&m[626]&m[627])|(m[621]&m[624]&~m[625]&m[626]&m[627])|(~m[621]&~m[624]&m[625]&m[626]&m[627])|(m[621]&~m[624]&m[625]&m[626]&m[627])|(m[621]&m[624]&m[625]&m[626]&m[627]));
    m[628] = (((m[626]&~m[629]&~m[630]&~m[631]&~m[632])|(~m[626]&~m[629]&~m[630]&m[631]&~m[632])|(m[626]&m[629]&~m[630]&m[631]&~m[632])|(m[626]&~m[629]&m[630]&m[631]&~m[632])|(~m[626]&m[629]&~m[630]&~m[631]&m[632])|(~m[626]&~m[629]&m[630]&~m[631]&m[632])|(m[626]&m[629]&m[630]&~m[631]&m[632])|(~m[626]&m[629]&m[630]&m[631]&m[632]))&UnbiasedRNG[20])|((m[626]&~m[629]&~m[630]&m[631]&~m[632])|(~m[626]&~m[629]&~m[630]&~m[631]&m[632])|(m[626]&~m[629]&~m[630]&~m[631]&m[632])|(m[626]&m[629]&~m[630]&~m[631]&m[632])|(m[626]&~m[629]&m[630]&~m[631]&m[632])|(~m[626]&~m[629]&~m[630]&m[631]&m[632])|(m[626]&~m[629]&~m[630]&m[631]&m[632])|(~m[626]&m[629]&~m[630]&m[631]&m[632])|(m[626]&m[629]&~m[630]&m[631]&m[632])|(~m[626]&~m[629]&m[630]&m[631]&m[632])|(m[626]&~m[629]&m[630]&m[631]&m[632])|(m[626]&m[629]&m[630]&m[631]&m[632]));
    m[633] = (((m[391]&~m[634]&~m[635]&~m[636]&~m[637])|(~m[391]&~m[634]&~m[635]&m[636]&~m[637])|(m[391]&m[634]&~m[635]&m[636]&~m[637])|(m[391]&~m[634]&m[635]&m[636]&~m[637])|(~m[391]&m[634]&~m[635]&~m[636]&m[637])|(~m[391]&~m[634]&m[635]&~m[636]&m[637])|(m[391]&m[634]&m[635]&~m[636]&m[637])|(~m[391]&m[634]&m[635]&m[636]&m[637]))&UnbiasedRNG[21])|((m[391]&~m[634]&~m[635]&m[636]&~m[637])|(~m[391]&~m[634]&~m[635]&~m[636]&m[637])|(m[391]&~m[634]&~m[635]&~m[636]&m[637])|(m[391]&m[634]&~m[635]&~m[636]&m[637])|(m[391]&~m[634]&m[635]&~m[636]&m[637])|(~m[391]&~m[634]&~m[635]&m[636]&m[637])|(m[391]&~m[634]&~m[635]&m[636]&m[637])|(~m[391]&m[634]&~m[635]&m[636]&m[637])|(m[391]&m[634]&~m[635]&m[636]&m[637])|(~m[391]&~m[634]&m[635]&m[636]&m[637])|(m[391]&~m[634]&m[635]&m[636]&m[637])|(m[391]&m[634]&m[635]&m[636]&m[637]));
    m[638] = (((m[636]&~m[639]&~m[640]&~m[641]&~m[642])|(~m[636]&~m[639]&~m[640]&m[641]&~m[642])|(m[636]&m[639]&~m[640]&m[641]&~m[642])|(m[636]&~m[639]&m[640]&m[641]&~m[642])|(~m[636]&m[639]&~m[640]&~m[641]&m[642])|(~m[636]&~m[639]&m[640]&~m[641]&m[642])|(m[636]&m[639]&m[640]&~m[641]&m[642])|(~m[636]&m[639]&m[640]&m[641]&m[642]))&UnbiasedRNG[22])|((m[636]&~m[639]&~m[640]&m[641]&~m[642])|(~m[636]&~m[639]&~m[640]&~m[641]&m[642])|(m[636]&~m[639]&~m[640]&~m[641]&m[642])|(m[636]&m[639]&~m[640]&~m[641]&m[642])|(m[636]&~m[639]&m[640]&~m[641]&m[642])|(~m[636]&~m[639]&~m[640]&m[641]&m[642])|(m[636]&~m[639]&~m[640]&m[641]&m[642])|(~m[636]&m[639]&~m[640]&m[641]&m[642])|(m[636]&m[639]&~m[640]&m[641]&m[642])|(~m[636]&~m[639]&m[640]&m[641]&m[642])|(m[636]&~m[639]&m[640]&m[641]&m[642])|(m[636]&m[639]&m[640]&m[641]&m[642]));
    m[643] = (((m[641]&~m[644]&~m[645]&~m[646]&~m[647])|(~m[641]&~m[644]&~m[645]&m[646]&~m[647])|(m[641]&m[644]&~m[645]&m[646]&~m[647])|(m[641]&~m[644]&m[645]&m[646]&~m[647])|(~m[641]&m[644]&~m[645]&~m[646]&m[647])|(~m[641]&~m[644]&m[645]&~m[646]&m[647])|(m[641]&m[644]&m[645]&~m[646]&m[647])|(~m[641]&m[644]&m[645]&m[646]&m[647]))&UnbiasedRNG[23])|((m[641]&~m[644]&~m[645]&m[646]&~m[647])|(~m[641]&~m[644]&~m[645]&~m[646]&m[647])|(m[641]&~m[644]&~m[645]&~m[646]&m[647])|(m[641]&m[644]&~m[645]&~m[646]&m[647])|(m[641]&~m[644]&m[645]&~m[646]&m[647])|(~m[641]&~m[644]&~m[645]&m[646]&m[647])|(m[641]&~m[644]&~m[645]&m[646]&m[647])|(~m[641]&m[644]&~m[645]&m[646]&m[647])|(m[641]&m[644]&~m[645]&m[646]&m[647])|(~m[641]&~m[644]&m[645]&m[646]&m[647])|(m[641]&~m[644]&m[645]&m[646]&m[647])|(m[641]&m[644]&m[645]&m[646]&m[647]));
    m[648] = (((m[646]&~m[649]&~m[650]&~m[651]&~m[652])|(~m[646]&~m[649]&~m[650]&m[651]&~m[652])|(m[646]&m[649]&~m[650]&m[651]&~m[652])|(m[646]&~m[649]&m[650]&m[651]&~m[652])|(~m[646]&m[649]&~m[650]&~m[651]&m[652])|(~m[646]&~m[649]&m[650]&~m[651]&m[652])|(m[646]&m[649]&m[650]&~m[651]&m[652])|(~m[646]&m[649]&m[650]&m[651]&m[652]))&UnbiasedRNG[24])|((m[646]&~m[649]&~m[650]&m[651]&~m[652])|(~m[646]&~m[649]&~m[650]&~m[651]&m[652])|(m[646]&~m[649]&~m[650]&~m[651]&m[652])|(m[646]&m[649]&~m[650]&~m[651]&m[652])|(m[646]&~m[649]&m[650]&~m[651]&m[652])|(~m[646]&~m[649]&~m[650]&m[651]&m[652])|(m[646]&~m[649]&~m[650]&m[651]&m[652])|(~m[646]&m[649]&~m[650]&m[651]&m[652])|(m[646]&m[649]&~m[650]&m[651]&m[652])|(~m[646]&~m[649]&m[650]&m[651]&m[652])|(m[646]&~m[649]&m[650]&m[651]&m[652])|(m[646]&m[649]&m[650]&m[651]&m[652]));
    m[653] = (((m[651]&~m[654]&~m[655]&~m[656]&~m[657])|(~m[651]&~m[654]&~m[655]&m[656]&~m[657])|(m[651]&m[654]&~m[655]&m[656]&~m[657])|(m[651]&~m[654]&m[655]&m[656]&~m[657])|(~m[651]&m[654]&~m[655]&~m[656]&m[657])|(~m[651]&~m[654]&m[655]&~m[656]&m[657])|(m[651]&m[654]&m[655]&~m[656]&m[657])|(~m[651]&m[654]&m[655]&m[656]&m[657]))&UnbiasedRNG[25])|((m[651]&~m[654]&~m[655]&m[656]&~m[657])|(~m[651]&~m[654]&~m[655]&~m[656]&m[657])|(m[651]&~m[654]&~m[655]&~m[656]&m[657])|(m[651]&m[654]&~m[655]&~m[656]&m[657])|(m[651]&~m[654]&m[655]&~m[656]&m[657])|(~m[651]&~m[654]&~m[655]&m[656]&m[657])|(m[651]&~m[654]&~m[655]&m[656]&m[657])|(~m[651]&m[654]&~m[655]&m[656]&m[657])|(m[651]&m[654]&~m[655]&m[656]&m[657])|(~m[651]&~m[654]&m[655]&m[656]&m[657])|(m[651]&~m[654]&m[655]&m[656]&m[657])|(m[651]&m[654]&m[655]&m[656]&m[657]));
    m[658] = (((m[656]&~m[659]&~m[660]&~m[661]&~m[662])|(~m[656]&~m[659]&~m[660]&m[661]&~m[662])|(m[656]&m[659]&~m[660]&m[661]&~m[662])|(m[656]&~m[659]&m[660]&m[661]&~m[662])|(~m[656]&m[659]&~m[660]&~m[661]&m[662])|(~m[656]&~m[659]&m[660]&~m[661]&m[662])|(m[656]&m[659]&m[660]&~m[661]&m[662])|(~m[656]&m[659]&m[660]&m[661]&m[662]))&UnbiasedRNG[26])|((m[656]&~m[659]&~m[660]&m[661]&~m[662])|(~m[656]&~m[659]&~m[660]&~m[661]&m[662])|(m[656]&~m[659]&~m[660]&~m[661]&m[662])|(m[656]&m[659]&~m[660]&~m[661]&m[662])|(m[656]&~m[659]&m[660]&~m[661]&m[662])|(~m[656]&~m[659]&~m[660]&m[661]&m[662])|(m[656]&~m[659]&~m[660]&m[661]&m[662])|(~m[656]&m[659]&~m[660]&m[661]&m[662])|(m[656]&m[659]&~m[660]&m[661]&m[662])|(~m[656]&~m[659]&m[660]&m[661]&m[662])|(m[656]&~m[659]&m[660]&m[661]&m[662])|(m[656]&m[659]&m[660]&m[661]&m[662]));
    m[663] = (((m[661]&~m[664]&~m[665]&~m[666]&~m[667])|(~m[661]&~m[664]&~m[665]&m[666]&~m[667])|(m[661]&m[664]&~m[665]&m[666]&~m[667])|(m[661]&~m[664]&m[665]&m[666]&~m[667])|(~m[661]&m[664]&~m[665]&~m[666]&m[667])|(~m[661]&~m[664]&m[665]&~m[666]&m[667])|(m[661]&m[664]&m[665]&~m[666]&m[667])|(~m[661]&m[664]&m[665]&m[666]&m[667]))&UnbiasedRNG[27])|((m[661]&~m[664]&~m[665]&m[666]&~m[667])|(~m[661]&~m[664]&~m[665]&~m[666]&m[667])|(m[661]&~m[664]&~m[665]&~m[666]&m[667])|(m[661]&m[664]&~m[665]&~m[666]&m[667])|(m[661]&~m[664]&m[665]&~m[666]&m[667])|(~m[661]&~m[664]&~m[665]&m[666]&m[667])|(m[661]&~m[664]&~m[665]&m[666]&m[667])|(~m[661]&m[664]&~m[665]&m[666]&m[667])|(m[661]&m[664]&~m[665]&m[666]&m[667])|(~m[661]&~m[664]&m[665]&m[666]&m[667])|(m[661]&~m[664]&m[665]&m[666]&m[667])|(m[661]&m[664]&m[665]&m[666]&m[667]));
    m[668] = (((m[392]&~m[669]&~m[670]&~m[671]&~m[672])|(~m[392]&~m[669]&~m[670]&m[671]&~m[672])|(m[392]&m[669]&~m[670]&m[671]&~m[672])|(m[392]&~m[669]&m[670]&m[671]&~m[672])|(~m[392]&m[669]&~m[670]&~m[671]&m[672])|(~m[392]&~m[669]&m[670]&~m[671]&m[672])|(m[392]&m[669]&m[670]&~m[671]&m[672])|(~m[392]&m[669]&m[670]&m[671]&m[672]))&UnbiasedRNG[28])|((m[392]&~m[669]&~m[670]&m[671]&~m[672])|(~m[392]&~m[669]&~m[670]&~m[671]&m[672])|(m[392]&~m[669]&~m[670]&~m[671]&m[672])|(m[392]&m[669]&~m[670]&~m[671]&m[672])|(m[392]&~m[669]&m[670]&~m[671]&m[672])|(~m[392]&~m[669]&~m[670]&m[671]&m[672])|(m[392]&~m[669]&~m[670]&m[671]&m[672])|(~m[392]&m[669]&~m[670]&m[671]&m[672])|(m[392]&m[669]&~m[670]&m[671]&m[672])|(~m[392]&~m[669]&m[670]&m[671]&m[672])|(m[392]&~m[669]&m[670]&m[671]&m[672])|(m[392]&m[669]&m[670]&m[671]&m[672]));
    m[673] = (((m[671]&~m[674]&~m[675]&~m[676]&~m[677])|(~m[671]&~m[674]&~m[675]&m[676]&~m[677])|(m[671]&m[674]&~m[675]&m[676]&~m[677])|(m[671]&~m[674]&m[675]&m[676]&~m[677])|(~m[671]&m[674]&~m[675]&~m[676]&m[677])|(~m[671]&~m[674]&m[675]&~m[676]&m[677])|(m[671]&m[674]&m[675]&~m[676]&m[677])|(~m[671]&m[674]&m[675]&m[676]&m[677]))&UnbiasedRNG[29])|((m[671]&~m[674]&~m[675]&m[676]&~m[677])|(~m[671]&~m[674]&~m[675]&~m[676]&m[677])|(m[671]&~m[674]&~m[675]&~m[676]&m[677])|(m[671]&m[674]&~m[675]&~m[676]&m[677])|(m[671]&~m[674]&m[675]&~m[676]&m[677])|(~m[671]&~m[674]&~m[675]&m[676]&m[677])|(m[671]&~m[674]&~m[675]&m[676]&m[677])|(~m[671]&m[674]&~m[675]&m[676]&m[677])|(m[671]&m[674]&~m[675]&m[676]&m[677])|(~m[671]&~m[674]&m[675]&m[676]&m[677])|(m[671]&~m[674]&m[675]&m[676]&m[677])|(m[671]&m[674]&m[675]&m[676]&m[677]));
    m[678] = (((m[676]&~m[679]&~m[680]&~m[681]&~m[682])|(~m[676]&~m[679]&~m[680]&m[681]&~m[682])|(m[676]&m[679]&~m[680]&m[681]&~m[682])|(m[676]&~m[679]&m[680]&m[681]&~m[682])|(~m[676]&m[679]&~m[680]&~m[681]&m[682])|(~m[676]&~m[679]&m[680]&~m[681]&m[682])|(m[676]&m[679]&m[680]&~m[681]&m[682])|(~m[676]&m[679]&m[680]&m[681]&m[682]))&UnbiasedRNG[30])|((m[676]&~m[679]&~m[680]&m[681]&~m[682])|(~m[676]&~m[679]&~m[680]&~m[681]&m[682])|(m[676]&~m[679]&~m[680]&~m[681]&m[682])|(m[676]&m[679]&~m[680]&~m[681]&m[682])|(m[676]&~m[679]&m[680]&~m[681]&m[682])|(~m[676]&~m[679]&~m[680]&m[681]&m[682])|(m[676]&~m[679]&~m[680]&m[681]&m[682])|(~m[676]&m[679]&~m[680]&m[681]&m[682])|(m[676]&m[679]&~m[680]&m[681]&m[682])|(~m[676]&~m[679]&m[680]&m[681]&m[682])|(m[676]&~m[679]&m[680]&m[681]&m[682])|(m[676]&m[679]&m[680]&m[681]&m[682]));
    m[683] = (((m[681]&~m[684]&~m[685]&~m[686]&~m[687])|(~m[681]&~m[684]&~m[685]&m[686]&~m[687])|(m[681]&m[684]&~m[685]&m[686]&~m[687])|(m[681]&~m[684]&m[685]&m[686]&~m[687])|(~m[681]&m[684]&~m[685]&~m[686]&m[687])|(~m[681]&~m[684]&m[685]&~m[686]&m[687])|(m[681]&m[684]&m[685]&~m[686]&m[687])|(~m[681]&m[684]&m[685]&m[686]&m[687]))&UnbiasedRNG[31])|((m[681]&~m[684]&~m[685]&m[686]&~m[687])|(~m[681]&~m[684]&~m[685]&~m[686]&m[687])|(m[681]&~m[684]&~m[685]&~m[686]&m[687])|(m[681]&m[684]&~m[685]&~m[686]&m[687])|(m[681]&~m[684]&m[685]&~m[686]&m[687])|(~m[681]&~m[684]&~m[685]&m[686]&m[687])|(m[681]&~m[684]&~m[685]&m[686]&m[687])|(~m[681]&m[684]&~m[685]&m[686]&m[687])|(m[681]&m[684]&~m[685]&m[686]&m[687])|(~m[681]&~m[684]&m[685]&m[686]&m[687])|(m[681]&~m[684]&m[685]&m[686]&m[687])|(m[681]&m[684]&m[685]&m[686]&m[687]));
    m[688] = (((m[686]&~m[689]&~m[690]&~m[691]&~m[692])|(~m[686]&~m[689]&~m[690]&m[691]&~m[692])|(m[686]&m[689]&~m[690]&m[691]&~m[692])|(m[686]&~m[689]&m[690]&m[691]&~m[692])|(~m[686]&m[689]&~m[690]&~m[691]&m[692])|(~m[686]&~m[689]&m[690]&~m[691]&m[692])|(m[686]&m[689]&m[690]&~m[691]&m[692])|(~m[686]&m[689]&m[690]&m[691]&m[692]))&UnbiasedRNG[32])|((m[686]&~m[689]&~m[690]&m[691]&~m[692])|(~m[686]&~m[689]&~m[690]&~m[691]&m[692])|(m[686]&~m[689]&~m[690]&~m[691]&m[692])|(m[686]&m[689]&~m[690]&~m[691]&m[692])|(m[686]&~m[689]&m[690]&~m[691]&m[692])|(~m[686]&~m[689]&~m[690]&m[691]&m[692])|(m[686]&~m[689]&~m[690]&m[691]&m[692])|(~m[686]&m[689]&~m[690]&m[691]&m[692])|(m[686]&m[689]&~m[690]&m[691]&m[692])|(~m[686]&~m[689]&m[690]&m[691]&m[692])|(m[686]&~m[689]&m[690]&m[691]&m[692])|(m[686]&m[689]&m[690]&m[691]&m[692]));
    m[693] = (((m[691]&~m[694]&~m[695]&~m[696]&~m[697])|(~m[691]&~m[694]&~m[695]&m[696]&~m[697])|(m[691]&m[694]&~m[695]&m[696]&~m[697])|(m[691]&~m[694]&m[695]&m[696]&~m[697])|(~m[691]&m[694]&~m[695]&~m[696]&m[697])|(~m[691]&~m[694]&m[695]&~m[696]&m[697])|(m[691]&m[694]&m[695]&~m[696]&m[697])|(~m[691]&m[694]&m[695]&m[696]&m[697]))&UnbiasedRNG[33])|((m[691]&~m[694]&~m[695]&m[696]&~m[697])|(~m[691]&~m[694]&~m[695]&~m[696]&m[697])|(m[691]&~m[694]&~m[695]&~m[696]&m[697])|(m[691]&m[694]&~m[695]&~m[696]&m[697])|(m[691]&~m[694]&m[695]&~m[696]&m[697])|(~m[691]&~m[694]&~m[695]&m[696]&m[697])|(m[691]&~m[694]&~m[695]&m[696]&m[697])|(~m[691]&m[694]&~m[695]&m[696]&m[697])|(m[691]&m[694]&~m[695]&m[696]&m[697])|(~m[691]&~m[694]&m[695]&m[696]&m[697])|(m[691]&~m[694]&m[695]&m[696]&m[697])|(m[691]&m[694]&m[695]&m[696]&m[697]));
    m[698] = (((m[696]&~m[699]&~m[700]&~m[701]&~m[702])|(~m[696]&~m[699]&~m[700]&m[701]&~m[702])|(m[696]&m[699]&~m[700]&m[701]&~m[702])|(m[696]&~m[699]&m[700]&m[701]&~m[702])|(~m[696]&m[699]&~m[700]&~m[701]&m[702])|(~m[696]&~m[699]&m[700]&~m[701]&m[702])|(m[696]&m[699]&m[700]&~m[701]&m[702])|(~m[696]&m[699]&m[700]&m[701]&m[702]))&UnbiasedRNG[34])|((m[696]&~m[699]&~m[700]&m[701]&~m[702])|(~m[696]&~m[699]&~m[700]&~m[701]&m[702])|(m[696]&~m[699]&~m[700]&~m[701]&m[702])|(m[696]&m[699]&~m[700]&~m[701]&m[702])|(m[696]&~m[699]&m[700]&~m[701]&m[702])|(~m[696]&~m[699]&~m[700]&m[701]&m[702])|(m[696]&~m[699]&~m[700]&m[701]&m[702])|(~m[696]&m[699]&~m[700]&m[701]&m[702])|(m[696]&m[699]&~m[700]&m[701]&m[702])|(~m[696]&~m[699]&m[700]&m[701]&m[702])|(m[696]&~m[699]&m[700]&m[701]&m[702])|(m[696]&m[699]&m[700]&m[701]&m[702]));
    m[703] = (((m[701]&~m[704]&~m[705]&~m[706]&~m[707])|(~m[701]&~m[704]&~m[705]&m[706]&~m[707])|(m[701]&m[704]&~m[705]&m[706]&~m[707])|(m[701]&~m[704]&m[705]&m[706]&~m[707])|(~m[701]&m[704]&~m[705]&~m[706]&m[707])|(~m[701]&~m[704]&m[705]&~m[706]&m[707])|(m[701]&m[704]&m[705]&~m[706]&m[707])|(~m[701]&m[704]&m[705]&m[706]&m[707]))&UnbiasedRNG[35])|((m[701]&~m[704]&~m[705]&m[706]&~m[707])|(~m[701]&~m[704]&~m[705]&~m[706]&m[707])|(m[701]&~m[704]&~m[705]&~m[706]&m[707])|(m[701]&m[704]&~m[705]&~m[706]&m[707])|(m[701]&~m[704]&m[705]&~m[706]&m[707])|(~m[701]&~m[704]&~m[705]&m[706]&m[707])|(m[701]&~m[704]&~m[705]&m[706]&m[707])|(~m[701]&m[704]&~m[705]&m[706]&m[707])|(m[701]&m[704]&~m[705]&m[706]&m[707])|(~m[701]&~m[704]&m[705]&m[706]&m[707])|(m[701]&~m[704]&m[705]&m[706]&m[707])|(m[701]&m[704]&m[705]&m[706]&m[707]));
    m[708] = (((m[393]&~m[709]&~m[710]&~m[711]&~m[712])|(~m[393]&~m[709]&~m[710]&m[711]&~m[712])|(m[393]&m[709]&~m[710]&m[711]&~m[712])|(m[393]&~m[709]&m[710]&m[711]&~m[712])|(~m[393]&m[709]&~m[710]&~m[711]&m[712])|(~m[393]&~m[709]&m[710]&~m[711]&m[712])|(m[393]&m[709]&m[710]&~m[711]&m[712])|(~m[393]&m[709]&m[710]&m[711]&m[712]))&UnbiasedRNG[36])|((m[393]&~m[709]&~m[710]&m[711]&~m[712])|(~m[393]&~m[709]&~m[710]&~m[711]&m[712])|(m[393]&~m[709]&~m[710]&~m[711]&m[712])|(m[393]&m[709]&~m[710]&~m[711]&m[712])|(m[393]&~m[709]&m[710]&~m[711]&m[712])|(~m[393]&~m[709]&~m[710]&m[711]&m[712])|(m[393]&~m[709]&~m[710]&m[711]&m[712])|(~m[393]&m[709]&~m[710]&m[711]&m[712])|(m[393]&m[709]&~m[710]&m[711]&m[712])|(~m[393]&~m[709]&m[710]&m[711]&m[712])|(m[393]&~m[709]&m[710]&m[711]&m[712])|(m[393]&m[709]&m[710]&m[711]&m[712]));
    m[713] = (((m[711]&~m[714]&~m[715]&~m[716]&~m[717])|(~m[711]&~m[714]&~m[715]&m[716]&~m[717])|(m[711]&m[714]&~m[715]&m[716]&~m[717])|(m[711]&~m[714]&m[715]&m[716]&~m[717])|(~m[711]&m[714]&~m[715]&~m[716]&m[717])|(~m[711]&~m[714]&m[715]&~m[716]&m[717])|(m[711]&m[714]&m[715]&~m[716]&m[717])|(~m[711]&m[714]&m[715]&m[716]&m[717]))&UnbiasedRNG[37])|((m[711]&~m[714]&~m[715]&m[716]&~m[717])|(~m[711]&~m[714]&~m[715]&~m[716]&m[717])|(m[711]&~m[714]&~m[715]&~m[716]&m[717])|(m[711]&m[714]&~m[715]&~m[716]&m[717])|(m[711]&~m[714]&m[715]&~m[716]&m[717])|(~m[711]&~m[714]&~m[715]&m[716]&m[717])|(m[711]&~m[714]&~m[715]&m[716]&m[717])|(~m[711]&m[714]&~m[715]&m[716]&m[717])|(m[711]&m[714]&~m[715]&m[716]&m[717])|(~m[711]&~m[714]&m[715]&m[716]&m[717])|(m[711]&~m[714]&m[715]&m[716]&m[717])|(m[711]&m[714]&m[715]&m[716]&m[717]));
    m[718] = (((m[716]&~m[719]&~m[720]&~m[721]&~m[722])|(~m[716]&~m[719]&~m[720]&m[721]&~m[722])|(m[716]&m[719]&~m[720]&m[721]&~m[722])|(m[716]&~m[719]&m[720]&m[721]&~m[722])|(~m[716]&m[719]&~m[720]&~m[721]&m[722])|(~m[716]&~m[719]&m[720]&~m[721]&m[722])|(m[716]&m[719]&m[720]&~m[721]&m[722])|(~m[716]&m[719]&m[720]&m[721]&m[722]))&UnbiasedRNG[38])|((m[716]&~m[719]&~m[720]&m[721]&~m[722])|(~m[716]&~m[719]&~m[720]&~m[721]&m[722])|(m[716]&~m[719]&~m[720]&~m[721]&m[722])|(m[716]&m[719]&~m[720]&~m[721]&m[722])|(m[716]&~m[719]&m[720]&~m[721]&m[722])|(~m[716]&~m[719]&~m[720]&m[721]&m[722])|(m[716]&~m[719]&~m[720]&m[721]&m[722])|(~m[716]&m[719]&~m[720]&m[721]&m[722])|(m[716]&m[719]&~m[720]&m[721]&m[722])|(~m[716]&~m[719]&m[720]&m[721]&m[722])|(m[716]&~m[719]&m[720]&m[721]&m[722])|(m[716]&m[719]&m[720]&m[721]&m[722]));
    m[723] = (((m[721]&~m[724]&~m[725]&~m[726]&~m[727])|(~m[721]&~m[724]&~m[725]&m[726]&~m[727])|(m[721]&m[724]&~m[725]&m[726]&~m[727])|(m[721]&~m[724]&m[725]&m[726]&~m[727])|(~m[721]&m[724]&~m[725]&~m[726]&m[727])|(~m[721]&~m[724]&m[725]&~m[726]&m[727])|(m[721]&m[724]&m[725]&~m[726]&m[727])|(~m[721]&m[724]&m[725]&m[726]&m[727]))&UnbiasedRNG[39])|((m[721]&~m[724]&~m[725]&m[726]&~m[727])|(~m[721]&~m[724]&~m[725]&~m[726]&m[727])|(m[721]&~m[724]&~m[725]&~m[726]&m[727])|(m[721]&m[724]&~m[725]&~m[726]&m[727])|(m[721]&~m[724]&m[725]&~m[726]&m[727])|(~m[721]&~m[724]&~m[725]&m[726]&m[727])|(m[721]&~m[724]&~m[725]&m[726]&m[727])|(~m[721]&m[724]&~m[725]&m[726]&m[727])|(m[721]&m[724]&~m[725]&m[726]&m[727])|(~m[721]&~m[724]&m[725]&m[726]&m[727])|(m[721]&~m[724]&m[725]&m[726]&m[727])|(m[721]&m[724]&m[725]&m[726]&m[727]));
    m[728] = (((m[726]&~m[729]&~m[730]&~m[731]&~m[732])|(~m[726]&~m[729]&~m[730]&m[731]&~m[732])|(m[726]&m[729]&~m[730]&m[731]&~m[732])|(m[726]&~m[729]&m[730]&m[731]&~m[732])|(~m[726]&m[729]&~m[730]&~m[731]&m[732])|(~m[726]&~m[729]&m[730]&~m[731]&m[732])|(m[726]&m[729]&m[730]&~m[731]&m[732])|(~m[726]&m[729]&m[730]&m[731]&m[732]))&UnbiasedRNG[40])|((m[726]&~m[729]&~m[730]&m[731]&~m[732])|(~m[726]&~m[729]&~m[730]&~m[731]&m[732])|(m[726]&~m[729]&~m[730]&~m[731]&m[732])|(m[726]&m[729]&~m[730]&~m[731]&m[732])|(m[726]&~m[729]&m[730]&~m[731]&m[732])|(~m[726]&~m[729]&~m[730]&m[731]&m[732])|(m[726]&~m[729]&~m[730]&m[731]&m[732])|(~m[726]&m[729]&~m[730]&m[731]&m[732])|(m[726]&m[729]&~m[730]&m[731]&m[732])|(~m[726]&~m[729]&m[730]&m[731]&m[732])|(m[726]&~m[729]&m[730]&m[731]&m[732])|(m[726]&m[729]&m[730]&m[731]&m[732]));
    m[733] = (((m[731]&~m[734]&~m[735]&~m[736]&~m[737])|(~m[731]&~m[734]&~m[735]&m[736]&~m[737])|(m[731]&m[734]&~m[735]&m[736]&~m[737])|(m[731]&~m[734]&m[735]&m[736]&~m[737])|(~m[731]&m[734]&~m[735]&~m[736]&m[737])|(~m[731]&~m[734]&m[735]&~m[736]&m[737])|(m[731]&m[734]&m[735]&~m[736]&m[737])|(~m[731]&m[734]&m[735]&m[736]&m[737]))&UnbiasedRNG[41])|((m[731]&~m[734]&~m[735]&m[736]&~m[737])|(~m[731]&~m[734]&~m[735]&~m[736]&m[737])|(m[731]&~m[734]&~m[735]&~m[736]&m[737])|(m[731]&m[734]&~m[735]&~m[736]&m[737])|(m[731]&~m[734]&m[735]&~m[736]&m[737])|(~m[731]&~m[734]&~m[735]&m[736]&m[737])|(m[731]&~m[734]&~m[735]&m[736]&m[737])|(~m[731]&m[734]&~m[735]&m[736]&m[737])|(m[731]&m[734]&~m[735]&m[736]&m[737])|(~m[731]&~m[734]&m[735]&m[736]&m[737])|(m[731]&~m[734]&m[735]&m[736]&m[737])|(m[731]&m[734]&m[735]&m[736]&m[737]));
    m[738] = (((m[736]&~m[739]&~m[740]&~m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&m[741]&~m[742])|(m[736]&m[739]&~m[740]&m[741]&~m[742])|(m[736]&~m[739]&m[740]&m[741]&~m[742])|(~m[736]&m[739]&~m[740]&~m[741]&m[742])|(~m[736]&~m[739]&m[740]&~m[741]&m[742])|(m[736]&m[739]&m[740]&~m[741]&m[742])|(~m[736]&m[739]&m[740]&m[741]&m[742]))&UnbiasedRNG[42])|((m[736]&~m[739]&~m[740]&m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&m[740]&~m[741]&m[742])|(~m[736]&~m[739]&~m[740]&m[741]&m[742])|(m[736]&~m[739]&~m[740]&m[741]&m[742])|(~m[736]&m[739]&~m[740]&m[741]&m[742])|(m[736]&m[739]&~m[740]&m[741]&m[742])|(~m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&m[739]&m[740]&m[741]&m[742]));
    m[743] = (((m[741]&~m[744]&~m[745]&~m[746]&~m[747])|(~m[741]&~m[744]&~m[745]&m[746]&~m[747])|(m[741]&m[744]&~m[745]&m[746]&~m[747])|(m[741]&~m[744]&m[745]&m[746]&~m[747])|(~m[741]&m[744]&~m[745]&~m[746]&m[747])|(~m[741]&~m[744]&m[745]&~m[746]&m[747])|(m[741]&m[744]&m[745]&~m[746]&m[747])|(~m[741]&m[744]&m[745]&m[746]&m[747]))&UnbiasedRNG[43])|((m[741]&~m[744]&~m[745]&m[746]&~m[747])|(~m[741]&~m[744]&~m[745]&~m[746]&m[747])|(m[741]&~m[744]&~m[745]&~m[746]&m[747])|(m[741]&m[744]&~m[745]&~m[746]&m[747])|(m[741]&~m[744]&m[745]&~m[746]&m[747])|(~m[741]&~m[744]&~m[745]&m[746]&m[747])|(m[741]&~m[744]&~m[745]&m[746]&m[747])|(~m[741]&m[744]&~m[745]&m[746]&m[747])|(m[741]&m[744]&~m[745]&m[746]&m[747])|(~m[741]&~m[744]&m[745]&m[746]&m[747])|(m[741]&~m[744]&m[745]&m[746]&m[747])|(m[741]&m[744]&m[745]&m[746]&m[747]));
    m[748] = (((m[746]&~m[749]&~m[750]&~m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&m[751]&~m[752])|(m[746]&m[749]&~m[750]&m[751]&~m[752])|(m[746]&~m[749]&m[750]&m[751]&~m[752])|(~m[746]&m[749]&~m[750]&~m[751]&m[752])|(~m[746]&~m[749]&m[750]&~m[751]&m[752])|(m[746]&m[749]&m[750]&~m[751]&m[752])|(~m[746]&m[749]&m[750]&m[751]&m[752]))&UnbiasedRNG[44])|((m[746]&~m[749]&~m[750]&m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&m[750]&~m[751]&m[752])|(~m[746]&~m[749]&~m[750]&m[751]&m[752])|(m[746]&~m[749]&~m[750]&m[751]&m[752])|(~m[746]&m[749]&~m[750]&m[751]&m[752])|(m[746]&m[749]&~m[750]&m[751]&m[752])|(~m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&m[749]&m[750]&m[751]&m[752]));
    m[753] = (((m[394]&~m[754]&~m[755]&~m[756]&~m[757])|(~m[394]&~m[754]&~m[755]&m[756]&~m[757])|(m[394]&m[754]&~m[755]&m[756]&~m[757])|(m[394]&~m[754]&m[755]&m[756]&~m[757])|(~m[394]&m[754]&~m[755]&~m[756]&m[757])|(~m[394]&~m[754]&m[755]&~m[756]&m[757])|(m[394]&m[754]&m[755]&~m[756]&m[757])|(~m[394]&m[754]&m[755]&m[756]&m[757]))&UnbiasedRNG[45])|((m[394]&~m[754]&~m[755]&m[756]&~m[757])|(~m[394]&~m[754]&~m[755]&~m[756]&m[757])|(m[394]&~m[754]&~m[755]&~m[756]&m[757])|(m[394]&m[754]&~m[755]&~m[756]&m[757])|(m[394]&~m[754]&m[755]&~m[756]&m[757])|(~m[394]&~m[754]&~m[755]&m[756]&m[757])|(m[394]&~m[754]&~m[755]&m[756]&m[757])|(~m[394]&m[754]&~m[755]&m[756]&m[757])|(m[394]&m[754]&~m[755]&m[756]&m[757])|(~m[394]&~m[754]&m[755]&m[756]&m[757])|(m[394]&~m[754]&m[755]&m[756]&m[757])|(m[394]&m[754]&m[755]&m[756]&m[757]));
    m[758] = (((m[756]&~m[759]&~m[760]&~m[761]&~m[762])|(~m[756]&~m[759]&~m[760]&m[761]&~m[762])|(m[756]&m[759]&~m[760]&m[761]&~m[762])|(m[756]&~m[759]&m[760]&m[761]&~m[762])|(~m[756]&m[759]&~m[760]&~m[761]&m[762])|(~m[756]&~m[759]&m[760]&~m[761]&m[762])|(m[756]&m[759]&m[760]&~m[761]&m[762])|(~m[756]&m[759]&m[760]&m[761]&m[762]))&UnbiasedRNG[46])|((m[756]&~m[759]&~m[760]&m[761]&~m[762])|(~m[756]&~m[759]&~m[760]&~m[761]&m[762])|(m[756]&~m[759]&~m[760]&~m[761]&m[762])|(m[756]&m[759]&~m[760]&~m[761]&m[762])|(m[756]&~m[759]&m[760]&~m[761]&m[762])|(~m[756]&~m[759]&~m[760]&m[761]&m[762])|(m[756]&~m[759]&~m[760]&m[761]&m[762])|(~m[756]&m[759]&~m[760]&m[761]&m[762])|(m[756]&m[759]&~m[760]&m[761]&m[762])|(~m[756]&~m[759]&m[760]&m[761]&m[762])|(m[756]&~m[759]&m[760]&m[761]&m[762])|(m[756]&m[759]&m[760]&m[761]&m[762]));
    m[763] = (((m[761]&~m[764]&~m[765]&~m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&m[766]&~m[767])|(m[761]&m[764]&~m[765]&m[766]&~m[767])|(m[761]&~m[764]&m[765]&m[766]&~m[767])|(~m[761]&m[764]&~m[765]&~m[766]&m[767])|(~m[761]&~m[764]&m[765]&~m[766]&m[767])|(m[761]&m[764]&m[765]&~m[766]&m[767])|(~m[761]&m[764]&m[765]&m[766]&m[767]))&UnbiasedRNG[47])|((m[761]&~m[764]&~m[765]&m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&m[765]&~m[766]&m[767])|(~m[761]&~m[764]&~m[765]&m[766]&m[767])|(m[761]&~m[764]&~m[765]&m[766]&m[767])|(~m[761]&m[764]&~m[765]&m[766]&m[767])|(m[761]&m[764]&~m[765]&m[766]&m[767])|(~m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&m[764]&m[765]&m[766]&m[767]));
    m[768] = (((m[766]&~m[769]&~m[770]&~m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&m[771]&~m[772])|(m[766]&m[769]&~m[770]&m[771]&~m[772])|(m[766]&~m[769]&m[770]&m[771]&~m[772])|(~m[766]&m[769]&~m[770]&~m[771]&m[772])|(~m[766]&~m[769]&m[770]&~m[771]&m[772])|(m[766]&m[769]&m[770]&~m[771]&m[772])|(~m[766]&m[769]&m[770]&m[771]&m[772]))&UnbiasedRNG[48])|((m[766]&~m[769]&~m[770]&m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&m[770]&~m[771]&m[772])|(~m[766]&~m[769]&~m[770]&m[771]&m[772])|(m[766]&~m[769]&~m[770]&m[771]&m[772])|(~m[766]&m[769]&~m[770]&m[771]&m[772])|(m[766]&m[769]&~m[770]&m[771]&m[772])|(~m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&m[769]&m[770]&m[771]&m[772]));
    m[773] = (((m[771]&~m[774]&~m[775]&~m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&m[776]&~m[777])|(m[771]&m[774]&~m[775]&m[776]&~m[777])|(m[771]&~m[774]&m[775]&m[776]&~m[777])|(~m[771]&m[774]&~m[775]&~m[776]&m[777])|(~m[771]&~m[774]&m[775]&~m[776]&m[777])|(m[771]&m[774]&m[775]&~m[776]&m[777])|(~m[771]&m[774]&m[775]&m[776]&m[777]))&UnbiasedRNG[49])|((m[771]&~m[774]&~m[775]&m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&m[775]&~m[776]&m[777])|(~m[771]&~m[774]&~m[775]&m[776]&m[777])|(m[771]&~m[774]&~m[775]&m[776]&m[777])|(~m[771]&m[774]&~m[775]&m[776]&m[777])|(m[771]&m[774]&~m[775]&m[776]&m[777])|(~m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&m[774]&m[775]&m[776]&m[777]));
    m[778] = (((m[776]&~m[779]&~m[780]&~m[781]&~m[782])|(~m[776]&~m[779]&~m[780]&m[781]&~m[782])|(m[776]&m[779]&~m[780]&m[781]&~m[782])|(m[776]&~m[779]&m[780]&m[781]&~m[782])|(~m[776]&m[779]&~m[780]&~m[781]&m[782])|(~m[776]&~m[779]&m[780]&~m[781]&m[782])|(m[776]&m[779]&m[780]&~m[781]&m[782])|(~m[776]&m[779]&m[780]&m[781]&m[782]))&UnbiasedRNG[50])|((m[776]&~m[779]&~m[780]&m[781]&~m[782])|(~m[776]&~m[779]&~m[780]&~m[781]&m[782])|(m[776]&~m[779]&~m[780]&~m[781]&m[782])|(m[776]&m[779]&~m[780]&~m[781]&m[782])|(m[776]&~m[779]&m[780]&~m[781]&m[782])|(~m[776]&~m[779]&~m[780]&m[781]&m[782])|(m[776]&~m[779]&~m[780]&m[781]&m[782])|(~m[776]&m[779]&~m[780]&m[781]&m[782])|(m[776]&m[779]&~m[780]&m[781]&m[782])|(~m[776]&~m[779]&m[780]&m[781]&m[782])|(m[776]&~m[779]&m[780]&m[781]&m[782])|(m[776]&m[779]&m[780]&m[781]&m[782]));
    m[783] = (((m[781]&~m[784]&~m[785]&~m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&m[786]&~m[787])|(m[781]&m[784]&~m[785]&m[786]&~m[787])|(m[781]&~m[784]&m[785]&m[786]&~m[787])|(~m[781]&m[784]&~m[785]&~m[786]&m[787])|(~m[781]&~m[784]&m[785]&~m[786]&m[787])|(m[781]&m[784]&m[785]&~m[786]&m[787])|(~m[781]&m[784]&m[785]&m[786]&m[787]))&UnbiasedRNG[51])|((m[781]&~m[784]&~m[785]&m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&m[785]&~m[786]&m[787])|(~m[781]&~m[784]&~m[785]&m[786]&m[787])|(m[781]&~m[784]&~m[785]&m[786]&m[787])|(~m[781]&m[784]&~m[785]&m[786]&m[787])|(m[781]&m[784]&~m[785]&m[786]&m[787])|(~m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&m[784]&m[785]&m[786]&m[787]));
    m[788] = (((m[786]&~m[789]&~m[790]&~m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&m[791]&~m[792])|(m[786]&m[789]&~m[790]&m[791]&~m[792])|(m[786]&~m[789]&m[790]&m[791]&~m[792])|(~m[786]&m[789]&~m[790]&~m[791]&m[792])|(~m[786]&~m[789]&m[790]&~m[791]&m[792])|(m[786]&m[789]&m[790]&~m[791]&m[792])|(~m[786]&m[789]&m[790]&m[791]&m[792]))&UnbiasedRNG[52])|((m[786]&~m[789]&~m[790]&m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&m[790]&~m[791]&m[792])|(~m[786]&~m[789]&~m[790]&m[791]&m[792])|(m[786]&~m[789]&~m[790]&m[791]&m[792])|(~m[786]&m[789]&~m[790]&m[791]&m[792])|(m[786]&m[789]&~m[790]&m[791]&m[792])|(~m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&m[789]&m[790]&m[791]&m[792]));
    m[793] = (((m[791]&~m[794]&~m[795]&~m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&m[796]&~m[797])|(m[791]&m[794]&~m[795]&m[796]&~m[797])|(m[791]&~m[794]&m[795]&m[796]&~m[797])|(~m[791]&m[794]&~m[795]&~m[796]&m[797])|(~m[791]&~m[794]&m[795]&~m[796]&m[797])|(m[791]&m[794]&m[795]&~m[796]&m[797])|(~m[791]&m[794]&m[795]&m[796]&m[797]))&UnbiasedRNG[53])|((m[791]&~m[794]&~m[795]&m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&m[795]&~m[796]&m[797])|(~m[791]&~m[794]&~m[795]&m[796]&m[797])|(m[791]&~m[794]&~m[795]&m[796]&m[797])|(~m[791]&m[794]&~m[795]&m[796]&m[797])|(m[791]&m[794]&~m[795]&m[796]&m[797])|(~m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&m[794]&m[795]&m[796]&m[797]));
    m[798] = (((m[796]&~m[799]&~m[800]&~m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&m[801]&~m[802])|(m[796]&m[799]&~m[800]&m[801]&~m[802])|(m[796]&~m[799]&m[800]&m[801]&~m[802])|(~m[796]&m[799]&~m[800]&~m[801]&m[802])|(~m[796]&~m[799]&m[800]&~m[801]&m[802])|(m[796]&m[799]&m[800]&~m[801]&m[802])|(~m[796]&m[799]&m[800]&m[801]&m[802]))&UnbiasedRNG[54])|((m[796]&~m[799]&~m[800]&m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&m[800]&~m[801]&m[802])|(~m[796]&~m[799]&~m[800]&m[801]&m[802])|(m[796]&~m[799]&~m[800]&m[801]&m[802])|(~m[796]&m[799]&~m[800]&m[801]&m[802])|(m[796]&m[799]&~m[800]&m[801]&m[802])|(~m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&m[799]&m[800]&m[801]&m[802]));
    m[803] = (((m[395]&~m[804]&~m[805]&~m[806]&~m[807])|(~m[395]&~m[804]&~m[805]&m[806]&~m[807])|(m[395]&m[804]&~m[805]&m[806]&~m[807])|(m[395]&~m[804]&m[805]&m[806]&~m[807])|(~m[395]&m[804]&~m[805]&~m[806]&m[807])|(~m[395]&~m[804]&m[805]&~m[806]&m[807])|(m[395]&m[804]&m[805]&~m[806]&m[807])|(~m[395]&m[804]&m[805]&m[806]&m[807]))&UnbiasedRNG[55])|((m[395]&~m[804]&~m[805]&m[806]&~m[807])|(~m[395]&~m[804]&~m[805]&~m[806]&m[807])|(m[395]&~m[804]&~m[805]&~m[806]&m[807])|(m[395]&m[804]&~m[805]&~m[806]&m[807])|(m[395]&~m[804]&m[805]&~m[806]&m[807])|(~m[395]&~m[804]&~m[805]&m[806]&m[807])|(m[395]&~m[804]&~m[805]&m[806]&m[807])|(~m[395]&m[804]&~m[805]&m[806]&m[807])|(m[395]&m[804]&~m[805]&m[806]&m[807])|(~m[395]&~m[804]&m[805]&m[806]&m[807])|(m[395]&~m[804]&m[805]&m[806]&m[807])|(m[395]&m[804]&m[805]&m[806]&m[807]));
    m[808] = (((m[806]&~m[809]&~m[810]&~m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&m[811]&~m[812])|(m[806]&m[809]&~m[810]&m[811]&~m[812])|(m[806]&~m[809]&m[810]&m[811]&~m[812])|(~m[806]&m[809]&~m[810]&~m[811]&m[812])|(~m[806]&~m[809]&m[810]&~m[811]&m[812])|(m[806]&m[809]&m[810]&~m[811]&m[812])|(~m[806]&m[809]&m[810]&m[811]&m[812]))&UnbiasedRNG[56])|((m[806]&~m[809]&~m[810]&m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&m[810]&~m[811]&m[812])|(~m[806]&~m[809]&~m[810]&m[811]&m[812])|(m[806]&~m[809]&~m[810]&m[811]&m[812])|(~m[806]&m[809]&~m[810]&m[811]&m[812])|(m[806]&m[809]&~m[810]&m[811]&m[812])|(~m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&m[809]&m[810]&m[811]&m[812]));
    m[813] = (((m[811]&~m[814]&~m[815]&~m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&m[816]&~m[817])|(m[811]&m[814]&~m[815]&m[816]&~m[817])|(m[811]&~m[814]&m[815]&m[816]&~m[817])|(~m[811]&m[814]&~m[815]&~m[816]&m[817])|(~m[811]&~m[814]&m[815]&~m[816]&m[817])|(m[811]&m[814]&m[815]&~m[816]&m[817])|(~m[811]&m[814]&m[815]&m[816]&m[817]))&UnbiasedRNG[57])|((m[811]&~m[814]&~m[815]&m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&m[815]&~m[816]&m[817])|(~m[811]&~m[814]&~m[815]&m[816]&m[817])|(m[811]&~m[814]&~m[815]&m[816]&m[817])|(~m[811]&m[814]&~m[815]&m[816]&m[817])|(m[811]&m[814]&~m[815]&m[816]&m[817])|(~m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&m[814]&m[815]&m[816]&m[817]));
    m[818] = (((m[816]&~m[819]&~m[820]&~m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&m[821]&~m[822])|(m[816]&m[819]&~m[820]&m[821]&~m[822])|(m[816]&~m[819]&m[820]&m[821]&~m[822])|(~m[816]&m[819]&~m[820]&~m[821]&m[822])|(~m[816]&~m[819]&m[820]&~m[821]&m[822])|(m[816]&m[819]&m[820]&~m[821]&m[822])|(~m[816]&m[819]&m[820]&m[821]&m[822]))&UnbiasedRNG[58])|((m[816]&~m[819]&~m[820]&m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&m[820]&~m[821]&m[822])|(~m[816]&~m[819]&~m[820]&m[821]&m[822])|(m[816]&~m[819]&~m[820]&m[821]&m[822])|(~m[816]&m[819]&~m[820]&m[821]&m[822])|(m[816]&m[819]&~m[820]&m[821]&m[822])|(~m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&m[819]&m[820]&m[821]&m[822]));
    m[823] = (((m[821]&~m[824]&~m[825]&~m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&m[826]&~m[827])|(m[821]&m[824]&~m[825]&m[826]&~m[827])|(m[821]&~m[824]&m[825]&m[826]&~m[827])|(~m[821]&m[824]&~m[825]&~m[826]&m[827])|(~m[821]&~m[824]&m[825]&~m[826]&m[827])|(m[821]&m[824]&m[825]&~m[826]&m[827])|(~m[821]&m[824]&m[825]&m[826]&m[827]))&UnbiasedRNG[59])|((m[821]&~m[824]&~m[825]&m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&m[825]&~m[826]&m[827])|(~m[821]&~m[824]&~m[825]&m[826]&m[827])|(m[821]&~m[824]&~m[825]&m[826]&m[827])|(~m[821]&m[824]&~m[825]&m[826]&m[827])|(m[821]&m[824]&~m[825]&m[826]&m[827])|(~m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&m[824]&m[825]&m[826]&m[827]));
    m[828] = (((m[826]&~m[829]&~m[830]&~m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&m[831]&~m[832])|(m[826]&m[829]&~m[830]&m[831]&~m[832])|(m[826]&~m[829]&m[830]&m[831]&~m[832])|(~m[826]&m[829]&~m[830]&~m[831]&m[832])|(~m[826]&~m[829]&m[830]&~m[831]&m[832])|(m[826]&m[829]&m[830]&~m[831]&m[832])|(~m[826]&m[829]&m[830]&m[831]&m[832]))&UnbiasedRNG[60])|((m[826]&~m[829]&~m[830]&m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&m[830]&~m[831]&m[832])|(~m[826]&~m[829]&~m[830]&m[831]&m[832])|(m[826]&~m[829]&~m[830]&m[831]&m[832])|(~m[826]&m[829]&~m[830]&m[831]&m[832])|(m[826]&m[829]&~m[830]&m[831]&m[832])|(~m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&m[829]&m[830]&m[831]&m[832]));
    m[833] = (((m[831]&~m[834]&~m[835]&~m[836]&~m[837])|(~m[831]&~m[834]&~m[835]&m[836]&~m[837])|(m[831]&m[834]&~m[835]&m[836]&~m[837])|(m[831]&~m[834]&m[835]&m[836]&~m[837])|(~m[831]&m[834]&~m[835]&~m[836]&m[837])|(~m[831]&~m[834]&m[835]&~m[836]&m[837])|(m[831]&m[834]&m[835]&~m[836]&m[837])|(~m[831]&m[834]&m[835]&m[836]&m[837]))&UnbiasedRNG[61])|((m[831]&~m[834]&~m[835]&m[836]&~m[837])|(~m[831]&~m[834]&~m[835]&~m[836]&m[837])|(m[831]&~m[834]&~m[835]&~m[836]&m[837])|(m[831]&m[834]&~m[835]&~m[836]&m[837])|(m[831]&~m[834]&m[835]&~m[836]&m[837])|(~m[831]&~m[834]&~m[835]&m[836]&m[837])|(m[831]&~m[834]&~m[835]&m[836]&m[837])|(~m[831]&m[834]&~m[835]&m[836]&m[837])|(m[831]&m[834]&~m[835]&m[836]&m[837])|(~m[831]&~m[834]&m[835]&m[836]&m[837])|(m[831]&~m[834]&m[835]&m[836]&m[837])|(m[831]&m[834]&m[835]&m[836]&m[837]));
    m[838] = (((m[836]&~m[839]&~m[840]&~m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&m[841]&~m[842])|(m[836]&m[839]&~m[840]&m[841]&~m[842])|(m[836]&~m[839]&m[840]&m[841]&~m[842])|(~m[836]&m[839]&~m[840]&~m[841]&m[842])|(~m[836]&~m[839]&m[840]&~m[841]&m[842])|(m[836]&m[839]&m[840]&~m[841]&m[842])|(~m[836]&m[839]&m[840]&m[841]&m[842]))&UnbiasedRNG[62])|((m[836]&~m[839]&~m[840]&m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&m[840]&~m[841]&m[842])|(~m[836]&~m[839]&~m[840]&m[841]&m[842])|(m[836]&~m[839]&~m[840]&m[841]&m[842])|(~m[836]&m[839]&~m[840]&m[841]&m[842])|(m[836]&m[839]&~m[840]&m[841]&m[842])|(~m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&m[839]&m[840]&m[841]&m[842]));
    m[843] = (((m[841]&~m[844]&~m[845]&~m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&m[846]&~m[847])|(m[841]&m[844]&~m[845]&m[846]&~m[847])|(m[841]&~m[844]&m[845]&m[846]&~m[847])|(~m[841]&m[844]&~m[845]&~m[846]&m[847])|(~m[841]&~m[844]&m[845]&~m[846]&m[847])|(m[841]&m[844]&m[845]&~m[846]&m[847])|(~m[841]&m[844]&m[845]&m[846]&m[847]))&UnbiasedRNG[63])|((m[841]&~m[844]&~m[845]&m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&m[845]&~m[846]&m[847])|(~m[841]&~m[844]&~m[845]&m[846]&m[847])|(m[841]&~m[844]&~m[845]&m[846]&m[847])|(~m[841]&m[844]&~m[845]&m[846]&m[847])|(m[841]&m[844]&~m[845]&m[846]&m[847])|(~m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&m[844]&m[845]&m[846]&m[847]));
    m[848] = (((m[846]&~m[849]&~m[850]&~m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&m[851]&~m[852])|(m[846]&m[849]&~m[850]&m[851]&~m[852])|(m[846]&~m[849]&m[850]&m[851]&~m[852])|(~m[846]&m[849]&~m[850]&~m[851]&m[852])|(~m[846]&~m[849]&m[850]&~m[851]&m[852])|(m[846]&m[849]&m[850]&~m[851]&m[852])|(~m[846]&m[849]&m[850]&m[851]&m[852]))&UnbiasedRNG[64])|((m[846]&~m[849]&~m[850]&m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&m[850]&~m[851]&m[852])|(~m[846]&~m[849]&~m[850]&m[851]&m[852])|(m[846]&~m[849]&~m[850]&m[851]&m[852])|(~m[846]&m[849]&~m[850]&m[851]&m[852])|(m[846]&m[849]&~m[850]&m[851]&m[852])|(~m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&m[849]&m[850]&m[851]&m[852]));
    m[853] = (((m[851]&~m[854]&~m[855]&~m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&m[856]&~m[857])|(m[851]&m[854]&~m[855]&m[856]&~m[857])|(m[851]&~m[854]&m[855]&m[856]&~m[857])|(~m[851]&m[854]&~m[855]&~m[856]&m[857])|(~m[851]&~m[854]&m[855]&~m[856]&m[857])|(m[851]&m[854]&m[855]&~m[856]&m[857])|(~m[851]&m[854]&m[855]&m[856]&m[857]))&UnbiasedRNG[65])|((m[851]&~m[854]&~m[855]&m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&m[855]&~m[856]&m[857])|(~m[851]&~m[854]&~m[855]&m[856]&m[857])|(m[851]&~m[854]&~m[855]&m[856]&m[857])|(~m[851]&m[854]&~m[855]&m[856]&m[857])|(m[851]&m[854]&~m[855]&m[856]&m[857])|(~m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&m[854]&m[855]&m[856]&m[857]));
    m[863] = (((m[861]&~m[864]&~m[865]&~m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&m[866]&~m[867])|(m[861]&m[864]&~m[865]&m[866]&~m[867])|(m[861]&~m[864]&m[865]&m[866]&~m[867])|(~m[861]&m[864]&~m[865]&~m[866]&m[867])|(~m[861]&~m[864]&m[865]&~m[866]&m[867])|(m[861]&m[864]&m[865]&~m[866]&m[867])|(~m[861]&m[864]&m[865]&m[866]&m[867]))&UnbiasedRNG[66])|((m[861]&~m[864]&~m[865]&m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&m[865]&~m[866]&m[867])|(~m[861]&~m[864]&~m[865]&m[866]&m[867])|(m[861]&~m[864]&~m[865]&m[866]&m[867])|(~m[861]&m[864]&~m[865]&m[866]&m[867])|(m[861]&m[864]&~m[865]&m[866]&m[867])|(~m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&m[864]&m[865]&m[866]&m[867]));
    m[868] = (((m[866]&~m[869]&~m[870]&~m[871]&~m[872])|(~m[866]&~m[869]&~m[870]&m[871]&~m[872])|(m[866]&m[869]&~m[870]&m[871]&~m[872])|(m[866]&~m[869]&m[870]&m[871]&~m[872])|(~m[866]&m[869]&~m[870]&~m[871]&m[872])|(~m[866]&~m[869]&m[870]&~m[871]&m[872])|(m[866]&m[869]&m[870]&~m[871]&m[872])|(~m[866]&m[869]&m[870]&m[871]&m[872]))&UnbiasedRNG[67])|((m[866]&~m[869]&~m[870]&m[871]&~m[872])|(~m[866]&~m[869]&~m[870]&~m[871]&m[872])|(m[866]&~m[869]&~m[870]&~m[871]&m[872])|(m[866]&m[869]&~m[870]&~m[871]&m[872])|(m[866]&~m[869]&m[870]&~m[871]&m[872])|(~m[866]&~m[869]&~m[870]&m[871]&m[872])|(m[866]&~m[869]&~m[870]&m[871]&m[872])|(~m[866]&m[869]&~m[870]&m[871]&m[872])|(m[866]&m[869]&~m[870]&m[871]&m[872])|(~m[866]&~m[869]&m[870]&m[871]&m[872])|(m[866]&~m[869]&m[870]&m[871]&m[872])|(m[866]&m[869]&m[870]&m[871]&m[872]));
    m[873] = (((m[871]&~m[874]&~m[875]&~m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&m[876]&~m[877])|(m[871]&m[874]&~m[875]&m[876]&~m[877])|(m[871]&~m[874]&m[875]&m[876]&~m[877])|(~m[871]&m[874]&~m[875]&~m[876]&m[877])|(~m[871]&~m[874]&m[875]&~m[876]&m[877])|(m[871]&m[874]&m[875]&~m[876]&m[877])|(~m[871]&m[874]&m[875]&m[876]&m[877]))&UnbiasedRNG[68])|((m[871]&~m[874]&~m[875]&m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&m[875]&~m[876]&m[877])|(~m[871]&~m[874]&~m[875]&m[876]&m[877])|(m[871]&~m[874]&~m[875]&m[876]&m[877])|(~m[871]&m[874]&~m[875]&m[876]&m[877])|(m[871]&m[874]&~m[875]&m[876]&m[877])|(~m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&m[874]&m[875]&m[876]&m[877]));
    m[878] = (((m[876]&~m[879]&~m[880]&~m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&m[881]&~m[882])|(m[876]&m[879]&~m[880]&m[881]&~m[882])|(m[876]&~m[879]&m[880]&m[881]&~m[882])|(~m[876]&m[879]&~m[880]&~m[881]&m[882])|(~m[876]&~m[879]&m[880]&~m[881]&m[882])|(m[876]&m[879]&m[880]&~m[881]&m[882])|(~m[876]&m[879]&m[880]&m[881]&m[882]))&UnbiasedRNG[69])|((m[876]&~m[879]&~m[880]&m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&m[880]&~m[881]&m[882])|(~m[876]&~m[879]&~m[880]&m[881]&m[882])|(m[876]&~m[879]&~m[880]&m[881]&m[882])|(~m[876]&m[879]&~m[880]&m[881]&m[882])|(m[876]&m[879]&~m[880]&m[881]&m[882])|(~m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&m[879]&m[880]&m[881]&m[882]));
    m[883] = (((m[881]&~m[884]&~m[885]&~m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&m[886]&~m[887])|(m[881]&m[884]&~m[885]&m[886]&~m[887])|(m[881]&~m[884]&m[885]&m[886]&~m[887])|(~m[881]&m[884]&~m[885]&~m[886]&m[887])|(~m[881]&~m[884]&m[885]&~m[886]&m[887])|(m[881]&m[884]&m[885]&~m[886]&m[887])|(~m[881]&m[884]&m[885]&m[886]&m[887]))&UnbiasedRNG[70])|((m[881]&~m[884]&~m[885]&m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&m[885]&~m[886]&m[887])|(~m[881]&~m[884]&~m[885]&m[886]&m[887])|(m[881]&~m[884]&~m[885]&m[886]&m[887])|(~m[881]&m[884]&~m[885]&m[886]&m[887])|(m[881]&m[884]&~m[885]&m[886]&m[887])|(~m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&m[884]&m[885]&m[886]&m[887]));
    m[888] = (((m[886]&~m[889]&~m[890]&~m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&m[891]&~m[892])|(m[886]&m[889]&~m[890]&m[891]&~m[892])|(m[886]&~m[889]&m[890]&m[891]&~m[892])|(~m[886]&m[889]&~m[890]&~m[891]&m[892])|(~m[886]&~m[889]&m[890]&~m[891]&m[892])|(m[886]&m[889]&m[890]&~m[891]&m[892])|(~m[886]&m[889]&m[890]&m[891]&m[892]))&UnbiasedRNG[71])|((m[886]&~m[889]&~m[890]&m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&m[890]&~m[891]&m[892])|(~m[886]&~m[889]&~m[890]&m[891]&m[892])|(m[886]&~m[889]&~m[890]&m[891]&m[892])|(~m[886]&m[889]&~m[890]&m[891]&m[892])|(m[886]&m[889]&~m[890]&m[891]&m[892])|(~m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&m[889]&m[890]&m[891]&m[892]));
    m[893] = (((m[891]&~m[894]&~m[895]&~m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&m[896]&~m[897])|(m[891]&m[894]&~m[895]&m[896]&~m[897])|(m[891]&~m[894]&m[895]&m[896]&~m[897])|(~m[891]&m[894]&~m[895]&~m[896]&m[897])|(~m[891]&~m[894]&m[895]&~m[896]&m[897])|(m[891]&m[894]&m[895]&~m[896]&m[897])|(~m[891]&m[894]&m[895]&m[896]&m[897]))&UnbiasedRNG[72])|((m[891]&~m[894]&~m[895]&m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&m[895]&~m[896]&m[897])|(~m[891]&~m[894]&~m[895]&m[896]&m[897])|(m[891]&~m[894]&~m[895]&m[896]&m[897])|(~m[891]&m[894]&~m[895]&m[896]&m[897])|(m[891]&m[894]&~m[895]&m[896]&m[897])|(~m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&m[894]&m[895]&m[896]&m[897]));
    m[898] = (((m[896]&~m[899]&~m[900]&~m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&m[901]&~m[902])|(m[896]&m[899]&~m[900]&m[901]&~m[902])|(m[896]&~m[899]&m[900]&m[901]&~m[902])|(~m[896]&m[899]&~m[900]&~m[901]&m[902])|(~m[896]&~m[899]&m[900]&~m[901]&m[902])|(m[896]&m[899]&m[900]&~m[901]&m[902])|(~m[896]&m[899]&m[900]&m[901]&m[902]))&UnbiasedRNG[73])|((m[896]&~m[899]&~m[900]&m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&m[900]&~m[901]&m[902])|(~m[896]&~m[899]&~m[900]&m[901]&m[902])|(m[896]&~m[899]&~m[900]&m[901]&m[902])|(~m[896]&m[899]&~m[900]&m[901]&m[902])|(m[896]&m[899]&~m[900]&m[901]&m[902])|(~m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&m[899]&m[900]&m[901]&m[902]));
    m[903] = (((m[901]&~m[904]&~m[905]&~m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&m[906]&~m[907])|(m[901]&m[904]&~m[905]&m[906]&~m[907])|(m[901]&~m[904]&m[905]&m[906]&~m[907])|(~m[901]&m[904]&~m[905]&~m[906]&m[907])|(~m[901]&~m[904]&m[905]&~m[906]&m[907])|(m[901]&m[904]&m[905]&~m[906]&m[907])|(~m[901]&m[904]&m[905]&m[906]&m[907]))&UnbiasedRNG[74])|((m[901]&~m[904]&~m[905]&m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&m[905]&~m[906]&m[907])|(~m[901]&~m[904]&~m[905]&m[906]&m[907])|(m[901]&~m[904]&~m[905]&m[906]&m[907])|(~m[901]&m[904]&~m[905]&m[906]&m[907])|(m[901]&m[904]&~m[905]&m[906]&m[907])|(~m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&m[904]&m[905]&m[906]&m[907]));
    m[908] = (((m[906]&~m[909]&~m[910]&~m[911]&~m[912])|(~m[906]&~m[909]&~m[910]&m[911]&~m[912])|(m[906]&m[909]&~m[910]&m[911]&~m[912])|(m[906]&~m[909]&m[910]&m[911]&~m[912])|(~m[906]&m[909]&~m[910]&~m[911]&m[912])|(~m[906]&~m[909]&m[910]&~m[911]&m[912])|(m[906]&m[909]&m[910]&~m[911]&m[912])|(~m[906]&m[909]&m[910]&m[911]&m[912]))&UnbiasedRNG[75])|((m[906]&~m[909]&~m[910]&m[911]&~m[912])|(~m[906]&~m[909]&~m[910]&~m[911]&m[912])|(m[906]&~m[909]&~m[910]&~m[911]&m[912])|(m[906]&m[909]&~m[910]&~m[911]&m[912])|(m[906]&~m[909]&m[910]&~m[911]&m[912])|(~m[906]&~m[909]&~m[910]&m[911]&m[912])|(m[906]&~m[909]&~m[910]&m[911]&m[912])|(~m[906]&m[909]&~m[910]&m[911]&m[912])|(m[906]&m[909]&~m[910]&m[911]&m[912])|(~m[906]&~m[909]&m[910]&m[911]&m[912])|(m[906]&~m[909]&m[910]&m[911]&m[912])|(m[906]&m[909]&m[910]&m[911]&m[912]));
    m[913] = (((m[862]&~m[914]&~m[915]&~m[916]&~m[917])|(~m[862]&~m[914]&~m[915]&m[916]&~m[917])|(m[862]&m[914]&~m[915]&m[916]&~m[917])|(m[862]&~m[914]&m[915]&m[916]&~m[917])|(~m[862]&m[914]&~m[915]&~m[916]&m[917])|(~m[862]&~m[914]&m[915]&~m[916]&m[917])|(m[862]&m[914]&m[915]&~m[916]&m[917])|(~m[862]&m[914]&m[915]&m[916]&m[917]))&UnbiasedRNG[76])|((m[862]&~m[914]&~m[915]&m[916]&~m[917])|(~m[862]&~m[914]&~m[915]&~m[916]&m[917])|(m[862]&~m[914]&~m[915]&~m[916]&m[917])|(m[862]&m[914]&~m[915]&~m[916]&m[917])|(m[862]&~m[914]&m[915]&~m[916]&m[917])|(~m[862]&~m[914]&~m[915]&m[916]&m[917])|(m[862]&~m[914]&~m[915]&m[916]&m[917])|(~m[862]&m[914]&~m[915]&m[916]&m[917])|(m[862]&m[914]&~m[915]&m[916]&m[917])|(~m[862]&~m[914]&m[915]&m[916]&m[917])|(m[862]&~m[914]&m[915]&m[916]&m[917])|(m[862]&m[914]&m[915]&m[916]&m[917]));
    m[918] = (((m[916]&~m[919]&~m[920]&~m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&m[921]&~m[922])|(m[916]&m[919]&~m[920]&m[921]&~m[922])|(m[916]&~m[919]&m[920]&m[921]&~m[922])|(~m[916]&m[919]&~m[920]&~m[921]&m[922])|(~m[916]&~m[919]&m[920]&~m[921]&m[922])|(m[916]&m[919]&m[920]&~m[921]&m[922])|(~m[916]&m[919]&m[920]&m[921]&m[922]))&UnbiasedRNG[77])|((m[916]&~m[919]&~m[920]&m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&m[920]&~m[921]&m[922])|(~m[916]&~m[919]&~m[920]&m[921]&m[922])|(m[916]&~m[919]&~m[920]&m[921]&m[922])|(~m[916]&m[919]&~m[920]&m[921]&m[922])|(m[916]&m[919]&~m[920]&m[921]&m[922])|(~m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&m[919]&m[920]&m[921]&m[922]));
    m[923] = (((m[921]&~m[924]&~m[925]&~m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&m[926]&~m[927])|(m[921]&m[924]&~m[925]&m[926]&~m[927])|(m[921]&~m[924]&m[925]&m[926]&~m[927])|(~m[921]&m[924]&~m[925]&~m[926]&m[927])|(~m[921]&~m[924]&m[925]&~m[926]&m[927])|(m[921]&m[924]&m[925]&~m[926]&m[927])|(~m[921]&m[924]&m[925]&m[926]&m[927]))&UnbiasedRNG[78])|((m[921]&~m[924]&~m[925]&m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&m[925]&~m[926]&m[927])|(~m[921]&~m[924]&~m[925]&m[926]&m[927])|(m[921]&~m[924]&~m[925]&m[926]&m[927])|(~m[921]&m[924]&~m[925]&m[926]&m[927])|(m[921]&m[924]&~m[925]&m[926]&m[927])|(~m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&m[924]&m[925]&m[926]&m[927]));
    m[928] = (((m[926]&~m[929]&~m[930]&~m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&m[931]&~m[932])|(m[926]&m[929]&~m[930]&m[931]&~m[932])|(m[926]&~m[929]&m[930]&m[931]&~m[932])|(~m[926]&m[929]&~m[930]&~m[931]&m[932])|(~m[926]&~m[929]&m[930]&~m[931]&m[932])|(m[926]&m[929]&m[930]&~m[931]&m[932])|(~m[926]&m[929]&m[930]&m[931]&m[932]))&UnbiasedRNG[79])|((m[926]&~m[929]&~m[930]&m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&m[930]&~m[931]&m[932])|(~m[926]&~m[929]&~m[930]&m[931]&m[932])|(m[926]&~m[929]&~m[930]&m[931]&m[932])|(~m[926]&m[929]&~m[930]&m[931]&m[932])|(m[926]&m[929]&~m[930]&m[931]&m[932])|(~m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&m[929]&m[930]&m[931]&m[932]));
    m[933] = (((m[931]&~m[934]&~m[935]&~m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&m[936]&~m[937])|(m[931]&m[934]&~m[935]&m[936]&~m[937])|(m[931]&~m[934]&m[935]&m[936]&~m[937])|(~m[931]&m[934]&~m[935]&~m[936]&m[937])|(~m[931]&~m[934]&m[935]&~m[936]&m[937])|(m[931]&m[934]&m[935]&~m[936]&m[937])|(~m[931]&m[934]&m[935]&m[936]&m[937]))&UnbiasedRNG[80])|((m[931]&~m[934]&~m[935]&m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&m[935]&~m[936]&m[937])|(~m[931]&~m[934]&~m[935]&m[936]&m[937])|(m[931]&~m[934]&~m[935]&m[936]&m[937])|(~m[931]&m[934]&~m[935]&m[936]&m[937])|(m[931]&m[934]&~m[935]&m[936]&m[937])|(~m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&m[934]&m[935]&m[936]&m[937]));
    m[938] = (((m[936]&~m[939]&~m[940]&~m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&m[941]&~m[942])|(m[936]&m[939]&~m[940]&m[941]&~m[942])|(m[936]&~m[939]&m[940]&m[941]&~m[942])|(~m[936]&m[939]&~m[940]&~m[941]&m[942])|(~m[936]&~m[939]&m[940]&~m[941]&m[942])|(m[936]&m[939]&m[940]&~m[941]&m[942])|(~m[936]&m[939]&m[940]&m[941]&m[942]))&UnbiasedRNG[81])|((m[936]&~m[939]&~m[940]&m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&m[940]&~m[941]&m[942])|(~m[936]&~m[939]&~m[940]&m[941]&m[942])|(m[936]&~m[939]&~m[940]&m[941]&m[942])|(~m[936]&m[939]&~m[940]&m[941]&m[942])|(m[936]&m[939]&~m[940]&m[941]&m[942])|(~m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&m[939]&m[940]&m[941]&m[942]));
    m[943] = (((m[941]&~m[944]&~m[945]&~m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&m[946]&~m[947])|(m[941]&m[944]&~m[945]&m[946]&~m[947])|(m[941]&~m[944]&m[945]&m[946]&~m[947])|(~m[941]&m[944]&~m[945]&~m[946]&m[947])|(~m[941]&~m[944]&m[945]&~m[946]&m[947])|(m[941]&m[944]&m[945]&~m[946]&m[947])|(~m[941]&m[944]&m[945]&m[946]&m[947]))&UnbiasedRNG[82])|((m[941]&~m[944]&~m[945]&m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&m[945]&~m[946]&m[947])|(~m[941]&~m[944]&~m[945]&m[946]&m[947])|(m[941]&~m[944]&~m[945]&m[946]&m[947])|(~m[941]&m[944]&~m[945]&m[946]&m[947])|(m[941]&m[944]&~m[945]&m[946]&m[947])|(~m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&m[944]&m[945]&m[946]&m[947]));
    m[948] = (((m[946]&~m[949]&~m[950]&~m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&m[951]&~m[952])|(m[946]&m[949]&~m[950]&m[951]&~m[952])|(m[946]&~m[949]&m[950]&m[951]&~m[952])|(~m[946]&m[949]&~m[950]&~m[951]&m[952])|(~m[946]&~m[949]&m[950]&~m[951]&m[952])|(m[946]&m[949]&m[950]&~m[951]&m[952])|(~m[946]&m[949]&m[950]&m[951]&m[952]))&UnbiasedRNG[83])|((m[946]&~m[949]&~m[950]&m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&m[950]&~m[951]&m[952])|(~m[946]&~m[949]&~m[950]&m[951]&m[952])|(m[946]&~m[949]&~m[950]&m[951]&m[952])|(~m[946]&m[949]&~m[950]&m[951]&m[952])|(m[946]&m[949]&~m[950]&m[951]&m[952])|(~m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&m[949]&m[950]&m[951]&m[952]));
    m[953] = (((m[951]&~m[954]&~m[955]&~m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&m[956]&~m[957])|(m[951]&m[954]&~m[955]&m[956]&~m[957])|(m[951]&~m[954]&m[955]&m[956]&~m[957])|(~m[951]&m[954]&~m[955]&~m[956]&m[957])|(~m[951]&~m[954]&m[955]&~m[956]&m[957])|(m[951]&m[954]&m[955]&~m[956]&m[957])|(~m[951]&m[954]&m[955]&m[956]&m[957]))&UnbiasedRNG[84])|((m[951]&~m[954]&~m[955]&m[956]&~m[957])|(~m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&~m[955]&~m[956]&m[957])|(m[951]&m[954]&~m[955]&~m[956]&m[957])|(m[951]&~m[954]&m[955]&~m[956]&m[957])|(~m[951]&~m[954]&~m[955]&m[956]&m[957])|(m[951]&~m[954]&~m[955]&m[956]&m[957])|(~m[951]&m[954]&~m[955]&m[956]&m[957])|(m[951]&m[954]&~m[955]&m[956]&m[957])|(~m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&~m[954]&m[955]&m[956]&m[957])|(m[951]&m[954]&m[955]&m[956]&m[957]));
    m[958] = (((m[956]&~m[959]&~m[960]&~m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&m[961]&~m[962])|(m[956]&m[959]&~m[960]&m[961]&~m[962])|(m[956]&~m[959]&m[960]&m[961]&~m[962])|(~m[956]&m[959]&~m[960]&~m[961]&m[962])|(~m[956]&~m[959]&m[960]&~m[961]&m[962])|(m[956]&m[959]&m[960]&~m[961]&m[962])|(~m[956]&m[959]&m[960]&m[961]&m[962]))&UnbiasedRNG[85])|((m[956]&~m[959]&~m[960]&m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&m[960]&~m[961]&m[962])|(~m[956]&~m[959]&~m[960]&m[961]&m[962])|(m[956]&~m[959]&~m[960]&m[961]&m[962])|(~m[956]&m[959]&~m[960]&m[961]&m[962])|(m[956]&m[959]&~m[960]&m[961]&m[962])|(~m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&m[959]&m[960]&m[961]&m[962]));
    m[963] = (((m[917]&~m[964]&~m[965]&~m[966]&~m[967])|(~m[917]&~m[964]&~m[965]&m[966]&~m[967])|(m[917]&m[964]&~m[965]&m[966]&~m[967])|(m[917]&~m[964]&m[965]&m[966]&~m[967])|(~m[917]&m[964]&~m[965]&~m[966]&m[967])|(~m[917]&~m[964]&m[965]&~m[966]&m[967])|(m[917]&m[964]&m[965]&~m[966]&m[967])|(~m[917]&m[964]&m[965]&m[966]&m[967]))&UnbiasedRNG[86])|((m[917]&~m[964]&~m[965]&m[966]&~m[967])|(~m[917]&~m[964]&~m[965]&~m[966]&m[967])|(m[917]&~m[964]&~m[965]&~m[966]&m[967])|(m[917]&m[964]&~m[965]&~m[966]&m[967])|(m[917]&~m[964]&m[965]&~m[966]&m[967])|(~m[917]&~m[964]&~m[965]&m[966]&m[967])|(m[917]&~m[964]&~m[965]&m[966]&m[967])|(~m[917]&m[964]&~m[965]&m[966]&m[967])|(m[917]&m[964]&~m[965]&m[966]&m[967])|(~m[917]&~m[964]&m[965]&m[966]&m[967])|(m[917]&~m[964]&m[965]&m[966]&m[967])|(m[917]&m[964]&m[965]&m[966]&m[967]));
    m[968] = (((m[966]&~m[969]&~m[970]&~m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&m[971]&~m[972])|(m[966]&m[969]&~m[970]&m[971]&~m[972])|(m[966]&~m[969]&m[970]&m[971]&~m[972])|(~m[966]&m[969]&~m[970]&~m[971]&m[972])|(~m[966]&~m[969]&m[970]&~m[971]&m[972])|(m[966]&m[969]&m[970]&~m[971]&m[972])|(~m[966]&m[969]&m[970]&m[971]&m[972]))&UnbiasedRNG[87])|((m[966]&~m[969]&~m[970]&m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&m[970]&~m[971]&m[972])|(~m[966]&~m[969]&~m[970]&m[971]&m[972])|(m[966]&~m[969]&~m[970]&m[971]&m[972])|(~m[966]&m[969]&~m[970]&m[971]&m[972])|(m[966]&m[969]&~m[970]&m[971]&m[972])|(~m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&m[969]&m[970]&m[971]&m[972]));
    m[973] = (((m[971]&~m[974]&~m[975]&~m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&m[976]&~m[977])|(m[971]&m[974]&~m[975]&m[976]&~m[977])|(m[971]&~m[974]&m[975]&m[976]&~m[977])|(~m[971]&m[974]&~m[975]&~m[976]&m[977])|(~m[971]&~m[974]&m[975]&~m[976]&m[977])|(m[971]&m[974]&m[975]&~m[976]&m[977])|(~m[971]&m[974]&m[975]&m[976]&m[977]))&UnbiasedRNG[88])|((m[971]&~m[974]&~m[975]&m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&m[975]&~m[976]&m[977])|(~m[971]&~m[974]&~m[975]&m[976]&m[977])|(m[971]&~m[974]&~m[975]&m[976]&m[977])|(~m[971]&m[974]&~m[975]&m[976]&m[977])|(m[971]&m[974]&~m[975]&m[976]&m[977])|(~m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&m[974]&m[975]&m[976]&m[977]));
    m[978] = (((m[976]&~m[979]&~m[980]&~m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&m[981]&~m[982])|(m[976]&m[979]&~m[980]&m[981]&~m[982])|(m[976]&~m[979]&m[980]&m[981]&~m[982])|(~m[976]&m[979]&~m[980]&~m[981]&m[982])|(~m[976]&~m[979]&m[980]&~m[981]&m[982])|(m[976]&m[979]&m[980]&~m[981]&m[982])|(~m[976]&m[979]&m[980]&m[981]&m[982]))&UnbiasedRNG[89])|((m[976]&~m[979]&~m[980]&m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&m[980]&~m[981]&m[982])|(~m[976]&~m[979]&~m[980]&m[981]&m[982])|(m[976]&~m[979]&~m[980]&m[981]&m[982])|(~m[976]&m[979]&~m[980]&m[981]&m[982])|(m[976]&m[979]&~m[980]&m[981]&m[982])|(~m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&m[979]&m[980]&m[981]&m[982]));
    m[983] = (((m[981]&~m[984]&~m[985]&~m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&m[986]&~m[987])|(m[981]&m[984]&~m[985]&m[986]&~m[987])|(m[981]&~m[984]&m[985]&m[986]&~m[987])|(~m[981]&m[984]&~m[985]&~m[986]&m[987])|(~m[981]&~m[984]&m[985]&~m[986]&m[987])|(m[981]&m[984]&m[985]&~m[986]&m[987])|(~m[981]&m[984]&m[985]&m[986]&m[987]))&UnbiasedRNG[90])|((m[981]&~m[984]&~m[985]&m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&m[985]&~m[986]&m[987])|(~m[981]&~m[984]&~m[985]&m[986]&m[987])|(m[981]&~m[984]&~m[985]&m[986]&m[987])|(~m[981]&m[984]&~m[985]&m[986]&m[987])|(m[981]&m[984]&~m[985]&m[986]&m[987])|(~m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&m[984]&m[985]&m[986]&m[987]));
    m[988] = (((m[986]&~m[989]&~m[990]&~m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&m[991]&~m[992])|(m[986]&m[989]&~m[990]&m[991]&~m[992])|(m[986]&~m[989]&m[990]&m[991]&~m[992])|(~m[986]&m[989]&~m[990]&~m[991]&m[992])|(~m[986]&~m[989]&m[990]&~m[991]&m[992])|(m[986]&m[989]&m[990]&~m[991]&m[992])|(~m[986]&m[989]&m[990]&m[991]&m[992]))&UnbiasedRNG[91])|((m[986]&~m[989]&~m[990]&m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&m[990]&~m[991]&m[992])|(~m[986]&~m[989]&~m[990]&m[991]&m[992])|(m[986]&~m[989]&~m[990]&m[991]&m[992])|(~m[986]&m[989]&~m[990]&m[991]&m[992])|(m[986]&m[989]&~m[990]&m[991]&m[992])|(~m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&m[989]&m[990]&m[991]&m[992]));
    m[993] = (((m[991]&~m[994]&~m[995]&~m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&m[996]&~m[997])|(m[991]&m[994]&~m[995]&m[996]&~m[997])|(m[991]&~m[994]&m[995]&m[996]&~m[997])|(~m[991]&m[994]&~m[995]&~m[996]&m[997])|(~m[991]&~m[994]&m[995]&~m[996]&m[997])|(m[991]&m[994]&m[995]&~m[996]&m[997])|(~m[991]&m[994]&m[995]&m[996]&m[997]))&UnbiasedRNG[92])|((m[991]&~m[994]&~m[995]&m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&m[995]&~m[996]&m[997])|(~m[991]&~m[994]&~m[995]&m[996]&m[997])|(m[991]&~m[994]&~m[995]&m[996]&m[997])|(~m[991]&m[994]&~m[995]&m[996]&m[997])|(m[991]&m[994]&~m[995]&m[996]&m[997])|(~m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&m[994]&m[995]&m[996]&m[997]));
    m[998] = (((m[996]&~m[999]&~m[1000]&~m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&~m[1002])|(~m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&m[999]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[93])|((m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&m[999]&m[1000]&m[1001]&m[1002]));
    m[1003] = (((m[1001]&~m[1004]&~m[1005]&~m[1006]&~m[1007])|(~m[1001]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(m[1001]&m[1004]&~m[1005]&m[1006]&~m[1007])|(m[1001]&~m[1004]&m[1005]&m[1006]&~m[1007])|(~m[1001]&m[1004]&~m[1005]&~m[1006]&m[1007])|(~m[1001]&~m[1004]&m[1005]&~m[1006]&m[1007])|(m[1001]&m[1004]&m[1005]&~m[1006]&m[1007])|(~m[1001]&m[1004]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[94])|((m[1001]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(~m[1001]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[1001]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[1001]&m[1004]&~m[1005]&~m[1006]&m[1007])|(m[1001]&~m[1004]&m[1005]&~m[1006]&m[1007])|(~m[1001]&~m[1004]&~m[1005]&m[1006]&m[1007])|(m[1001]&~m[1004]&~m[1005]&m[1006]&m[1007])|(~m[1001]&m[1004]&~m[1005]&m[1006]&m[1007])|(m[1001]&m[1004]&~m[1005]&m[1006]&m[1007])|(~m[1001]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[1001]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[1001]&m[1004]&m[1005]&m[1006]&m[1007]));
    m[1008] = (((m[967]&~m[1009]&~m[1010]&~m[1011]&~m[1012])|(~m[967]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(m[967]&m[1009]&~m[1010]&m[1011]&~m[1012])|(m[967]&~m[1009]&m[1010]&m[1011]&~m[1012])|(~m[967]&m[1009]&~m[1010]&~m[1011]&m[1012])|(~m[967]&~m[1009]&m[1010]&~m[1011]&m[1012])|(m[967]&m[1009]&m[1010]&~m[1011]&m[1012])|(~m[967]&m[1009]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[95])|((m[967]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(~m[967]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[967]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[967]&m[1009]&~m[1010]&~m[1011]&m[1012])|(m[967]&~m[1009]&m[1010]&~m[1011]&m[1012])|(~m[967]&~m[1009]&~m[1010]&m[1011]&m[1012])|(m[967]&~m[1009]&~m[1010]&m[1011]&m[1012])|(~m[967]&m[1009]&~m[1010]&m[1011]&m[1012])|(m[967]&m[1009]&~m[1010]&m[1011]&m[1012])|(~m[967]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[967]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[967]&m[1009]&m[1010]&m[1011]&m[1012]));
    m[1013] = (((m[1011]&~m[1014]&~m[1015]&~m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&~m[1017])|(~m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[96])|((m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&m[1016]&m[1017]));
    m[1018] = (((m[1016]&~m[1019]&~m[1020]&~m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&~m[1022])|(~m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[97])|((m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&m[1021]&m[1022]));
    m[1023] = (((m[1021]&~m[1024]&~m[1025]&~m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&~m[1027])|(~m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[98])|((m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&m[1026]&m[1027]));
    m[1028] = (((m[1026]&~m[1029]&~m[1030]&~m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&~m[1032])|(~m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[99])|((m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&m[1031]&m[1032]));
    m[1033] = (((m[1031]&~m[1034]&~m[1035]&~m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&~m[1037])|(~m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&m[1034]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[100])|((m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&m[1036]&m[1037]));
    m[1038] = (((m[1036]&~m[1039]&~m[1040]&~m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&~m[1042])|(~m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[101])|((m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&m[1041]&m[1042]));
    m[1043] = (((m[1041]&~m[1044]&~m[1045]&~m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&~m[1047])|(~m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[102])|((m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&m[1046]&m[1047]));
    m[1048] = (((m[1012]&~m[1049]&~m[1050]&~m[1051]&~m[1052])|(~m[1012]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1012]&m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1012]&~m[1049]&m[1050]&m[1051]&~m[1052])|(~m[1012]&m[1049]&~m[1050]&~m[1051]&m[1052])|(~m[1012]&~m[1049]&m[1050]&~m[1051]&m[1052])|(m[1012]&m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1012]&m[1049]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[103])|((m[1012]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(~m[1012]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1012]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1012]&m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1012]&~m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1012]&~m[1049]&~m[1050]&m[1051]&m[1052])|(m[1012]&~m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1012]&m[1049]&~m[1050]&m[1051]&m[1052])|(m[1012]&m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1012]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1012]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1012]&m[1049]&m[1050]&m[1051]&m[1052]));
    m[1053] = (((m[1051]&~m[1054]&~m[1055]&~m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&~m[1057])|(~m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[104])|((m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&m[1056]&m[1057]));
    m[1058] = (((m[1056]&~m[1059]&~m[1060]&~m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&~m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&~m[1062])|(~m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&m[1059]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[105])|((m[1056]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(~m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&~m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&~m[1061]&m[1062])|(~m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&~m[1060]&m[1061]&m[1062])|(~m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[1056]&m[1059]&m[1060]&m[1061]&m[1062]));
    m[1063] = (((m[1061]&~m[1064]&~m[1065]&~m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&~m[1067])|(~m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[106])|((m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&m[1066]&m[1067]));
    m[1068] = (((m[1066]&~m[1069]&~m[1070]&~m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&~m[1072])|(~m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&m[1069]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[107])|((m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&m[1071]&m[1072]));
    m[1073] = (((m[1071]&~m[1074]&~m[1075]&~m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&~m[1077])|(~m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[108])|((m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&m[1076]&m[1077]));
    m[1078] = (((m[1076]&~m[1079]&~m[1080]&~m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&~m[1082])|(~m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[109])|((m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&m[1081]&m[1082]));
    m[1083] = (((m[1052]&~m[1084]&~m[1085]&~m[1086]&~m[1087])|(~m[1052]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1052]&m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1052]&~m[1084]&m[1085]&m[1086]&~m[1087])|(~m[1052]&m[1084]&~m[1085]&~m[1086]&m[1087])|(~m[1052]&~m[1084]&m[1085]&~m[1086]&m[1087])|(m[1052]&m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1052]&m[1084]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[110])|((m[1052]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(~m[1052]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1052]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1052]&m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1052]&~m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1052]&~m[1084]&~m[1085]&m[1086]&m[1087])|(m[1052]&~m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1052]&m[1084]&~m[1085]&m[1086]&m[1087])|(m[1052]&m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1052]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1052]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1052]&m[1084]&m[1085]&m[1086]&m[1087]));
    m[1088] = (((m[1086]&~m[1089]&~m[1090]&~m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&~m[1092])|(~m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[111])|((m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&m[1091]&m[1092]));
    m[1093] = (((m[1091]&~m[1094]&~m[1095]&~m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&~m[1097])|(~m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[112])|((m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&m[1096]&m[1097]));
    m[1098] = (((m[1096]&~m[1099]&~m[1100]&~m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&~m[1102])|(~m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[113])|((m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&m[1101]&m[1102]));
    m[1103] = (((m[1101]&~m[1104]&~m[1105]&~m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&~m[1107])|(~m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[114])|((m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&m[1106]&m[1107]));
    m[1108] = (((m[1106]&~m[1109]&~m[1110]&~m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&~m[1112])|(~m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&m[1109]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[115])|((m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&m[1111]&m[1112]));
    m[1113] = (((m[1087]&~m[1114]&~m[1115]&~m[1116]&~m[1117])|(~m[1087]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1087]&m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1087]&~m[1114]&m[1115]&m[1116]&~m[1117])|(~m[1087]&m[1114]&~m[1115]&~m[1116]&m[1117])|(~m[1087]&~m[1114]&m[1115]&~m[1116]&m[1117])|(m[1087]&m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1087]&m[1114]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[116])|((m[1087]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(~m[1087]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1087]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1087]&m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1087]&~m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1087]&~m[1114]&~m[1115]&m[1116]&m[1117])|(m[1087]&~m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1087]&m[1114]&~m[1115]&m[1116]&m[1117])|(m[1087]&m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1087]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1087]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1087]&m[1114]&m[1115]&m[1116]&m[1117]));
    m[1118] = (((m[1116]&~m[1119]&~m[1120]&~m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&~m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&~m[1122])|(~m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&m[1119]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[117])|((m[1116]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(~m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&~m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&~m[1121]&m[1122])|(~m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&~m[1120]&m[1121]&m[1122])|(~m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[1116]&m[1119]&m[1120]&m[1121]&m[1122]));
    m[1123] = (((m[1121]&~m[1124]&~m[1125]&~m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&~m[1127])|(~m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[118])|((m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&m[1126]&m[1127]));
    m[1128] = (((m[1126]&~m[1129]&~m[1130]&~m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&~m[1132])|(~m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[119])|((m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&m[1131]&m[1132]));
    m[1133] = (((m[1131]&~m[1134]&~m[1135]&~m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&~m[1137])|(~m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[120])|((m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&m[1136]&m[1137]));
    m[1138] = (((m[1117]&~m[1139]&~m[1140]&~m[1141]&~m[1142])|(~m[1117]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1117]&m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1117]&~m[1139]&m[1140]&m[1141]&~m[1142])|(~m[1117]&m[1139]&~m[1140]&~m[1141]&m[1142])|(~m[1117]&~m[1139]&m[1140]&~m[1141]&m[1142])|(m[1117]&m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1117]&m[1139]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[121])|((m[1117]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(~m[1117]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1117]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1117]&m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1117]&~m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1117]&~m[1139]&~m[1140]&m[1141]&m[1142])|(m[1117]&~m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1117]&m[1139]&~m[1140]&m[1141]&m[1142])|(m[1117]&m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1117]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1117]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1117]&m[1139]&m[1140]&m[1141]&m[1142]));
    m[1143] = (((m[1141]&~m[1144]&~m[1145]&~m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&~m[1147])|(~m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[122])|((m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&m[1146]&m[1147]));
    m[1148] = (((m[1146]&~m[1149]&~m[1150]&~m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&~m[1152])|(~m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[123])|((m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&m[1151]&m[1152]));
    m[1153] = (((m[1151]&~m[1154]&~m[1155]&~m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&~m[1157])|(~m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&m[1154]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[124])|((m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&m[1156]&m[1157]));
    m[1158] = (((m[1142]&~m[1159]&~m[1160]&~m[1161]&~m[1162])|(~m[1142]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1142]&m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1142]&~m[1159]&m[1160]&m[1161]&~m[1162])|(~m[1142]&m[1159]&~m[1160]&~m[1161]&m[1162])|(~m[1142]&~m[1159]&m[1160]&~m[1161]&m[1162])|(m[1142]&m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1142]&m[1159]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[125])|((m[1142]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(~m[1142]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1142]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1142]&m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1142]&~m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1142]&~m[1159]&~m[1160]&m[1161]&m[1162])|(m[1142]&~m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1142]&m[1159]&~m[1160]&m[1161]&m[1162])|(m[1142]&m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1142]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1142]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1142]&m[1159]&m[1160]&m[1161]&m[1162]));
    m[1163] = (((m[1161]&~m[1164]&~m[1165]&~m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&~m[1167])|(~m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[126])|((m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&m[1166]&m[1167]));
    m[1168] = (((m[1166]&~m[1169]&~m[1170]&~m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&~m[1172])|(~m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[127])|((m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&m[1171]&m[1172]));
    m[1173] = (((m[1162]&~m[1174]&~m[1175]&~m[1176]&~m[1177])|(~m[1162]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1162]&m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1162]&~m[1174]&m[1175]&m[1176]&~m[1177])|(~m[1162]&m[1174]&~m[1175]&~m[1176]&m[1177])|(~m[1162]&~m[1174]&m[1175]&~m[1176]&m[1177])|(m[1162]&m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1162]&m[1174]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[128])|((m[1162]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(~m[1162]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1162]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1162]&m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1162]&~m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1162]&~m[1174]&~m[1175]&m[1176]&m[1177])|(m[1162]&~m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1162]&m[1174]&~m[1175]&m[1176]&m[1177])|(m[1162]&m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1162]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1162]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1162]&m[1174]&m[1175]&m[1176]&m[1177]));
    m[1178] = (((m[1176]&~m[1179]&~m[1180]&~m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&~m[1182])|(~m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[129])|((m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&m[1181]&m[1182]));
    m[1183] = (((m[1177]&~m[1184]&~m[1185]&~m[1186]&~m[1187])|(~m[1177]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1177]&m[1184]&~m[1185]&m[1186]&~m[1187])|(m[1177]&~m[1184]&m[1185]&m[1186]&~m[1187])|(~m[1177]&m[1184]&~m[1185]&~m[1186]&m[1187])|(~m[1177]&~m[1184]&m[1185]&~m[1186]&m[1187])|(m[1177]&m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1177]&m[1184]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[130])|((m[1177]&~m[1184]&~m[1185]&m[1186]&~m[1187])|(~m[1177]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1177]&~m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1177]&m[1184]&~m[1185]&~m[1186]&m[1187])|(m[1177]&~m[1184]&m[1185]&~m[1186]&m[1187])|(~m[1177]&~m[1184]&~m[1185]&m[1186]&m[1187])|(m[1177]&~m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1177]&m[1184]&~m[1185]&m[1186]&m[1187])|(m[1177]&m[1184]&~m[1185]&m[1186]&m[1187])|(~m[1177]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1177]&~m[1184]&m[1185]&m[1186]&m[1187])|(m[1177]&m[1184]&m[1185]&m[1186]&m[1187]));
end

always @(posedge color1_clk) begin
    m[24] = (((m[0]&m[96]&~m[97]&~m[98]&~m[99])|(m[0]&~m[96]&m[97]&~m[98]&~m[99])|(~m[0]&m[96]&m[97]&~m[98]&~m[99])|(m[0]&~m[96]&~m[97]&m[98]&~m[99])|(~m[0]&m[96]&~m[97]&m[98]&~m[99])|(~m[0]&~m[96]&m[97]&m[98]&~m[99])|(m[0]&~m[96]&~m[97]&~m[98]&m[99])|(~m[0]&m[96]&~m[97]&~m[98]&m[99])|(~m[0]&~m[96]&m[97]&~m[98]&m[99])|(~m[0]&~m[96]&~m[97]&m[98]&m[99]))&BiasedRNG[168])|(((m[0]&m[96]&m[97]&~m[98]&~m[99])|(m[0]&m[96]&~m[97]&m[98]&~m[99])|(m[0]&~m[96]&m[97]&m[98]&~m[99])|(~m[0]&m[96]&m[97]&m[98]&~m[99])|(m[0]&m[96]&~m[97]&~m[98]&m[99])|(m[0]&~m[96]&m[97]&~m[98]&m[99])|(~m[0]&m[96]&m[97]&~m[98]&m[99])|(m[0]&~m[96]&~m[97]&m[98]&m[99])|(~m[0]&m[96]&~m[97]&m[98]&m[99])|(~m[0]&~m[96]&m[97]&m[98]&m[99]))&~BiasedRNG[168])|((m[0]&m[96]&m[97]&m[98]&~m[99])|(m[0]&m[96]&m[97]&~m[98]&m[99])|(m[0]&m[96]&~m[97]&m[98]&m[99])|(m[0]&~m[96]&m[97]&m[98]&m[99])|(~m[0]&m[96]&m[97]&m[98]&m[99])|(m[0]&m[96]&m[97]&m[98]&m[99]));
    m[25] = (((m[0]&m[100]&~m[101]&~m[102]&~m[103])|(m[0]&~m[100]&m[101]&~m[102]&~m[103])|(~m[0]&m[100]&m[101]&~m[102]&~m[103])|(m[0]&~m[100]&~m[101]&m[102]&~m[103])|(~m[0]&m[100]&~m[101]&m[102]&~m[103])|(~m[0]&~m[100]&m[101]&m[102]&~m[103])|(m[0]&~m[100]&~m[101]&~m[102]&m[103])|(~m[0]&m[100]&~m[101]&~m[102]&m[103])|(~m[0]&~m[100]&m[101]&~m[102]&m[103])|(~m[0]&~m[100]&~m[101]&m[102]&m[103]))&BiasedRNG[169])|(((m[0]&m[100]&m[101]&~m[102]&~m[103])|(m[0]&m[100]&~m[101]&m[102]&~m[103])|(m[0]&~m[100]&m[101]&m[102]&~m[103])|(~m[0]&m[100]&m[101]&m[102]&~m[103])|(m[0]&m[100]&~m[101]&~m[102]&m[103])|(m[0]&~m[100]&m[101]&~m[102]&m[103])|(~m[0]&m[100]&m[101]&~m[102]&m[103])|(m[0]&~m[100]&~m[101]&m[102]&m[103])|(~m[0]&m[100]&~m[101]&m[102]&m[103])|(~m[0]&~m[100]&m[101]&m[102]&m[103]))&~BiasedRNG[169])|((m[0]&m[100]&m[101]&m[102]&~m[103])|(m[0]&m[100]&m[101]&~m[102]&m[103])|(m[0]&m[100]&~m[101]&m[102]&m[103])|(m[0]&~m[100]&m[101]&m[102]&m[103])|(~m[0]&m[100]&m[101]&m[102]&m[103])|(m[0]&m[100]&m[101]&m[102]&m[103]));
    m[26] = (((m[0]&m[104]&~m[105]&~m[106]&~m[107])|(m[0]&~m[104]&m[105]&~m[106]&~m[107])|(~m[0]&m[104]&m[105]&~m[106]&~m[107])|(m[0]&~m[104]&~m[105]&m[106]&~m[107])|(~m[0]&m[104]&~m[105]&m[106]&~m[107])|(~m[0]&~m[104]&m[105]&m[106]&~m[107])|(m[0]&~m[104]&~m[105]&~m[106]&m[107])|(~m[0]&m[104]&~m[105]&~m[106]&m[107])|(~m[0]&~m[104]&m[105]&~m[106]&m[107])|(~m[0]&~m[104]&~m[105]&m[106]&m[107]))&BiasedRNG[170])|(((m[0]&m[104]&m[105]&~m[106]&~m[107])|(m[0]&m[104]&~m[105]&m[106]&~m[107])|(m[0]&~m[104]&m[105]&m[106]&~m[107])|(~m[0]&m[104]&m[105]&m[106]&~m[107])|(m[0]&m[104]&~m[105]&~m[106]&m[107])|(m[0]&~m[104]&m[105]&~m[106]&m[107])|(~m[0]&m[104]&m[105]&~m[106]&m[107])|(m[0]&~m[104]&~m[105]&m[106]&m[107])|(~m[0]&m[104]&~m[105]&m[106]&m[107])|(~m[0]&~m[104]&m[105]&m[106]&m[107]))&~BiasedRNG[170])|((m[0]&m[104]&m[105]&m[106]&~m[107])|(m[0]&m[104]&m[105]&~m[106]&m[107])|(m[0]&m[104]&~m[105]&m[106]&m[107])|(m[0]&~m[104]&m[105]&m[106]&m[107])|(~m[0]&m[104]&m[105]&m[106]&m[107])|(m[0]&m[104]&m[105]&m[106]&m[107]));
    m[27] = (((m[1]&m[108]&~m[109]&~m[110]&~m[111])|(m[1]&~m[108]&m[109]&~m[110]&~m[111])|(~m[1]&m[108]&m[109]&~m[110]&~m[111])|(m[1]&~m[108]&~m[109]&m[110]&~m[111])|(~m[1]&m[108]&~m[109]&m[110]&~m[111])|(~m[1]&~m[108]&m[109]&m[110]&~m[111])|(m[1]&~m[108]&~m[109]&~m[110]&m[111])|(~m[1]&m[108]&~m[109]&~m[110]&m[111])|(~m[1]&~m[108]&m[109]&~m[110]&m[111])|(~m[1]&~m[108]&~m[109]&m[110]&m[111]))&BiasedRNG[171])|(((m[1]&m[108]&m[109]&~m[110]&~m[111])|(m[1]&m[108]&~m[109]&m[110]&~m[111])|(m[1]&~m[108]&m[109]&m[110]&~m[111])|(~m[1]&m[108]&m[109]&m[110]&~m[111])|(m[1]&m[108]&~m[109]&~m[110]&m[111])|(m[1]&~m[108]&m[109]&~m[110]&m[111])|(~m[1]&m[108]&m[109]&~m[110]&m[111])|(m[1]&~m[108]&~m[109]&m[110]&m[111])|(~m[1]&m[108]&~m[109]&m[110]&m[111])|(~m[1]&~m[108]&m[109]&m[110]&m[111]))&~BiasedRNG[171])|((m[1]&m[108]&m[109]&m[110]&~m[111])|(m[1]&m[108]&m[109]&~m[110]&m[111])|(m[1]&m[108]&~m[109]&m[110]&m[111])|(m[1]&~m[108]&m[109]&m[110]&m[111])|(~m[1]&m[108]&m[109]&m[110]&m[111])|(m[1]&m[108]&m[109]&m[110]&m[111]));
    m[28] = (((m[1]&m[112]&~m[113]&~m[114]&~m[115])|(m[1]&~m[112]&m[113]&~m[114]&~m[115])|(~m[1]&m[112]&m[113]&~m[114]&~m[115])|(m[1]&~m[112]&~m[113]&m[114]&~m[115])|(~m[1]&m[112]&~m[113]&m[114]&~m[115])|(~m[1]&~m[112]&m[113]&m[114]&~m[115])|(m[1]&~m[112]&~m[113]&~m[114]&m[115])|(~m[1]&m[112]&~m[113]&~m[114]&m[115])|(~m[1]&~m[112]&m[113]&~m[114]&m[115])|(~m[1]&~m[112]&~m[113]&m[114]&m[115]))&BiasedRNG[172])|(((m[1]&m[112]&m[113]&~m[114]&~m[115])|(m[1]&m[112]&~m[113]&m[114]&~m[115])|(m[1]&~m[112]&m[113]&m[114]&~m[115])|(~m[1]&m[112]&m[113]&m[114]&~m[115])|(m[1]&m[112]&~m[113]&~m[114]&m[115])|(m[1]&~m[112]&m[113]&~m[114]&m[115])|(~m[1]&m[112]&m[113]&~m[114]&m[115])|(m[1]&~m[112]&~m[113]&m[114]&m[115])|(~m[1]&m[112]&~m[113]&m[114]&m[115])|(~m[1]&~m[112]&m[113]&m[114]&m[115]))&~BiasedRNG[172])|((m[1]&m[112]&m[113]&m[114]&~m[115])|(m[1]&m[112]&m[113]&~m[114]&m[115])|(m[1]&m[112]&~m[113]&m[114]&m[115])|(m[1]&~m[112]&m[113]&m[114]&m[115])|(~m[1]&m[112]&m[113]&m[114]&m[115])|(m[1]&m[112]&m[113]&m[114]&m[115]));
    m[29] = (((m[1]&m[116]&~m[117]&~m[118]&~m[119])|(m[1]&~m[116]&m[117]&~m[118]&~m[119])|(~m[1]&m[116]&m[117]&~m[118]&~m[119])|(m[1]&~m[116]&~m[117]&m[118]&~m[119])|(~m[1]&m[116]&~m[117]&m[118]&~m[119])|(~m[1]&~m[116]&m[117]&m[118]&~m[119])|(m[1]&~m[116]&~m[117]&~m[118]&m[119])|(~m[1]&m[116]&~m[117]&~m[118]&m[119])|(~m[1]&~m[116]&m[117]&~m[118]&m[119])|(~m[1]&~m[116]&~m[117]&m[118]&m[119]))&BiasedRNG[173])|(((m[1]&m[116]&m[117]&~m[118]&~m[119])|(m[1]&m[116]&~m[117]&m[118]&~m[119])|(m[1]&~m[116]&m[117]&m[118]&~m[119])|(~m[1]&m[116]&m[117]&m[118]&~m[119])|(m[1]&m[116]&~m[117]&~m[118]&m[119])|(m[1]&~m[116]&m[117]&~m[118]&m[119])|(~m[1]&m[116]&m[117]&~m[118]&m[119])|(m[1]&~m[116]&~m[117]&m[118]&m[119])|(~m[1]&m[116]&~m[117]&m[118]&m[119])|(~m[1]&~m[116]&m[117]&m[118]&m[119]))&~BiasedRNG[173])|((m[1]&m[116]&m[117]&m[118]&~m[119])|(m[1]&m[116]&m[117]&~m[118]&m[119])|(m[1]&m[116]&~m[117]&m[118]&m[119])|(m[1]&~m[116]&m[117]&m[118]&m[119])|(~m[1]&m[116]&m[117]&m[118]&m[119])|(m[1]&m[116]&m[117]&m[118]&m[119]));
    m[30] = (((m[2]&m[120]&~m[121]&~m[122]&~m[123])|(m[2]&~m[120]&m[121]&~m[122]&~m[123])|(~m[2]&m[120]&m[121]&~m[122]&~m[123])|(m[2]&~m[120]&~m[121]&m[122]&~m[123])|(~m[2]&m[120]&~m[121]&m[122]&~m[123])|(~m[2]&~m[120]&m[121]&m[122]&~m[123])|(m[2]&~m[120]&~m[121]&~m[122]&m[123])|(~m[2]&m[120]&~m[121]&~m[122]&m[123])|(~m[2]&~m[120]&m[121]&~m[122]&m[123])|(~m[2]&~m[120]&~m[121]&m[122]&m[123]))&BiasedRNG[174])|(((m[2]&m[120]&m[121]&~m[122]&~m[123])|(m[2]&m[120]&~m[121]&m[122]&~m[123])|(m[2]&~m[120]&m[121]&m[122]&~m[123])|(~m[2]&m[120]&m[121]&m[122]&~m[123])|(m[2]&m[120]&~m[121]&~m[122]&m[123])|(m[2]&~m[120]&m[121]&~m[122]&m[123])|(~m[2]&m[120]&m[121]&~m[122]&m[123])|(m[2]&~m[120]&~m[121]&m[122]&m[123])|(~m[2]&m[120]&~m[121]&m[122]&m[123])|(~m[2]&~m[120]&m[121]&m[122]&m[123]))&~BiasedRNG[174])|((m[2]&m[120]&m[121]&m[122]&~m[123])|(m[2]&m[120]&m[121]&~m[122]&m[123])|(m[2]&m[120]&~m[121]&m[122]&m[123])|(m[2]&~m[120]&m[121]&m[122]&m[123])|(~m[2]&m[120]&m[121]&m[122]&m[123])|(m[2]&m[120]&m[121]&m[122]&m[123]));
    m[31] = (((m[2]&m[124]&~m[125]&~m[126]&~m[127])|(m[2]&~m[124]&m[125]&~m[126]&~m[127])|(~m[2]&m[124]&m[125]&~m[126]&~m[127])|(m[2]&~m[124]&~m[125]&m[126]&~m[127])|(~m[2]&m[124]&~m[125]&m[126]&~m[127])|(~m[2]&~m[124]&m[125]&m[126]&~m[127])|(m[2]&~m[124]&~m[125]&~m[126]&m[127])|(~m[2]&m[124]&~m[125]&~m[126]&m[127])|(~m[2]&~m[124]&m[125]&~m[126]&m[127])|(~m[2]&~m[124]&~m[125]&m[126]&m[127]))&BiasedRNG[175])|(((m[2]&m[124]&m[125]&~m[126]&~m[127])|(m[2]&m[124]&~m[125]&m[126]&~m[127])|(m[2]&~m[124]&m[125]&m[126]&~m[127])|(~m[2]&m[124]&m[125]&m[126]&~m[127])|(m[2]&m[124]&~m[125]&~m[126]&m[127])|(m[2]&~m[124]&m[125]&~m[126]&m[127])|(~m[2]&m[124]&m[125]&~m[126]&m[127])|(m[2]&~m[124]&~m[125]&m[126]&m[127])|(~m[2]&m[124]&~m[125]&m[126]&m[127])|(~m[2]&~m[124]&m[125]&m[126]&m[127]))&~BiasedRNG[175])|((m[2]&m[124]&m[125]&m[126]&~m[127])|(m[2]&m[124]&m[125]&~m[126]&m[127])|(m[2]&m[124]&~m[125]&m[126]&m[127])|(m[2]&~m[124]&m[125]&m[126]&m[127])|(~m[2]&m[124]&m[125]&m[126]&m[127])|(m[2]&m[124]&m[125]&m[126]&m[127]));
    m[32] = (((m[2]&m[128]&~m[129]&~m[130]&~m[131])|(m[2]&~m[128]&m[129]&~m[130]&~m[131])|(~m[2]&m[128]&m[129]&~m[130]&~m[131])|(m[2]&~m[128]&~m[129]&m[130]&~m[131])|(~m[2]&m[128]&~m[129]&m[130]&~m[131])|(~m[2]&~m[128]&m[129]&m[130]&~m[131])|(m[2]&~m[128]&~m[129]&~m[130]&m[131])|(~m[2]&m[128]&~m[129]&~m[130]&m[131])|(~m[2]&~m[128]&m[129]&~m[130]&m[131])|(~m[2]&~m[128]&~m[129]&m[130]&m[131]))&BiasedRNG[176])|(((m[2]&m[128]&m[129]&~m[130]&~m[131])|(m[2]&m[128]&~m[129]&m[130]&~m[131])|(m[2]&~m[128]&m[129]&m[130]&~m[131])|(~m[2]&m[128]&m[129]&m[130]&~m[131])|(m[2]&m[128]&~m[129]&~m[130]&m[131])|(m[2]&~m[128]&m[129]&~m[130]&m[131])|(~m[2]&m[128]&m[129]&~m[130]&m[131])|(m[2]&~m[128]&~m[129]&m[130]&m[131])|(~m[2]&m[128]&~m[129]&m[130]&m[131])|(~m[2]&~m[128]&m[129]&m[130]&m[131]))&~BiasedRNG[176])|((m[2]&m[128]&m[129]&m[130]&~m[131])|(m[2]&m[128]&m[129]&~m[130]&m[131])|(m[2]&m[128]&~m[129]&m[130]&m[131])|(m[2]&~m[128]&m[129]&m[130]&m[131])|(~m[2]&m[128]&m[129]&m[130]&m[131])|(m[2]&m[128]&m[129]&m[130]&m[131]));
    m[33] = (((m[3]&m[132]&~m[133]&~m[134]&~m[135])|(m[3]&~m[132]&m[133]&~m[134]&~m[135])|(~m[3]&m[132]&m[133]&~m[134]&~m[135])|(m[3]&~m[132]&~m[133]&m[134]&~m[135])|(~m[3]&m[132]&~m[133]&m[134]&~m[135])|(~m[3]&~m[132]&m[133]&m[134]&~m[135])|(m[3]&~m[132]&~m[133]&~m[134]&m[135])|(~m[3]&m[132]&~m[133]&~m[134]&m[135])|(~m[3]&~m[132]&m[133]&~m[134]&m[135])|(~m[3]&~m[132]&~m[133]&m[134]&m[135]))&BiasedRNG[177])|(((m[3]&m[132]&m[133]&~m[134]&~m[135])|(m[3]&m[132]&~m[133]&m[134]&~m[135])|(m[3]&~m[132]&m[133]&m[134]&~m[135])|(~m[3]&m[132]&m[133]&m[134]&~m[135])|(m[3]&m[132]&~m[133]&~m[134]&m[135])|(m[3]&~m[132]&m[133]&~m[134]&m[135])|(~m[3]&m[132]&m[133]&~m[134]&m[135])|(m[3]&~m[132]&~m[133]&m[134]&m[135])|(~m[3]&m[132]&~m[133]&m[134]&m[135])|(~m[3]&~m[132]&m[133]&m[134]&m[135]))&~BiasedRNG[177])|((m[3]&m[132]&m[133]&m[134]&~m[135])|(m[3]&m[132]&m[133]&~m[134]&m[135])|(m[3]&m[132]&~m[133]&m[134]&m[135])|(m[3]&~m[132]&m[133]&m[134]&m[135])|(~m[3]&m[132]&m[133]&m[134]&m[135])|(m[3]&m[132]&m[133]&m[134]&m[135]));
    m[34] = (((m[3]&m[136]&~m[137]&~m[138]&~m[139])|(m[3]&~m[136]&m[137]&~m[138]&~m[139])|(~m[3]&m[136]&m[137]&~m[138]&~m[139])|(m[3]&~m[136]&~m[137]&m[138]&~m[139])|(~m[3]&m[136]&~m[137]&m[138]&~m[139])|(~m[3]&~m[136]&m[137]&m[138]&~m[139])|(m[3]&~m[136]&~m[137]&~m[138]&m[139])|(~m[3]&m[136]&~m[137]&~m[138]&m[139])|(~m[3]&~m[136]&m[137]&~m[138]&m[139])|(~m[3]&~m[136]&~m[137]&m[138]&m[139]))&BiasedRNG[178])|(((m[3]&m[136]&m[137]&~m[138]&~m[139])|(m[3]&m[136]&~m[137]&m[138]&~m[139])|(m[3]&~m[136]&m[137]&m[138]&~m[139])|(~m[3]&m[136]&m[137]&m[138]&~m[139])|(m[3]&m[136]&~m[137]&~m[138]&m[139])|(m[3]&~m[136]&m[137]&~m[138]&m[139])|(~m[3]&m[136]&m[137]&~m[138]&m[139])|(m[3]&~m[136]&~m[137]&m[138]&m[139])|(~m[3]&m[136]&~m[137]&m[138]&m[139])|(~m[3]&~m[136]&m[137]&m[138]&m[139]))&~BiasedRNG[178])|((m[3]&m[136]&m[137]&m[138]&~m[139])|(m[3]&m[136]&m[137]&~m[138]&m[139])|(m[3]&m[136]&~m[137]&m[138]&m[139])|(m[3]&~m[136]&m[137]&m[138]&m[139])|(~m[3]&m[136]&m[137]&m[138]&m[139])|(m[3]&m[136]&m[137]&m[138]&m[139]));
    m[35] = (((m[3]&m[140]&~m[141]&~m[142]&~m[143])|(m[3]&~m[140]&m[141]&~m[142]&~m[143])|(~m[3]&m[140]&m[141]&~m[142]&~m[143])|(m[3]&~m[140]&~m[141]&m[142]&~m[143])|(~m[3]&m[140]&~m[141]&m[142]&~m[143])|(~m[3]&~m[140]&m[141]&m[142]&~m[143])|(m[3]&~m[140]&~m[141]&~m[142]&m[143])|(~m[3]&m[140]&~m[141]&~m[142]&m[143])|(~m[3]&~m[140]&m[141]&~m[142]&m[143])|(~m[3]&~m[140]&~m[141]&m[142]&m[143]))&BiasedRNG[179])|(((m[3]&m[140]&m[141]&~m[142]&~m[143])|(m[3]&m[140]&~m[141]&m[142]&~m[143])|(m[3]&~m[140]&m[141]&m[142]&~m[143])|(~m[3]&m[140]&m[141]&m[142]&~m[143])|(m[3]&m[140]&~m[141]&~m[142]&m[143])|(m[3]&~m[140]&m[141]&~m[142]&m[143])|(~m[3]&m[140]&m[141]&~m[142]&m[143])|(m[3]&~m[140]&~m[141]&m[142]&m[143])|(~m[3]&m[140]&~m[141]&m[142]&m[143])|(~m[3]&~m[140]&m[141]&m[142]&m[143]))&~BiasedRNG[179])|((m[3]&m[140]&m[141]&m[142]&~m[143])|(m[3]&m[140]&m[141]&~m[142]&m[143])|(m[3]&m[140]&~m[141]&m[142]&m[143])|(m[3]&~m[140]&m[141]&m[142]&m[143])|(~m[3]&m[140]&m[141]&m[142]&m[143])|(m[3]&m[140]&m[141]&m[142]&m[143]));
    m[36] = (((m[4]&m[144]&~m[145]&~m[146]&~m[147])|(m[4]&~m[144]&m[145]&~m[146]&~m[147])|(~m[4]&m[144]&m[145]&~m[146]&~m[147])|(m[4]&~m[144]&~m[145]&m[146]&~m[147])|(~m[4]&m[144]&~m[145]&m[146]&~m[147])|(~m[4]&~m[144]&m[145]&m[146]&~m[147])|(m[4]&~m[144]&~m[145]&~m[146]&m[147])|(~m[4]&m[144]&~m[145]&~m[146]&m[147])|(~m[4]&~m[144]&m[145]&~m[146]&m[147])|(~m[4]&~m[144]&~m[145]&m[146]&m[147]))&BiasedRNG[180])|(((m[4]&m[144]&m[145]&~m[146]&~m[147])|(m[4]&m[144]&~m[145]&m[146]&~m[147])|(m[4]&~m[144]&m[145]&m[146]&~m[147])|(~m[4]&m[144]&m[145]&m[146]&~m[147])|(m[4]&m[144]&~m[145]&~m[146]&m[147])|(m[4]&~m[144]&m[145]&~m[146]&m[147])|(~m[4]&m[144]&m[145]&~m[146]&m[147])|(m[4]&~m[144]&~m[145]&m[146]&m[147])|(~m[4]&m[144]&~m[145]&m[146]&m[147])|(~m[4]&~m[144]&m[145]&m[146]&m[147]))&~BiasedRNG[180])|((m[4]&m[144]&m[145]&m[146]&~m[147])|(m[4]&m[144]&m[145]&~m[146]&m[147])|(m[4]&m[144]&~m[145]&m[146]&m[147])|(m[4]&~m[144]&m[145]&m[146]&m[147])|(~m[4]&m[144]&m[145]&m[146]&m[147])|(m[4]&m[144]&m[145]&m[146]&m[147]));
    m[37] = (((m[4]&m[148]&~m[149]&~m[150]&~m[151])|(m[4]&~m[148]&m[149]&~m[150]&~m[151])|(~m[4]&m[148]&m[149]&~m[150]&~m[151])|(m[4]&~m[148]&~m[149]&m[150]&~m[151])|(~m[4]&m[148]&~m[149]&m[150]&~m[151])|(~m[4]&~m[148]&m[149]&m[150]&~m[151])|(m[4]&~m[148]&~m[149]&~m[150]&m[151])|(~m[4]&m[148]&~m[149]&~m[150]&m[151])|(~m[4]&~m[148]&m[149]&~m[150]&m[151])|(~m[4]&~m[148]&~m[149]&m[150]&m[151]))&BiasedRNG[181])|(((m[4]&m[148]&m[149]&~m[150]&~m[151])|(m[4]&m[148]&~m[149]&m[150]&~m[151])|(m[4]&~m[148]&m[149]&m[150]&~m[151])|(~m[4]&m[148]&m[149]&m[150]&~m[151])|(m[4]&m[148]&~m[149]&~m[150]&m[151])|(m[4]&~m[148]&m[149]&~m[150]&m[151])|(~m[4]&m[148]&m[149]&~m[150]&m[151])|(m[4]&~m[148]&~m[149]&m[150]&m[151])|(~m[4]&m[148]&~m[149]&m[150]&m[151])|(~m[4]&~m[148]&m[149]&m[150]&m[151]))&~BiasedRNG[181])|((m[4]&m[148]&m[149]&m[150]&~m[151])|(m[4]&m[148]&m[149]&~m[150]&m[151])|(m[4]&m[148]&~m[149]&m[150]&m[151])|(m[4]&~m[148]&m[149]&m[150]&m[151])|(~m[4]&m[148]&m[149]&m[150]&m[151])|(m[4]&m[148]&m[149]&m[150]&m[151]));
    m[38] = (((m[4]&m[152]&~m[153]&~m[154]&~m[155])|(m[4]&~m[152]&m[153]&~m[154]&~m[155])|(~m[4]&m[152]&m[153]&~m[154]&~m[155])|(m[4]&~m[152]&~m[153]&m[154]&~m[155])|(~m[4]&m[152]&~m[153]&m[154]&~m[155])|(~m[4]&~m[152]&m[153]&m[154]&~m[155])|(m[4]&~m[152]&~m[153]&~m[154]&m[155])|(~m[4]&m[152]&~m[153]&~m[154]&m[155])|(~m[4]&~m[152]&m[153]&~m[154]&m[155])|(~m[4]&~m[152]&~m[153]&m[154]&m[155]))&BiasedRNG[182])|(((m[4]&m[152]&m[153]&~m[154]&~m[155])|(m[4]&m[152]&~m[153]&m[154]&~m[155])|(m[4]&~m[152]&m[153]&m[154]&~m[155])|(~m[4]&m[152]&m[153]&m[154]&~m[155])|(m[4]&m[152]&~m[153]&~m[154]&m[155])|(m[4]&~m[152]&m[153]&~m[154]&m[155])|(~m[4]&m[152]&m[153]&~m[154]&m[155])|(m[4]&~m[152]&~m[153]&m[154]&m[155])|(~m[4]&m[152]&~m[153]&m[154]&m[155])|(~m[4]&~m[152]&m[153]&m[154]&m[155]))&~BiasedRNG[182])|((m[4]&m[152]&m[153]&m[154]&~m[155])|(m[4]&m[152]&m[153]&~m[154]&m[155])|(m[4]&m[152]&~m[153]&m[154]&m[155])|(m[4]&~m[152]&m[153]&m[154]&m[155])|(~m[4]&m[152]&m[153]&m[154]&m[155])|(m[4]&m[152]&m[153]&m[154]&m[155]));
    m[39] = (((m[5]&m[156]&~m[157]&~m[158]&~m[159])|(m[5]&~m[156]&m[157]&~m[158]&~m[159])|(~m[5]&m[156]&m[157]&~m[158]&~m[159])|(m[5]&~m[156]&~m[157]&m[158]&~m[159])|(~m[5]&m[156]&~m[157]&m[158]&~m[159])|(~m[5]&~m[156]&m[157]&m[158]&~m[159])|(m[5]&~m[156]&~m[157]&~m[158]&m[159])|(~m[5]&m[156]&~m[157]&~m[158]&m[159])|(~m[5]&~m[156]&m[157]&~m[158]&m[159])|(~m[5]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[183])|(((m[5]&m[156]&m[157]&~m[158]&~m[159])|(m[5]&m[156]&~m[157]&m[158]&~m[159])|(m[5]&~m[156]&m[157]&m[158]&~m[159])|(~m[5]&m[156]&m[157]&m[158]&~m[159])|(m[5]&m[156]&~m[157]&~m[158]&m[159])|(m[5]&~m[156]&m[157]&~m[158]&m[159])|(~m[5]&m[156]&m[157]&~m[158]&m[159])|(m[5]&~m[156]&~m[157]&m[158]&m[159])|(~m[5]&m[156]&~m[157]&m[158]&m[159])|(~m[5]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[183])|((m[5]&m[156]&m[157]&m[158]&~m[159])|(m[5]&m[156]&m[157]&~m[158]&m[159])|(m[5]&m[156]&~m[157]&m[158]&m[159])|(m[5]&~m[156]&m[157]&m[158]&m[159])|(~m[5]&m[156]&m[157]&m[158]&m[159])|(m[5]&m[156]&m[157]&m[158]&m[159]));
    m[40] = (((m[5]&m[160]&~m[161]&~m[162]&~m[163])|(m[5]&~m[160]&m[161]&~m[162]&~m[163])|(~m[5]&m[160]&m[161]&~m[162]&~m[163])|(m[5]&~m[160]&~m[161]&m[162]&~m[163])|(~m[5]&m[160]&~m[161]&m[162]&~m[163])|(~m[5]&~m[160]&m[161]&m[162]&~m[163])|(m[5]&~m[160]&~m[161]&~m[162]&m[163])|(~m[5]&m[160]&~m[161]&~m[162]&m[163])|(~m[5]&~m[160]&m[161]&~m[162]&m[163])|(~m[5]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[184])|(((m[5]&m[160]&m[161]&~m[162]&~m[163])|(m[5]&m[160]&~m[161]&m[162]&~m[163])|(m[5]&~m[160]&m[161]&m[162]&~m[163])|(~m[5]&m[160]&m[161]&m[162]&~m[163])|(m[5]&m[160]&~m[161]&~m[162]&m[163])|(m[5]&~m[160]&m[161]&~m[162]&m[163])|(~m[5]&m[160]&m[161]&~m[162]&m[163])|(m[5]&~m[160]&~m[161]&m[162]&m[163])|(~m[5]&m[160]&~m[161]&m[162]&m[163])|(~m[5]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[184])|((m[5]&m[160]&m[161]&m[162]&~m[163])|(m[5]&m[160]&m[161]&~m[162]&m[163])|(m[5]&m[160]&~m[161]&m[162]&m[163])|(m[5]&~m[160]&m[161]&m[162]&m[163])|(~m[5]&m[160]&m[161]&m[162]&m[163])|(m[5]&m[160]&m[161]&m[162]&m[163]));
    m[41] = (((m[5]&m[164]&~m[165]&~m[166]&~m[167])|(m[5]&~m[164]&m[165]&~m[166]&~m[167])|(~m[5]&m[164]&m[165]&~m[166]&~m[167])|(m[5]&~m[164]&~m[165]&m[166]&~m[167])|(~m[5]&m[164]&~m[165]&m[166]&~m[167])|(~m[5]&~m[164]&m[165]&m[166]&~m[167])|(m[5]&~m[164]&~m[165]&~m[166]&m[167])|(~m[5]&m[164]&~m[165]&~m[166]&m[167])|(~m[5]&~m[164]&m[165]&~m[166]&m[167])|(~m[5]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[185])|(((m[5]&m[164]&m[165]&~m[166]&~m[167])|(m[5]&m[164]&~m[165]&m[166]&~m[167])|(m[5]&~m[164]&m[165]&m[166]&~m[167])|(~m[5]&m[164]&m[165]&m[166]&~m[167])|(m[5]&m[164]&~m[165]&~m[166]&m[167])|(m[5]&~m[164]&m[165]&~m[166]&m[167])|(~m[5]&m[164]&m[165]&~m[166]&m[167])|(m[5]&~m[164]&~m[165]&m[166]&m[167])|(~m[5]&m[164]&~m[165]&m[166]&m[167])|(~m[5]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[185])|((m[5]&m[164]&m[165]&m[166]&~m[167])|(m[5]&m[164]&m[165]&~m[166]&m[167])|(m[5]&m[164]&~m[165]&m[166]&m[167])|(m[5]&~m[164]&m[165]&m[166]&m[167])|(~m[5]&m[164]&m[165]&m[166]&m[167])|(m[5]&m[164]&m[165]&m[166]&m[167]));
    m[42] = (((m[6]&m[168]&~m[169]&~m[170]&~m[171])|(m[6]&~m[168]&m[169]&~m[170]&~m[171])|(~m[6]&m[168]&m[169]&~m[170]&~m[171])|(m[6]&~m[168]&~m[169]&m[170]&~m[171])|(~m[6]&m[168]&~m[169]&m[170]&~m[171])|(~m[6]&~m[168]&m[169]&m[170]&~m[171])|(m[6]&~m[168]&~m[169]&~m[170]&m[171])|(~m[6]&m[168]&~m[169]&~m[170]&m[171])|(~m[6]&~m[168]&m[169]&~m[170]&m[171])|(~m[6]&~m[168]&~m[169]&m[170]&m[171]))&BiasedRNG[186])|(((m[6]&m[168]&m[169]&~m[170]&~m[171])|(m[6]&m[168]&~m[169]&m[170]&~m[171])|(m[6]&~m[168]&m[169]&m[170]&~m[171])|(~m[6]&m[168]&m[169]&m[170]&~m[171])|(m[6]&m[168]&~m[169]&~m[170]&m[171])|(m[6]&~m[168]&m[169]&~m[170]&m[171])|(~m[6]&m[168]&m[169]&~m[170]&m[171])|(m[6]&~m[168]&~m[169]&m[170]&m[171])|(~m[6]&m[168]&~m[169]&m[170]&m[171])|(~m[6]&~m[168]&m[169]&m[170]&m[171]))&~BiasedRNG[186])|((m[6]&m[168]&m[169]&m[170]&~m[171])|(m[6]&m[168]&m[169]&~m[170]&m[171])|(m[6]&m[168]&~m[169]&m[170]&m[171])|(m[6]&~m[168]&m[169]&m[170]&m[171])|(~m[6]&m[168]&m[169]&m[170]&m[171])|(m[6]&m[168]&m[169]&m[170]&m[171]));
    m[43] = (((m[6]&m[172]&~m[173]&~m[174]&~m[175])|(m[6]&~m[172]&m[173]&~m[174]&~m[175])|(~m[6]&m[172]&m[173]&~m[174]&~m[175])|(m[6]&~m[172]&~m[173]&m[174]&~m[175])|(~m[6]&m[172]&~m[173]&m[174]&~m[175])|(~m[6]&~m[172]&m[173]&m[174]&~m[175])|(m[6]&~m[172]&~m[173]&~m[174]&m[175])|(~m[6]&m[172]&~m[173]&~m[174]&m[175])|(~m[6]&~m[172]&m[173]&~m[174]&m[175])|(~m[6]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[187])|(((m[6]&m[172]&m[173]&~m[174]&~m[175])|(m[6]&m[172]&~m[173]&m[174]&~m[175])|(m[6]&~m[172]&m[173]&m[174]&~m[175])|(~m[6]&m[172]&m[173]&m[174]&~m[175])|(m[6]&m[172]&~m[173]&~m[174]&m[175])|(m[6]&~m[172]&m[173]&~m[174]&m[175])|(~m[6]&m[172]&m[173]&~m[174]&m[175])|(m[6]&~m[172]&~m[173]&m[174]&m[175])|(~m[6]&m[172]&~m[173]&m[174]&m[175])|(~m[6]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[187])|((m[6]&m[172]&m[173]&m[174]&~m[175])|(m[6]&m[172]&m[173]&~m[174]&m[175])|(m[6]&m[172]&~m[173]&m[174]&m[175])|(m[6]&~m[172]&m[173]&m[174]&m[175])|(~m[6]&m[172]&m[173]&m[174]&m[175])|(m[6]&m[172]&m[173]&m[174]&m[175]));
    m[44] = (((m[6]&m[176]&~m[177]&~m[178]&~m[179])|(m[6]&~m[176]&m[177]&~m[178]&~m[179])|(~m[6]&m[176]&m[177]&~m[178]&~m[179])|(m[6]&~m[176]&~m[177]&m[178]&~m[179])|(~m[6]&m[176]&~m[177]&m[178]&~m[179])|(~m[6]&~m[176]&m[177]&m[178]&~m[179])|(m[6]&~m[176]&~m[177]&~m[178]&m[179])|(~m[6]&m[176]&~m[177]&~m[178]&m[179])|(~m[6]&~m[176]&m[177]&~m[178]&m[179])|(~m[6]&~m[176]&~m[177]&m[178]&m[179]))&BiasedRNG[188])|(((m[6]&m[176]&m[177]&~m[178]&~m[179])|(m[6]&m[176]&~m[177]&m[178]&~m[179])|(m[6]&~m[176]&m[177]&m[178]&~m[179])|(~m[6]&m[176]&m[177]&m[178]&~m[179])|(m[6]&m[176]&~m[177]&~m[178]&m[179])|(m[6]&~m[176]&m[177]&~m[178]&m[179])|(~m[6]&m[176]&m[177]&~m[178]&m[179])|(m[6]&~m[176]&~m[177]&m[178]&m[179])|(~m[6]&m[176]&~m[177]&m[178]&m[179])|(~m[6]&~m[176]&m[177]&m[178]&m[179]))&~BiasedRNG[188])|((m[6]&m[176]&m[177]&m[178]&~m[179])|(m[6]&m[176]&m[177]&~m[178]&m[179])|(m[6]&m[176]&~m[177]&m[178]&m[179])|(m[6]&~m[176]&m[177]&m[178]&m[179])|(~m[6]&m[176]&m[177]&m[178]&m[179])|(m[6]&m[176]&m[177]&m[178]&m[179]));
    m[45] = (((m[7]&m[180]&~m[181]&~m[182]&~m[183])|(m[7]&~m[180]&m[181]&~m[182]&~m[183])|(~m[7]&m[180]&m[181]&~m[182]&~m[183])|(m[7]&~m[180]&~m[181]&m[182]&~m[183])|(~m[7]&m[180]&~m[181]&m[182]&~m[183])|(~m[7]&~m[180]&m[181]&m[182]&~m[183])|(m[7]&~m[180]&~m[181]&~m[182]&m[183])|(~m[7]&m[180]&~m[181]&~m[182]&m[183])|(~m[7]&~m[180]&m[181]&~m[182]&m[183])|(~m[7]&~m[180]&~m[181]&m[182]&m[183]))&BiasedRNG[189])|(((m[7]&m[180]&m[181]&~m[182]&~m[183])|(m[7]&m[180]&~m[181]&m[182]&~m[183])|(m[7]&~m[180]&m[181]&m[182]&~m[183])|(~m[7]&m[180]&m[181]&m[182]&~m[183])|(m[7]&m[180]&~m[181]&~m[182]&m[183])|(m[7]&~m[180]&m[181]&~m[182]&m[183])|(~m[7]&m[180]&m[181]&~m[182]&m[183])|(m[7]&~m[180]&~m[181]&m[182]&m[183])|(~m[7]&m[180]&~m[181]&m[182]&m[183])|(~m[7]&~m[180]&m[181]&m[182]&m[183]))&~BiasedRNG[189])|((m[7]&m[180]&m[181]&m[182]&~m[183])|(m[7]&m[180]&m[181]&~m[182]&m[183])|(m[7]&m[180]&~m[181]&m[182]&m[183])|(m[7]&~m[180]&m[181]&m[182]&m[183])|(~m[7]&m[180]&m[181]&m[182]&m[183])|(m[7]&m[180]&m[181]&m[182]&m[183]));
    m[46] = (((m[7]&m[184]&~m[185]&~m[186]&~m[187])|(m[7]&~m[184]&m[185]&~m[186]&~m[187])|(~m[7]&m[184]&m[185]&~m[186]&~m[187])|(m[7]&~m[184]&~m[185]&m[186]&~m[187])|(~m[7]&m[184]&~m[185]&m[186]&~m[187])|(~m[7]&~m[184]&m[185]&m[186]&~m[187])|(m[7]&~m[184]&~m[185]&~m[186]&m[187])|(~m[7]&m[184]&~m[185]&~m[186]&m[187])|(~m[7]&~m[184]&m[185]&~m[186]&m[187])|(~m[7]&~m[184]&~m[185]&m[186]&m[187]))&BiasedRNG[190])|(((m[7]&m[184]&m[185]&~m[186]&~m[187])|(m[7]&m[184]&~m[185]&m[186]&~m[187])|(m[7]&~m[184]&m[185]&m[186]&~m[187])|(~m[7]&m[184]&m[185]&m[186]&~m[187])|(m[7]&m[184]&~m[185]&~m[186]&m[187])|(m[7]&~m[184]&m[185]&~m[186]&m[187])|(~m[7]&m[184]&m[185]&~m[186]&m[187])|(m[7]&~m[184]&~m[185]&m[186]&m[187])|(~m[7]&m[184]&~m[185]&m[186]&m[187])|(~m[7]&~m[184]&m[185]&m[186]&m[187]))&~BiasedRNG[190])|((m[7]&m[184]&m[185]&m[186]&~m[187])|(m[7]&m[184]&m[185]&~m[186]&m[187])|(m[7]&m[184]&~m[185]&m[186]&m[187])|(m[7]&~m[184]&m[185]&m[186]&m[187])|(~m[7]&m[184]&m[185]&m[186]&m[187])|(m[7]&m[184]&m[185]&m[186]&m[187]));
    m[47] = (((m[7]&m[188]&~m[189]&~m[190]&~m[191])|(m[7]&~m[188]&m[189]&~m[190]&~m[191])|(~m[7]&m[188]&m[189]&~m[190]&~m[191])|(m[7]&~m[188]&~m[189]&m[190]&~m[191])|(~m[7]&m[188]&~m[189]&m[190]&~m[191])|(~m[7]&~m[188]&m[189]&m[190]&~m[191])|(m[7]&~m[188]&~m[189]&~m[190]&m[191])|(~m[7]&m[188]&~m[189]&~m[190]&m[191])|(~m[7]&~m[188]&m[189]&~m[190]&m[191])|(~m[7]&~m[188]&~m[189]&m[190]&m[191]))&BiasedRNG[191])|(((m[7]&m[188]&m[189]&~m[190]&~m[191])|(m[7]&m[188]&~m[189]&m[190]&~m[191])|(m[7]&~m[188]&m[189]&m[190]&~m[191])|(~m[7]&m[188]&m[189]&m[190]&~m[191])|(m[7]&m[188]&~m[189]&~m[190]&m[191])|(m[7]&~m[188]&m[189]&~m[190]&m[191])|(~m[7]&m[188]&m[189]&~m[190]&m[191])|(m[7]&~m[188]&~m[189]&m[190]&m[191])|(~m[7]&m[188]&~m[189]&m[190]&m[191])|(~m[7]&~m[188]&m[189]&m[190]&m[191]))&~BiasedRNG[191])|((m[7]&m[188]&m[189]&m[190]&~m[191])|(m[7]&m[188]&m[189]&~m[190]&m[191])|(m[7]&m[188]&~m[189]&m[190]&m[191])|(m[7]&~m[188]&m[189]&m[190]&m[191])|(~m[7]&m[188]&m[189]&m[190]&m[191])|(m[7]&m[188]&m[189]&m[190]&m[191]));
    m[48] = (((m[8]&m[192]&~m[193]&~m[194]&~m[195])|(m[8]&~m[192]&m[193]&~m[194]&~m[195])|(~m[8]&m[192]&m[193]&~m[194]&~m[195])|(m[8]&~m[192]&~m[193]&m[194]&~m[195])|(~m[8]&m[192]&~m[193]&m[194]&~m[195])|(~m[8]&~m[192]&m[193]&m[194]&~m[195])|(m[8]&~m[192]&~m[193]&~m[194]&m[195])|(~m[8]&m[192]&~m[193]&~m[194]&m[195])|(~m[8]&~m[192]&m[193]&~m[194]&m[195])|(~m[8]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[192])|(((m[8]&m[192]&m[193]&~m[194]&~m[195])|(m[8]&m[192]&~m[193]&m[194]&~m[195])|(m[8]&~m[192]&m[193]&m[194]&~m[195])|(~m[8]&m[192]&m[193]&m[194]&~m[195])|(m[8]&m[192]&~m[193]&~m[194]&m[195])|(m[8]&~m[192]&m[193]&~m[194]&m[195])|(~m[8]&m[192]&m[193]&~m[194]&m[195])|(m[8]&~m[192]&~m[193]&m[194]&m[195])|(~m[8]&m[192]&~m[193]&m[194]&m[195])|(~m[8]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[192])|((m[8]&m[192]&m[193]&m[194]&~m[195])|(m[8]&m[192]&m[193]&~m[194]&m[195])|(m[8]&m[192]&~m[193]&m[194]&m[195])|(m[8]&~m[192]&m[193]&m[194]&m[195])|(~m[8]&m[192]&m[193]&m[194]&m[195])|(m[8]&m[192]&m[193]&m[194]&m[195]));
    m[49] = (((m[8]&m[196]&~m[197]&~m[198]&~m[199])|(m[8]&~m[196]&m[197]&~m[198]&~m[199])|(~m[8]&m[196]&m[197]&~m[198]&~m[199])|(m[8]&~m[196]&~m[197]&m[198]&~m[199])|(~m[8]&m[196]&~m[197]&m[198]&~m[199])|(~m[8]&~m[196]&m[197]&m[198]&~m[199])|(m[8]&~m[196]&~m[197]&~m[198]&m[199])|(~m[8]&m[196]&~m[197]&~m[198]&m[199])|(~m[8]&~m[196]&m[197]&~m[198]&m[199])|(~m[8]&~m[196]&~m[197]&m[198]&m[199]))&BiasedRNG[193])|(((m[8]&m[196]&m[197]&~m[198]&~m[199])|(m[8]&m[196]&~m[197]&m[198]&~m[199])|(m[8]&~m[196]&m[197]&m[198]&~m[199])|(~m[8]&m[196]&m[197]&m[198]&~m[199])|(m[8]&m[196]&~m[197]&~m[198]&m[199])|(m[8]&~m[196]&m[197]&~m[198]&m[199])|(~m[8]&m[196]&m[197]&~m[198]&m[199])|(m[8]&~m[196]&~m[197]&m[198]&m[199])|(~m[8]&m[196]&~m[197]&m[198]&m[199])|(~m[8]&~m[196]&m[197]&m[198]&m[199]))&~BiasedRNG[193])|((m[8]&m[196]&m[197]&m[198]&~m[199])|(m[8]&m[196]&m[197]&~m[198]&m[199])|(m[8]&m[196]&~m[197]&m[198]&m[199])|(m[8]&~m[196]&m[197]&m[198]&m[199])|(~m[8]&m[196]&m[197]&m[198]&m[199])|(m[8]&m[196]&m[197]&m[198]&m[199]));
    m[50] = (((m[8]&m[200]&~m[201]&~m[202]&~m[203])|(m[8]&~m[200]&m[201]&~m[202]&~m[203])|(~m[8]&m[200]&m[201]&~m[202]&~m[203])|(m[8]&~m[200]&~m[201]&m[202]&~m[203])|(~m[8]&m[200]&~m[201]&m[202]&~m[203])|(~m[8]&~m[200]&m[201]&m[202]&~m[203])|(m[8]&~m[200]&~m[201]&~m[202]&m[203])|(~m[8]&m[200]&~m[201]&~m[202]&m[203])|(~m[8]&~m[200]&m[201]&~m[202]&m[203])|(~m[8]&~m[200]&~m[201]&m[202]&m[203]))&BiasedRNG[194])|(((m[8]&m[200]&m[201]&~m[202]&~m[203])|(m[8]&m[200]&~m[201]&m[202]&~m[203])|(m[8]&~m[200]&m[201]&m[202]&~m[203])|(~m[8]&m[200]&m[201]&m[202]&~m[203])|(m[8]&m[200]&~m[201]&~m[202]&m[203])|(m[8]&~m[200]&m[201]&~m[202]&m[203])|(~m[8]&m[200]&m[201]&~m[202]&m[203])|(m[8]&~m[200]&~m[201]&m[202]&m[203])|(~m[8]&m[200]&~m[201]&m[202]&m[203])|(~m[8]&~m[200]&m[201]&m[202]&m[203]))&~BiasedRNG[194])|((m[8]&m[200]&m[201]&m[202]&~m[203])|(m[8]&m[200]&m[201]&~m[202]&m[203])|(m[8]&m[200]&~m[201]&m[202]&m[203])|(m[8]&~m[200]&m[201]&m[202]&m[203])|(~m[8]&m[200]&m[201]&m[202]&m[203])|(m[8]&m[200]&m[201]&m[202]&m[203]));
    m[51] = (((m[9]&m[204]&~m[205]&~m[206]&~m[207])|(m[9]&~m[204]&m[205]&~m[206]&~m[207])|(~m[9]&m[204]&m[205]&~m[206]&~m[207])|(m[9]&~m[204]&~m[205]&m[206]&~m[207])|(~m[9]&m[204]&~m[205]&m[206]&~m[207])|(~m[9]&~m[204]&m[205]&m[206]&~m[207])|(m[9]&~m[204]&~m[205]&~m[206]&m[207])|(~m[9]&m[204]&~m[205]&~m[206]&m[207])|(~m[9]&~m[204]&m[205]&~m[206]&m[207])|(~m[9]&~m[204]&~m[205]&m[206]&m[207]))&BiasedRNG[195])|(((m[9]&m[204]&m[205]&~m[206]&~m[207])|(m[9]&m[204]&~m[205]&m[206]&~m[207])|(m[9]&~m[204]&m[205]&m[206]&~m[207])|(~m[9]&m[204]&m[205]&m[206]&~m[207])|(m[9]&m[204]&~m[205]&~m[206]&m[207])|(m[9]&~m[204]&m[205]&~m[206]&m[207])|(~m[9]&m[204]&m[205]&~m[206]&m[207])|(m[9]&~m[204]&~m[205]&m[206]&m[207])|(~m[9]&m[204]&~m[205]&m[206]&m[207])|(~m[9]&~m[204]&m[205]&m[206]&m[207]))&~BiasedRNG[195])|((m[9]&m[204]&m[205]&m[206]&~m[207])|(m[9]&m[204]&m[205]&~m[206]&m[207])|(m[9]&m[204]&~m[205]&m[206]&m[207])|(m[9]&~m[204]&m[205]&m[206]&m[207])|(~m[9]&m[204]&m[205]&m[206]&m[207])|(m[9]&m[204]&m[205]&m[206]&m[207]));
    m[52] = (((m[9]&m[208]&~m[209]&~m[210]&~m[211])|(m[9]&~m[208]&m[209]&~m[210]&~m[211])|(~m[9]&m[208]&m[209]&~m[210]&~m[211])|(m[9]&~m[208]&~m[209]&m[210]&~m[211])|(~m[9]&m[208]&~m[209]&m[210]&~m[211])|(~m[9]&~m[208]&m[209]&m[210]&~m[211])|(m[9]&~m[208]&~m[209]&~m[210]&m[211])|(~m[9]&m[208]&~m[209]&~m[210]&m[211])|(~m[9]&~m[208]&m[209]&~m[210]&m[211])|(~m[9]&~m[208]&~m[209]&m[210]&m[211]))&BiasedRNG[196])|(((m[9]&m[208]&m[209]&~m[210]&~m[211])|(m[9]&m[208]&~m[209]&m[210]&~m[211])|(m[9]&~m[208]&m[209]&m[210]&~m[211])|(~m[9]&m[208]&m[209]&m[210]&~m[211])|(m[9]&m[208]&~m[209]&~m[210]&m[211])|(m[9]&~m[208]&m[209]&~m[210]&m[211])|(~m[9]&m[208]&m[209]&~m[210]&m[211])|(m[9]&~m[208]&~m[209]&m[210]&m[211])|(~m[9]&m[208]&~m[209]&m[210]&m[211])|(~m[9]&~m[208]&m[209]&m[210]&m[211]))&~BiasedRNG[196])|((m[9]&m[208]&m[209]&m[210]&~m[211])|(m[9]&m[208]&m[209]&~m[210]&m[211])|(m[9]&m[208]&~m[209]&m[210]&m[211])|(m[9]&~m[208]&m[209]&m[210]&m[211])|(~m[9]&m[208]&m[209]&m[210]&m[211])|(m[9]&m[208]&m[209]&m[210]&m[211]));
    m[53] = (((m[9]&m[212]&~m[213]&~m[214]&~m[215])|(m[9]&~m[212]&m[213]&~m[214]&~m[215])|(~m[9]&m[212]&m[213]&~m[214]&~m[215])|(m[9]&~m[212]&~m[213]&m[214]&~m[215])|(~m[9]&m[212]&~m[213]&m[214]&~m[215])|(~m[9]&~m[212]&m[213]&m[214]&~m[215])|(m[9]&~m[212]&~m[213]&~m[214]&m[215])|(~m[9]&m[212]&~m[213]&~m[214]&m[215])|(~m[9]&~m[212]&m[213]&~m[214]&m[215])|(~m[9]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[197])|(((m[9]&m[212]&m[213]&~m[214]&~m[215])|(m[9]&m[212]&~m[213]&m[214]&~m[215])|(m[9]&~m[212]&m[213]&m[214]&~m[215])|(~m[9]&m[212]&m[213]&m[214]&~m[215])|(m[9]&m[212]&~m[213]&~m[214]&m[215])|(m[9]&~m[212]&m[213]&~m[214]&m[215])|(~m[9]&m[212]&m[213]&~m[214]&m[215])|(m[9]&~m[212]&~m[213]&m[214]&m[215])|(~m[9]&m[212]&~m[213]&m[214]&m[215])|(~m[9]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[197])|((m[9]&m[212]&m[213]&m[214]&~m[215])|(m[9]&m[212]&m[213]&~m[214]&m[215])|(m[9]&m[212]&~m[213]&m[214]&m[215])|(m[9]&~m[212]&m[213]&m[214]&m[215])|(~m[9]&m[212]&m[213]&m[214]&m[215])|(m[9]&m[212]&m[213]&m[214]&m[215]));
    m[54] = (((m[10]&m[216]&~m[217]&~m[218]&~m[219])|(m[10]&~m[216]&m[217]&~m[218]&~m[219])|(~m[10]&m[216]&m[217]&~m[218]&~m[219])|(m[10]&~m[216]&~m[217]&m[218]&~m[219])|(~m[10]&m[216]&~m[217]&m[218]&~m[219])|(~m[10]&~m[216]&m[217]&m[218]&~m[219])|(m[10]&~m[216]&~m[217]&~m[218]&m[219])|(~m[10]&m[216]&~m[217]&~m[218]&m[219])|(~m[10]&~m[216]&m[217]&~m[218]&m[219])|(~m[10]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[198])|(((m[10]&m[216]&m[217]&~m[218]&~m[219])|(m[10]&m[216]&~m[217]&m[218]&~m[219])|(m[10]&~m[216]&m[217]&m[218]&~m[219])|(~m[10]&m[216]&m[217]&m[218]&~m[219])|(m[10]&m[216]&~m[217]&~m[218]&m[219])|(m[10]&~m[216]&m[217]&~m[218]&m[219])|(~m[10]&m[216]&m[217]&~m[218]&m[219])|(m[10]&~m[216]&~m[217]&m[218]&m[219])|(~m[10]&m[216]&~m[217]&m[218]&m[219])|(~m[10]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[198])|((m[10]&m[216]&m[217]&m[218]&~m[219])|(m[10]&m[216]&m[217]&~m[218]&m[219])|(m[10]&m[216]&~m[217]&m[218]&m[219])|(m[10]&~m[216]&m[217]&m[218]&m[219])|(~m[10]&m[216]&m[217]&m[218]&m[219])|(m[10]&m[216]&m[217]&m[218]&m[219]));
    m[55] = (((m[10]&m[220]&~m[221]&~m[222]&~m[223])|(m[10]&~m[220]&m[221]&~m[222]&~m[223])|(~m[10]&m[220]&m[221]&~m[222]&~m[223])|(m[10]&~m[220]&~m[221]&m[222]&~m[223])|(~m[10]&m[220]&~m[221]&m[222]&~m[223])|(~m[10]&~m[220]&m[221]&m[222]&~m[223])|(m[10]&~m[220]&~m[221]&~m[222]&m[223])|(~m[10]&m[220]&~m[221]&~m[222]&m[223])|(~m[10]&~m[220]&m[221]&~m[222]&m[223])|(~m[10]&~m[220]&~m[221]&m[222]&m[223]))&BiasedRNG[199])|(((m[10]&m[220]&m[221]&~m[222]&~m[223])|(m[10]&m[220]&~m[221]&m[222]&~m[223])|(m[10]&~m[220]&m[221]&m[222]&~m[223])|(~m[10]&m[220]&m[221]&m[222]&~m[223])|(m[10]&m[220]&~m[221]&~m[222]&m[223])|(m[10]&~m[220]&m[221]&~m[222]&m[223])|(~m[10]&m[220]&m[221]&~m[222]&m[223])|(m[10]&~m[220]&~m[221]&m[222]&m[223])|(~m[10]&m[220]&~m[221]&m[222]&m[223])|(~m[10]&~m[220]&m[221]&m[222]&m[223]))&~BiasedRNG[199])|((m[10]&m[220]&m[221]&m[222]&~m[223])|(m[10]&m[220]&m[221]&~m[222]&m[223])|(m[10]&m[220]&~m[221]&m[222]&m[223])|(m[10]&~m[220]&m[221]&m[222]&m[223])|(~m[10]&m[220]&m[221]&m[222]&m[223])|(m[10]&m[220]&m[221]&m[222]&m[223]));
    m[56] = (((m[10]&m[224]&~m[225]&~m[226]&~m[227])|(m[10]&~m[224]&m[225]&~m[226]&~m[227])|(~m[10]&m[224]&m[225]&~m[226]&~m[227])|(m[10]&~m[224]&~m[225]&m[226]&~m[227])|(~m[10]&m[224]&~m[225]&m[226]&~m[227])|(~m[10]&~m[224]&m[225]&m[226]&~m[227])|(m[10]&~m[224]&~m[225]&~m[226]&m[227])|(~m[10]&m[224]&~m[225]&~m[226]&m[227])|(~m[10]&~m[224]&m[225]&~m[226]&m[227])|(~m[10]&~m[224]&~m[225]&m[226]&m[227]))&BiasedRNG[200])|(((m[10]&m[224]&m[225]&~m[226]&~m[227])|(m[10]&m[224]&~m[225]&m[226]&~m[227])|(m[10]&~m[224]&m[225]&m[226]&~m[227])|(~m[10]&m[224]&m[225]&m[226]&~m[227])|(m[10]&m[224]&~m[225]&~m[226]&m[227])|(m[10]&~m[224]&m[225]&~m[226]&m[227])|(~m[10]&m[224]&m[225]&~m[226]&m[227])|(m[10]&~m[224]&~m[225]&m[226]&m[227])|(~m[10]&m[224]&~m[225]&m[226]&m[227])|(~m[10]&~m[224]&m[225]&m[226]&m[227]))&~BiasedRNG[200])|((m[10]&m[224]&m[225]&m[226]&~m[227])|(m[10]&m[224]&m[225]&~m[226]&m[227])|(m[10]&m[224]&~m[225]&m[226]&m[227])|(m[10]&~m[224]&m[225]&m[226]&m[227])|(~m[10]&m[224]&m[225]&m[226]&m[227])|(m[10]&m[224]&m[225]&m[226]&m[227]));
    m[57] = (((m[11]&m[228]&~m[229]&~m[230]&~m[231])|(m[11]&~m[228]&m[229]&~m[230]&~m[231])|(~m[11]&m[228]&m[229]&~m[230]&~m[231])|(m[11]&~m[228]&~m[229]&m[230]&~m[231])|(~m[11]&m[228]&~m[229]&m[230]&~m[231])|(~m[11]&~m[228]&m[229]&m[230]&~m[231])|(m[11]&~m[228]&~m[229]&~m[230]&m[231])|(~m[11]&m[228]&~m[229]&~m[230]&m[231])|(~m[11]&~m[228]&m[229]&~m[230]&m[231])|(~m[11]&~m[228]&~m[229]&m[230]&m[231]))&BiasedRNG[201])|(((m[11]&m[228]&m[229]&~m[230]&~m[231])|(m[11]&m[228]&~m[229]&m[230]&~m[231])|(m[11]&~m[228]&m[229]&m[230]&~m[231])|(~m[11]&m[228]&m[229]&m[230]&~m[231])|(m[11]&m[228]&~m[229]&~m[230]&m[231])|(m[11]&~m[228]&m[229]&~m[230]&m[231])|(~m[11]&m[228]&m[229]&~m[230]&m[231])|(m[11]&~m[228]&~m[229]&m[230]&m[231])|(~m[11]&m[228]&~m[229]&m[230]&m[231])|(~m[11]&~m[228]&m[229]&m[230]&m[231]))&~BiasedRNG[201])|((m[11]&m[228]&m[229]&m[230]&~m[231])|(m[11]&m[228]&m[229]&~m[230]&m[231])|(m[11]&m[228]&~m[229]&m[230]&m[231])|(m[11]&~m[228]&m[229]&m[230]&m[231])|(~m[11]&m[228]&m[229]&m[230]&m[231])|(m[11]&m[228]&m[229]&m[230]&m[231]));
    m[58] = (((m[11]&m[232]&~m[233]&~m[234]&~m[235])|(m[11]&~m[232]&m[233]&~m[234]&~m[235])|(~m[11]&m[232]&m[233]&~m[234]&~m[235])|(m[11]&~m[232]&~m[233]&m[234]&~m[235])|(~m[11]&m[232]&~m[233]&m[234]&~m[235])|(~m[11]&~m[232]&m[233]&m[234]&~m[235])|(m[11]&~m[232]&~m[233]&~m[234]&m[235])|(~m[11]&m[232]&~m[233]&~m[234]&m[235])|(~m[11]&~m[232]&m[233]&~m[234]&m[235])|(~m[11]&~m[232]&~m[233]&m[234]&m[235]))&BiasedRNG[202])|(((m[11]&m[232]&m[233]&~m[234]&~m[235])|(m[11]&m[232]&~m[233]&m[234]&~m[235])|(m[11]&~m[232]&m[233]&m[234]&~m[235])|(~m[11]&m[232]&m[233]&m[234]&~m[235])|(m[11]&m[232]&~m[233]&~m[234]&m[235])|(m[11]&~m[232]&m[233]&~m[234]&m[235])|(~m[11]&m[232]&m[233]&~m[234]&m[235])|(m[11]&~m[232]&~m[233]&m[234]&m[235])|(~m[11]&m[232]&~m[233]&m[234]&m[235])|(~m[11]&~m[232]&m[233]&m[234]&m[235]))&~BiasedRNG[202])|((m[11]&m[232]&m[233]&m[234]&~m[235])|(m[11]&m[232]&m[233]&~m[234]&m[235])|(m[11]&m[232]&~m[233]&m[234]&m[235])|(m[11]&~m[232]&m[233]&m[234]&m[235])|(~m[11]&m[232]&m[233]&m[234]&m[235])|(m[11]&m[232]&m[233]&m[234]&m[235]));
    m[59] = (((m[11]&m[236]&~m[237]&~m[238]&~m[239])|(m[11]&~m[236]&m[237]&~m[238]&~m[239])|(~m[11]&m[236]&m[237]&~m[238]&~m[239])|(m[11]&~m[236]&~m[237]&m[238]&~m[239])|(~m[11]&m[236]&~m[237]&m[238]&~m[239])|(~m[11]&~m[236]&m[237]&m[238]&~m[239])|(m[11]&~m[236]&~m[237]&~m[238]&m[239])|(~m[11]&m[236]&~m[237]&~m[238]&m[239])|(~m[11]&~m[236]&m[237]&~m[238]&m[239])|(~m[11]&~m[236]&~m[237]&m[238]&m[239]))&BiasedRNG[203])|(((m[11]&m[236]&m[237]&~m[238]&~m[239])|(m[11]&m[236]&~m[237]&m[238]&~m[239])|(m[11]&~m[236]&m[237]&m[238]&~m[239])|(~m[11]&m[236]&m[237]&m[238]&~m[239])|(m[11]&m[236]&~m[237]&~m[238]&m[239])|(m[11]&~m[236]&m[237]&~m[238]&m[239])|(~m[11]&m[236]&m[237]&~m[238]&m[239])|(m[11]&~m[236]&~m[237]&m[238]&m[239])|(~m[11]&m[236]&~m[237]&m[238]&m[239])|(~m[11]&~m[236]&m[237]&m[238]&m[239]))&~BiasedRNG[203])|((m[11]&m[236]&m[237]&m[238]&~m[239])|(m[11]&m[236]&m[237]&~m[238]&m[239])|(m[11]&m[236]&~m[237]&m[238]&m[239])|(m[11]&~m[236]&m[237]&m[238]&m[239])|(~m[11]&m[236]&m[237]&m[238]&m[239])|(m[11]&m[236]&m[237]&m[238]&m[239]));
    m[60] = (((m[12]&m[240]&~m[241]&~m[242]&~m[243])|(m[12]&~m[240]&m[241]&~m[242]&~m[243])|(~m[12]&m[240]&m[241]&~m[242]&~m[243])|(m[12]&~m[240]&~m[241]&m[242]&~m[243])|(~m[12]&m[240]&~m[241]&m[242]&~m[243])|(~m[12]&~m[240]&m[241]&m[242]&~m[243])|(m[12]&~m[240]&~m[241]&~m[242]&m[243])|(~m[12]&m[240]&~m[241]&~m[242]&m[243])|(~m[12]&~m[240]&m[241]&~m[242]&m[243])|(~m[12]&~m[240]&~m[241]&m[242]&m[243]))&BiasedRNG[204])|(((m[12]&m[240]&m[241]&~m[242]&~m[243])|(m[12]&m[240]&~m[241]&m[242]&~m[243])|(m[12]&~m[240]&m[241]&m[242]&~m[243])|(~m[12]&m[240]&m[241]&m[242]&~m[243])|(m[12]&m[240]&~m[241]&~m[242]&m[243])|(m[12]&~m[240]&m[241]&~m[242]&m[243])|(~m[12]&m[240]&m[241]&~m[242]&m[243])|(m[12]&~m[240]&~m[241]&m[242]&m[243])|(~m[12]&m[240]&~m[241]&m[242]&m[243])|(~m[12]&~m[240]&m[241]&m[242]&m[243]))&~BiasedRNG[204])|((m[12]&m[240]&m[241]&m[242]&~m[243])|(m[12]&m[240]&m[241]&~m[242]&m[243])|(m[12]&m[240]&~m[241]&m[242]&m[243])|(m[12]&~m[240]&m[241]&m[242]&m[243])|(~m[12]&m[240]&m[241]&m[242]&m[243])|(m[12]&m[240]&m[241]&m[242]&m[243]));
    m[61] = (((m[12]&m[244]&~m[245]&~m[246]&~m[247])|(m[12]&~m[244]&m[245]&~m[246]&~m[247])|(~m[12]&m[244]&m[245]&~m[246]&~m[247])|(m[12]&~m[244]&~m[245]&m[246]&~m[247])|(~m[12]&m[244]&~m[245]&m[246]&~m[247])|(~m[12]&~m[244]&m[245]&m[246]&~m[247])|(m[12]&~m[244]&~m[245]&~m[246]&m[247])|(~m[12]&m[244]&~m[245]&~m[246]&m[247])|(~m[12]&~m[244]&m[245]&~m[246]&m[247])|(~m[12]&~m[244]&~m[245]&m[246]&m[247]))&BiasedRNG[205])|(((m[12]&m[244]&m[245]&~m[246]&~m[247])|(m[12]&m[244]&~m[245]&m[246]&~m[247])|(m[12]&~m[244]&m[245]&m[246]&~m[247])|(~m[12]&m[244]&m[245]&m[246]&~m[247])|(m[12]&m[244]&~m[245]&~m[246]&m[247])|(m[12]&~m[244]&m[245]&~m[246]&m[247])|(~m[12]&m[244]&m[245]&~m[246]&m[247])|(m[12]&~m[244]&~m[245]&m[246]&m[247])|(~m[12]&m[244]&~m[245]&m[246]&m[247])|(~m[12]&~m[244]&m[245]&m[246]&m[247]))&~BiasedRNG[205])|((m[12]&m[244]&m[245]&m[246]&~m[247])|(m[12]&m[244]&m[245]&~m[246]&m[247])|(m[12]&m[244]&~m[245]&m[246]&m[247])|(m[12]&~m[244]&m[245]&m[246]&m[247])|(~m[12]&m[244]&m[245]&m[246]&m[247])|(m[12]&m[244]&m[245]&m[246]&m[247]));
    m[62] = (((m[12]&m[248]&~m[249]&~m[250]&~m[251])|(m[12]&~m[248]&m[249]&~m[250]&~m[251])|(~m[12]&m[248]&m[249]&~m[250]&~m[251])|(m[12]&~m[248]&~m[249]&m[250]&~m[251])|(~m[12]&m[248]&~m[249]&m[250]&~m[251])|(~m[12]&~m[248]&m[249]&m[250]&~m[251])|(m[12]&~m[248]&~m[249]&~m[250]&m[251])|(~m[12]&m[248]&~m[249]&~m[250]&m[251])|(~m[12]&~m[248]&m[249]&~m[250]&m[251])|(~m[12]&~m[248]&~m[249]&m[250]&m[251]))&BiasedRNG[206])|(((m[12]&m[248]&m[249]&~m[250]&~m[251])|(m[12]&m[248]&~m[249]&m[250]&~m[251])|(m[12]&~m[248]&m[249]&m[250]&~m[251])|(~m[12]&m[248]&m[249]&m[250]&~m[251])|(m[12]&m[248]&~m[249]&~m[250]&m[251])|(m[12]&~m[248]&m[249]&~m[250]&m[251])|(~m[12]&m[248]&m[249]&~m[250]&m[251])|(m[12]&~m[248]&~m[249]&m[250]&m[251])|(~m[12]&m[248]&~m[249]&m[250]&m[251])|(~m[12]&~m[248]&m[249]&m[250]&m[251]))&~BiasedRNG[206])|((m[12]&m[248]&m[249]&m[250]&~m[251])|(m[12]&m[248]&m[249]&~m[250]&m[251])|(m[12]&m[248]&~m[249]&m[250]&m[251])|(m[12]&~m[248]&m[249]&m[250]&m[251])|(~m[12]&m[248]&m[249]&m[250]&m[251])|(m[12]&m[248]&m[249]&m[250]&m[251]));
    m[63] = (((m[13]&m[252]&~m[253]&~m[254]&~m[255])|(m[13]&~m[252]&m[253]&~m[254]&~m[255])|(~m[13]&m[252]&m[253]&~m[254]&~m[255])|(m[13]&~m[252]&~m[253]&m[254]&~m[255])|(~m[13]&m[252]&~m[253]&m[254]&~m[255])|(~m[13]&~m[252]&m[253]&m[254]&~m[255])|(m[13]&~m[252]&~m[253]&~m[254]&m[255])|(~m[13]&m[252]&~m[253]&~m[254]&m[255])|(~m[13]&~m[252]&m[253]&~m[254]&m[255])|(~m[13]&~m[252]&~m[253]&m[254]&m[255]))&BiasedRNG[207])|(((m[13]&m[252]&m[253]&~m[254]&~m[255])|(m[13]&m[252]&~m[253]&m[254]&~m[255])|(m[13]&~m[252]&m[253]&m[254]&~m[255])|(~m[13]&m[252]&m[253]&m[254]&~m[255])|(m[13]&m[252]&~m[253]&~m[254]&m[255])|(m[13]&~m[252]&m[253]&~m[254]&m[255])|(~m[13]&m[252]&m[253]&~m[254]&m[255])|(m[13]&~m[252]&~m[253]&m[254]&m[255])|(~m[13]&m[252]&~m[253]&m[254]&m[255])|(~m[13]&~m[252]&m[253]&m[254]&m[255]))&~BiasedRNG[207])|((m[13]&m[252]&m[253]&m[254]&~m[255])|(m[13]&m[252]&m[253]&~m[254]&m[255])|(m[13]&m[252]&~m[253]&m[254]&m[255])|(m[13]&~m[252]&m[253]&m[254]&m[255])|(~m[13]&m[252]&m[253]&m[254]&m[255])|(m[13]&m[252]&m[253]&m[254]&m[255]));
    m[64] = (((m[13]&m[256]&~m[257]&~m[258]&~m[259])|(m[13]&~m[256]&m[257]&~m[258]&~m[259])|(~m[13]&m[256]&m[257]&~m[258]&~m[259])|(m[13]&~m[256]&~m[257]&m[258]&~m[259])|(~m[13]&m[256]&~m[257]&m[258]&~m[259])|(~m[13]&~m[256]&m[257]&m[258]&~m[259])|(m[13]&~m[256]&~m[257]&~m[258]&m[259])|(~m[13]&m[256]&~m[257]&~m[258]&m[259])|(~m[13]&~m[256]&m[257]&~m[258]&m[259])|(~m[13]&~m[256]&~m[257]&m[258]&m[259]))&BiasedRNG[208])|(((m[13]&m[256]&m[257]&~m[258]&~m[259])|(m[13]&m[256]&~m[257]&m[258]&~m[259])|(m[13]&~m[256]&m[257]&m[258]&~m[259])|(~m[13]&m[256]&m[257]&m[258]&~m[259])|(m[13]&m[256]&~m[257]&~m[258]&m[259])|(m[13]&~m[256]&m[257]&~m[258]&m[259])|(~m[13]&m[256]&m[257]&~m[258]&m[259])|(m[13]&~m[256]&~m[257]&m[258]&m[259])|(~m[13]&m[256]&~m[257]&m[258]&m[259])|(~m[13]&~m[256]&m[257]&m[258]&m[259]))&~BiasedRNG[208])|((m[13]&m[256]&m[257]&m[258]&~m[259])|(m[13]&m[256]&m[257]&~m[258]&m[259])|(m[13]&m[256]&~m[257]&m[258]&m[259])|(m[13]&~m[256]&m[257]&m[258]&m[259])|(~m[13]&m[256]&m[257]&m[258]&m[259])|(m[13]&m[256]&m[257]&m[258]&m[259]));
    m[65] = (((m[13]&m[260]&~m[261]&~m[262]&~m[263])|(m[13]&~m[260]&m[261]&~m[262]&~m[263])|(~m[13]&m[260]&m[261]&~m[262]&~m[263])|(m[13]&~m[260]&~m[261]&m[262]&~m[263])|(~m[13]&m[260]&~m[261]&m[262]&~m[263])|(~m[13]&~m[260]&m[261]&m[262]&~m[263])|(m[13]&~m[260]&~m[261]&~m[262]&m[263])|(~m[13]&m[260]&~m[261]&~m[262]&m[263])|(~m[13]&~m[260]&m[261]&~m[262]&m[263])|(~m[13]&~m[260]&~m[261]&m[262]&m[263]))&BiasedRNG[209])|(((m[13]&m[260]&m[261]&~m[262]&~m[263])|(m[13]&m[260]&~m[261]&m[262]&~m[263])|(m[13]&~m[260]&m[261]&m[262]&~m[263])|(~m[13]&m[260]&m[261]&m[262]&~m[263])|(m[13]&m[260]&~m[261]&~m[262]&m[263])|(m[13]&~m[260]&m[261]&~m[262]&m[263])|(~m[13]&m[260]&m[261]&~m[262]&m[263])|(m[13]&~m[260]&~m[261]&m[262]&m[263])|(~m[13]&m[260]&~m[261]&m[262]&m[263])|(~m[13]&~m[260]&m[261]&m[262]&m[263]))&~BiasedRNG[209])|((m[13]&m[260]&m[261]&m[262]&~m[263])|(m[13]&m[260]&m[261]&~m[262]&m[263])|(m[13]&m[260]&~m[261]&m[262]&m[263])|(m[13]&~m[260]&m[261]&m[262]&m[263])|(~m[13]&m[260]&m[261]&m[262]&m[263])|(m[13]&m[260]&m[261]&m[262]&m[263]));
    m[66] = (((m[14]&m[264]&~m[265]&~m[266]&~m[267])|(m[14]&~m[264]&m[265]&~m[266]&~m[267])|(~m[14]&m[264]&m[265]&~m[266]&~m[267])|(m[14]&~m[264]&~m[265]&m[266]&~m[267])|(~m[14]&m[264]&~m[265]&m[266]&~m[267])|(~m[14]&~m[264]&m[265]&m[266]&~m[267])|(m[14]&~m[264]&~m[265]&~m[266]&m[267])|(~m[14]&m[264]&~m[265]&~m[266]&m[267])|(~m[14]&~m[264]&m[265]&~m[266]&m[267])|(~m[14]&~m[264]&~m[265]&m[266]&m[267]))&BiasedRNG[210])|(((m[14]&m[264]&m[265]&~m[266]&~m[267])|(m[14]&m[264]&~m[265]&m[266]&~m[267])|(m[14]&~m[264]&m[265]&m[266]&~m[267])|(~m[14]&m[264]&m[265]&m[266]&~m[267])|(m[14]&m[264]&~m[265]&~m[266]&m[267])|(m[14]&~m[264]&m[265]&~m[266]&m[267])|(~m[14]&m[264]&m[265]&~m[266]&m[267])|(m[14]&~m[264]&~m[265]&m[266]&m[267])|(~m[14]&m[264]&~m[265]&m[266]&m[267])|(~m[14]&~m[264]&m[265]&m[266]&m[267]))&~BiasedRNG[210])|((m[14]&m[264]&m[265]&m[266]&~m[267])|(m[14]&m[264]&m[265]&~m[266]&m[267])|(m[14]&m[264]&~m[265]&m[266]&m[267])|(m[14]&~m[264]&m[265]&m[266]&m[267])|(~m[14]&m[264]&m[265]&m[266]&m[267])|(m[14]&m[264]&m[265]&m[266]&m[267]));
    m[67] = (((m[14]&m[268]&~m[269]&~m[270]&~m[271])|(m[14]&~m[268]&m[269]&~m[270]&~m[271])|(~m[14]&m[268]&m[269]&~m[270]&~m[271])|(m[14]&~m[268]&~m[269]&m[270]&~m[271])|(~m[14]&m[268]&~m[269]&m[270]&~m[271])|(~m[14]&~m[268]&m[269]&m[270]&~m[271])|(m[14]&~m[268]&~m[269]&~m[270]&m[271])|(~m[14]&m[268]&~m[269]&~m[270]&m[271])|(~m[14]&~m[268]&m[269]&~m[270]&m[271])|(~m[14]&~m[268]&~m[269]&m[270]&m[271]))&BiasedRNG[211])|(((m[14]&m[268]&m[269]&~m[270]&~m[271])|(m[14]&m[268]&~m[269]&m[270]&~m[271])|(m[14]&~m[268]&m[269]&m[270]&~m[271])|(~m[14]&m[268]&m[269]&m[270]&~m[271])|(m[14]&m[268]&~m[269]&~m[270]&m[271])|(m[14]&~m[268]&m[269]&~m[270]&m[271])|(~m[14]&m[268]&m[269]&~m[270]&m[271])|(m[14]&~m[268]&~m[269]&m[270]&m[271])|(~m[14]&m[268]&~m[269]&m[270]&m[271])|(~m[14]&~m[268]&m[269]&m[270]&m[271]))&~BiasedRNG[211])|((m[14]&m[268]&m[269]&m[270]&~m[271])|(m[14]&m[268]&m[269]&~m[270]&m[271])|(m[14]&m[268]&~m[269]&m[270]&m[271])|(m[14]&~m[268]&m[269]&m[270]&m[271])|(~m[14]&m[268]&m[269]&m[270]&m[271])|(m[14]&m[268]&m[269]&m[270]&m[271]));
    m[68] = (((m[14]&m[272]&~m[273]&~m[274]&~m[275])|(m[14]&~m[272]&m[273]&~m[274]&~m[275])|(~m[14]&m[272]&m[273]&~m[274]&~m[275])|(m[14]&~m[272]&~m[273]&m[274]&~m[275])|(~m[14]&m[272]&~m[273]&m[274]&~m[275])|(~m[14]&~m[272]&m[273]&m[274]&~m[275])|(m[14]&~m[272]&~m[273]&~m[274]&m[275])|(~m[14]&m[272]&~m[273]&~m[274]&m[275])|(~m[14]&~m[272]&m[273]&~m[274]&m[275])|(~m[14]&~m[272]&~m[273]&m[274]&m[275]))&BiasedRNG[212])|(((m[14]&m[272]&m[273]&~m[274]&~m[275])|(m[14]&m[272]&~m[273]&m[274]&~m[275])|(m[14]&~m[272]&m[273]&m[274]&~m[275])|(~m[14]&m[272]&m[273]&m[274]&~m[275])|(m[14]&m[272]&~m[273]&~m[274]&m[275])|(m[14]&~m[272]&m[273]&~m[274]&m[275])|(~m[14]&m[272]&m[273]&~m[274]&m[275])|(m[14]&~m[272]&~m[273]&m[274]&m[275])|(~m[14]&m[272]&~m[273]&m[274]&m[275])|(~m[14]&~m[272]&m[273]&m[274]&m[275]))&~BiasedRNG[212])|((m[14]&m[272]&m[273]&m[274]&~m[275])|(m[14]&m[272]&m[273]&~m[274]&m[275])|(m[14]&m[272]&~m[273]&m[274]&m[275])|(m[14]&~m[272]&m[273]&m[274]&m[275])|(~m[14]&m[272]&m[273]&m[274]&m[275])|(m[14]&m[272]&m[273]&m[274]&m[275]));
    m[69] = (((m[15]&m[276]&~m[277]&~m[278]&~m[279])|(m[15]&~m[276]&m[277]&~m[278]&~m[279])|(~m[15]&m[276]&m[277]&~m[278]&~m[279])|(m[15]&~m[276]&~m[277]&m[278]&~m[279])|(~m[15]&m[276]&~m[277]&m[278]&~m[279])|(~m[15]&~m[276]&m[277]&m[278]&~m[279])|(m[15]&~m[276]&~m[277]&~m[278]&m[279])|(~m[15]&m[276]&~m[277]&~m[278]&m[279])|(~m[15]&~m[276]&m[277]&~m[278]&m[279])|(~m[15]&~m[276]&~m[277]&m[278]&m[279]))&BiasedRNG[213])|(((m[15]&m[276]&m[277]&~m[278]&~m[279])|(m[15]&m[276]&~m[277]&m[278]&~m[279])|(m[15]&~m[276]&m[277]&m[278]&~m[279])|(~m[15]&m[276]&m[277]&m[278]&~m[279])|(m[15]&m[276]&~m[277]&~m[278]&m[279])|(m[15]&~m[276]&m[277]&~m[278]&m[279])|(~m[15]&m[276]&m[277]&~m[278]&m[279])|(m[15]&~m[276]&~m[277]&m[278]&m[279])|(~m[15]&m[276]&~m[277]&m[278]&m[279])|(~m[15]&~m[276]&m[277]&m[278]&m[279]))&~BiasedRNG[213])|((m[15]&m[276]&m[277]&m[278]&~m[279])|(m[15]&m[276]&m[277]&~m[278]&m[279])|(m[15]&m[276]&~m[277]&m[278]&m[279])|(m[15]&~m[276]&m[277]&m[278]&m[279])|(~m[15]&m[276]&m[277]&m[278]&m[279])|(m[15]&m[276]&m[277]&m[278]&m[279]));
    m[70] = (((m[15]&m[280]&~m[281]&~m[282]&~m[283])|(m[15]&~m[280]&m[281]&~m[282]&~m[283])|(~m[15]&m[280]&m[281]&~m[282]&~m[283])|(m[15]&~m[280]&~m[281]&m[282]&~m[283])|(~m[15]&m[280]&~m[281]&m[282]&~m[283])|(~m[15]&~m[280]&m[281]&m[282]&~m[283])|(m[15]&~m[280]&~m[281]&~m[282]&m[283])|(~m[15]&m[280]&~m[281]&~m[282]&m[283])|(~m[15]&~m[280]&m[281]&~m[282]&m[283])|(~m[15]&~m[280]&~m[281]&m[282]&m[283]))&BiasedRNG[214])|(((m[15]&m[280]&m[281]&~m[282]&~m[283])|(m[15]&m[280]&~m[281]&m[282]&~m[283])|(m[15]&~m[280]&m[281]&m[282]&~m[283])|(~m[15]&m[280]&m[281]&m[282]&~m[283])|(m[15]&m[280]&~m[281]&~m[282]&m[283])|(m[15]&~m[280]&m[281]&~m[282]&m[283])|(~m[15]&m[280]&m[281]&~m[282]&m[283])|(m[15]&~m[280]&~m[281]&m[282]&m[283])|(~m[15]&m[280]&~m[281]&m[282]&m[283])|(~m[15]&~m[280]&m[281]&m[282]&m[283]))&~BiasedRNG[214])|((m[15]&m[280]&m[281]&m[282]&~m[283])|(m[15]&m[280]&m[281]&~m[282]&m[283])|(m[15]&m[280]&~m[281]&m[282]&m[283])|(m[15]&~m[280]&m[281]&m[282]&m[283])|(~m[15]&m[280]&m[281]&m[282]&m[283])|(m[15]&m[280]&m[281]&m[282]&m[283]));
    m[71] = (((m[15]&m[284]&~m[285]&~m[286]&~m[287])|(m[15]&~m[284]&m[285]&~m[286]&~m[287])|(~m[15]&m[284]&m[285]&~m[286]&~m[287])|(m[15]&~m[284]&~m[285]&m[286]&~m[287])|(~m[15]&m[284]&~m[285]&m[286]&~m[287])|(~m[15]&~m[284]&m[285]&m[286]&~m[287])|(m[15]&~m[284]&~m[285]&~m[286]&m[287])|(~m[15]&m[284]&~m[285]&~m[286]&m[287])|(~m[15]&~m[284]&m[285]&~m[286]&m[287])|(~m[15]&~m[284]&~m[285]&m[286]&m[287]))&BiasedRNG[215])|(((m[15]&m[284]&m[285]&~m[286]&~m[287])|(m[15]&m[284]&~m[285]&m[286]&~m[287])|(m[15]&~m[284]&m[285]&m[286]&~m[287])|(~m[15]&m[284]&m[285]&m[286]&~m[287])|(m[15]&m[284]&~m[285]&~m[286]&m[287])|(m[15]&~m[284]&m[285]&~m[286]&m[287])|(~m[15]&m[284]&m[285]&~m[286]&m[287])|(m[15]&~m[284]&~m[285]&m[286]&m[287])|(~m[15]&m[284]&~m[285]&m[286]&m[287])|(~m[15]&~m[284]&m[285]&m[286]&m[287]))&~BiasedRNG[215])|((m[15]&m[284]&m[285]&m[286]&~m[287])|(m[15]&m[284]&m[285]&~m[286]&m[287])|(m[15]&m[284]&~m[285]&m[286]&m[287])|(m[15]&~m[284]&m[285]&m[286]&m[287])|(~m[15]&m[284]&m[285]&m[286]&m[287])|(m[15]&m[284]&m[285]&m[286]&m[287]));
    m[72] = (((m[16]&m[288]&~m[289]&~m[290]&~m[291])|(m[16]&~m[288]&m[289]&~m[290]&~m[291])|(~m[16]&m[288]&m[289]&~m[290]&~m[291])|(m[16]&~m[288]&~m[289]&m[290]&~m[291])|(~m[16]&m[288]&~m[289]&m[290]&~m[291])|(~m[16]&~m[288]&m[289]&m[290]&~m[291])|(m[16]&~m[288]&~m[289]&~m[290]&m[291])|(~m[16]&m[288]&~m[289]&~m[290]&m[291])|(~m[16]&~m[288]&m[289]&~m[290]&m[291])|(~m[16]&~m[288]&~m[289]&m[290]&m[291]))&BiasedRNG[216])|(((m[16]&m[288]&m[289]&~m[290]&~m[291])|(m[16]&m[288]&~m[289]&m[290]&~m[291])|(m[16]&~m[288]&m[289]&m[290]&~m[291])|(~m[16]&m[288]&m[289]&m[290]&~m[291])|(m[16]&m[288]&~m[289]&~m[290]&m[291])|(m[16]&~m[288]&m[289]&~m[290]&m[291])|(~m[16]&m[288]&m[289]&~m[290]&m[291])|(m[16]&~m[288]&~m[289]&m[290]&m[291])|(~m[16]&m[288]&~m[289]&m[290]&m[291])|(~m[16]&~m[288]&m[289]&m[290]&m[291]))&~BiasedRNG[216])|((m[16]&m[288]&m[289]&m[290]&~m[291])|(m[16]&m[288]&m[289]&~m[290]&m[291])|(m[16]&m[288]&~m[289]&m[290]&m[291])|(m[16]&~m[288]&m[289]&m[290]&m[291])|(~m[16]&m[288]&m[289]&m[290]&m[291])|(m[16]&m[288]&m[289]&m[290]&m[291]));
    m[73] = (((m[16]&m[292]&~m[293]&~m[294]&~m[295])|(m[16]&~m[292]&m[293]&~m[294]&~m[295])|(~m[16]&m[292]&m[293]&~m[294]&~m[295])|(m[16]&~m[292]&~m[293]&m[294]&~m[295])|(~m[16]&m[292]&~m[293]&m[294]&~m[295])|(~m[16]&~m[292]&m[293]&m[294]&~m[295])|(m[16]&~m[292]&~m[293]&~m[294]&m[295])|(~m[16]&m[292]&~m[293]&~m[294]&m[295])|(~m[16]&~m[292]&m[293]&~m[294]&m[295])|(~m[16]&~m[292]&~m[293]&m[294]&m[295]))&BiasedRNG[217])|(((m[16]&m[292]&m[293]&~m[294]&~m[295])|(m[16]&m[292]&~m[293]&m[294]&~m[295])|(m[16]&~m[292]&m[293]&m[294]&~m[295])|(~m[16]&m[292]&m[293]&m[294]&~m[295])|(m[16]&m[292]&~m[293]&~m[294]&m[295])|(m[16]&~m[292]&m[293]&~m[294]&m[295])|(~m[16]&m[292]&m[293]&~m[294]&m[295])|(m[16]&~m[292]&~m[293]&m[294]&m[295])|(~m[16]&m[292]&~m[293]&m[294]&m[295])|(~m[16]&~m[292]&m[293]&m[294]&m[295]))&~BiasedRNG[217])|((m[16]&m[292]&m[293]&m[294]&~m[295])|(m[16]&m[292]&m[293]&~m[294]&m[295])|(m[16]&m[292]&~m[293]&m[294]&m[295])|(m[16]&~m[292]&m[293]&m[294]&m[295])|(~m[16]&m[292]&m[293]&m[294]&m[295])|(m[16]&m[292]&m[293]&m[294]&m[295]));
    m[74] = (((m[16]&m[296]&~m[297]&~m[298]&~m[299])|(m[16]&~m[296]&m[297]&~m[298]&~m[299])|(~m[16]&m[296]&m[297]&~m[298]&~m[299])|(m[16]&~m[296]&~m[297]&m[298]&~m[299])|(~m[16]&m[296]&~m[297]&m[298]&~m[299])|(~m[16]&~m[296]&m[297]&m[298]&~m[299])|(m[16]&~m[296]&~m[297]&~m[298]&m[299])|(~m[16]&m[296]&~m[297]&~m[298]&m[299])|(~m[16]&~m[296]&m[297]&~m[298]&m[299])|(~m[16]&~m[296]&~m[297]&m[298]&m[299]))&BiasedRNG[218])|(((m[16]&m[296]&m[297]&~m[298]&~m[299])|(m[16]&m[296]&~m[297]&m[298]&~m[299])|(m[16]&~m[296]&m[297]&m[298]&~m[299])|(~m[16]&m[296]&m[297]&m[298]&~m[299])|(m[16]&m[296]&~m[297]&~m[298]&m[299])|(m[16]&~m[296]&m[297]&~m[298]&m[299])|(~m[16]&m[296]&m[297]&~m[298]&m[299])|(m[16]&~m[296]&~m[297]&m[298]&m[299])|(~m[16]&m[296]&~m[297]&m[298]&m[299])|(~m[16]&~m[296]&m[297]&m[298]&m[299]))&~BiasedRNG[218])|((m[16]&m[296]&m[297]&m[298]&~m[299])|(m[16]&m[296]&m[297]&~m[298]&m[299])|(m[16]&m[296]&~m[297]&m[298]&m[299])|(m[16]&~m[296]&m[297]&m[298]&m[299])|(~m[16]&m[296]&m[297]&m[298]&m[299])|(m[16]&m[296]&m[297]&m[298]&m[299]));
    m[75] = (((m[17]&m[300]&~m[301]&~m[302]&~m[303])|(m[17]&~m[300]&m[301]&~m[302]&~m[303])|(~m[17]&m[300]&m[301]&~m[302]&~m[303])|(m[17]&~m[300]&~m[301]&m[302]&~m[303])|(~m[17]&m[300]&~m[301]&m[302]&~m[303])|(~m[17]&~m[300]&m[301]&m[302]&~m[303])|(m[17]&~m[300]&~m[301]&~m[302]&m[303])|(~m[17]&m[300]&~m[301]&~m[302]&m[303])|(~m[17]&~m[300]&m[301]&~m[302]&m[303])|(~m[17]&~m[300]&~m[301]&m[302]&m[303]))&BiasedRNG[219])|(((m[17]&m[300]&m[301]&~m[302]&~m[303])|(m[17]&m[300]&~m[301]&m[302]&~m[303])|(m[17]&~m[300]&m[301]&m[302]&~m[303])|(~m[17]&m[300]&m[301]&m[302]&~m[303])|(m[17]&m[300]&~m[301]&~m[302]&m[303])|(m[17]&~m[300]&m[301]&~m[302]&m[303])|(~m[17]&m[300]&m[301]&~m[302]&m[303])|(m[17]&~m[300]&~m[301]&m[302]&m[303])|(~m[17]&m[300]&~m[301]&m[302]&m[303])|(~m[17]&~m[300]&m[301]&m[302]&m[303]))&~BiasedRNG[219])|((m[17]&m[300]&m[301]&m[302]&~m[303])|(m[17]&m[300]&m[301]&~m[302]&m[303])|(m[17]&m[300]&~m[301]&m[302]&m[303])|(m[17]&~m[300]&m[301]&m[302]&m[303])|(~m[17]&m[300]&m[301]&m[302]&m[303])|(m[17]&m[300]&m[301]&m[302]&m[303]));
    m[76] = (((m[17]&m[304]&~m[305]&~m[306]&~m[307])|(m[17]&~m[304]&m[305]&~m[306]&~m[307])|(~m[17]&m[304]&m[305]&~m[306]&~m[307])|(m[17]&~m[304]&~m[305]&m[306]&~m[307])|(~m[17]&m[304]&~m[305]&m[306]&~m[307])|(~m[17]&~m[304]&m[305]&m[306]&~m[307])|(m[17]&~m[304]&~m[305]&~m[306]&m[307])|(~m[17]&m[304]&~m[305]&~m[306]&m[307])|(~m[17]&~m[304]&m[305]&~m[306]&m[307])|(~m[17]&~m[304]&~m[305]&m[306]&m[307]))&BiasedRNG[220])|(((m[17]&m[304]&m[305]&~m[306]&~m[307])|(m[17]&m[304]&~m[305]&m[306]&~m[307])|(m[17]&~m[304]&m[305]&m[306]&~m[307])|(~m[17]&m[304]&m[305]&m[306]&~m[307])|(m[17]&m[304]&~m[305]&~m[306]&m[307])|(m[17]&~m[304]&m[305]&~m[306]&m[307])|(~m[17]&m[304]&m[305]&~m[306]&m[307])|(m[17]&~m[304]&~m[305]&m[306]&m[307])|(~m[17]&m[304]&~m[305]&m[306]&m[307])|(~m[17]&~m[304]&m[305]&m[306]&m[307]))&~BiasedRNG[220])|((m[17]&m[304]&m[305]&m[306]&~m[307])|(m[17]&m[304]&m[305]&~m[306]&m[307])|(m[17]&m[304]&~m[305]&m[306]&m[307])|(m[17]&~m[304]&m[305]&m[306]&m[307])|(~m[17]&m[304]&m[305]&m[306]&m[307])|(m[17]&m[304]&m[305]&m[306]&m[307]));
    m[77] = (((m[17]&m[308]&~m[309]&~m[310]&~m[311])|(m[17]&~m[308]&m[309]&~m[310]&~m[311])|(~m[17]&m[308]&m[309]&~m[310]&~m[311])|(m[17]&~m[308]&~m[309]&m[310]&~m[311])|(~m[17]&m[308]&~m[309]&m[310]&~m[311])|(~m[17]&~m[308]&m[309]&m[310]&~m[311])|(m[17]&~m[308]&~m[309]&~m[310]&m[311])|(~m[17]&m[308]&~m[309]&~m[310]&m[311])|(~m[17]&~m[308]&m[309]&~m[310]&m[311])|(~m[17]&~m[308]&~m[309]&m[310]&m[311]))&BiasedRNG[221])|(((m[17]&m[308]&m[309]&~m[310]&~m[311])|(m[17]&m[308]&~m[309]&m[310]&~m[311])|(m[17]&~m[308]&m[309]&m[310]&~m[311])|(~m[17]&m[308]&m[309]&m[310]&~m[311])|(m[17]&m[308]&~m[309]&~m[310]&m[311])|(m[17]&~m[308]&m[309]&~m[310]&m[311])|(~m[17]&m[308]&m[309]&~m[310]&m[311])|(m[17]&~m[308]&~m[309]&m[310]&m[311])|(~m[17]&m[308]&~m[309]&m[310]&m[311])|(~m[17]&~m[308]&m[309]&m[310]&m[311]))&~BiasedRNG[221])|((m[17]&m[308]&m[309]&m[310]&~m[311])|(m[17]&m[308]&m[309]&~m[310]&m[311])|(m[17]&m[308]&~m[309]&m[310]&m[311])|(m[17]&~m[308]&m[309]&m[310]&m[311])|(~m[17]&m[308]&m[309]&m[310]&m[311])|(m[17]&m[308]&m[309]&m[310]&m[311]));
    m[78] = (((m[18]&m[312]&~m[313]&~m[314]&~m[315])|(m[18]&~m[312]&m[313]&~m[314]&~m[315])|(~m[18]&m[312]&m[313]&~m[314]&~m[315])|(m[18]&~m[312]&~m[313]&m[314]&~m[315])|(~m[18]&m[312]&~m[313]&m[314]&~m[315])|(~m[18]&~m[312]&m[313]&m[314]&~m[315])|(m[18]&~m[312]&~m[313]&~m[314]&m[315])|(~m[18]&m[312]&~m[313]&~m[314]&m[315])|(~m[18]&~m[312]&m[313]&~m[314]&m[315])|(~m[18]&~m[312]&~m[313]&m[314]&m[315]))&BiasedRNG[222])|(((m[18]&m[312]&m[313]&~m[314]&~m[315])|(m[18]&m[312]&~m[313]&m[314]&~m[315])|(m[18]&~m[312]&m[313]&m[314]&~m[315])|(~m[18]&m[312]&m[313]&m[314]&~m[315])|(m[18]&m[312]&~m[313]&~m[314]&m[315])|(m[18]&~m[312]&m[313]&~m[314]&m[315])|(~m[18]&m[312]&m[313]&~m[314]&m[315])|(m[18]&~m[312]&~m[313]&m[314]&m[315])|(~m[18]&m[312]&~m[313]&m[314]&m[315])|(~m[18]&~m[312]&m[313]&m[314]&m[315]))&~BiasedRNG[222])|((m[18]&m[312]&m[313]&m[314]&~m[315])|(m[18]&m[312]&m[313]&~m[314]&m[315])|(m[18]&m[312]&~m[313]&m[314]&m[315])|(m[18]&~m[312]&m[313]&m[314]&m[315])|(~m[18]&m[312]&m[313]&m[314]&m[315])|(m[18]&m[312]&m[313]&m[314]&m[315]));
    m[79] = (((m[18]&m[316]&~m[317]&~m[318]&~m[319])|(m[18]&~m[316]&m[317]&~m[318]&~m[319])|(~m[18]&m[316]&m[317]&~m[318]&~m[319])|(m[18]&~m[316]&~m[317]&m[318]&~m[319])|(~m[18]&m[316]&~m[317]&m[318]&~m[319])|(~m[18]&~m[316]&m[317]&m[318]&~m[319])|(m[18]&~m[316]&~m[317]&~m[318]&m[319])|(~m[18]&m[316]&~m[317]&~m[318]&m[319])|(~m[18]&~m[316]&m[317]&~m[318]&m[319])|(~m[18]&~m[316]&~m[317]&m[318]&m[319]))&BiasedRNG[223])|(((m[18]&m[316]&m[317]&~m[318]&~m[319])|(m[18]&m[316]&~m[317]&m[318]&~m[319])|(m[18]&~m[316]&m[317]&m[318]&~m[319])|(~m[18]&m[316]&m[317]&m[318]&~m[319])|(m[18]&m[316]&~m[317]&~m[318]&m[319])|(m[18]&~m[316]&m[317]&~m[318]&m[319])|(~m[18]&m[316]&m[317]&~m[318]&m[319])|(m[18]&~m[316]&~m[317]&m[318]&m[319])|(~m[18]&m[316]&~m[317]&m[318]&m[319])|(~m[18]&~m[316]&m[317]&m[318]&m[319]))&~BiasedRNG[223])|((m[18]&m[316]&m[317]&m[318]&~m[319])|(m[18]&m[316]&m[317]&~m[318]&m[319])|(m[18]&m[316]&~m[317]&m[318]&m[319])|(m[18]&~m[316]&m[317]&m[318]&m[319])|(~m[18]&m[316]&m[317]&m[318]&m[319])|(m[18]&m[316]&m[317]&m[318]&m[319]));
    m[80] = (((m[18]&m[320]&~m[321]&~m[322]&~m[323])|(m[18]&~m[320]&m[321]&~m[322]&~m[323])|(~m[18]&m[320]&m[321]&~m[322]&~m[323])|(m[18]&~m[320]&~m[321]&m[322]&~m[323])|(~m[18]&m[320]&~m[321]&m[322]&~m[323])|(~m[18]&~m[320]&m[321]&m[322]&~m[323])|(m[18]&~m[320]&~m[321]&~m[322]&m[323])|(~m[18]&m[320]&~m[321]&~m[322]&m[323])|(~m[18]&~m[320]&m[321]&~m[322]&m[323])|(~m[18]&~m[320]&~m[321]&m[322]&m[323]))&BiasedRNG[224])|(((m[18]&m[320]&m[321]&~m[322]&~m[323])|(m[18]&m[320]&~m[321]&m[322]&~m[323])|(m[18]&~m[320]&m[321]&m[322]&~m[323])|(~m[18]&m[320]&m[321]&m[322]&~m[323])|(m[18]&m[320]&~m[321]&~m[322]&m[323])|(m[18]&~m[320]&m[321]&~m[322]&m[323])|(~m[18]&m[320]&m[321]&~m[322]&m[323])|(m[18]&~m[320]&~m[321]&m[322]&m[323])|(~m[18]&m[320]&~m[321]&m[322]&m[323])|(~m[18]&~m[320]&m[321]&m[322]&m[323]))&~BiasedRNG[224])|((m[18]&m[320]&m[321]&m[322]&~m[323])|(m[18]&m[320]&m[321]&~m[322]&m[323])|(m[18]&m[320]&~m[321]&m[322]&m[323])|(m[18]&~m[320]&m[321]&m[322]&m[323])|(~m[18]&m[320]&m[321]&m[322]&m[323])|(m[18]&m[320]&m[321]&m[322]&m[323]));
    m[81] = (((m[19]&m[324]&~m[325]&~m[326]&~m[327])|(m[19]&~m[324]&m[325]&~m[326]&~m[327])|(~m[19]&m[324]&m[325]&~m[326]&~m[327])|(m[19]&~m[324]&~m[325]&m[326]&~m[327])|(~m[19]&m[324]&~m[325]&m[326]&~m[327])|(~m[19]&~m[324]&m[325]&m[326]&~m[327])|(m[19]&~m[324]&~m[325]&~m[326]&m[327])|(~m[19]&m[324]&~m[325]&~m[326]&m[327])|(~m[19]&~m[324]&m[325]&~m[326]&m[327])|(~m[19]&~m[324]&~m[325]&m[326]&m[327]))&BiasedRNG[225])|(((m[19]&m[324]&m[325]&~m[326]&~m[327])|(m[19]&m[324]&~m[325]&m[326]&~m[327])|(m[19]&~m[324]&m[325]&m[326]&~m[327])|(~m[19]&m[324]&m[325]&m[326]&~m[327])|(m[19]&m[324]&~m[325]&~m[326]&m[327])|(m[19]&~m[324]&m[325]&~m[326]&m[327])|(~m[19]&m[324]&m[325]&~m[326]&m[327])|(m[19]&~m[324]&~m[325]&m[326]&m[327])|(~m[19]&m[324]&~m[325]&m[326]&m[327])|(~m[19]&~m[324]&m[325]&m[326]&m[327]))&~BiasedRNG[225])|((m[19]&m[324]&m[325]&m[326]&~m[327])|(m[19]&m[324]&m[325]&~m[326]&m[327])|(m[19]&m[324]&~m[325]&m[326]&m[327])|(m[19]&~m[324]&m[325]&m[326]&m[327])|(~m[19]&m[324]&m[325]&m[326]&m[327])|(m[19]&m[324]&m[325]&m[326]&m[327]));
    m[82] = (((m[19]&m[328]&~m[329]&~m[330]&~m[331])|(m[19]&~m[328]&m[329]&~m[330]&~m[331])|(~m[19]&m[328]&m[329]&~m[330]&~m[331])|(m[19]&~m[328]&~m[329]&m[330]&~m[331])|(~m[19]&m[328]&~m[329]&m[330]&~m[331])|(~m[19]&~m[328]&m[329]&m[330]&~m[331])|(m[19]&~m[328]&~m[329]&~m[330]&m[331])|(~m[19]&m[328]&~m[329]&~m[330]&m[331])|(~m[19]&~m[328]&m[329]&~m[330]&m[331])|(~m[19]&~m[328]&~m[329]&m[330]&m[331]))&BiasedRNG[226])|(((m[19]&m[328]&m[329]&~m[330]&~m[331])|(m[19]&m[328]&~m[329]&m[330]&~m[331])|(m[19]&~m[328]&m[329]&m[330]&~m[331])|(~m[19]&m[328]&m[329]&m[330]&~m[331])|(m[19]&m[328]&~m[329]&~m[330]&m[331])|(m[19]&~m[328]&m[329]&~m[330]&m[331])|(~m[19]&m[328]&m[329]&~m[330]&m[331])|(m[19]&~m[328]&~m[329]&m[330]&m[331])|(~m[19]&m[328]&~m[329]&m[330]&m[331])|(~m[19]&~m[328]&m[329]&m[330]&m[331]))&~BiasedRNG[226])|((m[19]&m[328]&m[329]&m[330]&~m[331])|(m[19]&m[328]&m[329]&~m[330]&m[331])|(m[19]&m[328]&~m[329]&m[330]&m[331])|(m[19]&~m[328]&m[329]&m[330]&m[331])|(~m[19]&m[328]&m[329]&m[330]&m[331])|(m[19]&m[328]&m[329]&m[330]&m[331]));
    m[83] = (((m[19]&m[332]&~m[333]&~m[334]&~m[335])|(m[19]&~m[332]&m[333]&~m[334]&~m[335])|(~m[19]&m[332]&m[333]&~m[334]&~m[335])|(m[19]&~m[332]&~m[333]&m[334]&~m[335])|(~m[19]&m[332]&~m[333]&m[334]&~m[335])|(~m[19]&~m[332]&m[333]&m[334]&~m[335])|(m[19]&~m[332]&~m[333]&~m[334]&m[335])|(~m[19]&m[332]&~m[333]&~m[334]&m[335])|(~m[19]&~m[332]&m[333]&~m[334]&m[335])|(~m[19]&~m[332]&~m[333]&m[334]&m[335]))&BiasedRNG[227])|(((m[19]&m[332]&m[333]&~m[334]&~m[335])|(m[19]&m[332]&~m[333]&m[334]&~m[335])|(m[19]&~m[332]&m[333]&m[334]&~m[335])|(~m[19]&m[332]&m[333]&m[334]&~m[335])|(m[19]&m[332]&~m[333]&~m[334]&m[335])|(m[19]&~m[332]&m[333]&~m[334]&m[335])|(~m[19]&m[332]&m[333]&~m[334]&m[335])|(m[19]&~m[332]&~m[333]&m[334]&m[335])|(~m[19]&m[332]&~m[333]&m[334]&m[335])|(~m[19]&~m[332]&m[333]&m[334]&m[335]))&~BiasedRNG[227])|((m[19]&m[332]&m[333]&m[334]&~m[335])|(m[19]&m[332]&m[333]&~m[334]&m[335])|(m[19]&m[332]&~m[333]&m[334]&m[335])|(m[19]&~m[332]&m[333]&m[334]&m[335])|(~m[19]&m[332]&m[333]&m[334]&m[335])|(m[19]&m[332]&m[333]&m[334]&m[335]));
    m[84] = (((m[20]&m[336]&~m[337]&~m[338]&~m[339])|(m[20]&~m[336]&m[337]&~m[338]&~m[339])|(~m[20]&m[336]&m[337]&~m[338]&~m[339])|(m[20]&~m[336]&~m[337]&m[338]&~m[339])|(~m[20]&m[336]&~m[337]&m[338]&~m[339])|(~m[20]&~m[336]&m[337]&m[338]&~m[339])|(m[20]&~m[336]&~m[337]&~m[338]&m[339])|(~m[20]&m[336]&~m[337]&~m[338]&m[339])|(~m[20]&~m[336]&m[337]&~m[338]&m[339])|(~m[20]&~m[336]&~m[337]&m[338]&m[339]))&BiasedRNG[228])|(((m[20]&m[336]&m[337]&~m[338]&~m[339])|(m[20]&m[336]&~m[337]&m[338]&~m[339])|(m[20]&~m[336]&m[337]&m[338]&~m[339])|(~m[20]&m[336]&m[337]&m[338]&~m[339])|(m[20]&m[336]&~m[337]&~m[338]&m[339])|(m[20]&~m[336]&m[337]&~m[338]&m[339])|(~m[20]&m[336]&m[337]&~m[338]&m[339])|(m[20]&~m[336]&~m[337]&m[338]&m[339])|(~m[20]&m[336]&~m[337]&m[338]&m[339])|(~m[20]&~m[336]&m[337]&m[338]&m[339]))&~BiasedRNG[228])|((m[20]&m[336]&m[337]&m[338]&~m[339])|(m[20]&m[336]&m[337]&~m[338]&m[339])|(m[20]&m[336]&~m[337]&m[338]&m[339])|(m[20]&~m[336]&m[337]&m[338]&m[339])|(~m[20]&m[336]&m[337]&m[338]&m[339])|(m[20]&m[336]&m[337]&m[338]&m[339]));
    m[85] = (((m[20]&m[340]&~m[341]&~m[342]&~m[343])|(m[20]&~m[340]&m[341]&~m[342]&~m[343])|(~m[20]&m[340]&m[341]&~m[342]&~m[343])|(m[20]&~m[340]&~m[341]&m[342]&~m[343])|(~m[20]&m[340]&~m[341]&m[342]&~m[343])|(~m[20]&~m[340]&m[341]&m[342]&~m[343])|(m[20]&~m[340]&~m[341]&~m[342]&m[343])|(~m[20]&m[340]&~m[341]&~m[342]&m[343])|(~m[20]&~m[340]&m[341]&~m[342]&m[343])|(~m[20]&~m[340]&~m[341]&m[342]&m[343]))&BiasedRNG[229])|(((m[20]&m[340]&m[341]&~m[342]&~m[343])|(m[20]&m[340]&~m[341]&m[342]&~m[343])|(m[20]&~m[340]&m[341]&m[342]&~m[343])|(~m[20]&m[340]&m[341]&m[342]&~m[343])|(m[20]&m[340]&~m[341]&~m[342]&m[343])|(m[20]&~m[340]&m[341]&~m[342]&m[343])|(~m[20]&m[340]&m[341]&~m[342]&m[343])|(m[20]&~m[340]&~m[341]&m[342]&m[343])|(~m[20]&m[340]&~m[341]&m[342]&m[343])|(~m[20]&~m[340]&m[341]&m[342]&m[343]))&~BiasedRNG[229])|((m[20]&m[340]&m[341]&m[342]&~m[343])|(m[20]&m[340]&m[341]&~m[342]&m[343])|(m[20]&m[340]&~m[341]&m[342]&m[343])|(m[20]&~m[340]&m[341]&m[342]&m[343])|(~m[20]&m[340]&m[341]&m[342]&m[343])|(m[20]&m[340]&m[341]&m[342]&m[343]));
    m[86] = (((m[20]&m[344]&~m[345]&~m[346]&~m[347])|(m[20]&~m[344]&m[345]&~m[346]&~m[347])|(~m[20]&m[344]&m[345]&~m[346]&~m[347])|(m[20]&~m[344]&~m[345]&m[346]&~m[347])|(~m[20]&m[344]&~m[345]&m[346]&~m[347])|(~m[20]&~m[344]&m[345]&m[346]&~m[347])|(m[20]&~m[344]&~m[345]&~m[346]&m[347])|(~m[20]&m[344]&~m[345]&~m[346]&m[347])|(~m[20]&~m[344]&m[345]&~m[346]&m[347])|(~m[20]&~m[344]&~m[345]&m[346]&m[347]))&BiasedRNG[230])|(((m[20]&m[344]&m[345]&~m[346]&~m[347])|(m[20]&m[344]&~m[345]&m[346]&~m[347])|(m[20]&~m[344]&m[345]&m[346]&~m[347])|(~m[20]&m[344]&m[345]&m[346]&~m[347])|(m[20]&m[344]&~m[345]&~m[346]&m[347])|(m[20]&~m[344]&m[345]&~m[346]&m[347])|(~m[20]&m[344]&m[345]&~m[346]&m[347])|(m[20]&~m[344]&~m[345]&m[346]&m[347])|(~m[20]&m[344]&~m[345]&m[346]&m[347])|(~m[20]&~m[344]&m[345]&m[346]&m[347]))&~BiasedRNG[230])|((m[20]&m[344]&m[345]&m[346]&~m[347])|(m[20]&m[344]&m[345]&~m[346]&m[347])|(m[20]&m[344]&~m[345]&m[346]&m[347])|(m[20]&~m[344]&m[345]&m[346]&m[347])|(~m[20]&m[344]&m[345]&m[346]&m[347])|(m[20]&m[344]&m[345]&m[346]&m[347]));
    m[87] = (((m[21]&m[348]&~m[349]&~m[350]&~m[351])|(m[21]&~m[348]&m[349]&~m[350]&~m[351])|(~m[21]&m[348]&m[349]&~m[350]&~m[351])|(m[21]&~m[348]&~m[349]&m[350]&~m[351])|(~m[21]&m[348]&~m[349]&m[350]&~m[351])|(~m[21]&~m[348]&m[349]&m[350]&~m[351])|(m[21]&~m[348]&~m[349]&~m[350]&m[351])|(~m[21]&m[348]&~m[349]&~m[350]&m[351])|(~m[21]&~m[348]&m[349]&~m[350]&m[351])|(~m[21]&~m[348]&~m[349]&m[350]&m[351]))&BiasedRNG[231])|(((m[21]&m[348]&m[349]&~m[350]&~m[351])|(m[21]&m[348]&~m[349]&m[350]&~m[351])|(m[21]&~m[348]&m[349]&m[350]&~m[351])|(~m[21]&m[348]&m[349]&m[350]&~m[351])|(m[21]&m[348]&~m[349]&~m[350]&m[351])|(m[21]&~m[348]&m[349]&~m[350]&m[351])|(~m[21]&m[348]&m[349]&~m[350]&m[351])|(m[21]&~m[348]&~m[349]&m[350]&m[351])|(~m[21]&m[348]&~m[349]&m[350]&m[351])|(~m[21]&~m[348]&m[349]&m[350]&m[351]))&~BiasedRNG[231])|((m[21]&m[348]&m[349]&m[350]&~m[351])|(m[21]&m[348]&m[349]&~m[350]&m[351])|(m[21]&m[348]&~m[349]&m[350]&m[351])|(m[21]&~m[348]&m[349]&m[350]&m[351])|(~m[21]&m[348]&m[349]&m[350]&m[351])|(m[21]&m[348]&m[349]&m[350]&m[351]));
    m[88] = (((m[21]&m[352]&~m[353]&~m[354]&~m[355])|(m[21]&~m[352]&m[353]&~m[354]&~m[355])|(~m[21]&m[352]&m[353]&~m[354]&~m[355])|(m[21]&~m[352]&~m[353]&m[354]&~m[355])|(~m[21]&m[352]&~m[353]&m[354]&~m[355])|(~m[21]&~m[352]&m[353]&m[354]&~m[355])|(m[21]&~m[352]&~m[353]&~m[354]&m[355])|(~m[21]&m[352]&~m[353]&~m[354]&m[355])|(~m[21]&~m[352]&m[353]&~m[354]&m[355])|(~m[21]&~m[352]&~m[353]&m[354]&m[355]))&BiasedRNG[232])|(((m[21]&m[352]&m[353]&~m[354]&~m[355])|(m[21]&m[352]&~m[353]&m[354]&~m[355])|(m[21]&~m[352]&m[353]&m[354]&~m[355])|(~m[21]&m[352]&m[353]&m[354]&~m[355])|(m[21]&m[352]&~m[353]&~m[354]&m[355])|(m[21]&~m[352]&m[353]&~m[354]&m[355])|(~m[21]&m[352]&m[353]&~m[354]&m[355])|(m[21]&~m[352]&~m[353]&m[354]&m[355])|(~m[21]&m[352]&~m[353]&m[354]&m[355])|(~m[21]&~m[352]&m[353]&m[354]&m[355]))&~BiasedRNG[232])|((m[21]&m[352]&m[353]&m[354]&~m[355])|(m[21]&m[352]&m[353]&~m[354]&m[355])|(m[21]&m[352]&~m[353]&m[354]&m[355])|(m[21]&~m[352]&m[353]&m[354]&m[355])|(~m[21]&m[352]&m[353]&m[354]&m[355])|(m[21]&m[352]&m[353]&m[354]&m[355]));
    m[89] = (((m[21]&m[356]&~m[357]&~m[358]&~m[359])|(m[21]&~m[356]&m[357]&~m[358]&~m[359])|(~m[21]&m[356]&m[357]&~m[358]&~m[359])|(m[21]&~m[356]&~m[357]&m[358]&~m[359])|(~m[21]&m[356]&~m[357]&m[358]&~m[359])|(~m[21]&~m[356]&m[357]&m[358]&~m[359])|(m[21]&~m[356]&~m[357]&~m[358]&m[359])|(~m[21]&m[356]&~m[357]&~m[358]&m[359])|(~m[21]&~m[356]&m[357]&~m[358]&m[359])|(~m[21]&~m[356]&~m[357]&m[358]&m[359]))&BiasedRNG[233])|(((m[21]&m[356]&m[357]&~m[358]&~m[359])|(m[21]&m[356]&~m[357]&m[358]&~m[359])|(m[21]&~m[356]&m[357]&m[358]&~m[359])|(~m[21]&m[356]&m[357]&m[358]&~m[359])|(m[21]&m[356]&~m[357]&~m[358]&m[359])|(m[21]&~m[356]&m[357]&~m[358]&m[359])|(~m[21]&m[356]&m[357]&~m[358]&m[359])|(m[21]&~m[356]&~m[357]&m[358]&m[359])|(~m[21]&m[356]&~m[357]&m[358]&m[359])|(~m[21]&~m[356]&m[357]&m[358]&m[359]))&~BiasedRNG[233])|((m[21]&m[356]&m[357]&m[358]&~m[359])|(m[21]&m[356]&m[357]&~m[358]&m[359])|(m[21]&m[356]&~m[357]&m[358]&m[359])|(m[21]&~m[356]&m[357]&m[358]&m[359])|(~m[21]&m[356]&m[357]&m[358]&m[359])|(m[21]&m[356]&m[357]&m[358]&m[359]));
    m[90] = (((m[22]&m[360]&~m[361]&~m[362]&~m[363])|(m[22]&~m[360]&m[361]&~m[362]&~m[363])|(~m[22]&m[360]&m[361]&~m[362]&~m[363])|(m[22]&~m[360]&~m[361]&m[362]&~m[363])|(~m[22]&m[360]&~m[361]&m[362]&~m[363])|(~m[22]&~m[360]&m[361]&m[362]&~m[363])|(m[22]&~m[360]&~m[361]&~m[362]&m[363])|(~m[22]&m[360]&~m[361]&~m[362]&m[363])|(~m[22]&~m[360]&m[361]&~m[362]&m[363])|(~m[22]&~m[360]&~m[361]&m[362]&m[363]))&BiasedRNG[234])|(((m[22]&m[360]&m[361]&~m[362]&~m[363])|(m[22]&m[360]&~m[361]&m[362]&~m[363])|(m[22]&~m[360]&m[361]&m[362]&~m[363])|(~m[22]&m[360]&m[361]&m[362]&~m[363])|(m[22]&m[360]&~m[361]&~m[362]&m[363])|(m[22]&~m[360]&m[361]&~m[362]&m[363])|(~m[22]&m[360]&m[361]&~m[362]&m[363])|(m[22]&~m[360]&~m[361]&m[362]&m[363])|(~m[22]&m[360]&~m[361]&m[362]&m[363])|(~m[22]&~m[360]&m[361]&m[362]&m[363]))&~BiasedRNG[234])|((m[22]&m[360]&m[361]&m[362]&~m[363])|(m[22]&m[360]&m[361]&~m[362]&m[363])|(m[22]&m[360]&~m[361]&m[362]&m[363])|(m[22]&~m[360]&m[361]&m[362]&m[363])|(~m[22]&m[360]&m[361]&m[362]&m[363])|(m[22]&m[360]&m[361]&m[362]&m[363]));
    m[91] = (((m[22]&m[364]&~m[365]&~m[366]&~m[367])|(m[22]&~m[364]&m[365]&~m[366]&~m[367])|(~m[22]&m[364]&m[365]&~m[366]&~m[367])|(m[22]&~m[364]&~m[365]&m[366]&~m[367])|(~m[22]&m[364]&~m[365]&m[366]&~m[367])|(~m[22]&~m[364]&m[365]&m[366]&~m[367])|(m[22]&~m[364]&~m[365]&~m[366]&m[367])|(~m[22]&m[364]&~m[365]&~m[366]&m[367])|(~m[22]&~m[364]&m[365]&~m[366]&m[367])|(~m[22]&~m[364]&~m[365]&m[366]&m[367]))&BiasedRNG[235])|(((m[22]&m[364]&m[365]&~m[366]&~m[367])|(m[22]&m[364]&~m[365]&m[366]&~m[367])|(m[22]&~m[364]&m[365]&m[366]&~m[367])|(~m[22]&m[364]&m[365]&m[366]&~m[367])|(m[22]&m[364]&~m[365]&~m[366]&m[367])|(m[22]&~m[364]&m[365]&~m[366]&m[367])|(~m[22]&m[364]&m[365]&~m[366]&m[367])|(m[22]&~m[364]&~m[365]&m[366]&m[367])|(~m[22]&m[364]&~m[365]&m[366]&m[367])|(~m[22]&~m[364]&m[365]&m[366]&m[367]))&~BiasedRNG[235])|((m[22]&m[364]&m[365]&m[366]&~m[367])|(m[22]&m[364]&m[365]&~m[366]&m[367])|(m[22]&m[364]&~m[365]&m[366]&m[367])|(m[22]&~m[364]&m[365]&m[366]&m[367])|(~m[22]&m[364]&m[365]&m[366]&m[367])|(m[22]&m[364]&m[365]&m[366]&m[367]));
    m[92] = (((m[22]&m[368]&~m[369]&~m[370]&~m[371])|(m[22]&~m[368]&m[369]&~m[370]&~m[371])|(~m[22]&m[368]&m[369]&~m[370]&~m[371])|(m[22]&~m[368]&~m[369]&m[370]&~m[371])|(~m[22]&m[368]&~m[369]&m[370]&~m[371])|(~m[22]&~m[368]&m[369]&m[370]&~m[371])|(m[22]&~m[368]&~m[369]&~m[370]&m[371])|(~m[22]&m[368]&~m[369]&~m[370]&m[371])|(~m[22]&~m[368]&m[369]&~m[370]&m[371])|(~m[22]&~m[368]&~m[369]&m[370]&m[371]))&BiasedRNG[236])|(((m[22]&m[368]&m[369]&~m[370]&~m[371])|(m[22]&m[368]&~m[369]&m[370]&~m[371])|(m[22]&~m[368]&m[369]&m[370]&~m[371])|(~m[22]&m[368]&m[369]&m[370]&~m[371])|(m[22]&m[368]&~m[369]&~m[370]&m[371])|(m[22]&~m[368]&m[369]&~m[370]&m[371])|(~m[22]&m[368]&m[369]&~m[370]&m[371])|(m[22]&~m[368]&~m[369]&m[370]&m[371])|(~m[22]&m[368]&~m[369]&m[370]&m[371])|(~m[22]&~m[368]&m[369]&m[370]&m[371]))&~BiasedRNG[236])|((m[22]&m[368]&m[369]&m[370]&~m[371])|(m[22]&m[368]&m[369]&~m[370]&m[371])|(m[22]&m[368]&~m[369]&m[370]&m[371])|(m[22]&~m[368]&m[369]&m[370]&m[371])|(~m[22]&m[368]&m[369]&m[370]&m[371])|(m[22]&m[368]&m[369]&m[370]&m[371]));
    m[93] = (((m[23]&m[372]&~m[373]&~m[374]&~m[375])|(m[23]&~m[372]&m[373]&~m[374]&~m[375])|(~m[23]&m[372]&m[373]&~m[374]&~m[375])|(m[23]&~m[372]&~m[373]&m[374]&~m[375])|(~m[23]&m[372]&~m[373]&m[374]&~m[375])|(~m[23]&~m[372]&m[373]&m[374]&~m[375])|(m[23]&~m[372]&~m[373]&~m[374]&m[375])|(~m[23]&m[372]&~m[373]&~m[374]&m[375])|(~m[23]&~m[372]&m[373]&~m[374]&m[375])|(~m[23]&~m[372]&~m[373]&m[374]&m[375]))&BiasedRNG[237])|(((m[23]&m[372]&m[373]&~m[374]&~m[375])|(m[23]&m[372]&~m[373]&m[374]&~m[375])|(m[23]&~m[372]&m[373]&m[374]&~m[375])|(~m[23]&m[372]&m[373]&m[374]&~m[375])|(m[23]&m[372]&~m[373]&~m[374]&m[375])|(m[23]&~m[372]&m[373]&~m[374]&m[375])|(~m[23]&m[372]&m[373]&~m[374]&m[375])|(m[23]&~m[372]&~m[373]&m[374]&m[375])|(~m[23]&m[372]&~m[373]&m[374]&m[375])|(~m[23]&~m[372]&m[373]&m[374]&m[375]))&~BiasedRNG[237])|((m[23]&m[372]&m[373]&m[374]&~m[375])|(m[23]&m[372]&m[373]&~m[374]&m[375])|(m[23]&m[372]&~m[373]&m[374]&m[375])|(m[23]&~m[372]&m[373]&m[374]&m[375])|(~m[23]&m[372]&m[373]&m[374]&m[375])|(m[23]&m[372]&m[373]&m[374]&m[375]));
    m[94] = (((m[23]&m[376]&~m[377]&~m[378]&~m[379])|(m[23]&~m[376]&m[377]&~m[378]&~m[379])|(~m[23]&m[376]&m[377]&~m[378]&~m[379])|(m[23]&~m[376]&~m[377]&m[378]&~m[379])|(~m[23]&m[376]&~m[377]&m[378]&~m[379])|(~m[23]&~m[376]&m[377]&m[378]&~m[379])|(m[23]&~m[376]&~m[377]&~m[378]&m[379])|(~m[23]&m[376]&~m[377]&~m[378]&m[379])|(~m[23]&~m[376]&m[377]&~m[378]&m[379])|(~m[23]&~m[376]&~m[377]&m[378]&m[379]))&BiasedRNG[238])|(((m[23]&m[376]&m[377]&~m[378]&~m[379])|(m[23]&m[376]&~m[377]&m[378]&~m[379])|(m[23]&~m[376]&m[377]&m[378]&~m[379])|(~m[23]&m[376]&m[377]&m[378]&~m[379])|(m[23]&m[376]&~m[377]&~m[378]&m[379])|(m[23]&~m[376]&m[377]&~m[378]&m[379])|(~m[23]&m[376]&m[377]&~m[378]&m[379])|(m[23]&~m[376]&~m[377]&m[378]&m[379])|(~m[23]&m[376]&~m[377]&m[378]&m[379])|(~m[23]&~m[376]&m[377]&m[378]&m[379]))&~BiasedRNG[238])|((m[23]&m[376]&m[377]&m[378]&~m[379])|(m[23]&m[376]&m[377]&~m[378]&m[379])|(m[23]&m[376]&~m[377]&m[378]&m[379])|(m[23]&~m[376]&m[377]&m[378]&m[379])|(~m[23]&m[376]&m[377]&m[378]&m[379])|(m[23]&m[376]&m[377]&m[378]&m[379]));
    m[95] = (((m[23]&m[380]&~m[381]&~m[382]&~m[383])|(m[23]&~m[380]&m[381]&~m[382]&~m[383])|(~m[23]&m[380]&m[381]&~m[382]&~m[383])|(m[23]&~m[380]&~m[381]&m[382]&~m[383])|(~m[23]&m[380]&~m[381]&m[382]&~m[383])|(~m[23]&~m[380]&m[381]&m[382]&~m[383])|(m[23]&~m[380]&~m[381]&~m[382]&m[383])|(~m[23]&m[380]&~m[381]&~m[382]&m[383])|(~m[23]&~m[380]&m[381]&~m[382]&m[383])|(~m[23]&~m[380]&~m[381]&m[382]&m[383]))&BiasedRNG[239])|(((m[23]&m[380]&m[381]&~m[382]&~m[383])|(m[23]&m[380]&~m[381]&m[382]&~m[383])|(m[23]&~m[380]&m[381]&m[382]&~m[383])|(~m[23]&m[380]&m[381]&m[382]&~m[383])|(m[23]&m[380]&~m[381]&~m[382]&m[383])|(m[23]&~m[380]&m[381]&~m[382]&m[383])|(~m[23]&m[380]&m[381]&~m[382]&m[383])|(m[23]&~m[380]&~m[381]&m[382]&m[383])|(~m[23]&m[380]&~m[381]&m[382]&m[383])|(~m[23]&~m[380]&m[381]&m[382]&m[383]))&~BiasedRNG[239])|((m[23]&m[380]&m[381]&m[382]&~m[383])|(m[23]&m[380]&m[381]&~m[382]&m[383])|(m[23]&m[380]&~m[381]&m[382]&m[383])|(m[23]&~m[380]&m[381]&m[382]&m[383])|(~m[23]&m[380]&m[381]&m[382]&m[383])|(m[23]&m[380]&m[381]&m[382]&m[383]));
    m[385] = (((m[108]&~m[241]&m[528])|(~m[108]&m[241]&m[528]))&BiasedRNG[240])|(((m[108]&m[241]&~m[528]))&~BiasedRNG[240])|((m[108]&m[241]&m[528]));
    m[386] = (((m[120]&~m[242]&m[533])|(~m[120]&m[242]&m[533]))&BiasedRNG[241])|(((m[120]&m[242]&~m[533]))&~BiasedRNG[241])|((m[120]&m[242]&m[533]));
    m[387] = (((m[132]&~m[243]&m[543])|(~m[132]&m[243]&m[543]))&BiasedRNG[242])|(((m[132]&m[243]&~m[543]))&~BiasedRNG[242])|((m[132]&m[243]&m[543]));
    m[388] = (((m[144]&~m[244]&m[558])|(~m[144]&m[244]&m[558]))&BiasedRNG[243])|(((m[144]&m[244]&~m[558]))&~BiasedRNG[243])|((m[144]&m[244]&m[558]));
    m[389] = (((m[156]&~m[245]&m[578])|(~m[156]&m[245]&m[578]))&BiasedRNG[244])|(((m[156]&m[245]&~m[578]))&~BiasedRNG[244])|((m[156]&m[245]&m[578]));
    m[390] = (((m[168]&~m[246]&m[603])|(~m[168]&m[246]&m[603]))&BiasedRNG[245])|(((m[168]&m[246]&~m[603]))&~BiasedRNG[245])|((m[168]&m[246]&m[603]));
    m[391] = (((m[180]&~m[247]&m[633])|(~m[180]&m[247]&m[633]))&BiasedRNG[246])|(((m[180]&m[247]&~m[633]))&~BiasedRNG[246])|((m[180]&m[247]&m[633]));
    m[392] = (((m[192]&~m[248]&m[668])|(~m[192]&m[248]&m[668]))&BiasedRNG[247])|(((m[192]&m[248]&~m[668]))&~BiasedRNG[247])|((m[192]&m[248]&m[668]));
    m[393] = (((m[204]&~m[249]&m[708])|(~m[204]&m[249]&m[708]))&BiasedRNG[248])|(((m[204]&m[249]&~m[708]))&~BiasedRNG[248])|((m[204]&m[249]&m[708]));
    m[394] = (((m[216]&~m[250]&m[753])|(~m[216]&m[250]&m[753]))&BiasedRNG[249])|(((m[216]&m[250]&~m[753]))&~BiasedRNG[249])|((m[216]&m[250]&m[753]));
    m[395] = (((m[228]&~m[251]&m[803])|(~m[228]&m[251]&m[803]))&BiasedRNG[250])|(((m[228]&m[251]&~m[803]))&~BiasedRNG[250])|((m[228]&m[251]&m[803]));
    m[396] = (((m[97]&~m[252]&m[529])|(~m[97]&m[252]&m[529]))&BiasedRNG[251])|(((m[97]&m[252]&~m[529]))&~BiasedRNG[251])|((m[97]&m[252]&m[529]));
    m[397] = (((m[109]&~m[253]&m[534])|(~m[109]&m[253]&m[534]))&BiasedRNG[252])|(((m[109]&m[253]&~m[534]))&~BiasedRNG[252])|((m[109]&m[253]&m[534]));
    m[398] = (((m[121]&~m[254]&m[544])|(~m[121]&m[254]&m[544]))&BiasedRNG[253])|(((m[121]&m[254]&~m[544]))&~BiasedRNG[253])|((m[121]&m[254]&m[544]));
    m[399] = (((m[133]&~m[255]&m[559])|(~m[133]&m[255]&m[559]))&BiasedRNG[254])|(((m[133]&m[255]&~m[559]))&~BiasedRNG[254])|((m[133]&m[255]&m[559]));
    m[400] = (((m[145]&~m[256]&m[579])|(~m[145]&m[256]&m[579]))&BiasedRNG[255])|(((m[145]&m[256]&~m[579]))&~BiasedRNG[255])|((m[145]&m[256]&m[579]));
    m[401] = (((m[157]&~m[257]&m[604])|(~m[157]&m[257]&m[604]))&BiasedRNG[256])|(((m[157]&m[257]&~m[604]))&~BiasedRNG[256])|((m[157]&m[257]&m[604]));
    m[402] = (((m[169]&~m[258]&m[634])|(~m[169]&m[258]&m[634]))&BiasedRNG[257])|(((m[169]&m[258]&~m[634]))&~BiasedRNG[257])|((m[169]&m[258]&m[634]));
    m[403] = (((m[181]&~m[259]&m[669])|(~m[181]&m[259]&m[669]))&BiasedRNG[258])|(((m[181]&m[259]&~m[669]))&~BiasedRNG[258])|((m[181]&m[259]&m[669]));
    m[404] = (((m[193]&~m[260]&m[709])|(~m[193]&m[260]&m[709]))&BiasedRNG[259])|(((m[193]&m[260]&~m[709]))&~BiasedRNG[259])|((m[193]&m[260]&m[709]));
    m[405] = (((m[205]&~m[261]&m[754])|(~m[205]&m[261]&m[754]))&BiasedRNG[260])|(((m[205]&m[261]&~m[754]))&~BiasedRNG[260])|((m[205]&m[261]&m[754]));
    m[406] = (((m[217]&~m[262]&m[804])|(~m[217]&m[262]&m[804]))&BiasedRNG[261])|(((m[217]&m[262]&~m[804]))&~BiasedRNG[261])|((m[217]&m[262]&m[804]));
    m[407] = (((m[229]&~m[263]&m[859])|(~m[229]&m[263]&m[859]))&BiasedRNG[262])|(((m[229]&m[263]&~m[859]))&~BiasedRNG[262])|((m[229]&m[263]&m[859]));
    m[408] = (((m[98]&~m[264]&m[539])|(~m[98]&m[264]&m[539]))&BiasedRNG[263])|(((m[98]&m[264]&~m[539]))&~BiasedRNG[263])|((m[98]&m[264]&m[539]));
    m[409] = (((m[110]&~m[265]&m[549])|(~m[110]&m[265]&m[549]))&BiasedRNG[264])|(((m[110]&m[265]&~m[549]))&~BiasedRNG[264])|((m[110]&m[265]&m[549]));
    m[410] = (((m[122]&~m[266]&m[564])|(~m[122]&m[266]&m[564]))&BiasedRNG[265])|(((m[122]&m[266]&~m[564]))&~BiasedRNG[265])|((m[122]&m[266]&m[564]));
    m[411] = (((m[134]&~m[267]&m[584])|(~m[134]&m[267]&m[584]))&BiasedRNG[266])|(((m[134]&m[267]&~m[584]))&~BiasedRNG[266])|((m[134]&m[267]&m[584]));
    m[412] = (((m[146]&~m[268]&m[609])|(~m[146]&m[268]&m[609]))&BiasedRNG[267])|(((m[146]&m[268]&~m[609]))&~BiasedRNG[267])|((m[146]&m[268]&m[609]));
    m[413] = (((m[158]&~m[269]&m[639])|(~m[158]&m[269]&m[639]))&BiasedRNG[268])|(((m[158]&m[269]&~m[639]))&~BiasedRNG[268])|((m[158]&m[269]&m[639]));
    m[414] = (((m[170]&~m[270]&m[674])|(~m[170]&m[270]&m[674]))&BiasedRNG[269])|(((m[170]&m[270]&~m[674]))&~BiasedRNG[269])|((m[170]&m[270]&m[674]));
    m[415] = (((m[182]&~m[271]&m[714])|(~m[182]&m[271]&m[714]))&BiasedRNG[270])|(((m[182]&m[271]&~m[714]))&~BiasedRNG[270])|((m[182]&m[271]&m[714]));
    m[416] = (((m[194]&~m[272]&m[759])|(~m[194]&m[272]&m[759]))&BiasedRNG[271])|(((m[194]&m[272]&~m[759]))&~BiasedRNG[271])|((m[194]&m[272]&m[759]));
    m[417] = (((m[206]&~m[273]&m[809])|(~m[206]&m[273]&m[809]))&BiasedRNG[272])|(((m[206]&m[273]&~m[809]))&~BiasedRNG[272])|((m[206]&m[273]&m[809]));
    m[418] = (((m[218]&~m[274]&m[864])|(~m[218]&m[274]&m[864]))&BiasedRNG[273])|(((m[218]&m[274]&~m[864]))&~BiasedRNG[273])|((m[218]&m[274]&m[864]));
    m[419] = (((m[230]&~m[275]&m[914])|(~m[230]&m[275]&m[914]))&BiasedRNG[274])|(((m[230]&m[275]&~m[914]))&~BiasedRNG[274])|((m[230]&m[275]&m[914]));
    m[420] = (((m[99]&~m[276]&m[554])|(~m[99]&m[276]&m[554]))&BiasedRNG[275])|(((m[99]&m[276]&~m[554]))&~BiasedRNG[275])|((m[99]&m[276]&m[554]));
    m[421] = (((m[111]&~m[277]&m[569])|(~m[111]&m[277]&m[569]))&BiasedRNG[276])|(((m[111]&m[277]&~m[569]))&~BiasedRNG[276])|((m[111]&m[277]&m[569]));
    m[422] = (((m[123]&~m[278]&m[589])|(~m[123]&m[278]&m[589]))&BiasedRNG[277])|(((m[123]&m[278]&~m[589]))&~BiasedRNG[277])|((m[123]&m[278]&m[589]));
    m[423] = (((m[135]&~m[279]&m[614])|(~m[135]&m[279]&m[614]))&BiasedRNG[278])|(((m[135]&m[279]&~m[614]))&~BiasedRNG[278])|((m[135]&m[279]&m[614]));
    m[424] = (((m[147]&~m[280]&m[644])|(~m[147]&m[280]&m[644]))&BiasedRNG[279])|(((m[147]&m[280]&~m[644]))&~BiasedRNG[279])|((m[147]&m[280]&m[644]));
    m[425] = (((m[159]&~m[281]&m[679])|(~m[159]&m[281]&m[679]))&BiasedRNG[280])|(((m[159]&m[281]&~m[679]))&~BiasedRNG[280])|((m[159]&m[281]&m[679]));
    m[426] = (((m[171]&~m[282]&m[719])|(~m[171]&m[282]&m[719]))&BiasedRNG[281])|(((m[171]&m[282]&~m[719]))&~BiasedRNG[281])|((m[171]&m[282]&m[719]));
    m[427] = (((m[183]&~m[283]&m[764])|(~m[183]&m[283]&m[764]))&BiasedRNG[282])|(((m[183]&m[283]&~m[764]))&~BiasedRNG[282])|((m[183]&m[283]&m[764]));
    m[428] = (((m[195]&~m[284]&m[814])|(~m[195]&m[284]&m[814]))&BiasedRNG[283])|(((m[195]&m[284]&~m[814]))&~BiasedRNG[283])|((m[195]&m[284]&m[814]));
    m[429] = (((m[207]&~m[285]&m[869])|(~m[207]&m[285]&m[869]))&BiasedRNG[284])|(((m[207]&m[285]&~m[869]))&~BiasedRNG[284])|((m[207]&m[285]&m[869]));
    m[430] = (((m[219]&~m[286]&m[919])|(~m[219]&m[286]&m[919]))&BiasedRNG[285])|(((m[219]&m[286]&~m[919]))&~BiasedRNG[285])|((m[219]&m[286]&m[919]));
    m[431] = (((m[231]&~m[287]&m[964])|(~m[231]&m[287]&m[964]))&BiasedRNG[286])|(((m[231]&m[287]&~m[964]))&~BiasedRNG[286])|((m[231]&m[287]&m[964]));
    m[432] = (((m[100]&~m[288]&m[574])|(~m[100]&m[288]&m[574]))&BiasedRNG[287])|(((m[100]&m[288]&~m[574]))&~BiasedRNG[287])|((m[100]&m[288]&m[574]));
    m[433] = (((m[112]&~m[289]&m[594])|(~m[112]&m[289]&m[594]))&BiasedRNG[288])|(((m[112]&m[289]&~m[594]))&~BiasedRNG[288])|((m[112]&m[289]&m[594]));
    m[434] = (((m[124]&~m[290]&m[619])|(~m[124]&m[290]&m[619]))&BiasedRNG[289])|(((m[124]&m[290]&~m[619]))&~BiasedRNG[289])|((m[124]&m[290]&m[619]));
    m[435] = (((m[136]&~m[291]&m[649])|(~m[136]&m[291]&m[649]))&BiasedRNG[290])|(((m[136]&m[291]&~m[649]))&~BiasedRNG[290])|((m[136]&m[291]&m[649]));
    m[436] = (((m[148]&~m[292]&m[684])|(~m[148]&m[292]&m[684]))&BiasedRNG[291])|(((m[148]&m[292]&~m[684]))&~BiasedRNG[291])|((m[148]&m[292]&m[684]));
    m[437] = (((m[160]&~m[293]&m[724])|(~m[160]&m[293]&m[724]))&BiasedRNG[292])|(((m[160]&m[293]&~m[724]))&~BiasedRNG[292])|((m[160]&m[293]&m[724]));
    m[438] = (((m[172]&~m[294]&m[769])|(~m[172]&m[294]&m[769]))&BiasedRNG[293])|(((m[172]&m[294]&~m[769]))&~BiasedRNG[293])|((m[172]&m[294]&m[769]));
    m[439] = (((m[184]&~m[295]&m[819])|(~m[184]&m[295]&m[819]))&BiasedRNG[294])|(((m[184]&m[295]&~m[819]))&~BiasedRNG[294])|((m[184]&m[295]&m[819]));
    m[440] = (((m[196]&~m[296]&m[874])|(~m[196]&m[296]&m[874]))&BiasedRNG[295])|(((m[196]&m[296]&~m[874]))&~BiasedRNG[295])|((m[196]&m[296]&m[874]));
    m[441] = (((m[208]&~m[297]&m[924])|(~m[208]&m[297]&m[924]))&BiasedRNG[296])|(((m[208]&m[297]&~m[924]))&~BiasedRNG[296])|((m[208]&m[297]&m[924]));
    m[442] = (((m[220]&~m[298]&m[969])|(~m[220]&m[298]&m[969]))&BiasedRNG[297])|(((m[220]&m[298]&~m[969]))&~BiasedRNG[297])|((m[220]&m[298]&m[969]));
    m[443] = (((m[232]&~m[299]&m[1009])|(~m[232]&m[299]&m[1009]))&BiasedRNG[298])|(((m[232]&m[299]&~m[1009]))&~BiasedRNG[298])|((m[232]&m[299]&m[1009]));
    m[444] = (((m[101]&~m[300]&m[599])|(~m[101]&m[300]&m[599]))&BiasedRNG[299])|(((m[101]&m[300]&~m[599]))&~BiasedRNG[299])|((m[101]&m[300]&m[599]));
    m[445] = (((m[113]&~m[301]&m[624])|(~m[113]&m[301]&m[624]))&BiasedRNG[300])|(((m[113]&m[301]&~m[624]))&~BiasedRNG[300])|((m[113]&m[301]&m[624]));
    m[446] = (((m[125]&~m[302]&m[654])|(~m[125]&m[302]&m[654]))&BiasedRNG[301])|(((m[125]&m[302]&~m[654]))&~BiasedRNG[301])|((m[125]&m[302]&m[654]));
    m[447] = (((m[137]&~m[303]&m[689])|(~m[137]&m[303]&m[689]))&BiasedRNG[302])|(((m[137]&m[303]&~m[689]))&~BiasedRNG[302])|((m[137]&m[303]&m[689]));
    m[448] = (((m[149]&~m[304]&m[729])|(~m[149]&m[304]&m[729]))&BiasedRNG[303])|(((m[149]&m[304]&~m[729]))&~BiasedRNG[303])|((m[149]&m[304]&m[729]));
    m[449] = (((m[161]&~m[305]&m[774])|(~m[161]&m[305]&m[774]))&BiasedRNG[304])|(((m[161]&m[305]&~m[774]))&~BiasedRNG[304])|((m[161]&m[305]&m[774]));
    m[450] = (((m[173]&~m[306]&m[824])|(~m[173]&m[306]&m[824]))&BiasedRNG[305])|(((m[173]&m[306]&~m[824]))&~BiasedRNG[305])|((m[173]&m[306]&m[824]));
    m[451] = (((m[185]&~m[307]&m[879])|(~m[185]&m[307]&m[879]))&BiasedRNG[306])|(((m[185]&m[307]&~m[879]))&~BiasedRNG[306])|((m[185]&m[307]&m[879]));
    m[452] = (((m[197]&~m[308]&m[929])|(~m[197]&m[308]&m[929]))&BiasedRNG[307])|(((m[197]&m[308]&~m[929]))&~BiasedRNG[307])|((m[197]&m[308]&m[929]));
    m[453] = (((m[209]&~m[309]&m[974])|(~m[209]&m[309]&m[974]))&BiasedRNG[308])|(((m[209]&m[309]&~m[974]))&~BiasedRNG[308])|((m[209]&m[309]&m[974]));
    m[454] = (((m[221]&~m[310]&m[1014])|(~m[221]&m[310]&m[1014]))&BiasedRNG[309])|(((m[221]&m[310]&~m[1014]))&~BiasedRNG[309])|((m[221]&m[310]&m[1014]));
    m[455] = (((m[233]&~m[311]&m[1049])|(~m[233]&m[311]&m[1049]))&BiasedRNG[310])|(((m[233]&m[311]&~m[1049]))&~BiasedRNG[310])|((m[233]&m[311]&m[1049]));
    m[456] = (((m[102]&~m[312]&m[629])|(~m[102]&m[312]&m[629]))&BiasedRNG[311])|(((m[102]&m[312]&~m[629]))&~BiasedRNG[311])|((m[102]&m[312]&m[629]));
    m[457] = (((m[114]&~m[313]&m[659])|(~m[114]&m[313]&m[659]))&BiasedRNG[312])|(((m[114]&m[313]&~m[659]))&~BiasedRNG[312])|((m[114]&m[313]&m[659]));
    m[458] = (((m[126]&~m[314]&m[694])|(~m[126]&m[314]&m[694]))&BiasedRNG[313])|(((m[126]&m[314]&~m[694]))&~BiasedRNG[313])|((m[126]&m[314]&m[694]));
    m[459] = (((m[138]&~m[315]&m[734])|(~m[138]&m[315]&m[734]))&BiasedRNG[314])|(((m[138]&m[315]&~m[734]))&~BiasedRNG[314])|((m[138]&m[315]&m[734]));
    m[460] = (((m[150]&~m[316]&m[779])|(~m[150]&m[316]&m[779]))&BiasedRNG[315])|(((m[150]&m[316]&~m[779]))&~BiasedRNG[315])|((m[150]&m[316]&m[779]));
    m[461] = (((m[162]&~m[317]&m[829])|(~m[162]&m[317]&m[829]))&BiasedRNG[316])|(((m[162]&m[317]&~m[829]))&~BiasedRNG[316])|((m[162]&m[317]&m[829]));
    m[462] = (((m[174]&~m[318]&m[884])|(~m[174]&m[318]&m[884]))&BiasedRNG[317])|(((m[174]&m[318]&~m[884]))&~BiasedRNG[317])|((m[174]&m[318]&m[884]));
    m[463] = (((m[186]&~m[319]&m[934])|(~m[186]&m[319]&m[934]))&BiasedRNG[318])|(((m[186]&m[319]&~m[934]))&~BiasedRNG[318])|((m[186]&m[319]&m[934]));
    m[464] = (((m[198]&~m[320]&m[979])|(~m[198]&m[320]&m[979]))&BiasedRNG[319])|(((m[198]&m[320]&~m[979]))&~BiasedRNG[319])|((m[198]&m[320]&m[979]));
    m[465] = (((m[210]&~m[321]&m[1019])|(~m[210]&m[321]&m[1019]))&BiasedRNG[320])|(((m[210]&m[321]&~m[1019]))&~BiasedRNG[320])|((m[210]&m[321]&m[1019]));
    m[466] = (((m[222]&~m[322]&m[1054])|(~m[222]&m[322]&m[1054]))&BiasedRNG[321])|(((m[222]&m[322]&~m[1054]))&~BiasedRNG[321])|((m[222]&m[322]&m[1054]));
    m[467] = (((m[234]&~m[323]&m[1084])|(~m[234]&m[323]&m[1084]))&BiasedRNG[322])|(((m[234]&m[323]&~m[1084]))&~BiasedRNG[322])|((m[234]&m[323]&m[1084]));
    m[468] = (((m[103]&~m[324]&m[664])|(~m[103]&m[324]&m[664]))&BiasedRNG[323])|(((m[103]&m[324]&~m[664]))&~BiasedRNG[323])|((m[103]&m[324]&m[664]));
    m[469] = (((m[115]&~m[325]&m[699])|(~m[115]&m[325]&m[699]))&BiasedRNG[324])|(((m[115]&m[325]&~m[699]))&~BiasedRNG[324])|((m[115]&m[325]&m[699]));
    m[470] = (((m[127]&~m[326]&m[739])|(~m[127]&m[326]&m[739]))&BiasedRNG[325])|(((m[127]&m[326]&~m[739]))&~BiasedRNG[325])|((m[127]&m[326]&m[739]));
    m[471] = (((m[139]&~m[327]&m[784])|(~m[139]&m[327]&m[784]))&BiasedRNG[326])|(((m[139]&m[327]&~m[784]))&~BiasedRNG[326])|((m[139]&m[327]&m[784]));
    m[472] = (((m[151]&~m[328]&m[834])|(~m[151]&m[328]&m[834]))&BiasedRNG[327])|(((m[151]&m[328]&~m[834]))&~BiasedRNG[327])|((m[151]&m[328]&m[834]));
    m[473] = (((m[163]&~m[329]&m[889])|(~m[163]&m[329]&m[889]))&BiasedRNG[328])|(((m[163]&m[329]&~m[889]))&~BiasedRNG[328])|((m[163]&m[329]&m[889]));
    m[474] = (((m[175]&~m[330]&m[939])|(~m[175]&m[330]&m[939]))&BiasedRNG[329])|(((m[175]&m[330]&~m[939]))&~BiasedRNG[329])|((m[175]&m[330]&m[939]));
    m[475] = (((m[187]&~m[331]&m[984])|(~m[187]&m[331]&m[984]))&BiasedRNG[330])|(((m[187]&m[331]&~m[984]))&~BiasedRNG[330])|((m[187]&m[331]&m[984]));
    m[476] = (((m[199]&~m[332]&m[1024])|(~m[199]&m[332]&m[1024]))&BiasedRNG[331])|(((m[199]&m[332]&~m[1024]))&~BiasedRNG[331])|((m[199]&m[332]&m[1024]));
    m[477] = (((m[211]&~m[333]&m[1059])|(~m[211]&m[333]&m[1059]))&BiasedRNG[332])|(((m[211]&m[333]&~m[1059]))&~BiasedRNG[332])|((m[211]&m[333]&m[1059]));
    m[478] = (((m[223]&~m[334]&m[1089])|(~m[223]&m[334]&m[1089]))&BiasedRNG[333])|(((m[223]&m[334]&~m[1089]))&~BiasedRNG[333])|((m[223]&m[334]&m[1089]));
    m[479] = (((m[235]&~m[335]&m[1114])|(~m[235]&m[335]&m[1114]))&BiasedRNG[334])|(((m[235]&m[335]&~m[1114]))&~BiasedRNG[334])|((m[235]&m[335]&m[1114]));
    m[480] = (((m[104]&~m[336]&m[704])|(~m[104]&m[336]&m[704]))&BiasedRNG[335])|(((m[104]&m[336]&~m[704]))&~BiasedRNG[335])|((m[104]&m[336]&m[704]));
    m[481] = (((m[116]&~m[337]&m[744])|(~m[116]&m[337]&m[744]))&BiasedRNG[336])|(((m[116]&m[337]&~m[744]))&~BiasedRNG[336])|((m[116]&m[337]&m[744]));
    m[482] = (((m[128]&~m[338]&m[789])|(~m[128]&m[338]&m[789]))&BiasedRNG[337])|(((m[128]&m[338]&~m[789]))&~BiasedRNG[337])|((m[128]&m[338]&m[789]));
    m[483] = (((m[140]&~m[339]&m[839])|(~m[140]&m[339]&m[839]))&BiasedRNG[338])|(((m[140]&m[339]&~m[839]))&~BiasedRNG[338])|((m[140]&m[339]&m[839]));
    m[484] = (((m[152]&~m[340]&m[894])|(~m[152]&m[340]&m[894]))&BiasedRNG[339])|(((m[152]&m[340]&~m[894]))&~BiasedRNG[339])|((m[152]&m[340]&m[894]));
    m[485] = (((m[164]&~m[341]&m[944])|(~m[164]&m[341]&m[944]))&BiasedRNG[340])|(((m[164]&m[341]&~m[944]))&~BiasedRNG[340])|((m[164]&m[341]&m[944]));
    m[486] = (((m[176]&~m[342]&m[989])|(~m[176]&m[342]&m[989]))&BiasedRNG[341])|(((m[176]&m[342]&~m[989]))&~BiasedRNG[341])|((m[176]&m[342]&m[989]));
    m[487] = (((m[188]&~m[343]&m[1029])|(~m[188]&m[343]&m[1029]))&BiasedRNG[342])|(((m[188]&m[343]&~m[1029]))&~BiasedRNG[342])|((m[188]&m[343]&m[1029]));
    m[488] = (((m[200]&~m[344]&m[1064])|(~m[200]&m[344]&m[1064]))&BiasedRNG[343])|(((m[200]&m[344]&~m[1064]))&~BiasedRNG[343])|((m[200]&m[344]&m[1064]));
    m[489] = (((m[212]&~m[345]&m[1094])|(~m[212]&m[345]&m[1094]))&BiasedRNG[344])|(((m[212]&m[345]&~m[1094]))&~BiasedRNG[344])|((m[212]&m[345]&m[1094]));
    m[490] = (((m[224]&~m[346]&m[1119])|(~m[224]&m[346]&m[1119]))&BiasedRNG[345])|(((m[224]&m[346]&~m[1119]))&~BiasedRNG[345])|((m[224]&m[346]&m[1119]));
    m[491] = (((m[236]&~m[347]&m[1139])|(~m[236]&m[347]&m[1139]))&BiasedRNG[346])|(((m[236]&m[347]&~m[1139]))&~BiasedRNG[346])|((m[236]&m[347]&m[1139]));
    m[492] = (((m[105]&~m[348]&m[749])|(~m[105]&m[348]&m[749]))&BiasedRNG[347])|(((m[105]&m[348]&~m[749]))&~BiasedRNG[347])|((m[105]&m[348]&m[749]));
    m[493] = (((m[117]&~m[349]&m[794])|(~m[117]&m[349]&m[794]))&BiasedRNG[348])|(((m[117]&m[349]&~m[794]))&~BiasedRNG[348])|((m[117]&m[349]&m[794]));
    m[494] = (((m[129]&~m[350]&m[844])|(~m[129]&m[350]&m[844]))&BiasedRNG[349])|(((m[129]&m[350]&~m[844]))&~BiasedRNG[349])|((m[129]&m[350]&m[844]));
    m[495] = (((m[141]&~m[351]&m[899])|(~m[141]&m[351]&m[899]))&BiasedRNG[350])|(((m[141]&m[351]&~m[899]))&~BiasedRNG[350])|((m[141]&m[351]&m[899]));
    m[496] = (((m[153]&~m[352]&m[949])|(~m[153]&m[352]&m[949]))&BiasedRNG[351])|(((m[153]&m[352]&~m[949]))&~BiasedRNG[351])|((m[153]&m[352]&m[949]));
    m[497] = (((m[165]&~m[353]&m[994])|(~m[165]&m[353]&m[994]))&BiasedRNG[352])|(((m[165]&m[353]&~m[994]))&~BiasedRNG[352])|((m[165]&m[353]&m[994]));
    m[498] = (((m[177]&~m[354]&m[1034])|(~m[177]&m[354]&m[1034]))&BiasedRNG[353])|(((m[177]&m[354]&~m[1034]))&~BiasedRNG[353])|((m[177]&m[354]&m[1034]));
    m[499] = (((m[189]&~m[355]&m[1069])|(~m[189]&m[355]&m[1069]))&BiasedRNG[354])|(((m[189]&m[355]&~m[1069]))&~BiasedRNG[354])|((m[189]&m[355]&m[1069]));
    m[500] = (((m[201]&~m[356]&m[1099])|(~m[201]&m[356]&m[1099]))&BiasedRNG[355])|(((m[201]&m[356]&~m[1099]))&~BiasedRNG[355])|((m[201]&m[356]&m[1099]));
    m[501] = (((m[213]&~m[357]&m[1124])|(~m[213]&m[357]&m[1124]))&BiasedRNG[356])|(((m[213]&m[357]&~m[1124]))&~BiasedRNG[356])|((m[213]&m[357]&m[1124]));
    m[502] = (((m[225]&~m[358]&m[1144])|(~m[225]&m[358]&m[1144]))&BiasedRNG[357])|(((m[225]&m[358]&~m[1144]))&~BiasedRNG[357])|((m[225]&m[358]&m[1144]));
    m[503] = (((m[237]&~m[359]&m[1159])|(~m[237]&m[359]&m[1159]))&BiasedRNG[358])|(((m[237]&m[359]&~m[1159]))&~BiasedRNG[358])|((m[237]&m[359]&m[1159]));
    m[504] = (((m[106]&~m[360]&m[799])|(~m[106]&m[360]&m[799]))&BiasedRNG[359])|(((m[106]&m[360]&~m[799]))&~BiasedRNG[359])|((m[106]&m[360]&m[799]));
    m[505] = (((m[118]&~m[361]&m[849])|(~m[118]&m[361]&m[849]))&BiasedRNG[360])|(((m[118]&m[361]&~m[849]))&~BiasedRNG[360])|((m[118]&m[361]&m[849]));
    m[506] = (((m[130]&~m[362]&m[904])|(~m[130]&m[362]&m[904]))&BiasedRNG[361])|(((m[130]&m[362]&~m[904]))&~BiasedRNG[361])|((m[130]&m[362]&m[904]));
    m[507] = (((m[142]&~m[363]&m[954])|(~m[142]&m[363]&m[954]))&BiasedRNG[362])|(((m[142]&m[363]&~m[954]))&~BiasedRNG[362])|((m[142]&m[363]&m[954]));
    m[508] = (((m[154]&~m[364]&m[999])|(~m[154]&m[364]&m[999]))&BiasedRNG[363])|(((m[154]&m[364]&~m[999]))&~BiasedRNG[363])|((m[154]&m[364]&m[999]));
    m[509] = (((m[166]&~m[365]&m[1039])|(~m[166]&m[365]&m[1039]))&BiasedRNG[364])|(((m[166]&m[365]&~m[1039]))&~BiasedRNG[364])|((m[166]&m[365]&m[1039]));
    m[510] = (((m[178]&~m[366]&m[1074])|(~m[178]&m[366]&m[1074]))&BiasedRNG[365])|(((m[178]&m[366]&~m[1074]))&~BiasedRNG[365])|((m[178]&m[366]&m[1074]));
    m[511] = (((m[190]&~m[367]&m[1104])|(~m[190]&m[367]&m[1104]))&BiasedRNG[366])|(((m[190]&m[367]&~m[1104]))&~BiasedRNG[366])|((m[190]&m[367]&m[1104]));
    m[512] = (((m[202]&~m[368]&m[1129])|(~m[202]&m[368]&m[1129]))&BiasedRNG[367])|(((m[202]&m[368]&~m[1129]))&~BiasedRNG[367])|((m[202]&m[368]&m[1129]));
    m[513] = (((m[214]&~m[369]&m[1149])|(~m[214]&m[369]&m[1149]))&BiasedRNG[368])|(((m[214]&m[369]&~m[1149]))&~BiasedRNG[368])|((m[214]&m[369]&m[1149]));
    m[514] = (((m[226]&~m[370]&m[1164])|(~m[226]&m[370]&m[1164]))&BiasedRNG[369])|(((m[226]&m[370]&~m[1164]))&~BiasedRNG[369])|((m[226]&m[370]&m[1164]));
    m[515] = (((m[238]&~m[371]&m[1174])|(~m[238]&m[371]&m[1174]))&BiasedRNG[370])|(((m[238]&m[371]&~m[1174]))&~BiasedRNG[370])|((m[238]&m[371]&m[1174]));
    m[516] = (((m[107]&~m[372]&m[854])|(~m[107]&m[372]&m[854]))&BiasedRNG[371])|(((m[107]&m[372]&~m[854]))&~BiasedRNG[371])|((m[107]&m[372]&m[854]));
    m[517] = (((m[119]&~m[373]&m[909])|(~m[119]&m[373]&m[909]))&BiasedRNG[372])|(((m[119]&m[373]&~m[909]))&~BiasedRNG[372])|((m[119]&m[373]&m[909]));
    m[518] = (((m[131]&~m[374]&m[959])|(~m[131]&m[374]&m[959]))&BiasedRNG[373])|(((m[131]&m[374]&~m[959]))&~BiasedRNG[373])|((m[131]&m[374]&m[959]));
    m[519] = (((m[143]&~m[375]&m[1004])|(~m[143]&m[375]&m[1004]))&BiasedRNG[374])|(((m[143]&m[375]&~m[1004]))&~BiasedRNG[374])|((m[143]&m[375]&m[1004]));
    m[520] = (((m[155]&~m[376]&m[1044])|(~m[155]&m[376]&m[1044]))&BiasedRNG[375])|(((m[155]&m[376]&~m[1044]))&~BiasedRNG[375])|((m[155]&m[376]&m[1044]));
    m[521] = (((m[167]&~m[377]&m[1079])|(~m[167]&m[377]&m[1079]))&BiasedRNG[376])|(((m[167]&m[377]&~m[1079]))&~BiasedRNG[376])|((m[167]&m[377]&m[1079]));
    m[522] = (((m[179]&~m[378]&m[1109])|(~m[179]&m[378]&m[1109]))&BiasedRNG[377])|(((m[179]&m[378]&~m[1109]))&~BiasedRNG[377])|((m[179]&m[378]&m[1109]));
    m[523] = (((m[191]&~m[379]&m[1134])|(~m[191]&m[379]&m[1134]))&BiasedRNG[378])|(((m[191]&m[379]&~m[1134]))&~BiasedRNG[378])|((m[191]&m[379]&m[1134]));
    m[524] = (((m[203]&~m[380]&m[1154])|(~m[203]&m[380]&m[1154]))&BiasedRNG[379])|(((m[203]&m[380]&~m[1154]))&~BiasedRNG[379])|((m[203]&m[380]&m[1154]));
    m[525] = (((m[215]&~m[381]&m[1169])|(~m[215]&m[381]&m[1169]))&BiasedRNG[380])|(((m[215]&m[381]&~m[1169]))&~BiasedRNG[380])|((m[215]&m[381]&m[1169]));
    m[526] = (((m[227]&~m[382]&m[1179])|(~m[227]&m[382]&m[1179]))&BiasedRNG[381])|(((m[227]&m[382]&~m[1179]))&~BiasedRNG[381])|((m[227]&m[382]&m[1179]));
    m[527] = (((m[239]&~m[383]&m[1184])|(~m[239]&m[383]&m[1184]))&BiasedRNG[382])|(((m[239]&m[383]&~m[1184]))&~BiasedRNG[382])|((m[239]&m[383]&m[1184]));
    m[535] = (((m[532]&~m[533]&~m[534]&~m[536]&~m[537])|(~m[532]&~m[533]&~m[534]&m[536]&~m[537])|(m[532]&m[533]&~m[534]&m[536]&~m[537])|(m[532]&~m[533]&m[534]&m[536]&~m[537])|(~m[532]&m[533]&~m[534]&~m[536]&m[537])|(~m[532]&~m[533]&m[534]&~m[536]&m[537])|(m[532]&m[533]&m[534]&~m[536]&m[537])|(~m[532]&m[533]&m[534]&m[536]&m[537]))&UnbiasedRNG[131])|((m[532]&~m[533]&~m[534]&m[536]&~m[537])|(~m[532]&~m[533]&~m[534]&~m[536]&m[537])|(m[532]&~m[533]&~m[534]&~m[536]&m[537])|(m[532]&m[533]&~m[534]&~m[536]&m[537])|(m[532]&~m[533]&m[534]&~m[536]&m[537])|(~m[532]&~m[533]&~m[534]&m[536]&m[537])|(m[532]&~m[533]&~m[534]&m[536]&m[537])|(~m[532]&m[533]&~m[534]&m[536]&m[537])|(m[532]&m[533]&~m[534]&m[536]&m[537])|(~m[532]&~m[533]&m[534]&m[536]&m[537])|(m[532]&~m[533]&m[534]&m[536]&m[537])|(m[532]&m[533]&m[534]&m[536]&m[537]));
    m[545] = (((m[537]&~m[543]&~m[544]&~m[546]&~m[547])|(~m[537]&~m[543]&~m[544]&m[546]&~m[547])|(m[537]&m[543]&~m[544]&m[546]&~m[547])|(m[537]&~m[543]&m[544]&m[546]&~m[547])|(~m[537]&m[543]&~m[544]&~m[546]&m[547])|(~m[537]&~m[543]&m[544]&~m[546]&m[547])|(m[537]&m[543]&m[544]&~m[546]&m[547])|(~m[537]&m[543]&m[544]&m[546]&m[547]))&UnbiasedRNG[132])|((m[537]&~m[543]&~m[544]&m[546]&~m[547])|(~m[537]&~m[543]&~m[544]&~m[546]&m[547])|(m[537]&~m[543]&~m[544]&~m[546]&m[547])|(m[537]&m[543]&~m[544]&~m[546]&m[547])|(m[537]&~m[543]&m[544]&~m[546]&m[547])|(~m[537]&~m[543]&~m[544]&m[546]&m[547])|(m[537]&~m[543]&~m[544]&m[546]&m[547])|(~m[537]&m[543]&~m[544]&m[546]&m[547])|(m[537]&m[543]&~m[544]&m[546]&m[547])|(~m[537]&~m[543]&m[544]&m[546]&m[547])|(m[537]&~m[543]&m[544]&m[546]&m[547])|(m[537]&m[543]&m[544]&m[546]&m[547]));
    m[550] = (((m[542]&~m[548]&~m[549]&~m[551]&~m[552])|(~m[542]&~m[548]&~m[549]&m[551]&~m[552])|(m[542]&m[548]&~m[549]&m[551]&~m[552])|(m[542]&~m[548]&m[549]&m[551]&~m[552])|(~m[542]&m[548]&~m[549]&~m[551]&m[552])|(~m[542]&~m[548]&m[549]&~m[551]&m[552])|(m[542]&m[548]&m[549]&~m[551]&m[552])|(~m[542]&m[548]&m[549]&m[551]&m[552]))&UnbiasedRNG[133])|((m[542]&~m[548]&~m[549]&m[551]&~m[552])|(~m[542]&~m[548]&~m[549]&~m[551]&m[552])|(m[542]&~m[548]&~m[549]&~m[551]&m[552])|(m[542]&m[548]&~m[549]&~m[551]&m[552])|(m[542]&~m[548]&m[549]&~m[551]&m[552])|(~m[542]&~m[548]&~m[549]&m[551]&m[552])|(m[542]&~m[548]&~m[549]&m[551]&m[552])|(~m[542]&m[548]&~m[549]&m[551]&m[552])|(m[542]&m[548]&~m[549]&m[551]&m[552])|(~m[542]&~m[548]&m[549]&m[551]&m[552])|(m[542]&~m[548]&m[549]&m[551]&m[552])|(m[542]&m[548]&m[549]&m[551]&m[552]));
    m[560] = (((m[547]&~m[558]&~m[559]&~m[561]&~m[562])|(~m[547]&~m[558]&~m[559]&m[561]&~m[562])|(m[547]&m[558]&~m[559]&m[561]&~m[562])|(m[547]&~m[558]&m[559]&m[561]&~m[562])|(~m[547]&m[558]&~m[559]&~m[561]&m[562])|(~m[547]&~m[558]&m[559]&~m[561]&m[562])|(m[547]&m[558]&m[559]&~m[561]&m[562])|(~m[547]&m[558]&m[559]&m[561]&m[562]))&UnbiasedRNG[134])|((m[547]&~m[558]&~m[559]&m[561]&~m[562])|(~m[547]&~m[558]&~m[559]&~m[561]&m[562])|(m[547]&~m[558]&~m[559]&~m[561]&m[562])|(m[547]&m[558]&~m[559]&~m[561]&m[562])|(m[547]&~m[558]&m[559]&~m[561]&m[562])|(~m[547]&~m[558]&~m[559]&m[561]&m[562])|(m[547]&~m[558]&~m[559]&m[561]&m[562])|(~m[547]&m[558]&~m[559]&m[561]&m[562])|(m[547]&m[558]&~m[559]&m[561]&m[562])|(~m[547]&~m[558]&m[559]&m[561]&m[562])|(m[547]&~m[558]&m[559]&m[561]&m[562])|(m[547]&m[558]&m[559]&m[561]&m[562]));
    m[565] = (((m[552]&~m[563]&~m[564]&~m[566]&~m[567])|(~m[552]&~m[563]&~m[564]&m[566]&~m[567])|(m[552]&m[563]&~m[564]&m[566]&~m[567])|(m[552]&~m[563]&m[564]&m[566]&~m[567])|(~m[552]&m[563]&~m[564]&~m[566]&m[567])|(~m[552]&~m[563]&m[564]&~m[566]&m[567])|(m[552]&m[563]&m[564]&~m[566]&m[567])|(~m[552]&m[563]&m[564]&m[566]&m[567]))&UnbiasedRNG[135])|((m[552]&~m[563]&~m[564]&m[566]&~m[567])|(~m[552]&~m[563]&~m[564]&~m[566]&m[567])|(m[552]&~m[563]&~m[564]&~m[566]&m[567])|(m[552]&m[563]&~m[564]&~m[566]&m[567])|(m[552]&~m[563]&m[564]&~m[566]&m[567])|(~m[552]&~m[563]&~m[564]&m[566]&m[567])|(m[552]&~m[563]&~m[564]&m[566]&m[567])|(~m[552]&m[563]&~m[564]&m[566]&m[567])|(m[552]&m[563]&~m[564]&m[566]&m[567])|(~m[552]&~m[563]&m[564]&m[566]&m[567])|(m[552]&~m[563]&m[564]&m[566]&m[567])|(m[552]&m[563]&m[564]&m[566]&m[567]));
    m[570] = (((m[557]&~m[568]&~m[569]&~m[571]&~m[572])|(~m[557]&~m[568]&~m[569]&m[571]&~m[572])|(m[557]&m[568]&~m[569]&m[571]&~m[572])|(m[557]&~m[568]&m[569]&m[571]&~m[572])|(~m[557]&m[568]&~m[569]&~m[571]&m[572])|(~m[557]&~m[568]&m[569]&~m[571]&m[572])|(m[557]&m[568]&m[569]&~m[571]&m[572])|(~m[557]&m[568]&m[569]&m[571]&m[572]))&UnbiasedRNG[136])|((m[557]&~m[568]&~m[569]&m[571]&~m[572])|(~m[557]&~m[568]&~m[569]&~m[571]&m[572])|(m[557]&~m[568]&~m[569]&~m[571]&m[572])|(m[557]&m[568]&~m[569]&~m[571]&m[572])|(m[557]&~m[568]&m[569]&~m[571]&m[572])|(~m[557]&~m[568]&~m[569]&m[571]&m[572])|(m[557]&~m[568]&~m[569]&m[571]&m[572])|(~m[557]&m[568]&~m[569]&m[571]&m[572])|(m[557]&m[568]&~m[569]&m[571]&m[572])|(~m[557]&~m[568]&m[569]&m[571]&m[572])|(m[557]&~m[568]&m[569]&m[571]&m[572])|(m[557]&m[568]&m[569]&m[571]&m[572]));
    m[580] = (((m[562]&~m[578]&~m[579]&~m[581]&~m[582])|(~m[562]&~m[578]&~m[579]&m[581]&~m[582])|(m[562]&m[578]&~m[579]&m[581]&~m[582])|(m[562]&~m[578]&m[579]&m[581]&~m[582])|(~m[562]&m[578]&~m[579]&~m[581]&m[582])|(~m[562]&~m[578]&m[579]&~m[581]&m[582])|(m[562]&m[578]&m[579]&~m[581]&m[582])|(~m[562]&m[578]&m[579]&m[581]&m[582]))&UnbiasedRNG[137])|((m[562]&~m[578]&~m[579]&m[581]&~m[582])|(~m[562]&~m[578]&~m[579]&~m[581]&m[582])|(m[562]&~m[578]&~m[579]&~m[581]&m[582])|(m[562]&m[578]&~m[579]&~m[581]&m[582])|(m[562]&~m[578]&m[579]&~m[581]&m[582])|(~m[562]&~m[578]&~m[579]&m[581]&m[582])|(m[562]&~m[578]&~m[579]&m[581]&m[582])|(~m[562]&m[578]&~m[579]&m[581]&m[582])|(m[562]&m[578]&~m[579]&m[581]&m[582])|(~m[562]&~m[578]&m[579]&m[581]&m[582])|(m[562]&~m[578]&m[579]&m[581]&m[582])|(m[562]&m[578]&m[579]&m[581]&m[582]));
    m[585] = (((m[567]&~m[583]&~m[584]&~m[586]&~m[587])|(~m[567]&~m[583]&~m[584]&m[586]&~m[587])|(m[567]&m[583]&~m[584]&m[586]&~m[587])|(m[567]&~m[583]&m[584]&m[586]&~m[587])|(~m[567]&m[583]&~m[584]&~m[586]&m[587])|(~m[567]&~m[583]&m[584]&~m[586]&m[587])|(m[567]&m[583]&m[584]&~m[586]&m[587])|(~m[567]&m[583]&m[584]&m[586]&m[587]))&UnbiasedRNG[138])|((m[567]&~m[583]&~m[584]&m[586]&~m[587])|(~m[567]&~m[583]&~m[584]&~m[586]&m[587])|(m[567]&~m[583]&~m[584]&~m[586]&m[587])|(m[567]&m[583]&~m[584]&~m[586]&m[587])|(m[567]&~m[583]&m[584]&~m[586]&m[587])|(~m[567]&~m[583]&~m[584]&m[586]&m[587])|(m[567]&~m[583]&~m[584]&m[586]&m[587])|(~m[567]&m[583]&~m[584]&m[586]&m[587])|(m[567]&m[583]&~m[584]&m[586]&m[587])|(~m[567]&~m[583]&m[584]&m[586]&m[587])|(m[567]&~m[583]&m[584]&m[586]&m[587])|(m[567]&m[583]&m[584]&m[586]&m[587]));
    m[590] = (((m[572]&~m[588]&~m[589]&~m[591]&~m[592])|(~m[572]&~m[588]&~m[589]&m[591]&~m[592])|(m[572]&m[588]&~m[589]&m[591]&~m[592])|(m[572]&~m[588]&m[589]&m[591]&~m[592])|(~m[572]&m[588]&~m[589]&~m[591]&m[592])|(~m[572]&~m[588]&m[589]&~m[591]&m[592])|(m[572]&m[588]&m[589]&~m[591]&m[592])|(~m[572]&m[588]&m[589]&m[591]&m[592]))&UnbiasedRNG[139])|((m[572]&~m[588]&~m[589]&m[591]&~m[592])|(~m[572]&~m[588]&~m[589]&~m[591]&m[592])|(m[572]&~m[588]&~m[589]&~m[591]&m[592])|(m[572]&m[588]&~m[589]&~m[591]&m[592])|(m[572]&~m[588]&m[589]&~m[591]&m[592])|(~m[572]&~m[588]&~m[589]&m[591]&m[592])|(m[572]&~m[588]&~m[589]&m[591]&m[592])|(~m[572]&m[588]&~m[589]&m[591]&m[592])|(m[572]&m[588]&~m[589]&m[591]&m[592])|(~m[572]&~m[588]&m[589]&m[591]&m[592])|(m[572]&~m[588]&m[589]&m[591]&m[592])|(m[572]&m[588]&m[589]&m[591]&m[592]));
    m[595] = (((m[577]&~m[593]&~m[594]&~m[596]&~m[597])|(~m[577]&~m[593]&~m[594]&m[596]&~m[597])|(m[577]&m[593]&~m[594]&m[596]&~m[597])|(m[577]&~m[593]&m[594]&m[596]&~m[597])|(~m[577]&m[593]&~m[594]&~m[596]&m[597])|(~m[577]&~m[593]&m[594]&~m[596]&m[597])|(m[577]&m[593]&m[594]&~m[596]&m[597])|(~m[577]&m[593]&m[594]&m[596]&m[597]))&UnbiasedRNG[140])|((m[577]&~m[593]&~m[594]&m[596]&~m[597])|(~m[577]&~m[593]&~m[594]&~m[596]&m[597])|(m[577]&~m[593]&~m[594]&~m[596]&m[597])|(m[577]&m[593]&~m[594]&~m[596]&m[597])|(m[577]&~m[593]&m[594]&~m[596]&m[597])|(~m[577]&~m[593]&~m[594]&m[596]&m[597])|(m[577]&~m[593]&~m[594]&m[596]&m[597])|(~m[577]&m[593]&~m[594]&m[596]&m[597])|(m[577]&m[593]&~m[594]&m[596]&m[597])|(~m[577]&~m[593]&m[594]&m[596]&m[597])|(m[577]&~m[593]&m[594]&m[596]&m[597])|(m[577]&m[593]&m[594]&m[596]&m[597]));
    m[605] = (((m[582]&~m[603]&~m[604]&~m[606]&~m[607])|(~m[582]&~m[603]&~m[604]&m[606]&~m[607])|(m[582]&m[603]&~m[604]&m[606]&~m[607])|(m[582]&~m[603]&m[604]&m[606]&~m[607])|(~m[582]&m[603]&~m[604]&~m[606]&m[607])|(~m[582]&~m[603]&m[604]&~m[606]&m[607])|(m[582]&m[603]&m[604]&~m[606]&m[607])|(~m[582]&m[603]&m[604]&m[606]&m[607]))&UnbiasedRNG[141])|((m[582]&~m[603]&~m[604]&m[606]&~m[607])|(~m[582]&~m[603]&~m[604]&~m[606]&m[607])|(m[582]&~m[603]&~m[604]&~m[606]&m[607])|(m[582]&m[603]&~m[604]&~m[606]&m[607])|(m[582]&~m[603]&m[604]&~m[606]&m[607])|(~m[582]&~m[603]&~m[604]&m[606]&m[607])|(m[582]&~m[603]&~m[604]&m[606]&m[607])|(~m[582]&m[603]&~m[604]&m[606]&m[607])|(m[582]&m[603]&~m[604]&m[606]&m[607])|(~m[582]&~m[603]&m[604]&m[606]&m[607])|(m[582]&~m[603]&m[604]&m[606]&m[607])|(m[582]&m[603]&m[604]&m[606]&m[607]));
    m[610] = (((m[587]&~m[608]&~m[609]&~m[611]&~m[612])|(~m[587]&~m[608]&~m[609]&m[611]&~m[612])|(m[587]&m[608]&~m[609]&m[611]&~m[612])|(m[587]&~m[608]&m[609]&m[611]&~m[612])|(~m[587]&m[608]&~m[609]&~m[611]&m[612])|(~m[587]&~m[608]&m[609]&~m[611]&m[612])|(m[587]&m[608]&m[609]&~m[611]&m[612])|(~m[587]&m[608]&m[609]&m[611]&m[612]))&UnbiasedRNG[142])|((m[587]&~m[608]&~m[609]&m[611]&~m[612])|(~m[587]&~m[608]&~m[609]&~m[611]&m[612])|(m[587]&~m[608]&~m[609]&~m[611]&m[612])|(m[587]&m[608]&~m[609]&~m[611]&m[612])|(m[587]&~m[608]&m[609]&~m[611]&m[612])|(~m[587]&~m[608]&~m[609]&m[611]&m[612])|(m[587]&~m[608]&~m[609]&m[611]&m[612])|(~m[587]&m[608]&~m[609]&m[611]&m[612])|(m[587]&m[608]&~m[609]&m[611]&m[612])|(~m[587]&~m[608]&m[609]&m[611]&m[612])|(m[587]&~m[608]&m[609]&m[611]&m[612])|(m[587]&m[608]&m[609]&m[611]&m[612]));
    m[615] = (((m[592]&~m[613]&~m[614]&~m[616]&~m[617])|(~m[592]&~m[613]&~m[614]&m[616]&~m[617])|(m[592]&m[613]&~m[614]&m[616]&~m[617])|(m[592]&~m[613]&m[614]&m[616]&~m[617])|(~m[592]&m[613]&~m[614]&~m[616]&m[617])|(~m[592]&~m[613]&m[614]&~m[616]&m[617])|(m[592]&m[613]&m[614]&~m[616]&m[617])|(~m[592]&m[613]&m[614]&m[616]&m[617]))&UnbiasedRNG[143])|((m[592]&~m[613]&~m[614]&m[616]&~m[617])|(~m[592]&~m[613]&~m[614]&~m[616]&m[617])|(m[592]&~m[613]&~m[614]&~m[616]&m[617])|(m[592]&m[613]&~m[614]&~m[616]&m[617])|(m[592]&~m[613]&m[614]&~m[616]&m[617])|(~m[592]&~m[613]&~m[614]&m[616]&m[617])|(m[592]&~m[613]&~m[614]&m[616]&m[617])|(~m[592]&m[613]&~m[614]&m[616]&m[617])|(m[592]&m[613]&~m[614]&m[616]&m[617])|(~m[592]&~m[613]&m[614]&m[616]&m[617])|(m[592]&~m[613]&m[614]&m[616]&m[617])|(m[592]&m[613]&m[614]&m[616]&m[617]));
    m[620] = (((m[597]&~m[618]&~m[619]&~m[621]&~m[622])|(~m[597]&~m[618]&~m[619]&m[621]&~m[622])|(m[597]&m[618]&~m[619]&m[621]&~m[622])|(m[597]&~m[618]&m[619]&m[621]&~m[622])|(~m[597]&m[618]&~m[619]&~m[621]&m[622])|(~m[597]&~m[618]&m[619]&~m[621]&m[622])|(m[597]&m[618]&m[619]&~m[621]&m[622])|(~m[597]&m[618]&m[619]&m[621]&m[622]))&UnbiasedRNG[144])|((m[597]&~m[618]&~m[619]&m[621]&~m[622])|(~m[597]&~m[618]&~m[619]&~m[621]&m[622])|(m[597]&~m[618]&~m[619]&~m[621]&m[622])|(m[597]&m[618]&~m[619]&~m[621]&m[622])|(m[597]&~m[618]&m[619]&~m[621]&m[622])|(~m[597]&~m[618]&~m[619]&m[621]&m[622])|(m[597]&~m[618]&~m[619]&m[621]&m[622])|(~m[597]&m[618]&~m[619]&m[621]&m[622])|(m[597]&m[618]&~m[619]&m[621]&m[622])|(~m[597]&~m[618]&m[619]&m[621]&m[622])|(m[597]&~m[618]&m[619]&m[621]&m[622])|(m[597]&m[618]&m[619]&m[621]&m[622]));
    m[625] = (((m[602]&~m[623]&~m[624]&~m[626]&~m[627])|(~m[602]&~m[623]&~m[624]&m[626]&~m[627])|(m[602]&m[623]&~m[624]&m[626]&~m[627])|(m[602]&~m[623]&m[624]&m[626]&~m[627])|(~m[602]&m[623]&~m[624]&~m[626]&m[627])|(~m[602]&~m[623]&m[624]&~m[626]&m[627])|(m[602]&m[623]&m[624]&~m[626]&m[627])|(~m[602]&m[623]&m[624]&m[626]&m[627]))&UnbiasedRNG[145])|((m[602]&~m[623]&~m[624]&m[626]&~m[627])|(~m[602]&~m[623]&~m[624]&~m[626]&m[627])|(m[602]&~m[623]&~m[624]&~m[626]&m[627])|(m[602]&m[623]&~m[624]&~m[626]&m[627])|(m[602]&~m[623]&m[624]&~m[626]&m[627])|(~m[602]&~m[623]&~m[624]&m[626]&m[627])|(m[602]&~m[623]&~m[624]&m[626]&m[627])|(~m[602]&m[623]&~m[624]&m[626]&m[627])|(m[602]&m[623]&~m[624]&m[626]&m[627])|(~m[602]&~m[623]&m[624]&m[626]&m[627])|(m[602]&~m[623]&m[624]&m[626]&m[627])|(m[602]&m[623]&m[624]&m[626]&m[627]));
    m[635] = (((m[607]&~m[633]&~m[634]&~m[636]&~m[637])|(~m[607]&~m[633]&~m[634]&m[636]&~m[637])|(m[607]&m[633]&~m[634]&m[636]&~m[637])|(m[607]&~m[633]&m[634]&m[636]&~m[637])|(~m[607]&m[633]&~m[634]&~m[636]&m[637])|(~m[607]&~m[633]&m[634]&~m[636]&m[637])|(m[607]&m[633]&m[634]&~m[636]&m[637])|(~m[607]&m[633]&m[634]&m[636]&m[637]))&UnbiasedRNG[146])|((m[607]&~m[633]&~m[634]&m[636]&~m[637])|(~m[607]&~m[633]&~m[634]&~m[636]&m[637])|(m[607]&~m[633]&~m[634]&~m[636]&m[637])|(m[607]&m[633]&~m[634]&~m[636]&m[637])|(m[607]&~m[633]&m[634]&~m[636]&m[637])|(~m[607]&~m[633]&~m[634]&m[636]&m[637])|(m[607]&~m[633]&~m[634]&m[636]&m[637])|(~m[607]&m[633]&~m[634]&m[636]&m[637])|(m[607]&m[633]&~m[634]&m[636]&m[637])|(~m[607]&~m[633]&m[634]&m[636]&m[637])|(m[607]&~m[633]&m[634]&m[636]&m[637])|(m[607]&m[633]&m[634]&m[636]&m[637]));
    m[640] = (((m[612]&~m[638]&~m[639]&~m[641]&~m[642])|(~m[612]&~m[638]&~m[639]&m[641]&~m[642])|(m[612]&m[638]&~m[639]&m[641]&~m[642])|(m[612]&~m[638]&m[639]&m[641]&~m[642])|(~m[612]&m[638]&~m[639]&~m[641]&m[642])|(~m[612]&~m[638]&m[639]&~m[641]&m[642])|(m[612]&m[638]&m[639]&~m[641]&m[642])|(~m[612]&m[638]&m[639]&m[641]&m[642]))&UnbiasedRNG[147])|((m[612]&~m[638]&~m[639]&m[641]&~m[642])|(~m[612]&~m[638]&~m[639]&~m[641]&m[642])|(m[612]&~m[638]&~m[639]&~m[641]&m[642])|(m[612]&m[638]&~m[639]&~m[641]&m[642])|(m[612]&~m[638]&m[639]&~m[641]&m[642])|(~m[612]&~m[638]&~m[639]&m[641]&m[642])|(m[612]&~m[638]&~m[639]&m[641]&m[642])|(~m[612]&m[638]&~m[639]&m[641]&m[642])|(m[612]&m[638]&~m[639]&m[641]&m[642])|(~m[612]&~m[638]&m[639]&m[641]&m[642])|(m[612]&~m[638]&m[639]&m[641]&m[642])|(m[612]&m[638]&m[639]&m[641]&m[642]));
    m[645] = (((m[617]&~m[643]&~m[644]&~m[646]&~m[647])|(~m[617]&~m[643]&~m[644]&m[646]&~m[647])|(m[617]&m[643]&~m[644]&m[646]&~m[647])|(m[617]&~m[643]&m[644]&m[646]&~m[647])|(~m[617]&m[643]&~m[644]&~m[646]&m[647])|(~m[617]&~m[643]&m[644]&~m[646]&m[647])|(m[617]&m[643]&m[644]&~m[646]&m[647])|(~m[617]&m[643]&m[644]&m[646]&m[647]))&UnbiasedRNG[148])|((m[617]&~m[643]&~m[644]&m[646]&~m[647])|(~m[617]&~m[643]&~m[644]&~m[646]&m[647])|(m[617]&~m[643]&~m[644]&~m[646]&m[647])|(m[617]&m[643]&~m[644]&~m[646]&m[647])|(m[617]&~m[643]&m[644]&~m[646]&m[647])|(~m[617]&~m[643]&~m[644]&m[646]&m[647])|(m[617]&~m[643]&~m[644]&m[646]&m[647])|(~m[617]&m[643]&~m[644]&m[646]&m[647])|(m[617]&m[643]&~m[644]&m[646]&m[647])|(~m[617]&~m[643]&m[644]&m[646]&m[647])|(m[617]&~m[643]&m[644]&m[646]&m[647])|(m[617]&m[643]&m[644]&m[646]&m[647]));
    m[650] = (((m[622]&~m[648]&~m[649]&~m[651]&~m[652])|(~m[622]&~m[648]&~m[649]&m[651]&~m[652])|(m[622]&m[648]&~m[649]&m[651]&~m[652])|(m[622]&~m[648]&m[649]&m[651]&~m[652])|(~m[622]&m[648]&~m[649]&~m[651]&m[652])|(~m[622]&~m[648]&m[649]&~m[651]&m[652])|(m[622]&m[648]&m[649]&~m[651]&m[652])|(~m[622]&m[648]&m[649]&m[651]&m[652]))&UnbiasedRNG[149])|((m[622]&~m[648]&~m[649]&m[651]&~m[652])|(~m[622]&~m[648]&~m[649]&~m[651]&m[652])|(m[622]&~m[648]&~m[649]&~m[651]&m[652])|(m[622]&m[648]&~m[649]&~m[651]&m[652])|(m[622]&~m[648]&m[649]&~m[651]&m[652])|(~m[622]&~m[648]&~m[649]&m[651]&m[652])|(m[622]&~m[648]&~m[649]&m[651]&m[652])|(~m[622]&m[648]&~m[649]&m[651]&m[652])|(m[622]&m[648]&~m[649]&m[651]&m[652])|(~m[622]&~m[648]&m[649]&m[651]&m[652])|(m[622]&~m[648]&m[649]&m[651]&m[652])|(m[622]&m[648]&m[649]&m[651]&m[652]));
    m[655] = (((m[627]&~m[653]&~m[654]&~m[656]&~m[657])|(~m[627]&~m[653]&~m[654]&m[656]&~m[657])|(m[627]&m[653]&~m[654]&m[656]&~m[657])|(m[627]&~m[653]&m[654]&m[656]&~m[657])|(~m[627]&m[653]&~m[654]&~m[656]&m[657])|(~m[627]&~m[653]&m[654]&~m[656]&m[657])|(m[627]&m[653]&m[654]&~m[656]&m[657])|(~m[627]&m[653]&m[654]&m[656]&m[657]))&UnbiasedRNG[150])|((m[627]&~m[653]&~m[654]&m[656]&~m[657])|(~m[627]&~m[653]&~m[654]&~m[656]&m[657])|(m[627]&~m[653]&~m[654]&~m[656]&m[657])|(m[627]&m[653]&~m[654]&~m[656]&m[657])|(m[627]&~m[653]&m[654]&~m[656]&m[657])|(~m[627]&~m[653]&~m[654]&m[656]&m[657])|(m[627]&~m[653]&~m[654]&m[656]&m[657])|(~m[627]&m[653]&~m[654]&m[656]&m[657])|(m[627]&m[653]&~m[654]&m[656]&m[657])|(~m[627]&~m[653]&m[654]&m[656]&m[657])|(m[627]&~m[653]&m[654]&m[656]&m[657])|(m[627]&m[653]&m[654]&m[656]&m[657]));
    m[660] = (((m[632]&~m[658]&~m[659]&~m[661]&~m[662])|(~m[632]&~m[658]&~m[659]&m[661]&~m[662])|(m[632]&m[658]&~m[659]&m[661]&~m[662])|(m[632]&~m[658]&m[659]&m[661]&~m[662])|(~m[632]&m[658]&~m[659]&~m[661]&m[662])|(~m[632]&~m[658]&m[659]&~m[661]&m[662])|(m[632]&m[658]&m[659]&~m[661]&m[662])|(~m[632]&m[658]&m[659]&m[661]&m[662]))&UnbiasedRNG[151])|((m[632]&~m[658]&~m[659]&m[661]&~m[662])|(~m[632]&~m[658]&~m[659]&~m[661]&m[662])|(m[632]&~m[658]&~m[659]&~m[661]&m[662])|(m[632]&m[658]&~m[659]&~m[661]&m[662])|(m[632]&~m[658]&m[659]&~m[661]&m[662])|(~m[632]&~m[658]&~m[659]&m[661]&m[662])|(m[632]&~m[658]&~m[659]&m[661]&m[662])|(~m[632]&m[658]&~m[659]&m[661]&m[662])|(m[632]&m[658]&~m[659]&m[661]&m[662])|(~m[632]&~m[658]&m[659]&m[661]&m[662])|(m[632]&~m[658]&m[659]&m[661]&m[662])|(m[632]&m[658]&m[659]&m[661]&m[662]));
    m[670] = (((m[637]&~m[668]&~m[669]&~m[671]&~m[672])|(~m[637]&~m[668]&~m[669]&m[671]&~m[672])|(m[637]&m[668]&~m[669]&m[671]&~m[672])|(m[637]&~m[668]&m[669]&m[671]&~m[672])|(~m[637]&m[668]&~m[669]&~m[671]&m[672])|(~m[637]&~m[668]&m[669]&~m[671]&m[672])|(m[637]&m[668]&m[669]&~m[671]&m[672])|(~m[637]&m[668]&m[669]&m[671]&m[672]))&UnbiasedRNG[152])|((m[637]&~m[668]&~m[669]&m[671]&~m[672])|(~m[637]&~m[668]&~m[669]&~m[671]&m[672])|(m[637]&~m[668]&~m[669]&~m[671]&m[672])|(m[637]&m[668]&~m[669]&~m[671]&m[672])|(m[637]&~m[668]&m[669]&~m[671]&m[672])|(~m[637]&~m[668]&~m[669]&m[671]&m[672])|(m[637]&~m[668]&~m[669]&m[671]&m[672])|(~m[637]&m[668]&~m[669]&m[671]&m[672])|(m[637]&m[668]&~m[669]&m[671]&m[672])|(~m[637]&~m[668]&m[669]&m[671]&m[672])|(m[637]&~m[668]&m[669]&m[671]&m[672])|(m[637]&m[668]&m[669]&m[671]&m[672]));
    m[675] = (((m[642]&~m[673]&~m[674]&~m[676]&~m[677])|(~m[642]&~m[673]&~m[674]&m[676]&~m[677])|(m[642]&m[673]&~m[674]&m[676]&~m[677])|(m[642]&~m[673]&m[674]&m[676]&~m[677])|(~m[642]&m[673]&~m[674]&~m[676]&m[677])|(~m[642]&~m[673]&m[674]&~m[676]&m[677])|(m[642]&m[673]&m[674]&~m[676]&m[677])|(~m[642]&m[673]&m[674]&m[676]&m[677]))&UnbiasedRNG[153])|((m[642]&~m[673]&~m[674]&m[676]&~m[677])|(~m[642]&~m[673]&~m[674]&~m[676]&m[677])|(m[642]&~m[673]&~m[674]&~m[676]&m[677])|(m[642]&m[673]&~m[674]&~m[676]&m[677])|(m[642]&~m[673]&m[674]&~m[676]&m[677])|(~m[642]&~m[673]&~m[674]&m[676]&m[677])|(m[642]&~m[673]&~m[674]&m[676]&m[677])|(~m[642]&m[673]&~m[674]&m[676]&m[677])|(m[642]&m[673]&~m[674]&m[676]&m[677])|(~m[642]&~m[673]&m[674]&m[676]&m[677])|(m[642]&~m[673]&m[674]&m[676]&m[677])|(m[642]&m[673]&m[674]&m[676]&m[677]));
    m[680] = (((m[647]&~m[678]&~m[679]&~m[681]&~m[682])|(~m[647]&~m[678]&~m[679]&m[681]&~m[682])|(m[647]&m[678]&~m[679]&m[681]&~m[682])|(m[647]&~m[678]&m[679]&m[681]&~m[682])|(~m[647]&m[678]&~m[679]&~m[681]&m[682])|(~m[647]&~m[678]&m[679]&~m[681]&m[682])|(m[647]&m[678]&m[679]&~m[681]&m[682])|(~m[647]&m[678]&m[679]&m[681]&m[682]))&UnbiasedRNG[154])|((m[647]&~m[678]&~m[679]&m[681]&~m[682])|(~m[647]&~m[678]&~m[679]&~m[681]&m[682])|(m[647]&~m[678]&~m[679]&~m[681]&m[682])|(m[647]&m[678]&~m[679]&~m[681]&m[682])|(m[647]&~m[678]&m[679]&~m[681]&m[682])|(~m[647]&~m[678]&~m[679]&m[681]&m[682])|(m[647]&~m[678]&~m[679]&m[681]&m[682])|(~m[647]&m[678]&~m[679]&m[681]&m[682])|(m[647]&m[678]&~m[679]&m[681]&m[682])|(~m[647]&~m[678]&m[679]&m[681]&m[682])|(m[647]&~m[678]&m[679]&m[681]&m[682])|(m[647]&m[678]&m[679]&m[681]&m[682]));
    m[685] = (((m[652]&~m[683]&~m[684]&~m[686]&~m[687])|(~m[652]&~m[683]&~m[684]&m[686]&~m[687])|(m[652]&m[683]&~m[684]&m[686]&~m[687])|(m[652]&~m[683]&m[684]&m[686]&~m[687])|(~m[652]&m[683]&~m[684]&~m[686]&m[687])|(~m[652]&~m[683]&m[684]&~m[686]&m[687])|(m[652]&m[683]&m[684]&~m[686]&m[687])|(~m[652]&m[683]&m[684]&m[686]&m[687]))&UnbiasedRNG[155])|((m[652]&~m[683]&~m[684]&m[686]&~m[687])|(~m[652]&~m[683]&~m[684]&~m[686]&m[687])|(m[652]&~m[683]&~m[684]&~m[686]&m[687])|(m[652]&m[683]&~m[684]&~m[686]&m[687])|(m[652]&~m[683]&m[684]&~m[686]&m[687])|(~m[652]&~m[683]&~m[684]&m[686]&m[687])|(m[652]&~m[683]&~m[684]&m[686]&m[687])|(~m[652]&m[683]&~m[684]&m[686]&m[687])|(m[652]&m[683]&~m[684]&m[686]&m[687])|(~m[652]&~m[683]&m[684]&m[686]&m[687])|(m[652]&~m[683]&m[684]&m[686]&m[687])|(m[652]&m[683]&m[684]&m[686]&m[687]));
    m[690] = (((m[657]&~m[688]&~m[689]&~m[691]&~m[692])|(~m[657]&~m[688]&~m[689]&m[691]&~m[692])|(m[657]&m[688]&~m[689]&m[691]&~m[692])|(m[657]&~m[688]&m[689]&m[691]&~m[692])|(~m[657]&m[688]&~m[689]&~m[691]&m[692])|(~m[657]&~m[688]&m[689]&~m[691]&m[692])|(m[657]&m[688]&m[689]&~m[691]&m[692])|(~m[657]&m[688]&m[689]&m[691]&m[692]))&UnbiasedRNG[156])|((m[657]&~m[688]&~m[689]&m[691]&~m[692])|(~m[657]&~m[688]&~m[689]&~m[691]&m[692])|(m[657]&~m[688]&~m[689]&~m[691]&m[692])|(m[657]&m[688]&~m[689]&~m[691]&m[692])|(m[657]&~m[688]&m[689]&~m[691]&m[692])|(~m[657]&~m[688]&~m[689]&m[691]&m[692])|(m[657]&~m[688]&~m[689]&m[691]&m[692])|(~m[657]&m[688]&~m[689]&m[691]&m[692])|(m[657]&m[688]&~m[689]&m[691]&m[692])|(~m[657]&~m[688]&m[689]&m[691]&m[692])|(m[657]&~m[688]&m[689]&m[691]&m[692])|(m[657]&m[688]&m[689]&m[691]&m[692]));
    m[695] = (((m[662]&~m[693]&~m[694]&~m[696]&~m[697])|(~m[662]&~m[693]&~m[694]&m[696]&~m[697])|(m[662]&m[693]&~m[694]&m[696]&~m[697])|(m[662]&~m[693]&m[694]&m[696]&~m[697])|(~m[662]&m[693]&~m[694]&~m[696]&m[697])|(~m[662]&~m[693]&m[694]&~m[696]&m[697])|(m[662]&m[693]&m[694]&~m[696]&m[697])|(~m[662]&m[693]&m[694]&m[696]&m[697]))&UnbiasedRNG[157])|((m[662]&~m[693]&~m[694]&m[696]&~m[697])|(~m[662]&~m[693]&~m[694]&~m[696]&m[697])|(m[662]&~m[693]&~m[694]&~m[696]&m[697])|(m[662]&m[693]&~m[694]&~m[696]&m[697])|(m[662]&~m[693]&m[694]&~m[696]&m[697])|(~m[662]&~m[693]&~m[694]&m[696]&m[697])|(m[662]&~m[693]&~m[694]&m[696]&m[697])|(~m[662]&m[693]&~m[694]&m[696]&m[697])|(m[662]&m[693]&~m[694]&m[696]&m[697])|(~m[662]&~m[693]&m[694]&m[696]&m[697])|(m[662]&~m[693]&m[694]&m[696]&m[697])|(m[662]&m[693]&m[694]&m[696]&m[697]));
    m[700] = (((m[667]&~m[698]&~m[699]&~m[701]&~m[702])|(~m[667]&~m[698]&~m[699]&m[701]&~m[702])|(m[667]&m[698]&~m[699]&m[701]&~m[702])|(m[667]&~m[698]&m[699]&m[701]&~m[702])|(~m[667]&m[698]&~m[699]&~m[701]&m[702])|(~m[667]&~m[698]&m[699]&~m[701]&m[702])|(m[667]&m[698]&m[699]&~m[701]&m[702])|(~m[667]&m[698]&m[699]&m[701]&m[702]))&UnbiasedRNG[158])|((m[667]&~m[698]&~m[699]&m[701]&~m[702])|(~m[667]&~m[698]&~m[699]&~m[701]&m[702])|(m[667]&~m[698]&~m[699]&~m[701]&m[702])|(m[667]&m[698]&~m[699]&~m[701]&m[702])|(m[667]&~m[698]&m[699]&~m[701]&m[702])|(~m[667]&~m[698]&~m[699]&m[701]&m[702])|(m[667]&~m[698]&~m[699]&m[701]&m[702])|(~m[667]&m[698]&~m[699]&m[701]&m[702])|(m[667]&m[698]&~m[699]&m[701]&m[702])|(~m[667]&~m[698]&m[699]&m[701]&m[702])|(m[667]&~m[698]&m[699]&m[701]&m[702])|(m[667]&m[698]&m[699]&m[701]&m[702]));
    m[710] = (((m[672]&~m[708]&~m[709]&~m[711]&~m[712])|(~m[672]&~m[708]&~m[709]&m[711]&~m[712])|(m[672]&m[708]&~m[709]&m[711]&~m[712])|(m[672]&~m[708]&m[709]&m[711]&~m[712])|(~m[672]&m[708]&~m[709]&~m[711]&m[712])|(~m[672]&~m[708]&m[709]&~m[711]&m[712])|(m[672]&m[708]&m[709]&~m[711]&m[712])|(~m[672]&m[708]&m[709]&m[711]&m[712]))&UnbiasedRNG[159])|((m[672]&~m[708]&~m[709]&m[711]&~m[712])|(~m[672]&~m[708]&~m[709]&~m[711]&m[712])|(m[672]&~m[708]&~m[709]&~m[711]&m[712])|(m[672]&m[708]&~m[709]&~m[711]&m[712])|(m[672]&~m[708]&m[709]&~m[711]&m[712])|(~m[672]&~m[708]&~m[709]&m[711]&m[712])|(m[672]&~m[708]&~m[709]&m[711]&m[712])|(~m[672]&m[708]&~m[709]&m[711]&m[712])|(m[672]&m[708]&~m[709]&m[711]&m[712])|(~m[672]&~m[708]&m[709]&m[711]&m[712])|(m[672]&~m[708]&m[709]&m[711]&m[712])|(m[672]&m[708]&m[709]&m[711]&m[712]));
    m[715] = (((m[677]&~m[713]&~m[714]&~m[716]&~m[717])|(~m[677]&~m[713]&~m[714]&m[716]&~m[717])|(m[677]&m[713]&~m[714]&m[716]&~m[717])|(m[677]&~m[713]&m[714]&m[716]&~m[717])|(~m[677]&m[713]&~m[714]&~m[716]&m[717])|(~m[677]&~m[713]&m[714]&~m[716]&m[717])|(m[677]&m[713]&m[714]&~m[716]&m[717])|(~m[677]&m[713]&m[714]&m[716]&m[717]))&UnbiasedRNG[160])|((m[677]&~m[713]&~m[714]&m[716]&~m[717])|(~m[677]&~m[713]&~m[714]&~m[716]&m[717])|(m[677]&~m[713]&~m[714]&~m[716]&m[717])|(m[677]&m[713]&~m[714]&~m[716]&m[717])|(m[677]&~m[713]&m[714]&~m[716]&m[717])|(~m[677]&~m[713]&~m[714]&m[716]&m[717])|(m[677]&~m[713]&~m[714]&m[716]&m[717])|(~m[677]&m[713]&~m[714]&m[716]&m[717])|(m[677]&m[713]&~m[714]&m[716]&m[717])|(~m[677]&~m[713]&m[714]&m[716]&m[717])|(m[677]&~m[713]&m[714]&m[716]&m[717])|(m[677]&m[713]&m[714]&m[716]&m[717]));
    m[720] = (((m[682]&~m[718]&~m[719]&~m[721]&~m[722])|(~m[682]&~m[718]&~m[719]&m[721]&~m[722])|(m[682]&m[718]&~m[719]&m[721]&~m[722])|(m[682]&~m[718]&m[719]&m[721]&~m[722])|(~m[682]&m[718]&~m[719]&~m[721]&m[722])|(~m[682]&~m[718]&m[719]&~m[721]&m[722])|(m[682]&m[718]&m[719]&~m[721]&m[722])|(~m[682]&m[718]&m[719]&m[721]&m[722]))&UnbiasedRNG[161])|((m[682]&~m[718]&~m[719]&m[721]&~m[722])|(~m[682]&~m[718]&~m[719]&~m[721]&m[722])|(m[682]&~m[718]&~m[719]&~m[721]&m[722])|(m[682]&m[718]&~m[719]&~m[721]&m[722])|(m[682]&~m[718]&m[719]&~m[721]&m[722])|(~m[682]&~m[718]&~m[719]&m[721]&m[722])|(m[682]&~m[718]&~m[719]&m[721]&m[722])|(~m[682]&m[718]&~m[719]&m[721]&m[722])|(m[682]&m[718]&~m[719]&m[721]&m[722])|(~m[682]&~m[718]&m[719]&m[721]&m[722])|(m[682]&~m[718]&m[719]&m[721]&m[722])|(m[682]&m[718]&m[719]&m[721]&m[722]));
    m[725] = (((m[687]&~m[723]&~m[724]&~m[726]&~m[727])|(~m[687]&~m[723]&~m[724]&m[726]&~m[727])|(m[687]&m[723]&~m[724]&m[726]&~m[727])|(m[687]&~m[723]&m[724]&m[726]&~m[727])|(~m[687]&m[723]&~m[724]&~m[726]&m[727])|(~m[687]&~m[723]&m[724]&~m[726]&m[727])|(m[687]&m[723]&m[724]&~m[726]&m[727])|(~m[687]&m[723]&m[724]&m[726]&m[727]))&UnbiasedRNG[162])|((m[687]&~m[723]&~m[724]&m[726]&~m[727])|(~m[687]&~m[723]&~m[724]&~m[726]&m[727])|(m[687]&~m[723]&~m[724]&~m[726]&m[727])|(m[687]&m[723]&~m[724]&~m[726]&m[727])|(m[687]&~m[723]&m[724]&~m[726]&m[727])|(~m[687]&~m[723]&~m[724]&m[726]&m[727])|(m[687]&~m[723]&~m[724]&m[726]&m[727])|(~m[687]&m[723]&~m[724]&m[726]&m[727])|(m[687]&m[723]&~m[724]&m[726]&m[727])|(~m[687]&~m[723]&m[724]&m[726]&m[727])|(m[687]&~m[723]&m[724]&m[726]&m[727])|(m[687]&m[723]&m[724]&m[726]&m[727]));
    m[730] = (((m[692]&~m[728]&~m[729]&~m[731]&~m[732])|(~m[692]&~m[728]&~m[729]&m[731]&~m[732])|(m[692]&m[728]&~m[729]&m[731]&~m[732])|(m[692]&~m[728]&m[729]&m[731]&~m[732])|(~m[692]&m[728]&~m[729]&~m[731]&m[732])|(~m[692]&~m[728]&m[729]&~m[731]&m[732])|(m[692]&m[728]&m[729]&~m[731]&m[732])|(~m[692]&m[728]&m[729]&m[731]&m[732]))&UnbiasedRNG[163])|((m[692]&~m[728]&~m[729]&m[731]&~m[732])|(~m[692]&~m[728]&~m[729]&~m[731]&m[732])|(m[692]&~m[728]&~m[729]&~m[731]&m[732])|(m[692]&m[728]&~m[729]&~m[731]&m[732])|(m[692]&~m[728]&m[729]&~m[731]&m[732])|(~m[692]&~m[728]&~m[729]&m[731]&m[732])|(m[692]&~m[728]&~m[729]&m[731]&m[732])|(~m[692]&m[728]&~m[729]&m[731]&m[732])|(m[692]&m[728]&~m[729]&m[731]&m[732])|(~m[692]&~m[728]&m[729]&m[731]&m[732])|(m[692]&~m[728]&m[729]&m[731]&m[732])|(m[692]&m[728]&m[729]&m[731]&m[732]));
    m[735] = (((m[697]&~m[733]&~m[734]&~m[736]&~m[737])|(~m[697]&~m[733]&~m[734]&m[736]&~m[737])|(m[697]&m[733]&~m[734]&m[736]&~m[737])|(m[697]&~m[733]&m[734]&m[736]&~m[737])|(~m[697]&m[733]&~m[734]&~m[736]&m[737])|(~m[697]&~m[733]&m[734]&~m[736]&m[737])|(m[697]&m[733]&m[734]&~m[736]&m[737])|(~m[697]&m[733]&m[734]&m[736]&m[737]))&UnbiasedRNG[164])|((m[697]&~m[733]&~m[734]&m[736]&~m[737])|(~m[697]&~m[733]&~m[734]&~m[736]&m[737])|(m[697]&~m[733]&~m[734]&~m[736]&m[737])|(m[697]&m[733]&~m[734]&~m[736]&m[737])|(m[697]&~m[733]&m[734]&~m[736]&m[737])|(~m[697]&~m[733]&~m[734]&m[736]&m[737])|(m[697]&~m[733]&~m[734]&m[736]&m[737])|(~m[697]&m[733]&~m[734]&m[736]&m[737])|(m[697]&m[733]&~m[734]&m[736]&m[737])|(~m[697]&~m[733]&m[734]&m[736]&m[737])|(m[697]&~m[733]&m[734]&m[736]&m[737])|(m[697]&m[733]&m[734]&m[736]&m[737]));
    m[740] = (((m[702]&~m[738]&~m[739]&~m[741]&~m[742])|(~m[702]&~m[738]&~m[739]&m[741]&~m[742])|(m[702]&m[738]&~m[739]&m[741]&~m[742])|(m[702]&~m[738]&m[739]&m[741]&~m[742])|(~m[702]&m[738]&~m[739]&~m[741]&m[742])|(~m[702]&~m[738]&m[739]&~m[741]&m[742])|(m[702]&m[738]&m[739]&~m[741]&m[742])|(~m[702]&m[738]&m[739]&m[741]&m[742]))&UnbiasedRNG[165])|((m[702]&~m[738]&~m[739]&m[741]&~m[742])|(~m[702]&~m[738]&~m[739]&~m[741]&m[742])|(m[702]&~m[738]&~m[739]&~m[741]&m[742])|(m[702]&m[738]&~m[739]&~m[741]&m[742])|(m[702]&~m[738]&m[739]&~m[741]&m[742])|(~m[702]&~m[738]&~m[739]&m[741]&m[742])|(m[702]&~m[738]&~m[739]&m[741]&m[742])|(~m[702]&m[738]&~m[739]&m[741]&m[742])|(m[702]&m[738]&~m[739]&m[741]&m[742])|(~m[702]&~m[738]&m[739]&m[741]&m[742])|(m[702]&~m[738]&m[739]&m[741]&m[742])|(m[702]&m[738]&m[739]&m[741]&m[742]));
    m[745] = (((m[707]&~m[743]&~m[744]&~m[746]&~m[747])|(~m[707]&~m[743]&~m[744]&m[746]&~m[747])|(m[707]&m[743]&~m[744]&m[746]&~m[747])|(m[707]&~m[743]&m[744]&m[746]&~m[747])|(~m[707]&m[743]&~m[744]&~m[746]&m[747])|(~m[707]&~m[743]&m[744]&~m[746]&m[747])|(m[707]&m[743]&m[744]&~m[746]&m[747])|(~m[707]&m[743]&m[744]&m[746]&m[747]))&UnbiasedRNG[166])|((m[707]&~m[743]&~m[744]&m[746]&~m[747])|(~m[707]&~m[743]&~m[744]&~m[746]&m[747])|(m[707]&~m[743]&~m[744]&~m[746]&m[747])|(m[707]&m[743]&~m[744]&~m[746]&m[747])|(m[707]&~m[743]&m[744]&~m[746]&m[747])|(~m[707]&~m[743]&~m[744]&m[746]&m[747])|(m[707]&~m[743]&~m[744]&m[746]&m[747])|(~m[707]&m[743]&~m[744]&m[746]&m[747])|(m[707]&m[743]&~m[744]&m[746]&m[747])|(~m[707]&~m[743]&m[744]&m[746]&m[747])|(m[707]&~m[743]&m[744]&m[746]&m[747])|(m[707]&m[743]&m[744]&m[746]&m[747]));
    m[755] = (((m[712]&~m[753]&~m[754]&~m[756]&~m[757])|(~m[712]&~m[753]&~m[754]&m[756]&~m[757])|(m[712]&m[753]&~m[754]&m[756]&~m[757])|(m[712]&~m[753]&m[754]&m[756]&~m[757])|(~m[712]&m[753]&~m[754]&~m[756]&m[757])|(~m[712]&~m[753]&m[754]&~m[756]&m[757])|(m[712]&m[753]&m[754]&~m[756]&m[757])|(~m[712]&m[753]&m[754]&m[756]&m[757]))&UnbiasedRNG[167])|((m[712]&~m[753]&~m[754]&m[756]&~m[757])|(~m[712]&~m[753]&~m[754]&~m[756]&m[757])|(m[712]&~m[753]&~m[754]&~m[756]&m[757])|(m[712]&m[753]&~m[754]&~m[756]&m[757])|(m[712]&~m[753]&m[754]&~m[756]&m[757])|(~m[712]&~m[753]&~m[754]&m[756]&m[757])|(m[712]&~m[753]&~m[754]&m[756]&m[757])|(~m[712]&m[753]&~m[754]&m[756]&m[757])|(m[712]&m[753]&~m[754]&m[756]&m[757])|(~m[712]&~m[753]&m[754]&m[756]&m[757])|(m[712]&~m[753]&m[754]&m[756]&m[757])|(m[712]&m[753]&m[754]&m[756]&m[757]));
    m[760] = (((m[717]&~m[758]&~m[759]&~m[761]&~m[762])|(~m[717]&~m[758]&~m[759]&m[761]&~m[762])|(m[717]&m[758]&~m[759]&m[761]&~m[762])|(m[717]&~m[758]&m[759]&m[761]&~m[762])|(~m[717]&m[758]&~m[759]&~m[761]&m[762])|(~m[717]&~m[758]&m[759]&~m[761]&m[762])|(m[717]&m[758]&m[759]&~m[761]&m[762])|(~m[717]&m[758]&m[759]&m[761]&m[762]))&UnbiasedRNG[168])|((m[717]&~m[758]&~m[759]&m[761]&~m[762])|(~m[717]&~m[758]&~m[759]&~m[761]&m[762])|(m[717]&~m[758]&~m[759]&~m[761]&m[762])|(m[717]&m[758]&~m[759]&~m[761]&m[762])|(m[717]&~m[758]&m[759]&~m[761]&m[762])|(~m[717]&~m[758]&~m[759]&m[761]&m[762])|(m[717]&~m[758]&~m[759]&m[761]&m[762])|(~m[717]&m[758]&~m[759]&m[761]&m[762])|(m[717]&m[758]&~m[759]&m[761]&m[762])|(~m[717]&~m[758]&m[759]&m[761]&m[762])|(m[717]&~m[758]&m[759]&m[761]&m[762])|(m[717]&m[758]&m[759]&m[761]&m[762]));
    m[765] = (((m[722]&~m[763]&~m[764]&~m[766]&~m[767])|(~m[722]&~m[763]&~m[764]&m[766]&~m[767])|(m[722]&m[763]&~m[764]&m[766]&~m[767])|(m[722]&~m[763]&m[764]&m[766]&~m[767])|(~m[722]&m[763]&~m[764]&~m[766]&m[767])|(~m[722]&~m[763]&m[764]&~m[766]&m[767])|(m[722]&m[763]&m[764]&~m[766]&m[767])|(~m[722]&m[763]&m[764]&m[766]&m[767]))&UnbiasedRNG[169])|((m[722]&~m[763]&~m[764]&m[766]&~m[767])|(~m[722]&~m[763]&~m[764]&~m[766]&m[767])|(m[722]&~m[763]&~m[764]&~m[766]&m[767])|(m[722]&m[763]&~m[764]&~m[766]&m[767])|(m[722]&~m[763]&m[764]&~m[766]&m[767])|(~m[722]&~m[763]&~m[764]&m[766]&m[767])|(m[722]&~m[763]&~m[764]&m[766]&m[767])|(~m[722]&m[763]&~m[764]&m[766]&m[767])|(m[722]&m[763]&~m[764]&m[766]&m[767])|(~m[722]&~m[763]&m[764]&m[766]&m[767])|(m[722]&~m[763]&m[764]&m[766]&m[767])|(m[722]&m[763]&m[764]&m[766]&m[767]));
    m[770] = (((m[727]&~m[768]&~m[769]&~m[771]&~m[772])|(~m[727]&~m[768]&~m[769]&m[771]&~m[772])|(m[727]&m[768]&~m[769]&m[771]&~m[772])|(m[727]&~m[768]&m[769]&m[771]&~m[772])|(~m[727]&m[768]&~m[769]&~m[771]&m[772])|(~m[727]&~m[768]&m[769]&~m[771]&m[772])|(m[727]&m[768]&m[769]&~m[771]&m[772])|(~m[727]&m[768]&m[769]&m[771]&m[772]))&UnbiasedRNG[170])|((m[727]&~m[768]&~m[769]&m[771]&~m[772])|(~m[727]&~m[768]&~m[769]&~m[771]&m[772])|(m[727]&~m[768]&~m[769]&~m[771]&m[772])|(m[727]&m[768]&~m[769]&~m[771]&m[772])|(m[727]&~m[768]&m[769]&~m[771]&m[772])|(~m[727]&~m[768]&~m[769]&m[771]&m[772])|(m[727]&~m[768]&~m[769]&m[771]&m[772])|(~m[727]&m[768]&~m[769]&m[771]&m[772])|(m[727]&m[768]&~m[769]&m[771]&m[772])|(~m[727]&~m[768]&m[769]&m[771]&m[772])|(m[727]&~m[768]&m[769]&m[771]&m[772])|(m[727]&m[768]&m[769]&m[771]&m[772]));
    m[775] = (((m[732]&~m[773]&~m[774]&~m[776]&~m[777])|(~m[732]&~m[773]&~m[774]&m[776]&~m[777])|(m[732]&m[773]&~m[774]&m[776]&~m[777])|(m[732]&~m[773]&m[774]&m[776]&~m[777])|(~m[732]&m[773]&~m[774]&~m[776]&m[777])|(~m[732]&~m[773]&m[774]&~m[776]&m[777])|(m[732]&m[773]&m[774]&~m[776]&m[777])|(~m[732]&m[773]&m[774]&m[776]&m[777]))&UnbiasedRNG[171])|((m[732]&~m[773]&~m[774]&m[776]&~m[777])|(~m[732]&~m[773]&~m[774]&~m[776]&m[777])|(m[732]&~m[773]&~m[774]&~m[776]&m[777])|(m[732]&m[773]&~m[774]&~m[776]&m[777])|(m[732]&~m[773]&m[774]&~m[776]&m[777])|(~m[732]&~m[773]&~m[774]&m[776]&m[777])|(m[732]&~m[773]&~m[774]&m[776]&m[777])|(~m[732]&m[773]&~m[774]&m[776]&m[777])|(m[732]&m[773]&~m[774]&m[776]&m[777])|(~m[732]&~m[773]&m[774]&m[776]&m[777])|(m[732]&~m[773]&m[774]&m[776]&m[777])|(m[732]&m[773]&m[774]&m[776]&m[777]));
    m[780] = (((m[737]&~m[778]&~m[779]&~m[781]&~m[782])|(~m[737]&~m[778]&~m[779]&m[781]&~m[782])|(m[737]&m[778]&~m[779]&m[781]&~m[782])|(m[737]&~m[778]&m[779]&m[781]&~m[782])|(~m[737]&m[778]&~m[779]&~m[781]&m[782])|(~m[737]&~m[778]&m[779]&~m[781]&m[782])|(m[737]&m[778]&m[779]&~m[781]&m[782])|(~m[737]&m[778]&m[779]&m[781]&m[782]))&UnbiasedRNG[172])|((m[737]&~m[778]&~m[779]&m[781]&~m[782])|(~m[737]&~m[778]&~m[779]&~m[781]&m[782])|(m[737]&~m[778]&~m[779]&~m[781]&m[782])|(m[737]&m[778]&~m[779]&~m[781]&m[782])|(m[737]&~m[778]&m[779]&~m[781]&m[782])|(~m[737]&~m[778]&~m[779]&m[781]&m[782])|(m[737]&~m[778]&~m[779]&m[781]&m[782])|(~m[737]&m[778]&~m[779]&m[781]&m[782])|(m[737]&m[778]&~m[779]&m[781]&m[782])|(~m[737]&~m[778]&m[779]&m[781]&m[782])|(m[737]&~m[778]&m[779]&m[781]&m[782])|(m[737]&m[778]&m[779]&m[781]&m[782]));
    m[785] = (((m[742]&~m[783]&~m[784]&~m[786]&~m[787])|(~m[742]&~m[783]&~m[784]&m[786]&~m[787])|(m[742]&m[783]&~m[784]&m[786]&~m[787])|(m[742]&~m[783]&m[784]&m[786]&~m[787])|(~m[742]&m[783]&~m[784]&~m[786]&m[787])|(~m[742]&~m[783]&m[784]&~m[786]&m[787])|(m[742]&m[783]&m[784]&~m[786]&m[787])|(~m[742]&m[783]&m[784]&m[786]&m[787]))&UnbiasedRNG[173])|((m[742]&~m[783]&~m[784]&m[786]&~m[787])|(~m[742]&~m[783]&~m[784]&~m[786]&m[787])|(m[742]&~m[783]&~m[784]&~m[786]&m[787])|(m[742]&m[783]&~m[784]&~m[786]&m[787])|(m[742]&~m[783]&m[784]&~m[786]&m[787])|(~m[742]&~m[783]&~m[784]&m[786]&m[787])|(m[742]&~m[783]&~m[784]&m[786]&m[787])|(~m[742]&m[783]&~m[784]&m[786]&m[787])|(m[742]&m[783]&~m[784]&m[786]&m[787])|(~m[742]&~m[783]&m[784]&m[786]&m[787])|(m[742]&~m[783]&m[784]&m[786]&m[787])|(m[742]&m[783]&m[784]&m[786]&m[787]));
    m[790] = (((m[747]&~m[788]&~m[789]&~m[791]&~m[792])|(~m[747]&~m[788]&~m[789]&m[791]&~m[792])|(m[747]&m[788]&~m[789]&m[791]&~m[792])|(m[747]&~m[788]&m[789]&m[791]&~m[792])|(~m[747]&m[788]&~m[789]&~m[791]&m[792])|(~m[747]&~m[788]&m[789]&~m[791]&m[792])|(m[747]&m[788]&m[789]&~m[791]&m[792])|(~m[747]&m[788]&m[789]&m[791]&m[792]))&UnbiasedRNG[174])|((m[747]&~m[788]&~m[789]&m[791]&~m[792])|(~m[747]&~m[788]&~m[789]&~m[791]&m[792])|(m[747]&~m[788]&~m[789]&~m[791]&m[792])|(m[747]&m[788]&~m[789]&~m[791]&m[792])|(m[747]&~m[788]&m[789]&~m[791]&m[792])|(~m[747]&~m[788]&~m[789]&m[791]&m[792])|(m[747]&~m[788]&~m[789]&m[791]&m[792])|(~m[747]&m[788]&~m[789]&m[791]&m[792])|(m[747]&m[788]&~m[789]&m[791]&m[792])|(~m[747]&~m[788]&m[789]&m[791]&m[792])|(m[747]&~m[788]&m[789]&m[791]&m[792])|(m[747]&m[788]&m[789]&m[791]&m[792]));
    m[795] = (((m[752]&~m[793]&~m[794]&~m[796]&~m[797])|(~m[752]&~m[793]&~m[794]&m[796]&~m[797])|(m[752]&m[793]&~m[794]&m[796]&~m[797])|(m[752]&~m[793]&m[794]&m[796]&~m[797])|(~m[752]&m[793]&~m[794]&~m[796]&m[797])|(~m[752]&~m[793]&m[794]&~m[796]&m[797])|(m[752]&m[793]&m[794]&~m[796]&m[797])|(~m[752]&m[793]&m[794]&m[796]&m[797]))&UnbiasedRNG[175])|((m[752]&~m[793]&~m[794]&m[796]&~m[797])|(~m[752]&~m[793]&~m[794]&~m[796]&m[797])|(m[752]&~m[793]&~m[794]&~m[796]&m[797])|(m[752]&m[793]&~m[794]&~m[796]&m[797])|(m[752]&~m[793]&m[794]&~m[796]&m[797])|(~m[752]&~m[793]&~m[794]&m[796]&m[797])|(m[752]&~m[793]&~m[794]&m[796]&m[797])|(~m[752]&m[793]&~m[794]&m[796]&m[797])|(m[752]&m[793]&~m[794]&m[796]&m[797])|(~m[752]&~m[793]&m[794]&m[796]&m[797])|(m[752]&~m[793]&m[794]&m[796]&m[797])|(m[752]&m[793]&m[794]&m[796]&m[797]));
    m[805] = (((m[757]&~m[803]&~m[804]&~m[806]&~m[807])|(~m[757]&~m[803]&~m[804]&m[806]&~m[807])|(m[757]&m[803]&~m[804]&m[806]&~m[807])|(m[757]&~m[803]&m[804]&m[806]&~m[807])|(~m[757]&m[803]&~m[804]&~m[806]&m[807])|(~m[757]&~m[803]&m[804]&~m[806]&m[807])|(m[757]&m[803]&m[804]&~m[806]&m[807])|(~m[757]&m[803]&m[804]&m[806]&m[807]))&UnbiasedRNG[176])|((m[757]&~m[803]&~m[804]&m[806]&~m[807])|(~m[757]&~m[803]&~m[804]&~m[806]&m[807])|(m[757]&~m[803]&~m[804]&~m[806]&m[807])|(m[757]&m[803]&~m[804]&~m[806]&m[807])|(m[757]&~m[803]&m[804]&~m[806]&m[807])|(~m[757]&~m[803]&~m[804]&m[806]&m[807])|(m[757]&~m[803]&~m[804]&m[806]&m[807])|(~m[757]&m[803]&~m[804]&m[806]&m[807])|(m[757]&m[803]&~m[804]&m[806]&m[807])|(~m[757]&~m[803]&m[804]&m[806]&m[807])|(m[757]&~m[803]&m[804]&m[806]&m[807])|(m[757]&m[803]&m[804]&m[806]&m[807]));
    m[810] = (((m[762]&~m[808]&~m[809]&~m[811]&~m[812])|(~m[762]&~m[808]&~m[809]&m[811]&~m[812])|(m[762]&m[808]&~m[809]&m[811]&~m[812])|(m[762]&~m[808]&m[809]&m[811]&~m[812])|(~m[762]&m[808]&~m[809]&~m[811]&m[812])|(~m[762]&~m[808]&m[809]&~m[811]&m[812])|(m[762]&m[808]&m[809]&~m[811]&m[812])|(~m[762]&m[808]&m[809]&m[811]&m[812]))&UnbiasedRNG[177])|((m[762]&~m[808]&~m[809]&m[811]&~m[812])|(~m[762]&~m[808]&~m[809]&~m[811]&m[812])|(m[762]&~m[808]&~m[809]&~m[811]&m[812])|(m[762]&m[808]&~m[809]&~m[811]&m[812])|(m[762]&~m[808]&m[809]&~m[811]&m[812])|(~m[762]&~m[808]&~m[809]&m[811]&m[812])|(m[762]&~m[808]&~m[809]&m[811]&m[812])|(~m[762]&m[808]&~m[809]&m[811]&m[812])|(m[762]&m[808]&~m[809]&m[811]&m[812])|(~m[762]&~m[808]&m[809]&m[811]&m[812])|(m[762]&~m[808]&m[809]&m[811]&m[812])|(m[762]&m[808]&m[809]&m[811]&m[812]));
    m[815] = (((m[767]&~m[813]&~m[814]&~m[816]&~m[817])|(~m[767]&~m[813]&~m[814]&m[816]&~m[817])|(m[767]&m[813]&~m[814]&m[816]&~m[817])|(m[767]&~m[813]&m[814]&m[816]&~m[817])|(~m[767]&m[813]&~m[814]&~m[816]&m[817])|(~m[767]&~m[813]&m[814]&~m[816]&m[817])|(m[767]&m[813]&m[814]&~m[816]&m[817])|(~m[767]&m[813]&m[814]&m[816]&m[817]))&UnbiasedRNG[178])|((m[767]&~m[813]&~m[814]&m[816]&~m[817])|(~m[767]&~m[813]&~m[814]&~m[816]&m[817])|(m[767]&~m[813]&~m[814]&~m[816]&m[817])|(m[767]&m[813]&~m[814]&~m[816]&m[817])|(m[767]&~m[813]&m[814]&~m[816]&m[817])|(~m[767]&~m[813]&~m[814]&m[816]&m[817])|(m[767]&~m[813]&~m[814]&m[816]&m[817])|(~m[767]&m[813]&~m[814]&m[816]&m[817])|(m[767]&m[813]&~m[814]&m[816]&m[817])|(~m[767]&~m[813]&m[814]&m[816]&m[817])|(m[767]&~m[813]&m[814]&m[816]&m[817])|(m[767]&m[813]&m[814]&m[816]&m[817]));
    m[820] = (((m[772]&~m[818]&~m[819]&~m[821]&~m[822])|(~m[772]&~m[818]&~m[819]&m[821]&~m[822])|(m[772]&m[818]&~m[819]&m[821]&~m[822])|(m[772]&~m[818]&m[819]&m[821]&~m[822])|(~m[772]&m[818]&~m[819]&~m[821]&m[822])|(~m[772]&~m[818]&m[819]&~m[821]&m[822])|(m[772]&m[818]&m[819]&~m[821]&m[822])|(~m[772]&m[818]&m[819]&m[821]&m[822]))&UnbiasedRNG[179])|((m[772]&~m[818]&~m[819]&m[821]&~m[822])|(~m[772]&~m[818]&~m[819]&~m[821]&m[822])|(m[772]&~m[818]&~m[819]&~m[821]&m[822])|(m[772]&m[818]&~m[819]&~m[821]&m[822])|(m[772]&~m[818]&m[819]&~m[821]&m[822])|(~m[772]&~m[818]&~m[819]&m[821]&m[822])|(m[772]&~m[818]&~m[819]&m[821]&m[822])|(~m[772]&m[818]&~m[819]&m[821]&m[822])|(m[772]&m[818]&~m[819]&m[821]&m[822])|(~m[772]&~m[818]&m[819]&m[821]&m[822])|(m[772]&~m[818]&m[819]&m[821]&m[822])|(m[772]&m[818]&m[819]&m[821]&m[822]));
    m[825] = (((m[777]&~m[823]&~m[824]&~m[826]&~m[827])|(~m[777]&~m[823]&~m[824]&m[826]&~m[827])|(m[777]&m[823]&~m[824]&m[826]&~m[827])|(m[777]&~m[823]&m[824]&m[826]&~m[827])|(~m[777]&m[823]&~m[824]&~m[826]&m[827])|(~m[777]&~m[823]&m[824]&~m[826]&m[827])|(m[777]&m[823]&m[824]&~m[826]&m[827])|(~m[777]&m[823]&m[824]&m[826]&m[827]))&UnbiasedRNG[180])|((m[777]&~m[823]&~m[824]&m[826]&~m[827])|(~m[777]&~m[823]&~m[824]&~m[826]&m[827])|(m[777]&~m[823]&~m[824]&~m[826]&m[827])|(m[777]&m[823]&~m[824]&~m[826]&m[827])|(m[777]&~m[823]&m[824]&~m[826]&m[827])|(~m[777]&~m[823]&~m[824]&m[826]&m[827])|(m[777]&~m[823]&~m[824]&m[826]&m[827])|(~m[777]&m[823]&~m[824]&m[826]&m[827])|(m[777]&m[823]&~m[824]&m[826]&m[827])|(~m[777]&~m[823]&m[824]&m[826]&m[827])|(m[777]&~m[823]&m[824]&m[826]&m[827])|(m[777]&m[823]&m[824]&m[826]&m[827]));
    m[830] = (((m[782]&~m[828]&~m[829]&~m[831]&~m[832])|(~m[782]&~m[828]&~m[829]&m[831]&~m[832])|(m[782]&m[828]&~m[829]&m[831]&~m[832])|(m[782]&~m[828]&m[829]&m[831]&~m[832])|(~m[782]&m[828]&~m[829]&~m[831]&m[832])|(~m[782]&~m[828]&m[829]&~m[831]&m[832])|(m[782]&m[828]&m[829]&~m[831]&m[832])|(~m[782]&m[828]&m[829]&m[831]&m[832]))&UnbiasedRNG[181])|((m[782]&~m[828]&~m[829]&m[831]&~m[832])|(~m[782]&~m[828]&~m[829]&~m[831]&m[832])|(m[782]&~m[828]&~m[829]&~m[831]&m[832])|(m[782]&m[828]&~m[829]&~m[831]&m[832])|(m[782]&~m[828]&m[829]&~m[831]&m[832])|(~m[782]&~m[828]&~m[829]&m[831]&m[832])|(m[782]&~m[828]&~m[829]&m[831]&m[832])|(~m[782]&m[828]&~m[829]&m[831]&m[832])|(m[782]&m[828]&~m[829]&m[831]&m[832])|(~m[782]&~m[828]&m[829]&m[831]&m[832])|(m[782]&~m[828]&m[829]&m[831]&m[832])|(m[782]&m[828]&m[829]&m[831]&m[832]));
    m[835] = (((m[787]&~m[833]&~m[834]&~m[836]&~m[837])|(~m[787]&~m[833]&~m[834]&m[836]&~m[837])|(m[787]&m[833]&~m[834]&m[836]&~m[837])|(m[787]&~m[833]&m[834]&m[836]&~m[837])|(~m[787]&m[833]&~m[834]&~m[836]&m[837])|(~m[787]&~m[833]&m[834]&~m[836]&m[837])|(m[787]&m[833]&m[834]&~m[836]&m[837])|(~m[787]&m[833]&m[834]&m[836]&m[837]))&UnbiasedRNG[182])|((m[787]&~m[833]&~m[834]&m[836]&~m[837])|(~m[787]&~m[833]&~m[834]&~m[836]&m[837])|(m[787]&~m[833]&~m[834]&~m[836]&m[837])|(m[787]&m[833]&~m[834]&~m[836]&m[837])|(m[787]&~m[833]&m[834]&~m[836]&m[837])|(~m[787]&~m[833]&~m[834]&m[836]&m[837])|(m[787]&~m[833]&~m[834]&m[836]&m[837])|(~m[787]&m[833]&~m[834]&m[836]&m[837])|(m[787]&m[833]&~m[834]&m[836]&m[837])|(~m[787]&~m[833]&m[834]&m[836]&m[837])|(m[787]&~m[833]&m[834]&m[836]&m[837])|(m[787]&m[833]&m[834]&m[836]&m[837]));
    m[840] = (((m[792]&~m[838]&~m[839]&~m[841]&~m[842])|(~m[792]&~m[838]&~m[839]&m[841]&~m[842])|(m[792]&m[838]&~m[839]&m[841]&~m[842])|(m[792]&~m[838]&m[839]&m[841]&~m[842])|(~m[792]&m[838]&~m[839]&~m[841]&m[842])|(~m[792]&~m[838]&m[839]&~m[841]&m[842])|(m[792]&m[838]&m[839]&~m[841]&m[842])|(~m[792]&m[838]&m[839]&m[841]&m[842]))&UnbiasedRNG[183])|((m[792]&~m[838]&~m[839]&m[841]&~m[842])|(~m[792]&~m[838]&~m[839]&~m[841]&m[842])|(m[792]&~m[838]&~m[839]&~m[841]&m[842])|(m[792]&m[838]&~m[839]&~m[841]&m[842])|(m[792]&~m[838]&m[839]&~m[841]&m[842])|(~m[792]&~m[838]&~m[839]&m[841]&m[842])|(m[792]&~m[838]&~m[839]&m[841]&m[842])|(~m[792]&m[838]&~m[839]&m[841]&m[842])|(m[792]&m[838]&~m[839]&m[841]&m[842])|(~m[792]&~m[838]&m[839]&m[841]&m[842])|(m[792]&~m[838]&m[839]&m[841]&m[842])|(m[792]&m[838]&m[839]&m[841]&m[842]));
    m[845] = (((m[797]&~m[843]&~m[844]&~m[846]&~m[847])|(~m[797]&~m[843]&~m[844]&m[846]&~m[847])|(m[797]&m[843]&~m[844]&m[846]&~m[847])|(m[797]&~m[843]&m[844]&m[846]&~m[847])|(~m[797]&m[843]&~m[844]&~m[846]&m[847])|(~m[797]&~m[843]&m[844]&~m[846]&m[847])|(m[797]&m[843]&m[844]&~m[846]&m[847])|(~m[797]&m[843]&m[844]&m[846]&m[847]))&UnbiasedRNG[184])|((m[797]&~m[843]&~m[844]&m[846]&~m[847])|(~m[797]&~m[843]&~m[844]&~m[846]&m[847])|(m[797]&~m[843]&~m[844]&~m[846]&m[847])|(m[797]&m[843]&~m[844]&~m[846]&m[847])|(m[797]&~m[843]&m[844]&~m[846]&m[847])|(~m[797]&~m[843]&~m[844]&m[846]&m[847])|(m[797]&~m[843]&~m[844]&m[846]&m[847])|(~m[797]&m[843]&~m[844]&m[846]&m[847])|(m[797]&m[843]&~m[844]&m[846]&m[847])|(~m[797]&~m[843]&m[844]&m[846]&m[847])|(m[797]&~m[843]&m[844]&m[846]&m[847])|(m[797]&m[843]&m[844]&m[846]&m[847]));
    m[850] = (((m[802]&~m[848]&~m[849]&~m[851]&~m[852])|(~m[802]&~m[848]&~m[849]&m[851]&~m[852])|(m[802]&m[848]&~m[849]&m[851]&~m[852])|(m[802]&~m[848]&m[849]&m[851]&~m[852])|(~m[802]&m[848]&~m[849]&~m[851]&m[852])|(~m[802]&~m[848]&m[849]&~m[851]&m[852])|(m[802]&m[848]&m[849]&~m[851]&m[852])|(~m[802]&m[848]&m[849]&m[851]&m[852]))&UnbiasedRNG[185])|((m[802]&~m[848]&~m[849]&m[851]&~m[852])|(~m[802]&~m[848]&~m[849]&~m[851]&m[852])|(m[802]&~m[848]&~m[849]&~m[851]&m[852])|(m[802]&m[848]&~m[849]&~m[851]&m[852])|(m[802]&~m[848]&m[849]&~m[851]&m[852])|(~m[802]&~m[848]&~m[849]&m[851]&m[852])|(m[802]&~m[848]&~m[849]&m[851]&m[852])|(~m[802]&m[848]&~m[849]&m[851]&m[852])|(m[802]&m[848]&~m[849]&m[851]&m[852])|(~m[802]&~m[848]&m[849]&m[851]&m[852])|(m[802]&~m[848]&m[849]&m[851]&m[852])|(m[802]&m[848]&m[849]&m[851]&m[852]));
    m[860] = (((m[807]&~m[858]&~m[859]&~m[861]&~m[862])|(~m[807]&~m[858]&~m[859]&m[861]&~m[862])|(m[807]&m[858]&~m[859]&m[861]&~m[862])|(m[807]&~m[858]&m[859]&m[861]&~m[862])|(~m[807]&m[858]&~m[859]&~m[861]&m[862])|(~m[807]&~m[858]&m[859]&~m[861]&m[862])|(m[807]&m[858]&m[859]&~m[861]&m[862])|(~m[807]&m[858]&m[859]&m[861]&m[862]))&UnbiasedRNG[186])|((m[807]&~m[858]&~m[859]&m[861]&~m[862])|(~m[807]&~m[858]&~m[859]&~m[861]&m[862])|(m[807]&~m[858]&~m[859]&~m[861]&m[862])|(m[807]&m[858]&~m[859]&~m[861]&m[862])|(m[807]&~m[858]&m[859]&~m[861]&m[862])|(~m[807]&~m[858]&~m[859]&m[861]&m[862])|(m[807]&~m[858]&~m[859]&m[861]&m[862])|(~m[807]&m[858]&~m[859]&m[861]&m[862])|(m[807]&m[858]&~m[859]&m[861]&m[862])|(~m[807]&~m[858]&m[859]&m[861]&m[862])|(m[807]&~m[858]&m[859]&m[861]&m[862])|(m[807]&m[858]&m[859]&m[861]&m[862]));
    m[865] = (((m[812]&~m[863]&~m[864]&~m[866]&~m[867])|(~m[812]&~m[863]&~m[864]&m[866]&~m[867])|(m[812]&m[863]&~m[864]&m[866]&~m[867])|(m[812]&~m[863]&m[864]&m[866]&~m[867])|(~m[812]&m[863]&~m[864]&~m[866]&m[867])|(~m[812]&~m[863]&m[864]&~m[866]&m[867])|(m[812]&m[863]&m[864]&~m[866]&m[867])|(~m[812]&m[863]&m[864]&m[866]&m[867]))&UnbiasedRNG[187])|((m[812]&~m[863]&~m[864]&m[866]&~m[867])|(~m[812]&~m[863]&~m[864]&~m[866]&m[867])|(m[812]&~m[863]&~m[864]&~m[866]&m[867])|(m[812]&m[863]&~m[864]&~m[866]&m[867])|(m[812]&~m[863]&m[864]&~m[866]&m[867])|(~m[812]&~m[863]&~m[864]&m[866]&m[867])|(m[812]&~m[863]&~m[864]&m[866]&m[867])|(~m[812]&m[863]&~m[864]&m[866]&m[867])|(m[812]&m[863]&~m[864]&m[866]&m[867])|(~m[812]&~m[863]&m[864]&m[866]&m[867])|(m[812]&~m[863]&m[864]&m[866]&m[867])|(m[812]&m[863]&m[864]&m[866]&m[867]));
    m[870] = (((m[817]&~m[868]&~m[869]&~m[871]&~m[872])|(~m[817]&~m[868]&~m[869]&m[871]&~m[872])|(m[817]&m[868]&~m[869]&m[871]&~m[872])|(m[817]&~m[868]&m[869]&m[871]&~m[872])|(~m[817]&m[868]&~m[869]&~m[871]&m[872])|(~m[817]&~m[868]&m[869]&~m[871]&m[872])|(m[817]&m[868]&m[869]&~m[871]&m[872])|(~m[817]&m[868]&m[869]&m[871]&m[872]))&UnbiasedRNG[188])|((m[817]&~m[868]&~m[869]&m[871]&~m[872])|(~m[817]&~m[868]&~m[869]&~m[871]&m[872])|(m[817]&~m[868]&~m[869]&~m[871]&m[872])|(m[817]&m[868]&~m[869]&~m[871]&m[872])|(m[817]&~m[868]&m[869]&~m[871]&m[872])|(~m[817]&~m[868]&~m[869]&m[871]&m[872])|(m[817]&~m[868]&~m[869]&m[871]&m[872])|(~m[817]&m[868]&~m[869]&m[871]&m[872])|(m[817]&m[868]&~m[869]&m[871]&m[872])|(~m[817]&~m[868]&m[869]&m[871]&m[872])|(m[817]&~m[868]&m[869]&m[871]&m[872])|(m[817]&m[868]&m[869]&m[871]&m[872]));
    m[875] = (((m[822]&~m[873]&~m[874]&~m[876]&~m[877])|(~m[822]&~m[873]&~m[874]&m[876]&~m[877])|(m[822]&m[873]&~m[874]&m[876]&~m[877])|(m[822]&~m[873]&m[874]&m[876]&~m[877])|(~m[822]&m[873]&~m[874]&~m[876]&m[877])|(~m[822]&~m[873]&m[874]&~m[876]&m[877])|(m[822]&m[873]&m[874]&~m[876]&m[877])|(~m[822]&m[873]&m[874]&m[876]&m[877]))&UnbiasedRNG[189])|((m[822]&~m[873]&~m[874]&m[876]&~m[877])|(~m[822]&~m[873]&~m[874]&~m[876]&m[877])|(m[822]&~m[873]&~m[874]&~m[876]&m[877])|(m[822]&m[873]&~m[874]&~m[876]&m[877])|(m[822]&~m[873]&m[874]&~m[876]&m[877])|(~m[822]&~m[873]&~m[874]&m[876]&m[877])|(m[822]&~m[873]&~m[874]&m[876]&m[877])|(~m[822]&m[873]&~m[874]&m[876]&m[877])|(m[822]&m[873]&~m[874]&m[876]&m[877])|(~m[822]&~m[873]&m[874]&m[876]&m[877])|(m[822]&~m[873]&m[874]&m[876]&m[877])|(m[822]&m[873]&m[874]&m[876]&m[877]));
    m[880] = (((m[827]&~m[878]&~m[879]&~m[881]&~m[882])|(~m[827]&~m[878]&~m[879]&m[881]&~m[882])|(m[827]&m[878]&~m[879]&m[881]&~m[882])|(m[827]&~m[878]&m[879]&m[881]&~m[882])|(~m[827]&m[878]&~m[879]&~m[881]&m[882])|(~m[827]&~m[878]&m[879]&~m[881]&m[882])|(m[827]&m[878]&m[879]&~m[881]&m[882])|(~m[827]&m[878]&m[879]&m[881]&m[882]))&UnbiasedRNG[190])|((m[827]&~m[878]&~m[879]&m[881]&~m[882])|(~m[827]&~m[878]&~m[879]&~m[881]&m[882])|(m[827]&~m[878]&~m[879]&~m[881]&m[882])|(m[827]&m[878]&~m[879]&~m[881]&m[882])|(m[827]&~m[878]&m[879]&~m[881]&m[882])|(~m[827]&~m[878]&~m[879]&m[881]&m[882])|(m[827]&~m[878]&~m[879]&m[881]&m[882])|(~m[827]&m[878]&~m[879]&m[881]&m[882])|(m[827]&m[878]&~m[879]&m[881]&m[882])|(~m[827]&~m[878]&m[879]&m[881]&m[882])|(m[827]&~m[878]&m[879]&m[881]&m[882])|(m[827]&m[878]&m[879]&m[881]&m[882]));
    m[885] = (((m[832]&~m[883]&~m[884]&~m[886]&~m[887])|(~m[832]&~m[883]&~m[884]&m[886]&~m[887])|(m[832]&m[883]&~m[884]&m[886]&~m[887])|(m[832]&~m[883]&m[884]&m[886]&~m[887])|(~m[832]&m[883]&~m[884]&~m[886]&m[887])|(~m[832]&~m[883]&m[884]&~m[886]&m[887])|(m[832]&m[883]&m[884]&~m[886]&m[887])|(~m[832]&m[883]&m[884]&m[886]&m[887]))&UnbiasedRNG[191])|((m[832]&~m[883]&~m[884]&m[886]&~m[887])|(~m[832]&~m[883]&~m[884]&~m[886]&m[887])|(m[832]&~m[883]&~m[884]&~m[886]&m[887])|(m[832]&m[883]&~m[884]&~m[886]&m[887])|(m[832]&~m[883]&m[884]&~m[886]&m[887])|(~m[832]&~m[883]&~m[884]&m[886]&m[887])|(m[832]&~m[883]&~m[884]&m[886]&m[887])|(~m[832]&m[883]&~m[884]&m[886]&m[887])|(m[832]&m[883]&~m[884]&m[886]&m[887])|(~m[832]&~m[883]&m[884]&m[886]&m[887])|(m[832]&~m[883]&m[884]&m[886]&m[887])|(m[832]&m[883]&m[884]&m[886]&m[887]));
    m[890] = (((m[837]&~m[888]&~m[889]&~m[891]&~m[892])|(~m[837]&~m[888]&~m[889]&m[891]&~m[892])|(m[837]&m[888]&~m[889]&m[891]&~m[892])|(m[837]&~m[888]&m[889]&m[891]&~m[892])|(~m[837]&m[888]&~m[889]&~m[891]&m[892])|(~m[837]&~m[888]&m[889]&~m[891]&m[892])|(m[837]&m[888]&m[889]&~m[891]&m[892])|(~m[837]&m[888]&m[889]&m[891]&m[892]))&UnbiasedRNG[192])|((m[837]&~m[888]&~m[889]&m[891]&~m[892])|(~m[837]&~m[888]&~m[889]&~m[891]&m[892])|(m[837]&~m[888]&~m[889]&~m[891]&m[892])|(m[837]&m[888]&~m[889]&~m[891]&m[892])|(m[837]&~m[888]&m[889]&~m[891]&m[892])|(~m[837]&~m[888]&~m[889]&m[891]&m[892])|(m[837]&~m[888]&~m[889]&m[891]&m[892])|(~m[837]&m[888]&~m[889]&m[891]&m[892])|(m[837]&m[888]&~m[889]&m[891]&m[892])|(~m[837]&~m[888]&m[889]&m[891]&m[892])|(m[837]&~m[888]&m[889]&m[891]&m[892])|(m[837]&m[888]&m[889]&m[891]&m[892]));
    m[895] = (((m[842]&~m[893]&~m[894]&~m[896]&~m[897])|(~m[842]&~m[893]&~m[894]&m[896]&~m[897])|(m[842]&m[893]&~m[894]&m[896]&~m[897])|(m[842]&~m[893]&m[894]&m[896]&~m[897])|(~m[842]&m[893]&~m[894]&~m[896]&m[897])|(~m[842]&~m[893]&m[894]&~m[896]&m[897])|(m[842]&m[893]&m[894]&~m[896]&m[897])|(~m[842]&m[893]&m[894]&m[896]&m[897]))&UnbiasedRNG[193])|((m[842]&~m[893]&~m[894]&m[896]&~m[897])|(~m[842]&~m[893]&~m[894]&~m[896]&m[897])|(m[842]&~m[893]&~m[894]&~m[896]&m[897])|(m[842]&m[893]&~m[894]&~m[896]&m[897])|(m[842]&~m[893]&m[894]&~m[896]&m[897])|(~m[842]&~m[893]&~m[894]&m[896]&m[897])|(m[842]&~m[893]&~m[894]&m[896]&m[897])|(~m[842]&m[893]&~m[894]&m[896]&m[897])|(m[842]&m[893]&~m[894]&m[896]&m[897])|(~m[842]&~m[893]&m[894]&m[896]&m[897])|(m[842]&~m[893]&m[894]&m[896]&m[897])|(m[842]&m[893]&m[894]&m[896]&m[897]));
    m[900] = (((m[847]&~m[898]&~m[899]&~m[901]&~m[902])|(~m[847]&~m[898]&~m[899]&m[901]&~m[902])|(m[847]&m[898]&~m[899]&m[901]&~m[902])|(m[847]&~m[898]&m[899]&m[901]&~m[902])|(~m[847]&m[898]&~m[899]&~m[901]&m[902])|(~m[847]&~m[898]&m[899]&~m[901]&m[902])|(m[847]&m[898]&m[899]&~m[901]&m[902])|(~m[847]&m[898]&m[899]&m[901]&m[902]))&UnbiasedRNG[194])|((m[847]&~m[898]&~m[899]&m[901]&~m[902])|(~m[847]&~m[898]&~m[899]&~m[901]&m[902])|(m[847]&~m[898]&~m[899]&~m[901]&m[902])|(m[847]&m[898]&~m[899]&~m[901]&m[902])|(m[847]&~m[898]&m[899]&~m[901]&m[902])|(~m[847]&~m[898]&~m[899]&m[901]&m[902])|(m[847]&~m[898]&~m[899]&m[901]&m[902])|(~m[847]&m[898]&~m[899]&m[901]&m[902])|(m[847]&m[898]&~m[899]&m[901]&m[902])|(~m[847]&~m[898]&m[899]&m[901]&m[902])|(m[847]&~m[898]&m[899]&m[901]&m[902])|(m[847]&m[898]&m[899]&m[901]&m[902]));
    m[905] = (((m[852]&~m[903]&~m[904]&~m[906]&~m[907])|(~m[852]&~m[903]&~m[904]&m[906]&~m[907])|(m[852]&m[903]&~m[904]&m[906]&~m[907])|(m[852]&~m[903]&m[904]&m[906]&~m[907])|(~m[852]&m[903]&~m[904]&~m[906]&m[907])|(~m[852]&~m[903]&m[904]&~m[906]&m[907])|(m[852]&m[903]&m[904]&~m[906]&m[907])|(~m[852]&m[903]&m[904]&m[906]&m[907]))&UnbiasedRNG[195])|((m[852]&~m[903]&~m[904]&m[906]&~m[907])|(~m[852]&~m[903]&~m[904]&~m[906]&m[907])|(m[852]&~m[903]&~m[904]&~m[906]&m[907])|(m[852]&m[903]&~m[904]&~m[906]&m[907])|(m[852]&~m[903]&m[904]&~m[906]&m[907])|(~m[852]&~m[903]&~m[904]&m[906]&m[907])|(m[852]&~m[903]&~m[904]&m[906]&m[907])|(~m[852]&m[903]&~m[904]&m[906]&m[907])|(m[852]&m[903]&~m[904]&m[906]&m[907])|(~m[852]&~m[903]&m[904]&m[906]&m[907])|(m[852]&~m[903]&m[904]&m[906]&m[907])|(m[852]&m[903]&m[904]&m[906]&m[907]));
    m[910] = (((m[857]&~m[908]&~m[909]&~m[911]&~m[912])|(~m[857]&~m[908]&~m[909]&m[911]&~m[912])|(m[857]&m[908]&~m[909]&m[911]&~m[912])|(m[857]&~m[908]&m[909]&m[911]&~m[912])|(~m[857]&m[908]&~m[909]&~m[911]&m[912])|(~m[857]&~m[908]&m[909]&~m[911]&m[912])|(m[857]&m[908]&m[909]&~m[911]&m[912])|(~m[857]&m[908]&m[909]&m[911]&m[912]))&UnbiasedRNG[196])|((m[857]&~m[908]&~m[909]&m[911]&~m[912])|(~m[857]&~m[908]&~m[909]&~m[911]&m[912])|(m[857]&~m[908]&~m[909]&~m[911]&m[912])|(m[857]&m[908]&~m[909]&~m[911]&m[912])|(m[857]&~m[908]&m[909]&~m[911]&m[912])|(~m[857]&~m[908]&~m[909]&m[911]&m[912])|(m[857]&~m[908]&~m[909]&m[911]&m[912])|(~m[857]&m[908]&~m[909]&m[911]&m[912])|(m[857]&m[908]&~m[909]&m[911]&m[912])|(~m[857]&~m[908]&m[909]&m[911]&m[912])|(m[857]&~m[908]&m[909]&m[911]&m[912])|(m[857]&m[908]&m[909]&m[911]&m[912]));
    m[915] = (((m[867]&~m[913]&~m[914]&~m[916]&~m[917])|(~m[867]&~m[913]&~m[914]&m[916]&~m[917])|(m[867]&m[913]&~m[914]&m[916]&~m[917])|(m[867]&~m[913]&m[914]&m[916]&~m[917])|(~m[867]&m[913]&~m[914]&~m[916]&m[917])|(~m[867]&~m[913]&m[914]&~m[916]&m[917])|(m[867]&m[913]&m[914]&~m[916]&m[917])|(~m[867]&m[913]&m[914]&m[916]&m[917]))&UnbiasedRNG[197])|((m[867]&~m[913]&~m[914]&m[916]&~m[917])|(~m[867]&~m[913]&~m[914]&~m[916]&m[917])|(m[867]&~m[913]&~m[914]&~m[916]&m[917])|(m[867]&m[913]&~m[914]&~m[916]&m[917])|(m[867]&~m[913]&m[914]&~m[916]&m[917])|(~m[867]&~m[913]&~m[914]&m[916]&m[917])|(m[867]&~m[913]&~m[914]&m[916]&m[917])|(~m[867]&m[913]&~m[914]&m[916]&m[917])|(m[867]&m[913]&~m[914]&m[916]&m[917])|(~m[867]&~m[913]&m[914]&m[916]&m[917])|(m[867]&~m[913]&m[914]&m[916]&m[917])|(m[867]&m[913]&m[914]&m[916]&m[917]));
    m[920] = (((m[872]&~m[918]&~m[919]&~m[921]&~m[922])|(~m[872]&~m[918]&~m[919]&m[921]&~m[922])|(m[872]&m[918]&~m[919]&m[921]&~m[922])|(m[872]&~m[918]&m[919]&m[921]&~m[922])|(~m[872]&m[918]&~m[919]&~m[921]&m[922])|(~m[872]&~m[918]&m[919]&~m[921]&m[922])|(m[872]&m[918]&m[919]&~m[921]&m[922])|(~m[872]&m[918]&m[919]&m[921]&m[922]))&UnbiasedRNG[198])|((m[872]&~m[918]&~m[919]&m[921]&~m[922])|(~m[872]&~m[918]&~m[919]&~m[921]&m[922])|(m[872]&~m[918]&~m[919]&~m[921]&m[922])|(m[872]&m[918]&~m[919]&~m[921]&m[922])|(m[872]&~m[918]&m[919]&~m[921]&m[922])|(~m[872]&~m[918]&~m[919]&m[921]&m[922])|(m[872]&~m[918]&~m[919]&m[921]&m[922])|(~m[872]&m[918]&~m[919]&m[921]&m[922])|(m[872]&m[918]&~m[919]&m[921]&m[922])|(~m[872]&~m[918]&m[919]&m[921]&m[922])|(m[872]&~m[918]&m[919]&m[921]&m[922])|(m[872]&m[918]&m[919]&m[921]&m[922]));
    m[925] = (((m[877]&~m[923]&~m[924]&~m[926]&~m[927])|(~m[877]&~m[923]&~m[924]&m[926]&~m[927])|(m[877]&m[923]&~m[924]&m[926]&~m[927])|(m[877]&~m[923]&m[924]&m[926]&~m[927])|(~m[877]&m[923]&~m[924]&~m[926]&m[927])|(~m[877]&~m[923]&m[924]&~m[926]&m[927])|(m[877]&m[923]&m[924]&~m[926]&m[927])|(~m[877]&m[923]&m[924]&m[926]&m[927]))&UnbiasedRNG[199])|((m[877]&~m[923]&~m[924]&m[926]&~m[927])|(~m[877]&~m[923]&~m[924]&~m[926]&m[927])|(m[877]&~m[923]&~m[924]&~m[926]&m[927])|(m[877]&m[923]&~m[924]&~m[926]&m[927])|(m[877]&~m[923]&m[924]&~m[926]&m[927])|(~m[877]&~m[923]&~m[924]&m[926]&m[927])|(m[877]&~m[923]&~m[924]&m[926]&m[927])|(~m[877]&m[923]&~m[924]&m[926]&m[927])|(m[877]&m[923]&~m[924]&m[926]&m[927])|(~m[877]&~m[923]&m[924]&m[926]&m[927])|(m[877]&~m[923]&m[924]&m[926]&m[927])|(m[877]&m[923]&m[924]&m[926]&m[927]));
    m[930] = (((m[882]&~m[928]&~m[929]&~m[931]&~m[932])|(~m[882]&~m[928]&~m[929]&m[931]&~m[932])|(m[882]&m[928]&~m[929]&m[931]&~m[932])|(m[882]&~m[928]&m[929]&m[931]&~m[932])|(~m[882]&m[928]&~m[929]&~m[931]&m[932])|(~m[882]&~m[928]&m[929]&~m[931]&m[932])|(m[882]&m[928]&m[929]&~m[931]&m[932])|(~m[882]&m[928]&m[929]&m[931]&m[932]))&UnbiasedRNG[200])|((m[882]&~m[928]&~m[929]&m[931]&~m[932])|(~m[882]&~m[928]&~m[929]&~m[931]&m[932])|(m[882]&~m[928]&~m[929]&~m[931]&m[932])|(m[882]&m[928]&~m[929]&~m[931]&m[932])|(m[882]&~m[928]&m[929]&~m[931]&m[932])|(~m[882]&~m[928]&~m[929]&m[931]&m[932])|(m[882]&~m[928]&~m[929]&m[931]&m[932])|(~m[882]&m[928]&~m[929]&m[931]&m[932])|(m[882]&m[928]&~m[929]&m[931]&m[932])|(~m[882]&~m[928]&m[929]&m[931]&m[932])|(m[882]&~m[928]&m[929]&m[931]&m[932])|(m[882]&m[928]&m[929]&m[931]&m[932]));
    m[935] = (((m[887]&~m[933]&~m[934]&~m[936]&~m[937])|(~m[887]&~m[933]&~m[934]&m[936]&~m[937])|(m[887]&m[933]&~m[934]&m[936]&~m[937])|(m[887]&~m[933]&m[934]&m[936]&~m[937])|(~m[887]&m[933]&~m[934]&~m[936]&m[937])|(~m[887]&~m[933]&m[934]&~m[936]&m[937])|(m[887]&m[933]&m[934]&~m[936]&m[937])|(~m[887]&m[933]&m[934]&m[936]&m[937]))&UnbiasedRNG[201])|((m[887]&~m[933]&~m[934]&m[936]&~m[937])|(~m[887]&~m[933]&~m[934]&~m[936]&m[937])|(m[887]&~m[933]&~m[934]&~m[936]&m[937])|(m[887]&m[933]&~m[934]&~m[936]&m[937])|(m[887]&~m[933]&m[934]&~m[936]&m[937])|(~m[887]&~m[933]&~m[934]&m[936]&m[937])|(m[887]&~m[933]&~m[934]&m[936]&m[937])|(~m[887]&m[933]&~m[934]&m[936]&m[937])|(m[887]&m[933]&~m[934]&m[936]&m[937])|(~m[887]&~m[933]&m[934]&m[936]&m[937])|(m[887]&~m[933]&m[934]&m[936]&m[937])|(m[887]&m[933]&m[934]&m[936]&m[937]));
    m[940] = (((m[892]&~m[938]&~m[939]&~m[941]&~m[942])|(~m[892]&~m[938]&~m[939]&m[941]&~m[942])|(m[892]&m[938]&~m[939]&m[941]&~m[942])|(m[892]&~m[938]&m[939]&m[941]&~m[942])|(~m[892]&m[938]&~m[939]&~m[941]&m[942])|(~m[892]&~m[938]&m[939]&~m[941]&m[942])|(m[892]&m[938]&m[939]&~m[941]&m[942])|(~m[892]&m[938]&m[939]&m[941]&m[942]))&UnbiasedRNG[202])|((m[892]&~m[938]&~m[939]&m[941]&~m[942])|(~m[892]&~m[938]&~m[939]&~m[941]&m[942])|(m[892]&~m[938]&~m[939]&~m[941]&m[942])|(m[892]&m[938]&~m[939]&~m[941]&m[942])|(m[892]&~m[938]&m[939]&~m[941]&m[942])|(~m[892]&~m[938]&~m[939]&m[941]&m[942])|(m[892]&~m[938]&~m[939]&m[941]&m[942])|(~m[892]&m[938]&~m[939]&m[941]&m[942])|(m[892]&m[938]&~m[939]&m[941]&m[942])|(~m[892]&~m[938]&m[939]&m[941]&m[942])|(m[892]&~m[938]&m[939]&m[941]&m[942])|(m[892]&m[938]&m[939]&m[941]&m[942]));
    m[945] = (((m[897]&~m[943]&~m[944]&~m[946]&~m[947])|(~m[897]&~m[943]&~m[944]&m[946]&~m[947])|(m[897]&m[943]&~m[944]&m[946]&~m[947])|(m[897]&~m[943]&m[944]&m[946]&~m[947])|(~m[897]&m[943]&~m[944]&~m[946]&m[947])|(~m[897]&~m[943]&m[944]&~m[946]&m[947])|(m[897]&m[943]&m[944]&~m[946]&m[947])|(~m[897]&m[943]&m[944]&m[946]&m[947]))&UnbiasedRNG[203])|((m[897]&~m[943]&~m[944]&m[946]&~m[947])|(~m[897]&~m[943]&~m[944]&~m[946]&m[947])|(m[897]&~m[943]&~m[944]&~m[946]&m[947])|(m[897]&m[943]&~m[944]&~m[946]&m[947])|(m[897]&~m[943]&m[944]&~m[946]&m[947])|(~m[897]&~m[943]&~m[944]&m[946]&m[947])|(m[897]&~m[943]&~m[944]&m[946]&m[947])|(~m[897]&m[943]&~m[944]&m[946]&m[947])|(m[897]&m[943]&~m[944]&m[946]&m[947])|(~m[897]&~m[943]&m[944]&m[946]&m[947])|(m[897]&~m[943]&m[944]&m[946]&m[947])|(m[897]&m[943]&m[944]&m[946]&m[947]));
    m[950] = (((m[902]&~m[948]&~m[949]&~m[951]&~m[952])|(~m[902]&~m[948]&~m[949]&m[951]&~m[952])|(m[902]&m[948]&~m[949]&m[951]&~m[952])|(m[902]&~m[948]&m[949]&m[951]&~m[952])|(~m[902]&m[948]&~m[949]&~m[951]&m[952])|(~m[902]&~m[948]&m[949]&~m[951]&m[952])|(m[902]&m[948]&m[949]&~m[951]&m[952])|(~m[902]&m[948]&m[949]&m[951]&m[952]))&UnbiasedRNG[204])|((m[902]&~m[948]&~m[949]&m[951]&~m[952])|(~m[902]&~m[948]&~m[949]&~m[951]&m[952])|(m[902]&~m[948]&~m[949]&~m[951]&m[952])|(m[902]&m[948]&~m[949]&~m[951]&m[952])|(m[902]&~m[948]&m[949]&~m[951]&m[952])|(~m[902]&~m[948]&~m[949]&m[951]&m[952])|(m[902]&~m[948]&~m[949]&m[951]&m[952])|(~m[902]&m[948]&~m[949]&m[951]&m[952])|(m[902]&m[948]&~m[949]&m[951]&m[952])|(~m[902]&~m[948]&m[949]&m[951]&m[952])|(m[902]&~m[948]&m[949]&m[951]&m[952])|(m[902]&m[948]&m[949]&m[951]&m[952]));
    m[955] = (((m[907]&~m[953]&~m[954]&~m[956]&~m[957])|(~m[907]&~m[953]&~m[954]&m[956]&~m[957])|(m[907]&m[953]&~m[954]&m[956]&~m[957])|(m[907]&~m[953]&m[954]&m[956]&~m[957])|(~m[907]&m[953]&~m[954]&~m[956]&m[957])|(~m[907]&~m[953]&m[954]&~m[956]&m[957])|(m[907]&m[953]&m[954]&~m[956]&m[957])|(~m[907]&m[953]&m[954]&m[956]&m[957]))&UnbiasedRNG[205])|((m[907]&~m[953]&~m[954]&m[956]&~m[957])|(~m[907]&~m[953]&~m[954]&~m[956]&m[957])|(m[907]&~m[953]&~m[954]&~m[956]&m[957])|(m[907]&m[953]&~m[954]&~m[956]&m[957])|(m[907]&~m[953]&m[954]&~m[956]&m[957])|(~m[907]&~m[953]&~m[954]&m[956]&m[957])|(m[907]&~m[953]&~m[954]&m[956]&m[957])|(~m[907]&m[953]&~m[954]&m[956]&m[957])|(m[907]&m[953]&~m[954]&m[956]&m[957])|(~m[907]&~m[953]&m[954]&m[956]&m[957])|(m[907]&~m[953]&m[954]&m[956]&m[957])|(m[907]&m[953]&m[954]&m[956]&m[957]));
    m[960] = (((m[912]&~m[958]&~m[959]&~m[961]&~m[962])|(~m[912]&~m[958]&~m[959]&m[961]&~m[962])|(m[912]&m[958]&~m[959]&m[961]&~m[962])|(m[912]&~m[958]&m[959]&m[961]&~m[962])|(~m[912]&m[958]&~m[959]&~m[961]&m[962])|(~m[912]&~m[958]&m[959]&~m[961]&m[962])|(m[912]&m[958]&m[959]&~m[961]&m[962])|(~m[912]&m[958]&m[959]&m[961]&m[962]))&UnbiasedRNG[206])|((m[912]&~m[958]&~m[959]&m[961]&~m[962])|(~m[912]&~m[958]&~m[959]&~m[961]&m[962])|(m[912]&~m[958]&~m[959]&~m[961]&m[962])|(m[912]&m[958]&~m[959]&~m[961]&m[962])|(m[912]&~m[958]&m[959]&~m[961]&m[962])|(~m[912]&~m[958]&~m[959]&m[961]&m[962])|(m[912]&~m[958]&~m[959]&m[961]&m[962])|(~m[912]&m[958]&~m[959]&m[961]&m[962])|(m[912]&m[958]&~m[959]&m[961]&m[962])|(~m[912]&~m[958]&m[959]&m[961]&m[962])|(m[912]&~m[958]&m[959]&m[961]&m[962])|(m[912]&m[958]&m[959]&m[961]&m[962]));
    m[965] = (((m[922]&~m[963]&~m[964]&~m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&m[966]&~m[967])|(m[922]&m[963]&~m[964]&m[966]&~m[967])|(m[922]&~m[963]&m[964]&m[966]&~m[967])|(~m[922]&m[963]&~m[964]&~m[966]&m[967])|(~m[922]&~m[963]&m[964]&~m[966]&m[967])|(m[922]&m[963]&m[964]&~m[966]&m[967])|(~m[922]&m[963]&m[964]&m[966]&m[967]))&UnbiasedRNG[207])|((m[922]&~m[963]&~m[964]&m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&m[964]&~m[966]&m[967])|(~m[922]&~m[963]&~m[964]&m[966]&m[967])|(m[922]&~m[963]&~m[964]&m[966]&m[967])|(~m[922]&m[963]&~m[964]&m[966]&m[967])|(m[922]&m[963]&~m[964]&m[966]&m[967])|(~m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&m[963]&m[964]&m[966]&m[967]));
    m[970] = (((m[927]&~m[968]&~m[969]&~m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&m[971]&~m[972])|(m[927]&m[968]&~m[969]&m[971]&~m[972])|(m[927]&~m[968]&m[969]&m[971]&~m[972])|(~m[927]&m[968]&~m[969]&~m[971]&m[972])|(~m[927]&~m[968]&m[969]&~m[971]&m[972])|(m[927]&m[968]&m[969]&~m[971]&m[972])|(~m[927]&m[968]&m[969]&m[971]&m[972]))&UnbiasedRNG[208])|((m[927]&~m[968]&~m[969]&m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&m[969]&~m[971]&m[972])|(~m[927]&~m[968]&~m[969]&m[971]&m[972])|(m[927]&~m[968]&~m[969]&m[971]&m[972])|(~m[927]&m[968]&~m[969]&m[971]&m[972])|(m[927]&m[968]&~m[969]&m[971]&m[972])|(~m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&m[968]&m[969]&m[971]&m[972]));
    m[975] = (((m[932]&~m[973]&~m[974]&~m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&m[976]&~m[977])|(m[932]&m[973]&~m[974]&m[976]&~m[977])|(m[932]&~m[973]&m[974]&m[976]&~m[977])|(~m[932]&m[973]&~m[974]&~m[976]&m[977])|(~m[932]&~m[973]&m[974]&~m[976]&m[977])|(m[932]&m[973]&m[974]&~m[976]&m[977])|(~m[932]&m[973]&m[974]&m[976]&m[977]))&UnbiasedRNG[209])|((m[932]&~m[973]&~m[974]&m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&m[974]&~m[976]&m[977])|(~m[932]&~m[973]&~m[974]&m[976]&m[977])|(m[932]&~m[973]&~m[974]&m[976]&m[977])|(~m[932]&m[973]&~m[974]&m[976]&m[977])|(m[932]&m[973]&~m[974]&m[976]&m[977])|(~m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&m[973]&m[974]&m[976]&m[977]));
    m[980] = (((m[937]&~m[978]&~m[979]&~m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&m[981]&~m[982])|(m[937]&m[978]&~m[979]&m[981]&~m[982])|(m[937]&~m[978]&m[979]&m[981]&~m[982])|(~m[937]&m[978]&~m[979]&~m[981]&m[982])|(~m[937]&~m[978]&m[979]&~m[981]&m[982])|(m[937]&m[978]&m[979]&~m[981]&m[982])|(~m[937]&m[978]&m[979]&m[981]&m[982]))&UnbiasedRNG[210])|((m[937]&~m[978]&~m[979]&m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&m[979]&~m[981]&m[982])|(~m[937]&~m[978]&~m[979]&m[981]&m[982])|(m[937]&~m[978]&~m[979]&m[981]&m[982])|(~m[937]&m[978]&~m[979]&m[981]&m[982])|(m[937]&m[978]&~m[979]&m[981]&m[982])|(~m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&m[978]&m[979]&m[981]&m[982]));
    m[985] = (((m[942]&~m[983]&~m[984]&~m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&m[986]&~m[987])|(m[942]&m[983]&~m[984]&m[986]&~m[987])|(m[942]&~m[983]&m[984]&m[986]&~m[987])|(~m[942]&m[983]&~m[984]&~m[986]&m[987])|(~m[942]&~m[983]&m[984]&~m[986]&m[987])|(m[942]&m[983]&m[984]&~m[986]&m[987])|(~m[942]&m[983]&m[984]&m[986]&m[987]))&UnbiasedRNG[211])|((m[942]&~m[983]&~m[984]&m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&m[984]&~m[986]&m[987])|(~m[942]&~m[983]&~m[984]&m[986]&m[987])|(m[942]&~m[983]&~m[984]&m[986]&m[987])|(~m[942]&m[983]&~m[984]&m[986]&m[987])|(m[942]&m[983]&~m[984]&m[986]&m[987])|(~m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&m[983]&m[984]&m[986]&m[987]));
    m[990] = (((m[947]&~m[988]&~m[989]&~m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&m[991]&~m[992])|(m[947]&m[988]&~m[989]&m[991]&~m[992])|(m[947]&~m[988]&m[989]&m[991]&~m[992])|(~m[947]&m[988]&~m[989]&~m[991]&m[992])|(~m[947]&~m[988]&m[989]&~m[991]&m[992])|(m[947]&m[988]&m[989]&~m[991]&m[992])|(~m[947]&m[988]&m[989]&m[991]&m[992]))&UnbiasedRNG[212])|((m[947]&~m[988]&~m[989]&m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&m[989]&~m[991]&m[992])|(~m[947]&~m[988]&~m[989]&m[991]&m[992])|(m[947]&~m[988]&~m[989]&m[991]&m[992])|(~m[947]&m[988]&~m[989]&m[991]&m[992])|(m[947]&m[988]&~m[989]&m[991]&m[992])|(~m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&m[988]&m[989]&m[991]&m[992]));
    m[995] = (((m[952]&~m[993]&~m[994]&~m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&m[996]&~m[997])|(m[952]&m[993]&~m[994]&m[996]&~m[997])|(m[952]&~m[993]&m[994]&m[996]&~m[997])|(~m[952]&m[993]&~m[994]&~m[996]&m[997])|(~m[952]&~m[993]&m[994]&~m[996]&m[997])|(m[952]&m[993]&m[994]&~m[996]&m[997])|(~m[952]&m[993]&m[994]&m[996]&m[997]))&UnbiasedRNG[213])|((m[952]&~m[993]&~m[994]&m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&m[994]&~m[996]&m[997])|(~m[952]&~m[993]&~m[994]&m[996]&m[997])|(m[952]&~m[993]&~m[994]&m[996]&m[997])|(~m[952]&m[993]&~m[994]&m[996]&m[997])|(m[952]&m[993]&~m[994]&m[996]&m[997])|(~m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&m[993]&m[994]&m[996]&m[997]));
    m[1000] = (((m[957]&~m[998]&~m[999]&~m[1001]&~m[1002])|(~m[957]&~m[998]&~m[999]&m[1001]&~m[1002])|(m[957]&m[998]&~m[999]&m[1001]&~m[1002])|(m[957]&~m[998]&m[999]&m[1001]&~m[1002])|(~m[957]&m[998]&~m[999]&~m[1001]&m[1002])|(~m[957]&~m[998]&m[999]&~m[1001]&m[1002])|(m[957]&m[998]&m[999]&~m[1001]&m[1002])|(~m[957]&m[998]&m[999]&m[1001]&m[1002]))&UnbiasedRNG[214])|((m[957]&~m[998]&~m[999]&m[1001]&~m[1002])|(~m[957]&~m[998]&~m[999]&~m[1001]&m[1002])|(m[957]&~m[998]&~m[999]&~m[1001]&m[1002])|(m[957]&m[998]&~m[999]&~m[1001]&m[1002])|(m[957]&~m[998]&m[999]&~m[1001]&m[1002])|(~m[957]&~m[998]&~m[999]&m[1001]&m[1002])|(m[957]&~m[998]&~m[999]&m[1001]&m[1002])|(~m[957]&m[998]&~m[999]&m[1001]&m[1002])|(m[957]&m[998]&~m[999]&m[1001]&m[1002])|(~m[957]&~m[998]&m[999]&m[1001]&m[1002])|(m[957]&~m[998]&m[999]&m[1001]&m[1002])|(m[957]&m[998]&m[999]&m[1001]&m[1002]));
    m[1005] = (((m[962]&~m[1003]&~m[1004]&~m[1006]&~m[1007])|(~m[962]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(m[962]&m[1003]&~m[1004]&m[1006]&~m[1007])|(m[962]&~m[1003]&m[1004]&m[1006]&~m[1007])|(~m[962]&m[1003]&~m[1004]&~m[1006]&m[1007])|(~m[962]&~m[1003]&m[1004]&~m[1006]&m[1007])|(m[962]&m[1003]&m[1004]&~m[1006]&m[1007])|(~m[962]&m[1003]&m[1004]&m[1006]&m[1007]))&UnbiasedRNG[215])|((m[962]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(~m[962]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[962]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[962]&m[1003]&~m[1004]&~m[1006]&m[1007])|(m[962]&~m[1003]&m[1004]&~m[1006]&m[1007])|(~m[962]&~m[1003]&~m[1004]&m[1006]&m[1007])|(m[962]&~m[1003]&~m[1004]&m[1006]&m[1007])|(~m[962]&m[1003]&~m[1004]&m[1006]&m[1007])|(m[962]&m[1003]&~m[1004]&m[1006]&m[1007])|(~m[962]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[962]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[962]&m[1003]&m[1004]&m[1006]&m[1007]));
    m[1010] = (((m[972]&~m[1008]&~m[1009]&~m[1011]&~m[1012])|(~m[972]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(m[972]&m[1008]&~m[1009]&m[1011]&~m[1012])|(m[972]&~m[1008]&m[1009]&m[1011]&~m[1012])|(~m[972]&m[1008]&~m[1009]&~m[1011]&m[1012])|(~m[972]&~m[1008]&m[1009]&~m[1011]&m[1012])|(m[972]&m[1008]&m[1009]&~m[1011]&m[1012])|(~m[972]&m[1008]&m[1009]&m[1011]&m[1012]))&UnbiasedRNG[216])|((m[972]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(~m[972]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[972]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[972]&m[1008]&~m[1009]&~m[1011]&m[1012])|(m[972]&~m[1008]&m[1009]&~m[1011]&m[1012])|(~m[972]&~m[1008]&~m[1009]&m[1011]&m[1012])|(m[972]&~m[1008]&~m[1009]&m[1011]&m[1012])|(~m[972]&m[1008]&~m[1009]&m[1011]&m[1012])|(m[972]&m[1008]&~m[1009]&m[1011]&m[1012])|(~m[972]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[972]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[972]&m[1008]&m[1009]&m[1011]&m[1012]));
    m[1015] = (((m[977]&~m[1013]&~m[1014]&~m[1016]&~m[1017])|(~m[977]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(m[977]&m[1013]&~m[1014]&m[1016]&~m[1017])|(m[977]&~m[1013]&m[1014]&m[1016]&~m[1017])|(~m[977]&m[1013]&~m[1014]&~m[1016]&m[1017])|(~m[977]&~m[1013]&m[1014]&~m[1016]&m[1017])|(m[977]&m[1013]&m[1014]&~m[1016]&m[1017])|(~m[977]&m[1013]&m[1014]&m[1016]&m[1017]))&UnbiasedRNG[217])|((m[977]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(~m[977]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[977]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[977]&m[1013]&~m[1014]&~m[1016]&m[1017])|(m[977]&~m[1013]&m[1014]&~m[1016]&m[1017])|(~m[977]&~m[1013]&~m[1014]&m[1016]&m[1017])|(m[977]&~m[1013]&~m[1014]&m[1016]&m[1017])|(~m[977]&m[1013]&~m[1014]&m[1016]&m[1017])|(m[977]&m[1013]&~m[1014]&m[1016]&m[1017])|(~m[977]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[977]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[977]&m[1013]&m[1014]&m[1016]&m[1017]));
    m[1020] = (((m[982]&~m[1018]&~m[1019]&~m[1021]&~m[1022])|(~m[982]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(m[982]&m[1018]&~m[1019]&m[1021]&~m[1022])|(m[982]&~m[1018]&m[1019]&m[1021]&~m[1022])|(~m[982]&m[1018]&~m[1019]&~m[1021]&m[1022])|(~m[982]&~m[1018]&m[1019]&~m[1021]&m[1022])|(m[982]&m[1018]&m[1019]&~m[1021]&m[1022])|(~m[982]&m[1018]&m[1019]&m[1021]&m[1022]))&UnbiasedRNG[218])|((m[982]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(~m[982]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[982]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[982]&m[1018]&~m[1019]&~m[1021]&m[1022])|(m[982]&~m[1018]&m[1019]&~m[1021]&m[1022])|(~m[982]&~m[1018]&~m[1019]&m[1021]&m[1022])|(m[982]&~m[1018]&~m[1019]&m[1021]&m[1022])|(~m[982]&m[1018]&~m[1019]&m[1021]&m[1022])|(m[982]&m[1018]&~m[1019]&m[1021]&m[1022])|(~m[982]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[982]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[982]&m[1018]&m[1019]&m[1021]&m[1022]));
    m[1025] = (((m[987]&~m[1023]&~m[1024]&~m[1026]&~m[1027])|(~m[987]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(m[987]&m[1023]&~m[1024]&m[1026]&~m[1027])|(m[987]&~m[1023]&m[1024]&m[1026]&~m[1027])|(~m[987]&m[1023]&~m[1024]&~m[1026]&m[1027])|(~m[987]&~m[1023]&m[1024]&~m[1026]&m[1027])|(m[987]&m[1023]&m[1024]&~m[1026]&m[1027])|(~m[987]&m[1023]&m[1024]&m[1026]&m[1027]))&UnbiasedRNG[219])|((m[987]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(~m[987]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[987]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[987]&m[1023]&~m[1024]&~m[1026]&m[1027])|(m[987]&~m[1023]&m[1024]&~m[1026]&m[1027])|(~m[987]&~m[1023]&~m[1024]&m[1026]&m[1027])|(m[987]&~m[1023]&~m[1024]&m[1026]&m[1027])|(~m[987]&m[1023]&~m[1024]&m[1026]&m[1027])|(m[987]&m[1023]&~m[1024]&m[1026]&m[1027])|(~m[987]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[987]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[987]&m[1023]&m[1024]&m[1026]&m[1027]));
    m[1030] = (((m[992]&~m[1028]&~m[1029]&~m[1031]&~m[1032])|(~m[992]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(m[992]&m[1028]&~m[1029]&m[1031]&~m[1032])|(m[992]&~m[1028]&m[1029]&m[1031]&~m[1032])|(~m[992]&m[1028]&~m[1029]&~m[1031]&m[1032])|(~m[992]&~m[1028]&m[1029]&~m[1031]&m[1032])|(m[992]&m[1028]&m[1029]&~m[1031]&m[1032])|(~m[992]&m[1028]&m[1029]&m[1031]&m[1032]))&UnbiasedRNG[220])|((m[992]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(~m[992]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[992]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[992]&m[1028]&~m[1029]&~m[1031]&m[1032])|(m[992]&~m[1028]&m[1029]&~m[1031]&m[1032])|(~m[992]&~m[1028]&~m[1029]&m[1031]&m[1032])|(m[992]&~m[1028]&~m[1029]&m[1031]&m[1032])|(~m[992]&m[1028]&~m[1029]&m[1031]&m[1032])|(m[992]&m[1028]&~m[1029]&m[1031]&m[1032])|(~m[992]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[992]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[992]&m[1028]&m[1029]&m[1031]&m[1032]));
    m[1035] = (((m[997]&~m[1033]&~m[1034]&~m[1036]&~m[1037])|(~m[997]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(m[997]&m[1033]&~m[1034]&m[1036]&~m[1037])|(m[997]&~m[1033]&m[1034]&m[1036]&~m[1037])|(~m[997]&m[1033]&~m[1034]&~m[1036]&m[1037])|(~m[997]&~m[1033]&m[1034]&~m[1036]&m[1037])|(m[997]&m[1033]&m[1034]&~m[1036]&m[1037])|(~m[997]&m[1033]&m[1034]&m[1036]&m[1037]))&UnbiasedRNG[221])|((m[997]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(~m[997]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[997]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[997]&m[1033]&~m[1034]&~m[1036]&m[1037])|(m[997]&~m[1033]&m[1034]&~m[1036]&m[1037])|(~m[997]&~m[1033]&~m[1034]&m[1036]&m[1037])|(m[997]&~m[1033]&~m[1034]&m[1036]&m[1037])|(~m[997]&m[1033]&~m[1034]&m[1036]&m[1037])|(m[997]&m[1033]&~m[1034]&m[1036]&m[1037])|(~m[997]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[997]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[997]&m[1033]&m[1034]&m[1036]&m[1037]));
    m[1040] = (((m[1002]&~m[1038]&~m[1039]&~m[1041]&~m[1042])|(~m[1002]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1002]&m[1038]&~m[1039]&m[1041]&~m[1042])|(m[1002]&~m[1038]&m[1039]&m[1041]&~m[1042])|(~m[1002]&m[1038]&~m[1039]&~m[1041]&m[1042])|(~m[1002]&~m[1038]&m[1039]&~m[1041]&m[1042])|(m[1002]&m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1002]&m[1038]&m[1039]&m[1041]&m[1042]))&UnbiasedRNG[222])|((m[1002]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(~m[1002]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1002]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1002]&m[1038]&~m[1039]&~m[1041]&m[1042])|(m[1002]&~m[1038]&m[1039]&~m[1041]&m[1042])|(~m[1002]&~m[1038]&~m[1039]&m[1041]&m[1042])|(m[1002]&~m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1002]&m[1038]&~m[1039]&m[1041]&m[1042])|(m[1002]&m[1038]&~m[1039]&m[1041]&m[1042])|(~m[1002]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1002]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[1002]&m[1038]&m[1039]&m[1041]&m[1042]));
    m[1045] = (((m[1007]&~m[1043]&~m[1044]&~m[1046]&~m[1047])|(~m[1007]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1007]&m[1043]&~m[1044]&m[1046]&~m[1047])|(m[1007]&~m[1043]&m[1044]&m[1046]&~m[1047])|(~m[1007]&m[1043]&~m[1044]&~m[1046]&m[1047])|(~m[1007]&~m[1043]&m[1044]&~m[1046]&m[1047])|(m[1007]&m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1007]&m[1043]&m[1044]&m[1046]&m[1047]))&UnbiasedRNG[223])|((m[1007]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(~m[1007]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1007]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1007]&m[1043]&~m[1044]&~m[1046]&m[1047])|(m[1007]&~m[1043]&m[1044]&~m[1046]&m[1047])|(~m[1007]&~m[1043]&~m[1044]&m[1046]&m[1047])|(m[1007]&~m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1007]&m[1043]&~m[1044]&m[1046]&m[1047])|(m[1007]&m[1043]&~m[1044]&m[1046]&m[1047])|(~m[1007]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1007]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[1007]&m[1043]&m[1044]&m[1046]&m[1047]));
    m[1050] = (((m[1017]&~m[1048]&~m[1049]&~m[1051]&~m[1052])|(~m[1017]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1017]&m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1017]&~m[1048]&m[1049]&m[1051]&~m[1052])|(~m[1017]&m[1048]&~m[1049]&~m[1051]&m[1052])|(~m[1017]&~m[1048]&m[1049]&~m[1051]&m[1052])|(m[1017]&m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1017]&m[1048]&m[1049]&m[1051]&m[1052]))&UnbiasedRNG[224])|((m[1017]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(~m[1017]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1017]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1017]&m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1017]&~m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1017]&~m[1048]&~m[1049]&m[1051]&m[1052])|(m[1017]&~m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1017]&m[1048]&~m[1049]&m[1051]&m[1052])|(m[1017]&m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1017]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1017]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1017]&m[1048]&m[1049]&m[1051]&m[1052]));
    m[1055] = (((m[1022]&~m[1053]&~m[1054]&~m[1056]&~m[1057])|(~m[1022]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1022]&m[1053]&~m[1054]&m[1056]&~m[1057])|(m[1022]&~m[1053]&m[1054]&m[1056]&~m[1057])|(~m[1022]&m[1053]&~m[1054]&~m[1056]&m[1057])|(~m[1022]&~m[1053]&m[1054]&~m[1056]&m[1057])|(m[1022]&m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1022]&m[1053]&m[1054]&m[1056]&m[1057]))&UnbiasedRNG[225])|((m[1022]&~m[1053]&~m[1054]&m[1056]&~m[1057])|(~m[1022]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1022]&~m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1022]&m[1053]&~m[1054]&~m[1056]&m[1057])|(m[1022]&~m[1053]&m[1054]&~m[1056]&m[1057])|(~m[1022]&~m[1053]&~m[1054]&m[1056]&m[1057])|(m[1022]&~m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1022]&m[1053]&~m[1054]&m[1056]&m[1057])|(m[1022]&m[1053]&~m[1054]&m[1056]&m[1057])|(~m[1022]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1022]&~m[1053]&m[1054]&m[1056]&m[1057])|(m[1022]&m[1053]&m[1054]&m[1056]&m[1057]));
    m[1060] = (((m[1027]&~m[1058]&~m[1059]&~m[1061]&~m[1062])|(~m[1027]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1027]&m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1027]&~m[1058]&m[1059]&m[1061]&~m[1062])|(~m[1027]&m[1058]&~m[1059]&~m[1061]&m[1062])|(~m[1027]&~m[1058]&m[1059]&~m[1061]&m[1062])|(m[1027]&m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1027]&m[1058]&m[1059]&m[1061]&m[1062]))&UnbiasedRNG[226])|((m[1027]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(~m[1027]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1027]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1027]&m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1027]&~m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1027]&~m[1058]&~m[1059]&m[1061]&m[1062])|(m[1027]&~m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1027]&m[1058]&~m[1059]&m[1061]&m[1062])|(m[1027]&m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1027]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1027]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1027]&m[1058]&m[1059]&m[1061]&m[1062]));
    m[1065] = (((m[1032]&~m[1063]&~m[1064]&~m[1066]&~m[1067])|(~m[1032]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1032]&m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1032]&~m[1063]&m[1064]&m[1066]&~m[1067])|(~m[1032]&m[1063]&~m[1064]&~m[1066]&m[1067])|(~m[1032]&~m[1063]&m[1064]&~m[1066]&m[1067])|(m[1032]&m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1032]&m[1063]&m[1064]&m[1066]&m[1067]))&UnbiasedRNG[227])|((m[1032]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(~m[1032]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1032]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1032]&m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1032]&~m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1032]&~m[1063]&~m[1064]&m[1066]&m[1067])|(m[1032]&~m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1032]&m[1063]&~m[1064]&m[1066]&m[1067])|(m[1032]&m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1032]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1032]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1032]&m[1063]&m[1064]&m[1066]&m[1067]));
    m[1070] = (((m[1037]&~m[1068]&~m[1069]&~m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&~m[1072])|(~m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&m[1068]&m[1069]&m[1071]&m[1072]))&UnbiasedRNG[228])|((m[1037]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(~m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1037]&m[1068]&m[1069]&m[1071]&m[1072]));
    m[1075] = (((m[1042]&~m[1073]&~m[1074]&~m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&~m[1077])|(~m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&m[1073]&m[1074]&m[1076]&m[1077]))&UnbiasedRNG[229])|((m[1042]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(~m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1042]&m[1073]&m[1074]&m[1076]&m[1077]));
    m[1080] = (((m[1047]&~m[1078]&~m[1079]&~m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&~m[1082])|(~m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&m[1078]&m[1079]&m[1081]&m[1082]))&UnbiasedRNG[230])|((m[1047]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(~m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1047]&m[1078]&m[1079]&m[1081]&m[1082]));
    m[1085] = (((m[1057]&~m[1083]&~m[1084]&~m[1086]&~m[1087])|(~m[1057]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1057]&m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1057]&~m[1083]&m[1084]&m[1086]&~m[1087])|(~m[1057]&m[1083]&~m[1084]&~m[1086]&m[1087])|(~m[1057]&~m[1083]&m[1084]&~m[1086]&m[1087])|(m[1057]&m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1057]&m[1083]&m[1084]&m[1086]&m[1087]))&UnbiasedRNG[231])|((m[1057]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(~m[1057]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1057]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1057]&m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1057]&~m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1057]&~m[1083]&~m[1084]&m[1086]&m[1087])|(m[1057]&~m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1057]&m[1083]&~m[1084]&m[1086]&m[1087])|(m[1057]&m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1057]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1057]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1057]&m[1083]&m[1084]&m[1086]&m[1087]));
    m[1090] = (((m[1062]&~m[1088]&~m[1089]&~m[1091]&~m[1092])|(~m[1062]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1062]&m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1062]&~m[1088]&m[1089]&m[1091]&~m[1092])|(~m[1062]&m[1088]&~m[1089]&~m[1091]&m[1092])|(~m[1062]&~m[1088]&m[1089]&~m[1091]&m[1092])|(m[1062]&m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1062]&m[1088]&m[1089]&m[1091]&m[1092]))&UnbiasedRNG[232])|((m[1062]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(~m[1062]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1062]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1062]&m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1062]&~m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1062]&~m[1088]&~m[1089]&m[1091]&m[1092])|(m[1062]&~m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1062]&m[1088]&~m[1089]&m[1091]&m[1092])|(m[1062]&m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1062]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1062]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1062]&m[1088]&m[1089]&m[1091]&m[1092]));
    m[1095] = (((m[1067]&~m[1093]&~m[1094]&~m[1096]&~m[1097])|(~m[1067]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1067]&m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1067]&~m[1093]&m[1094]&m[1096]&~m[1097])|(~m[1067]&m[1093]&~m[1094]&~m[1096]&m[1097])|(~m[1067]&~m[1093]&m[1094]&~m[1096]&m[1097])|(m[1067]&m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1067]&m[1093]&m[1094]&m[1096]&m[1097]))&UnbiasedRNG[233])|((m[1067]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(~m[1067]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1067]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1067]&m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1067]&~m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1067]&~m[1093]&~m[1094]&m[1096]&m[1097])|(m[1067]&~m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1067]&m[1093]&~m[1094]&m[1096]&m[1097])|(m[1067]&m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1067]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1067]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1067]&m[1093]&m[1094]&m[1096]&m[1097]));
    m[1100] = (((m[1072]&~m[1098]&~m[1099]&~m[1101]&~m[1102])|(~m[1072]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1072]&m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1072]&~m[1098]&m[1099]&m[1101]&~m[1102])|(~m[1072]&m[1098]&~m[1099]&~m[1101]&m[1102])|(~m[1072]&~m[1098]&m[1099]&~m[1101]&m[1102])|(m[1072]&m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1072]&m[1098]&m[1099]&m[1101]&m[1102]))&UnbiasedRNG[234])|((m[1072]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(~m[1072]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1072]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1072]&m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1072]&~m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1072]&~m[1098]&~m[1099]&m[1101]&m[1102])|(m[1072]&~m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1072]&m[1098]&~m[1099]&m[1101]&m[1102])|(m[1072]&m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1072]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1072]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1072]&m[1098]&m[1099]&m[1101]&m[1102]));
    m[1105] = (((m[1077]&~m[1103]&~m[1104]&~m[1106]&~m[1107])|(~m[1077]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1077]&m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1077]&~m[1103]&m[1104]&m[1106]&~m[1107])|(~m[1077]&m[1103]&~m[1104]&~m[1106]&m[1107])|(~m[1077]&~m[1103]&m[1104]&~m[1106]&m[1107])|(m[1077]&m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1077]&m[1103]&m[1104]&m[1106]&m[1107]))&UnbiasedRNG[235])|((m[1077]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(~m[1077]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1077]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1077]&m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1077]&~m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1077]&~m[1103]&~m[1104]&m[1106]&m[1107])|(m[1077]&~m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1077]&m[1103]&~m[1104]&m[1106]&m[1107])|(m[1077]&m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1077]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1077]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1077]&m[1103]&m[1104]&m[1106]&m[1107]));
    m[1110] = (((m[1082]&~m[1108]&~m[1109]&~m[1111]&~m[1112])|(~m[1082]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1082]&m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1082]&~m[1108]&m[1109]&m[1111]&~m[1112])|(~m[1082]&m[1108]&~m[1109]&~m[1111]&m[1112])|(~m[1082]&~m[1108]&m[1109]&~m[1111]&m[1112])|(m[1082]&m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1082]&m[1108]&m[1109]&m[1111]&m[1112]))&UnbiasedRNG[236])|((m[1082]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(~m[1082]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1082]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1082]&m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1082]&~m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1082]&~m[1108]&~m[1109]&m[1111]&m[1112])|(m[1082]&~m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1082]&m[1108]&~m[1109]&m[1111]&m[1112])|(m[1082]&m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1082]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1082]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1082]&m[1108]&m[1109]&m[1111]&m[1112]));
    m[1115] = (((m[1092]&~m[1113]&~m[1114]&~m[1116]&~m[1117])|(~m[1092]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1092]&m[1113]&~m[1114]&m[1116]&~m[1117])|(m[1092]&~m[1113]&m[1114]&m[1116]&~m[1117])|(~m[1092]&m[1113]&~m[1114]&~m[1116]&m[1117])|(~m[1092]&~m[1113]&m[1114]&~m[1116]&m[1117])|(m[1092]&m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1092]&m[1113]&m[1114]&m[1116]&m[1117]))&UnbiasedRNG[237])|((m[1092]&~m[1113]&~m[1114]&m[1116]&~m[1117])|(~m[1092]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1092]&~m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1092]&m[1113]&~m[1114]&~m[1116]&m[1117])|(m[1092]&~m[1113]&m[1114]&~m[1116]&m[1117])|(~m[1092]&~m[1113]&~m[1114]&m[1116]&m[1117])|(m[1092]&~m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1092]&m[1113]&~m[1114]&m[1116]&m[1117])|(m[1092]&m[1113]&~m[1114]&m[1116]&m[1117])|(~m[1092]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1092]&~m[1113]&m[1114]&m[1116]&m[1117])|(m[1092]&m[1113]&m[1114]&m[1116]&m[1117]));
    m[1120] = (((m[1097]&~m[1118]&~m[1119]&~m[1121]&~m[1122])|(~m[1097]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1097]&m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1097]&~m[1118]&m[1119]&m[1121]&~m[1122])|(~m[1097]&m[1118]&~m[1119]&~m[1121]&m[1122])|(~m[1097]&~m[1118]&m[1119]&~m[1121]&m[1122])|(m[1097]&m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1097]&m[1118]&m[1119]&m[1121]&m[1122]))&UnbiasedRNG[238])|((m[1097]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(~m[1097]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1097]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1097]&m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1097]&~m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1097]&~m[1118]&~m[1119]&m[1121]&m[1122])|(m[1097]&~m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1097]&m[1118]&~m[1119]&m[1121]&m[1122])|(m[1097]&m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1097]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1097]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1097]&m[1118]&m[1119]&m[1121]&m[1122]));
    m[1125] = (((m[1102]&~m[1123]&~m[1124]&~m[1126]&~m[1127])|(~m[1102]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1102]&m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1102]&~m[1123]&m[1124]&m[1126]&~m[1127])|(~m[1102]&m[1123]&~m[1124]&~m[1126]&m[1127])|(~m[1102]&~m[1123]&m[1124]&~m[1126]&m[1127])|(m[1102]&m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1102]&m[1123]&m[1124]&m[1126]&m[1127]))&UnbiasedRNG[239])|((m[1102]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(~m[1102]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1102]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1102]&m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1102]&~m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1102]&~m[1123]&~m[1124]&m[1126]&m[1127])|(m[1102]&~m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1102]&m[1123]&~m[1124]&m[1126]&m[1127])|(m[1102]&m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1102]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1102]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1102]&m[1123]&m[1124]&m[1126]&m[1127]));
    m[1130] = (((m[1107]&~m[1128]&~m[1129]&~m[1131]&~m[1132])|(~m[1107]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1107]&m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1107]&~m[1128]&m[1129]&m[1131]&~m[1132])|(~m[1107]&m[1128]&~m[1129]&~m[1131]&m[1132])|(~m[1107]&~m[1128]&m[1129]&~m[1131]&m[1132])|(m[1107]&m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1107]&m[1128]&m[1129]&m[1131]&m[1132]))&UnbiasedRNG[240])|((m[1107]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(~m[1107]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1107]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1107]&m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1107]&~m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1107]&~m[1128]&~m[1129]&m[1131]&m[1132])|(m[1107]&~m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1107]&m[1128]&~m[1129]&m[1131]&m[1132])|(m[1107]&m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1107]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1107]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1107]&m[1128]&m[1129]&m[1131]&m[1132]));
    m[1135] = (((m[1112]&~m[1133]&~m[1134]&~m[1136]&~m[1137])|(~m[1112]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1112]&m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1112]&~m[1133]&m[1134]&m[1136]&~m[1137])|(~m[1112]&m[1133]&~m[1134]&~m[1136]&m[1137])|(~m[1112]&~m[1133]&m[1134]&~m[1136]&m[1137])|(m[1112]&m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1112]&m[1133]&m[1134]&m[1136]&m[1137]))&UnbiasedRNG[241])|((m[1112]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(~m[1112]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1112]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1112]&m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1112]&~m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1112]&~m[1133]&~m[1134]&m[1136]&m[1137])|(m[1112]&~m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1112]&m[1133]&~m[1134]&m[1136]&m[1137])|(m[1112]&m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1112]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1112]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1112]&m[1133]&m[1134]&m[1136]&m[1137]));
    m[1140] = (((m[1122]&~m[1138]&~m[1139]&~m[1141]&~m[1142])|(~m[1122]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1122]&m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1122]&~m[1138]&m[1139]&m[1141]&~m[1142])|(~m[1122]&m[1138]&~m[1139]&~m[1141]&m[1142])|(~m[1122]&~m[1138]&m[1139]&~m[1141]&m[1142])|(m[1122]&m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1122]&m[1138]&m[1139]&m[1141]&m[1142]))&UnbiasedRNG[242])|((m[1122]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(~m[1122]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1122]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1122]&m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1122]&~m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1122]&~m[1138]&~m[1139]&m[1141]&m[1142])|(m[1122]&~m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1122]&m[1138]&~m[1139]&m[1141]&m[1142])|(m[1122]&m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1122]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1122]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1122]&m[1138]&m[1139]&m[1141]&m[1142]));
    m[1145] = (((m[1127]&~m[1143]&~m[1144]&~m[1146]&~m[1147])|(~m[1127]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1127]&m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1127]&~m[1143]&m[1144]&m[1146]&~m[1147])|(~m[1127]&m[1143]&~m[1144]&~m[1146]&m[1147])|(~m[1127]&~m[1143]&m[1144]&~m[1146]&m[1147])|(m[1127]&m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1127]&m[1143]&m[1144]&m[1146]&m[1147]))&UnbiasedRNG[243])|((m[1127]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(~m[1127]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1127]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1127]&m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1127]&~m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1127]&~m[1143]&~m[1144]&m[1146]&m[1147])|(m[1127]&~m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1127]&m[1143]&~m[1144]&m[1146]&m[1147])|(m[1127]&m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1127]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1127]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1127]&m[1143]&m[1144]&m[1146]&m[1147]));
    m[1150] = (((m[1132]&~m[1148]&~m[1149]&~m[1151]&~m[1152])|(~m[1132]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1132]&m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1132]&~m[1148]&m[1149]&m[1151]&~m[1152])|(~m[1132]&m[1148]&~m[1149]&~m[1151]&m[1152])|(~m[1132]&~m[1148]&m[1149]&~m[1151]&m[1152])|(m[1132]&m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1132]&m[1148]&m[1149]&m[1151]&m[1152]))&UnbiasedRNG[244])|((m[1132]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(~m[1132]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1132]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1132]&m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1132]&~m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1132]&~m[1148]&~m[1149]&m[1151]&m[1152])|(m[1132]&~m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1132]&m[1148]&~m[1149]&m[1151]&m[1152])|(m[1132]&m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1132]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1132]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1132]&m[1148]&m[1149]&m[1151]&m[1152]));
    m[1155] = (((m[1137]&~m[1153]&~m[1154]&~m[1156]&~m[1157])|(~m[1137]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1137]&m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1137]&~m[1153]&m[1154]&m[1156]&~m[1157])|(~m[1137]&m[1153]&~m[1154]&~m[1156]&m[1157])|(~m[1137]&~m[1153]&m[1154]&~m[1156]&m[1157])|(m[1137]&m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1137]&m[1153]&m[1154]&m[1156]&m[1157]))&UnbiasedRNG[245])|((m[1137]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(~m[1137]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1137]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1137]&m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1137]&~m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1137]&~m[1153]&~m[1154]&m[1156]&m[1157])|(m[1137]&~m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1137]&m[1153]&~m[1154]&m[1156]&m[1157])|(m[1137]&m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1137]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1137]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1137]&m[1153]&m[1154]&m[1156]&m[1157]));
    m[1160] = (((m[1147]&~m[1158]&~m[1159]&~m[1161]&~m[1162])|(~m[1147]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1147]&m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1147]&~m[1158]&m[1159]&m[1161]&~m[1162])|(~m[1147]&m[1158]&~m[1159]&~m[1161]&m[1162])|(~m[1147]&~m[1158]&m[1159]&~m[1161]&m[1162])|(m[1147]&m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1147]&m[1158]&m[1159]&m[1161]&m[1162]))&UnbiasedRNG[246])|((m[1147]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(~m[1147]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1147]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1147]&m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1147]&~m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1147]&~m[1158]&~m[1159]&m[1161]&m[1162])|(m[1147]&~m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1147]&m[1158]&~m[1159]&m[1161]&m[1162])|(m[1147]&m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1147]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1147]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1147]&m[1158]&m[1159]&m[1161]&m[1162]));
    m[1165] = (((m[1152]&~m[1163]&~m[1164]&~m[1166]&~m[1167])|(~m[1152]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1152]&m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1152]&~m[1163]&m[1164]&m[1166]&~m[1167])|(~m[1152]&m[1163]&~m[1164]&~m[1166]&m[1167])|(~m[1152]&~m[1163]&m[1164]&~m[1166]&m[1167])|(m[1152]&m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1152]&m[1163]&m[1164]&m[1166]&m[1167]))&UnbiasedRNG[247])|((m[1152]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(~m[1152]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1152]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1152]&m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1152]&~m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1152]&~m[1163]&~m[1164]&m[1166]&m[1167])|(m[1152]&~m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1152]&m[1163]&~m[1164]&m[1166]&m[1167])|(m[1152]&m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1152]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1152]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1152]&m[1163]&m[1164]&m[1166]&m[1167]));
    m[1170] = (((m[1157]&~m[1168]&~m[1169]&~m[1171]&~m[1172])|(~m[1157]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1157]&m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1157]&~m[1168]&m[1169]&m[1171]&~m[1172])|(~m[1157]&m[1168]&~m[1169]&~m[1171]&m[1172])|(~m[1157]&~m[1168]&m[1169]&~m[1171]&m[1172])|(m[1157]&m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1157]&m[1168]&m[1169]&m[1171]&m[1172]))&UnbiasedRNG[248])|((m[1157]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(~m[1157]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1157]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1157]&m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1157]&~m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1157]&~m[1168]&~m[1169]&m[1171]&m[1172])|(m[1157]&~m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1157]&m[1168]&~m[1169]&m[1171]&m[1172])|(m[1157]&m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1157]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1157]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1157]&m[1168]&m[1169]&m[1171]&m[1172]));
    m[1175] = (((m[1167]&~m[1173]&~m[1174]&~m[1176]&~m[1177])|(~m[1167]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1167]&m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1167]&~m[1173]&m[1174]&m[1176]&~m[1177])|(~m[1167]&m[1173]&~m[1174]&~m[1176]&m[1177])|(~m[1167]&~m[1173]&m[1174]&~m[1176]&m[1177])|(m[1167]&m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1167]&m[1173]&m[1174]&m[1176]&m[1177]))&UnbiasedRNG[249])|((m[1167]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(~m[1167]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1167]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1167]&m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1167]&~m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1167]&~m[1173]&~m[1174]&m[1176]&m[1177])|(m[1167]&~m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1167]&m[1173]&~m[1174]&m[1176]&m[1177])|(m[1167]&m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1167]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1167]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1167]&m[1173]&m[1174]&m[1176]&m[1177]));
    m[1180] = (((m[1172]&~m[1178]&~m[1179]&~m[1181]&~m[1182])|(~m[1172]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1172]&m[1178]&~m[1179]&m[1181]&~m[1182])|(m[1172]&~m[1178]&m[1179]&m[1181]&~m[1182])|(~m[1172]&m[1178]&~m[1179]&~m[1181]&m[1182])|(~m[1172]&~m[1178]&m[1179]&~m[1181]&m[1182])|(m[1172]&m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1172]&m[1178]&m[1179]&m[1181]&m[1182]))&UnbiasedRNG[250])|((m[1172]&~m[1178]&~m[1179]&m[1181]&~m[1182])|(~m[1172]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1172]&~m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1172]&m[1178]&~m[1179]&~m[1181]&m[1182])|(m[1172]&~m[1178]&m[1179]&~m[1181]&m[1182])|(~m[1172]&~m[1178]&~m[1179]&m[1181]&m[1182])|(m[1172]&~m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1172]&m[1178]&~m[1179]&m[1181]&m[1182])|(m[1172]&m[1178]&~m[1179]&m[1181]&m[1182])|(~m[1172]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1172]&~m[1178]&m[1179]&m[1181]&m[1182])|(m[1172]&m[1178]&m[1179]&m[1181]&m[1182]));
    m[1185] = (((m[1182]&~m[1183]&~m[1184]&~m[1186]&~m[1187])|(~m[1182]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1182]&m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1182]&~m[1183]&m[1184]&m[1186]&~m[1187])|(~m[1182]&m[1183]&~m[1184]&~m[1186]&m[1187])|(~m[1182]&~m[1183]&m[1184]&~m[1186]&m[1187])|(m[1182]&m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1182]&m[1183]&m[1184]&m[1186]&m[1187]))&UnbiasedRNG[251])|((m[1182]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(~m[1182]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1182]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1182]&m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1182]&~m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1182]&~m[1183]&~m[1184]&m[1186]&m[1187])|(m[1182]&~m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1182]&m[1183]&~m[1184]&m[1186]&m[1187])|(m[1182]&m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1182]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1182]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1182]&m[1183]&m[1184]&m[1186]&m[1187]));
end

always @(posedge color2_clk) begin
    m[240] = (((~m[60]&~m[96]&~m[384])|(m[60]&m[96]&~m[384]))&BiasedRNG[383])|(((m[60]&~m[96]&~m[384])|(~m[60]&m[96]&m[384]))&~BiasedRNG[383])|((~m[60]&~m[96]&m[384])|(m[60]&~m[96]&m[384])|(m[60]&m[96]&m[384]));
    m[241] = (((~m[60]&~m[108]&~m[385])|(m[60]&m[108]&~m[385]))&BiasedRNG[384])|(((m[60]&~m[108]&~m[385])|(~m[60]&m[108]&m[385]))&~BiasedRNG[384])|((~m[60]&~m[108]&m[385])|(m[60]&~m[108]&m[385])|(m[60]&m[108]&m[385]));
    m[242] = (((~m[60]&~m[120]&~m[386])|(m[60]&m[120]&~m[386]))&BiasedRNG[385])|(((m[60]&~m[120]&~m[386])|(~m[60]&m[120]&m[386]))&~BiasedRNG[385])|((~m[60]&~m[120]&m[386])|(m[60]&~m[120]&m[386])|(m[60]&m[120]&m[386]));
    m[243] = (((~m[60]&~m[132]&~m[387])|(m[60]&m[132]&~m[387]))&BiasedRNG[386])|(((m[60]&~m[132]&~m[387])|(~m[60]&m[132]&m[387]))&~BiasedRNG[386])|((~m[60]&~m[132]&m[387])|(m[60]&~m[132]&m[387])|(m[60]&m[132]&m[387]));
    m[244] = (((~m[61]&~m[144]&~m[388])|(m[61]&m[144]&~m[388]))&BiasedRNG[387])|(((m[61]&~m[144]&~m[388])|(~m[61]&m[144]&m[388]))&~BiasedRNG[387])|((~m[61]&~m[144]&m[388])|(m[61]&~m[144]&m[388])|(m[61]&m[144]&m[388]));
    m[245] = (((~m[61]&~m[156]&~m[389])|(m[61]&m[156]&~m[389]))&BiasedRNG[388])|(((m[61]&~m[156]&~m[389])|(~m[61]&m[156]&m[389]))&~BiasedRNG[388])|((~m[61]&~m[156]&m[389])|(m[61]&~m[156]&m[389])|(m[61]&m[156]&m[389]));
    m[246] = (((~m[61]&~m[168]&~m[390])|(m[61]&m[168]&~m[390]))&BiasedRNG[389])|(((m[61]&~m[168]&~m[390])|(~m[61]&m[168]&m[390]))&~BiasedRNG[389])|((~m[61]&~m[168]&m[390])|(m[61]&~m[168]&m[390])|(m[61]&m[168]&m[390]));
    m[247] = (((~m[61]&~m[180]&~m[391])|(m[61]&m[180]&~m[391]))&BiasedRNG[390])|(((m[61]&~m[180]&~m[391])|(~m[61]&m[180]&m[391]))&~BiasedRNG[390])|((~m[61]&~m[180]&m[391])|(m[61]&~m[180]&m[391])|(m[61]&m[180]&m[391]));
    m[248] = (((~m[62]&~m[192]&~m[392])|(m[62]&m[192]&~m[392]))&BiasedRNG[391])|(((m[62]&~m[192]&~m[392])|(~m[62]&m[192]&m[392]))&~BiasedRNG[391])|((~m[62]&~m[192]&m[392])|(m[62]&~m[192]&m[392])|(m[62]&m[192]&m[392]));
    m[249] = (((~m[62]&~m[204]&~m[393])|(m[62]&m[204]&~m[393]))&BiasedRNG[392])|(((m[62]&~m[204]&~m[393])|(~m[62]&m[204]&m[393]))&~BiasedRNG[392])|((~m[62]&~m[204]&m[393])|(m[62]&~m[204]&m[393])|(m[62]&m[204]&m[393]));
    m[250] = (((~m[62]&~m[216]&~m[394])|(m[62]&m[216]&~m[394]))&BiasedRNG[393])|(((m[62]&~m[216]&~m[394])|(~m[62]&m[216]&m[394]))&~BiasedRNG[393])|((~m[62]&~m[216]&m[394])|(m[62]&~m[216]&m[394])|(m[62]&m[216]&m[394]));
    m[251] = (((~m[62]&~m[228]&~m[395])|(m[62]&m[228]&~m[395]))&BiasedRNG[394])|(((m[62]&~m[228]&~m[395])|(~m[62]&m[228]&m[395]))&~BiasedRNG[394])|((~m[62]&~m[228]&m[395])|(m[62]&~m[228]&m[395])|(m[62]&m[228]&m[395]));
    m[252] = (((~m[63]&~m[97]&~m[396])|(m[63]&m[97]&~m[396]))&BiasedRNG[395])|(((m[63]&~m[97]&~m[396])|(~m[63]&m[97]&m[396]))&~BiasedRNG[395])|((~m[63]&~m[97]&m[396])|(m[63]&~m[97]&m[396])|(m[63]&m[97]&m[396]));
    m[253] = (((~m[63]&~m[109]&~m[397])|(m[63]&m[109]&~m[397]))&BiasedRNG[396])|(((m[63]&~m[109]&~m[397])|(~m[63]&m[109]&m[397]))&~BiasedRNG[396])|((~m[63]&~m[109]&m[397])|(m[63]&~m[109]&m[397])|(m[63]&m[109]&m[397]));
    m[254] = (((~m[63]&~m[121]&~m[398])|(m[63]&m[121]&~m[398]))&BiasedRNG[397])|(((m[63]&~m[121]&~m[398])|(~m[63]&m[121]&m[398]))&~BiasedRNG[397])|((~m[63]&~m[121]&m[398])|(m[63]&~m[121]&m[398])|(m[63]&m[121]&m[398]));
    m[255] = (((~m[63]&~m[133]&~m[399])|(m[63]&m[133]&~m[399]))&BiasedRNG[398])|(((m[63]&~m[133]&~m[399])|(~m[63]&m[133]&m[399]))&~BiasedRNG[398])|((~m[63]&~m[133]&m[399])|(m[63]&~m[133]&m[399])|(m[63]&m[133]&m[399]));
    m[256] = (((~m[64]&~m[145]&~m[400])|(m[64]&m[145]&~m[400]))&BiasedRNG[399])|(((m[64]&~m[145]&~m[400])|(~m[64]&m[145]&m[400]))&~BiasedRNG[399])|((~m[64]&~m[145]&m[400])|(m[64]&~m[145]&m[400])|(m[64]&m[145]&m[400]));
    m[257] = (((~m[64]&~m[157]&~m[401])|(m[64]&m[157]&~m[401]))&BiasedRNG[400])|(((m[64]&~m[157]&~m[401])|(~m[64]&m[157]&m[401]))&~BiasedRNG[400])|((~m[64]&~m[157]&m[401])|(m[64]&~m[157]&m[401])|(m[64]&m[157]&m[401]));
    m[258] = (((~m[64]&~m[169]&~m[402])|(m[64]&m[169]&~m[402]))&BiasedRNG[401])|(((m[64]&~m[169]&~m[402])|(~m[64]&m[169]&m[402]))&~BiasedRNG[401])|((~m[64]&~m[169]&m[402])|(m[64]&~m[169]&m[402])|(m[64]&m[169]&m[402]));
    m[259] = (((~m[64]&~m[181]&~m[403])|(m[64]&m[181]&~m[403]))&BiasedRNG[402])|(((m[64]&~m[181]&~m[403])|(~m[64]&m[181]&m[403]))&~BiasedRNG[402])|((~m[64]&~m[181]&m[403])|(m[64]&~m[181]&m[403])|(m[64]&m[181]&m[403]));
    m[260] = (((~m[65]&~m[193]&~m[404])|(m[65]&m[193]&~m[404]))&BiasedRNG[403])|(((m[65]&~m[193]&~m[404])|(~m[65]&m[193]&m[404]))&~BiasedRNG[403])|((~m[65]&~m[193]&m[404])|(m[65]&~m[193]&m[404])|(m[65]&m[193]&m[404]));
    m[261] = (((~m[65]&~m[205]&~m[405])|(m[65]&m[205]&~m[405]))&BiasedRNG[404])|(((m[65]&~m[205]&~m[405])|(~m[65]&m[205]&m[405]))&~BiasedRNG[404])|((~m[65]&~m[205]&m[405])|(m[65]&~m[205]&m[405])|(m[65]&m[205]&m[405]));
    m[262] = (((~m[65]&~m[217]&~m[406])|(m[65]&m[217]&~m[406]))&BiasedRNG[405])|(((m[65]&~m[217]&~m[406])|(~m[65]&m[217]&m[406]))&~BiasedRNG[405])|((~m[65]&~m[217]&m[406])|(m[65]&~m[217]&m[406])|(m[65]&m[217]&m[406]));
    m[263] = (((~m[65]&~m[229]&~m[407])|(m[65]&m[229]&~m[407]))&BiasedRNG[406])|(((m[65]&~m[229]&~m[407])|(~m[65]&m[229]&m[407]))&~BiasedRNG[406])|((~m[65]&~m[229]&m[407])|(m[65]&~m[229]&m[407])|(m[65]&m[229]&m[407]));
    m[264] = (((~m[66]&~m[98]&~m[408])|(m[66]&m[98]&~m[408]))&BiasedRNG[407])|(((m[66]&~m[98]&~m[408])|(~m[66]&m[98]&m[408]))&~BiasedRNG[407])|((~m[66]&~m[98]&m[408])|(m[66]&~m[98]&m[408])|(m[66]&m[98]&m[408]));
    m[265] = (((~m[66]&~m[110]&~m[409])|(m[66]&m[110]&~m[409]))&BiasedRNG[408])|(((m[66]&~m[110]&~m[409])|(~m[66]&m[110]&m[409]))&~BiasedRNG[408])|((~m[66]&~m[110]&m[409])|(m[66]&~m[110]&m[409])|(m[66]&m[110]&m[409]));
    m[266] = (((~m[66]&~m[122]&~m[410])|(m[66]&m[122]&~m[410]))&BiasedRNG[409])|(((m[66]&~m[122]&~m[410])|(~m[66]&m[122]&m[410]))&~BiasedRNG[409])|((~m[66]&~m[122]&m[410])|(m[66]&~m[122]&m[410])|(m[66]&m[122]&m[410]));
    m[267] = (((~m[66]&~m[134]&~m[411])|(m[66]&m[134]&~m[411]))&BiasedRNG[410])|(((m[66]&~m[134]&~m[411])|(~m[66]&m[134]&m[411]))&~BiasedRNG[410])|((~m[66]&~m[134]&m[411])|(m[66]&~m[134]&m[411])|(m[66]&m[134]&m[411]));
    m[268] = (((~m[67]&~m[146]&~m[412])|(m[67]&m[146]&~m[412]))&BiasedRNG[411])|(((m[67]&~m[146]&~m[412])|(~m[67]&m[146]&m[412]))&~BiasedRNG[411])|((~m[67]&~m[146]&m[412])|(m[67]&~m[146]&m[412])|(m[67]&m[146]&m[412]));
    m[269] = (((~m[67]&~m[158]&~m[413])|(m[67]&m[158]&~m[413]))&BiasedRNG[412])|(((m[67]&~m[158]&~m[413])|(~m[67]&m[158]&m[413]))&~BiasedRNG[412])|((~m[67]&~m[158]&m[413])|(m[67]&~m[158]&m[413])|(m[67]&m[158]&m[413]));
    m[270] = (((~m[67]&~m[170]&~m[414])|(m[67]&m[170]&~m[414]))&BiasedRNG[413])|(((m[67]&~m[170]&~m[414])|(~m[67]&m[170]&m[414]))&~BiasedRNG[413])|((~m[67]&~m[170]&m[414])|(m[67]&~m[170]&m[414])|(m[67]&m[170]&m[414]));
    m[271] = (((~m[67]&~m[182]&~m[415])|(m[67]&m[182]&~m[415]))&BiasedRNG[414])|(((m[67]&~m[182]&~m[415])|(~m[67]&m[182]&m[415]))&~BiasedRNG[414])|((~m[67]&~m[182]&m[415])|(m[67]&~m[182]&m[415])|(m[67]&m[182]&m[415]));
    m[272] = (((~m[68]&~m[194]&~m[416])|(m[68]&m[194]&~m[416]))&BiasedRNG[415])|(((m[68]&~m[194]&~m[416])|(~m[68]&m[194]&m[416]))&~BiasedRNG[415])|((~m[68]&~m[194]&m[416])|(m[68]&~m[194]&m[416])|(m[68]&m[194]&m[416]));
    m[273] = (((~m[68]&~m[206]&~m[417])|(m[68]&m[206]&~m[417]))&BiasedRNG[416])|(((m[68]&~m[206]&~m[417])|(~m[68]&m[206]&m[417]))&~BiasedRNG[416])|((~m[68]&~m[206]&m[417])|(m[68]&~m[206]&m[417])|(m[68]&m[206]&m[417]));
    m[274] = (((~m[68]&~m[218]&~m[418])|(m[68]&m[218]&~m[418]))&BiasedRNG[417])|(((m[68]&~m[218]&~m[418])|(~m[68]&m[218]&m[418]))&~BiasedRNG[417])|((~m[68]&~m[218]&m[418])|(m[68]&~m[218]&m[418])|(m[68]&m[218]&m[418]));
    m[275] = (((~m[68]&~m[230]&~m[419])|(m[68]&m[230]&~m[419]))&BiasedRNG[418])|(((m[68]&~m[230]&~m[419])|(~m[68]&m[230]&m[419]))&~BiasedRNG[418])|((~m[68]&~m[230]&m[419])|(m[68]&~m[230]&m[419])|(m[68]&m[230]&m[419]));
    m[276] = (((~m[69]&~m[99]&~m[420])|(m[69]&m[99]&~m[420]))&BiasedRNG[419])|(((m[69]&~m[99]&~m[420])|(~m[69]&m[99]&m[420]))&~BiasedRNG[419])|((~m[69]&~m[99]&m[420])|(m[69]&~m[99]&m[420])|(m[69]&m[99]&m[420]));
    m[277] = (((~m[69]&~m[111]&~m[421])|(m[69]&m[111]&~m[421]))&BiasedRNG[420])|(((m[69]&~m[111]&~m[421])|(~m[69]&m[111]&m[421]))&~BiasedRNG[420])|((~m[69]&~m[111]&m[421])|(m[69]&~m[111]&m[421])|(m[69]&m[111]&m[421]));
    m[278] = (((~m[69]&~m[123]&~m[422])|(m[69]&m[123]&~m[422]))&BiasedRNG[421])|(((m[69]&~m[123]&~m[422])|(~m[69]&m[123]&m[422]))&~BiasedRNG[421])|((~m[69]&~m[123]&m[422])|(m[69]&~m[123]&m[422])|(m[69]&m[123]&m[422]));
    m[279] = (((~m[69]&~m[135]&~m[423])|(m[69]&m[135]&~m[423]))&BiasedRNG[422])|(((m[69]&~m[135]&~m[423])|(~m[69]&m[135]&m[423]))&~BiasedRNG[422])|((~m[69]&~m[135]&m[423])|(m[69]&~m[135]&m[423])|(m[69]&m[135]&m[423]));
    m[280] = (((~m[70]&~m[147]&~m[424])|(m[70]&m[147]&~m[424]))&BiasedRNG[423])|(((m[70]&~m[147]&~m[424])|(~m[70]&m[147]&m[424]))&~BiasedRNG[423])|((~m[70]&~m[147]&m[424])|(m[70]&~m[147]&m[424])|(m[70]&m[147]&m[424]));
    m[281] = (((~m[70]&~m[159]&~m[425])|(m[70]&m[159]&~m[425]))&BiasedRNG[424])|(((m[70]&~m[159]&~m[425])|(~m[70]&m[159]&m[425]))&~BiasedRNG[424])|((~m[70]&~m[159]&m[425])|(m[70]&~m[159]&m[425])|(m[70]&m[159]&m[425]));
    m[282] = (((~m[70]&~m[171]&~m[426])|(m[70]&m[171]&~m[426]))&BiasedRNG[425])|(((m[70]&~m[171]&~m[426])|(~m[70]&m[171]&m[426]))&~BiasedRNG[425])|((~m[70]&~m[171]&m[426])|(m[70]&~m[171]&m[426])|(m[70]&m[171]&m[426]));
    m[283] = (((~m[70]&~m[183]&~m[427])|(m[70]&m[183]&~m[427]))&BiasedRNG[426])|(((m[70]&~m[183]&~m[427])|(~m[70]&m[183]&m[427]))&~BiasedRNG[426])|((~m[70]&~m[183]&m[427])|(m[70]&~m[183]&m[427])|(m[70]&m[183]&m[427]));
    m[284] = (((~m[71]&~m[195]&~m[428])|(m[71]&m[195]&~m[428]))&BiasedRNG[427])|(((m[71]&~m[195]&~m[428])|(~m[71]&m[195]&m[428]))&~BiasedRNG[427])|((~m[71]&~m[195]&m[428])|(m[71]&~m[195]&m[428])|(m[71]&m[195]&m[428]));
    m[285] = (((~m[71]&~m[207]&~m[429])|(m[71]&m[207]&~m[429]))&BiasedRNG[428])|(((m[71]&~m[207]&~m[429])|(~m[71]&m[207]&m[429]))&~BiasedRNG[428])|((~m[71]&~m[207]&m[429])|(m[71]&~m[207]&m[429])|(m[71]&m[207]&m[429]));
    m[286] = (((~m[71]&~m[219]&~m[430])|(m[71]&m[219]&~m[430]))&BiasedRNG[429])|(((m[71]&~m[219]&~m[430])|(~m[71]&m[219]&m[430]))&~BiasedRNG[429])|((~m[71]&~m[219]&m[430])|(m[71]&~m[219]&m[430])|(m[71]&m[219]&m[430]));
    m[287] = (((~m[71]&~m[231]&~m[431])|(m[71]&m[231]&~m[431]))&BiasedRNG[430])|(((m[71]&~m[231]&~m[431])|(~m[71]&m[231]&m[431]))&~BiasedRNG[430])|((~m[71]&~m[231]&m[431])|(m[71]&~m[231]&m[431])|(m[71]&m[231]&m[431]));
    m[288] = (((~m[72]&~m[100]&~m[432])|(m[72]&m[100]&~m[432]))&BiasedRNG[431])|(((m[72]&~m[100]&~m[432])|(~m[72]&m[100]&m[432]))&~BiasedRNG[431])|((~m[72]&~m[100]&m[432])|(m[72]&~m[100]&m[432])|(m[72]&m[100]&m[432]));
    m[289] = (((~m[72]&~m[112]&~m[433])|(m[72]&m[112]&~m[433]))&BiasedRNG[432])|(((m[72]&~m[112]&~m[433])|(~m[72]&m[112]&m[433]))&~BiasedRNG[432])|((~m[72]&~m[112]&m[433])|(m[72]&~m[112]&m[433])|(m[72]&m[112]&m[433]));
    m[290] = (((~m[72]&~m[124]&~m[434])|(m[72]&m[124]&~m[434]))&BiasedRNG[433])|(((m[72]&~m[124]&~m[434])|(~m[72]&m[124]&m[434]))&~BiasedRNG[433])|((~m[72]&~m[124]&m[434])|(m[72]&~m[124]&m[434])|(m[72]&m[124]&m[434]));
    m[291] = (((~m[72]&~m[136]&~m[435])|(m[72]&m[136]&~m[435]))&BiasedRNG[434])|(((m[72]&~m[136]&~m[435])|(~m[72]&m[136]&m[435]))&~BiasedRNG[434])|((~m[72]&~m[136]&m[435])|(m[72]&~m[136]&m[435])|(m[72]&m[136]&m[435]));
    m[292] = (((~m[73]&~m[148]&~m[436])|(m[73]&m[148]&~m[436]))&BiasedRNG[435])|(((m[73]&~m[148]&~m[436])|(~m[73]&m[148]&m[436]))&~BiasedRNG[435])|((~m[73]&~m[148]&m[436])|(m[73]&~m[148]&m[436])|(m[73]&m[148]&m[436]));
    m[293] = (((~m[73]&~m[160]&~m[437])|(m[73]&m[160]&~m[437]))&BiasedRNG[436])|(((m[73]&~m[160]&~m[437])|(~m[73]&m[160]&m[437]))&~BiasedRNG[436])|((~m[73]&~m[160]&m[437])|(m[73]&~m[160]&m[437])|(m[73]&m[160]&m[437]));
    m[294] = (((~m[73]&~m[172]&~m[438])|(m[73]&m[172]&~m[438]))&BiasedRNG[437])|(((m[73]&~m[172]&~m[438])|(~m[73]&m[172]&m[438]))&~BiasedRNG[437])|((~m[73]&~m[172]&m[438])|(m[73]&~m[172]&m[438])|(m[73]&m[172]&m[438]));
    m[295] = (((~m[73]&~m[184]&~m[439])|(m[73]&m[184]&~m[439]))&BiasedRNG[438])|(((m[73]&~m[184]&~m[439])|(~m[73]&m[184]&m[439]))&~BiasedRNG[438])|((~m[73]&~m[184]&m[439])|(m[73]&~m[184]&m[439])|(m[73]&m[184]&m[439]));
    m[296] = (((~m[74]&~m[196]&~m[440])|(m[74]&m[196]&~m[440]))&BiasedRNG[439])|(((m[74]&~m[196]&~m[440])|(~m[74]&m[196]&m[440]))&~BiasedRNG[439])|((~m[74]&~m[196]&m[440])|(m[74]&~m[196]&m[440])|(m[74]&m[196]&m[440]));
    m[297] = (((~m[74]&~m[208]&~m[441])|(m[74]&m[208]&~m[441]))&BiasedRNG[440])|(((m[74]&~m[208]&~m[441])|(~m[74]&m[208]&m[441]))&~BiasedRNG[440])|((~m[74]&~m[208]&m[441])|(m[74]&~m[208]&m[441])|(m[74]&m[208]&m[441]));
    m[298] = (((~m[74]&~m[220]&~m[442])|(m[74]&m[220]&~m[442]))&BiasedRNG[441])|(((m[74]&~m[220]&~m[442])|(~m[74]&m[220]&m[442]))&~BiasedRNG[441])|((~m[74]&~m[220]&m[442])|(m[74]&~m[220]&m[442])|(m[74]&m[220]&m[442]));
    m[299] = (((~m[74]&~m[232]&~m[443])|(m[74]&m[232]&~m[443]))&BiasedRNG[442])|(((m[74]&~m[232]&~m[443])|(~m[74]&m[232]&m[443]))&~BiasedRNG[442])|((~m[74]&~m[232]&m[443])|(m[74]&~m[232]&m[443])|(m[74]&m[232]&m[443]));
    m[300] = (((~m[75]&~m[101]&~m[444])|(m[75]&m[101]&~m[444]))&BiasedRNG[443])|(((m[75]&~m[101]&~m[444])|(~m[75]&m[101]&m[444]))&~BiasedRNG[443])|((~m[75]&~m[101]&m[444])|(m[75]&~m[101]&m[444])|(m[75]&m[101]&m[444]));
    m[301] = (((~m[75]&~m[113]&~m[445])|(m[75]&m[113]&~m[445]))&BiasedRNG[444])|(((m[75]&~m[113]&~m[445])|(~m[75]&m[113]&m[445]))&~BiasedRNG[444])|((~m[75]&~m[113]&m[445])|(m[75]&~m[113]&m[445])|(m[75]&m[113]&m[445]));
    m[302] = (((~m[75]&~m[125]&~m[446])|(m[75]&m[125]&~m[446]))&BiasedRNG[445])|(((m[75]&~m[125]&~m[446])|(~m[75]&m[125]&m[446]))&~BiasedRNG[445])|((~m[75]&~m[125]&m[446])|(m[75]&~m[125]&m[446])|(m[75]&m[125]&m[446]));
    m[303] = (((~m[75]&~m[137]&~m[447])|(m[75]&m[137]&~m[447]))&BiasedRNG[446])|(((m[75]&~m[137]&~m[447])|(~m[75]&m[137]&m[447]))&~BiasedRNG[446])|((~m[75]&~m[137]&m[447])|(m[75]&~m[137]&m[447])|(m[75]&m[137]&m[447]));
    m[304] = (((~m[76]&~m[149]&~m[448])|(m[76]&m[149]&~m[448]))&BiasedRNG[447])|(((m[76]&~m[149]&~m[448])|(~m[76]&m[149]&m[448]))&~BiasedRNG[447])|((~m[76]&~m[149]&m[448])|(m[76]&~m[149]&m[448])|(m[76]&m[149]&m[448]));
    m[305] = (((~m[76]&~m[161]&~m[449])|(m[76]&m[161]&~m[449]))&BiasedRNG[448])|(((m[76]&~m[161]&~m[449])|(~m[76]&m[161]&m[449]))&~BiasedRNG[448])|((~m[76]&~m[161]&m[449])|(m[76]&~m[161]&m[449])|(m[76]&m[161]&m[449]));
    m[306] = (((~m[76]&~m[173]&~m[450])|(m[76]&m[173]&~m[450]))&BiasedRNG[449])|(((m[76]&~m[173]&~m[450])|(~m[76]&m[173]&m[450]))&~BiasedRNG[449])|((~m[76]&~m[173]&m[450])|(m[76]&~m[173]&m[450])|(m[76]&m[173]&m[450]));
    m[307] = (((~m[76]&~m[185]&~m[451])|(m[76]&m[185]&~m[451]))&BiasedRNG[450])|(((m[76]&~m[185]&~m[451])|(~m[76]&m[185]&m[451]))&~BiasedRNG[450])|((~m[76]&~m[185]&m[451])|(m[76]&~m[185]&m[451])|(m[76]&m[185]&m[451]));
    m[308] = (((~m[77]&~m[197]&~m[452])|(m[77]&m[197]&~m[452]))&BiasedRNG[451])|(((m[77]&~m[197]&~m[452])|(~m[77]&m[197]&m[452]))&~BiasedRNG[451])|((~m[77]&~m[197]&m[452])|(m[77]&~m[197]&m[452])|(m[77]&m[197]&m[452]));
    m[309] = (((~m[77]&~m[209]&~m[453])|(m[77]&m[209]&~m[453]))&BiasedRNG[452])|(((m[77]&~m[209]&~m[453])|(~m[77]&m[209]&m[453]))&~BiasedRNG[452])|((~m[77]&~m[209]&m[453])|(m[77]&~m[209]&m[453])|(m[77]&m[209]&m[453]));
    m[310] = (((~m[77]&~m[221]&~m[454])|(m[77]&m[221]&~m[454]))&BiasedRNG[453])|(((m[77]&~m[221]&~m[454])|(~m[77]&m[221]&m[454]))&~BiasedRNG[453])|((~m[77]&~m[221]&m[454])|(m[77]&~m[221]&m[454])|(m[77]&m[221]&m[454]));
    m[311] = (((~m[77]&~m[233]&~m[455])|(m[77]&m[233]&~m[455]))&BiasedRNG[454])|(((m[77]&~m[233]&~m[455])|(~m[77]&m[233]&m[455]))&~BiasedRNG[454])|((~m[77]&~m[233]&m[455])|(m[77]&~m[233]&m[455])|(m[77]&m[233]&m[455]));
    m[312] = (((~m[78]&~m[102]&~m[456])|(m[78]&m[102]&~m[456]))&BiasedRNG[455])|(((m[78]&~m[102]&~m[456])|(~m[78]&m[102]&m[456]))&~BiasedRNG[455])|((~m[78]&~m[102]&m[456])|(m[78]&~m[102]&m[456])|(m[78]&m[102]&m[456]));
    m[313] = (((~m[78]&~m[114]&~m[457])|(m[78]&m[114]&~m[457]))&BiasedRNG[456])|(((m[78]&~m[114]&~m[457])|(~m[78]&m[114]&m[457]))&~BiasedRNG[456])|((~m[78]&~m[114]&m[457])|(m[78]&~m[114]&m[457])|(m[78]&m[114]&m[457]));
    m[314] = (((~m[78]&~m[126]&~m[458])|(m[78]&m[126]&~m[458]))&BiasedRNG[457])|(((m[78]&~m[126]&~m[458])|(~m[78]&m[126]&m[458]))&~BiasedRNG[457])|((~m[78]&~m[126]&m[458])|(m[78]&~m[126]&m[458])|(m[78]&m[126]&m[458]));
    m[315] = (((~m[78]&~m[138]&~m[459])|(m[78]&m[138]&~m[459]))&BiasedRNG[458])|(((m[78]&~m[138]&~m[459])|(~m[78]&m[138]&m[459]))&~BiasedRNG[458])|((~m[78]&~m[138]&m[459])|(m[78]&~m[138]&m[459])|(m[78]&m[138]&m[459]));
    m[316] = (((~m[79]&~m[150]&~m[460])|(m[79]&m[150]&~m[460]))&BiasedRNG[459])|(((m[79]&~m[150]&~m[460])|(~m[79]&m[150]&m[460]))&~BiasedRNG[459])|((~m[79]&~m[150]&m[460])|(m[79]&~m[150]&m[460])|(m[79]&m[150]&m[460]));
    m[317] = (((~m[79]&~m[162]&~m[461])|(m[79]&m[162]&~m[461]))&BiasedRNG[460])|(((m[79]&~m[162]&~m[461])|(~m[79]&m[162]&m[461]))&~BiasedRNG[460])|((~m[79]&~m[162]&m[461])|(m[79]&~m[162]&m[461])|(m[79]&m[162]&m[461]));
    m[318] = (((~m[79]&~m[174]&~m[462])|(m[79]&m[174]&~m[462]))&BiasedRNG[461])|(((m[79]&~m[174]&~m[462])|(~m[79]&m[174]&m[462]))&~BiasedRNG[461])|((~m[79]&~m[174]&m[462])|(m[79]&~m[174]&m[462])|(m[79]&m[174]&m[462]));
    m[319] = (((~m[79]&~m[186]&~m[463])|(m[79]&m[186]&~m[463]))&BiasedRNG[462])|(((m[79]&~m[186]&~m[463])|(~m[79]&m[186]&m[463]))&~BiasedRNG[462])|((~m[79]&~m[186]&m[463])|(m[79]&~m[186]&m[463])|(m[79]&m[186]&m[463]));
    m[320] = (((~m[80]&~m[198]&~m[464])|(m[80]&m[198]&~m[464]))&BiasedRNG[463])|(((m[80]&~m[198]&~m[464])|(~m[80]&m[198]&m[464]))&~BiasedRNG[463])|((~m[80]&~m[198]&m[464])|(m[80]&~m[198]&m[464])|(m[80]&m[198]&m[464]));
    m[321] = (((~m[80]&~m[210]&~m[465])|(m[80]&m[210]&~m[465]))&BiasedRNG[464])|(((m[80]&~m[210]&~m[465])|(~m[80]&m[210]&m[465]))&~BiasedRNG[464])|((~m[80]&~m[210]&m[465])|(m[80]&~m[210]&m[465])|(m[80]&m[210]&m[465]));
    m[322] = (((~m[80]&~m[222]&~m[466])|(m[80]&m[222]&~m[466]))&BiasedRNG[465])|(((m[80]&~m[222]&~m[466])|(~m[80]&m[222]&m[466]))&~BiasedRNG[465])|((~m[80]&~m[222]&m[466])|(m[80]&~m[222]&m[466])|(m[80]&m[222]&m[466]));
    m[323] = (((~m[80]&~m[234]&~m[467])|(m[80]&m[234]&~m[467]))&BiasedRNG[466])|(((m[80]&~m[234]&~m[467])|(~m[80]&m[234]&m[467]))&~BiasedRNG[466])|((~m[80]&~m[234]&m[467])|(m[80]&~m[234]&m[467])|(m[80]&m[234]&m[467]));
    m[324] = (((~m[81]&~m[103]&~m[468])|(m[81]&m[103]&~m[468]))&BiasedRNG[467])|(((m[81]&~m[103]&~m[468])|(~m[81]&m[103]&m[468]))&~BiasedRNG[467])|((~m[81]&~m[103]&m[468])|(m[81]&~m[103]&m[468])|(m[81]&m[103]&m[468]));
    m[325] = (((~m[81]&~m[115]&~m[469])|(m[81]&m[115]&~m[469]))&BiasedRNG[468])|(((m[81]&~m[115]&~m[469])|(~m[81]&m[115]&m[469]))&~BiasedRNG[468])|((~m[81]&~m[115]&m[469])|(m[81]&~m[115]&m[469])|(m[81]&m[115]&m[469]));
    m[326] = (((~m[81]&~m[127]&~m[470])|(m[81]&m[127]&~m[470]))&BiasedRNG[469])|(((m[81]&~m[127]&~m[470])|(~m[81]&m[127]&m[470]))&~BiasedRNG[469])|((~m[81]&~m[127]&m[470])|(m[81]&~m[127]&m[470])|(m[81]&m[127]&m[470]));
    m[327] = (((~m[81]&~m[139]&~m[471])|(m[81]&m[139]&~m[471]))&BiasedRNG[470])|(((m[81]&~m[139]&~m[471])|(~m[81]&m[139]&m[471]))&~BiasedRNG[470])|((~m[81]&~m[139]&m[471])|(m[81]&~m[139]&m[471])|(m[81]&m[139]&m[471]));
    m[328] = (((~m[82]&~m[151]&~m[472])|(m[82]&m[151]&~m[472]))&BiasedRNG[471])|(((m[82]&~m[151]&~m[472])|(~m[82]&m[151]&m[472]))&~BiasedRNG[471])|((~m[82]&~m[151]&m[472])|(m[82]&~m[151]&m[472])|(m[82]&m[151]&m[472]));
    m[329] = (((~m[82]&~m[163]&~m[473])|(m[82]&m[163]&~m[473]))&BiasedRNG[472])|(((m[82]&~m[163]&~m[473])|(~m[82]&m[163]&m[473]))&~BiasedRNG[472])|((~m[82]&~m[163]&m[473])|(m[82]&~m[163]&m[473])|(m[82]&m[163]&m[473]));
    m[330] = (((~m[82]&~m[175]&~m[474])|(m[82]&m[175]&~m[474]))&BiasedRNG[473])|(((m[82]&~m[175]&~m[474])|(~m[82]&m[175]&m[474]))&~BiasedRNG[473])|((~m[82]&~m[175]&m[474])|(m[82]&~m[175]&m[474])|(m[82]&m[175]&m[474]));
    m[331] = (((~m[82]&~m[187]&~m[475])|(m[82]&m[187]&~m[475]))&BiasedRNG[474])|(((m[82]&~m[187]&~m[475])|(~m[82]&m[187]&m[475]))&~BiasedRNG[474])|((~m[82]&~m[187]&m[475])|(m[82]&~m[187]&m[475])|(m[82]&m[187]&m[475]));
    m[332] = (((~m[83]&~m[199]&~m[476])|(m[83]&m[199]&~m[476]))&BiasedRNG[475])|(((m[83]&~m[199]&~m[476])|(~m[83]&m[199]&m[476]))&~BiasedRNG[475])|((~m[83]&~m[199]&m[476])|(m[83]&~m[199]&m[476])|(m[83]&m[199]&m[476]));
    m[333] = (((~m[83]&~m[211]&~m[477])|(m[83]&m[211]&~m[477]))&BiasedRNG[476])|(((m[83]&~m[211]&~m[477])|(~m[83]&m[211]&m[477]))&~BiasedRNG[476])|((~m[83]&~m[211]&m[477])|(m[83]&~m[211]&m[477])|(m[83]&m[211]&m[477]));
    m[334] = (((~m[83]&~m[223]&~m[478])|(m[83]&m[223]&~m[478]))&BiasedRNG[477])|(((m[83]&~m[223]&~m[478])|(~m[83]&m[223]&m[478]))&~BiasedRNG[477])|((~m[83]&~m[223]&m[478])|(m[83]&~m[223]&m[478])|(m[83]&m[223]&m[478]));
    m[335] = (((~m[83]&~m[235]&~m[479])|(m[83]&m[235]&~m[479]))&BiasedRNG[478])|(((m[83]&~m[235]&~m[479])|(~m[83]&m[235]&m[479]))&~BiasedRNG[478])|((~m[83]&~m[235]&m[479])|(m[83]&~m[235]&m[479])|(m[83]&m[235]&m[479]));
    m[336] = (((~m[84]&~m[104]&~m[480])|(m[84]&m[104]&~m[480]))&BiasedRNG[479])|(((m[84]&~m[104]&~m[480])|(~m[84]&m[104]&m[480]))&~BiasedRNG[479])|((~m[84]&~m[104]&m[480])|(m[84]&~m[104]&m[480])|(m[84]&m[104]&m[480]));
    m[337] = (((~m[84]&~m[116]&~m[481])|(m[84]&m[116]&~m[481]))&BiasedRNG[480])|(((m[84]&~m[116]&~m[481])|(~m[84]&m[116]&m[481]))&~BiasedRNG[480])|((~m[84]&~m[116]&m[481])|(m[84]&~m[116]&m[481])|(m[84]&m[116]&m[481]));
    m[338] = (((~m[84]&~m[128]&~m[482])|(m[84]&m[128]&~m[482]))&BiasedRNG[481])|(((m[84]&~m[128]&~m[482])|(~m[84]&m[128]&m[482]))&~BiasedRNG[481])|((~m[84]&~m[128]&m[482])|(m[84]&~m[128]&m[482])|(m[84]&m[128]&m[482]));
    m[339] = (((~m[84]&~m[140]&~m[483])|(m[84]&m[140]&~m[483]))&BiasedRNG[482])|(((m[84]&~m[140]&~m[483])|(~m[84]&m[140]&m[483]))&~BiasedRNG[482])|((~m[84]&~m[140]&m[483])|(m[84]&~m[140]&m[483])|(m[84]&m[140]&m[483]));
    m[340] = (((~m[85]&~m[152]&~m[484])|(m[85]&m[152]&~m[484]))&BiasedRNG[483])|(((m[85]&~m[152]&~m[484])|(~m[85]&m[152]&m[484]))&~BiasedRNG[483])|((~m[85]&~m[152]&m[484])|(m[85]&~m[152]&m[484])|(m[85]&m[152]&m[484]));
    m[341] = (((~m[85]&~m[164]&~m[485])|(m[85]&m[164]&~m[485]))&BiasedRNG[484])|(((m[85]&~m[164]&~m[485])|(~m[85]&m[164]&m[485]))&~BiasedRNG[484])|((~m[85]&~m[164]&m[485])|(m[85]&~m[164]&m[485])|(m[85]&m[164]&m[485]));
    m[342] = (((~m[85]&~m[176]&~m[486])|(m[85]&m[176]&~m[486]))&BiasedRNG[485])|(((m[85]&~m[176]&~m[486])|(~m[85]&m[176]&m[486]))&~BiasedRNG[485])|((~m[85]&~m[176]&m[486])|(m[85]&~m[176]&m[486])|(m[85]&m[176]&m[486]));
    m[343] = (((~m[85]&~m[188]&~m[487])|(m[85]&m[188]&~m[487]))&BiasedRNG[486])|(((m[85]&~m[188]&~m[487])|(~m[85]&m[188]&m[487]))&~BiasedRNG[486])|((~m[85]&~m[188]&m[487])|(m[85]&~m[188]&m[487])|(m[85]&m[188]&m[487]));
    m[344] = (((~m[86]&~m[200]&~m[488])|(m[86]&m[200]&~m[488]))&BiasedRNG[487])|(((m[86]&~m[200]&~m[488])|(~m[86]&m[200]&m[488]))&~BiasedRNG[487])|((~m[86]&~m[200]&m[488])|(m[86]&~m[200]&m[488])|(m[86]&m[200]&m[488]));
    m[345] = (((~m[86]&~m[212]&~m[489])|(m[86]&m[212]&~m[489]))&BiasedRNG[488])|(((m[86]&~m[212]&~m[489])|(~m[86]&m[212]&m[489]))&~BiasedRNG[488])|((~m[86]&~m[212]&m[489])|(m[86]&~m[212]&m[489])|(m[86]&m[212]&m[489]));
    m[346] = (((~m[86]&~m[224]&~m[490])|(m[86]&m[224]&~m[490]))&BiasedRNG[489])|(((m[86]&~m[224]&~m[490])|(~m[86]&m[224]&m[490]))&~BiasedRNG[489])|((~m[86]&~m[224]&m[490])|(m[86]&~m[224]&m[490])|(m[86]&m[224]&m[490]));
    m[347] = (((~m[86]&~m[236]&~m[491])|(m[86]&m[236]&~m[491]))&BiasedRNG[490])|(((m[86]&~m[236]&~m[491])|(~m[86]&m[236]&m[491]))&~BiasedRNG[490])|((~m[86]&~m[236]&m[491])|(m[86]&~m[236]&m[491])|(m[86]&m[236]&m[491]));
    m[348] = (((~m[87]&~m[105]&~m[492])|(m[87]&m[105]&~m[492]))&BiasedRNG[491])|(((m[87]&~m[105]&~m[492])|(~m[87]&m[105]&m[492]))&~BiasedRNG[491])|((~m[87]&~m[105]&m[492])|(m[87]&~m[105]&m[492])|(m[87]&m[105]&m[492]));
    m[349] = (((~m[87]&~m[117]&~m[493])|(m[87]&m[117]&~m[493]))&BiasedRNG[492])|(((m[87]&~m[117]&~m[493])|(~m[87]&m[117]&m[493]))&~BiasedRNG[492])|((~m[87]&~m[117]&m[493])|(m[87]&~m[117]&m[493])|(m[87]&m[117]&m[493]));
    m[350] = (((~m[87]&~m[129]&~m[494])|(m[87]&m[129]&~m[494]))&BiasedRNG[493])|(((m[87]&~m[129]&~m[494])|(~m[87]&m[129]&m[494]))&~BiasedRNG[493])|((~m[87]&~m[129]&m[494])|(m[87]&~m[129]&m[494])|(m[87]&m[129]&m[494]));
    m[351] = (((~m[87]&~m[141]&~m[495])|(m[87]&m[141]&~m[495]))&BiasedRNG[494])|(((m[87]&~m[141]&~m[495])|(~m[87]&m[141]&m[495]))&~BiasedRNG[494])|((~m[87]&~m[141]&m[495])|(m[87]&~m[141]&m[495])|(m[87]&m[141]&m[495]));
    m[352] = (((~m[88]&~m[153]&~m[496])|(m[88]&m[153]&~m[496]))&BiasedRNG[495])|(((m[88]&~m[153]&~m[496])|(~m[88]&m[153]&m[496]))&~BiasedRNG[495])|((~m[88]&~m[153]&m[496])|(m[88]&~m[153]&m[496])|(m[88]&m[153]&m[496]));
    m[353] = (((~m[88]&~m[165]&~m[497])|(m[88]&m[165]&~m[497]))&BiasedRNG[496])|(((m[88]&~m[165]&~m[497])|(~m[88]&m[165]&m[497]))&~BiasedRNG[496])|((~m[88]&~m[165]&m[497])|(m[88]&~m[165]&m[497])|(m[88]&m[165]&m[497]));
    m[354] = (((~m[88]&~m[177]&~m[498])|(m[88]&m[177]&~m[498]))&BiasedRNG[497])|(((m[88]&~m[177]&~m[498])|(~m[88]&m[177]&m[498]))&~BiasedRNG[497])|((~m[88]&~m[177]&m[498])|(m[88]&~m[177]&m[498])|(m[88]&m[177]&m[498]));
    m[355] = (((~m[88]&~m[189]&~m[499])|(m[88]&m[189]&~m[499]))&BiasedRNG[498])|(((m[88]&~m[189]&~m[499])|(~m[88]&m[189]&m[499]))&~BiasedRNG[498])|((~m[88]&~m[189]&m[499])|(m[88]&~m[189]&m[499])|(m[88]&m[189]&m[499]));
    m[356] = (((~m[89]&~m[201]&~m[500])|(m[89]&m[201]&~m[500]))&BiasedRNG[499])|(((m[89]&~m[201]&~m[500])|(~m[89]&m[201]&m[500]))&~BiasedRNG[499])|((~m[89]&~m[201]&m[500])|(m[89]&~m[201]&m[500])|(m[89]&m[201]&m[500]));
    m[357] = (((~m[89]&~m[213]&~m[501])|(m[89]&m[213]&~m[501]))&BiasedRNG[500])|(((m[89]&~m[213]&~m[501])|(~m[89]&m[213]&m[501]))&~BiasedRNG[500])|((~m[89]&~m[213]&m[501])|(m[89]&~m[213]&m[501])|(m[89]&m[213]&m[501]));
    m[358] = (((~m[89]&~m[225]&~m[502])|(m[89]&m[225]&~m[502]))&BiasedRNG[501])|(((m[89]&~m[225]&~m[502])|(~m[89]&m[225]&m[502]))&~BiasedRNG[501])|((~m[89]&~m[225]&m[502])|(m[89]&~m[225]&m[502])|(m[89]&m[225]&m[502]));
    m[359] = (((~m[89]&~m[237]&~m[503])|(m[89]&m[237]&~m[503]))&BiasedRNG[502])|(((m[89]&~m[237]&~m[503])|(~m[89]&m[237]&m[503]))&~BiasedRNG[502])|((~m[89]&~m[237]&m[503])|(m[89]&~m[237]&m[503])|(m[89]&m[237]&m[503]));
    m[360] = (((~m[90]&~m[106]&~m[504])|(m[90]&m[106]&~m[504]))&BiasedRNG[503])|(((m[90]&~m[106]&~m[504])|(~m[90]&m[106]&m[504]))&~BiasedRNG[503])|((~m[90]&~m[106]&m[504])|(m[90]&~m[106]&m[504])|(m[90]&m[106]&m[504]));
    m[361] = (((~m[90]&~m[118]&~m[505])|(m[90]&m[118]&~m[505]))&BiasedRNG[504])|(((m[90]&~m[118]&~m[505])|(~m[90]&m[118]&m[505]))&~BiasedRNG[504])|((~m[90]&~m[118]&m[505])|(m[90]&~m[118]&m[505])|(m[90]&m[118]&m[505]));
    m[362] = (((~m[90]&~m[130]&~m[506])|(m[90]&m[130]&~m[506]))&BiasedRNG[505])|(((m[90]&~m[130]&~m[506])|(~m[90]&m[130]&m[506]))&~BiasedRNG[505])|((~m[90]&~m[130]&m[506])|(m[90]&~m[130]&m[506])|(m[90]&m[130]&m[506]));
    m[363] = (((~m[90]&~m[142]&~m[507])|(m[90]&m[142]&~m[507]))&BiasedRNG[506])|(((m[90]&~m[142]&~m[507])|(~m[90]&m[142]&m[507]))&~BiasedRNG[506])|((~m[90]&~m[142]&m[507])|(m[90]&~m[142]&m[507])|(m[90]&m[142]&m[507]));
    m[364] = (((~m[91]&~m[154]&~m[508])|(m[91]&m[154]&~m[508]))&BiasedRNG[507])|(((m[91]&~m[154]&~m[508])|(~m[91]&m[154]&m[508]))&~BiasedRNG[507])|((~m[91]&~m[154]&m[508])|(m[91]&~m[154]&m[508])|(m[91]&m[154]&m[508]));
    m[365] = (((~m[91]&~m[166]&~m[509])|(m[91]&m[166]&~m[509]))&BiasedRNG[508])|(((m[91]&~m[166]&~m[509])|(~m[91]&m[166]&m[509]))&~BiasedRNG[508])|((~m[91]&~m[166]&m[509])|(m[91]&~m[166]&m[509])|(m[91]&m[166]&m[509]));
    m[366] = (((~m[91]&~m[178]&~m[510])|(m[91]&m[178]&~m[510]))&BiasedRNG[509])|(((m[91]&~m[178]&~m[510])|(~m[91]&m[178]&m[510]))&~BiasedRNG[509])|((~m[91]&~m[178]&m[510])|(m[91]&~m[178]&m[510])|(m[91]&m[178]&m[510]));
    m[367] = (((~m[91]&~m[190]&~m[511])|(m[91]&m[190]&~m[511]))&BiasedRNG[510])|(((m[91]&~m[190]&~m[511])|(~m[91]&m[190]&m[511]))&~BiasedRNG[510])|((~m[91]&~m[190]&m[511])|(m[91]&~m[190]&m[511])|(m[91]&m[190]&m[511]));
    m[368] = (((~m[92]&~m[202]&~m[512])|(m[92]&m[202]&~m[512]))&BiasedRNG[511])|(((m[92]&~m[202]&~m[512])|(~m[92]&m[202]&m[512]))&~BiasedRNG[511])|((~m[92]&~m[202]&m[512])|(m[92]&~m[202]&m[512])|(m[92]&m[202]&m[512]));
    m[369] = (((~m[92]&~m[214]&~m[513])|(m[92]&m[214]&~m[513]))&BiasedRNG[512])|(((m[92]&~m[214]&~m[513])|(~m[92]&m[214]&m[513]))&~BiasedRNG[512])|((~m[92]&~m[214]&m[513])|(m[92]&~m[214]&m[513])|(m[92]&m[214]&m[513]));
    m[370] = (((~m[92]&~m[226]&~m[514])|(m[92]&m[226]&~m[514]))&BiasedRNG[513])|(((m[92]&~m[226]&~m[514])|(~m[92]&m[226]&m[514]))&~BiasedRNG[513])|((~m[92]&~m[226]&m[514])|(m[92]&~m[226]&m[514])|(m[92]&m[226]&m[514]));
    m[371] = (((~m[92]&~m[238]&~m[515])|(m[92]&m[238]&~m[515]))&BiasedRNG[514])|(((m[92]&~m[238]&~m[515])|(~m[92]&m[238]&m[515]))&~BiasedRNG[514])|((~m[92]&~m[238]&m[515])|(m[92]&~m[238]&m[515])|(m[92]&m[238]&m[515]));
    m[372] = (((~m[93]&~m[107]&~m[516])|(m[93]&m[107]&~m[516]))&BiasedRNG[515])|(((m[93]&~m[107]&~m[516])|(~m[93]&m[107]&m[516]))&~BiasedRNG[515])|((~m[93]&~m[107]&m[516])|(m[93]&~m[107]&m[516])|(m[93]&m[107]&m[516]));
    m[373] = (((~m[93]&~m[119]&~m[517])|(m[93]&m[119]&~m[517]))&BiasedRNG[516])|(((m[93]&~m[119]&~m[517])|(~m[93]&m[119]&m[517]))&~BiasedRNG[516])|((~m[93]&~m[119]&m[517])|(m[93]&~m[119]&m[517])|(m[93]&m[119]&m[517]));
    m[374] = (((~m[93]&~m[131]&~m[518])|(m[93]&m[131]&~m[518]))&BiasedRNG[517])|(((m[93]&~m[131]&~m[518])|(~m[93]&m[131]&m[518]))&~BiasedRNG[517])|((~m[93]&~m[131]&m[518])|(m[93]&~m[131]&m[518])|(m[93]&m[131]&m[518]));
    m[375] = (((~m[93]&~m[143]&~m[519])|(m[93]&m[143]&~m[519]))&BiasedRNG[518])|(((m[93]&~m[143]&~m[519])|(~m[93]&m[143]&m[519]))&~BiasedRNG[518])|((~m[93]&~m[143]&m[519])|(m[93]&~m[143]&m[519])|(m[93]&m[143]&m[519]));
    m[376] = (((~m[94]&~m[155]&~m[520])|(m[94]&m[155]&~m[520]))&BiasedRNG[519])|(((m[94]&~m[155]&~m[520])|(~m[94]&m[155]&m[520]))&~BiasedRNG[519])|((~m[94]&~m[155]&m[520])|(m[94]&~m[155]&m[520])|(m[94]&m[155]&m[520]));
    m[377] = (((~m[94]&~m[167]&~m[521])|(m[94]&m[167]&~m[521]))&BiasedRNG[520])|(((m[94]&~m[167]&~m[521])|(~m[94]&m[167]&m[521]))&~BiasedRNG[520])|((~m[94]&~m[167]&m[521])|(m[94]&~m[167]&m[521])|(m[94]&m[167]&m[521]));
    m[378] = (((~m[94]&~m[179]&~m[522])|(m[94]&m[179]&~m[522]))&BiasedRNG[521])|(((m[94]&~m[179]&~m[522])|(~m[94]&m[179]&m[522]))&~BiasedRNG[521])|((~m[94]&~m[179]&m[522])|(m[94]&~m[179]&m[522])|(m[94]&m[179]&m[522]));
    m[379] = (((~m[94]&~m[191]&~m[523])|(m[94]&m[191]&~m[523]))&BiasedRNG[522])|(((m[94]&~m[191]&~m[523])|(~m[94]&m[191]&m[523]))&~BiasedRNG[522])|((~m[94]&~m[191]&m[523])|(m[94]&~m[191]&m[523])|(m[94]&m[191]&m[523]));
    m[380] = (((~m[95]&~m[203]&~m[524])|(m[95]&m[203]&~m[524]))&BiasedRNG[523])|(((m[95]&~m[203]&~m[524])|(~m[95]&m[203]&m[524]))&~BiasedRNG[523])|((~m[95]&~m[203]&m[524])|(m[95]&~m[203]&m[524])|(m[95]&m[203]&m[524]));
    m[381] = (((~m[95]&~m[215]&~m[525])|(m[95]&m[215]&~m[525]))&BiasedRNG[524])|(((m[95]&~m[215]&~m[525])|(~m[95]&m[215]&m[525]))&~BiasedRNG[524])|((~m[95]&~m[215]&m[525])|(m[95]&~m[215]&m[525])|(m[95]&m[215]&m[525]));
    m[382] = (((~m[95]&~m[227]&~m[526])|(m[95]&m[227]&~m[526]))&BiasedRNG[525])|(((m[95]&~m[227]&~m[526])|(~m[95]&m[227]&m[526]))&~BiasedRNG[525])|((~m[95]&~m[227]&m[526])|(m[95]&~m[227]&m[526])|(m[95]&m[227]&m[526]));
    m[383] = (((~m[95]&~m[239]&~m[527])|(m[95]&m[239]&~m[527]))&BiasedRNG[526])|(((m[95]&~m[239]&~m[527])|(~m[95]&m[239]&m[527]))&~BiasedRNG[526])|((~m[95]&~m[239]&m[527])|(m[95]&~m[239]&m[527])|(m[95]&m[239]&m[527]));
    m[529] = (((m[396]&~m[528]&~m[530]&~m[531]&~m[532])|(~m[396]&~m[528]&~m[530]&m[531]&~m[532])|(m[396]&m[528]&~m[530]&m[531]&~m[532])|(m[396]&~m[528]&m[530]&m[531]&~m[532])|(~m[396]&m[528]&~m[530]&~m[531]&m[532])|(~m[396]&~m[528]&m[530]&~m[531]&m[532])|(m[396]&m[528]&m[530]&~m[531]&m[532])|(~m[396]&m[528]&m[530]&m[531]&m[532]))&UnbiasedRNG[252])|((m[396]&~m[528]&~m[530]&m[531]&~m[532])|(~m[396]&~m[528]&~m[530]&~m[531]&m[532])|(m[396]&~m[528]&~m[530]&~m[531]&m[532])|(m[396]&m[528]&~m[530]&~m[531]&m[532])|(m[396]&~m[528]&m[530]&~m[531]&m[532])|(~m[396]&~m[528]&~m[530]&m[531]&m[532])|(m[396]&~m[528]&~m[530]&m[531]&m[532])|(~m[396]&m[528]&~m[530]&m[531]&m[532])|(m[396]&m[528]&~m[530]&m[531]&m[532])|(~m[396]&~m[528]&m[530]&m[531]&m[532])|(m[396]&~m[528]&m[530]&m[531]&m[532])|(m[396]&m[528]&m[530]&m[531]&m[532]));
    m[534] = (((m[397]&~m[533]&~m[535]&~m[536]&~m[537])|(~m[397]&~m[533]&~m[535]&m[536]&~m[537])|(m[397]&m[533]&~m[535]&m[536]&~m[537])|(m[397]&~m[533]&m[535]&m[536]&~m[537])|(~m[397]&m[533]&~m[535]&~m[536]&m[537])|(~m[397]&~m[533]&m[535]&~m[536]&m[537])|(m[397]&m[533]&m[535]&~m[536]&m[537])|(~m[397]&m[533]&m[535]&m[536]&m[537]))&UnbiasedRNG[253])|((m[397]&~m[533]&~m[535]&m[536]&~m[537])|(~m[397]&~m[533]&~m[535]&~m[536]&m[537])|(m[397]&~m[533]&~m[535]&~m[536]&m[537])|(m[397]&m[533]&~m[535]&~m[536]&m[537])|(m[397]&~m[533]&m[535]&~m[536]&m[537])|(~m[397]&~m[533]&~m[535]&m[536]&m[537])|(m[397]&~m[533]&~m[535]&m[536]&m[537])|(~m[397]&m[533]&~m[535]&m[536]&m[537])|(m[397]&m[533]&~m[535]&m[536]&m[537])|(~m[397]&~m[533]&m[535]&m[536]&m[537])|(m[397]&~m[533]&m[535]&m[536]&m[537])|(m[397]&m[533]&m[535]&m[536]&m[537]));
    m[539] = (((m[408]&~m[538]&~m[540]&~m[541]&~m[542])|(~m[408]&~m[538]&~m[540]&m[541]&~m[542])|(m[408]&m[538]&~m[540]&m[541]&~m[542])|(m[408]&~m[538]&m[540]&m[541]&~m[542])|(~m[408]&m[538]&~m[540]&~m[541]&m[542])|(~m[408]&~m[538]&m[540]&~m[541]&m[542])|(m[408]&m[538]&m[540]&~m[541]&m[542])|(~m[408]&m[538]&m[540]&m[541]&m[542]))&UnbiasedRNG[254])|((m[408]&~m[538]&~m[540]&m[541]&~m[542])|(~m[408]&~m[538]&~m[540]&~m[541]&m[542])|(m[408]&~m[538]&~m[540]&~m[541]&m[542])|(m[408]&m[538]&~m[540]&~m[541]&m[542])|(m[408]&~m[538]&m[540]&~m[541]&m[542])|(~m[408]&~m[538]&~m[540]&m[541]&m[542])|(m[408]&~m[538]&~m[540]&m[541]&m[542])|(~m[408]&m[538]&~m[540]&m[541]&m[542])|(m[408]&m[538]&~m[540]&m[541]&m[542])|(~m[408]&~m[538]&m[540]&m[541]&m[542])|(m[408]&~m[538]&m[540]&m[541]&m[542])|(m[408]&m[538]&m[540]&m[541]&m[542]));
    m[544] = (((m[398]&~m[543]&~m[545]&~m[546]&~m[547])|(~m[398]&~m[543]&~m[545]&m[546]&~m[547])|(m[398]&m[543]&~m[545]&m[546]&~m[547])|(m[398]&~m[543]&m[545]&m[546]&~m[547])|(~m[398]&m[543]&~m[545]&~m[546]&m[547])|(~m[398]&~m[543]&m[545]&~m[546]&m[547])|(m[398]&m[543]&m[545]&~m[546]&m[547])|(~m[398]&m[543]&m[545]&m[546]&m[547]))&UnbiasedRNG[255])|((m[398]&~m[543]&~m[545]&m[546]&~m[547])|(~m[398]&~m[543]&~m[545]&~m[546]&m[547])|(m[398]&~m[543]&~m[545]&~m[546]&m[547])|(m[398]&m[543]&~m[545]&~m[546]&m[547])|(m[398]&~m[543]&m[545]&~m[546]&m[547])|(~m[398]&~m[543]&~m[545]&m[546]&m[547])|(m[398]&~m[543]&~m[545]&m[546]&m[547])|(~m[398]&m[543]&~m[545]&m[546]&m[547])|(m[398]&m[543]&~m[545]&m[546]&m[547])|(~m[398]&~m[543]&m[545]&m[546]&m[547])|(m[398]&~m[543]&m[545]&m[546]&m[547])|(m[398]&m[543]&m[545]&m[546]&m[547]));
    m[549] = (((m[409]&~m[548]&~m[550]&~m[551]&~m[552])|(~m[409]&~m[548]&~m[550]&m[551]&~m[552])|(m[409]&m[548]&~m[550]&m[551]&~m[552])|(m[409]&~m[548]&m[550]&m[551]&~m[552])|(~m[409]&m[548]&~m[550]&~m[551]&m[552])|(~m[409]&~m[548]&m[550]&~m[551]&m[552])|(m[409]&m[548]&m[550]&~m[551]&m[552])|(~m[409]&m[548]&m[550]&m[551]&m[552]))&UnbiasedRNG[256])|((m[409]&~m[548]&~m[550]&m[551]&~m[552])|(~m[409]&~m[548]&~m[550]&~m[551]&m[552])|(m[409]&~m[548]&~m[550]&~m[551]&m[552])|(m[409]&m[548]&~m[550]&~m[551]&m[552])|(m[409]&~m[548]&m[550]&~m[551]&m[552])|(~m[409]&~m[548]&~m[550]&m[551]&m[552])|(m[409]&~m[548]&~m[550]&m[551]&m[552])|(~m[409]&m[548]&~m[550]&m[551]&m[552])|(m[409]&m[548]&~m[550]&m[551]&m[552])|(~m[409]&~m[548]&m[550]&m[551]&m[552])|(m[409]&~m[548]&m[550]&m[551]&m[552])|(m[409]&m[548]&m[550]&m[551]&m[552]));
    m[554] = (((m[420]&~m[553]&~m[555]&~m[556]&~m[557])|(~m[420]&~m[553]&~m[555]&m[556]&~m[557])|(m[420]&m[553]&~m[555]&m[556]&~m[557])|(m[420]&~m[553]&m[555]&m[556]&~m[557])|(~m[420]&m[553]&~m[555]&~m[556]&m[557])|(~m[420]&~m[553]&m[555]&~m[556]&m[557])|(m[420]&m[553]&m[555]&~m[556]&m[557])|(~m[420]&m[553]&m[555]&m[556]&m[557]))&UnbiasedRNG[257])|((m[420]&~m[553]&~m[555]&m[556]&~m[557])|(~m[420]&~m[553]&~m[555]&~m[556]&m[557])|(m[420]&~m[553]&~m[555]&~m[556]&m[557])|(m[420]&m[553]&~m[555]&~m[556]&m[557])|(m[420]&~m[553]&m[555]&~m[556]&m[557])|(~m[420]&~m[553]&~m[555]&m[556]&m[557])|(m[420]&~m[553]&~m[555]&m[556]&m[557])|(~m[420]&m[553]&~m[555]&m[556]&m[557])|(m[420]&m[553]&~m[555]&m[556]&m[557])|(~m[420]&~m[553]&m[555]&m[556]&m[557])|(m[420]&~m[553]&m[555]&m[556]&m[557])|(m[420]&m[553]&m[555]&m[556]&m[557]));
    m[559] = (((m[399]&~m[558]&~m[560]&~m[561]&~m[562])|(~m[399]&~m[558]&~m[560]&m[561]&~m[562])|(m[399]&m[558]&~m[560]&m[561]&~m[562])|(m[399]&~m[558]&m[560]&m[561]&~m[562])|(~m[399]&m[558]&~m[560]&~m[561]&m[562])|(~m[399]&~m[558]&m[560]&~m[561]&m[562])|(m[399]&m[558]&m[560]&~m[561]&m[562])|(~m[399]&m[558]&m[560]&m[561]&m[562]))&UnbiasedRNG[258])|((m[399]&~m[558]&~m[560]&m[561]&~m[562])|(~m[399]&~m[558]&~m[560]&~m[561]&m[562])|(m[399]&~m[558]&~m[560]&~m[561]&m[562])|(m[399]&m[558]&~m[560]&~m[561]&m[562])|(m[399]&~m[558]&m[560]&~m[561]&m[562])|(~m[399]&~m[558]&~m[560]&m[561]&m[562])|(m[399]&~m[558]&~m[560]&m[561]&m[562])|(~m[399]&m[558]&~m[560]&m[561]&m[562])|(m[399]&m[558]&~m[560]&m[561]&m[562])|(~m[399]&~m[558]&m[560]&m[561]&m[562])|(m[399]&~m[558]&m[560]&m[561]&m[562])|(m[399]&m[558]&m[560]&m[561]&m[562]));
    m[564] = (((m[410]&~m[563]&~m[565]&~m[566]&~m[567])|(~m[410]&~m[563]&~m[565]&m[566]&~m[567])|(m[410]&m[563]&~m[565]&m[566]&~m[567])|(m[410]&~m[563]&m[565]&m[566]&~m[567])|(~m[410]&m[563]&~m[565]&~m[566]&m[567])|(~m[410]&~m[563]&m[565]&~m[566]&m[567])|(m[410]&m[563]&m[565]&~m[566]&m[567])|(~m[410]&m[563]&m[565]&m[566]&m[567]))&UnbiasedRNG[259])|((m[410]&~m[563]&~m[565]&m[566]&~m[567])|(~m[410]&~m[563]&~m[565]&~m[566]&m[567])|(m[410]&~m[563]&~m[565]&~m[566]&m[567])|(m[410]&m[563]&~m[565]&~m[566]&m[567])|(m[410]&~m[563]&m[565]&~m[566]&m[567])|(~m[410]&~m[563]&~m[565]&m[566]&m[567])|(m[410]&~m[563]&~m[565]&m[566]&m[567])|(~m[410]&m[563]&~m[565]&m[566]&m[567])|(m[410]&m[563]&~m[565]&m[566]&m[567])|(~m[410]&~m[563]&m[565]&m[566]&m[567])|(m[410]&~m[563]&m[565]&m[566]&m[567])|(m[410]&m[563]&m[565]&m[566]&m[567]));
    m[569] = (((m[421]&~m[568]&~m[570]&~m[571]&~m[572])|(~m[421]&~m[568]&~m[570]&m[571]&~m[572])|(m[421]&m[568]&~m[570]&m[571]&~m[572])|(m[421]&~m[568]&m[570]&m[571]&~m[572])|(~m[421]&m[568]&~m[570]&~m[571]&m[572])|(~m[421]&~m[568]&m[570]&~m[571]&m[572])|(m[421]&m[568]&m[570]&~m[571]&m[572])|(~m[421]&m[568]&m[570]&m[571]&m[572]))&UnbiasedRNG[260])|((m[421]&~m[568]&~m[570]&m[571]&~m[572])|(~m[421]&~m[568]&~m[570]&~m[571]&m[572])|(m[421]&~m[568]&~m[570]&~m[571]&m[572])|(m[421]&m[568]&~m[570]&~m[571]&m[572])|(m[421]&~m[568]&m[570]&~m[571]&m[572])|(~m[421]&~m[568]&~m[570]&m[571]&m[572])|(m[421]&~m[568]&~m[570]&m[571]&m[572])|(~m[421]&m[568]&~m[570]&m[571]&m[572])|(m[421]&m[568]&~m[570]&m[571]&m[572])|(~m[421]&~m[568]&m[570]&m[571]&m[572])|(m[421]&~m[568]&m[570]&m[571]&m[572])|(m[421]&m[568]&m[570]&m[571]&m[572]));
    m[574] = (((m[432]&~m[573]&~m[575]&~m[576]&~m[577])|(~m[432]&~m[573]&~m[575]&m[576]&~m[577])|(m[432]&m[573]&~m[575]&m[576]&~m[577])|(m[432]&~m[573]&m[575]&m[576]&~m[577])|(~m[432]&m[573]&~m[575]&~m[576]&m[577])|(~m[432]&~m[573]&m[575]&~m[576]&m[577])|(m[432]&m[573]&m[575]&~m[576]&m[577])|(~m[432]&m[573]&m[575]&m[576]&m[577]))&UnbiasedRNG[261])|((m[432]&~m[573]&~m[575]&m[576]&~m[577])|(~m[432]&~m[573]&~m[575]&~m[576]&m[577])|(m[432]&~m[573]&~m[575]&~m[576]&m[577])|(m[432]&m[573]&~m[575]&~m[576]&m[577])|(m[432]&~m[573]&m[575]&~m[576]&m[577])|(~m[432]&~m[573]&~m[575]&m[576]&m[577])|(m[432]&~m[573]&~m[575]&m[576]&m[577])|(~m[432]&m[573]&~m[575]&m[576]&m[577])|(m[432]&m[573]&~m[575]&m[576]&m[577])|(~m[432]&~m[573]&m[575]&m[576]&m[577])|(m[432]&~m[573]&m[575]&m[576]&m[577])|(m[432]&m[573]&m[575]&m[576]&m[577]));
    m[579] = (((m[400]&~m[578]&~m[580]&~m[581]&~m[582])|(~m[400]&~m[578]&~m[580]&m[581]&~m[582])|(m[400]&m[578]&~m[580]&m[581]&~m[582])|(m[400]&~m[578]&m[580]&m[581]&~m[582])|(~m[400]&m[578]&~m[580]&~m[581]&m[582])|(~m[400]&~m[578]&m[580]&~m[581]&m[582])|(m[400]&m[578]&m[580]&~m[581]&m[582])|(~m[400]&m[578]&m[580]&m[581]&m[582]))&UnbiasedRNG[262])|((m[400]&~m[578]&~m[580]&m[581]&~m[582])|(~m[400]&~m[578]&~m[580]&~m[581]&m[582])|(m[400]&~m[578]&~m[580]&~m[581]&m[582])|(m[400]&m[578]&~m[580]&~m[581]&m[582])|(m[400]&~m[578]&m[580]&~m[581]&m[582])|(~m[400]&~m[578]&~m[580]&m[581]&m[582])|(m[400]&~m[578]&~m[580]&m[581]&m[582])|(~m[400]&m[578]&~m[580]&m[581]&m[582])|(m[400]&m[578]&~m[580]&m[581]&m[582])|(~m[400]&~m[578]&m[580]&m[581]&m[582])|(m[400]&~m[578]&m[580]&m[581]&m[582])|(m[400]&m[578]&m[580]&m[581]&m[582]));
    m[584] = (((m[411]&~m[583]&~m[585]&~m[586]&~m[587])|(~m[411]&~m[583]&~m[585]&m[586]&~m[587])|(m[411]&m[583]&~m[585]&m[586]&~m[587])|(m[411]&~m[583]&m[585]&m[586]&~m[587])|(~m[411]&m[583]&~m[585]&~m[586]&m[587])|(~m[411]&~m[583]&m[585]&~m[586]&m[587])|(m[411]&m[583]&m[585]&~m[586]&m[587])|(~m[411]&m[583]&m[585]&m[586]&m[587]))&UnbiasedRNG[263])|((m[411]&~m[583]&~m[585]&m[586]&~m[587])|(~m[411]&~m[583]&~m[585]&~m[586]&m[587])|(m[411]&~m[583]&~m[585]&~m[586]&m[587])|(m[411]&m[583]&~m[585]&~m[586]&m[587])|(m[411]&~m[583]&m[585]&~m[586]&m[587])|(~m[411]&~m[583]&~m[585]&m[586]&m[587])|(m[411]&~m[583]&~m[585]&m[586]&m[587])|(~m[411]&m[583]&~m[585]&m[586]&m[587])|(m[411]&m[583]&~m[585]&m[586]&m[587])|(~m[411]&~m[583]&m[585]&m[586]&m[587])|(m[411]&~m[583]&m[585]&m[586]&m[587])|(m[411]&m[583]&m[585]&m[586]&m[587]));
    m[589] = (((m[422]&~m[588]&~m[590]&~m[591]&~m[592])|(~m[422]&~m[588]&~m[590]&m[591]&~m[592])|(m[422]&m[588]&~m[590]&m[591]&~m[592])|(m[422]&~m[588]&m[590]&m[591]&~m[592])|(~m[422]&m[588]&~m[590]&~m[591]&m[592])|(~m[422]&~m[588]&m[590]&~m[591]&m[592])|(m[422]&m[588]&m[590]&~m[591]&m[592])|(~m[422]&m[588]&m[590]&m[591]&m[592]))&UnbiasedRNG[264])|((m[422]&~m[588]&~m[590]&m[591]&~m[592])|(~m[422]&~m[588]&~m[590]&~m[591]&m[592])|(m[422]&~m[588]&~m[590]&~m[591]&m[592])|(m[422]&m[588]&~m[590]&~m[591]&m[592])|(m[422]&~m[588]&m[590]&~m[591]&m[592])|(~m[422]&~m[588]&~m[590]&m[591]&m[592])|(m[422]&~m[588]&~m[590]&m[591]&m[592])|(~m[422]&m[588]&~m[590]&m[591]&m[592])|(m[422]&m[588]&~m[590]&m[591]&m[592])|(~m[422]&~m[588]&m[590]&m[591]&m[592])|(m[422]&~m[588]&m[590]&m[591]&m[592])|(m[422]&m[588]&m[590]&m[591]&m[592]));
    m[594] = (((m[433]&~m[593]&~m[595]&~m[596]&~m[597])|(~m[433]&~m[593]&~m[595]&m[596]&~m[597])|(m[433]&m[593]&~m[595]&m[596]&~m[597])|(m[433]&~m[593]&m[595]&m[596]&~m[597])|(~m[433]&m[593]&~m[595]&~m[596]&m[597])|(~m[433]&~m[593]&m[595]&~m[596]&m[597])|(m[433]&m[593]&m[595]&~m[596]&m[597])|(~m[433]&m[593]&m[595]&m[596]&m[597]))&UnbiasedRNG[265])|((m[433]&~m[593]&~m[595]&m[596]&~m[597])|(~m[433]&~m[593]&~m[595]&~m[596]&m[597])|(m[433]&~m[593]&~m[595]&~m[596]&m[597])|(m[433]&m[593]&~m[595]&~m[596]&m[597])|(m[433]&~m[593]&m[595]&~m[596]&m[597])|(~m[433]&~m[593]&~m[595]&m[596]&m[597])|(m[433]&~m[593]&~m[595]&m[596]&m[597])|(~m[433]&m[593]&~m[595]&m[596]&m[597])|(m[433]&m[593]&~m[595]&m[596]&m[597])|(~m[433]&~m[593]&m[595]&m[596]&m[597])|(m[433]&~m[593]&m[595]&m[596]&m[597])|(m[433]&m[593]&m[595]&m[596]&m[597]));
    m[599] = (((m[444]&~m[598]&~m[600]&~m[601]&~m[602])|(~m[444]&~m[598]&~m[600]&m[601]&~m[602])|(m[444]&m[598]&~m[600]&m[601]&~m[602])|(m[444]&~m[598]&m[600]&m[601]&~m[602])|(~m[444]&m[598]&~m[600]&~m[601]&m[602])|(~m[444]&~m[598]&m[600]&~m[601]&m[602])|(m[444]&m[598]&m[600]&~m[601]&m[602])|(~m[444]&m[598]&m[600]&m[601]&m[602]))&UnbiasedRNG[266])|((m[444]&~m[598]&~m[600]&m[601]&~m[602])|(~m[444]&~m[598]&~m[600]&~m[601]&m[602])|(m[444]&~m[598]&~m[600]&~m[601]&m[602])|(m[444]&m[598]&~m[600]&~m[601]&m[602])|(m[444]&~m[598]&m[600]&~m[601]&m[602])|(~m[444]&~m[598]&~m[600]&m[601]&m[602])|(m[444]&~m[598]&~m[600]&m[601]&m[602])|(~m[444]&m[598]&~m[600]&m[601]&m[602])|(m[444]&m[598]&~m[600]&m[601]&m[602])|(~m[444]&~m[598]&m[600]&m[601]&m[602])|(m[444]&~m[598]&m[600]&m[601]&m[602])|(m[444]&m[598]&m[600]&m[601]&m[602]));
    m[604] = (((m[401]&~m[603]&~m[605]&~m[606]&~m[607])|(~m[401]&~m[603]&~m[605]&m[606]&~m[607])|(m[401]&m[603]&~m[605]&m[606]&~m[607])|(m[401]&~m[603]&m[605]&m[606]&~m[607])|(~m[401]&m[603]&~m[605]&~m[606]&m[607])|(~m[401]&~m[603]&m[605]&~m[606]&m[607])|(m[401]&m[603]&m[605]&~m[606]&m[607])|(~m[401]&m[603]&m[605]&m[606]&m[607]))&UnbiasedRNG[267])|((m[401]&~m[603]&~m[605]&m[606]&~m[607])|(~m[401]&~m[603]&~m[605]&~m[606]&m[607])|(m[401]&~m[603]&~m[605]&~m[606]&m[607])|(m[401]&m[603]&~m[605]&~m[606]&m[607])|(m[401]&~m[603]&m[605]&~m[606]&m[607])|(~m[401]&~m[603]&~m[605]&m[606]&m[607])|(m[401]&~m[603]&~m[605]&m[606]&m[607])|(~m[401]&m[603]&~m[605]&m[606]&m[607])|(m[401]&m[603]&~m[605]&m[606]&m[607])|(~m[401]&~m[603]&m[605]&m[606]&m[607])|(m[401]&~m[603]&m[605]&m[606]&m[607])|(m[401]&m[603]&m[605]&m[606]&m[607]));
    m[609] = (((m[412]&~m[608]&~m[610]&~m[611]&~m[612])|(~m[412]&~m[608]&~m[610]&m[611]&~m[612])|(m[412]&m[608]&~m[610]&m[611]&~m[612])|(m[412]&~m[608]&m[610]&m[611]&~m[612])|(~m[412]&m[608]&~m[610]&~m[611]&m[612])|(~m[412]&~m[608]&m[610]&~m[611]&m[612])|(m[412]&m[608]&m[610]&~m[611]&m[612])|(~m[412]&m[608]&m[610]&m[611]&m[612]))&UnbiasedRNG[268])|((m[412]&~m[608]&~m[610]&m[611]&~m[612])|(~m[412]&~m[608]&~m[610]&~m[611]&m[612])|(m[412]&~m[608]&~m[610]&~m[611]&m[612])|(m[412]&m[608]&~m[610]&~m[611]&m[612])|(m[412]&~m[608]&m[610]&~m[611]&m[612])|(~m[412]&~m[608]&~m[610]&m[611]&m[612])|(m[412]&~m[608]&~m[610]&m[611]&m[612])|(~m[412]&m[608]&~m[610]&m[611]&m[612])|(m[412]&m[608]&~m[610]&m[611]&m[612])|(~m[412]&~m[608]&m[610]&m[611]&m[612])|(m[412]&~m[608]&m[610]&m[611]&m[612])|(m[412]&m[608]&m[610]&m[611]&m[612]));
    m[614] = (((m[423]&~m[613]&~m[615]&~m[616]&~m[617])|(~m[423]&~m[613]&~m[615]&m[616]&~m[617])|(m[423]&m[613]&~m[615]&m[616]&~m[617])|(m[423]&~m[613]&m[615]&m[616]&~m[617])|(~m[423]&m[613]&~m[615]&~m[616]&m[617])|(~m[423]&~m[613]&m[615]&~m[616]&m[617])|(m[423]&m[613]&m[615]&~m[616]&m[617])|(~m[423]&m[613]&m[615]&m[616]&m[617]))&UnbiasedRNG[269])|((m[423]&~m[613]&~m[615]&m[616]&~m[617])|(~m[423]&~m[613]&~m[615]&~m[616]&m[617])|(m[423]&~m[613]&~m[615]&~m[616]&m[617])|(m[423]&m[613]&~m[615]&~m[616]&m[617])|(m[423]&~m[613]&m[615]&~m[616]&m[617])|(~m[423]&~m[613]&~m[615]&m[616]&m[617])|(m[423]&~m[613]&~m[615]&m[616]&m[617])|(~m[423]&m[613]&~m[615]&m[616]&m[617])|(m[423]&m[613]&~m[615]&m[616]&m[617])|(~m[423]&~m[613]&m[615]&m[616]&m[617])|(m[423]&~m[613]&m[615]&m[616]&m[617])|(m[423]&m[613]&m[615]&m[616]&m[617]));
    m[619] = (((m[434]&~m[618]&~m[620]&~m[621]&~m[622])|(~m[434]&~m[618]&~m[620]&m[621]&~m[622])|(m[434]&m[618]&~m[620]&m[621]&~m[622])|(m[434]&~m[618]&m[620]&m[621]&~m[622])|(~m[434]&m[618]&~m[620]&~m[621]&m[622])|(~m[434]&~m[618]&m[620]&~m[621]&m[622])|(m[434]&m[618]&m[620]&~m[621]&m[622])|(~m[434]&m[618]&m[620]&m[621]&m[622]))&UnbiasedRNG[270])|((m[434]&~m[618]&~m[620]&m[621]&~m[622])|(~m[434]&~m[618]&~m[620]&~m[621]&m[622])|(m[434]&~m[618]&~m[620]&~m[621]&m[622])|(m[434]&m[618]&~m[620]&~m[621]&m[622])|(m[434]&~m[618]&m[620]&~m[621]&m[622])|(~m[434]&~m[618]&~m[620]&m[621]&m[622])|(m[434]&~m[618]&~m[620]&m[621]&m[622])|(~m[434]&m[618]&~m[620]&m[621]&m[622])|(m[434]&m[618]&~m[620]&m[621]&m[622])|(~m[434]&~m[618]&m[620]&m[621]&m[622])|(m[434]&~m[618]&m[620]&m[621]&m[622])|(m[434]&m[618]&m[620]&m[621]&m[622]));
    m[624] = (((m[445]&~m[623]&~m[625]&~m[626]&~m[627])|(~m[445]&~m[623]&~m[625]&m[626]&~m[627])|(m[445]&m[623]&~m[625]&m[626]&~m[627])|(m[445]&~m[623]&m[625]&m[626]&~m[627])|(~m[445]&m[623]&~m[625]&~m[626]&m[627])|(~m[445]&~m[623]&m[625]&~m[626]&m[627])|(m[445]&m[623]&m[625]&~m[626]&m[627])|(~m[445]&m[623]&m[625]&m[626]&m[627]))&UnbiasedRNG[271])|((m[445]&~m[623]&~m[625]&m[626]&~m[627])|(~m[445]&~m[623]&~m[625]&~m[626]&m[627])|(m[445]&~m[623]&~m[625]&~m[626]&m[627])|(m[445]&m[623]&~m[625]&~m[626]&m[627])|(m[445]&~m[623]&m[625]&~m[626]&m[627])|(~m[445]&~m[623]&~m[625]&m[626]&m[627])|(m[445]&~m[623]&~m[625]&m[626]&m[627])|(~m[445]&m[623]&~m[625]&m[626]&m[627])|(m[445]&m[623]&~m[625]&m[626]&m[627])|(~m[445]&~m[623]&m[625]&m[626]&m[627])|(m[445]&~m[623]&m[625]&m[626]&m[627])|(m[445]&m[623]&m[625]&m[626]&m[627]));
    m[629] = (((m[456]&~m[628]&~m[630]&~m[631]&~m[632])|(~m[456]&~m[628]&~m[630]&m[631]&~m[632])|(m[456]&m[628]&~m[630]&m[631]&~m[632])|(m[456]&~m[628]&m[630]&m[631]&~m[632])|(~m[456]&m[628]&~m[630]&~m[631]&m[632])|(~m[456]&~m[628]&m[630]&~m[631]&m[632])|(m[456]&m[628]&m[630]&~m[631]&m[632])|(~m[456]&m[628]&m[630]&m[631]&m[632]))&UnbiasedRNG[272])|((m[456]&~m[628]&~m[630]&m[631]&~m[632])|(~m[456]&~m[628]&~m[630]&~m[631]&m[632])|(m[456]&~m[628]&~m[630]&~m[631]&m[632])|(m[456]&m[628]&~m[630]&~m[631]&m[632])|(m[456]&~m[628]&m[630]&~m[631]&m[632])|(~m[456]&~m[628]&~m[630]&m[631]&m[632])|(m[456]&~m[628]&~m[630]&m[631]&m[632])|(~m[456]&m[628]&~m[630]&m[631]&m[632])|(m[456]&m[628]&~m[630]&m[631]&m[632])|(~m[456]&~m[628]&m[630]&m[631]&m[632])|(m[456]&~m[628]&m[630]&m[631]&m[632])|(m[456]&m[628]&m[630]&m[631]&m[632]));
    m[634] = (((m[402]&~m[633]&~m[635]&~m[636]&~m[637])|(~m[402]&~m[633]&~m[635]&m[636]&~m[637])|(m[402]&m[633]&~m[635]&m[636]&~m[637])|(m[402]&~m[633]&m[635]&m[636]&~m[637])|(~m[402]&m[633]&~m[635]&~m[636]&m[637])|(~m[402]&~m[633]&m[635]&~m[636]&m[637])|(m[402]&m[633]&m[635]&~m[636]&m[637])|(~m[402]&m[633]&m[635]&m[636]&m[637]))&UnbiasedRNG[273])|((m[402]&~m[633]&~m[635]&m[636]&~m[637])|(~m[402]&~m[633]&~m[635]&~m[636]&m[637])|(m[402]&~m[633]&~m[635]&~m[636]&m[637])|(m[402]&m[633]&~m[635]&~m[636]&m[637])|(m[402]&~m[633]&m[635]&~m[636]&m[637])|(~m[402]&~m[633]&~m[635]&m[636]&m[637])|(m[402]&~m[633]&~m[635]&m[636]&m[637])|(~m[402]&m[633]&~m[635]&m[636]&m[637])|(m[402]&m[633]&~m[635]&m[636]&m[637])|(~m[402]&~m[633]&m[635]&m[636]&m[637])|(m[402]&~m[633]&m[635]&m[636]&m[637])|(m[402]&m[633]&m[635]&m[636]&m[637]));
    m[639] = (((m[413]&~m[638]&~m[640]&~m[641]&~m[642])|(~m[413]&~m[638]&~m[640]&m[641]&~m[642])|(m[413]&m[638]&~m[640]&m[641]&~m[642])|(m[413]&~m[638]&m[640]&m[641]&~m[642])|(~m[413]&m[638]&~m[640]&~m[641]&m[642])|(~m[413]&~m[638]&m[640]&~m[641]&m[642])|(m[413]&m[638]&m[640]&~m[641]&m[642])|(~m[413]&m[638]&m[640]&m[641]&m[642]))&UnbiasedRNG[274])|((m[413]&~m[638]&~m[640]&m[641]&~m[642])|(~m[413]&~m[638]&~m[640]&~m[641]&m[642])|(m[413]&~m[638]&~m[640]&~m[641]&m[642])|(m[413]&m[638]&~m[640]&~m[641]&m[642])|(m[413]&~m[638]&m[640]&~m[641]&m[642])|(~m[413]&~m[638]&~m[640]&m[641]&m[642])|(m[413]&~m[638]&~m[640]&m[641]&m[642])|(~m[413]&m[638]&~m[640]&m[641]&m[642])|(m[413]&m[638]&~m[640]&m[641]&m[642])|(~m[413]&~m[638]&m[640]&m[641]&m[642])|(m[413]&~m[638]&m[640]&m[641]&m[642])|(m[413]&m[638]&m[640]&m[641]&m[642]));
    m[644] = (((m[424]&~m[643]&~m[645]&~m[646]&~m[647])|(~m[424]&~m[643]&~m[645]&m[646]&~m[647])|(m[424]&m[643]&~m[645]&m[646]&~m[647])|(m[424]&~m[643]&m[645]&m[646]&~m[647])|(~m[424]&m[643]&~m[645]&~m[646]&m[647])|(~m[424]&~m[643]&m[645]&~m[646]&m[647])|(m[424]&m[643]&m[645]&~m[646]&m[647])|(~m[424]&m[643]&m[645]&m[646]&m[647]))&UnbiasedRNG[275])|((m[424]&~m[643]&~m[645]&m[646]&~m[647])|(~m[424]&~m[643]&~m[645]&~m[646]&m[647])|(m[424]&~m[643]&~m[645]&~m[646]&m[647])|(m[424]&m[643]&~m[645]&~m[646]&m[647])|(m[424]&~m[643]&m[645]&~m[646]&m[647])|(~m[424]&~m[643]&~m[645]&m[646]&m[647])|(m[424]&~m[643]&~m[645]&m[646]&m[647])|(~m[424]&m[643]&~m[645]&m[646]&m[647])|(m[424]&m[643]&~m[645]&m[646]&m[647])|(~m[424]&~m[643]&m[645]&m[646]&m[647])|(m[424]&~m[643]&m[645]&m[646]&m[647])|(m[424]&m[643]&m[645]&m[646]&m[647]));
    m[649] = (((m[435]&~m[648]&~m[650]&~m[651]&~m[652])|(~m[435]&~m[648]&~m[650]&m[651]&~m[652])|(m[435]&m[648]&~m[650]&m[651]&~m[652])|(m[435]&~m[648]&m[650]&m[651]&~m[652])|(~m[435]&m[648]&~m[650]&~m[651]&m[652])|(~m[435]&~m[648]&m[650]&~m[651]&m[652])|(m[435]&m[648]&m[650]&~m[651]&m[652])|(~m[435]&m[648]&m[650]&m[651]&m[652]))&UnbiasedRNG[276])|((m[435]&~m[648]&~m[650]&m[651]&~m[652])|(~m[435]&~m[648]&~m[650]&~m[651]&m[652])|(m[435]&~m[648]&~m[650]&~m[651]&m[652])|(m[435]&m[648]&~m[650]&~m[651]&m[652])|(m[435]&~m[648]&m[650]&~m[651]&m[652])|(~m[435]&~m[648]&~m[650]&m[651]&m[652])|(m[435]&~m[648]&~m[650]&m[651]&m[652])|(~m[435]&m[648]&~m[650]&m[651]&m[652])|(m[435]&m[648]&~m[650]&m[651]&m[652])|(~m[435]&~m[648]&m[650]&m[651]&m[652])|(m[435]&~m[648]&m[650]&m[651]&m[652])|(m[435]&m[648]&m[650]&m[651]&m[652]));
    m[654] = (((m[446]&~m[653]&~m[655]&~m[656]&~m[657])|(~m[446]&~m[653]&~m[655]&m[656]&~m[657])|(m[446]&m[653]&~m[655]&m[656]&~m[657])|(m[446]&~m[653]&m[655]&m[656]&~m[657])|(~m[446]&m[653]&~m[655]&~m[656]&m[657])|(~m[446]&~m[653]&m[655]&~m[656]&m[657])|(m[446]&m[653]&m[655]&~m[656]&m[657])|(~m[446]&m[653]&m[655]&m[656]&m[657]))&UnbiasedRNG[277])|((m[446]&~m[653]&~m[655]&m[656]&~m[657])|(~m[446]&~m[653]&~m[655]&~m[656]&m[657])|(m[446]&~m[653]&~m[655]&~m[656]&m[657])|(m[446]&m[653]&~m[655]&~m[656]&m[657])|(m[446]&~m[653]&m[655]&~m[656]&m[657])|(~m[446]&~m[653]&~m[655]&m[656]&m[657])|(m[446]&~m[653]&~m[655]&m[656]&m[657])|(~m[446]&m[653]&~m[655]&m[656]&m[657])|(m[446]&m[653]&~m[655]&m[656]&m[657])|(~m[446]&~m[653]&m[655]&m[656]&m[657])|(m[446]&~m[653]&m[655]&m[656]&m[657])|(m[446]&m[653]&m[655]&m[656]&m[657]));
    m[659] = (((m[457]&~m[658]&~m[660]&~m[661]&~m[662])|(~m[457]&~m[658]&~m[660]&m[661]&~m[662])|(m[457]&m[658]&~m[660]&m[661]&~m[662])|(m[457]&~m[658]&m[660]&m[661]&~m[662])|(~m[457]&m[658]&~m[660]&~m[661]&m[662])|(~m[457]&~m[658]&m[660]&~m[661]&m[662])|(m[457]&m[658]&m[660]&~m[661]&m[662])|(~m[457]&m[658]&m[660]&m[661]&m[662]))&UnbiasedRNG[278])|((m[457]&~m[658]&~m[660]&m[661]&~m[662])|(~m[457]&~m[658]&~m[660]&~m[661]&m[662])|(m[457]&~m[658]&~m[660]&~m[661]&m[662])|(m[457]&m[658]&~m[660]&~m[661]&m[662])|(m[457]&~m[658]&m[660]&~m[661]&m[662])|(~m[457]&~m[658]&~m[660]&m[661]&m[662])|(m[457]&~m[658]&~m[660]&m[661]&m[662])|(~m[457]&m[658]&~m[660]&m[661]&m[662])|(m[457]&m[658]&~m[660]&m[661]&m[662])|(~m[457]&~m[658]&m[660]&m[661]&m[662])|(m[457]&~m[658]&m[660]&m[661]&m[662])|(m[457]&m[658]&m[660]&m[661]&m[662]));
    m[664] = (((m[468]&~m[663]&~m[665]&~m[666]&~m[667])|(~m[468]&~m[663]&~m[665]&m[666]&~m[667])|(m[468]&m[663]&~m[665]&m[666]&~m[667])|(m[468]&~m[663]&m[665]&m[666]&~m[667])|(~m[468]&m[663]&~m[665]&~m[666]&m[667])|(~m[468]&~m[663]&m[665]&~m[666]&m[667])|(m[468]&m[663]&m[665]&~m[666]&m[667])|(~m[468]&m[663]&m[665]&m[666]&m[667]))&UnbiasedRNG[279])|((m[468]&~m[663]&~m[665]&m[666]&~m[667])|(~m[468]&~m[663]&~m[665]&~m[666]&m[667])|(m[468]&~m[663]&~m[665]&~m[666]&m[667])|(m[468]&m[663]&~m[665]&~m[666]&m[667])|(m[468]&~m[663]&m[665]&~m[666]&m[667])|(~m[468]&~m[663]&~m[665]&m[666]&m[667])|(m[468]&~m[663]&~m[665]&m[666]&m[667])|(~m[468]&m[663]&~m[665]&m[666]&m[667])|(m[468]&m[663]&~m[665]&m[666]&m[667])|(~m[468]&~m[663]&m[665]&m[666]&m[667])|(m[468]&~m[663]&m[665]&m[666]&m[667])|(m[468]&m[663]&m[665]&m[666]&m[667]));
    m[669] = (((m[403]&~m[668]&~m[670]&~m[671]&~m[672])|(~m[403]&~m[668]&~m[670]&m[671]&~m[672])|(m[403]&m[668]&~m[670]&m[671]&~m[672])|(m[403]&~m[668]&m[670]&m[671]&~m[672])|(~m[403]&m[668]&~m[670]&~m[671]&m[672])|(~m[403]&~m[668]&m[670]&~m[671]&m[672])|(m[403]&m[668]&m[670]&~m[671]&m[672])|(~m[403]&m[668]&m[670]&m[671]&m[672]))&UnbiasedRNG[280])|((m[403]&~m[668]&~m[670]&m[671]&~m[672])|(~m[403]&~m[668]&~m[670]&~m[671]&m[672])|(m[403]&~m[668]&~m[670]&~m[671]&m[672])|(m[403]&m[668]&~m[670]&~m[671]&m[672])|(m[403]&~m[668]&m[670]&~m[671]&m[672])|(~m[403]&~m[668]&~m[670]&m[671]&m[672])|(m[403]&~m[668]&~m[670]&m[671]&m[672])|(~m[403]&m[668]&~m[670]&m[671]&m[672])|(m[403]&m[668]&~m[670]&m[671]&m[672])|(~m[403]&~m[668]&m[670]&m[671]&m[672])|(m[403]&~m[668]&m[670]&m[671]&m[672])|(m[403]&m[668]&m[670]&m[671]&m[672]));
    m[674] = (((m[414]&~m[673]&~m[675]&~m[676]&~m[677])|(~m[414]&~m[673]&~m[675]&m[676]&~m[677])|(m[414]&m[673]&~m[675]&m[676]&~m[677])|(m[414]&~m[673]&m[675]&m[676]&~m[677])|(~m[414]&m[673]&~m[675]&~m[676]&m[677])|(~m[414]&~m[673]&m[675]&~m[676]&m[677])|(m[414]&m[673]&m[675]&~m[676]&m[677])|(~m[414]&m[673]&m[675]&m[676]&m[677]))&UnbiasedRNG[281])|((m[414]&~m[673]&~m[675]&m[676]&~m[677])|(~m[414]&~m[673]&~m[675]&~m[676]&m[677])|(m[414]&~m[673]&~m[675]&~m[676]&m[677])|(m[414]&m[673]&~m[675]&~m[676]&m[677])|(m[414]&~m[673]&m[675]&~m[676]&m[677])|(~m[414]&~m[673]&~m[675]&m[676]&m[677])|(m[414]&~m[673]&~m[675]&m[676]&m[677])|(~m[414]&m[673]&~m[675]&m[676]&m[677])|(m[414]&m[673]&~m[675]&m[676]&m[677])|(~m[414]&~m[673]&m[675]&m[676]&m[677])|(m[414]&~m[673]&m[675]&m[676]&m[677])|(m[414]&m[673]&m[675]&m[676]&m[677]));
    m[679] = (((m[425]&~m[678]&~m[680]&~m[681]&~m[682])|(~m[425]&~m[678]&~m[680]&m[681]&~m[682])|(m[425]&m[678]&~m[680]&m[681]&~m[682])|(m[425]&~m[678]&m[680]&m[681]&~m[682])|(~m[425]&m[678]&~m[680]&~m[681]&m[682])|(~m[425]&~m[678]&m[680]&~m[681]&m[682])|(m[425]&m[678]&m[680]&~m[681]&m[682])|(~m[425]&m[678]&m[680]&m[681]&m[682]))&UnbiasedRNG[282])|((m[425]&~m[678]&~m[680]&m[681]&~m[682])|(~m[425]&~m[678]&~m[680]&~m[681]&m[682])|(m[425]&~m[678]&~m[680]&~m[681]&m[682])|(m[425]&m[678]&~m[680]&~m[681]&m[682])|(m[425]&~m[678]&m[680]&~m[681]&m[682])|(~m[425]&~m[678]&~m[680]&m[681]&m[682])|(m[425]&~m[678]&~m[680]&m[681]&m[682])|(~m[425]&m[678]&~m[680]&m[681]&m[682])|(m[425]&m[678]&~m[680]&m[681]&m[682])|(~m[425]&~m[678]&m[680]&m[681]&m[682])|(m[425]&~m[678]&m[680]&m[681]&m[682])|(m[425]&m[678]&m[680]&m[681]&m[682]));
    m[684] = (((m[436]&~m[683]&~m[685]&~m[686]&~m[687])|(~m[436]&~m[683]&~m[685]&m[686]&~m[687])|(m[436]&m[683]&~m[685]&m[686]&~m[687])|(m[436]&~m[683]&m[685]&m[686]&~m[687])|(~m[436]&m[683]&~m[685]&~m[686]&m[687])|(~m[436]&~m[683]&m[685]&~m[686]&m[687])|(m[436]&m[683]&m[685]&~m[686]&m[687])|(~m[436]&m[683]&m[685]&m[686]&m[687]))&UnbiasedRNG[283])|((m[436]&~m[683]&~m[685]&m[686]&~m[687])|(~m[436]&~m[683]&~m[685]&~m[686]&m[687])|(m[436]&~m[683]&~m[685]&~m[686]&m[687])|(m[436]&m[683]&~m[685]&~m[686]&m[687])|(m[436]&~m[683]&m[685]&~m[686]&m[687])|(~m[436]&~m[683]&~m[685]&m[686]&m[687])|(m[436]&~m[683]&~m[685]&m[686]&m[687])|(~m[436]&m[683]&~m[685]&m[686]&m[687])|(m[436]&m[683]&~m[685]&m[686]&m[687])|(~m[436]&~m[683]&m[685]&m[686]&m[687])|(m[436]&~m[683]&m[685]&m[686]&m[687])|(m[436]&m[683]&m[685]&m[686]&m[687]));
    m[689] = (((m[447]&~m[688]&~m[690]&~m[691]&~m[692])|(~m[447]&~m[688]&~m[690]&m[691]&~m[692])|(m[447]&m[688]&~m[690]&m[691]&~m[692])|(m[447]&~m[688]&m[690]&m[691]&~m[692])|(~m[447]&m[688]&~m[690]&~m[691]&m[692])|(~m[447]&~m[688]&m[690]&~m[691]&m[692])|(m[447]&m[688]&m[690]&~m[691]&m[692])|(~m[447]&m[688]&m[690]&m[691]&m[692]))&UnbiasedRNG[284])|((m[447]&~m[688]&~m[690]&m[691]&~m[692])|(~m[447]&~m[688]&~m[690]&~m[691]&m[692])|(m[447]&~m[688]&~m[690]&~m[691]&m[692])|(m[447]&m[688]&~m[690]&~m[691]&m[692])|(m[447]&~m[688]&m[690]&~m[691]&m[692])|(~m[447]&~m[688]&~m[690]&m[691]&m[692])|(m[447]&~m[688]&~m[690]&m[691]&m[692])|(~m[447]&m[688]&~m[690]&m[691]&m[692])|(m[447]&m[688]&~m[690]&m[691]&m[692])|(~m[447]&~m[688]&m[690]&m[691]&m[692])|(m[447]&~m[688]&m[690]&m[691]&m[692])|(m[447]&m[688]&m[690]&m[691]&m[692]));
    m[694] = (((m[458]&~m[693]&~m[695]&~m[696]&~m[697])|(~m[458]&~m[693]&~m[695]&m[696]&~m[697])|(m[458]&m[693]&~m[695]&m[696]&~m[697])|(m[458]&~m[693]&m[695]&m[696]&~m[697])|(~m[458]&m[693]&~m[695]&~m[696]&m[697])|(~m[458]&~m[693]&m[695]&~m[696]&m[697])|(m[458]&m[693]&m[695]&~m[696]&m[697])|(~m[458]&m[693]&m[695]&m[696]&m[697]))&UnbiasedRNG[285])|((m[458]&~m[693]&~m[695]&m[696]&~m[697])|(~m[458]&~m[693]&~m[695]&~m[696]&m[697])|(m[458]&~m[693]&~m[695]&~m[696]&m[697])|(m[458]&m[693]&~m[695]&~m[696]&m[697])|(m[458]&~m[693]&m[695]&~m[696]&m[697])|(~m[458]&~m[693]&~m[695]&m[696]&m[697])|(m[458]&~m[693]&~m[695]&m[696]&m[697])|(~m[458]&m[693]&~m[695]&m[696]&m[697])|(m[458]&m[693]&~m[695]&m[696]&m[697])|(~m[458]&~m[693]&m[695]&m[696]&m[697])|(m[458]&~m[693]&m[695]&m[696]&m[697])|(m[458]&m[693]&m[695]&m[696]&m[697]));
    m[699] = (((m[469]&~m[698]&~m[700]&~m[701]&~m[702])|(~m[469]&~m[698]&~m[700]&m[701]&~m[702])|(m[469]&m[698]&~m[700]&m[701]&~m[702])|(m[469]&~m[698]&m[700]&m[701]&~m[702])|(~m[469]&m[698]&~m[700]&~m[701]&m[702])|(~m[469]&~m[698]&m[700]&~m[701]&m[702])|(m[469]&m[698]&m[700]&~m[701]&m[702])|(~m[469]&m[698]&m[700]&m[701]&m[702]))&UnbiasedRNG[286])|((m[469]&~m[698]&~m[700]&m[701]&~m[702])|(~m[469]&~m[698]&~m[700]&~m[701]&m[702])|(m[469]&~m[698]&~m[700]&~m[701]&m[702])|(m[469]&m[698]&~m[700]&~m[701]&m[702])|(m[469]&~m[698]&m[700]&~m[701]&m[702])|(~m[469]&~m[698]&~m[700]&m[701]&m[702])|(m[469]&~m[698]&~m[700]&m[701]&m[702])|(~m[469]&m[698]&~m[700]&m[701]&m[702])|(m[469]&m[698]&~m[700]&m[701]&m[702])|(~m[469]&~m[698]&m[700]&m[701]&m[702])|(m[469]&~m[698]&m[700]&m[701]&m[702])|(m[469]&m[698]&m[700]&m[701]&m[702]));
    m[704] = (((m[480]&~m[703]&~m[705]&~m[706]&~m[707])|(~m[480]&~m[703]&~m[705]&m[706]&~m[707])|(m[480]&m[703]&~m[705]&m[706]&~m[707])|(m[480]&~m[703]&m[705]&m[706]&~m[707])|(~m[480]&m[703]&~m[705]&~m[706]&m[707])|(~m[480]&~m[703]&m[705]&~m[706]&m[707])|(m[480]&m[703]&m[705]&~m[706]&m[707])|(~m[480]&m[703]&m[705]&m[706]&m[707]))&UnbiasedRNG[287])|((m[480]&~m[703]&~m[705]&m[706]&~m[707])|(~m[480]&~m[703]&~m[705]&~m[706]&m[707])|(m[480]&~m[703]&~m[705]&~m[706]&m[707])|(m[480]&m[703]&~m[705]&~m[706]&m[707])|(m[480]&~m[703]&m[705]&~m[706]&m[707])|(~m[480]&~m[703]&~m[705]&m[706]&m[707])|(m[480]&~m[703]&~m[705]&m[706]&m[707])|(~m[480]&m[703]&~m[705]&m[706]&m[707])|(m[480]&m[703]&~m[705]&m[706]&m[707])|(~m[480]&~m[703]&m[705]&m[706]&m[707])|(m[480]&~m[703]&m[705]&m[706]&m[707])|(m[480]&m[703]&m[705]&m[706]&m[707]));
    m[709] = (((m[404]&~m[708]&~m[710]&~m[711]&~m[712])|(~m[404]&~m[708]&~m[710]&m[711]&~m[712])|(m[404]&m[708]&~m[710]&m[711]&~m[712])|(m[404]&~m[708]&m[710]&m[711]&~m[712])|(~m[404]&m[708]&~m[710]&~m[711]&m[712])|(~m[404]&~m[708]&m[710]&~m[711]&m[712])|(m[404]&m[708]&m[710]&~m[711]&m[712])|(~m[404]&m[708]&m[710]&m[711]&m[712]))&UnbiasedRNG[288])|((m[404]&~m[708]&~m[710]&m[711]&~m[712])|(~m[404]&~m[708]&~m[710]&~m[711]&m[712])|(m[404]&~m[708]&~m[710]&~m[711]&m[712])|(m[404]&m[708]&~m[710]&~m[711]&m[712])|(m[404]&~m[708]&m[710]&~m[711]&m[712])|(~m[404]&~m[708]&~m[710]&m[711]&m[712])|(m[404]&~m[708]&~m[710]&m[711]&m[712])|(~m[404]&m[708]&~m[710]&m[711]&m[712])|(m[404]&m[708]&~m[710]&m[711]&m[712])|(~m[404]&~m[708]&m[710]&m[711]&m[712])|(m[404]&~m[708]&m[710]&m[711]&m[712])|(m[404]&m[708]&m[710]&m[711]&m[712]));
    m[714] = (((m[415]&~m[713]&~m[715]&~m[716]&~m[717])|(~m[415]&~m[713]&~m[715]&m[716]&~m[717])|(m[415]&m[713]&~m[715]&m[716]&~m[717])|(m[415]&~m[713]&m[715]&m[716]&~m[717])|(~m[415]&m[713]&~m[715]&~m[716]&m[717])|(~m[415]&~m[713]&m[715]&~m[716]&m[717])|(m[415]&m[713]&m[715]&~m[716]&m[717])|(~m[415]&m[713]&m[715]&m[716]&m[717]))&UnbiasedRNG[289])|((m[415]&~m[713]&~m[715]&m[716]&~m[717])|(~m[415]&~m[713]&~m[715]&~m[716]&m[717])|(m[415]&~m[713]&~m[715]&~m[716]&m[717])|(m[415]&m[713]&~m[715]&~m[716]&m[717])|(m[415]&~m[713]&m[715]&~m[716]&m[717])|(~m[415]&~m[713]&~m[715]&m[716]&m[717])|(m[415]&~m[713]&~m[715]&m[716]&m[717])|(~m[415]&m[713]&~m[715]&m[716]&m[717])|(m[415]&m[713]&~m[715]&m[716]&m[717])|(~m[415]&~m[713]&m[715]&m[716]&m[717])|(m[415]&~m[713]&m[715]&m[716]&m[717])|(m[415]&m[713]&m[715]&m[716]&m[717]));
    m[719] = (((m[426]&~m[718]&~m[720]&~m[721]&~m[722])|(~m[426]&~m[718]&~m[720]&m[721]&~m[722])|(m[426]&m[718]&~m[720]&m[721]&~m[722])|(m[426]&~m[718]&m[720]&m[721]&~m[722])|(~m[426]&m[718]&~m[720]&~m[721]&m[722])|(~m[426]&~m[718]&m[720]&~m[721]&m[722])|(m[426]&m[718]&m[720]&~m[721]&m[722])|(~m[426]&m[718]&m[720]&m[721]&m[722]))&UnbiasedRNG[290])|((m[426]&~m[718]&~m[720]&m[721]&~m[722])|(~m[426]&~m[718]&~m[720]&~m[721]&m[722])|(m[426]&~m[718]&~m[720]&~m[721]&m[722])|(m[426]&m[718]&~m[720]&~m[721]&m[722])|(m[426]&~m[718]&m[720]&~m[721]&m[722])|(~m[426]&~m[718]&~m[720]&m[721]&m[722])|(m[426]&~m[718]&~m[720]&m[721]&m[722])|(~m[426]&m[718]&~m[720]&m[721]&m[722])|(m[426]&m[718]&~m[720]&m[721]&m[722])|(~m[426]&~m[718]&m[720]&m[721]&m[722])|(m[426]&~m[718]&m[720]&m[721]&m[722])|(m[426]&m[718]&m[720]&m[721]&m[722]));
    m[724] = (((m[437]&~m[723]&~m[725]&~m[726]&~m[727])|(~m[437]&~m[723]&~m[725]&m[726]&~m[727])|(m[437]&m[723]&~m[725]&m[726]&~m[727])|(m[437]&~m[723]&m[725]&m[726]&~m[727])|(~m[437]&m[723]&~m[725]&~m[726]&m[727])|(~m[437]&~m[723]&m[725]&~m[726]&m[727])|(m[437]&m[723]&m[725]&~m[726]&m[727])|(~m[437]&m[723]&m[725]&m[726]&m[727]))&UnbiasedRNG[291])|((m[437]&~m[723]&~m[725]&m[726]&~m[727])|(~m[437]&~m[723]&~m[725]&~m[726]&m[727])|(m[437]&~m[723]&~m[725]&~m[726]&m[727])|(m[437]&m[723]&~m[725]&~m[726]&m[727])|(m[437]&~m[723]&m[725]&~m[726]&m[727])|(~m[437]&~m[723]&~m[725]&m[726]&m[727])|(m[437]&~m[723]&~m[725]&m[726]&m[727])|(~m[437]&m[723]&~m[725]&m[726]&m[727])|(m[437]&m[723]&~m[725]&m[726]&m[727])|(~m[437]&~m[723]&m[725]&m[726]&m[727])|(m[437]&~m[723]&m[725]&m[726]&m[727])|(m[437]&m[723]&m[725]&m[726]&m[727]));
    m[729] = (((m[448]&~m[728]&~m[730]&~m[731]&~m[732])|(~m[448]&~m[728]&~m[730]&m[731]&~m[732])|(m[448]&m[728]&~m[730]&m[731]&~m[732])|(m[448]&~m[728]&m[730]&m[731]&~m[732])|(~m[448]&m[728]&~m[730]&~m[731]&m[732])|(~m[448]&~m[728]&m[730]&~m[731]&m[732])|(m[448]&m[728]&m[730]&~m[731]&m[732])|(~m[448]&m[728]&m[730]&m[731]&m[732]))&UnbiasedRNG[292])|((m[448]&~m[728]&~m[730]&m[731]&~m[732])|(~m[448]&~m[728]&~m[730]&~m[731]&m[732])|(m[448]&~m[728]&~m[730]&~m[731]&m[732])|(m[448]&m[728]&~m[730]&~m[731]&m[732])|(m[448]&~m[728]&m[730]&~m[731]&m[732])|(~m[448]&~m[728]&~m[730]&m[731]&m[732])|(m[448]&~m[728]&~m[730]&m[731]&m[732])|(~m[448]&m[728]&~m[730]&m[731]&m[732])|(m[448]&m[728]&~m[730]&m[731]&m[732])|(~m[448]&~m[728]&m[730]&m[731]&m[732])|(m[448]&~m[728]&m[730]&m[731]&m[732])|(m[448]&m[728]&m[730]&m[731]&m[732]));
    m[734] = (((m[459]&~m[733]&~m[735]&~m[736]&~m[737])|(~m[459]&~m[733]&~m[735]&m[736]&~m[737])|(m[459]&m[733]&~m[735]&m[736]&~m[737])|(m[459]&~m[733]&m[735]&m[736]&~m[737])|(~m[459]&m[733]&~m[735]&~m[736]&m[737])|(~m[459]&~m[733]&m[735]&~m[736]&m[737])|(m[459]&m[733]&m[735]&~m[736]&m[737])|(~m[459]&m[733]&m[735]&m[736]&m[737]))&UnbiasedRNG[293])|((m[459]&~m[733]&~m[735]&m[736]&~m[737])|(~m[459]&~m[733]&~m[735]&~m[736]&m[737])|(m[459]&~m[733]&~m[735]&~m[736]&m[737])|(m[459]&m[733]&~m[735]&~m[736]&m[737])|(m[459]&~m[733]&m[735]&~m[736]&m[737])|(~m[459]&~m[733]&~m[735]&m[736]&m[737])|(m[459]&~m[733]&~m[735]&m[736]&m[737])|(~m[459]&m[733]&~m[735]&m[736]&m[737])|(m[459]&m[733]&~m[735]&m[736]&m[737])|(~m[459]&~m[733]&m[735]&m[736]&m[737])|(m[459]&~m[733]&m[735]&m[736]&m[737])|(m[459]&m[733]&m[735]&m[736]&m[737]));
    m[739] = (((m[470]&~m[738]&~m[740]&~m[741]&~m[742])|(~m[470]&~m[738]&~m[740]&m[741]&~m[742])|(m[470]&m[738]&~m[740]&m[741]&~m[742])|(m[470]&~m[738]&m[740]&m[741]&~m[742])|(~m[470]&m[738]&~m[740]&~m[741]&m[742])|(~m[470]&~m[738]&m[740]&~m[741]&m[742])|(m[470]&m[738]&m[740]&~m[741]&m[742])|(~m[470]&m[738]&m[740]&m[741]&m[742]))&UnbiasedRNG[294])|((m[470]&~m[738]&~m[740]&m[741]&~m[742])|(~m[470]&~m[738]&~m[740]&~m[741]&m[742])|(m[470]&~m[738]&~m[740]&~m[741]&m[742])|(m[470]&m[738]&~m[740]&~m[741]&m[742])|(m[470]&~m[738]&m[740]&~m[741]&m[742])|(~m[470]&~m[738]&~m[740]&m[741]&m[742])|(m[470]&~m[738]&~m[740]&m[741]&m[742])|(~m[470]&m[738]&~m[740]&m[741]&m[742])|(m[470]&m[738]&~m[740]&m[741]&m[742])|(~m[470]&~m[738]&m[740]&m[741]&m[742])|(m[470]&~m[738]&m[740]&m[741]&m[742])|(m[470]&m[738]&m[740]&m[741]&m[742]));
    m[744] = (((m[481]&~m[743]&~m[745]&~m[746]&~m[747])|(~m[481]&~m[743]&~m[745]&m[746]&~m[747])|(m[481]&m[743]&~m[745]&m[746]&~m[747])|(m[481]&~m[743]&m[745]&m[746]&~m[747])|(~m[481]&m[743]&~m[745]&~m[746]&m[747])|(~m[481]&~m[743]&m[745]&~m[746]&m[747])|(m[481]&m[743]&m[745]&~m[746]&m[747])|(~m[481]&m[743]&m[745]&m[746]&m[747]))&UnbiasedRNG[295])|((m[481]&~m[743]&~m[745]&m[746]&~m[747])|(~m[481]&~m[743]&~m[745]&~m[746]&m[747])|(m[481]&~m[743]&~m[745]&~m[746]&m[747])|(m[481]&m[743]&~m[745]&~m[746]&m[747])|(m[481]&~m[743]&m[745]&~m[746]&m[747])|(~m[481]&~m[743]&~m[745]&m[746]&m[747])|(m[481]&~m[743]&~m[745]&m[746]&m[747])|(~m[481]&m[743]&~m[745]&m[746]&m[747])|(m[481]&m[743]&~m[745]&m[746]&m[747])|(~m[481]&~m[743]&m[745]&m[746]&m[747])|(m[481]&~m[743]&m[745]&m[746]&m[747])|(m[481]&m[743]&m[745]&m[746]&m[747]));
    m[749] = (((m[492]&~m[748]&~m[750]&~m[751]&~m[752])|(~m[492]&~m[748]&~m[750]&m[751]&~m[752])|(m[492]&m[748]&~m[750]&m[751]&~m[752])|(m[492]&~m[748]&m[750]&m[751]&~m[752])|(~m[492]&m[748]&~m[750]&~m[751]&m[752])|(~m[492]&~m[748]&m[750]&~m[751]&m[752])|(m[492]&m[748]&m[750]&~m[751]&m[752])|(~m[492]&m[748]&m[750]&m[751]&m[752]))&UnbiasedRNG[296])|((m[492]&~m[748]&~m[750]&m[751]&~m[752])|(~m[492]&~m[748]&~m[750]&~m[751]&m[752])|(m[492]&~m[748]&~m[750]&~m[751]&m[752])|(m[492]&m[748]&~m[750]&~m[751]&m[752])|(m[492]&~m[748]&m[750]&~m[751]&m[752])|(~m[492]&~m[748]&~m[750]&m[751]&m[752])|(m[492]&~m[748]&~m[750]&m[751]&m[752])|(~m[492]&m[748]&~m[750]&m[751]&m[752])|(m[492]&m[748]&~m[750]&m[751]&m[752])|(~m[492]&~m[748]&m[750]&m[751]&m[752])|(m[492]&~m[748]&m[750]&m[751]&m[752])|(m[492]&m[748]&m[750]&m[751]&m[752]));
    m[754] = (((m[405]&~m[753]&~m[755]&~m[756]&~m[757])|(~m[405]&~m[753]&~m[755]&m[756]&~m[757])|(m[405]&m[753]&~m[755]&m[756]&~m[757])|(m[405]&~m[753]&m[755]&m[756]&~m[757])|(~m[405]&m[753]&~m[755]&~m[756]&m[757])|(~m[405]&~m[753]&m[755]&~m[756]&m[757])|(m[405]&m[753]&m[755]&~m[756]&m[757])|(~m[405]&m[753]&m[755]&m[756]&m[757]))&UnbiasedRNG[297])|((m[405]&~m[753]&~m[755]&m[756]&~m[757])|(~m[405]&~m[753]&~m[755]&~m[756]&m[757])|(m[405]&~m[753]&~m[755]&~m[756]&m[757])|(m[405]&m[753]&~m[755]&~m[756]&m[757])|(m[405]&~m[753]&m[755]&~m[756]&m[757])|(~m[405]&~m[753]&~m[755]&m[756]&m[757])|(m[405]&~m[753]&~m[755]&m[756]&m[757])|(~m[405]&m[753]&~m[755]&m[756]&m[757])|(m[405]&m[753]&~m[755]&m[756]&m[757])|(~m[405]&~m[753]&m[755]&m[756]&m[757])|(m[405]&~m[753]&m[755]&m[756]&m[757])|(m[405]&m[753]&m[755]&m[756]&m[757]));
    m[759] = (((m[416]&~m[758]&~m[760]&~m[761]&~m[762])|(~m[416]&~m[758]&~m[760]&m[761]&~m[762])|(m[416]&m[758]&~m[760]&m[761]&~m[762])|(m[416]&~m[758]&m[760]&m[761]&~m[762])|(~m[416]&m[758]&~m[760]&~m[761]&m[762])|(~m[416]&~m[758]&m[760]&~m[761]&m[762])|(m[416]&m[758]&m[760]&~m[761]&m[762])|(~m[416]&m[758]&m[760]&m[761]&m[762]))&UnbiasedRNG[298])|((m[416]&~m[758]&~m[760]&m[761]&~m[762])|(~m[416]&~m[758]&~m[760]&~m[761]&m[762])|(m[416]&~m[758]&~m[760]&~m[761]&m[762])|(m[416]&m[758]&~m[760]&~m[761]&m[762])|(m[416]&~m[758]&m[760]&~m[761]&m[762])|(~m[416]&~m[758]&~m[760]&m[761]&m[762])|(m[416]&~m[758]&~m[760]&m[761]&m[762])|(~m[416]&m[758]&~m[760]&m[761]&m[762])|(m[416]&m[758]&~m[760]&m[761]&m[762])|(~m[416]&~m[758]&m[760]&m[761]&m[762])|(m[416]&~m[758]&m[760]&m[761]&m[762])|(m[416]&m[758]&m[760]&m[761]&m[762]));
    m[764] = (((m[427]&~m[763]&~m[765]&~m[766]&~m[767])|(~m[427]&~m[763]&~m[765]&m[766]&~m[767])|(m[427]&m[763]&~m[765]&m[766]&~m[767])|(m[427]&~m[763]&m[765]&m[766]&~m[767])|(~m[427]&m[763]&~m[765]&~m[766]&m[767])|(~m[427]&~m[763]&m[765]&~m[766]&m[767])|(m[427]&m[763]&m[765]&~m[766]&m[767])|(~m[427]&m[763]&m[765]&m[766]&m[767]))&UnbiasedRNG[299])|((m[427]&~m[763]&~m[765]&m[766]&~m[767])|(~m[427]&~m[763]&~m[765]&~m[766]&m[767])|(m[427]&~m[763]&~m[765]&~m[766]&m[767])|(m[427]&m[763]&~m[765]&~m[766]&m[767])|(m[427]&~m[763]&m[765]&~m[766]&m[767])|(~m[427]&~m[763]&~m[765]&m[766]&m[767])|(m[427]&~m[763]&~m[765]&m[766]&m[767])|(~m[427]&m[763]&~m[765]&m[766]&m[767])|(m[427]&m[763]&~m[765]&m[766]&m[767])|(~m[427]&~m[763]&m[765]&m[766]&m[767])|(m[427]&~m[763]&m[765]&m[766]&m[767])|(m[427]&m[763]&m[765]&m[766]&m[767]));
    m[769] = (((m[438]&~m[768]&~m[770]&~m[771]&~m[772])|(~m[438]&~m[768]&~m[770]&m[771]&~m[772])|(m[438]&m[768]&~m[770]&m[771]&~m[772])|(m[438]&~m[768]&m[770]&m[771]&~m[772])|(~m[438]&m[768]&~m[770]&~m[771]&m[772])|(~m[438]&~m[768]&m[770]&~m[771]&m[772])|(m[438]&m[768]&m[770]&~m[771]&m[772])|(~m[438]&m[768]&m[770]&m[771]&m[772]))&UnbiasedRNG[300])|((m[438]&~m[768]&~m[770]&m[771]&~m[772])|(~m[438]&~m[768]&~m[770]&~m[771]&m[772])|(m[438]&~m[768]&~m[770]&~m[771]&m[772])|(m[438]&m[768]&~m[770]&~m[771]&m[772])|(m[438]&~m[768]&m[770]&~m[771]&m[772])|(~m[438]&~m[768]&~m[770]&m[771]&m[772])|(m[438]&~m[768]&~m[770]&m[771]&m[772])|(~m[438]&m[768]&~m[770]&m[771]&m[772])|(m[438]&m[768]&~m[770]&m[771]&m[772])|(~m[438]&~m[768]&m[770]&m[771]&m[772])|(m[438]&~m[768]&m[770]&m[771]&m[772])|(m[438]&m[768]&m[770]&m[771]&m[772]));
    m[774] = (((m[449]&~m[773]&~m[775]&~m[776]&~m[777])|(~m[449]&~m[773]&~m[775]&m[776]&~m[777])|(m[449]&m[773]&~m[775]&m[776]&~m[777])|(m[449]&~m[773]&m[775]&m[776]&~m[777])|(~m[449]&m[773]&~m[775]&~m[776]&m[777])|(~m[449]&~m[773]&m[775]&~m[776]&m[777])|(m[449]&m[773]&m[775]&~m[776]&m[777])|(~m[449]&m[773]&m[775]&m[776]&m[777]))&UnbiasedRNG[301])|((m[449]&~m[773]&~m[775]&m[776]&~m[777])|(~m[449]&~m[773]&~m[775]&~m[776]&m[777])|(m[449]&~m[773]&~m[775]&~m[776]&m[777])|(m[449]&m[773]&~m[775]&~m[776]&m[777])|(m[449]&~m[773]&m[775]&~m[776]&m[777])|(~m[449]&~m[773]&~m[775]&m[776]&m[777])|(m[449]&~m[773]&~m[775]&m[776]&m[777])|(~m[449]&m[773]&~m[775]&m[776]&m[777])|(m[449]&m[773]&~m[775]&m[776]&m[777])|(~m[449]&~m[773]&m[775]&m[776]&m[777])|(m[449]&~m[773]&m[775]&m[776]&m[777])|(m[449]&m[773]&m[775]&m[776]&m[777]));
    m[779] = (((m[460]&~m[778]&~m[780]&~m[781]&~m[782])|(~m[460]&~m[778]&~m[780]&m[781]&~m[782])|(m[460]&m[778]&~m[780]&m[781]&~m[782])|(m[460]&~m[778]&m[780]&m[781]&~m[782])|(~m[460]&m[778]&~m[780]&~m[781]&m[782])|(~m[460]&~m[778]&m[780]&~m[781]&m[782])|(m[460]&m[778]&m[780]&~m[781]&m[782])|(~m[460]&m[778]&m[780]&m[781]&m[782]))&UnbiasedRNG[302])|((m[460]&~m[778]&~m[780]&m[781]&~m[782])|(~m[460]&~m[778]&~m[780]&~m[781]&m[782])|(m[460]&~m[778]&~m[780]&~m[781]&m[782])|(m[460]&m[778]&~m[780]&~m[781]&m[782])|(m[460]&~m[778]&m[780]&~m[781]&m[782])|(~m[460]&~m[778]&~m[780]&m[781]&m[782])|(m[460]&~m[778]&~m[780]&m[781]&m[782])|(~m[460]&m[778]&~m[780]&m[781]&m[782])|(m[460]&m[778]&~m[780]&m[781]&m[782])|(~m[460]&~m[778]&m[780]&m[781]&m[782])|(m[460]&~m[778]&m[780]&m[781]&m[782])|(m[460]&m[778]&m[780]&m[781]&m[782]));
    m[784] = (((m[471]&~m[783]&~m[785]&~m[786]&~m[787])|(~m[471]&~m[783]&~m[785]&m[786]&~m[787])|(m[471]&m[783]&~m[785]&m[786]&~m[787])|(m[471]&~m[783]&m[785]&m[786]&~m[787])|(~m[471]&m[783]&~m[785]&~m[786]&m[787])|(~m[471]&~m[783]&m[785]&~m[786]&m[787])|(m[471]&m[783]&m[785]&~m[786]&m[787])|(~m[471]&m[783]&m[785]&m[786]&m[787]))&UnbiasedRNG[303])|((m[471]&~m[783]&~m[785]&m[786]&~m[787])|(~m[471]&~m[783]&~m[785]&~m[786]&m[787])|(m[471]&~m[783]&~m[785]&~m[786]&m[787])|(m[471]&m[783]&~m[785]&~m[786]&m[787])|(m[471]&~m[783]&m[785]&~m[786]&m[787])|(~m[471]&~m[783]&~m[785]&m[786]&m[787])|(m[471]&~m[783]&~m[785]&m[786]&m[787])|(~m[471]&m[783]&~m[785]&m[786]&m[787])|(m[471]&m[783]&~m[785]&m[786]&m[787])|(~m[471]&~m[783]&m[785]&m[786]&m[787])|(m[471]&~m[783]&m[785]&m[786]&m[787])|(m[471]&m[783]&m[785]&m[786]&m[787]));
    m[789] = (((m[482]&~m[788]&~m[790]&~m[791]&~m[792])|(~m[482]&~m[788]&~m[790]&m[791]&~m[792])|(m[482]&m[788]&~m[790]&m[791]&~m[792])|(m[482]&~m[788]&m[790]&m[791]&~m[792])|(~m[482]&m[788]&~m[790]&~m[791]&m[792])|(~m[482]&~m[788]&m[790]&~m[791]&m[792])|(m[482]&m[788]&m[790]&~m[791]&m[792])|(~m[482]&m[788]&m[790]&m[791]&m[792]))&UnbiasedRNG[304])|((m[482]&~m[788]&~m[790]&m[791]&~m[792])|(~m[482]&~m[788]&~m[790]&~m[791]&m[792])|(m[482]&~m[788]&~m[790]&~m[791]&m[792])|(m[482]&m[788]&~m[790]&~m[791]&m[792])|(m[482]&~m[788]&m[790]&~m[791]&m[792])|(~m[482]&~m[788]&~m[790]&m[791]&m[792])|(m[482]&~m[788]&~m[790]&m[791]&m[792])|(~m[482]&m[788]&~m[790]&m[791]&m[792])|(m[482]&m[788]&~m[790]&m[791]&m[792])|(~m[482]&~m[788]&m[790]&m[791]&m[792])|(m[482]&~m[788]&m[790]&m[791]&m[792])|(m[482]&m[788]&m[790]&m[791]&m[792]));
    m[794] = (((m[493]&~m[793]&~m[795]&~m[796]&~m[797])|(~m[493]&~m[793]&~m[795]&m[796]&~m[797])|(m[493]&m[793]&~m[795]&m[796]&~m[797])|(m[493]&~m[793]&m[795]&m[796]&~m[797])|(~m[493]&m[793]&~m[795]&~m[796]&m[797])|(~m[493]&~m[793]&m[795]&~m[796]&m[797])|(m[493]&m[793]&m[795]&~m[796]&m[797])|(~m[493]&m[793]&m[795]&m[796]&m[797]))&UnbiasedRNG[305])|((m[493]&~m[793]&~m[795]&m[796]&~m[797])|(~m[493]&~m[793]&~m[795]&~m[796]&m[797])|(m[493]&~m[793]&~m[795]&~m[796]&m[797])|(m[493]&m[793]&~m[795]&~m[796]&m[797])|(m[493]&~m[793]&m[795]&~m[796]&m[797])|(~m[493]&~m[793]&~m[795]&m[796]&m[797])|(m[493]&~m[793]&~m[795]&m[796]&m[797])|(~m[493]&m[793]&~m[795]&m[796]&m[797])|(m[493]&m[793]&~m[795]&m[796]&m[797])|(~m[493]&~m[793]&m[795]&m[796]&m[797])|(m[493]&~m[793]&m[795]&m[796]&m[797])|(m[493]&m[793]&m[795]&m[796]&m[797]));
    m[799] = (((m[504]&~m[798]&~m[800]&~m[801]&~m[802])|(~m[504]&~m[798]&~m[800]&m[801]&~m[802])|(m[504]&m[798]&~m[800]&m[801]&~m[802])|(m[504]&~m[798]&m[800]&m[801]&~m[802])|(~m[504]&m[798]&~m[800]&~m[801]&m[802])|(~m[504]&~m[798]&m[800]&~m[801]&m[802])|(m[504]&m[798]&m[800]&~m[801]&m[802])|(~m[504]&m[798]&m[800]&m[801]&m[802]))&UnbiasedRNG[306])|((m[504]&~m[798]&~m[800]&m[801]&~m[802])|(~m[504]&~m[798]&~m[800]&~m[801]&m[802])|(m[504]&~m[798]&~m[800]&~m[801]&m[802])|(m[504]&m[798]&~m[800]&~m[801]&m[802])|(m[504]&~m[798]&m[800]&~m[801]&m[802])|(~m[504]&~m[798]&~m[800]&m[801]&m[802])|(m[504]&~m[798]&~m[800]&m[801]&m[802])|(~m[504]&m[798]&~m[800]&m[801]&m[802])|(m[504]&m[798]&~m[800]&m[801]&m[802])|(~m[504]&~m[798]&m[800]&m[801]&m[802])|(m[504]&~m[798]&m[800]&m[801]&m[802])|(m[504]&m[798]&m[800]&m[801]&m[802]));
    m[804] = (((m[406]&~m[803]&~m[805]&~m[806]&~m[807])|(~m[406]&~m[803]&~m[805]&m[806]&~m[807])|(m[406]&m[803]&~m[805]&m[806]&~m[807])|(m[406]&~m[803]&m[805]&m[806]&~m[807])|(~m[406]&m[803]&~m[805]&~m[806]&m[807])|(~m[406]&~m[803]&m[805]&~m[806]&m[807])|(m[406]&m[803]&m[805]&~m[806]&m[807])|(~m[406]&m[803]&m[805]&m[806]&m[807]))&UnbiasedRNG[307])|((m[406]&~m[803]&~m[805]&m[806]&~m[807])|(~m[406]&~m[803]&~m[805]&~m[806]&m[807])|(m[406]&~m[803]&~m[805]&~m[806]&m[807])|(m[406]&m[803]&~m[805]&~m[806]&m[807])|(m[406]&~m[803]&m[805]&~m[806]&m[807])|(~m[406]&~m[803]&~m[805]&m[806]&m[807])|(m[406]&~m[803]&~m[805]&m[806]&m[807])|(~m[406]&m[803]&~m[805]&m[806]&m[807])|(m[406]&m[803]&~m[805]&m[806]&m[807])|(~m[406]&~m[803]&m[805]&m[806]&m[807])|(m[406]&~m[803]&m[805]&m[806]&m[807])|(m[406]&m[803]&m[805]&m[806]&m[807]));
    m[809] = (((m[417]&~m[808]&~m[810]&~m[811]&~m[812])|(~m[417]&~m[808]&~m[810]&m[811]&~m[812])|(m[417]&m[808]&~m[810]&m[811]&~m[812])|(m[417]&~m[808]&m[810]&m[811]&~m[812])|(~m[417]&m[808]&~m[810]&~m[811]&m[812])|(~m[417]&~m[808]&m[810]&~m[811]&m[812])|(m[417]&m[808]&m[810]&~m[811]&m[812])|(~m[417]&m[808]&m[810]&m[811]&m[812]))&UnbiasedRNG[308])|((m[417]&~m[808]&~m[810]&m[811]&~m[812])|(~m[417]&~m[808]&~m[810]&~m[811]&m[812])|(m[417]&~m[808]&~m[810]&~m[811]&m[812])|(m[417]&m[808]&~m[810]&~m[811]&m[812])|(m[417]&~m[808]&m[810]&~m[811]&m[812])|(~m[417]&~m[808]&~m[810]&m[811]&m[812])|(m[417]&~m[808]&~m[810]&m[811]&m[812])|(~m[417]&m[808]&~m[810]&m[811]&m[812])|(m[417]&m[808]&~m[810]&m[811]&m[812])|(~m[417]&~m[808]&m[810]&m[811]&m[812])|(m[417]&~m[808]&m[810]&m[811]&m[812])|(m[417]&m[808]&m[810]&m[811]&m[812]));
    m[814] = (((m[428]&~m[813]&~m[815]&~m[816]&~m[817])|(~m[428]&~m[813]&~m[815]&m[816]&~m[817])|(m[428]&m[813]&~m[815]&m[816]&~m[817])|(m[428]&~m[813]&m[815]&m[816]&~m[817])|(~m[428]&m[813]&~m[815]&~m[816]&m[817])|(~m[428]&~m[813]&m[815]&~m[816]&m[817])|(m[428]&m[813]&m[815]&~m[816]&m[817])|(~m[428]&m[813]&m[815]&m[816]&m[817]))&UnbiasedRNG[309])|((m[428]&~m[813]&~m[815]&m[816]&~m[817])|(~m[428]&~m[813]&~m[815]&~m[816]&m[817])|(m[428]&~m[813]&~m[815]&~m[816]&m[817])|(m[428]&m[813]&~m[815]&~m[816]&m[817])|(m[428]&~m[813]&m[815]&~m[816]&m[817])|(~m[428]&~m[813]&~m[815]&m[816]&m[817])|(m[428]&~m[813]&~m[815]&m[816]&m[817])|(~m[428]&m[813]&~m[815]&m[816]&m[817])|(m[428]&m[813]&~m[815]&m[816]&m[817])|(~m[428]&~m[813]&m[815]&m[816]&m[817])|(m[428]&~m[813]&m[815]&m[816]&m[817])|(m[428]&m[813]&m[815]&m[816]&m[817]));
    m[819] = (((m[439]&~m[818]&~m[820]&~m[821]&~m[822])|(~m[439]&~m[818]&~m[820]&m[821]&~m[822])|(m[439]&m[818]&~m[820]&m[821]&~m[822])|(m[439]&~m[818]&m[820]&m[821]&~m[822])|(~m[439]&m[818]&~m[820]&~m[821]&m[822])|(~m[439]&~m[818]&m[820]&~m[821]&m[822])|(m[439]&m[818]&m[820]&~m[821]&m[822])|(~m[439]&m[818]&m[820]&m[821]&m[822]))&UnbiasedRNG[310])|((m[439]&~m[818]&~m[820]&m[821]&~m[822])|(~m[439]&~m[818]&~m[820]&~m[821]&m[822])|(m[439]&~m[818]&~m[820]&~m[821]&m[822])|(m[439]&m[818]&~m[820]&~m[821]&m[822])|(m[439]&~m[818]&m[820]&~m[821]&m[822])|(~m[439]&~m[818]&~m[820]&m[821]&m[822])|(m[439]&~m[818]&~m[820]&m[821]&m[822])|(~m[439]&m[818]&~m[820]&m[821]&m[822])|(m[439]&m[818]&~m[820]&m[821]&m[822])|(~m[439]&~m[818]&m[820]&m[821]&m[822])|(m[439]&~m[818]&m[820]&m[821]&m[822])|(m[439]&m[818]&m[820]&m[821]&m[822]));
    m[824] = (((m[450]&~m[823]&~m[825]&~m[826]&~m[827])|(~m[450]&~m[823]&~m[825]&m[826]&~m[827])|(m[450]&m[823]&~m[825]&m[826]&~m[827])|(m[450]&~m[823]&m[825]&m[826]&~m[827])|(~m[450]&m[823]&~m[825]&~m[826]&m[827])|(~m[450]&~m[823]&m[825]&~m[826]&m[827])|(m[450]&m[823]&m[825]&~m[826]&m[827])|(~m[450]&m[823]&m[825]&m[826]&m[827]))&UnbiasedRNG[311])|((m[450]&~m[823]&~m[825]&m[826]&~m[827])|(~m[450]&~m[823]&~m[825]&~m[826]&m[827])|(m[450]&~m[823]&~m[825]&~m[826]&m[827])|(m[450]&m[823]&~m[825]&~m[826]&m[827])|(m[450]&~m[823]&m[825]&~m[826]&m[827])|(~m[450]&~m[823]&~m[825]&m[826]&m[827])|(m[450]&~m[823]&~m[825]&m[826]&m[827])|(~m[450]&m[823]&~m[825]&m[826]&m[827])|(m[450]&m[823]&~m[825]&m[826]&m[827])|(~m[450]&~m[823]&m[825]&m[826]&m[827])|(m[450]&~m[823]&m[825]&m[826]&m[827])|(m[450]&m[823]&m[825]&m[826]&m[827]));
    m[829] = (((m[461]&~m[828]&~m[830]&~m[831]&~m[832])|(~m[461]&~m[828]&~m[830]&m[831]&~m[832])|(m[461]&m[828]&~m[830]&m[831]&~m[832])|(m[461]&~m[828]&m[830]&m[831]&~m[832])|(~m[461]&m[828]&~m[830]&~m[831]&m[832])|(~m[461]&~m[828]&m[830]&~m[831]&m[832])|(m[461]&m[828]&m[830]&~m[831]&m[832])|(~m[461]&m[828]&m[830]&m[831]&m[832]))&UnbiasedRNG[312])|((m[461]&~m[828]&~m[830]&m[831]&~m[832])|(~m[461]&~m[828]&~m[830]&~m[831]&m[832])|(m[461]&~m[828]&~m[830]&~m[831]&m[832])|(m[461]&m[828]&~m[830]&~m[831]&m[832])|(m[461]&~m[828]&m[830]&~m[831]&m[832])|(~m[461]&~m[828]&~m[830]&m[831]&m[832])|(m[461]&~m[828]&~m[830]&m[831]&m[832])|(~m[461]&m[828]&~m[830]&m[831]&m[832])|(m[461]&m[828]&~m[830]&m[831]&m[832])|(~m[461]&~m[828]&m[830]&m[831]&m[832])|(m[461]&~m[828]&m[830]&m[831]&m[832])|(m[461]&m[828]&m[830]&m[831]&m[832]));
    m[834] = (((m[472]&~m[833]&~m[835]&~m[836]&~m[837])|(~m[472]&~m[833]&~m[835]&m[836]&~m[837])|(m[472]&m[833]&~m[835]&m[836]&~m[837])|(m[472]&~m[833]&m[835]&m[836]&~m[837])|(~m[472]&m[833]&~m[835]&~m[836]&m[837])|(~m[472]&~m[833]&m[835]&~m[836]&m[837])|(m[472]&m[833]&m[835]&~m[836]&m[837])|(~m[472]&m[833]&m[835]&m[836]&m[837]))&UnbiasedRNG[313])|((m[472]&~m[833]&~m[835]&m[836]&~m[837])|(~m[472]&~m[833]&~m[835]&~m[836]&m[837])|(m[472]&~m[833]&~m[835]&~m[836]&m[837])|(m[472]&m[833]&~m[835]&~m[836]&m[837])|(m[472]&~m[833]&m[835]&~m[836]&m[837])|(~m[472]&~m[833]&~m[835]&m[836]&m[837])|(m[472]&~m[833]&~m[835]&m[836]&m[837])|(~m[472]&m[833]&~m[835]&m[836]&m[837])|(m[472]&m[833]&~m[835]&m[836]&m[837])|(~m[472]&~m[833]&m[835]&m[836]&m[837])|(m[472]&~m[833]&m[835]&m[836]&m[837])|(m[472]&m[833]&m[835]&m[836]&m[837]));
    m[839] = (((m[483]&~m[838]&~m[840]&~m[841]&~m[842])|(~m[483]&~m[838]&~m[840]&m[841]&~m[842])|(m[483]&m[838]&~m[840]&m[841]&~m[842])|(m[483]&~m[838]&m[840]&m[841]&~m[842])|(~m[483]&m[838]&~m[840]&~m[841]&m[842])|(~m[483]&~m[838]&m[840]&~m[841]&m[842])|(m[483]&m[838]&m[840]&~m[841]&m[842])|(~m[483]&m[838]&m[840]&m[841]&m[842]))&UnbiasedRNG[314])|((m[483]&~m[838]&~m[840]&m[841]&~m[842])|(~m[483]&~m[838]&~m[840]&~m[841]&m[842])|(m[483]&~m[838]&~m[840]&~m[841]&m[842])|(m[483]&m[838]&~m[840]&~m[841]&m[842])|(m[483]&~m[838]&m[840]&~m[841]&m[842])|(~m[483]&~m[838]&~m[840]&m[841]&m[842])|(m[483]&~m[838]&~m[840]&m[841]&m[842])|(~m[483]&m[838]&~m[840]&m[841]&m[842])|(m[483]&m[838]&~m[840]&m[841]&m[842])|(~m[483]&~m[838]&m[840]&m[841]&m[842])|(m[483]&~m[838]&m[840]&m[841]&m[842])|(m[483]&m[838]&m[840]&m[841]&m[842]));
    m[844] = (((m[494]&~m[843]&~m[845]&~m[846]&~m[847])|(~m[494]&~m[843]&~m[845]&m[846]&~m[847])|(m[494]&m[843]&~m[845]&m[846]&~m[847])|(m[494]&~m[843]&m[845]&m[846]&~m[847])|(~m[494]&m[843]&~m[845]&~m[846]&m[847])|(~m[494]&~m[843]&m[845]&~m[846]&m[847])|(m[494]&m[843]&m[845]&~m[846]&m[847])|(~m[494]&m[843]&m[845]&m[846]&m[847]))&UnbiasedRNG[315])|((m[494]&~m[843]&~m[845]&m[846]&~m[847])|(~m[494]&~m[843]&~m[845]&~m[846]&m[847])|(m[494]&~m[843]&~m[845]&~m[846]&m[847])|(m[494]&m[843]&~m[845]&~m[846]&m[847])|(m[494]&~m[843]&m[845]&~m[846]&m[847])|(~m[494]&~m[843]&~m[845]&m[846]&m[847])|(m[494]&~m[843]&~m[845]&m[846]&m[847])|(~m[494]&m[843]&~m[845]&m[846]&m[847])|(m[494]&m[843]&~m[845]&m[846]&m[847])|(~m[494]&~m[843]&m[845]&m[846]&m[847])|(m[494]&~m[843]&m[845]&m[846]&m[847])|(m[494]&m[843]&m[845]&m[846]&m[847]));
    m[849] = (((m[505]&~m[848]&~m[850]&~m[851]&~m[852])|(~m[505]&~m[848]&~m[850]&m[851]&~m[852])|(m[505]&m[848]&~m[850]&m[851]&~m[852])|(m[505]&~m[848]&m[850]&m[851]&~m[852])|(~m[505]&m[848]&~m[850]&~m[851]&m[852])|(~m[505]&~m[848]&m[850]&~m[851]&m[852])|(m[505]&m[848]&m[850]&~m[851]&m[852])|(~m[505]&m[848]&m[850]&m[851]&m[852]))&UnbiasedRNG[316])|((m[505]&~m[848]&~m[850]&m[851]&~m[852])|(~m[505]&~m[848]&~m[850]&~m[851]&m[852])|(m[505]&~m[848]&~m[850]&~m[851]&m[852])|(m[505]&m[848]&~m[850]&~m[851]&m[852])|(m[505]&~m[848]&m[850]&~m[851]&m[852])|(~m[505]&~m[848]&~m[850]&m[851]&m[852])|(m[505]&~m[848]&~m[850]&m[851]&m[852])|(~m[505]&m[848]&~m[850]&m[851]&m[852])|(m[505]&m[848]&~m[850]&m[851]&m[852])|(~m[505]&~m[848]&m[850]&m[851]&m[852])|(m[505]&~m[848]&m[850]&m[851]&m[852])|(m[505]&m[848]&m[850]&m[851]&m[852]));
    m[854] = (((m[516]&~m[853]&~m[855]&~m[856]&~m[857])|(~m[516]&~m[853]&~m[855]&m[856]&~m[857])|(m[516]&m[853]&~m[855]&m[856]&~m[857])|(m[516]&~m[853]&m[855]&m[856]&~m[857])|(~m[516]&m[853]&~m[855]&~m[856]&m[857])|(~m[516]&~m[853]&m[855]&~m[856]&m[857])|(m[516]&m[853]&m[855]&~m[856]&m[857])|(~m[516]&m[853]&m[855]&m[856]&m[857]))&UnbiasedRNG[317])|((m[516]&~m[853]&~m[855]&m[856]&~m[857])|(~m[516]&~m[853]&~m[855]&~m[856]&m[857])|(m[516]&~m[853]&~m[855]&~m[856]&m[857])|(m[516]&m[853]&~m[855]&~m[856]&m[857])|(m[516]&~m[853]&m[855]&~m[856]&m[857])|(~m[516]&~m[853]&~m[855]&m[856]&m[857])|(m[516]&~m[853]&~m[855]&m[856]&m[857])|(~m[516]&m[853]&~m[855]&m[856]&m[857])|(m[516]&m[853]&~m[855]&m[856]&m[857])|(~m[516]&~m[853]&m[855]&m[856]&m[857])|(m[516]&~m[853]&m[855]&m[856]&m[857])|(m[516]&m[853]&m[855]&m[856]&m[857]));
    m[859] = (((m[407]&~m[858]&~m[860]&~m[861]&~m[862])|(~m[407]&~m[858]&~m[860]&m[861]&~m[862])|(m[407]&m[858]&~m[860]&m[861]&~m[862])|(m[407]&~m[858]&m[860]&m[861]&~m[862])|(~m[407]&m[858]&~m[860]&~m[861]&m[862])|(~m[407]&~m[858]&m[860]&~m[861]&m[862])|(m[407]&m[858]&m[860]&~m[861]&m[862])|(~m[407]&m[858]&m[860]&m[861]&m[862]))&UnbiasedRNG[318])|((m[407]&~m[858]&~m[860]&m[861]&~m[862])|(~m[407]&~m[858]&~m[860]&~m[861]&m[862])|(m[407]&~m[858]&~m[860]&~m[861]&m[862])|(m[407]&m[858]&~m[860]&~m[861]&m[862])|(m[407]&~m[858]&m[860]&~m[861]&m[862])|(~m[407]&~m[858]&~m[860]&m[861]&m[862])|(m[407]&~m[858]&~m[860]&m[861]&m[862])|(~m[407]&m[858]&~m[860]&m[861]&m[862])|(m[407]&m[858]&~m[860]&m[861]&m[862])|(~m[407]&~m[858]&m[860]&m[861]&m[862])|(m[407]&~m[858]&m[860]&m[861]&m[862])|(m[407]&m[858]&m[860]&m[861]&m[862]));
    m[864] = (((m[418]&~m[863]&~m[865]&~m[866]&~m[867])|(~m[418]&~m[863]&~m[865]&m[866]&~m[867])|(m[418]&m[863]&~m[865]&m[866]&~m[867])|(m[418]&~m[863]&m[865]&m[866]&~m[867])|(~m[418]&m[863]&~m[865]&~m[866]&m[867])|(~m[418]&~m[863]&m[865]&~m[866]&m[867])|(m[418]&m[863]&m[865]&~m[866]&m[867])|(~m[418]&m[863]&m[865]&m[866]&m[867]))&UnbiasedRNG[319])|((m[418]&~m[863]&~m[865]&m[866]&~m[867])|(~m[418]&~m[863]&~m[865]&~m[866]&m[867])|(m[418]&~m[863]&~m[865]&~m[866]&m[867])|(m[418]&m[863]&~m[865]&~m[866]&m[867])|(m[418]&~m[863]&m[865]&~m[866]&m[867])|(~m[418]&~m[863]&~m[865]&m[866]&m[867])|(m[418]&~m[863]&~m[865]&m[866]&m[867])|(~m[418]&m[863]&~m[865]&m[866]&m[867])|(m[418]&m[863]&~m[865]&m[866]&m[867])|(~m[418]&~m[863]&m[865]&m[866]&m[867])|(m[418]&~m[863]&m[865]&m[866]&m[867])|(m[418]&m[863]&m[865]&m[866]&m[867]));
    m[869] = (((m[429]&~m[868]&~m[870]&~m[871]&~m[872])|(~m[429]&~m[868]&~m[870]&m[871]&~m[872])|(m[429]&m[868]&~m[870]&m[871]&~m[872])|(m[429]&~m[868]&m[870]&m[871]&~m[872])|(~m[429]&m[868]&~m[870]&~m[871]&m[872])|(~m[429]&~m[868]&m[870]&~m[871]&m[872])|(m[429]&m[868]&m[870]&~m[871]&m[872])|(~m[429]&m[868]&m[870]&m[871]&m[872]))&UnbiasedRNG[320])|((m[429]&~m[868]&~m[870]&m[871]&~m[872])|(~m[429]&~m[868]&~m[870]&~m[871]&m[872])|(m[429]&~m[868]&~m[870]&~m[871]&m[872])|(m[429]&m[868]&~m[870]&~m[871]&m[872])|(m[429]&~m[868]&m[870]&~m[871]&m[872])|(~m[429]&~m[868]&~m[870]&m[871]&m[872])|(m[429]&~m[868]&~m[870]&m[871]&m[872])|(~m[429]&m[868]&~m[870]&m[871]&m[872])|(m[429]&m[868]&~m[870]&m[871]&m[872])|(~m[429]&~m[868]&m[870]&m[871]&m[872])|(m[429]&~m[868]&m[870]&m[871]&m[872])|(m[429]&m[868]&m[870]&m[871]&m[872]));
    m[874] = (((m[440]&~m[873]&~m[875]&~m[876]&~m[877])|(~m[440]&~m[873]&~m[875]&m[876]&~m[877])|(m[440]&m[873]&~m[875]&m[876]&~m[877])|(m[440]&~m[873]&m[875]&m[876]&~m[877])|(~m[440]&m[873]&~m[875]&~m[876]&m[877])|(~m[440]&~m[873]&m[875]&~m[876]&m[877])|(m[440]&m[873]&m[875]&~m[876]&m[877])|(~m[440]&m[873]&m[875]&m[876]&m[877]))&UnbiasedRNG[321])|((m[440]&~m[873]&~m[875]&m[876]&~m[877])|(~m[440]&~m[873]&~m[875]&~m[876]&m[877])|(m[440]&~m[873]&~m[875]&~m[876]&m[877])|(m[440]&m[873]&~m[875]&~m[876]&m[877])|(m[440]&~m[873]&m[875]&~m[876]&m[877])|(~m[440]&~m[873]&~m[875]&m[876]&m[877])|(m[440]&~m[873]&~m[875]&m[876]&m[877])|(~m[440]&m[873]&~m[875]&m[876]&m[877])|(m[440]&m[873]&~m[875]&m[876]&m[877])|(~m[440]&~m[873]&m[875]&m[876]&m[877])|(m[440]&~m[873]&m[875]&m[876]&m[877])|(m[440]&m[873]&m[875]&m[876]&m[877]));
    m[879] = (((m[451]&~m[878]&~m[880]&~m[881]&~m[882])|(~m[451]&~m[878]&~m[880]&m[881]&~m[882])|(m[451]&m[878]&~m[880]&m[881]&~m[882])|(m[451]&~m[878]&m[880]&m[881]&~m[882])|(~m[451]&m[878]&~m[880]&~m[881]&m[882])|(~m[451]&~m[878]&m[880]&~m[881]&m[882])|(m[451]&m[878]&m[880]&~m[881]&m[882])|(~m[451]&m[878]&m[880]&m[881]&m[882]))&UnbiasedRNG[322])|((m[451]&~m[878]&~m[880]&m[881]&~m[882])|(~m[451]&~m[878]&~m[880]&~m[881]&m[882])|(m[451]&~m[878]&~m[880]&~m[881]&m[882])|(m[451]&m[878]&~m[880]&~m[881]&m[882])|(m[451]&~m[878]&m[880]&~m[881]&m[882])|(~m[451]&~m[878]&~m[880]&m[881]&m[882])|(m[451]&~m[878]&~m[880]&m[881]&m[882])|(~m[451]&m[878]&~m[880]&m[881]&m[882])|(m[451]&m[878]&~m[880]&m[881]&m[882])|(~m[451]&~m[878]&m[880]&m[881]&m[882])|(m[451]&~m[878]&m[880]&m[881]&m[882])|(m[451]&m[878]&m[880]&m[881]&m[882]));
    m[884] = (((m[462]&~m[883]&~m[885]&~m[886]&~m[887])|(~m[462]&~m[883]&~m[885]&m[886]&~m[887])|(m[462]&m[883]&~m[885]&m[886]&~m[887])|(m[462]&~m[883]&m[885]&m[886]&~m[887])|(~m[462]&m[883]&~m[885]&~m[886]&m[887])|(~m[462]&~m[883]&m[885]&~m[886]&m[887])|(m[462]&m[883]&m[885]&~m[886]&m[887])|(~m[462]&m[883]&m[885]&m[886]&m[887]))&UnbiasedRNG[323])|((m[462]&~m[883]&~m[885]&m[886]&~m[887])|(~m[462]&~m[883]&~m[885]&~m[886]&m[887])|(m[462]&~m[883]&~m[885]&~m[886]&m[887])|(m[462]&m[883]&~m[885]&~m[886]&m[887])|(m[462]&~m[883]&m[885]&~m[886]&m[887])|(~m[462]&~m[883]&~m[885]&m[886]&m[887])|(m[462]&~m[883]&~m[885]&m[886]&m[887])|(~m[462]&m[883]&~m[885]&m[886]&m[887])|(m[462]&m[883]&~m[885]&m[886]&m[887])|(~m[462]&~m[883]&m[885]&m[886]&m[887])|(m[462]&~m[883]&m[885]&m[886]&m[887])|(m[462]&m[883]&m[885]&m[886]&m[887]));
    m[889] = (((m[473]&~m[888]&~m[890]&~m[891]&~m[892])|(~m[473]&~m[888]&~m[890]&m[891]&~m[892])|(m[473]&m[888]&~m[890]&m[891]&~m[892])|(m[473]&~m[888]&m[890]&m[891]&~m[892])|(~m[473]&m[888]&~m[890]&~m[891]&m[892])|(~m[473]&~m[888]&m[890]&~m[891]&m[892])|(m[473]&m[888]&m[890]&~m[891]&m[892])|(~m[473]&m[888]&m[890]&m[891]&m[892]))&UnbiasedRNG[324])|((m[473]&~m[888]&~m[890]&m[891]&~m[892])|(~m[473]&~m[888]&~m[890]&~m[891]&m[892])|(m[473]&~m[888]&~m[890]&~m[891]&m[892])|(m[473]&m[888]&~m[890]&~m[891]&m[892])|(m[473]&~m[888]&m[890]&~m[891]&m[892])|(~m[473]&~m[888]&~m[890]&m[891]&m[892])|(m[473]&~m[888]&~m[890]&m[891]&m[892])|(~m[473]&m[888]&~m[890]&m[891]&m[892])|(m[473]&m[888]&~m[890]&m[891]&m[892])|(~m[473]&~m[888]&m[890]&m[891]&m[892])|(m[473]&~m[888]&m[890]&m[891]&m[892])|(m[473]&m[888]&m[890]&m[891]&m[892]));
    m[894] = (((m[484]&~m[893]&~m[895]&~m[896]&~m[897])|(~m[484]&~m[893]&~m[895]&m[896]&~m[897])|(m[484]&m[893]&~m[895]&m[896]&~m[897])|(m[484]&~m[893]&m[895]&m[896]&~m[897])|(~m[484]&m[893]&~m[895]&~m[896]&m[897])|(~m[484]&~m[893]&m[895]&~m[896]&m[897])|(m[484]&m[893]&m[895]&~m[896]&m[897])|(~m[484]&m[893]&m[895]&m[896]&m[897]))&UnbiasedRNG[325])|((m[484]&~m[893]&~m[895]&m[896]&~m[897])|(~m[484]&~m[893]&~m[895]&~m[896]&m[897])|(m[484]&~m[893]&~m[895]&~m[896]&m[897])|(m[484]&m[893]&~m[895]&~m[896]&m[897])|(m[484]&~m[893]&m[895]&~m[896]&m[897])|(~m[484]&~m[893]&~m[895]&m[896]&m[897])|(m[484]&~m[893]&~m[895]&m[896]&m[897])|(~m[484]&m[893]&~m[895]&m[896]&m[897])|(m[484]&m[893]&~m[895]&m[896]&m[897])|(~m[484]&~m[893]&m[895]&m[896]&m[897])|(m[484]&~m[893]&m[895]&m[896]&m[897])|(m[484]&m[893]&m[895]&m[896]&m[897]));
    m[899] = (((m[495]&~m[898]&~m[900]&~m[901]&~m[902])|(~m[495]&~m[898]&~m[900]&m[901]&~m[902])|(m[495]&m[898]&~m[900]&m[901]&~m[902])|(m[495]&~m[898]&m[900]&m[901]&~m[902])|(~m[495]&m[898]&~m[900]&~m[901]&m[902])|(~m[495]&~m[898]&m[900]&~m[901]&m[902])|(m[495]&m[898]&m[900]&~m[901]&m[902])|(~m[495]&m[898]&m[900]&m[901]&m[902]))&UnbiasedRNG[326])|((m[495]&~m[898]&~m[900]&m[901]&~m[902])|(~m[495]&~m[898]&~m[900]&~m[901]&m[902])|(m[495]&~m[898]&~m[900]&~m[901]&m[902])|(m[495]&m[898]&~m[900]&~m[901]&m[902])|(m[495]&~m[898]&m[900]&~m[901]&m[902])|(~m[495]&~m[898]&~m[900]&m[901]&m[902])|(m[495]&~m[898]&~m[900]&m[901]&m[902])|(~m[495]&m[898]&~m[900]&m[901]&m[902])|(m[495]&m[898]&~m[900]&m[901]&m[902])|(~m[495]&~m[898]&m[900]&m[901]&m[902])|(m[495]&~m[898]&m[900]&m[901]&m[902])|(m[495]&m[898]&m[900]&m[901]&m[902]));
    m[904] = (((m[506]&~m[903]&~m[905]&~m[906]&~m[907])|(~m[506]&~m[903]&~m[905]&m[906]&~m[907])|(m[506]&m[903]&~m[905]&m[906]&~m[907])|(m[506]&~m[903]&m[905]&m[906]&~m[907])|(~m[506]&m[903]&~m[905]&~m[906]&m[907])|(~m[506]&~m[903]&m[905]&~m[906]&m[907])|(m[506]&m[903]&m[905]&~m[906]&m[907])|(~m[506]&m[903]&m[905]&m[906]&m[907]))&UnbiasedRNG[327])|((m[506]&~m[903]&~m[905]&m[906]&~m[907])|(~m[506]&~m[903]&~m[905]&~m[906]&m[907])|(m[506]&~m[903]&~m[905]&~m[906]&m[907])|(m[506]&m[903]&~m[905]&~m[906]&m[907])|(m[506]&~m[903]&m[905]&~m[906]&m[907])|(~m[506]&~m[903]&~m[905]&m[906]&m[907])|(m[506]&~m[903]&~m[905]&m[906]&m[907])|(~m[506]&m[903]&~m[905]&m[906]&m[907])|(m[506]&m[903]&~m[905]&m[906]&m[907])|(~m[506]&~m[903]&m[905]&m[906]&m[907])|(m[506]&~m[903]&m[905]&m[906]&m[907])|(m[506]&m[903]&m[905]&m[906]&m[907]));
    m[909] = (((m[517]&~m[908]&~m[910]&~m[911]&~m[912])|(~m[517]&~m[908]&~m[910]&m[911]&~m[912])|(m[517]&m[908]&~m[910]&m[911]&~m[912])|(m[517]&~m[908]&m[910]&m[911]&~m[912])|(~m[517]&m[908]&~m[910]&~m[911]&m[912])|(~m[517]&~m[908]&m[910]&~m[911]&m[912])|(m[517]&m[908]&m[910]&~m[911]&m[912])|(~m[517]&m[908]&m[910]&m[911]&m[912]))&UnbiasedRNG[328])|((m[517]&~m[908]&~m[910]&m[911]&~m[912])|(~m[517]&~m[908]&~m[910]&~m[911]&m[912])|(m[517]&~m[908]&~m[910]&~m[911]&m[912])|(m[517]&m[908]&~m[910]&~m[911]&m[912])|(m[517]&~m[908]&m[910]&~m[911]&m[912])|(~m[517]&~m[908]&~m[910]&m[911]&m[912])|(m[517]&~m[908]&~m[910]&m[911]&m[912])|(~m[517]&m[908]&~m[910]&m[911]&m[912])|(m[517]&m[908]&~m[910]&m[911]&m[912])|(~m[517]&~m[908]&m[910]&m[911]&m[912])|(m[517]&~m[908]&m[910]&m[911]&m[912])|(m[517]&m[908]&m[910]&m[911]&m[912]));
    m[914] = (((m[419]&~m[913]&~m[915]&~m[916]&~m[917])|(~m[419]&~m[913]&~m[915]&m[916]&~m[917])|(m[419]&m[913]&~m[915]&m[916]&~m[917])|(m[419]&~m[913]&m[915]&m[916]&~m[917])|(~m[419]&m[913]&~m[915]&~m[916]&m[917])|(~m[419]&~m[913]&m[915]&~m[916]&m[917])|(m[419]&m[913]&m[915]&~m[916]&m[917])|(~m[419]&m[913]&m[915]&m[916]&m[917]))&UnbiasedRNG[329])|((m[419]&~m[913]&~m[915]&m[916]&~m[917])|(~m[419]&~m[913]&~m[915]&~m[916]&m[917])|(m[419]&~m[913]&~m[915]&~m[916]&m[917])|(m[419]&m[913]&~m[915]&~m[916]&m[917])|(m[419]&~m[913]&m[915]&~m[916]&m[917])|(~m[419]&~m[913]&~m[915]&m[916]&m[917])|(m[419]&~m[913]&~m[915]&m[916]&m[917])|(~m[419]&m[913]&~m[915]&m[916]&m[917])|(m[419]&m[913]&~m[915]&m[916]&m[917])|(~m[419]&~m[913]&m[915]&m[916]&m[917])|(m[419]&~m[913]&m[915]&m[916]&m[917])|(m[419]&m[913]&m[915]&m[916]&m[917]));
    m[919] = (((m[430]&~m[918]&~m[920]&~m[921]&~m[922])|(~m[430]&~m[918]&~m[920]&m[921]&~m[922])|(m[430]&m[918]&~m[920]&m[921]&~m[922])|(m[430]&~m[918]&m[920]&m[921]&~m[922])|(~m[430]&m[918]&~m[920]&~m[921]&m[922])|(~m[430]&~m[918]&m[920]&~m[921]&m[922])|(m[430]&m[918]&m[920]&~m[921]&m[922])|(~m[430]&m[918]&m[920]&m[921]&m[922]))&UnbiasedRNG[330])|((m[430]&~m[918]&~m[920]&m[921]&~m[922])|(~m[430]&~m[918]&~m[920]&~m[921]&m[922])|(m[430]&~m[918]&~m[920]&~m[921]&m[922])|(m[430]&m[918]&~m[920]&~m[921]&m[922])|(m[430]&~m[918]&m[920]&~m[921]&m[922])|(~m[430]&~m[918]&~m[920]&m[921]&m[922])|(m[430]&~m[918]&~m[920]&m[921]&m[922])|(~m[430]&m[918]&~m[920]&m[921]&m[922])|(m[430]&m[918]&~m[920]&m[921]&m[922])|(~m[430]&~m[918]&m[920]&m[921]&m[922])|(m[430]&~m[918]&m[920]&m[921]&m[922])|(m[430]&m[918]&m[920]&m[921]&m[922]));
    m[924] = (((m[441]&~m[923]&~m[925]&~m[926]&~m[927])|(~m[441]&~m[923]&~m[925]&m[926]&~m[927])|(m[441]&m[923]&~m[925]&m[926]&~m[927])|(m[441]&~m[923]&m[925]&m[926]&~m[927])|(~m[441]&m[923]&~m[925]&~m[926]&m[927])|(~m[441]&~m[923]&m[925]&~m[926]&m[927])|(m[441]&m[923]&m[925]&~m[926]&m[927])|(~m[441]&m[923]&m[925]&m[926]&m[927]))&UnbiasedRNG[331])|((m[441]&~m[923]&~m[925]&m[926]&~m[927])|(~m[441]&~m[923]&~m[925]&~m[926]&m[927])|(m[441]&~m[923]&~m[925]&~m[926]&m[927])|(m[441]&m[923]&~m[925]&~m[926]&m[927])|(m[441]&~m[923]&m[925]&~m[926]&m[927])|(~m[441]&~m[923]&~m[925]&m[926]&m[927])|(m[441]&~m[923]&~m[925]&m[926]&m[927])|(~m[441]&m[923]&~m[925]&m[926]&m[927])|(m[441]&m[923]&~m[925]&m[926]&m[927])|(~m[441]&~m[923]&m[925]&m[926]&m[927])|(m[441]&~m[923]&m[925]&m[926]&m[927])|(m[441]&m[923]&m[925]&m[926]&m[927]));
    m[929] = (((m[452]&~m[928]&~m[930]&~m[931]&~m[932])|(~m[452]&~m[928]&~m[930]&m[931]&~m[932])|(m[452]&m[928]&~m[930]&m[931]&~m[932])|(m[452]&~m[928]&m[930]&m[931]&~m[932])|(~m[452]&m[928]&~m[930]&~m[931]&m[932])|(~m[452]&~m[928]&m[930]&~m[931]&m[932])|(m[452]&m[928]&m[930]&~m[931]&m[932])|(~m[452]&m[928]&m[930]&m[931]&m[932]))&UnbiasedRNG[332])|((m[452]&~m[928]&~m[930]&m[931]&~m[932])|(~m[452]&~m[928]&~m[930]&~m[931]&m[932])|(m[452]&~m[928]&~m[930]&~m[931]&m[932])|(m[452]&m[928]&~m[930]&~m[931]&m[932])|(m[452]&~m[928]&m[930]&~m[931]&m[932])|(~m[452]&~m[928]&~m[930]&m[931]&m[932])|(m[452]&~m[928]&~m[930]&m[931]&m[932])|(~m[452]&m[928]&~m[930]&m[931]&m[932])|(m[452]&m[928]&~m[930]&m[931]&m[932])|(~m[452]&~m[928]&m[930]&m[931]&m[932])|(m[452]&~m[928]&m[930]&m[931]&m[932])|(m[452]&m[928]&m[930]&m[931]&m[932]));
    m[934] = (((m[463]&~m[933]&~m[935]&~m[936]&~m[937])|(~m[463]&~m[933]&~m[935]&m[936]&~m[937])|(m[463]&m[933]&~m[935]&m[936]&~m[937])|(m[463]&~m[933]&m[935]&m[936]&~m[937])|(~m[463]&m[933]&~m[935]&~m[936]&m[937])|(~m[463]&~m[933]&m[935]&~m[936]&m[937])|(m[463]&m[933]&m[935]&~m[936]&m[937])|(~m[463]&m[933]&m[935]&m[936]&m[937]))&UnbiasedRNG[333])|((m[463]&~m[933]&~m[935]&m[936]&~m[937])|(~m[463]&~m[933]&~m[935]&~m[936]&m[937])|(m[463]&~m[933]&~m[935]&~m[936]&m[937])|(m[463]&m[933]&~m[935]&~m[936]&m[937])|(m[463]&~m[933]&m[935]&~m[936]&m[937])|(~m[463]&~m[933]&~m[935]&m[936]&m[937])|(m[463]&~m[933]&~m[935]&m[936]&m[937])|(~m[463]&m[933]&~m[935]&m[936]&m[937])|(m[463]&m[933]&~m[935]&m[936]&m[937])|(~m[463]&~m[933]&m[935]&m[936]&m[937])|(m[463]&~m[933]&m[935]&m[936]&m[937])|(m[463]&m[933]&m[935]&m[936]&m[937]));
    m[939] = (((m[474]&~m[938]&~m[940]&~m[941]&~m[942])|(~m[474]&~m[938]&~m[940]&m[941]&~m[942])|(m[474]&m[938]&~m[940]&m[941]&~m[942])|(m[474]&~m[938]&m[940]&m[941]&~m[942])|(~m[474]&m[938]&~m[940]&~m[941]&m[942])|(~m[474]&~m[938]&m[940]&~m[941]&m[942])|(m[474]&m[938]&m[940]&~m[941]&m[942])|(~m[474]&m[938]&m[940]&m[941]&m[942]))&UnbiasedRNG[334])|((m[474]&~m[938]&~m[940]&m[941]&~m[942])|(~m[474]&~m[938]&~m[940]&~m[941]&m[942])|(m[474]&~m[938]&~m[940]&~m[941]&m[942])|(m[474]&m[938]&~m[940]&~m[941]&m[942])|(m[474]&~m[938]&m[940]&~m[941]&m[942])|(~m[474]&~m[938]&~m[940]&m[941]&m[942])|(m[474]&~m[938]&~m[940]&m[941]&m[942])|(~m[474]&m[938]&~m[940]&m[941]&m[942])|(m[474]&m[938]&~m[940]&m[941]&m[942])|(~m[474]&~m[938]&m[940]&m[941]&m[942])|(m[474]&~m[938]&m[940]&m[941]&m[942])|(m[474]&m[938]&m[940]&m[941]&m[942]));
    m[944] = (((m[485]&~m[943]&~m[945]&~m[946]&~m[947])|(~m[485]&~m[943]&~m[945]&m[946]&~m[947])|(m[485]&m[943]&~m[945]&m[946]&~m[947])|(m[485]&~m[943]&m[945]&m[946]&~m[947])|(~m[485]&m[943]&~m[945]&~m[946]&m[947])|(~m[485]&~m[943]&m[945]&~m[946]&m[947])|(m[485]&m[943]&m[945]&~m[946]&m[947])|(~m[485]&m[943]&m[945]&m[946]&m[947]))&UnbiasedRNG[335])|((m[485]&~m[943]&~m[945]&m[946]&~m[947])|(~m[485]&~m[943]&~m[945]&~m[946]&m[947])|(m[485]&~m[943]&~m[945]&~m[946]&m[947])|(m[485]&m[943]&~m[945]&~m[946]&m[947])|(m[485]&~m[943]&m[945]&~m[946]&m[947])|(~m[485]&~m[943]&~m[945]&m[946]&m[947])|(m[485]&~m[943]&~m[945]&m[946]&m[947])|(~m[485]&m[943]&~m[945]&m[946]&m[947])|(m[485]&m[943]&~m[945]&m[946]&m[947])|(~m[485]&~m[943]&m[945]&m[946]&m[947])|(m[485]&~m[943]&m[945]&m[946]&m[947])|(m[485]&m[943]&m[945]&m[946]&m[947]));
    m[949] = (((m[496]&~m[948]&~m[950]&~m[951]&~m[952])|(~m[496]&~m[948]&~m[950]&m[951]&~m[952])|(m[496]&m[948]&~m[950]&m[951]&~m[952])|(m[496]&~m[948]&m[950]&m[951]&~m[952])|(~m[496]&m[948]&~m[950]&~m[951]&m[952])|(~m[496]&~m[948]&m[950]&~m[951]&m[952])|(m[496]&m[948]&m[950]&~m[951]&m[952])|(~m[496]&m[948]&m[950]&m[951]&m[952]))&UnbiasedRNG[336])|((m[496]&~m[948]&~m[950]&m[951]&~m[952])|(~m[496]&~m[948]&~m[950]&~m[951]&m[952])|(m[496]&~m[948]&~m[950]&~m[951]&m[952])|(m[496]&m[948]&~m[950]&~m[951]&m[952])|(m[496]&~m[948]&m[950]&~m[951]&m[952])|(~m[496]&~m[948]&~m[950]&m[951]&m[952])|(m[496]&~m[948]&~m[950]&m[951]&m[952])|(~m[496]&m[948]&~m[950]&m[951]&m[952])|(m[496]&m[948]&~m[950]&m[951]&m[952])|(~m[496]&~m[948]&m[950]&m[951]&m[952])|(m[496]&~m[948]&m[950]&m[951]&m[952])|(m[496]&m[948]&m[950]&m[951]&m[952]));
    m[954] = (((m[507]&~m[953]&~m[955]&~m[956]&~m[957])|(~m[507]&~m[953]&~m[955]&m[956]&~m[957])|(m[507]&m[953]&~m[955]&m[956]&~m[957])|(m[507]&~m[953]&m[955]&m[956]&~m[957])|(~m[507]&m[953]&~m[955]&~m[956]&m[957])|(~m[507]&~m[953]&m[955]&~m[956]&m[957])|(m[507]&m[953]&m[955]&~m[956]&m[957])|(~m[507]&m[953]&m[955]&m[956]&m[957]))&UnbiasedRNG[337])|((m[507]&~m[953]&~m[955]&m[956]&~m[957])|(~m[507]&~m[953]&~m[955]&~m[956]&m[957])|(m[507]&~m[953]&~m[955]&~m[956]&m[957])|(m[507]&m[953]&~m[955]&~m[956]&m[957])|(m[507]&~m[953]&m[955]&~m[956]&m[957])|(~m[507]&~m[953]&~m[955]&m[956]&m[957])|(m[507]&~m[953]&~m[955]&m[956]&m[957])|(~m[507]&m[953]&~m[955]&m[956]&m[957])|(m[507]&m[953]&~m[955]&m[956]&m[957])|(~m[507]&~m[953]&m[955]&m[956]&m[957])|(m[507]&~m[953]&m[955]&m[956]&m[957])|(m[507]&m[953]&m[955]&m[956]&m[957]));
    m[959] = (((m[518]&~m[958]&~m[960]&~m[961]&~m[962])|(~m[518]&~m[958]&~m[960]&m[961]&~m[962])|(m[518]&m[958]&~m[960]&m[961]&~m[962])|(m[518]&~m[958]&m[960]&m[961]&~m[962])|(~m[518]&m[958]&~m[960]&~m[961]&m[962])|(~m[518]&~m[958]&m[960]&~m[961]&m[962])|(m[518]&m[958]&m[960]&~m[961]&m[962])|(~m[518]&m[958]&m[960]&m[961]&m[962]))&UnbiasedRNG[338])|((m[518]&~m[958]&~m[960]&m[961]&~m[962])|(~m[518]&~m[958]&~m[960]&~m[961]&m[962])|(m[518]&~m[958]&~m[960]&~m[961]&m[962])|(m[518]&m[958]&~m[960]&~m[961]&m[962])|(m[518]&~m[958]&m[960]&~m[961]&m[962])|(~m[518]&~m[958]&~m[960]&m[961]&m[962])|(m[518]&~m[958]&~m[960]&m[961]&m[962])|(~m[518]&m[958]&~m[960]&m[961]&m[962])|(m[518]&m[958]&~m[960]&m[961]&m[962])|(~m[518]&~m[958]&m[960]&m[961]&m[962])|(m[518]&~m[958]&m[960]&m[961]&m[962])|(m[518]&m[958]&m[960]&m[961]&m[962]));
    m[964] = (((m[431]&~m[963]&~m[965]&~m[966]&~m[967])|(~m[431]&~m[963]&~m[965]&m[966]&~m[967])|(m[431]&m[963]&~m[965]&m[966]&~m[967])|(m[431]&~m[963]&m[965]&m[966]&~m[967])|(~m[431]&m[963]&~m[965]&~m[966]&m[967])|(~m[431]&~m[963]&m[965]&~m[966]&m[967])|(m[431]&m[963]&m[965]&~m[966]&m[967])|(~m[431]&m[963]&m[965]&m[966]&m[967]))&UnbiasedRNG[339])|((m[431]&~m[963]&~m[965]&m[966]&~m[967])|(~m[431]&~m[963]&~m[965]&~m[966]&m[967])|(m[431]&~m[963]&~m[965]&~m[966]&m[967])|(m[431]&m[963]&~m[965]&~m[966]&m[967])|(m[431]&~m[963]&m[965]&~m[966]&m[967])|(~m[431]&~m[963]&~m[965]&m[966]&m[967])|(m[431]&~m[963]&~m[965]&m[966]&m[967])|(~m[431]&m[963]&~m[965]&m[966]&m[967])|(m[431]&m[963]&~m[965]&m[966]&m[967])|(~m[431]&~m[963]&m[965]&m[966]&m[967])|(m[431]&~m[963]&m[965]&m[966]&m[967])|(m[431]&m[963]&m[965]&m[966]&m[967]));
    m[969] = (((m[442]&~m[968]&~m[970]&~m[971]&~m[972])|(~m[442]&~m[968]&~m[970]&m[971]&~m[972])|(m[442]&m[968]&~m[970]&m[971]&~m[972])|(m[442]&~m[968]&m[970]&m[971]&~m[972])|(~m[442]&m[968]&~m[970]&~m[971]&m[972])|(~m[442]&~m[968]&m[970]&~m[971]&m[972])|(m[442]&m[968]&m[970]&~m[971]&m[972])|(~m[442]&m[968]&m[970]&m[971]&m[972]))&UnbiasedRNG[340])|((m[442]&~m[968]&~m[970]&m[971]&~m[972])|(~m[442]&~m[968]&~m[970]&~m[971]&m[972])|(m[442]&~m[968]&~m[970]&~m[971]&m[972])|(m[442]&m[968]&~m[970]&~m[971]&m[972])|(m[442]&~m[968]&m[970]&~m[971]&m[972])|(~m[442]&~m[968]&~m[970]&m[971]&m[972])|(m[442]&~m[968]&~m[970]&m[971]&m[972])|(~m[442]&m[968]&~m[970]&m[971]&m[972])|(m[442]&m[968]&~m[970]&m[971]&m[972])|(~m[442]&~m[968]&m[970]&m[971]&m[972])|(m[442]&~m[968]&m[970]&m[971]&m[972])|(m[442]&m[968]&m[970]&m[971]&m[972]));
    m[974] = (((m[453]&~m[973]&~m[975]&~m[976]&~m[977])|(~m[453]&~m[973]&~m[975]&m[976]&~m[977])|(m[453]&m[973]&~m[975]&m[976]&~m[977])|(m[453]&~m[973]&m[975]&m[976]&~m[977])|(~m[453]&m[973]&~m[975]&~m[976]&m[977])|(~m[453]&~m[973]&m[975]&~m[976]&m[977])|(m[453]&m[973]&m[975]&~m[976]&m[977])|(~m[453]&m[973]&m[975]&m[976]&m[977]))&UnbiasedRNG[341])|((m[453]&~m[973]&~m[975]&m[976]&~m[977])|(~m[453]&~m[973]&~m[975]&~m[976]&m[977])|(m[453]&~m[973]&~m[975]&~m[976]&m[977])|(m[453]&m[973]&~m[975]&~m[976]&m[977])|(m[453]&~m[973]&m[975]&~m[976]&m[977])|(~m[453]&~m[973]&~m[975]&m[976]&m[977])|(m[453]&~m[973]&~m[975]&m[976]&m[977])|(~m[453]&m[973]&~m[975]&m[976]&m[977])|(m[453]&m[973]&~m[975]&m[976]&m[977])|(~m[453]&~m[973]&m[975]&m[976]&m[977])|(m[453]&~m[973]&m[975]&m[976]&m[977])|(m[453]&m[973]&m[975]&m[976]&m[977]));
    m[979] = (((m[464]&~m[978]&~m[980]&~m[981]&~m[982])|(~m[464]&~m[978]&~m[980]&m[981]&~m[982])|(m[464]&m[978]&~m[980]&m[981]&~m[982])|(m[464]&~m[978]&m[980]&m[981]&~m[982])|(~m[464]&m[978]&~m[980]&~m[981]&m[982])|(~m[464]&~m[978]&m[980]&~m[981]&m[982])|(m[464]&m[978]&m[980]&~m[981]&m[982])|(~m[464]&m[978]&m[980]&m[981]&m[982]))&UnbiasedRNG[342])|((m[464]&~m[978]&~m[980]&m[981]&~m[982])|(~m[464]&~m[978]&~m[980]&~m[981]&m[982])|(m[464]&~m[978]&~m[980]&~m[981]&m[982])|(m[464]&m[978]&~m[980]&~m[981]&m[982])|(m[464]&~m[978]&m[980]&~m[981]&m[982])|(~m[464]&~m[978]&~m[980]&m[981]&m[982])|(m[464]&~m[978]&~m[980]&m[981]&m[982])|(~m[464]&m[978]&~m[980]&m[981]&m[982])|(m[464]&m[978]&~m[980]&m[981]&m[982])|(~m[464]&~m[978]&m[980]&m[981]&m[982])|(m[464]&~m[978]&m[980]&m[981]&m[982])|(m[464]&m[978]&m[980]&m[981]&m[982]));
    m[984] = (((m[475]&~m[983]&~m[985]&~m[986]&~m[987])|(~m[475]&~m[983]&~m[985]&m[986]&~m[987])|(m[475]&m[983]&~m[985]&m[986]&~m[987])|(m[475]&~m[983]&m[985]&m[986]&~m[987])|(~m[475]&m[983]&~m[985]&~m[986]&m[987])|(~m[475]&~m[983]&m[985]&~m[986]&m[987])|(m[475]&m[983]&m[985]&~m[986]&m[987])|(~m[475]&m[983]&m[985]&m[986]&m[987]))&UnbiasedRNG[343])|((m[475]&~m[983]&~m[985]&m[986]&~m[987])|(~m[475]&~m[983]&~m[985]&~m[986]&m[987])|(m[475]&~m[983]&~m[985]&~m[986]&m[987])|(m[475]&m[983]&~m[985]&~m[986]&m[987])|(m[475]&~m[983]&m[985]&~m[986]&m[987])|(~m[475]&~m[983]&~m[985]&m[986]&m[987])|(m[475]&~m[983]&~m[985]&m[986]&m[987])|(~m[475]&m[983]&~m[985]&m[986]&m[987])|(m[475]&m[983]&~m[985]&m[986]&m[987])|(~m[475]&~m[983]&m[985]&m[986]&m[987])|(m[475]&~m[983]&m[985]&m[986]&m[987])|(m[475]&m[983]&m[985]&m[986]&m[987]));
    m[989] = (((m[486]&~m[988]&~m[990]&~m[991]&~m[992])|(~m[486]&~m[988]&~m[990]&m[991]&~m[992])|(m[486]&m[988]&~m[990]&m[991]&~m[992])|(m[486]&~m[988]&m[990]&m[991]&~m[992])|(~m[486]&m[988]&~m[990]&~m[991]&m[992])|(~m[486]&~m[988]&m[990]&~m[991]&m[992])|(m[486]&m[988]&m[990]&~m[991]&m[992])|(~m[486]&m[988]&m[990]&m[991]&m[992]))&UnbiasedRNG[344])|((m[486]&~m[988]&~m[990]&m[991]&~m[992])|(~m[486]&~m[988]&~m[990]&~m[991]&m[992])|(m[486]&~m[988]&~m[990]&~m[991]&m[992])|(m[486]&m[988]&~m[990]&~m[991]&m[992])|(m[486]&~m[988]&m[990]&~m[991]&m[992])|(~m[486]&~m[988]&~m[990]&m[991]&m[992])|(m[486]&~m[988]&~m[990]&m[991]&m[992])|(~m[486]&m[988]&~m[990]&m[991]&m[992])|(m[486]&m[988]&~m[990]&m[991]&m[992])|(~m[486]&~m[988]&m[990]&m[991]&m[992])|(m[486]&~m[988]&m[990]&m[991]&m[992])|(m[486]&m[988]&m[990]&m[991]&m[992]));
    m[994] = (((m[497]&~m[993]&~m[995]&~m[996]&~m[997])|(~m[497]&~m[993]&~m[995]&m[996]&~m[997])|(m[497]&m[993]&~m[995]&m[996]&~m[997])|(m[497]&~m[993]&m[995]&m[996]&~m[997])|(~m[497]&m[993]&~m[995]&~m[996]&m[997])|(~m[497]&~m[993]&m[995]&~m[996]&m[997])|(m[497]&m[993]&m[995]&~m[996]&m[997])|(~m[497]&m[993]&m[995]&m[996]&m[997]))&UnbiasedRNG[345])|((m[497]&~m[993]&~m[995]&m[996]&~m[997])|(~m[497]&~m[993]&~m[995]&~m[996]&m[997])|(m[497]&~m[993]&~m[995]&~m[996]&m[997])|(m[497]&m[993]&~m[995]&~m[996]&m[997])|(m[497]&~m[993]&m[995]&~m[996]&m[997])|(~m[497]&~m[993]&~m[995]&m[996]&m[997])|(m[497]&~m[993]&~m[995]&m[996]&m[997])|(~m[497]&m[993]&~m[995]&m[996]&m[997])|(m[497]&m[993]&~m[995]&m[996]&m[997])|(~m[497]&~m[993]&m[995]&m[996]&m[997])|(m[497]&~m[993]&m[995]&m[996]&m[997])|(m[497]&m[993]&m[995]&m[996]&m[997]));
    m[999] = (((m[508]&~m[998]&~m[1000]&~m[1001]&~m[1002])|(~m[508]&~m[998]&~m[1000]&m[1001]&~m[1002])|(m[508]&m[998]&~m[1000]&m[1001]&~m[1002])|(m[508]&~m[998]&m[1000]&m[1001]&~m[1002])|(~m[508]&m[998]&~m[1000]&~m[1001]&m[1002])|(~m[508]&~m[998]&m[1000]&~m[1001]&m[1002])|(m[508]&m[998]&m[1000]&~m[1001]&m[1002])|(~m[508]&m[998]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[346])|((m[508]&~m[998]&~m[1000]&m[1001]&~m[1002])|(~m[508]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[508]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[508]&m[998]&~m[1000]&~m[1001]&m[1002])|(m[508]&~m[998]&m[1000]&~m[1001]&m[1002])|(~m[508]&~m[998]&~m[1000]&m[1001]&m[1002])|(m[508]&~m[998]&~m[1000]&m[1001]&m[1002])|(~m[508]&m[998]&~m[1000]&m[1001]&m[1002])|(m[508]&m[998]&~m[1000]&m[1001]&m[1002])|(~m[508]&~m[998]&m[1000]&m[1001]&m[1002])|(m[508]&~m[998]&m[1000]&m[1001]&m[1002])|(m[508]&m[998]&m[1000]&m[1001]&m[1002]));
    m[1004] = (((m[519]&~m[1003]&~m[1005]&~m[1006]&~m[1007])|(~m[519]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(m[519]&m[1003]&~m[1005]&m[1006]&~m[1007])|(m[519]&~m[1003]&m[1005]&m[1006]&~m[1007])|(~m[519]&m[1003]&~m[1005]&~m[1006]&m[1007])|(~m[519]&~m[1003]&m[1005]&~m[1006]&m[1007])|(m[519]&m[1003]&m[1005]&~m[1006]&m[1007])|(~m[519]&m[1003]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[347])|((m[519]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(~m[519]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[519]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[519]&m[1003]&~m[1005]&~m[1006]&m[1007])|(m[519]&~m[1003]&m[1005]&~m[1006]&m[1007])|(~m[519]&~m[1003]&~m[1005]&m[1006]&m[1007])|(m[519]&~m[1003]&~m[1005]&m[1006]&m[1007])|(~m[519]&m[1003]&~m[1005]&m[1006]&m[1007])|(m[519]&m[1003]&~m[1005]&m[1006]&m[1007])|(~m[519]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[519]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[519]&m[1003]&m[1005]&m[1006]&m[1007]));
    m[1009] = (((m[443]&~m[1008]&~m[1010]&~m[1011]&~m[1012])|(~m[443]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(m[443]&m[1008]&~m[1010]&m[1011]&~m[1012])|(m[443]&~m[1008]&m[1010]&m[1011]&~m[1012])|(~m[443]&m[1008]&~m[1010]&~m[1011]&m[1012])|(~m[443]&~m[1008]&m[1010]&~m[1011]&m[1012])|(m[443]&m[1008]&m[1010]&~m[1011]&m[1012])|(~m[443]&m[1008]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[348])|((m[443]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(~m[443]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[443]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[443]&m[1008]&~m[1010]&~m[1011]&m[1012])|(m[443]&~m[1008]&m[1010]&~m[1011]&m[1012])|(~m[443]&~m[1008]&~m[1010]&m[1011]&m[1012])|(m[443]&~m[1008]&~m[1010]&m[1011]&m[1012])|(~m[443]&m[1008]&~m[1010]&m[1011]&m[1012])|(m[443]&m[1008]&~m[1010]&m[1011]&m[1012])|(~m[443]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[443]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[443]&m[1008]&m[1010]&m[1011]&m[1012]));
    m[1014] = (((m[454]&~m[1013]&~m[1015]&~m[1016]&~m[1017])|(~m[454]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(m[454]&m[1013]&~m[1015]&m[1016]&~m[1017])|(m[454]&~m[1013]&m[1015]&m[1016]&~m[1017])|(~m[454]&m[1013]&~m[1015]&~m[1016]&m[1017])|(~m[454]&~m[1013]&m[1015]&~m[1016]&m[1017])|(m[454]&m[1013]&m[1015]&~m[1016]&m[1017])|(~m[454]&m[1013]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[349])|((m[454]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(~m[454]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[454]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[454]&m[1013]&~m[1015]&~m[1016]&m[1017])|(m[454]&~m[1013]&m[1015]&~m[1016]&m[1017])|(~m[454]&~m[1013]&~m[1015]&m[1016]&m[1017])|(m[454]&~m[1013]&~m[1015]&m[1016]&m[1017])|(~m[454]&m[1013]&~m[1015]&m[1016]&m[1017])|(m[454]&m[1013]&~m[1015]&m[1016]&m[1017])|(~m[454]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[454]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[454]&m[1013]&m[1015]&m[1016]&m[1017]));
    m[1019] = (((m[465]&~m[1018]&~m[1020]&~m[1021]&~m[1022])|(~m[465]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(m[465]&m[1018]&~m[1020]&m[1021]&~m[1022])|(m[465]&~m[1018]&m[1020]&m[1021]&~m[1022])|(~m[465]&m[1018]&~m[1020]&~m[1021]&m[1022])|(~m[465]&~m[1018]&m[1020]&~m[1021]&m[1022])|(m[465]&m[1018]&m[1020]&~m[1021]&m[1022])|(~m[465]&m[1018]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[350])|((m[465]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(~m[465]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[465]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[465]&m[1018]&~m[1020]&~m[1021]&m[1022])|(m[465]&~m[1018]&m[1020]&~m[1021]&m[1022])|(~m[465]&~m[1018]&~m[1020]&m[1021]&m[1022])|(m[465]&~m[1018]&~m[1020]&m[1021]&m[1022])|(~m[465]&m[1018]&~m[1020]&m[1021]&m[1022])|(m[465]&m[1018]&~m[1020]&m[1021]&m[1022])|(~m[465]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[465]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[465]&m[1018]&m[1020]&m[1021]&m[1022]));
    m[1024] = (((m[476]&~m[1023]&~m[1025]&~m[1026]&~m[1027])|(~m[476]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(m[476]&m[1023]&~m[1025]&m[1026]&~m[1027])|(m[476]&~m[1023]&m[1025]&m[1026]&~m[1027])|(~m[476]&m[1023]&~m[1025]&~m[1026]&m[1027])|(~m[476]&~m[1023]&m[1025]&~m[1026]&m[1027])|(m[476]&m[1023]&m[1025]&~m[1026]&m[1027])|(~m[476]&m[1023]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[351])|((m[476]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(~m[476]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[476]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[476]&m[1023]&~m[1025]&~m[1026]&m[1027])|(m[476]&~m[1023]&m[1025]&~m[1026]&m[1027])|(~m[476]&~m[1023]&~m[1025]&m[1026]&m[1027])|(m[476]&~m[1023]&~m[1025]&m[1026]&m[1027])|(~m[476]&m[1023]&~m[1025]&m[1026]&m[1027])|(m[476]&m[1023]&~m[1025]&m[1026]&m[1027])|(~m[476]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[476]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[476]&m[1023]&m[1025]&m[1026]&m[1027]));
    m[1029] = (((m[487]&~m[1028]&~m[1030]&~m[1031]&~m[1032])|(~m[487]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(m[487]&m[1028]&~m[1030]&m[1031]&~m[1032])|(m[487]&~m[1028]&m[1030]&m[1031]&~m[1032])|(~m[487]&m[1028]&~m[1030]&~m[1031]&m[1032])|(~m[487]&~m[1028]&m[1030]&~m[1031]&m[1032])|(m[487]&m[1028]&m[1030]&~m[1031]&m[1032])|(~m[487]&m[1028]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[352])|((m[487]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(~m[487]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[487]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[487]&m[1028]&~m[1030]&~m[1031]&m[1032])|(m[487]&~m[1028]&m[1030]&~m[1031]&m[1032])|(~m[487]&~m[1028]&~m[1030]&m[1031]&m[1032])|(m[487]&~m[1028]&~m[1030]&m[1031]&m[1032])|(~m[487]&m[1028]&~m[1030]&m[1031]&m[1032])|(m[487]&m[1028]&~m[1030]&m[1031]&m[1032])|(~m[487]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[487]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[487]&m[1028]&m[1030]&m[1031]&m[1032]));
    m[1034] = (((m[498]&~m[1033]&~m[1035]&~m[1036]&~m[1037])|(~m[498]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(m[498]&m[1033]&~m[1035]&m[1036]&~m[1037])|(m[498]&~m[1033]&m[1035]&m[1036]&~m[1037])|(~m[498]&m[1033]&~m[1035]&~m[1036]&m[1037])|(~m[498]&~m[1033]&m[1035]&~m[1036]&m[1037])|(m[498]&m[1033]&m[1035]&~m[1036]&m[1037])|(~m[498]&m[1033]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[353])|((m[498]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(~m[498]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[498]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[498]&m[1033]&~m[1035]&~m[1036]&m[1037])|(m[498]&~m[1033]&m[1035]&~m[1036]&m[1037])|(~m[498]&~m[1033]&~m[1035]&m[1036]&m[1037])|(m[498]&~m[1033]&~m[1035]&m[1036]&m[1037])|(~m[498]&m[1033]&~m[1035]&m[1036]&m[1037])|(m[498]&m[1033]&~m[1035]&m[1036]&m[1037])|(~m[498]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[498]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[498]&m[1033]&m[1035]&m[1036]&m[1037]));
    m[1039] = (((m[509]&~m[1038]&~m[1040]&~m[1041]&~m[1042])|(~m[509]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(m[509]&m[1038]&~m[1040]&m[1041]&~m[1042])|(m[509]&~m[1038]&m[1040]&m[1041]&~m[1042])|(~m[509]&m[1038]&~m[1040]&~m[1041]&m[1042])|(~m[509]&~m[1038]&m[1040]&~m[1041]&m[1042])|(m[509]&m[1038]&m[1040]&~m[1041]&m[1042])|(~m[509]&m[1038]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[354])|((m[509]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(~m[509]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[509]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[509]&m[1038]&~m[1040]&~m[1041]&m[1042])|(m[509]&~m[1038]&m[1040]&~m[1041]&m[1042])|(~m[509]&~m[1038]&~m[1040]&m[1041]&m[1042])|(m[509]&~m[1038]&~m[1040]&m[1041]&m[1042])|(~m[509]&m[1038]&~m[1040]&m[1041]&m[1042])|(m[509]&m[1038]&~m[1040]&m[1041]&m[1042])|(~m[509]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[509]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[509]&m[1038]&m[1040]&m[1041]&m[1042]));
    m[1044] = (((m[520]&~m[1043]&~m[1045]&~m[1046]&~m[1047])|(~m[520]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(m[520]&m[1043]&~m[1045]&m[1046]&~m[1047])|(m[520]&~m[1043]&m[1045]&m[1046]&~m[1047])|(~m[520]&m[1043]&~m[1045]&~m[1046]&m[1047])|(~m[520]&~m[1043]&m[1045]&~m[1046]&m[1047])|(m[520]&m[1043]&m[1045]&~m[1046]&m[1047])|(~m[520]&m[1043]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[355])|((m[520]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(~m[520]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[520]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[520]&m[1043]&~m[1045]&~m[1046]&m[1047])|(m[520]&~m[1043]&m[1045]&~m[1046]&m[1047])|(~m[520]&~m[1043]&~m[1045]&m[1046]&m[1047])|(m[520]&~m[1043]&~m[1045]&m[1046]&m[1047])|(~m[520]&m[1043]&~m[1045]&m[1046]&m[1047])|(m[520]&m[1043]&~m[1045]&m[1046]&m[1047])|(~m[520]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[520]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[520]&m[1043]&m[1045]&m[1046]&m[1047]));
    m[1049] = (((m[455]&~m[1048]&~m[1050]&~m[1051]&~m[1052])|(~m[455]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(m[455]&m[1048]&~m[1050]&m[1051]&~m[1052])|(m[455]&~m[1048]&m[1050]&m[1051]&~m[1052])|(~m[455]&m[1048]&~m[1050]&~m[1051]&m[1052])|(~m[455]&~m[1048]&m[1050]&~m[1051]&m[1052])|(m[455]&m[1048]&m[1050]&~m[1051]&m[1052])|(~m[455]&m[1048]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[356])|((m[455]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(~m[455]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[455]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[455]&m[1048]&~m[1050]&~m[1051]&m[1052])|(m[455]&~m[1048]&m[1050]&~m[1051]&m[1052])|(~m[455]&~m[1048]&~m[1050]&m[1051]&m[1052])|(m[455]&~m[1048]&~m[1050]&m[1051]&m[1052])|(~m[455]&m[1048]&~m[1050]&m[1051]&m[1052])|(m[455]&m[1048]&~m[1050]&m[1051]&m[1052])|(~m[455]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[455]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[455]&m[1048]&m[1050]&m[1051]&m[1052]));
    m[1054] = (((m[466]&~m[1053]&~m[1055]&~m[1056]&~m[1057])|(~m[466]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(m[466]&m[1053]&~m[1055]&m[1056]&~m[1057])|(m[466]&~m[1053]&m[1055]&m[1056]&~m[1057])|(~m[466]&m[1053]&~m[1055]&~m[1056]&m[1057])|(~m[466]&~m[1053]&m[1055]&~m[1056]&m[1057])|(m[466]&m[1053]&m[1055]&~m[1056]&m[1057])|(~m[466]&m[1053]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[357])|((m[466]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(~m[466]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[466]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[466]&m[1053]&~m[1055]&~m[1056]&m[1057])|(m[466]&~m[1053]&m[1055]&~m[1056]&m[1057])|(~m[466]&~m[1053]&~m[1055]&m[1056]&m[1057])|(m[466]&~m[1053]&~m[1055]&m[1056]&m[1057])|(~m[466]&m[1053]&~m[1055]&m[1056]&m[1057])|(m[466]&m[1053]&~m[1055]&m[1056]&m[1057])|(~m[466]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[466]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[466]&m[1053]&m[1055]&m[1056]&m[1057]));
    m[1059] = (((m[477]&~m[1058]&~m[1060]&~m[1061]&~m[1062])|(~m[477]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(m[477]&m[1058]&~m[1060]&m[1061]&~m[1062])|(m[477]&~m[1058]&m[1060]&m[1061]&~m[1062])|(~m[477]&m[1058]&~m[1060]&~m[1061]&m[1062])|(~m[477]&~m[1058]&m[1060]&~m[1061]&m[1062])|(m[477]&m[1058]&m[1060]&~m[1061]&m[1062])|(~m[477]&m[1058]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[358])|((m[477]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(~m[477]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[477]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[477]&m[1058]&~m[1060]&~m[1061]&m[1062])|(m[477]&~m[1058]&m[1060]&~m[1061]&m[1062])|(~m[477]&~m[1058]&~m[1060]&m[1061]&m[1062])|(m[477]&~m[1058]&~m[1060]&m[1061]&m[1062])|(~m[477]&m[1058]&~m[1060]&m[1061]&m[1062])|(m[477]&m[1058]&~m[1060]&m[1061]&m[1062])|(~m[477]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[477]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[477]&m[1058]&m[1060]&m[1061]&m[1062]));
    m[1064] = (((m[488]&~m[1063]&~m[1065]&~m[1066]&~m[1067])|(~m[488]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(m[488]&m[1063]&~m[1065]&m[1066]&~m[1067])|(m[488]&~m[1063]&m[1065]&m[1066]&~m[1067])|(~m[488]&m[1063]&~m[1065]&~m[1066]&m[1067])|(~m[488]&~m[1063]&m[1065]&~m[1066]&m[1067])|(m[488]&m[1063]&m[1065]&~m[1066]&m[1067])|(~m[488]&m[1063]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[359])|((m[488]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(~m[488]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[488]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[488]&m[1063]&~m[1065]&~m[1066]&m[1067])|(m[488]&~m[1063]&m[1065]&~m[1066]&m[1067])|(~m[488]&~m[1063]&~m[1065]&m[1066]&m[1067])|(m[488]&~m[1063]&~m[1065]&m[1066]&m[1067])|(~m[488]&m[1063]&~m[1065]&m[1066]&m[1067])|(m[488]&m[1063]&~m[1065]&m[1066]&m[1067])|(~m[488]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[488]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[488]&m[1063]&m[1065]&m[1066]&m[1067]));
    m[1069] = (((m[499]&~m[1068]&~m[1070]&~m[1071]&~m[1072])|(~m[499]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(m[499]&m[1068]&~m[1070]&m[1071]&~m[1072])|(m[499]&~m[1068]&m[1070]&m[1071]&~m[1072])|(~m[499]&m[1068]&~m[1070]&~m[1071]&m[1072])|(~m[499]&~m[1068]&m[1070]&~m[1071]&m[1072])|(m[499]&m[1068]&m[1070]&~m[1071]&m[1072])|(~m[499]&m[1068]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[360])|((m[499]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(~m[499]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[499]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[499]&m[1068]&~m[1070]&~m[1071]&m[1072])|(m[499]&~m[1068]&m[1070]&~m[1071]&m[1072])|(~m[499]&~m[1068]&~m[1070]&m[1071]&m[1072])|(m[499]&~m[1068]&~m[1070]&m[1071]&m[1072])|(~m[499]&m[1068]&~m[1070]&m[1071]&m[1072])|(m[499]&m[1068]&~m[1070]&m[1071]&m[1072])|(~m[499]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[499]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[499]&m[1068]&m[1070]&m[1071]&m[1072]));
    m[1074] = (((m[510]&~m[1073]&~m[1075]&~m[1076]&~m[1077])|(~m[510]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(m[510]&m[1073]&~m[1075]&m[1076]&~m[1077])|(m[510]&~m[1073]&m[1075]&m[1076]&~m[1077])|(~m[510]&m[1073]&~m[1075]&~m[1076]&m[1077])|(~m[510]&~m[1073]&m[1075]&~m[1076]&m[1077])|(m[510]&m[1073]&m[1075]&~m[1076]&m[1077])|(~m[510]&m[1073]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[361])|((m[510]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(~m[510]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[510]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[510]&m[1073]&~m[1075]&~m[1076]&m[1077])|(m[510]&~m[1073]&m[1075]&~m[1076]&m[1077])|(~m[510]&~m[1073]&~m[1075]&m[1076]&m[1077])|(m[510]&~m[1073]&~m[1075]&m[1076]&m[1077])|(~m[510]&m[1073]&~m[1075]&m[1076]&m[1077])|(m[510]&m[1073]&~m[1075]&m[1076]&m[1077])|(~m[510]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[510]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[510]&m[1073]&m[1075]&m[1076]&m[1077]));
    m[1079] = (((m[521]&~m[1078]&~m[1080]&~m[1081]&~m[1082])|(~m[521]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(m[521]&m[1078]&~m[1080]&m[1081]&~m[1082])|(m[521]&~m[1078]&m[1080]&m[1081]&~m[1082])|(~m[521]&m[1078]&~m[1080]&~m[1081]&m[1082])|(~m[521]&~m[1078]&m[1080]&~m[1081]&m[1082])|(m[521]&m[1078]&m[1080]&~m[1081]&m[1082])|(~m[521]&m[1078]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[362])|((m[521]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(~m[521]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[521]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[521]&m[1078]&~m[1080]&~m[1081]&m[1082])|(m[521]&~m[1078]&m[1080]&~m[1081]&m[1082])|(~m[521]&~m[1078]&~m[1080]&m[1081]&m[1082])|(m[521]&~m[1078]&~m[1080]&m[1081]&m[1082])|(~m[521]&m[1078]&~m[1080]&m[1081]&m[1082])|(m[521]&m[1078]&~m[1080]&m[1081]&m[1082])|(~m[521]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[521]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[521]&m[1078]&m[1080]&m[1081]&m[1082]));
    m[1084] = (((m[467]&~m[1083]&~m[1085]&~m[1086]&~m[1087])|(~m[467]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(m[467]&m[1083]&~m[1085]&m[1086]&~m[1087])|(m[467]&~m[1083]&m[1085]&m[1086]&~m[1087])|(~m[467]&m[1083]&~m[1085]&~m[1086]&m[1087])|(~m[467]&~m[1083]&m[1085]&~m[1086]&m[1087])|(m[467]&m[1083]&m[1085]&~m[1086]&m[1087])|(~m[467]&m[1083]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[363])|((m[467]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(~m[467]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[467]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[467]&m[1083]&~m[1085]&~m[1086]&m[1087])|(m[467]&~m[1083]&m[1085]&~m[1086]&m[1087])|(~m[467]&~m[1083]&~m[1085]&m[1086]&m[1087])|(m[467]&~m[1083]&~m[1085]&m[1086]&m[1087])|(~m[467]&m[1083]&~m[1085]&m[1086]&m[1087])|(m[467]&m[1083]&~m[1085]&m[1086]&m[1087])|(~m[467]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[467]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[467]&m[1083]&m[1085]&m[1086]&m[1087]));
    m[1089] = (((m[478]&~m[1088]&~m[1090]&~m[1091]&~m[1092])|(~m[478]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(m[478]&m[1088]&~m[1090]&m[1091]&~m[1092])|(m[478]&~m[1088]&m[1090]&m[1091]&~m[1092])|(~m[478]&m[1088]&~m[1090]&~m[1091]&m[1092])|(~m[478]&~m[1088]&m[1090]&~m[1091]&m[1092])|(m[478]&m[1088]&m[1090]&~m[1091]&m[1092])|(~m[478]&m[1088]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[364])|((m[478]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(~m[478]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[478]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[478]&m[1088]&~m[1090]&~m[1091]&m[1092])|(m[478]&~m[1088]&m[1090]&~m[1091]&m[1092])|(~m[478]&~m[1088]&~m[1090]&m[1091]&m[1092])|(m[478]&~m[1088]&~m[1090]&m[1091]&m[1092])|(~m[478]&m[1088]&~m[1090]&m[1091]&m[1092])|(m[478]&m[1088]&~m[1090]&m[1091]&m[1092])|(~m[478]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[478]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[478]&m[1088]&m[1090]&m[1091]&m[1092]));
    m[1094] = (((m[489]&~m[1093]&~m[1095]&~m[1096]&~m[1097])|(~m[489]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(m[489]&m[1093]&~m[1095]&m[1096]&~m[1097])|(m[489]&~m[1093]&m[1095]&m[1096]&~m[1097])|(~m[489]&m[1093]&~m[1095]&~m[1096]&m[1097])|(~m[489]&~m[1093]&m[1095]&~m[1096]&m[1097])|(m[489]&m[1093]&m[1095]&~m[1096]&m[1097])|(~m[489]&m[1093]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[365])|((m[489]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(~m[489]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[489]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[489]&m[1093]&~m[1095]&~m[1096]&m[1097])|(m[489]&~m[1093]&m[1095]&~m[1096]&m[1097])|(~m[489]&~m[1093]&~m[1095]&m[1096]&m[1097])|(m[489]&~m[1093]&~m[1095]&m[1096]&m[1097])|(~m[489]&m[1093]&~m[1095]&m[1096]&m[1097])|(m[489]&m[1093]&~m[1095]&m[1096]&m[1097])|(~m[489]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[489]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[489]&m[1093]&m[1095]&m[1096]&m[1097]));
    m[1099] = (((m[500]&~m[1098]&~m[1100]&~m[1101]&~m[1102])|(~m[500]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(m[500]&m[1098]&~m[1100]&m[1101]&~m[1102])|(m[500]&~m[1098]&m[1100]&m[1101]&~m[1102])|(~m[500]&m[1098]&~m[1100]&~m[1101]&m[1102])|(~m[500]&~m[1098]&m[1100]&~m[1101]&m[1102])|(m[500]&m[1098]&m[1100]&~m[1101]&m[1102])|(~m[500]&m[1098]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[366])|((m[500]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(~m[500]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[500]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[500]&m[1098]&~m[1100]&~m[1101]&m[1102])|(m[500]&~m[1098]&m[1100]&~m[1101]&m[1102])|(~m[500]&~m[1098]&~m[1100]&m[1101]&m[1102])|(m[500]&~m[1098]&~m[1100]&m[1101]&m[1102])|(~m[500]&m[1098]&~m[1100]&m[1101]&m[1102])|(m[500]&m[1098]&~m[1100]&m[1101]&m[1102])|(~m[500]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[500]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[500]&m[1098]&m[1100]&m[1101]&m[1102]));
    m[1104] = (((m[511]&~m[1103]&~m[1105]&~m[1106]&~m[1107])|(~m[511]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(m[511]&m[1103]&~m[1105]&m[1106]&~m[1107])|(m[511]&~m[1103]&m[1105]&m[1106]&~m[1107])|(~m[511]&m[1103]&~m[1105]&~m[1106]&m[1107])|(~m[511]&~m[1103]&m[1105]&~m[1106]&m[1107])|(m[511]&m[1103]&m[1105]&~m[1106]&m[1107])|(~m[511]&m[1103]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[367])|((m[511]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(~m[511]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[511]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[511]&m[1103]&~m[1105]&~m[1106]&m[1107])|(m[511]&~m[1103]&m[1105]&~m[1106]&m[1107])|(~m[511]&~m[1103]&~m[1105]&m[1106]&m[1107])|(m[511]&~m[1103]&~m[1105]&m[1106]&m[1107])|(~m[511]&m[1103]&~m[1105]&m[1106]&m[1107])|(m[511]&m[1103]&~m[1105]&m[1106]&m[1107])|(~m[511]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[511]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[511]&m[1103]&m[1105]&m[1106]&m[1107]));
    m[1109] = (((m[522]&~m[1108]&~m[1110]&~m[1111]&~m[1112])|(~m[522]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(m[522]&m[1108]&~m[1110]&m[1111]&~m[1112])|(m[522]&~m[1108]&m[1110]&m[1111]&~m[1112])|(~m[522]&m[1108]&~m[1110]&~m[1111]&m[1112])|(~m[522]&~m[1108]&m[1110]&~m[1111]&m[1112])|(m[522]&m[1108]&m[1110]&~m[1111]&m[1112])|(~m[522]&m[1108]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[368])|((m[522]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(~m[522]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[522]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[522]&m[1108]&~m[1110]&~m[1111]&m[1112])|(m[522]&~m[1108]&m[1110]&~m[1111]&m[1112])|(~m[522]&~m[1108]&~m[1110]&m[1111]&m[1112])|(m[522]&~m[1108]&~m[1110]&m[1111]&m[1112])|(~m[522]&m[1108]&~m[1110]&m[1111]&m[1112])|(m[522]&m[1108]&~m[1110]&m[1111]&m[1112])|(~m[522]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[522]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[522]&m[1108]&m[1110]&m[1111]&m[1112]));
    m[1114] = (((m[479]&~m[1113]&~m[1115]&~m[1116]&~m[1117])|(~m[479]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(m[479]&m[1113]&~m[1115]&m[1116]&~m[1117])|(m[479]&~m[1113]&m[1115]&m[1116]&~m[1117])|(~m[479]&m[1113]&~m[1115]&~m[1116]&m[1117])|(~m[479]&~m[1113]&m[1115]&~m[1116]&m[1117])|(m[479]&m[1113]&m[1115]&~m[1116]&m[1117])|(~m[479]&m[1113]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[369])|((m[479]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(~m[479]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[479]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[479]&m[1113]&~m[1115]&~m[1116]&m[1117])|(m[479]&~m[1113]&m[1115]&~m[1116]&m[1117])|(~m[479]&~m[1113]&~m[1115]&m[1116]&m[1117])|(m[479]&~m[1113]&~m[1115]&m[1116]&m[1117])|(~m[479]&m[1113]&~m[1115]&m[1116]&m[1117])|(m[479]&m[1113]&~m[1115]&m[1116]&m[1117])|(~m[479]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[479]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[479]&m[1113]&m[1115]&m[1116]&m[1117]));
    m[1119] = (((m[490]&~m[1118]&~m[1120]&~m[1121]&~m[1122])|(~m[490]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(m[490]&m[1118]&~m[1120]&m[1121]&~m[1122])|(m[490]&~m[1118]&m[1120]&m[1121]&~m[1122])|(~m[490]&m[1118]&~m[1120]&~m[1121]&m[1122])|(~m[490]&~m[1118]&m[1120]&~m[1121]&m[1122])|(m[490]&m[1118]&m[1120]&~m[1121]&m[1122])|(~m[490]&m[1118]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[370])|((m[490]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(~m[490]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[490]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[490]&m[1118]&~m[1120]&~m[1121]&m[1122])|(m[490]&~m[1118]&m[1120]&~m[1121]&m[1122])|(~m[490]&~m[1118]&~m[1120]&m[1121]&m[1122])|(m[490]&~m[1118]&~m[1120]&m[1121]&m[1122])|(~m[490]&m[1118]&~m[1120]&m[1121]&m[1122])|(m[490]&m[1118]&~m[1120]&m[1121]&m[1122])|(~m[490]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[490]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[490]&m[1118]&m[1120]&m[1121]&m[1122]));
    m[1124] = (((m[501]&~m[1123]&~m[1125]&~m[1126]&~m[1127])|(~m[501]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(m[501]&m[1123]&~m[1125]&m[1126]&~m[1127])|(m[501]&~m[1123]&m[1125]&m[1126]&~m[1127])|(~m[501]&m[1123]&~m[1125]&~m[1126]&m[1127])|(~m[501]&~m[1123]&m[1125]&~m[1126]&m[1127])|(m[501]&m[1123]&m[1125]&~m[1126]&m[1127])|(~m[501]&m[1123]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[371])|((m[501]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(~m[501]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[501]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[501]&m[1123]&~m[1125]&~m[1126]&m[1127])|(m[501]&~m[1123]&m[1125]&~m[1126]&m[1127])|(~m[501]&~m[1123]&~m[1125]&m[1126]&m[1127])|(m[501]&~m[1123]&~m[1125]&m[1126]&m[1127])|(~m[501]&m[1123]&~m[1125]&m[1126]&m[1127])|(m[501]&m[1123]&~m[1125]&m[1126]&m[1127])|(~m[501]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[501]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[501]&m[1123]&m[1125]&m[1126]&m[1127]));
    m[1129] = (((m[512]&~m[1128]&~m[1130]&~m[1131]&~m[1132])|(~m[512]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(m[512]&m[1128]&~m[1130]&m[1131]&~m[1132])|(m[512]&~m[1128]&m[1130]&m[1131]&~m[1132])|(~m[512]&m[1128]&~m[1130]&~m[1131]&m[1132])|(~m[512]&~m[1128]&m[1130]&~m[1131]&m[1132])|(m[512]&m[1128]&m[1130]&~m[1131]&m[1132])|(~m[512]&m[1128]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[372])|((m[512]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(~m[512]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[512]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[512]&m[1128]&~m[1130]&~m[1131]&m[1132])|(m[512]&~m[1128]&m[1130]&~m[1131]&m[1132])|(~m[512]&~m[1128]&~m[1130]&m[1131]&m[1132])|(m[512]&~m[1128]&~m[1130]&m[1131]&m[1132])|(~m[512]&m[1128]&~m[1130]&m[1131]&m[1132])|(m[512]&m[1128]&~m[1130]&m[1131]&m[1132])|(~m[512]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[512]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[512]&m[1128]&m[1130]&m[1131]&m[1132]));
    m[1134] = (((m[523]&~m[1133]&~m[1135]&~m[1136]&~m[1137])|(~m[523]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(m[523]&m[1133]&~m[1135]&m[1136]&~m[1137])|(m[523]&~m[1133]&m[1135]&m[1136]&~m[1137])|(~m[523]&m[1133]&~m[1135]&~m[1136]&m[1137])|(~m[523]&~m[1133]&m[1135]&~m[1136]&m[1137])|(m[523]&m[1133]&m[1135]&~m[1136]&m[1137])|(~m[523]&m[1133]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[373])|((m[523]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(~m[523]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[523]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[523]&m[1133]&~m[1135]&~m[1136]&m[1137])|(m[523]&~m[1133]&m[1135]&~m[1136]&m[1137])|(~m[523]&~m[1133]&~m[1135]&m[1136]&m[1137])|(m[523]&~m[1133]&~m[1135]&m[1136]&m[1137])|(~m[523]&m[1133]&~m[1135]&m[1136]&m[1137])|(m[523]&m[1133]&~m[1135]&m[1136]&m[1137])|(~m[523]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[523]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[523]&m[1133]&m[1135]&m[1136]&m[1137]));
    m[1139] = (((m[491]&~m[1138]&~m[1140]&~m[1141]&~m[1142])|(~m[491]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(m[491]&m[1138]&~m[1140]&m[1141]&~m[1142])|(m[491]&~m[1138]&m[1140]&m[1141]&~m[1142])|(~m[491]&m[1138]&~m[1140]&~m[1141]&m[1142])|(~m[491]&~m[1138]&m[1140]&~m[1141]&m[1142])|(m[491]&m[1138]&m[1140]&~m[1141]&m[1142])|(~m[491]&m[1138]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[374])|((m[491]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(~m[491]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[491]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[491]&m[1138]&~m[1140]&~m[1141]&m[1142])|(m[491]&~m[1138]&m[1140]&~m[1141]&m[1142])|(~m[491]&~m[1138]&~m[1140]&m[1141]&m[1142])|(m[491]&~m[1138]&~m[1140]&m[1141]&m[1142])|(~m[491]&m[1138]&~m[1140]&m[1141]&m[1142])|(m[491]&m[1138]&~m[1140]&m[1141]&m[1142])|(~m[491]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[491]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[491]&m[1138]&m[1140]&m[1141]&m[1142]));
    m[1144] = (((m[502]&~m[1143]&~m[1145]&~m[1146]&~m[1147])|(~m[502]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(m[502]&m[1143]&~m[1145]&m[1146]&~m[1147])|(m[502]&~m[1143]&m[1145]&m[1146]&~m[1147])|(~m[502]&m[1143]&~m[1145]&~m[1146]&m[1147])|(~m[502]&~m[1143]&m[1145]&~m[1146]&m[1147])|(m[502]&m[1143]&m[1145]&~m[1146]&m[1147])|(~m[502]&m[1143]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[375])|((m[502]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(~m[502]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[502]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[502]&m[1143]&~m[1145]&~m[1146]&m[1147])|(m[502]&~m[1143]&m[1145]&~m[1146]&m[1147])|(~m[502]&~m[1143]&~m[1145]&m[1146]&m[1147])|(m[502]&~m[1143]&~m[1145]&m[1146]&m[1147])|(~m[502]&m[1143]&~m[1145]&m[1146]&m[1147])|(m[502]&m[1143]&~m[1145]&m[1146]&m[1147])|(~m[502]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[502]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[502]&m[1143]&m[1145]&m[1146]&m[1147]));
    m[1149] = (((m[513]&~m[1148]&~m[1150]&~m[1151]&~m[1152])|(~m[513]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(m[513]&m[1148]&~m[1150]&m[1151]&~m[1152])|(m[513]&~m[1148]&m[1150]&m[1151]&~m[1152])|(~m[513]&m[1148]&~m[1150]&~m[1151]&m[1152])|(~m[513]&~m[1148]&m[1150]&~m[1151]&m[1152])|(m[513]&m[1148]&m[1150]&~m[1151]&m[1152])|(~m[513]&m[1148]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[376])|((m[513]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(~m[513]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[513]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[513]&m[1148]&~m[1150]&~m[1151]&m[1152])|(m[513]&~m[1148]&m[1150]&~m[1151]&m[1152])|(~m[513]&~m[1148]&~m[1150]&m[1151]&m[1152])|(m[513]&~m[1148]&~m[1150]&m[1151]&m[1152])|(~m[513]&m[1148]&~m[1150]&m[1151]&m[1152])|(m[513]&m[1148]&~m[1150]&m[1151]&m[1152])|(~m[513]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[513]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[513]&m[1148]&m[1150]&m[1151]&m[1152]));
    m[1154] = (((m[524]&~m[1153]&~m[1155]&~m[1156]&~m[1157])|(~m[524]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(m[524]&m[1153]&~m[1155]&m[1156]&~m[1157])|(m[524]&~m[1153]&m[1155]&m[1156]&~m[1157])|(~m[524]&m[1153]&~m[1155]&~m[1156]&m[1157])|(~m[524]&~m[1153]&m[1155]&~m[1156]&m[1157])|(m[524]&m[1153]&m[1155]&~m[1156]&m[1157])|(~m[524]&m[1153]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[377])|((m[524]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(~m[524]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[524]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[524]&m[1153]&~m[1155]&~m[1156]&m[1157])|(m[524]&~m[1153]&m[1155]&~m[1156]&m[1157])|(~m[524]&~m[1153]&~m[1155]&m[1156]&m[1157])|(m[524]&~m[1153]&~m[1155]&m[1156]&m[1157])|(~m[524]&m[1153]&~m[1155]&m[1156]&m[1157])|(m[524]&m[1153]&~m[1155]&m[1156]&m[1157])|(~m[524]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[524]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[524]&m[1153]&m[1155]&m[1156]&m[1157]));
    m[1159] = (((m[503]&~m[1158]&~m[1160]&~m[1161]&~m[1162])|(~m[503]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(m[503]&m[1158]&~m[1160]&m[1161]&~m[1162])|(m[503]&~m[1158]&m[1160]&m[1161]&~m[1162])|(~m[503]&m[1158]&~m[1160]&~m[1161]&m[1162])|(~m[503]&~m[1158]&m[1160]&~m[1161]&m[1162])|(m[503]&m[1158]&m[1160]&~m[1161]&m[1162])|(~m[503]&m[1158]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[378])|((m[503]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(~m[503]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[503]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[503]&m[1158]&~m[1160]&~m[1161]&m[1162])|(m[503]&~m[1158]&m[1160]&~m[1161]&m[1162])|(~m[503]&~m[1158]&~m[1160]&m[1161]&m[1162])|(m[503]&~m[1158]&~m[1160]&m[1161]&m[1162])|(~m[503]&m[1158]&~m[1160]&m[1161]&m[1162])|(m[503]&m[1158]&~m[1160]&m[1161]&m[1162])|(~m[503]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[503]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[503]&m[1158]&m[1160]&m[1161]&m[1162]));
    m[1164] = (((m[514]&~m[1163]&~m[1165]&~m[1166]&~m[1167])|(~m[514]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(m[514]&m[1163]&~m[1165]&m[1166]&~m[1167])|(m[514]&~m[1163]&m[1165]&m[1166]&~m[1167])|(~m[514]&m[1163]&~m[1165]&~m[1166]&m[1167])|(~m[514]&~m[1163]&m[1165]&~m[1166]&m[1167])|(m[514]&m[1163]&m[1165]&~m[1166]&m[1167])|(~m[514]&m[1163]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[379])|((m[514]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(~m[514]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[514]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[514]&m[1163]&~m[1165]&~m[1166]&m[1167])|(m[514]&~m[1163]&m[1165]&~m[1166]&m[1167])|(~m[514]&~m[1163]&~m[1165]&m[1166]&m[1167])|(m[514]&~m[1163]&~m[1165]&m[1166]&m[1167])|(~m[514]&m[1163]&~m[1165]&m[1166]&m[1167])|(m[514]&m[1163]&~m[1165]&m[1166]&m[1167])|(~m[514]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[514]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[514]&m[1163]&m[1165]&m[1166]&m[1167]));
    m[1169] = (((m[525]&~m[1168]&~m[1170]&~m[1171]&~m[1172])|(~m[525]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(m[525]&m[1168]&~m[1170]&m[1171]&~m[1172])|(m[525]&~m[1168]&m[1170]&m[1171]&~m[1172])|(~m[525]&m[1168]&~m[1170]&~m[1171]&m[1172])|(~m[525]&~m[1168]&m[1170]&~m[1171]&m[1172])|(m[525]&m[1168]&m[1170]&~m[1171]&m[1172])|(~m[525]&m[1168]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[380])|((m[525]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(~m[525]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[525]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[525]&m[1168]&~m[1170]&~m[1171]&m[1172])|(m[525]&~m[1168]&m[1170]&~m[1171]&m[1172])|(~m[525]&~m[1168]&~m[1170]&m[1171]&m[1172])|(m[525]&~m[1168]&~m[1170]&m[1171]&m[1172])|(~m[525]&m[1168]&~m[1170]&m[1171]&m[1172])|(m[525]&m[1168]&~m[1170]&m[1171]&m[1172])|(~m[525]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[525]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[525]&m[1168]&m[1170]&m[1171]&m[1172]));
    m[1174] = (((m[515]&~m[1173]&~m[1175]&~m[1176]&~m[1177])|(~m[515]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(m[515]&m[1173]&~m[1175]&m[1176]&~m[1177])|(m[515]&~m[1173]&m[1175]&m[1176]&~m[1177])|(~m[515]&m[1173]&~m[1175]&~m[1176]&m[1177])|(~m[515]&~m[1173]&m[1175]&~m[1176]&m[1177])|(m[515]&m[1173]&m[1175]&~m[1176]&m[1177])|(~m[515]&m[1173]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[381])|((m[515]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(~m[515]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[515]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[515]&m[1173]&~m[1175]&~m[1176]&m[1177])|(m[515]&~m[1173]&m[1175]&~m[1176]&m[1177])|(~m[515]&~m[1173]&~m[1175]&m[1176]&m[1177])|(m[515]&~m[1173]&~m[1175]&m[1176]&m[1177])|(~m[515]&m[1173]&~m[1175]&m[1176]&m[1177])|(m[515]&m[1173]&~m[1175]&m[1176]&m[1177])|(~m[515]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[515]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[515]&m[1173]&m[1175]&m[1176]&m[1177]));
    m[1179] = (((m[526]&~m[1178]&~m[1180]&~m[1181]&~m[1182])|(~m[526]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(m[526]&m[1178]&~m[1180]&m[1181]&~m[1182])|(m[526]&~m[1178]&m[1180]&m[1181]&~m[1182])|(~m[526]&m[1178]&~m[1180]&~m[1181]&m[1182])|(~m[526]&~m[1178]&m[1180]&~m[1181]&m[1182])|(m[526]&m[1178]&m[1180]&~m[1181]&m[1182])|(~m[526]&m[1178]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[382])|((m[526]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(~m[526]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[526]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[526]&m[1178]&~m[1180]&~m[1181]&m[1182])|(m[526]&~m[1178]&m[1180]&~m[1181]&m[1182])|(~m[526]&~m[1178]&~m[1180]&m[1181]&m[1182])|(m[526]&~m[1178]&~m[1180]&m[1181]&m[1182])|(~m[526]&m[1178]&~m[1180]&m[1181]&m[1182])|(m[526]&m[1178]&~m[1180]&m[1181]&m[1182])|(~m[526]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[526]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[526]&m[1178]&m[1180]&m[1181]&m[1182]));
    m[1184] = (((m[527]&~m[1183]&~m[1185]&~m[1186]&~m[1187])|(~m[527]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(m[527]&m[1183]&~m[1185]&m[1186]&~m[1187])|(m[527]&~m[1183]&m[1185]&m[1186]&~m[1187])|(~m[527]&m[1183]&~m[1185]&~m[1186]&m[1187])|(~m[527]&~m[1183]&m[1185]&~m[1186]&m[1187])|(m[527]&m[1183]&m[1185]&~m[1186]&m[1187])|(~m[527]&m[1183]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[383])|((m[527]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(~m[527]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[527]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[527]&m[1183]&~m[1185]&~m[1186]&m[1187])|(m[527]&~m[1183]&m[1185]&~m[1186]&m[1187])|(~m[527]&~m[1183]&~m[1185]&m[1186]&m[1187])|(m[527]&~m[1183]&~m[1185]&m[1186]&m[1187])|(~m[527]&m[1183]&~m[1185]&m[1186]&m[1187])|(m[527]&m[1183]&~m[1185]&m[1186]&m[1187])|(~m[527]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[527]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[527]&m[1183]&m[1185]&m[1186]&m[1187]));
end

always @(posedge color3_clk) begin
    m[536] = (((m[533]&~m[534]&~m[535]&~m[537]&~m[538])|(~m[533]&m[534]&~m[535]&~m[537]&~m[538])|(~m[533]&~m[534]&m[535]&~m[537]&~m[538])|(m[533]&m[534]&m[535]&m[537]&~m[538])|(~m[533]&~m[534]&~m[535]&~m[537]&m[538])|(m[533]&m[534]&~m[535]&m[537]&m[538])|(m[533]&~m[534]&m[535]&m[537]&m[538])|(~m[533]&m[534]&m[535]&m[537]&m[538]))&UnbiasedRNG[384])|((m[533]&m[534]&~m[535]&~m[537]&~m[538])|(m[533]&~m[534]&m[535]&~m[537]&~m[538])|(~m[533]&m[534]&m[535]&~m[537]&~m[538])|(m[533]&m[534]&m[535]&~m[537]&~m[538])|(m[533]&~m[534]&~m[535]&~m[537]&m[538])|(~m[533]&m[534]&~m[535]&~m[537]&m[538])|(m[533]&m[534]&~m[535]&~m[537]&m[538])|(~m[533]&~m[534]&m[535]&~m[537]&m[538])|(m[533]&~m[534]&m[535]&~m[537]&m[538])|(~m[533]&m[534]&m[535]&~m[537]&m[538])|(m[533]&m[534]&m[535]&~m[537]&m[538])|(m[533]&m[534]&m[535]&m[537]&m[538]));
    m[546] = (((m[543]&~m[544]&~m[545]&~m[547]&~m[548])|(~m[543]&m[544]&~m[545]&~m[547]&~m[548])|(~m[543]&~m[544]&m[545]&~m[547]&~m[548])|(m[543]&m[544]&m[545]&m[547]&~m[548])|(~m[543]&~m[544]&~m[545]&~m[547]&m[548])|(m[543]&m[544]&~m[545]&m[547]&m[548])|(m[543]&~m[544]&m[545]&m[547]&m[548])|(~m[543]&m[544]&m[545]&m[547]&m[548]))&UnbiasedRNG[385])|((m[543]&m[544]&~m[545]&~m[547]&~m[548])|(m[543]&~m[544]&m[545]&~m[547]&~m[548])|(~m[543]&m[544]&m[545]&~m[547]&~m[548])|(m[543]&m[544]&m[545]&~m[547]&~m[548])|(m[543]&~m[544]&~m[545]&~m[547]&m[548])|(~m[543]&m[544]&~m[545]&~m[547]&m[548])|(m[543]&m[544]&~m[545]&~m[547]&m[548])|(~m[543]&~m[544]&m[545]&~m[547]&m[548])|(m[543]&~m[544]&m[545]&~m[547]&m[548])|(~m[543]&m[544]&m[545]&~m[547]&m[548])|(m[543]&m[544]&m[545]&~m[547]&m[548])|(m[543]&m[544]&m[545]&m[547]&m[548]));
    m[551] = (((m[548]&~m[549]&~m[550]&~m[552]&~m[553])|(~m[548]&m[549]&~m[550]&~m[552]&~m[553])|(~m[548]&~m[549]&m[550]&~m[552]&~m[553])|(m[548]&m[549]&m[550]&m[552]&~m[553])|(~m[548]&~m[549]&~m[550]&~m[552]&m[553])|(m[548]&m[549]&~m[550]&m[552]&m[553])|(m[548]&~m[549]&m[550]&m[552]&m[553])|(~m[548]&m[549]&m[550]&m[552]&m[553]))&UnbiasedRNG[386])|((m[548]&m[549]&~m[550]&~m[552]&~m[553])|(m[548]&~m[549]&m[550]&~m[552]&~m[553])|(~m[548]&m[549]&m[550]&~m[552]&~m[553])|(m[548]&m[549]&m[550]&~m[552]&~m[553])|(m[548]&~m[549]&~m[550]&~m[552]&m[553])|(~m[548]&m[549]&~m[550]&~m[552]&m[553])|(m[548]&m[549]&~m[550]&~m[552]&m[553])|(~m[548]&~m[549]&m[550]&~m[552]&m[553])|(m[548]&~m[549]&m[550]&~m[552]&m[553])|(~m[548]&m[549]&m[550]&~m[552]&m[553])|(m[548]&m[549]&m[550]&~m[552]&m[553])|(m[548]&m[549]&m[550]&m[552]&m[553]));
    m[561] = (((m[558]&~m[559]&~m[560]&~m[562]&~m[563])|(~m[558]&m[559]&~m[560]&~m[562]&~m[563])|(~m[558]&~m[559]&m[560]&~m[562]&~m[563])|(m[558]&m[559]&m[560]&m[562]&~m[563])|(~m[558]&~m[559]&~m[560]&~m[562]&m[563])|(m[558]&m[559]&~m[560]&m[562]&m[563])|(m[558]&~m[559]&m[560]&m[562]&m[563])|(~m[558]&m[559]&m[560]&m[562]&m[563]))&UnbiasedRNG[387])|((m[558]&m[559]&~m[560]&~m[562]&~m[563])|(m[558]&~m[559]&m[560]&~m[562]&~m[563])|(~m[558]&m[559]&m[560]&~m[562]&~m[563])|(m[558]&m[559]&m[560]&~m[562]&~m[563])|(m[558]&~m[559]&~m[560]&~m[562]&m[563])|(~m[558]&m[559]&~m[560]&~m[562]&m[563])|(m[558]&m[559]&~m[560]&~m[562]&m[563])|(~m[558]&~m[559]&m[560]&~m[562]&m[563])|(m[558]&~m[559]&m[560]&~m[562]&m[563])|(~m[558]&m[559]&m[560]&~m[562]&m[563])|(m[558]&m[559]&m[560]&~m[562]&m[563])|(m[558]&m[559]&m[560]&m[562]&m[563]));
    m[566] = (((m[563]&~m[564]&~m[565]&~m[567]&~m[568])|(~m[563]&m[564]&~m[565]&~m[567]&~m[568])|(~m[563]&~m[564]&m[565]&~m[567]&~m[568])|(m[563]&m[564]&m[565]&m[567]&~m[568])|(~m[563]&~m[564]&~m[565]&~m[567]&m[568])|(m[563]&m[564]&~m[565]&m[567]&m[568])|(m[563]&~m[564]&m[565]&m[567]&m[568])|(~m[563]&m[564]&m[565]&m[567]&m[568]))&UnbiasedRNG[388])|((m[563]&m[564]&~m[565]&~m[567]&~m[568])|(m[563]&~m[564]&m[565]&~m[567]&~m[568])|(~m[563]&m[564]&m[565]&~m[567]&~m[568])|(m[563]&m[564]&m[565]&~m[567]&~m[568])|(m[563]&~m[564]&~m[565]&~m[567]&m[568])|(~m[563]&m[564]&~m[565]&~m[567]&m[568])|(m[563]&m[564]&~m[565]&~m[567]&m[568])|(~m[563]&~m[564]&m[565]&~m[567]&m[568])|(m[563]&~m[564]&m[565]&~m[567]&m[568])|(~m[563]&m[564]&m[565]&~m[567]&m[568])|(m[563]&m[564]&m[565]&~m[567]&m[568])|(m[563]&m[564]&m[565]&m[567]&m[568]));
    m[571] = (((m[568]&~m[569]&~m[570]&~m[572]&~m[573])|(~m[568]&m[569]&~m[570]&~m[572]&~m[573])|(~m[568]&~m[569]&m[570]&~m[572]&~m[573])|(m[568]&m[569]&m[570]&m[572]&~m[573])|(~m[568]&~m[569]&~m[570]&~m[572]&m[573])|(m[568]&m[569]&~m[570]&m[572]&m[573])|(m[568]&~m[569]&m[570]&m[572]&m[573])|(~m[568]&m[569]&m[570]&m[572]&m[573]))&UnbiasedRNG[389])|((m[568]&m[569]&~m[570]&~m[572]&~m[573])|(m[568]&~m[569]&m[570]&~m[572]&~m[573])|(~m[568]&m[569]&m[570]&~m[572]&~m[573])|(m[568]&m[569]&m[570]&~m[572]&~m[573])|(m[568]&~m[569]&~m[570]&~m[572]&m[573])|(~m[568]&m[569]&~m[570]&~m[572]&m[573])|(m[568]&m[569]&~m[570]&~m[572]&m[573])|(~m[568]&~m[569]&m[570]&~m[572]&m[573])|(m[568]&~m[569]&m[570]&~m[572]&m[573])|(~m[568]&m[569]&m[570]&~m[572]&m[573])|(m[568]&m[569]&m[570]&~m[572]&m[573])|(m[568]&m[569]&m[570]&m[572]&m[573]));
    m[581] = (((m[578]&~m[579]&~m[580]&~m[582]&~m[583])|(~m[578]&m[579]&~m[580]&~m[582]&~m[583])|(~m[578]&~m[579]&m[580]&~m[582]&~m[583])|(m[578]&m[579]&m[580]&m[582]&~m[583])|(~m[578]&~m[579]&~m[580]&~m[582]&m[583])|(m[578]&m[579]&~m[580]&m[582]&m[583])|(m[578]&~m[579]&m[580]&m[582]&m[583])|(~m[578]&m[579]&m[580]&m[582]&m[583]))&UnbiasedRNG[390])|((m[578]&m[579]&~m[580]&~m[582]&~m[583])|(m[578]&~m[579]&m[580]&~m[582]&~m[583])|(~m[578]&m[579]&m[580]&~m[582]&~m[583])|(m[578]&m[579]&m[580]&~m[582]&~m[583])|(m[578]&~m[579]&~m[580]&~m[582]&m[583])|(~m[578]&m[579]&~m[580]&~m[582]&m[583])|(m[578]&m[579]&~m[580]&~m[582]&m[583])|(~m[578]&~m[579]&m[580]&~m[582]&m[583])|(m[578]&~m[579]&m[580]&~m[582]&m[583])|(~m[578]&m[579]&m[580]&~m[582]&m[583])|(m[578]&m[579]&m[580]&~m[582]&m[583])|(m[578]&m[579]&m[580]&m[582]&m[583]));
    m[586] = (((m[583]&~m[584]&~m[585]&~m[587]&~m[588])|(~m[583]&m[584]&~m[585]&~m[587]&~m[588])|(~m[583]&~m[584]&m[585]&~m[587]&~m[588])|(m[583]&m[584]&m[585]&m[587]&~m[588])|(~m[583]&~m[584]&~m[585]&~m[587]&m[588])|(m[583]&m[584]&~m[585]&m[587]&m[588])|(m[583]&~m[584]&m[585]&m[587]&m[588])|(~m[583]&m[584]&m[585]&m[587]&m[588]))&UnbiasedRNG[391])|((m[583]&m[584]&~m[585]&~m[587]&~m[588])|(m[583]&~m[584]&m[585]&~m[587]&~m[588])|(~m[583]&m[584]&m[585]&~m[587]&~m[588])|(m[583]&m[584]&m[585]&~m[587]&~m[588])|(m[583]&~m[584]&~m[585]&~m[587]&m[588])|(~m[583]&m[584]&~m[585]&~m[587]&m[588])|(m[583]&m[584]&~m[585]&~m[587]&m[588])|(~m[583]&~m[584]&m[585]&~m[587]&m[588])|(m[583]&~m[584]&m[585]&~m[587]&m[588])|(~m[583]&m[584]&m[585]&~m[587]&m[588])|(m[583]&m[584]&m[585]&~m[587]&m[588])|(m[583]&m[584]&m[585]&m[587]&m[588]));
    m[591] = (((m[588]&~m[589]&~m[590]&~m[592]&~m[593])|(~m[588]&m[589]&~m[590]&~m[592]&~m[593])|(~m[588]&~m[589]&m[590]&~m[592]&~m[593])|(m[588]&m[589]&m[590]&m[592]&~m[593])|(~m[588]&~m[589]&~m[590]&~m[592]&m[593])|(m[588]&m[589]&~m[590]&m[592]&m[593])|(m[588]&~m[589]&m[590]&m[592]&m[593])|(~m[588]&m[589]&m[590]&m[592]&m[593]))&UnbiasedRNG[392])|((m[588]&m[589]&~m[590]&~m[592]&~m[593])|(m[588]&~m[589]&m[590]&~m[592]&~m[593])|(~m[588]&m[589]&m[590]&~m[592]&~m[593])|(m[588]&m[589]&m[590]&~m[592]&~m[593])|(m[588]&~m[589]&~m[590]&~m[592]&m[593])|(~m[588]&m[589]&~m[590]&~m[592]&m[593])|(m[588]&m[589]&~m[590]&~m[592]&m[593])|(~m[588]&~m[589]&m[590]&~m[592]&m[593])|(m[588]&~m[589]&m[590]&~m[592]&m[593])|(~m[588]&m[589]&m[590]&~m[592]&m[593])|(m[588]&m[589]&m[590]&~m[592]&m[593])|(m[588]&m[589]&m[590]&m[592]&m[593]));
    m[596] = (((m[593]&~m[594]&~m[595]&~m[597]&~m[598])|(~m[593]&m[594]&~m[595]&~m[597]&~m[598])|(~m[593]&~m[594]&m[595]&~m[597]&~m[598])|(m[593]&m[594]&m[595]&m[597]&~m[598])|(~m[593]&~m[594]&~m[595]&~m[597]&m[598])|(m[593]&m[594]&~m[595]&m[597]&m[598])|(m[593]&~m[594]&m[595]&m[597]&m[598])|(~m[593]&m[594]&m[595]&m[597]&m[598]))&UnbiasedRNG[393])|((m[593]&m[594]&~m[595]&~m[597]&~m[598])|(m[593]&~m[594]&m[595]&~m[597]&~m[598])|(~m[593]&m[594]&m[595]&~m[597]&~m[598])|(m[593]&m[594]&m[595]&~m[597]&~m[598])|(m[593]&~m[594]&~m[595]&~m[597]&m[598])|(~m[593]&m[594]&~m[595]&~m[597]&m[598])|(m[593]&m[594]&~m[595]&~m[597]&m[598])|(~m[593]&~m[594]&m[595]&~m[597]&m[598])|(m[593]&~m[594]&m[595]&~m[597]&m[598])|(~m[593]&m[594]&m[595]&~m[597]&m[598])|(m[593]&m[594]&m[595]&~m[597]&m[598])|(m[593]&m[594]&m[595]&m[597]&m[598]));
    m[606] = (((m[603]&~m[604]&~m[605]&~m[607]&~m[608])|(~m[603]&m[604]&~m[605]&~m[607]&~m[608])|(~m[603]&~m[604]&m[605]&~m[607]&~m[608])|(m[603]&m[604]&m[605]&m[607]&~m[608])|(~m[603]&~m[604]&~m[605]&~m[607]&m[608])|(m[603]&m[604]&~m[605]&m[607]&m[608])|(m[603]&~m[604]&m[605]&m[607]&m[608])|(~m[603]&m[604]&m[605]&m[607]&m[608]))&UnbiasedRNG[394])|((m[603]&m[604]&~m[605]&~m[607]&~m[608])|(m[603]&~m[604]&m[605]&~m[607]&~m[608])|(~m[603]&m[604]&m[605]&~m[607]&~m[608])|(m[603]&m[604]&m[605]&~m[607]&~m[608])|(m[603]&~m[604]&~m[605]&~m[607]&m[608])|(~m[603]&m[604]&~m[605]&~m[607]&m[608])|(m[603]&m[604]&~m[605]&~m[607]&m[608])|(~m[603]&~m[604]&m[605]&~m[607]&m[608])|(m[603]&~m[604]&m[605]&~m[607]&m[608])|(~m[603]&m[604]&m[605]&~m[607]&m[608])|(m[603]&m[604]&m[605]&~m[607]&m[608])|(m[603]&m[604]&m[605]&m[607]&m[608]));
    m[611] = (((m[608]&~m[609]&~m[610]&~m[612]&~m[613])|(~m[608]&m[609]&~m[610]&~m[612]&~m[613])|(~m[608]&~m[609]&m[610]&~m[612]&~m[613])|(m[608]&m[609]&m[610]&m[612]&~m[613])|(~m[608]&~m[609]&~m[610]&~m[612]&m[613])|(m[608]&m[609]&~m[610]&m[612]&m[613])|(m[608]&~m[609]&m[610]&m[612]&m[613])|(~m[608]&m[609]&m[610]&m[612]&m[613]))&UnbiasedRNG[395])|((m[608]&m[609]&~m[610]&~m[612]&~m[613])|(m[608]&~m[609]&m[610]&~m[612]&~m[613])|(~m[608]&m[609]&m[610]&~m[612]&~m[613])|(m[608]&m[609]&m[610]&~m[612]&~m[613])|(m[608]&~m[609]&~m[610]&~m[612]&m[613])|(~m[608]&m[609]&~m[610]&~m[612]&m[613])|(m[608]&m[609]&~m[610]&~m[612]&m[613])|(~m[608]&~m[609]&m[610]&~m[612]&m[613])|(m[608]&~m[609]&m[610]&~m[612]&m[613])|(~m[608]&m[609]&m[610]&~m[612]&m[613])|(m[608]&m[609]&m[610]&~m[612]&m[613])|(m[608]&m[609]&m[610]&m[612]&m[613]));
    m[616] = (((m[613]&~m[614]&~m[615]&~m[617]&~m[618])|(~m[613]&m[614]&~m[615]&~m[617]&~m[618])|(~m[613]&~m[614]&m[615]&~m[617]&~m[618])|(m[613]&m[614]&m[615]&m[617]&~m[618])|(~m[613]&~m[614]&~m[615]&~m[617]&m[618])|(m[613]&m[614]&~m[615]&m[617]&m[618])|(m[613]&~m[614]&m[615]&m[617]&m[618])|(~m[613]&m[614]&m[615]&m[617]&m[618]))&UnbiasedRNG[396])|((m[613]&m[614]&~m[615]&~m[617]&~m[618])|(m[613]&~m[614]&m[615]&~m[617]&~m[618])|(~m[613]&m[614]&m[615]&~m[617]&~m[618])|(m[613]&m[614]&m[615]&~m[617]&~m[618])|(m[613]&~m[614]&~m[615]&~m[617]&m[618])|(~m[613]&m[614]&~m[615]&~m[617]&m[618])|(m[613]&m[614]&~m[615]&~m[617]&m[618])|(~m[613]&~m[614]&m[615]&~m[617]&m[618])|(m[613]&~m[614]&m[615]&~m[617]&m[618])|(~m[613]&m[614]&m[615]&~m[617]&m[618])|(m[613]&m[614]&m[615]&~m[617]&m[618])|(m[613]&m[614]&m[615]&m[617]&m[618]));
    m[621] = (((m[618]&~m[619]&~m[620]&~m[622]&~m[623])|(~m[618]&m[619]&~m[620]&~m[622]&~m[623])|(~m[618]&~m[619]&m[620]&~m[622]&~m[623])|(m[618]&m[619]&m[620]&m[622]&~m[623])|(~m[618]&~m[619]&~m[620]&~m[622]&m[623])|(m[618]&m[619]&~m[620]&m[622]&m[623])|(m[618]&~m[619]&m[620]&m[622]&m[623])|(~m[618]&m[619]&m[620]&m[622]&m[623]))&UnbiasedRNG[397])|((m[618]&m[619]&~m[620]&~m[622]&~m[623])|(m[618]&~m[619]&m[620]&~m[622]&~m[623])|(~m[618]&m[619]&m[620]&~m[622]&~m[623])|(m[618]&m[619]&m[620]&~m[622]&~m[623])|(m[618]&~m[619]&~m[620]&~m[622]&m[623])|(~m[618]&m[619]&~m[620]&~m[622]&m[623])|(m[618]&m[619]&~m[620]&~m[622]&m[623])|(~m[618]&~m[619]&m[620]&~m[622]&m[623])|(m[618]&~m[619]&m[620]&~m[622]&m[623])|(~m[618]&m[619]&m[620]&~m[622]&m[623])|(m[618]&m[619]&m[620]&~m[622]&m[623])|(m[618]&m[619]&m[620]&m[622]&m[623]));
    m[626] = (((m[623]&~m[624]&~m[625]&~m[627]&~m[628])|(~m[623]&m[624]&~m[625]&~m[627]&~m[628])|(~m[623]&~m[624]&m[625]&~m[627]&~m[628])|(m[623]&m[624]&m[625]&m[627]&~m[628])|(~m[623]&~m[624]&~m[625]&~m[627]&m[628])|(m[623]&m[624]&~m[625]&m[627]&m[628])|(m[623]&~m[624]&m[625]&m[627]&m[628])|(~m[623]&m[624]&m[625]&m[627]&m[628]))&UnbiasedRNG[398])|((m[623]&m[624]&~m[625]&~m[627]&~m[628])|(m[623]&~m[624]&m[625]&~m[627]&~m[628])|(~m[623]&m[624]&m[625]&~m[627]&~m[628])|(m[623]&m[624]&m[625]&~m[627]&~m[628])|(m[623]&~m[624]&~m[625]&~m[627]&m[628])|(~m[623]&m[624]&~m[625]&~m[627]&m[628])|(m[623]&m[624]&~m[625]&~m[627]&m[628])|(~m[623]&~m[624]&m[625]&~m[627]&m[628])|(m[623]&~m[624]&m[625]&~m[627]&m[628])|(~m[623]&m[624]&m[625]&~m[627]&m[628])|(m[623]&m[624]&m[625]&~m[627]&m[628])|(m[623]&m[624]&m[625]&m[627]&m[628]));
    m[636] = (((m[633]&~m[634]&~m[635]&~m[637]&~m[638])|(~m[633]&m[634]&~m[635]&~m[637]&~m[638])|(~m[633]&~m[634]&m[635]&~m[637]&~m[638])|(m[633]&m[634]&m[635]&m[637]&~m[638])|(~m[633]&~m[634]&~m[635]&~m[637]&m[638])|(m[633]&m[634]&~m[635]&m[637]&m[638])|(m[633]&~m[634]&m[635]&m[637]&m[638])|(~m[633]&m[634]&m[635]&m[637]&m[638]))&UnbiasedRNG[399])|((m[633]&m[634]&~m[635]&~m[637]&~m[638])|(m[633]&~m[634]&m[635]&~m[637]&~m[638])|(~m[633]&m[634]&m[635]&~m[637]&~m[638])|(m[633]&m[634]&m[635]&~m[637]&~m[638])|(m[633]&~m[634]&~m[635]&~m[637]&m[638])|(~m[633]&m[634]&~m[635]&~m[637]&m[638])|(m[633]&m[634]&~m[635]&~m[637]&m[638])|(~m[633]&~m[634]&m[635]&~m[637]&m[638])|(m[633]&~m[634]&m[635]&~m[637]&m[638])|(~m[633]&m[634]&m[635]&~m[637]&m[638])|(m[633]&m[634]&m[635]&~m[637]&m[638])|(m[633]&m[634]&m[635]&m[637]&m[638]));
    m[641] = (((m[638]&~m[639]&~m[640]&~m[642]&~m[643])|(~m[638]&m[639]&~m[640]&~m[642]&~m[643])|(~m[638]&~m[639]&m[640]&~m[642]&~m[643])|(m[638]&m[639]&m[640]&m[642]&~m[643])|(~m[638]&~m[639]&~m[640]&~m[642]&m[643])|(m[638]&m[639]&~m[640]&m[642]&m[643])|(m[638]&~m[639]&m[640]&m[642]&m[643])|(~m[638]&m[639]&m[640]&m[642]&m[643]))&UnbiasedRNG[400])|((m[638]&m[639]&~m[640]&~m[642]&~m[643])|(m[638]&~m[639]&m[640]&~m[642]&~m[643])|(~m[638]&m[639]&m[640]&~m[642]&~m[643])|(m[638]&m[639]&m[640]&~m[642]&~m[643])|(m[638]&~m[639]&~m[640]&~m[642]&m[643])|(~m[638]&m[639]&~m[640]&~m[642]&m[643])|(m[638]&m[639]&~m[640]&~m[642]&m[643])|(~m[638]&~m[639]&m[640]&~m[642]&m[643])|(m[638]&~m[639]&m[640]&~m[642]&m[643])|(~m[638]&m[639]&m[640]&~m[642]&m[643])|(m[638]&m[639]&m[640]&~m[642]&m[643])|(m[638]&m[639]&m[640]&m[642]&m[643]));
    m[646] = (((m[643]&~m[644]&~m[645]&~m[647]&~m[648])|(~m[643]&m[644]&~m[645]&~m[647]&~m[648])|(~m[643]&~m[644]&m[645]&~m[647]&~m[648])|(m[643]&m[644]&m[645]&m[647]&~m[648])|(~m[643]&~m[644]&~m[645]&~m[647]&m[648])|(m[643]&m[644]&~m[645]&m[647]&m[648])|(m[643]&~m[644]&m[645]&m[647]&m[648])|(~m[643]&m[644]&m[645]&m[647]&m[648]))&UnbiasedRNG[401])|((m[643]&m[644]&~m[645]&~m[647]&~m[648])|(m[643]&~m[644]&m[645]&~m[647]&~m[648])|(~m[643]&m[644]&m[645]&~m[647]&~m[648])|(m[643]&m[644]&m[645]&~m[647]&~m[648])|(m[643]&~m[644]&~m[645]&~m[647]&m[648])|(~m[643]&m[644]&~m[645]&~m[647]&m[648])|(m[643]&m[644]&~m[645]&~m[647]&m[648])|(~m[643]&~m[644]&m[645]&~m[647]&m[648])|(m[643]&~m[644]&m[645]&~m[647]&m[648])|(~m[643]&m[644]&m[645]&~m[647]&m[648])|(m[643]&m[644]&m[645]&~m[647]&m[648])|(m[643]&m[644]&m[645]&m[647]&m[648]));
    m[651] = (((m[648]&~m[649]&~m[650]&~m[652]&~m[653])|(~m[648]&m[649]&~m[650]&~m[652]&~m[653])|(~m[648]&~m[649]&m[650]&~m[652]&~m[653])|(m[648]&m[649]&m[650]&m[652]&~m[653])|(~m[648]&~m[649]&~m[650]&~m[652]&m[653])|(m[648]&m[649]&~m[650]&m[652]&m[653])|(m[648]&~m[649]&m[650]&m[652]&m[653])|(~m[648]&m[649]&m[650]&m[652]&m[653]))&UnbiasedRNG[402])|((m[648]&m[649]&~m[650]&~m[652]&~m[653])|(m[648]&~m[649]&m[650]&~m[652]&~m[653])|(~m[648]&m[649]&m[650]&~m[652]&~m[653])|(m[648]&m[649]&m[650]&~m[652]&~m[653])|(m[648]&~m[649]&~m[650]&~m[652]&m[653])|(~m[648]&m[649]&~m[650]&~m[652]&m[653])|(m[648]&m[649]&~m[650]&~m[652]&m[653])|(~m[648]&~m[649]&m[650]&~m[652]&m[653])|(m[648]&~m[649]&m[650]&~m[652]&m[653])|(~m[648]&m[649]&m[650]&~m[652]&m[653])|(m[648]&m[649]&m[650]&~m[652]&m[653])|(m[648]&m[649]&m[650]&m[652]&m[653]));
    m[656] = (((m[653]&~m[654]&~m[655]&~m[657]&~m[658])|(~m[653]&m[654]&~m[655]&~m[657]&~m[658])|(~m[653]&~m[654]&m[655]&~m[657]&~m[658])|(m[653]&m[654]&m[655]&m[657]&~m[658])|(~m[653]&~m[654]&~m[655]&~m[657]&m[658])|(m[653]&m[654]&~m[655]&m[657]&m[658])|(m[653]&~m[654]&m[655]&m[657]&m[658])|(~m[653]&m[654]&m[655]&m[657]&m[658]))&UnbiasedRNG[403])|((m[653]&m[654]&~m[655]&~m[657]&~m[658])|(m[653]&~m[654]&m[655]&~m[657]&~m[658])|(~m[653]&m[654]&m[655]&~m[657]&~m[658])|(m[653]&m[654]&m[655]&~m[657]&~m[658])|(m[653]&~m[654]&~m[655]&~m[657]&m[658])|(~m[653]&m[654]&~m[655]&~m[657]&m[658])|(m[653]&m[654]&~m[655]&~m[657]&m[658])|(~m[653]&~m[654]&m[655]&~m[657]&m[658])|(m[653]&~m[654]&m[655]&~m[657]&m[658])|(~m[653]&m[654]&m[655]&~m[657]&m[658])|(m[653]&m[654]&m[655]&~m[657]&m[658])|(m[653]&m[654]&m[655]&m[657]&m[658]));
    m[661] = (((m[658]&~m[659]&~m[660]&~m[662]&~m[663])|(~m[658]&m[659]&~m[660]&~m[662]&~m[663])|(~m[658]&~m[659]&m[660]&~m[662]&~m[663])|(m[658]&m[659]&m[660]&m[662]&~m[663])|(~m[658]&~m[659]&~m[660]&~m[662]&m[663])|(m[658]&m[659]&~m[660]&m[662]&m[663])|(m[658]&~m[659]&m[660]&m[662]&m[663])|(~m[658]&m[659]&m[660]&m[662]&m[663]))&UnbiasedRNG[404])|((m[658]&m[659]&~m[660]&~m[662]&~m[663])|(m[658]&~m[659]&m[660]&~m[662]&~m[663])|(~m[658]&m[659]&m[660]&~m[662]&~m[663])|(m[658]&m[659]&m[660]&~m[662]&~m[663])|(m[658]&~m[659]&~m[660]&~m[662]&m[663])|(~m[658]&m[659]&~m[660]&~m[662]&m[663])|(m[658]&m[659]&~m[660]&~m[662]&m[663])|(~m[658]&~m[659]&m[660]&~m[662]&m[663])|(m[658]&~m[659]&m[660]&~m[662]&m[663])|(~m[658]&m[659]&m[660]&~m[662]&m[663])|(m[658]&m[659]&m[660]&~m[662]&m[663])|(m[658]&m[659]&m[660]&m[662]&m[663]));
    m[671] = (((m[668]&~m[669]&~m[670]&~m[672]&~m[673])|(~m[668]&m[669]&~m[670]&~m[672]&~m[673])|(~m[668]&~m[669]&m[670]&~m[672]&~m[673])|(m[668]&m[669]&m[670]&m[672]&~m[673])|(~m[668]&~m[669]&~m[670]&~m[672]&m[673])|(m[668]&m[669]&~m[670]&m[672]&m[673])|(m[668]&~m[669]&m[670]&m[672]&m[673])|(~m[668]&m[669]&m[670]&m[672]&m[673]))&UnbiasedRNG[405])|((m[668]&m[669]&~m[670]&~m[672]&~m[673])|(m[668]&~m[669]&m[670]&~m[672]&~m[673])|(~m[668]&m[669]&m[670]&~m[672]&~m[673])|(m[668]&m[669]&m[670]&~m[672]&~m[673])|(m[668]&~m[669]&~m[670]&~m[672]&m[673])|(~m[668]&m[669]&~m[670]&~m[672]&m[673])|(m[668]&m[669]&~m[670]&~m[672]&m[673])|(~m[668]&~m[669]&m[670]&~m[672]&m[673])|(m[668]&~m[669]&m[670]&~m[672]&m[673])|(~m[668]&m[669]&m[670]&~m[672]&m[673])|(m[668]&m[669]&m[670]&~m[672]&m[673])|(m[668]&m[669]&m[670]&m[672]&m[673]));
    m[676] = (((m[673]&~m[674]&~m[675]&~m[677]&~m[678])|(~m[673]&m[674]&~m[675]&~m[677]&~m[678])|(~m[673]&~m[674]&m[675]&~m[677]&~m[678])|(m[673]&m[674]&m[675]&m[677]&~m[678])|(~m[673]&~m[674]&~m[675]&~m[677]&m[678])|(m[673]&m[674]&~m[675]&m[677]&m[678])|(m[673]&~m[674]&m[675]&m[677]&m[678])|(~m[673]&m[674]&m[675]&m[677]&m[678]))&UnbiasedRNG[406])|((m[673]&m[674]&~m[675]&~m[677]&~m[678])|(m[673]&~m[674]&m[675]&~m[677]&~m[678])|(~m[673]&m[674]&m[675]&~m[677]&~m[678])|(m[673]&m[674]&m[675]&~m[677]&~m[678])|(m[673]&~m[674]&~m[675]&~m[677]&m[678])|(~m[673]&m[674]&~m[675]&~m[677]&m[678])|(m[673]&m[674]&~m[675]&~m[677]&m[678])|(~m[673]&~m[674]&m[675]&~m[677]&m[678])|(m[673]&~m[674]&m[675]&~m[677]&m[678])|(~m[673]&m[674]&m[675]&~m[677]&m[678])|(m[673]&m[674]&m[675]&~m[677]&m[678])|(m[673]&m[674]&m[675]&m[677]&m[678]));
    m[681] = (((m[678]&~m[679]&~m[680]&~m[682]&~m[683])|(~m[678]&m[679]&~m[680]&~m[682]&~m[683])|(~m[678]&~m[679]&m[680]&~m[682]&~m[683])|(m[678]&m[679]&m[680]&m[682]&~m[683])|(~m[678]&~m[679]&~m[680]&~m[682]&m[683])|(m[678]&m[679]&~m[680]&m[682]&m[683])|(m[678]&~m[679]&m[680]&m[682]&m[683])|(~m[678]&m[679]&m[680]&m[682]&m[683]))&UnbiasedRNG[407])|((m[678]&m[679]&~m[680]&~m[682]&~m[683])|(m[678]&~m[679]&m[680]&~m[682]&~m[683])|(~m[678]&m[679]&m[680]&~m[682]&~m[683])|(m[678]&m[679]&m[680]&~m[682]&~m[683])|(m[678]&~m[679]&~m[680]&~m[682]&m[683])|(~m[678]&m[679]&~m[680]&~m[682]&m[683])|(m[678]&m[679]&~m[680]&~m[682]&m[683])|(~m[678]&~m[679]&m[680]&~m[682]&m[683])|(m[678]&~m[679]&m[680]&~m[682]&m[683])|(~m[678]&m[679]&m[680]&~m[682]&m[683])|(m[678]&m[679]&m[680]&~m[682]&m[683])|(m[678]&m[679]&m[680]&m[682]&m[683]));
    m[686] = (((m[683]&~m[684]&~m[685]&~m[687]&~m[688])|(~m[683]&m[684]&~m[685]&~m[687]&~m[688])|(~m[683]&~m[684]&m[685]&~m[687]&~m[688])|(m[683]&m[684]&m[685]&m[687]&~m[688])|(~m[683]&~m[684]&~m[685]&~m[687]&m[688])|(m[683]&m[684]&~m[685]&m[687]&m[688])|(m[683]&~m[684]&m[685]&m[687]&m[688])|(~m[683]&m[684]&m[685]&m[687]&m[688]))&UnbiasedRNG[408])|((m[683]&m[684]&~m[685]&~m[687]&~m[688])|(m[683]&~m[684]&m[685]&~m[687]&~m[688])|(~m[683]&m[684]&m[685]&~m[687]&~m[688])|(m[683]&m[684]&m[685]&~m[687]&~m[688])|(m[683]&~m[684]&~m[685]&~m[687]&m[688])|(~m[683]&m[684]&~m[685]&~m[687]&m[688])|(m[683]&m[684]&~m[685]&~m[687]&m[688])|(~m[683]&~m[684]&m[685]&~m[687]&m[688])|(m[683]&~m[684]&m[685]&~m[687]&m[688])|(~m[683]&m[684]&m[685]&~m[687]&m[688])|(m[683]&m[684]&m[685]&~m[687]&m[688])|(m[683]&m[684]&m[685]&m[687]&m[688]));
    m[691] = (((m[688]&~m[689]&~m[690]&~m[692]&~m[693])|(~m[688]&m[689]&~m[690]&~m[692]&~m[693])|(~m[688]&~m[689]&m[690]&~m[692]&~m[693])|(m[688]&m[689]&m[690]&m[692]&~m[693])|(~m[688]&~m[689]&~m[690]&~m[692]&m[693])|(m[688]&m[689]&~m[690]&m[692]&m[693])|(m[688]&~m[689]&m[690]&m[692]&m[693])|(~m[688]&m[689]&m[690]&m[692]&m[693]))&UnbiasedRNG[409])|((m[688]&m[689]&~m[690]&~m[692]&~m[693])|(m[688]&~m[689]&m[690]&~m[692]&~m[693])|(~m[688]&m[689]&m[690]&~m[692]&~m[693])|(m[688]&m[689]&m[690]&~m[692]&~m[693])|(m[688]&~m[689]&~m[690]&~m[692]&m[693])|(~m[688]&m[689]&~m[690]&~m[692]&m[693])|(m[688]&m[689]&~m[690]&~m[692]&m[693])|(~m[688]&~m[689]&m[690]&~m[692]&m[693])|(m[688]&~m[689]&m[690]&~m[692]&m[693])|(~m[688]&m[689]&m[690]&~m[692]&m[693])|(m[688]&m[689]&m[690]&~m[692]&m[693])|(m[688]&m[689]&m[690]&m[692]&m[693]));
    m[696] = (((m[693]&~m[694]&~m[695]&~m[697]&~m[698])|(~m[693]&m[694]&~m[695]&~m[697]&~m[698])|(~m[693]&~m[694]&m[695]&~m[697]&~m[698])|(m[693]&m[694]&m[695]&m[697]&~m[698])|(~m[693]&~m[694]&~m[695]&~m[697]&m[698])|(m[693]&m[694]&~m[695]&m[697]&m[698])|(m[693]&~m[694]&m[695]&m[697]&m[698])|(~m[693]&m[694]&m[695]&m[697]&m[698]))&UnbiasedRNG[410])|((m[693]&m[694]&~m[695]&~m[697]&~m[698])|(m[693]&~m[694]&m[695]&~m[697]&~m[698])|(~m[693]&m[694]&m[695]&~m[697]&~m[698])|(m[693]&m[694]&m[695]&~m[697]&~m[698])|(m[693]&~m[694]&~m[695]&~m[697]&m[698])|(~m[693]&m[694]&~m[695]&~m[697]&m[698])|(m[693]&m[694]&~m[695]&~m[697]&m[698])|(~m[693]&~m[694]&m[695]&~m[697]&m[698])|(m[693]&~m[694]&m[695]&~m[697]&m[698])|(~m[693]&m[694]&m[695]&~m[697]&m[698])|(m[693]&m[694]&m[695]&~m[697]&m[698])|(m[693]&m[694]&m[695]&m[697]&m[698]));
    m[701] = (((m[698]&~m[699]&~m[700]&~m[702]&~m[703])|(~m[698]&m[699]&~m[700]&~m[702]&~m[703])|(~m[698]&~m[699]&m[700]&~m[702]&~m[703])|(m[698]&m[699]&m[700]&m[702]&~m[703])|(~m[698]&~m[699]&~m[700]&~m[702]&m[703])|(m[698]&m[699]&~m[700]&m[702]&m[703])|(m[698]&~m[699]&m[700]&m[702]&m[703])|(~m[698]&m[699]&m[700]&m[702]&m[703]))&UnbiasedRNG[411])|((m[698]&m[699]&~m[700]&~m[702]&~m[703])|(m[698]&~m[699]&m[700]&~m[702]&~m[703])|(~m[698]&m[699]&m[700]&~m[702]&~m[703])|(m[698]&m[699]&m[700]&~m[702]&~m[703])|(m[698]&~m[699]&~m[700]&~m[702]&m[703])|(~m[698]&m[699]&~m[700]&~m[702]&m[703])|(m[698]&m[699]&~m[700]&~m[702]&m[703])|(~m[698]&~m[699]&m[700]&~m[702]&m[703])|(m[698]&~m[699]&m[700]&~m[702]&m[703])|(~m[698]&m[699]&m[700]&~m[702]&m[703])|(m[698]&m[699]&m[700]&~m[702]&m[703])|(m[698]&m[699]&m[700]&m[702]&m[703]));
    m[711] = (((m[708]&~m[709]&~m[710]&~m[712]&~m[713])|(~m[708]&m[709]&~m[710]&~m[712]&~m[713])|(~m[708]&~m[709]&m[710]&~m[712]&~m[713])|(m[708]&m[709]&m[710]&m[712]&~m[713])|(~m[708]&~m[709]&~m[710]&~m[712]&m[713])|(m[708]&m[709]&~m[710]&m[712]&m[713])|(m[708]&~m[709]&m[710]&m[712]&m[713])|(~m[708]&m[709]&m[710]&m[712]&m[713]))&UnbiasedRNG[412])|((m[708]&m[709]&~m[710]&~m[712]&~m[713])|(m[708]&~m[709]&m[710]&~m[712]&~m[713])|(~m[708]&m[709]&m[710]&~m[712]&~m[713])|(m[708]&m[709]&m[710]&~m[712]&~m[713])|(m[708]&~m[709]&~m[710]&~m[712]&m[713])|(~m[708]&m[709]&~m[710]&~m[712]&m[713])|(m[708]&m[709]&~m[710]&~m[712]&m[713])|(~m[708]&~m[709]&m[710]&~m[712]&m[713])|(m[708]&~m[709]&m[710]&~m[712]&m[713])|(~m[708]&m[709]&m[710]&~m[712]&m[713])|(m[708]&m[709]&m[710]&~m[712]&m[713])|(m[708]&m[709]&m[710]&m[712]&m[713]));
    m[716] = (((m[713]&~m[714]&~m[715]&~m[717]&~m[718])|(~m[713]&m[714]&~m[715]&~m[717]&~m[718])|(~m[713]&~m[714]&m[715]&~m[717]&~m[718])|(m[713]&m[714]&m[715]&m[717]&~m[718])|(~m[713]&~m[714]&~m[715]&~m[717]&m[718])|(m[713]&m[714]&~m[715]&m[717]&m[718])|(m[713]&~m[714]&m[715]&m[717]&m[718])|(~m[713]&m[714]&m[715]&m[717]&m[718]))&UnbiasedRNG[413])|((m[713]&m[714]&~m[715]&~m[717]&~m[718])|(m[713]&~m[714]&m[715]&~m[717]&~m[718])|(~m[713]&m[714]&m[715]&~m[717]&~m[718])|(m[713]&m[714]&m[715]&~m[717]&~m[718])|(m[713]&~m[714]&~m[715]&~m[717]&m[718])|(~m[713]&m[714]&~m[715]&~m[717]&m[718])|(m[713]&m[714]&~m[715]&~m[717]&m[718])|(~m[713]&~m[714]&m[715]&~m[717]&m[718])|(m[713]&~m[714]&m[715]&~m[717]&m[718])|(~m[713]&m[714]&m[715]&~m[717]&m[718])|(m[713]&m[714]&m[715]&~m[717]&m[718])|(m[713]&m[714]&m[715]&m[717]&m[718]));
    m[721] = (((m[718]&~m[719]&~m[720]&~m[722]&~m[723])|(~m[718]&m[719]&~m[720]&~m[722]&~m[723])|(~m[718]&~m[719]&m[720]&~m[722]&~m[723])|(m[718]&m[719]&m[720]&m[722]&~m[723])|(~m[718]&~m[719]&~m[720]&~m[722]&m[723])|(m[718]&m[719]&~m[720]&m[722]&m[723])|(m[718]&~m[719]&m[720]&m[722]&m[723])|(~m[718]&m[719]&m[720]&m[722]&m[723]))&UnbiasedRNG[414])|((m[718]&m[719]&~m[720]&~m[722]&~m[723])|(m[718]&~m[719]&m[720]&~m[722]&~m[723])|(~m[718]&m[719]&m[720]&~m[722]&~m[723])|(m[718]&m[719]&m[720]&~m[722]&~m[723])|(m[718]&~m[719]&~m[720]&~m[722]&m[723])|(~m[718]&m[719]&~m[720]&~m[722]&m[723])|(m[718]&m[719]&~m[720]&~m[722]&m[723])|(~m[718]&~m[719]&m[720]&~m[722]&m[723])|(m[718]&~m[719]&m[720]&~m[722]&m[723])|(~m[718]&m[719]&m[720]&~m[722]&m[723])|(m[718]&m[719]&m[720]&~m[722]&m[723])|(m[718]&m[719]&m[720]&m[722]&m[723]));
    m[726] = (((m[723]&~m[724]&~m[725]&~m[727]&~m[728])|(~m[723]&m[724]&~m[725]&~m[727]&~m[728])|(~m[723]&~m[724]&m[725]&~m[727]&~m[728])|(m[723]&m[724]&m[725]&m[727]&~m[728])|(~m[723]&~m[724]&~m[725]&~m[727]&m[728])|(m[723]&m[724]&~m[725]&m[727]&m[728])|(m[723]&~m[724]&m[725]&m[727]&m[728])|(~m[723]&m[724]&m[725]&m[727]&m[728]))&UnbiasedRNG[415])|((m[723]&m[724]&~m[725]&~m[727]&~m[728])|(m[723]&~m[724]&m[725]&~m[727]&~m[728])|(~m[723]&m[724]&m[725]&~m[727]&~m[728])|(m[723]&m[724]&m[725]&~m[727]&~m[728])|(m[723]&~m[724]&~m[725]&~m[727]&m[728])|(~m[723]&m[724]&~m[725]&~m[727]&m[728])|(m[723]&m[724]&~m[725]&~m[727]&m[728])|(~m[723]&~m[724]&m[725]&~m[727]&m[728])|(m[723]&~m[724]&m[725]&~m[727]&m[728])|(~m[723]&m[724]&m[725]&~m[727]&m[728])|(m[723]&m[724]&m[725]&~m[727]&m[728])|(m[723]&m[724]&m[725]&m[727]&m[728]));
    m[731] = (((m[728]&~m[729]&~m[730]&~m[732]&~m[733])|(~m[728]&m[729]&~m[730]&~m[732]&~m[733])|(~m[728]&~m[729]&m[730]&~m[732]&~m[733])|(m[728]&m[729]&m[730]&m[732]&~m[733])|(~m[728]&~m[729]&~m[730]&~m[732]&m[733])|(m[728]&m[729]&~m[730]&m[732]&m[733])|(m[728]&~m[729]&m[730]&m[732]&m[733])|(~m[728]&m[729]&m[730]&m[732]&m[733]))&UnbiasedRNG[416])|((m[728]&m[729]&~m[730]&~m[732]&~m[733])|(m[728]&~m[729]&m[730]&~m[732]&~m[733])|(~m[728]&m[729]&m[730]&~m[732]&~m[733])|(m[728]&m[729]&m[730]&~m[732]&~m[733])|(m[728]&~m[729]&~m[730]&~m[732]&m[733])|(~m[728]&m[729]&~m[730]&~m[732]&m[733])|(m[728]&m[729]&~m[730]&~m[732]&m[733])|(~m[728]&~m[729]&m[730]&~m[732]&m[733])|(m[728]&~m[729]&m[730]&~m[732]&m[733])|(~m[728]&m[729]&m[730]&~m[732]&m[733])|(m[728]&m[729]&m[730]&~m[732]&m[733])|(m[728]&m[729]&m[730]&m[732]&m[733]));
    m[736] = (((m[733]&~m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&~m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&m[737]&~m[738])|(~m[733]&~m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&m[737]&m[738])|(m[733]&~m[734]&m[735]&m[737]&m[738])|(~m[733]&m[734]&m[735]&m[737]&m[738]))&UnbiasedRNG[417])|((m[733]&m[734]&~m[735]&~m[737]&~m[738])|(m[733]&~m[734]&m[735]&~m[737]&~m[738])|(~m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&~m[734]&~m[735]&~m[737]&m[738])|(~m[733]&m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&~m[737]&m[738])|(~m[733]&~m[734]&m[735]&~m[737]&m[738])|(m[733]&~m[734]&m[735]&~m[737]&m[738])|(~m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&m[737]&m[738]));
    m[741] = (((m[738]&~m[739]&~m[740]&~m[742]&~m[743])|(~m[738]&m[739]&~m[740]&~m[742]&~m[743])|(~m[738]&~m[739]&m[740]&~m[742]&~m[743])|(m[738]&m[739]&m[740]&m[742]&~m[743])|(~m[738]&~m[739]&~m[740]&~m[742]&m[743])|(m[738]&m[739]&~m[740]&m[742]&m[743])|(m[738]&~m[739]&m[740]&m[742]&m[743])|(~m[738]&m[739]&m[740]&m[742]&m[743]))&UnbiasedRNG[418])|((m[738]&m[739]&~m[740]&~m[742]&~m[743])|(m[738]&~m[739]&m[740]&~m[742]&~m[743])|(~m[738]&m[739]&m[740]&~m[742]&~m[743])|(m[738]&m[739]&m[740]&~m[742]&~m[743])|(m[738]&~m[739]&~m[740]&~m[742]&m[743])|(~m[738]&m[739]&~m[740]&~m[742]&m[743])|(m[738]&m[739]&~m[740]&~m[742]&m[743])|(~m[738]&~m[739]&m[740]&~m[742]&m[743])|(m[738]&~m[739]&m[740]&~m[742]&m[743])|(~m[738]&m[739]&m[740]&~m[742]&m[743])|(m[738]&m[739]&m[740]&~m[742]&m[743])|(m[738]&m[739]&m[740]&m[742]&m[743]));
    m[746] = (((m[743]&~m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&~m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&m[747]&~m[748])|(~m[743]&~m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&m[747]&m[748])|(m[743]&~m[744]&m[745]&m[747]&m[748])|(~m[743]&m[744]&m[745]&m[747]&m[748]))&UnbiasedRNG[419])|((m[743]&m[744]&~m[745]&~m[747]&~m[748])|(m[743]&~m[744]&m[745]&~m[747]&~m[748])|(~m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&~m[744]&~m[745]&~m[747]&m[748])|(~m[743]&m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&~m[747]&m[748])|(~m[743]&~m[744]&m[745]&~m[747]&m[748])|(m[743]&~m[744]&m[745]&~m[747]&m[748])|(~m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&m[747]&m[748]));
    m[756] = (((m[753]&~m[754]&~m[755]&~m[757]&~m[758])|(~m[753]&m[754]&~m[755]&~m[757]&~m[758])|(~m[753]&~m[754]&m[755]&~m[757]&~m[758])|(m[753]&m[754]&m[755]&m[757]&~m[758])|(~m[753]&~m[754]&~m[755]&~m[757]&m[758])|(m[753]&m[754]&~m[755]&m[757]&m[758])|(m[753]&~m[754]&m[755]&m[757]&m[758])|(~m[753]&m[754]&m[755]&m[757]&m[758]))&UnbiasedRNG[420])|((m[753]&m[754]&~m[755]&~m[757]&~m[758])|(m[753]&~m[754]&m[755]&~m[757]&~m[758])|(~m[753]&m[754]&m[755]&~m[757]&~m[758])|(m[753]&m[754]&m[755]&~m[757]&~m[758])|(m[753]&~m[754]&~m[755]&~m[757]&m[758])|(~m[753]&m[754]&~m[755]&~m[757]&m[758])|(m[753]&m[754]&~m[755]&~m[757]&m[758])|(~m[753]&~m[754]&m[755]&~m[757]&m[758])|(m[753]&~m[754]&m[755]&~m[757]&m[758])|(~m[753]&m[754]&m[755]&~m[757]&m[758])|(m[753]&m[754]&m[755]&~m[757]&m[758])|(m[753]&m[754]&m[755]&m[757]&m[758]));
    m[761] = (((m[758]&~m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&~m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&m[762]&~m[763])|(~m[758]&~m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&m[762]&m[763])|(m[758]&~m[759]&m[760]&m[762]&m[763])|(~m[758]&m[759]&m[760]&m[762]&m[763]))&UnbiasedRNG[421])|((m[758]&m[759]&~m[760]&~m[762]&~m[763])|(m[758]&~m[759]&m[760]&~m[762]&~m[763])|(~m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&~m[759]&~m[760]&~m[762]&m[763])|(~m[758]&m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&~m[762]&m[763])|(~m[758]&~m[759]&m[760]&~m[762]&m[763])|(m[758]&~m[759]&m[760]&~m[762]&m[763])|(~m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&m[762]&m[763]));
    m[766] = (((m[763]&~m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&~m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&m[767]&~m[768])|(~m[763]&~m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&m[767]&m[768])|(m[763]&~m[764]&m[765]&m[767]&m[768])|(~m[763]&m[764]&m[765]&m[767]&m[768]))&UnbiasedRNG[422])|((m[763]&m[764]&~m[765]&~m[767]&~m[768])|(m[763]&~m[764]&m[765]&~m[767]&~m[768])|(~m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&~m[764]&~m[765]&~m[767]&m[768])|(~m[763]&m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&~m[767]&m[768])|(~m[763]&~m[764]&m[765]&~m[767]&m[768])|(m[763]&~m[764]&m[765]&~m[767]&m[768])|(~m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&m[767]&m[768]));
    m[771] = (((m[768]&~m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&~m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&m[772]&~m[773])|(~m[768]&~m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&m[772]&m[773])|(m[768]&~m[769]&m[770]&m[772]&m[773])|(~m[768]&m[769]&m[770]&m[772]&m[773]))&UnbiasedRNG[423])|((m[768]&m[769]&~m[770]&~m[772]&~m[773])|(m[768]&~m[769]&m[770]&~m[772]&~m[773])|(~m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&~m[769]&~m[770]&~m[772]&m[773])|(~m[768]&m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&~m[772]&m[773])|(~m[768]&~m[769]&m[770]&~m[772]&m[773])|(m[768]&~m[769]&m[770]&~m[772]&m[773])|(~m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&m[772]&m[773]));
    m[776] = (((m[773]&~m[774]&~m[775]&~m[777]&~m[778])|(~m[773]&m[774]&~m[775]&~m[777]&~m[778])|(~m[773]&~m[774]&m[775]&~m[777]&~m[778])|(m[773]&m[774]&m[775]&m[777]&~m[778])|(~m[773]&~m[774]&~m[775]&~m[777]&m[778])|(m[773]&m[774]&~m[775]&m[777]&m[778])|(m[773]&~m[774]&m[775]&m[777]&m[778])|(~m[773]&m[774]&m[775]&m[777]&m[778]))&UnbiasedRNG[424])|((m[773]&m[774]&~m[775]&~m[777]&~m[778])|(m[773]&~m[774]&m[775]&~m[777]&~m[778])|(~m[773]&m[774]&m[775]&~m[777]&~m[778])|(m[773]&m[774]&m[775]&~m[777]&~m[778])|(m[773]&~m[774]&~m[775]&~m[777]&m[778])|(~m[773]&m[774]&~m[775]&~m[777]&m[778])|(m[773]&m[774]&~m[775]&~m[777]&m[778])|(~m[773]&~m[774]&m[775]&~m[777]&m[778])|(m[773]&~m[774]&m[775]&~m[777]&m[778])|(~m[773]&m[774]&m[775]&~m[777]&m[778])|(m[773]&m[774]&m[775]&~m[777]&m[778])|(m[773]&m[774]&m[775]&m[777]&m[778]));
    m[781] = (((m[778]&~m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&~m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&m[782]&~m[783])|(~m[778]&~m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&m[782]&m[783])|(m[778]&~m[779]&m[780]&m[782]&m[783])|(~m[778]&m[779]&m[780]&m[782]&m[783]))&UnbiasedRNG[425])|((m[778]&m[779]&~m[780]&~m[782]&~m[783])|(m[778]&~m[779]&m[780]&~m[782]&~m[783])|(~m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&~m[779]&~m[780]&~m[782]&m[783])|(~m[778]&m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&~m[782]&m[783])|(~m[778]&~m[779]&m[780]&~m[782]&m[783])|(m[778]&~m[779]&m[780]&~m[782]&m[783])|(~m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&m[782]&m[783]));
    m[786] = (((m[783]&~m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&~m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&m[787]&~m[788])|(~m[783]&~m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&m[787]&m[788])|(m[783]&~m[784]&m[785]&m[787]&m[788])|(~m[783]&m[784]&m[785]&m[787]&m[788]))&UnbiasedRNG[426])|((m[783]&m[784]&~m[785]&~m[787]&~m[788])|(m[783]&~m[784]&m[785]&~m[787]&~m[788])|(~m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&~m[784]&~m[785]&~m[787]&m[788])|(~m[783]&m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&~m[787]&m[788])|(~m[783]&~m[784]&m[785]&~m[787]&m[788])|(m[783]&~m[784]&m[785]&~m[787]&m[788])|(~m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&m[787]&m[788]));
    m[791] = (((m[788]&~m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&~m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&m[792]&~m[793])|(~m[788]&~m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&m[792]&m[793])|(m[788]&~m[789]&m[790]&m[792]&m[793])|(~m[788]&m[789]&m[790]&m[792]&m[793]))&UnbiasedRNG[427])|((m[788]&m[789]&~m[790]&~m[792]&~m[793])|(m[788]&~m[789]&m[790]&~m[792]&~m[793])|(~m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&~m[789]&~m[790]&~m[792]&m[793])|(~m[788]&m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&~m[792]&m[793])|(~m[788]&~m[789]&m[790]&~m[792]&m[793])|(m[788]&~m[789]&m[790]&~m[792]&m[793])|(~m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&m[792]&m[793]));
    m[796] = (((m[793]&~m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&~m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&m[797]&~m[798])|(~m[793]&~m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&m[797]&m[798])|(m[793]&~m[794]&m[795]&m[797]&m[798])|(~m[793]&m[794]&m[795]&m[797]&m[798]))&UnbiasedRNG[428])|((m[793]&m[794]&~m[795]&~m[797]&~m[798])|(m[793]&~m[794]&m[795]&~m[797]&~m[798])|(~m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&~m[794]&~m[795]&~m[797]&m[798])|(~m[793]&m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&~m[797]&m[798])|(~m[793]&~m[794]&m[795]&~m[797]&m[798])|(m[793]&~m[794]&m[795]&~m[797]&m[798])|(~m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&m[797]&m[798]));
    m[806] = (((m[803]&~m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&~m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&m[807]&~m[808])|(~m[803]&~m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&m[807]&m[808])|(m[803]&~m[804]&m[805]&m[807]&m[808])|(~m[803]&m[804]&m[805]&m[807]&m[808]))&UnbiasedRNG[429])|((m[803]&m[804]&~m[805]&~m[807]&~m[808])|(m[803]&~m[804]&m[805]&~m[807]&~m[808])|(~m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&~m[804]&~m[805]&~m[807]&m[808])|(~m[803]&m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&~m[807]&m[808])|(~m[803]&~m[804]&m[805]&~m[807]&m[808])|(m[803]&~m[804]&m[805]&~m[807]&m[808])|(~m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&m[807]&m[808]));
    m[811] = (((m[808]&~m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&~m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&m[812]&~m[813])|(~m[808]&~m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&m[812]&m[813])|(m[808]&~m[809]&m[810]&m[812]&m[813])|(~m[808]&m[809]&m[810]&m[812]&m[813]))&UnbiasedRNG[430])|((m[808]&m[809]&~m[810]&~m[812]&~m[813])|(m[808]&~m[809]&m[810]&~m[812]&~m[813])|(~m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&~m[809]&~m[810]&~m[812]&m[813])|(~m[808]&m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&~m[812]&m[813])|(~m[808]&~m[809]&m[810]&~m[812]&m[813])|(m[808]&~m[809]&m[810]&~m[812]&m[813])|(~m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&m[812]&m[813]));
    m[816] = (((m[813]&~m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&~m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&m[817]&~m[818])|(~m[813]&~m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&m[817]&m[818])|(m[813]&~m[814]&m[815]&m[817]&m[818])|(~m[813]&m[814]&m[815]&m[817]&m[818]))&UnbiasedRNG[431])|((m[813]&m[814]&~m[815]&~m[817]&~m[818])|(m[813]&~m[814]&m[815]&~m[817]&~m[818])|(~m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&~m[814]&~m[815]&~m[817]&m[818])|(~m[813]&m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&~m[817]&m[818])|(~m[813]&~m[814]&m[815]&~m[817]&m[818])|(m[813]&~m[814]&m[815]&~m[817]&m[818])|(~m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&m[817]&m[818]));
    m[821] = (((m[818]&~m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&~m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&m[822]&~m[823])|(~m[818]&~m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&m[822]&m[823])|(m[818]&~m[819]&m[820]&m[822]&m[823])|(~m[818]&m[819]&m[820]&m[822]&m[823]))&UnbiasedRNG[432])|((m[818]&m[819]&~m[820]&~m[822]&~m[823])|(m[818]&~m[819]&m[820]&~m[822]&~m[823])|(~m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&~m[819]&~m[820]&~m[822]&m[823])|(~m[818]&m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&~m[822]&m[823])|(~m[818]&~m[819]&m[820]&~m[822]&m[823])|(m[818]&~m[819]&m[820]&~m[822]&m[823])|(~m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&m[822]&m[823]));
    m[826] = (((m[823]&~m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&~m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&m[827]&~m[828])|(~m[823]&~m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&m[827]&m[828])|(m[823]&~m[824]&m[825]&m[827]&m[828])|(~m[823]&m[824]&m[825]&m[827]&m[828]))&UnbiasedRNG[433])|((m[823]&m[824]&~m[825]&~m[827]&~m[828])|(m[823]&~m[824]&m[825]&~m[827]&~m[828])|(~m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&~m[824]&~m[825]&~m[827]&m[828])|(~m[823]&m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&~m[827]&m[828])|(~m[823]&~m[824]&m[825]&~m[827]&m[828])|(m[823]&~m[824]&m[825]&~m[827]&m[828])|(~m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&m[827]&m[828]));
    m[831] = (((m[828]&~m[829]&~m[830]&~m[832]&~m[833])|(~m[828]&m[829]&~m[830]&~m[832]&~m[833])|(~m[828]&~m[829]&m[830]&~m[832]&~m[833])|(m[828]&m[829]&m[830]&m[832]&~m[833])|(~m[828]&~m[829]&~m[830]&~m[832]&m[833])|(m[828]&m[829]&~m[830]&m[832]&m[833])|(m[828]&~m[829]&m[830]&m[832]&m[833])|(~m[828]&m[829]&m[830]&m[832]&m[833]))&UnbiasedRNG[434])|((m[828]&m[829]&~m[830]&~m[832]&~m[833])|(m[828]&~m[829]&m[830]&~m[832]&~m[833])|(~m[828]&m[829]&m[830]&~m[832]&~m[833])|(m[828]&m[829]&m[830]&~m[832]&~m[833])|(m[828]&~m[829]&~m[830]&~m[832]&m[833])|(~m[828]&m[829]&~m[830]&~m[832]&m[833])|(m[828]&m[829]&~m[830]&~m[832]&m[833])|(~m[828]&~m[829]&m[830]&~m[832]&m[833])|(m[828]&~m[829]&m[830]&~m[832]&m[833])|(~m[828]&m[829]&m[830]&~m[832]&m[833])|(m[828]&m[829]&m[830]&~m[832]&m[833])|(m[828]&m[829]&m[830]&m[832]&m[833]));
    m[836] = (((m[833]&~m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&~m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&m[837]&~m[838])|(~m[833]&~m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&m[837]&m[838])|(m[833]&~m[834]&m[835]&m[837]&m[838])|(~m[833]&m[834]&m[835]&m[837]&m[838]))&UnbiasedRNG[435])|((m[833]&m[834]&~m[835]&~m[837]&~m[838])|(m[833]&~m[834]&m[835]&~m[837]&~m[838])|(~m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&~m[834]&~m[835]&~m[837]&m[838])|(~m[833]&m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&~m[837]&m[838])|(~m[833]&~m[834]&m[835]&~m[837]&m[838])|(m[833]&~m[834]&m[835]&~m[837]&m[838])|(~m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&m[837]&m[838]));
    m[841] = (((m[838]&~m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&~m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&m[842]&~m[843])|(~m[838]&~m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&m[842]&m[843])|(m[838]&~m[839]&m[840]&m[842]&m[843])|(~m[838]&m[839]&m[840]&m[842]&m[843]))&UnbiasedRNG[436])|((m[838]&m[839]&~m[840]&~m[842]&~m[843])|(m[838]&~m[839]&m[840]&~m[842]&~m[843])|(~m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&~m[839]&~m[840]&~m[842]&m[843])|(~m[838]&m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&~m[842]&m[843])|(~m[838]&~m[839]&m[840]&~m[842]&m[843])|(m[838]&~m[839]&m[840]&~m[842]&m[843])|(~m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&m[842]&m[843]));
    m[846] = (((m[843]&~m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&~m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&m[847]&~m[848])|(~m[843]&~m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&m[847]&m[848])|(m[843]&~m[844]&m[845]&m[847]&m[848])|(~m[843]&m[844]&m[845]&m[847]&m[848]))&UnbiasedRNG[437])|((m[843]&m[844]&~m[845]&~m[847]&~m[848])|(m[843]&~m[844]&m[845]&~m[847]&~m[848])|(~m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&~m[844]&~m[845]&~m[847]&m[848])|(~m[843]&m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&~m[847]&m[848])|(~m[843]&~m[844]&m[845]&~m[847]&m[848])|(m[843]&~m[844]&m[845]&~m[847]&m[848])|(~m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&m[847]&m[848]));
    m[851] = (((m[848]&~m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&~m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&m[852]&~m[853])|(~m[848]&~m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&m[852]&m[853])|(m[848]&~m[849]&m[850]&m[852]&m[853])|(~m[848]&m[849]&m[850]&m[852]&m[853]))&UnbiasedRNG[438])|((m[848]&m[849]&~m[850]&~m[852]&~m[853])|(m[848]&~m[849]&m[850]&~m[852]&~m[853])|(~m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&~m[849]&~m[850]&~m[852]&m[853])|(~m[848]&m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&~m[852]&m[853])|(~m[848]&~m[849]&m[850]&~m[852]&m[853])|(m[848]&~m[849]&m[850]&~m[852]&m[853])|(~m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&m[852]&m[853]));
    m[861] = (((m[858]&~m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&~m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&m[862]&~m[863])|(~m[858]&~m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&m[862]&m[863])|(m[858]&~m[859]&m[860]&m[862]&m[863])|(~m[858]&m[859]&m[860]&m[862]&m[863]))&UnbiasedRNG[439])|((m[858]&m[859]&~m[860]&~m[862]&~m[863])|(m[858]&~m[859]&m[860]&~m[862]&~m[863])|(~m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&~m[859]&~m[860]&~m[862]&m[863])|(~m[858]&m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&~m[862]&m[863])|(~m[858]&~m[859]&m[860]&~m[862]&m[863])|(m[858]&~m[859]&m[860]&~m[862]&m[863])|(~m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&m[862]&m[863]));
    m[866] = (((m[863]&~m[864]&~m[865]&~m[867]&~m[868])|(~m[863]&m[864]&~m[865]&~m[867]&~m[868])|(~m[863]&~m[864]&m[865]&~m[867]&~m[868])|(m[863]&m[864]&m[865]&m[867]&~m[868])|(~m[863]&~m[864]&~m[865]&~m[867]&m[868])|(m[863]&m[864]&~m[865]&m[867]&m[868])|(m[863]&~m[864]&m[865]&m[867]&m[868])|(~m[863]&m[864]&m[865]&m[867]&m[868]))&UnbiasedRNG[440])|((m[863]&m[864]&~m[865]&~m[867]&~m[868])|(m[863]&~m[864]&m[865]&~m[867]&~m[868])|(~m[863]&m[864]&m[865]&~m[867]&~m[868])|(m[863]&m[864]&m[865]&~m[867]&~m[868])|(m[863]&~m[864]&~m[865]&~m[867]&m[868])|(~m[863]&m[864]&~m[865]&~m[867]&m[868])|(m[863]&m[864]&~m[865]&~m[867]&m[868])|(~m[863]&~m[864]&m[865]&~m[867]&m[868])|(m[863]&~m[864]&m[865]&~m[867]&m[868])|(~m[863]&m[864]&m[865]&~m[867]&m[868])|(m[863]&m[864]&m[865]&~m[867]&m[868])|(m[863]&m[864]&m[865]&m[867]&m[868]));
    m[871] = (((m[868]&~m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&~m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&m[872]&~m[873])|(~m[868]&~m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&m[872]&m[873])|(m[868]&~m[869]&m[870]&m[872]&m[873])|(~m[868]&m[869]&m[870]&m[872]&m[873]))&UnbiasedRNG[441])|((m[868]&m[869]&~m[870]&~m[872]&~m[873])|(m[868]&~m[869]&m[870]&~m[872]&~m[873])|(~m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&~m[869]&~m[870]&~m[872]&m[873])|(~m[868]&m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&~m[872]&m[873])|(~m[868]&~m[869]&m[870]&~m[872]&m[873])|(m[868]&~m[869]&m[870]&~m[872]&m[873])|(~m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&m[872]&m[873]));
    m[876] = (((m[873]&~m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&~m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&m[877]&~m[878])|(~m[873]&~m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&m[877]&m[878])|(m[873]&~m[874]&m[875]&m[877]&m[878])|(~m[873]&m[874]&m[875]&m[877]&m[878]))&UnbiasedRNG[442])|((m[873]&m[874]&~m[875]&~m[877]&~m[878])|(m[873]&~m[874]&m[875]&~m[877]&~m[878])|(~m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&~m[874]&~m[875]&~m[877]&m[878])|(~m[873]&m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&~m[877]&m[878])|(~m[873]&~m[874]&m[875]&~m[877]&m[878])|(m[873]&~m[874]&m[875]&~m[877]&m[878])|(~m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&m[877]&m[878]));
    m[881] = (((m[878]&~m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&~m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&m[882]&~m[883])|(~m[878]&~m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&m[882]&m[883])|(m[878]&~m[879]&m[880]&m[882]&m[883])|(~m[878]&m[879]&m[880]&m[882]&m[883]))&UnbiasedRNG[443])|((m[878]&m[879]&~m[880]&~m[882]&~m[883])|(m[878]&~m[879]&m[880]&~m[882]&~m[883])|(~m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&~m[879]&~m[880]&~m[882]&m[883])|(~m[878]&m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&~m[882]&m[883])|(~m[878]&~m[879]&m[880]&~m[882]&m[883])|(m[878]&~m[879]&m[880]&~m[882]&m[883])|(~m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&m[882]&m[883]));
    m[886] = (((m[883]&~m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&~m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&m[887]&~m[888])|(~m[883]&~m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&m[887]&m[888])|(m[883]&~m[884]&m[885]&m[887]&m[888])|(~m[883]&m[884]&m[885]&m[887]&m[888]))&UnbiasedRNG[444])|((m[883]&m[884]&~m[885]&~m[887]&~m[888])|(m[883]&~m[884]&m[885]&~m[887]&~m[888])|(~m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&~m[884]&~m[885]&~m[887]&m[888])|(~m[883]&m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&~m[887]&m[888])|(~m[883]&~m[884]&m[885]&~m[887]&m[888])|(m[883]&~m[884]&m[885]&~m[887]&m[888])|(~m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&m[887]&m[888]));
    m[891] = (((m[888]&~m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&~m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&m[892]&~m[893])|(~m[888]&~m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&m[892]&m[893])|(m[888]&~m[889]&m[890]&m[892]&m[893])|(~m[888]&m[889]&m[890]&m[892]&m[893]))&UnbiasedRNG[445])|((m[888]&m[889]&~m[890]&~m[892]&~m[893])|(m[888]&~m[889]&m[890]&~m[892]&~m[893])|(~m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&~m[889]&~m[890]&~m[892]&m[893])|(~m[888]&m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&~m[892]&m[893])|(~m[888]&~m[889]&m[890]&~m[892]&m[893])|(m[888]&~m[889]&m[890]&~m[892]&m[893])|(~m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&m[892]&m[893]));
    m[896] = (((m[893]&~m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&~m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&m[897]&~m[898])|(~m[893]&~m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&m[897]&m[898])|(m[893]&~m[894]&m[895]&m[897]&m[898])|(~m[893]&m[894]&m[895]&m[897]&m[898]))&UnbiasedRNG[446])|((m[893]&m[894]&~m[895]&~m[897]&~m[898])|(m[893]&~m[894]&m[895]&~m[897]&~m[898])|(~m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&~m[894]&~m[895]&~m[897]&m[898])|(~m[893]&m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&~m[897]&m[898])|(~m[893]&~m[894]&m[895]&~m[897]&m[898])|(m[893]&~m[894]&m[895]&~m[897]&m[898])|(~m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&m[897]&m[898]));
    m[901] = (((m[898]&~m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&~m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&m[902]&~m[903])|(~m[898]&~m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&m[902]&m[903])|(m[898]&~m[899]&m[900]&m[902]&m[903])|(~m[898]&m[899]&m[900]&m[902]&m[903]))&UnbiasedRNG[447])|((m[898]&m[899]&~m[900]&~m[902]&~m[903])|(m[898]&~m[899]&m[900]&~m[902]&~m[903])|(~m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&~m[899]&~m[900]&~m[902]&m[903])|(~m[898]&m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&~m[902]&m[903])|(~m[898]&~m[899]&m[900]&~m[902]&m[903])|(m[898]&~m[899]&m[900]&~m[902]&m[903])|(~m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&m[902]&m[903]));
    m[906] = (((m[903]&~m[904]&~m[905]&~m[907]&~m[908])|(~m[903]&m[904]&~m[905]&~m[907]&~m[908])|(~m[903]&~m[904]&m[905]&~m[907]&~m[908])|(m[903]&m[904]&m[905]&m[907]&~m[908])|(~m[903]&~m[904]&~m[905]&~m[907]&m[908])|(m[903]&m[904]&~m[905]&m[907]&m[908])|(m[903]&~m[904]&m[905]&m[907]&m[908])|(~m[903]&m[904]&m[905]&m[907]&m[908]))&UnbiasedRNG[448])|((m[903]&m[904]&~m[905]&~m[907]&~m[908])|(m[903]&~m[904]&m[905]&~m[907]&~m[908])|(~m[903]&m[904]&m[905]&~m[907]&~m[908])|(m[903]&m[904]&m[905]&~m[907]&~m[908])|(m[903]&~m[904]&~m[905]&~m[907]&m[908])|(~m[903]&m[904]&~m[905]&~m[907]&m[908])|(m[903]&m[904]&~m[905]&~m[907]&m[908])|(~m[903]&~m[904]&m[905]&~m[907]&m[908])|(m[903]&~m[904]&m[905]&~m[907]&m[908])|(~m[903]&m[904]&m[905]&~m[907]&m[908])|(m[903]&m[904]&m[905]&~m[907]&m[908])|(m[903]&m[904]&m[905]&m[907]&m[908]));
    m[916] = (((m[913]&~m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&~m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&m[917]&~m[918])|(~m[913]&~m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&m[917]&m[918])|(m[913]&~m[914]&m[915]&m[917]&m[918])|(~m[913]&m[914]&m[915]&m[917]&m[918]))&UnbiasedRNG[449])|((m[913]&m[914]&~m[915]&~m[917]&~m[918])|(m[913]&~m[914]&m[915]&~m[917]&~m[918])|(~m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&~m[914]&~m[915]&~m[917]&m[918])|(~m[913]&m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&~m[917]&m[918])|(~m[913]&~m[914]&m[915]&~m[917]&m[918])|(m[913]&~m[914]&m[915]&~m[917]&m[918])|(~m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&m[917]&m[918]));
    m[921] = (((m[918]&~m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&~m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&m[922]&~m[923])|(~m[918]&~m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&m[922]&m[923])|(m[918]&~m[919]&m[920]&m[922]&m[923])|(~m[918]&m[919]&m[920]&m[922]&m[923]))&UnbiasedRNG[450])|((m[918]&m[919]&~m[920]&~m[922]&~m[923])|(m[918]&~m[919]&m[920]&~m[922]&~m[923])|(~m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&~m[919]&~m[920]&~m[922]&m[923])|(~m[918]&m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&~m[922]&m[923])|(~m[918]&~m[919]&m[920]&~m[922]&m[923])|(m[918]&~m[919]&m[920]&~m[922]&m[923])|(~m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&m[922]&m[923]));
    m[926] = (((m[923]&~m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&~m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&m[927]&~m[928])|(~m[923]&~m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&m[927]&m[928])|(m[923]&~m[924]&m[925]&m[927]&m[928])|(~m[923]&m[924]&m[925]&m[927]&m[928]))&UnbiasedRNG[451])|((m[923]&m[924]&~m[925]&~m[927]&~m[928])|(m[923]&~m[924]&m[925]&~m[927]&~m[928])|(~m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&~m[924]&~m[925]&~m[927]&m[928])|(~m[923]&m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&~m[927]&m[928])|(~m[923]&~m[924]&m[925]&~m[927]&m[928])|(m[923]&~m[924]&m[925]&~m[927]&m[928])|(~m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&m[927]&m[928]));
    m[931] = (((m[928]&~m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&~m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&m[932]&~m[933])|(~m[928]&~m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&m[932]&m[933])|(m[928]&~m[929]&m[930]&m[932]&m[933])|(~m[928]&m[929]&m[930]&m[932]&m[933]))&UnbiasedRNG[452])|((m[928]&m[929]&~m[930]&~m[932]&~m[933])|(m[928]&~m[929]&m[930]&~m[932]&~m[933])|(~m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&~m[929]&~m[930]&~m[932]&m[933])|(~m[928]&m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&~m[932]&m[933])|(~m[928]&~m[929]&m[930]&~m[932]&m[933])|(m[928]&~m[929]&m[930]&~m[932]&m[933])|(~m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&m[932]&m[933]));
    m[936] = (((m[933]&~m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&~m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&m[937]&~m[938])|(~m[933]&~m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&m[937]&m[938])|(m[933]&~m[934]&m[935]&m[937]&m[938])|(~m[933]&m[934]&m[935]&m[937]&m[938]))&UnbiasedRNG[453])|((m[933]&m[934]&~m[935]&~m[937]&~m[938])|(m[933]&~m[934]&m[935]&~m[937]&~m[938])|(~m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&~m[934]&~m[935]&~m[937]&m[938])|(~m[933]&m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&~m[937]&m[938])|(~m[933]&~m[934]&m[935]&~m[937]&m[938])|(m[933]&~m[934]&m[935]&~m[937]&m[938])|(~m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&m[937]&m[938]));
    m[941] = (((m[938]&~m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&~m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&m[942]&~m[943])|(~m[938]&~m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&m[942]&m[943])|(m[938]&~m[939]&m[940]&m[942]&m[943])|(~m[938]&m[939]&m[940]&m[942]&m[943]))&UnbiasedRNG[454])|((m[938]&m[939]&~m[940]&~m[942]&~m[943])|(m[938]&~m[939]&m[940]&~m[942]&~m[943])|(~m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&~m[939]&~m[940]&~m[942]&m[943])|(~m[938]&m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&~m[942]&m[943])|(~m[938]&~m[939]&m[940]&~m[942]&m[943])|(m[938]&~m[939]&m[940]&~m[942]&m[943])|(~m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&m[942]&m[943]));
    m[946] = (((m[943]&~m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&~m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&m[947]&~m[948])|(~m[943]&~m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&m[947]&m[948])|(m[943]&~m[944]&m[945]&m[947]&m[948])|(~m[943]&m[944]&m[945]&m[947]&m[948]))&UnbiasedRNG[455])|((m[943]&m[944]&~m[945]&~m[947]&~m[948])|(m[943]&~m[944]&m[945]&~m[947]&~m[948])|(~m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&~m[944]&~m[945]&~m[947]&m[948])|(~m[943]&m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&~m[947]&m[948])|(~m[943]&~m[944]&m[945]&~m[947]&m[948])|(m[943]&~m[944]&m[945]&~m[947]&m[948])|(~m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&m[947]&m[948]));
    m[951] = (((m[948]&~m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&m[949]&~m[950]&~m[952]&~m[953])|(~m[948]&~m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&m[952]&~m[953])|(~m[948]&~m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&m[952]&m[953])|(m[948]&~m[949]&m[950]&m[952]&m[953])|(~m[948]&m[949]&m[950]&m[952]&m[953]))&UnbiasedRNG[456])|((m[948]&m[949]&~m[950]&~m[952]&~m[953])|(m[948]&~m[949]&m[950]&~m[952]&~m[953])|(~m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&m[949]&m[950]&~m[952]&~m[953])|(m[948]&~m[949]&~m[950]&~m[952]&m[953])|(~m[948]&m[949]&~m[950]&~m[952]&m[953])|(m[948]&m[949]&~m[950]&~m[952]&m[953])|(~m[948]&~m[949]&m[950]&~m[952]&m[953])|(m[948]&~m[949]&m[950]&~m[952]&m[953])|(~m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&~m[952]&m[953])|(m[948]&m[949]&m[950]&m[952]&m[953]));
    m[956] = (((m[953]&~m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&~m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&m[957]&~m[958])|(~m[953]&~m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&m[957]&m[958])|(m[953]&~m[954]&m[955]&m[957]&m[958])|(~m[953]&m[954]&m[955]&m[957]&m[958]))&UnbiasedRNG[457])|((m[953]&m[954]&~m[955]&~m[957]&~m[958])|(m[953]&~m[954]&m[955]&~m[957]&~m[958])|(~m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&~m[954]&~m[955]&~m[957]&m[958])|(~m[953]&m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&~m[957]&m[958])|(~m[953]&~m[954]&m[955]&~m[957]&m[958])|(m[953]&~m[954]&m[955]&~m[957]&m[958])|(~m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&m[957]&m[958]));
    m[966] = (((m[963]&~m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&~m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&m[967]&~m[968])|(~m[963]&~m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&m[967]&m[968])|(m[963]&~m[964]&m[965]&m[967]&m[968])|(~m[963]&m[964]&m[965]&m[967]&m[968]))&UnbiasedRNG[458])|((m[963]&m[964]&~m[965]&~m[967]&~m[968])|(m[963]&~m[964]&m[965]&~m[967]&~m[968])|(~m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&~m[964]&~m[965]&~m[967]&m[968])|(~m[963]&m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&~m[967]&m[968])|(~m[963]&~m[964]&m[965]&~m[967]&m[968])|(m[963]&~m[964]&m[965]&~m[967]&m[968])|(~m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&m[967]&m[968]));
    m[971] = (((m[968]&~m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&~m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&m[972]&~m[973])|(~m[968]&~m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&m[972]&m[973])|(m[968]&~m[969]&m[970]&m[972]&m[973])|(~m[968]&m[969]&m[970]&m[972]&m[973]))&UnbiasedRNG[459])|((m[968]&m[969]&~m[970]&~m[972]&~m[973])|(m[968]&~m[969]&m[970]&~m[972]&~m[973])|(~m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&~m[969]&~m[970]&~m[972]&m[973])|(~m[968]&m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&~m[972]&m[973])|(~m[968]&~m[969]&m[970]&~m[972]&m[973])|(m[968]&~m[969]&m[970]&~m[972]&m[973])|(~m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&m[972]&m[973]));
    m[976] = (((m[973]&~m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&~m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&m[977]&~m[978])|(~m[973]&~m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&m[977]&m[978])|(m[973]&~m[974]&m[975]&m[977]&m[978])|(~m[973]&m[974]&m[975]&m[977]&m[978]))&UnbiasedRNG[460])|((m[973]&m[974]&~m[975]&~m[977]&~m[978])|(m[973]&~m[974]&m[975]&~m[977]&~m[978])|(~m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&~m[974]&~m[975]&~m[977]&m[978])|(~m[973]&m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&~m[977]&m[978])|(~m[973]&~m[974]&m[975]&~m[977]&m[978])|(m[973]&~m[974]&m[975]&~m[977]&m[978])|(~m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&m[977]&m[978]));
    m[981] = (((m[978]&~m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&~m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&m[982]&~m[983])|(~m[978]&~m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&m[982]&m[983])|(m[978]&~m[979]&m[980]&m[982]&m[983])|(~m[978]&m[979]&m[980]&m[982]&m[983]))&UnbiasedRNG[461])|((m[978]&m[979]&~m[980]&~m[982]&~m[983])|(m[978]&~m[979]&m[980]&~m[982]&~m[983])|(~m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&~m[979]&~m[980]&~m[982]&m[983])|(~m[978]&m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&~m[982]&m[983])|(~m[978]&~m[979]&m[980]&~m[982]&m[983])|(m[978]&~m[979]&m[980]&~m[982]&m[983])|(~m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&m[982]&m[983]));
    m[986] = (((m[983]&~m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&~m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&m[987]&~m[988])|(~m[983]&~m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&m[987]&m[988])|(m[983]&~m[984]&m[985]&m[987]&m[988])|(~m[983]&m[984]&m[985]&m[987]&m[988]))&UnbiasedRNG[462])|((m[983]&m[984]&~m[985]&~m[987]&~m[988])|(m[983]&~m[984]&m[985]&~m[987]&~m[988])|(~m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&~m[984]&~m[985]&~m[987]&m[988])|(~m[983]&m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&~m[987]&m[988])|(~m[983]&~m[984]&m[985]&~m[987]&m[988])|(m[983]&~m[984]&m[985]&~m[987]&m[988])|(~m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&m[987]&m[988]));
    m[991] = (((m[988]&~m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&~m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&m[992]&~m[993])|(~m[988]&~m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&m[992]&m[993])|(m[988]&~m[989]&m[990]&m[992]&m[993])|(~m[988]&m[989]&m[990]&m[992]&m[993]))&UnbiasedRNG[463])|((m[988]&m[989]&~m[990]&~m[992]&~m[993])|(m[988]&~m[989]&m[990]&~m[992]&~m[993])|(~m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&~m[989]&~m[990]&~m[992]&m[993])|(~m[988]&m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&~m[992]&m[993])|(~m[988]&~m[989]&m[990]&~m[992]&m[993])|(m[988]&~m[989]&m[990]&~m[992]&m[993])|(~m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&m[992]&m[993]));
    m[996] = (((m[993]&~m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&~m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&m[997]&~m[998])|(~m[993]&~m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&m[997]&m[998])|(m[993]&~m[994]&m[995]&m[997]&m[998])|(~m[993]&m[994]&m[995]&m[997]&m[998]))&UnbiasedRNG[464])|((m[993]&m[994]&~m[995]&~m[997]&~m[998])|(m[993]&~m[994]&m[995]&~m[997]&~m[998])|(~m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&~m[994]&~m[995]&~m[997]&m[998])|(~m[993]&m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&~m[997]&m[998])|(~m[993]&~m[994]&m[995]&~m[997]&m[998])|(m[993]&~m[994]&m[995]&~m[997]&m[998])|(~m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&m[997]&m[998]));
    m[1001] = (((m[998]&~m[999]&~m[1000]&~m[1002]&~m[1003])|(~m[998]&m[999]&~m[1000]&~m[1002]&~m[1003])|(~m[998]&~m[999]&m[1000]&~m[1002]&~m[1003])|(m[998]&m[999]&m[1000]&m[1002]&~m[1003])|(~m[998]&~m[999]&~m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&~m[1000]&m[1002]&m[1003])|(m[998]&~m[999]&m[1000]&m[1002]&m[1003])|(~m[998]&m[999]&m[1000]&m[1002]&m[1003]))&UnbiasedRNG[465])|((m[998]&m[999]&~m[1000]&~m[1002]&~m[1003])|(m[998]&~m[999]&m[1000]&~m[1002]&~m[1003])|(~m[998]&m[999]&m[1000]&~m[1002]&~m[1003])|(m[998]&m[999]&m[1000]&~m[1002]&~m[1003])|(m[998]&~m[999]&~m[1000]&~m[1002]&m[1003])|(~m[998]&m[999]&~m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&~m[1000]&~m[1002]&m[1003])|(~m[998]&~m[999]&m[1000]&~m[1002]&m[1003])|(m[998]&~m[999]&m[1000]&~m[1002]&m[1003])|(~m[998]&m[999]&m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&m[1000]&~m[1002]&m[1003])|(m[998]&m[999]&m[1000]&m[1002]&m[1003]));
    m[1011] = (((m[1008]&~m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&~m[1013])|(~m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))&UnbiasedRNG[466])|((m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&m[1013]));
    m[1016] = (((m[1013]&~m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&~m[1018])|(~m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))&UnbiasedRNG[467])|((m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&m[1018]));
    m[1021] = (((m[1018]&~m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&~m[1023])|(~m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))&UnbiasedRNG[468])|((m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&m[1023]));
    m[1026] = (((m[1023]&~m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&~m[1028])|(~m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))&UnbiasedRNG[469])|((m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&m[1028]));
    m[1031] = (((m[1028]&~m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&~m[1033])|(~m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&m[1032]&m[1033]))&UnbiasedRNG[470])|((m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&m[1033]));
    m[1036] = (((m[1033]&~m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&~m[1038])|(~m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))&UnbiasedRNG[471])|((m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&m[1038]));
    m[1041] = (((m[1038]&~m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&~m[1043])|(~m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))&UnbiasedRNG[472])|((m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&m[1043]));
    m[1051] = (((m[1048]&~m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&~m[1053])|(~m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))&UnbiasedRNG[473])|((m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&m[1053]));
    m[1056] = (((m[1053]&~m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&~m[1058])|(~m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&m[1057]&m[1058]))&UnbiasedRNG[474])|((m[1053]&m[1054]&~m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&~m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&~m[1058])|(m[1053]&~m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&~m[1055]&~m[1057]&m[1058])|(~m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&~m[1054]&m[1055]&~m[1057]&m[1058])|(~m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&~m[1057]&m[1058])|(m[1053]&m[1054]&m[1055]&m[1057]&m[1058]));
    m[1061] = (((m[1058]&~m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&~m[1063])|(~m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))&UnbiasedRNG[475])|((m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&m[1063]));
    m[1066] = (((m[1063]&~m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&~m[1068])|(~m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&m[1067]&m[1068]))&UnbiasedRNG[476])|((m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&m[1068]));
    m[1071] = (((m[1068]&~m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&~m[1073])|(~m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))&UnbiasedRNG[477])|((m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&m[1073]));
    m[1076] = (((m[1073]&~m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&~m[1078])|(~m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))&UnbiasedRNG[478])|((m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&m[1078]));
    m[1086] = (((m[1083]&~m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&~m[1088])|(~m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))&UnbiasedRNG[479])|((m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&m[1088]));
    m[1091] = (((m[1088]&~m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&~m[1093])|(~m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))&UnbiasedRNG[480])|((m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&m[1093]));
    m[1096] = (((m[1093]&~m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&~m[1098])|(~m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))&UnbiasedRNG[481])|((m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&m[1098]));
    m[1101] = (((m[1098]&~m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&~m[1103])|(~m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))&UnbiasedRNG[482])|((m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&m[1103]));
    m[1106] = (((m[1103]&~m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&~m[1108])|(~m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&m[1107]&m[1108]))&UnbiasedRNG[483])|((m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&m[1108]));
    m[1116] = (((m[1113]&~m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&~m[1118])|(~m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&m[1117]&m[1118]))&UnbiasedRNG[484])|((m[1113]&m[1114]&~m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&~m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&~m[1118])|(m[1113]&~m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&~m[1115]&~m[1117]&m[1118])|(~m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&~m[1114]&m[1115]&~m[1117]&m[1118])|(~m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&~m[1117]&m[1118])|(m[1113]&m[1114]&m[1115]&m[1117]&m[1118]));
    m[1121] = (((m[1118]&~m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&~m[1123])|(~m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))&UnbiasedRNG[485])|((m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&m[1123]));
    m[1126] = (((m[1123]&~m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&~m[1128])|(~m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))&UnbiasedRNG[486])|((m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&m[1128]));
    m[1131] = (((m[1128]&~m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&~m[1133])|(~m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))&UnbiasedRNG[487])|((m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&m[1133]));
    m[1141] = (((m[1138]&~m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&~m[1143])|(~m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))&UnbiasedRNG[488])|((m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&m[1143]));
    m[1146] = (((m[1143]&~m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&~m[1148])|(~m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))&UnbiasedRNG[489])|((m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&m[1148]));
    m[1151] = (((m[1148]&~m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&~m[1153])|(~m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&m[1152]&m[1153]))&UnbiasedRNG[490])|((m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&m[1153]));
    m[1161] = (((m[1158]&~m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&~m[1163])|(~m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))&UnbiasedRNG[491])|((m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&m[1163]));
    m[1166] = (((m[1163]&~m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&~m[1168])|(~m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))&UnbiasedRNG[492])|((m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&m[1168]));
    m[1176] = (((m[1173]&~m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&~m[1178])|(~m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))&UnbiasedRNG[493])|((m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&m[1178]));
end

always @(posedge color4_clk) begin
    m[532] = (((m[528]&~m[529]&~m[530]&~m[531]&~m[535])|(~m[528]&m[529]&~m[530]&~m[531]&~m[535])|(~m[528]&~m[529]&m[530]&~m[531]&~m[535])|(m[528]&m[529]&~m[530]&m[531]&~m[535])|(m[528]&~m[529]&m[530]&m[531]&~m[535])|(~m[528]&m[529]&m[530]&m[531]&~m[535]))&BiasedRNG[527])|(((m[528]&~m[529]&~m[530]&~m[531]&m[535])|(~m[528]&m[529]&~m[530]&~m[531]&m[535])|(~m[528]&~m[529]&m[530]&~m[531]&m[535])|(m[528]&m[529]&~m[530]&m[531]&m[535])|(m[528]&~m[529]&m[530]&m[531]&m[535])|(~m[528]&m[529]&m[530]&m[531]&m[535]))&~BiasedRNG[527])|((m[528]&m[529]&~m[530]&~m[531]&~m[535])|(m[528]&~m[529]&m[530]&~m[531]&~m[535])|(~m[528]&m[529]&m[530]&~m[531]&~m[535])|(m[528]&m[529]&m[530]&~m[531]&~m[535])|(m[528]&m[529]&m[530]&m[531]&~m[535])|(m[528]&m[529]&~m[530]&~m[531]&m[535])|(m[528]&~m[529]&m[530]&~m[531]&m[535])|(~m[528]&m[529]&m[530]&~m[531]&m[535])|(m[528]&m[529]&m[530]&~m[531]&m[535])|(m[528]&m[529]&m[530]&m[531]&m[535]));
    m[537] = (((m[533]&~m[534]&~m[535]&~m[536]&~m[545])|(~m[533]&m[534]&~m[535]&~m[536]&~m[545])|(~m[533]&~m[534]&m[535]&~m[536]&~m[545])|(m[533]&m[534]&~m[535]&m[536]&~m[545])|(m[533]&~m[534]&m[535]&m[536]&~m[545])|(~m[533]&m[534]&m[535]&m[536]&~m[545]))&BiasedRNG[528])|(((m[533]&~m[534]&~m[535]&~m[536]&m[545])|(~m[533]&m[534]&~m[535]&~m[536]&m[545])|(~m[533]&~m[534]&m[535]&~m[536]&m[545])|(m[533]&m[534]&~m[535]&m[536]&m[545])|(m[533]&~m[534]&m[535]&m[536]&m[545])|(~m[533]&m[534]&m[535]&m[536]&m[545]))&~BiasedRNG[528])|((m[533]&m[534]&~m[535]&~m[536]&~m[545])|(m[533]&~m[534]&m[535]&~m[536]&~m[545])|(~m[533]&m[534]&m[535]&~m[536]&~m[545])|(m[533]&m[534]&m[535]&~m[536]&~m[545])|(m[533]&m[534]&m[535]&m[536]&~m[545])|(m[533]&m[534]&~m[535]&~m[536]&m[545])|(m[533]&~m[534]&m[535]&~m[536]&m[545])|(~m[533]&m[534]&m[535]&~m[536]&m[545])|(m[533]&m[534]&m[535]&~m[536]&m[545])|(m[533]&m[534]&m[535]&m[536]&m[545]));
    m[542] = (((m[538]&~m[539]&~m[540]&~m[541]&~m[550])|(~m[538]&m[539]&~m[540]&~m[541]&~m[550])|(~m[538]&~m[539]&m[540]&~m[541]&~m[550])|(m[538]&m[539]&~m[540]&m[541]&~m[550])|(m[538]&~m[539]&m[540]&m[541]&~m[550])|(~m[538]&m[539]&m[540]&m[541]&~m[550]))&BiasedRNG[529])|(((m[538]&~m[539]&~m[540]&~m[541]&m[550])|(~m[538]&m[539]&~m[540]&~m[541]&m[550])|(~m[538]&~m[539]&m[540]&~m[541]&m[550])|(m[538]&m[539]&~m[540]&m[541]&m[550])|(m[538]&~m[539]&m[540]&m[541]&m[550])|(~m[538]&m[539]&m[540]&m[541]&m[550]))&~BiasedRNG[529])|((m[538]&m[539]&~m[540]&~m[541]&~m[550])|(m[538]&~m[539]&m[540]&~m[541]&~m[550])|(~m[538]&m[539]&m[540]&~m[541]&~m[550])|(m[538]&m[539]&m[540]&~m[541]&~m[550])|(m[538]&m[539]&m[540]&m[541]&~m[550])|(m[538]&m[539]&~m[540]&~m[541]&m[550])|(m[538]&~m[539]&m[540]&~m[541]&m[550])|(~m[538]&m[539]&m[540]&~m[541]&m[550])|(m[538]&m[539]&m[540]&~m[541]&m[550])|(m[538]&m[539]&m[540]&m[541]&m[550]));
    m[547] = (((m[543]&~m[544]&~m[545]&~m[546]&~m[560])|(~m[543]&m[544]&~m[545]&~m[546]&~m[560])|(~m[543]&~m[544]&m[545]&~m[546]&~m[560])|(m[543]&m[544]&~m[545]&m[546]&~m[560])|(m[543]&~m[544]&m[545]&m[546]&~m[560])|(~m[543]&m[544]&m[545]&m[546]&~m[560]))&BiasedRNG[530])|(((m[543]&~m[544]&~m[545]&~m[546]&m[560])|(~m[543]&m[544]&~m[545]&~m[546]&m[560])|(~m[543]&~m[544]&m[545]&~m[546]&m[560])|(m[543]&m[544]&~m[545]&m[546]&m[560])|(m[543]&~m[544]&m[545]&m[546]&m[560])|(~m[543]&m[544]&m[545]&m[546]&m[560]))&~BiasedRNG[530])|((m[543]&m[544]&~m[545]&~m[546]&~m[560])|(m[543]&~m[544]&m[545]&~m[546]&~m[560])|(~m[543]&m[544]&m[545]&~m[546]&~m[560])|(m[543]&m[544]&m[545]&~m[546]&~m[560])|(m[543]&m[544]&m[545]&m[546]&~m[560])|(m[543]&m[544]&~m[545]&~m[546]&m[560])|(m[543]&~m[544]&m[545]&~m[546]&m[560])|(~m[543]&m[544]&m[545]&~m[546]&m[560])|(m[543]&m[544]&m[545]&~m[546]&m[560])|(m[543]&m[544]&m[545]&m[546]&m[560]));
    m[552] = (((m[548]&~m[549]&~m[550]&~m[551]&~m[565])|(~m[548]&m[549]&~m[550]&~m[551]&~m[565])|(~m[548]&~m[549]&m[550]&~m[551]&~m[565])|(m[548]&m[549]&~m[550]&m[551]&~m[565])|(m[548]&~m[549]&m[550]&m[551]&~m[565])|(~m[548]&m[549]&m[550]&m[551]&~m[565]))&BiasedRNG[531])|(((m[548]&~m[549]&~m[550]&~m[551]&m[565])|(~m[548]&m[549]&~m[550]&~m[551]&m[565])|(~m[548]&~m[549]&m[550]&~m[551]&m[565])|(m[548]&m[549]&~m[550]&m[551]&m[565])|(m[548]&~m[549]&m[550]&m[551]&m[565])|(~m[548]&m[549]&m[550]&m[551]&m[565]))&~BiasedRNG[531])|((m[548]&m[549]&~m[550]&~m[551]&~m[565])|(m[548]&~m[549]&m[550]&~m[551]&~m[565])|(~m[548]&m[549]&m[550]&~m[551]&~m[565])|(m[548]&m[549]&m[550]&~m[551]&~m[565])|(m[548]&m[549]&m[550]&m[551]&~m[565])|(m[548]&m[549]&~m[550]&~m[551]&m[565])|(m[548]&~m[549]&m[550]&~m[551]&m[565])|(~m[548]&m[549]&m[550]&~m[551]&m[565])|(m[548]&m[549]&m[550]&~m[551]&m[565])|(m[548]&m[549]&m[550]&m[551]&m[565]));
    m[557] = (((m[553]&~m[554]&~m[555]&~m[556]&~m[570])|(~m[553]&m[554]&~m[555]&~m[556]&~m[570])|(~m[553]&~m[554]&m[555]&~m[556]&~m[570])|(m[553]&m[554]&~m[555]&m[556]&~m[570])|(m[553]&~m[554]&m[555]&m[556]&~m[570])|(~m[553]&m[554]&m[555]&m[556]&~m[570]))&BiasedRNG[532])|(((m[553]&~m[554]&~m[555]&~m[556]&m[570])|(~m[553]&m[554]&~m[555]&~m[556]&m[570])|(~m[553]&~m[554]&m[555]&~m[556]&m[570])|(m[553]&m[554]&~m[555]&m[556]&m[570])|(m[553]&~m[554]&m[555]&m[556]&m[570])|(~m[553]&m[554]&m[555]&m[556]&m[570]))&~BiasedRNG[532])|((m[553]&m[554]&~m[555]&~m[556]&~m[570])|(m[553]&~m[554]&m[555]&~m[556]&~m[570])|(~m[553]&m[554]&m[555]&~m[556]&~m[570])|(m[553]&m[554]&m[555]&~m[556]&~m[570])|(m[553]&m[554]&m[555]&m[556]&~m[570])|(m[553]&m[554]&~m[555]&~m[556]&m[570])|(m[553]&~m[554]&m[555]&~m[556]&m[570])|(~m[553]&m[554]&m[555]&~m[556]&m[570])|(m[553]&m[554]&m[555]&~m[556]&m[570])|(m[553]&m[554]&m[555]&m[556]&m[570]));
    m[562] = (((m[558]&~m[559]&~m[560]&~m[561]&~m[580])|(~m[558]&m[559]&~m[560]&~m[561]&~m[580])|(~m[558]&~m[559]&m[560]&~m[561]&~m[580])|(m[558]&m[559]&~m[560]&m[561]&~m[580])|(m[558]&~m[559]&m[560]&m[561]&~m[580])|(~m[558]&m[559]&m[560]&m[561]&~m[580]))&BiasedRNG[533])|(((m[558]&~m[559]&~m[560]&~m[561]&m[580])|(~m[558]&m[559]&~m[560]&~m[561]&m[580])|(~m[558]&~m[559]&m[560]&~m[561]&m[580])|(m[558]&m[559]&~m[560]&m[561]&m[580])|(m[558]&~m[559]&m[560]&m[561]&m[580])|(~m[558]&m[559]&m[560]&m[561]&m[580]))&~BiasedRNG[533])|((m[558]&m[559]&~m[560]&~m[561]&~m[580])|(m[558]&~m[559]&m[560]&~m[561]&~m[580])|(~m[558]&m[559]&m[560]&~m[561]&~m[580])|(m[558]&m[559]&m[560]&~m[561]&~m[580])|(m[558]&m[559]&m[560]&m[561]&~m[580])|(m[558]&m[559]&~m[560]&~m[561]&m[580])|(m[558]&~m[559]&m[560]&~m[561]&m[580])|(~m[558]&m[559]&m[560]&~m[561]&m[580])|(m[558]&m[559]&m[560]&~m[561]&m[580])|(m[558]&m[559]&m[560]&m[561]&m[580]));
    m[567] = (((m[563]&~m[564]&~m[565]&~m[566]&~m[585])|(~m[563]&m[564]&~m[565]&~m[566]&~m[585])|(~m[563]&~m[564]&m[565]&~m[566]&~m[585])|(m[563]&m[564]&~m[565]&m[566]&~m[585])|(m[563]&~m[564]&m[565]&m[566]&~m[585])|(~m[563]&m[564]&m[565]&m[566]&~m[585]))&BiasedRNG[534])|(((m[563]&~m[564]&~m[565]&~m[566]&m[585])|(~m[563]&m[564]&~m[565]&~m[566]&m[585])|(~m[563]&~m[564]&m[565]&~m[566]&m[585])|(m[563]&m[564]&~m[565]&m[566]&m[585])|(m[563]&~m[564]&m[565]&m[566]&m[585])|(~m[563]&m[564]&m[565]&m[566]&m[585]))&~BiasedRNG[534])|((m[563]&m[564]&~m[565]&~m[566]&~m[585])|(m[563]&~m[564]&m[565]&~m[566]&~m[585])|(~m[563]&m[564]&m[565]&~m[566]&~m[585])|(m[563]&m[564]&m[565]&~m[566]&~m[585])|(m[563]&m[564]&m[565]&m[566]&~m[585])|(m[563]&m[564]&~m[565]&~m[566]&m[585])|(m[563]&~m[564]&m[565]&~m[566]&m[585])|(~m[563]&m[564]&m[565]&~m[566]&m[585])|(m[563]&m[564]&m[565]&~m[566]&m[585])|(m[563]&m[564]&m[565]&m[566]&m[585]));
    m[572] = (((m[568]&~m[569]&~m[570]&~m[571]&~m[590])|(~m[568]&m[569]&~m[570]&~m[571]&~m[590])|(~m[568]&~m[569]&m[570]&~m[571]&~m[590])|(m[568]&m[569]&~m[570]&m[571]&~m[590])|(m[568]&~m[569]&m[570]&m[571]&~m[590])|(~m[568]&m[569]&m[570]&m[571]&~m[590]))&BiasedRNG[535])|(((m[568]&~m[569]&~m[570]&~m[571]&m[590])|(~m[568]&m[569]&~m[570]&~m[571]&m[590])|(~m[568]&~m[569]&m[570]&~m[571]&m[590])|(m[568]&m[569]&~m[570]&m[571]&m[590])|(m[568]&~m[569]&m[570]&m[571]&m[590])|(~m[568]&m[569]&m[570]&m[571]&m[590]))&~BiasedRNG[535])|((m[568]&m[569]&~m[570]&~m[571]&~m[590])|(m[568]&~m[569]&m[570]&~m[571]&~m[590])|(~m[568]&m[569]&m[570]&~m[571]&~m[590])|(m[568]&m[569]&m[570]&~m[571]&~m[590])|(m[568]&m[569]&m[570]&m[571]&~m[590])|(m[568]&m[569]&~m[570]&~m[571]&m[590])|(m[568]&~m[569]&m[570]&~m[571]&m[590])|(~m[568]&m[569]&m[570]&~m[571]&m[590])|(m[568]&m[569]&m[570]&~m[571]&m[590])|(m[568]&m[569]&m[570]&m[571]&m[590]));
    m[577] = (((m[573]&~m[574]&~m[575]&~m[576]&~m[595])|(~m[573]&m[574]&~m[575]&~m[576]&~m[595])|(~m[573]&~m[574]&m[575]&~m[576]&~m[595])|(m[573]&m[574]&~m[575]&m[576]&~m[595])|(m[573]&~m[574]&m[575]&m[576]&~m[595])|(~m[573]&m[574]&m[575]&m[576]&~m[595]))&BiasedRNG[536])|(((m[573]&~m[574]&~m[575]&~m[576]&m[595])|(~m[573]&m[574]&~m[575]&~m[576]&m[595])|(~m[573]&~m[574]&m[575]&~m[576]&m[595])|(m[573]&m[574]&~m[575]&m[576]&m[595])|(m[573]&~m[574]&m[575]&m[576]&m[595])|(~m[573]&m[574]&m[575]&m[576]&m[595]))&~BiasedRNG[536])|((m[573]&m[574]&~m[575]&~m[576]&~m[595])|(m[573]&~m[574]&m[575]&~m[576]&~m[595])|(~m[573]&m[574]&m[575]&~m[576]&~m[595])|(m[573]&m[574]&m[575]&~m[576]&~m[595])|(m[573]&m[574]&m[575]&m[576]&~m[595])|(m[573]&m[574]&~m[575]&~m[576]&m[595])|(m[573]&~m[574]&m[575]&~m[576]&m[595])|(~m[573]&m[574]&m[575]&~m[576]&m[595])|(m[573]&m[574]&m[575]&~m[576]&m[595])|(m[573]&m[574]&m[575]&m[576]&m[595]));
    m[582] = (((m[578]&~m[579]&~m[580]&~m[581]&~m[605])|(~m[578]&m[579]&~m[580]&~m[581]&~m[605])|(~m[578]&~m[579]&m[580]&~m[581]&~m[605])|(m[578]&m[579]&~m[580]&m[581]&~m[605])|(m[578]&~m[579]&m[580]&m[581]&~m[605])|(~m[578]&m[579]&m[580]&m[581]&~m[605]))&BiasedRNG[537])|(((m[578]&~m[579]&~m[580]&~m[581]&m[605])|(~m[578]&m[579]&~m[580]&~m[581]&m[605])|(~m[578]&~m[579]&m[580]&~m[581]&m[605])|(m[578]&m[579]&~m[580]&m[581]&m[605])|(m[578]&~m[579]&m[580]&m[581]&m[605])|(~m[578]&m[579]&m[580]&m[581]&m[605]))&~BiasedRNG[537])|((m[578]&m[579]&~m[580]&~m[581]&~m[605])|(m[578]&~m[579]&m[580]&~m[581]&~m[605])|(~m[578]&m[579]&m[580]&~m[581]&~m[605])|(m[578]&m[579]&m[580]&~m[581]&~m[605])|(m[578]&m[579]&m[580]&m[581]&~m[605])|(m[578]&m[579]&~m[580]&~m[581]&m[605])|(m[578]&~m[579]&m[580]&~m[581]&m[605])|(~m[578]&m[579]&m[580]&~m[581]&m[605])|(m[578]&m[579]&m[580]&~m[581]&m[605])|(m[578]&m[579]&m[580]&m[581]&m[605]));
    m[587] = (((m[583]&~m[584]&~m[585]&~m[586]&~m[610])|(~m[583]&m[584]&~m[585]&~m[586]&~m[610])|(~m[583]&~m[584]&m[585]&~m[586]&~m[610])|(m[583]&m[584]&~m[585]&m[586]&~m[610])|(m[583]&~m[584]&m[585]&m[586]&~m[610])|(~m[583]&m[584]&m[585]&m[586]&~m[610]))&BiasedRNG[538])|(((m[583]&~m[584]&~m[585]&~m[586]&m[610])|(~m[583]&m[584]&~m[585]&~m[586]&m[610])|(~m[583]&~m[584]&m[585]&~m[586]&m[610])|(m[583]&m[584]&~m[585]&m[586]&m[610])|(m[583]&~m[584]&m[585]&m[586]&m[610])|(~m[583]&m[584]&m[585]&m[586]&m[610]))&~BiasedRNG[538])|((m[583]&m[584]&~m[585]&~m[586]&~m[610])|(m[583]&~m[584]&m[585]&~m[586]&~m[610])|(~m[583]&m[584]&m[585]&~m[586]&~m[610])|(m[583]&m[584]&m[585]&~m[586]&~m[610])|(m[583]&m[584]&m[585]&m[586]&~m[610])|(m[583]&m[584]&~m[585]&~m[586]&m[610])|(m[583]&~m[584]&m[585]&~m[586]&m[610])|(~m[583]&m[584]&m[585]&~m[586]&m[610])|(m[583]&m[584]&m[585]&~m[586]&m[610])|(m[583]&m[584]&m[585]&m[586]&m[610]));
    m[592] = (((m[588]&~m[589]&~m[590]&~m[591]&~m[615])|(~m[588]&m[589]&~m[590]&~m[591]&~m[615])|(~m[588]&~m[589]&m[590]&~m[591]&~m[615])|(m[588]&m[589]&~m[590]&m[591]&~m[615])|(m[588]&~m[589]&m[590]&m[591]&~m[615])|(~m[588]&m[589]&m[590]&m[591]&~m[615]))&BiasedRNG[539])|(((m[588]&~m[589]&~m[590]&~m[591]&m[615])|(~m[588]&m[589]&~m[590]&~m[591]&m[615])|(~m[588]&~m[589]&m[590]&~m[591]&m[615])|(m[588]&m[589]&~m[590]&m[591]&m[615])|(m[588]&~m[589]&m[590]&m[591]&m[615])|(~m[588]&m[589]&m[590]&m[591]&m[615]))&~BiasedRNG[539])|((m[588]&m[589]&~m[590]&~m[591]&~m[615])|(m[588]&~m[589]&m[590]&~m[591]&~m[615])|(~m[588]&m[589]&m[590]&~m[591]&~m[615])|(m[588]&m[589]&m[590]&~m[591]&~m[615])|(m[588]&m[589]&m[590]&m[591]&~m[615])|(m[588]&m[589]&~m[590]&~m[591]&m[615])|(m[588]&~m[589]&m[590]&~m[591]&m[615])|(~m[588]&m[589]&m[590]&~m[591]&m[615])|(m[588]&m[589]&m[590]&~m[591]&m[615])|(m[588]&m[589]&m[590]&m[591]&m[615]));
    m[597] = (((m[593]&~m[594]&~m[595]&~m[596]&~m[620])|(~m[593]&m[594]&~m[595]&~m[596]&~m[620])|(~m[593]&~m[594]&m[595]&~m[596]&~m[620])|(m[593]&m[594]&~m[595]&m[596]&~m[620])|(m[593]&~m[594]&m[595]&m[596]&~m[620])|(~m[593]&m[594]&m[595]&m[596]&~m[620]))&BiasedRNG[540])|(((m[593]&~m[594]&~m[595]&~m[596]&m[620])|(~m[593]&m[594]&~m[595]&~m[596]&m[620])|(~m[593]&~m[594]&m[595]&~m[596]&m[620])|(m[593]&m[594]&~m[595]&m[596]&m[620])|(m[593]&~m[594]&m[595]&m[596]&m[620])|(~m[593]&m[594]&m[595]&m[596]&m[620]))&~BiasedRNG[540])|((m[593]&m[594]&~m[595]&~m[596]&~m[620])|(m[593]&~m[594]&m[595]&~m[596]&~m[620])|(~m[593]&m[594]&m[595]&~m[596]&~m[620])|(m[593]&m[594]&m[595]&~m[596]&~m[620])|(m[593]&m[594]&m[595]&m[596]&~m[620])|(m[593]&m[594]&~m[595]&~m[596]&m[620])|(m[593]&~m[594]&m[595]&~m[596]&m[620])|(~m[593]&m[594]&m[595]&~m[596]&m[620])|(m[593]&m[594]&m[595]&~m[596]&m[620])|(m[593]&m[594]&m[595]&m[596]&m[620]));
    m[602] = (((m[598]&~m[599]&~m[600]&~m[601]&~m[625])|(~m[598]&m[599]&~m[600]&~m[601]&~m[625])|(~m[598]&~m[599]&m[600]&~m[601]&~m[625])|(m[598]&m[599]&~m[600]&m[601]&~m[625])|(m[598]&~m[599]&m[600]&m[601]&~m[625])|(~m[598]&m[599]&m[600]&m[601]&~m[625]))&BiasedRNG[541])|(((m[598]&~m[599]&~m[600]&~m[601]&m[625])|(~m[598]&m[599]&~m[600]&~m[601]&m[625])|(~m[598]&~m[599]&m[600]&~m[601]&m[625])|(m[598]&m[599]&~m[600]&m[601]&m[625])|(m[598]&~m[599]&m[600]&m[601]&m[625])|(~m[598]&m[599]&m[600]&m[601]&m[625]))&~BiasedRNG[541])|((m[598]&m[599]&~m[600]&~m[601]&~m[625])|(m[598]&~m[599]&m[600]&~m[601]&~m[625])|(~m[598]&m[599]&m[600]&~m[601]&~m[625])|(m[598]&m[599]&m[600]&~m[601]&~m[625])|(m[598]&m[599]&m[600]&m[601]&~m[625])|(m[598]&m[599]&~m[600]&~m[601]&m[625])|(m[598]&~m[599]&m[600]&~m[601]&m[625])|(~m[598]&m[599]&m[600]&~m[601]&m[625])|(m[598]&m[599]&m[600]&~m[601]&m[625])|(m[598]&m[599]&m[600]&m[601]&m[625]));
    m[607] = (((m[603]&~m[604]&~m[605]&~m[606]&~m[635])|(~m[603]&m[604]&~m[605]&~m[606]&~m[635])|(~m[603]&~m[604]&m[605]&~m[606]&~m[635])|(m[603]&m[604]&~m[605]&m[606]&~m[635])|(m[603]&~m[604]&m[605]&m[606]&~m[635])|(~m[603]&m[604]&m[605]&m[606]&~m[635]))&BiasedRNG[542])|(((m[603]&~m[604]&~m[605]&~m[606]&m[635])|(~m[603]&m[604]&~m[605]&~m[606]&m[635])|(~m[603]&~m[604]&m[605]&~m[606]&m[635])|(m[603]&m[604]&~m[605]&m[606]&m[635])|(m[603]&~m[604]&m[605]&m[606]&m[635])|(~m[603]&m[604]&m[605]&m[606]&m[635]))&~BiasedRNG[542])|((m[603]&m[604]&~m[605]&~m[606]&~m[635])|(m[603]&~m[604]&m[605]&~m[606]&~m[635])|(~m[603]&m[604]&m[605]&~m[606]&~m[635])|(m[603]&m[604]&m[605]&~m[606]&~m[635])|(m[603]&m[604]&m[605]&m[606]&~m[635])|(m[603]&m[604]&~m[605]&~m[606]&m[635])|(m[603]&~m[604]&m[605]&~m[606]&m[635])|(~m[603]&m[604]&m[605]&~m[606]&m[635])|(m[603]&m[604]&m[605]&~m[606]&m[635])|(m[603]&m[604]&m[605]&m[606]&m[635]));
    m[612] = (((m[608]&~m[609]&~m[610]&~m[611]&~m[640])|(~m[608]&m[609]&~m[610]&~m[611]&~m[640])|(~m[608]&~m[609]&m[610]&~m[611]&~m[640])|(m[608]&m[609]&~m[610]&m[611]&~m[640])|(m[608]&~m[609]&m[610]&m[611]&~m[640])|(~m[608]&m[609]&m[610]&m[611]&~m[640]))&BiasedRNG[543])|(((m[608]&~m[609]&~m[610]&~m[611]&m[640])|(~m[608]&m[609]&~m[610]&~m[611]&m[640])|(~m[608]&~m[609]&m[610]&~m[611]&m[640])|(m[608]&m[609]&~m[610]&m[611]&m[640])|(m[608]&~m[609]&m[610]&m[611]&m[640])|(~m[608]&m[609]&m[610]&m[611]&m[640]))&~BiasedRNG[543])|((m[608]&m[609]&~m[610]&~m[611]&~m[640])|(m[608]&~m[609]&m[610]&~m[611]&~m[640])|(~m[608]&m[609]&m[610]&~m[611]&~m[640])|(m[608]&m[609]&m[610]&~m[611]&~m[640])|(m[608]&m[609]&m[610]&m[611]&~m[640])|(m[608]&m[609]&~m[610]&~m[611]&m[640])|(m[608]&~m[609]&m[610]&~m[611]&m[640])|(~m[608]&m[609]&m[610]&~m[611]&m[640])|(m[608]&m[609]&m[610]&~m[611]&m[640])|(m[608]&m[609]&m[610]&m[611]&m[640]));
    m[617] = (((m[613]&~m[614]&~m[615]&~m[616]&~m[645])|(~m[613]&m[614]&~m[615]&~m[616]&~m[645])|(~m[613]&~m[614]&m[615]&~m[616]&~m[645])|(m[613]&m[614]&~m[615]&m[616]&~m[645])|(m[613]&~m[614]&m[615]&m[616]&~m[645])|(~m[613]&m[614]&m[615]&m[616]&~m[645]))&BiasedRNG[544])|(((m[613]&~m[614]&~m[615]&~m[616]&m[645])|(~m[613]&m[614]&~m[615]&~m[616]&m[645])|(~m[613]&~m[614]&m[615]&~m[616]&m[645])|(m[613]&m[614]&~m[615]&m[616]&m[645])|(m[613]&~m[614]&m[615]&m[616]&m[645])|(~m[613]&m[614]&m[615]&m[616]&m[645]))&~BiasedRNG[544])|((m[613]&m[614]&~m[615]&~m[616]&~m[645])|(m[613]&~m[614]&m[615]&~m[616]&~m[645])|(~m[613]&m[614]&m[615]&~m[616]&~m[645])|(m[613]&m[614]&m[615]&~m[616]&~m[645])|(m[613]&m[614]&m[615]&m[616]&~m[645])|(m[613]&m[614]&~m[615]&~m[616]&m[645])|(m[613]&~m[614]&m[615]&~m[616]&m[645])|(~m[613]&m[614]&m[615]&~m[616]&m[645])|(m[613]&m[614]&m[615]&~m[616]&m[645])|(m[613]&m[614]&m[615]&m[616]&m[645]));
    m[622] = (((m[618]&~m[619]&~m[620]&~m[621]&~m[650])|(~m[618]&m[619]&~m[620]&~m[621]&~m[650])|(~m[618]&~m[619]&m[620]&~m[621]&~m[650])|(m[618]&m[619]&~m[620]&m[621]&~m[650])|(m[618]&~m[619]&m[620]&m[621]&~m[650])|(~m[618]&m[619]&m[620]&m[621]&~m[650]))&BiasedRNG[545])|(((m[618]&~m[619]&~m[620]&~m[621]&m[650])|(~m[618]&m[619]&~m[620]&~m[621]&m[650])|(~m[618]&~m[619]&m[620]&~m[621]&m[650])|(m[618]&m[619]&~m[620]&m[621]&m[650])|(m[618]&~m[619]&m[620]&m[621]&m[650])|(~m[618]&m[619]&m[620]&m[621]&m[650]))&~BiasedRNG[545])|((m[618]&m[619]&~m[620]&~m[621]&~m[650])|(m[618]&~m[619]&m[620]&~m[621]&~m[650])|(~m[618]&m[619]&m[620]&~m[621]&~m[650])|(m[618]&m[619]&m[620]&~m[621]&~m[650])|(m[618]&m[619]&m[620]&m[621]&~m[650])|(m[618]&m[619]&~m[620]&~m[621]&m[650])|(m[618]&~m[619]&m[620]&~m[621]&m[650])|(~m[618]&m[619]&m[620]&~m[621]&m[650])|(m[618]&m[619]&m[620]&~m[621]&m[650])|(m[618]&m[619]&m[620]&m[621]&m[650]));
    m[627] = (((m[623]&~m[624]&~m[625]&~m[626]&~m[655])|(~m[623]&m[624]&~m[625]&~m[626]&~m[655])|(~m[623]&~m[624]&m[625]&~m[626]&~m[655])|(m[623]&m[624]&~m[625]&m[626]&~m[655])|(m[623]&~m[624]&m[625]&m[626]&~m[655])|(~m[623]&m[624]&m[625]&m[626]&~m[655]))&BiasedRNG[546])|(((m[623]&~m[624]&~m[625]&~m[626]&m[655])|(~m[623]&m[624]&~m[625]&~m[626]&m[655])|(~m[623]&~m[624]&m[625]&~m[626]&m[655])|(m[623]&m[624]&~m[625]&m[626]&m[655])|(m[623]&~m[624]&m[625]&m[626]&m[655])|(~m[623]&m[624]&m[625]&m[626]&m[655]))&~BiasedRNG[546])|((m[623]&m[624]&~m[625]&~m[626]&~m[655])|(m[623]&~m[624]&m[625]&~m[626]&~m[655])|(~m[623]&m[624]&m[625]&~m[626]&~m[655])|(m[623]&m[624]&m[625]&~m[626]&~m[655])|(m[623]&m[624]&m[625]&m[626]&~m[655])|(m[623]&m[624]&~m[625]&~m[626]&m[655])|(m[623]&~m[624]&m[625]&~m[626]&m[655])|(~m[623]&m[624]&m[625]&~m[626]&m[655])|(m[623]&m[624]&m[625]&~m[626]&m[655])|(m[623]&m[624]&m[625]&m[626]&m[655]));
    m[632] = (((m[628]&~m[629]&~m[630]&~m[631]&~m[660])|(~m[628]&m[629]&~m[630]&~m[631]&~m[660])|(~m[628]&~m[629]&m[630]&~m[631]&~m[660])|(m[628]&m[629]&~m[630]&m[631]&~m[660])|(m[628]&~m[629]&m[630]&m[631]&~m[660])|(~m[628]&m[629]&m[630]&m[631]&~m[660]))&BiasedRNG[547])|(((m[628]&~m[629]&~m[630]&~m[631]&m[660])|(~m[628]&m[629]&~m[630]&~m[631]&m[660])|(~m[628]&~m[629]&m[630]&~m[631]&m[660])|(m[628]&m[629]&~m[630]&m[631]&m[660])|(m[628]&~m[629]&m[630]&m[631]&m[660])|(~m[628]&m[629]&m[630]&m[631]&m[660]))&~BiasedRNG[547])|((m[628]&m[629]&~m[630]&~m[631]&~m[660])|(m[628]&~m[629]&m[630]&~m[631]&~m[660])|(~m[628]&m[629]&m[630]&~m[631]&~m[660])|(m[628]&m[629]&m[630]&~m[631]&~m[660])|(m[628]&m[629]&m[630]&m[631]&~m[660])|(m[628]&m[629]&~m[630]&~m[631]&m[660])|(m[628]&~m[629]&m[630]&~m[631]&m[660])|(~m[628]&m[629]&m[630]&~m[631]&m[660])|(m[628]&m[629]&m[630]&~m[631]&m[660])|(m[628]&m[629]&m[630]&m[631]&m[660]));
    m[637] = (((m[633]&~m[634]&~m[635]&~m[636]&~m[670])|(~m[633]&m[634]&~m[635]&~m[636]&~m[670])|(~m[633]&~m[634]&m[635]&~m[636]&~m[670])|(m[633]&m[634]&~m[635]&m[636]&~m[670])|(m[633]&~m[634]&m[635]&m[636]&~m[670])|(~m[633]&m[634]&m[635]&m[636]&~m[670]))&BiasedRNG[548])|(((m[633]&~m[634]&~m[635]&~m[636]&m[670])|(~m[633]&m[634]&~m[635]&~m[636]&m[670])|(~m[633]&~m[634]&m[635]&~m[636]&m[670])|(m[633]&m[634]&~m[635]&m[636]&m[670])|(m[633]&~m[634]&m[635]&m[636]&m[670])|(~m[633]&m[634]&m[635]&m[636]&m[670]))&~BiasedRNG[548])|((m[633]&m[634]&~m[635]&~m[636]&~m[670])|(m[633]&~m[634]&m[635]&~m[636]&~m[670])|(~m[633]&m[634]&m[635]&~m[636]&~m[670])|(m[633]&m[634]&m[635]&~m[636]&~m[670])|(m[633]&m[634]&m[635]&m[636]&~m[670])|(m[633]&m[634]&~m[635]&~m[636]&m[670])|(m[633]&~m[634]&m[635]&~m[636]&m[670])|(~m[633]&m[634]&m[635]&~m[636]&m[670])|(m[633]&m[634]&m[635]&~m[636]&m[670])|(m[633]&m[634]&m[635]&m[636]&m[670]));
    m[642] = (((m[638]&~m[639]&~m[640]&~m[641]&~m[675])|(~m[638]&m[639]&~m[640]&~m[641]&~m[675])|(~m[638]&~m[639]&m[640]&~m[641]&~m[675])|(m[638]&m[639]&~m[640]&m[641]&~m[675])|(m[638]&~m[639]&m[640]&m[641]&~m[675])|(~m[638]&m[639]&m[640]&m[641]&~m[675]))&BiasedRNG[549])|(((m[638]&~m[639]&~m[640]&~m[641]&m[675])|(~m[638]&m[639]&~m[640]&~m[641]&m[675])|(~m[638]&~m[639]&m[640]&~m[641]&m[675])|(m[638]&m[639]&~m[640]&m[641]&m[675])|(m[638]&~m[639]&m[640]&m[641]&m[675])|(~m[638]&m[639]&m[640]&m[641]&m[675]))&~BiasedRNG[549])|((m[638]&m[639]&~m[640]&~m[641]&~m[675])|(m[638]&~m[639]&m[640]&~m[641]&~m[675])|(~m[638]&m[639]&m[640]&~m[641]&~m[675])|(m[638]&m[639]&m[640]&~m[641]&~m[675])|(m[638]&m[639]&m[640]&m[641]&~m[675])|(m[638]&m[639]&~m[640]&~m[641]&m[675])|(m[638]&~m[639]&m[640]&~m[641]&m[675])|(~m[638]&m[639]&m[640]&~m[641]&m[675])|(m[638]&m[639]&m[640]&~m[641]&m[675])|(m[638]&m[639]&m[640]&m[641]&m[675]));
    m[647] = (((m[643]&~m[644]&~m[645]&~m[646]&~m[680])|(~m[643]&m[644]&~m[645]&~m[646]&~m[680])|(~m[643]&~m[644]&m[645]&~m[646]&~m[680])|(m[643]&m[644]&~m[645]&m[646]&~m[680])|(m[643]&~m[644]&m[645]&m[646]&~m[680])|(~m[643]&m[644]&m[645]&m[646]&~m[680]))&BiasedRNG[550])|(((m[643]&~m[644]&~m[645]&~m[646]&m[680])|(~m[643]&m[644]&~m[645]&~m[646]&m[680])|(~m[643]&~m[644]&m[645]&~m[646]&m[680])|(m[643]&m[644]&~m[645]&m[646]&m[680])|(m[643]&~m[644]&m[645]&m[646]&m[680])|(~m[643]&m[644]&m[645]&m[646]&m[680]))&~BiasedRNG[550])|((m[643]&m[644]&~m[645]&~m[646]&~m[680])|(m[643]&~m[644]&m[645]&~m[646]&~m[680])|(~m[643]&m[644]&m[645]&~m[646]&~m[680])|(m[643]&m[644]&m[645]&~m[646]&~m[680])|(m[643]&m[644]&m[645]&m[646]&~m[680])|(m[643]&m[644]&~m[645]&~m[646]&m[680])|(m[643]&~m[644]&m[645]&~m[646]&m[680])|(~m[643]&m[644]&m[645]&~m[646]&m[680])|(m[643]&m[644]&m[645]&~m[646]&m[680])|(m[643]&m[644]&m[645]&m[646]&m[680]));
    m[652] = (((m[648]&~m[649]&~m[650]&~m[651]&~m[685])|(~m[648]&m[649]&~m[650]&~m[651]&~m[685])|(~m[648]&~m[649]&m[650]&~m[651]&~m[685])|(m[648]&m[649]&~m[650]&m[651]&~m[685])|(m[648]&~m[649]&m[650]&m[651]&~m[685])|(~m[648]&m[649]&m[650]&m[651]&~m[685]))&BiasedRNG[551])|(((m[648]&~m[649]&~m[650]&~m[651]&m[685])|(~m[648]&m[649]&~m[650]&~m[651]&m[685])|(~m[648]&~m[649]&m[650]&~m[651]&m[685])|(m[648]&m[649]&~m[650]&m[651]&m[685])|(m[648]&~m[649]&m[650]&m[651]&m[685])|(~m[648]&m[649]&m[650]&m[651]&m[685]))&~BiasedRNG[551])|((m[648]&m[649]&~m[650]&~m[651]&~m[685])|(m[648]&~m[649]&m[650]&~m[651]&~m[685])|(~m[648]&m[649]&m[650]&~m[651]&~m[685])|(m[648]&m[649]&m[650]&~m[651]&~m[685])|(m[648]&m[649]&m[650]&m[651]&~m[685])|(m[648]&m[649]&~m[650]&~m[651]&m[685])|(m[648]&~m[649]&m[650]&~m[651]&m[685])|(~m[648]&m[649]&m[650]&~m[651]&m[685])|(m[648]&m[649]&m[650]&~m[651]&m[685])|(m[648]&m[649]&m[650]&m[651]&m[685]));
    m[657] = (((m[653]&~m[654]&~m[655]&~m[656]&~m[690])|(~m[653]&m[654]&~m[655]&~m[656]&~m[690])|(~m[653]&~m[654]&m[655]&~m[656]&~m[690])|(m[653]&m[654]&~m[655]&m[656]&~m[690])|(m[653]&~m[654]&m[655]&m[656]&~m[690])|(~m[653]&m[654]&m[655]&m[656]&~m[690]))&BiasedRNG[552])|(((m[653]&~m[654]&~m[655]&~m[656]&m[690])|(~m[653]&m[654]&~m[655]&~m[656]&m[690])|(~m[653]&~m[654]&m[655]&~m[656]&m[690])|(m[653]&m[654]&~m[655]&m[656]&m[690])|(m[653]&~m[654]&m[655]&m[656]&m[690])|(~m[653]&m[654]&m[655]&m[656]&m[690]))&~BiasedRNG[552])|((m[653]&m[654]&~m[655]&~m[656]&~m[690])|(m[653]&~m[654]&m[655]&~m[656]&~m[690])|(~m[653]&m[654]&m[655]&~m[656]&~m[690])|(m[653]&m[654]&m[655]&~m[656]&~m[690])|(m[653]&m[654]&m[655]&m[656]&~m[690])|(m[653]&m[654]&~m[655]&~m[656]&m[690])|(m[653]&~m[654]&m[655]&~m[656]&m[690])|(~m[653]&m[654]&m[655]&~m[656]&m[690])|(m[653]&m[654]&m[655]&~m[656]&m[690])|(m[653]&m[654]&m[655]&m[656]&m[690]));
    m[662] = (((m[658]&~m[659]&~m[660]&~m[661]&~m[695])|(~m[658]&m[659]&~m[660]&~m[661]&~m[695])|(~m[658]&~m[659]&m[660]&~m[661]&~m[695])|(m[658]&m[659]&~m[660]&m[661]&~m[695])|(m[658]&~m[659]&m[660]&m[661]&~m[695])|(~m[658]&m[659]&m[660]&m[661]&~m[695]))&BiasedRNG[553])|(((m[658]&~m[659]&~m[660]&~m[661]&m[695])|(~m[658]&m[659]&~m[660]&~m[661]&m[695])|(~m[658]&~m[659]&m[660]&~m[661]&m[695])|(m[658]&m[659]&~m[660]&m[661]&m[695])|(m[658]&~m[659]&m[660]&m[661]&m[695])|(~m[658]&m[659]&m[660]&m[661]&m[695]))&~BiasedRNG[553])|((m[658]&m[659]&~m[660]&~m[661]&~m[695])|(m[658]&~m[659]&m[660]&~m[661]&~m[695])|(~m[658]&m[659]&m[660]&~m[661]&~m[695])|(m[658]&m[659]&m[660]&~m[661]&~m[695])|(m[658]&m[659]&m[660]&m[661]&~m[695])|(m[658]&m[659]&~m[660]&~m[661]&m[695])|(m[658]&~m[659]&m[660]&~m[661]&m[695])|(~m[658]&m[659]&m[660]&~m[661]&m[695])|(m[658]&m[659]&m[660]&~m[661]&m[695])|(m[658]&m[659]&m[660]&m[661]&m[695]));
    m[667] = (((m[663]&~m[664]&~m[665]&~m[666]&~m[700])|(~m[663]&m[664]&~m[665]&~m[666]&~m[700])|(~m[663]&~m[664]&m[665]&~m[666]&~m[700])|(m[663]&m[664]&~m[665]&m[666]&~m[700])|(m[663]&~m[664]&m[665]&m[666]&~m[700])|(~m[663]&m[664]&m[665]&m[666]&~m[700]))&BiasedRNG[554])|(((m[663]&~m[664]&~m[665]&~m[666]&m[700])|(~m[663]&m[664]&~m[665]&~m[666]&m[700])|(~m[663]&~m[664]&m[665]&~m[666]&m[700])|(m[663]&m[664]&~m[665]&m[666]&m[700])|(m[663]&~m[664]&m[665]&m[666]&m[700])|(~m[663]&m[664]&m[665]&m[666]&m[700]))&~BiasedRNG[554])|((m[663]&m[664]&~m[665]&~m[666]&~m[700])|(m[663]&~m[664]&m[665]&~m[666]&~m[700])|(~m[663]&m[664]&m[665]&~m[666]&~m[700])|(m[663]&m[664]&m[665]&~m[666]&~m[700])|(m[663]&m[664]&m[665]&m[666]&~m[700])|(m[663]&m[664]&~m[665]&~m[666]&m[700])|(m[663]&~m[664]&m[665]&~m[666]&m[700])|(~m[663]&m[664]&m[665]&~m[666]&m[700])|(m[663]&m[664]&m[665]&~m[666]&m[700])|(m[663]&m[664]&m[665]&m[666]&m[700]));
    m[672] = (((m[668]&~m[669]&~m[670]&~m[671]&~m[710])|(~m[668]&m[669]&~m[670]&~m[671]&~m[710])|(~m[668]&~m[669]&m[670]&~m[671]&~m[710])|(m[668]&m[669]&~m[670]&m[671]&~m[710])|(m[668]&~m[669]&m[670]&m[671]&~m[710])|(~m[668]&m[669]&m[670]&m[671]&~m[710]))&BiasedRNG[555])|(((m[668]&~m[669]&~m[670]&~m[671]&m[710])|(~m[668]&m[669]&~m[670]&~m[671]&m[710])|(~m[668]&~m[669]&m[670]&~m[671]&m[710])|(m[668]&m[669]&~m[670]&m[671]&m[710])|(m[668]&~m[669]&m[670]&m[671]&m[710])|(~m[668]&m[669]&m[670]&m[671]&m[710]))&~BiasedRNG[555])|((m[668]&m[669]&~m[670]&~m[671]&~m[710])|(m[668]&~m[669]&m[670]&~m[671]&~m[710])|(~m[668]&m[669]&m[670]&~m[671]&~m[710])|(m[668]&m[669]&m[670]&~m[671]&~m[710])|(m[668]&m[669]&m[670]&m[671]&~m[710])|(m[668]&m[669]&~m[670]&~m[671]&m[710])|(m[668]&~m[669]&m[670]&~m[671]&m[710])|(~m[668]&m[669]&m[670]&~m[671]&m[710])|(m[668]&m[669]&m[670]&~m[671]&m[710])|(m[668]&m[669]&m[670]&m[671]&m[710]));
    m[677] = (((m[673]&~m[674]&~m[675]&~m[676]&~m[715])|(~m[673]&m[674]&~m[675]&~m[676]&~m[715])|(~m[673]&~m[674]&m[675]&~m[676]&~m[715])|(m[673]&m[674]&~m[675]&m[676]&~m[715])|(m[673]&~m[674]&m[675]&m[676]&~m[715])|(~m[673]&m[674]&m[675]&m[676]&~m[715]))&BiasedRNG[556])|(((m[673]&~m[674]&~m[675]&~m[676]&m[715])|(~m[673]&m[674]&~m[675]&~m[676]&m[715])|(~m[673]&~m[674]&m[675]&~m[676]&m[715])|(m[673]&m[674]&~m[675]&m[676]&m[715])|(m[673]&~m[674]&m[675]&m[676]&m[715])|(~m[673]&m[674]&m[675]&m[676]&m[715]))&~BiasedRNG[556])|((m[673]&m[674]&~m[675]&~m[676]&~m[715])|(m[673]&~m[674]&m[675]&~m[676]&~m[715])|(~m[673]&m[674]&m[675]&~m[676]&~m[715])|(m[673]&m[674]&m[675]&~m[676]&~m[715])|(m[673]&m[674]&m[675]&m[676]&~m[715])|(m[673]&m[674]&~m[675]&~m[676]&m[715])|(m[673]&~m[674]&m[675]&~m[676]&m[715])|(~m[673]&m[674]&m[675]&~m[676]&m[715])|(m[673]&m[674]&m[675]&~m[676]&m[715])|(m[673]&m[674]&m[675]&m[676]&m[715]));
    m[682] = (((m[678]&~m[679]&~m[680]&~m[681]&~m[720])|(~m[678]&m[679]&~m[680]&~m[681]&~m[720])|(~m[678]&~m[679]&m[680]&~m[681]&~m[720])|(m[678]&m[679]&~m[680]&m[681]&~m[720])|(m[678]&~m[679]&m[680]&m[681]&~m[720])|(~m[678]&m[679]&m[680]&m[681]&~m[720]))&BiasedRNG[557])|(((m[678]&~m[679]&~m[680]&~m[681]&m[720])|(~m[678]&m[679]&~m[680]&~m[681]&m[720])|(~m[678]&~m[679]&m[680]&~m[681]&m[720])|(m[678]&m[679]&~m[680]&m[681]&m[720])|(m[678]&~m[679]&m[680]&m[681]&m[720])|(~m[678]&m[679]&m[680]&m[681]&m[720]))&~BiasedRNG[557])|((m[678]&m[679]&~m[680]&~m[681]&~m[720])|(m[678]&~m[679]&m[680]&~m[681]&~m[720])|(~m[678]&m[679]&m[680]&~m[681]&~m[720])|(m[678]&m[679]&m[680]&~m[681]&~m[720])|(m[678]&m[679]&m[680]&m[681]&~m[720])|(m[678]&m[679]&~m[680]&~m[681]&m[720])|(m[678]&~m[679]&m[680]&~m[681]&m[720])|(~m[678]&m[679]&m[680]&~m[681]&m[720])|(m[678]&m[679]&m[680]&~m[681]&m[720])|(m[678]&m[679]&m[680]&m[681]&m[720]));
    m[687] = (((m[683]&~m[684]&~m[685]&~m[686]&~m[725])|(~m[683]&m[684]&~m[685]&~m[686]&~m[725])|(~m[683]&~m[684]&m[685]&~m[686]&~m[725])|(m[683]&m[684]&~m[685]&m[686]&~m[725])|(m[683]&~m[684]&m[685]&m[686]&~m[725])|(~m[683]&m[684]&m[685]&m[686]&~m[725]))&BiasedRNG[558])|(((m[683]&~m[684]&~m[685]&~m[686]&m[725])|(~m[683]&m[684]&~m[685]&~m[686]&m[725])|(~m[683]&~m[684]&m[685]&~m[686]&m[725])|(m[683]&m[684]&~m[685]&m[686]&m[725])|(m[683]&~m[684]&m[685]&m[686]&m[725])|(~m[683]&m[684]&m[685]&m[686]&m[725]))&~BiasedRNG[558])|((m[683]&m[684]&~m[685]&~m[686]&~m[725])|(m[683]&~m[684]&m[685]&~m[686]&~m[725])|(~m[683]&m[684]&m[685]&~m[686]&~m[725])|(m[683]&m[684]&m[685]&~m[686]&~m[725])|(m[683]&m[684]&m[685]&m[686]&~m[725])|(m[683]&m[684]&~m[685]&~m[686]&m[725])|(m[683]&~m[684]&m[685]&~m[686]&m[725])|(~m[683]&m[684]&m[685]&~m[686]&m[725])|(m[683]&m[684]&m[685]&~m[686]&m[725])|(m[683]&m[684]&m[685]&m[686]&m[725]));
    m[692] = (((m[688]&~m[689]&~m[690]&~m[691]&~m[730])|(~m[688]&m[689]&~m[690]&~m[691]&~m[730])|(~m[688]&~m[689]&m[690]&~m[691]&~m[730])|(m[688]&m[689]&~m[690]&m[691]&~m[730])|(m[688]&~m[689]&m[690]&m[691]&~m[730])|(~m[688]&m[689]&m[690]&m[691]&~m[730]))&BiasedRNG[559])|(((m[688]&~m[689]&~m[690]&~m[691]&m[730])|(~m[688]&m[689]&~m[690]&~m[691]&m[730])|(~m[688]&~m[689]&m[690]&~m[691]&m[730])|(m[688]&m[689]&~m[690]&m[691]&m[730])|(m[688]&~m[689]&m[690]&m[691]&m[730])|(~m[688]&m[689]&m[690]&m[691]&m[730]))&~BiasedRNG[559])|((m[688]&m[689]&~m[690]&~m[691]&~m[730])|(m[688]&~m[689]&m[690]&~m[691]&~m[730])|(~m[688]&m[689]&m[690]&~m[691]&~m[730])|(m[688]&m[689]&m[690]&~m[691]&~m[730])|(m[688]&m[689]&m[690]&m[691]&~m[730])|(m[688]&m[689]&~m[690]&~m[691]&m[730])|(m[688]&~m[689]&m[690]&~m[691]&m[730])|(~m[688]&m[689]&m[690]&~m[691]&m[730])|(m[688]&m[689]&m[690]&~m[691]&m[730])|(m[688]&m[689]&m[690]&m[691]&m[730]));
    m[697] = (((m[693]&~m[694]&~m[695]&~m[696]&~m[735])|(~m[693]&m[694]&~m[695]&~m[696]&~m[735])|(~m[693]&~m[694]&m[695]&~m[696]&~m[735])|(m[693]&m[694]&~m[695]&m[696]&~m[735])|(m[693]&~m[694]&m[695]&m[696]&~m[735])|(~m[693]&m[694]&m[695]&m[696]&~m[735]))&BiasedRNG[560])|(((m[693]&~m[694]&~m[695]&~m[696]&m[735])|(~m[693]&m[694]&~m[695]&~m[696]&m[735])|(~m[693]&~m[694]&m[695]&~m[696]&m[735])|(m[693]&m[694]&~m[695]&m[696]&m[735])|(m[693]&~m[694]&m[695]&m[696]&m[735])|(~m[693]&m[694]&m[695]&m[696]&m[735]))&~BiasedRNG[560])|((m[693]&m[694]&~m[695]&~m[696]&~m[735])|(m[693]&~m[694]&m[695]&~m[696]&~m[735])|(~m[693]&m[694]&m[695]&~m[696]&~m[735])|(m[693]&m[694]&m[695]&~m[696]&~m[735])|(m[693]&m[694]&m[695]&m[696]&~m[735])|(m[693]&m[694]&~m[695]&~m[696]&m[735])|(m[693]&~m[694]&m[695]&~m[696]&m[735])|(~m[693]&m[694]&m[695]&~m[696]&m[735])|(m[693]&m[694]&m[695]&~m[696]&m[735])|(m[693]&m[694]&m[695]&m[696]&m[735]));
    m[702] = (((m[698]&~m[699]&~m[700]&~m[701]&~m[740])|(~m[698]&m[699]&~m[700]&~m[701]&~m[740])|(~m[698]&~m[699]&m[700]&~m[701]&~m[740])|(m[698]&m[699]&~m[700]&m[701]&~m[740])|(m[698]&~m[699]&m[700]&m[701]&~m[740])|(~m[698]&m[699]&m[700]&m[701]&~m[740]))&BiasedRNG[561])|(((m[698]&~m[699]&~m[700]&~m[701]&m[740])|(~m[698]&m[699]&~m[700]&~m[701]&m[740])|(~m[698]&~m[699]&m[700]&~m[701]&m[740])|(m[698]&m[699]&~m[700]&m[701]&m[740])|(m[698]&~m[699]&m[700]&m[701]&m[740])|(~m[698]&m[699]&m[700]&m[701]&m[740]))&~BiasedRNG[561])|((m[698]&m[699]&~m[700]&~m[701]&~m[740])|(m[698]&~m[699]&m[700]&~m[701]&~m[740])|(~m[698]&m[699]&m[700]&~m[701]&~m[740])|(m[698]&m[699]&m[700]&~m[701]&~m[740])|(m[698]&m[699]&m[700]&m[701]&~m[740])|(m[698]&m[699]&~m[700]&~m[701]&m[740])|(m[698]&~m[699]&m[700]&~m[701]&m[740])|(~m[698]&m[699]&m[700]&~m[701]&m[740])|(m[698]&m[699]&m[700]&~m[701]&m[740])|(m[698]&m[699]&m[700]&m[701]&m[740]));
    m[707] = (((m[703]&~m[704]&~m[705]&~m[706]&~m[745])|(~m[703]&m[704]&~m[705]&~m[706]&~m[745])|(~m[703]&~m[704]&m[705]&~m[706]&~m[745])|(m[703]&m[704]&~m[705]&m[706]&~m[745])|(m[703]&~m[704]&m[705]&m[706]&~m[745])|(~m[703]&m[704]&m[705]&m[706]&~m[745]))&BiasedRNG[562])|(((m[703]&~m[704]&~m[705]&~m[706]&m[745])|(~m[703]&m[704]&~m[705]&~m[706]&m[745])|(~m[703]&~m[704]&m[705]&~m[706]&m[745])|(m[703]&m[704]&~m[705]&m[706]&m[745])|(m[703]&~m[704]&m[705]&m[706]&m[745])|(~m[703]&m[704]&m[705]&m[706]&m[745]))&~BiasedRNG[562])|((m[703]&m[704]&~m[705]&~m[706]&~m[745])|(m[703]&~m[704]&m[705]&~m[706]&~m[745])|(~m[703]&m[704]&m[705]&~m[706]&~m[745])|(m[703]&m[704]&m[705]&~m[706]&~m[745])|(m[703]&m[704]&m[705]&m[706]&~m[745])|(m[703]&m[704]&~m[705]&~m[706]&m[745])|(m[703]&~m[704]&m[705]&~m[706]&m[745])|(~m[703]&m[704]&m[705]&~m[706]&m[745])|(m[703]&m[704]&m[705]&~m[706]&m[745])|(m[703]&m[704]&m[705]&m[706]&m[745]));
    m[712] = (((m[708]&~m[709]&~m[710]&~m[711]&~m[755])|(~m[708]&m[709]&~m[710]&~m[711]&~m[755])|(~m[708]&~m[709]&m[710]&~m[711]&~m[755])|(m[708]&m[709]&~m[710]&m[711]&~m[755])|(m[708]&~m[709]&m[710]&m[711]&~m[755])|(~m[708]&m[709]&m[710]&m[711]&~m[755]))&BiasedRNG[563])|(((m[708]&~m[709]&~m[710]&~m[711]&m[755])|(~m[708]&m[709]&~m[710]&~m[711]&m[755])|(~m[708]&~m[709]&m[710]&~m[711]&m[755])|(m[708]&m[709]&~m[710]&m[711]&m[755])|(m[708]&~m[709]&m[710]&m[711]&m[755])|(~m[708]&m[709]&m[710]&m[711]&m[755]))&~BiasedRNG[563])|((m[708]&m[709]&~m[710]&~m[711]&~m[755])|(m[708]&~m[709]&m[710]&~m[711]&~m[755])|(~m[708]&m[709]&m[710]&~m[711]&~m[755])|(m[708]&m[709]&m[710]&~m[711]&~m[755])|(m[708]&m[709]&m[710]&m[711]&~m[755])|(m[708]&m[709]&~m[710]&~m[711]&m[755])|(m[708]&~m[709]&m[710]&~m[711]&m[755])|(~m[708]&m[709]&m[710]&~m[711]&m[755])|(m[708]&m[709]&m[710]&~m[711]&m[755])|(m[708]&m[709]&m[710]&m[711]&m[755]));
    m[717] = (((m[713]&~m[714]&~m[715]&~m[716]&~m[760])|(~m[713]&m[714]&~m[715]&~m[716]&~m[760])|(~m[713]&~m[714]&m[715]&~m[716]&~m[760])|(m[713]&m[714]&~m[715]&m[716]&~m[760])|(m[713]&~m[714]&m[715]&m[716]&~m[760])|(~m[713]&m[714]&m[715]&m[716]&~m[760]))&BiasedRNG[564])|(((m[713]&~m[714]&~m[715]&~m[716]&m[760])|(~m[713]&m[714]&~m[715]&~m[716]&m[760])|(~m[713]&~m[714]&m[715]&~m[716]&m[760])|(m[713]&m[714]&~m[715]&m[716]&m[760])|(m[713]&~m[714]&m[715]&m[716]&m[760])|(~m[713]&m[714]&m[715]&m[716]&m[760]))&~BiasedRNG[564])|((m[713]&m[714]&~m[715]&~m[716]&~m[760])|(m[713]&~m[714]&m[715]&~m[716]&~m[760])|(~m[713]&m[714]&m[715]&~m[716]&~m[760])|(m[713]&m[714]&m[715]&~m[716]&~m[760])|(m[713]&m[714]&m[715]&m[716]&~m[760])|(m[713]&m[714]&~m[715]&~m[716]&m[760])|(m[713]&~m[714]&m[715]&~m[716]&m[760])|(~m[713]&m[714]&m[715]&~m[716]&m[760])|(m[713]&m[714]&m[715]&~m[716]&m[760])|(m[713]&m[714]&m[715]&m[716]&m[760]));
    m[722] = (((m[718]&~m[719]&~m[720]&~m[721]&~m[765])|(~m[718]&m[719]&~m[720]&~m[721]&~m[765])|(~m[718]&~m[719]&m[720]&~m[721]&~m[765])|(m[718]&m[719]&~m[720]&m[721]&~m[765])|(m[718]&~m[719]&m[720]&m[721]&~m[765])|(~m[718]&m[719]&m[720]&m[721]&~m[765]))&BiasedRNG[565])|(((m[718]&~m[719]&~m[720]&~m[721]&m[765])|(~m[718]&m[719]&~m[720]&~m[721]&m[765])|(~m[718]&~m[719]&m[720]&~m[721]&m[765])|(m[718]&m[719]&~m[720]&m[721]&m[765])|(m[718]&~m[719]&m[720]&m[721]&m[765])|(~m[718]&m[719]&m[720]&m[721]&m[765]))&~BiasedRNG[565])|((m[718]&m[719]&~m[720]&~m[721]&~m[765])|(m[718]&~m[719]&m[720]&~m[721]&~m[765])|(~m[718]&m[719]&m[720]&~m[721]&~m[765])|(m[718]&m[719]&m[720]&~m[721]&~m[765])|(m[718]&m[719]&m[720]&m[721]&~m[765])|(m[718]&m[719]&~m[720]&~m[721]&m[765])|(m[718]&~m[719]&m[720]&~m[721]&m[765])|(~m[718]&m[719]&m[720]&~m[721]&m[765])|(m[718]&m[719]&m[720]&~m[721]&m[765])|(m[718]&m[719]&m[720]&m[721]&m[765]));
    m[727] = (((m[723]&~m[724]&~m[725]&~m[726]&~m[770])|(~m[723]&m[724]&~m[725]&~m[726]&~m[770])|(~m[723]&~m[724]&m[725]&~m[726]&~m[770])|(m[723]&m[724]&~m[725]&m[726]&~m[770])|(m[723]&~m[724]&m[725]&m[726]&~m[770])|(~m[723]&m[724]&m[725]&m[726]&~m[770]))&BiasedRNG[566])|(((m[723]&~m[724]&~m[725]&~m[726]&m[770])|(~m[723]&m[724]&~m[725]&~m[726]&m[770])|(~m[723]&~m[724]&m[725]&~m[726]&m[770])|(m[723]&m[724]&~m[725]&m[726]&m[770])|(m[723]&~m[724]&m[725]&m[726]&m[770])|(~m[723]&m[724]&m[725]&m[726]&m[770]))&~BiasedRNG[566])|((m[723]&m[724]&~m[725]&~m[726]&~m[770])|(m[723]&~m[724]&m[725]&~m[726]&~m[770])|(~m[723]&m[724]&m[725]&~m[726]&~m[770])|(m[723]&m[724]&m[725]&~m[726]&~m[770])|(m[723]&m[724]&m[725]&m[726]&~m[770])|(m[723]&m[724]&~m[725]&~m[726]&m[770])|(m[723]&~m[724]&m[725]&~m[726]&m[770])|(~m[723]&m[724]&m[725]&~m[726]&m[770])|(m[723]&m[724]&m[725]&~m[726]&m[770])|(m[723]&m[724]&m[725]&m[726]&m[770]));
    m[732] = (((m[728]&~m[729]&~m[730]&~m[731]&~m[775])|(~m[728]&m[729]&~m[730]&~m[731]&~m[775])|(~m[728]&~m[729]&m[730]&~m[731]&~m[775])|(m[728]&m[729]&~m[730]&m[731]&~m[775])|(m[728]&~m[729]&m[730]&m[731]&~m[775])|(~m[728]&m[729]&m[730]&m[731]&~m[775]))&BiasedRNG[567])|(((m[728]&~m[729]&~m[730]&~m[731]&m[775])|(~m[728]&m[729]&~m[730]&~m[731]&m[775])|(~m[728]&~m[729]&m[730]&~m[731]&m[775])|(m[728]&m[729]&~m[730]&m[731]&m[775])|(m[728]&~m[729]&m[730]&m[731]&m[775])|(~m[728]&m[729]&m[730]&m[731]&m[775]))&~BiasedRNG[567])|((m[728]&m[729]&~m[730]&~m[731]&~m[775])|(m[728]&~m[729]&m[730]&~m[731]&~m[775])|(~m[728]&m[729]&m[730]&~m[731]&~m[775])|(m[728]&m[729]&m[730]&~m[731]&~m[775])|(m[728]&m[729]&m[730]&m[731]&~m[775])|(m[728]&m[729]&~m[730]&~m[731]&m[775])|(m[728]&~m[729]&m[730]&~m[731]&m[775])|(~m[728]&m[729]&m[730]&~m[731]&m[775])|(m[728]&m[729]&m[730]&~m[731]&m[775])|(m[728]&m[729]&m[730]&m[731]&m[775]));
    m[737] = (((m[733]&~m[734]&~m[735]&~m[736]&~m[780])|(~m[733]&m[734]&~m[735]&~m[736]&~m[780])|(~m[733]&~m[734]&m[735]&~m[736]&~m[780])|(m[733]&m[734]&~m[735]&m[736]&~m[780])|(m[733]&~m[734]&m[735]&m[736]&~m[780])|(~m[733]&m[734]&m[735]&m[736]&~m[780]))&BiasedRNG[568])|(((m[733]&~m[734]&~m[735]&~m[736]&m[780])|(~m[733]&m[734]&~m[735]&~m[736]&m[780])|(~m[733]&~m[734]&m[735]&~m[736]&m[780])|(m[733]&m[734]&~m[735]&m[736]&m[780])|(m[733]&~m[734]&m[735]&m[736]&m[780])|(~m[733]&m[734]&m[735]&m[736]&m[780]))&~BiasedRNG[568])|((m[733]&m[734]&~m[735]&~m[736]&~m[780])|(m[733]&~m[734]&m[735]&~m[736]&~m[780])|(~m[733]&m[734]&m[735]&~m[736]&~m[780])|(m[733]&m[734]&m[735]&~m[736]&~m[780])|(m[733]&m[734]&m[735]&m[736]&~m[780])|(m[733]&m[734]&~m[735]&~m[736]&m[780])|(m[733]&~m[734]&m[735]&~m[736]&m[780])|(~m[733]&m[734]&m[735]&~m[736]&m[780])|(m[733]&m[734]&m[735]&~m[736]&m[780])|(m[733]&m[734]&m[735]&m[736]&m[780]));
    m[742] = (((m[738]&~m[739]&~m[740]&~m[741]&~m[785])|(~m[738]&m[739]&~m[740]&~m[741]&~m[785])|(~m[738]&~m[739]&m[740]&~m[741]&~m[785])|(m[738]&m[739]&~m[740]&m[741]&~m[785])|(m[738]&~m[739]&m[740]&m[741]&~m[785])|(~m[738]&m[739]&m[740]&m[741]&~m[785]))&BiasedRNG[569])|(((m[738]&~m[739]&~m[740]&~m[741]&m[785])|(~m[738]&m[739]&~m[740]&~m[741]&m[785])|(~m[738]&~m[739]&m[740]&~m[741]&m[785])|(m[738]&m[739]&~m[740]&m[741]&m[785])|(m[738]&~m[739]&m[740]&m[741]&m[785])|(~m[738]&m[739]&m[740]&m[741]&m[785]))&~BiasedRNG[569])|((m[738]&m[739]&~m[740]&~m[741]&~m[785])|(m[738]&~m[739]&m[740]&~m[741]&~m[785])|(~m[738]&m[739]&m[740]&~m[741]&~m[785])|(m[738]&m[739]&m[740]&~m[741]&~m[785])|(m[738]&m[739]&m[740]&m[741]&~m[785])|(m[738]&m[739]&~m[740]&~m[741]&m[785])|(m[738]&~m[739]&m[740]&~m[741]&m[785])|(~m[738]&m[739]&m[740]&~m[741]&m[785])|(m[738]&m[739]&m[740]&~m[741]&m[785])|(m[738]&m[739]&m[740]&m[741]&m[785]));
    m[747] = (((m[743]&~m[744]&~m[745]&~m[746]&~m[790])|(~m[743]&m[744]&~m[745]&~m[746]&~m[790])|(~m[743]&~m[744]&m[745]&~m[746]&~m[790])|(m[743]&m[744]&~m[745]&m[746]&~m[790])|(m[743]&~m[744]&m[745]&m[746]&~m[790])|(~m[743]&m[744]&m[745]&m[746]&~m[790]))&BiasedRNG[570])|(((m[743]&~m[744]&~m[745]&~m[746]&m[790])|(~m[743]&m[744]&~m[745]&~m[746]&m[790])|(~m[743]&~m[744]&m[745]&~m[746]&m[790])|(m[743]&m[744]&~m[745]&m[746]&m[790])|(m[743]&~m[744]&m[745]&m[746]&m[790])|(~m[743]&m[744]&m[745]&m[746]&m[790]))&~BiasedRNG[570])|((m[743]&m[744]&~m[745]&~m[746]&~m[790])|(m[743]&~m[744]&m[745]&~m[746]&~m[790])|(~m[743]&m[744]&m[745]&~m[746]&~m[790])|(m[743]&m[744]&m[745]&~m[746]&~m[790])|(m[743]&m[744]&m[745]&m[746]&~m[790])|(m[743]&m[744]&~m[745]&~m[746]&m[790])|(m[743]&~m[744]&m[745]&~m[746]&m[790])|(~m[743]&m[744]&m[745]&~m[746]&m[790])|(m[743]&m[744]&m[745]&~m[746]&m[790])|(m[743]&m[744]&m[745]&m[746]&m[790]));
    m[752] = (((m[748]&~m[749]&~m[750]&~m[751]&~m[795])|(~m[748]&m[749]&~m[750]&~m[751]&~m[795])|(~m[748]&~m[749]&m[750]&~m[751]&~m[795])|(m[748]&m[749]&~m[750]&m[751]&~m[795])|(m[748]&~m[749]&m[750]&m[751]&~m[795])|(~m[748]&m[749]&m[750]&m[751]&~m[795]))&BiasedRNG[571])|(((m[748]&~m[749]&~m[750]&~m[751]&m[795])|(~m[748]&m[749]&~m[750]&~m[751]&m[795])|(~m[748]&~m[749]&m[750]&~m[751]&m[795])|(m[748]&m[749]&~m[750]&m[751]&m[795])|(m[748]&~m[749]&m[750]&m[751]&m[795])|(~m[748]&m[749]&m[750]&m[751]&m[795]))&~BiasedRNG[571])|((m[748]&m[749]&~m[750]&~m[751]&~m[795])|(m[748]&~m[749]&m[750]&~m[751]&~m[795])|(~m[748]&m[749]&m[750]&~m[751]&~m[795])|(m[748]&m[749]&m[750]&~m[751]&~m[795])|(m[748]&m[749]&m[750]&m[751]&~m[795])|(m[748]&m[749]&~m[750]&~m[751]&m[795])|(m[748]&~m[749]&m[750]&~m[751]&m[795])|(~m[748]&m[749]&m[750]&~m[751]&m[795])|(m[748]&m[749]&m[750]&~m[751]&m[795])|(m[748]&m[749]&m[750]&m[751]&m[795]));
    m[757] = (((m[753]&~m[754]&~m[755]&~m[756]&~m[805])|(~m[753]&m[754]&~m[755]&~m[756]&~m[805])|(~m[753]&~m[754]&m[755]&~m[756]&~m[805])|(m[753]&m[754]&~m[755]&m[756]&~m[805])|(m[753]&~m[754]&m[755]&m[756]&~m[805])|(~m[753]&m[754]&m[755]&m[756]&~m[805]))&BiasedRNG[572])|(((m[753]&~m[754]&~m[755]&~m[756]&m[805])|(~m[753]&m[754]&~m[755]&~m[756]&m[805])|(~m[753]&~m[754]&m[755]&~m[756]&m[805])|(m[753]&m[754]&~m[755]&m[756]&m[805])|(m[753]&~m[754]&m[755]&m[756]&m[805])|(~m[753]&m[754]&m[755]&m[756]&m[805]))&~BiasedRNG[572])|((m[753]&m[754]&~m[755]&~m[756]&~m[805])|(m[753]&~m[754]&m[755]&~m[756]&~m[805])|(~m[753]&m[754]&m[755]&~m[756]&~m[805])|(m[753]&m[754]&m[755]&~m[756]&~m[805])|(m[753]&m[754]&m[755]&m[756]&~m[805])|(m[753]&m[754]&~m[755]&~m[756]&m[805])|(m[753]&~m[754]&m[755]&~m[756]&m[805])|(~m[753]&m[754]&m[755]&~m[756]&m[805])|(m[753]&m[754]&m[755]&~m[756]&m[805])|(m[753]&m[754]&m[755]&m[756]&m[805]));
    m[762] = (((m[758]&~m[759]&~m[760]&~m[761]&~m[810])|(~m[758]&m[759]&~m[760]&~m[761]&~m[810])|(~m[758]&~m[759]&m[760]&~m[761]&~m[810])|(m[758]&m[759]&~m[760]&m[761]&~m[810])|(m[758]&~m[759]&m[760]&m[761]&~m[810])|(~m[758]&m[759]&m[760]&m[761]&~m[810]))&BiasedRNG[573])|(((m[758]&~m[759]&~m[760]&~m[761]&m[810])|(~m[758]&m[759]&~m[760]&~m[761]&m[810])|(~m[758]&~m[759]&m[760]&~m[761]&m[810])|(m[758]&m[759]&~m[760]&m[761]&m[810])|(m[758]&~m[759]&m[760]&m[761]&m[810])|(~m[758]&m[759]&m[760]&m[761]&m[810]))&~BiasedRNG[573])|((m[758]&m[759]&~m[760]&~m[761]&~m[810])|(m[758]&~m[759]&m[760]&~m[761]&~m[810])|(~m[758]&m[759]&m[760]&~m[761]&~m[810])|(m[758]&m[759]&m[760]&~m[761]&~m[810])|(m[758]&m[759]&m[760]&m[761]&~m[810])|(m[758]&m[759]&~m[760]&~m[761]&m[810])|(m[758]&~m[759]&m[760]&~m[761]&m[810])|(~m[758]&m[759]&m[760]&~m[761]&m[810])|(m[758]&m[759]&m[760]&~m[761]&m[810])|(m[758]&m[759]&m[760]&m[761]&m[810]));
    m[767] = (((m[763]&~m[764]&~m[765]&~m[766]&~m[815])|(~m[763]&m[764]&~m[765]&~m[766]&~m[815])|(~m[763]&~m[764]&m[765]&~m[766]&~m[815])|(m[763]&m[764]&~m[765]&m[766]&~m[815])|(m[763]&~m[764]&m[765]&m[766]&~m[815])|(~m[763]&m[764]&m[765]&m[766]&~m[815]))&BiasedRNG[574])|(((m[763]&~m[764]&~m[765]&~m[766]&m[815])|(~m[763]&m[764]&~m[765]&~m[766]&m[815])|(~m[763]&~m[764]&m[765]&~m[766]&m[815])|(m[763]&m[764]&~m[765]&m[766]&m[815])|(m[763]&~m[764]&m[765]&m[766]&m[815])|(~m[763]&m[764]&m[765]&m[766]&m[815]))&~BiasedRNG[574])|((m[763]&m[764]&~m[765]&~m[766]&~m[815])|(m[763]&~m[764]&m[765]&~m[766]&~m[815])|(~m[763]&m[764]&m[765]&~m[766]&~m[815])|(m[763]&m[764]&m[765]&~m[766]&~m[815])|(m[763]&m[764]&m[765]&m[766]&~m[815])|(m[763]&m[764]&~m[765]&~m[766]&m[815])|(m[763]&~m[764]&m[765]&~m[766]&m[815])|(~m[763]&m[764]&m[765]&~m[766]&m[815])|(m[763]&m[764]&m[765]&~m[766]&m[815])|(m[763]&m[764]&m[765]&m[766]&m[815]));
    m[772] = (((m[768]&~m[769]&~m[770]&~m[771]&~m[820])|(~m[768]&m[769]&~m[770]&~m[771]&~m[820])|(~m[768]&~m[769]&m[770]&~m[771]&~m[820])|(m[768]&m[769]&~m[770]&m[771]&~m[820])|(m[768]&~m[769]&m[770]&m[771]&~m[820])|(~m[768]&m[769]&m[770]&m[771]&~m[820]))&BiasedRNG[575])|(((m[768]&~m[769]&~m[770]&~m[771]&m[820])|(~m[768]&m[769]&~m[770]&~m[771]&m[820])|(~m[768]&~m[769]&m[770]&~m[771]&m[820])|(m[768]&m[769]&~m[770]&m[771]&m[820])|(m[768]&~m[769]&m[770]&m[771]&m[820])|(~m[768]&m[769]&m[770]&m[771]&m[820]))&~BiasedRNG[575])|((m[768]&m[769]&~m[770]&~m[771]&~m[820])|(m[768]&~m[769]&m[770]&~m[771]&~m[820])|(~m[768]&m[769]&m[770]&~m[771]&~m[820])|(m[768]&m[769]&m[770]&~m[771]&~m[820])|(m[768]&m[769]&m[770]&m[771]&~m[820])|(m[768]&m[769]&~m[770]&~m[771]&m[820])|(m[768]&~m[769]&m[770]&~m[771]&m[820])|(~m[768]&m[769]&m[770]&~m[771]&m[820])|(m[768]&m[769]&m[770]&~m[771]&m[820])|(m[768]&m[769]&m[770]&m[771]&m[820]));
    m[777] = (((m[773]&~m[774]&~m[775]&~m[776]&~m[825])|(~m[773]&m[774]&~m[775]&~m[776]&~m[825])|(~m[773]&~m[774]&m[775]&~m[776]&~m[825])|(m[773]&m[774]&~m[775]&m[776]&~m[825])|(m[773]&~m[774]&m[775]&m[776]&~m[825])|(~m[773]&m[774]&m[775]&m[776]&~m[825]))&BiasedRNG[576])|(((m[773]&~m[774]&~m[775]&~m[776]&m[825])|(~m[773]&m[774]&~m[775]&~m[776]&m[825])|(~m[773]&~m[774]&m[775]&~m[776]&m[825])|(m[773]&m[774]&~m[775]&m[776]&m[825])|(m[773]&~m[774]&m[775]&m[776]&m[825])|(~m[773]&m[774]&m[775]&m[776]&m[825]))&~BiasedRNG[576])|((m[773]&m[774]&~m[775]&~m[776]&~m[825])|(m[773]&~m[774]&m[775]&~m[776]&~m[825])|(~m[773]&m[774]&m[775]&~m[776]&~m[825])|(m[773]&m[774]&m[775]&~m[776]&~m[825])|(m[773]&m[774]&m[775]&m[776]&~m[825])|(m[773]&m[774]&~m[775]&~m[776]&m[825])|(m[773]&~m[774]&m[775]&~m[776]&m[825])|(~m[773]&m[774]&m[775]&~m[776]&m[825])|(m[773]&m[774]&m[775]&~m[776]&m[825])|(m[773]&m[774]&m[775]&m[776]&m[825]));
    m[782] = (((m[778]&~m[779]&~m[780]&~m[781]&~m[830])|(~m[778]&m[779]&~m[780]&~m[781]&~m[830])|(~m[778]&~m[779]&m[780]&~m[781]&~m[830])|(m[778]&m[779]&~m[780]&m[781]&~m[830])|(m[778]&~m[779]&m[780]&m[781]&~m[830])|(~m[778]&m[779]&m[780]&m[781]&~m[830]))&BiasedRNG[577])|(((m[778]&~m[779]&~m[780]&~m[781]&m[830])|(~m[778]&m[779]&~m[780]&~m[781]&m[830])|(~m[778]&~m[779]&m[780]&~m[781]&m[830])|(m[778]&m[779]&~m[780]&m[781]&m[830])|(m[778]&~m[779]&m[780]&m[781]&m[830])|(~m[778]&m[779]&m[780]&m[781]&m[830]))&~BiasedRNG[577])|((m[778]&m[779]&~m[780]&~m[781]&~m[830])|(m[778]&~m[779]&m[780]&~m[781]&~m[830])|(~m[778]&m[779]&m[780]&~m[781]&~m[830])|(m[778]&m[779]&m[780]&~m[781]&~m[830])|(m[778]&m[779]&m[780]&m[781]&~m[830])|(m[778]&m[779]&~m[780]&~m[781]&m[830])|(m[778]&~m[779]&m[780]&~m[781]&m[830])|(~m[778]&m[779]&m[780]&~m[781]&m[830])|(m[778]&m[779]&m[780]&~m[781]&m[830])|(m[778]&m[779]&m[780]&m[781]&m[830]));
    m[787] = (((m[783]&~m[784]&~m[785]&~m[786]&~m[835])|(~m[783]&m[784]&~m[785]&~m[786]&~m[835])|(~m[783]&~m[784]&m[785]&~m[786]&~m[835])|(m[783]&m[784]&~m[785]&m[786]&~m[835])|(m[783]&~m[784]&m[785]&m[786]&~m[835])|(~m[783]&m[784]&m[785]&m[786]&~m[835]))&BiasedRNG[578])|(((m[783]&~m[784]&~m[785]&~m[786]&m[835])|(~m[783]&m[784]&~m[785]&~m[786]&m[835])|(~m[783]&~m[784]&m[785]&~m[786]&m[835])|(m[783]&m[784]&~m[785]&m[786]&m[835])|(m[783]&~m[784]&m[785]&m[786]&m[835])|(~m[783]&m[784]&m[785]&m[786]&m[835]))&~BiasedRNG[578])|((m[783]&m[784]&~m[785]&~m[786]&~m[835])|(m[783]&~m[784]&m[785]&~m[786]&~m[835])|(~m[783]&m[784]&m[785]&~m[786]&~m[835])|(m[783]&m[784]&m[785]&~m[786]&~m[835])|(m[783]&m[784]&m[785]&m[786]&~m[835])|(m[783]&m[784]&~m[785]&~m[786]&m[835])|(m[783]&~m[784]&m[785]&~m[786]&m[835])|(~m[783]&m[784]&m[785]&~m[786]&m[835])|(m[783]&m[784]&m[785]&~m[786]&m[835])|(m[783]&m[784]&m[785]&m[786]&m[835]));
    m[792] = (((m[788]&~m[789]&~m[790]&~m[791]&~m[840])|(~m[788]&m[789]&~m[790]&~m[791]&~m[840])|(~m[788]&~m[789]&m[790]&~m[791]&~m[840])|(m[788]&m[789]&~m[790]&m[791]&~m[840])|(m[788]&~m[789]&m[790]&m[791]&~m[840])|(~m[788]&m[789]&m[790]&m[791]&~m[840]))&BiasedRNG[579])|(((m[788]&~m[789]&~m[790]&~m[791]&m[840])|(~m[788]&m[789]&~m[790]&~m[791]&m[840])|(~m[788]&~m[789]&m[790]&~m[791]&m[840])|(m[788]&m[789]&~m[790]&m[791]&m[840])|(m[788]&~m[789]&m[790]&m[791]&m[840])|(~m[788]&m[789]&m[790]&m[791]&m[840]))&~BiasedRNG[579])|((m[788]&m[789]&~m[790]&~m[791]&~m[840])|(m[788]&~m[789]&m[790]&~m[791]&~m[840])|(~m[788]&m[789]&m[790]&~m[791]&~m[840])|(m[788]&m[789]&m[790]&~m[791]&~m[840])|(m[788]&m[789]&m[790]&m[791]&~m[840])|(m[788]&m[789]&~m[790]&~m[791]&m[840])|(m[788]&~m[789]&m[790]&~m[791]&m[840])|(~m[788]&m[789]&m[790]&~m[791]&m[840])|(m[788]&m[789]&m[790]&~m[791]&m[840])|(m[788]&m[789]&m[790]&m[791]&m[840]));
    m[797] = (((m[793]&~m[794]&~m[795]&~m[796]&~m[845])|(~m[793]&m[794]&~m[795]&~m[796]&~m[845])|(~m[793]&~m[794]&m[795]&~m[796]&~m[845])|(m[793]&m[794]&~m[795]&m[796]&~m[845])|(m[793]&~m[794]&m[795]&m[796]&~m[845])|(~m[793]&m[794]&m[795]&m[796]&~m[845]))&BiasedRNG[580])|(((m[793]&~m[794]&~m[795]&~m[796]&m[845])|(~m[793]&m[794]&~m[795]&~m[796]&m[845])|(~m[793]&~m[794]&m[795]&~m[796]&m[845])|(m[793]&m[794]&~m[795]&m[796]&m[845])|(m[793]&~m[794]&m[795]&m[796]&m[845])|(~m[793]&m[794]&m[795]&m[796]&m[845]))&~BiasedRNG[580])|((m[793]&m[794]&~m[795]&~m[796]&~m[845])|(m[793]&~m[794]&m[795]&~m[796]&~m[845])|(~m[793]&m[794]&m[795]&~m[796]&~m[845])|(m[793]&m[794]&m[795]&~m[796]&~m[845])|(m[793]&m[794]&m[795]&m[796]&~m[845])|(m[793]&m[794]&~m[795]&~m[796]&m[845])|(m[793]&~m[794]&m[795]&~m[796]&m[845])|(~m[793]&m[794]&m[795]&~m[796]&m[845])|(m[793]&m[794]&m[795]&~m[796]&m[845])|(m[793]&m[794]&m[795]&m[796]&m[845]));
    m[802] = (((m[798]&~m[799]&~m[800]&~m[801]&~m[850])|(~m[798]&m[799]&~m[800]&~m[801]&~m[850])|(~m[798]&~m[799]&m[800]&~m[801]&~m[850])|(m[798]&m[799]&~m[800]&m[801]&~m[850])|(m[798]&~m[799]&m[800]&m[801]&~m[850])|(~m[798]&m[799]&m[800]&m[801]&~m[850]))&BiasedRNG[581])|(((m[798]&~m[799]&~m[800]&~m[801]&m[850])|(~m[798]&m[799]&~m[800]&~m[801]&m[850])|(~m[798]&~m[799]&m[800]&~m[801]&m[850])|(m[798]&m[799]&~m[800]&m[801]&m[850])|(m[798]&~m[799]&m[800]&m[801]&m[850])|(~m[798]&m[799]&m[800]&m[801]&m[850]))&~BiasedRNG[581])|((m[798]&m[799]&~m[800]&~m[801]&~m[850])|(m[798]&~m[799]&m[800]&~m[801]&~m[850])|(~m[798]&m[799]&m[800]&~m[801]&~m[850])|(m[798]&m[799]&m[800]&~m[801]&~m[850])|(m[798]&m[799]&m[800]&m[801]&~m[850])|(m[798]&m[799]&~m[800]&~m[801]&m[850])|(m[798]&~m[799]&m[800]&~m[801]&m[850])|(~m[798]&m[799]&m[800]&~m[801]&m[850])|(m[798]&m[799]&m[800]&~m[801]&m[850])|(m[798]&m[799]&m[800]&m[801]&m[850]));
    m[807] = (((m[803]&~m[804]&~m[805]&~m[806]&~m[860])|(~m[803]&m[804]&~m[805]&~m[806]&~m[860])|(~m[803]&~m[804]&m[805]&~m[806]&~m[860])|(m[803]&m[804]&~m[805]&m[806]&~m[860])|(m[803]&~m[804]&m[805]&m[806]&~m[860])|(~m[803]&m[804]&m[805]&m[806]&~m[860]))&BiasedRNG[582])|(((m[803]&~m[804]&~m[805]&~m[806]&m[860])|(~m[803]&m[804]&~m[805]&~m[806]&m[860])|(~m[803]&~m[804]&m[805]&~m[806]&m[860])|(m[803]&m[804]&~m[805]&m[806]&m[860])|(m[803]&~m[804]&m[805]&m[806]&m[860])|(~m[803]&m[804]&m[805]&m[806]&m[860]))&~BiasedRNG[582])|((m[803]&m[804]&~m[805]&~m[806]&~m[860])|(m[803]&~m[804]&m[805]&~m[806]&~m[860])|(~m[803]&m[804]&m[805]&~m[806]&~m[860])|(m[803]&m[804]&m[805]&~m[806]&~m[860])|(m[803]&m[804]&m[805]&m[806]&~m[860])|(m[803]&m[804]&~m[805]&~m[806]&m[860])|(m[803]&~m[804]&m[805]&~m[806]&m[860])|(~m[803]&m[804]&m[805]&~m[806]&m[860])|(m[803]&m[804]&m[805]&~m[806]&m[860])|(m[803]&m[804]&m[805]&m[806]&m[860]));
    m[812] = (((m[808]&~m[809]&~m[810]&~m[811]&~m[865])|(~m[808]&m[809]&~m[810]&~m[811]&~m[865])|(~m[808]&~m[809]&m[810]&~m[811]&~m[865])|(m[808]&m[809]&~m[810]&m[811]&~m[865])|(m[808]&~m[809]&m[810]&m[811]&~m[865])|(~m[808]&m[809]&m[810]&m[811]&~m[865]))&BiasedRNG[583])|(((m[808]&~m[809]&~m[810]&~m[811]&m[865])|(~m[808]&m[809]&~m[810]&~m[811]&m[865])|(~m[808]&~m[809]&m[810]&~m[811]&m[865])|(m[808]&m[809]&~m[810]&m[811]&m[865])|(m[808]&~m[809]&m[810]&m[811]&m[865])|(~m[808]&m[809]&m[810]&m[811]&m[865]))&~BiasedRNG[583])|((m[808]&m[809]&~m[810]&~m[811]&~m[865])|(m[808]&~m[809]&m[810]&~m[811]&~m[865])|(~m[808]&m[809]&m[810]&~m[811]&~m[865])|(m[808]&m[809]&m[810]&~m[811]&~m[865])|(m[808]&m[809]&m[810]&m[811]&~m[865])|(m[808]&m[809]&~m[810]&~m[811]&m[865])|(m[808]&~m[809]&m[810]&~m[811]&m[865])|(~m[808]&m[809]&m[810]&~m[811]&m[865])|(m[808]&m[809]&m[810]&~m[811]&m[865])|(m[808]&m[809]&m[810]&m[811]&m[865]));
    m[817] = (((m[813]&~m[814]&~m[815]&~m[816]&~m[870])|(~m[813]&m[814]&~m[815]&~m[816]&~m[870])|(~m[813]&~m[814]&m[815]&~m[816]&~m[870])|(m[813]&m[814]&~m[815]&m[816]&~m[870])|(m[813]&~m[814]&m[815]&m[816]&~m[870])|(~m[813]&m[814]&m[815]&m[816]&~m[870]))&BiasedRNG[584])|(((m[813]&~m[814]&~m[815]&~m[816]&m[870])|(~m[813]&m[814]&~m[815]&~m[816]&m[870])|(~m[813]&~m[814]&m[815]&~m[816]&m[870])|(m[813]&m[814]&~m[815]&m[816]&m[870])|(m[813]&~m[814]&m[815]&m[816]&m[870])|(~m[813]&m[814]&m[815]&m[816]&m[870]))&~BiasedRNG[584])|((m[813]&m[814]&~m[815]&~m[816]&~m[870])|(m[813]&~m[814]&m[815]&~m[816]&~m[870])|(~m[813]&m[814]&m[815]&~m[816]&~m[870])|(m[813]&m[814]&m[815]&~m[816]&~m[870])|(m[813]&m[814]&m[815]&m[816]&~m[870])|(m[813]&m[814]&~m[815]&~m[816]&m[870])|(m[813]&~m[814]&m[815]&~m[816]&m[870])|(~m[813]&m[814]&m[815]&~m[816]&m[870])|(m[813]&m[814]&m[815]&~m[816]&m[870])|(m[813]&m[814]&m[815]&m[816]&m[870]));
    m[822] = (((m[818]&~m[819]&~m[820]&~m[821]&~m[875])|(~m[818]&m[819]&~m[820]&~m[821]&~m[875])|(~m[818]&~m[819]&m[820]&~m[821]&~m[875])|(m[818]&m[819]&~m[820]&m[821]&~m[875])|(m[818]&~m[819]&m[820]&m[821]&~m[875])|(~m[818]&m[819]&m[820]&m[821]&~m[875]))&BiasedRNG[585])|(((m[818]&~m[819]&~m[820]&~m[821]&m[875])|(~m[818]&m[819]&~m[820]&~m[821]&m[875])|(~m[818]&~m[819]&m[820]&~m[821]&m[875])|(m[818]&m[819]&~m[820]&m[821]&m[875])|(m[818]&~m[819]&m[820]&m[821]&m[875])|(~m[818]&m[819]&m[820]&m[821]&m[875]))&~BiasedRNG[585])|((m[818]&m[819]&~m[820]&~m[821]&~m[875])|(m[818]&~m[819]&m[820]&~m[821]&~m[875])|(~m[818]&m[819]&m[820]&~m[821]&~m[875])|(m[818]&m[819]&m[820]&~m[821]&~m[875])|(m[818]&m[819]&m[820]&m[821]&~m[875])|(m[818]&m[819]&~m[820]&~m[821]&m[875])|(m[818]&~m[819]&m[820]&~m[821]&m[875])|(~m[818]&m[819]&m[820]&~m[821]&m[875])|(m[818]&m[819]&m[820]&~m[821]&m[875])|(m[818]&m[819]&m[820]&m[821]&m[875]));
    m[827] = (((m[823]&~m[824]&~m[825]&~m[826]&~m[880])|(~m[823]&m[824]&~m[825]&~m[826]&~m[880])|(~m[823]&~m[824]&m[825]&~m[826]&~m[880])|(m[823]&m[824]&~m[825]&m[826]&~m[880])|(m[823]&~m[824]&m[825]&m[826]&~m[880])|(~m[823]&m[824]&m[825]&m[826]&~m[880]))&BiasedRNG[586])|(((m[823]&~m[824]&~m[825]&~m[826]&m[880])|(~m[823]&m[824]&~m[825]&~m[826]&m[880])|(~m[823]&~m[824]&m[825]&~m[826]&m[880])|(m[823]&m[824]&~m[825]&m[826]&m[880])|(m[823]&~m[824]&m[825]&m[826]&m[880])|(~m[823]&m[824]&m[825]&m[826]&m[880]))&~BiasedRNG[586])|((m[823]&m[824]&~m[825]&~m[826]&~m[880])|(m[823]&~m[824]&m[825]&~m[826]&~m[880])|(~m[823]&m[824]&m[825]&~m[826]&~m[880])|(m[823]&m[824]&m[825]&~m[826]&~m[880])|(m[823]&m[824]&m[825]&m[826]&~m[880])|(m[823]&m[824]&~m[825]&~m[826]&m[880])|(m[823]&~m[824]&m[825]&~m[826]&m[880])|(~m[823]&m[824]&m[825]&~m[826]&m[880])|(m[823]&m[824]&m[825]&~m[826]&m[880])|(m[823]&m[824]&m[825]&m[826]&m[880]));
    m[832] = (((m[828]&~m[829]&~m[830]&~m[831]&~m[885])|(~m[828]&m[829]&~m[830]&~m[831]&~m[885])|(~m[828]&~m[829]&m[830]&~m[831]&~m[885])|(m[828]&m[829]&~m[830]&m[831]&~m[885])|(m[828]&~m[829]&m[830]&m[831]&~m[885])|(~m[828]&m[829]&m[830]&m[831]&~m[885]))&BiasedRNG[587])|(((m[828]&~m[829]&~m[830]&~m[831]&m[885])|(~m[828]&m[829]&~m[830]&~m[831]&m[885])|(~m[828]&~m[829]&m[830]&~m[831]&m[885])|(m[828]&m[829]&~m[830]&m[831]&m[885])|(m[828]&~m[829]&m[830]&m[831]&m[885])|(~m[828]&m[829]&m[830]&m[831]&m[885]))&~BiasedRNG[587])|((m[828]&m[829]&~m[830]&~m[831]&~m[885])|(m[828]&~m[829]&m[830]&~m[831]&~m[885])|(~m[828]&m[829]&m[830]&~m[831]&~m[885])|(m[828]&m[829]&m[830]&~m[831]&~m[885])|(m[828]&m[829]&m[830]&m[831]&~m[885])|(m[828]&m[829]&~m[830]&~m[831]&m[885])|(m[828]&~m[829]&m[830]&~m[831]&m[885])|(~m[828]&m[829]&m[830]&~m[831]&m[885])|(m[828]&m[829]&m[830]&~m[831]&m[885])|(m[828]&m[829]&m[830]&m[831]&m[885]));
    m[837] = (((m[833]&~m[834]&~m[835]&~m[836]&~m[890])|(~m[833]&m[834]&~m[835]&~m[836]&~m[890])|(~m[833]&~m[834]&m[835]&~m[836]&~m[890])|(m[833]&m[834]&~m[835]&m[836]&~m[890])|(m[833]&~m[834]&m[835]&m[836]&~m[890])|(~m[833]&m[834]&m[835]&m[836]&~m[890]))&BiasedRNG[588])|(((m[833]&~m[834]&~m[835]&~m[836]&m[890])|(~m[833]&m[834]&~m[835]&~m[836]&m[890])|(~m[833]&~m[834]&m[835]&~m[836]&m[890])|(m[833]&m[834]&~m[835]&m[836]&m[890])|(m[833]&~m[834]&m[835]&m[836]&m[890])|(~m[833]&m[834]&m[835]&m[836]&m[890]))&~BiasedRNG[588])|((m[833]&m[834]&~m[835]&~m[836]&~m[890])|(m[833]&~m[834]&m[835]&~m[836]&~m[890])|(~m[833]&m[834]&m[835]&~m[836]&~m[890])|(m[833]&m[834]&m[835]&~m[836]&~m[890])|(m[833]&m[834]&m[835]&m[836]&~m[890])|(m[833]&m[834]&~m[835]&~m[836]&m[890])|(m[833]&~m[834]&m[835]&~m[836]&m[890])|(~m[833]&m[834]&m[835]&~m[836]&m[890])|(m[833]&m[834]&m[835]&~m[836]&m[890])|(m[833]&m[834]&m[835]&m[836]&m[890]));
    m[842] = (((m[838]&~m[839]&~m[840]&~m[841]&~m[895])|(~m[838]&m[839]&~m[840]&~m[841]&~m[895])|(~m[838]&~m[839]&m[840]&~m[841]&~m[895])|(m[838]&m[839]&~m[840]&m[841]&~m[895])|(m[838]&~m[839]&m[840]&m[841]&~m[895])|(~m[838]&m[839]&m[840]&m[841]&~m[895]))&BiasedRNG[589])|(((m[838]&~m[839]&~m[840]&~m[841]&m[895])|(~m[838]&m[839]&~m[840]&~m[841]&m[895])|(~m[838]&~m[839]&m[840]&~m[841]&m[895])|(m[838]&m[839]&~m[840]&m[841]&m[895])|(m[838]&~m[839]&m[840]&m[841]&m[895])|(~m[838]&m[839]&m[840]&m[841]&m[895]))&~BiasedRNG[589])|((m[838]&m[839]&~m[840]&~m[841]&~m[895])|(m[838]&~m[839]&m[840]&~m[841]&~m[895])|(~m[838]&m[839]&m[840]&~m[841]&~m[895])|(m[838]&m[839]&m[840]&~m[841]&~m[895])|(m[838]&m[839]&m[840]&m[841]&~m[895])|(m[838]&m[839]&~m[840]&~m[841]&m[895])|(m[838]&~m[839]&m[840]&~m[841]&m[895])|(~m[838]&m[839]&m[840]&~m[841]&m[895])|(m[838]&m[839]&m[840]&~m[841]&m[895])|(m[838]&m[839]&m[840]&m[841]&m[895]));
    m[847] = (((m[843]&~m[844]&~m[845]&~m[846]&~m[900])|(~m[843]&m[844]&~m[845]&~m[846]&~m[900])|(~m[843]&~m[844]&m[845]&~m[846]&~m[900])|(m[843]&m[844]&~m[845]&m[846]&~m[900])|(m[843]&~m[844]&m[845]&m[846]&~m[900])|(~m[843]&m[844]&m[845]&m[846]&~m[900]))&BiasedRNG[590])|(((m[843]&~m[844]&~m[845]&~m[846]&m[900])|(~m[843]&m[844]&~m[845]&~m[846]&m[900])|(~m[843]&~m[844]&m[845]&~m[846]&m[900])|(m[843]&m[844]&~m[845]&m[846]&m[900])|(m[843]&~m[844]&m[845]&m[846]&m[900])|(~m[843]&m[844]&m[845]&m[846]&m[900]))&~BiasedRNG[590])|((m[843]&m[844]&~m[845]&~m[846]&~m[900])|(m[843]&~m[844]&m[845]&~m[846]&~m[900])|(~m[843]&m[844]&m[845]&~m[846]&~m[900])|(m[843]&m[844]&m[845]&~m[846]&~m[900])|(m[843]&m[844]&m[845]&m[846]&~m[900])|(m[843]&m[844]&~m[845]&~m[846]&m[900])|(m[843]&~m[844]&m[845]&~m[846]&m[900])|(~m[843]&m[844]&m[845]&~m[846]&m[900])|(m[843]&m[844]&m[845]&~m[846]&m[900])|(m[843]&m[844]&m[845]&m[846]&m[900]));
    m[852] = (((m[848]&~m[849]&~m[850]&~m[851]&~m[905])|(~m[848]&m[849]&~m[850]&~m[851]&~m[905])|(~m[848]&~m[849]&m[850]&~m[851]&~m[905])|(m[848]&m[849]&~m[850]&m[851]&~m[905])|(m[848]&~m[849]&m[850]&m[851]&~m[905])|(~m[848]&m[849]&m[850]&m[851]&~m[905]))&BiasedRNG[591])|(((m[848]&~m[849]&~m[850]&~m[851]&m[905])|(~m[848]&m[849]&~m[850]&~m[851]&m[905])|(~m[848]&~m[849]&m[850]&~m[851]&m[905])|(m[848]&m[849]&~m[850]&m[851]&m[905])|(m[848]&~m[849]&m[850]&m[851]&m[905])|(~m[848]&m[849]&m[850]&m[851]&m[905]))&~BiasedRNG[591])|((m[848]&m[849]&~m[850]&~m[851]&~m[905])|(m[848]&~m[849]&m[850]&~m[851]&~m[905])|(~m[848]&m[849]&m[850]&~m[851]&~m[905])|(m[848]&m[849]&m[850]&~m[851]&~m[905])|(m[848]&m[849]&m[850]&m[851]&~m[905])|(m[848]&m[849]&~m[850]&~m[851]&m[905])|(m[848]&~m[849]&m[850]&~m[851]&m[905])|(~m[848]&m[849]&m[850]&~m[851]&m[905])|(m[848]&m[849]&m[850]&~m[851]&m[905])|(m[848]&m[849]&m[850]&m[851]&m[905]));
    m[857] = (((m[853]&~m[854]&~m[855]&~m[856]&~m[910])|(~m[853]&m[854]&~m[855]&~m[856]&~m[910])|(~m[853]&~m[854]&m[855]&~m[856]&~m[910])|(m[853]&m[854]&~m[855]&m[856]&~m[910])|(m[853]&~m[854]&m[855]&m[856]&~m[910])|(~m[853]&m[854]&m[855]&m[856]&~m[910]))&BiasedRNG[592])|(((m[853]&~m[854]&~m[855]&~m[856]&m[910])|(~m[853]&m[854]&~m[855]&~m[856]&m[910])|(~m[853]&~m[854]&m[855]&~m[856]&m[910])|(m[853]&m[854]&~m[855]&m[856]&m[910])|(m[853]&~m[854]&m[855]&m[856]&m[910])|(~m[853]&m[854]&m[855]&m[856]&m[910]))&~BiasedRNG[592])|((m[853]&m[854]&~m[855]&~m[856]&~m[910])|(m[853]&~m[854]&m[855]&~m[856]&~m[910])|(~m[853]&m[854]&m[855]&~m[856]&~m[910])|(m[853]&m[854]&m[855]&~m[856]&~m[910])|(m[853]&m[854]&m[855]&m[856]&~m[910])|(m[853]&m[854]&~m[855]&~m[856]&m[910])|(m[853]&~m[854]&m[855]&~m[856]&m[910])|(~m[853]&m[854]&m[855]&~m[856]&m[910])|(m[853]&m[854]&m[855]&~m[856]&m[910])|(m[853]&m[854]&m[855]&m[856]&m[910]));
    m[862] = (((m[858]&~m[859]&~m[860]&~m[861]&~m[913])|(~m[858]&m[859]&~m[860]&~m[861]&~m[913])|(~m[858]&~m[859]&m[860]&~m[861]&~m[913])|(m[858]&m[859]&~m[860]&m[861]&~m[913])|(m[858]&~m[859]&m[860]&m[861]&~m[913])|(~m[858]&m[859]&m[860]&m[861]&~m[913]))&BiasedRNG[593])|(((m[858]&~m[859]&~m[860]&~m[861]&m[913])|(~m[858]&m[859]&~m[860]&~m[861]&m[913])|(~m[858]&~m[859]&m[860]&~m[861]&m[913])|(m[858]&m[859]&~m[860]&m[861]&m[913])|(m[858]&~m[859]&m[860]&m[861]&m[913])|(~m[858]&m[859]&m[860]&m[861]&m[913]))&~BiasedRNG[593])|((m[858]&m[859]&~m[860]&~m[861]&~m[913])|(m[858]&~m[859]&m[860]&~m[861]&~m[913])|(~m[858]&m[859]&m[860]&~m[861]&~m[913])|(m[858]&m[859]&m[860]&~m[861]&~m[913])|(m[858]&m[859]&m[860]&m[861]&~m[913])|(m[858]&m[859]&~m[860]&~m[861]&m[913])|(m[858]&~m[859]&m[860]&~m[861]&m[913])|(~m[858]&m[859]&m[860]&~m[861]&m[913])|(m[858]&m[859]&m[860]&~m[861]&m[913])|(m[858]&m[859]&m[860]&m[861]&m[913]));
    m[867] = (((m[863]&~m[864]&~m[865]&~m[866]&~m[915])|(~m[863]&m[864]&~m[865]&~m[866]&~m[915])|(~m[863]&~m[864]&m[865]&~m[866]&~m[915])|(m[863]&m[864]&~m[865]&m[866]&~m[915])|(m[863]&~m[864]&m[865]&m[866]&~m[915])|(~m[863]&m[864]&m[865]&m[866]&~m[915]))&BiasedRNG[594])|(((m[863]&~m[864]&~m[865]&~m[866]&m[915])|(~m[863]&m[864]&~m[865]&~m[866]&m[915])|(~m[863]&~m[864]&m[865]&~m[866]&m[915])|(m[863]&m[864]&~m[865]&m[866]&m[915])|(m[863]&~m[864]&m[865]&m[866]&m[915])|(~m[863]&m[864]&m[865]&m[866]&m[915]))&~BiasedRNG[594])|((m[863]&m[864]&~m[865]&~m[866]&~m[915])|(m[863]&~m[864]&m[865]&~m[866]&~m[915])|(~m[863]&m[864]&m[865]&~m[866]&~m[915])|(m[863]&m[864]&m[865]&~m[866]&~m[915])|(m[863]&m[864]&m[865]&m[866]&~m[915])|(m[863]&m[864]&~m[865]&~m[866]&m[915])|(m[863]&~m[864]&m[865]&~m[866]&m[915])|(~m[863]&m[864]&m[865]&~m[866]&m[915])|(m[863]&m[864]&m[865]&~m[866]&m[915])|(m[863]&m[864]&m[865]&m[866]&m[915]));
    m[872] = (((m[868]&~m[869]&~m[870]&~m[871]&~m[920])|(~m[868]&m[869]&~m[870]&~m[871]&~m[920])|(~m[868]&~m[869]&m[870]&~m[871]&~m[920])|(m[868]&m[869]&~m[870]&m[871]&~m[920])|(m[868]&~m[869]&m[870]&m[871]&~m[920])|(~m[868]&m[869]&m[870]&m[871]&~m[920]))&BiasedRNG[595])|(((m[868]&~m[869]&~m[870]&~m[871]&m[920])|(~m[868]&m[869]&~m[870]&~m[871]&m[920])|(~m[868]&~m[869]&m[870]&~m[871]&m[920])|(m[868]&m[869]&~m[870]&m[871]&m[920])|(m[868]&~m[869]&m[870]&m[871]&m[920])|(~m[868]&m[869]&m[870]&m[871]&m[920]))&~BiasedRNG[595])|((m[868]&m[869]&~m[870]&~m[871]&~m[920])|(m[868]&~m[869]&m[870]&~m[871]&~m[920])|(~m[868]&m[869]&m[870]&~m[871]&~m[920])|(m[868]&m[869]&m[870]&~m[871]&~m[920])|(m[868]&m[869]&m[870]&m[871]&~m[920])|(m[868]&m[869]&~m[870]&~m[871]&m[920])|(m[868]&~m[869]&m[870]&~m[871]&m[920])|(~m[868]&m[869]&m[870]&~m[871]&m[920])|(m[868]&m[869]&m[870]&~m[871]&m[920])|(m[868]&m[869]&m[870]&m[871]&m[920]));
    m[877] = (((m[873]&~m[874]&~m[875]&~m[876]&~m[925])|(~m[873]&m[874]&~m[875]&~m[876]&~m[925])|(~m[873]&~m[874]&m[875]&~m[876]&~m[925])|(m[873]&m[874]&~m[875]&m[876]&~m[925])|(m[873]&~m[874]&m[875]&m[876]&~m[925])|(~m[873]&m[874]&m[875]&m[876]&~m[925]))&BiasedRNG[596])|(((m[873]&~m[874]&~m[875]&~m[876]&m[925])|(~m[873]&m[874]&~m[875]&~m[876]&m[925])|(~m[873]&~m[874]&m[875]&~m[876]&m[925])|(m[873]&m[874]&~m[875]&m[876]&m[925])|(m[873]&~m[874]&m[875]&m[876]&m[925])|(~m[873]&m[874]&m[875]&m[876]&m[925]))&~BiasedRNG[596])|((m[873]&m[874]&~m[875]&~m[876]&~m[925])|(m[873]&~m[874]&m[875]&~m[876]&~m[925])|(~m[873]&m[874]&m[875]&~m[876]&~m[925])|(m[873]&m[874]&m[875]&~m[876]&~m[925])|(m[873]&m[874]&m[875]&m[876]&~m[925])|(m[873]&m[874]&~m[875]&~m[876]&m[925])|(m[873]&~m[874]&m[875]&~m[876]&m[925])|(~m[873]&m[874]&m[875]&~m[876]&m[925])|(m[873]&m[874]&m[875]&~m[876]&m[925])|(m[873]&m[874]&m[875]&m[876]&m[925]));
    m[882] = (((m[878]&~m[879]&~m[880]&~m[881]&~m[930])|(~m[878]&m[879]&~m[880]&~m[881]&~m[930])|(~m[878]&~m[879]&m[880]&~m[881]&~m[930])|(m[878]&m[879]&~m[880]&m[881]&~m[930])|(m[878]&~m[879]&m[880]&m[881]&~m[930])|(~m[878]&m[879]&m[880]&m[881]&~m[930]))&BiasedRNG[597])|(((m[878]&~m[879]&~m[880]&~m[881]&m[930])|(~m[878]&m[879]&~m[880]&~m[881]&m[930])|(~m[878]&~m[879]&m[880]&~m[881]&m[930])|(m[878]&m[879]&~m[880]&m[881]&m[930])|(m[878]&~m[879]&m[880]&m[881]&m[930])|(~m[878]&m[879]&m[880]&m[881]&m[930]))&~BiasedRNG[597])|((m[878]&m[879]&~m[880]&~m[881]&~m[930])|(m[878]&~m[879]&m[880]&~m[881]&~m[930])|(~m[878]&m[879]&m[880]&~m[881]&~m[930])|(m[878]&m[879]&m[880]&~m[881]&~m[930])|(m[878]&m[879]&m[880]&m[881]&~m[930])|(m[878]&m[879]&~m[880]&~m[881]&m[930])|(m[878]&~m[879]&m[880]&~m[881]&m[930])|(~m[878]&m[879]&m[880]&~m[881]&m[930])|(m[878]&m[879]&m[880]&~m[881]&m[930])|(m[878]&m[879]&m[880]&m[881]&m[930]));
    m[887] = (((m[883]&~m[884]&~m[885]&~m[886]&~m[935])|(~m[883]&m[884]&~m[885]&~m[886]&~m[935])|(~m[883]&~m[884]&m[885]&~m[886]&~m[935])|(m[883]&m[884]&~m[885]&m[886]&~m[935])|(m[883]&~m[884]&m[885]&m[886]&~m[935])|(~m[883]&m[884]&m[885]&m[886]&~m[935]))&BiasedRNG[598])|(((m[883]&~m[884]&~m[885]&~m[886]&m[935])|(~m[883]&m[884]&~m[885]&~m[886]&m[935])|(~m[883]&~m[884]&m[885]&~m[886]&m[935])|(m[883]&m[884]&~m[885]&m[886]&m[935])|(m[883]&~m[884]&m[885]&m[886]&m[935])|(~m[883]&m[884]&m[885]&m[886]&m[935]))&~BiasedRNG[598])|((m[883]&m[884]&~m[885]&~m[886]&~m[935])|(m[883]&~m[884]&m[885]&~m[886]&~m[935])|(~m[883]&m[884]&m[885]&~m[886]&~m[935])|(m[883]&m[884]&m[885]&~m[886]&~m[935])|(m[883]&m[884]&m[885]&m[886]&~m[935])|(m[883]&m[884]&~m[885]&~m[886]&m[935])|(m[883]&~m[884]&m[885]&~m[886]&m[935])|(~m[883]&m[884]&m[885]&~m[886]&m[935])|(m[883]&m[884]&m[885]&~m[886]&m[935])|(m[883]&m[884]&m[885]&m[886]&m[935]));
    m[892] = (((m[888]&~m[889]&~m[890]&~m[891]&~m[940])|(~m[888]&m[889]&~m[890]&~m[891]&~m[940])|(~m[888]&~m[889]&m[890]&~m[891]&~m[940])|(m[888]&m[889]&~m[890]&m[891]&~m[940])|(m[888]&~m[889]&m[890]&m[891]&~m[940])|(~m[888]&m[889]&m[890]&m[891]&~m[940]))&BiasedRNG[599])|(((m[888]&~m[889]&~m[890]&~m[891]&m[940])|(~m[888]&m[889]&~m[890]&~m[891]&m[940])|(~m[888]&~m[889]&m[890]&~m[891]&m[940])|(m[888]&m[889]&~m[890]&m[891]&m[940])|(m[888]&~m[889]&m[890]&m[891]&m[940])|(~m[888]&m[889]&m[890]&m[891]&m[940]))&~BiasedRNG[599])|((m[888]&m[889]&~m[890]&~m[891]&~m[940])|(m[888]&~m[889]&m[890]&~m[891]&~m[940])|(~m[888]&m[889]&m[890]&~m[891]&~m[940])|(m[888]&m[889]&m[890]&~m[891]&~m[940])|(m[888]&m[889]&m[890]&m[891]&~m[940])|(m[888]&m[889]&~m[890]&~m[891]&m[940])|(m[888]&~m[889]&m[890]&~m[891]&m[940])|(~m[888]&m[889]&m[890]&~m[891]&m[940])|(m[888]&m[889]&m[890]&~m[891]&m[940])|(m[888]&m[889]&m[890]&m[891]&m[940]));
    m[897] = (((m[893]&~m[894]&~m[895]&~m[896]&~m[945])|(~m[893]&m[894]&~m[895]&~m[896]&~m[945])|(~m[893]&~m[894]&m[895]&~m[896]&~m[945])|(m[893]&m[894]&~m[895]&m[896]&~m[945])|(m[893]&~m[894]&m[895]&m[896]&~m[945])|(~m[893]&m[894]&m[895]&m[896]&~m[945]))&BiasedRNG[600])|(((m[893]&~m[894]&~m[895]&~m[896]&m[945])|(~m[893]&m[894]&~m[895]&~m[896]&m[945])|(~m[893]&~m[894]&m[895]&~m[896]&m[945])|(m[893]&m[894]&~m[895]&m[896]&m[945])|(m[893]&~m[894]&m[895]&m[896]&m[945])|(~m[893]&m[894]&m[895]&m[896]&m[945]))&~BiasedRNG[600])|((m[893]&m[894]&~m[895]&~m[896]&~m[945])|(m[893]&~m[894]&m[895]&~m[896]&~m[945])|(~m[893]&m[894]&m[895]&~m[896]&~m[945])|(m[893]&m[894]&m[895]&~m[896]&~m[945])|(m[893]&m[894]&m[895]&m[896]&~m[945])|(m[893]&m[894]&~m[895]&~m[896]&m[945])|(m[893]&~m[894]&m[895]&~m[896]&m[945])|(~m[893]&m[894]&m[895]&~m[896]&m[945])|(m[893]&m[894]&m[895]&~m[896]&m[945])|(m[893]&m[894]&m[895]&m[896]&m[945]));
    m[902] = (((m[898]&~m[899]&~m[900]&~m[901]&~m[950])|(~m[898]&m[899]&~m[900]&~m[901]&~m[950])|(~m[898]&~m[899]&m[900]&~m[901]&~m[950])|(m[898]&m[899]&~m[900]&m[901]&~m[950])|(m[898]&~m[899]&m[900]&m[901]&~m[950])|(~m[898]&m[899]&m[900]&m[901]&~m[950]))&BiasedRNG[601])|(((m[898]&~m[899]&~m[900]&~m[901]&m[950])|(~m[898]&m[899]&~m[900]&~m[901]&m[950])|(~m[898]&~m[899]&m[900]&~m[901]&m[950])|(m[898]&m[899]&~m[900]&m[901]&m[950])|(m[898]&~m[899]&m[900]&m[901]&m[950])|(~m[898]&m[899]&m[900]&m[901]&m[950]))&~BiasedRNG[601])|((m[898]&m[899]&~m[900]&~m[901]&~m[950])|(m[898]&~m[899]&m[900]&~m[901]&~m[950])|(~m[898]&m[899]&m[900]&~m[901]&~m[950])|(m[898]&m[899]&m[900]&~m[901]&~m[950])|(m[898]&m[899]&m[900]&m[901]&~m[950])|(m[898]&m[899]&~m[900]&~m[901]&m[950])|(m[898]&~m[899]&m[900]&~m[901]&m[950])|(~m[898]&m[899]&m[900]&~m[901]&m[950])|(m[898]&m[899]&m[900]&~m[901]&m[950])|(m[898]&m[899]&m[900]&m[901]&m[950]));
    m[907] = (((m[903]&~m[904]&~m[905]&~m[906]&~m[955])|(~m[903]&m[904]&~m[905]&~m[906]&~m[955])|(~m[903]&~m[904]&m[905]&~m[906]&~m[955])|(m[903]&m[904]&~m[905]&m[906]&~m[955])|(m[903]&~m[904]&m[905]&m[906]&~m[955])|(~m[903]&m[904]&m[905]&m[906]&~m[955]))&BiasedRNG[602])|(((m[903]&~m[904]&~m[905]&~m[906]&m[955])|(~m[903]&m[904]&~m[905]&~m[906]&m[955])|(~m[903]&~m[904]&m[905]&~m[906]&m[955])|(m[903]&m[904]&~m[905]&m[906]&m[955])|(m[903]&~m[904]&m[905]&m[906]&m[955])|(~m[903]&m[904]&m[905]&m[906]&m[955]))&~BiasedRNG[602])|((m[903]&m[904]&~m[905]&~m[906]&~m[955])|(m[903]&~m[904]&m[905]&~m[906]&~m[955])|(~m[903]&m[904]&m[905]&~m[906]&~m[955])|(m[903]&m[904]&m[905]&~m[906]&~m[955])|(m[903]&m[904]&m[905]&m[906]&~m[955])|(m[903]&m[904]&~m[905]&~m[906]&m[955])|(m[903]&~m[904]&m[905]&~m[906]&m[955])|(~m[903]&m[904]&m[905]&~m[906]&m[955])|(m[903]&m[904]&m[905]&~m[906]&m[955])|(m[903]&m[904]&m[905]&m[906]&m[955]));
    m[912] = (((m[908]&~m[909]&~m[910]&~m[911]&~m[960])|(~m[908]&m[909]&~m[910]&~m[911]&~m[960])|(~m[908]&~m[909]&m[910]&~m[911]&~m[960])|(m[908]&m[909]&~m[910]&m[911]&~m[960])|(m[908]&~m[909]&m[910]&m[911]&~m[960])|(~m[908]&m[909]&m[910]&m[911]&~m[960]))&BiasedRNG[603])|(((m[908]&~m[909]&~m[910]&~m[911]&m[960])|(~m[908]&m[909]&~m[910]&~m[911]&m[960])|(~m[908]&~m[909]&m[910]&~m[911]&m[960])|(m[908]&m[909]&~m[910]&m[911]&m[960])|(m[908]&~m[909]&m[910]&m[911]&m[960])|(~m[908]&m[909]&m[910]&m[911]&m[960]))&~BiasedRNG[603])|((m[908]&m[909]&~m[910]&~m[911]&~m[960])|(m[908]&~m[909]&m[910]&~m[911]&~m[960])|(~m[908]&m[909]&m[910]&~m[911]&~m[960])|(m[908]&m[909]&m[910]&~m[911]&~m[960])|(m[908]&m[909]&m[910]&m[911]&~m[960])|(m[908]&m[909]&~m[910]&~m[911]&m[960])|(m[908]&~m[909]&m[910]&~m[911]&m[960])|(~m[908]&m[909]&m[910]&~m[911]&m[960])|(m[908]&m[909]&m[910]&~m[911]&m[960])|(m[908]&m[909]&m[910]&m[911]&m[960]));
    m[917] = (((m[913]&~m[914]&~m[915]&~m[916]&~m[963])|(~m[913]&m[914]&~m[915]&~m[916]&~m[963])|(~m[913]&~m[914]&m[915]&~m[916]&~m[963])|(m[913]&m[914]&~m[915]&m[916]&~m[963])|(m[913]&~m[914]&m[915]&m[916]&~m[963])|(~m[913]&m[914]&m[915]&m[916]&~m[963]))&BiasedRNG[604])|(((m[913]&~m[914]&~m[915]&~m[916]&m[963])|(~m[913]&m[914]&~m[915]&~m[916]&m[963])|(~m[913]&~m[914]&m[915]&~m[916]&m[963])|(m[913]&m[914]&~m[915]&m[916]&m[963])|(m[913]&~m[914]&m[915]&m[916]&m[963])|(~m[913]&m[914]&m[915]&m[916]&m[963]))&~BiasedRNG[604])|((m[913]&m[914]&~m[915]&~m[916]&~m[963])|(m[913]&~m[914]&m[915]&~m[916]&~m[963])|(~m[913]&m[914]&m[915]&~m[916]&~m[963])|(m[913]&m[914]&m[915]&~m[916]&~m[963])|(m[913]&m[914]&m[915]&m[916]&~m[963])|(m[913]&m[914]&~m[915]&~m[916]&m[963])|(m[913]&~m[914]&m[915]&~m[916]&m[963])|(~m[913]&m[914]&m[915]&~m[916]&m[963])|(m[913]&m[914]&m[915]&~m[916]&m[963])|(m[913]&m[914]&m[915]&m[916]&m[963]));
    m[922] = (((m[918]&~m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&~m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&~m[920]&m[921]&~m[965])|(m[918]&~m[919]&m[920]&m[921]&~m[965])|(~m[918]&m[919]&m[920]&m[921]&~m[965]))&BiasedRNG[605])|(((m[918]&~m[919]&~m[920]&~m[921]&m[965])|(~m[918]&m[919]&~m[920]&~m[921]&m[965])|(~m[918]&~m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&~m[920]&m[921]&m[965])|(m[918]&~m[919]&m[920]&m[921]&m[965])|(~m[918]&m[919]&m[920]&m[921]&m[965]))&~BiasedRNG[605])|((m[918]&m[919]&~m[920]&~m[921]&~m[965])|(m[918]&~m[919]&m[920]&~m[921]&~m[965])|(~m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&m[921]&~m[965])|(m[918]&m[919]&~m[920]&~m[921]&m[965])|(m[918]&~m[919]&m[920]&~m[921]&m[965])|(~m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&m[921]&m[965]));
    m[927] = (((m[923]&~m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&~m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&~m[925]&m[926]&~m[970])|(m[923]&~m[924]&m[925]&m[926]&~m[970])|(~m[923]&m[924]&m[925]&m[926]&~m[970]))&BiasedRNG[606])|(((m[923]&~m[924]&~m[925]&~m[926]&m[970])|(~m[923]&m[924]&~m[925]&~m[926]&m[970])|(~m[923]&~m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&~m[925]&m[926]&m[970])|(m[923]&~m[924]&m[925]&m[926]&m[970])|(~m[923]&m[924]&m[925]&m[926]&m[970]))&~BiasedRNG[606])|((m[923]&m[924]&~m[925]&~m[926]&~m[970])|(m[923]&~m[924]&m[925]&~m[926]&~m[970])|(~m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&m[926]&~m[970])|(m[923]&m[924]&~m[925]&~m[926]&m[970])|(m[923]&~m[924]&m[925]&~m[926]&m[970])|(~m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&m[926]&m[970]));
    m[932] = (((m[928]&~m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&~m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&~m[930]&m[931]&~m[975])|(m[928]&~m[929]&m[930]&m[931]&~m[975])|(~m[928]&m[929]&m[930]&m[931]&~m[975]))&BiasedRNG[607])|(((m[928]&~m[929]&~m[930]&~m[931]&m[975])|(~m[928]&m[929]&~m[930]&~m[931]&m[975])|(~m[928]&~m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&~m[930]&m[931]&m[975])|(m[928]&~m[929]&m[930]&m[931]&m[975])|(~m[928]&m[929]&m[930]&m[931]&m[975]))&~BiasedRNG[607])|((m[928]&m[929]&~m[930]&~m[931]&~m[975])|(m[928]&~m[929]&m[930]&~m[931]&~m[975])|(~m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&m[931]&~m[975])|(m[928]&m[929]&~m[930]&~m[931]&m[975])|(m[928]&~m[929]&m[930]&~m[931]&m[975])|(~m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&m[931]&m[975]));
    m[937] = (((m[933]&~m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&~m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&~m[935]&m[936]&~m[980])|(m[933]&~m[934]&m[935]&m[936]&~m[980])|(~m[933]&m[934]&m[935]&m[936]&~m[980]))&BiasedRNG[608])|(((m[933]&~m[934]&~m[935]&~m[936]&m[980])|(~m[933]&m[934]&~m[935]&~m[936]&m[980])|(~m[933]&~m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&~m[935]&m[936]&m[980])|(m[933]&~m[934]&m[935]&m[936]&m[980])|(~m[933]&m[934]&m[935]&m[936]&m[980]))&~BiasedRNG[608])|((m[933]&m[934]&~m[935]&~m[936]&~m[980])|(m[933]&~m[934]&m[935]&~m[936]&~m[980])|(~m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&m[936]&~m[980])|(m[933]&m[934]&~m[935]&~m[936]&m[980])|(m[933]&~m[934]&m[935]&~m[936]&m[980])|(~m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&m[936]&m[980]));
    m[942] = (((m[938]&~m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&~m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&~m[940]&m[941]&~m[985])|(m[938]&~m[939]&m[940]&m[941]&~m[985])|(~m[938]&m[939]&m[940]&m[941]&~m[985]))&BiasedRNG[609])|(((m[938]&~m[939]&~m[940]&~m[941]&m[985])|(~m[938]&m[939]&~m[940]&~m[941]&m[985])|(~m[938]&~m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&~m[940]&m[941]&m[985])|(m[938]&~m[939]&m[940]&m[941]&m[985])|(~m[938]&m[939]&m[940]&m[941]&m[985]))&~BiasedRNG[609])|((m[938]&m[939]&~m[940]&~m[941]&~m[985])|(m[938]&~m[939]&m[940]&~m[941]&~m[985])|(~m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&m[941]&~m[985])|(m[938]&m[939]&~m[940]&~m[941]&m[985])|(m[938]&~m[939]&m[940]&~m[941]&m[985])|(~m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&m[941]&m[985]));
    m[947] = (((m[943]&~m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&~m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&~m[945]&m[946]&~m[990])|(m[943]&~m[944]&m[945]&m[946]&~m[990])|(~m[943]&m[944]&m[945]&m[946]&~m[990]))&BiasedRNG[610])|(((m[943]&~m[944]&~m[945]&~m[946]&m[990])|(~m[943]&m[944]&~m[945]&~m[946]&m[990])|(~m[943]&~m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&~m[945]&m[946]&m[990])|(m[943]&~m[944]&m[945]&m[946]&m[990])|(~m[943]&m[944]&m[945]&m[946]&m[990]))&~BiasedRNG[610])|((m[943]&m[944]&~m[945]&~m[946]&~m[990])|(m[943]&~m[944]&m[945]&~m[946]&~m[990])|(~m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&m[946]&~m[990])|(m[943]&m[944]&~m[945]&~m[946]&m[990])|(m[943]&~m[944]&m[945]&~m[946]&m[990])|(~m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&m[946]&m[990]));
    m[952] = (((m[948]&~m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&~m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&~m[950]&m[951]&~m[995])|(m[948]&~m[949]&m[950]&m[951]&~m[995])|(~m[948]&m[949]&m[950]&m[951]&~m[995]))&BiasedRNG[611])|(((m[948]&~m[949]&~m[950]&~m[951]&m[995])|(~m[948]&m[949]&~m[950]&~m[951]&m[995])|(~m[948]&~m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&~m[950]&m[951]&m[995])|(m[948]&~m[949]&m[950]&m[951]&m[995])|(~m[948]&m[949]&m[950]&m[951]&m[995]))&~BiasedRNG[611])|((m[948]&m[949]&~m[950]&~m[951]&~m[995])|(m[948]&~m[949]&m[950]&~m[951]&~m[995])|(~m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&m[951]&~m[995])|(m[948]&m[949]&~m[950]&~m[951]&m[995])|(m[948]&~m[949]&m[950]&~m[951]&m[995])|(~m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&m[951]&m[995]));
    m[957] = (((m[953]&~m[954]&~m[955]&~m[956]&~m[1000])|(~m[953]&m[954]&~m[955]&~m[956]&~m[1000])|(~m[953]&~m[954]&m[955]&~m[956]&~m[1000])|(m[953]&m[954]&~m[955]&m[956]&~m[1000])|(m[953]&~m[954]&m[955]&m[956]&~m[1000])|(~m[953]&m[954]&m[955]&m[956]&~m[1000]))&BiasedRNG[612])|(((m[953]&~m[954]&~m[955]&~m[956]&m[1000])|(~m[953]&m[954]&~m[955]&~m[956]&m[1000])|(~m[953]&~m[954]&m[955]&~m[956]&m[1000])|(m[953]&m[954]&~m[955]&m[956]&m[1000])|(m[953]&~m[954]&m[955]&m[956]&m[1000])|(~m[953]&m[954]&m[955]&m[956]&m[1000]))&~BiasedRNG[612])|((m[953]&m[954]&~m[955]&~m[956]&~m[1000])|(m[953]&~m[954]&m[955]&~m[956]&~m[1000])|(~m[953]&m[954]&m[955]&~m[956]&~m[1000])|(m[953]&m[954]&m[955]&~m[956]&~m[1000])|(m[953]&m[954]&m[955]&m[956]&~m[1000])|(m[953]&m[954]&~m[955]&~m[956]&m[1000])|(m[953]&~m[954]&m[955]&~m[956]&m[1000])|(~m[953]&m[954]&m[955]&~m[956]&m[1000])|(m[953]&m[954]&m[955]&~m[956]&m[1000])|(m[953]&m[954]&m[955]&m[956]&m[1000]));
    m[962] = (((m[958]&~m[959]&~m[960]&~m[961]&~m[1005])|(~m[958]&m[959]&~m[960]&~m[961]&~m[1005])|(~m[958]&~m[959]&m[960]&~m[961]&~m[1005])|(m[958]&m[959]&~m[960]&m[961]&~m[1005])|(m[958]&~m[959]&m[960]&m[961]&~m[1005])|(~m[958]&m[959]&m[960]&m[961]&~m[1005]))&BiasedRNG[613])|(((m[958]&~m[959]&~m[960]&~m[961]&m[1005])|(~m[958]&m[959]&~m[960]&~m[961]&m[1005])|(~m[958]&~m[959]&m[960]&~m[961]&m[1005])|(m[958]&m[959]&~m[960]&m[961]&m[1005])|(m[958]&~m[959]&m[960]&m[961]&m[1005])|(~m[958]&m[959]&m[960]&m[961]&m[1005]))&~BiasedRNG[613])|((m[958]&m[959]&~m[960]&~m[961]&~m[1005])|(m[958]&~m[959]&m[960]&~m[961]&~m[1005])|(~m[958]&m[959]&m[960]&~m[961]&~m[1005])|(m[958]&m[959]&m[960]&~m[961]&~m[1005])|(m[958]&m[959]&m[960]&m[961]&~m[1005])|(m[958]&m[959]&~m[960]&~m[961]&m[1005])|(m[958]&~m[959]&m[960]&~m[961]&m[1005])|(~m[958]&m[959]&m[960]&~m[961]&m[1005])|(m[958]&m[959]&m[960]&~m[961]&m[1005])|(m[958]&m[959]&m[960]&m[961]&m[1005]));
    m[967] = (((m[963]&~m[964]&~m[965]&~m[966]&~m[1008])|(~m[963]&m[964]&~m[965]&~m[966]&~m[1008])|(~m[963]&~m[964]&m[965]&~m[966]&~m[1008])|(m[963]&m[964]&~m[965]&m[966]&~m[1008])|(m[963]&~m[964]&m[965]&m[966]&~m[1008])|(~m[963]&m[964]&m[965]&m[966]&~m[1008]))&BiasedRNG[614])|(((m[963]&~m[964]&~m[965]&~m[966]&m[1008])|(~m[963]&m[964]&~m[965]&~m[966]&m[1008])|(~m[963]&~m[964]&m[965]&~m[966]&m[1008])|(m[963]&m[964]&~m[965]&m[966]&m[1008])|(m[963]&~m[964]&m[965]&m[966]&m[1008])|(~m[963]&m[964]&m[965]&m[966]&m[1008]))&~BiasedRNG[614])|((m[963]&m[964]&~m[965]&~m[966]&~m[1008])|(m[963]&~m[964]&m[965]&~m[966]&~m[1008])|(~m[963]&m[964]&m[965]&~m[966]&~m[1008])|(m[963]&m[964]&m[965]&~m[966]&~m[1008])|(m[963]&m[964]&m[965]&m[966]&~m[1008])|(m[963]&m[964]&~m[965]&~m[966]&m[1008])|(m[963]&~m[964]&m[965]&~m[966]&m[1008])|(~m[963]&m[964]&m[965]&~m[966]&m[1008])|(m[963]&m[964]&m[965]&~m[966]&m[1008])|(m[963]&m[964]&m[965]&m[966]&m[1008]));
    m[972] = (((m[968]&~m[969]&~m[970]&~m[971]&~m[1010])|(~m[968]&m[969]&~m[970]&~m[971]&~m[1010])|(~m[968]&~m[969]&m[970]&~m[971]&~m[1010])|(m[968]&m[969]&~m[970]&m[971]&~m[1010])|(m[968]&~m[969]&m[970]&m[971]&~m[1010])|(~m[968]&m[969]&m[970]&m[971]&~m[1010]))&BiasedRNG[615])|(((m[968]&~m[969]&~m[970]&~m[971]&m[1010])|(~m[968]&m[969]&~m[970]&~m[971]&m[1010])|(~m[968]&~m[969]&m[970]&~m[971]&m[1010])|(m[968]&m[969]&~m[970]&m[971]&m[1010])|(m[968]&~m[969]&m[970]&m[971]&m[1010])|(~m[968]&m[969]&m[970]&m[971]&m[1010]))&~BiasedRNG[615])|((m[968]&m[969]&~m[970]&~m[971]&~m[1010])|(m[968]&~m[969]&m[970]&~m[971]&~m[1010])|(~m[968]&m[969]&m[970]&~m[971]&~m[1010])|(m[968]&m[969]&m[970]&~m[971]&~m[1010])|(m[968]&m[969]&m[970]&m[971]&~m[1010])|(m[968]&m[969]&~m[970]&~m[971]&m[1010])|(m[968]&~m[969]&m[970]&~m[971]&m[1010])|(~m[968]&m[969]&m[970]&~m[971]&m[1010])|(m[968]&m[969]&m[970]&~m[971]&m[1010])|(m[968]&m[969]&m[970]&m[971]&m[1010]));
    m[977] = (((m[973]&~m[974]&~m[975]&~m[976]&~m[1015])|(~m[973]&m[974]&~m[975]&~m[976]&~m[1015])|(~m[973]&~m[974]&m[975]&~m[976]&~m[1015])|(m[973]&m[974]&~m[975]&m[976]&~m[1015])|(m[973]&~m[974]&m[975]&m[976]&~m[1015])|(~m[973]&m[974]&m[975]&m[976]&~m[1015]))&BiasedRNG[616])|(((m[973]&~m[974]&~m[975]&~m[976]&m[1015])|(~m[973]&m[974]&~m[975]&~m[976]&m[1015])|(~m[973]&~m[974]&m[975]&~m[976]&m[1015])|(m[973]&m[974]&~m[975]&m[976]&m[1015])|(m[973]&~m[974]&m[975]&m[976]&m[1015])|(~m[973]&m[974]&m[975]&m[976]&m[1015]))&~BiasedRNG[616])|((m[973]&m[974]&~m[975]&~m[976]&~m[1015])|(m[973]&~m[974]&m[975]&~m[976]&~m[1015])|(~m[973]&m[974]&m[975]&~m[976]&~m[1015])|(m[973]&m[974]&m[975]&~m[976]&~m[1015])|(m[973]&m[974]&m[975]&m[976]&~m[1015])|(m[973]&m[974]&~m[975]&~m[976]&m[1015])|(m[973]&~m[974]&m[975]&~m[976]&m[1015])|(~m[973]&m[974]&m[975]&~m[976]&m[1015])|(m[973]&m[974]&m[975]&~m[976]&m[1015])|(m[973]&m[974]&m[975]&m[976]&m[1015]));
    m[982] = (((m[978]&~m[979]&~m[980]&~m[981]&~m[1020])|(~m[978]&m[979]&~m[980]&~m[981]&~m[1020])|(~m[978]&~m[979]&m[980]&~m[981]&~m[1020])|(m[978]&m[979]&~m[980]&m[981]&~m[1020])|(m[978]&~m[979]&m[980]&m[981]&~m[1020])|(~m[978]&m[979]&m[980]&m[981]&~m[1020]))&BiasedRNG[617])|(((m[978]&~m[979]&~m[980]&~m[981]&m[1020])|(~m[978]&m[979]&~m[980]&~m[981]&m[1020])|(~m[978]&~m[979]&m[980]&~m[981]&m[1020])|(m[978]&m[979]&~m[980]&m[981]&m[1020])|(m[978]&~m[979]&m[980]&m[981]&m[1020])|(~m[978]&m[979]&m[980]&m[981]&m[1020]))&~BiasedRNG[617])|((m[978]&m[979]&~m[980]&~m[981]&~m[1020])|(m[978]&~m[979]&m[980]&~m[981]&~m[1020])|(~m[978]&m[979]&m[980]&~m[981]&~m[1020])|(m[978]&m[979]&m[980]&~m[981]&~m[1020])|(m[978]&m[979]&m[980]&m[981]&~m[1020])|(m[978]&m[979]&~m[980]&~m[981]&m[1020])|(m[978]&~m[979]&m[980]&~m[981]&m[1020])|(~m[978]&m[979]&m[980]&~m[981]&m[1020])|(m[978]&m[979]&m[980]&~m[981]&m[1020])|(m[978]&m[979]&m[980]&m[981]&m[1020]));
    m[987] = (((m[983]&~m[984]&~m[985]&~m[986]&~m[1025])|(~m[983]&m[984]&~m[985]&~m[986]&~m[1025])|(~m[983]&~m[984]&m[985]&~m[986]&~m[1025])|(m[983]&m[984]&~m[985]&m[986]&~m[1025])|(m[983]&~m[984]&m[985]&m[986]&~m[1025])|(~m[983]&m[984]&m[985]&m[986]&~m[1025]))&BiasedRNG[618])|(((m[983]&~m[984]&~m[985]&~m[986]&m[1025])|(~m[983]&m[984]&~m[985]&~m[986]&m[1025])|(~m[983]&~m[984]&m[985]&~m[986]&m[1025])|(m[983]&m[984]&~m[985]&m[986]&m[1025])|(m[983]&~m[984]&m[985]&m[986]&m[1025])|(~m[983]&m[984]&m[985]&m[986]&m[1025]))&~BiasedRNG[618])|((m[983]&m[984]&~m[985]&~m[986]&~m[1025])|(m[983]&~m[984]&m[985]&~m[986]&~m[1025])|(~m[983]&m[984]&m[985]&~m[986]&~m[1025])|(m[983]&m[984]&m[985]&~m[986]&~m[1025])|(m[983]&m[984]&m[985]&m[986]&~m[1025])|(m[983]&m[984]&~m[985]&~m[986]&m[1025])|(m[983]&~m[984]&m[985]&~m[986]&m[1025])|(~m[983]&m[984]&m[985]&~m[986]&m[1025])|(m[983]&m[984]&m[985]&~m[986]&m[1025])|(m[983]&m[984]&m[985]&m[986]&m[1025]));
    m[992] = (((m[988]&~m[989]&~m[990]&~m[991]&~m[1030])|(~m[988]&m[989]&~m[990]&~m[991]&~m[1030])|(~m[988]&~m[989]&m[990]&~m[991]&~m[1030])|(m[988]&m[989]&~m[990]&m[991]&~m[1030])|(m[988]&~m[989]&m[990]&m[991]&~m[1030])|(~m[988]&m[989]&m[990]&m[991]&~m[1030]))&BiasedRNG[619])|(((m[988]&~m[989]&~m[990]&~m[991]&m[1030])|(~m[988]&m[989]&~m[990]&~m[991]&m[1030])|(~m[988]&~m[989]&m[990]&~m[991]&m[1030])|(m[988]&m[989]&~m[990]&m[991]&m[1030])|(m[988]&~m[989]&m[990]&m[991]&m[1030])|(~m[988]&m[989]&m[990]&m[991]&m[1030]))&~BiasedRNG[619])|((m[988]&m[989]&~m[990]&~m[991]&~m[1030])|(m[988]&~m[989]&m[990]&~m[991]&~m[1030])|(~m[988]&m[989]&m[990]&~m[991]&~m[1030])|(m[988]&m[989]&m[990]&~m[991]&~m[1030])|(m[988]&m[989]&m[990]&m[991]&~m[1030])|(m[988]&m[989]&~m[990]&~m[991]&m[1030])|(m[988]&~m[989]&m[990]&~m[991]&m[1030])|(~m[988]&m[989]&m[990]&~m[991]&m[1030])|(m[988]&m[989]&m[990]&~m[991]&m[1030])|(m[988]&m[989]&m[990]&m[991]&m[1030]));
    m[997] = (((m[993]&~m[994]&~m[995]&~m[996]&~m[1035])|(~m[993]&m[994]&~m[995]&~m[996]&~m[1035])|(~m[993]&~m[994]&m[995]&~m[996]&~m[1035])|(m[993]&m[994]&~m[995]&m[996]&~m[1035])|(m[993]&~m[994]&m[995]&m[996]&~m[1035])|(~m[993]&m[994]&m[995]&m[996]&~m[1035]))&BiasedRNG[620])|(((m[993]&~m[994]&~m[995]&~m[996]&m[1035])|(~m[993]&m[994]&~m[995]&~m[996]&m[1035])|(~m[993]&~m[994]&m[995]&~m[996]&m[1035])|(m[993]&m[994]&~m[995]&m[996]&m[1035])|(m[993]&~m[994]&m[995]&m[996]&m[1035])|(~m[993]&m[994]&m[995]&m[996]&m[1035]))&~BiasedRNG[620])|((m[993]&m[994]&~m[995]&~m[996]&~m[1035])|(m[993]&~m[994]&m[995]&~m[996]&~m[1035])|(~m[993]&m[994]&m[995]&~m[996]&~m[1035])|(m[993]&m[994]&m[995]&~m[996]&~m[1035])|(m[993]&m[994]&m[995]&m[996]&~m[1035])|(m[993]&m[994]&~m[995]&~m[996]&m[1035])|(m[993]&~m[994]&m[995]&~m[996]&m[1035])|(~m[993]&m[994]&m[995]&~m[996]&m[1035])|(m[993]&m[994]&m[995]&~m[996]&m[1035])|(m[993]&m[994]&m[995]&m[996]&m[1035]));
    m[1002] = (((m[998]&~m[999]&~m[1000]&~m[1001]&~m[1040])|(~m[998]&m[999]&~m[1000]&~m[1001]&~m[1040])|(~m[998]&~m[999]&m[1000]&~m[1001]&~m[1040])|(m[998]&m[999]&~m[1000]&m[1001]&~m[1040])|(m[998]&~m[999]&m[1000]&m[1001]&~m[1040])|(~m[998]&m[999]&m[1000]&m[1001]&~m[1040]))&BiasedRNG[621])|(((m[998]&~m[999]&~m[1000]&~m[1001]&m[1040])|(~m[998]&m[999]&~m[1000]&~m[1001]&m[1040])|(~m[998]&~m[999]&m[1000]&~m[1001]&m[1040])|(m[998]&m[999]&~m[1000]&m[1001]&m[1040])|(m[998]&~m[999]&m[1000]&m[1001]&m[1040])|(~m[998]&m[999]&m[1000]&m[1001]&m[1040]))&~BiasedRNG[621])|((m[998]&m[999]&~m[1000]&~m[1001]&~m[1040])|(m[998]&~m[999]&m[1000]&~m[1001]&~m[1040])|(~m[998]&m[999]&m[1000]&~m[1001]&~m[1040])|(m[998]&m[999]&m[1000]&~m[1001]&~m[1040])|(m[998]&m[999]&m[1000]&m[1001]&~m[1040])|(m[998]&m[999]&~m[1000]&~m[1001]&m[1040])|(m[998]&~m[999]&m[1000]&~m[1001]&m[1040])|(~m[998]&m[999]&m[1000]&~m[1001]&m[1040])|(m[998]&m[999]&m[1000]&~m[1001]&m[1040])|(m[998]&m[999]&m[1000]&m[1001]&m[1040]));
    m[1007] = (((m[1003]&~m[1004]&~m[1005]&~m[1006]&~m[1045])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1045])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1045])|(m[1003]&m[1004]&~m[1005]&m[1006]&~m[1045])|(m[1003]&~m[1004]&m[1005]&m[1006]&~m[1045])|(~m[1003]&m[1004]&m[1005]&m[1006]&~m[1045]))&BiasedRNG[622])|(((m[1003]&~m[1004]&~m[1005]&~m[1006]&m[1045])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&m[1045])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&m[1045])|(m[1003]&m[1004]&~m[1005]&m[1006]&m[1045])|(m[1003]&~m[1004]&m[1005]&m[1006]&m[1045])|(~m[1003]&m[1004]&m[1005]&m[1006]&m[1045]))&~BiasedRNG[622])|((m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1045])|(m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1045])|(~m[1003]&m[1004]&m[1005]&~m[1006]&~m[1045])|(m[1003]&m[1004]&m[1005]&~m[1006]&~m[1045])|(m[1003]&m[1004]&m[1005]&m[1006]&~m[1045])|(m[1003]&m[1004]&~m[1005]&~m[1006]&m[1045])|(m[1003]&~m[1004]&m[1005]&~m[1006]&m[1045])|(~m[1003]&m[1004]&m[1005]&~m[1006]&m[1045])|(m[1003]&m[1004]&m[1005]&~m[1006]&m[1045])|(m[1003]&m[1004]&m[1005]&m[1006]&m[1045]));
    m[1012] = (((m[1008]&~m[1009]&~m[1010]&~m[1011]&~m[1048])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1048])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1048])|(m[1008]&m[1009]&~m[1010]&m[1011]&~m[1048])|(m[1008]&~m[1009]&m[1010]&m[1011]&~m[1048])|(~m[1008]&m[1009]&m[1010]&m[1011]&~m[1048]))&BiasedRNG[623])|(((m[1008]&~m[1009]&~m[1010]&~m[1011]&m[1048])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&m[1048])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&m[1048])|(m[1008]&m[1009]&~m[1010]&m[1011]&m[1048])|(m[1008]&~m[1009]&m[1010]&m[1011]&m[1048])|(~m[1008]&m[1009]&m[1010]&m[1011]&m[1048]))&~BiasedRNG[623])|((m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1048])|(m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1048])|(~m[1008]&m[1009]&m[1010]&~m[1011]&~m[1048])|(m[1008]&m[1009]&m[1010]&~m[1011]&~m[1048])|(m[1008]&m[1009]&m[1010]&m[1011]&~m[1048])|(m[1008]&m[1009]&~m[1010]&~m[1011]&m[1048])|(m[1008]&~m[1009]&m[1010]&~m[1011]&m[1048])|(~m[1008]&m[1009]&m[1010]&~m[1011]&m[1048])|(m[1008]&m[1009]&m[1010]&~m[1011]&m[1048])|(m[1008]&m[1009]&m[1010]&m[1011]&m[1048]));
    m[1017] = (((m[1013]&~m[1014]&~m[1015]&~m[1016]&~m[1050])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1050])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1050])|(m[1013]&m[1014]&~m[1015]&m[1016]&~m[1050])|(m[1013]&~m[1014]&m[1015]&m[1016]&~m[1050])|(~m[1013]&m[1014]&m[1015]&m[1016]&~m[1050]))&BiasedRNG[624])|(((m[1013]&~m[1014]&~m[1015]&~m[1016]&m[1050])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&m[1050])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&m[1050])|(m[1013]&m[1014]&~m[1015]&m[1016]&m[1050])|(m[1013]&~m[1014]&m[1015]&m[1016]&m[1050])|(~m[1013]&m[1014]&m[1015]&m[1016]&m[1050]))&~BiasedRNG[624])|((m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1050])|(m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1050])|(~m[1013]&m[1014]&m[1015]&~m[1016]&~m[1050])|(m[1013]&m[1014]&m[1015]&~m[1016]&~m[1050])|(m[1013]&m[1014]&m[1015]&m[1016]&~m[1050])|(m[1013]&m[1014]&~m[1015]&~m[1016]&m[1050])|(m[1013]&~m[1014]&m[1015]&~m[1016]&m[1050])|(~m[1013]&m[1014]&m[1015]&~m[1016]&m[1050])|(m[1013]&m[1014]&m[1015]&~m[1016]&m[1050])|(m[1013]&m[1014]&m[1015]&m[1016]&m[1050]));
    m[1022] = (((m[1018]&~m[1019]&~m[1020]&~m[1021]&~m[1055])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1055])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1055])|(m[1018]&m[1019]&~m[1020]&m[1021]&~m[1055])|(m[1018]&~m[1019]&m[1020]&m[1021]&~m[1055])|(~m[1018]&m[1019]&m[1020]&m[1021]&~m[1055]))&BiasedRNG[625])|(((m[1018]&~m[1019]&~m[1020]&~m[1021]&m[1055])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&m[1055])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&m[1055])|(m[1018]&m[1019]&~m[1020]&m[1021]&m[1055])|(m[1018]&~m[1019]&m[1020]&m[1021]&m[1055])|(~m[1018]&m[1019]&m[1020]&m[1021]&m[1055]))&~BiasedRNG[625])|((m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1055])|(m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1055])|(~m[1018]&m[1019]&m[1020]&~m[1021]&~m[1055])|(m[1018]&m[1019]&m[1020]&~m[1021]&~m[1055])|(m[1018]&m[1019]&m[1020]&m[1021]&~m[1055])|(m[1018]&m[1019]&~m[1020]&~m[1021]&m[1055])|(m[1018]&~m[1019]&m[1020]&~m[1021]&m[1055])|(~m[1018]&m[1019]&m[1020]&~m[1021]&m[1055])|(m[1018]&m[1019]&m[1020]&~m[1021]&m[1055])|(m[1018]&m[1019]&m[1020]&m[1021]&m[1055]));
    m[1027] = (((m[1023]&~m[1024]&~m[1025]&~m[1026]&~m[1060])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1060])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1060])|(m[1023]&m[1024]&~m[1025]&m[1026]&~m[1060])|(m[1023]&~m[1024]&m[1025]&m[1026]&~m[1060])|(~m[1023]&m[1024]&m[1025]&m[1026]&~m[1060]))&BiasedRNG[626])|(((m[1023]&~m[1024]&~m[1025]&~m[1026]&m[1060])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&m[1060])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&m[1060])|(m[1023]&m[1024]&~m[1025]&m[1026]&m[1060])|(m[1023]&~m[1024]&m[1025]&m[1026]&m[1060])|(~m[1023]&m[1024]&m[1025]&m[1026]&m[1060]))&~BiasedRNG[626])|((m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1060])|(m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1060])|(~m[1023]&m[1024]&m[1025]&~m[1026]&~m[1060])|(m[1023]&m[1024]&m[1025]&~m[1026]&~m[1060])|(m[1023]&m[1024]&m[1025]&m[1026]&~m[1060])|(m[1023]&m[1024]&~m[1025]&~m[1026]&m[1060])|(m[1023]&~m[1024]&m[1025]&~m[1026]&m[1060])|(~m[1023]&m[1024]&m[1025]&~m[1026]&m[1060])|(m[1023]&m[1024]&m[1025]&~m[1026]&m[1060])|(m[1023]&m[1024]&m[1025]&m[1026]&m[1060]));
    m[1032] = (((m[1028]&~m[1029]&~m[1030]&~m[1031]&~m[1065])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1065])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1065])|(m[1028]&m[1029]&~m[1030]&m[1031]&~m[1065])|(m[1028]&~m[1029]&m[1030]&m[1031]&~m[1065])|(~m[1028]&m[1029]&m[1030]&m[1031]&~m[1065]))&BiasedRNG[627])|(((m[1028]&~m[1029]&~m[1030]&~m[1031]&m[1065])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&m[1065])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&m[1065])|(m[1028]&m[1029]&~m[1030]&m[1031]&m[1065])|(m[1028]&~m[1029]&m[1030]&m[1031]&m[1065])|(~m[1028]&m[1029]&m[1030]&m[1031]&m[1065]))&~BiasedRNG[627])|((m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1065])|(m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1065])|(~m[1028]&m[1029]&m[1030]&~m[1031]&~m[1065])|(m[1028]&m[1029]&m[1030]&~m[1031]&~m[1065])|(m[1028]&m[1029]&m[1030]&m[1031]&~m[1065])|(m[1028]&m[1029]&~m[1030]&~m[1031]&m[1065])|(m[1028]&~m[1029]&m[1030]&~m[1031]&m[1065])|(~m[1028]&m[1029]&m[1030]&~m[1031]&m[1065])|(m[1028]&m[1029]&m[1030]&~m[1031]&m[1065])|(m[1028]&m[1029]&m[1030]&m[1031]&m[1065]));
    m[1037] = (((m[1033]&~m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&~m[1070]))&BiasedRNG[628])|(((m[1033]&~m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&~m[1035]&m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&m[1036]&m[1070]))&~BiasedRNG[628])|((m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&~m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&~m[1070])|(m[1033]&m[1034]&~m[1035]&~m[1036]&m[1070])|(m[1033]&~m[1034]&m[1035]&~m[1036]&m[1070])|(~m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&~m[1036]&m[1070])|(m[1033]&m[1034]&m[1035]&m[1036]&m[1070]));
    m[1042] = (((m[1038]&~m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&~m[1075]))&BiasedRNG[629])|(((m[1038]&~m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&~m[1040]&m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&m[1041]&m[1075]))&~BiasedRNG[629])|((m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&~m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&~m[1075])|(m[1038]&m[1039]&~m[1040]&~m[1041]&m[1075])|(m[1038]&~m[1039]&m[1040]&~m[1041]&m[1075])|(~m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&~m[1041]&m[1075])|(m[1038]&m[1039]&m[1040]&m[1041]&m[1075]));
    m[1047] = (((m[1043]&~m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&~m[1080]))&BiasedRNG[630])|(((m[1043]&~m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&~m[1045]&m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&m[1046]&m[1080]))&~BiasedRNG[630])|((m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&~m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&~m[1080])|(m[1043]&m[1044]&~m[1045]&~m[1046]&m[1080])|(m[1043]&~m[1044]&m[1045]&~m[1046]&m[1080])|(~m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&~m[1046]&m[1080])|(m[1043]&m[1044]&m[1045]&m[1046]&m[1080]));
    m[1052] = (((m[1048]&~m[1049]&~m[1050]&~m[1051]&~m[1083])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1083])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1083])|(m[1048]&m[1049]&~m[1050]&m[1051]&~m[1083])|(m[1048]&~m[1049]&m[1050]&m[1051]&~m[1083])|(~m[1048]&m[1049]&m[1050]&m[1051]&~m[1083]))&BiasedRNG[631])|(((m[1048]&~m[1049]&~m[1050]&~m[1051]&m[1083])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&m[1083])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&m[1083])|(m[1048]&m[1049]&~m[1050]&m[1051]&m[1083])|(m[1048]&~m[1049]&m[1050]&m[1051]&m[1083])|(~m[1048]&m[1049]&m[1050]&m[1051]&m[1083]))&~BiasedRNG[631])|((m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1083])|(m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1083])|(~m[1048]&m[1049]&m[1050]&~m[1051]&~m[1083])|(m[1048]&m[1049]&m[1050]&~m[1051]&~m[1083])|(m[1048]&m[1049]&m[1050]&m[1051]&~m[1083])|(m[1048]&m[1049]&~m[1050]&~m[1051]&m[1083])|(m[1048]&~m[1049]&m[1050]&~m[1051]&m[1083])|(~m[1048]&m[1049]&m[1050]&~m[1051]&m[1083])|(m[1048]&m[1049]&m[1050]&~m[1051]&m[1083])|(m[1048]&m[1049]&m[1050]&m[1051]&m[1083]));
    m[1057] = (((m[1053]&~m[1054]&~m[1055]&~m[1056]&~m[1085])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1085])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1085])|(m[1053]&m[1054]&~m[1055]&m[1056]&~m[1085])|(m[1053]&~m[1054]&m[1055]&m[1056]&~m[1085])|(~m[1053]&m[1054]&m[1055]&m[1056]&~m[1085]))&BiasedRNG[632])|(((m[1053]&~m[1054]&~m[1055]&~m[1056]&m[1085])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&m[1085])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&m[1085])|(m[1053]&m[1054]&~m[1055]&m[1056]&m[1085])|(m[1053]&~m[1054]&m[1055]&m[1056]&m[1085])|(~m[1053]&m[1054]&m[1055]&m[1056]&m[1085]))&~BiasedRNG[632])|((m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1085])|(m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1085])|(~m[1053]&m[1054]&m[1055]&~m[1056]&~m[1085])|(m[1053]&m[1054]&m[1055]&~m[1056]&~m[1085])|(m[1053]&m[1054]&m[1055]&m[1056]&~m[1085])|(m[1053]&m[1054]&~m[1055]&~m[1056]&m[1085])|(m[1053]&~m[1054]&m[1055]&~m[1056]&m[1085])|(~m[1053]&m[1054]&m[1055]&~m[1056]&m[1085])|(m[1053]&m[1054]&m[1055]&~m[1056]&m[1085])|(m[1053]&m[1054]&m[1055]&m[1056]&m[1085]));
    m[1062] = (((m[1058]&~m[1059]&~m[1060]&~m[1061]&~m[1090])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1090])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1090])|(m[1058]&m[1059]&~m[1060]&m[1061]&~m[1090])|(m[1058]&~m[1059]&m[1060]&m[1061]&~m[1090])|(~m[1058]&m[1059]&m[1060]&m[1061]&~m[1090]))&BiasedRNG[633])|(((m[1058]&~m[1059]&~m[1060]&~m[1061]&m[1090])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&m[1090])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&m[1090])|(m[1058]&m[1059]&~m[1060]&m[1061]&m[1090])|(m[1058]&~m[1059]&m[1060]&m[1061]&m[1090])|(~m[1058]&m[1059]&m[1060]&m[1061]&m[1090]))&~BiasedRNG[633])|((m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1090])|(m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1090])|(~m[1058]&m[1059]&m[1060]&~m[1061]&~m[1090])|(m[1058]&m[1059]&m[1060]&~m[1061]&~m[1090])|(m[1058]&m[1059]&m[1060]&m[1061]&~m[1090])|(m[1058]&m[1059]&~m[1060]&~m[1061]&m[1090])|(m[1058]&~m[1059]&m[1060]&~m[1061]&m[1090])|(~m[1058]&m[1059]&m[1060]&~m[1061]&m[1090])|(m[1058]&m[1059]&m[1060]&~m[1061]&m[1090])|(m[1058]&m[1059]&m[1060]&m[1061]&m[1090]));
    m[1067] = (((m[1063]&~m[1064]&~m[1065]&~m[1066]&~m[1095])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1095])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1095])|(m[1063]&m[1064]&~m[1065]&m[1066]&~m[1095])|(m[1063]&~m[1064]&m[1065]&m[1066]&~m[1095])|(~m[1063]&m[1064]&m[1065]&m[1066]&~m[1095]))&BiasedRNG[634])|(((m[1063]&~m[1064]&~m[1065]&~m[1066]&m[1095])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&m[1095])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&m[1095])|(m[1063]&m[1064]&~m[1065]&m[1066]&m[1095])|(m[1063]&~m[1064]&m[1065]&m[1066]&m[1095])|(~m[1063]&m[1064]&m[1065]&m[1066]&m[1095]))&~BiasedRNG[634])|((m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1095])|(m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1095])|(~m[1063]&m[1064]&m[1065]&~m[1066]&~m[1095])|(m[1063]&m[1064]&m[1065]&~m[1066]&~m[1095])|(m[1063]&m[1064]&m[1065]&m[1066]&~m[1095])|(m[1063]&m[1064]&~m[1065]&~m[1066]&m[1095])|(m[1063]&~m[1064]&m[1065]&~m[1066]&m[1095])|(~m[1063]&m[1064]&m[1065]&~m[1066]&m[1095])|(m[1063]&m[1064]&m[1065]&~m[1066]&m[1095])|(m[1063]&m[1064]&m[1065]&m[1066]&m[1095]));
    m[1072] = (((m[1068]&~m[1069]&~m[1070]&~m[1071]&~m[1100])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1100])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1100])|(m[1068]&m[1069]&~m[1070]&m[1071]&~m[1100])|(m[1068]&~m[1069]&m[1070]&m[1071]&~m[1100])|(~m[1068]&m[1069]&m[1070]&m[1071]&~m[1100]))&BiasedRNG[635])|(((m[1068]&~m[1069]&~m[1070]&~m[1071]&m[1100])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&m[1100])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&m[1100])|(m[1068]&m[1069]&~m[1070]&m[1071]&m[1100])|(m[1068]&~m[1069]&m[1070]&m[1071]&m[1100])|(~m[1068]&m[1069]&m[1070]&m[1071]&m[1100]))&~BiasedRNG[635])|((m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1100])|(m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1100])|(~m[1068]&m[1069]&m[1070]&~m[1071]&~m[1100])|(m[1068]&m[1069]&m[1070]&~m[1071]&~m[1100])|(m[1068]&m[1069]&m[1070]&m[1071]&~m[1100])|(m[1068]&m[1069]&~m[1070]&~m[1071]&m[1100])|(m[1068]&~m[1069]&m[1070]&~m[1071]&m[1100])|(~m[1068]&m[1069]&m[1070]&~m[1071]&m[1100])|(m[1068]&m[1069]&m[1070]&~m[1071]&m[1100])|(m[1068]&m[1069]&m[1070]&m[1071]&m[1100]));
    m[1077] = (((m[1073]&~m[1074]&~m[1075]&~m[1076]&~m[1105])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1105])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1105])|(m[1073]&m[1074]&~m[1075]&m[1076]&~m[1105])|(m[1073]&~m[1074]&m[1075]&m[1076]&~m[1105])|(~m[1073]&m[1074]&m[1075]&m[1076]&~m[1105]))&BiasedRNG[636])|(((m[1073]&~m[1074]&~m[1075]&~m[1076]&m[1105])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&m[1105])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&m[1105])|(m[1073]&m[1074]&~m[1075]&m[1076]&m[1105])|(m[1073]&~m[1074]&m[1075]&m[1076]&m[1105])|(~m[1073]&m[1074]&m[1075]&m[1076]&m[1105]))&~BiasedRNG[636])|((m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1105])|(m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1105])|(~m[1073]&m[1074]&m[1075]&~m[1076]&~m[1105])|(m[1073]&m[1074]&m[1075]&~m[1076]&~m[1105])|(m[1073]&m[1074]&m[1075]&m[1076]&~m[1105])|(m[1073]&m[1074]&~m[1075]&~m[1076]&m[1105])|(m[1073]&~m[1074]&m[1075]&~m[1076]&m[1105])|(~m[1073]&m[1074]&m[1075]&~m[1076]&m[1105])|(m[1073]&m[1074]&m[1075]&~m[1076]&m[1105])|(m[1073]&m[1074]&m[1075]&m[1076]&m[1105]));
    m[1082] = (((m[1078]&~m[1079]&~m[1080]&~m[1081]&~m[1110])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1110])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1110])|(m[1078]&m[1079]&~m[1080]&m[1081]&~m[1110])|(m[1078]&~m[1079]&m[1080]&m[1081]&~m[1110])|(~m[1078]&m[1079]&m[1080]&m[1081]&~m[1110]))&BiasedRNG[637])|(((m[1078]&~m[1079]&~m[1080]&~m[1081]&m[1110])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&m[1110])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&m[1110])|(m[1078]&m[1079]&~m[1080]&m[1081]&m[1110])|(m[1078]&~m[1079]&m[1080]&m[1081]&m[1110])|(~m[1078]&m[1079]&m[1080]&m[1081]&m[1110]))&~BiasedRNG[637])|((m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1110])|(m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1110])|(~m[1078]&m[1079]&m[1080]&~m[1081]&~m[1110])|(m[1078]&m[1079]&m[1080]&~m[1081]&~m[1110])|(m[1078]&m[1079]&m[1080]&m[1081]&~m[1110])|(m[1078]&m[1079]&~m[1080]&~m[1081]&m[1110])|(m[1078]&~m[1079]&m[1080]&~m[1081]&m[1110])|(~m[1078]&m[1079]&m[1080]&~m[1081]&m[1110])|(m[1078]&m[1079]&m[1080]&~m[1081]&m[1110])|(m[1078]&m[1079]&m[1080]&m[1081]&m[1110]));
    m[1087] = (((m[1083]&~m[1084]&~m[1085]&~m[1086]&~m[1113])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1113])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1113])|(m[1083]&m[1084]&~m[1085]&m[1086]&~m[1113])|(m[1083]&~m[1084]&m[1085]&m[1086]&~m[1113])|(~m[1083]&m[1084]&m[1085]&m[1086]&~m[1113]))&BiasedRNG[638])|(((m[1083]&~m[1084]&~m[1085]&~m[1086]&m[1113])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&m[1113])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&m[1113])|(m[1083]&m[1084]&~m[1085]&m[1086]&m[1113])|(m[1083]&~m[1084]&m[1085]&m[1086]&m[1113])|(~m[1083]&m[1084]&m[1085]&m[1086]&m[1113]))&~BiasedRNG[638])|((m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1113])|(m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1113])|(~m[1083]&m[1084]&m[1085]&~m[1086]&~m[1113])|(m[1083]&m[1084]&m[1085]&~m[1086]&~m[1113])|(m[1083]&m[1084]&m[1085]&m[1086]&~m[1113])|(m[1083]&m[1084]&~m[1085]&~m[1086]&m[1113])|(m[1083]&~m[1084]&m[1085]&~m[1086]&m[1113])|(~m[1083]&m[1084]&m[1085]&~m[1086]&m[1113])|(m[1083]&m[1084]&m[1085]&~m[1086]&m[1113])|(m[1083]&m[1084]&m[1085]&m[1086]&m[1113]));
    m[1092] = (((m[1088]&~m[1089]&~m[1090]&~m[1091]&~m[1115])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1115])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1115])|(m[1088]&m[1089]&~m[1090]&m[1091]&~m[1115])|(m[1088]&~m[1089]&m[1090]&m[1091]&~m[1115])|(~m[1088]&m[1089]&m[1090]&m[1091]&~m[1115]))&BiasedRNG[639])|(((m[1088]&~m[1089]&~m[1090]&~m[1091]&m[1115])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&m[1115])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&m[1115])|(m[1088]&m[1089]&~m[1090]&m[1091]&m[1115])|(m[1088]&~m[1089]&m[1090]&m[1091]&m[1115])|(~m[1088]&m[1089]&m[1090]&m[1091]&m[1115]))&~BiasedRNG[639])|((m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1115])|(m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1115])|(~m[1088]&m[1089]&m[1090]&~m[1091]&~m[1115])|(m[1088]&m[1089]&m[1090]&~m[1091]&~m[1115])|(m[1088]&m[1089]&m[1090]&m[1091]&~m[1115])|(m[1088]&m[1089]&~m[1090]&~m[1091]&m[1115])|(m[1088]&~m[1089]&m[1090]&~m[1091]&m[1115])|(~m[1088]&m[1089]&m[1090]&~m[1091]&m[1115])|(m[1088]&m[1089]&m[1090]&~m[1091]&m[1115])|(m[1088]&m[1089]&m[1090]&m[1091]&m[1115]));
    m[1097] = (((m[1093]&~m[1094]&~m[1095]&~m[1096]&~m[1120])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1120])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1120])|(m[1093]&m[1094]&~m[1095]&m[1096]&~m[1120])|(m[1093]&~m[1094]&m[1095]&m[1096]&~m[1120])|(~m[1093]&m[1094]&m[1095]&m[1096]&~m[1120]))&BiasedRNG[640])|(((m[1093]&~m[1094]&~m[1095]&~m[1096]&m[1120])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&m[1120])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&m[1120])|(m[1093]&m[1094]&~m[1095]&m[1096]&m[1120])|(m[1093]&~m[1094]&m[1095]&m[1096]&m[1120])|(~m[1093]&m[1094]&m[1095]&m[1096]&m[1120]))&~BiasedRNG[640])|((m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1120])|(m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1120])|(~m[1093]&m[1094]&m[1095]&~m[1096]&~m[1120])|(m[1093]&m[1094]&m[1095]&~m[1096]&~m[1120])|(m[1093]&m[1094]&m[1095]&m[1096]&~m[1120])|(m[1093]&m[1094]&~m[1095]&~m[1096]&m[1120])|(m[1093]&~m[1094]&m[1095]&~m[1096]&m[1120])|(~m[1093]&m[1094]&m[1095]&~m[1096]&m[1120])|(m[1093]&m[1094]&m[1095]&~m[1096]&m[1120])|(m[1093]&m[1094]&m[1095]&m[1096]&m[1120]));
    m[1102] = (((m[1098]&~m[1099]&~m[1100]&~m[1101]&~m[1125])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1125])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1125])|(m[1098]&m[1099]&~m[1100]&m[1101]&~m[1125])|(m[1098]&~m[1099]&m[1100]&m[1101]&~m[1125])|(~m[1098]&m[1099]&m[1100]&m[1101]&~m[1125]))&BiasedRNG[641])|(((m[1098]&~m[1099]&~m[1100]&~m[1101]&m[1125])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&m[1125])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&m[1125])|(m[1098]&m[1099]&~m[1100]&m[1101]&m[1125])|(m[1098]&~m[1099]&m[1100]&m[1101]&m[1125])|(~m[1098]&m[1099]&m[1100]&m[1101]&m[1125]))&~BiasedRNG[641])|((m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1125])|(m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1125])|(~m[1098]&m[1099]&m[1100]&~m[1101]&~m[1125])|(m[1098]&m[1099]&m[1100]&~m[1101]&~m[1125])|(m[1098]&m[1099]&m[1100]&m[1101]&~m[1125])|(m[1098]&m[1099]&~m[1100]&~m[1101]&m[1125])|(m[1098]&~m[1099]&m[1100]&~m[1101]&m[1125])|(~m[1098]&m[1099]&m[1100]&~m[1101]&m[1125])|(m[1098]&m[1099]&m[1100]&~m[1101]&m[1125])|(m[1098]&m[1099]&m[1100]&m[1101]&m[1125]));
    m[1107] = (((m[1103]&~m[1104]&~m[1105]&~m[1106]&~m[1130])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1130])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1130])|(m[1103]&m[1104]&~m[1105]&m[1106]&~m[1130])|(m[1103]&~m[1104]&m[1105]&m[1106]&~m[1130])|(~m[1103]&m[1104]&m[1105]&m[1106]&~m[1130]))&BiasedRNG[642])|(((m[1103]&~m[1104]&~m[1105]&~m[1106]&m[1130])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&m[1130])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&m[1130])|(m[1103]&m[1104]&~m[1105]&m[1106]&m[1130])|(m[1103]&~m[1104]&m[1105]&m[1106]&m[1130])|(~m[1103]&m[1104]&m[1105]&m[1106]&m[1130]))&~BiasedRNG[642])|((m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1130])|(m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1130])|(~m[1103]&m[1104]&m[1105]&~m[1106]&~m[1130])|(m[1103]&m[1104]&m[1105]&~m[1106]&~m[1130])|(m[1103]&m[1104]&m[1105]&m[1106]&~m[1130])|(m[1103]&m[1104]&~m[1105]&~m[1106]&m[1130])|(m[1103]&~m[1104]&m[1105]&~m[1106]&m[1130])|(~m[1103]&m[1104]&m[1105]&~m[1106]&m[1130])|(m[1103]&m[1104]&m[1105]&~m[1106]&m[1130])|(m[1103]&m[1104]&m[1105]&m[1106]&m[1130]));
    m[1112] = (((m[1108]&~m[1109]&~m[1110]&~m[1111]&~m[1135])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1135])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1135])|(m[1108]&m[1109]&~m[1110]&m[1111]&~m[1135])|(m[1108]&~m[1109]&m[1110]&m[1111]&~m[1135])|(~m[1108]&m[1109]&m[1110]&m[1111]&~m[1135]))&BiasedRNG[643])|(((m[1108]&~m[1109]&~m[1110]&~m[1111]&m[1135])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&m[1135])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&m[1135])|(m[1108]&m[1109]&~m[1110]&m[1111]&m[1135])|(m[1108]&~m[1109]&m[1110]&m[1111]&m[1135])|(~m[1108]&m[1109]&m[1110]&m[1111]&m[1135]))&~BiasedRNG[643])|((m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1135])|(m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1135])|(~m[1108]&m[1109]&m[1110]&~m[1111]&~m[1135])|(m[1108]&m[1109]&m[1110]&~m[1111]&~m[1135])|(m[1108]&m[1109]&m[1110]&m[1111]&~m[1135])|(m[1108]&m[1109]&~m[1110]&~m[1111]&m[1135])|(m[1108]&~m[1109]&m[1110]&~m[1111]&m[1135])|(~m[1108]&m[1109]&m[1110]&~m[1111]&m[1135])|(m[1108]&m[1109]&m[1110]&~m[1111]&m[1135])|(m[1108]&m[1109]&m[1110]&m[1111]&m[1135]));
    m[1117] = (((m[1113]&~m[1114]&~m[1115]&~m[1116]&~m[1138])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1138])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1138])|(m[1113]&m[1114]&~m[1115]&m[1116]&~m[1138])|(m[1113]&~m[1114]&m[1115]&m[1116]&~m[1138])|(~m[1113]&m[1114]&m[1115]&m[1116]&~m[1138]))&BiasedRNG[644])|(((m[1113]&~m[1114]&~m[1115]&~m[1116]&m[1138])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&m[1138])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&m[1138])|(m[1113]&m[1114]&~m[1115]&m[1116]&m[1138])|(m[1113]&~m[1114]&m[1115]&m[1116]&m[1138])|(~m[1113]&m[1114]&m[1115]&m[1116]&m[1138]))&~BiasedRNG[644])|((m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1138])|(m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1138])|(~m[1113]&m[1114]&m[1115]&~m[1116]&~m[1138])|(m[1113]&m[1114]&m[1115]&~m[1116]&~m[1138])|(m[1113]&m[1114]&m[1115]&m[1116]&~m[1138])|(m[1113]&m[1114]&~m[1115]&~m[1116]&m[1138])|(m[1113]&~m[1114]&m[1115]&~m[1116]&m[1138])|(~m[1113]&m[1114]&m[1115]&~m[1116]&m[1138])|(m[1113]&m[1114]&m[1115]&~m[1116]&m[1138])|(m[1113]&m[1114]&m[1115]&m[1116]&m[1138]));
    m[1122] = (((m[1118]&~m[1119]&~m[1120]&~m[1121]&~m[1140])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1140])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1140])|(m[1118]&m[1119]&~m[1120]&m[1121]&~m[1140])|(m[1118]&~m[1119]&m[1120]&m[1121]&~m[1140])|(~m[1118]&m[1119]&m[1120]&m[1121]&~m[1140]))&BiasedRNG[645])|(((m[1118]&~m[1119]&~m[1120]&~m[1121]&m[1140])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&m[1140])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&m[1140])|(m[1118]&m[1119]&~m[1120]&m[1121]&m[1140])|(m[1118]&~m[1119]&m[1120]&m[1121]&m[1140])|(~m[1118]&m[1119]&m[1120]&m[1121]&m[1140]))&~BiasedRNG[645])|((m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1140])|(m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1140])|(~m[1118]&m[1119]&m[1120]&~m[1121]&~m[1140])|(m[1118]&m[1119]&m[1120]&~m[1121]&~m[1140])|(m[1118]&m[1119]&m[1120]&m[1121]&~m[1140])|(m[1118]&m[1119]&~m[1120]&~m[1121]&m[1140])|(m[1118]&~m[1119]&m[1120]&~m[1121]&m[1140])|(~m[1118]&m[1119]&m[1120]&~m[1121]&m[1140])|(m[1118]&m[1119]&m[1120]&~m[1121]&m[1140])|(m[1118]&m[1119]&m[1120]&m[1121]&m[1140]));
    m[1127] = (((m[1123]&~m[1124]&~m[1125]&~m[1126]&~m[1145])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1145])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1145])|(m[1123]&m[1124]&~m[1125]&m[1126]&~m[1145])|(m[1123]&~m[1124]&m[1125]&m[1126]&~m[1145])|(~m[1123]&m[1124]&m[1125]&m[1126]&~m[1145]))&BiasedRNG[646])|(((m[1123]&~m[1124]&~m[1125]&~m[1126]&m[1145])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&m[1145])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&m[1145])|(m[1123]&m[1124]&~m[1125]&m[1126]&m[1145])|(m[1123]&~m[1124]&m[1125]&m[1126]&m[1145])|(~m[1123]&m[1124]&m[1125]&m[1126]&m[1145]))&~BiasedRNG[646])|((m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1145])|(m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1145])|(~m[1123]&m[1124]&m[1125]&~m[1126]&~m[1145])|(m[1123]&m[1124]&m[1125]&~m[1126]&~m[1145])|(m[1123]&m[1124]&m[1125]&m[1126]&~m[1145])|(m[1123]&m[1124]&~m[1125]&~m[1126]&m[1145])|(m[1123]&~m[1124]&m[1125]&~m[1126]&m[1145])|(~m[1123]&m[1124]&m[1125]&~m[1126]&m[1145])|(m[1123]&m[1124]&m[1125]&~m[1126]&m[1145])|(m[1123]&m[1124]&m[1125]&m[1126]&m[1145]));
    m[1132] = (((m[1128]&~m[1129]&~m[1130]&~m[1131]&~m[1150])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1150])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1150])|(m[1128]&m[1129]&~m[1130]&m[1131]&~m[1150])|(m[1128]&~m[1129]&m[1130]&m[1131]&~m[1150])|(~m[1128]&m[1129]&m[1130]&m[1131]&~m[1150]))&BiasedRNG[647])|(((m[1128]&~m[1129]&~m[1130]&~m[1131]&m[1150])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&m[1150])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&m[1150])|(m[1128]&m[1129]&~m[1130]&m[1131]&m[1150])|(m[1128]&~m[1129]&m[1130]&m[1131]&m[1150])|(~m[1128]&m[1129]&m[1130]&m[1131]&m[1150]))&~BiasedRNG[647])|((m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1150])|(m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1150])|(~m[1128]&m[1129]&m[1130]&~m[1131]&~m[1150])|(m[1128]&m[1129]&m[1130]&~m[1131]&~m[1150])|(m[1128]&m[1129]&m[1130]&m[1131]&~m[1150])|(m[1128]&m[1129]&~m[1130]&~m[1131]&m[1150])|(m[1128]&~m[1129]&m[1130]&~m[1131]&m[1150])|(~m[1128]&m[1129]&m[1130]&~m[1131]&m[1150])|(m[1128]&m[1129]&m[1130]&~m[1131]&m[1150])|(m[1128]&m[1129]&m[1130]&m[1131]&m[1150]));
    m[1137] = (((m[1133]&~m[1134]&~m[1135]&~m[1136]&~m[1155])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1155])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1155])|(m[1133]&m[1134]&~m[1135]&m[1136]&~m[1155])|(m[1133]&~m[1134]&m[1135]&m[1136]&~m[1155])|(~m[1133]&m[1134]&m[1135]&m[1136]&~m[1155]))&BiasedRNG[648])|(((m[1133]&~m[1134]&~m[1135]&~m[1136]&m[1155])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&m[1155])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&m[1155])|(m[1133]&m[1134]&~m[1135]&m[1136]&m[1155])|(m[1133]&~m[1134]&m[1135]&m[1136]&m[1155])|(~m[1133]&m[1134]&m[1135]&m[1136]&m[1155]))&~BiasedRNG[648])|((m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1155])|(m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1155])|(~m[1133]&m[1134]&m[1135]&~m[1136]&~m[1155])|(m[1133]&m[1134]&m[1135]&~m[1136]&~m[1155])|(m[1133]&m[1134]&m[1135]&m[1136]&~m[1155])|(m[1133]&m[1134]&~m[1135]&~m[1136]&m[1155])|(m[1133]&~m[1134]&m[1135]&~m[1136]&m[1155])|(~m[1133]&m[1134]&m[1135]&~m[1136]&m[1155])|(m[1133]&m[1134]&m[1135]&~m[1136]&m[1155])|(m[1133]&m[1134]&m[1135]&m[1136]&m[1155]));
    m[1142] = (((m[1138]&~m[1139]&~m[1140]&~m[1141]&~m[1158])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1158])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1158])|(m[1138]&m[1139]&~m[1140]&m[1141]&~m[1158])|(m[1138]&~m[1139]&m[1140]&m[1141]&~m[1158])|(~m[1138]&m[1139]&m[1140]&m[1141]&~m[1158]))&BiasedRNG[649])|(((m[1138]&~m[1139]&~m[1140]&~m[1141]&m[1158])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&m[1158])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&m[1158])|(m[1138]&m[1139]&~m[1140]&m[1141]&m[1158])|(m[1138]&~m[1139]&m[1140]&m[1141]&m[1158])|(~m[1138]&m[1139]&m[1140]&m[1141]&m[1158]))&~BiasedRNG[649])|((m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1158])|(m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1158])|(~m[1138]&m[1139]&m[1140]&~m[1141]&~m[1158])|(m[1138]&m[1139]&m[1140]&~m[1141]&~m[1158])|(m[1138]&m[1139]&m[1140]&m[1141]&~m[1158])|(m[1138]&m[1139]&~m[1140]&~m[1141]&m[1158])|(m[1138]&~m[1139]&m[1140]&~m[1141]&m[1158])|(~m[1138]&m[1139]&m[1140]&~m[1141]&m[1158])|(m[1138]&m[1139]&m[1140]&~m[1141]&m[1158])|(m[1138]&m[1139]&m[1140]&m[1141]&m[1158]));
    m[1147] = (((m[1143]&~m[1144]&~m[1145]&~m[1146]&~m[1160])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1160])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1160])|(m[1143]&m[1144]&~m[1145]&m[1146]&~m[1160])|(m[1143]&~m[1144]&m[1145]&m[1146]&~m[1160])|(~m[1143]&m[1144]&m[1145]&m[1146]&~m[1160]))&BiasedRNG[650])|(((m[1143]&~m[1144]&~m[1145]&~m[1146]&m[1160])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&m[1160])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&m[1160])|(m[1143]&m[1144]&~m[1145]&m[1146]&m[1160])|(m[1143]&~m[1144]&m[1145]&m[1146]&m[1160])|(~m[1143]&m[1144]&m[1145]&m[1146]&m[1160]))&~BiasedRNG[650])|((m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1160])|(m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1160])|(~m[1143]&m[1144]&m[1145]&~m[1146]&~m[1160])|(m[1143]&m[1144]&m[1145]&~m[1146]&~m[1160])|(m[1143]&m[1144]&m[1145]&m[1146]&~m[1160])|(m[1143]&m[1144]&~m[1145]&~m[1146]&m[1160])|(m[1143]&~m[1144]&m[1145]&~m[1146]&m[1160])|(~m[1143]&m[1144]&m[1145]&~m[1146]&m[1160])|(m[1143]&m[1144]&m[1145]&~m[1146]&m[1160])|(m[1143]&m[1144]&m[1145]&m[1146]&m[1160]));
    m[1152] = (((m[1148]&~m[1149]&~m[1150]&~m[1151]&~m[1165])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1165])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1165])|(m[1148]&m[1149]&~m[1150]&m[1151]&~m[1165])|(m[1148]&~m[1149]&m[1150]&m[1151]&~m[1165])|(~m[1148]&m[1149]&m[1150]&m[1151]&~m[1165]))&BiasedRNG[651])|(((m[1148]&~m[1149]&~m[1150]&~m[1151]&m[1165])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&m[1165])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&m[1165])|(m[1148]&m[1149]&~m[1150]&m[1151]&m[1165])|(m[1148]&~m[1149]&m[1150]&m[1151]&m[1165])|(~m[1148]&m[1149]&m[1150]&m[1151]&m[1165]))&~BiasedRNG[651])|((m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1165])|(m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1165])|(~m[1148]&m[1149]&m[1150]&~m[1151]&~m[1165])|(m[1148]&m[1149]&m[1150]&~m[1151]&~m[1165])|(m[1148]&m[1149]&m[1150]&m[1151]&~m[1165])|(m[1148]&m[1149]&~m[1150]&~m[1151]&m[1165])|(m[1148]&~m[1149]&m[1150]&~m[1151]&m[1165])|(~m[1148]&m[1149]&m[1150]&~m[1151]&m[1165])|(m[1148]&m[1149]&m[1150]&~m[1151]&m[1165])|(m[1148]&m[1149]&m[1150]&m[1151]&m[1165]));
    m[1157] = (((m[1153]&~m[1154]&~m[1155]&~m[1156]&~m[1170])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1170])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1170])|(m[1153]&m[1154]&~m[1155]&m[1156]&~m[1170])|(m[1153]&~m[1154]&m[1155]&m[1156]&~m[1170])|(~m[1153]&m[1154]&m[1155]&m[1156]&~m[1170]))&BiasedRNG[652])|(((m[1153]&~m[1154]&~m[1155]&~m[1156]&m[1170])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&m[1170])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&m[1170])|(m[1153]&m[1154]&~m[1155]&m[1156]&m[1170])|(m[1153]&~m[1154]&m[1155]&m[1156]&m[1170])|(~m[1153]&m[1154]&m[1155]&m[1156]&m[1170]))&~BiasedRNG[652])|((m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1170])|(m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1170])|(~m[1153]&m[1154]&m[1155]&~m[1156]&~m[1170])|(m[1153]&m[1154]&m[1155]&~m[1156]&~m[1170])|(m[1153]&m[1154]&m[1155]&m[1156]&~m[1170])|(m[1153]&m[1154]&~m[1155]&~m[1156]&m[1170])|(m[1153]&~m[1154]&m[1155]&~m[1156]&m[1170])|(~m[1153]&m[1154]&m[1155]&~m[1156]&m[1170])|(m[1153]&m[1154]&m[1155]&~m[1156]&m[1170])|(m[1153]&m[1154]&m[1155]&m[1156]&m[1170]));
    m[1162] = (((m[1158]&~m[1159]&~m[1160]&~m[1161]&~m[1173])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1173])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1173])|(m[1158]&m[1159]&~m[1160]&m[1161]&~m[1173])|(m[1158]&~m[1159]&m[1160]&m[1161]&~m[1173])|(~m[1158]&m[1159]&m[1160]&m[1161]&~m[1173]))&BiasedRNG[653])|(((m[1158]&~m[1159]&~m[1160]&~m[1161]&m[1173])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&m[1173])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&m[1173])|(m[1158]&m[1159]&~m[1160]&m[1161]&m[1173])|(m[1158]&~m[1159]&m[1160]&m[1161]&m[1173])|(~m[1158]&m[1159]&m[1160]&m[1161]&m[1173]))&~BiasedRNG[653])|((m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1173])|(m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1173])|(~m[1158]&m[1159]&m[1160]&~m[1161]&~m[1173])|(m[1158]&m[1159]&m[1160]&~m[1161]&~m[1173])|(m[1158]&m[1159]&m[1160]&m[1161]&~m[1173])|(m[1158]&m[1159]&~m[1160]&~m[1161]&m[1173])|(m[1158]&~m[1159]&m[1160]&~m[1161]&m[1173])|(~m[1158]&m[1159]&m[1160]&~m[1161]&m[1173])|(m[1158]&m[1159]&m[1160]&~m[1161]&m[1173])|(m[1158]&m[1159]&m[1160]&m[1161]&m[1173]));
    m[1167] = (((m[1163]&~m[1164]&~m[1165]&~m[1166]&~m[1175])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1175])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1175])|(m[1163]&m[1164]&~m[1165]&m[1166]&~m[1175])|(m[1163]&~m[1164]&m[1165]&m[1166]&~m[1175])|(~m[1163]&m[1164]&m[1165]&m[1166]&~m[1175]))&BiasedRNG[654])|(((m[1163]&~m[1164]&~m[1165]&~m[1166]&m[1175])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&m[1175])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&m[1175])|(m[1163]&m[1164]&~m[1165]&m[1166]&m[1175])|(m[1163]&~m[1164]&m[1165]&m[1166]&m[1175])|(~m[1163]&m[1164]&m[1165]&m[1166]&m[1175]))&~BiasedRNG[654])|((m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1175])|(m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1175])|(~m[1163]&m[1164]&m[1165]&~m[1166]&~m[1175])|(m[1163]&m[1164]&m[1165]&~m[1166]&~m[1175])|(m[1163]&m[1164]&m[1165]&m[1166]&~m[1175])|(m[1163]&m[1164]&~m[1165]&~m[1166]&m[1175])|(m[1163]&~m[1164]&m[1165]&~m[1166]&m[1175])|(~m[1163]&m[1164]&m[1165]&~m[1166]&m[1175])|(m[1163]&m[1164]&m[1165]&~m[1166]&m[1175])|(m[1163]&m[1164]&m[1165]&m[1166]&m[1175]));
    m[1172] = (((m[1168]&~m[1169]&~m[1170]&~m[1171]&~m[1180])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1180])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1180])|(m[1168]&m[1169]&~m[1170]&m[1171]&~m[1180])|(m[1168]&~m[1169]&m[1170]&m[1171]&~m[1180])|(~m[1168]&m[1169]&m[1170]&m[1171]&~m[1180]))&BiasedRNG[655])|(((m[1168]&~m[1169]&~m[1170]&~m[1171]&m[1180])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&m[1180])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&m[1180])|(m[1168]&m[1169]&~m[1170]&m[1171]&m[1180])|(m[1168]&~m[1169]&m[1170]&m[1171]&m[1180])|(~m[1168]&m[1169]&m[1170]&m[1171]&m[1180]))&~BiasedRNG[655])|((m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1180])|(m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1180])|(~m[1168]&m[1169]&m[1170]&~m[1171]&~m[1180])|(m[1168]&m[1169]&m[1170]&~m[1171]&~m[1180])|(m[1168]&m[1169]&m[1170]&m[1171]&~m[1180])|(m[1168]&m[1169]&~m[1170]&~m[1171]&m[1180])|(m[1168]&~m[1169]&m[1170]&~m[1171]&m[1180])|(~m[1168]&m[1169]&m[1170]&~m[1171]&m[1180])|(m[1168]&m[1169]&m[1170]&~m[1171]&m[1180])|(m[1168]&m[1169]&m[1170]&m[1171]&m[1180]));
    m[1177] = (((m[1173]&~m[1174]&~m[1175]&~m[1176]&~m[1183])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1183])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1183])|(m[1173]&m[1174]&~m[1175]&m[1176]&~m[1183])|(m[1173]&~m[1174]&m[1175]&m[1176]&~m[1183])|(~m[1173]&m[1174]&m[1175]&m[1176]&~m[1183]))&BiasedRNG[656])|(((m[1173]&~m[1174]&~m[1175]&~m[1176]&m[1183])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&m[1183])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&m[1183])|(m[1173]&m[1174]&~m[1175]&m[1176]&m[1183])|(m[1173]&~m[1174]&m[1175]&m[1176]&m[1183])|(~m[1173]&m[1174]&m[1175]&m[1176]&m[1183]))&~BiasedRNG[656])|((m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1183])|(m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1183])|(~m[1173]&m[1174]&m[1175]&~m[1176]&~m[1183])|(m[1173]&m[1174]&m[1175]&~m[1176]&~m[1183])|(m[1173]&m[1174]&m[1175]&m[1176]&~m[1183])|(m[1173]&m[1174]&~m[1175]&~m[1176]&m[1183])|(m[1173]&~m[1174]&m[1175]&~m[1176]&m[1183])|(~m[1173]&m[1174]&m[1175]&~m[1176]&m[1183])|(m[1173]&m[1174]&m[1175]&~m[1176]&m[1183])|(m[1173]&m[1174]&m[1175]&m[1176]&m[1183]));
    m[1182] = (((m[1178]&~m[1179]&~m[1180]&~m[1181]&~m[1185])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1185])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1185])|(m[1178]&m[1179]&~m[1180]&m[1181]&~m[1185])|(m[1178]&~m[1179]&m[1180]&m[1181]&~m[1185])|(~m[1178]&m[1179]&m[1180]&m[1181]&~m[1185]))&BiasedRNG[657])|(((m[1178]&~m[1179]&~m[1180]&~m[1181]&m[1185])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&m[1185])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&m[1185])|(m[1178]&m[1179]&~m[1180]&m[1181]&m[1185])|(m[1178]&~m[1179]&m[1180]&m[1181]&m[1185])|(~m[1178]&m[1179]&m[1180]&m[1181]&m[1185]))&~BiasedRNG[657])|((m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1185])|(m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1185])|(~m[1178]&m[1179]&m[1180]&~m[1181]&~m[1185])|(m[1178]&m[1179]&m[1180]&~m[1181]&~m[1185])|(m[1178]&m[1179]&m[1180]&m[1181]&~m[1185])|(m[1178]&m[1179]&~m[1180]&~m[1181]&m[1185])|(m[1178]&~m[1179]&m[1180]&~m[1181]&m[1185])|(~m[1178]&m[1179]&m[1180]&~m[1181]&m[1185])|(m[1178]&m[1179]&m[1180]&~m[1181]&m[1185])|(m[1178]&m[1179]&m[1180]&m[1181]&m[1185]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[717]&LFSRcolor0[445]&LFSRcolor0[579]&LFSRcolor0[731]);
    BiasedRNG[1] = (LFSRcolor0[656]&LFSRcolor0[265]&LFSRcolor0[594]&LFSRcolor0[349]);
    BiasedRNG[2] = (LFSRcolor0[308]&LFSRcolor0[325]&LFSRcolor0[678]&LFSRcolor0[214]);
    BiasedRNG[3] = (LFSRcolor0[12]&LFSRcolor0[373]&LFSRcolor0[718]&LFSRcolor0[45]);
    BiasedRNG[4] = (LFSRcolor0[140]&LFSRcolor0[564]&LFSRcolor0[498]&LFSRcolor0[813]);
    BiasedRNG[5] = (LFSRcolor0[281]&LFSRcolor0[478]&LFSRcolor0[183]&LFSRcolor0[379]);
    BiasedRNG[6] = (LFSRcolor0[198]&LFSRcolor0[290]&LFSRcolor0[738]&LFSRcolor0[82]);
    BiasedRNG[7] = (LFSRcolor0[416]&LFSRcolor0[737]&LFSRcolor0[417]&LFSRcolor0[289]);
    BiasedRNG[8] = (LFSRcolor0[115]&LFSRcolor0[427]&LFSRcolor0[704]&LFSRcolor0[272]);
    BiasedRNG[9] = (LFSRcolor0[617]&LFSRcolor0[152]&LFSRcolor0[602]&LFSRcolor0[740]);
    BiasedRNG[10] = (LFSRcolor0[228]&LFSRcolor0[173]&LFSRcolor0[295]&LFSRcolor0[565]);
    BiasedRNG[11] = (LFSRcolor0[673]&LFSRcolor0[22]&LFSRcolor0[283]&LFSRcolor0[707]);
    BiasedRNG[12] = (LFSRcolor0[613]&LFSRcolor0[596]&LFSRcolor0[4]&LFSRcolor0[772]);
    BiasedRNG[13] = (LFSRcolor0[441]&LFSRcolor0[48]&LFSRcolor0[165]&LFSRcolor0[159]);
    BiasedRNG[14] = (LFSRcolor0[79]&LFSRcolor0[729]&LFSRcolor0[382]&LFSRcolor0[149]);
    BiasedRNG[15] = (LFSRcolor0[284]&LFSRcolor0[476]&LFSRcolor0[288]&LFSRcolor0[8]);
    BiasedRNG[16] = (LFSRcolor0[491]&LFSRcolor0[642]&LFSRcolor0[218]&LFSRcolor0[741]);
    BiasedRNG[17] = (LFSRcolor0[213]&LFSRcolor0[57]&LFSRcolor0[628]&LFSRcolor0[697]);
    BiasedRNG[18] = (LFSRcolor0[589]&LFSRcolor0[392]&LFSRcolor0[111]&LFSRcolor0[812]);
    BiasedRNG[19] = (LFSRcolor0[473]&LFSRcolor0[107]&LFSRcolor0[610]&LFSRcolor0[7]);
    BiasedRNG[20] = (LFSRcolor0[612]&LFSRcolor0[541]&LFSRcolor0[771]&LFSRcolor0[181]);
    BiasedRNG[21] = (LFSRcolor0[355]&LFSRcolor0[654]&LFSRcolor0[224]&LFSRcolor0[160]);
    BiasedRNG[22] = (LFSRcolor0[62]&LFSRcolor0[102]&LFSRcolor0[703]&LFSRcolor0[301]);
    BiasedRNG[23] = (LFSRcolor0[2]&LFSRcolor0[465]&LFSRcolor0[637]&LFSRcolor0[547]);
    BiasedRNG[24] = (LFSRcolor0[614]&LFSRcolor0[650]&LFSRcolor0[609]&LFSRcolor0[815]);
    BiasedRNG[25] = (LFSRcolor0[517]&LFSRcolor0[626]&LFSRcolor0[627]&LFSRcolor0[639]);
    BiasedRNG[26] = (LFSRcolor0[229]&LFSRcolor0[53]&LFSRcolor0[116]&LFSRcolor0[568]);
    BiasedRNG[27] = (LFSRcolor0[636]&LFSRcolor0[180]&LFSRcolor0[665]&LFSRcolor0[35]);
    BiasedRNG[28] = (LFSRcolor0[543]&LFSRcolor0[775]&LFSRcolor0[822]&LFSRcolor0[825]);
    BiasedRNG[29] = (LFSRcolor0[254]&LFSRcolor0[350]&LFSRcolor0[384]&LFSRcolor0[693]);
    BiasedRNG[30] = (LFSRcolor0[477]&LFSRcolor0[511]&LFSRcolor0[506]&LFSRcolor0[16]);
    BiasedRNG[31] = (LFSRcolor0[555]&LFSRcolor0[575]&LFSRcolor0[279]&LFSRcolor0[250]);
    BiasedRNG[32] = (LFSRcolor0[578]&LFSRcolor0[385]&LFSRcolor0[37]&LFSRcolor0[209]);
    BiasedRNG[33] = (LFSRcolor0[194]&LFSRcolor0[127]&LFSRcolor0[546]&LFSRcolor0[178]);
    BiasedRNG[34] = (LFSRcolor0[234]&LFSRcolor0[54]&LFSRcolor0[788]&LFSRcolor0[606]);
    BiasedRNG[35] = (LFSRcolor0[719]&LFSRcolor0[155]&LFSRcolor0[527]&LFSRcolor0[138]);
    BiasedRNG[36] = (LFSRcolor0[273]&LFSRcolor0[27]&LFSRcolor0[197]&LFSRcolor0[317]);
    BiasedRNG[37] = (LFSRcolor0[646]&LFSRcolor0[466]&LFSRcolor0[507]&LFSRcolor0[817]);
    BiasedRNG[38] = (LFSRcolor0[368]&LFSRcolor0[657]&LFSRcolor0[302]&LFSRcolor0[455]);
    BiasedRNG[39] = (LFSRcolor0[109]&LFSRcolor0[691]&LFSRcolor0[294]&LFSRcolor0[563]);
    BiasedRNG[40] = (LFSRcolor0[200]&LFSRcolor0[19]&LFSRcolor0[514]&LFSRcolor0[413]);
    BiasedRNG[41] = (LFSRcolor0[408]&LFSRcolor0[595]&LFSRcolor0[526]&LFSRcolor0[409]);
    BiasedRNG[42] = (LFSRcolor0[130]&LFSRcolor0[715]&LFSRcolor0[461]&LFSRcolor0[632]);
    BiasedRNG[43] = (LFSRcolor0[81]&LFSRcolor0[341]&LFSRcolor0[488]&LFSRcolor0[63]);
    BiasedRNG[44] = (LFSRcolor0[649]&LFSRcolor0[347]&LFSRcolor0[403]&LFSRcolor0[597]);
    BiasedRNG[45] = (LFSRcolor0[390]&LFSRcolor0[275]&LFSRcolor0[810]&LFSRcolor0[635]);
    BiasedRNG[46] = (LFSRcolor0[332]&LFSRcolor0[93]&LFSRcolor0[169]&LFSRcolor0[502]);
    BiasedRNG[47] = (LFSRcolor0[803]&LFSRcolor0[58]&LFSRcolor0[588]&LFSRcolor0[97]);
    BiasedRNG[48] = (LFSRcolor0[467]&LFSRcolor0[201]&LFSRcolor0[3]&LFSRcolor0[365]);
    BiasedRNG[49] = (LFSRcolor0[779]&LFSRcolor0[651]&LFSRcolor0[443]&LFSRcolor0[510]);
    BiasedRNG[50] = (LFSRcolor0[136]&LFSRcolor0[792]&LFSRcolor0[106]&LFSRcolor0[687]);
    BiasedRNG[51] = (LFSRcolor0[126]&LFSRcolor0[730]&LFSRcolor0[560]&LFSRcolor0[383]);
    BiasedRNG[52] = (LFSRcolor0[141]&LFSRcolor0[363]&LFSRcolor0[278]&LFSRcolor0[780]);
    BiasedRNG[53] = (LFSRcolor0[168]&LFSRcolor0[464]&LFSRcolor0[804]&LFSRcolor0[211]);
    BiasedRNG[54] = (LFSRcolor0[501]&LFSRcolor0[745]&LFSRcolor0[348]&LFSRcolor0[118]);
    BiasedRNG[55] = (LFSRcolor0[240]&LFSRcolor0[611]&LFSRcolor0[816]&LFSRcolor0[196]);
    BiasedRNG[56] = (LFSRcolor0[333]&LFSRcolor0[519]&LFSRcolor0[330]&LFSRcolor0[397]);
    BiasedRNG[57] = (LFSRcolor0[262]&LFSRcolor0[454]&LFSRcolor0[346]&LFSRcolor0[667]);
    BiasedRNG[58] = (LFSRcolor0[40]&LFSRcolor0[216]&LFSRcolor0[619]&LFSRcolor0[672]);
    BiasedRNG[59] = (LFSRcolor0[695]&LFSRcolor0[468]&LFSRcolor0[68]&LFSRcolor0[700]);
    BiasedRNG[60] = (LFSRcolor0[344]&LFSRcolor0[791]&LFSRcolor0[758]&LFSRcolor0[753]);
    BiasedRNG[61] = (LFSRcolor0[566]&LFSRcolor0[584]&LFSRcolor0[376]&LFSRcolor0[472]);
    BiasedRNG[62] = (LFSRcolor0[545]&LFSRcolor0[266]&LFSRcolor0[6]&LFSRcolor0[193]);
    BiasedRNG[63] = (LFSRcolor0[182]&LFSRcolor0[324]&LFSRcolor0[735]&LFSRcolor0[720]);
    BiasedRNG[64] = (LFSRcolor0[648]&LFSRcolor0[76]&LFSRcolor0[342]&LFSRcolor0[61]);
    BiasedRNG[65] = (LFSRcolor0[43]&LFSRcolor0[688]&LFSRcolor0[179]&LFSRcolor0[259]);
    BiasedRNG[66] = (LFSRcolor0[334]&LFSRcolor0[251]&LFSRcolor0[487]&LFSRcolor0[559]);
    BiasedRNG[67] = (LFSRcolor0[258]&LFSRcolor0[686]&LFSRcolor0[674]&LFSRcolor0[551]);
    BiasedRNG[68] = (LFSRcolor0[826]&LFSRcolor0[659]&LFSRcolor0[131]&LFSRcolor0[257]);
    BiasedRNG[69] = (LFSRcolor0[503]&LFSRcolor0[83]&LFSRcolor0[204]&LFSRcolor0[299]);
    BiasedRNG[70] = (LFSRcolor0[742]&LFSRcolor0[696]&LFSRcolor0[357]&LFSRcolor0[99]);
    BiasedRNG[71] = (LFSRcolor0[580]&LFSRcolor0[795]&LFSRcolor0[354]&LFSRcolor0[129]);
    BiasedRNG[72] = (LFSRcolor0[371]&LFSRcolor0[798]&LFSRcolor0[429]&LFSRcolor0[329]);
    BiasedRNG[73] = (LFSRcolor0[335]&LFSRcolor0[680]&LFSRcolor0[244]&LFSRcolor0[142]);
    BiasedRNG[74] = (LFSRcolor0[103]&LFSRcolor0[664]&LFSRcolor0[78]&LFSRcolor0[490]);
    BiasedRNG[75] = (LFSRcolor0[743]&LFSRcolor0[399]&LFSRcolor0[653]&LFSRcolor0[360]);
    BiasedRNG[76] = (LFSRcolor0[34]&LFSRcolor0[442]&LFSRcolor0[540]&LFSRcolor0[727]);
    BiasedRNG[77] = (LFSRcolor0[402]&LFSRcolor0[679]&LFSRcolor0[55]&LFSRcolor0[774]);
    BiasedRNG[78] = (LFSRcolor0[261]&LFSRcolor0[31]&LFSRcolor0[14]&LFSRcolor0[814]);
    BiasedRNG[79] = (LFSRcolor0[135]&LFSRcolor0[367]&LFSRcolor0[361]&LFSRcolor0[625]);
    BiasedRNG[80] = (LFSRcolor0[549]&LFSRcolor0[634]&LFSRcolor0[377]&LFSRcolor0[684]);
    BiasedRNG[81] = (LFSRcolor0[358]&LFSRcolor0[827]&LFSRcolor0[42]&LFSRcolor0[431]);
    BiasedRNG[82] = (LFSRcolor0[191]&LFSRcolor0[794]&LFSRcolor0[437]&LFSRcolor0[799]);
    BiasedRNG[83] = (LFSRcolor0[438]&LFSRcolor0[46]&LFSRcolor0[702]&LFSRcolor0[486]);
    BiasedRNG[84] = (LFSRcolor0[556]&LFSRcolor0[428]&LFSRcolor0[203]&LFSRcolor0[762]);
    BiasedRNG[85] = (LFSRcolor0[100]&LFSRcolor0[227]&LFSRcolor0[336]&LFSRcolor0[132]);
    BiasedRNG[86] = (LFSRcolor0[425]&LFSRcolor0[415]&LFSRcolor0[577]&LFSRcolor0[600]);
    BiasedRNG[87] = (LFSRcolor0[806]&LFSRcolor0[542]&LFSRcolor0[424]&LFSRcolor0[529]);
    BiasedRNG[88] = (LFSRcolor0[450]&LFSRcolor0[808]&LFSRcolor0[393]&LFSRcolor0[67]);
    BiasedRNG[89] = (LFSRcolor0[489]&LFSRcolor0[215]&LFSRcolor0[444]&LFSRcolor0[448]);
    BiasedRNG[90] = (LFSRcolor0[120]&LFSRcolor0[148]&LFSRcolor0[352]&LFSRcolor0[471]);
    BiasedRNG[91] = (LFSRcolor0[158]&LFSRcolor0[154]&LFSRcolor0[426]&LFSRcolor0[1]);
    BiasedRNG[92] = (LFSRcolor0[112]&LFSRcolor0[459]&LFSRcolor0[247]&LFSRcolor0[692]);
    BiasedRNG[93] = (LFSRcolor0[96]&LFSRcolor0[570]&LFSRcolor0[207]&LFSRcolor0[494]);
    BiasedRNG[94] = (LFSRcolor0[561]&LFSRcolor0[91]&LFSRcolor0[446]&LFSRcolor0[496]);
    BiasedRNG[95] = (LFSRcolor0[604]&LFSRcolor0[189]&LFSRcolor0[92]&LFSRcolor0[356]);
    BiasedRNG[96] = (LFSRcolor0[671]&LFSRcolor0[230]&LFSRcolor0[447]&LFSRcolor0[469]);
    BiasedRNG[97] = (LFSRcolor0[391]&LFSRcolor0[765]&LFSRcolor0[71]&LFSRcolor0[789]);
    BiasedRNG[98] = (LFSRcolor0[282]&LFSRcolor0[624]&LFSRcolor0[499]&LFSRcolor0[509]);
    BiasedRNG[99] = (LFSRcolor0[768]&LFSRcolor0[137]&LFSRcolor0[122]&LFSRcolor0[643]);
    BiasedRNG[100] = (LFSRcolor0[353]&LFSRcolor0[313]&LFSRcolor0[456]&LFSRcolor0[733]);
    BiasedRNG[101] = (LFSRcolor0[726]&LFSRcolor0[421]&LFSRcolor0[668]&LFSRcolor0[492]);
    BiasedRNG[102] = (LFSRcolor0[407]&LFSRcolor0[184]&LFSRcolor0[245]&LFSRcolor0[269]);
    BiasedRNG[103] = (LFSRcolor0[315]&LFSRcolor0[33]&LFSRcolor0[94]&LFSRcolor0[114]);
    BiasedRNG[104] = (LFSRcolor0[801]&LFSRcolor0[818]&LFSRcolor0[552]&LFSRcolor0[508]);
    BiasedRNG[105] = (LFSRcolor0[422]&LFSRcolor0[359]&LFSRcolor0[108]&LFSRcolor0[188]);
    BiasedRNG[106] = (LFSRcolor0[481]&LFSRcolor0[764]&LFSRcolor0[593]&LFSRcolor0[493]);
    BiasedRNG[107] = (LFSRcolor0[21]&LFSRcolor0[260]&LFSRcolor0[474]&LFSRcolor0[264]);
    BiasedRNG[108] = (LFSRcolor0[750]&LFSRcolor0[633]&LFSRcolor0[323]&LFSRcolor0[297]);
    BiasedRNG[109] = (LFSRcolor0[404]&LFSRcolor0[144]&LFSRcolor0[398]&LFSRcolor0[756]);
    BiasedRNG[110] = (LFSRcolor0[72]&LFSRcolor0[291]&LFSRcolor0[309]&LFSRcolor0[746]);
    BiasedRNG[111] = (LFSRcolor0[760]&LFSRcolor0[318]&LFSRcolor0[694]&LFSRcolor0[823]);
    BiasedRNG[112] = (LFSRcolor0[88]&LFSRcolor0[146]&LFSRcolor0[17]&LFSRcolor0[134]);
    BiasedRNG[113] = (LFSRcolor0[232]&LFSRcolor0[708]&LFSRcolor0[212]&LFSRcolor0[725]);
    BiasedRNG[114] = (LFSRcolor0[669]&LFSRcolor0[713]&LFSRcolor0[802]&LFSRcolor0[195]);
    BiasedRNG[115] = (LFSRcolor0[769]&LFSRcolor0[396]&LFSRcolor0[9]&LFSRcolor0[716]);
    BiasedRNG[116] = (LFSRcolor0[145]&LFSRcolor0[710]&LFSRcolor0[620]&LFSRcolor0[581]);
    BiasedRNG[117] = (LFSRcolor0[414]&LFSRcolor0[143]&LFSRcolor0[161]&LFSRcolor0[10]);
    BiasedRNG[118] = (LFSRcolor0[513]&LFSRcolor0[366]&LFSRcolor0[386]&LFSRcolor0[766]);
    BiasedRNG[119] = (LFSRcolor0[734]&LFSRcolor0[711]&LFSRcolor0[231]&LFSRcolor0[598]);
    BiasedRNG[120] = (LFSRcolor0[453]&LFSRcolor0[548]&LFSRcolor0[380]&LFSRcolor0[66]);
    BiasedRNG[121] = (LFSRcolor0[370]&LFSRcolor0[483]&LFSRcolor0[412]&LFSRcolor0[343]);
    BiasedRNG[122] = (LFSRcolor0[435]&LFSRcolor0[418]&LFSRcolor0[463]&LFSRcolor0[268]);
    BiasedRNG[123] = (LFSRcolor0[721]&LFSRcolor0[5]&LFSRcolor0[246]&LFSRcolor0[85]);
    BiasedRNG[124] = (LFSRcolor0[185]&LFSRcolor0[248]&LFSRcolor0[172]&LFSRcolor0[623]);
    BiasedRNG[125] = (LFSRcolor0[328]&LFSRcolor0[150]&LFSRcolor0[75]&LFSRcolor0[186]);
    BiasedRNG[126] = (LFSRcolor0[755]&LFSRcolor0[306]&LFSRcolor0[652]&LFSRcolor0[401]);
    BiasedRNG[127] = (LFSRcolor0[553]&LFSRcolor0[90]&LFSRcolor0[378]&LFSRcolor0[29]);
    BiasedRNG[128] = (LFSRcolor0[629]&LFSRcolor0[293]&LFSRcolor0[52]&LFSRcolor0[759]);
    BiasedRNG[129] = (LFSRcolor0[23]&LFSRcolor0[809]&LFSRcolor0[521]&LFSRcolor0[436]);
    BiasedRNG[130] = (LFSRcolor0[777]&LFSRcolor0[670]&LFSRcolor0[783]&LFSRcolor0[658]);
    BiasedRNG[131] = (LFSRcolor0[56]&LFSRcolor0[319]&LFSRcolor0[534]&LFSRcolor0[701]);
    BiasedRNG[132] = (LFSRcolor0[572]&LFSRcolor0[28]&LFSRcolor0[757]&LFSRcolor0[124]);
    BiasedRNG[133] = (LFSRcolor0[233]&LFSRcolor0[533]&LFSRcolor0[790]&LFSRcolor0[221]);
    BiasedRNG[134] = (LFSRcolor0[562]&LFSRcolor0[15]&LFSRcolor0[631]&LFSRcolor0[683]);
    BiasedRNG[135] = (LFSRcolor0[175]&LFSRcolor0[661]&LFSRcolor0[167]&LFSRcolor0[223]);
    BiasedRNG[136] = (LFSRcolor0[249]&LFSRcolor0[410]&LFSRcolor0[110]&LFSRcolor0[274]);
    BiasedRNG[137] = (LFSRcolor0[322]&LFSRcolor0[89]&LFSRcolor0[252]&LFSRcolor0[515]);
    BiasedRNG[138] = (LFSRcolor0[119]&LFSRcolor0[312]&LFSRcolor0[400]&LFSRcolor0[205]);
    BiasedRNG[139] = (LFSRcolor0[24]&LFSRcolor0[782]&LFSRcolor0[381]&LFSRcolor0[225]);
    BiasedRNG[140] = (LFSRcolor0[495]&LFSRcolor0[699]&LFSRcolor0[11]&LFSRcolor0[420]);
    BiasedRNG[141] = (LFSRcolor0[287]&LFSRcolor0[87]&LFSRcolor0[44]&LFSRcolor0[538]);
    BiasedRNG[142] = (LFSRcolor0[739]&LFSRcolor0[387]&LFSRcolor0[267]&LFSRcolor0[25]);
    BiasedRNG[143] = (LFSRcolor0[77]&LFSRcolor0[754]&LFSRcolor0[583]&LFSRcolor0[586]);
    BiasedRNG[144] = (LFSRcolor0[292]&LFSRcolor0[199]&LFSRcolor0[300]&LFSRcolor0[239]);
    BiasedRNG[145] = (LFSRcolor0[752]&LFSRcolor0[226]&LFSRcolor0[571]&LFSRcolor0[217]);
    BiasedRNG[146] = (LFSRcolor0[337]&LFSRcolor0[767]&LFSRcolor0[74]&LFSRcolor0[485]);
    BiasedRNG[147] = (LFSRcolor0[36]&LFSRcolor0[162]&LFSRcolor0[395]&LFSRcolor0[104]);
    BiasedRNG[148] = (LFSRcolor0[528]&LFSRcolor0[480]&LFSRcolor0[615]&LFSRcolor0[452]);
    BiasedRNG[149] = (LFSRcolor0[190]&LFSRcolor0[60]&LFSRcolor0[523]&LFSRcolor0[327]);
    BiasedRNG[150] = (LFSRcolor0[69]&LFSRcolor0[187]&LFSRcolor0[20]&LFSRcolor0[64]);
    BiasedRNG[151] = (LFSRcolor0[440]&LFSRcolor0[153]&LFSRcolor0[800]&LFSRcolor0[537]);
    BiasedRNG[152] = (LFSRcolor0[811]&LFSRcolor0[535]&LFSRcolor0[98]&LFSRcolor0[423]);
    BiasedRNG[153] = (LFSRcolor0[339]&LFSRcolor0[263]&LFSRcolor0[73]&LFSRcolor0[640]);
    BiasedRNG[154] = (LFSRcolor0[554]&LFSRcolor0[220]&LFSRcolor0[210]&LFSRcolor0[164]);
    BiasedRNG[155] = (LFSRcolor0[505]&LFSRcolor0[723]&LFSRcolor0[394]&LFSRcolor0[298]);
    BiasedRNG[156] = (LFSRcolor0[235]&LFSRcolor0[222]&LFSRcolor0[470]&LFSRcolor0[84]);
    BiasedRNG[157] = (LFSRcolor0[388]&LFSRcolor0[13]&LFSRcolor0[585]&LFSRcolor0[573]);
    BiasedRNG[158] = (LFSRcolor0[47]&LFSRcolor0[277]&LFSRcolor0[574]&LFSRcolor0[321]);
    BiasedRNG[159] = (LFSRcolor0[787]&LFSRcolor0[525]&LFSRcolor0[590]&LFSRcolor0[500]);
    BiasedRNG[160] = (LFSRcolor0[592]&LFSRcolor0[732]&LFSRcolor0[616]&LFSRcolor0[530]);
    BiasedRNG[161] = (LFSRcolor0[151]&LFSRcolor0[747]&LFSRcolor0[728]&LFSRcolor0[237]);
    BiasedRNG[162] = (LFSRcolor0[340]&LFSRcolor0[819]&LFSRcolor0[736]&LFSRcolor0[176]);
    BiasedRNG[163] = (LFSRcolor0[722]&LFSRcolor0[238]&LFSRcolor0[80]&LFSRcolor0[128]);
    BiasedRNG[164] = (LFSRcolor0[177]&LFSRcolor0[796]&LFSRcolor0[689]&LFSRcolor0[457]);
    BiasedRNG[165] = (LFSRcolor0[280]&LFSRcolor0[320]&LFSRcolor0[520]&LFSRcolor0[785]);
    BiasedRNG[166] = (LFSRcolor0[311]&LFSRcolor0[139]&LFSRcolor0[698]&LFSRcolor0[163]);
    BiasedRNG[167] = (LFSRcolor0[641]&LFSRcolor0[18]&LFSRcolor0[125]&LFSRcolor0[630]);
    UnbiasedRNG[0] = LFSRcolor0[430];
    UnbiasedRNG[1] = LFSRcolor0[389];
    UnbiasedRNG[2] = LFSRcolor0[824];
    UnbiasedRNG[3] = LFSRcolor0[645];
    UnbiasedRNG[4] = LFSRcolor0[662];
    UnbiasedRNG[5] = LFSRcolor0[550];
    UnbiasedRNG[6] = LFSRcolor0[458];
    UnbiasedRNG[7] = LFSRcolor0[601];
    UnbiasedRNG[8] = LFSRcolor0[567];
    UnbiasedRNG[9] = LFSRcolor0[603];
    UnbiasedRNG[10] = LFSRcolor0[576];
    UnbiasedRNG[11] = LFSRcolor0[86];
    UnbiasedRNG[12] = LFSRcolor0[676];
    UnbiasedRNG[13] = LFSRcolor0[305];
    UnbiasedRNG[14] = LFSRcolor0[123];
    UnbiasedRNG[15] = LFSRcolor0[326];
    UnbiasedRNG[16] = LFSRcolor0[105];
    UnbiasedRNG[17] = LFSRcolor0[532];
    UnbiasedRNG[18] = LFSRcolor0[433];
    UnbiasedRNG[19] = LFSRcolor0[536];
    UnbiasedRNG[20] = LFSRcolor0[605];
    UnbiasedRNG[21] = LFSRcolor0[362];
    UnbiasedRNG[22] = LFSRcolor0[714];
    UnbiasedRNG[23] = LFSRcolor0[30];
    UnbiasedRNG[24] = LFSRcolor0[582];
    UnbiasedRNG[25] = LFSRcolor0[460];
    UnbiasedRNG[26] = LFSRcolor0[451];
    UnbiasedRNG[27] = LFSRcolor0[434];
    UnbiasedRNG[28] = LFSRcolor0[374];
    UnbiasedRNG[29] = LFSRcolor0[807];
    UnbiasedRNG[30] = LFSRcolor0[462];
    UnbiasedRNG[31] = LFSRcolor0[202];
    UnbiasedRNG[32] = LFSRcolor0[206];
    UnbiasedRNG[33] = LFSRcolor0[351];
    UnbiasedRNG[34] = LFSRcolor0[763];
    UnbiasedRNG[35] = LFSRcolor0[638];
    UnbiasedRNG[36] = LFSRcolor0[608];
    UnbiasedRNG[37] = LFSRcolor0[419];
    UnbiasedRNG[38] = LFSRcolor0[770];
    UnbiasedRNG[39] = LFSRcolor0[32];
    UnbiasedRNG[40] = LFSRcolor0[26];
    UnbiasedRNG[41] = LFSRcolor0[706];
    UnbiasedRNG[42] = LFSRcolor0[793];
    UnbiasedRNG[43] = LFSRcolor0[773];
    UnbiasedRNG[44] = LFSRcolor0[797];
    UnbiasedRNG[45] = LFSRcolor0[406];
    UnbiasedRNG[46] = LFSRcolor0[484];
    UnbiasedRNG[47] = LFSRcolor0[121];
    UnbiasedRNG[48] = LFSRcolor0[156];
    UnbiasedRNG[49] = LFSRcolor0[712];
    UnbiasedRNG[50] = LFSRcolor0[682];
    UnbiasedRNG[51] = LFSRcolor0[236];
    UnbiasedRNG[52] = LFSRcolor0[784];
    UnbiasedRNG[53] = LFSRcolor0[50];
    UnbiasedRNG[54] = LFSRcolor0[497];
    UnbiasedRNG[55] = LFSRcolor0[690];
    UnbiasedRNG[56] = LFSRcolor0[558];
    UnbiasedRNG[57] = LFSRcolor0[411];
    UnbiasedRNG[58] = LFSRcolor0[405];
    UnbiasedRNG[59] = LFSRcolor0[271];
    UnbiasedRNG[60] = LFSRcolor0[705];
    UnbiasedRNG[61] = LFSRcolor0[345];
    UnbiasedRNG[62] = LFSRcolor0[724];
    UnbiasedRNG[63] = LFSRcolor0[644];
    UnbiasedRNG[64] = LFSRcolor0[518];
    UnbiasedRNG[65] = LFSRcolor0[524];
    UnbiasedRNG[66] = LFSRcolor0[557];
    UnbiasedRNG[67] = LFSRcolor0[622];
    UnbiasedRNG[68] = LFSRcolor0[338];
    UnbiasedRNG[69] = LFSRcolor0[41];
    UnbiasedRNG[70] = LFSRcolor0[675];
    UnbiasedRNG[71] = LFSRcolor0[117];
    UnbiasedRNG[72] = LFSRcolor0[647];
    UnbiasedRNG[73] = LFSRcolor0[482];
    UnbiasedRNG[74] = LFSRcolor0[296];
    UnbiasedRNG[75] = LFSRcolor0[49];
    UnbiasedRNG[76] = LFSRcolor0[314];
    UnbiasedRNG[77] = LFSRcolor0[59];
    UnbiasedRNG[78] = LFSRcolor0[776];
    UnbiasedRNG[79] = LFSRcolor0[303];
    UnbiasedRNG[80] = LFSRcolor0[171];
    UnbiasedRNG[81] = LFSRcolor0[504];
    UnbiasedRNG[82] = LFSRcolor0[157];
    UnbiasedRNG[83] = LFSRcolor0[544];
    UnbiasedRNG[84] = LFSRcolor0[786];
    UnbiasedRNG[85] = LFSRcolor0[113];
    UnbiasedRNG[86] = LFSRcolor0[587];
    UnbiasedRNG[87] = LFSRcolor0[101];
    UnbiasedRNG[88] = LFSRcolor0[39];
    UnbiasedRNG[89] = LFSRcolor0[621];
    UnbiasedRNG[90] = LFSRcolor0[748];
    UnbiasedRNG[91] = LFSRcolor0[531];
    UnbiasedRNG[92] = LFSRcolor0[255];
    UnbiasedRNG[93] = LFSRcolor0[432];
    UnbiasedRNG[94] = LFSRcolor0[479];
    UnbiasedRNG[95] = LFSRcolor0[364];
    UnbiasedRNG[96] = LFSRcolor0[805];
    UnbiasedRNG[97] = LFSRcolor0[316];
    UnbiasedRNG[98] = LFSRcolor0[65];
    UnbiasedRNG[99] = LFSRcolor0[660];
    UnbiasedRNG[100] = LFSRcolor0[285];
    UnbiasedRNG[101] = LFSRcolor0[375];
    UnbiasedRNG[102] = LFSRcolor0[219];
    UnbiasedRNG[103] = LFSRcolor0[242];
    UnbiasedRNG[104] = LFSRcolor0[512];
    UnbiasedRNG[105] = LFSRcolor0[539];
    UnbiasedRNG[106] = LFSRcolor0[253];
    UnbiasedRNG[107] = LFSRcolor0[208];
    UnbiasedRNG[108] = LFSRcolor0[663];
    UnbiasedRNG[109] = LFSRcolor0[439];
    UnbiasedRNG[110] = LFSRcolor0[276];
    UnbiasedRNG[111] = LFSRcolor0[681];
    UnbiasedRNG[112] = LFSRcolor0[820];
    UnbiasedRNG[113] = LFSRcolor0[270];
    UnbiasedRNG[114] = LFSRcolor0[522];
    UnbiasedRNG[115] = LFSRcolor0[599];
    UnbiasedRNG[116] = LFSRcolor0[744];
    UnbiasedRNG[117] = LFSRcolor0[761];
    UnbiasedRNG[118] = LFSRcolor0[38];
    UnbiasedRNG[119] = LFSRcolor0[310];
    UnbiasedRNG[120] = LFSRcolor0[70];
    UnbiasedRNG[121] = LFSRcolor0[170];
    UnbiasedRNG[122] = LFSRcolor0[821];
    UnbiasedRNG[123] = LFSRcolor0[174];
    UnbiasedRNG[124] = LFSRcolor0[243];
    UnbiasedRNG[125] = LFSRcolor0[286];
    UnbiasedRNG[126] = LFSRcolor0[241];
    UnbiasedRNG[127] = LFSRcolor0[372];
    UnbiasedRNG[128] = LFSRcolor0[256];
    UnbiasedRNG[129] = LFSRcolor0[607];
    UnbiasedRNG[130] = LFSRcolor0[666];
end

always @(posedge color0_clk) begin
    BiasedRNG[168] = (LFSRcolor1[929]&LFSRcolor1[411]&LFSRcolor1[969]&LFSRcolor1[280]);
    BiasedRNG[169] = (LFSRcolor1[697]&LFSRcolor1[948]&LFSRcolor1[11]&LFSRcolor1[558]);
    BiasedRNG[170] = (LFSRcolor1[572]&LFSRcolor1[71]&LFSRcolor1[958]&LFSRcolor1[767]);
    BiasedRNG[171] = (LFSRcolor1[830]&LFSRcolor1[839]&LFSRcolor1[462]&LFSRcolor1[573]);
    BiasedRNG[172] = (LFSRcolor1[775]&LFSRcolor1[170]&LFSRcolor1[457]&LFSRcolor1[33]);
    BiasedRNG[173] = (LFSRcolor1[679]&LFSRcolor1[478]&LFSRcolor1[203]&LFSRcolor1[984]);
    BiasedRNG[174] = (LFSRcolor1[685]&LFSRcolor1[1001]&LFSRcolor1[901]&LFSRcolor1[379]);
    BiasedRNG[175] = (LFSRcolor1[502]&LFSRcolor1[646]&LFSRcolor1[922]&LFSRcolor1[0]);
    BiasedRNG[176] = (LFSRcolor1[737]&LFSRcolor1[731]&LFSRcolor1[119]&LFSRcolor1[317]);
    BiasedRNG[177] = (LFSRcolor1[145]&LFSRcolor1[431]&LFSRcolor1[136]&LFSRcolor1[348]);
    BiasedRNG[178] = (LFSRcolor1[628]&LFSRcolor1[950]&LFSRcolor1[754]&LFSRcolor1[470]);
    BiasedRNG[179] = (LFSRcolor1[230]&LFSRcolor1[916]&LFSRcolor1[568]&LFSRcolor1[963]);
    BiasedRNG[180] = (LFSRcolor1[882]&LFSRcolor1[113]&LFSRcolor1[930]&LFSRcolor1[437]);
    BiasedRNG[181] = (LFSRcolor1[135]&LFSRcolor1[279]&LFSRcolor1[32]&LFSRcolor1[425]);
    BiasedRNG[182] = (LFSRcolor1[523]&LFSRcolor1[710]&LFSRcolor1[68]&LFSRcolor1[131]);
    BiasedRNG[183] = (LFSRcolor1[555]&LFSRcolor1[757]&LFSRcolor1[427]&LFSRcolor1[387]);
    BiasedRNG[184] = (LFSRcolor1[407]&LFSRcolor1[400]&LFSRcolor1[726]&LFSRcolor1[197]);
    BiasedRNG[185] = (LFSRcolor1[966]&LFSRcolor1[816]&LFSRcolor1[385]&LFSRcolor1[994]);
    BiasedRNG[186] = (LFSRcolor1[349]&LFSRcolor1[388]&LFSRcolor1[911]&LFSRcolor1[567]);
    BiasedRNG[187] = (LFSRcolor1[786]&LFSRcolor1[159]&LFSRcolor1[458]&LFSRcolor1[305]);
    BiasedRNG[188] = (LFSRcolor1[643]&LFSRcolor1[408]&LFSRcolor1[73]&LFSRcolor1[964]);
    BiasedRNG[189] = (LFSRcolor1[917]&LFSRcolor1[1006]&LFSRcolor1[753]&LFSRcolor1[673]);
    BiasedRNG[190] = (LFSRcolor1[188]&LFSRcolor1[869]&LFSRcolor1[968]&LFSRcolor1[121]);
    BiasedRNG[191] = (LFSRcolor1[689]&LFSRcolor1[722]&LFSRcolor1[1008]&LFSRcolor1[863]);
    BiasedRNG[192] = (LFSRcolor1[819]&LFSRcolor1[320]&LFSRcolor1[115]&LFSRcolor1[93]);
    BiasedRNG[193] = (LFSRcolor1[552]&LFSRcolor1[465]&LFSRcolor1[608]&LFSRcolor1[727]);
    BiasedRNG[194] = (LFSRcolor1[51]&LFSRcolor1[933]&LFSRcolor1[978]&LFSRcolor1[971]);
    BiasedRNG[195] = (LFSRcolor1[625]&LFSRcolor1[401]&LFSRcolor1[541]&LFSRcolor1[189]);
    BiasedRNG[196] = (LFSRcolor1[504]&LFSRcolor1[820]&LFSRcolor1[972]&LFSRcolor1[584]);
    BiasedRNG[197] = (LFSRcolor1[690]&LFSRcolor1[238]&LFSRcolor1[947]&LFSRcolor1[663]);
    BiasedRNG[198] = (LFSRcolor1[773]&LFSRcolor1[133]&LFSRcolor1[490]&LFSRcolor1[103]);
    BiasedRNG[199] = (LFSRcolor1[324]&LFSRcolor1[840]&LFSRcolor1[294]&LFSRcolor1[199]);
    BiasedRNG[200] = (LFSRcolor1[870]&LFSRcolor1[709]&LFSRcolor1[733]&LFSRcolor1[879]);
    BiasedRNG[201] = (LFSRcolor1[758]&LFSRcolor1[311]&LFSRcolor1[307]&LFSRcolor1[798]);
    BiasedRNG[202] = (LFSRcolor1[707]&LFSRcolor1[474]&LFSRcolor1[406]&LFSRcolor1[376]);
    BiasedRNG[203] = (LFSRcolor1[50]&LFSRcolor1[168]&LFSRcolor1[662]&LFSRcolor1[214]);
    BiasedRNG[204] = (LFSRcolor1[480]&LFSRcolor1[600]&LFSRcolor1[67]&LFSRcolor1[62]);
    BiasedRNG[205] = (LFSRcolor1[506]&LFSRcolor1[973]&LFSRcolor1[479]&LFSRcolor1[614]);
    BiasedRNG[206] = (LFSRcolor1[355]&LFSRcolor1[866]&LFSRcolor1[8]&LFSRcolor1[418]);
    BiasedRNG[207] = (LFSRcolor1[546]&LFSRcolor1[191]&LFSRcolor1[501]&LFSRcolor1[249]);
    BiasedRNG[208] = (LFSRcolor1[29]&LFSRcolor1[992]&LFSRcolor1[509]&LFSRcolor1[769]);
    BiasedRNG[209] = (LFSRcolor1[977]&LFSRcolor1[398]&LFSRcolor1[6]&LFSRcolor1[629]);
    BiasedRNG[210] = (LFSRcolor1[43]&LFSRcolor1[993]&LFSRcolor1[615]&LFSRcolor1[485]);
    BiasedRNG[211] = (LFSRcolor1[642]&LFSRcolor1[120]&LFSRcolor1[245]&LFSRcolor1[239]);
    BiasedRNG[212] = (LFSRcolor1[678]&LFSRcolor1[659]&LFSRcolor1[261]&LFSRcolor1[291]);
    BiasedRNG[213] = (LFSRcolor1[335]&LFSRcolor1[783]&LFSRcolor1[301]&LFSRcolor1[326]);
    BiasedRNG[214] = (LFSRcolor1[723]&LFSRcolor1[953]&LFSRcolor1[591]&LFSRcolor1[809]);
    BiasedRNG[215] = (LFSRcolor1[276]&LFSRcolor1[828]&LFSRcolor1[684]&LFSRcolor1[47]);
    BiasedRNG[216] = (LFSRcolor1[599]&LFSRcolor1[414]&LFSRcolor1[652]&LFSRcolor1[27]);
    BiasedRNG[217] = (LFSRcolor1[875]&LFSRcolor1[477]&LFSRcolor1[702]&LFSRcolor1[207]);
    BiasedRNG[218] = (LFSRcolor1[434]&LFSRcolor1[80]&LFSRcolor1[21]&LFSRcolor1[905]);
    BiasedRNG[219] = (LFSRcolor1[63]&LFSRcolor1[999]&LFSRcolor1[799]&LFSRcolor1[30]);
    BiasedRNG[220] = (LFSRcolor1[915]&LFSRcolor1[393]&LFSRcolor1[475]&LFSRcolor1[868]);
    BiasedRNG[221] = (LFSRcolor1[272]&LFSRcolor1[186]&LFSRcolor1[692]&LFSRcolor1[210]);
    BiasedRNG[222] = (LFSRcolor1[794]&LFSRcolor1[653]&LFSRcolor1[37]&LFSRcolor1[461]);
    BiasedRNG[223] = (LFSRcolor1[196]&LFSRcolor1[871]&LFSRcolor1[821]&LFSRcolor1[126]);
    BiasedRNG[224] = (LFSRcolor1[842]&LFSRcolor1[476]&LFSRcolor1[817]&LFSRcolor1[499]);
    BiasedRNG[225] = (LFSRcolor1[25]&LFSRcolor1[565]&LFSRcolor1[35]&LFSRcolor1[101]);
    BiasedRNG[226] = (LFSRcolor1[764]&LFSRcolor1[654]&LFSRcolor1[246]&LFSRcolor1[534]);
    BiasedRNG[227] = (LFSRcolor1[811]&LFSRcolor1[708]&LFSRcolor1[900]&LFSRcolor1[149]);
    BiasedRNG[228] = (LFSRcolor1[296]&LFSRcolor1[281]&LFSRcolor1[826]&LFSRcolor1[666]);
    BiasedRNG[229] = (LFSRcolor1[560]&LFSRcolor1[127]&LFSRcolor1[537]&LFSRcolor1[996]);
    BiasedRNG[230] = (LFSRcolor1[651]&LFSRcolor1[74]&LFSRcolor1[396]&LFSRcolor1[303]);
    BiasedRNG[231] = (LFSRcolor1[162]&LFSRcolor1[638]&LFSRcolor1[656]&LFSRcolor1[138]);
    BiasedRNG[232] = (LFSRcolor1[374]&LFSRcolor1[645]&LFSRcolor1[384]&LFSRcolor1[227]);
    BiasedRNG[233] = (LFSRcolor1[175]&LFSRcolor1[766]&LFSRcolor1[902]&LFSRcolor1[83]);
    BiasedRNG[234] = (LFSRcolor1[267]&LFSRcolor1[39]&LFSRcolor1[420]&LFSRcolor1[661]);
    BiasedRNG[235] = (LFSRcolor1[890]&LFSRcolor1[446]&LFSRcolor1[522]&LFSRcolor1[248]);
    BiasedRNG[236] = (LFSRcolor1[95]&LFSRcolor1[460]&LFSRcolor1[117]&LFSRcolor1[386]);
    BiasedRNG[237] = (LFSRcolor1[157]&LFSRcolor1[329]&LFSRcolor1[150]&LFSRcolor1[782]);
    BiasedRNG[238] = (LFSRcolor1[853]&LFSRcolor1[545]&LFSRcolor1[527]&LFSRcolor1[891]);
    BiasedRNG[239] = (LFSRcolor1[432]&LFSRcolor1[834]&LFSRcolor1[743]&LFSRcolor1[728]);
    BiasedRNG[240] = (LFSRcolor1[424]&LFSRcolor1[854]&LFSRcolor1[185]&LFSRcolor1[332]);
    BiasedRNG[241] = (LFSRcolor1[56]&LFSRcolor1[951]&LFSRcolor1[601]&LFSRcolor1[985]);
    BiasedRNG[242] = (LFSRcolor1[212]&LFSRcolor1[206]&LFSRcolor1[466]&LFSRcolor1[9]);
    BiasedRNG[243] = (LFSRcolor1[862]&LFSRcolor1[221]&LFSRcolor1[410]&LFSRcolor1[626]);
    BiasedRNG[244] = (LFSRcolor1[293]&LFSRcolor1[176]&LFSRcolor1[359]&LFSRcolor1[974]);
    BiasedRNG[245] = (LFSRcolor1[832]&LFSRcolor1[780]&LFSRcolor1[213]&LFSRcolor1[397]);
    BiasedRNG[246] = (LFSRcolor1[445]&LFSRcolor1[192]&LFSRcolor1[580]&LFSRcolor1[333]);
    BiasedRNG[247] = (LFSRcolor1[4]&LFSRcolor1[287]&LFSRcolor1[104]&LFSRcolor1[945]);
    BiasedRNG[248] = (LFSRcolor1[621]&LFSRcolor1[229]&LFSRcolor1[718]&LFSRcolor1[865]);
    BiasedRNG[249] = (LFSRcolor1[430]&LFSRcolor1[703]&LFSRcolor1[128]&LFSRcolor1[624]);
    BiasedRNG[250] = (LFSRcolor1[378]&LFSRcolor1[389]&LFSRcolor1[613]&LFSRcolor1[90]);
    BiasedRNG[251] = (LFSRcolor1[551]&LFSRcolor1[680]&LFSRcolor1[169]&LFSRcolor1[451]);
    BiasedRNG[252] = (LFSRcolor1[838]&LFSRcolor1[464]&LFSRcolor1[695]&LFSRcolor1[837]);
    BiasedRNG[253] = (LFSRcolor1[807]&LFSRcolor1[943]&LFSRcolor1[639]&LFSRcolor1[899]);
    BiasedRNG[254] = (LFSRcolor1[776]&LFSRcolor1[706]&LFSRcolor1[511]&LFSRcolor1[140]);
    BiasedRNG[255] = (LFSRcolor1[72]&LFSRcolor1[306]&LFSRcolor1[589]&LFSRcolor1[729]);
    BiasedRNG[256] = (LFSRcolor1[1002]&LFSRcolor1[97]&LFSRcolor1[561]&LFSRcolor1[880]);
    BiasedRNG[257] = (LFSRcolor1[322]&LFSRcolor1[741]&LFSRcolor1[756]&LFSRcolor1[841]);
    BiasedRNG[258] = (LFSRcolor1[677]&LFSRcolor1[264]&LFSRcolor1[934]&LFSRcolor1[98]);
    BiasedRNG[259] = (LFSRcolor1[403]&LFSRcolor1[236]&LFSRcolor1[931]&LFSRcolor1[228]);
    BiasedRNG[260] = (LFSRcolor1[713]&LFSRcolor1[524]&LFSRcolor1[177]&LFSRcolor1[777]);
    BiasedRNG[261] = (LFSRcolor1[328]&LFSRcolor1[740]&LFSRcolor1[835]&LFSRcolor1[790]);
    BiasedRNG[262] = (LFSRcolor1[231]&LFSRcolor1[277]&LFSRcolor1[129]&LFSRcolor1[260]);
    BiasedRNG[263] = (LFSRcolor1[1010]&LFSRcolor1[314]&LFSRcolor1[350]&LFSRcolor1[763]);
    BiasedRNG[264] = (LFSRcolor1[627]&LFSRcolor1[873]&LFSRcolor1[361]&LFSRcolor1[299]);
    BiasedRNG[265] = (LFSRcolor1[513]&LFSRcolor1[347]&LFSRcolor1[636]&LFSRcolor1[57]);
    BiasedRNG[266] = (LFSRcolor1[919]&LFSRcolor1[59]&LFSRcolor1[944]&LFSRcolor1[796]);
    BiasedRNG[267] = (LFSRcolor1[793]&LFSRcolor1[346]&LFSRcolor1[60]&LFSRcolor1[918]);
    BiasedRNG[268] = (LFSRcolor1[70]&LFSRcolor1[247]&LFSRcolor1[507]&LFSRcolor1[193]);
    BiasedRNG[269] = (LFSRcolor1[909]&LFSRcolor1[172]&LFSRcolor1[49]&LFSRcolor1[467]);
    BiasedRNG[270] = (LFSRcolor1[520]&LFSRcolor1[941]&LFSRcolor1[473]&LFSRcolor1[982]);
    BiasedRNG[271] = (LFSRcolor1[141]&LFSRcolor1[488]&LFSRcolor1[89]&LFSRcolor1[855]);
    BiasedRNG[272] = (LFSRcolor1[298]&LFSRcolor1[925]&LFSRcolor1[559]&LFSRcolor1[803]);
    BiasedRNG[273] = (LFSRcolor1[536]&LFSRcolor1[547]&LFSRcolor1[691]&LFSRcolor1[886]);
    BiasedRNG[274] = (LFSRcolor1[539]&LFSRcolor1[368]&LFSRcolor1[698]&LFSRcolor1[575]);
    BiasedRNG[275] = (LFSRcolor1[438]&LFSRcolor1[1000]&LFSRcolor1[372]&LFSRcolor1[288]);
    BiasedRNG[276] = (LFSRcolor1[269]&LFSRcolor1[275]&LFSRcolor1[455]&LFSRcolor1[700]);
    BiasedRNG[277] = (LFSRcolor1[570]&LFSRcolor1[381]&LFSRcolor1[779]&LFSRcolor1[557]);
    BiasedRNG[278] = (LFSRcolor1[864]&LFSRcolor1[577]&LFSRcolor1[949]&LFSRcolor1[883]);
    BiasedRNG[279] = (LFSRcolor1[18]&LFSRcolor1[459]&LFSRcolor1[491]&LFSRcolor1[42]);
    BiasedRNG[280] = (LFSRcolor1[631]&LFSRcolor1[954]&LFSRcolor1[562]&LFSRcolor1[789]);
    BiasedRNG[281] = (LFSRcolor1[237]&LFSRcolor1[694]&LFSRcolor1[576]&LFSRcolor1[844]);
    BiasedRNG[282] = (LFSRcolor1[123]&LFSRcolor1[734]&LFSRcolor1[144]&LFSRcolor1[156]);
    BiasedRNG[283] = (LFSRcolor1[851]&LFSRcolor1[531]&LFSRcolor1[812]&LFSRcolor1[549]);
    BiasedRNG[284] = (LFSRcolor1[748]&LFSRcolor1[858]&LFSRcolor1[990]&LFSRcolor1[153]);
    BiasedRNG[285] = (LFSRcolor1[923]&LFSRcolor1[223]&LFSRcolor1[111]&LFSRcolor1[340]);
    BiasedRNG[286] = (LFSRcolor1[250]&LFSRcolor1[612]&LFSRcolor1[112]&LFSRcolor1[716]);
    BiasedRNG[287] = (LFSRcolor1[152]&LFSRcolor1[79]&LFSRcolor1[976]&LFSRcolor1[334]);
    BiasedRNG[288] = (LFSRcolor1[166]&LFSRcolor1[518]&LFSRcolor1[184]&LFSRcolor1[271]);
    BiasedRNG[289] = (LFSRcolor1[970]&LFSRcolor1[927]&LFSRcolor1[668]&LFSRcolor1[772]);
    BiasedRNG[290] = (LFSRcolor1[265]&LFSRcolor1[898]&LFSRcolor1[224]&LFSRcolor1[146]);
    BiasedRNG[291] = (LFSRcolor1[845]&LFSRcolor1[472]&LFSRcolor1[17]&LFSRcolor1[525]);
    BiasedRNG[292] = (LFSRcolor1[132]&LFSRcolor1[380]&LFSRcolor1[382]&LFSRcolor1[856]);
    BiasedRNG[293] = (LFSRcolor1[96]&LFSRcolor1[910]&LFSRcolor1[495]&LFSRcolor1[282]);
    BiasedRNG[294] = (LFSRcolor1[337]&LFSRcolor1[961]&LFSRcolor1[183]&LFSRcolor1[163]);
    BiasedRNG[295] = (LFSRcolor1[658]&LFSRcolor1[440]&LFSRcolor1[671]&LFSRcolor1[492]);
    BiasedRNG[296] = (LFSRcolor1[771]&LFSRcolor1[313]&LFSRcolor1[226]&LFSRcolor1[124]);
    BiasedRNG[297] = (LFSRcolor1[699]&LFSRcolor1[308]&LFSRcolor1[234]&LFSRcolor1[998]);
    BiasedRNG[298] = (LFSRcolor1[967]&LFSRcolor1[394]&LFSRcolor1[521]&LFSRcolor1[715]);
    BiasedRNG[299] = (LFSRcolor1[579]&LFSRcolor1[92]&LFSRcolor1[717]&LFSRcolor1[500]);
    BiasedRNG[300] = (LFSRcolor1[481]&LFSRcolor1[241]&LFSRcolor1[563]&LFSRcolor1[38]);
    BiasedRNG[301] = (LFSRcolor1[366]&LFSRcolor1[395]&LFSRcolor1[443]&LFSRcolor1[489]);
    BiasedRNG[302] = (LFSRcolor1[938]&LFSRcolor1[921]&LFSRcolor1[22]&LFSRcolor1[924]);
    BiasedRNG[303] = (LFSRcolor1[920]&LFSRcolor1[423]&LFSRcolor1[202]&LFSRcolor1[218]);
    BiasedRNG[304] = (LFSRcolor1[530]&LFSRcolor1[704]&LFSRcolor1[894]&LFSRcolor1[161]);
    BiasedRNG[305] = (LFSRcolor1[884]&LFSRcolor1[510]&LFSRcolor1[55]&LFSRcolor1[893]);
    BiasedRNG[306] = (LFSRcolor1[583]&LFSRcolor1[788]&LFSRcolor1[981]&LFSRcolor1[928]);
    BiasedRNG[307] = (LFSRcolor1[848]&LFSRcolor1[219]&LFSRcolor1[892]&LFSRcolor1[532]);
    BiasedRNG[308] = (LFSRcolor1[94]&LFSRcolor1[897]&LFSRcolor1[182]&LFSRcolor1[860]);
    BiasedRNG[309] = (LFSRcolor1[23]&LFSRcolor1[399]&LFSRcolor1[676]&LFSRcolor1[913]);
    BiasedRNG[310] = (LFSRcolor1[266]&LFSRcolor1[160]&LFSRcolor1[327]&LFSRcolor1[339]);
    BiasedRNG[311] = (LFSRcolor1[956]&LFSRcolor1[304]&LFSRcolor1[211]&LFSRcolor1[20]);
    BiasedRNG[312] = (LFSRcolor1[450]&LFSRcolor1[58]&LFSRcolor1[1]&LFSRcolor1[665]);
    BiasedRNG[313] = (LFSRcolor1[825]&LFSRcolor1[31]&LFSRcolor1[371]&LFSRcolor1[233]);
    BiasedRNG[314] = (LFSRcolor1[484]&LFSRcolor1[528]&LFSRcolor1[914]&LFSRcolor1[818]);
    BiasedRNG[315] = (LFSRcolor1[975]&LFSRcolor1[877]&LFSRcolor1[297]&LFSRcolor1[362]);
    BiasedRNG[316] = (LFSRcolor1[957]&LFSRcolor1[962]&LFSRcolor1[309]&LFSRcolor1[77]);
    BiasedRNG[317] = (LFSRcolor1[822]&LFSRcolor1[363]&LFSRcolor1[810]&LFSRcolor1[15]);
    BiasedRNG[318] = (LFSRcolor1[40]&LFSRcolor1[610]&LFSRcolor1[831]&LFSRcolor1[632]);
    BiasedRNG[319] = (LFSRcolor1[609]&LFSRcolor1[526]&LFSRcolor1[667]&LFSRcolor1[720]);
    BiasedRNG[320] = (LFSRcolor1[1003]&LFSRcolor1[785]&LFSRcolor1[587]&LFSRcolor1[553]);
    BiasedRNG[321] = (LFSRcolor1[604]&LFSRcolor1[289]&LFSRcolor1[813]&LFSRcolor1[849]);
    BiasedRNG[322] = (LFSRcolor1[730]&LFSRcolor1[711]&LFSRcolor1[415]&LFSRcolor1[597]);
    BiasedRNG[323] = (LFSRcolor1[419]&LFSRcolor1[180]&LFSRcolor1[496]&LFSRcolor1[542]);
    BiasedRNG[324] = (LFSRcolor1[486]&LFSRcolor1[745]&LFSRcolor1[417]&LFSRcolor1[158]);
    BiasedRNG[325] = (LFSRcolor1[505]&LFSRcolor1[588]&LFSRcolor1[300]&LFSRcolor1[257]);
    BiasedRNG[326] = (LFSRcolor1[377]&LFSRcolor1[44]&LFSRcolor1[174]&LFSRcolor1[686]);
    BiasedRNG[327] = (LFSRcolor1[617]&LFSRcolor1[498]&LFSRcolor1[660]&LFSRcolor1[354]);
    BiasedRNG[328] = (LFSRcolor1[874]&LFSRcolor1[742]&LFSRcolor1[540]&LFSRcolor1[118]);
    BiasedRNG[329] = (LFSRcolor1[338]&LFSRcolor1[755]&LFSRcolor1[12]&LFSRcolor1[187]);
    BiasedRNG[330] = (LFSRcolor1[787]&LFSRcolor1[290]&LFSRcolor1[980]&LFSRcolor1[114]);
    BiasedRNG[331] = (LFSRcolor1[318]&LFSRcolor1[548]&LFSRcolor1[669]&LFSRcolor1[323]);
    BiasedRNG[332] = (LFSRcolor1[942]&LFSRcolor1[402]&LFSRcolor1[696]&LFSRcolor1[635]);
    BiasedRNG[333] = (LFSRcolor1[955]&LFSRcolor1[791]&LFSRcolor1[302]&LFSRcolor1[806]);
    BiasedRNG[334] = (LFSRcolor1[352]&LFSRcolor1[341]&LFSRcolor1[752]&LFSRcolor1[404]);
    BiasedRNG[335] = (LFSRcolor1[564]&LFSRcolor1[253]&LFSRcolor1[738]&LFSRcolor1[171]);
    BiasedRNG[336] = (LFSRcolor1[208]&LFSRcolor1[543]&LFSRcolor1[634]&LFSRcolor1[286]);
    BiasedRNG[337] = (LFSRcolor1[142]&LFSRcolor1[76]&LFSRcolor1[887]&LFSRcolor1[284]);
    BiasedRNG[338] = (LFSRcolor1[179]&LFSRcolor1[13]&LFSRcolor1[657]&LFSRcolor1[315]);
    BiasedRNG[339] = (LFSRcolor1[781]&LFSRcolor1[538]&LFSRcolor1[19]&LFSRcolor1[108]);
    BiasedRNG[340] = (LFSRcolor1[529]&LFSRcolor1[497]&LFSRcolor1[225]&LFSRcolor1[392]);
    BiasedRNG[341] = (LFSRcolor1[217]&LFSRcolor1[2]&LFSRcolor1[683]&LFSRcolor1[468]);
    BiasedRNG[342] = (LFSRcolor1[48]&LFSRcolor1[321]&LFSRcolor1[109]&LFSRcolor1[82]);
    BiasedRNG[343] = (LFSRcolor1[439]&LFSRcolor1[595]&LFSRcolor1[827]&LFSRcolor1[672]);
    BiasedRNG[344] = (LFSRcolor1[343]&LFSRcolor1[34]&LFSRcolor1[907]&LFSRcolor1[198]);
    BiasedRNG[345] = (LFSRcolor1[797]&LFSRcolor1[566]&LFSRcolor1[421]&LFSRcolor1[391]);
    BiasedRNG[346] = (LFSRcolor1[78]&LFSRcolor1[997]&LFSRcolor1[122]&LFSRcolor1[778]);
    BiasedRNG[347] = (LFSRcolor1[846]&LFSRcolor1[453]&LFSRcolor1[201]&LFSRcolor1[65]);
    BiasedRNG[348] = (LFSRcolor1[751]&LFSRcolor1[620]&LFSRcolor1[768]&LFSRcolor1[370]);
    BiasedRNG[349] = (LFSRcolor1[165]&LFSRcolor1[833]&LFSRcolor1[721]&LFSRcolor1[155]);
    BiasedRNG[350] = (LFSRcolor1[824]&LFSRcolor1[965]&LFSRcolor1[759]&LFSRcolor1[220]);
    BiasedRNG[351] = (LFSRcolor1[618]&LFSRcolor1[16]&LFSRcolor1[749]&LFSRcolor1[10]);
    BiasedRNG[352] = (LFSRcolor1[843]&LFSRcolor1[316]&LFSRcolor1[61]&LFSRcolor1[554]);
    BiasedRNG[353] = (LFSRcolor1[268]&LFSRcolor1[650]&LFSRcolor1[606]&LFSRcolor1[983]);
    BiasedRNG[354] = (LFSRcolor1[173]&LFSRcolor1[147]&LFSRcolor1[383]&LFSRcolor1[448]);
    BiasedRNG[355] = (LFSRcolor1[829]&LFSRcolor1[582]&LFSRcolor1[881]&LFSRcolor1[75]);
    BiasedRNG[356] = (LFSRcolor1[493]&LFSRcolor1[7]&LFSRcolor1[857]&LFSRcolor1[369]);
    BiasedRNG[357] = (LFSRcolor1[876]&LFSRcolor1[750]&LFSRcolor1[116]&LFSRcolor1[53]);
    BiasedRNG[358] = (LFSRcolor1[805]&LFSRcolor1[784]&LFSRcolor1[342]&LFSRcolor1[88]);
    BiasedRNG[359] = (LFSRcolor1[514]&LFSRcolor1[508]&LFSRcolor1[312]&LFSRcolor1[487]);
    BiasedRNG[360] = (LFSRcolor1[205]&LFSRcolor1[774]&LFSRcolor1[295]&LFSRcolor1[878]);
    BiasedRNG[361] = (LFSRcolor1[435]&LFSRcolor1[655]&LFSRcolor1[895]&LFSRcolor1[619]);
    BiasedRNG[362] = (LFSRcolor1[991]&LFSRcolor1[623]&LFSRcolor1[390]&LFSRcolor1[336]);
    BiasedRNG[363] = (LFSRcolor1[447]&LFSRcolor1[649]&LFSRcolor1[515]&LFSRcolor1[167]);
    BiasedRNG[364] = (LFSRcolor1[412]&LFSRcolor1[263]&LFSRcolor1[682]&LFSRcolor1[344]);
    BiasedRNG[365] = (LFSRcolor1[674]&LFSRcolor1[940]&LFSRcolor1[194]&LFSRcolor1[102]);
    BiasedRNG[366] = (LFSRcolor1[952]&LFSRcolor1[181]&LFSRcolor1[283]&LFSRcolor1[517]);
    BiasedRNG[367] = (LFSRcolor1[594]&LFSRcolor1[814]&LFSRcolor1[232]&LFSRcolor1[190]);
    BiasedRNG[368] = (LFSRcolor1[64]&LFSRcolor1[442]&LFSRcolor1[867]&LFSRcolor1[195]);
    BiasedRNG[369] = (LFSRcolor1[252]&LFSRcolor1[54]&LFSRcolor1[251]&LFSRcolor1[747]);
    BiasedRNG[370] = (LFSRcolor1[216]&LFSRcolor1[360]&LFSRcolor1[148]&LFSRcolor1[852]);
    BiasedRNG[371] = (LFSRcolor1[240]&LFSRcolor1[746]&LFSRcolor1[735]&LFSRcolor1[243]);
    BiasedRNG[372] = (LFSRcolor1[375]&LFSRcolor1[544]&LFSRcolor1[242]&LFSRcolor1[593]);
    BiasedRNG[373] = (LFSRcolor1[936]&LFSRcolor1[256]&LFSRcolor1[906]&LFSRcolor1[770]);
    BiasedRNG[374] = (LFSRcolor1[178]&LFSRcolor1[130]&LFSRcolor1[52]&LFSRcolor1[761]);
    BiasedRNG[375] = (LFSRcolor1[765]&LFSRcolor1[585]&LFSRcolor1[644]&LFSRcolor1[416]);
    BiasedRNG[376] = (LFSRcolor1[714]&LFSRcolor1[959]&LFSRcolor1[648]&LFSRcolor1[28]);
    BiasedRNG[377] = (LFSRcolor1[215]&LFSRcolor1[872]&LFSRcolor1[353]&LFSRcolor1[744]);
    BiasedRNG[378] = (LFSRcolor1[69]&LFSRcolor1[847]&LFSRcolor1[762]&LFSRcolor1[452]);
    BiasedRNG[379] = (LFSRcolor1[262]&LFSRcolor1[712]&LFSRcolor1[641]&LFSRcolor1[413]);
    BiasedRNG[380] = (LFSRcolor1[637]&LFSRcolor1[926]&LFSRcolor1[45]&LFSRcolor1[693]);
    BiasedRNG[381] = (LFSRcolor1[235]&LFSRcolor1[633]&LFSRcolor1[405]&LFSRcolor1[889]);
    BiasedRNG[382] = (LFSRcolor1[244]&LFSRcolor1[802]&LFSRcolor1[351]&LFSRcolor1[850]);
    UnbiasedRNG[131] = LFSRcolor1[26];
    UnbiasedRNG[132] = LFSRcolor1[105];
    UnbiasedRNG[133] = LFSRcolor1[804];
    UnbiasedRNG[134] = LFSRcolor1[571];
    UnbiasedRNG[135] = LFSRcolor1[800];
    UnbiasedRNG[136] = LFSRcolor1[285];
    UnbiasedRNG[137] = LFSRcolor1[134];
    UnbiasedRNG[138] = LFSRcolor1[139];
    UnbiasedRNG[139] = LFSRcolor1[512];
    UnbiasedRNG[140] = LFSRcolor1[908];
    UnbiasedRNG[141] = LFSRcolor1[436];
    UnbiasedRNG[142] = LFSRcolor1[106];
    UnbiasedRNG[143] = LFSRcolor1[687];
    UnbiasedRNG[144] = LFSRcolor1[273];
    UnbiasedRNG[145] = LFSRcolor1[701];
    UnbiasedRNG[146] = LFSRcolor1[100];
    UnbiasedRNG[147] = LFSRcolor1[795];
    UnbiasedRNG[148] = LFSRcolor1[815];
    UnbiasedRNG[149] = LFSRcolor1[603];
    UnbiasedRNG[150] = LFSRcolor1[519];
    UnbiasedRNG[151] = LFSRcolor1[939];
    UnbiasedRNG[152] = LFSRcolor1[935];
    UnbiasedRNG[153] = LFSRcolor1[454];
    UnbiasedRNG[154] = LFSRcolor1[91];
    UnbiasedRNG[155] = LFSRcolor1[979];
    UnbiasedRNG[156] = LFSRcolor1[107];
    UnbiasedRNG[157] = LFSRcolor1[590];
    UnbiasedRNG[158] = LFSRcolor1[471];
    UnbiasedRNG[159] = LFSRcolor1[556];
    UnbiasedRNG[160] = LFSRcolor1[428];
    UnbiasedRNG[161] = LFSRcolor1[373];
    UnbiasedRNG[162] = LFSRcolor1[125];
    UnbiasedRNG[163] = LFSRcolor1[449];
    UnbiasedRNG[164] = LFSRcolor1[1011];
    UnbiasedRNG[165] = LFSRcolor1[640];
    UnbiasedRNG[166] = LFSRcolor1[664];
    UnbiasedRNG[167] = LFSRcolor1[688];
    UnbiasedRNG[168] = LFSRcolor1[357];
    UnbiasedRNG[169] = LFSRcolor1[1005];
    UnbiasedRNG[170] = LFSRcolor1[885];
    UnbiasedRNG[171] = LFSRcolor1[331];
    UnbiasedRNG[172] = LFSRcolor1[630];
    UnbiasedRNG[173] = LFSRcolor1[719];
    UnbiasedRNG[174] = LFSRcolor1[586];
    UnbiasedRNG[175] = LFSRcolor1[255];
    UnbiasedRNG[176] = LFSRcolor1[903];
    UnbiasedRNG[177] = LFSRcolor1[808];
    UnbiasedRNG[178] = LFSRcolor1[705];
    UnbiasedRNG[179] = LFSRcolor1[482];
    UnbiasedRNG[180] = LFSRcolor1[861];
    UnbiasedRNG[181] = LFSRcolor1[81];
    UnbiasedRNG[182] = LFSRcolor1[592];
    UnbiasedRNG[183] = LFSRcolor1[611];
    UnbiasedRNG[184] = LFSRcolor1[732];
    UnbiasedRNG[185] = LFSRcolor1[319];
    UnbiasedRNG[186] = LFSRcolor1[516];
    UnbiasedRNG[187] = LFSRcolor1[681];
    UnbiasedRNG[188] = LFSRcolor1[607];
    UnbiasedRNG[189] = LFSRcolor1[912];
    UnbiasedRNG[190] = LFSRcolor1[278];
    UnbiasedRNG[191] = LFSRcolor1[310];
    UnbiasedRNG[192] = LFSRcolor1[143];
    UnbiasedRNG[193] = LFSRcolor1[550];
    UnbiasedRNG[194] = LFSRcolor1[99];
    UnbiasedRNG[195] = LFSRcolor1[736];
    UnbiasedRNG[196] = LFSRcolor1[87];
    UnbiasedRNG[197] = LFSRcolor1[330];
    UnbiasedRNG[198] = LFSRcolor1[946];
    UnbiasedRNG[199] = LFSRcolor1[988];
    UnbiasedRNG[200] = LFSRcolor1[85];
    UnbiasedRNG[201] = LFSRcolor1[960];
    UnbiasedRNG[202] = LFSRcolor1[483];
    UnbiasedRNG[203] = LFSRcolor1[456];
    UnbiasedRNG[204] = LFSRcolor1[3];
    UnbiasedRNG[205] = LFSRcolor1[41];
    UnbiasedRNG[206] = LFSRcolor1[24];
    UnbiasedRNG[207] = LFSRcolor1[429];
    UnbiasedRNG[208] = LFSRcolor1[602];
    UnbiasedRNG[209] = LFSRcolor1[605];
    UnbiasedRNG[210] = LFSRcolor1[358];
    UnbiasedRNG[211] = LFSRcolor1[535];
    UnbiasedRNG[212] = LFSRcolor1[164];
    UnbiasedRNG[213] = LFSRcolor1[36];
    UnbiasedRNG[214] = LFSRcolor1[274];
    UnbiasedRNG[215] = LFSRcolor1[367];
    UnbiasedRNG[216] = LFSRcolor1[989];
    UnbiasedRNG[217] = LFSRcolor1[670];
    UnbiasedRNG[218] = LFSRcolor1[292];
    UnbiasedRNG[219] = LFSRcolor1[503];
    UnbiasedRNG[220] = LFSRcolor1[904];
    UnbiasedRNG[221] = LFSRcolor1[801];
    UnbiasedRNG[222] = LFSRcolor1[578];
    UnbiasedRNG[223] = LFSRcolor1[937];
    UnbiasedRNG[224] = LFSRcolor1[739];
    UnbiasedRNG[225] = LFSRcolor1[5];
    UnbiasedRNG[226] = LFSRcolor1[84];
    UnbiasedRNG[227] = LFSRcolor1[1009];
    UnbiasedRNG[228] = LFSRcolor1[581];
    UnbiasedRNG[229] = LFSRcolor1[270];
    UnbiasedRNG[230] = LFSRcolor1[200];
    UnbiasedRNG[231] = LFSRcolor1[836];
    UnbiasedRNG[232] = LFSRcolor1[254];
    UnbiasedRNG[233] = LFSRcolor1[995];
    UnbiasedRNG[234] = LFSRcolor1[433];
    UnbiasedRNG[235] = LFSRcolor1[469];
    UnbiasedRNG[236] = LFSRcolor1[426];
    UnbiasedRNG[237] = LFSRcolor1[365];
    UnbiasedRNG[238] = LFSRcolor1[259];
    UnbiasedRNG[239] = LFSRcolor1[1004];
    UnbiasedRNG[240] = LFSRcolor1[151];
    UnbiasedRNG[241] = LFSRcolor1[986];
    UnbiasedRNG[242] = LFSRcolor1[345];
    UnbiasedRNG[243] = LFSRcolor1[888];
    UnbiasedRNG[244] = LFSRcolor1[932];
    UnbiasedRNG[245] = LFSRcolor1[616];
    UnbiasedRNG[246] = LFSRcolor1[258];
    UnbiasedRNG[247] = LFSRcolor1[422];
    UnbiasedRNG[248] = LFSRcolor1[444];
    UnbiasedRNG[249] = LFSRcolor1[222];
    UnbiasedRNG[250] = LFSRcolor1[896];
    UnbiasedRNG[251] = LFSRcolor1[598];
end

always @(posedge color1_clk) begin
    BiasedRNG[383] = (LFSRcolor2[687]&LFSRcolor2[257]&LFSRcolor2[640]&LFSRcolor2[389]);
    BiasedRNG[384] = (LFSRcolor2[468]&LFSRcolor2[362]&LFSRcolor2[444]&LFSRcolor2[394]);
    BiasedRNG[385] = (LFSRcolor2[18]&LFSRcolor2[466]&LFSRcolor2[7]&LFSRcolor2[304]);
    BiasedRNG[386] = (LFSRcolor2[547]&LFSRcolor2[470]&LFSRcolor2[583]&LFSRcolor2[88]);
    BiasedRNG[387] = (LFSRcolor2[663]&LFSRcolor2[115]&LFSRcolor2[669]&LFSRcolor2[524]);
    BiasedRNG[388] = (LFSRcolor2[729]&LFSRcolor2[731]&LFSRcolor2[249]&LFSRcolor2[483]);
    BiasedRNG[389] = (LFSRcolor2[485]&LFSRcolor2[232]&LFSRcolor2[691]&LFSRcolor2[89]);
    BiasedRNG[390] = (LFSRcolor2[653]&LFSRcolor2[529]&LFSRcolor2[322]&LFSRcolor2[78]);
    BiasedRNG[391] = (LFSRcolor2[591]&LFSRcolor2[544]&LFSRcolor2[572]&LFSRcolor2[301]);
    BiasedRNG[392] = (LFSRcolor2[621]&LFSRcolor2[278]&LFSRcolor2[719]&LFSRcolor2[221]);
    BiasedRNG[393] = (LFSRcolor2[343]&LFSRcolor2[460]&LFSRcolor2[37]&LFSRcolor2[271]);
    BiasedRNG[394] = (LFSRcolor2[47]&LFSRcolor2[712]&LFSRcolor2[623]&LFSRcolor2[610]);
    BiasedRNG[395] = (LFSRcolor2[146]&LFSRcolor2[596]&LFSRcolor2[505]&LFSRcolor2[335]);
    BiasedRNG[396] = (LFSRcolor2[361]&LFSRcolor2[536]&LFSRcolor2[388]&LFSRcolor2[298]);
    BiasedRNG[397] = (LFSRcolor2[262]&LFSRcolor2[274]&LFSRcolor2[540]&LFSRcolor2[573]);
    BiasedRNG[398] = (LFSRcolor2[49]&LFSRcolor2[254]&LFSRcolor2[179]&LFSRcolor2[287]);
    BiasedRNG[399] = (LFSRcolor2[332]&LFSRcolor2[369]&LFSRcolor2[399]&LFSRcolor2[725]);
    BiasedRNG[400] = (LFSRcolor2[395]&LFSRcolor2[341]&LFSRcolor2[122]&LFSRcolor2[80]);
    BiasedRNG[401] = (LFSRcolor2[720]&LFSRcolor2[109]&LFSRcolor2[21]&LFSRcolor2[68]);
    BiasedRNG[402] = (LFSRcolor2[512]&LFSRcolor2[513]&LFSRcolor2[345]&LFSRcolor2[225]);
    BiasedRNG[403] = (LFSRcolor2[484]&LFSRcolor2[127]&LFSRcolor2[15]&LFSRcolor2[387]);
    BiasedRNG[404] = (LFSRcolor2[417]&LFSRcolor2[502]&LFSRcolor2[420]&LFSRcolor2[693]);
    BiasedRNG[405] = (LFSRcolor2[283]&LFSRcolor2[715]&LFSRcolor2[405]&LFSRcolor2[134]);
    BiasedRNG[406] = (LFSRcolor2[282]&LFSRcolor2[527]&LFSRcolor2[154]&LFSRcolor2[377]);
    BiasedRNG[407] = (LFSRcolor2[448]&LFSRcolor2[550]&LFSRcolor2[275]&LFSRcolor2[279]);
    BiasedRNG[408] = (LFSRcolor2[519]&LFSRcolor2[722]&LFSRcolor2[201]&LFSRcolor2[239]);
    BiasedRNG[409] = (LFSRcolor2[251]&LFSRcolor2[557]&LFSRcolor2[160]&LFSRcolor2[514]);
    BiasedRNG[410] = (LFSRcolor2[704]&LFSRcolor2[62]&LFSRcolor2[14]&LFSRcolor2[609]);
    BiasedRNG[411] = (LFSRcolor2[36]&LFSRcolor2[656]&LFSRcolor2[503]&LFSRcolor2[622]);
    BiasedRNG[412] = (LFSRcolor2[29]&LFSRcolor2[507]&LFSRcolor2[213]&LFSRcolor2[414]);
    BiasedRNG[413] = (LFSRcolor2[321]&LFSRcolor2[569]&LFSRcolor2[229]&LFSRcolor2[495]);
    BiasedRNG[414] = (LFSRcolor2[517]&LFSRcolor2[351]&LFSRcolor2[545]&LFSRcolor2[159]);
    BiasedRNG[415] = (LFSRcolor2[624]&LFSRcolor2[546]&LFSRcolor2[651]&LFSRcolor2[595]);
    BiasedRNG[416] = (LFSRcolor2[73]&LFSRcolor2[446]&LFSRcolor2[218]&LFSRcolor2[305]);
    BiasedRNG[417] = (LFSRcolor2[222]&LFSRcolor2[53]&LFSRcolor2[401]&LFSRcolor2[376]);
    BiasedRNG[418] = (LFSRcolor2[72]&LFSRcolor2[358]&LFSRcolor2[188]&LFSRcolor2[327]);
    BiasedRNG[419] = (LFSRcolor2[342]&LFSRcolor2[698]&LFSRcolor2[105]&LFSRcolor2[506]);
    BiasedRNG[420] = (LFSRcolor2[593]&LFSRcolor2[328]&LFSRcolor2[183]&LFSRcolor2[598]);
    BiasedRNG[421] = (LFSRcolor2[685]&LFSRcolor2[701]&LFSRcolor2[289]&LFSRcolor2[120]);
    BiasedRNG[422] = (LFSRcolor2[141]&LFSRcolor2[148]&LFSRcolor2[60]&LFSRcolor2[390]);
    BiasedRNG[423] = (LFSRcolor2[734]&LFSRcolor2[566]&LFSRcolor2[379]&LFSRcolor2[13]);
    BiasedRNG[424] = (LFSRcolor2[235]&LFSRcolor2[579]&LFSRcolor2[404]&LFSRcolor2[438]);
    BiasedRNG[425] = (LFSRcolor2[186]&LFSRcolor2[373]&LFSRcolor2[469]&LFSRcolor2[299]);
    BiasedRNG[426] = (LFSRcolor2[184]&LFSRcolor2[486]&LFSRcolor2[578]&LFSRcolor2[646]);
    BiasedRNG[427] = (LFSRcolor2[331]&LFSRcolor2[34]&LFSRcolor2[110]&LFSRcolor2[392]);
    BiasedRNG[428] = (LFSRcolor2[463]&LFSRcolor2[632]&LFSRcolor2[518]&LFSRcolor2[581]);
    BiasedRNG[429] = (LFSRcolor2[692]&LFSRcolor2[384]&LFSRcolor2[368]&LFSRcolor2[592]);
    BiasedRNG[430] = (LFSRcolor2[189]&LFSRcolor2[348]&LFSRcolor2[398]&LFSRcolor2[676]);
    BiasedRNG[431] = (LFSRcolor2[534]&LFSRcolor2[167]&LFSRcolor2[560]&LFSRcolor2[733]);
    BiasedRNG[432] = (LFSRcolor2[385]&LFSRcolor2[474]&LFSRcolor2[268]&LFSRcolor2[106]);
    BiasedRNG[433] = (LFSRcolor2[2]&LFSRcolor2[454]&LFSRcolor2[310]&LFSRcolor2[69]);
    BiasedRNG[434] = (LFSRcolor2[261]&LFSRcolor2[346]&LFSRcolor2[24]&LFSRcolor2[292]);
    BiasedRNG[435] = (LFSRcolor2[638]&LFSRcolor2[207]&LFSRcolor2[95]&LFSRcolor2[599]);
    BiasedRNG[436] = (LFSRcolor2[363]&LFSRcolor2[678]&LFSRcolor2[732]&LFSRcolor2[175]);
    BiasedRNG[437] = (LFSRcolor2[433]&LFSRcolor2[288]&LFSRcolor2[137]&LFSRcolor2[264]);
    BiasedRNG[438] = (LFSRcolor2[216]&LFSRcolor2[586]&LFSRcolor2[138]&LFSRcolor2[238]);
    BiasedRNG[439] = (LFSRcolor2[217]&LFSRcolor2[119]&LFSRcolor2[567]&LFSRcolor2[728]);
    BiasedRNG[440] = (LFSRcolor2[50]&LFSRcolor2[449]&LFSRcolor2[10]&LFSRcolor2[453]);
    BiasedRNG[441] = (LFSRcolor2[172]&LFSRcolor2[41]&LFSRcolor2[125]&LFSRcolor2[627]);
    BiasedRNG[442] = (LFSRcolor2[462]&LFSRcolor2[614]&LFSRcolor2[481]&LFSRcolor2[0]);
    BiasedRNG[443] = (LFSRcolor2[380]&LFSRcolor2[608]&LFSRcolor2[190]&LFSRcolor2[334]);
    BiasedRNG[444] = (LFSRcolor2[93]&LFSRcolor2[199]&LFSRcolor2[489]&LFSRcolor2[402]);
    BiasedRNG[445] = (LFSRcolor2[30]&LFSRcolor2[163]&LFSRcolor2[451]&LFSRcolor2[90]);
    BiasedRNG[446] = (LFSRcolor2[639]&LFSRcolor2[22]&LFSRcolor2[510]&LFSRcolor2[382]);
    BiasedRNG[447] = (LFSRcolor2[236]&LFSRcolor2[674]&LFSRcolor2[83]&LFSRcolor2[226]);
    BiasedRNG[448] = (LFSRcolor2[250]&LFSRcolor2[237]&LFSRcolor2[422]&LFSRcolor2[25]);
    BiasedRNG[449] = (LFSRcolor2[65]&LFSRcolor2[530]&LFSRcolor2[683]&LFSRcolor2[473]);
    BiasedRNG[450] = (LFSRcolor2[475]&LFSRcolor2[708]&LFSRcolor2[185]&LFSRcolor2[714]);
    BiasedRNG[451] = (LFSRcolor2[147]&LFSRcolor2[675]&LFSRcolor2[124]&LFSRcolor2[272]);
    BiasedRNG[452] = (LFSRcolor2[253]&LFSRcolor2[12]&LFSRcolor2[492]&LFSRcolor2[594]);
    BiasedRNG[453] = (LFSRcolor2[241]&LFSRcolor2[370]&LFSRcolor2[352]&LFSRcolor2[57]);
    BiasedRNG[454] = (LFSRcolor2[295]&LFSRcolor2[56]&LFSRcolor2[690]&LFSRcolor2[723]);
    BiasedRNG[455] = (LFSRcolor2[657]&LFSRcolor2[108]&LFSRcolor2[58]&LFSRcolor2[494]);
    BiasedRNG[456] = (LFSRcolor2[19]&LFSRcolor2[46]&LFSRcolor2[20]&LFSRcolor2[457]);
    BiasedRNG[457] = (LFSRcolor2[700]&LFSRcolor2[168]&LFSRcolor2[558]&LFSRcolor2[317]);
    BiasedRNG[458] = (LFSRcolor2[612]&LFSRcolor2[166]&LFSRcolor2[447]&LFSRcolor2[315]);
    BiasedRNG[459] = (LFSRcolor2[45]&LFSRcolor2[16]&LFSRcolor2[350]&LFSRcolor2[613]);
    BiasedRNG[460] = (LFSRcolor2[430]&LFSRcolor2[114]&LFSRcolor2[620]&LFSRcolor2[531]);
    BiasedRNG[461] = (LFSRcolor2[490]&LFSRcolor2[198]&LFSRcolor2[411]&LFSRcolor2[244]);
    BiasedRNG[462] = (LFSRcolor2[607]&LFSRcolor2[590]&LFSRcolor2[314]&LFSRcolor2[383]);
    BiasedRNG[463] = (LFSRcolor2[143]&LFSRcolor2[554]&LFSRcolor2[192]&LFSRcolor2[455]);
    BiasedRNG[464] = (LFSRcolor2[145]&LFSRcolor2[630]&LFSRcolor2[353]&LFSRcolor2[568]);
    BiasedRNG[465] = (LFSRcolor2[498]&LFSRcolor2[206]&LFSRcolor2[391]&LFSRcolor2[55]);
    BiasedRNG[466] = (LFSRcolor2[703]&LFSRcolor2[323]&LFSRcolor2[587]&LFSRcolor2[709]);
    BiasedRNG[467] = (LFSRcolor2[316]&LFSRcolor2[458]&LFSRcolor2[427]&LFSRcolor2[717]);
    BiasedRNG[468] = (LFSRcolor2[79]&LFSRcolor2[176]&LFSRcolor2[500]&LFSRcolor2[688]);
    BiasedRNG[469] = (LFSRcolor2[445]&LFSRcolor2[480]&LFSRcolor2[35]&LFSRcolor2[107]);
    BiasedRNG[470] = (LFSRcolor2[707]&LFSRcolor2[629]&LFSRcolor2[215]&LFSRcolor2[360]);
    BiasedRNG[471] = (LFSRcolor2[559]&LFSRcolor2[336]&LFSRcolor2[425]&LFSRcolor2[718]);
    BiasedRNG[472] = (LFSRcolor2[574]&LFSRcolor2[59]&LFSRcolor2[27]&LFSRcolor2[170]);
    BiasedRNG[473] = (LFSRcolor2[270]&LFSRcolor2[666]&LFSRcolor2[280]&LFSRcolor2[464]);
    BiasedRNG[474] = (LFSRcolor2[482]&LFSRcolor2[496]&LFSRcolor2[618]&LFSRcolor2[397]);
    BiasedRNG[475] = (LFSRcolor2[523]&LFSRcolor2[511]&LFSRcolor2[180]&LFSRcolor2[372]);
    BiasedRNG[476] = (LFSRcolor2[165]&LFSRcolor2[601]&LFSRcolor2[726]&LFSRcolor2[245]);
    BiasedRNG[477] = (LFSRcolor2[296]&LFSRcolor2[171]&LFSRcolor2[585]&LFSRcolor2[477]);
    BiasedRNG[478] = (LFSRcolor2[428]&LFSRcolor2[219]&LFSRcolor2[98]&LFSRcolor2[431]);
    BiasedRNG[479] = (LFSRcolor2[349]&LFSRcolor2[96]&LFSRcolor2[509]&LFSRcolor2[61]);
    BiasedRNG[480] = (LFSRcolor2[265]&LFSRcolor2[374]&LFSRcolor2[424]&LFSRcolor2[682]);
    BiasedRNG[481] = (LFSRcolor2[230]&LFSRcolor2[64]&LFSRcolor2[164]&LFSRcolor2[713]);
    BiasedRNG[482] = (LFSRcolor2[689]&LFSRcolor2[319]&LFSRcolor2[126]&LFSRcolor2[603]);
    BiasedRNG[483] = (LFSRcolor2[302]&LFSRcolor2[410]&LFSRcolor2[626]&LFSRcolor2[366]);
    BiasedRNG[484] = (LFSRcolor2[308]&LFSRcolor2[193]&LFSRcolor2[129]&LFSRcolor2[312]);
    BiasedRNG[485] = (LFSRcolor2[408]&LFSRcolor2[727]&LFSRcolor2[220]&LFSRcolor2[340]);
    BiasedRNG[486] = (LFSRcolor2[409]&LFSRcolor2[161]&LFSRcolor2[641]&LFSRcolor2[52]);
    BiasedRNG[487] = (LFSRcolor2[429]&LFSRcolor2[28]&LFSRcolor2[670]&LFSRcolor2[354]);
    BiasedRNG[488] = (LFSRcolor2[619]&LFSRcolor2[602]&LFSRcolor2[537]&LFSRcolor2[548]);
    BiasedRNG[489] = (LFSRcolor2[82]&LFSRcolor2[3]&LFSRcolor2[87]&LFSRcolor2[673]);
    BiasedRNG[490] = (LFSRcolor2[660]&LFSRcolor2[681]&LFSRcolor2[247]&LFSRcolor2[227]);
    BiasedRNG[491] = (LFSRcolor2[307]&LFSRcolor2[400]&LFSRcolor2[256]&LFSRcolor2[679]);
    BiasedRNG[492] = (LFSRcolor2[695]&LFSRcolor2[575]&LFSRcolor2[40]&LFSRcolor2[309]);
    BiasedRNG[493] = (LFSRcolor2[655]&LFSRcolor2[85]&LFSRcolor2[576]&LFSRcolor2[234]);
    BiasedRNG[494] = (LFSRcolor2[456]&LFSRcolor2[205]&LFSRcolor2[258]&LFSRcolor2[442]);
    BiasedRNG[495] = (LFSRcolor2[538]&LFSRcolor2[128]&LFSRcolor2[246]&LFSRcolor2[111]);
    BiasedRNG[496] = (LFSRcolor2[515]&LFSRcolor2[303]&LFSRcolor2[665]&LFSRcolor2[8]);
    BiasedRNG[497] = (LFSRcolor2[135]&LFSRcolor2[671]&LFSRcolor2[441]&LFSRcolor2[604]);
    BiasedRNG[498] = (LFSRcolor2[344]&LFSRcolor2[471]&LFSRcolor2[1]&LFSRcolor2[92]);
    BiasedRNG[499] = (LFSRcolor2[541]&LFSRcolor2[615]&LFSRcolor2[224]&LFSRcolor2[664]);
    BiasedRNG[500] = (LFSRcolor2[76]&LFSRcolor2[437]&LFSRcolor2[631]&LFSRcolor2[320]);
    BiasedRNG[501] = (LFSRcolor2[371]&LFSRcolor2[347]&LFSRcolor2[294]&LFSRcolor2[313]);
    BiasedRNG[502] = (LFSRcolor2[633]&LFSRcolor2[71]&LFSRcolor2[104]&LFSRcolor2[606]);
    BiasedRNG[503] = (LFSRcolor2[195]&LFSRcolor2[493]&LFSRcolor2[597]&LFSRcolor2[357]);
    BiasedRNG[504] = (LFSRcolor2[476]&LFSRcolor2[499]&LFSRcolor2[333]&LFSRcolor2[231]);
    BiasedRNG[505] = (LFSRcolor2[66]&LFSRcolor2[26]&LFSRcolor2[259]&LFSRcolor2[43]);
    BiasedRNG[506] = (LFSRcolor2[325]&LFSRcolor2[11]&LFSRcolor2[152]&LFSRcolor2[209]);
    BiasedRNG[507] = (LFSRcolor2[121]&LFSRcolor2[23]&LFSRcolor2[616]&LFSRcolor2[210]);
    BiasedRNG[508] = (LFSRcolor2[648]&LFSRcolor2[600]&LFSRcolor2[521]&LFSRcolor2[552]);
    BiasedRNG[509] = (LFSRcolor2[696]&LFSRcolor2[101]&LFSRcolor2[644]&LFSRcolor2[605]);
    BiasedRNG[510] = (LFSRcolor2[407]&LFSRcolor2[423]&LFSRcolor2[324]&LFSRcolor2[418]);
    BiasedRNG[511] = (LFSRcolor2[434]&LFSRcolor2[203]&LFSRcolor2[240]&LFSRcolor2[577]);
    BiasedRNG[512] = (LFSRcolor2[684]&LFSRcolor2[549]&LFSRcolor2[202]&LFSRcolor2[565]);
    BiasedRNG[513] = (LFSRcolor2[266]&LFSRcolor2[501]&LFSRcolor2[628]&LFSRcolor2[6]);
    BiasedRNG[514] = (LFSRcolor2[588]&LFSRcolor2[532]&LFSRcolor2[223]&LFSRcolor2[412]);
    BiasedRNG[515] = (LFSRcolor2[539]&LFSRcolor2[637]&LFSRcolor2[543]&LFSRcolor2[582]);
    BiasedRNG[516] = (LFSRcolor2[716]&LFSRcolor2[617]&LFSRcolor2[381]&LFSRcolor2[467]);
    BiasedRNG[517] = (LFSRcolor2[100]&LFSRcolor2[267]&LFSRcolor2[155]&LFSRcolor2[39]);
    BiasedRNG[518] = (LFSRcolor2[564]&LFSRcolor2[136]&LFSRcolor2[367]&LFSRcolor2[200]);
    BiasedRNG[519] = (LFSRcolor2[416]&LFSRcolor2[625]&LFSRcolor2[661]&LFSRcolor2[158]);
    BiasedRNG[520] = (LFSRcolor2[97]&LFSRcolor2[556]&LFSRcolor2[702]&LFSRcolor2[436]);
    BiasedRNG[521] = (LFSRcolor2[33]&LFSRcolor2[263]&LFSRcolor2[17]&LFSRcolor2[730]);
    BiasedRNG[522] = (LFSRcolor2[77]&LFSRcolor2[339]&LFSRcolor2[144]&LFSRcolor2[584]);
    BiasedRNG[523] = (LFSRcolor2[103]&LFSRcolor2[406]&LFSRcolor2[306]&LFSRcolor2[551]);
    BiasedRNG[524] = (LFSRcolor2[635]&LFSRcolor2[139]&LFSRcolor2[153]&LFSRcolor2[243]);
    BiasedRNG[525] = (LFSRcolor2[443]&LFSRcolor2[113]&LFSRcolor2[706]&LFSRcolor2[658]);
    BiasedRNG[526] = (LFSRcolor2[553]&LFSRcolor2[140]&LFSRcolor2[649]&LFSRcolor2[132]);
    UnbiasedRNG[252] = LFSRcolor2[580];
    UnbiasedRNG[253] = LFSRcolor2[130];
    UnbiasedRNG[254] = LFSRcolor2[735];
    UnbiasedRNG[255] = LFSRcolor2[214];
    UnbiasedRNG[256] = LFSRcolor2[461];
    UnbiasedRNG[257] = LFSRcolor2[705];
    UnbiasedRNG[258] = LFSRcolor2[432];
    UnbiasedRNG[259] = LFSRcolor2[94];
    UnbiasedRNG[260] = LFSRcolor2[149];
    UnbiasedRNG[261] = LFSRcolor2[291];
    UnbiasedRNG[262] = LFSRcolor2[162];
    UnbiasedRNG[263] = LFSRcolor2[277];
    UnbiasedRNG[264] = LFSRcolor2[74];
    UnbiasedRNG[265] = LFSRcolor2[326];
    UnbiasedRNG[266] = LFSRcolor2[285];
    UnbiasedRNG[267] = LFSRcolor2[208];
    UnbiasedRNG[268] = LFSRcolor2[636];
    UnbiasedRNG[269] = LFSRcolor2[355];
    UnbiasedRNG[270] = LFSRcolor2[450];
    UnbiasedRNG[271] = LFSRcolor2[415];
    UnbiasedRNG[272] = LFSRcolor2[652];
    UnbiasedRNG[273] = LFSRcolor2[570];
    UnbiasedRNG[274] = LFSRcolor2[150];
    UnbiasedRNG[275] = LFSRcolor2[38];
    UnbiasedRNG[276] = LFSRcolor2[131];
    UnbiasedRNG[277] = LFSRcolor2[99];
    UnbiasedRNG[278] = LFSRcolor2[365];
    UnbiasedRNG[279] = LFSRcolor2[102];
    UnbiasedRNG[280] = LFSRcolor2[504];
    UnbiasedRNG[281] = LFSRcolor2[194];
    UnbiasedRNG[282] = LFSRcolor2[290];
    UnbiasedRNG[283] = LFSRcolor2[421];
    UnbiasedRNG[284] = LFSRcolor2[459];
    UnbiasedRNG[285] = LFSRcolor2[522];
    UnbiasedRNG[286] = LFSRcolor2[710];
    UnbiasedRNG[287] = LFSRcolor2[44];
    UnbiasedRNG[288] = LFSRcolor2[276];
    UnbiasedRNG[289] = LFSRcolor2[465];
    UnbiasedRNG[290] = LFSRcolor2[157];
    UnbiasedRNG[291] = LFSRcolor2[711];
    UnbiasedRNG[292] = LFSRcolor2[211];
    UnbiasedRNG[293] = LFSRcolor2[31];
    UnbiasedRNG[294] = LFSRcolor2[284];
    UnbiasedRNG[295] = LFSRcolor2[123];
    UnbiasedRNG[296] = LFSRcolor2[252];
    UnbiasedRNG[297] = LFSRcolor2[356];
    UnbiasedRNG[298] = LFSRcolor2[571];
    UnbiasedRNG[299] = LFSRcolor2[174];
    UnbiasedRNG[300] = LFSRcolor2[497];
    UnbiasedRNG[301] = LFSRcolor2[699];
    UnbiasedRNG[302] = LFSRcolor2[488];
    UnbiasedRNG[303] = LFSRcolor2[668];
    UnbiasedRNG[304] = LFSRcolor2[338];
    UnbiasedRNG[305] = LFSRcolor2[151];
    UnbiasedRNG[306] = LFSRcolor2[386];
    UnbiasedRNG[307] = LFSRcolor2[4];
    UnbiasedRNG[308] = LFSRcolor2[330];
    UnbiasedRNG[309] = LFSRcolor2[142];
    UnbiasedRNG[310] = LFSRcolor2[112];
    UnbiasedRNG[311] = LFSRcolor2[403];
    UnbiasedRNG[312] = LFSRcolor2[75];
    UnbiasedRNG[313] = LFSRcolor2[228];
    UnbiasedRNG[314] = LFSRcolor2[589];
    UnbiasedRNG[315] = LFSRcolor2[659];
    UnbiasedRNG[316] = LFSRcolor2[694];
    UnbiasedRNG[317] = LFSRcolor2[187];
    UnbiasedRNG[318] = LFSRcolor2[260];
    UnbiasedRNG[319] = LFSRcolor2[178];
    UnbiasedRNG[320] = LFSRcolor2[440];
    UnbiasedRNG[321] = LFSRcolor2[542];
    UnbiasedRNG[322] = LFSRcolor2[478];
    UnbiasedRNG[323] = LFSRcolor2[182];
    UnbiasedRNG[324] = LFSRcolor2[269];
    UnbiasedRNG[325] = LFSRcolor2[197];
    UnbiasedRNG[326] = LFSRcolor2[196];
    UnbiasedRNG[327] = LFSRcolor2[70];
    UnbiasedRNG[328] = LFSRcolor2[535];
    UnbiasedRNG[329] = LFSRcolor2[117];
    UnbiasedRNG[330] = LFSRcolor2[48];
    UnbiasedRNG[331] = LFSRcolor2[32];
    UnbiasedRNG[332] = LFSRcolor2[212];
    UnbiasedRNG[333] = LFSRcolor2[611];
    UnbiasedRNG[334] = LFSRcolor2[645];
    UnbiasedRNG[335] = LFSRcolor2[318];
    UnbiasedRNG[336] = LFSRcolor2[364];
    UnbiasedRNG[337] = LFSRcolor2[525];
    UnbiasedRNG[338] = LFSRcolor2[91];
    UnbiasedRNG[339] = LFSRcolor2[281];
    UnbiasedRNG[340] = LFSRcolor2[248];
    UnbiasedRNG[341] = LFSRcolor2[156];
    UnbiasedRNG[342] = LFSRcolor2[5];
    UnbiasedRNG[343] = LFSRcolor2[84];
    UnbiasedRNG[344] = LFSRcolor2[516];
    UnbiasedRNG[345] = LFSRcolor2[311];
    UnbiasedRNG[346] = LFSRcolor2[472];
    UnbiasedRNG[347] = LFSRcolor2[520];
    UnbiasedRNG[348] = LFSRcolor2[359];
    UnbiasedRNG[349] = LFSRcolor2[233];
    UnbiasedRNG[350] = LFSRcolor2[9];
    UnbiasedRNG[351] = LFSRcolor2[378];
    UnbiasedRNG[352] = LFSRcolor2[491];
    UnbiasedRNG[353] = LFSRcolor2[393];
    UnbiasedRNG[354] = LFSRcolor2[533];
    UnbiasedRNG[355] = LFSRcolor2[396];
    UnbiasedRNG[356] = LFSRcolor2[118];
    UnbiasedRNG[357] = LFSRcolor2[562];
    UnbiasedRNG[358] = LFSRcolor2[286];
    UnbiasedRNG[359] = LFSRcolor2[555];
    UnbiasedRNG[360] = LFSRcolor2[300];
    UnbiasedRNG[361] = LFSRcolor2[528];
    UnbiasedRNG[362] = LFSRcolor2[654];
    UnbiasedRNG[363] = LFSRcolor2[721];
    UnbiasedRNG[364] = LFSRcolor2[329];
    UnbiasedRNG[365] = LFSRcolor2[561];
    UnbiasedRNG[366] = LFSRcolor2[487];
    UnbiasedRNG[367] = LFSRcolor2[204];
    UnbiasedRNG[368] = LFSRcolor2[563];
    UnbiasedRNG[369] = LFSRcolor2[435];
    UnbiasedRNG[370] = LFSRcolor2[173];
    UnbiasedRNG[371] = LFSRcolor2[634];
    UnbiasedRNG[372] = LFSRcolor2[686];
    UnbiasedRNG[373] = LFSRcolor2[375];
    UnbiasedRNG[374] = LFSRcolor2[647];
    UnbiasedRNG[375] = LFSRcolor2[242];
    UnbiasedRNG[376] = LFSRcolor2[667];
    UnbiasedRNG[377] = LFSRcolor2[439];
    UnbiasedRNG[378] = LFSRcolor2[116];
    UnbiasedRNG[379] = LFSRcolor2[337];
    UnbiasedRNG[380] = LFSRcolor2[643];
    UnbiasedRNG[381] = LFSRcolor2[724];
    UnbiasedRNG[382] = LFSRcolor2[181];
    UnbiasedRNG[383] = LFSRcolor2[650];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[384] = LFSRcolor3[24];
    UnbiasedRNG[385] = LFSRcolor3[47];
    UnbiasedRNG[386] = LFSRcolor3[53];
    UnbiasedRNG[387] = LFSRcolor3[58];
    UnbiasedRNG[388] = LFSRcolor3[67];
    UnbiasedRNG[389] = LFSRcolor3[86];
    UnbiasedRNG[390] = LFSRcolor3[84];
    UnbiasedRNG[391] = LFSRcolor3[79];
    UnbiasedRNG[392] = LFSRcolor3[132];
    UnbiasedRNG[393] = LFSRcolor3[117];
    UnbiasedRNG[394] = LFSRcolor3[80];
    UnbiasedRNG[395] = LFSRcolor3[90];
    UnbiasedRNG[396] = LFSRcolor3[66];
    UnbiasedRNG[397] = LFSRcolor3[61];
    UnbiasedRNG[398] = LFSRcolor3[129];
    UnbiasedRNG[399] = LFSRcolor3[63];
    UnbiasedRNG[400] = LFSRcolor3[20];
    UnbiasedRNG[401] = LFSRcolor3[38];
    UnbiasedRNG[402] = LFSRcolor3[78];
    UnbiasedRNG[403] = LFSRcolor3[121];
    UnbiasedRNG[404] = LFSRcolor3[21];
    UnbiasedRNG[405] = LFSRcolor3[88];
    UnbiasedRNG[406] = LFSRcolor3[16];
    UnbiasedRNG[407] = LFSRcolor3[124];
    UnbiasedRNG[408] = LFSRcolor3[87];
    UnbiasedRNG[409] = LFSRcolor3[59];
    UnbiasedRNG[410] = LFSRcolor3[92];
    UnbiasedRNG[411] = LFSRcolor3[11];
    UnbiasedRNG[412] = LFSRcolor3[39];
    UnbiasedRNG[413] = LFSRcolor3[33];
    UnbiasedRNG[414] = LFSRcolor3[54];
    UnbiasedRNG[415] = LFSRcolor3[70];
    UnbiasedRNG[416] = LFSRcolor3[85];
    UnbiasedRNG[417] = LFSRcolor3[49];
    UnbiasedRNG[418] = LFSRcolor3[97];
    UnbiasedRNG[419] = LFSRcolor3[30];
    UnbiasedRNG[420] = LFSRcolor3[13];
    UnbiasedRNG[421] = LFSRcolor3[62];
    UnbiasedRNG[422] = LFSRcolor3[116];
    UnbiasedRNG[423] = LFSRcolor3[114];
    UnbiasedRNG[424] = LFSRcolor3[8];
    UnbiasedRNG[425] = LFSRcolor3[89];
    UnbiasedRNG[426] = LFSRcolor3[37];
    UnbiasedRNG[427] = LFSRcolor3[73];
    UnbiasedRNG[428] = LFSRcolor3[130];
    UnbiasedRNG[429] = LFSRcolor3[125];
    UnbiasedRNG[430] = LFSRcolor3[109];
    UnbiasedRNG[431] = LFSRcolor3[95];
    UnbiasedRNG[432] = LFSRcolor3[17];
    UnbiasedRNG[433] = LFSRcolor3[94];
    UnbiasedRNG[434] = LFSRcolor3[56];
    UnbiasedRNG[435] = LFSRcolor3[6];
    UnbiasedRNG[436] = LFSRcolor3[55];
    UnbiasedRNG[437] = LFSRcolor3[101];
    UnbiasedRNG[438] = LFSRcolor3[43];
    UnbiasedRNG[439] = LFSRcolor3[118];
    UnbiasedRNG[440] = LFSRcolor3[10];
    UnbiasedRNG[441] = LFSRcolor3[83];
    UnbiasedRNG[442] = LFSRcolor3[60];
    UnbiasedRNG[443] = LFSRcolor3[122];
    UnbiasedRNG[444] = LFSRcolor3[9];
    UnbiasedRNG[445] = LFSRcolor3[71];
    UnbiasedRNG[446] = LFSRcolor3[34];
    UnbiasedRNG[447] = LFSRcolor3[110];
    UnbiasedRNG[448] = LFSRcolor3[15];
    UnbiasedRNG[449] = LFSRcolor3[127];
    UnbiasedRNG[450] = LFSRcolor3[131];
    UnbiasedRNG[451] = LFSRcolor3[137];
    UnbiasedRNG[452] = LFSRcolor3[36];
    UnbiasedRNG[453] = LFSRcolor3[72];
    UnbiasedRNG[454] = LFSRcolor3[100];
    UnbiasedRNG[455] = LFSRcolor3[112];
    UnbiasedRNG[456] = LFSRcolor3[104];
    UnbiasedRNG[457] = LFSRcolor3[7];
    UnbiasedRNG[458] = LFSRcolor3[102];
    UnbiasedRNG[459] = LFSRcolor3[76];
    UnbiasedRNG[460] = LFSRcolor3[111];
    UnbiasedRNG[461] = LFSRcolor3[29];
    UnbiasedRNG[462] = LFSRcolor3[32];
    UnbiasedRNG[463] = LFSRcolor3[133];
    UnbiasedRNG[464] = LFSRcolor3[51];
    UnbiasedRNG[465] = LFSRcolor3[12];
    UnbiasedRNG[466] = LFSRcolor3[107];
    UnbiasedRNG[467] = LFSRcolor3[40];
    UnbiasedRNG[468] = LFSRcolor3[135];
    UnbiasedRNG[469] = LFSRcolor3[98];
    UnbiasedRNG[470] = LFSRcolor3[81];
    UnbiasedRNG[471] = LFSRcolor3[68];
    UnbiasedRNG[472] = LFSRcolor3[113];
    UnbiasedRNG[473] = LFSRcolor3[57];
    UnbiasedRNG[474] = LFSRcolor3[123];
    UnbiasedRNG[475] = LFSRcolor3[77];
    UnbiasedRNG[476] = LFSRcolor3[74];
    UnbiasedRNG[477] = LFSRcolor3[65];
    UnbiasedRNG[478] = LFSRcolor3[0];
    UnbiasedRNG[479] = LFSRcolor3[31];
    UnbiasedRNG[480] = LFSRcolor3[64];
    UnbiasedRNG[481] = LFSRcolor3[22];
    UnbiasedRNG[482] = LFSRcolor3[18];
    UnbiasedRNG[483] = LFSRcolor3[3];
    UnbiasedRNG[484] = LFSRcolor3[4];
    UnbiasedRNG[485] = LFSRcolor3[28];
    UnbiasedRNG[486] = LFSRcolor3[126];
    UnbiasedRNG[487] = LFSRcolor3[120];
    UnbiasedRNG[488] = LFSRcolor3[106];
    UnbiasedRNG[489] = LFSRcolor3[75];
    UnbiasedRNG[490] = LFSRcolor3[108];
    UnbiasedRNG[491] = LFSRcolor3[23];
    UnbiasedRNG[492] = LFSRcolor3[25];
    UnbiasedRNG[493] = LFSRcolor3[69];
end

always @(posedge color3_clk) begin
    BiasedRNG[527] = (LFSRcolor4[315]&LFSRcolor4[381]&LFSRcolor4[86]&LFSRcolor4[179]);
    BiasedRNG[528] = (LFSRcolor4[438]&LFSRcolor4[134]&LFSRcolor4[121]&LFSRcolor4[255]);
    BiasedRNG[529] = (LFSRcolor4[73]&LFSRcolor4[378]&LFSRcolor4[480]&LFSRcolor4[372]);
    BiasedRNG[530] = (LFSRcolor4[403]&LFSRcolor4[549]&LFSRcolor4[230]&LFSRcolor4[478]);
    BiasedRNG[531] = (LFSRcolor4[495]&LFSRcolor4[289]&LFSRcolor4[368]&LFSRcolor4[504]);
    BiasedRNG[532] = (LFSRcolor4[456]&LFSRcolor4[386]&LFSRcolor4[226]&LFSRcolor4[200]);
    BiasedRNG[533] = (LFSRcolor4[419]&LFSRcolor4[461]&LFSRcolor4[281]&LFSRcolor4[514]);
    BiasedRNG[534] = (LFSRcolor4[95]&LFSRcolor4[135]&LFSRcolor4[380]&LFSRcolor4[435]);
    BiasedRNG[535] = (LFSRcolor4[307]&LFSRcolor4[327]&LFSRcolor4[223]&LFSRcolor4[191]);
    BiasedRNG[536] = (LFSRcolor4[244]&LFSRcolor4[228]&LFSRcolor4[36]&LFSRcolor4[241]);
    BiasedRNG[537] = (LFSRcolor4[9]&LFSRcolor4[334]&LFSRcolor4[11]&LFSRcolor4[515]);
    BiasedRNG[538] = (LFSRcolor4[526]&LFSRcolor4[274]&LFSRcolor4[321]&LFSRcolor4[217]);
    BiasedRNG[539] = (LFSRcolor4[489]&LFSRcolor4[306]&LFSRcolor4[220]&LFSRcolor4[261]);
    BiasedRNG[540] = (LFSRcolor4[376]&LFSRcolor4[311]&LFSRcolor4[172]&LFSRcolor4[117]);
    BiasedRNG[541] = (LFSRcolor4[264]&LFSRcolor4[488]&LFSRcolor4[151]&LFSRcolor4[432]);
    BiasedRNG[542] = (LFSRcolor4[523]&LFSRcolor4[115]&LFSRcolor4[490]&LFSRcolor4[104]);
    BiasedRNG[543] = (LFSRcolor4[393]&LFSRcolor4[347]&LFSRcolor4[519]&LFSRcolor4[229]);
    BiasedRNG[544] = (LFSRcolor4[145]&LFSRcolor4[340]&LFSRcolor4[253]&LFSRcolor4[87]);
    BiasedRNG[545] = (LFSRcolor4[149]&LFSRcolor4[80]&LFSRcolor4[518]&LFSRcolor4[85]);
    BiasedRNG[546] = (LFSRcolor4[90]&LFSRcolor4[257]&LFSRcolor4[502]&LFSRcolor4[328]);
    BiasedRNG[547] = (LFSRcolor4[129]&LFSRcolor4[444]&LFSRcolor4[28]&LFSRcolor4[47]);
    BiasedRNG[548] = (LFSRcolor4[152]&LFSRcolor4[430]&LFSRcolor4[199]&LFSRcolor4[537]);
    BiasedRNG[549] = (LFSRcolor4[18]&LFSRcolor4[467]&LFSRcolor4[455]&LFSRcolor4[351]);
    BiasedRNG[550] = (LFSRcolor4[12]&LFSRcolor4[57]&LFSRcolor4[81]&LFSRcolor4[114]);
    BiasedRNG[551] = (LFSRcolor4[123]&LFSRcolor4[130]&LFSRcolor4[548]&LFSRcolor4[99]);
    BiasedRNG[552] = (LFSRcolor4[431]&LFSRcolor4[182]&LFSRcolor4[366]&LFSRcolor4[63]);
    BiasedRNG[553] = (LFSRcolor4[450]&LFSRcolor4[337]&LFSRcolor4[269]&LFSRcolor4[240]);
    BiasedRNG[554] = (LFSRcolor4[24]&LFSRcolor4[43]&LFSRcolor4[246]&LFSRcolor4[379]);
    BiasedRNG[555] = (LFSRcolor4[391]&LFSRcolor4[541]&LFSRcolor4[292]&LFSRcolor4[4]);
    BiasedRNG[556] = (LFSRcolor4[466]&LFSRcolor4[139]&LFSRcolor4[109]&LFSRcolor4[155]);
    BiasedRNG[557] = (LFSRcolor4[493]&LFSRcolor4[446]&LFSRcolor4[338]&LFSRcolor4[184]);
    BiasedRNG[558] = (LFSRcolor4[396]&LFSRcolor4[300]&LFSRcolor4[440]&LFSRcolor4[325]);
    BiasedRNG[559] = (LFSRcolor4[454]&LFSRcolor4[336]&LFSRcolor4[205]&LFSRcolor4[89]);
    BiasedRNG[560] = (LFSRcolor4[165]&LFSRcolor4[206]&LFSRcolor4[163]&LFSRcolor4[245]);
    BiasedRNG[561] = (LFSRcolor4[288]&LFSRcolor4[210]&LFSRcolor4[40]&LFSRcolor4[276]);
    BiasedRNG[562] = (LFSRcolor4[160]&LFSRcolor4[247]&LFSRcolor4[237]&LFSRcolor4[124]);
    BiasedRNG[563] = (LFSRcolor4[355]&LFSRcolor4[5]&LFSRcolor4[439]&LFSRcolor4[271]);
    BiasedRNG[564] = (LFSRcolor4[437]&LFSRcolor4[293]&LFSRcolor4[481]&LFSRcolor4[539]);
    BiasedRNG[565] = (LFSRcolor4[428]&LFSRcolor4[322]&LFSRcolor4[512]&LFSRcolor4[301]);
    BiasedRNG[566] = (LFSRcolor4[74]&LFSRcolor4[256]&LFSRcolor4[103]&LFSRcolor4[75]);
    BiasedRNG[567] = (LFSRcolor4[522]&LFSRcolor4[285]&LFSRcolor4[547]&LFSRcolor4[98]);
    BiasedRNG[568] = (LFSRcolor4[542]&LFSRcolor4[61]&LFSRcolor4[38]&LFSRcolor4[110]);
    BiasedRNG[569] = (LFSRcolor4[303]&LFSRcolor4[330]&LFSRcolor4[318]&LFSRcolor4[116]);
    BiasedRNG[570] = (LFSRcolor4[387]&LFSRcolor4[362]&LFSRcolor4[320]&LFSRcolor4[411]);
    BiasedRNG[571] = (LFSRcolor4[383]&LFSRcolor4[350]&LFSRcolor4[23]&LFSRcolor4[279]);
    BiasedRNG[572] = (LFSRcolor4[180]&LFSRcolor4[166]&LFSRcolor4[389]&LFSRcolor4[238]);
    BiasedRNG[573] = (LFSRcolor4[239]&LFSRcolor4[232]&LFSRcolor4[453]&LFSRcolor4[55]);
    BiasedRNG[574] = (LFSRcolor4[176]&LFSRcolor4[187]&LFSRcolor4[272]&LFSRcolor4[249]);
    BiasedRNG[575] = (LFSRcolor4[529]&LFSRcolor4[499]&LFSRcolor4[221]&LFSRcolor4[308]);
    BiasedRNG[576] = (LFSRcolor4[359]&LFSRcolor4[390]&LFSRcolor4[234]&LFSRcolor4[305]);
    BiasedRNG[577] = (LFSRcolor4[349]&LFSRcolor4[445]&LFSRcolor4[296]&LFSRcolor4[120]);
    BiasedRNG[578] = (LFSRcolor4[452]&LFSRcolor4[26]&LFSRcolor4[544]&LFSRcolor4[510]);
    BiasedRNG[579] = (LFSRcolor4[105]&LFSRcolor4[302]&LFSRcolor4[363]&LFSRcolor4[270]);
    BiasedRNG[580] = (LFSRcolor4[100]&LFSRcolor4[106]&LFSRcolor4[500]&LFSRcolor4[10]);
    BiasedRNG[581] = (LFSRcolor4[319]&LFSRcolor4[209]&LFSRcolor4[339]&LFSRcolor4[97]);
    BiasedRNG[582] = (LFSRcolor4[375]&LFSRcolor4[146]&LFSRcolor4[516]&LFSRcolor4[398]);
    BiasedRNG[583] = (LFSRcolor4[231]&LFSRcolor4[496]&LFSRcolor4[314]&LFSRcolor4[344]);
    BiasedRNG[584] = (LFSRcolor4[233]&LFSRcolor4[15]&LFSRcolor4[304]&LFSRcolor4[227]);
    BiasedRNG[585] = (LFSRcolor4[400]&LFSRcolor4[528]&LFSRcolor4[41]&LFSRcolor4[298]);
    BiasedRNG[586] = (LFSRcolor4[33]&LFSRcolor4[243]&LFSRcolor4[345]&LFSRcolor4[25]);
    BiasedRNG[587] = (LFSRcolor4[51]&LFSRcolor4[62]&LFSRcolor4[125]&LFSRcolor4[513]);
    BiasedRNG[588] = (LFSRcolor4[260]&LFSRcolor4[458]&LFSRcolor4[35]&LFSRcolor4[353]);
    BiasedRNG[589] = (LFSRcolor4[189]&LFSRcolor4[472]&LFSRcolor4[13]&LFSRcolor4[477]);
    BiasedRNG[590] = (LFSRcolor4[72]&LFSRcolor4[471]&LFSRcolor4[408]&LFSRcolor4[364]);
    BiasedRNG[591] = (LFSRcolor4[164]&LFSRcolor4[201]&LFSRcolor4[282]&LFSRcolor4[6]);
    BiasedRNG[592] = (LFSRcolor4[333]&LFSRcolor4[39]&LFSRcolor4[20]&LFSRcolor4[262]);
    BiasedRNG[593] = (LFSRcolor4[317]&LFSRcolor4[460]&LFSRcolor4[69]&LFSRcolor4[384]);
    BiasedRNG[594] = (LFSRcolor4[422]&LFSRcolor4[434]&LFSRcolor4[31]&LFSRcolor4[170]);
    BiasedRNG[595] = (LFSRcolor4[491]&LFSRcolor4[49]&LFSRcolor4[235]&LFSRcolor4[204]);
    BiasedRNG[596] = (LFSRcolor4[132]&LFSRcolor4[348]&LFSRcolor4[1]&LFSRcolor4[248]);
    BiasedRNG[597] = (LFSRcolor4[53]&LFSRcolor4[113]&LFSRcolor4[331]&LFSRcolor4[148]);
    BiasedRNG[598] = (LFSRcolor4[476]&LFSRcolor4[520]&LFSRcolor4[420]&LFSRcolor4[326]);
    BiasedRNG[599] = (LFSRcolor4[259]&LFSRcolor4[533]&LFSRcolor4[50]&LFSRcolor4[154]);
    BiasedRNG[600] = (LFSRcolor4[250]&LFSRcolor4[413]&LFSRcolor4[190]&LFSRcolor4[147]);
    BiasedRNG[601] = (LFSRcolor4[162]&LFSRcolor4[225]&LFSRcolor4[354]&LFSRcolor4[212]);
    BiasedRNG[602] = (LFSRcolor4[425]&LFSRcolor4[291]&LFSRcolor4[37]&LFSRcolor4[102]);
    BiasedRNG[603] = (LFSRcolor4[59]&LFSRcolor4[8]&LFSRcolor4[268]&LFSRcolor4[335]);
    BiasedRNG[604] = (LFSRcolor4[183]&LFSRcolor4[214]&LFSRcolor4[483]&LFSRcolor4[3]);
    BiasedRNG[605] = (LFSRcolor4[297]&LFSRcolor4[96]&LFSRcolor4[382]&LFSRcolor4[527]);
    BiasedRNG[606] = (LFSRcolor4[169]&LFSRcolor4[409]&LFSRcolor4[361]&LFSRcolor4[508]);
    BiasedRNG[607] = (LFSRcolor4[505]&LFSRcolor4[136]&LFSRcolor4[76]&LFSRcolor4[545]);
    BiasedRNG[608] = (LFSRcolor4[436]&LFSRcolor4[119]&LFSRcolor4[356]&LFSRcolor4[93]);
    BiasedRNG[609] = (LFSRcolor4[392]&LFSRcolor4[524]&LFSRcolor4[46]&LFSRcolor4[459]);
    BiasedRNG[610] = (LFSRcolor4[58]&LFSRcolor4[198]&LFSRcolor4[222]&LFSRcolor4[138]);
    BiasedRNG[611] = (LFSRcolor4[91]&LFSRcolor4[373]&LFSRcolor4[468]&LFSRcolor4[507]);
    BiasedRNG[612] = (LFSRcolor4[211]&LFSRcolor4[429]&LFSRcolor4[126]&LFSRcolor4[487]);
    BiasedRNG[613] = (LFSRcolor4[342]&LFSRcolor4[194]&LFSRcolor4[112]&LFSRcolor4[27]);
    BiasedRNG[614] = (LFSRcolor4[290]&LFSRcolor4[142]&LFSRcolor4[143]&LFSRcolor4[192]);
    BiasedRNG[615] = (LFSRcolor4[405]&LFSRcolor4[399]&LFSRcolor4[341]&LFSRcolor4[70]);
    BiasedRNG[616] = (LFSRcolor4[309]&LFSRcolor4[60]&LFSRcolor4[406]&LFSRcolor4[484]);
    BiasedRNG[617] = (LFSRcolor4[543]&LFSRcolor4[7]&LFSRcolor4[67]&LFSRcolor4[216]);
    BiasedRNG[618] = (LFSRcolor4[343]&LFSRcolor4[423]&LFSRcolor4[42]&LFSRcolor4[178]);
    BiasedRNG[619] = (LFSRcolor4[407]&LFSRcolor4[118]&LFSRcolor4[153]&LFSRcolor4[127]);
    BiasedRNG[620] = (LFSRcolor4[498]&LFSRcolor4[202]&LFSRcolor4[538]&LFSRcolor4[157]);
    BiasedRNG[621] = (LFSRcolor4[394]&LFSRcolor4[492]&LFSRcolor4[218]&LFSRcolor4[174]);
    BiasedRNG[622] = (LFSRcolor4[357]&LFSRcolor4[32]&LFSRcolor4[365]&LFSRcolor4[417]);
    BiasedRNG[623] = (LFSRcolor4[224]&LFSRcolor4[287]&LFSRcolor4[48]&LFSRcolor4[457]);
    BiasedRNG[624] = (LFSRcolor4[286]&LFSRcolor4[208]&LFSRcolor4[448]&LFSRcolor4[283]);
    BiasedRNG[625] = (LFSRcolor4[128]&LFSRcolor4[82]&LFSRcolor4[203]&LFSRcolor4[280]);
    BiasedRNG[626] = (LFSRcolor4[275]&LFSRcolor4[385]&LFSRcolor4[509]&LFSRcolor4[273]);
    BiasedRNG[627] = (LFSRcolor4[265]&LFSRcolor4[486]&LFSRcolor4[517]&LFSRcolor4[316]);
    BiasedRNG[628] = (LFSRcolor4[52]&LFSRcolor4[441]&LFSRcolor4[137]&LFSRcolor4[150]);
    BiasedRNG[629] = (LFSRcolor4[371]&LFSRcolor4[2]&LFSRcolor4[482]&LFSRcolor4[101]);
    BiasedRNG[630] = (LFSRcolor4[140]&LFSRcolor4[94]&LFSRcolor4[479]&LFSRcolor4[107]);
    BiasedRNG[631] = (LFSRcolor4[277]&LFSRcolor4[158]&LFSRcolor4[108]&LFSRcolor4[219]);
    BiasedRNG[632] = (LFSRcolor4[401]&LFSRcolor4[294]&LFSRcolor4[177]&LFSRcolor4[16]);
    BiasedRNG[633] = (LFSRcolor4[535]&LFSRcolor4[474]&LFSRcolor4[195]&LFSRcolor4[71]);
    BiasedRNG[634] = (LFSRcolor4[278]&LFSRcolor4[83]&LFSRcolor4[186]&LFSRcolor4[323]);
    BiasedRNG[635] = (LFSRcolor4[242]&LFSRcolor4[530]&LFSRcolor4[254]&LFSRcolor4[284]);
    BiasedRNG[636] = (LFSRcolor4[196]&LFSRcolor4[133]&LFSRcolor4[92]&LFSRcolor4[131]);
    BiasedRNG[637] = (LFSRcolor4[410]&LFSRcolor4[144]&LFSRcolor4[370]&LFSRcolor4[171]);
    BiasedRNG[638] = (LFSRcolor4[213]&LFSRcolor4[45]&LFSRcolor4[84]&LFSRcolor4[426]);
    BiasedRNG[639] = (LFSRcolor4[402]&LFSRcolor4[68]&LFSRcolor4[193]&LFSRcolor4[421]);
    BiasedRNG[640] = (LFSRcolor4[346]&LFSRcolor4[44]&LFSRcolor4[473]&LFSRcolor4[540]);
    BiasedRNG[641] = (LFSRcolor4[332]&LFSRcolor4[197]&LFSRcolor4[464]&LFSRcolor4[159]);
    BiasedRNG[642] = (LFSRcolor4[310]&LFSRcolor4[21]&LFSRcolor4[251]&LFSRcolor4[451]);
    BiasedRNG[643] = (LFSRcolor4[536]&LFSRcolor4[470]&LFSRcolor4[207]&LFSRcolor4[22]);
    BiasedRNG[644] = (LFSRcolor4[122]&LFSRcolor4[497]&LFSRcolor4[433]&LFSRcolor4[14]);
    BiasedRNG[645] = (LFSRcolor4[551]&LFSRcolor4[449]&LFSRcolor4[374]&LFSRcolor4[377]);
    BiasedRNG[646] = (LFSRcolor4[29]&LFSRcolor4[56]&LFSRcolor4[531]&LFSRcolor4[78]);
    BiasedRNG[647] = (LFSRcolor4[427]&LFSRcolor4[65]&LFSRcolor4[188]&LFSRcolor4[447]);
    BiasedRNG[648] = (LFSRcolor4[181]&LFSRcolor4[534]&LFSRcolor4[503]&LFSRcolor4[79]);
    BiasedRNG[649] = (LFSRcolor4[485]&LFSRcolor4[173]&LFSRcolor4[532]&LFSRcolor4[267]);
    BiasedRNG[650] = (LFSRcolor4[324]&LFSRcolor4[329]&LFSRcolor4[521]&LFSRcolor4[0]);
    BiasedRNG[651] = (LFSRcolor4[550]&LFSRcolor4[506]&LFSRcolor4[358]&LFSRcolor4[367]);
    BiasedRNG[652] = (LFSRcolor4[295]&LFSRcolor4[215]&LFSRcolor4[352]&LFSRcolor4[175]);
    BiasedRNG[653] = (LFSRcolor4[369]&LFSRcolor4[19]&LFSRcolor4[111]&LFSRcolor4[185]);
    BiasedRNG[654] = (LFSRcolor4[236]&LFSRcolor4[418]&LFSRcolor4[424]&LFSRcolor4[525]);
    BiasedRNG[655] = (LFSRcolor4[412]&LFSRcolor4[443]&LFSRcolor4[141]&LFSRcolor4[77]);
    BiasedRNG[656] = (LFSRcolor4[263]&LFSRcolor4[415]&LFSRcolor4[266]&LFSRcolor4[388]);
    BiasedRNG[657] = (LFSRcolor4[313]&LFSRcolor4[312]&LFSRcolor4[469]&LFSRcolor4[511]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule