//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [37:0] counter;
initial counter = 38'b0;
reg [19:0] solution;
reg [19:0] solution_check;
wire [19:0] solution_set;
initial solution_check = 20'b11110100000111101111;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
reg [0:779] InitCond;
reg run;
wire [413:0] LFSRcolor0;
wire [551:0] LFSRcolor1;
wire [413:0] LFSRcolor2;
wire [91:0] LFSRcolor3;
wire [275:0] LFSRcolor4;
reg [427:0] BiasedRNG;       //For I=+/-1 cases
reg [351:0] UnbiasedRNG;   //For I=0 cases
reg [0:809] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[260] = 1'b1;
initial m[363] = 1'b1;
initial m[373] = 1'b1;
initial m[388] = 1'b1;
initial m[408] = 1'b0;
initial m[433] = 1'b1;
initial m[463] = 1'b1;
initial m[498] = 1'b1;
initial m[538] = 1'b1;
initial m[583] = 1'b0;
initial m[628] = 1'b0;
initial m[668] = 1'b0;
initial m[703] = 1'b0;
initial m[733] = 1'b0;
initial m[758] = 1'b1;
initial m[778] = 1'b0;
initial m[793] = 1'b1;
initial m[803] = 1'b1;
initial m[808] = 1'b1;
initial m[809] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[362] = 1'b0;
initial m[372] = 1'b0;
initial m[387] = 1'b0;
initial m[407] = 1'b0;
initial m[432] = 1'b0;
initial m[462] = 1'b0;
initial m[497] = 1'b0;
initial m[537] = 1'b0;
initial m[582] = 1'b0;
initial m[585] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
//To control whether the system runs or resets using VIO and counter:
always @(posedge sample_clk) begin
    if (reset) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 20'b0;
        failure = 1'b0;
        solution_check = solution_set;
        m[260] = solution_set[0];
        m[363] = solution_set[1];
        m[373] = solution_set[2];
        m[388] = solution_set[3];
        m[408] = solution_set[4];
        m[433] = solution_set[5];
        m[463] = solution_set[6];
        m[498] = solution_set[7];
        m[538] = solution_set[8];
        m[583] = solution_set[9];
        m[628] = solution_set[10];
        m[668] = solution_set[11];
        m[703] = solution_set[12];
        m[733] = solution_set[13];
        m[758] = solution_set[14];
        m[778] = solution_set[15];
        m[793] = solution_set[16];
        m[803] = solution_set[17];
        m[808] = solution_set[18];
        m[809] = solution_set[19];
    end else if (solution_flag) begin
        run = 1'b0;
        counter = 38'b0;
        solution = 20'b0;
        failure = 1'b0;
    end else if (counter < 38'b11111111111111111111111111111111111111) begin
        if (counter == 1) begin
            InitCond[0] = UnbiasedRNG[0];
            InitCond[1] = UnbiasedRNG[1];
            InitCond[2] = UnbiasedRNG[2];
            InitCond[3] = UnbiasedRNG[3];
            InitCond[4] = UnbiasedRNG[4];
            InitCond[5] = UnbiasedRNG[5];
            InitCond[6] = UnbiasedRNG[6];
            InitCond[7] = UnbiasedRNG[7];
            InitCond[8] = UnbiasedRNG[8];
            InitCond[9] = UnbiasedRNG[9];
            InitCond[10] = UnbiasedRNG[10];
            InitCond[11] = UnbiasedRNG[11];
            InitCond[12] = UnbiasedRNG[12];
            InitCond[13] = UnbiasedRNG[13];
            InitCond[14] = UnbiasedRNG[14];
            InitCond[15] = UnbiasedRNG[15];
            InitCond[16] = UnbiasedRNG[16];
            InitCond[17] = UnbiasedRNG[17];
            InitCond[18] = UnbiasedRNG[18];
            InitCond[19] = UnbiasedRNG[19];
            InitCond[20] = UnbiasedRNG[20];
            InitCond[21] = UnbiasedRNG[21];
            InitCond[22] = UnbiasedRNG[22];
            InitCond[23] = UnbiasedRNG[23];
            InitCond[24] = UnbiasedRNG[24];
            InitCond[25] = UnbiasedRNG[25];
            InitCond[26] = UnbiasedRNG[26];
            InitCond[27] = UnbiasedRNG[27];
            InitCond[28] = UnbiasedRNG[28];
            InitCond[29] = UnbiasedRNG[29];
            InitCond[30] = UnbiasedRNG[30];
            InitCond[31] = UnbiasedRNG[31];
            InitCond[32] = UnbiasedRNG[32];
            InitCond[33] = UnbiasedRNG[33];
            InitCond[34] = UnbiasedRNG[34];
            InitCond[35] = UnbiasedRNG[35];
            InitCond[36] = UnbiasedRNG[36];
            InitCond[37] = UnbiasedRNG[37];
            InitCond[38] = UnbiasedRNG[38];
            InitCond[39] = UnbiasedRNG[39];
            InitCond[40] = UnbiasedRNG[40];
            InitCond[41] = UnbiasedRNG[41];
            InitCond[42] = UnbiasedRNG[42];
            InitCond[43] = UnbiasedRNG[43];
            InitCond[44] = UnbiasedRNG[44];
            InitCond[45] = UnbiasedRNG[45];
            InitCond[46] = UnbiasedRNG[46];
            InitCond[47] = UnbiasedRNG[47];
            InitCond[48] = UnbiasedRNG[48];
            InitCond[49] = UnbiasedRNG[49];
            InitCond[50] = UnbiasedRNG[50];
            InitCond[51] = UnbiasedRNG[51];
            InitCond[52] = UnbiasedRNG[52];
            InitCond[53] = UnbiasedRNG[53];
            InitCond[54] = UnbiasedRNG[54];
            InitCond[55] = UnbiasedRNG[55];
            InitCond[56] = UnbiasedRNG[56];
            InitCond[57] = UnbiasedRNG[57];
            InitCond[58] = UnbiasedRNG[58];
            InitCond[59] = UnbiasedRNG[59];
            InitCond[60] = UnbiasedRNG[60];
            InitCond[61] = UnbiasedRNG[61];
            InitCond[62] = UnbiasedRNG[62];
            InitCond[63] = UnbiasedRNG[63];
            InitCond[64] = UnbiasedRNG[64];
            InitCond[65] = UnbiasedRNG[65];
            InitCond[66] = UnbiasedRNG[66];
            InitCond[67] = UnbiasedRNG[67];
            InitCond[68] = UnbiasedRNG[68];
            InitCond[69] = UnbiasedRNG[69];
            InitCond[70] = UnbiasedRNG[70];
            InitCond[71] = UnbiasedRNG[71];
            InitCond[72] = UnbiasedRNG[72];
            InitCond[73] = UnbiasedRNG[73];
            InitCond[74] = UnbiasedRNG[74];
            InitCond[75] = UnbiasedRNG[75];
            InitCond[76] = UnbiasedRNG[76];
            InitCond[77] = UnbiasedRNG[77];
            InitCond[78] = UnbiasedRNG[78];
            InitCond[79] = UnbiasedRNG[79];
            InitCond[80] = UnbiasedRNG[80];
            InitCond[81] = UnbiasedRNG[81];
            InitCond[82] = UnbiasedRNG[82];
            InitCond[83] = UnbiasedRNG[83];
            InitCond[84] = UnbiasedRNG[84];
            InitCond[85] = UnbiasedRNG[85];
            InitCond[86] = UnbiasedRNG[86];
            InitCond[87] = UnbiasedRNG[87];
            InitCond[88] = UnbiasedRNG[88];
            InitCond[89] = UnbiasedRNG[89];
            InitCond[90] = UnbiasedRNG[90];
            InitCond[91] = UnbiasedRNG[91];
            InitCond[92] = UnbiasedRNG[92];
            InitCond[93] = UnbiasedRNG[93];
            InitCond[94] = UnbiasedRNG[94];
            InitCond[95] = UnbiasedRNG[95];
            InitCond[96] = UnbiasedRNG[96];
            InitCond[97] = UnbiasedRNG[97];
            InitCond[98] = UnbiasedRNG[98];
            InitCond[99] = UnbiasedRNG[99];
            InitCond[100] = UnbiasedRNG[100];
            InitCond[101] = UnbiasedRNG[101];
            InitCond[102] = UnbiasedRNG[102];
            InitCond[103] = UnbiasedRNG[103];
            InitCond[104] = UnbiasedRNG[104];
            InitCond[105] = UnbiasedRNG[105];
            InitCond[106] = UnbiasedRNG[106];
            InitCond[107] = UnbiasedRNG[107];
            InitCond[108] = UnbiasedRNG[108];
            InitCond[109] = UnbiasedRNG[109];
            InitCond[110] = UnbiasedRNG[110];
            InitCond[111] = UnbiasedRNG[111];
            InitCond[112] = UnbiasedRNG[112];
            InitCond[113] = UnbiasedRNG[113];
            InitCond[114] = UnbiasedRNG[114];
            InitCond[115] = UnbiasedRNG[115];
            InitCond[116] = UnbiasedRNG[116];
            InitCond[117] = UnbiasedRNG[117];
            InitCond[118] = UnbiasedRNG[118];
            InitCond[119] = UnbiasedRNG[119];
            InitCond[120] = UnbiasedRNG[120];
            InitCond[121] = UnbiasedRNG[121];
            InitCond[122] = UnbiasedRNG[122];
            InitCond[123] = UnbiasedRNG[123];
            InitCond[124] = UnbiasedRNG[124];
            InitCond[125] = UnbiasedRNG[125];
            InitCond[126] = UnbiasedRNG[126];
            InitCond[127] = UnbiasedRNG[127];
            InitCond[128] = UnbiasedRNG[128];
            InitCond[129] = UnbiasedRNG[129];
            InitCond[130] = UnbiasedRNG[130];
            InitCond[131] = UnbiasedRNG[131];
            InitCond[132] = UnbiasedRNG[132];
            InitCond[133] = UnbiasedRNG[133];
            InitCond[134] = UnbiasedRNG[134];
            InitCond[135] = UnbiasedRNG[135];
            InitCond[136] = UnbiasedRNG[136];
            InitCond[137] = UnbiasedRNG[137];
            InitCond[138] = UnbiasedRNG[138];
            InitCond[139] = UnbiasedRNG[139];
            InitCond[140] = UnbiasedRNG[140];
            InitCond[141] = UnbiasedRNG[141];
            InitCond[142] = UnbiasedRNG[142];
            InitCond[143] = UnbiasedRNG[143];
            InitCond[144] = UnbiasedRNG[144];
            InitCond[145] = UnbiasedRNG[145];
            InitCond[146] = UnbiasedRNG[146];
            InitCond[147] = UnbiasedRNG[147];
            InitCond[148] = UnbiasedRNG[148];
            InitCond[149] = UnbiasedRNG[149];
            InitCond[150] = UnbiasedRNG[150];
            InitCond[151] = UnbiasedRNG[151];
            InitCond[152] = UnbiasedRNG[152];
            InitCond[153] = UnbiasedRNG[153];
            InitCond[154] = UnbiasedRNG[154];
            InitCond[155] = UnbiasedRNG[155];
            InitCond[156] = UnbiasedRNG[156];
            InitCond[157] = UnbiasedRNG[157];
            InitCond[158] = UnbiasedRNG[158];
            InitCond[159] = UnbiasedRNG[159];
            InitCond[160] = UnbiasedRNG[160];
            InitCond[161] = UnbiasedRNG[161];
            InitCond[162] = UnbiasedRNG[162];
            InitCond[163] = UnbiasedRNG[163];
            InitCond[164] = UnbiasedRNG[164];
            InitCond[165] = UnbiasedRNG[165];
            InitCond[166] = UnbiasedRNG[166];
            InitCond[167] = UnbiasedRNG[167];
            InitCond[168] = UnbiasedRNG[168];
            InitCond[169] = UnbiasedRNG[169];
            InitCond[170] = UnbiasedRNG[170];
            InitCond[171] = UnbiasedRNG[171];
            InitCond[172] = UnbiasedRNG[172];
            InitCond[173] = UnbiasedRNG[173];
            InitCond[174] = UnbiasedRNG[174];
            InitCond[175] = UnbiasedRNG[175];
            InitCond[176] = UnbiasedRNG[176];
            InitCond[177] = UnbiasedRNG[177];
            InitCond[178] = UnbiasedRNG[178];
            InitCond[179] = UnbiasedRNG[179];
            InitCond[180] = UnbiasedRNG[180];
            InitCond[181] = UnbiasedRNG[181];
            InitCond[182] = UnbiasedRNG[182];
            InitCond[183] = UnbiasedRNG[183];
            InitCond[184] = UnbiasedRNG[184];
            InitCond[185] = UnbiasedRNG[185];
            InitCond[186] = UnbiasedRNG[186];
            InitCond[187] = UnbiasedRNG[187];
            InitCond[188] = UnbiasedRNG[188];
            InitCond[189] = UnbiasedRNG[189];
            InitCond[190] = UnbiasedRNG[190];
            InitCond[191] = UnbiasedRNG[191];
            InitCond[192] = UnbiasedRNG[192];
            InitCond[193] = UnbiasedRNG[193];
            InitCond[194] = UnbiasedRNG[194];
            InitCond[195] = UnbiasedRNG[195];
            InitCond[196] = UnbiasedRNG[196];
            InitCond[197] = UnbiasedRNG[197];
            InitCond[198] = UnbiasedRNG[198];
            InitCond[199] = UnbiasedRNG[199];
            InitCond[200] = UnbiasedRNG[200];
            InitCond[201] = UnbiasedRNG[201];
            InitCond[202] = UnbiasedRNG[202];
            InitCond[203] = UnbiasedRNG[203];
            InitCond[204] = UnbiasedRNG[204];
            InitCond[205] = UnbiasedRNG[205];
            InitCond[206] = UnbiasedRNG[206];
            InitCond[207] = UnbiasedRNG[207];
            InitCond[208] = UnbiasedRNG[208];
            InitCond[209] = UnbiasedRNG[209];
            InitCond[210] = UnbiasedRNG[210];
            InitCond[211] = UnbiasedRNG[211];
            InitCond[212] = UnbiasedRNG[212];
            InitCond[213] = UnbiasedRNG[213];
            InitCond[214] = UnbiasedRNG[214];
            InitCond[215] = UnbiasedRNG[215];
            InitCond[216] = UnbiasedRNG[216];
            InitCond[217] = UnbiasedRNG[217];
            InitCond[218] = UnbiasedRNG[218];
            InitCond[219] = UnbiasedRNG[219];
            InitCond[220] = UnbiasedRNG[220];
            InitCond[221] = UnbiasedRNG[221];
            InitCond[222] = UnbiasedRNG[222];
            InitCond[223] = UnbiasedRNG[223];
            InitCond[224] = UnbiasedRNG[224];
            InitCond[225] = UnbiasedRNG[225];
            InitCond[226] = UnbiasedRNG[226];
            InitCond[227] = UnbiasedRNG[227];
            InitCond[228] = UnbiasedRNG[228];
            InitCond[229] = UnbiasedRNG[229];
            InitCond[230] = UnbiasedRNG[230];
            InitCond[231] = UnbiasedRNG[231];
            InitCond[232] = UnbiasedRNG[232];
            InitCond[233] = UnbiasedRNG[233];
            InitCond[234] = UnbiasedRNG[234];
            InitCond[235] = UnbiasedRNG[235];
            InitCond[236] = UnbiasedRNG[236];
            InitCond[237] = UnbiasedRNG[237];
            InitCond[238] = UnbiasedRNG[238];
            InitCond[239] = UnbiasedRNG[239];
            InitCond[240] = UnbiasedRNG[240];
            InitCond[241] = UnbiasedRNG[241];
            InitCond[242] = UnbiasedRNG[242];
            InitCond[243] = UnbiasedRNG[243];
            InitCond[244] = UnbiasedRNG[244];
            InitCond[245] = UnbiasedRNG[245];
            InitCond[246] = UnbiasedRNG[246];
            InitCond[247] = UnbiasedRNG[247];
            InitCond[248] = UnbiasedRNG[248];
            InitCond[249] = UnbiasedRNG[249];
            InitCond[250] = UnbiasedRNG[250];
            InitCond[251] = UnbiasedRNG[251];
            InitCond[252] = UnbiasedRNG[252];
            InitCond[253] = UnbiasedRNG[253];
            InitCond[254] = UnbiasedRNG[254];
            InitCond[255] = UnbiasedRNG[255];
            InitCond[256] = UnbiasedRNG[256];
            InitCond[257] = UnbiasedRNG[257];
            InitCond[258] = UnbiasedRNG[258];
            InitCond[259] = UnbiasedRNG[259];
            InitCond[260] = UnbiasedRNG[260];
            InitCond[261] = UnbiasedRNG[261];
            InitCond[262] = UnbiasedRNG[262];
            InitCond[263] = UnbiasedRNG[263];
            InitCond[264] = UnbiasedRNG[264];
            InitCond[265] = UnbiasedRNG[265];
            InitCond[266] = UnbiasedRNG[266];
            InitCond[267] = UnbiasedRNG[267];
            InitCond[268] = UnbiasedRNG[268];
            InitCond[269] = UnbiasedRNG[269];
            InitCond[270] = UnbiasedRNG[270];
            InitCond[271] = UnbiasedRNG[271];
            InitCond[272] = UnbiasedRNG[272];
            InitCond[273] = UnbiasedRNG[273];
            InitCond[274] = UnbiasedRNG[274];
            InitCond[275] = UnbiasedRNG[275];
            InitCond[276] = UnbiasedRNG[276];
            InitCond[277] = UnbiasedRNG[277];
            InitCond[278] = UnbiasedRNG[278];
            InitCond[279] = UnbiasedRNG[279];
            InitCond[280] = UnbiasedRNG[280];
            InitCond[281] = UnbiasedRNG[281];
            InitCond[282] = UnbiasedRNG[282];
            InitCond[283] = UnbiasedRNG[283];
            InitCond[284] = UnbiasedRNG[284];
            InitCond[285] = UnbiasedRNG[285];
            InitCond[286] = UnbiasedRNG[286];
            InitCond[287] = UnbiasedRNG[287];
            InitCond[288] = UnbiasedRNG[288];
            InitCond[289] = UnbiasedRNG[289];
            InitCond[290] = UnbiasedRNG[290];
            InitCond[291] = UnbiasedRNG[291];
            InitCond[292] = UnbiasedRNG[292];
            InitCond[293] = UnbiasedRNG[293];
            InitCond[294] = UnbiasedRNG[294];
            InitCond[295] = UnbiasedRNG[295];
            InitCond[296] = UnbiasedRNG[296];
            InitCond[297] = UnbiasedRNG[297];
            InitCond[298] = UnbiasedRNG[298];
            InitCond[299] = UnbiasedRNG[299];
            InitCond[300] = UnbiasedRNG[300];
            InitCond[301] = UnbiasedRNG[301];
            InitCond[302] = UnbiasedRNG[302];
            InitCond[303] = UnbiasedRNG[303];
            InitCond[304] = UnbiasedRNG[304];
            InitCond[305] = UnbiasedRNG[305];
            InitCond[306] = UnbiasedRNG[306];
            InitCond[307] = UnbiasedRNG[307];
            InitCond[308] = UnbiasedRNG[308];
            InitCond[309] = UnbiasedRNG[309];
            InitCond[310] = UnbiasedRNG[310];
            InitCond[311] = UnbiasedRNG[311];
            InitCond[312] = UnbiasedRNG[312];
            InitCond[313] = UnbiasedRNG[313];
            InitCond[314] = UnbiasedRNG[314];
            InitCond[315] = UnbiasedRNG[315];
            InitCond[316] = UnbiasedRNG[316];
            InitCond[317] = UnbiasedRNG[317];
            InitCond[318] = UnbiasedRNG[318];
            InitCond[319] = UnbiasedRNG[319];
            InitCond[320] = UnbiasedRNG[320];
            InitCond[321] = UnbiasedRNG[321];
            InitCond[322] = UnbiasedRNG[322];
            InitCond[323] = UnbiasedRNG[323];
            InitCond[324] = UnbiasedRNG[324];
            InitCond[325] = UnbiasedRNG[325];
            InitCond[326] = UnbiasedRNG[326];
            InitCond[327] = UnbiasedRNG[327];
            InitCond[328] = UnbiasedRNG[328];
            InitCond[329] = UnbiasedRNG[329];
            InitCond[330] = UnbiasedRNG[330];
            InitCond[331] = UnbiasedRNG[331];
            InitCond[332] = UnbiasedRNG[332];
            InitCond[333] = UnbiasedRNG[333];
            InitCond[334] = UnbiasedRNG[334];
            InitCond[335] = UnbiasedRNG[335];
            InitCond[336] = UnbiasedRNG[336];
            InitCond[337] = UnbiasedRNG[337];
            InitCond[338] = UnbiasedRNG[338];
            InitCond[339] = UnbiasedRNG[339];
            InitCond[340] = UnbiasedRNG[340];
            InitCond[341] = UnbiasedRNG[341];
            InitCond[342] = UnbiasedRNG[342];
            InitCond[343] = UnbiasedRNG[343];
            InitCond[344] = UnbiasedRNG[344];
            InitCond[345] = UnbiasedRNG[345];
            InitCond[346] = UnbiasedRNG[346];
            InitCond[347] = UnbiasedRNG[347];
            InitCond[348] = UnbiasedRNG[348];
            InitCond[349] = UnbiasedRNG[349];
            InitCond[350] = UnbiasedRNG[350];
            InitCond[351] = UnbiasedRNG[351];
        end
        else if (counter == 2) begin
            InitCond[352] = UnbiasedRNG[0];
            InitCond[353] = UnbiasedRNG[1];
            InitCond[354] = UnbiasedRNG[2];
            InitCond[355] = UnbiasedRNG[3];
            InitCond[356] = UnbiasedRNG[4];
            InitCond[357] = UnbiasedRNG[5];
            InitCond[358] = UnbiasedRNG[6];
            InitCond[359] = UnbiasedRNG[7];
            InitCond[360] = UnbiasedRNG[8];
            InitCond[361] = UnbiasedRNG[9];
            InitCond[362] = UnbiasedRNG[10];
            InitCond[363] = UnbiasedRNG[11];
            InitCond[364] = UnbiasedRNG[12];
            InitCond[365] = UnbiasedRNG[13];
            InitCond[366] = UnbiasedRNG[14];
            InitCond[367] = UnbiasedRNG[15];
            InitCond[368] = UnbiasedRNG[16];
            InitCond[369] = UnbiasedRNG[17];
            InitCond[370] = UnbiasedRNG[18];
            InitCond[371] = UnbiasedRNG[19];
            InitCond[372] = UnbiasedRNG[20];
            InitCond[373] = UnbiasedRNG[21];
            InitCond[374] = UnbiasedRNG[22];
            InitCond[375] = UnbiasedRNG[23];
            InitCond[376] = UnbiasedRNG[24];
            InitCond[377] = UnbiasedRNG[25];
            InitCond[378] = UnbiasedRNG[26];
            InitCond[379] = UnbiasedRNG[27];
            InitCond[380] = UnbiasedRNG[28];
            InitCond[381] = UnbiasedRNG[29];
            InitCond[382] = UnbiasedRNG[30];
            InitCond[383] = UnbiasedRNG[31];
            InitCond[384] = UnbiasedRNG[32];
            InitCond[385] = UnbiasedRNG[33];
            InitCond[386] = UnbiasedRNG[34];
            InitCond[387] = UnbiasedRNG[35];
            InitCond[388] = UnbiasedRNG[36];
            InitCond[389] = UnbiasedRNG[37];
            InitCond[390] = UnbiasedRNG[38];
            InitCond[391] = UnbiasedRNG[39];
            InitCond[392] = UnbiasedRNG[40];
            InitCond[393] = UnbiasedRNG[41];
            InitCond[394] = UnbiasedRNG[42];
            InitCond[395] = UnbiasedRNG[43];
            InitCond[396] = UnbiasedRNG[44];
            InitCond[397] = UnbiasedRNG[45];
            InitCond[398] = UnbiasedRNG[46];
            InitCond[399] = UnbiasedRNG[47];
            InitCond[400] = UnbiasedRNG[48];
            InitCond[401] = UnbiasedRNG[49];
            InitCond[402] = UnbiasedRNG[50];
            InitCond[403] = UnbiasedRNG[51];
            InitCond[404] = UnbiasedRNG[52];
            InitCond[405] = UnbiasedRNG[53];
            InitCond[406] = UnbiasedRNG[54];
            InitCond[407] = UnbiasedRNG[55];
            InitCond[408] = UnbiasedRNG[56];
            InitCond[409] = UnbiasedRNG[57];
            InitCond[410] = UnbiasedRNG[58];
            InitCond[411] = UnbiasedRNG[59];
            InitCond[412] = UnbiasedRNG[60];
            InitCond[413] = UnbiasedRNG[61];
            InitCond[414] = UnbiasedRNG[62];
            InitCond[415] = UnbiasedRNG[63];
            InitCond[416] = UnbiasedRNG[64];
            InitCond[417] = UnbiasedRNG[65];
            InitCond[418] = UnbiasedRNG[66];
            InitCond[419] = UnbiasedRNG[67];
            InitCond[420] = UnbiasedRNG[68];
            InitCond[421] = UnbiasedRNG[69];
            InitCond[422] = UnbiasedRNG[70];
            InitCond[423] = UnbiasedRNG[71];
            InitCond[424] = UnbiasedRNG[72];
            InitCond[425] = UnbiasedRNG[73];
            InitCond[426] = UnbiasedRNG[74];
            InitCond[427] = UnbiasedRNG[75];
            InitCond[428] = UnbiasedRNG[76];
            InitCond[429] = UnbiasedRNG[77];
            InitCond[430] = UnbiasedRNG[78];
            InitCond[431] = UnbiasedRNG[79];
            InitCond[432] = UnbiasedRNG[80];
            InitCond[433] = UnbiasedRNG[81];
            InitCond[434] = UnbiasedRNG[82];
            InitCond[435] = UnbiasedRNG[83];
            InitCond[436] = UnbiasedRNG[84];
            InitCond[437] = UnbiasedRNG[85];
            InitCond[438] = UnbiasedRNG[86];
            InitCond[439] = UnbiasedRNG[87];
            InitCond[440] = UnbiasedRNG[88];
            InitCond[441] = UnbiasedRNG[89];
            InitCond[442] = UnbiasedRNG[90];
            InitCond[443] = UnbiasedRNG[91];
            InitCond[444] = UnbiasedRNG[92];
            InitCond[445] = UnbiasedRNG[93];
            InitCond[446] = UnbiasedRNG[94];
            InitCond[447] = UnbiasedRNG[95];
            InitCond[448] = UnbiasedRNG[96];
            InitCond[449] = UnbiasedRNG[97];
            InitCond[450] = UnbiasedRNG[98];
            InitCond[451] = UnbiasedRNG[99];
            InitCond[452] = UnbiasedRNG[100];
            InitCond[453] = UnbiasedRNG[101];
            InitCond[454] = UnbiasedRNG[102];
            InitCond[455] = UnbiasedRNG[103];
            InitCond[456] = UnbiasedRNG[104];
            InitCond[457] = UnbiasedRNG[105];
            InitCond[458] = UnbiasedRNG[106];
            InitCond[459] = UnbiasedRNG[107];
            InitCond[460] = UnbiasedRNG[108];
            InitCond[461] = UnbiasedRNG[109];
            InitCond[462] = UnbiasedRNG[110];
            InitCond[463] = UnbiasedRNG[111];
            InitCond[464] = UnbiasedRNG[112];
            InitCond[465] = UnbiasedRNG[113];
            InitCond[466] = UnbiasedRNG[114];
            InitCond[467] = UnbiasedRNG[115];
            InitCond[468] = UnbiasedRNG[116];
            InitCond[469] = UnbiasedRNG[117];
            InitCond[470] = UnbiasedRNG[118];
            InitCond[471] = UnbiasedRNG[119];
            InitCond[472] = UnbiasedRNG[120];
            InitCond[473] = UnbiasedRNG[121];
            InitCond[474] = UnbiasedRNG[122];
            InitCond[475] = UnbiasedRNG[123];
            InitCond[476] = UnbiasedRNG[124];
            InitCond[477] = UnbiasedRNG[125];
            InitCond[478] = UnbiasedRNG[126];
            InitCond[479] = UnbiasedRNG[127];
            InitCond[480] = UnbiasedRNG[128];
            InitCond[481] = UnbiasedRNG[129];
            InitCond[482] = UnbiasedRNG[130];
            InitCond[483] = UnbiasedRNG[131];
            InitCond[484] = UnbiasedRNG[132];
            InitCond[485] = UnbiasedRNG[133];
            InitCond[486] = UnbiasedRNG[134];
            InitCond[487] = UnbiasedRNG[135];
            InitCond[488] = UnbiasedRNG[136];
            InitCond[489] = UnbiasedRNG[137];
            InitCond[490] = UnbiasedRNG[138];
            InitCond[491] = UnbiasedRNG[139];
            InitCond[492] = UnbiasedRNG[140];
            InitCond[493] = UnbiasedRNG[141];
            InitCond[494] = UnbiasedRNG[142];
            InitCond[495] = UnbiasedRNG[143];
            InitCond[496] = UnbiasedRNG[144];
            InitCond[497] = UnbiasedRNG[145];
            InitCond[498] = UnbiasedRNG[146];
            InitCond[499] = UnbiasedRNG[147];
            InitCond[500] = UnbiasedRNG[148];
            InitCond[501] = UnbiasedRNG[149];
            InitCond[502] = UnbiasedRNG[150];
            InitCond[503] = UnbiasedRNG[151];
            InitCond[504] = UnbiasedRNG[152];
            InitCond[505] = UnbiasedRNG[153];
            InitCond[506] = UnbiasedRNG[154];
            InitCond[507] = UnbiasedRNG[155];
            InitCond[508] = UnbiasedRNG[156];
            InitCond[509] = UnbiasedRNG[157];
            InitCond[510] = UnbiasedRNG[158];
            InitCond[511] = UnbiasedRNG[159];
            InitCond[512] = UnbiasedRNG[160];
            InitCond[513] = UnbiasedRNG[161];
            InitCond[514] = UnbiasedRNG[162];
            InitCond[515] = UnbiasedRNG[163];
            InitCond[516] = UnbiasedRNG[164];
            InitCond[517] = UnbiasedRNG[165];
            InitCond[518] = UnbiasedRNG[166];
            InitCond[519] = UnbiasedRNG[167];
            InitCond[520] = UnbiasedRNG[168];
            InitCond[521] = UnbiasedRNG[169];
            InitCond[522] = UnbiasedRNG[170];
            InitCond[523] = UnbiasedRNG[171];
            InitCond[524] = UnbiasedRNG[172];
            InitCond[525] = UnbiasedRNG[173];
            InitCond[526] = UnbiasedRNG[174];
            InitCond[527] = UnbiasedRNG[175];
            InitCond[528] = UnbiasedRNG[176];
            InitCond[529] = UnbiasedRNG[177];
            InitCond[530] = UnbiasedRNG[178];
            InitCond[531] = UnbiasedRNG[179];
            InitCond[532] = UnbiasedRNG[180];
            InitCond[533] = UnbiasedRNG[181];
            InitCond[534] = UnbiasedRNG[182];
            InitCond[535] = UnbiasedRNG[183];
            InitCond[536] = UnbiasedRNG[184];
            InitCond[537] = UnbiasedRNG[185];
            InitCond[538] = UnbiasedRNG[186];
            InitCond[539] = UnbiasedRNG[187];
            InitCond[540] = UnbiasedRNG[188];
            InitCond[541] = UnbiasedRNG[189];
            InitCond[542] = UnbiasedRNG[190];
            InitCond[543] = UnbiasedRNG[191];
            InitCond[544] = UnbiasedRNG[192];
            InitCond[545] = UnbiasedRNG[193];
            InitCond[546] = UnbiasedRNG[194];
            InitCond[547] = UnbiasedRNG[195];
            InitCond[548] = UnbiasedRNG[196];
            InitCond[549] = UnbiasedRNG[197];
            InitCond[550] = UnbiasedRNG[198];
            InitCond[551] = UnbiasedRNG[199];
            InitCond[552] = UnbiasedRNG[200];
            InitCond[553] = UnbiasedRNG[201];
            InitCond[554] = UnbiasedRNG[202];
            InitCond[555] = UnbiasedRNG[203];
            InitCond[556] = UnbiasedRNG[204];
            InitCond[557] = UnbiasedRNG[205];
            InitCond[558] = UnbiasedRNG[206];
            InitCond[559] = UnbiasedRNG[207];
            InitCond[560] = UnbiasedRNG[208];
            InitCond[561] = UnbiasedRNG[209];
            InitCond[562] = UnbiasedRNG[210];
            InitCond[563] = UnbiasedRNG[211];
            InitCond[564] = UnbiasedRNG[212];
            InitCond[565] = UnbiasedRNG[213];
            InitCond[566] = UnbiasedRNG[214];
            InitCond[567] = UnbiasedRNG[215];
            InitCond[568] = UnbiasedRNG[216];
            InitCond[569] = UnbiasedRNG[217];
            InitCond[570] = UnbiasedRNG[218];
            InitCond[571] = UnbiasedRNG[219];
            InitCond[572] = UnbiasedRNG[220];
            InitCond[573] = UnbiasedRNG[221];
            InitCond[574] = UnbiasedRNG[222];
            InitCond[575] = UnbiasedRNG[223];
            InitCond[576] = UnbiasedRNG[224];
            InitCond[577] = UnbiasedRNG[225];
            InitCond[578] = UnbiasedRNG[226];
            InitCond[579] = UnbiasedRNG[227];
            InitCond[580] = UnbiasedRNG[228];
            InitCond[581] = UnbiasedRNG[229];
            InitCond[582] = UnbiasedRNG[230];
            InitCond[583] = UnbiasedRNG[231];
            InitCond[584] = UnbiasedRNG[232];
            InitCond[585] = UnbiasedRNG[233];
            InitCond[586] = UnbiasedRNG[234];
            InitCond[587] = UnbiasedRNG[235];
            InitCond[588] = UnbiasedRNG[236];
            InitCond[589] = UnbiasedRNG[237];
            InitCond[590] = UnbiasedRNG[238];
            InitCond[591] = UnbiasedRNG[239];
            InitCond[592] = UnbiasedRNG[240];
            InitCond[593] = UnbiasedRNG[241];
            InitCond[594] = UnbiasedRNG[242];
            InitCond[595] = UnbiasedRNG[243];
            InitCond[596] = UnbiasedRNG[244];
            InitCond[597] = UnbiasedRNG[245];
            InitCond[598] = UnbiasedRNG[246];
            InitCond[599] = UnbiasedRNG[247];
            InitCond[600] = UnbiasedRNG[248];
            InitCond[601] = UnbiasedRNG[249];
            InitCond[602] = UnbiasedRNG[250];
            InitCond[603] = UnbiasedRNG[251];
            InitCond[604] = UnbiasedRNG[252];
            InitCond[605] = UnbiasedRNG[253];
            InitCond[606] = UnbiasedRNG[254];
            InitCond[607] = UnbiasedRNG[255];
            InitCond[608] = UnbiasedRNG[256];
            InitCond[609] = UnbiasedRNG[257];
            InitCond[610] = UnbiasedRNG[258];
            InitCond[611] = UnbiasedRNG[259];
            InitCond[612] = UnbiasedRNG[260];
            InitCond[613] = UnbiasedRNG[261];
            InitCond[614] = UnbiasedRNG[262];
            InitCond[615] = UnbiasedRNG[263];
            InitCond[616] = UnbiasedRNG[264];
            InitCond[617] = UnbiasedRNG[265];
            InitCond[618] = UnbiasedRNG[266];
            InitCond[619] = UnbiasedRNG[267];
            InitCond[620] = UnbiasedRNG[268];
            InitCond[621] = UnbiasedRNG[269];
            InitCond[622] = UnbiasedRNG[270];
            InitCond[623] = UnbiasedRNG[271];
            InitCond[624] = UnbiasedRNG[272];
            InitCond[625] = UnbiasedRNG[273];
            InitCond[626] = UnbiasedRNG[274];
            InitCond[627] = UnbiasedRNG[275];
            InitCond[628] = UnbiasedRNG[276];
            InitCond[629] = UnbiasedRNG[277];
            InitCond[630] = UnbiasedRNG[278];
            InitCond[631] = UnbiasedRNG[279];
            InitCond[632] = UnbiasedRNG[280];
            InitCond[633] = UnbiasedRNG[281];
            InitCond[634] = UnbiasedRNG[282];
            InitCond[635] = UnbiasedRNG[283];
            InitCond[636] = UnbiasedRNG[284];
            InitCond[637] = UnbiasedRNG[285];
            InitCond[638] = UnbiasedRNG[286];
            InitCond[639] = UnbiasedRNG[287];
            InitCond[640] = UnbiasedRNG[288];
            InitCond[641] = UnbiasedRNG[289];
            InitCond[642] = UnbiasedRNG[290];
            InitCond[643] = UnbiasedRNG[291];
            InitCond[644] = UnbiasedRNG[292];
            InitCond[645] = UnbiasedRNG[293];
            InitCond[646] = UnbiasedRNG[294];
            InitCond[647] = UnbiasedRNG[295];
            InitCond[648] = UnbiasedRNG[296];
            InitCond[649] = UnbiasedRNG[297];
            InitCond[650] = UnbiasedRNG[298];
            InitCond[651] = UnbiasedRNG[299];
            InitCond[652] = UnbiasedRNG[300];
            InitCond[653] = UnbiasedRNG[301];
            InitCond[654] = UnbiasedRNG[302];
            InitCond[655] = UnbiasedRNG[303];
            InitCond[656] = UnbiasedRNG[304];
            InitCond[657] = UnbiasedRNG[305];
            InitCond[658] = UnbiasedRNG[306];
            InitCond[659] = UnbiasedRNG[307];
            InitCond[660] = UnbiasedRNG[308];
            InitCond[661] = UnbiasedRNG[309];
            InitCond[662] = UnbiasedRNG[310];
            InitCond[663] = UnbiasedRNG[311];
            InitCond[664] = UnbiasedRNG[312];
            InitCond[665] = UnbiasedRNG[313];
            InitCond[666] = UnbiasedRNG[314];
            InitCond[667] = UnbiasedRNG[315];
            InitCond[668] = UnbiasedRNG[316];
            InitCond[669] = UnbiasedRNG[317];
            InitCond[670] = UnbiasedRNG[318];
            InitCond[671] = UnbiasedRNG[319];
            InitCond[672] = UnbiasedRNG[320];
            InitCond[673] = UnbiasedRNG[321];
            InitCond[674] = UnbiasedRNG[322];
            InitCond[675] = UnbiasedRNG[323];
            InitCond[676] = UnbiasedRNG[324];
            InitCond[677] = UnbiasedRNG[325];
            InitCond[678] = UnbiasedRNG[326];
            InitCond[679] = UnbiasedRNG[327];
            InitCond[680] = UnbiasedRNG[328];
            InitCond[681] = UnbiasedRNG[329];
            InitCond[682] = UnbiasedRNG[330];
            InitCond[683] = UnbiasedRNG[331];
            InitCond[684] = UnbiasedRNG[332];
            InitCond[685] = UnbiasedRNG[333];
            InitCond[686] = UnbiasedRNG[334];
            InitCond[687] = UnbiasedRNG[335];
            InitCond[688] = UnbiasedRNG[336];
            InitCond[689] = UnbiasedRNG[337];
            InitCond[690] = UnbiasedRNG[338];
            InitCond[691] = UnbiasedRNG[339];
            InitCond[692] = UnbiasedRNG[340];
            InitCond[693] = UnbiasedRNG[341];
            InitCond[694] = UnbiasedRNG[342];
            InitCond[695] = UnbiasedRNG[343];
            InitCond[696] = UnbiasedRNG[344];
            InitCond[697] = UnbiasedRNG[345];
            InitCond[698] = UnbiasedRNG[346];
            InitCond[699] = UnbiasedRNG[347];
            InitCond[700] = UnbiasedRNG[348];
            InitCond[701] = UnbiasedRNG[349];
            InitCond[702] = UnbiasedRNG[350];
            InitCond[703] = UnbiasedRNG[351];
        end
        else if (counter == 3) begin
            InitCond[704] = UnbiasedRNG[0];
            InitCond[705] = UnbiasedRNG[1];
            InitCond[706] = UnbiasedRNG[2];
            InitCond[707] = UnbiasedRNG[3];
            InitCond[708] = UnbiasedRNG[4];
            InitCond[709] = UnbiasedRNG[5];
            InitCond[710] = UnbiasedRNG[6];
            InitCond[711] = UnbiasedRNG[7];
            InitCond[712] = UnbiasedRNG[8];
            InitCond[713] = UnbiasedRNG[9];
            InitCond[714] = UnbiasedRNG[10];
            InitCond[715] = UnbiasedRNG[11];
            InitCond[716] = UnbiasedRNG[12];
            InitCond[717] = UnbiasedRNG[13];
            InitCond[718] = UnbiasedRNG[14];
            InitCond[719] = UnbiasedRNG[15];
            InitCond[720] = UnbiasedRNG[16];
            InitCond[721] = UnbiasedRNG[17];
            InitCond[722] = UnbiasedRNG[18];
            InitCond[723] = UnbiasedRNG[19];
            InitCond[724] = UnbiasedRNG[20];
            InitCond[725] = UnbiasedRNG[21];
            InitCond[726] = UnbiasedRNG[22];
            InitCond[727] = UnbiasedRNG[23];
            InitCond[728] = UnbiasedRNG[24];
            InitCond[729] = UnbiasedRNG[25];
            InitCond[730] = UnbiasedRNG[26];
            InitCond[731] = UnbiasedRNG[27];
            InitCond[732] = UnbiasedRNG[28];
            InitCond[733] = UnbiasedRNG[29];
            InitCond[734] = UnbiasedRNG[30];
            InitCond[735] = UnbiasedRNG[31];
            InitCond[736] = UnbiasedRNG[32];
            InitCond[737] = UnbiasedRNG[33];
            InitCond[738] = UnbiasedRNG[34];
            InitCond[739] = UnbiasedRNG[35];
            InitCond[740] = UnbiasedRNG[36];
            InitCond[741] = UnbiasedRNG[37];
            InitCond[742] = UnbiasedRNG[38];
            InitCond[743] = UnbiasedRNG[39];
            InitCond[744] = UnbiasedRNG[40];
            InitCond[745] = UnbiasedRNG[41];
            InitCond[746] = UnbiasedRNG[42];
            InitCond[747] = UnbiasedRNG[43];
            InitCond[748] = UnbiasedRNG[44];
            InitCond[749] = UnbiasedRNG[45];
            InitCond[750] = UnbiasedRNG[46];
            InitCond[751] = UnbiasedRNG[47];
            InitCond[752] = UnbiasedRNG[48];
            InitCond[753] = UnbiasedRNG[49];
            InitCond[754] = UnbiasedRNG[50];
            InitCond[755] = UnbiasedRNG[51];
            InitCond[756] = UnbiasedRNG[52];
            InitCond[757] = UnbiasedRNG[53];
            InitCond[758] = UnbiasedRNG[54];
            InitCond[759] = UnbiasedRNG[55];
            InitCond[760] = UnbiasedRNG[56];
            InitCond[761] = UnbiasedRNG[57];
            InitCond[762] = UnbiasedRNG[58];
            InitCond[763] = UnbiasedRNG[59];
            InitCond[764] = UnbiasedRNG[60];
            InitCond[765] = UnbiasedRNG[61];
            InitCond[766] = UnbiasedRNG[62];
            InitCond[767] = UnbiasedRNG[63];
            InitCond[768] = UnbiasedRNG[64];
            InitCond[769] = UnbiasedRNG[65];
            InitCond[770] = UnbiasedRNG[66];
            InitCond[771] = UnbiasedRNG[67];
            InitCond[772] = UnbiasedRNG[68];
            InitCond[773] = UnbiasedRNG[69];
            InitCond[774] = UnbiasedRNG[70];
            InitCond[775] = UnbiasedRNG[71];
            InitCond[776] = UnbiasedRNG[72];
            InitCond[777] = UnbiasedRNG[73];
            InitCond[778] = UnbiasedRNG[74];
            InitCond[779] = UnbiasedRNG[75];
        end
        else if (counter==5)
            run = 1'b1;
        counter = counter+38'b1;
        solution = {m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[19],m[18],m[17],m[16],m[15],m[14],m[13],m[12],m[11],m[10]};
    end else begin 
        counter = 38'b0;
        failure = 1'b1;
        run = 1'b0;
    end
end

//To measure on only the last step using ILA:
always @(negedge sample_clk) begin
    if (solution_flag)
        solution_flag = 1'b0;
    else if ((run & (solution == solution_check)) | failure)
        solution_flag = 1'b1;
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = run?((((m[20]&m[21]&~m[60]&~m[61])|(m[20]&~m[21]&m[60]&~m[61])|(~m[20]&m[21]&m[60]&~m[61])|(m[20]&~m[21]&~m[60]&m[61])|(~m[20]&m[21]&~m[60]&m[61])|(~m[20]&~m[21]&m[60]&m[61]))&UnbiasedRNG[0])|((m[20]&m[21]&m[60]&~m[61])|(m[20]&m[21]&~m[60]&m[61])|(m[20]&~m[21]&m[60]&m[61])|(~m[20]&m[21]&m[60]&m[61])|(m[20]&m[21]&m[60]&m[61]))):InitCond[0];
    m[1] = run?((((m[22]&m[23]&~m[70]&~m[71])|(m[22]&~m[23]&m[70]&~m[71])|(~m[22]&m[23]&m[70]&~m[71])|(m[22]&~m[23]&~m[70]&m[71])|(~m[22]&m[23]&~m[70]&m[71])|(~m[22]&~m[23]&m[70]&m[71]))&UnbiasedRNG[1])|((m[22]&m[23]&m[70]&~m[71])|(m[22]&m[23]&~m[70]&m[71])|(m[22]&~m[23]&m[70]&m[71])|(~m[22]&m[23]&m[70]&m[71])|(m[22]&m[23]&m[70]&m[71]))):InitCond[1];
    m[2] = run?((((m[24]&m[25]&~m[80]&~m[81])|(m[24]&~m[25]&m[80]&~m[81])|(~m[24]&m[25]&m[80]&~m[81])|(m[24]&~m[25]&~m[80]&m[81])|(~m[24]&m[25]&~m[80]&m[81])|(~m[24]&~m[25]&m[80]&m[81]))&UnbiasedRNG[2])|((m[24]&m[25]&m[80]&~m[81])|(m[24]&m[25]&~m[80]&m[81])|(m[24]&~m[25]&m[80]&m[81])|(~m[24]&m[25]&m[80]&m[81])|(m[24]&m[25]&m[80]&m[81]))):InitCond[2];
    m[3] = run?((((m[26]&m[27]&~m[90]&~m[91])|(m[26]&~m[27]&m[90]&~m[91])|(~m[26]&m[27]&m[90]&~m[91])|(m[26]&~m[27]&~m[90]&m[91])|(~m[26]&m[27]&~m[90]&m[91])|(~m[26]&~m[27]&m[90]&m[91]))&UnbiasedRNG[3])|((m[26]&m[27]&m[90]&~m[91])|(m[26]&m[27]&~m[90]&m[91])|(m[26]&~m[27]&m[90]&m[91])|(~m[26]&m[27]&m[90]&m[91])|(m[26]&m[27]&m[90]&m[91]))):InitCond[3];
    m[4] = run?((((m[28]&m[29]&~m[100]&~m[101])|(m[28]&~m[29]&m[100]&~m[101])|(~m[28]&m[29]&m[100]&~m[101])|(m[28]&~m[29]&~m[100]&m[101])|(~m[28]&m[29]&~m[100]&m[101])|(~m[28]&~m[29]&m[100]&m[101]))&UnbiasedRNG[4])|((m[28]&m[29]&m[100]&~m[101])|(m[28]&m[29]&~m[100]&m[101])|(m[28]&~m[29]&m[100]&m[101])|(~m[28]&m[29]&m[100]&m[101])|(m[28]&m[29]&m[100]&m[101]))):InitCond[4];
    m[5] = run?((((m[30]&m[31]&~m[110]&~m[111])|(m[30]&~m[31]&m[110]&~m[111])|(~m[30]&m[31]&m[110]&~m[111])|(m[30]&~m[31]&~m[110]&m[111])|(~m[30]&m[31]&~m[110]&m[111])|(~m[30]&~m[31]&m[110]&m[111]))&UnbiasedRNG[5])|((m[30]&m[31]&m[110]&~m[111])|(m[30]&m[31]&~m[110]&m[111])|(m[30]&~m[31]&m[110]&m[111])|(~m[30]&m[31]&m[110]&m[111])|(m[30]&m[31]&m[110]&m[111]))):InitCond[5];
    m[6] = run?((((m[32]&m[33]&~m[120]&~m[121])|(m[32]&~m[33]&m[120]&~m[121])|(~m[32]&m[33]&m[120]&~m[121])|(m[32]&~m[33]&~m[120]&m[121])|(~m[32]&m[33]&~m[120]&m[121])|(~m[32]&~m[33]&m[120]&m[121]))&UnbiasedRNG[6])|((m[32]&m[33]&m[120]&~m[121])|(m[32]&m[33]&~m[120]&m[121])|(m[32]&~m[33]&m[120]&m[121])|(~m[32]&m[33]&m[120]&m[121])|(m[32]&m[33]&m[120]&m[121]))):InitCond[6];
    m[7] = run?((((m[34]&m[35]&~m[130]&~m[131])|(m[34]&~m[35]&m[130]&~m[131])|(~m[34]&m[35]&m[130]&~m[131])|(m[34]&~m[35]&~m[130]&m[131])|(~m[34]&m[35]&~m[130]&m[131])|(~m[34]&~m[35]&m[130]&m[131]))&UnbiasedRNG[7])|((m[34]&m[35]&m[130]&~m[131])|(m[34]&m[35]&~m[130]&m[131])|(m[34]&~m[35]&m[130]&m[131])|(~m[34]&m[35]&m[130]&m[131])|(m[34]&m[35]&m[130]&m[131]))):InitCond[7];
    m[8] = run?((((m[36]&m[37]&~m[140]&~m[141])|(m[36]&~m[37]&m[140]&~m[141])|(~m[36]&m[37]&m[140]&~m[141])|(m[36]&~m[37]&~m[140]&m[141])|(~m[36]&m[37]&~m[140]&m[141])|(~m[36]&~m[37]&m[140]&m[141]))&UnbiasedRNG[8])|((m[36]&m[37]&m[140]&~m[141])|(m[36]&m[37]&~m[140]&m[141])|(m[36]&~m[37]&m[140]&m[141])|(~m[36]&m[37]&m[140]&m[141])|(m[36]&m[37]&m[140]&m[141]))):InitCond[8];
    m[9] = run?((((m[38]&m[39]&~m[150]&~m[151])|(m[38]&~m[39]&m[150]&~m[151])|(~m[38]&m[39]&m[150]&~m[151])|(m[38]&~m[39]&~m[150]&m[151])|(~m[38]&m[39]&~m[150]&m[151])|(~m[38]&~m[39]&m[150]&m[151]))&UnbiasedRNG[9])|((m[38]&m[39]&m[150]&~m[151])|(m[38]&m[39]&~m[150]&m[151])|(m[38]&~m[39]&m[150]&m[151])|(~m[38]&m[39]&m[150]&m[151])|(m[38]&m[39]&m[150]&m[151]))):InitCond[9];
    m[10] = run?((((m[40]&m[41]&~m[160]&~m[161])|(m[40]&~m[41]&m[160]&~m[161])|(~m[40]&m[41]&m[160]&~m[161])|(m[40]&~m[41]&~m[160]&m[161])|(~m[40]&m[41]&~m[160]&m[161])|(~m[40]&~m[41]&m[160]&m[161]))&UnbiasedRNG[10])|((m[40]&m[41]&m[160]&~m[161])|(m[40]&m[41]&~m[160]&m[161])|(m[40]&~m[41]&m[160]&m[161])|(~m[40]&m[41]&m[160]&m[161])|(m[40]&m[41]&m[160]&m[161]))):InitCond[10];
    m[11] = run?((((m[42]&m[43]&~m[170]&~m[171])|(m[42]&~m[43]&m[170]&~m[171])|(~m[42]&m[43]&m[170]&~m[171])|(m[42]&~m[43]&~m[170]&m[171])|(~m[42]&m[43]&~m[170]&m[171])|(~m[42]&~m[43]&m[170]&m[171]))&UnbiasedRNG[11])|((m[42]&m[43]&m[170]&~m[171])|(m[42]&m[43]&~m[170]&m[171])|(m[42]&~m[43]&m[170]&m[171])|(~m[42]&m[43]&m[170]&m[171])|(m[42]&m[43]&m[170]&m[171]))):InitCond[11];
    m[12] = run?((((m[44]&m[45]&~m[180]&~m[181])|(m[44]&~m[45]&m[180]&~m[181])|(~m[44]&m[45]&m[180]&~m[181])|(m[44]&~m[45]&~m[180]&m[181])|(~m[44]&m[45]&~m[180]&m[181])|(~m[44]&~m[45]&m[180]&m[181]))&UnbiasedRNG[12])|((m[44]&m[45]&m[180]&~m[181])|(m[44]&m[45]&~m[180]&m[181])|(m[44]&~m[45]&m[180]&m[181])|(~m[44]&m[45]&m[180]&m[181])|(m[44]&m[45]&m[180]&m[181]))):InitCond[12];
    m[13] = run?((((m[46]&m[47]&~m[190]&~m[191])|(m[46]&~m[47]&m[190]&~m[191])|(~m[46]&m[47]&m[190]&~m[191])|(m[46]&~m[47]&~m[190]&m[191])|(~m[46]&m[47]&~m[190]&m[191])|(~m[46]&~m[47]&m[190]&m[191]))&UnbiasedRNG[13])|((m[46]&m[47]&m[190]&~m[191])|(m[46]&m[47]&~m[190]&m[191])|(m[46]&~m[47]&m[190]&m[191])|(~m[46]&m[47]&m[190]&m[191])|(m[46]&m[47]&m[190]&m[191]))):InitCond[13];
    m[14] = run?((((m[48]&m[49]&~m[200]&~m[201])|(m[48]&~m[49]&m[200]&~m[201])|(~m[48]&m[49]&m[200]&~m[201])|(m[48]&~m[49]&~m[200]&m[201])|(~m[48]&m[49]&~m[200]&m[201])|(~m[48]&~m[49]&m[200]&m[201]))&UnbiasedRNG[14])|((m[48]&m[49]&m[200]&~m[201])|(m[48]&m[49]&~m[200]&m[201])|(m[48]&~m[49]&m[200]&m[201])|(~m[48]&m[49]&m[200]&m[201])|(m[48]&m[49]&m[200]&m[201]))):InitCond[14];
    m[15] = run?((((m[50]&m[51]&~m[210]&~m[211])|(m[50]&~m[51]&m[210]&~m[211])|(~m[50]&m[51]&m[210]&~m[211])|(m[50]&~m[51]&~m[210]&m[211])|(~m[50]&m[51]&~m[210]&m[211])|(~m[50]&~m[51]&m[210]&m[211]))&UnbiasedRNG[15])|((m[50]&m[51]&m[210]&~m[211])|(m[50]&m[51]&~m[210]&m[211])|(m[50]&~m[51]&m[210]&m[211])|(~m[50]&m[51]&m[210]&m[211])|(m[50]&m[51]&m[210]&m[211]))):InitCond[15];
    m[16] = run?((((m[52]&m[53]&~m[220]&~m[221])|(m[52]&~m[53]&m[220]&~m[221])|(~m[52]&m[53]&m[220]&~m[221])|(m[52]&~m[53]&~m[220]&m[221])|(~m[52]&m[53]&~m[220]&m[221])|(~m[52]&~m[53]&m[220]&m[221]))&UnbiasedRNG[16])|((m[52]&m[53]&m[220]&~m[221])|(m[52]&m[53]&~m[220]&m[221])|(m[52]&~m[53]&m[220]&m[221])|(~m[52]&m[53]&m[220]&m[221])|(m[52]&m[53]&m[220]&m[221]))):InitCond[16];
    m[17] = run?((((m[54]&m[55]&~m[230]&~m[231])|(m[54]&~m[55]&m[230]&~m[231])|(~m[54]&m[55]&m[230]&~m[231])|(m[54]&~m[55]&~m[230]&m[231])|(~m[54]&m[55]&~m[230]&m[231])|(~m[54]&~m[55]&m[230]&m[231]))&UnbiasedRNG[17])|((m[54]&m[55]&m[230]&~m[231])|(m[54]&m[55]&~m[230]&m[231])|(m[54]&~m[55]&m[230]&m[231])|(~m[54]&m[55]&m[230]&m[231])|(m[54]&m[55]&m[230]&m[231]))):InitCond[17];
    m[18] = run?((((m[56]&m[57]&~m[240]&~m[241])|(m[56]&~m[57]&m[240]&~m[241])|(~m[56]&m[57]&m[240]&~m[241])|(m[56]&~m[57]&~m[240]&m[241])|(~m[56]&m[57]&~m[240]&m[241])|(~m[56]&~m[57]&m[240]&m[241]))&UnbiasedRNG[18])|((m[56]&m[57]&m[240]&~m[241])|(m[56]&m[57]&~m[240]&m[241])|(m[56]&~m[57]&m[240]&m[241])|(~m[56]&m[57]&m[240]&m[241])|(m[56]&m[57]&m[240]&m[241]))):InitCond[18];
    m[19] = run?((((m[58]&m[59]&~m[250]&~m[251])|(m[58]&~m[59]&m[250]&~m[251])|(~m[58]&m[59]&m[250]&~m[251])|(m[58]&~m[59]&~m[250]&m[251])|(~m[58]&m[59]&~m[250]&m[251])|(~m[58]&~m[59]&m[250]&m[251]))&UnbiasedRNG[19])|((m[58]&m[59]&m[250]&~m[251])|(m[58]&m[59]&~m[250]&m[251])|(m[58]&~m[59]&m[250]&m[251])|(~m[58]&m[59]&m[250]&m[251])|(m[58]&m[59]&m[250]&m[251]))):InitCond[19];
    m[62] = run?((((~m[20]&~m[180]&~m[280])|(m[20]&m[180]&~m[280]))&BiasedRNG[0])|(((m[20]&~m[180]&~m[280])|(~m[20]&m[180]&m[280]))&~BiasedRNG[0])|((~m[20]&~m[180]&m[280])|(m[20]&~m[180]&m[280])|(m[20]&m[180]&m[280]))):InitCond[20];
    m[63] = run?((((~m[20]&~m[190]&~m[290])|(m[20]&m[190]&~m[290]))&BiasedRNG[1])|(((m[20]&~m[190]&~m[290])|(~m[20]&m[190]&m[290]))&~BiasedRNG[1])|((~m[20]&~m[190]&m[290])|(m[20]&~m[190]&m[290])|(m[20]&m[190]&m[290]))):InitCond[21];
    m[64] = run?((((~m[20]&~m[200]&~m[300])|(m[20]&m[200]&~m[300]))&BiasedRNG[2])|(((m[20]&~m[200]&~m[300])|(~m[20]&m[200]&m[300]))&~BiasedRNG[2])|((~m[20]&~m[200]&m[300])|(m[20]&~m[200]&m[300])|(m[20]&m[200]&m[300]))):InitCond[22];
    m[65] = run?((((~m[20]&~m[210]&~m[310])|(m[20]&m[210]&~m[310]))&BiasedRNG[3])|(((m[20]&~m[210]&~m[310])|(~m[20]&m[210]&m[310]))&~BiasedRNG[3])|((~m[20]&~m[210]&m[310])|(m[20]&~m[210]&m[310])|(m[20]&m[210]&m[310]))):InitCond[23];
    m[66] = run?((((~m[21]&~m[220]&~m[320])|(m[21]&m[220]&~m[320]))&BiasedRNG[4])|(((m[21]&~m[220]&~m[320])|(~m[21]&m[220]&m[320]))&~BiasedRNG[4])|((~m[21]&~m[220]&m[320])|(m[21]&~m[220]&m[320])|(m[21]&m[220]&m[320]))):InitCond[24];
    m[67] = run?((((~m[21]&~m[230]&~m[330])|(m[21]&m[230]&~m[330]))&BiasedRNG[5])|(((m[21]&~m[230]&~m[330])|(~m[21]&m[230]&m[330]))&~BiasedRNG[5])|((~m[21]&~m[230]&m[330])|(m[21]&~m[230]&m[330])|(m[21]&m[230]&m[330]))):InitCond[25];
    m[68] = run?((((~m[21]&~m[240]&~m[340])|(m[21]&m[240]&~m[340]))&BiasedRNG[6])|(((m[21]&~m[240]&~m[340])|(~m[21]&m[240]&m[340]))&~BiasedRNG[6])|((~m[21]&~m[240]&m[340])|(m[21]&~m[240]&m[340])|(m[21]&m[240]&m[340]))):InitCond[26];
    m[69] = run?((((~m[21]&~m[250]&~m[350])|(m[21]&m[250]&~m[350]))&BiasedRNG[7])|(((m[21]&~m[250]&~m[350])|(~m[21]&m[250]&m[350]))&~BiasedRNG[7])|((~m[21]&~m[250]&m[350])|(m[21]&~m[250]&m[350])|(m[21]&m[250]&m[350]))):InitCond[27];
    m[72] = run?((((~m[22]&~m[181]&~m[281])|(m[22]&m[181]&~m[281]))&BiasedRNG[8])|(((m[22]&~m[181]&~m[281])|(~m[22]&m[181]&m[281]))&~BiasedRNG[8])|((~m[22]&~m[181]&m[281])|(m[22]&~m[181]&m[281])|(m[22]&m[181]&m[281]))):InitCond[28];
    m[73] = run?((((~m[22]&~m[191]&~m[291])|(m[22]&m[191]&~m[291]))&BiasedRNG[9])|(((m[22]&~m[191]&~m[291])|(~m[22]&m[191]&m[291]))&~BiasedRNG[9])|((~m[22]&~m[191]&m[291])|(m[22]&~m[191]&m[291])|(m[22]&m[191]&m[291]))):InitCond[29];
    m[74] = run?((((~m[22]&~m[201]&~m[301])|(m[22]&m[201]&~m[301]))&BiasedRNG[10])|(((m[22]&~m[201]&~m[301])|(~m[22]&m[201]&m[301]))&~BiasedRNG[10])|((~m[22]&~m[201]&m[301])|(m[22]&~m[201]&m[301])|(m[22]&m[201]&m[301]))):InitCond[30];
    m[75] = run?((((~m[22]&~m[211]&~m[311])|(m[22]&m[211]&~m[311]))&BiasedRNG[11])|(((m[22]&~m[211]&~m[311])|(~m[22]&m[211]&m[311]))&~BiasedRNG[11])|((~m[22]&~m[211]&m[311])|(m[22]&~m[211]&m[311])|(m[22]&m[211]&m[311]))):InitCond[31];
    m[76] = run?((((~m[23]&~m[221]&~m[321])|(m[23]&m[221]&~m[321]))&BiasedRNG[12])|(((m[23]&~m[221]&~m[321])|(~m[23]&m[221]&m[321]))&~BiasedRNG[12])|((~m[23]&~m[221]&m[321])|(m[23]&~m[221]&m[321])|(m[23]&m[221]&m[321]))):InitCond[32];
    m[77] = run?((((~m[23]&~m[231]&~m[331])|(m[23]&m[231]&~m[331]))&BiasedRNG[13])|(((m[23]&~m[231]&~m[331])|(~m[23]&m[231]&m[331]))&~BiasedRNG[13])|((~m[23]&~m[231]&m[331])|(m[23]&~m[231]&m[331])|(m[23]&m[231]&m[331]))):InitCond[33];
    m[78] = run?((((~m[23]&~m[241]&~m[341])|(m[23]&m[241]&~m[341]))&BiasedRNG[14])|(((m[23]&~m[241]&~m[341])|(~m[23]&m[241]&m[341]))&~BiasedRNG[14])|((~m[23]&~m[241]&m[341])|(m[23]&~m[241]&m[341])|(m[23]&m[241]&m[341]))):InitCond[34];
    m[79] = run?((((~m[23]&~m[251]&~m[351])|(m[23]&m[251]&~m[351]))&BiasedRNG[15])|(((m[23]&~m[251]&~m[351])|(~m[23]&m[251]&m[351]))&~BiasedRNG[15])|((~m[23]&~m[251]&m[351])|(m[23]&~m[251]&m[351])|(m[23]&m[251]&m[351]))):InitCond[35];
    m[82] = run?((((~m[24]&~m[182]&~m[282])|(m[24]&m[182]&~m[282]))&BiasedRNG[16])|(((m[24]&~m[182]&~m[282])|(~m[24]&m[182]&m[282]))&~BiasedRNG[16])|((~m[24]&~m[182]&m[282])|(m[24]&~m[182]&m[282])|(m[24]&m[182]&m[282]))):InitCond[36];
    m[83] = run?((((~m[24]&~m[192]&~m[292])|(m[24]&m[192]&~m[292]))&BiasedRNG[17])|(((m[24]&~m[192]&~m[292])|(~m[24]&m[192]&m[292]))&~BiasedRNG[17])|((~m[24]&~m[192]&m[292])|(m[24]&~m[192]&m[292])|(m[24]&m[192]&m[292]))):InitCond[37];
    m[84] = run?((((~m[24]&~m[202]&~m[302])|(m[24]&m[202]&~m[302]))&BiasedRNG[18])|(((m[24]&~m[202]&~m[302])|(~m[24]&m[202]&m[302]))&~BiasedRNG[18])|((~m[24]&~m[202]&m[302])|(m[24]&~m[202]&m[302])|(m[24]&m[202]&m[302]))):InitCond[38];
    m[85] = run?((((~m[24]&~m[212]&~m[312])|(m[24]&m[212]&~m[312]))&BiasedRNG[19])|(((m[24]&~m[212]&~m[312])|(~m[24]&m[212]&m[312]))&~BiasedRNG[19])|((~m[24]&~m[212]&m[312])|(m[24]&~m[212]&m[312])|(m[24]&m[212]&m[312]))):InitCond[39];
    m[86] = run?((((~m[25]&~m[222]&~m[322])|(m[25]&m[222]&~m[322]))&BiasedRNG[20])|(((m[25]&~m[222]&~m[322])|(~m[25]&m[222]&m[322]))&~BiasedRNG[20])|((~m[25]&~m[222]&m[322])|(m[25]&~m[222]&m[322])|(m[25]&m[222]&m[322]))):InitCond[40];
    m[87] = run?((((~m[25]&~m[232]&~m[332])|(m[25]&m[232]&~m[332]))&BiasedRNG[21])|(((m[25]&~m[232]&~m[332])|(~m[25]&m[232]&m[332]))&~BiasedRNG[21])|((~m[25]&~m[232]&m[332])|(m[25]&~m[232]&m[332])|(m[25]&m[232]&m[332]))):InitCond[41];
    m[88] = run?((((~m[25]&~m[242]&~m[342])|(m[25]&m[242]&~m[342]))&BiasedRNG[22])|(((m[25]&~m[242]&~m[342])|(~m[25]&m[242]&m[342]))&~BiasedRNG[22])|((~m[25]&~m[242]&m[342])|(m[25]&~m[242]&m[342])|(m[25]&m[242]&m[342]))):InitCond[42];
    m[89] = run?((((~m[25]&~m[252]&~m[352])|(m[25]&m[252]&~m[352]))&BiasedRNG[23])|(((m[25]&~m[252]&~m[352])|(~m[25]&m[252]&m[352]))&~BiasedRNG[23])|((~m[25]&~m[252]&m[352])|(m[25]&~m[252]&m[352])|(m[25]&m[252]&m[352]))):InitCond[43];
    m[92] = run?((((~m[26]&~m[183]&~m[283])|(m[26]&m[183]&~m[283]))&BiasedRNG[24])|(((m[26]&~m[183]&~m[283])|(~m[26]&m[183]&m[283]))&~BiasedRNG[24])|((~m[26]&~m[183]&m[283])|(m[26]&~m[183]&m[283])|(m[26]&m[183]&m[283]))):InitCond[44];
    m[93] = run?((((~m[26]&~m[193]&~m[293])|(m[26]&m[193]&~m[293]))&BiasedRNG[25])|(((m[26]&~m[193]&~m[293])|(~m[26]&m[193]&m[293]))&~BiasedRNG[25])|((~m[26]&~m[193]&m[293])|(m[26]&~m[193]&m[293])|(m[26]&m[193]&m[293]))):InitCond[45];
    m[94] = run?((((~m[26]&~m[203]&~m[303])|(m[26]&m[203]&~m[303]))&BiasedRNG[26])|(((m[26]&~m[203]&~m[303])|(~m[26]&m[203]&m[303]))&~BiasedRNG[26])|((~m[26]&~m[203]&m[303])|(m[26]&~m[203]&m[303])|(m[26]&m[203]&m[303]))):InitCond[46];
    m[95] = run?((((~m[26]&~m[213]&~m[313])|(m[26]&m[213]&~m[313]))&BiasedRNG[27])|(((m[26]&~m[213]&~m[313])|(~m[26]&m[213]&m[313]))&~BiasedRNG[27])|((~m[26]&~m[213]&m[313])|(m[26]&~m[213]&m[313])|(m[26]&m[213]&m[313]))):InitCond[47];
    m[96] = run?((((~m[27]&~m[223]&~m[323])|(m[27]&m[223]&~m[323]))&BiasedRNG[28])|(((m[27]&~m[223]&~m[323])|(~m[27]&m[223]&m[323]))&~BiasedRNG[28])|((~m[27]&~m[223]&m[323])|(m[27]&~m[223]&m[323])|(m[27]&m[223]&m[323]))):InitCond[48];
    m[97] = run?((((~m[27]&~m[233]&~m[333])|(m[27]&m[233]&~m[333]))&BiasedRNG[29])|(((m[27]&~m[233]&~m[333])|(~m[27]&m[233]&m[333]))&~BiasedRNG[29])|((~m[27]&~m[233]&m[333])|(m[27]&~m[233]&m[333])|(m[27]&m[233]&m[333]))):InitCond[49];
    m[98] = run?((((~m[27]&~m[243]&~m[343])|(m[27]&m[243]&~m[343]))&BiasedRNG[30])|(((m[27]&~m[243]&~m[343])|(~m[27]&m[243]&m[343]))&~BiasedRNG[30])|((~m[27]&~m[243]&m[343])|(m[27]&~m[243]&m[343])|(m[27]&m[243]&m[343]))):InitCond[50];
    m[99] = run?((((~m[27]&~m[253]&~m[353])|(m[27]&m[253]&~m[353]))&BiasedRNG[31])|(((m[27]&~m[253]&~m[353])|(~m[27]&m[253]&m[353]))&~BiasedRNG[31])|((~m[27]&~m[253]&m[353])|(m[27]&~m[253]&m[353])|(m[27]&m[253]&m[353]))):InitCond[51];
    m[102] = run?((((~m[28]&~m[184]&~m[284])|(m[28]&m[184]&~m[284]))&BiasedRNG[32])|(((m[28]&~m[184]&~m[284])|(~m[28]&m[184]&m[284]))&~BiasedRNG[32])|((~m[28]&~m[184]&m[284])|(m[28]&~m[184]&m[284])|(m[28]&m[184]&m[284]))):InitCond[52];
    m[103] = run?((((~m[28]&~m[194]&~m[294])|(m[28]&m[194]&~m[294]))&BiasedRNG[33])|(((m[28]&~m[194]&~m[294])|(~m[28]&m[194]&m[294]))&~BiasedRNG[33])|((~m[28]&~m[194]&m[294])|(m[28]&~m[194]&m[294])|(m[28]&m[194]&m[294]))):InitCond[53];
    m[104] = run?((((~m[28]&~m[204]&~m[304])|(m[28]&m[204]&~m[304]))&BiasedRNG[34])|(((m[28]&~m[204]&~m[304])|(~m[28]&m[204]&m[304]))&~BiasedRNG[34])|((~m[28]&~m[204]&m[304])|(m[28]&~m[204]&m[304])|(m[28]&m[204]&m[304]))):InitCond[54];
    m[105] = run?((((~m[28]&~m[214]&~m[314])|(m[28]&m[214]&~m[314]))&BiasedRNG[35])|(((m[28]&~m[214]&~m[314])|(~m[28]&m[214]&m[314]))&~BiasedRNG[35])|((~m[28]&~m[214]&m[314])|(m[28]&~m[214]&m[314])|(m[28]&m[214]&m[314]))):InitCond[55];
    m[106] = run?((((~m[29]&~m[224]&~m[324])|(m[29]&m[224]&~m[324]))&BiasedRNG[36])|(((m[29]&~m[224]&~m[324])|(~m[29]&m[224]&m[324]))&~BiasedRNG[36])|((~m[29]&~m[224]&m[324])|(m[29]&~m[224]&m[324])|(m[29]&m[224]&m[324]))):InitCond[56];
    m[107] = run?((((~m[29]&~m[234]&~m[334])|(m[29]&m[234]&~m[334]))&BiasedRNG[37])|(((m[29]&~m[234]&~m[334])|(~m[29]&m[234]&m[334]))&~BiasedRNG[37])|((~m[29]&~m[234]&m[334])|(m[29]&~m[234]&m[334])|(m[29]&m[234]&m[334]))):InitCond[57];
    m[108] = run?((((~m[29]&~m[244]&~m[344])|(m[29]&m[244]&~m[344]))&BiasedRNG[38])|(((m[29]&~m[244]&~m[344])|(~m[29]&m[244]&m[344]))&~BiasedRNG[38])|((~m[29]&~m[244]&m[344])|(m[29]&~m[244]&m[344])|(m[29]&m[244]&m[344]))):InitCond[58];
    m[109] = run?((((~m[29]&~m[254]&~m[354])|(m[29]&m[254]&~m[354]))&BiasedRNG[39])|(((m[29]&~m[254]&~m[354])|(~m[29]&m[254]&m[354]))&~BiasedRNG[39])|((~m[29]&~m[254]&m[354])|(m[29]&~m[254]&m[354])|(m[29]&m[254]&m[354]))):InitCond[59];
    m[112] = run?((((~m[30]&~m[185]&~m[285])|(m[30]&m[185]&~m[285]))&BiasedRNG[40])|(((m[30]&~m[185]&~m[285])|(~m[30]&m[185]&m[285]))&~BiasedRNG[40])|((~m[30]&~m[185]&m[285])|(m[30]&~m[185]&m[285])|(m[30]&m[185]&m[285]))):InitCond[60];
    m[113] = run?((((~m[30]&~m[195]&~m[295])|(m[30]&m[195]&~m[295]))&BiasedRNG[41])|(((m[30]&~m[195]&~m[295])|(~m[30]&m[195]&m[295]))&~BiasedRNG[41])|((~m[30]&~m[195]&m[295])|(m[30]&~m[195]&m[295])|(m[30]&m[195]&m[295]))):InitCond[61];
    m[114] = run?((((~m[30]&~m[205]&~m[305])|(m[30]&m[205]&~m[305]))&BiasedRNG[42])|(((m[30]&~m[205]&~m[305])|(~m[30]&m[205]&m[305]))&~BiasedRNG[42])|((~m[30]&~m[205]&m[305])|(m[30]&~m[205]&m[305])|(m[30]&m[205]&m[305]))):InitCond[62];
    m[115] = run?((((~m[30]&~m[215]&~m[315])|(m[30]&m[215]&~m[315]))&BiasedRNG[43])|(((m[30]&~m[215]&~m[315])|(~m[30]&m[215]&m[315]))&~BiasedRNG[43])|((~m[30]&~m[215]&m[315])|(m[30]&~m[215]&m[315])|(m[30]&m[215]&m[315]))):InitCond[63];
    m[116] = run?((((~m[31]&~m[225]&~m[325])|(m[31]&m[225]&~m[325]))&BiasedRNG[44])|(((m[31]&~m[225]&~m[325])|(~m[31]&m[225]&m[325]))&~BiasedRNG[44])|((~m[31]&~m[225]&m[325])|(m[31]&~m[225]&m[325])|(m[31]&m[225]&m[325]))):InitCond[64];
    m[117] = run?((((~m[31]&~m[235]&~m[335])|(m[31]&m[235]&~m[335]))&BiasedRNG[45])|(((m[31]&~m[235]&~m[335])|(~m[31]&m[235]&m[335]))&~BiasedRNG[45])|((~m[31]&~m[235]&m[335])|(m[31]&~m[235]&m[335])|(m[31]&m[235]&m[335]))):InitCond[65];
    m[118] = run?((((~m[31]&~m[245]&~m[345])|(m[31]&m[245]&~m[345]))&BiasedRNG[46])|(((m[31]&~m[245]&~m[345])|(~m[31]&m[245]&m[345]))&~BiasedRNG[46])|((~m[31]&~m[245]&m[345])|(m[31]&~m[245]&m[345])|(m[31]&m[245]&m[345]))):InitCond[66];
    m[119] = run?((((~m[31]&~m[255]&~m[355])|(m[31]&m[255]&~m[355]))&BiasedRNG[47])|(((m[31]&~m[255]&~m[355])|(~m[31]&m[255]&m[355]))&~BiasedRNG[47])|((~m[31]&~m[255]&m[355])|(m[31]&~m[255]&m[355])|(m[31]&m[255]&m[355]))):InitCond[67];
    m[122] = run?((((~m[32]&~m[186]&~m[286])|(m[32]&m[186]&~m[286]))&BiasedRNG[48])|(((m[32]&~m[186]&~m[286])|(~m[32]&m[186]&m[286]))&~BiasedRNG[48])|((~m[32]&~m[186]&m[286])|(m[32]&~m[186]&m[286])|(m[32]&m[186]&m[286]))):InitCond[68];
    m[123] = run?((((~m[32]&~m[196]&~m[296])|(m[32]&m[196]&~m[296]))&BiasedRNG[49])|(((m[32]&~m[196]&~m[296])|(~m[32]&m[196]&m[296]))&~BiasedRNG[49])|((~m[32]&~m[196]&m[296])|(m[32]&~m[196]&m[296])|(m[32]&m[196]&m[296]))):InitCond[69];
    m[124] = run?((((~m[32]&~m[206]&~m[306])|(m[32]&m[206]&~m[306]))&BiasedRNG[50])|(((m[32]&~m[206]&~m[306])|(~m[32]&m[206]&m[306]))&~BiasedRNG[50])|((~m[32]&~m[206]&m[306])|(m[32]&~m[206]&m[306])|(m[32]&m[206]&m[306]))):InitCond[70];
    m[125] = run?((((~m[32]&~m[216]&~m[316])|(m[32]&m[216]&~m[316]))&BiasedRNG[51])|(((m[32]&~m[216]&~m[316])|(~m[32]&m[216]&m[316]))&~BiasedRNG[51])|((~m[32]&~m[216]&m[316])|(m[32]&~m[216]&m[316])|(m[32]&m[216]&m[316]))):InitCond[71];
    m[126] = run?((((~m[33]&~m[226]&~m[326])|(m[33]&m[226]&~m[326]))&BiasedRNG[52])|(((m[33]&~m[226]&~m[326])|(~m[33]&m[226]&m[326]))&~BiasedRNG[52])|((~m[33]&~m[226]&m[326])|(m[33]&~m[226]&m[326])|(m[33]&m[226]&m[326]))):InitCond[72];
    m[127] = run?((((~m[33]&~m[236]&~m[336])|(m[33]&m[236]&~m[336]))&BiasedRNG[53])|(((m[33]&~m[236]&~m[336])|(~m[33]&m[236]&m[336]))&~BiasedRNG[53])|((~m[33]&~m[236]&m[336])|(m[33]&~m[236]&m[336])|(m[33]&m[236]&m[336]))):InitCond[73];
    m[128] = run?((((~m[33]&~m[246]&~m[346])|(m[33]&m[246]&~m[346]))&BiasedRNG[54])|(((m[33]&~m[246]&~m[346])|(~m[33]&m[246]&m[346]))&~BiasedRNG[54])|((~m[33]&~m[246]&m[346])|(m[33]&~m[246]&m[346])|(m[33]&m[246]&m[346]))):InitCond[74];
    m[129] = run?((((~m[33]&~m[256]&~m[356])|(m[33]&m[256]&~m[356]))&BiasedRNG[55])|(((m[33]&~m[256]&~m[356])|(~m[33]&m[256]&m[356]))&~BiasedRNG[55])|((~m[33]&~m[256]&m[356])|(m[33]&~m[256]&m[356])|(m[33]&m[256]&m[356]))):InitCond[75];
    m[132] = run?((((~m[34]&~m[187]&~m[287])|(m[34]&m[187]&~m[287]))&BiasedRNG[56])|(((m[34]&~m[187]&~m[287])|(~m[34]&m[187]&m[287]))&~BiasedRNG[56])|((~m[34]&~m[187]&m[287])|(m[34]&~m[187]&m[287])|(m[34]&m[187]&m[287]))):InitCond[76];
    m[133] = run?((((~m[34]&~m[197]&~m[297])|(m[34]&m[197]&~m[297]))&BiasedRNG[57])|(((m[34]&~m[197]&~m[297])|(~m[34]&m[197]&m[297]))&~BiasedRNG[57])|((~m[34]&~m[197]&m[297])|(m[34]&~m[197]&m[297])|(m[34]&m[197]&m[297]))):InitCond[77];
    m[134] = run?((((~m[34]&~m[207]&~m[307])|(m[34]&m[207]&~m[307]))&BiasedRNG[58])|(((m[34]&~m[207]&~m[307])|(~m[34]&m[207]&m[307]))&~BiasedRNG[58])|((~m[34]&~m[207]&m[307])|(m[34]&~m[207]&m[307])|(m[34]&m[207]&m[307]))):InitCond[78];
    m[135] = run?((((~m[34]&~m[217]&~m[317])|(m[34]&m[217]&~m[317]))&BiasedRNG[59])|(((m[34]&~m[217]&~m[317])|(~m[34]&m[217]&m[317]))&~BiasedRNG[59])|((~m[34]&~m[217]&m[317])|(m[34]&~m[217]&m[317])|(m[34]&m[217]&m[317]))):InitCond[79];
    m[136] = run?((((~m[35]&~m[227]&~m[327])|(m[35]&m[227]&~m[327]))&BiasedRNG[60])|(((m[35]&~m[227]&~m[327])|(~m[35]&m[227]&m[327]))&~BiasedRNG[60])|((~m[35]&~m[227]&m[327])|(m[35]&~m[227]&m[327])|(m[35]&m[227]&m[327]))):InitCond[80];
    m[137] = run?((((~m[35]&~m[237]&~m[337])|(m[35]&m[237]&~m[337]))&BiasedRNG[61])|(((m[35]&~m[237]&~m[337])|(~m[35]&m[237]&m[337]))&~BiasedRNG[61])|((~m[35]&~m[237]&m[337])|(m[35]&~m[237]&m[337])|(m[35]&m[237]&m[337]))):InitCond[81];
    m[138] = run?((((~m[35]&~m[247]&~m[347])|(m[35]&m[247]&~m[347]))&BiasedRNG[62])|(((m[35]&~m[247]&~m[347])|(~m[35]&m[247]&m[347]))&~BiasedRNG[62])|((~m[35]&~m[247]&m[347])|(m[35]&~m[247]&m[347])|(m[35]&m[247]&m[347]))):InitCond[82];
    m[139] = run?((((~m[35]&~m[257]&~m[357])|(m[35]&m[257]&~m[357]))&BiasedRNG[63])|(((m[35]&~m[257]&~m[357])|(~m[35]&m[257]&m[357]))&~BiasedRNG[63])|((~m[35]&~m[257]&m[357])|(m[35]&~m[257]&m[357])|(m[35]&m[257]&m[357]))):InitCond[83];
    m[142] = run?((((~m[36]&~m[188]&~m[288])|(m[36]&m[188]&~m[288]))&BiasedRNG[64])|(((m[36]&~m[188]&~m[288])|(~m[36]&m[188]&m[288]))&~BiasedRNG[64])|((~m[36]&~m[188]&m[288])|(m[36]&~m[188]&m[288])|(m[36]&m[188]&m[288]))):InitCond[84];
    m[143] = run?((((~m[36]&~m[198]&~m[298])|(m[36]&m[198]&~m[298]))&BiasedRNG[65])|(((m[36]&~m[198]&~m[298])|(~m[36]&m[198]&m[298]))&~BiasedRNG[65])|((~m[36]&~m[198]&m[298])|(m[36]&~m[198]&m[298])|(m[36]&m[198]&m[298]))):InitCond[85];
    m[144] = run?((((~m[36]&~m[208]&~m[308])|(m[36]&m[208]&~m[308]))&BiasedRNG[66])|(((m[36]&~m[208]&~m[308])|(~m[36]&m[208]&m[308]))&~BiasedRNG[66])|((~m[36]&~m[208]&m[308])|(m[36]&~m[208]&m[308])|(m[36]&m[208]&m[308]))):InitCond[86];
    m[145] = run?((((~m[36]&~m[218]&~m[318])|(m[36]&m[218]&~m[318]))&BiasedRNG[67])|(((m[36]&~m[218]&~m[318])|(~m[36]&m[218]&m[318]))&~BiasedRNG[67])|((~m[36]&~m[218]&m[318])|(m[36]&~m[218]&m[318])|(m[36]&m[218]&m[318]))):InitCond[87];
    m[146] = run?((((~m[37]&~m[228]&~m[328])|(m[37]&m[228]&~m[328]))&BiasedRNG[68])|(((m[37]&~m[228]&~m[328])|(~m[37]&m[228]&m[328]))&~BiasedRNG[68])|((~m[37]&~m[228]&m[328])|(m[37]&~m[228]&m[328])|(m[37]&m[228]&m[328]))):InitCond[88];
    m[147] = run?((((~m[37]&~m[238]&~m[338])|(m[37]&m[238]&~m[338]))&BiasedRNG[69])|(((m[37]&~m[238]&~m[338])|(~m[37]&m[238]&m[338]))&~BiasedRNG[69])|((~m[37]&~m[238]&m[338])|(m[37]&~m[238]&m[338])|(m[37]&m[238]&m[338]))):InitCond[89];
    m[148] = run?((((~m[37]&~m[248]&~m[348])|(m[37]&m[248]&~m[348]))&BiasedRNG[70])|(((m[37]&~m[248]&~m[348])|(~m[37]&m[248]&m[348]))&~BiasedRNG[70])|((~m[37]&~m[248]&m[348])|(m[37]&~m[248]&m[348])|(m[37]&m[248]&m[348]))):InitCond[90];
    m[149] = run?((((~m[37]&~m[258]&~m[358])|(m[37]&m[258]&~m[358]))&BiasedRNG[71])|(((m[37]&~m[258]&~m[358])|(~m[37]&m[258]&m[358]))&~BiasedRNG[71])|((~m[37]&~m[258]&m[358])|(m[37]&~m[258]&m[358])|(m[37]&m[258]&m[358]))):InitCond[91];
    m[152] = run?((((~m[38]&~m[189]&~m[289])|(m[38]&m[189]&~m[289]))&BiasedRNG[72])|(((m[38]&~m[189]&~m[289])|(~m[38]&m[189]&m[289]))&~BiasedRNG[72])|((~m[38]&~m[189]&m[289])|(m[38]&~m[189]&m[289])|(m[38]&m[189]&m[289]))):InitCond[92];
    m[153] = run?((((~m[38]&~m[199]&~m[299])|(m[38]&m[199]&~m[299]))&BiasedRNG[73])|(((m[38]&~m[199]&~m[299])|(~m[38]&m[199]&m[299]))&~BiasedRNG[73])|((~m[38]&~m[199]&m[299])|(m[38]&~m[199]&m[299])|(m[38]&m[199]&m[299]))):InitCond[93];
    m[154] = run?((((~m[38]&~m[209]&~m[309])|(m[38]&m[209]&~m[309]))&BiasedRNG[74])|(((m[38]&~m[209]&~m[309])|(~m[38]&m[209]&m[309]))&~BiasedRNG[74])|((~m[38]&~m[209]&m[309])|(m[38]&~m[209]&m[309])|(m[38]&m[209]&m[309]))):InitCond[94];
    m[155] = run?((((~m[38]&~m[219]&~m[319])|(m[38]&m[219]&~m[319]))&BiasedRNG[75])|(((m[38]&~m[219]&~m[319])|(~m[38]&m[219]&m[319]))&~BiasedRNG[75])|((~m[38]&~m[219]&m[319])|(m[38]&~m[219]&m[319])|(m[38]&m[219]&m[319]))):InitCond[95];
    m[156] = run?((((~m[39]&~m[229]&~m[329])|(m[39]&m[229]&~m[329]))&BiasedRNG[76])|(((m[39]&~m[229]&~m[329])|(~m[39]&m[229]&m[329]))&~BiasedRNG[76])|((~m[39]&~m[229]&m[329])|(m[39]&~m[229]&m[329])|(m[39]&m[229]&m[329]))):InitCond[96];
    m[157] = run?((((~m[39]&~m[239]&~m[339])|(m[39]&m[239]&~m[339]))&BiasedRNG[77])|(((m[39]&~m[239]&~m[339])|(~m[39]&m[239]&m[339]))&~BiasedRNG[77])|((~m[39]&~m[239]&m[339])|(m[39]&~m[239]&m[339])|(m[39]&m[239]&m[339]))):InitCond[97];
    m[158] = run?((((~m[39]&~m[249]&~m[349])|(m[39]&m[249]&~m[349]))&BiasedRNG[78])|(((m[39]&~m[249]&~m[349])|(~m[39]&m[249]&m[349]))&~BiasedRNG[78])|((~m[39]&~m[249]&m[349])|(m[39]&~m[249]&m[349])|(m[39]&m[249]&m[349]))):InitCond[98];
    m[159] = run?((((~m[39]&~m[259]&~m[359])|(m[39]&m[259]&~m[359]))&BiasedRNG[79])|(((m[39]&~m[259]&~m[359])|(~m[39]&m[259]&m[359]))&~BiasedRNG[79])|((~m[39]&~m[259]&m[359])|(m[39]&~m[259]&m[359])|(m[39]&m[259]&m[359]))):InitCond[99];
    m[162] = run?((((~m[40]&~m[80]&~m[262])|(m[40]&m[80]&~m[262]))&BiasedRNG[80])|(((m[40]&~m[80]&~m[262])|(~m[40]&m[80]&m[262]))&~BiasedRNG[80])|((~m[40]&~m[80]&m[262])|(m[40]&~m[80]&m[262])|(m[40]&m[80]&m[262]))):InitCond[100];
    m[163] = run?((((~m[40]&~m[90]&~m[263])|(m[40]&m[90]&~m[263]))&BiasedRNG[81])|(((m[40]&~m[90]&~m[263])|(~m[40]&m[90]&m[263]))&~BiasedRNG[81])|((~m[40]&~m[90]&m[263])|(m[40]&~m[90]&m[263])|(m[40]&m[90]&m[263]))):InitCond[101];
    m[164] = run?((((~m[40]&~m[100]&~m[264])|(m[40]&m[100]&~m[264]))&BiasedRNG[82])|(((m[40]&~m[100]&~m[264])|(~m[40]&m[100]&m[264]))&~BiasedRNG[82])|((~m[40]&~m[100]&m[264])|(m[40]&~m[100]&m[264])|(m[40]&m[100]&m[264]))):InitCond[102];
    m[165] = run?((((~m[40]&~m[110]&~m[265])|(m[40]&m[110]&~m[265]))&BiasedRNG[83])|(((m[40]&~m[110]&~m[265])|(~m[40]&m[110]&m[265]))&~BiasedRNG[83])|((~m[40]&~m[110]&m[265])|(m[40]&~m[110]&m[265])|(m[40]&m[110]&m[265]))):InitCond[103];
    m[166] = run?((((~m[41]&~m[120]&~m[266])|(m[41]&m[120]&~m[266]))&BiasedRNG[84])|(((m[41]&~m[120]&~m[266])|(~m[41]&m[120]&m[266]))&~BiasedRNG[84])|((~m[41]&~m[120]&m[266])|(m[41]&~m[120]&m[266])|(m[41]&m[120]&m[266]))):InitCond[104];
    m[167] = run?((((~m[41]&~m[130]&~m[267])|(m[41]&m[130]&~m[267]))&BiasedRNG[85])|(((m[41]&~m[130]&~m[267])|(~m[41]&m[130]&m[267]))&~BiasedRNG[85])|((~m[41]&~m[130]&m[267])|(m[41]&~m[130]&m[267])|(m[41]&m[130]&m[267]))):InitCond[105];
    m[168] = run?((((~m[41]&~m[140]&~m[268])|(m[41]&m[140]&~m[268]))&BiasedRNG[86])|(((m[41]&~m[140]&~m[268])|(~m[41]&m[140]&m[268]))&~BiasedRNG[86])|((~m[41]&~m[140]&m[268])|(m[41]&~m[140]&m[268])|(m[41]&m[140]&m[268]))):InitCond[106];
    m[169] = run?((((~m[41]&~m[150]&~m[269])|(m[41]&m[150]&~m[269]))&BiasedRNG[87])|(((m[41]&~m[150]&~m[269])|(~m[41]&m[150]&m[269]))&~BiasedRNG[87])|((~m[41]&~m[150]&m[269])|(m[41]&~m[150]&m[269])|(m[41]&m[150]&m[269]))):InitCond[107];
    m[172] = run?((((~m[42]&~m[81]&~m[272])|(m[42]&m[81]&~m[272]))&BiasedRNG[88])|(((m[42]&~m[81]&~m[272])|(~m[42]&m[81]&m[272]))&~BiasedRNG[88])|((~m[42]&~m[81]&m[272])|(m[42]&~m[81]&m[272])|(m[42]&m[81]&m[272]))):InitCond[108];
    m[173] = run?((((~m[42]&~m[91]&~m[273])|(m[42]&m[91]&~m[273]))&BiasedRNG[89])|(((m[42]&~m[91]&~m[273])|(~m[42]&m[91]&m[273]))&~BiasedRNG[89])|((~m[42]&~m[91]&m[273])|(m[42]&~m[91]&m[273])|(m[42]&m[91]&m[273]))):InitCond[109];
    m[174] = run?((((~m[42]&~m[101]&~m[274])|(m[42]&m[101]&~m[274]))&BiasedRNG[90])|(((m[42]&~m[101]&~m[274])|(~m[42]&m[101]&m[274]))&~BiasedRNG[90])|((~m[42]&~m[101]&m[274])|(m[42]&~m[101]&m[274])|(m[42]&m[101]&m[274]))):InitCond[110];
    m[175] = run?((((~m[42]&~m[111]&~m[275])|(m[42]&m[111]&~m[275]))&BiasedRNG[91])|(((m[42]&~m[111]&~m[275])|(~m[42]&m[111]&m[275]))&~BiasedRNG[91])|((~m[42]&~m[111]&m[275])|(m[42]&~m[111]&m[275])|(m[42]&m[111]&m[275]))):InitCond[111];
    m[176] = run?((((~m[43]&~m[121]&~m[276])|(m[43]&m[121]&~m[276]))&BiasedRNG[92])|(((m[43]&~m[121]&~m[276])|(~m[43]&m[121]&m[276]))&~BiasedRNG[92])|((~m[43]&~m[121]&m[276])|(m[43]&~m[121]&m[276])|(m[43]&m[121]&m[276]))):InitCond[112];
    m[177] = run?((((~m[43]&~m[131]&~m[277])|(m[43]&m[131]&~m[277]))&BiasedRNG[93])|(((m[43]&~m[131]&~m[277])|(~m[43]&m[131]&m[277]))&~BiasedRNG[93])|((~m[43]&~m[131]&m[277])|(m[43]&~m[131]&m[277])|(m[43]&m[131]&m[277]))):InitCond[113];
    m[178] = run?((((~m[43]&~m[141]&~m[278])|(m[43]&m[141]&~m[278]))&BiasedRNG[94])|(((m[43]&~m[141]&~m[278])|(~m[43]&m[141]&m[278]))&~BiasedRNG[94])|((~m[43]&~m[141]&m[278])|(m[43]&~m[141]&m[278])|(m[43]&m[141]&m[278]))):InitCond[114];
    m[179] = run?((((~m[43]&~m[151]&~m[279])|(m[43]&m[151]&~m[279]))&BiasedRNG[95])|(((m[43]&~m[151]&~m[279])|(~m[43]&m[151]&m[279]))&~BiasedRNG[95])|((~m[43]&~m[151]&m[279])|(m[43]&~m[151]&m[279])|(m[43]&m[151]&m[279]))):InitCond[115];
    m[261] = run?((((m[70]&~m[161]&m[360])|(~m[70]&m[161]&m[360]))&BiasedRNG[96])|(((m[70]&m[161]&~m[360]))&~BiasedRNG[96])|((m[70]&m[161]&m[360]))):InitCond[116];
    m[270] = run?((((m[61]&~m[170]&m[361])|(~m[61]&m[170]&m[361]))&BiasedRNG[97])|(((m[61]&m[170]&~m[361]))&~BiasedRNG[97])|((m[61]&m[170]&m[361]))):InitCond[117];
    m[271] = run?((((m[71]&~m[171]&m[366])|(~m[71]&m[171]&m[366]))&BiasedRNG[98])|(((m[71]&m[171]&~m[366]))&~BiasedRNG[98])|((m[71]&m[171]&m[366]))):InitCond[118];
    m[365] = run?((((m[262]&~m[366]&~m[367]&~m[368]&~m[369])|(~m[262]&~m[366]&~m[367]&m[368]&~m[369])|(m[262]&m[366]&~m[367]&m[368]&~m[369])|(m[262]&~m[366]&m[367]&m[368]&~m[369])|(~m[262]&m[366]&~m[367]&~m[368]&m[369])|(~m[262]&~m[366]&m[367]&~m[368]&m[369])|(m[262]&m[366]&m[367]&~m[368]&m[369])|(~m[262]&m[366]&m[367]&m[368]&m[369]))&UnbiasedRNG[20])|((m[262]&~m[366]&~m[367]&m[368]&~m[369])|(~m[262]&~m[366]&~m[367]&~m[368]&m[369])|(m[262]&~m[366]&~m[367]&~m[368]&m[369])|(m[262]&m[366]&~m[367]&~m[368]&m[369])|(m[262]&~m[366]&m[367]&~m[368]&m[369])|(~m[262]&~m[366]&~m[367]&m[368]&m[369])|(m[262]&~m[366]&~m[367]&m[368]&m[369])|(~m[262]&m[366]&~m[367]&m[368]&m[369])|(m[262]&m[366]&~m[367]&m[368]&m[369])|(~m[262]&~m[366]&m[367]&m[368]&m[369])|(m[262]&~m[366]&m[367]&m[368]&m[369])|(m[262]&m[366]&m[367]&m[368]&m[369]))):InitCond[119];
    m[370] = run?((((m[368]&~m[371]&~m[372]&~m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&m[373]&~m[374])|(m[368]&m[371]&~m[372]&m[373]&~m[374])|(m[368]&~m[371]&m[372]&m[373]&~m[374])|(~m[368]&m[371]&~m[372]&~m[373]&m[374])|(~m[368]&~m[371]&m[372]&~m[373]&m[374])|(m[368]&m[371]&m[372]&~m[373]&m[374])|(~m[368]&m[371]&m[372]&m[373]&m[374]))&UnbiasedRNG[21])|((m[368]&~m[371]&~m[372]&m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&m[372]&~m[373]&m[374])|(~m[368]&~m[371]&~m[372]&m[373]&m[374])|(m[368]&~m[371]&~m[372]&m[373]&m[374])|(~m[368]&m[371]&~m[372]&m[373]&m[374])|(m[368]&m[371]&~m[372]&m[373]&m[374])|(~m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&m[371]&m[372]&m[373]&m[374]))):InitCond[120];
    m[375] = run?((((m[263]&~m[376]&~m[377]&~m[378]&~m[379])|(~m[263]&~m[376]&~m[377]&m[378]&~m[379])|(m[263]&m[376]&~m[377]&m[378]&~m[379])|(m[263]&~m[376]&m[377]&m[378]&~m[379])|(~m[263]&m[376]&~m[377]&~m[378]&m[379])|(~m[263]&~m[376]&m[377]&~m[378]&m[379])|(m[263]&m[376]&m[377]&~m[378]&m[379])|(~m[263]&m[376]&m[377]&m[378]&m[379]))&UnbiasedRNG[22])|((m[263]&~m[376]&~m[377]&m[378]&~m[379])|(~m[263]&~m[376]&~m[377]&~m[378]&m[379])|(m[263]&~m[376]&~m[377]&~m[378]&m[379])|(m[263]&m[376]&~m[377]&~m[378]&m[379])|(m[263]&~m[376]&m[377]&~m[378]&m[379])|(~m[263]&~m[376]&~m[377]&m[378]&m[379])|(m[263]&~m[376]&~m[377]&m[378]&m[379])|(~m[263]&m[376]&~m[377]&m[378]&m[379])|(m[263]&m[376]&~m[377]&m[378]&m[379])|(~m[263]&~m[376]&m[377]&m[378]&m[379])|(m[263]&~m[376]&m[377]&m[378]&m[379])|(m[263]&m[376]&m[377]&m[378]&m[379]))):InitCond[121];
    m[380] = run?((((m[378]&~m[381]&~m[382]&~m[383]&~m[384])|(~m[378]&~m[381]&~m[382]&m[383]&~m[384])|(m[378]&m[381]&~m[382]&m[383]&~m[384])|(m[378]&~m[381]&m[382]&m[383]&~m[384])|(~m[378]&m[381]&~m[382]&~m[383]&m[384])|(~m[378]&~m[381]&m[382]&~m[383]&m[384])|(m[378]&m[381]&m[382]&~m[383]&m[384])|(~m[378]&m[381]&m[382]&m[383]&m[384]))&UnbiasedRNG[23])|((m[378]&~m[381]&~m[382]&m[383]&~m[384])|(~m[378]&~m[381]&~m[382]&~m[383]&m[384])|(m[378]&~m[381]&~m[382]&~m[383]&m[384])|(m[378]&m[381]&~m[382]&~m[383]&m[384])|(m[378]&~m[381]&m[382]&~m[383]&m[384])|(~m[378]&~m[381]&~m[382]&m[383]&m[384])|(m[378]&~m[381]&~m[382]&m[383]&m[384])|(~m[378]&m[381]&~m[382]&m[383]&m[384])|(m[378]&m[381]&~m[382]&m[383]&m[384])|(~m[378]&~m[381]&m[382]&m[383]&m[384])|(m[378]&~m[381]&m[382]&m[383]&m[384])|(m[378]&m[381]&m[382]&m[383]&m[384]))):InitCond[122];
    m[385] = run?((((m[383]&~m[386]&~m[387]&~m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&m[388]&~m[389])|(m[383]&m[386]&~m[387]&m[388]&~m[389])|(m[383]&~m[386]&m[387]&m[388]&~m[389])|(~m[383]&m[386]&~m[387]&~m[388]&m[389])|(~m[383]&~m[386]&m[387]&~m[388]&m[389])|(m[383]&m[386]&m[387]&~m[388]&m[389])|(~m[383]&m[386]&m[387]&m[388]&m[389]))&UnbiasedRNG[24])|((m[383]&~m[386]&~m[387]&m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&m[387]&~m[388]&m[389])|(~m[383]&~m[386]&~m[387]&m[388]&m[389])|(m[383]&~m[386]&~m[387]&m[388]&m[389])|(~m[383]&m[386]&~m[387]&m[388]&m[389])|(m[383]&m[386]&~m[387]&m[388]&m[389])|(~m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&m[386]&m[387]&m[388]&m[389]))):InitCond[123];
    m[390] = run?((((m[264]&~m[391]&~m[392]&~m[393]&~m[394])|(~m[264]&~m[391]&~m[392]&m[393]&~m[394])|(m[264]&m[391]&~m[392]&m[393]&~m[394])|(m[264]&~m[391]&m[392]&m[393]&~m[394])|(~m[264]&m[391]&~m[392]&~m[393]&m[394])|(~m[264]&~m[391]&m[392]&~m[393]&m[394])|(m[264]&m[391]&m[392]&~m[393]&m[394])|(~m[264]&m[391]&m[392]&m[393]&m[394]))&UnbiasedRNG[25])|((m[264]&~m[391]&~m[392]&m[393]&~m[394])|(~m[264]&~m[391]&~m[392]&~m[393]&m[394])|(m[264]&~m[391]&~m[392]&~m[393]&m[394])|(m[264]&m[391]&~m[392]&~m[393]&m[394])|(m[264]&~m[391]&m[392]&~m[393]&m[394])|(~m[264]&~m[391]&~m[392]&m[393]&m[394])|(m[264]&~m[391]&~m[392]&m[393]&m[394])|(~m[264]&m[391]&~m[392]&m[393]&m[394])|(m[264]&m[391]&~m[392]&m[393]&m[394])|(~m[264]&~m[391]&m[392]&m[393]&m[394])|(m[264]&~m[391]&m[392]&m[393]&m[394])|(m[264]&m[391]&m[392]&m[393]&m[394]))):InitCond[124];
    m[395] = run?((((m[393]&~m[396]&~m[397]&~m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&m[398]&~m[399])|(m[393]&m[396]&~m[397]&m[398]&~m[399])|(m[393]&~m[396]&m[397]&m[398]&~m[399])|(~m[393]&m[396]&~m[397]&~m[398]&m[399])|(~m[393]&~m[396]&m[397]&~m[398]&m[399])|(m[393]&m[396]&m[397]&~m[398]&m[399])|(~m[393]&m[396]&m[397]&m[398]&m[399]))&UnbiasedRNG[26])|((m[393]&~m[396]&~m[397]&m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&m[397]&~m[398]&m[399])|(~m[393]&~m[396]&~m[397]&m[398]&m[399])|(m[393]&~m[396]&~m[397]&m[398]&m[399])|(~m[393]&m[396]&~m[397]&m[398]&m[399])|(m[393]&m[396]&~m[397]&m[398]&m[399])|(~m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&m[396]&m[397]&m[398]&m[399]))):InitCond[125];
    m[400] = run?((((m[398]&~m[401]&~m[402]&~m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&m[403]&~m[404])|(m[398]&m[401]&~m[402]&m[403]&~m[404])|(m[398]&~m[401]&m[402]&m[403]&~m[404])|(~m[398]&m[401]&~m[402]&~m[403]&m[404])|(~m[398]&~m[401]&m[402]&~m[403]&m[404])|(m[398]&m[401]&m[402]&~m[403]&m[404])|(~m[398]&m[401]&m[402]&m[403]&m[404]))&UnbiasedRNG[27])|((m[398]&~m[401]&~m[402]&m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&m[402]&~m[403]&m[404])|(~m[398]&~m[401]&~m[402]&m[403]&m[404])|(m[398]&~m[401]&~m[402]&m[403]&m[404])|(~m[398]&m[401]&~m[402]&m[403]&m[404])|(m[398]&m[401]&~m[402]&m[403]&m[404])|(~m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&m[401]&m[402]&m[403]&m[404]))):InitCond[126];
    m[405] = run?((((m[403]&~m[406]&~m[407]&~m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&m[408]&~m[409])|(m[403]&m[406]&~m[407]&m[408]&~m[409])|(m[403]&~m[406]&m[407]&m[408]&~m[409])|(~m[403]&m[406]&~m[407]&~m[408]&m[409])|(~m[403]&~m[406]&m[407]&~m[408]&m[409])|(m[403]&m[406]&m[407]&~m[408]&m[409])|(~m[403]&m[406]&m[407]&m[408]&m[409]))&UnbiasedRNG[28])|((m[403]&~m[406]&~m[407]&m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&m[407]&~m[408]&m[409])|(~m[403]&~m[406]&~m[407]&m[408]&m[409])|(m[403]&~m[406]&~m[407]&m[408]&m[409])|(~m[403]&m[406]&~m[407]&m[408]&m[409])|(m[403]&m[406]&~m[407]&m[408]&m[409])|(~m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&m[406]&m[407]&m[408]&m[409]))):InitCond[127];
    m[410] = run?((((m[265]&~m[411]&~m[412]&~m[413]&~m[414])|(~m[265]&~m[411]&~m[412]&m[413]&~m[414])|(m[265]&m[411]&~m[412]&m[413]&~m[414])|(m[265]&~m[411]&m[412]&m[413]&~m[414])|(~m[265]&m[411]&~m[412]&~m[413]&m[414])|(~m[265]&~m[411]&m[412]&~m[413]&m[414])|(m[265]&m[411]&m[412]&~m[413]&m[414])|(~m[265]&m[411]&m[412]&m[413]&m[414]))&UnbiasedRNG[29])|((m[265]&~m[411]&~m[412]&m[413]&~m[414])|(~m[265]&~m[411]&~m[412]&~m[413]&m[414])|(m[265]&~m[411]&~m[412]&~m[413]&m[414])|(m[265]&m[411]&~m[412]&~m[413]&m[414])|(m[265]&~m[411]&m[412]&~m[413]&m[414])|(~m[265]&~m[411]&~m[412]&m[413]&m[414])|(m[265]&~m[411]&~m[412]&m[413]&m[414])|(~m[265]&m[411]&~m[412]&m[413]&m[414])|(m[265]&m[411]&~m[412]&m[413]&m[414])|(~m[265]&~m[411]&m[412]&m[413]&m[414])|(m[265]&~m[411]&m[412]&m[413]&m[414])|(m[265]&m[411]&m[412]&m[413]&m[414]))):InitCond[128];
    m[415] = run?((((m[413]&~m[416]&~m[417]&~m[418]&~m[419])|(~m[413]&~m[416]&~m[417]&m[418]&~m[419])|(m[413]&m[416]&~m[417]&m[418]&~m[419])|(m[413]&~m[416]&m[417]&m[418]&~m[419])|(~m[413]&m[416]&~m[417]&~m[418]&m[419])|(~m[413]&~m[416]&m[417]&~m[418]&m[419])|(m[413]&m[416]&m[417]&~m[418]&m[419])|(~m[413]&m[416]&m[417]&m[418]&m[419]))&UnbiasedRNG[30])|((m[413]&~m[416]&~m[417]&m[418]&~m[419])|(~m[413]&~m[416]&~m[417]&~m[418]&m[419])|(m[413]&~m[416]&~m[417]&~m[418]&m[419])|(m[413]&m[416]&~m[417]&~m[418]&m[419])|(m[413]&~m[416]&m[417]&~m[418]&m[419])|(~m[413]&~m[416]&~m[417]&m[418]&m[419])|(m[413]&~m[416]&~m[417]&m[418]&m[419])|(~m[413]&m[416]&~m[417]&m[418]&m[419])|(m[413]&m[416]&~m[417]&m[418]&m[419])|(~m[413]&~m[416]&m[417]&m[418]&m[419])|(m[413]&~m[416]&m[417]&m[418]&m[419])|(m[413]&m[416]&m[417]&m[418]&m[419]))):InitCond[129];
    m[420] = run?((((m[418]&~m[421]&~m[422]&~m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&m[423]&~m[424])|(m[418]&m[421]&~m[422]&m[423]&~m[424])|(m[418]&~m[421]&m[422]&m[423]&~m[424])|(~m[418]&m[421]&~m[422]&~m[423]&m[424])|(~m[418]&~m[421]&m[422]&~m[423]&m[424])|(m[418]&m[421]&m[422]&~m[423]&m[424])|(~m[418]&m[421]&m[422]&m[423]&m[424]))&UnbiasedRNG[31])|((m[418]&~m[421]&~m[422]&m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&m[422]&~m[423]&m[424])|(~m[418]&~m[421]&~m[422]&m[423]&m[424])|(m[418]&~m[421]&~m[422]&m[423]&m[424])|(~m[418]&m[421]&~m[422]&m[423]&m[424])|(m[418]&m[421]&~m[422]&m[423]&m[424])|(~m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&m[421]&m[422]&m[423]&m[424]))):InitCond[130];
    m[425] = run?((((m[423]&~m[426]&~m[427]&~m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&m[428]&~m[429])|(m[423]&m[426]&~m[427]&m[428]&~m[429])|(m[423]&~m[426]&m[427]&m[428]&~m[429])|(~m[423]&m[426]&~m[427]&~m[428]&m[429])|(~m[423]&~m[426]&m[427]&~m[428]&m[429])|(m[423]&m[426]&m[427]&~m[428]&m[429])|(~m[423]&m[426]&m[427]&m[428]&m[429]))&UnbiasedRNG[32])|((m[423]&~m[426]&~m[427]&m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&m[427]&~m[428]&m[429])|(~m[423]&~m[426]&~m[427]&m[428]&m[429])|(m[423]&~m[426]&~m[427]&m[428]&m[429])|(~m[423]&m[426]&~m[427]&m[428]&m[429])|(m[423]&m[426]&~m[427]&m[428]&m[429])|(~m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&m[426]&m[427]&m[428]&m[429]))):InitCond[131];
    m[430] = run?((((m[428]&~m[431]&~m[432]&~m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&m[433]&~m[434])|(m[428]&m[431]&~m[432]&m[433]&~m[434])|(m[428]&~m[431]&m[432]&m[433]&~m[434])|(~m[428]&m[431]&~m[432]&~m[433]&m[434])|(~m[428]&~m[431]&m[432]&~m[433]&m[434])|(m[428]&m[431]&m[432]&~m[433]&m[434])|(~m[428]&m[431]&m[432]&m[433]&m[434]))&UnbiasedRNG[33])|((m[428]&~m[431]&~m[432]&m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&m[432]&~m[433]&m[434])|(~m[428]&~m[431]&~m[432]&m[433]&m[434])|(m[428]&~m[431]&~m[432]&m[433]&m[434])|(~m[428]&m[431]&~m[432]&m[433]&m[434])|(m[428]&m[431]&~m[432]&m[433]&m[434])|(~m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&m[431]&m[432]&m[433]&m[434]))):InitCond[132];
    m[435] = run?((((m[266]&~m[436]&~m[437]&~m[438]&~m[439])|(~m[266]&~m[436]&~m[437]&m[438]&~m[439])|(m[266]&m[436]&~m[437]&m[438]&~m[439])|(m[266]&~m[436]&m[437]&m[438]&~m[439])|(~m[266]&m[436]&~m[437]&~m[438]&m[439])|(~m[266]&~m[436]&m[437]&~m[438]&m[439])|(m[266]&m[436]&m[437]&~m[438]&m[439])|(~m[266]&m[436]&m[437]&m[438]&m[439]))&UnbiasedRNG[34])|((m[266]&~m[436]&~m[437]&m[438]&~m[439])|(~m[266]&~m[436]&~m[437]&~m[438]&m[439])|(m[266]&~m[436]&~m[437]&~m[438]&m[439])|(m[266]&m[436]&~m[437]&~m[438]&m[439])|(m[266]&~m[436]&m[437]&~m[438]&m[439])|(~m[266]&~m[436]&~m[437]&m[438]&m[439])|(m[266]&~m[436]&~m[437]&m[438]&m[439])|(~m[266]&m[436]&~m[437]&m[438]&m[439])|(m[266]&m[436]&~m[437]&m[438]&m[439])|(~m[266]&~m[436]&m[437]&m[438]&m[439])|(m[266]&~m[436]&m[437]&m[438]&m[439])|(m[266]&m[436]&m[437]&m[438]&m[439]))):InitCond[133];
    m[440] = run?((((m[438]&~m[441]&~m[442]&~m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&m[443]&~m[444])|(m[438]&m[441]&~m[442]&m[443]&~m[444])|(m[438]&~m[441]&m[442]&m[443]&~m[444])|(~m[438]&m[441]&~m[442]&~m[443]&m[444])|(~m[438]&~m[441]&m[442]&~m[443]&m[444])|(m[438]&m[441]&m[442]&~m[443]&m[444])|(~m[438]&m[441]&m[442]&m[443]&m[444]))&UnbiasedRNG[35])|((m[438]&~m[441]&~m[442]&m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&m[442]&~m[443]&m[444])|(~m[438]&~m[441]&~m[442]&m[443]&m[444])|(m[438]&~m[441]&~m[442]&m[443]&m[444])|(~m[438]&m[441]&~m[442]&m[443]&m[444])|(m[438]&m[441]&~m[442]&m[443]&m[444])|(~m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&m[441]&m[442]&m[443]&m[444]))):InitCond[134];
    m[445] = run?((((m[443]&~m[446]&~m[447]&~m[448]&~m[449])|(~m[443]&~m[446]&~m[447]&m[448]&~m[449])|(m[443]&m[446]&~m[447]&m[448]&~m[449])|(m[443]&~m[446]&m[447]&m[448]&~m[449])|(~m[443]&m[446]&~m[447]&~m[448]&m[449])|(~m[443]&~m[446]&m[447]&~m[448]&m[449])|(m[443]&m[446]&m[447]&~m[448]&m[449])|(~m[443]&m[446]&m[447]&m[448]&m[449]))&UnbiasedRNG[36])|((m[443]&~m[446]&~m[447]&m[448]&~m[449])|(~m[443]&~m[446]&~m[447]&~m[448]&m[449])|(m[443]&~m[446]&~m[447]&~m[448]&m[449])|(m[443]&m[446]&~m[447]&~m[448]&m[449])|(m[443]&~m[446]&m[447]&~m[448]&m[449])|(~m[443]&~m[446]&~m[447]&m[448]&m[449])|(m[443]&~m[446]&~m[447]&m[448]&m[449])|(~m[443]&m[446]&~m[447]&m[448]&m[449])|(m[443]&m[446]&~m[447]&m[448]&m[449])|(~m[443]&~m[446]&m[447]&m[448]&m[449])|(m[443]&~m[446]&m[447]&m[448]&m[449])|(m[443]&m[446]&m[447]&m[448]&m[449]))):InitCond[135];
    m[450] = run?((((m[448]&~m[451]&~m[452]&~m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&m[453]&~m[454])|(m[448]&m[451]&~m[452]&m[453]&~m[454])|(m[448]&~m[451]&m[452]&m[453]&~m[454])|(~m[448]&m[451]&~m[452]&~m[453]&m[454])|(~m[448]&~m[451]&m[452]&~m[453]&m[454])|(m[448]&m[451]&m[452]&~m[453]&m[454])|(~m[448]&m[451]&m[452]&m[453]&m[454]))&UnbiasedRNG[37])|((m[448]&~m[451]&~m[452]&m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&m[452]&~m[453]&m[454])|(~m[448]&~m[451]&~m[452]&m[453]&m[454])|(m[448]&~m[451]&~m[452]&m[453]&m[454])|(~m[448]&m[451]&~m[452]&m[453]&m[454])|(m[448]&m[451]&~m[452]&m[453]&m[454])|(~m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&m[451]&m[452]&m[453]&m[454]))):InitCond[136];
    m[455] = run?((((m[453]&~m[456]&~m[457]&~m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&m[458]&~m[459])|(m[453]&m[456]&~m[457]&m[458]&~m[459])|(m[453]&~m[456]&m[457]&m[458]&~m[459])|(~m[453]&m[456]&~m[457]&~m[458]&m[459])|(~m[453]&~m[456]&m[457]&~m[458]&m[459])|(m[453]&m[456]&m[457]&~m[458]&m[459])|(~m[453]&m[456]&m[457]&m[458]&m[459]))&UnbiasedRNG[38])|((m[453]&~m[456]&~m[457]&m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&m[457]&~m[458]&m[459])|(~m[453]&~m[456]&~m[457]&m[458]&m[459])|(m[453]&~m[456]&~m[457]&m[458]&m[459])|(~m[453]&m[456]&~m[457]&m[458]&m[459])|(m[453]&m[456]&~m[457]&m[458]&m[459])|(~m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&m[456]&m[457]&m[458]&m[459]))):InitCond[137];
    m[460] = run?((((m[458]&~m[461]&~m[462]&~m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&m[463]&~m[464])|(m[458]&m[461]&~m[462]&m[463]&~m[464])|(m[458]&~m[461]&m[462]&m[463]&~m[464])|(~m[458]&m[461]&~m[462]&~m[463]&m[464])|(~m[458]&~m[461]&m[462]&~m[463]&m[464])|(m[458]&m[461]&m[462]&~m[463]&m[464])|(~m[458]&m[461]&m[462]&m[463]&m[464]))&UnbiasedRNG[39])|((m[458]&~m[461]&~m[462]&m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&m[462]&~m[463]&m[464])|(~m[458]&~m[461]&~m[462]&m[463]&m[464])|(m[458]&~m[461]&~m[462]&m[463]&m[464])|(~m[458]&m[461]&~m[462]&m[463]&m[464])|(m[458]&m[461]&~m[462]&m[463]&m[464])|(~m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&m[461]&m[462]&m[463]&m[464]))):InitCond[138];
    m[465] = run?((((m[267]&~m[466]&~m[467]&~m[468]&~m[469])|(~m[267]&~m[466]&~m[467]&m[468]&~m[469])|(m[267]&m[466]&~m[467]&m[468]&~m[469])|(m[267]&~m[466]&m[467]&m[468]&~m[469])|(~m[267]&m[466]&~m[467]&~m[468]&m[469])|(~m[267]&~m[466]&m[467]&~m[468]&m[469])|(m[267]&m[466]&m[467]&~m[468]&m[469])|(~m[267]&m[466]&m[467]&m[468]&m[469]))&UnbiasedRNG[40])|((m[267]&~m[466]&~m[467]&m[468]&~m[469])|(~m[267]&~m[466]&~m[467]&~m[468]&m[469])|(m[267]&~m[466]&~m[467]&~m[468]&m[469])|(m[267]&m[466]&~m[467]&~m[468]&m[469])|(m[267]&~m[466]&m[467]&~m[468]&m[469])|(~m[267]&~m[466]&~m[467]&m[468]&m[469])|(m[267]&~m[466]&~m[467]&m[468]&m[469])|(~m[267]&m[466]&~m[467]&m[468]&m[469])|(m[267]&m[466]&~m[467]&m[468]&m[469])|(~m[267]&~m[466]&m[467]&m[468]&m[469])|(m[267]&~m[466]&m[467]&m[468]&m[469])|(m[267]&m[466]&m[467]&m[468]&m[469]))):InitCond[139];
    m[470] = run?((((m[468]&~m[471]&~m[472]&~m[473]&~m[474])|(~m[468]&~m[471]&~m[472]&m[473]&~m[474])|(m[468]&m[471]&~m[472]&m[473]&~m[474])|(m[468]&~m[471]&m[472]&m[473]&~m[474])|(~m[468]&m[471]&~m[472]&~m[473]&m[474])|(~m[468]&~m[471]&m[472]&~m[473]&m[474])|(m[468]&m[471]&m[472]&~m[473]&m[474])|(~m[468]&m[471]&m[472]&m[473]&m[474]))&UnbiasedRNG[41])|((m[468]&~m[471]&~m[472]&m[473]&~m[474])|(~m[468]&~m[471]&~m[472]&~m[473]&m[474])|(m[468]&~m[471]&~m[472]&~m[473]&m[474])|(m[468]&m[471]&~m[472]&~m[473]&m[474])|(m[468]&~m[471]&m[472]&~m[473]&m[474])|(~m[468]&~m[471]&~m[472]&m[473]&m[474])|(m[468]&~m[471]&~m[472]&m[473]&m[474])|(~m[468]&m[471]&~m[472]&m[473]&m[474])|(m[468]&m[471]&~m[472]&m[473]&m[474])|(~m[468]&~m[471]&m[472]&m[473]&m[474])|(m[468]&~m[471]&m[472]&m[473]&m[474])|(m[468]&m[471]&m[472]&m[473]&m[474]))):InitCond[140];
    m[475] = run?((((m[473]&~m[476]&~m[477]&~m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&m[478]&~m[479])|(m[473]&m[476]&~m[477]&m[478]&~m[479])|(m[473]&~m[476]&m[477]&m[478]&~m[479])|(~m[473]&m[476]&~m[477]&~m[478]&m[479])|(~m[473]&~m[476]&m[477]&~m[478]&m[479])|(m[473]&m[476]&m[477]&~m[478]&m[479])|(~m[473]&m[476]&m[477]&m[478]&m[479]))&UnbiasedRNG[42])|((m[473]&~m[476]&~m[477]&m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&m[477]&~m[478]&m[479])|(~m[473]&~m[476]&~m[477]&m[478]&m[479])|(m[473]&~m[476]&~m[477]&m[478]&m[479])|(~m[473]&m[476]&~m[477]&m[478]&m[479])|(m[473]&m[476]&~m[477]&m[478]&m[479])|(~m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&m[476]&m[477]&m[478]&m[479]))):InitCond[141];
    m[480] = run?((((m[478]&~m[481]&~m[482]&~m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&m[483]&~m[484])|(m[478]&m[481]&~m[482]&m[483]&~m[484])|(m[478]&~m[481]&m[482]&m[483]&~m[484])|(~m[478]&m[481]&~m[482]&~m[483]&m[484])|(~m[478]&~m[481]&m[482]&~m[483]&m[484])|(m[478]&m[481]&m[482]&~m[483]&m[484])|(~m[478]&m[481]&m[482]&m[483]&m[484]))&UnbiasedRNG[43])|((m[478]&~m[481]&~m[482]&m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&m[482]&~m[483]&m[484])|(~m[478]&~m[481]&~m[482]&m[483]&m[484])|(m[478]&~m[481]&~m[482]&m[483]&m[484])|(~m[478]&m[481]&~m[482]&m[483]&m[484])|(m[478]&m[481]&~m[482]&m[483]&m[484])|(~m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&m[481]&m[482]&m[483]&m[484]))):InitCond[142];
    m[485] = run?((((m[483]&~m[486]&~m[487]&~m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&m[488]&~m[489])|(m[483]&m[486]&~m[487]&m[488]&~m[489])|(m[483]&~m[486]&m[487]&m[488]&~m[489])|(~m[483]&m[486]&~m[487]&~m[488]&m[489])|(~m[483]&~m[486]&m[487]&~m[488]&m[489])|(m[483]&m[486]&m[487]&~m[488]&m[489])|(~m[483]&m[486]&m[487]&m[488]&m[489]))&UnbiasedRNG[44])|((m[483]&~m[486]&~m[487]&m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&m[487]&~m[488]&m[489])|(~m[483]&~m[486]&~m[487]&m[488]&m[489])|(m[483]&~m[486]&~m[487]&m[488]&m[489])|(~m[483]&m[486]&~m[487]&m[488]&m[489])|(m[483]&m[486]&~m[487]&m[488]&m[489])|(~m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&m[486]&m[487]&m[488]&m[489]))):InitCond[143];
    m[490] = run?((((m[488]&~m[491]&~m[492]&~m[493]&~m[494])|(~m[488]&~m[491]&~m[492]&m[493]&~m[494])|(m[488]&m[491]&~m[492]&m[493]&~m[494])|(m[488]&~m[491]&m[492]&m[493]&~m[494])|(~m[488]&m[491]&~m[492]&~m[493]&m[494])|(~m[488]&~m[491]&m[492]&~m[493]&m[494])|(m[488]&m[491]&m[492]&~m[493]&m[494])|(~m[488]&m[491]&m[492]&m[493]&m[494]))&UnbiasedRNG[45])|((m[488]&~m[491]&~m[492]&m[493]&~m[494])|(~m[488]&~m[491]&~m[492]&~m[493]&m[494])|(m[488]&~m[491]&~m[492]&~m[493]&m[494])|(m[488]&m[491]&~m[492]&~m[493]&m[494])|(m[488]&~m[491]&m[492]&~m[493]&m[494])|(~m[488]&~m[491]&~m[492]&m[493]&m[494])|(m[488]&~m[491]&~m[492]&m[493]&m[494])|(~m[488]&m[491]&~m[492]&m[493]&m[494])|(m[488]&m[491]&~m[492]&m[493]&m[494])|(~m[488]&~m[491]&m[492]&m[493]&m[494])|(m[488]&~m[491]&m[492]&m[493]&m[494])|(m[488]&m[491]&m[492]&m[493]&m[494]))):InitCond[144];
    m[495] = run?((((m[493]&~m[496]&~m[497]&~m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&m[498]&~m[499])|(m[493]&m[496]&~m[497]&m[498]&~m[499])|(m[493]&~m[496]&m[497]&m[498]&~m[499])|(~m[493]&m[496]&~m[497]&~m[498]&m[499])|(~m[493]&~m[496]&m[497]&~m[498]&m[499])|(m[493]&m[496]&m[497]&~m[498]&m[499])|(~m[493]&m[496]&m[497]&m[498]&m[499]))&UnbiasedRNG[46])|((m[493]&~m[496]&~m[497]&m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&m[497]&~m[498]&m[499])|(~m[493]&~m[496]&~m[497]&m[498]&m[499])|(m[493]&~m[496]&~m[497]&m[498]&m[499])|(~m[493]&m[496]&~m[497]&m[498]&m[499])|(m[493]&m[496]&~m[497]&m[498]&m[499])|(~m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&m[496]&m[497]&m[498]&m[499]))):InitCond[145];
    m[500] = run?((((m[268]&~m[501]&~m[502]&~m[503]&~m[504])|(~m[268]&~m[501]&~m[502]&m[503]&~m[504])|(m[268]&m[501]&~m[502]&m[503]&~m[504])|(m[268]&~m[501]&m[502]&m[503]&~m[504])|(~m[268]&m[501]&~m[502]&~m[503]&m[504])|(~m[268]&~m[501]&m[502]&~m[503]&m[504])|(m[268]&m[501]&m[502]&~m[503]&m[504])|(~m[268]&m[501]&m[502]&m[503]&m[504]))&UnbiasedRNG[47])|((m[268]&~m[501]&~m[502]&m[503]&~m[504])|(~m[268]&~m[501]&~m[502]&~m[503]&m[504])|(m[268]&~m[501]&~m[502]&~m[503]&m[504])|(m[268]&m[501]&~m[502]&~m[503]&m[504])|(m[268]&~m[501]&m[502]&~m[503]&m[504])|(~m[268]&~m[501]&~m[502]&m[503]&m[504])|(m[268]&~m[501]&~m[502]&m[503]&m[504])|(~m[268]&m[501]&~m[502]&m[503]&m[504])|(m[268]&m[501]&~m[502]&m[503]&m[504])|(~m[268]&~m[501]&m[502]&m[503]&m[504])|(m[268]&~m[501]&m[502]&m[503]&m[504])|(m[268]&m[501]&m[502]&m[503]&m[504]))):InitCond[146];
    m[505] = run?((((m[503]&~m[506]&~m[507]&~m[508]&~m[509])|(~m[503]&~m[506]&~m[507]&m[508]&~m[509])|(m[503]&m[506]&~m[507]&m[508]&~m[509])|(m[503]&~m[506]&m[507]&m[508]&~m[509])|(~m[503]&m[506]&~m[507]&~m[508]&m[509])|(~m[503]&~m[506]&m[507]&~m[508]&m[509])|(m[503]&m[506]&m[507]&~m[508]&m[509])|(~m[503]&m[506]&m[507]&m[508]&m[509]))&UnbiasedRNG[48])|((m[503]&~m[506]&~m[507]&m[508]&~m[509])|(~m[503]&~m[506]&~m[507]&~m[508]&m[509])|(m[503]&~m[506]&~m[507]&~m[508]&m[509])|(m[503]&m[506]&~m[507]&~m[508]&m[509])|(m[503]&~m[506]&m[507]&~m[508]&m[509])|(~m[503]&~m[506]&~m[507]&m[508]&m[509])|(m[503]&~m[506]&~m[507]&m[508]&m[509])|(~m[503]&m[506]&~m[507]&m[508]&m[509])|(m[503]&m[506]&~m[507]&m[508]&m[509])|(~m[503]&~m[506]&m[507]&m[508]&m[509])|(m[503]&~m[506]&m[507]&m[508]&m[509])|(m[503]&m[506]&m[507]&m[508]&m[509]))):InitCond[147];
    m[510] = run?((((m[508]&~m[511]&~m[512]&~m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&m[513]&~m[514])|(m[508]&m[511]&~m[512]&m[513]&~m[514])|(m[508]&~m[511]&m[512]&m[513]&~m[514])|(~m[508]&m[511]&~m[512]&~m[513]&m[514])|(~m[508]&~m[511]&m[512]&~m[513]&m[514])|(m[508]&m[511]&m[512]&~m[513]&m[514])|(~m[508]&m[511]&m[512]&m[513]&m[514]))&UnbiasedRNG[49])|((m[508]&~m[511]&~m[512]&m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&m[512]&~m[513]&m[514])|(~m[508]&~m[511]&~m[512]&m[513]&m[514])|(m[508]&~m[511]&~m[512]&m[513]&m[514])|(~m[508]&m[511]&~m[512]&m[513]&m[514])|(m[508]&m[511]&~m[512]&m[513]&m[514])|(~m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&m[511]&m[512]&m[513]&m[514]))):InitCond[148];
    m[515] = run?((((m[513]&~m[516]&~m[517]&~m[518]&~m[519])|(~m[513]&~m[516]&~m[517]&m[518]&~m[519])|(m[513]&m[516]&~m[517]&m[518]&~m[519])|(m[513]&~m[516]&m[517]&m[518]&~m[519])|(~m[513]&m[516]&~m[517]&~m[518]&m[519])|(~m[513]&~m[516]&m[517]&~m[518]&m[519])|(m[513]&m[516]&m[517]&~m[518]&m[519])|(~m[513]&m[516]&m[517]&m[518]&m[519]))&UnbiasedRNG[50])|((m[513]&~m[516]&~m[517]&m[518]&~m[519])|(~m[513]&~m[516]&~m[517]&~m[518]&m[519])|(m[513]&~m[516]&~m[517]&~m[518]&m[519])|(m[513]&m[516]&~m[517]&~m[518]&m[519])|(m[513]&~m[516]&m[517]&~m[518]&m[519])|(~m[513]&~m[516]&~m[517]&m[518]&m[519])|(m[513]&~m[516]&~m[517]&m[518]&m[519])|(~m[513]&m[516]&~m[517]&m[518]&m[519])|(m[513]&m[516]&~m[517]&m[518]&m[519])|(~m[513]&~m[516]&m[517]&m[518]&m[519])|(m[513]&~m[516]&m[517]&m[518]&m[519])|(m[513]&m[516]&m[517]&m[518]&m[519]))):InitCond[149];
    m[520] = run?((((m[518]&~m[521]&~m[522]&~m[523]&~m[524])|(~m[518]&~m[521]&~m[522]&m[523]&~m[524])|(m[518]&m[521]&~m[522]&m[523]&~m[524])|(m[518]&~m[521]&m[522]&m[523]&~m[524])|(~m[518]&m[521]&~m[522]&~m[523]&m[524])|(~m[518]&~m[521]&m[522]&~m[523]&m[524])|(m[518]&m[521]&m[522]&~m[523]&m[524])|(~m[518]&m[521]&m[522]&m[523]&m[524]))&UnbiasedRNG[51])|((m[518]&~m[521]&~m[522]&m[523]&~m[524])|(~m[518]&~m[521]&~m[522]&~m[523]&m[524])|(m[518]&~m[521]&~m[522]&~m[523]&m[524])|(m[518]&m[521]&~m[522]&~m[523]&m[524])|(m[518]&~m[521]&m[522]&~m[523]&m[524])|(~m[518]&~m[521]&~m[522]&m[523]&m[524])|(m[518]&~m[521]&~m[522]&m[523]&m[524])|(~m[518]&m[521]&~m[522]&m[523]&m[524])|(m[518]&m[521]&~m[522]&m[523]&m[524])|(~m[518]&~m[521]&m[522]&m[523]&m[524])|(m[518]&~m[521]&m[522]&m[523]&m[524])|(m[518]&m[521]&m[522]&m[523]&m[524]))):InitCond[150];
    m[525] = run?((((m[523]&~m[526]&~m[527]&~m[528]&~m[529])|(~m[523]&~m[526]&~m[527]&m[528]&~m[529])|(m[523]&m[526]&~m[527]&m[528]&~m[529])|(m[523]&~m[526]&m[527]&m[528]&~m[529])|(~m[523]&m[526]&~m[527]&~m[528]&m[529])|(~m[523]&~m[526]&m[527]&~m[528]&m[529])|(m[523]&m[526]&m[527]&~m[528]&m[529])|(~m[523]&m[526]&m[527]&m[528]&m[529]))&UnbiasedRNG[52])|((m[523]&~m[526]&~m[527]&m[528]&~m[529])|(~m[523]&~m[526]&~m[527]&~m[528]&m[529])|(m[523]&~m[526]&~m[527]&~m[528]&m[529])|(m[523]&m[526]&~m[527]&~m[528]&m[529])|(m[523]&~m[526]&m[527]&~m[528]&m[529])|(~m[523]&~m[526]&~m[527]&m[528]&m[529])|(m[523]&~m[526]&~m[527]&m[528]&m[529])|(~m[523]&m[526]&~m[527]&m[528]&m[529])|(m[523]&m[526]&~m[527]&m[528]&m[529])|(~m[523]&~m[526]&m[527]&m[528]&m[529])|(m[523]&~m[526]&m[527]&m[528]&m[529])|(m[523]&m[526]&m[527]&m[528]&m[529]))):InitCond[151];
    m[530] = run?((((m[528]&~m[531]&~m[532]&~m[533]&~m[534])|(~m[528]&~m[531]&~m[532]&m[533]&~m[534])|(m[528]&m[531]&~m[532]&m[533]&~m[534])|(m[528]&~m[531]&m[532]&m[533]&~m[534])|(~m[528]&m[531]&~m[532]&~m[533]&m[534])|(~m[528]&~m[531]&m[532]&~m[533]&m[534])|(m[528]&m[531]&m[532]&~m[533]&m[534])|(~m[528]&m[531]&m[532]&m[533]&m[534]))&UnbiasedRNG[53])|((m[528]&~m[531]&~m[532]&m[533]&~m[534])|(~m[528]&~m[531]&~m[532]&~m[533]&m[534])|(m[528]&~m[531]&~m[532]&~m[533]&m[534])|(m[528]&m[531]&~m[532]&~m[533]&m[534])|(m[528]&~m[531]&m[532]&~m[533]&m[534])|(~m[528]&~m[531]&~m[532]&m[533]&m[534])|(m[528]&~m[531]&~m[532]&m[533]&m[534])|(~m[528]&m[531]&~m[532]&m[533]&m[534])|(m[528]&m[531]&~m[532]&m[533]&m[534])|(~m[528]&~m[531]&m[532]&m[533]&m[534])|(m[528]&~m[531]&m[532]&m[533]&m[534])|(m[528]&m[531]&m[532]&m[533]&m[534]))):InitCond[152];
    m[535] = run?((((m[533]&~m[536]&~m[537]&~m[538]&~m[539])|(~m[533]&~m[536]&~m[537]&m[538]&~m[539])|(m[533]&m[536]&~m[537]&m[538]&~m[539])|(m[533]&~m[536]&m[537]&m[538]&~m[539])|(~m[533]&m[536]&~m[537]&~m[538]&m[539])|(~m[533]&~m[536]&m[537]&~m[538]&m[539])|(m[533]&m[536]&m[537]&~m[538]&m[539])|(~m[533]&m[536]&m[537]&m[538]&m[539]))&UnbiasedRNG[54])|((m[533]&~m[536]&~m[537]&m[538]&~m[539])|(~m[533]&~m[536]&~m[537]&~m[538]&m[539])|(m[533]&~m[536]&~m[537]&~m[538]&m[539])|(m[533]&m[536]&~m[537]&~m[538]&m[539])|(m[533]&~m[536]&m[537]&~m[538]&m[539])|(~m[533]&~m[536]&~m[537]&m[538]&m[539])|(m[533]&~m[536]&~m[537]&m[538]&m[539])|(~m[533]&m[536]&~m[537]&m[538]&m[539])|(m[533]&m[536]&~m[537]&m[538]&m[539])|(~m[533]&~m[536]&m[537]&m[538]&m[539])|(m[533]&~m[536]&m[537]&m[538]&m[539])|(m[533]&m[536]&m[537]&m[538]&m[539]))):InitCond[153];
    m[540] = run?((((m[269]&~m[541]&~m[542]&~m[543]&~m[544])|(~m[269]&~m[541]&~m[542]&m[543]&~m[544])|(m[269]&m[541]&~m[542]&m[543]&~m[544])|(m[269]&~m[541]&m[542]&m[543]&~m[544])|(~m[269]&m[541]&~m[542]&~m[543]&m[544])|(~m[269]&~m[541]&m[542]&~m[543]&m[544])|(m[269]&m[541]&m[542]&~m[543]&m[544])|(~m[269]&m[541]&m[542]&m[543]&m[544]))&UnbiasedRNG[55])|((m[269]&~m[541]&~m[542]&m[543]&~m[544])|(~m[269]&~m[541]&~m[542]&~m[543]&m[544])|(m[269]&~m[541]&~m[542]&~m[543]&m[544])|(m[269]&m[541]&~m[542]&~m[543]&m[544])|(m[269]&~m[541]&m[542]&~m[543]&m[544])|(~m[269]&~m[541]&~m[542]&m[543]&m[544])|(m[269]&~m[541]&~m[542]&m[543]&m[544])|(~m[269]&m[541]&~m[542]&m[543]&m[544])|(m[269]&m[541]&~m[542]&m[543]&m[544])|(~m[269]&~m[541]&m[542]&m[543]&m[544])|(m[269]&~m[541]&m[542]&m[543]&m[544])|(m[269]&m[541]&m[542]&m[543]&m[544]))):InitCond[154];
    m[545] = run?((((m[543]&~m[546]&~m[547]&~m[548]&~m[549])|(~m[543]&~m[546]&~m[547]&m[548]&~m[549])|(m[543]&m[546]&~m[547]&m[548]&~m[549])|(m[543]&~m[546]&m[547]&m[548]&~m[549])|(~m[543]&m[546]&~m[547]&~m[548]&m[549])|(~m[543]&~m[546]&m[547]&~m[548]&m[549])|(m[543]&m[546]&m[547]&~m[548]&m[549])|(~m[543]&m[546]&m[547]&m[548]&m[549]))&UnbiasedRNG[56])|((m[543]&~m[546]&~m[547]&m[548]&~m[549])|(~m[543]&~m[546]&~m[547]&~m[548]&m[549])|(m[543]&~m[546]&~m[547]&~m[548]&m[549])|(m[543]&m[546]&~m[547]&~m[548]&m[549])|(m[543]&~m[546]&m[547]&~m[548]&m[549])|(~m[543]&~m[546]&~m[547]&m[548]&m[549])|(m[543]&~m[546]&~m[547]&m[548]&m[549])|(~m[543]&m[546]&~m[547]&m[548]&m[549])|(m[543]&m[546]&~m[547]&m[548]&m[549])|(~m[543]&~m[546]&m[547]&m[548]&m[549])|(m[543]&~m[546]&m[547]&m[548]&m[549])|(m[543]&m[546]&m[547]&m[548]&m[549]))):InitCond[155];
    m[550] = run?((((m[548]&~m[551]&~m[552]&~m[553]&~m[554])|(~m[548]&~m[551]&~m[552]&m[553]&~m[554])|(m[548]&m[551]&~m[552]&m[553]&~m[554])|(m[548]&~m[551]&m[552]&m[553]&~m[554])|(~m[548]&m[551]&~m[552]&~m[553]&m[554])|(~m[548]&~m[551]&m[552]&~m[553]&m[554])|(m[548]&m[551]&m[552]&~m[553]&m[554])|(~m[548]&m[551]&m[552]&m[553]&m[554]))&UnbiasedRNG[57])|((m[548]&~m[551]&~m[552]&m[553]&~m[554])|(~m[548]&~m[551]&~m[552]&~m[553]&m[554])|(m[548]&~m[551]&~m[552]&~m[553]&m[554])|(m[548]&m[551]&~m[552]&~m[553]&m[554])|(m[548]&~m[551]&m[552]&~m[553]&m[554])|(~m[548]&~m[551]&~m[552]&m[553]&m[554])|(m[548]&~m[551]&~m[552]&m[553]&m[554])|(~m[548]&m[551]&~m[552]&m[553]&m[554])|(m[548]&m[551]&~m[552]&m[553]&m[554])|(~m[548]&~m[551]&m[552]&m[553]&m[554])|(m[548]&~m[551]&m[552]&m[553]&m[554])|(m[548]&m[551]&m[552]&m[553]&m[554]))):InitCond[156];
    m[555] = run?((((m[553]&~m[556]&~m[557]&~m[558]&~m[559])|(~m[553]&~m[556]&~m[557]&m[558]&~m[559])|(m[553]&m[556]&~m[557]&m[558]&~m[559])|(m[553]&~m[556]&m[557]&m[558]&~m[559])|(~m[553]&m[556]&~m[557]&~m[558]&m[559])|(~m[553]&~m[556]&m[557]&~m[558]&m[559])|(m[553]&m[556]&m[557]&~m[558]&m[559])|(~m[553]&m[556]&m[557]&m[558]&m[559]))&UnbiasedRNG[58])|((m[553]&~m[556]&~m[557]&m[558]&~m[559])|(~m[553]&~m[556]&~m[557]&~m[558]&m[559])|(m[553]&~m[556]&~m[557]&~m[558]&m[559])|(m[553]&m[556]&~m[557]&~m[558]&m[559])|(m[553]&~m[556]&m[557]&~m[558]&m[559])|(~m[553]&~m[556]&~m[557]&m[558]&m[559])|(m[553]&~m[556]&~m[557]&m[558]&m[559])|(~m[553]&m[556]&~m[557]&m[558]&m[559])|(m[553]&m[556]&~m[557]&m[558]&m[559])|(~m[553]&~m[556]&m[557]&m[558]&m[559])|(m[553]&~m[556]&m[557]&m[558]&m[559])|(m[553]&m[556]&m[557]&m[558]&m[559]))):InitCond[157];
    m[560] = run?((((m[558]&~m[561]&~m[562]&~m[563]&~m[564])|(~m[558]&~m[561]&~m[562]&m[563]&~m[564])|(m[558]&m[561]&~m[562]&m[563]&~m[564])|(m[558]&~m[561]&m[562]&m[563]&~m[564])|(~m[558]&m[561]&~m[562]&~m[563]&m[564])|(~m[558]&~m[561]&m[562]&~m[563]&m[564])|(m[558]&m[561]&m[562]&~m[563]&m[564])|(~m[558]&m[561]&m[562]&m[563]&m[564]))&UnbiasedRNG[59])|((m[558]&~m[561]&~m[562]&m[563]&~m[564])|(~m[558]&~m[561]&~m[562]&~m[563]&m[564])|(m[558]&~m[561]&~m[562]&~m[563]&m[564])|(m[558]&m[561]&~m[562]&~m[563]&m[564])|(m[558]&~m[561]&m[562]&~m[563]&m[564])|(~m[558]&~m[561]&~m[562]&m[563]&m[564])|(m[558]&~m[561]&~m[562]&m[563]&m[564])|(~m[558]&m[561]&~m[562]&m[563]&m[564])|(m[558]&m[561]&~m[562]&m[563]&m[564])|(~m[558]&~m[561]&m[562]&m[563]&m[564])|(m[558]&~m[561]&m[562]&m[563]&m[564])|(m[558]&m[561]&m[562]&m[563]&m[564]))):InitCond[158];
    m[565] = run?((((m[563]&~m[566]&~m[567]&~m[568]&~m[569])|(~m[563]&~m[566]&~m[567]&m[568]&~m[569])|(m[563]&m[566]&~m[567]&m[568]&~m[569])|(m[563]&~m[566]&m[567]&m[568]&~m[569])|(~m[563]&m[566]&~m[567]&~m[568]&m[569])|(~m[563]&~m[566]&m[567]&~m[568]&m[569])|(m[563]&m[566]&m[567]&~m[568]&m[569])|(~m[563]&m[566]&m[567]&m[568]&m[569]))&UnbiasedRNG[60])|((m[563]&~m[566]&~m[567]&m[568]&~m[569])|(~m[563]&~m[566]&~m[567]&~m[568]&m[569])|(m[563]&~m[566]&~m[567]&~m[568]&m[569])|(m[563]&m[566]&~m[567]&~m[568]&m[569])|(m[563]&~m[566]&m[567]&~m[568]&m[569])|(~m[563]&~m[566]&~m[567]&m[568]&m[569])|(m[563]&~m[566]&~m[567]&m[568]&m[569])|(~m[563]&m[566]&~m[567]&m[568]&m[569])|(m[563]&m[566]&~m[567]&m[568]&m[569])|(~m[563]&~m[566]&m[567]&m[568]&m[569])|(m[563]&~m[566]&m[567]&m[568]&m[569])|(m[563]&m[566]&m[567]&m[568]&m[569]))):InitCond[159];
    m[570] = run?((((m[568]&~m[571]&~m[572]&~m[573]&~m[574])|(~m[568]&~m[571]&~m[572]&m[573]&~m[574])|(m[568]&m[571]&~m[572]&m[573]&~m[574])|(m[568]&~m[571]&m[572]&m[573]&~m[574])|(~m[568]&m[571]&~m[572]&~m[573]&m[574])|(~m[568]&~m[571]&m[572]&~m[573]&m[574])|(m[568]&m[571]&m[572]&~m[573]&m[574])|(~m[568]&m[571]&m[572]&m[573]&m[574]))&UnbiasedRNG[61])|((m[568]&~m[571]&~m[572]&m[573]&~m[574])|(~m[568]&~m[571]&~m[572]&~m[573]&m[574])|(m[568]&~m[571]&~m[572]&~m[573]&m[574])|(m[568]&m[571]&~m[572]&~m[573]&m[574])|(m[568]&~m[571]&m[572]&~m[573]&m[574])|(~m[568]&~m[571]&~m[572]&m[573]&m[574])|(m[568]&~m[571]&~m[572]&m[573]&m[574])|(~m[568]&m[571]&~m[572]&m[573]&m[574])|(m[568]&m[571]&~m[572]&m[573]&m[574])|(~m[568]&~m[571]&m[572]&m[573]&m[574])|(m[568]&~m[571]&m[572]&m[573]&m[574])|(m[568]&m[571]&m[572]&m[573]&m[574]))):InitCond[160];
    m[575] = run?((((m[573]&~m[576]&~m[577]&~m[578]&~m[579])|(~m[573]&~m[576]&~m[577]&m[578]&~m[579])|(m[573]&m[576]&~m[577]&m[578]&~m[579])|(m[573]&~m[576]&m[577]&m[578]&~m[579])|(~m[573]&m[576]&~m[577]&~m[578]&m[579])|(~m[573]&~m[576]&m[577]&~m[578]&m[579])|(m[573]&m[576]&m[577]&~m[578]&m[579])|(~m[573]&m[576]&m[577]&m[578]&m[579]))&UnbiasedRNG[62])|((m[573]&~m[576]&~m[577]&m[578]&~m[579])|(~m[573]&~m[576]&~m[577]&~m[578]&m[579])|(m[573]&~m[576]&~m[577]&~m[578]&m[579])|(m[573]&m[576]&~m[577]&~m[578]&m[579])|(m[573]&~m[576]&m[577]&~m[578]&m[579])|(~m[573]&~m[576]&~m[577]&m[578]&m[579])|(m[573]&~m[576]&~m[577]&m[578]&m[579])|(~m[573]&m[576]&~m[577]&m[578]&m[579])|(m[573]&m[576]&~m[577]&m[578]&m[579])|(~m[573]&~m[576]&m[577]&m[578]&m[579])|(m[573]&~m[576]&m[577]&m[578]&m[579])|(m[573]&m[576]&m[577]&m[578]&m[579]))):InitCond[161];
    m[580] = run?((((m[578]&~m[581]&~m[582]&~m[583]&~m[584])|(~m[578]&~m[581]&~m[582]&m[583]&~m[584])|(m[578]&m[581]&~m[582]&m[583]&~m[584])|(m[578]&~m[581]&m[582]&m[583]&~m[584])|(~m[578]&m[581]&~m[582]&~m[583]&m[584])|(~m[578]&~m[581]&m[582]&~m[583]&m[584])|(m[578]&m[581]&m[582]&~m[583]&m[584])|(~m[578]&m[581]&m[582]&m[583]&m[584]))&UnbiasedRNG[63])|((m[578]&~m[581]&~m[582]&m[583]&~m[584])|(~m[578]&~m[581]&~m[582]&~m[583]&m[584])|(m[578]&~m[581]&~m[582]&~m[583]&m[584])|(m[578]&m[581]&~m[582]&~m[583]&m[584])|(m[578]&~m[581]&m[582]&~m[583]&m[584])|(~m[578]&~m[581]&~m[582]&m[583]&m[584])|(m[578]&~m[581]&~m[582]&m[583]&m[584])|(~m[578]&m[581]&~m[582]&m[583]&m[584])|(m[578]&m[581]&~m[582]&m[583]&m[584])|(~m[578]&~m[581]&m[582]&m[583]&m[584])|(m[578]&~m[581]&m[582]&m[583]&m[584])|(m[578]&m[581]&m[582]&m[583]&m[584]))):InitCond[162];
    m[590] = run?((((m[588]&~m[591]&~m[592]&~m[593]&~m[594])|(~m[588]&~m[591]&~m[592]&m[593]&~m[594])|(m[588]&m[591]&~m[592]&m[593]&~m[594])|(m[588]&~m[591]&m[592]&m[593]&~m[594])|(~m[588]&m[591]&~m[592]&~m[593]&m[594])|(~m[588]&~m[591]&m[592]&~m[593]&m[594])|(m[588]&m[591]&m[592]&~m[593]&m[594])|(~m[588]&m[591]&m[592]&m[593]&m[594]))&UnbiasedRNG[64])|((m[588]&~m[591]&~m[592]&m[593]&~m[594])|(~m[588]&~m[591]&~m[592]&~m[593]&m[594])|(m[588]&~m[591]&~m[592]&~m[593]&m[594])|(m[588]&m[591]&~m[592]&~m[593]&m[594])|(m[588]&~m[591]&m[592]&~m[593]&m[594])|(~m[588]&~m[591]&~m[592]&m[593]&m[594])|(m[588]&~m[591]&~m[592]&m[593]&m[594])|(~m[588]&m[591]&~m[592]&m[593]&m[594])|(m[588]&m[591]&~m[592]&m[593]&m[594])|(~m[588]&~m[591]&m[592]&m[593]&m[594])|(m[588]&~m[591]&m[592]&m[593]&m[594])|(m[588]&m[591]&m[592]&m[593]&m[594]))):InitCond[163];
    m[595] = run?((((m[593]&~m[596]&~m[597]&~m[598]&~m[599])|(~m[593]&~m[596]&~m[597]&m[598]&~m[599])|(m[593]&m[596]&~m[597]&m[598]&~m[599])|(m[593]&~m[596]&m[597]&m[598]&~m[599])|(~m[593]&m[596]&~m[597]&~m[598]&m[599])|(~m[593]&~m[596]&m[597]&~m[598]&m[599])|(m[593]&m[596]&m[597]&~m[598]&m[599])|(~m[593]&m[596]&m[597]&m[598]&m[599]))&UnbiasedRNG[65])|((m[593]&~m[596]&~m[597]&m[598]&~m[599])|(~m[593]&~m[596]&~m[597]&~m[598]&m[599])|(m[593]&~m[596]&~m[597]&~m[598]&m[599])|(m[593]&m[596]&~m[597]&~m[598]&m[599])|(m[593]&~m[596]&m[597]&~m[598]&m[599])|(~m[593]&~m[596]&~m[597]&m[598]&m[599])|(m[593]&~m[596]&~m[597]&m[598]&m[599])|(~m[593]&m[596]&~m[597]&m[598]&m[599])|(m[593]&m[596]&~m[597]&m[598]&m[599])|(~m[593]&~m[596]&m[597]&m[598]&m[599])|(m[593]&~m[596]&m[597]&m[598]&m[599])|(m[593]&m[596]&m[597]&m[598]&m[599]))):InitCond[164];
    m[600] = run?((((m[598]&~m[601]&~m[602]&~m[603]&~m[604])|(~m[598]&~m[601]&~m[602]&m[603]&~m[604])|(m[598]&m[601]&~m[602]&m[603]&~m[604])|(m[598]&~m[601]&m[602]&m[603]&~m[604])|(~m[598]&m[601]&~m[602]&~m[603]&m[604])|(~m[598]&~m[601]&m[602]&~m[603]&m[604])|(m[598]&m[601]&m[602]&~m[603]&m[604])|(~m[598]&m[601]&m[602]&m[603]&m[604]))&UnbiasedRNG[66])|((m[598]&~m[601]&~m[602]&m[603]&~m[604])|(~m[598]&~m[601]&~m[602]&~m[603]&m[604])|(m[598]&~m[601]&~m[602]&~m[603]&m[604])|(m[598]&m[601]&~m[602]&~m[603]&m[604])|(m[598]&~m[601]&m[602]&~m[603]&m[604])|(~m[598]&~m[601]&~m[602]&m[603]&m[604])|(m[598]&~m[601]&~m[602]&m[603]&m[604])|(~m[598]&m[601]&~m[602]&m[603]&m[604])|(m[598]&m[601]&~m[602]&m[603]&m[604])|(~m[598]&~m[601]&m[602]&m[603]&m[604])|(m[598]&~m[601]&m[602]&m[603]&m[604])|(m[598]&m[601]&m[602]&m[603]&m[604]))):InitCond[165];
    m[605] = run?((((m[603]&~m[606]&~m[607]&~m[608]&~m[609])|(~m[603]&~m[606]&~m[607]&m[608]&~m[609])|(m[603]&m[606]&~m[607]&m[608]&~m[609])|(m[603]&~m[606]&m[607]&m[608]&~m[609])|(~m[603]&m[606]&~m[607]&~m[608]&m[609])|(~m[603]&~m[606]&m[607]&~m[608]&m[609])|(m[603]&m[606]&m[607]&~m[608]&m[609])|(~m[603]&m[606]&m[607]&m[608]&m[609]))&UnbiasedRNG[67])|((m[603]&~m[606]&~m[607]&m[608]&~m[609])|(~m[603]&~m[606]&~m[607]&~m[608]&m[609])|(m[603]&~m[606]&~m[607]&~m[608]&m[609])|(m[603]&m[606]&~m[607]&~m[608]&m[609])|(m[603]&~m[606]&m[607]&~m[608]&m[609])|(~m[603]&~m[606]&~m[607]&m[608]&m[609])|(m[603]&~m[606]&~m[607]&m[608]&m[609])|(~m[603]&m[606]&~m[607]&m[608]&m[609])|(m[603]&m[606]&~m[607]&m[608]&m[609])|(~m[603]&~m[606]&m[607]&m[608]&m[609])|(m[603]&~m[606]&m[607]&m[608]&m[609])|(m[603]&m[606]&m[607]&m[608]&m[609]))):InitCond[166];
    m[610] = run?((((m[608]&~m[611]&~m[612]&~m[613]&~m[614])|(~m[608]&~m[611]&~m[612]&m[613]&~m[614])|(m[608]&m[611]&~m[612]&m[613]&~m[614])|(m[608]&~m[611]&m[612]&m[613]&~m[614])|(~m[608]&m[611]&~m[612]&~m[613]&m[614])|(~m[608]&~m[611]&m[612]&~m[613]&m[614])|(m[608]&m[611]&m[612]&~m[613]&m[614])|(~m[608]&m[611]&m[612]&m[613]&m[614]))&UnbiasedRNG[68])|((m[608]&~m[611]&~m[612]&m[613]&~m[614])|(~m[608]&~m[611]&~m[612]&~m[613]&m[614])|(m[608]&~m[611]&~m[612]&~m[613]&m[614])|(m[608]&m[611]&~m[612]&~m[613]&m[614])|(m[608]&~m[611]&m[612]&~m[613]&m[614])|(~m[608]&~m[611]&~m[612]&m[613]&m[614])|(m[608]&~m[611]&~m[612]&m[613]&m[614])|(~m[608]&m[611]&~m[612]&m[613]&m[614])|(m[608]&m[611]&~m[612]&m[613]&m[614])|(~m[608]&~m[611]&m[612]&m[613]&m[614])|(m[608]&~m[611]&m[612]&m[613]&m[614])|(m[608]&m[611]&m[612]&m[613]&m[614]))):InitCond[167];
    m[615] = run?((((m[613]&~m[616]&~m[617]&~m[618]&~m[619])|(~m[613]&~m[616]&~m[617]&m[618]&~m[619])|(m[613]&m[616]&~m[617]&m[618]&~m[619])|(m[613]&~m[616]&m[617]&m[618]&~m[619])|(~m[613]&m[616]&~m[617]&~m[618]&m[619])|(~m[613]&~m[616]&m[617]&~m[618]&m[619])|(m[613]&m[616]&m[617]&~m[618]&m[619])|(~m[613]&m[616]&m[617]&m[618]&m[619]))&UnbiasedRNG[69])|((m[613]&~m[616]&~m[617]&m[618]&~m[619])|(~m[613]&~m[616]&~m[617]&~m[618]&m[619])|(m[613]&~m[616]&~m[617]&~m[618]&m[619])|(m[613]&m[616]&~m[617]&~m[618]&m[619])|(m[613]&~m[616]&m[617]&~m[618]&m[619])|(~m[613]&~m[616]&~m[617]&m[618]&m[619])|(m[613]&~m[616]&~m[617]&m[618]&m[619])|(~m[613]&m[616]&~m[617]&m[618]&m[619])|(m[613]&m[616]&~m[617]&m[618]&m[619])|(~m[613]&~m[616]&m[617]&m[618]&m[619])|(m[613]&~m[616]&m[617]&m[618]&m[619])|(m[613]&m[616]&m[617]&m[618]&m[619]))):InitCond[168];
    m[620] = run?((((m[618]&~m[621]&~m[622]&~m[623]&~m[624])|(~m[618]&~m[621]&~m[622]&m[623]&~m[624])|(m[618]&m[621]&~m[622]&m[623]&~m[624])|(m[618]&~m[621]&m[622]&m[623]&~m[624])|(~m[618]&m[621]&~m[622]&~m[623]&m[624])|(~m[618]&~m[621]&m[622]&~m[623]&m[624])|(m[618]&m[621]&m[622]&~m[623]&m[624])|(~m[618]&m[621]&m[622]&m[623]&m[624]))&UnbiasedRNG[70])|((m[618]&~m[621]&~m[622]&m[623]&~m[624])|(~m[618]&~m[621]&~m[622]&~m[623]&m[624])|(m[618]&~m[621]&~m[622]&~m[623]&m[624])|(m[618]&m[621]&~m[622]&~m[623]&m[624])|(m[618]&~m[621]&m[622]&~m[623]&m[624])|(~m[618]&~m[621]&~m[622]&m[623]&m[624])|(m[618]&~m[621]&~m[622]&m[623]&m[624])|(~m[618]&m[621]&~m[622]&m[623]&m[624])|(m[618]&m[621]&~m[622]&m[623]&m[624])|(~m[618]&~m[621]&m[622]&m[623]&m[624])|(m[618]&~m[621]&m[622]&m[623]&m[624])|(m[618]&m[621]&m[622]&m[623]&m[624]))):InitCond[169];
    m[625] = run?((((m[623]&~m[626]&~m[627]&~m[628]&~m[629])|(~m[623]&~m[626]&~m[627]&m[628]&~m[629])|(m[623]&m[626]&~m[627]&m[628]&~m[629])|(m[623]&~m[626]&m[627]&m[628]&~m[629])|(~m[623]&m[626]&~m[627]&~m[628]&m[629])|(~m[623]&~m[626]&m[627]&~m[628]&m[629])|(m[623]&m[626]&m[627]&~m[628]&m[629])|(~m[623]&m[626]&m[627]&m[628]&m[629]))&UnbiasedRNG[71])|((m[623]&~m[626]&~m[627]&m[628]&~m[629])|(~m[623]&~m[626]&~m[627]&~m[628]&m[629])|(m[623]&~m[626]&~m[627]&~m[628]&m[629])|(m[623]&m[626]&~m[627]&~m[628]&m[629])|(m[623]&~m[626]&m[627]&~m[628]&m[629])|(~m[623]&~m[626]&~m[627]&m[628]&m[629])|(m[623]&~m[626]&~m[627]&m[628]&m[629])|(~m[623]&m[626]&~m[627]&m[628]&m[629])|(m[623]&m[626]&~m[627]&m[628]&m[629])|(~m[623]&~m[626]&m[627]&m[628]&m[629])|(m[623]&~m[626]&m[627]&m[628]&m[629])|(m[623]&m[626]&m[627]&m[628]&m[629]))):InitCond[170];
    m[630] = run?((((m[589]&~m[631]&~m[632]&~m[633]&~m[634])|(~m[589]&~m[631]&~m[632]&m[633]&~m[634])|(m[589]&m[631]&~m[632]&m[633]&~m[634])|(m[589]&~m[631]&m[632]&m[633]&~m[634])|(~m[589]&m[631]&~m[632]&~m[633]&m[634])|(~m[589]&~m[631]&m[632]&~m[633]&m[634])|(m[589]&m[631]&m[632]&~m[633]&m[634])|(~m[589]&m[631]&m[632]&m[633]&m[634]))&UnbiasedRNG[72])|((m[589]&~m[631]&~m[632]&m[633]&~m[634])|(~m[589]&~m[631]&~m[632]&~m[633]&m[634])|(m[589]&~m[631]&~m[632]&~m[633]&m[634])|(m[589]&m[631]&~m[632]&~m[633]&m[634])|(m[589]&~m[631]&m[632]&~m[633]&m[634])|(~m[589]&~m[631]&~m[632]&m[633]&m[634])|(m[589]&~m[631]&~m[632]&m[633]&m[634])|(~m[589]&m[631]&~m[632]&m[633]&m[634])|(m[589]&m[631]&~m[632]&m[633]&m[634])|(~m[589]&~m[631]&m[632]&m[633]&m[634])|(m[589]&~m[631]&m[632]&m[633]&m[634])|(m[589]&m[631]&m[632]&m[633]&m[634]))):InitCond[171];
    m[635] = run?((((m[633]&~m[636]&~m[637]&~m[638]&~m[639])|(~m[633]&~m[636]&~m[637]&m[638]&~m[639])|(m[633]&m[636]&~m[637]&m[638]&~m[639])|(m[633]&~m[636]&m[637]&m[638]&~m[639])|(~m[633]&m[636]&~m[637]&~m[638]&m[639])|(~m[633]&~m[636]&m[637]&~m[638]&m[639])|(m[633]&m[636]&m[637]&~m[638]&m[639])|(~m[633]&m[636]&m[637]&m[638]&m[639]))&UnbiasedRNG[73])|((m[633]&~m[636]&~m[637]&m[638]&~m[639])|(~m[633]&~m[636]&~m[637]&~m[638]&m[639])|(m[633]&~m[636]&~m[637]&~m[638]&m[639])|(m[633]&m[636]&~m[637]&~m[638]&m[639])|(m[633]&~m[636]&m[637]&~m[638]&m[639])|(~m[633]&~m[636]&~m[637]&m[638]&m[639])|(m[633]&~m[636]&~m[637]&m[638]&m[639])|(~m[633]&m[636]&~m[637]&m[638]&m[639])|(m[633]&m[636]&~m[637]&m[638]&m[639])|(~m[633]&~m[636]&m[637]&m[638]&m[639])|(m[633]&~m[636]&m[637]&m[638]&m[639])|(m[633]&m[636]&m[637]&m[638]&m[639]))):InitCond[172];
    m[640] = run?((((m[638]&~m[641]&~m[642]&~m[643]&~m[644])|(~m[638]&~m[641]&~m[642]&m[643]&~m[644])|(m[638]&m[641]&~m[642]&m[643]&~m[644])|(m[638]&~m[641]&m[642]&m[643]&~m[644])|(~m[638]&m[641]&~m[642]&~m[643]&m[644])|(~m[638]&~m[641]&m[642]&~m[643]&m[644])|(m[638]&m[641]&m[642]&~m[643]&m[644])|(~m[638]&m[641]&m[642]&m[643]&m[644]))&UnbiasedRNG[74])|((m[638]&~m[641]&~m[642]&m[643]&~m[644])|(~m[638]&~m[641]&~m[642]&~m[643]&m[644])|(m[638]&~m[641]&~m[642]&~m[643]&m[644])|(m[638]&m[641]&~m[642]&~m[643]&m[644])|(m[638]&~m[641]&m[642]&~m[643]&m[644])|(~m[638]&~m[641]&~m[642]&m[643]&m[644])|(m[638]&~m[641]&~m[642]&m[643]&m[644])|(~m[638]&m[641]&~m[642]&m[643]&m[644])|(m[638]&m[641]&~m[642]&m[643]&m[644])|(~m[638]&~m[641]&m[642]&m[643]&m[644])|(m[638]&~m[641]&m[642]&m[643]&m[644])|(m[638]&m[641]&m[642]&m[643]&m[644]))):InitCond[173];
    m[645] = run?((((m[643]&~m[646]&~m[647]&~m[648]&~m[649])|(~m[643]&~m[646]&~m[647]&m[648]&~m[649])|(m[643]&m[646]&~m[647]&m[648]&~m[649])|(m[643]&~m[646]&m[647]&m[648]&~m[649])|(~m[643]&m[646]&~m[647]&~m[648]&m[649])|(~m[643]&~m[646]&m[647]&~m[648]&m[649])|(m[643]&m[646]&m[647]&~m[648]&m[649])|(~m[643]&m[646]&m[647]&m[648]&m[649]))&UnbiasedRNG[75])|((m[643]&~m[646]&~m[647]&m[648]&~m[649])|(~m[643]&~m[646]&~m[647]&~m[648]&m[649])|(m[643]&~m[646]&~m[647]&~m[648]&m[649])|(m[643]&m[646]&~m[647]&~m[648]&m[649])|(m[643]&~m[646]&m[647]&~m[648]&m[649])|(~m[643]&~m[646]&~m[647]&m[648]&m[649])|(m[643]&~m[646]&~m[647]&m[648]&m[649])|(~m[643]&m[646]&~m[647]&m[648]&m[649])|(m[643]&m[646]&~m[647]&m[648]&m[649])|(~m[643]&~m[646]&m[647]&m[648]&m[649])|(m[643]&~m[646]&m[647]&m[648]&m[649])|(m[643]&m[646]&m[647]&m[648]&m[649]))):InitCond[174];
    m[650] = run?((((m[648]&~m[651]&~m[652]&~m[653]&~m[654])|(~m[648]&~m[651]&~m[652]&m[653]&~m[654])|(m[648]&m[651]&~m[652]&m[653]&~m[654])|(m[648]&~m[651]&m[652]&m[653]&~m[654])|(~m[648]&m[651]&~m[652]&~m[653]&m[654])|(~m[648]&~m[651]&m[652]&~m[653]&m[654])|(m[648]&m[651]&m[652]&~m[653]&m[654])|(~m[648]&m[651]&m[652]&m[653]&m[654]))&UnbiasedRNG[76])|((m[648]&~m[651]&~m[652]&m[653]&~m[654])|(~m[648]&~m[651]&~m[652]&~m[653]&m[654])|(m[648]&~m[651]&~m[652]&~m[653]&m[654])|(m[648]&m[651]&~m[652]&~m[653]&m[654])|(m[648]&~m[651]&m[652]&~m[653]&m[654])|(~m[648]&~m[651]&~m[652]&m[653]&m[654])|(m[648]&~m[651]&~m[652]&m[653]&m[654])|(~m[648]&m[651]&~m[652]&m[653]&m[654])|(m[648]&m[651]&~m[652]&m[653]&m[654])|(~m[648]&~m[651]&m[652]&m[653]&m[654])|(m[648]&~m[651]&m[652]&m[653]&m[654])|(m[648]&m[651]&m[652]&m[653]&m[654]))):InitCond[175];
    m[655] = run?((((m[653]&~m[656]&~m[657]&~m[658]&~m[659])|(~m[653]&~m[656]&~m[657]&m[658]&~m[659])|(m[653]&m[656]&~m[657]&m[658]&~m[659])|(m[653]&~m[656]&m[657]&m[658]&~m[659])|(~m[653]&m[656]&~m[657]&~m[658]&m[659])|(~m[653]&~m[656]&m[657]&~m[658]&m[659])|(m[653]&m[656]&m[657]&~m[658]&m[659])|(~m[653]&m[656]&m[657]&m[658]&m[659]))&UnbiasedRNG[77])|((m[653]&~m[656]&~m[657]&m[658]&~m[659])|(~m[653]&~m[656]&~m[657]&~m[658]&m[659])|(m[653]&~m[656]&~m[657]&~m[658]&m[659])|(m[653]&m[656]&~m[657]&~m[658]&m[659])|(m[653]&~m[656]&m[657]&~m[658]&m[659])|(~m[653]&~m[656]&~m[657]&m[658]&m[659])|(m[653]&~m[656]&~m[657]&m[658]&m[659])|(~m[653]&m[656]&~m[657]&m[658]&m[659])|(m[653]&m[656]&~m[657]&m[658]&m[659])|(~m[653]&~m[656]&m[657]&m[658]&m[659])|(m[653]&~m[656]&m[657]&m[658]&m[659])|(m[653]&m[656]&m[657]&m[658]&m[659]))):InitCond[176];
    m[660] = run?((((m[658]&~m[661]&~m[662]&~m[663]&~m[664])|(~m[658]&~m[661]&~m[662]&m[663]&~m[664])|(m[658]&m[661]&~m[662]&m[663]&~m[664])|(m[658]&~m[661]&m[662]&m[663]&~m[664])|(~m[658]&m[661]&~m[662]&~m[663]&m[664])|(~m[658]&~m[661]&m[662]&~m[663]&m[664])|(m[658]&m[661]&m[662]&~m[663]&m[664])|(~m[658]&m[661]&m[662]&m[663]&m[664]))&UnbiasedRNG[78])|((m[658]&~m[661]&~m[662]&m[663]&~m[664])|(~m[658]&~m[661]&~m[662]&~m[663]&m[664])|(m[658]&~m[661]&~m[662]&~m[663]&m[664])|(m[658]&m[661]&~m[662]&~m[663]&m[664])|(m[658]&~m[661]&m[662]&~m[663]&m[664])|(~m[658]&~m[661]&~m[662]&m[663]&m[664])|(m[658]&~m[661]&~m[662]&m[663]&m[664])|(~m[658]&m[661]&~m[662]&m[663]&m[664])|(m[658]&m[661]&~m[662]&m[663]&m[664])|(~m[658]&~m[661]&m[662]&m[663]&m[664])|(m[658]&~m[661]&m[662]&m[663]&m[664])|(m[658]&m[661]&m[662]&m[663]&m[664]))):InitCond[177];
    m[665] = run?((((m[663]&~m[666]&~m[667]&~m[668]&~m[669])|(~m[663]&~m[666]&~m[667]&m[668]&~m[669])|(m[663]&m[666]&~m[667]&m[668]&~m[669])|(m[663]&~m[666]&m[667]&m[668]&~m[669])|(~m[663]&m[666]&~m[667]&~m[668]&m[669])|(~m[663]&~m[666]&m[667]&~m[668]&m[669])|(m[663]&m[666]&m[667]&~m[668]&m[669])|(~m[663]&m[666]&m[667]&m[668]&m[669]))&UnbiasedRNG[79])|((m[663]&~m[666]&~m[667]&m[668]&~m[669])|(~m[663]&~m[666]&~m[667]&~m[668]&m[669])|(m[663]&~m[666]&~m[667]&~m[668]&m[669])|(m[663]&m[666]&~m[667]&~m[668]&m[669])|(m[663]&~m[666]&m[667]&~m[668]&m[669])|(~m[663]&~m[666]&~m[667]&m[668]&m[669])|(m[663]&~m[666]&~m[667]&m[668]&m[669])|(~m[663]&m[666]&~m[667]&m[668]&m[669])|(m[663]&m[666]&~m[667]&m[668]&m[669])|(~m[663]&~m[666]&m[667]&m[668]&m[669])|(m[663]&~m[666]&m[667]&m[668]&m[669])|(m[663]&m[666]&m[667]&m[668]&m[669]))):InitCond[178];
    m[670] = run?((((m[634]&~m[671]&~m[672]&~m[673]&~m[674])|(~m[634]&~m[671]&~m[672]&m[673]&~m[674])|(m[634]&m[671]&~m[672]&m[673]&~m[674])|(m[634]&~m[671]&m[672]&m[673]&~m[674])|(~m[634]&m[671]&~m[672]&~m[673]&m[674])|(~m[634]&~m[671]&m[672]&~m[673]&m[674])|(m[634]&m[671]&m[672]&~m[673]&m[674])|(~m[634]&m[671]&m[672]&m[673]&m[674]))&UnbiasedRNG[80])|((m[634]&~m[671]&~m[672]&m[673]&~m[674])|(~m[634]&~m[671]&~m[672]&~m[673]&m[674])|(m[634]&~m[671]&~m[672]&~m[673]&m[674])|(m[634]&m[671]&~m[672]&~m[673]&m[674])|(m[634]&~m[671]&m[672]&~m[673]&m[674])|(~m[634]&~m[671]&~m[672]&m[673]&m[674])|(m[634]&~m[671]&~m[672]&m[673]&m[674])|(~m[634]&m[671]&~m[672]&m[673]&m[674])|(m[634]&m[671]&~m[672]&m[673]&m[674])|(~m[634]&~m[671]&m[672]&m[673]&m[674])|(m[634]&~m[671]&m[672]&m[673]&m[674])|(m[634]&m[671]&m[672]&m[673]&m[674]))):InitCond[179];
    m[675] = run?((((m[673]&~m[676]&~m[677]&~m[678]&~m[679])|(~m[673]&~m[676]&~m[677]&m[678]&~m[679])|(m[673]&m[676]&~m[677]&m[678]&~m[679])|(m[673]&~m[676]&m[677]&m[678]&~m[679])|(~m[673]&m[676]&~m[677]&~m[678]&m[679])|(~m[673]&~m[676]&m[677]&~m[678]&m[679])|(m[673]&m[676]&m[677]&~m[678]&m[679])|(~m[673]&m[676]&m[677]&m[678]&m[679]))&UnbiasedRNG[81])|((m[673]&~m[676]&~m[677]&m[678]&~m[679])|(~m[673]&~m[676]&~m[677]&~m[678]&m[679])|(m[673]&~m[676]&~m[677]&~m[678]&m[679])|(m[673]&m[676]&~m[677]&~m[678]&m[679])|(m[673]&~m[676]&m[677]&~m[678]&m[679])|(~m[673]&~m[676]&~m[677]&m[678]&m[679])|(m[673]&~m[676]&~m[677]&m[678]&m[679])|(~m[673]&m[676]&~m[677]&m[678]&m[679])|(m[673]&m[676]&~m[677]&m[678]&m[679])|(~m[673]&~m[676]&m[677]&m[678]&m[679])|(m[673]&~m[676]&m[677]&m[678]&m[679])|(m[673]&m[676]&m[677]&m[678]&m[679]))):InitCond[180];
    m[680] = run?((((m[678]&~m[681]&~m[682]&~m[683]&~m[684])|(~m[678]&~m[681]&~m[682]&m[683]&~m[684])|(m[678]&m[681]&~m[682]&m[683]&~m[684])|(m[678]&~m[681]&m[682]&m[683]&~m[684])|(~m[678]&m[681]&~m[682]&~m[683]&m[684])|(~m[678]&~m[681]&m[682]&~m[683]&m[684])|(m[678]&m[681]&m[682]&~m[683]&m[684])|(~m[678]&m[681]&m[682]&m[683]&m[684]))&UnbiasedRNG[82])|((m[678]&~m[681]&~m[682]&m[683]&~m[684])|(~m[678]&~m[681]&~m[682]&~m[683]&m[684])|(m[678]&~m[681]&~m[682]&~m[683]&m[684])|(m[678]&m[681]&~m[682]&~m[683]&m[684])|(m[678]&~m[681]&m[682]&~m[683]&m[684])|(~m[678]&~m[681]&~m[682]&m[683]&m[684])|(m[678]&~m[681]&~m[682]&m[683]&m[684])|(~m[678]&m[681]&~m[682]&m[683]&m[684])|(m[678]&m[681]&~m[682]&m[683]&m[684])|(~m[678]&~m[681]&m[682]&m[683]&m[684])|(m[678]&~m[681]&m[682]&m[683]&m[684])|(m[678]&m[681]&m[682]&m[683]&m[684]))):InitCond[181];
    m[685] = run?((((m[683]&~m[686]&~m[687]&~m[688]&~m[689])|(~m[683]&~m[686]&~m[687]&m[688]&~m[689])|(m[683]&m[686]&~m[687]&m[688]&~m[689])|(m[683]&~m[686]&m[687]&m[688]&~m[689])|(~m[683]&m[686]&~m[687]&~m[688]&m[689])|(~m[683]&~m[686]&m[687]&~m[688]&m[689])|(m[683]&m[686]&m[687]&~m[688]&m[689])|(~m[683]&m[686]&m[687]&m[688]&m[689]))&UnbiasedRNG[83])|((m[683]&~m[686]&~m[687]&m[688]&~m[689])|(~m[683]&~m[686]&~m[687]&~m[688]&m[689])|(m[683]&~m[686]&~m[687]&~m[688]&m[689])|(m[683]&m[686]&~m[687]&~m[688]&m[689])|(m[683]&~m[686]&m[687]&~m[688]&m[689])|(~m[683]&~m[686]&~m[687]&m[688]&m[689])|(m[683]&~m[686]&~m[687]&m[688]&m[689])|(~m[683]&m[686]&~m[687]&m[688]&m[689])|(m[683]&m[686]&~m[687]&m[688]&m[689])|(~m[683]&~m[686]&m[687]&m[688]&m[689])|(m[683]&~m[686]&m[687]&m[688]&m[689])|(m[683]&m[686]&m[687]&m[688]&m[689]))):InitCond[182];
    m[690] = run?((((m[688]&~m[691]&~m[692]&~m[693]&~m[694])|(~m[688]&~m[691]&~m[692]&m[693]&~m[694])|(m[688]&m[691]&~m[692]&m[693]&~m[694])|(m[688]&~m[691]&m[692]&m[693]&~m[694])|(~m[688]&m[691]&~m[692]&~m[693]&m[694])|(~m[688]&~m[691]&m[692]&~m[693]&m[694])|(m[688]&m[691]&m[692]&~m[693]&m[694])|(~m[688]&m[691]&m[692]&m[693]&m[694]))&UnbiasedRNG[84])|((m[688]&~m[691]&~m[692]&m[693]&~m[694])|(~m[688]&~m[691]&~m[692]&~m[693]&m[694])|(m[688]&~m[691]&~m[692]&~m[693]&m[694])|(m[688]&m[691]&~m[692]&~m[693]&m[694])|(m[688]&~m[691]&m[692]&~m[693]&m[694])|(~m[688]&~m[691]&~m[692]&m[693]&m[694])|(m[688]&~m[691]&~m[692]&m[693]&m[694])|(~m[688]&m[691]&~m[692]&m[693]&m[694])|(m[688]&m[691]&~m[692]&m[693]&m[694])|(~m[688]&~m[691]&m[692]&m[693]&m[694])|(m[688]&~m[691]&m[692]&m[693]&m[694])|(m[688]&m[691]&m[692]&m[693]&m[694]))):InitCond[183];
    m[695] = run?((((m[693]&~m[696]&~m[697]&~m[698]&~m[699])|(~m[693]&~m[696]&~m[697]&m[698]&~m[699])|(m[693]&m[696]&~m[697]&m[698]&~m[699])|(m[693]&~m[696]&m[697]&m[698]&~m[699])|(~m[693]&m[696]&~m[697]&~m[698]&m[699])|(~m[693]&~m[696]&m[697]&~m[698]&m[699])|(m[693]&m[696]&m[697]&~m[698]&m[699])|(~m[693]&m[696]&m[697]&m[698]&m[699]))&UnbiasedRNG[85])|((m[693]&~m[696]&~m[697]&m[698]&~m[699])|(~m[693]&~m[696]&~m[697]&~m[698]&m[699])|(m[693]&~m[696]&~m[697]&~m[698]&m[699])|(m[693]&m[696]&~m[697]&~m[698]&m[699])|(m[693]&~m[696]&m[697]&~m[698]&m[699])|(~m[693]&~m[696]&~m[697]&m[698]&m[699])|(m[693]&~m[696]&~m[697]&m[698]&m[699])|(~m[693]&m[696]&~m[697]&m[698]&m[699])|(m[693]&m[696]&~m[697]&m[698]&m[699])|(~m[693]&~m[696]&m[697]&m[698]&m[699])|(m[693]&~m[696]&m[697]&m[698]&m[699])|(m[693]&m[696]&m[697]&m[698]&m[699]))):InitCond[184];
    m[700] = run?((((m[698]&~m[701]&~m[702]&~m[703]&~m[704])|(~m[698]&~m[701]&~m[702]&m[703]&~m[704])|(m[698]&m[701]&~m[702]&m[703]&~m[704])|(m[698]&~m[701]&m[702]&m[703]&~m[704])|(~m[698]&m[701]&~m[702]&~m[703]&m[704])|(~m[698]&~m[701]&m[702]&~m[703]&m[704])|(m[698]&m[701]&m[702]&~m[703]&m[704])|(~m[698]&m[701]&m[702]&m[703]&m[704]))&UnbiasedRNG[86])|((m[698]&~m[701]&~m[702]&m[703]&~m[704])|(~m[698]&~m[701]&~m[702]&~m[703]&m[704])|(m[698]&~m[701]&~m[702]&~m[703]&m[704])|(m[698]&m[701]&~m[702]&~m[703]&m[704])|(m[698]&~m[701]&m[702]&~m[703]&m[704])|(~m[698]&~m[701]&~m[702]&m[703]&m[704])|(m[698]&~m[701]&~m[702]&m[703]&m[704])|(~m[698]&m[701]&~m[702]&m[703]&m[704])|(m[698]&m[701]&~m[702]&m[703]&m[704])|(~m[698]&~m[701]&m[702]&m[703]&m[704])|(m[698]&~m[701]&m[702]&m[703]&m[704])|(m[698]&m[701]&m[702]&m[703]&m[704]))):InitCond[185];
    m[705] = run?((((m[674]&~m[706]&~m[707]&~m[708]&~m[709])|(~m[674]&~m[706]&~m[707]&m[708]&~m[709])|(m[674]&m[706]&~m[707]&m[708]&~m[709])|(m[674]&~m[706]&m[707]&m[708]&~m[709])|(~m[674]&m[706]&~m[707]&~m[708]&m[709])|(~m[674]&~m[706]&m[707]&~m[708]&m[709])|(m[674]&m[706]&m[707]&~m[708]&m[709])|(~m[674]&m[706]&m[707]&m[708]&m[709]))&UnbiasedRNG[87])|((m[674]&~m[706]&~m[707]&m[708]&~m[709])|(~m[674]&~m[706]&~m[707]&~m[708]&m[709])|(m[674]&~m[706]&~m[707]&~m[708]&m[709])|(m[674]&m[706]&~m[707]&~m[708]&m[709])|(m[674]&~m[706]&m[707]&~m[708]&m[709])|(~m[674]&~m[706]&~m[707]&m[708]&m[709])|(m[674]&~m[706]&~m[707]&m[708]&m[709])|(~m[674]&m[706]&~m[707]&m[708]&m[709])|(m[674]&m[706]&~m[707]&m[708]&m[709])|(~m[674]&~m[706]&m[707]&m[708]&m[709])|(m[674]&~m[706]&m[707]&m[708]&m[709])|(m[674]&m[706]&m[707]&m[708]&m[709]))):InitCond[186];
    m[710] = run?((((m[708]&~m[711]&~m[712]&~m[713]&~m[714])|(~m[708]&~m[711]&~m[712]&m[713]&~m[714])|(m[708]&m[711]&~m[712]&m[713]&~m[714])|(m[708]&~m[711]&m[712]&m[713]&~m[714])|(~m[708]&m[711]&~m[712]&~m[713]&m[714])|(~m[708]&~m[711]&m[712]&~m[713]&m[714])|(m[708]&m[711]&m[712]&~m[713]&m[714])|(~m[708]&m[711]&m[712]&m[713]&m[714]))&UnbiasedRNG[88])|((m[708]&~m[711]&~m[712]&m[713]&~m[714])|(~m[708]&~m[711]&~m[712]&~m[713]&m[714])|(m[708]&~m[711]&~m[712]&~m[713]&m[714])|(m[708]&m[711]&~m[712]&~m[713]&m[714])|(m[708]&~m[711]&m[712]&~m[713]&m[714])|(~m[708]&~m[711]&~m[712]&m[713]&m[714])|(m[708]&~m[711]&~m[712]&m[713]&m[714])|(~m[708]&m[711]&~m[712]&m[713]&m[714])|(m[708]&m[711]&~m[712]&m[713]&m[714])|(~m[708]&~m[711]&m[712]&m[713]&m[714])|(m[708]&~m[711]&m[712]&m[713]&m[714])|(m[708]&m[711]&m[712]&m[713]&m[714]))):InitCond[187];
    m[715] = run?((((m[713]&~m[716]&~m[717]&~m[718]&~m[719])|(~m[713]&~m[716]&~m[717]&m[718]&~m[719])|(m[713]&m[716]&~m[717]&m[718]&~m[719])|(m[713]&~m[716]&m[717]&m[718]&~m[719])|(~m[713]&m[716]&~m[717]&~m[718]&m[719])|(~m[713]&~m[716]&m[717]&~m[718]&m[719])|(m[713]&m[716]&m[717]&~m[718]&m[719])|(~m[713]&m[716]&m[717]&m[718]&m[719]))&UnbiasedRNG[89])|((m[713]&~m[716]&~m[717]&m[718]&~m[719])|(~m[713]&~m[716]&~m[717]&~m[718]&m[719])|(m[713]&~m[716]&~m[717]&~m[718]&m[719])|(m[713]&m[716]&~m[717]&~m[718]&m[719])|(m[713]&~m[716]&m[717]&~m[718]&m[719])|(~m[713]&~m[716]&~m[717]&m[718]&m[719])|(m[713]&~m[716]&~m[717]&m[718]&m[719])|(~m[713]&m[716]&~m[717]&m[718]&m[719])|(m[713]&m[716]&~m[717]&m[718]&m[719])|(~m[713]&~m[716]&m[717]&m[718]&m[719])|(m[713]&~m[716]&m[717]&m[718]&m[719])|(m[713]&m[716]&m[717]&m[718]&m[719]))):InitCond[188];
    m[720] = run?((((m[718]&~m[721]&~m[722]&~m[723]&~m[724])|(~m[718]&~m[721]&~m[722]&m[723]&~m[724])|(m[718]&m[721]&~m[722]&m[723]&~m[724])|(m[718]&~m[721]&m[722]&m[723]&~m[724])|(~m[718]&m[721]&~m[722]&~m[723]&m[724])|(~m[718]&~m[721]&m[722]&~m[723]&m[724])|(m[718]&m[721]&m[722]&~m[723]&m[724])|(~m[718]&m[721]&m[722]&m[723]&m[724]))&UnbiasedRNG[90])|((m[718]&~m[721]&~m[722]&m[723]&~m[724])|(~m[718]&~m[721]&~m[722]&~m[723]&m[724])|(m[718]&~m[721]&~m[722]&~m[723]&m[724])|(m[718]&m[721]&~m[722]&~m[723]&m[724])|(m[718]&~m[721]&m[722]&~m[723]&m[724])|(~m[718]&~m[721]&~m[722]&m[723]&m[724])|(m[718]&~m[721]&~m[722]&m[723]&m[724])|(~m[718]&m[721]&~m[722]&m[723]&m[724])|(m[718]&m[721]&~m[722]&m[723]&m[724])|(~m[718]&~m[721]&m[722]&m[723]&m[724])|(m[718]&~m[721]&m[722]&m[723]&m[724])|(m[718]&m[721]&m[722]&m[723]&m[724]))):InitCond[189];
    m[725] = run?((((m[723]&~m[726]&~m[727]&~m[728]&~m[729])|(~m[723]&~m[726]&~m[727]&m[728]&~m[729])|(m[723]&m[726]&~m[727]&m[728]&~m[729])|(m[723]&~m[726]&m[727]&m[728]&~m[729])|(~m[723]&m[726]&~m[727]&~m[728]&m[729])|(~m[723]&~m[726]&m[727]&~m[728]&m[729])|(m[723]&m[726]&m[727]&~m[728]&m[729])|(~m[723]&m[726]&m[727]&m[728]&m[729]))&UnbiasedRNG[91])|((m[723]&~m[726]&~m[727]&m[728]&~m[729])|(~m[723]&~m[726]&~m[727]&~m[728]&m[729])|(m[723]&~m[726]&~m[727]&~m[728]&m[729])|(m[723]&m[726]&~m[727]&~m[728]&m[729])|(m[723]&~m[726]&m[727]&~m[728]&m[729])|(~m[723]&~m[726]&~m[727]&m[728]&m[729])|(m[723]&~m[726]&~m[727]&m[728]&m[729])|(~m[723]&m[726]&~m[727]&m[728]&m[729])|(m[723]&m[726]&~m[727]&m[728]&m[729])|(~m[723]&~m[726]&m[727]&m[728]&m[729])|(m[723]&~m[726]&m[727]&m[728]&m[729])|(m[723]&m[726]&m[727]&m[728]&m[729]))):InitCond[190];
    m[730] = run?((((m[728]&~m[731]&~m[732]&~m[733]&~m[734])|(~m[728]&~m[731]&~m[732]&m[733]&~m[734])|(m[728]&m[731]&~m[732]&m[733]&~m[734])|(m[728]&~m[731]&m[732]&m[733]&~m[734])|(~m[728]&m[731]&~m[732]&~m[733]&m[734])|(~m[728]&~m[731]&m[732]&~m[733]&m[734])|(m[728]&m[731]&m[732]&~m[733]&m[734])|(~m[728]&m[731]&m[732]&m[733]&m[734]))&UnbiasedRNG[92])|((m[728]&~m[731]&~m[732]&m[733]&~m[734])|(~m[728]&~m[731]&~m[732]&~m[733]&m[734])|(m[728]&~m[731]&~m[732]&~m[733]&m[734])|(m[728]&m[731]&~m[732]&~m[733]&m[734])|(m[728]&~m[731]&m[732]&~m[733]&m[734])|(~m[728]&~m[731]&~m[732]&m[733]&m[734])|(m[728]&~m[731]&~m[732]&m[733]&m[734])|(~m[728]&m[731]&~m[732]&m[733]&m[734])|(m[728]&m[731]&~m[732]&m[733]&m[734])|(~m[728]&~m[731]&m[732]&m[733]&m[734])|(m[728]&~m[731]&m[732]&m[733]&m[734])|(m[728]&m[731]&m[732]&m[733]&m[734]))):InitCond[191];
    m[735] = run?((((m[709]&~m[736]&~m[737]&~m[738]&~m[739])|(~m[709]&~m[736]&~m[737]&m[738]&~m[739])|(m[709]&m[736]&~m[737]&m[738]&~m[739])|(m[709]&~m[736]&m[737]&m[738]&~m[739])|(~m[709]&m[736]&~m[737]&~m[738]&m[739])|(~m[709]&~m[736]&m[737]&~m[738]&m[739])|(m[709]&m[736]&m[737]&~m[738]&m[739])|(~m[709]&m[736]&m[737]&m[738]&m[739]))&UnbiasedRNG[93])|((m[709]&~m[736]&~m[737]&m[738]&~m[739])|(~m[709]&~m[736]&~m[737]&~m[738]&m[739])|(m[709]&~m[736]&~m[737]&~m[738]&m[739])|(m[709]&m[736]&~m[737]&~m[738]&m[739])|(m[709]&~m[736]&m[737]&~m[738]&m[739])|(~m[709]&~m[736]&~m[737]&m[738]&m[739])|(m[709]&~m[736]&~m[737]&m[738]&m[739])|(~m[709]&m[736]&~m[737]&m[738]&m[739])|(m[709]&m[736]&~m[737]&m[738]&m[739])|(~m[709]&~m[736]&m[737]&m[738]&m[739])|(m[709]&~m[736]&m[737]&m[738]&m[739])|(m[709]&m[736]&m[737]&m[738]&m[739]))):InitCond[192];
    m[740] = run?((((m[738]&~m[741]&~m[742]&~m[743]&~m[744])|(~m[738]&~m[741]&~m[742]&m[743]&~m[744])|(m[738]&m[741]&~m[742]&m[743]&~m[744])|(m[738]&~m[741]&m[742]&m[743]&~m[744])|(~m[738]&m[741]&~m[742]&~m[743]&m[744])|(~m[738]&~m[741]&m[742]&~m[743]&m[744])|(m[738]&m[741]&m[742]&~m[743]&m[744])|(~m[738]&m[741]&m[742]&m[743]&m[744]))&UnbiasedRNG[94])|((m[738]&~m[741]&~m[742]&m[743]&~m[744])|(~m[738]&~m[741]&~m[742]&~m[743]&m[744])|(m[738]&~m[741]&~m[742]&~m[743]&m[744])|(m[738]&m[741]&~m[742]&~m[743]&m[744])|(m[738]&~m[741]&m[742]&~m[743]&m[744])|(~m[738]&~m[741]&~m[742]&m[743]&m[744])|(m[738]&~m[741]&~m[742]&m[743]&m[744])|(~m[738]&m[741]&~m[742]&m[743]&m[744])|(m[738]&m[741]&~m[742]&m[743]&m[744])|(~m[738]&~m[741]&m[742]&m[743]&m[744])|(m[738]&~m[741]&m[742]&m[743]&m[744])|(m[738]&m[741]&m[742]&m[743]&m[744]))):InitCond[193];
    m[745] = run?((((m[743]&~m[746]&~m[747]&~m[748]&~m[749])|(~m[743]&~m[746]&~m[747]&m[748]&~m[749])|(m[743]&m[746]&~m[747]&m[748]&~m[749])|(m[743]&~m[746]&m[747]&m[748]&~m[749])|(~m[743]&m[746]&~m[747]&~m[748]&m[749])|(~m[743]&~m[746]&m[747]&~m[748]&m[749])|(m[743]&m[746]&m[747]&~m[748]&m[749])|(~m[743]&m[746]&m[747]&m[748]&m[749]))&UnbiasedRNG[95])|((m[743]&~m[746]&~m[747]&m[748]&~m[749])|(~m[743]&~m[746]&~m[747]&~m[748]&m[749])|(m[743]&~m[746]&~m[747]&~m[748]&m[749])|(m[743]&m[746]&~m[747]&~m[748]&m[749])|(m[743]&~m[746]&m[747]&~m[748]&m[749])|(~m[743]&~m[746]&~m[747]&m[748]&m[749])|(m[743]&~m[746]&~m[747]&m[748]&m[749])|(~m[743]&m[746]&~m[747]&m[748]&m[749])|(m[743]&m[746]&~m[747]&m[748]&m[749])|(~m[743]&~m[746]&m[747]&m[748]&m[749])|(m[743]&~m[746]&m[747]&m[748]&m[749])|(m[743]&m[746]&m[747]&m[748]&m[749]))):InitCond[194];
    m[750] = run?((((m[748]&~m[751]&~m[752]&~m[753]&~m[754])|(~m[748]&~m[751]&~m[752]&m[753]&~m[754])|(m[748]&m[751]&~m[752]&m[753]&~m[754])|(m[748]&~m[751]&m[752]&m[753]&~m[754])|(~m[748]&m[751]&~m[752]&~m[753]&m[754])|(~m[748]&~m[751]&m[752]&~m[753]&m[754])|(m[748]&m[751]&m[752]&~m[753]&m[754])|(~m[748]&m[751]&m[752]&m[753]&m[754]))&UnbiasedRNG[96])|((m[748]&~m[751]&~m[752]&m[753]&~m[754])|(~m[748]&~m[751]&~m[752]&~m[753]&m[754])|(m[748]&~m[751]&~m[752]&~m[753]&m[754])|(m[748]&m[751]&~m[752]&~m[753]&m[754])|(m[748]&~m[751]&m[752]&~m[753]&m[754])|(~m[748]&~m[751]&~m[752]&m[753]&m[754])|(m[748]&~m[751]&~m[752]&m[753]&m[754])|(~m[748]&m[751]&~m[752]&m[753]&m[754])|(m[748]&m[751]&~m[752]&m[753]&m[754])|(~m[748]&~m[751]&m[752]&m[753]&m[754])|(m[748]&~m[751]&m[752]&m[753]&m[754])|(m[748]&m[751]&m[752]&m[753]&m[754]))):InitCond[195];
    m[755] = run?((((m[753]&~m[756]&~m[757]&~m[758]&~m[759])|(~m[753]&~m[756]&~m[757]&m[758]&~m[759])|(m[753]&m[756]&~m[757]&m[758]&~m[759])|(m[753]&~m[756]&m[757]&m[758]&~m[759])|(~m[753]&m[756]&~m[757]&~m[758]&m[759])|(~m[753]&~m[756]&m[757]&~m[758]&m[759])|(m[753]&m[756]&m[757]&~m[758]&m[759])|(~m[753]&m[756]&m[757]&m[758]&m[759]))&UnbiasedRNG[97])|((m[753]&~m[756]&~m[757]&m[758]&~m[759])|(~m[753]&~m[756]&~m[757]&~m[758]&m[759])|(m[753]&~m[756]&~m[757]&~m[758]&m[759])|(m[753]&m[756]&~m[757]&~m[758]&m[759])|(m[753]&~m[756]&m[757]&~m[758]&m[759])|(~m[753]&~m[756]&~m[757]&m[758]&m[759])|(m[753]&~m[756]&~m[757]&m[758]&m[759])|(~m[753]&m[756]&~m[757]&m[758]&m[759])|(m[753]&m[756]&~m[757]&m[758]&m[759])|(~m[753]&~m[756]&m[757]&m[758]&m[759])|(m[753]&~m[756]&m[757]&m[758]&m[759])|(m[753]&m[756]&m[757]&m[758]&m[759]))):InitCond[196];
    m[760] = run?((((m[739]&~m[761]&~m[762]&~m[763]&~m[764])|(~m[739]&~m[761]&~m[762]&m[763]&~m[764])|(m[739]&m[761]&~m[762]&m[763]&~m[764])|(m[739]&~m[761]&m[762]&m[763]&~m[764])|(~m[739]&m[761]&~m[762]&~m[763]&m[764])|(~m[739]&~m[761]&m[762]&~m[763]&m[764])|(m[739]&m[761]&m[762]&~m[763]&m[764])|(~m[739]&m[761]&m[762]&m[763]&m[764]))&UnbiasedRNG[98])|((m[739]&~m[761]&~m[762]&m[763]&~m[764])|(~m[739]&~m[761]&~m[762]&~m[763]&m[764])|(m[739]&~m[761]&~m[762]&~m[763]&m[764])|(m[739]&m[761]&~m[762]&~m[763]&m[764])|(m[739]&~m[761]&m[762]&~m[763]&m[764])|(~m[739]&~m[761]&~m[762]&m[763]&m[764])|(m[739]&~m[761]&~m[762]&m[763]&m[764])|(~m[739]&m[761]&~m[762]&m[763]&m[764])|(m[739]&m[761]&~m[762]&m[763]&m[764])|(~m[739]&~m[761]&m[762]&m[763]&m[764])|(m[739]&~m[761]&m[762]&m[763]&m[764])|(m[739]&m[761]&m[762]&m[763]&m[764]))):InitCond[197];
    m[765] = run?((((m[763]&~m[766]&~m[767]&~m[768]&~m[769])|(~m[763]&~m[766]&~m[767]&m[768]&~m[769])|(m[763]&m[766]&~m[767]&m[768]&~m[769])|(m[763]&~m[766]&m[767]&m[768]&~m[769])|(~m[763]&m[766]&~m[767]&~m[768]&m[769])|(~m[763]&~m[766]&m[767]&~m[768]&m[769])|(m[763]&m[766]&m[767]&~m[768]&m[769])|(~m[763]&m[766]&m[767]&m[768]&m[769]))&UnbiasedRNG[99])|((m[763]&~m[766]&~m[767]&m[768]&~m[769])|(~m[763]&~m[766]&~m[767]&~m[768]&m[769])|(m[763]&~m[766]&~m[767]&~m[768]&m[769])|(m[763]&m[766]&~m[767]&~m[768]&m[769])|(m[763]&~m[766]&m[767]&~m[768]&m[769])|(~m[763]&~m[766]&~m[767]&m[768]&m[769])|(m[763]&~m[766]&~m[767]&m[768]&m[769])|(~m[763]&m[766]&~m[767]&m[768]&m[769])|(m[763]&m[766]&~m[767]&m[768]&m[769])|(~m[763]&~m[766]&m[767]&m[768]&m[769])|(m[763]&~m[766]&m[767]&m[768]&m[769])|(m[763]&m[766]&m[767]&m[768]&m[769]))):InitCond[198];
    m[770] = run?((((m[768]&~m[771]&~m[772]&~m[773]&~m[774])|(~m[768]&~m[771]&~m[772]&m[773]&~m[774])|(m[768]&m[771]&~m[772]&m[773]&~m[774])|(m[768]&~m[771]&m[772]&m[773]&~m[774])|(~m[768]&m[771]&~m[772]&~m[773]&m[774])|(~m[768]&~m[771]&m[772]&~m[773]&m[774])|(m[768]&m[771]&m[772]&~m[773]&m[774])|(~m[768]&m[771]&m[772]&m[773]&m[774]))&UnbiasedRNG[100])|((m[768]&~m[771]&~m[772]&m[773]&~m[774])|(~m[768]&~m[771]&~m[772]&~m[773]&m[774])|(m[768]&~m[771]&~m[772]&~m[773]&m[774])|(m[768]&m[771]&~m[772]&~m[773]&m[774])|(m[768]&~m[771]&m[772]&~m[773]&m[774])|(~m[768]&~m[771]&~m[772]&m[773]&m[774])|(m[768]&~m[771]&~m[772]&m[773]&m[774])|(~m[768]&m[771]&~m[772]&m[773]&m[774])|(m[768]&m[771]&~m[772]&m[773]&m[774])|(~m[768]&~m[771]&m[772]&m[773]&m[774])|(m[768]&~m[771]&m[772]&m[773]&m[774])|(m[768]&m[771]&m[772]&m[773]&m[774]))):InitCond[199];
    m[775] = run?((((m[773]&~m[776]&~m[777]&~m[778]&~m[779])|(~m[773]&~m[776]&~m[777]&m[778]&~m[779])|(m[773]&m[776]&~m[777]&m[778]&~m[779])|(m[773]&~m[776]&m[777]&m[778]&~m[779])|(~m[773]&m[776]&~m[777]&~m[778]&m[779])|(~m[773]&~m[776]&m[777]&~m[778]&m[779])|(m[773]&m[776]&m[777]&~m[778]&m[779])|(~m[773]&m[776]&m[777]&m[778]&m[779]))&UnbiasedRNG[101])|((m[773]&~m[776]&~m[777]&m[778]&~m[779])|(~m[773]&~m[776]&~m[777]&~m[778]&m[779])|(m[773]&~m[776]&~m[777]&~m[778]&m[779])|(m[773]&m[776]&~m[777]&~m[778]&m[779])|(m[773]&~m[776]&m[777]&~m[778]&m[779])|(~m[773]&~m[776]&~m[777]&m[778]&m[779])|(m[773]&~m[776]&~m[777]&m[778]&m[779])|(~m[773]&m[776]&~m[777]&m[778]&m[779])|(m[773]&m[776]&~m[777]&m[778]&m[779])|(~m[773]&~m[776]&m[777]&m[778]&m[779])|(m[773]&~m[776]&m[777]&m[778]&m[779])|(m[773]&m[776]&m[777]&m[778]&m[779]))):InitCond[200];
    m[780] = run?((((m[764]&~m[781]&~m[782]&~m[783]&~m[784])|(~m[764]&~m[781]&~m[782]&m[783]&~m[784])|(m[764]&m[781]&~m[782]&m[783]&~m[784])|(m[764]&~m[781]&m[782]&m[783]&~m[784])|(~m[764]&m[781]&~m[782]&~m[783]&m[784])|(~m[764]&~m[781]&m[782]&~m[783]&m[784])|(m[764]&m[781]&m[782]&~m[783]&m[784])|(~m[764]&m[781]&m[782]&m[783]&m[784]))&UnbiasedRNG[102])|((m[764]&~m[781]&~m[782]&m[783]&~m[784])|(~m[764]&~m[781]&~m[782]&~m[783]&m[784])|(m[764]&~m[781]&~m[782]&~m[783]&m[784])|(m[764]&m[781]&~m[782]&~m[783]&m[784])|(m[764]&~m[781]&m[782]&~m[783]&m[784])|(~m[764]&~m[781]&~m[782]&m[783]&m[784])|(m[764]&~m[781]&~m[782]&m[783]&m[784])|(~m[764]&m[781]&~m[782]&m[783]&m[784])|(m[764]&m[781]&~m[782]&m[783]&m[784])|(~m[764]&~m[781]&m[782]&m[783]&m[784])|(m[764]&~m[781]&m[782]&m[783]&m[784])|(m[764]&m[781]&m[782]&m[783]&m[784]))):InitCond[201];
    m[785] = run?((((m[783]&~m[786]&~m[787]&~m[788]&~m[789])|(~m[783]&~m[786]&~m[787]&m[788]&~m[789])|(m[783]&m[786]&~m[787]&m[788]&~m[789])|(m[783]&~m[786]&m[787]&m[788]&~m[789])|(~m[783]&m[786]&~m[787]&~m[788]&m[789])|(~m[783]&~m[786]&m[787]&~m[788]&m[789])|(m[783]&m[786]&m[787]&~m[788]&m[789])|(~m[783]&m[786]&m[787]&m[788]&m[789]))&UnbiasedRNG[103])|((m[783]&~m[786]&~m[787]&m[788]&~m[789])|(~m[783]&~m[786]&~m[787]&~m[788]&m[789])|(m[783]&~m[786]&~m[787]&~m[788]&m[789])|(m[783]&m[786]&~m[787]&~m[788]&m[789])|(m[783]&~m[786]&m[787]&~m[788]&m[789])|(~m[783]&~m[786]&~m[787]&m[788]&m[789])|(m[783]&~m[786]&~m[787]&m[788]&m[789])|(~m[783]&m[786]&~m[787]&m[788]&m[789])|(m[783]&m[786]&~m[787]&m[788]&m[789])|(~m[783]&~m[786]&m[787]&m[788]&m[789])|(m[783]&~m[786]&m[787]&m[788]&m[789])|(m[783]&m[786]&m[787]&m[788]&m[789]))):InitCond[202];
    m[790] = run?((((m[788]&~m[791]&~m[792]&~m[793]&~m[794])|(~m[788]&~m[791]&~m[792]&m[793]&~m[794])|(m[788]&m[791]&~m[792]&m[793]&~m[794])|(m[788]&~m[791]&m[792]&m[793]&~m[794])|(~m[788]&m[791]&~m[792]&~m[793]&m[794])|(~m[788]&~m[791]&m[792]&~m[793]&m[794])|(m[788]&m[791]&m[792]&~m[793]&m[794])|(~m[788]&m[791]&m[792]&m[793]&m[794]))&UnbiasedRNG[104])|((m[788]&~m[791]&~m[792]&m[793]&~m[794])|(~m[788]&~m[791]&~m[792]&~m[793]&m[794])|(m[788]&~m[791]&~m[792]&~m[793]&m[794])|(m[788]&m[791]&~m[792]&~m[793]&m[794])|(m[788]&~m[791]&m[792]&~m[793]&m[794])|(~m[788]&~m[791]&~m[792]&m[793]&m[794])|(m[788]&~m[791]&~m[792]&m[793]&m[794])|(~m[788]&m[791]&~m[792]&m[793]&m[794])|(m[788]&m[791]&~m[792]&m[793]&m[794])|(~m[788]&~m[791]&m[792]&m[793]&m[794])|(m[788]&~m[791]&m[792]&m[793]&m[794])|(m[788]&m[791]&m[792]&m[793]&m[794]))):InitCond[203];
    m[795] = run?((((m[784]&~m[796]&~m[797]&~m[798]&~m[799])|(~m[784]&~m[796]&~m[797]&m[798]&~m[799])|(m[784]&m[796]&~m[797]&m[798]&~m[799])|(m[784]&~m[796]&m[797]&m[798]&~m[799])|(~m[784]&m[796]&~m[797]&~m[798]&m[799])|(~m[784]&~m[796]&m[797]&~m[798]&m[799])|(m[784]&m[796]&m[797]&~m[798]&m[799])|(~m[784]&m[796]&m[797]&m[798]&m[799]))&UnbiasedRNG[105])|((m[784]&~m[796]&~m[797]&m[798]&~m[799])|(~m[784]&~m[796]&~m[797]&~m[798]&m[799])|(m[784]&~m[796]&~m[797]&~m[798]&m[799])|(m[784]&m[796]&~m[797]&~m[798]&m[799])|(m[784]&~m[796]&m[797]&~m[798]&m[799])|(~m[784]&~m[796]&~m[797]&m[798]&m[799])|(m[784]&~m[796]&~m[797]&m[798]&m[799])|(~m[784]&m[796]&~m[797]&m[798]&m[799])|(m[784]&m[796]&~m[797]&m[798]&m[799])|(~m[784]&~m[796]&m[797]&m[798]&m[799])|(m[784]&~m[796]&m[797]&m[798]&m[799])|(m[784]&m[796]&m[797]&m[798]&m[799]))):InitCond[204];
    m[800] = run?((((m[798]&~m[801]&~m[802]&~m[803]&~m[804])|(~m[798]&~m[801]&~m[802]&m[803]&~m[804])|(m[798]&m[801]&~m[802]&m[803]&~m[804])|(m[798]&~m[801]&m[802]&m[803]&~m[804])|(~m[798]&m[801]&~m[802]&~m[803]&m[804])|(~m[798]&~m[801]&m[802]&~m[803]&m[804])|(m[798]&m[801]&m[802]&~m[803]&m[804])|(~m[798]&m[801]&m[802]&m[803]&m[804]))&UnbiasedRNG[106])|((m[798]&~m[801]&~m[802]&m[803]&~m[804])|(~m[798]&~m[801]&~m[802]&~m[803]&m[804])|(m[798]&~m[801]&~m[802]&~m[803]&m[804])|(m[798]&m[801]&~m[802]&~m[803]&m[804])|(m[798]&~m[801]&m[802]&~m[803]&m[804])|(~m[798]&~m[801]&~m[802]&m[803]&m[804])|(m[798]&~m[801]&~m[802]&m[803]&m[804])|(~m[798]&m[801]&~m[802]&m[803]&m[804])|(m[798]&m[801]&~m[802]&m[803]&m[804])|(~m[798]&~m[801]&m[802]&m[803]&m[804])|(m[798]&~m[801]&m[802]&m[803]&m[804])|(m[798]&m[801]&m[802]&m[803]&m[804]))):InitCond[205];
    m[805] = run?((((m[799]&~m[806]&~m[807]&~m[808]&~m[809])|(~m[799]&~m[806]&~m[807]&m[808]&~m[809])|(m[799]&m[806]&~m[807]&m[808]&~m[809])|(m[799]&~m[806]&m[807]&m[808]&~m[809])|(~m[799]&m[806]&~m[807]&~m[808]&m[809])|(~m[799]&~m[806]&m[807]&~m[808]&m[809])|(m[799]&m[806]&m[807]&~m[808]&m[809])|(~m[799]&m[806]&m[807]&m[808]&m[809]))&UnbiasedRNG[107])|((m[799]&~m[806]&~m[807]&m[808]&~m[809])|(~m[799]&~m[806]&~m[807]&~m[808]&m[809])|(m[799]&~m[806]&~m[807]&~m[808]&m[809])|(m[799]&m[806]&~m[807]&~m[808]&m[809])|(m[799]&~m[806]&m[807]&~m[808]&m[809])|(~m[799]&~m[806]&~m[807]&m[808]&m[809])|(m[799]&~m[806]&~m[807]&m[808]&m[809])|(~m[799]&m[806]&~m[807]&m[808]&m[809])|(m[799]&m[806]&~m[807]&m[808]&m[809])|(~m[799]&~m[806]&m[807]&m[808]&m[809])|(m[799]&~m[806]&m[807]&m[808]&m[809])|(m[799]&m[806]&m[807]&m[808]&m[809]))):InitCond[206];
end

always @(posedge color1_clk) begin
    m[20] = run?((((m[0]&m[62]&~m[63]&~m[64]&~m[65])|(m[0]&~m[62]&m[63]&~m[64]&~m[65])|(~m[0]&m[62]&m[63]&~m[64]&~m[65])|(m[0]&~m[62]&~m[63]&m[64]&~m[65])|(~m[0]&m[62]&~m[63]&m[64]&~m[65])|(~m[0]&~m[62]&m[63]&m[64]&~m[65])|(m[0]&~m[62]&~m[63]&~m[64]&m[65])|(~m[0]&m[62]&~m[63]&~m[64]&m[65])|(~m[0]&~m[62]&m[63]&~m[64]&m[65])|(~m[0]&~m[62]&~m[63]&m[64]&m[65]))&BiasedRNG[99])|(((m[0]&m[62]&m[63]&~m[64]&~m[65])|(m[0]&m[62]&~m[63]&m[64]&~m[65])|(m[0]&~m[62]&m[63]&m[64]&~m[65])|(~m[0]&m[62]&m[63]&m[64]&~m[65])|(m[0]&m[62]&~m[63]&~m[64]&m[65])|(m[0]&~m[62]&m[63]&~m[64]&m[65])|(~m[0]&m[62]&m[63]&~m[64]&m[65])|(m[0]&~m[62]&~m[63]&m[64]&m[65])|(~m[0]&m[62]&~m[63]&m[64]&m[65])|(~m[0]&~m[62]&m[63]&m[64]&m[65]))&~BiasedRNG[99])|((m[0]&m[62]&m[63]&m[64]&~m[65])|(m[0]&m[62]&m[63]&~m[64]&m[65])|(m[0]&m[62]&~m[63]&m[64]&m[65])|(m[0]&~m[62]&m[63]&m[64]&m[65])|(~m[0]&m[62]&m[63]&m[64]&m[65])|(m[0]&m[62]&m[63]&m[64]&m[65]))):InitCond[207];
    m[21] = run?((((m[0]&m[66]&~m[67]&~m[68]&~m[69])|(m[0]&~m[66]&m[67]&~m[68]&~m[69])|(~m[0]&m[66]&m[67]&~m[68]&~m[69])|(m[0]&~m[66]&~m[67]&m[68]&~m[69])|(~m[0]&m[66]&~m[67]&m[68]&~m[69])|(~m[0]&~m[66]&m[67]&m[68]&~m[69])|(m[0]&~m[66]&~m[67]&~m[68]&m[69])|(~m[0]&m[66]&~m[67]&~m[68]&m[69])|(~m[0]&~m[66]&m[67]&~m[68]&m[69])|(~m[0]&~m[66]&~m[67]&m[68]&m[69]))&BiasedRNG[100])|(((m[0]&m[66]&m[67]&~m[68]&~m[69])|(m[0]&m[66]&~m[67]&m[68]&~m[69])|(m[0]&~m[66]&m[67]&m[68]&~m[69])|(~m[0]&m[66]&m[67]&m[68]&~m[69])|(m[0]&m[66]&~m[67]&~m[68]&m[69])|(m[0]&~m[66]&m[67]&~m[68]&m[69])|(~m[0]&m[66]&m[67]&~m[68]&m[69])|(m[0]&~m[66]&~m[67]&m[68]&m[69])|(~m[0]&m[66]&~m[67]&m[68]&m[69])|(~m[0]&~m[66]&m[67]&m[68]&m[69]))&~BiasedRNG[100])|((m[0]&m[66]&m[67]&m[68]&~m[69])|(m[0]&m[66]&m[67]&~m[68]&m[69])|(m[0]&m[66]&~m[67]&m[68]&m[69])|(m[0]&~m[66]&m[67]&m[68]&m[69])|(~m[0]&m[66]&m[67]&m[68]&m[69])|(m[0]&m[66]&m[67]&m[68]&m[69]))):InitCond[208];
    m[22] = run?((((m[1]&m[72]&~m[73]&~m[74]&~m[75])|(m[1]&~m[72]&m[73]&~m[74]&~m[75])|(~m[1]&m[72]&m[73]&~m[74]&~m[75])|(m[1]&~m[72]&~m[73]&m[74]&~m[75])|(~m[1]&m[72]&~m[73]&m[74]&~m[75])|(~m[1]&~m[72]&m[73]&m[74]&~m[75])|(m[1]&~m[72]&~m[73]&~m[74]&m[75])|(~m[1]&m[72]&~m[73]&~m[74]&m[75])|(~m[1]&~m[72]&m[73]&~m[74]&m[75])|(~m[1]&~m[72]&~m[73]&m[74]&m[75]))&BiasedRNG[101])|(((m[1]&m[72]&m[73]&~m[74]&~m[75])|(m[1]&m[72]&~m[73]&m[74]&~m[75])|(m[1]&~m[72]&m[73]&m[74]&~m[75])|(~m[1]&m[72]&m[73]&m[74]&~m[75])|(m[1]&m[72]&~m[73]&~m[74]&m[75])|(m[1]&~m[72]&m[73]&~m[74]&m[75])|(~m[1]&m[72]&m[73]&~m[74]&m[75])|(m[1]&~m[72]&~m[73]&m[74]&m[75])|(~m[1]&m[72]&~m[73]&m[74]&m[75])|(~m[1]&~m[72]&m[73]&m[74]&m[75]))&~BiasedRNG[101])|((m[1]&m[72]&m[73]&m[74]&~m[75])|(m[1]&m[72]&m[73]&~m[74]&m[75])|(m[1]&m[72]&~m[73]&m[74]&m[75])|(m[1]&~m[72]&m[73]&m[74]&m[75])|(~m[1]&m[72]&m[73]&m[74]&m[75])|(m[1]&m[72]&m[73]&m[74]&m[75]))):InitCond[209];
    m[23] = run?((((m[1]&m[76]&~m[77]&~m[78]&~m[79])|(m[1]&~m[76]&m[77]&~m[78]&~m[79])|(~m[1]&m[76]&m[77]&~m[78]&~m[79])|(m[1]&~m[76]&~m[77]&m[78]&~m[79])|(~m[1]&m[76]&~m[77]&m[78]&~m[79])|(~m[1]&~m[76]&m[77]&m[78]&~m[79])|(m[1]&~m[76]&~m[77]&~m[78]&m[79])|(~m[1]&m[76]&~m[77]&~m[78]&m[79])|(~m[1]&~m[76]&m[77]&~m[78]&m[79])|(~m[1]&~m[76]&~m[77]&m[78]&m[79]))&BiasedRNG[102])|(((m[1]&m[76]&m[77]&~m[78]&~m[79])|(m[1]&m[76]&~m[77]&m[78]&~m[79])|(m[1]&~m[76]&m[77]&m[78]&~m[79])|(~m[1]&m[76]&m[77]&m[78]&~m[79])|(m[1]&m[76]&~m[77]&~m[78]&m[79])|(m[1]&~m[76]&m[77]&~m[78]&m[79])|(~m[1]&m[76]&m[77]&~m[78]&m[79])|(m[1]&~m[76]&~m[77]&m[78]&m[79])|(~m[1]&m[76]&~m[77]&m[78]&m[79])|(~m[1]&~m[76]&m[77]&m[78]&m[79]))&~BiasedRNG[102])|((m[1]&m[76]&m[77]&m[78]&~m[79])|(m[1]&m[76]&m[77]&~m[78]&m[79])|(m[1]&m[76]&~m[77]&m[78]&m[79])|(m[1]&~m[76]&m[77]&m[78]&m[79])|(~m[1]&m[76]&m[77]&m[78]&m[79])|(m[1]&m[76]&m[77]&m[78]&m[79]))):InitCond[210];
    m[24] = run?((((m[2]&m[82]&~m[83]&~m[84]&~m[85])|(m[2]&~m[82]&m[83]&~m[84]&~m[85])|(~m[2]&m[82]&m[83]&~m[84]&~m[85])|(m[2]&~m[82]&~m[83]&m[84]&~m[85])|(~m[2]&m[82]&~m[83]&m[84]&~m[85])|(~m[2]&~m[82]&m[83]&m[84]&~m[85])|(m[2]&~m[82]&~m[83]&~m[84]&m[85])|(~m[2]&m[82]&~m[83]&~m[84]&m[85])|(~m[2]&~m[82]&m[83]&~m[84]&m[85])|(~m[2]&~m[82]&~m[83]&m[84]&m[85]))&BiasedRNG[103])|(((m[2]&m[82]&m[83]&~m[84]&~m[85])|(m[2]&m[82]&~m[83]&m[84]&~m[85])|(m[2]&~m[82]&m[83]&m[84]&~m[85])|(~m[2]&m[82]&m[83]&m[84]&~m[85])|(m[2]&m[82]&~m[83]&~m[84]&m[85])|(m[2]&~m[82]&m[83]&~m[84]&m[85])|(~m[2]&m[82]&m[83]&~m[84]&m[85])|(m[2]&~m[82]&~m[83]&m[84]&m[85])|(~m[2]&m[82]&~m[83]&m[84]&m[85])|(~m[2]&~m[82]&m[83]&m[84]&m[85]))&~BiasedRNG[103])|((m[2]&m[82]&m[83]&m[84]&~m[85])|(m[2]&m[82]&m[83]&~m[84]&m[85])|(m[2]&m[82]&~m[83]&m[84]&m[85])|(m[2]&~m[82]&m[83]&m[84]&m[85])|(~m[2]&m[82]&m[83]&m[84]&m[85])|(m[2]&m[82]&m[83]&m[84]&m[85]))):InitCond[211];
    m[25] = run?((((m[2]&m[86]&~m[87]&~m[88]&~m[89])|(m[2]&~m[86]&m[87]&~m[88]&~m[89])|(~m[2]&m[86]&m[87]&~m[88]&~m[89])|(m[2]&~m[86]&~m[87]&m[88]&~m[89])|(~m[2]&m[86]&~m[87]&m[88]&~m[89])|(~m[2]&~m[86]&m[87]&m[88]&~m[89])|(m[2]&~m[86]&~m[87]&~m[88]&m[89])|(~m[2]&m[86]&~m[87]&~m[88]&m[89])|(~m[2]&~m[86]&m[87]&~m[88]&m[89])|(~m[2]&~m[86]&~m[87]&m[88]&m[89]))&BiasedRNG[104])|(((m[2]&m[86]&m[87]&~m[88]&~m[89])|(m[2]&m[86]&~m[87]&m[88]&~m[89])|(m[2]&~m[86]&m[87]&m[88]&~m[89])|(~m[2]&m[86]&m[87]&m[88]&~m[89])|(m[2]&m[86]&~m[87]&~m[88]&m[89])|(m[2]&~m[86]&m[87]&~m[88]&m[89])|(~m[2]&m[86]&m[87]&~m[88]&m[89])|(m[2]&~m[86]&~m[87]&m[88]&m[89])|(~m[2]&m[86]&~m[87]&m[88]&m[89])|(~m[2]&~m[86]&m[87]&m[88]&m[89]))&~BiasedRNG[104])|((m[2]&m[86]&m[87]&m[88]&~m[89])|(m[2]&m[86]&m[87]&~m[88]&m[89])|(m[2]&m[86]&~m[87]&m[88]&m[89])|(m[2]&~m[86]&m[87]&m[88]&m[89])|(~m[2]&m[86]&m[87]&m[88]&m[89])|(m[2]&m[86]&m[87]&m[88]&m[89]))):InitCond[212];
    m[26] = run?((((m[3]&m[92]&~m[93]&~m[94]&~m[95])|(m[3]&~m[92]&m[93]&~m[94]&~m[95])|(~m[3]&m[92]&m[93]&~m[94]&~m[95])|(m[3]&~m[92]&~m[93]&m[94]&~m[95])|(~m[3]&m[92]&~m[93]&m[94]&~m[95])|(~m[3]&~m[92]&m[93]&m[94]&~m[95])|(m[3]&~m[92]&~m[93]&~m[94]&m[95])|(~m[3]&m[92]&~m[93]&~m[94]&m[95])|(~m[3]&~m[92]&m[93]&~m[94]&m[95])|(~m[3]&~m[92]&~m[93]&m[94]&m[95]))&BiasedRNG[105])|(((m[3]&m[92]&m[93]&~m[94]&~m[95])|(m[3]&m[92]&~m[93]&m[94]&~m[95])|(m[3]&~m[92]&m[93]&m[94]&~m[95])|(~m[3]&m[92]&m[93]&m[94]&~m[95])|(m[3]&m[92]&~m[93]&~m[94]&m[95])|(m[3]&~m[92]&m[93]&~m[94]&m[95])|(~m[3]&m[92]&m[93]&~m[94]&m[95])|(m[3]&~m[92]&~m[93]&m[94]&m[95])|(~m[3]&m[92]&~m[93]&m[94]&m[95])|(~m[3]&~m[92]&m[93]&m[94]&m[95]))&~BiasedRNG[105])|((m[3]&m[92]&m[93]&m[94]&~m[95])|(m[3]&m[92]&m[93]&~m[94]&m[95])|(m[3]&m[92]&~m[93]&m[94]&m[95])|(m[3]&~m[92]&m[93]&m[94]&m[95])|(~m[3]&m[92]&m[93]&m[94]&m[95])|(m[3]&m[92]&m[93]&m[94]&m[95]))):InitCond[213];
    m[27] = run?((((m[3]&m[96]&~m[97]&~m[98]&~m[99])|(m[3]&~m[96]&m[97]&~m[98]&~m[99])|(~m[3]&m[96]&m[97]&~m[98]&~m[99])|(m[3]&~m[96]&~m[97]&m[98]&~m[99])|(~m[3]&m[96]&~m[97]&m[98]&~m[99])|(~m[3]&~m[96]&m[97]&m[98]&~m[99])|(m[3]&~m[96]&~m[97]&~m[98]&m[99])|(~m[3]&m[96]&~m[97]&~m[98]&m[99])|(~m[3]&~m[96]&m[97]&~m[98]&m[99])|(~m[3]&~m[96]&~m[97]&m[98]&m[99]))&BiasedRNG[106])|(((m[3]&m[96]&m[97]&~m[98]&~m[99])|(m[3]&m[96]&~m[97]&m[98]&~m[99])|(m[3]&~m[96]&m[97]&m[98]&~m[99])|(~m[3]&m[96]&m[97]&m[98]&~m[99])|(m[3]&m[96]&~m[97]&~m[98]&m[99])|(m[3]&~m[96]&m[97]&~m[98]&m[99])|(~m[3]&m[96]&m[97]&~m[98]&m[99])|(m[3]&~m[96]&~m[97]&m[98]&m[99])|(~m[3]&m[96]&~m[97]&m[98]&m[99])|(~m[3]&~m[96]&m[97]&m[98]&m[99]))&~BiasedRNG[106])|((m[3]&m[96]&m[97]&m[98]&~m[99])|(m[3]&m[96]&m[97]&~m[98]&m[99])|(m[3]&m[96]&~m[97]&m[98]&m[99])|(m[3]&~m[96]&m[97]&m[98]&m[99])|(~m[3]&m[96]&m[97]&m[98]&m[99])|(m[3]&m[96]&m[97]&m[98]&m[99]))):InitCond[214];
    m[28] = run?((((m[4]&m[102]&~m[103]&~m[104]&~m[105])|(m[4]&~m[102]&m[103]&~m[104]&~m[105])|(~m[4]&m[102]&m[103]&~m[104]&~m[105])|(m[4]&~m[102]&~m[103]&m[104]&~m[105])|(~m[4]&m[102]&~m[103]&m[104]&~m[105])|(~m[4]&~m[102]&m[103]&m[104]&~m[105])|(m[4]&~m[102]&~m[103]&~m[104]&m[105])|(~m[4]&m[102]&~m[103]&~m[104]&m[105])|(~m[4]&~m[102]&m[103]&~m[104]&m[105])|(~m[4]&~m[102]&~m[103]&m[104]&m[105]))&BiasedRNG[107])|(((m[4]&m[102]&m[103]&~m[104]&~m[105])|(m[4]&m[102]&~m[103]&m[104]&~m[105])|(m[4]&~m[102]&m[103]&m[104]&~m[105])|(~m[4]&m[102]&m[103]&m[104]&~m[105])|(m[4]&m[102]&~m[103]&~m[104]&m[105])|(m[4]&~m[102]&m[103]&~m[104]&m[105])|(~m[4]&m[102]&m[103]&~m[104]&m[105])|(m[4]&~m[102]&~m[103]&m[104]&m[105])|(~m[4]&m[102]&~m[103]&m[104]&m[105])|(~m[4]&~m[102]&m[103]&m[104]&m[105]))&~BiasedRNG[107])|((m[4]&m[102]&m[103]&m[104]&~m[105])|(m[4]&m[102]&m[103]&~m[104]&m[105])|(m[4]&m[102]&~m[103]&m[104]&m[105])|(m[4]&~m[102]&m[103]&m[104]&m[105])|(~m[4]&m[102]&m[103]&m[104]&m[105])|(m[4]&m[102]&m[103]&m[104]&m[105]))):InitCond[215];
    m[29] = run?((((m[4]&m[106]&~m[107]&~m[108]&~m[109])|(m[4]&~m[106]&m[107]&~m[108]&~m[109])|(~m[4]&m[106]&m[107]&~m[108]&~m[109])|(m[4]&~m[106]&~m[107]&m[108]&~m[109])|(~m[4]&m[106]&~m[107]&m[108]&~m[109])|(~m[4]&~m[106]&m[107]&m[108]&~m[109])|(m[4]&~m[106]&~m[107]&~m[108]&m[109])|(~m[4]&m[106]&~m[107]&~m[108]&m[109])|(~m[4]&~m[106]&m[107]&~m[108]&m[109])|(~m[4]&~m[106]&~m[107]&m[108]&m[109]))&BiasedRNG[108])|(((m[4]&m[106]&m[107]&~m[108]&~m[109])|(m[4]&m[106]&~m[107]&m[108]&~m[109])|(m[4]&~m[106]&m[107]&m[108]&~m[109])|(~m[4]&m[106]&m[107]&m[108]&~m[109])|(m[4]&m[106]&~m[107]&~m[108]&m[109])|(m[4]&~m[106]&m[107]&~m[108]&m[109])|(~m[4]&m[106]&m[107]&~m[108]&m[109])|(m[4]&~m[106]&~m[107]&m[108]&m[109])|(~m[4]&m[106]&~m[107]&m[108]&m[109])|(~m[4]&~m[106]&m[107]&m[108]&m[109]))&~BiasedRNG[108])|((m[4]&m[106]&m[107]&m[108]&~m[109])|(m[4]&m[106]&m[107]&~m[108]&m[109])|(m[4]&m[106]&~m[107]&m[108]&m[109])|(m[4]&~m[106]&m[107]&m[108]&m[109])|(~m[4]&m[106]&m[107]&m[108]&m[109])|(m[4]&m[106]&m[107]&m[108]&m[109]))):InitCond[216];
    m[30] = run?((((m[5]&m[112]&~m[113]&~m[114]&~m[115])|(m[5]&~m[112]&m[113]&~m[114]&~m[115])|(~m[5]&m[112]&m[113]&~m[114]&~m[115])|(m[5]&~m[112]&~m[113]&m[114]&~m[115])|(~m[5]&m[112]&~m[113]&m[114]&~m[115])|(~m[5]&~m[112]&m[113]&m[114]&~m[115])|(m[5]&~m[112]&~m[113]&~m[114]&m[115])|(~m[5]&m[112]&~m[113]&~m[114]&m[115])|(~m[5]&~m[112]&m[113]&~m[114]&m[115])|(~m[5]&~m[112]&~m[113]&m[114]&m[115]))&BiasedRNG[109])|(((m[5]&m[112]&m[113]&~m[114]&~m[115])|(m[5]&m[112]&~m[113]&m[114]&~m[115])|(m[5]&~m[112]&m[113]&m[114]&~m[115])|(~m[5]&m[112]&m[113]&m[114]&~m[115])|(m[5]&m[112]&~m[113]&~m[114]&m[115])|(m[5]&~m[112]&m[113]&~m[114]&m[115])|(~m[5]&m[112]&m[113]&~m[114]&m[115])|(m[5]&~m[112]&~m[113]&m[114]&m[115])|(~m[5]&m[112]&~m[113]&m[114]&m[115])|(~m[5]&~m[112]&m[113]&m[114]&m[115]))&~BiasedRNG[109])|((m[5]&m[112]&m[113]&m[114]&~m[115])|(m[5]&m[112]&m[113]&~m[114]&m[115])|(m[5]&m[112]&~m[113]&m[114]&m[115])|(m[5]&~m[112]&m[113]&m[114]&m[115])|(~m[5]&m[112]&m[113]&m[114]&m[115])|(m[5]&m[112]&m[113]&m[114]&m[115]))):InitCond[217];
    m[31] = run?((((m[5]&m[116]&~m[117]&~m[118]&~m[119])|(m[5]&~m[116]&m[117]&~m[118]&~m[119])|(~m[5]&m[116]&m[117]&~m[118]&~m[119])|(m[5]&~m[116]&~m[117]&m[118]&~m[119])|(~m[5]&m[116]&~m[117]&m[118]&~m[119])|(~m[5]&~m[116]&m[117]&m[118]&~m[119])|(m[5]&~m[116]&~m[117]&~m[118]&m[119])|(~m[5]&m[116]&~m[117]&~m[118]&m[119])|(~m[5]&~m[116]&m[117]&~m[118]&m[119])|(~m[5]&~m[116]&~m[117]&m[118]&m[119]))&BiasedRNG[110])|(((m[5]&m[116]&m[117]&~m[118]&~m[119])|(m[5]&m[116]&~m[117]&m[118]&~m[119])|(m[5]&~m[116]&m[117]&m[118]&~m[119])|(~m[5]&m[116]&m[117]&m[118]&~m[119])|(m[5]&m[116]&~m[117]&~m[118]&m[119])|(m[5]&~m[116]&m[117]&~m[118]&m[119])|(~m[5]&m[116]&m[117]&~m[118]&m[119])|(m[5]&~m[116]&~m[117]&m[118]&m[119])|(~m[5]&m[116]&~m[117]&m[118]&m[119])|(~m[5]&~m[116]&m[117]&m[118]&m[119]))&~BiasedRNG[110])|((m[5]&m[116]&m[117]&m[118]&~m[119])|(m[5]&m[116]&m[117]&~m[118]&m[119])|(m[5]&m[116]&~m[117]&m[118]&m[119])|(m[5]&~m[116]&m[117]&m[118]&m[119])|(~m[5]&m[116]&m[117]&m[118]&m[119])|(m[5]&m[116]&m[117]&m[118]&m[119]))):InitCond[218];
    m[32] = run?((((m[6]&m[122]&~m[123]&~m[124]&~m[125])|(m[6]&~m[122]&m[123]&~m[124]&~m[125])|(~m[6]&m[122]&m[123]&~m[124]&~m[125])|(m[6]&~m[122]&~m[123]&m[124]&~m[125])|(~m[6]&m[122]&~m[123]&m[124]&~m[125])|(~m[6]&~m[122]&m[123]&m[124]&~m[125])|(m[6]&~m[122]&~m[123]&~m[124]&m[125])|(~m[6]&m[122]&~m[123]&~m[124]&m[125])|(~m[6]&~m[122]&m[123]&~m[124]&m[125])|(~m[6]&~m[122]&~m[123]&m[124]&m[125]))&BiasedRNG[111])|(((m[6]&m[122]&m[123]&~m[124]&~m[125])|(m[6]&m[122]&~m[123]&m[124]&~m[125])|(m[6]&~m[122]&m[123]&m[124]&~m[125])|(~m[6]&m[122]&m[123]&m[124]&~m[125])|(m[6]&m[122]&~m[123]&~m[124]&m[125])|(m[6]&~m[122]&m[123]&~m[124]&m[125])|(~m[6]&m[122]&m[123]&~m[124]&m[125])|(m[6]&~m[122]&~m[123]&m[124]&m[125])|(~m[6]&m[122]&~m[123]&m[124]&m[125])|(~m[6]&~m[122]&m[123]&m[124]&m[125]))&~BiasedRNG[111])|((m[6]&m[122]&m[123]&m[124]&~m[125])|(m[6]&m[122]&m[123]&~m[124]&m[125])|(m[6]&m[122]&~m[123]&m[124]&m[125])|(m[6]&~m[122]&m[123]&m[124]&m[125])|(~m[6]&m[122]&m[123]&m[124]&m[125])|(m[6]&m[122]&m[123]&m[124]&m[125]))):InitCond[219];
    m[33] = run?((((m[6]&m[126]&~m[127]&~m[128]&~m[129])|(m[6]&~m[126]&m[127]&~m[128]&~m[129])|(~m[6]&m[126]&m[127]&~m[128]&~m[129])|(m[6]&~m[126]&~m[127]&m[128]&~m[129])|(~m[6]&m[126]&~m[127]&m[128]&~m[129])|(~m[6]&~m[126]&m[127]&m[128]&~m[129])|(m[6]&~m[126]&~m[127]&~m[128]&m[129])|(~m[6]&m[126]&~m[127]&~m[128]&m[129])|(~m[6]&~m[126]&m[127]&~m[128]&m[129])|(~m[6]&~m[126]&~m[127]&m[128]&m[129]))&BiasedRNG[112])|(((m[6]&m[126]&m[127]&~m[128]&~m[129])|(m[6]&m[126]&~m[127]&m[128]&~m[129])|(m[6]&~m[126]&m[127]&m[128]&~m[129])|(~m[6]&m[126]&m[127]&m[128]&~m[129])|(m[6]&m[126]&~m[127]&~m[128]&m[129])|(m[6]&~m[126]&m[127]&~m[128]&m[129])|(~m[6]&m[126]&m[127]&~m[128]&m[129])|(m[6]&~m[126]&~m[127]&m[128]&m[129])|(~m[6]&m[126]&~m[127]&m[128]&m[129])|(~m[6]&~m[126]&m[127]&m[128]&m[129]))&~BiasedRNG[112])|((m[6]&m[126]&m[127]&m[128]&~m[129])|(m[6]&m[126]&m[127]&~m[128]&m[129])|(m[6]&m[126]&~m[127]&m[128]&m[129])|(m[6]&~m[126]&m[127]&m[128]&m[129])|(~m[6]&m[126]&m[127]&m[128]&m[129])|(m[6]&m[126]&m[127]&m[128]&m[129]))):InitCond[220];
    m[34] = run?((((m[7]&m[132]&~m[133]&~m[134]&~m[135])|(m[7]&~m[132]&m[133]&~m[134]&~m[135])|(~m[7]&m[132]&m[133]&~m[134]&~m[135])|(m[7]&~m[132]&~m[133]&m[134]&~m[135])|(~m[7]&m[132]&~m[133]&m[134]&~m[135])|(~m[7]&~m[132]&m[133]&m[134]&~m[135])|(m[7]&~m[132]&~m[133]&~m[134]&m[135])|(~m[7]&m[132]&~m[133]&~m[134]&m[135])|(~m[7]&~m[132]&m[133]&~m[134]&m[135])|(~m[7]&~m[132]&~m[133]&m[134]&m[135]))&BiasedRNG[113])|(((m[7]&m[132]&m[133]&~m[134]&~m[135])|(m[7]&m[132]&~m[133]&m[134]&~m[135])|(m[7]&~m[132]&m[133]&m[134]&~m[135])|(~m[7]&m[132]&m[133]&m[134]&~m[135])|(m[7]&m[132]&~m[133]&~m[134]&m[135])|(m[7]&~m[132]&m[133]&~m[134]&m[135])|(~m[7]&m[132]&m[133]&~m[134]&m[135])|(m[7]&~m[132]&~m[133]&m[134]&m[135])|(~m[7]&m[132]&~m[133]&m[134]&m[135])|(~m[7]&~m[132]&m[133]&m[134]&m[135]))&~BiasedRNG[113])|((m[7]&m[132]&m[133]&m[134]&~m[135])|(m[7]&m[132]&m[133]&~m[134]&m[135])|(m[7]&m[132]&~m[133]&m[134]&m[135])|(m[7]&~m[132]&m[133]&m[134]&m[135])|(~m[7]&m[132]&m[133]&m[134]&m[135])|(m[7]&m[132]&m[133]&m[134]&m[135]))):InitCond[221];
    m[35] = run?((((m[7]&m[136]&~m[137]&~m[138]&~m[139])|(m[7]&~m[136]&m[137]&~m[138]&~m[139])|(~m[7]&m[136]&m[137]&~m[138]&~m[139])|(m[7]&~m[136]&~m[137]&m[138]&~m[139])|(~m[7]&m[136]&~m[137]&m[138]&~m[139])|(~m[7]&~m[136]&m[137]&m[138]&~m[139])|(m[7]&~m[136]&~m[137]&~m[138]&m[139])|(~m[7]&m[136]&~m[137]&~m[138]&m[139])|(~m[7]&~m[136]&m[137]&~m[138]&m[139])|(~m[7]&~m[136]&~m[137]&m[138]&m[139]))&BiasedRNG[114])|(((m[7]&m[136]&m[137]&~m[138]&~m[139])|(m[7]&m[136]&~m[137]&m[138]&~m[139])|(m[7]&~m[136]&m[137]&m[138]&~m[139])|(~m[7]&m[136]&m[137]&m[138]&~m[139])|(m[7]&m[136]&~m[137]&~m[138]&m[139])|(m[7]&~m[136]&m[137]&~m[138]&m[139])|(~m[7]&m[136]&m[137]&~m[138]&m[139])|(m[7]&~m[136]&~m[137]&m[138]&m[139])|(~m[7]&m[136]&~m[137]&m[138]&m[139])|(~m[7]&~m[136]&m[137]&m[138]&m[139]))&~BiasedRNG[114])|((m[7]&m[136]&m[137]&m[138]&~m[139])|(m[7]&m[136]&m[137]&~m[138]&m[139])|(m[7]&m[136]&~m[137]&m[138]&m[139])|(m[7]&~m[136]&m[137]&m[138]&m[139])|(~m[7]&m[136]&m[137]&m[138]&m[139])|(m[7]&m[136]&m[137]&m[138]&m[139]))):InitCond[222];
    m[36] = run?((((m[8]&m[142]&~m[143]&~m[144]&~m[145])|(m[8]&~m[142]&m[143]&~m[144]&~m[145])|(~m[8]&m[142]&m[143]&~m[144]&~m[145])|(m[8]&~m[142]&~m[143]&m[144]&~m[145])|(~m[8]&m[142]&~m[143]&m[144]&~m[145])|(~m[8]&~m[142]&m[143]&m[144]&~m[145])|(m[8]&~m[142]&~m[143]&~m[144]&m[145])|(~m[8]&m[142]&~m[143]&~m[144]&m[145])|(~m[8]&~m[142]&m[143]&~m[144]&m[145])|(~m[8]&~m[142]&~m[143]&m[144]&m[145]))&BiasedRNG[115])|(((m[8]&m[142]&m[143]&~m[144]&~m[145])|(m[8]&m[142]&~m[143]&m[144]&~m[145])|(m[8]&~m[142]&m[143]&m[144]&~m[145])|(~m[8]&m[142]&m[143]&m[144]&~m[145])|(m[8]&m[142]&~m[143]&~m[144]&m[145])|(m[8]&~m[142]&m[143]&~m[144]&m[145])|(~m[8]&m[142]&m[143]&~m[144]&m[145])|(m[8]&~m[142]&~m[143]&m[144]&m[145])|(~m[8]&m[142]&~m[143]&m[144]&m[145])|(~m[8]&~m[142]&m[143]&m[144]&m[145]))&~BiasedRNG[115])|((m[8]&m[142]&m[143]&m[144]&~m[145])|(m[8]&m[142]&m[143]&~m[144]&m[145])|(m[8]&m[142]&~m[143]&m[144]&m[145])|(m[8]&~m[142]&m[143]&m[144]&m[145])|(~m[8]&m[142]&m[143]&m[144]&m[145])|(m[8]&m[142]&m[143]&m[144]&m[145]))):InitCond[223];
    m[37] = run?((((m[8]&m[146]&~m[147]&~m[148]&~m[149])|(m[8]&~m[146]&m[147]&~m[148]&~m[149])|(~m[8]&m[146]&m[147]&~m[148]&~m[149])|(m[8]&~m[146]&~m[147]&m[148]&~m[149])|(~m[8]&m[146]&~m[147]&m[148]&~m[149])|(~m[8]&~m[146]&m[147]&m[148]&~m[149])|(m[8]&~m[146]&~m[147]&~m[148]&m[149])|(~m[8]&m[146]&~m[147]&~m[148]&m[149])|(~m[8]&~m[146]&m[147]&~m[148]&m[149])|(~m[8]&~m[146]&~m[147]&m[148]&m[149]))&BiasedRNG[116])|(((m[8]&m[146]&m[147]&~m[148]&~m[149])|(m[8]&m[146]&~m[147]&m[148]&~m[149])|(m[8]&~m[146]&m[147]&m[148]&~m[149])|(~m[8]&m[146]&m[147]&m[148]&~m[149])|(m[8]&m[146]&~m[147]&~m[148]&m[149])|(m[8]&~m[146]&m[147]&~m[148]&m[149])|(~m[8]&m[146]&m[147]&~m[148]&m[149])|(m[8]&~m[146]&~m[147]&m[148]&m[149])|(~m[8]&m[146]&~m[147]&m[148]&m[149])|(~m[8]&~m[146]&m[147]&m[148]&m[149]))&~BiasedRNG[116])|((m[8]&m[146]&m[147]&m[148]&~m[149])|(m[8]&m[146]&m[147]&~m[148]&m[149])|(m[8]&m[146]&~m[147]&m[148]&m[149])|(m[8]&~m[146]&m[147]&m[148]&m[149])|(~m[8]&m[146]&m[147]&m[148]&m[149])|(m[8]&m[146]&m[147]&m[148]&m[149]))):InitCond[224];
    m[38] = run?((((m[9]&m[152]&~m[153]&~m[154]&~m[155])|(m[9]&~m[152]&m[153]&~m[154]&~m[155])|(~m[9]&m[152]&m[153]&~m[154]&~m[155])|(m[9]&~m[152]&~m[153]&m[154]&~m[155])|(~m[9]&m[152]&~m[153]&m[154]&~m[155])|(~m[9]&~m[152]&m[153]&m[154]&~m[155])|(m[9]&~m[152]&~m[153]&~m[154]&m[155])|(~m[9]&m[152]&~m[153]&~m[154]&m[155])|(~m[9]&~m[152]&m[153]&~m[154]&m[155])|(~m[9]&~m[152]&~m[153]&m[154]&m[155]))&BiasedRNG[117])|(((m[9]&m[152]&m[153]&~m[154]&~m[155])|(m[9]&m[152]&~m[153]&m[154]&~m[155])|(m[9]&~m[152]&m[153]&m[154]&~m[155])|(~m[9]&m[152]&m[153]&m[154]&~m[155])|(m[9]&m[152]&~m[153]&~m[154]&m[155])|(m[9]&~m[152]&m[153]&~m[154]&m[155])|(~m[9]&m[152]&m[153]&~m[154]&m[155])|(m[9]&~m[152]&~m[153]&m[154]&m[155])|(~m[9]&m[152]&~m[153]&m[154]&m[155])|(~m[9]&~m[152]&m[153]&m[154]&m[155]))&~BiasedRNG[117])|((m[9]&m[152]&m[153]&m[154]&~m[155])|(m[9]&m[152]&m[153]&~m[154]&m[155])|(m[9]&m[152]&~m[153]&m[154]&m[155])|(m[9]&~m[152]&m[153]&m[154]&m[155])|(~m[9]&m[152]&m[153]&m[154]&m[155])|(m[9]&m[152]&m[153]&m[154]&m[155]))):InitCond[225];
    m[39] = run?((((m[9]&m[156]&~m[157]&~m[158]&~m[159])|(m[9]&~m[156]&m[157]&~m[158]&~m[159])|(~m[9]&m[156]&m[157]&~m[158]&~m[159])|(m[9]&~m[156]&~m[157]&m[158]&~m[159])|(~m[9]&m[156]&~m[157]&m[158]&~m[159])|(~m[9]&~m[156]&m[157]&m[158]&~m[159])|(m[9]&~m[156]&~m[157]&~m[158]&m[159])|(~m[9]&m[156]&~m[157]&~m[158]&m[159])|(~m[9]&~m[156]&m[157]&~m[158]&m[159])|(~m[9]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[118])|(((m[9]&m[156]&m[157]&~m[158]&~m[159])|(m[9]&m[156]&~m[157]&m[158]&~m[159])|(m[9]&~m[156]&m[157]&m[158]&~m[159])|(~m[9]&m[156]&m[157]&m[158]&~m[159])|(m[9]&m[156]&~m[157]&~m[158]&m[159])|(m[9]&~m[156]&m[157]&~m[158]&m[159])|(~m[9]&m[156]&m[157]&~m[158]&m[159])|(m[9]&~m[156]&~m[157]&m[158]&m[159])|(~m[9]&m[156]&~m[157]&m[158]&m[159])|(~m[9]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[118])|((m[9]&m[156]&m[157]&m[158]&~m[159])|(m[9]&m[156]&m[157]&~m[158]&m[159])|(m[9]&m[156]&~m[157]&m[158]&m[159])|(m[9]&~m[156]&m[157]&m[158]&m[159])|(~m[9]&m[156]&m[157]&m[158]&m[159])|(m[9]&m[156]&m[157]&m[158]&m[159]))):InitCond[226];
    m[40] = run?((((m[10]&m[162]&~m[163]&~m[164]&~m[165])|(m[10]&~m[162]&m[163]&~m[164]&~m[165])|(~m[10]&m[162]&m[163]&~m[164]&~m[165])|(m[10]&~m[162]&~m[163]&m[164]&~m[165])|(~m[10]&m[162]&~m[163]&m[164]&~m[165])|(~m[10]&~m[162]&m[163]&m[164]&~m[165])|(m[10]&~m[162]&~m[163]&~m[164]&m[165])|(~m[10]&m[162]&~m[163]&~m[164]&m[165])|(~m[10]&~m[162]&m[163]&~m[164]&m[165])|(~m[10]&~m[162]&~m[163]&m[164]&m[165]))&BiasedRNG[119])|(((m[10]&m[162]&m[163]&~m[164]&~m[165])|(m[10]&m[162]&~m[163]&m[164]&~m[165])|(m[10]&~m[162]&m[163]&m[164]&~m[165])|(~m[10]&m[162]&m[163]&m[164]&~m[165])|(m[10]&m[162]&~m[163]&~m[164]&m[165])|(m[10]&~m[162]&m[163]&~m[164]&m[165])|(~m[10]&m[162]&m[163]&~m[164]&m[165])|(m[10]&~m[162]&~m[163]&m[164]&m[165])|(~m[10]&m[162]&~m[163]&m[164]&m[165])|(~m[10]&~m[162]&m[163]&m[164]&m[165]))&~BiasedRNG[119])|((m[10]&m[162]&m[163]&m[164]&~m[165])|(m[10]&m[162]&m[163]&~m[164]&m[165])|(m[10]&m[162]&~m[163]&m[164]&m[165])|(m[10]&~m[162]&m[163]&m[164]&m[165])|(~m[10]&m[162]&m[163]&m[164]&m[165])|(m[10]&m[162]&m[163]&m[164]&m[165]))):InitCond[227];
    m[41] = run?((((m[10]&m[166]&~m[167]&~m[168]&~m[169])|(m[10]&~m[166]&m[167]&~m[168]&~m[169])|(~m[10]&m[166]&m[167]&~m[168]&~m[169])|(m[10]&~m[166]&~m[167]&m[168]&~m[169])|(~m[10]&m[166]&~m[167]&m[168]&~m[169])|(~m[10]&~m[166]&m[167]&m[168]&~m[169])|(m[10]&~m[166]&~m[167]&~m[168]&m[169])|(~m[10]&m[166]&~m[167]&~m[168]&m[169])|(~m[10]&~m[166]&m[167]&~m[168]&m[169])|(~m[10]&~m[166]&~m[167]&m[168]&m[169]))&BiasedRNG[120])|(((m[10]&m[166]&m[167]&~m[168]&~m[169])|(m[10]&m[166]&~m[167]&m[168]&~m[169])|(m[10]&~m[166]&m[167]&m[168]&~m[169])|(~m[10]&m[166]&m[167]&m[168]&~m[169])|(m[10]&m[166]&~m[167]&~m[168]&m[169])|(m[10]&~m[166]&m[167]&~m[168]&m[169])|(~m[10]&m[166]&m[167]&~m[168]&m[169])|(m[10]&~m[166]&~m[167]&m[168]&m[169])|(~m[10]&m[166]&~m[167]&m[168]&m[169])|(~m[10]&~m[166]&m[167]&m[168]&m[169]))&~BiasedRNG[120])|((m[10]&m[166]&m[167]&m[168]&~m[169])|(m[10]&m[166]&m[167]&~m[168]&m[169])|(m[10]&m[166]&~m[167]&m[168]&m[169])|(m[10]&~m[166]&m[167]&m[168]&m[169])|(~m[10]&m[166]&m[167]&m[168]&m[169])|(m[10]&m[166]&m[167]&m[168]&m[169]))):InitCond[228];
    m[42] = run?((((m[11]&m[172]&~m[173]&~m[174]&~m[175])|(m[11]&~m[172]&m[173]&~m[174]&~m[175])|(~m[11]&m[172]&m[173]&~m[174]&~m[175])|(m[11]&~m[172]&~m[173]&m[174]&~m[175])|(~m[11]&m[172]&~m[173]&m[174]&~m[175])|(~m[11]&~m[172]&m[173]&m[174]&~m[175])|(m[11]&~m[172]&~m[173]&~m[174]&m[175])|(~m[11]&m[172]&~m[173]&~m[174]&m[175])|(~m[11]&~m[172]&m[173]&~m[174]&m[175])|(~m[11]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[121])|(((m[11]&m[172]&m[173]&~m[174]&~m[175])|(m[11]&m[172]&~m[173]&m[174]&~m[175])|(m[11]&~m[172]&m[173]&m[174]&~m[175])|(~m[11]&m[172]&m[173]&m[174]&~m[175])|(m[11]&m[172]&~m[173]&~m[174]&m[175])|(m[11]&~m[172]&m[173]&~m[174]&m[175])|(~m[11]&m[172]&m[173]&~m[174]&m[175])|(m[11]&~m[172]&~m[173]&m[174]&m[175])|(~m[11]&m[172]&~m[173]&m[174]&m[175])|(~m[11]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[121])|((m[11]&m[172]&m[173]&m[174]&~m[175])|(m[11]&m[172]&m[173]&~m[174]&m[175])|(m[11]&m[172]&~m[173]&m[174]&m[175])|(m[11]&~m[172]&m[173]&m[174]&m[175])|(~m[11]&m[172]&m[173]&m[174]&m[175])|(m[11]&m[172]&m[173]&m[174]&m[175]))):InitCond[229];
    m[43] = run?((((m[11]&m[176]&~m[177]&~m[178]&~m[179])|(m[11]&~m[176]&m[177]&~m[178]&~m[179])|(~m[11]&m[176]&m[177]&~m[178]&~m[179])|(m[11]&~m[176]&~m[177]&m[178]&~m[179])|(~m[11]&m[176]&~m[177]&m[178]&~m[179])|(~m[11]&~m[176]&m[177]&m[178]&~m[179])|(m[11]&~m[176]&~m[177]&~m[178]&m[179])|(~m[11]&m[176]&~m[177]&~m[178]&m[179])|(~m[11]&~m[176]&m[177]&~m[178]&m[179])|(~m[11]&~m[176]&~m[177]&m[178]&m[179]))&BiasedRNG[122])|(((m[11]&m[176]&m[177]&~m[178]&~m[179])|(m[11]&m[176]&~m[177]&m[178]&~m[179])|(m[11]&~m[176]&m[177]&m[178]&~m[179])|(~m[11]&m[176]&m[177]&m[178]&~m[179])|(m[11]&m[176]&~m[177]&~m[178]&m[179])|(m[11]&~m[176]&m[177]&~m[178]&m[179])|(~m[11]&m[176]&m[177]&~m[178]&m[179])|(m[11]&~m[176]&~m[177]&m[178]&m[179])|(~m[11]&m[176]&~m[177]&m[178]&m[179])|(~m[11]&~m[176]&m[177]&m[178]&m[179]))&~BiasedRNG[122])|((m[11]&m[176]&m[177]&m[178]&~m[179])|(m[11]&m[176]&m[177]&~m[178]&m[179])|(m[11]&m[176]&~m[177]&m[178]&m[179])|(m[11]&~m[176]&m[177]&m[178]&m[179])|(~m[11]&m[176]&m[177]&m[178]&m[179])|(m[11]&m[176]&m[177]&m[178]&m[179]))):InitCond[230];
    m[44] = run?((((m[12]&m[182]&~m[183]&~m[184]&~m[185])|(m[12]&~m[182]&m[183]&~m[184]&~m[185])|(~m[12]&m[182]&m[183]&~m[184]&~m[185])|(m[12]&~m[182]&~m[183]&m[184]&~m[185])|(~m[12]&m[182]&~m[183]&m[184]&~m[185])|(~m[12]&~m[182]&m[183]&m[184]&~m[185])|(m[12]&~m[182]&~m[183]&~m[184]&m[185])|(~m[12]&m[182]&~m[183]&~m[184]&m[185])|(~m[12]&~m[182]&m[183]&~m[184]&m[185])|(~m[12]&~m[182]&~m[183]&m[184]&m[185]))&BiasedRNG[123])|(((m[12]&m[182]&m[183]&~m[184]&~m[185])|(m[12]&m[182]&~m[183]&m[184]&~m[185])|(m[12]&~m[182]&m[183]&m[184]&~m[185])|(~m[12]&m[182]&m[183]&m[184]&~m[185])|(m[12]&m[182]&~m[183]&~m[184]&m[185])|(m[12]&~m[182]&m[183]&~m[184]&m[185])|(~m[12]&m[182]&m[183]&~m[184]&m[185])|(m[12]&~m[182]&~m[183]&m[184]&m[185])|(~m[12]&m[182]&~m[183]&m[184]&m[185])|(~m[12]&~m[182]&m[183]&m[184]&m[185]))&~BiasedRNG[123])|((m[12]&m[182]&m[183]&m[184]&~m[185])|(m[12]&m[182]&m[183]&~m[184]&m[185])|(m[12]&m[182]&~m[183]&m[184]&m[185])|(m[12]&~m[182]&m[183]&m[184]&m[185])|(~m[12]&m[182]&m[183]&m[184]&m[185])|(m[12]&m[182]&m[183]&m[184]&m[185]))):InitCond[231];
    m[45] = run?((((m[12]&m[186]&~m[187]&~m[188]&~m[189])|(m[12]&~m[186]&m[187]&~m[188]&~m[189])|(~m[12]&m[186]&m[187]&~m[188]&~m[189])|(m[12]&~m[186]&~m[187]&m[188]&~m[189])|(~m[12]&m[186]&~m[187]&m[188]&~m[189])|(~m[12]&~m[186]&m[187]&m[188]&~m[189])|(m[12]&~m[186]&~m[187]&~m[188]&m[189])|(~m[12]&m[186]&~m[187]&~m[188]&m[189])|(~m[12]&~m[186]&m[187]&~m[188]&m[189])|(~m[12]&~m[186]&~m[187]&m[188]&m[189]))&BiasedRNG[124])|(((m[12]&m[186]&m[187]&~m[188]&~m[189])|(m[12]&m[186]&~m[187]&m[188]&~m[189])|(m[12]&~m[186]&m[187]&m[188]&~m[189])|(~m[12]&m[186]&m[187]&m[188]&~m[189])|(m[12]&m[186]&~m[187]&~m[188]&m[189])|(m[12]&~m[186]&m[187]&~m[188]&m[189])|(~m[12]&m[186]&m[187]&~m[188]&m[189])|(m[12]&~m[186]&~m[187]&m[188]&m[189])|(~m[12]&m[186]&~m[187]&m[188]&m[189])|(~m[12]&~m[186]&m[187]&m[188]&m[189]))&~BiasedRNG[124])|((m[12]&m[186]&m[187]&m[188]&~m[189])|(m[12]&m[186]&m[187]&~m[188]&m[189])|(m[12]&m[186]&~m[187]&m[188]&m[189])|(m[12]&~m[186]&m[187]&m[188]&m[189])|(~m[12]&m[186]&m[187]&m[188]&m[189])|(m[12]&m[186]&m[187]&m[188]&m[189]))):InitCond[232];
    m[46] = run?((((m[13]&m[192]&~m[193]&~m[194]&~m[195])|(m[13]&~m[192]&m[193]&~m[194]&~m[195])|(~m[13]&m[192]&m[193]&~m[194]&~m[195])|(m[13]&~m[192]&~m[193]&m[194]&~m[195])|(~m[13]&m[192]&~m[193]&m[194]&~m[195])|(~m[13]&~m[192]&m[193]&m[194]&~m[195])|(m[13]&~m[192]&~m[193]&~m[194]&m[195])|(~m[13]&m[192]&~m[193]&~m[194]&m[195])|(~m[13]&~m[192]&m[193]&~m[194]&m[195])|(~m[13]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[125])|(((m[13]&m[192]&m[193]&~m[194]&~m[195])|(m[13]&m[192]&~m[193]&m[194]&~m[195])|(m[13]&~m[192]&m[193]&m[194]&~m[195])|(~m[13]&m[192]&m[193]&m[194]&~m[195])|(m[13]&m[192]&~m[193]&~m[194]&m[195])|(m[13]&~m[192]&m[193]&~m[194]&m[195])|(~m[13]&m[192]&m[193]&~m[194]&m[195])|(m[13]&~m[192]&~m[193]&m[194]&m[195])|(~m[13]&m[192]&~m[193]&m[194]&m[195])|(~m[13]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[125])|((m[13]&m[192]&m[193]&m[194]&~m[195])|(m[13]&m[192]&m[193]&~m[194]&m[195])|(m[13]&m[192]&~m[193]&m[194]&m[195])|(m[13]&~m[192]&m[193]&m[194]&m[195])|(~m[13]&m[192]&m[193]&m[194]&m[195])|(m[13]&m[192]&m[193]&m[194]&m[195]))):InitCond[233];
    m[47] = run?((((m[13]&m[196]&~m[197]&~m[198]&~m[199])|(m[13]&~m[196]&m[197]&~m[198]&~m[199])|(~m[13]&m[196]&m[197]&~m[198]&~m[199])|(m[13]&~m[196]&~m[197]&m[198]&~m[199])|(~m[13]&m[196]&~m[197]&m[198]&~m[199])|(~m[13]&~m[196]&m[197]&m[198]&~m[199])|(m[13]&~m[196]&~m[197]&~m[198]&m[199])|(~m[13]&m[196]&~m[197]&~m[198]&m[199])|(~m[13]&~m[196]&m[197]&~m[198]&m[199])|(~m[13]&~m[196]&~m[197]&m[198]&m[199]))&BiasedRNG[126])|(((m[13]&m[196]&m[197]&~m[198]&~m[199])|(m[13]&m[196]&~m[197]&m[198]&~m[199])|(m[13]&~m[196]&m[197]&m[198]&~m[199])|(~m[13]&m[196]&m[197]&m[198]&~m[199])|(m[13]&m[196]&~m[197]&~m[198]&m[199])|(m[13]&~m[196]&m[197]&~m[198]&m[199])|(~m[13]&m[196]&m[197]&~m[198]&m[199])|(m[13]&~m[196]&~m[197]&m[198]&m[199])|(~m[13]&m[196]&~m[197]&m[198]&m[199])|(~m[13]&~m[196]&m[197]&m[198]&m[199]))&~BiasedRNG[126])|((m[13]&m[196]&m[197]&m[198]&~m[199])|(m[13]&m[196]&m[197]&~m[198]&m[199])|(m[13]&m[196]&~m[197]&m[198]&m[199])|(m[13]&~m[196]&m[197]&m[198]&m[199])|(~m[13]&m[196]&m[197]&m[198]&m[199])|(m[13]&m[196]&m[197]&m[198]&m[199]))):InitCond[234];
    m[48] = run?((((m[14]&m[202]&~m[203]&~m[204]&~m[205])|(m[14]&~m[202]&m[203]&~m[204]&~m[205])|(~m[14]&m[202]&m[203]&~m[204]&~m[205])|(m[14]&~m[202]&~m[203]&m[204]&~m[205])|(~m[14]&m[202]&~m[203]&m[204]&~m[205])|(~m[14]&~m[202]&m[203]&m[204]&~m[205])|(m[14]&~m[202]&~m[203]&~m[204]&m[205])|(~m[14]&m[202]&~m[203]&~m[204]&m[205])|(~m[14]&~m[202]&m[203]&~m[204]&m[205])|(~m[14]&~m[202]&~m[203]&m[204]&m[205]))&BiasedRNG[127])|(((m[14]&m[202]&m[203]&~m[204]&~m[205])|(m[14]&m[202]&~m[203]&m[204]&~m[205])|(m[14]&~m[202]&m[203]&m[204]&~m[205])|(~m[14]&m[202]&m[203]&m[204]&~m[205])|(m[14]&m[202]&~m[203]&~m[204]&m[205])|(m[14]&~m[202]&m[203]&~m[204]&m[205])|(~m[14]&m[202]&m[203]&~m[204]&m[205])|(m[14]&~m[202]&~m[203]&m[204]&m[205])|(~m[14]&m[202]&~m[203]&m[204]&m[205])|(~m[14]&~m[202]&m[203]&m[204]&m[205]))&~BiasedRNG[127])|((m[14]&m[202]&m[203]&m[204]&~m[205])|(m[14]&m[202]&m[203]&~m[204]&m[205])|(m[14]&m[202]&~m[203]&m[204]&m[205])|(m[14]&~m[202]&m[203]&m[204]&m[205])|(~m[14]&m[202]&m[203]&m[204]&m[205])|(m[14]&m[202]&m[203]&m[204]&m[205]))):InitCond[235];
    m[49] = run?((((m[14]&m[206]&~m[207]&~m[208]&~m[209])|(m[14]&~m[206]&m[207]&~m[208]&~m[209])|(~m[14]&m[206]&m[207]&~m[208]&~m[209])|(m[14]&~m[206]&~m[207]&m[208]&~m[209])|(~m[14]&m[206]&~m[207]&m[208]&~m[209])|(~m[14]&~m[206]&m[207]&m[208]&~m[209])|(m[14]&~m[206]&~m[207]&~m[208]&m[209])|(~m[14]&m[206]&~m[207]&~m[208]&m[209])|(~m[14]&~m[206]&m[207]&~m[208]&m[209])|(~m[14]&~m[206]&~m[207]&m[208]&m[209]))&BiasedRNG[128])|(((m[14]&m[206]&m[207]&~m[208]&~m[209])|(m[14]&m[206]&~m[207]&m[208]&~m[209])|(m[14]&~m[206]&m[207]&m[208]&~m[209])|(~m[14]&m[206]&m[207]&m[208]&~m[209])|(m[14]&m[206]&~m[207]&~m[208]&m[209])|(m[14]&~m[206]&m[207]&~m[208]&m[209])|(~m[14]&m[206]&m[207]&~m[208]&m[209])|(m[14]&~m[206]&~m[207]&m[208]&m[209])|(~m[14]&m[206]&~m[207]&m[208]&m[209])|(~m[14]&~m[206]&m[207]&m[208]&m[209]))&~BiasedRNG[128])|((m[14]&m[206]&m[207]&m[208]&~m[209])|(m[14]&m[206]&m[207]&~m[208]&m[209])|(m[14]&m[206]&~m[207]&m[208]&m[209])|(m[14]&~m[206]&m[207]&m[208]&m[209])|(~m[14]&m[206]&m[207]&m[208]&m[209])|(m[14]&m[206]&m[207]&m[208]&m[209]))):InitCond[236];
    m[50] = run?((((m[15]&m[212]&~m[213]&~m[214]&~m[215])|(m[15]&~m[212]&m[213]&~m[214]&~m[215])|(~m[15]&m[212]&m[213]&~m[214]&~m[215])|(m[15]&~m[212]&~m[213]&m[214]&~m[215])|(~m[15]&m[212]&~m[213]&m[214]&~m[215])|(~m[15]&~m[212]&m[213]&m[214]&~m[215])|(m[15]&~m[212]&~m[213]&~m[214]&m[215])|(~m[15]&m[212]&~m[213]&~m[214]&m[215])|(~m[15]&~m[212]&m[213]&~m[214]&m[215])|(~m[15]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[129])|(((m[15]&m[212]&m[213]&~m[214]&~m[215])|(m[15]&m[212]&~m[213]&m[214]&~m[215])|(m[15]&~m[212]&m[213]&m[214]&~m[215])|(~m[15]&m[212]&m[213]&m[214]&~m[215])|(m[15]&m[212]&~m[213]&~m[214]&m[215])|(m[15]&~m[212]&m[213]&~m[214]&m[215])|(~m[15]&m[212]&m[213]&~m[214]&m[215])|(m[15]&~m[212]&~m[213]&m[214]&m[215])|(~m[15]&m[212]&~m[213]&m[214]&m[215])|(~m[15]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[129])|((m[15]&m[212]&m[213]&m[214]&~m[215])|(m[15]&m[212]&m[213]&~m[214]&m[215])|(m[15]&m[212]&~m[213]&m[214]&m[215])|(m[15]&~m[212]&m[213]&m[214]&m[215])|(~m[15]&m[212]&m[213]&m[214]&m[215])|(m[15]&m[212]&m[213]&m[214]&m[215]))):InitCond[237];
    m[51] = run?((((m[15]&m[216]&~m[217]&~m[218]&~m[219])|(m[15]&~m[216]&m[217]&~m[218]&~m[219])|(~m[15]&m[216]&m[217]&~m[218]&~m[219])|(m[15]&~m[216]&~m[217]&m[218]&~m[219])|(~m[15]&m[216]&~m[217]&m[218]&~m[219])|(~m[15]&~m[216]&m[217]&m[218]&~m[219])|(m[15]&~m[216]&~m[217]&~m[218]&m[219])|(~m[15]&m[216]&~m[217]&~m[218]&m[219])|(~m[15]&~m[216]&m[217]&~m[218]&m[219])|(~m[15]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[130])|(((m[15]&m[216]&m[217]&~m[218]&~m[219])|(m[15]&m[216]&~m[217]&m[218]&~m[219])|(m[15]&~m[216]&m[217]&m[218]&~m[219])|(~m[15]&m[216]&m[217]&m[218]&~m[219])|(m[15]&m[216]&~m[217]&~m[218]&m[219])|(m[15]&~m[216]&m[217]&~m[218]&m[219])|(~m[15]&m[216]&m[217]&~m[218]&m[219])|(m[15]&~m[216]&~m[217]&m[218]&m[219])|(~m[15]&m[216]&~m[217]&m[218]&m[219])|(~m[15]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[130])|((m[15]&m[216]&m[217]&m[218]&~m[219])|(m[15]&m[216]&m[217]&~m[218]&m[219])|(m[15]&m[216]&~m[217]&m[218]&m[219])|(m[15]&~m[216]&m[217]&m[218]&m[219])|(~m[15]&m[216]&m[217]&m[218]&m[219])|(m[15]&m[216]&m[217]&m[218]&m[219]))):InitCond[238];
    m[52] = run?((((m[16]&m[222]&~m[223]&~m[224]&~m[225])|(m[16]&~m[222]&m[223]&~m[224]&~m[225])|(~m[16]&m[222]&m[223]&~m[224]&~m[225])|(m[16]&~m[222]&~m[223]&m[224]&~m[225])|(~m[16]&m[222]&~m[223]&m[224]&~m[225])|(~m[16]&~m[222]&m[223]&m[224]&~m[225])|(m[16]&~m[222]&~m[223]&~m[224]&m[225])|(~m[16]&m[222]&~m[223]&~m[224]&m[225])|(~m[16]&~m[222]&m[223]&~m[224]&m[225])|(~m[16]&~m[222]&~m[223]&m[224]&m[225]))&BiasedRNG[131])|(((m[16]&m[222]&m[223]&~m[224]&~m[225])|(m[16]&m[222]&~m[223]&m[224]&~m[225])|(m[16]&~m[222]&m[223]&m[224]&~m[225])|(~m[16]&m[222]&m[223]&m[224]&~m[225])|(m[16]&m[222]&~m[223]&~m[224]&m[225])|(m[16]&~m[222]&m[223]&~m[224]&m[225])|(~m[16]&m[222]&m[223]&~m[224]&m[225])|(m[16]&~m[222]&~m[223]&m[224]&m[225])|(~m[16]&m[222]&~m[223]&m[224]&m[225])|(~m[16]&~m[222]&m[223]&m[224]&m[225]))&~BiasedRNG[131])|((m[16]&m[222]&m[223]&m[224]&~m[225])|(m[16]&m[222]&m[223]&~m[224]&m[225])|(m[16]&m[222]&~m[223]&m[224]&m[225])|(m[16]&~m[222]&m[223]&m[224]&m[225])|(~m[16]&m[222]&m[223]&m[224]&m[225])|(m[16]&m[222]&m[223]&m[224]&m[225]))):InitCond[239];
    m[53] = run?((((m[16]&m[226]&~m[227]&~m[228]&~m[229])|(m[16]&~m[226]&m[227]&~m[228]&~m[229])|(~m[16]&m[226]&m[227]&~m[228]&~m[229])|(m[16]&~m[226]&~m[227]&m[228]&~m[229])|(~m[16]&m[226]&~m[227]&m[228]&~m[229])|(~m[16]&~m[226]&m[227]&m[228]&~m[229])|(m[16]&~m[226]&~m[227]&~m[228]&m[229])|(~m[16]&m[226]&~m[227]&~m[228]&m[229])|(~m[16]&~m[226]&m[227]&~m[228]&m[229])|(~m[16]&~m[226]&~m[227]&m[228]&m[229]))&BiasedRNG[132])|(((m[16]&m[226]&m[227]&~m[228]&~m[229])|(m[16]&m[226]&~m[227]&m[228]&~m[229])|(m[16]&~m[226]&m[227]&m[228]&~m[229])|(~m[16]&m[226]&m[227]&m[228]&~m[229])|(m[16]&m[226]&~m[227]&~m[228]&m[229])|(m[16]&~m[226]&m[227]&~m[228]&m[229])|(~m[16]&m[226]&m[227]&~m[228]&m[229])|(m[16]&~m[226]&~m[227]&m[228]&m[229])|(~m[16]&m[226]&~m[227]&m[228]&m[229])|(~m[16]&~m[226]&m[227]&m[228]&m[229]))&~BiasedRNG[132])|((m[16]&m[226]&m[227]&m[228]&~m[229])|(m[16]&m[226]&m[227]&~m[228]&m[229])|(m[16]&m[226]&~m[227]&m[228]&m[229])|(m[16]&~m[226]&m[227]&m[228]&m[229])|(~m[16]&m[226]&m[227]&m[228]&m[229])|(m[16]&m[226]&m[227]&m[228]&m[229]))):InitCond[240];
    m[54] = run?((((m[17]&m[232]&~m[233]&~m[234]&~m[235])|(m[17]&~m[232]&m[233]&~m[234]&~m[235])|(~m[17]&m[232]&m[233]&~m[234]&~m[235])|(m[17]&~m[232]&~m[233]&m[234]&~m[235])|(~m[17]&m[232]&~m[233]&m[234]&~m[235])|(~m[17]&~m[232]&m[233]&m[234]&~m[235])|(m[17]&~m[232]&~m[233]&~m[234]&m[235])|(~m[17]&m[232]&~m[233]&~m[234]&m[235])|(~m[17]&~m[232]&m[233]&~m[234]&m[235])|(~m[17]&~m[232]&~m[233]&m[234]&m[235]))&BiasedRNG[133])|(((m[17]&m[232]&m[233]&~m[234]&~m[235])|(m[17]&m[232]&~m[233]&m[234]&~m[235])|(m[17]&~m[232]&m[233]&m[234]&~m[235])|(~m[17]&m[232]&m[233]&m[234]&~m[235])|(m[17]&m[232]&~m[233]&~m[234]&m[235])|(m[17]&~m[232]&m[233]&~m[234]&m[235])|(~m[17]&m[232]&m[233]&~m[234]&m[235])|(m[17]&~m[232]&~m[233]&m[234]&m[235])|(~m[17]&m[232]&~m[233]&m[234]&m[235])|(~m[17]&~m[232]&m[233]&m[234]&m[235]))&~BiasedRNG[133])|((m[17]&m[232]&m[233]&m[234]&~m[235])|(m[17]&m[232]&m[233]&~m[234]&m[235])|(m[17]&m[232]&~m[233]&m[234]&m[235])|(m[17]&~m[232]&m[233]&m[234]&m[235])|(~m[17]&m[232]&m[233]&m[234]&m[235])|(m[17]&m[232]&m[233]&m[234]&m[235]))):InitCond[241];
    m[55] = run?((((m[17]&m[236]&~m[237]&~m[238]&~m[239])|(m[17]&~m[236]&m[237]&~m[238]&~m[239])|(~m[17]&m[236]&m[237]&~m[238]&~m[239])|(m[17]&~m[236]&~m[237]&m[238]&~m[239])|(~m[17]&m[236]&~m[237]&m[238]&~m[239])|(~m[17]&~m[236]&m[237]&m[238]&~m[239])|(m[17]&~m[236]&~m[237]&~m[238]&m[239])|(~m[17]&m[236]&~m[237]&~m[238]&m[239])|(~m[17]&~m[236]&m[237]&~m[238]&m[239])|(~m[17]&~m[236]&~m[237]&m[238]&m[239]))&BiasedRNG[134])|(((m[17]&m[236]&m[237]&~m[238]&~m[239])|(m[17]&m[236]&~m[237]&m[238]&~m[239])|(m[17]&~m[236]&m[237]&m[238]&~m[239])|(~m[17]&m[236]&m[237]&m[238]&~m[239])|(m[17]&m[236]&~m[237]&~m[238]&m[239])|(m[17]&~m[236]&m[237]&~m[238]&m[239])|(~m[17]&m[236]&m[237]&~m[238]&m[239])|(m[17]&~m[236]&~m[237]&m[238]&m[239])|(~m[17]&m[236]&~m[237]&m[238]&m[239])|(~m[17]&~m[236]&m[237]&m[238]&m[239]))&~BiasedRNG[134])|((m[17]&m[236]&m[237]&m[238]&~m[239])|(m[17]&m[236]&m[237]&~m[238]&m[239])|(m[17]&m[236]&~m[237]&m[238]&m[239])|(m[17]&~m[236]&m[237]&m[238]&m[239])|(~m[17]&m[236]&m[237]&m[238]&m[239])|(m[17]&m[236]&m[237]&m[238]&m[239]))):InitCond[242];
    m[56] = run?((((m[18]&m[242]&~m[243]&~m[244]&~m[245])|(m[18]&~m[242]&m[243]&~m[244]&~m[245])|(~m[18]&m[242]&m[243]&~m[244]&~m[245])|(m[18]&~m[242]&~m[243]&m[244]&~m[245])|(~m[18]&m[242]&~m[243]&m[244]&~m[245])|(~m[18]&~m[242]&m[243]&m[244]&~m[245])|(m[18]&~m[242]&~m[243]&~m[244]&m[245])|(~m[18]&m[242]&~m[243]&~m[244]&m[245])|(~m[18]&~m[242]&m[243]&~m[244]&m[245])|(~m[18]&~m[242]&~m[243]&m[244]&m[245]))&BiasedRNG[135])|(((m[18]&m[242]&m[243]&~m[244]&~m[245])|(m[18]&m[242]&~m[243]&m[244]&~m[245])|(m[18]&~m[242]&m[243]&m[244]&~m[245])|(~m[18]&m[242]&m[243]&m[244]&~m[245])|(m[18]&m[242]&~m[243]&~m[244]&m[245])|(m[18]&~m[242]&m[243]&~m[244]&m[245])|(~m[18]&m[242]&m[243]&~m[244]&m[245])|(m[18]&~m[242]&~m[243]&m[244]&m[245])|(~m[18]&m[242]&~m[243]&m[244]&m[245])|(~m[18]&~m[242]&m[243]&m[244]&m[245]))&~BiasedRNG[135])|((m[18]&m[242]&m[243]&m[244]&~m[245])|(m[18]&m[242]&m[243]&~m[244]&m[245])|(m[18]&m[242]&~m[243]&m[244]&m[245])|(m[18]&~m[242]&m[243]&m[244]&m[245])|(~m[18]&m[242]&m[243]&m[244]&m[245])|(m[18]&m[242]&m[243]&m[244]&m[245]))):InitCond[243];
    m[57] = run?((((m[18]&m[246]&~m[247]&~m[248]&~m[249])|(m[18]&~m[246]&m[247]&~m[248]&~m[249])|(~m[18]&m[246]&m[247]&~m[248]&~m[249])|(m[18]&~m[246]&~m[247]&m[248]&~m[249])|(~m[18]&m[246]&~m[247]&m[248]&~m[249])|(~m[18]&~m[246]&m[247]&m[248]&~m[249])|(m[18]&~m[246]&~m[247]&~m[248]&m[249])|(~m[18]&m[246]&~m[247]&~m[248]&m[249])|(~m[18]&~m[246]&m[247]&~m[248]&m[249])|(~m[18]&~m[246]&~m[247]&m[248]&m[249]))&BiasedRNG[136])|(((m[18]&m[246]&m[247]&~m[248]&~m[249])|(m[18]&m[246]&~m[247]&m[248]&~m[249])|(m[18]&~m[246]&m[247]&m[248]&~m[249])|(~m[18]&m[246]&m[247]&m[248]&~m[249])|(m[18]&m[246]&~m[247]&~m[248]&m[249])|(m[18]&~m[246]&m[247]&~m[248]&m[249])|(~m[18]&m[246]&m[247]&~m[248]&m[249])|(m[18]&~m[246]&~m[247]&m[248]&m[249])|(~m[18]&m[246]&~m[247]&m[248]&m[249])|(~m[18]&~m[246]&m[247]&m[248]&m[249]))&~BiasedRNG[136])|((m[18]&m[246]&m[247]&m[248]&~m[249])|(m[18]&m[246]&m[247]&~m[248]&m[249])|(m[18]&m[246]&~m[247]&m[248]&m[249])|(m[18]&~m[246]&m[247]&m[248]&m[249])|(~m[18]&m[246]&m[247]&m[248]&m[249])|(m[18]&m[246]&m[247]&m[248]&m[249]))):InitCond[244];
    m[58] = run?((((m[19]&m[252]&~m[253]&~m[254]&~m[255])|(m[19]&~m[252]&m[253]&~m[254]&~m[255])|(~m[19]&m[252]&m[253]&~m[254]&~m[255])|(m[19]&~m[252]&~m[253]&m[254]&~m[255])|(~m[19]&m[252]&~m[253]&m[254]&~m[255])|(~m[19]&~m[252]&m[253]&m[254]&~m[255])|(m[19]&~m[252]&~m[253]&~m[254]&m[255])|(~m[19]&m[252]&~m[253]&~m[254]&m[255])|(~m[19]&~m[252]&m[253]&~m[254]&m[255])|(~m[19]&~m[252]&~m[253]&m[254]&m[255]))&BiasedRNG[137])|(((m[19]&m[252]&m[253]&~m[254]&~m[255])|(m[19]&m[252]&~m[253]&m[254]&~m[255])|(m[19]&~m[252]&m[253]&m[254]&~m[255])|(~m[19]&m[252]&m[253]&m[254]&~m[255])|(m[19]&m[252]&~m[253]&~m[254]&m[255])|(m[19]&~m[252]&m[253]&~m[254]&m[255])|(~m[19]&m[252]&m[253]&~m[254]&m[255])|(m[19]&~m[252]&~m[253]&m[254]&m[255])|(~m[19]&m[252]&~m[253]&m[254]&m[255])|(~m[19]&~m[252]&m[253]&m[254]&m[255]))&~BiasedRNG[137])|((m[19]&m[252]&m[253]&m[254]&~m[255])|(m[19]&m[252]&m[253]&~m[254]&m[255])|(m[19]&m[252]&~m[253]&m[254]&m[255])|(m[19]&~m[252]&m[253]&m[254]&m[255])|(~m[19]&m[252]&m[253]&m[254]&m[255])|(m[19]&m[252]&m[253]&m[254]&m[255]))):InitCond[245];
    m[59] = run?((((m[19]&m[256]&~m[257]&~m[258]&~m[259])|(m[19]&~m[256]&m[257]&~m[258]&~m[259])|(~m[19]&m[256]&m[257]&~m[258]&~m[259])|(m[19]&~m[256]&~m[257]&m[258]&~m[259])|(~m[19]&m[256]&~m[257]&m[258]&~m[259])|(~m[19]&~m[256]&m[257]&m[258]&~m[259])|(m[19]&~m[256]&~m[257]&~m[258]&m[259])|(~m[19]&m[256]&~m[257]&~m[258]&m[259])|(~m[19]&~m[256]&m[257]&~m[258]&m[259])|(~m[19]&~m[256]&~m[257]&m[258]&m[259]))&BiasedRNG[138])|(((m[19]&m[256]&m[257]&~m[258]&~m[259])|(m[19]&m[256]&~m[257]&m[258]&~m[259])|(m[19]&~m[256]&m[257]&m[258]&~m[259])|(~m[19]&m[256]&m[257]&m[258]&~m[259])|(m[19]&m[256]&~m[257]&~m[258]&m[259])|(m[19]&~m[256]&m[257]&~m[258]&m[259])|(~m[19]&m[256]&m[257]&~m[258]&m[259])|(m[19]&~m[256]&~m[257]&m[258]&m[259])|(~m[19]&m[256]&~m[257]&m[258]&m[259])|(~m[19]&~m[256]&m[257]&m[258]&m[259]))&~BiasedRNG[138])|((m[19]&m[256]&m[257]&m[258]&~m[259])|(m[19]&m[256]&m[257]&~m[258]&m[259])|(m[19]&m[256]&~m[257]&m[258]&m[259])|(m[19]&~m[256]&m[257]&m[258]&m[259])|(~m[19]&m[256]&m[257]&m[258]&m[259])|(m[19]&m[256]&m[257]&m[258]&m[259]))):InitCond[246];
    m[60] = run?((((~m[0]&~m[160]&~m[260])|(m[0]&m[160]&~m[260]))&BiasedRNG[139])|(((m[0]&~m[160]&~m[260])|(~m[0]&m[160]&m[260]))&~BiasedRNG[139])|((~m[0]&~m[160]&m[260])|(m[0]&~m[160]&m[260])|(m[0]&m[160]&m[260]))):InitCond[247];
    m[61] = run?((((~m[0]&~m[170]&~m[270])|(m[0]&m[170]&~m[270]))&BiasedRNG[140])|(((m[0]&~m[170]&~m[270])|(~m[0]&m[170]&m[270]))&~BiasedRNG[140])|((~m[0]&~m[170]&m[270])|(m[0]&~m[170]&m[270])|(m[0]&m[170]&m[270]))):InitCond[248];
    m[70] = run?((((~m[1]&~m[161]&~m[261])|(m[1]&m[161]&~m[261]))&BiasedRNG[141])|(((m[1]&~m[161]&~m[261])|(~m[1]&m[161]&m[261]))&~BiasedRNG[141])|((~m[1]&~m[161]&m[261])|(m[1]&~m[161]&m[261])|(m[1]&m[161]&m[261]))):InitCond[249];
    m[71] = run?((((~m[1]&~m[171]&~m[271])|(m[1]&m[171]&~m[271]))&BiasedRNG[142])|(((m[1]&~m[171]&~m[271])|(~m[1]&m[171]&m[271]))&~BiasedRNG[142])|((~m[1]&~m[171]&m[271])|(m[1]&~m[171]&m[271])|(m[1]&m[171]&m[271]))):InitCond[250];
    m[80] = run?((((~m[2]&~m[162]&~m[262])|(m[2]&m[162]&~m[262]))&BiasedRNG[143])|(((m[2]&~m[162]&~m[262])|(~m[2]&m[162]&m[262]))&~BiasedRNG[143])|((~m[2]&~m[162]&m[262])|(m[2]&~m[162]&m[262])|(m[2]&m[162]&m[262]))):InitCond[251];
    m[81] = run?((((~m[2]&~m[172]&~m[272])|(m[2]&m[172]&~m[272]))&BiasedRNG[144])|(((m[2]&~m[172]&~m[272])|(~m[2]&m[172]&m[272]))&~BiasedRNG[144])|((~m[2]&~m[172]&m[272])|(m[2]&~m[172]&m[272])|(m[2]&m[172]&m[272]))):InitCond[252];
    m[90] = run?((((~m[3]&~m[163]&~m[263])|(m[3]&m[163]&~m[263]))&BiasedRNG[145])|(((m[3]&~m[163]&~m[263])|(~m[3]&m[163]&m[263]))&~BiasedRNG[145])|((~m[3]&~m[163]&m[263])|(m[3]&~m[163]&m[263])|(m[3]&m[163]&m[263]))):InitCond[253];
    m[91] = run?((((~m[3]&~m[173]&~m[273])|(m[3]&m[173]&~m[273]))&BiasedRNG[146])|(((m[3]&~m[173]&~m[273])|(~m[3]&m[173]&m[273]))&~BiasedRNG[146])|((~m[3]&~m[173]&m[273])|(m[3]&~m[173]&m[273])|(m[3]&m[173]&m[273]))):InitCond[254];
    m[100] = run?((((~m[4]&~m[164]&~m[264])|(m[4]&m[164]&~m[264]))&BiasedRNG[147])|(((m[4]&~m[164]&~m[264])|(~m[4]&m[164]&m[264]))&~BiasedRNG[147])|((~m[4]&~m[164]&m[264])|(m[4]&~m[164]&m[264])|(m[4]&m[164]&m[264]))):InitCond[255];
    m[101] = run?((((~m[4]&~m[174]&~m[274])|(m[4]&m[174]&~m[274]))&BiasedRNG[148])|(((m[4]&~m[174]&~m[274])|(~m[4]&m[174]&m[274]))&~BiasedRNG[148])|((~m[4]&~m[174]&m[274])|(m[4]&~m[174]&m[274])|(m[4]&m[174]&m[274]))):InitCond[256];
    m[110] = run?((((~m[5]&~m[165]&~m[265])|(m[5]&m[165]&~m[265]))&BiasedRNG[149])|(((m[5]&~m[165]&~m[265])|(~m[5]&m[165]&m[265]))&~BiasedRNG[149])|((~m[5]&~m[165]&m[265])|(m[5]&~m[165]&m[265])|(m[5]&m[165]&m[265]))):InitCond[257];
    m[111] = run?((((~m[5]&~m[175]&~m[275])|(m[5]&m[175]&~m[275]))&BiasedRNG[150])|(((m[5]&~m[175]&~m[275])|(~m[5]&m[175]&m[275]))&~BiasedRNG[150])|((~m[5]&~m[175]&m[275])|(m[5]&~m[175]&m[275])|(m[5]&m[175]&m[275]))):InitCond[258];
    m[120] = run?((((~m[6]&~m[166]&~m[266])|(m[6]&m[166]&~m[266]))&BiasedRNG[151])|(((m[6]&~m[166]&~m[266])|(~m[6]&m[166]&m[266]))&~BiasedRNG[151])|((~m[6]&~m[166]&m[266])|(m[6]&~m[166]&m[266])|(m[6]&m[166]&m[266]))):InitCond[259];
    m[121] = run?((((~m[6]&~m[176]&~m[276])|(m[6]&m[176]&~m[276]))&BiasedRNG[152])|(((m[6]&~m[176]&~m[276])|(~m[6]&m[176]&m[276]))&~BiasedRNG[152])|((~m[6]&~m[176]&m[276])|(m[6]&~m[176]&m[276])|(m[6]&m[176]&m[276]))):InitCond[260];
    m[130] = run?((((~m[7]&~m[167]&~m[267])|(m[7]&m[167]&~m[267]))&BiasedRNG[153])|(((m[7]&~m[167]&~m[267])|(~m[7]&m[167]&m[267]))&~BiasedRNG[153])|((~m[7]&~m[167]&m[267])|(m[7]&~m[167]&m[267])|(m[7]&m[167]&m[267]))):InitCond[261];
    m[131] = run?((((~m[7]&~m[177]&~m[277])|(m[7]&m[177]&~m[277]))&BiasedRNG[154])|(((m[7]&~m[177]&~m[277])|(~m[7]&m[177]&m[277]))&~BiasedRNG[154])|((~m[7]&~m[177]&m[277])|(m[7]&~m[177]&m[277])|(m[7]&m[177]&m[277]))):InitCond[262];
    m[140] = run?((((~m[8]&~m[168]&~m[268])|(m[8]&m[168]&~m[268]))&BiasedRNG[155])|(((m[8]&~m[168]&~m[268])|(~m[8]&m[168]&m[268]))&~BiasedRNG[155])|((~m[8]&~m[168]&m[268])|(m[8]&~m[168]&m[268])|(m[8]&m[168]&m[268]))):InitCond[263];
    m[141] = run?((((~m[8]&~m[178]&~m[278])|(m[8]&m[178]&~m[278]))&BiasedRNG[156])|(((m[8]&~m[178]&~m[278])|(~m[8]&m[178]&m[278]))&~BiasedRNG[156])|((~m[8]&~m[178]&m[278])|(m[8]&~m[178]&m[278])|(m[8]&m[178]&m[278]))):InitCond[264];
    m[150] = run?((((~m[9]&~m[169]&~m[269])|(m[9]&m[169]&~m[269]))&BiasedRNG[157])|(((m[9]&~m[169]&~m[269])|(~m[9]&m[169]&m[269]))&~BiasedRNG[157])|((~m[9]&~m[169]&m[269])|(m[9]&~m[169]&m[269])|(m[9]&m[169]&m[269]))):InitCond[265];
    m[151] = run?((((~m[9]&~m[179]&~m[279])|(m[9]&m[179]&~m[279]))&BiasedRNG[158])|(((m[9]&~m[179]&~m[279])|(~m[9]&m[179]&m[279]))&~BiasedRNG[158])|((~m[9]&~m[179]&m[279])|(m[9]&~m[179]&m[279])|(m[9]&m[179]&m[279]))):InitCond[266];
    m[180] = run?((((~m[12]&~m[62]&~m[280])|(m[12]&m[62]&~m[280]))&BiasedRNG[159])|(((m[12]&~m[62]&~m[280])|(~m[12]&m[62]&m[280]))&~BiasedRNG[159])|((~m[12]&~m[62]&m[280])|(m[12]&~m[62]&m[280])|(m[12]&m[62]&m[280]))):InitCond[267];
    m[181] = run?((((~m[12]&~m[72]&~m[281])|(m[12]&m[72]&~m[281]))&BiasedRNG[160])|(((m[12]&~m[72]&~m[281])|(~m[12]&m[72]&m[281]))&~BiasedRNG[160])|((~m[12]&~m[72]&m[281])|(m[12]&~m[72]&m[281])|(m[12]&m[72]&m[281]))):InitCond[268];
    m[190] = run?((((~m[13]&~m[63]&~m[290])|(m[13]&m[63]&~m[290]))&BiasedRNG[161])|(((m[13]&~m[63]&~m[290])|(~m[13]&m[63]&m[290]))&~BiasedRNG[161])|((~m[13]&~m[63]&m[290])|(m[13]&~m[63]&m[290])|(m[13]&m[63]&m[290]))):InitCond[269];
    m[191] = run?((((~m[13]&~m[73]&~m[291])|(m[13]&m[73]&~m[291]))&BiasedRNG[162])|(((m[13]&~m[73]&~m[291])|(~m[13]&m[73]&m[291]))&~BiasedRNG[162])|((~m[13]&~m[73]&m[291])|(m[13]&~m[73]&m[291])|(m[13]&m[73]&m[291]))):InitCond[270];
    m[200] = run?((((~m[14]&~m[64]&~m[300])|(m[14]&m[64]&~m[300]))&BiasedRNG[163])|(((m[14]&~m[64]&~m[300])|(~m[14]&m[64]&m[300]))&~BiasedRNG[163])|((~m[14]&~m[64]&m[300])|(m[14]&~m[64]&m[300])|(m[14]&m[64]&m[300]))):InitCond[271];
    m[201] = run?((((~m[14]&~m[74]&~m[301])|(m[14]&m[74]&~m[301]))&BiasedRNG[164])|(((m[14]&~m[74]&~m[301])|(~m[14]&m[74]&m[301]))&~BiasedRNG[164])|((~m[14]&~m[74]&m[301])|(m[14]&~m[74]&m[301])|(m[14]&m[74]&m[301]))):InitCond[272];
    m[210] = run?((((~m[15]&~m[65]&~m[310])|(m[15]&m[65]&~m[310]))&BiasedRNG[165])|(((m[15]&~m[65]&~m[310])|(~m[15]&m[65]&m[310]))&~BiasedRNG[165])|((~m[15]&~m[65]&m[310])|(m[15]&~m[65]&m[310])|(m[15]&m[65]&m[310]))):InitCond[273];
    m[211] = run?((((~m[15]&~m[75]&~m[311])|(m[15]&m[75]&~m[311]))&BiasedRNG[166])|(((m[15]&~m[75]&~m[311])|(~m[15]&m[75]&m[311]))&~BiasedRNG[166])|((~m[15]&~m[75]&m[311])|(m[15]&~m[75]&m[311])|(m[15]&m[75]&m[311]))):InitCond[274];
    m[220] = run?((((~m[16]&~m[66]&~m[320])|(m[16]&m[66]&~m[320]))&BiasedRNG[167])|(((m[16]&~m[66]&~m[320])|(~m[16]&m[66]&m[320]))&~BiasedRNG[167])|((~m[16]&~m[66]&m[320])|(m[16]&~m[66]&m[320])|(m[16]&m[66]&m[320]))):InitCond[275];
    m[221] = run?((((~m[16]&~m[76]&~m[321])|(m[16]&m[76]&~m[321]))&BiasedRNG[168])|(((m[16]&~m[76]&~m[321])|(~m[16]&m[76]&m[321]))&~BiasedRNG[168])|((~m[16]&~m[76]&m[321])|(m[16]&~m[76]&m[321])|(m[16]&m[76]&m[321]))):InitCond[276];
    m[230] = run?((((~m[17]&~m[67]&~m[330])|(m[17]&m[67]&~m[330]))&BiasedRNG[169])|(((m[17]&~m[67]&~m[330])|(~m[17]&m[67]&m[330]))&~BiasedRNG[169])|((~m[17]&~m[67]&m[330])|(m[17]&~m[67]&m[330])|(m[17]&m[67]&m[330]))):InitCond[277];
    m[231] = run?((((~m[17]&~m[77]&~m[331])|(m[17]&m[77]&~m[331]))&BiasedRNG[170])|(((m[17]&~m[77]&~m[331])|(~m[17]&m[77]&m[331]))&~BiasedRNG[170])|((~m[17]&~m[77]&m[331])|(m[17]&~m[77]&m[331])|(m[17]&m[77]&m[331]))):InitCond[278];
    m[240] = run?((((~m[18]&~m[68]&~m[340])|(m[18]&m[68]&~m[340]))&BiasedRNG[171])|(((m[18]&~m[68]&~m[340])|(~m[18]&m[68]&m[340]))&~BiasedRNG[171])|((~m[18]&~m[68]&m[340])|(m[18]&~m[68]&m[340])|(m[18]&m[68]&m[340]))):InitCond[279];
    m[241] = run?((((~m[18]&~m[78]&~m[341])|(m[18]&m[78]&~m[341]))&BiasedRNG[172])|(((m[18]&~m[78]&~m[341])|(~m[18]&m[78]&m[341]))&~BiasedRNG[172])|((~m[18]&~m[78]&m[341])|(m[18]&~m[78]&m[341])|(m[18]&m[78]&m[341]))):InitCond[280];
    m[250] = run?((((~m[19]&~m[69]&~m[350])|(m[19]&m[69]&~m[350]))&BiasedRNG[173])|(((m[19]&~m[69]&~m[350])|(~m[19]&m[69]&m[350]))&~BiasedRNG[173])|((~m[19]&~m[69]&m[350])|(m[19]&~m[69]&m[350])|(m[19]&m[69]&m[350]))):InitCond[281];
    m[251] = run?((((~m[19]&~m[79]&~m[351])|(m[19]&m[79]&~m[351]))&BiasedRNG[174])|(((m[19]&~m[79]&~m[351])|(~m[19]&m[79]&m[351]))&~BiasedRNG[174])|((~m[19]&~m[79]&m[351])|(m[19]&~m[79]&m[351])|(m[19]&m[79]&m[351]))):InitCond[282];
    m[282] = run?((((m[82]&~m[182]&m[396])|(~m[82]&m[182]&m[396]))&BiasedRNG[175])|(((m[82]&m[182]&~m[396]))&~BiasedRNG[175])|((m[82]&m[182]&m[396]))):InitCond[283];
    m[283] = run?((((m[92]&~m[183]&m[416])|(~m[92]&m[183]&m[416]))&BiasedRNG[176])|(((m[92]&m[183]&~m[416]))&~BiasedRNG[176])|((m[92]&m[183]&m[416]))):InitCond[284];
    m[284] = run?((((m[102]&~m[184]&m[441])|(~m[102]&m[184]&m[441]))&BiasedRNG[177])|(((m[102]&m[184]&~m[441]))&~BiasedRNG[177])|((m[102]&m[184]&m[441]))):InitCond[285];
    m[285] = run?((((m[112]&~m[185]&m[471])|(~m[112]&m[185]&m[471]))&BiasedRNG[178])|(((m[112]&m[185]&~m[471]))&~BiasedRNG[178])|((m[112]&m[185]&m[471]))):InitCond[286];
    m[286] = run?((((m[122]&~m[186]&m[506])|(~m[122]&m[186]&m[506]))&BiasedRNG[179])|(((m[122]&m[186]&~m[506]))&~BiasedRNG[179])|((m[122]&m[186]&m[506]))):InitCond[287];
    m[287] = run?((((m[132]&~m[187]&m[546])|(~m[132]&m[187]&m[546]))&BiasedRNG[180])|(((m[132]&m[187]&~m[546]))&~BiasedRNG[180])|((m[132]&m[187]&m[546]))):InitCond[288];
    m[288] = run?((((m[142]&~m[188]&m[591])|(~m[142]&m[188]&m[591]))&BiasedRNG[181])|(((m[142]&m[188]&~m[591]))&~BiasedRNG[181])|((m[142]&m[188]&m[591]))):InitCond[289];
    m[289] = run?((((m[152]&~m[189]&m[631])|(~m[152]&m[189]&m[631]))&BiasedRNG[182])|(((m[152]&m[189]&~m[631]))&~BiasedRNG[182])|((m[152]&m[189]&m[631]))):InitCond[290];
    m[292] = run?((((m[83]&~m[192]&m[421])|(~m[83]&m[192]&m[421]))&BiasedRNG[183])|(((m[83]&m[192]&~m[421]))&~BiasedRNG[183])|((m[83]&m[192]&m[421]))):InitCond[291];
    m[293] = run?((((m[93]&~m[193]&m[446])|(~m[93]&m[193]&m[446]))&BiasedRNG[184])|(((m[93]&m[193]&~m[446]))&~BiasedRNG[184])|((m[93]&m[193]&m[446]))):InitCond[292];
    m[294] = run?((((m[103]&~m[194]&m[476])|(~m[103]&m[194]&m[476]))&BiasedRNG[185])|(((m[103]&m[194]&~m[476]))&~BiasedRNG[185])|((m[103]&m[194]&m[476]))):InitCond[293];
    m[295] = run?((((m[113]&~m[195]&m[511])|(~m[113]&m[195]&m[511]))&BiasedRNG[186])|(((m[113]&m[195]&~m[511]))&~BiasedRNG[186])|((m[113]&m[195]&m[511]))):InitCond[294];
    m[296] = run?((((m[123]&~m[196]&m[551])|(~m[123]&m[196]&m[551]))&BiasedRNG[187])|(((m[123]&m[196]&~m[551]))&~BiasedRNG[187])|((m[123]&m[196]&m[551]))):InitCond[295];
    m[297] = run?((((m[133]&~m[197]&m[596])|(~m[133]&m[197]&m[596]))&BiasedRNG[188])|(((m[133]&m[197]&~m[596]))&~BiasedRNG[188])|((m[133]&m[197]&m[596]))):InitCond[296];
    m[298] = run?((((m[143]&~m[198]&m[636])|(~m[143]&m[198]&m[636]))&BiasedRNG[189])|(((m[143]&m[198]&~m[636]))&~BiasedRNG[189])|((m[143]&m[198]&m[636]))):InitCond[297];
    m[299] = run?((((m[153]&~m[199]&m[671])|(~m[153]&m[199]&m[671]))&BiasedRNG[190])|(((m[153]&m[199]&~m[671]))&~BiasedRNG[190])|((m[153]&m[199]&m[671]))):InitCond[298];
    m[302] = run?((((m[84]&~m[202]&m[451])|(~m[84]&m[202]&m[451]))&BiasedRNG[191])|(((m[84]&m[202]&~m[451]))&~BiasedRNG[191])|((m[84]&m[202]&m[451]))):InitCond[299];
    m[303] = run?((((m[94]&~m[203]&m[481])|(~m[94]&m[203]&m[481]))&BiasedRNG[192])|(((m[94]&m[203]&~m[481]))&~BiasedRNG[192])|((m[94]&m[203]&m[481]))):InitCond[300];
    m[304] = run?((((m[104]&~m[204]&m[516])|(~m[104]&m[204]&m[516]))&BiasedRNG[193])|(((m[104]&m[204]&~m[516]))&~BiasedRNG[193])|((m[104]&m[204]&m[516]))):InitCond[301];
    m[305] = run?((((m[114]&~m[205]&m[556])|(~m[114]&m[205]&m[556]))&BiasedRNG[194])|(((m[114]&m[205]&~m[556]))&~BiasedRNG[194])|((m[114]&m[205]&m[556]))):InitCond[302];
    m[306] = run?((((m[124]&~m[206]&m[601])|(~m[124]&m[206]&m[601]))&BiasedRNG[195])|(((m[124]&m[206]&~m[601]))&~BiasedRNG[195])|((m[124]&m[206]&m[601]))):InitCond[303];
    m[307] = run?((((m[134]&~m[207]&m[641])|(~m[134]&m[207]&m[641]))&BiasedRNG[196])|(((m[134]&m[207]&~m[641]))&~BiasedRNG[196])|((m[134]&m[207]&m[641]))):InitCond[304];
    m[308] = run?((((m[144]&~m[208]&m[676])|(~m[144]&m[208]&m[676]))&BiasedRNG[197])|(((m[144]&m[208]&~m[676]))&~BiasedRNG[197])|((m[144]&m[208]&m[676]))):InitCond[305];
    m[309] = run?((((m[154]&~m[209]&m[706])|(~m[154]&m[209]&m[706]))&BiasedRNG[198])|(((m[154]&m[209]&~m[706]))&~BiasedRNG[198])|((m[154]&m[209]&m[706]))):InitCond[306];
    m[312] = run?((((m[85]&~m[212]&m[486])|(~m[85]&m[212]&m[486]))&BiasedRNG[199])|(((m[85]&m[212]&~m[486]))&~BiasedRNG[199])|((m[85]&m[212]&m[486]))):InitCond[307];
    m[313] = run?((((m[95]&~m[213]&m[521])|(~m[95]&m[213]&m[521]))&BiasedRNG[200])|(((m[95]&m[213]&~m[521]))&~BiasedRNG[200])|((m[95]&m[213]&m[521]))):InitCond[308];
    m[314] = run?((((m[105]&~m[214]&m[561])|(~m[105]&m[214]&m[561]))&BiasedRNG[201])|(((m[105]&m[214]&~m[561]))&~BiasedRNG[201])|((m[105]&m[214]&m[561]))):InitCond[309];
    m[315] = run?((((m[115]&~m[215]&m[606])|(~m[115]&m[215]&m[606]))&BiasedRNG[202])|(((m[115]&m[215]&~m[606]))&~BiasedRNG[202])|((m[115]&m[215]&m[606]))):InitCond[310];
    m[316] = run?((((m[125]&~m[216]&m[646])|(~m[125]&m[216]&m[646]))&BiasedRNG[203])|(((m[125]&m[216]&~m[646]))&~BiasedRNG[203])|((m[125]&m[216]&m[646]))):InitCond[311];
    m[317] = run?((((m[135]&~m[217]&m[681])|(~m[135]&m[217]&m[681]))&BiasedRNG[204])|(((m[135]&m[217]&~m[681]))&~BiasedRNG[204])|((m[135]&m[217]&m[681]))):InitCond[312];
    m[318] = run?((((m[145]&~m[218]&m[711])|(~m[145]&m[218]&m[711]))&BiasedRNG[205])|(((m[145]&m[218]&~m[711]))&~BiasedRNG[205])|((m[145]&m[218]&m[711]))):InitCond[313];
    m[319] = run?((((m[155]&~m[219]&m[736])|(~m[155]&m[219]&m[736]))&BiasedRNG[206])|(((m[155]&m[219]&~m[736]))&~BiasedRNG[206])|((m[155]&m[219]&m[736]))):InitCond[314];
    m[322] = run?((((m[86]&~m[222]&m[526])|(~m[86]&m[222]&m[526]))&BiasedRNG[207])|(((m[86]&m[222]&~m[526]))&~BiasedRNG[207])|((m[86]&m[222]&m[526]))):InitCond[315];
    m[323] = run?((((m[96]&~m[223]&m[566])|(~m[96]&m[223]&m[566]))&BiasedRNG[208])|(((m[96]&m[223]&~m[566]))&~BiasedRNG[208])|((m[96]&m[223]&m[566]))):InitCond[316];
    m[324] = run?((((m[106]&~m[224]&m[611])|(~m[106]&m[224]&m[611]))&BiasedRNG[209])|(((m[106]&m[224]&~m[611]))&~BiasedRNG[209])|((m[106]&m[224]&m[611]))):InitCond[317];
    m[325] = run?((((m[116]&~m[225]&m[651])|(~m[116]&m[225]&m[651]))&BiasedRNG[210])|(((m[116]&m[225]&~m[651]))&~BiasedRNG[210])|((m[116]&m[225]&m[651]))):InitCond[318];
    m[326] = run?((((m[126]&~m[226]&m[686])|(~m[126]&m[226]&m[686]))&BiasedRNG[211])|(((m[126]&m[226]&~m[686]))&~BiasedRNG[211])|((m[126]&m[226]&m[686]))):InitCond[319];
    m[327] = run?((((m[136]&~m[227]&m[716])|(~m[136]&m[227]&m[716]))&BiasedRNG[212])|(((m[136]&m[227]&~m[716]))&~BiasedRNG[212])|((m[136]&m[227]&m[716]))):InitCond[320];
    m[328] = run?((((m[146]&~m[228]&m[741])|(~m[146]&m[228]&m[741]))&BiasedRNG[213])|(((m[146]&m[228]&~m[741]))&~BiasedRNG[213])|((m[146]&m[228]&m[741]))):InitCond[321];
    m[329] = run?((((m[156]&~m[229]&m[761])|(~m[156]&m[229]&m[761]))&BiasedRNG[214])|(((m[156]&m[229]&~m[761]))&~BiasedRNG[214])|((m[156]&m[229]&m[761]))):InitCond[322];
    m[332] = run?((((m[87]&~m[232]&m[571])|(~m[87]&m[232]&m[571]))&BiasedRNG[215])|(((m[87]&m[232]&~m[571]))&~BiasedRNG[215])|((m[87]&m[232]&m[571]))):InitCond[323];
    m[333] = run?((((m[97]&~m[233]&m[616])|(~m[97]&m[233]&m[616]))&BiasedRNG[216])|(((m[97]&m[233]&~m[616]))&~BiasedRNG[216])|((m[97]&m[233]&m[616]))):InitCond[324];
    m[334] = run?((((m[107]&~m[234]&m[656])|(~m[107]&m[234]&m[656]))&BiasedRNG[217])|(((m[107]&m[234]&~m[656]))&~BiasedRNG[217])|((m[107]&m[234]&m[656]))):InitCond[325];
    m[335] = run?((((m[117]&~m[235]&m[691])|(~m[117]&m[235]&m[691]))&BiasedRNG[218])|(((m[117]&m[235]&~m[691]))&~BiasedRNG[218])|((m[117]&m[235]&m[691]))):InitCond[326];
    m[336] = run?((((m[127]&~m[236]&m[721])|(~m[127]&m[236]&m[721]))&BiasedRNG[219])|(((m[127]&m[236]&~m[721]))&~BiasedRNG[219])|((m[127]&m[236]&m[721]))):InitCond[327];
    m[337] = run?((((m[137]&~m[237]&m[746])|(~m[137]&m[237]&m[746]))&BiasedRNG[220])|(((m[137]&m[237]&~m[746]))&~BiasedRNG[220])|((m[137]&m[237]&m[746]))):InitCond[328];
    m[338] = run?((((m[147]&~m[238]&m[766])|(~m[147]&m[238]&m[766]))&BiasedRNG[221])|(((m[147]&m[238]&~m[766]))&~BiasedRNG[221])|((m[147]&m[238]&m[766]))):InitCond[329];
    m[339] = run?((((m[157]&~m[239]&m[781])|(~m[157]&m[239]&m[781]))&BiasedRNG[222])|(((m[157]&m[239]&~m[781]))&~BiasedRNG[222])|((m[157]&m[239]&m[781]))):InitCond[330];
    m[342] = run?((((m[88]&~m[242]&m[621])|(~m[88]&m[242]&m[621]))&BiasedRNG[223])|(((m[88]&m[242]&~m[621]))&~BiasedRNG[223])|((m[88]&m[242]&m[621]))):InitCond[331];
    m[343] = run?((((m[98]&~m[243]&m[661])|(~m[98]&m[243]&m[661]))&BiasedRNG[224])|(((m[98]&m[243]&~m[661]))&~BiasedRNG[224])|((m[98]&m[243]&m[661]))):InitCond[332];
    m[344] = run?((((m[108]&~m[244]&m[696])|(~m[108]&m[244]&m[696]))&BiasedRNG[225])|(((m[108]&m[244]&~m[696]))&~BiasedRNG[225])|((m[108]&m[244]&m[696]))):InitCond[333];
    m[345] = run?((((m[118]&~m[245]&m[726])|(~m[118]&m[245]&m[726]))&BiasedRNG[226])|(((m[118]&m[245]&~m[726]))&~BiasedRNG[226])|((m[118]&m[245]&m[726]))):InitCond[334];
    m[346] = run?((((m[128]&~m[246]&m[751])|(~m[128]&m[246]&m[751]))&BiasedRNG[227])|(((m[128]&m[246]&~m[751]))&~BiasedRNG[227])|((m[128]&m[246]&m[751]))):InitCond[335];
    m[347] = run?((((m[138]&~m[247]&m[771])|(~m[138]&m[247]&m[771]))&BiasedRNG[228])|(((m[138]&m[247]&~m[771]))&~BiasedRNG[228])|((m[138]&m[247]&m[771]))):InitCond[336];
    m[348] = run?((((m[148]&~m[248]&m[786])|(~m[148]&m[248]&m[786]))&BiasedRNG[229])|(((m[148]&m[248]&~m[786]))&~BiasedRNG[229])|((m[148]&m[248]&m[786]))):InitCond[337];
    m[349] = run?((((m[158]&~m[249]&m[796])|(~m[158]&m[249]&m[796]))&BiasedRNG[230])|(((m[158]&m[249]&~m[796]))&~BiasedRNG[230])|((m[158]&m[249]&m[796]))):InitCond[338];
    m[352] = run?((((m[89]&~m[252]&m[666])|(~m[89]&m[252]&m[666]))&BiasedRNG[231])|(((m[89]&m[252]&~m[666]))&~BiasedRNG[231])|((m[89]&m[252]&m[666]))):InitCond[339];
    m[353] = run?((((m[99]&~m[253]&m[701])|(~m[99]&m[253]&m[701]))&BiasedRNG[232])|(((m[99]&m[253]&~m[701]))&~BiasedRNG[232])|((m[99]&m[253]&m[701]))):InitCond[340];
    m[354] = run?((((m[109]&~m[254]&m[731])|(~m[109]&m[254]&m[731]))&BiasedRNG[233])|(((m[109]&m[254]&~m[731]))&~BiasedRNG[233])|((m[109]&m[254]&m[731]))):InitCond[341];
    m[355] = run?((((m[119]&~m[255]&m[756])|(~m[119]&m[255]&m[756]))&BiasedRNG[234])|(((m[119]&m[255]&~m[756]))&~BiasedRNG[234])|((m[119]&m[255]&m[756]))):InitCond[342];
    m[356] = run?((((m[129]&~m[256]&m[776])|(~m[129]&m[256]&m[776]))&BiasedRNG[235])|(((m[129]&m[256]&~m[776]))&~BiasedRNG[235])|((m[129]&m[256]&m[776]))):InitCond[343];
    m[357] = run?((((m[139]&~m[257]&m[791])|(~m[139]&m[257]&m[791]))&BiasedRNG[236])|(((m[139]&m[257]&~m[791]))&~BiasedRNG[236])|((m[139]&m[257]&m[791]))):InitCond[344];
    m[358] = run?((((m[149]&~m[258]&m[801])|(~m[149]&m[258]&m[801]))&BiasedRNG[237])|(((m[149]&m[258]&~m[801]))&~BiasedRNG[237])|((m[149]&m[258]&m[801]))):InitCond[345];
    m[359] = run?((((m[159]&~m[259]&m[806])|(~m[159]&m[259]&m[806]))&BiasedRNG[238])|(((m[159]&m[259]&~m[806]))&~BiasedRNG[238])|((m[159]&m[259]&m[806]))):InitCond[346];
    m[360] = run?((((m[261]&~m[361]&~m[362]&~m[363]&~m[364])|(~m[261]&~m[361]&~m[362]&m[363]&~m[364])|(m[261]&m[361]&~m[362]&m[363]&~m[364])|(m[261]&~m[361]&m[362]&m[363]&~m[364])|(~m[261]&m[361]&~m[362]&~m[363]&m[364])|(~m[261]&~m[361]&m[362]&~m[363]&m[364])|(m[261]&m[361]&m[362]&~m[363]&m[364])|(~m[261]&m[361]&m[362]&m[363]&m[364]))&UnbiasedRNG[108])|((m[261]&~m[361]&~m[362]&m[363]&~m[364])|(~m[261]&~m[361]&~m[362]&~m[363]&m[364])|(m[261]&~m[361]&~m[362]&~m[363]&m[364])|(m[261]&m[361]&~m[362]&~m[363]&m[364])|(m[261]&~m[361]&m[362]&~m[363]&m[364])|(~m[261]&~m[361]&~m[362]&m[363]&m[364])|(m[261]&~m[361]&~m[362]&m[363]&m[364])|(~m[261]&m[361]&~m[362]&m[363]&m[364])|(m[261]&m[361]&~m[362]&m[363]&m[364])|(~m[261]&~m[361]&m[362]&m[363]&m[364])|(m[261]&~m[361]&m[362]&m[363]&m[364])|(m[261]&m[361]&m[362]&m[363]&m[364]))):InitCond[347];
    m[366] = run?((((m[271]&~m[365]&~m[367]&~m[368]&~m[369])|(~m[271]&~m[365]&~m[367]&m[368]&~m[369])|(m[271]&m[365]&~m[367]&m[368]&~m[369])|(m[271]&~m[365]&m[367]&m[368]&~m[369])|(~m[271]&m[365]&~m[367]&~m[368]&m[369])|(~m[271]&~m[365]&m[367]&~m[368]&m[369])|(m[271]&m[365]&m[367]&~m[368]&m[369])|(~m[271]&m[365]&m[367]&m[368]&m[369]))&UnbiasedRNG[109])|((m[271]&~m[365]&~m[367]&m[368]&~m[369])|(~m[271]&~m[365]&~m[367]&~m[368]&m[369])|(m[271]&~m[365]&~m[367]&~m[368]&m[369])|(m[271]&m[365]&~m[367]&~m[368]&m[369])|(m[271]&~m[365]&m[367]&~m[368]&m[369])|(~m[271]&~m[365]&~m[367]&m[368]&m[369])|(m[271]&~m[365]&~m[367]&m[368]&m[369])|(~m[271]&m[365]&~m[367]&m[368]&m[369])|(m[271]&m[365]&~m[367]&m[368]&m[369])|(~m[271]&~m[365]&m[367]&m[368]&m[369])|(m[271]&~m[365]&m[367]&m[368]&m[369])|(m[271]&m[365]&m[367]&m[368]&m[369]))):InitCond[348];
    m[371] = run?((((m[280]&~m[370]&~m[372]&~m[373]&~m[374])|(~m[280]&~m[370]&~m[372]&m[373]&~m[374])|(m[280]&m[370]&~m[372]&m[373]&~m[374])|(m[280]&~m[370]&m[372]&m[373]&~m[374])|(~m[280]&m[370]&~m[372]&~m[373]&m[374])|(~m[280]&~m[370]&m[372]&~m[373]&m[374])|(m[280]&m[370]&m[372]&~m[373]&m[374])|(~m[280]&m[370]&m[372]&m[373]&m[374]))&UnbiasedRNG[110])|((m[280]&~m[370]&~m[372]&m[373]&~m[374])|(~m[280]&~m[370]&~m[372]&~m[373]&m[374])|(m[280]&~m[370]&~m[372]&~m[373]&m[374])|(m[280]&m[370]&~m[372]&~m[373]&m[374])|(m[280]&~m[370]&m[372]&~m[373]&m[374])|(~m[280]&~m[370]&~m[372]&m[373]&m[374])|(m[280]&~m[370]&~m[372]&m[373]&m[374])|(~m[280]&m[370]&~m[372]&m[373]&m[374])|(m[280]&m[370]&~m[372]&m[373]&m[374])|(~m[280]&~m[370]&m[372]&m[373]&m[374])|(m[280]&~m[370]&m[372]&m[373]&m[374])|(m[280]&m[370]&m[372]&m[373]&m[374]))):InitCond[349];
    m[376] = run?((((m[272]&~m[375]&~m[377]&~m[378]&~m[379])|(~m[272]&~m[375]&~m[377]&m[378]&~m[379])|(m[272]&m[375]&~m[377]&m[378]&~m[379])|(m[272]&~m[375]&m[377]&m[378]&~m[379])|(~m[272]&m[375]&~m[377]&~m[378]&m[379])|(~m[272]&~m[375]&m[377]&~m[378]&m[379])|(m[272]&m[375]&m[377]&~m[378]&m[379])|(~m[272]&m[375]&m[377]&m[378]&m[379]))&UnbiasedRNG[111])|((m[272]&~m[375]&~m[377]&m[378]&~m[379])|(~m[272]&~m[375]&~m[377]&~m[378]&m[379])|(m[272]&~m[375]&~m[377]&~m[378]&m[379])|(m[272]&m[375]&~m[377]&~m[378]&m[379])|(m[272]&~m[375]&m[377]&~m[378]&m[379])|(~m[272]&~m[375]&~m[377]&m[378]&m[379])|(m[272]&~m[375]&~m[377]&m[378]&m[379])|(~m[272]&m[375]&~m[377]&m[378]&m[379])|(m[272]&m[375]&~m[377]&m[378]&m[379])|(~m[272]&~m[375]&m[377]&m[378]&m[379])|(m[272]&~m[375]&m[377]&m[378]&m[379])|(m[272]&m[375]&m[377]&m[378]&m[379]))):InitCond[350];
    m[381] = run?((((m[281]&~m[380]&~m[382]&~m[383]&~m[384])|(~m[281]&~m[380]&~m[382]&m[383]&~m[384])|(m[281]&m[380]&~m[382]&m[383]&~m[384])|(m[281]&~m[380]&m[382]&m[383]&~m[384])|(~m[281]&m[380]&~m[382]&~m[383]&m[384])|(~m[281]&~m[380]&m[382]&~m[383]&m[384])|(m[281]&m[380]&m[382]&~m[383]&m[384])|(~m[281]&m[380]&m[382]&m[383]&m[384]))&UnbiasedRNG[112])|((m[281]&~m[380]&~m[382]&m[383]&~m[384])|(~m[281]&~m[380]&~m[382]&~m[383]&m[384])|(m[281]&~m[380]&~m[382]&~m[383]&m[384])|(m[281]&m[380]&~m[382]&~m[383]&m[384])|(m[281]&~m[380]&m[382]&~m[383]&m[384])|(~m[281]&~m[380]&~m[382]&m[383]&m[384])|(m[281]&~m[380]&~m[382]&m[383]&m[384])|(~m[281]&m[380]&~m[382]&m[383]&m[384])|(m[281]&m[380]&~m[382]&m[383]&m[384])|(~m[281]&~m[380]&m[382]&m[383]&m[384])|(m[281]&~m[380]&m[382]&m[383]&m[384])|(m[281]&m[380]&m[382]&m[383]&m[384]))):InitCond[351];
    m[386] = run?((((m[290]&~m[385]&~m[387]&~m[388]&~m[389])|(~m[290]&~m[385]&~m[387]&m[388]&~m[389])|(m[290]&m[385]&~m[387]&m[388]&~m[389])|(m[290]&~m[385]&m[387]&m[388]&~m[389])|(~m[290]&m[385]&~m[387]&~m[388]&m[389])|(~m[290]&~m[385]&m[387]&~m[388]&m[389])|(m[290]&m[385]&m[387]&~m[388]&m[389])|(~m[290]&m[385]&m[387]&m[388]&m[389]))&UnbiasedRNG[113])|((m[290]&~m[385]&~m[387]&m[388]&~m[389])|(~m[290]&~m[385]&~m[387]&~m[388]&m[389])|(m[290]&~m[385]&~m[387]&~m[388]&m[389])|(m[290]&m[385]&~m[387]&~m[388]&m[389])|(m[290]&~m[385]&m[387]&~m[388]&m[389])|(~m[290]&~m[385]&~m[387]&m[388]&m[389])|(m[290]&~m[385]&~m[387]&m[388]&m[389])|(~m[290]&m[385]&~m[387]&m[388]&m[389])|(m[290]&m[385]&~m[387]&m[388]&m[389])|(~m[290]&~m[385]&m[387]&m[388]&m[389])|(m[290]&~m[385]&m[387]&m[388]&m[389])|(m[290]&m[385]&m[387]&m[388]&m[389]))):InitCond[352];
    m[391] = run?((((m[273]&~m[390]&~m[392]&~m[393]&~m[394])|(~m[273]&~m[390]&~m[392]&m[393]&~m[394])|(m[273]&m[390]&~m[392]&m[393]&~m[394])|(m[273]&~m[390]&m[392]&m[393]&~m[394])|(~m[273]&m[390]&~m[392]&~m[393]&m[394])|(~m[273]&~m[390]&m[392]&~m[393]&m[394])|(m[273]&m[390]&m[392]&~m[393]&m[394])|(~m[273]&m[390]&m[392]&m[393]&m[394]))&UnbiasedRNG[114])|((m[273]&~m[390]&~m[392]&m[393]&~m[394])|(~m[273]&~m[390]&~m[392]&~m[393]&m[394])|(m[273]&~m[390]&~m[392]&~m[393]&m[394])|(m[273]&m[390]&~m[392]&~m[393]&m[394])|(m[273]&~m[390]&m[392]&~m[393]&m[394])|(~m[273]&~m[390]&~m[392]&m[393]&m[394])|(m[273]&~m[390]&~m[392]&m[393]&m[394])|(~m[273]&m[390]&~m[392]&m[393]&m[394])|(m[273]&m[390]&~m[392]&m[393]&m[394])|(~m[273]&~m[390]&m[392]&m[393]&m[394])|(m[273]&~m[390]&m[392]&m[393]&m[394])|(m[273]&m[390]&m[392]&m[393]&m[394]))):InitCond[353];
    m[397] = run?((((m[384]&~m[395]&~m[396]&~m[398]&~m[399])|(~m[384]&~m[395]&~m[396]&m[398]&~m[399])|(m[384]&m[395]&~m[396]&m[398]&~m[399])|(m[384]&~m[395]&m[396]&m[398]&~m[399])|(~m[384]&m[395]&~m[396]&~m[398]&m[399])|(~m[384]&~m[395]&m[396]&~m[398]&m[399])|(m[384]&m[395]&m[396]&~m[398]&m[399])|(~m[384]&m[395]&m[396]&m[398]&m[399]))&UnbiasedRNG[115])|((m[384]&~m[395]&~m[396]&m[398]&~m[399])|(~m[384]&~m[395]&~m[396]&~m[398]&m[399])|(m[384]&~m[395]&~m[396]&~m[398]&m[399])|(m[384]&m[395]&~m[396]&~m[398]&m[399])|(m[384]&~m[395]&m[396]&~m[398]&m[399])|(~m[384]&~m[395]&~m[396]&m[398]&m[399])|(m[384]&~m[395]&~m[396]&m[398]&m[399])|(~m[384]&m[395]&~m[396]&m[398]&m[399])|(m[384]&m[395]&~m[396]&m[398]&m[399])|(~m[384]&~m[395]&m[396]&m[398]&m[399])|(m[384]&~m[395]&m[396]&m[398]&m[399])|(m[384]&m[395]&m[396]&m[398]&m[399]))):InitCond[354];
    m[401] = run?((((m[291]&~m[400]&~m[402]&~m[403]&~m[404])|(~m[291]&~m[400]&~m[402]&m[403]&~m[404])|(m[291]&m[400]&~m[402]&m[403]&~m[404])|(m[291]&~m[400]&m[402]&m[403]&~m[404])|(~m[291]&m[400]&~m[402]&~m[403]&m[404])|(~m[291]&~m[400]&m[402]&~m[403]&m[404])|(m[291]&m[400]&m[402]&~m[403]&m[404])|(~m[291]&m[400]&m[402]&m[403]&m[404]))&UnbiasedRNG[116])|((m[291]&~m[400]&~m[402]&m[403]&~m[404])|(~m[291]&~m[400]&~m[402]&~m[403]&m[404])|(m[291]&~m[400]&~m[402]&~m[403]&m[404])|(m[291]&m[400]&~m[402]&~m[403]&m[404])|(m[291]&~m[400]&m[402]&~m[403]&m[404])|(~m[291]&~m[400]&~m[402]&m[403]&m[404])|(m[291]&~m[400]&~m[402]&m[403]&m[404])|(~m[291]&m[400]&~m[402]&m[403]&m[404])|(m[291]&m[400]&~m[402]&m[403]&m[404])|(~m[291]&~m[400]&m[402]&m[403]&m[404])|(m[291]&~m[400]&m[402]&m[403]&m[404])|(m[291]&m[400]&m[402]&m[403]&m[404]))):InitCond[355];
    m[406] = run?((((m[300]&~m[405]&~m[407]&~m[408]&~m[409])|(~m[300]&~m[405]&~m[407]&m[408]&~m[409])|(m[300]&m[405]&~m[407]&m[408]&~m[409])|(m[300]&~m[405]&m[407]&m[408]&~m[409])|(~m[300]&m[405]&~m[407]&~m[408]&m[409])|(~m[300]&~m[405]&m[407]&~m[408]&m[409])|(m[300]&m[405]&m[407]&~m[408]&m[409])|(~m[300]&m[405]&m[407]&m[408]&m[409]))&UnbiasedRNG[117])|((m[300]&~m[405]&~m[407]&m[408]&~m[409])|(~m[300]&~m[405]&~m[407]&~m[408]&m[409])|(m[300]&~m[405]&~m[407]&~m[408]&m[409])|(m[300]&m[405]&~m[407]&~m[408]&m[409])|(m[300]&~m[405]&m[407]&~m[408]&m[409])|(~m[300]&~m[405]&~m[407]&m[408]&m[409])|(m[300]&~m[405]&~m[407]&m[408]&m[409])|(~m[300]&m[405]&~m[407]&m[408]&m[409])|(m[300]&m[405]&~m[407]&m[408]&m[409])|(~m[300]&~m[405]&m[407]&m[408]&m[409])|(m[300]&~m[405]&m[407]&m[408]&m[409])|(m[300]&m[405]&m[407]&m[408]&m[409]))):InitCond[356];
    m[411] = run?((((m[274]&~m[410]&~m[412]&~m[413]&~m[414])|(~m[274]&~m[410]&~m[412]&m[413]&~m[414])|(m[274]&m[410]&~m[412]&m[413]&~m[414])|(m[274]&~m[410]&m[412]&m[413]&~m[414])|(~m[274]&m[410]&~m[412]&~m[413]&m[414])|(~m[274]&~m[410]&m[412]&~m[413]&m[414])|(m[274]&m[410]&m[412]&~m[413]&m[414])|(~m[274]&m[410]&m[412]&m[413]&m[414]))&UnbiasedRNG[118])|((m[274]&~m[410]&~m[412]&m[413]&~m[414])|(~m[274]&~m[410]&~m[412]&~m[413]&m[414])|(m[274]&~m[410]&~m[412]&~m[413]&m[414])|(m[274]&m[410]&~m[412]&~m[413]&m[414])|(m[274]&~m[410]&m[412]&~m[413]&m[414])|(~m[274]&~m[410]&~m[412]&m[413]&m[414])|(m[274]&~m[410]&~m[412]&m[413]&m[414])|(~m[274]&m[410]&~m[412]&m[413]&m[414])|(m[274]&m[410]&~m[412]&m[413]&m[414])|(~m[274]&~m[410]&m[412]&m[413]&m[414])|(m[274]&~m[410]&m[412]&m[413]&m[414])|(m[274]&m[410]&m[412]&m[413]&m[414]))):InitCond[357];
    m[417] = run?((((m[399]&~m[415]&~m[416]&~m[418]&~m[419])|(~m[399]&~m[415]&~m[416]&m[418]&~m[419])|(m[399]&m[415]&~m[416]&m[418]&~m[419])|(m[399]&~m[415]&m[416]&m[418]&~m[419])|(~m[399]&m[415]&~m[416]&~m[418]&m[419])|(~m[399]&~m[415]&m[416]&~m[418]&m[419])|(m[399]&m[415]&m[416]&~m[418]&m[419])|(~m[399]&m[415]&m[416]&m[418]&m[419]))&UnbiasedRNG[119])|((m[399]&~m[415]&~m[416]&m[418]&~m[419])|(~m[399]&~m[415]&~m[416]&~m[418]&m[419])|(m[399]&~m[415]&~m[416]&~m[418]&m[419])|(m[399]&m[415]&~m[416]&~m[418]&m[419])|(m[399]&~m[415]&m[416]&~m[418]&m[419])|(~m[399]&~m[415]&~m[416]&m[418]&m[419])|(m[399]&~m[415]&~m[416]&m[418]&m[419])|(~m[399]&m[415]&~m[416]&m[418]&m[419])|(m[399]&m[415]&~m[416]&m[418]&m[419])|(~m[399]&~m[415]&m[416]&m[418]&m[419])|(m[399]&~m[415]&m[416]&m[418]&m[419])|(m[399]&m[415]&m[416]&m[418]&m[419]))):InitCond[358];
    m[422] = run?((((m[404]&~m[420]&~m[421]&~m[423]&~m[424])|(~m[404]&~m[420]&~m[421]&m[423]&~m[424])|(m[404]&m[420]&~m[421]&m[423]&~m[424])|(m[404]&~m[420]&m[421]&m[423]&~m[424])|(~m[404]&m[420]&~m[421]&~m[423]&m[424])|(~m[404]&~m[420]&m[421]&~m[423]&m[424])|(m[404]&m[420]&m[421]&~m[423]&m[424])|(~m[404]&m[420]&m[421]&m[423]&m[424]))&UnbiasedRNG[120])|((m[404]&~m[420]&~m[421]&m[423]&~m[424])|(~m[404]&~m[420]&~m[421]&~m[423]&m[424])|(m[404]&~m[420]&~m[421]&~m[423]&m[424])|(m[404]&m[420]&~m[421]&~m[423]&m[424])|(m[404]&~m[420]&m[421]&~m[423]&m[424])|(~m[404]&~m[420]&~m[421]&m[423]&m[424])|(m[404]&~m[420]&~m[421]&m[423]&m[424])|(~m[404]&m[420]&~m[421]&m[423]&m[424])|(m[404]&m[420]&~m[421]&m[423]&m[424])|(~m[404]&~m[420]&m[421]&m[423]&m[424])|(m[404]&~m[420]&m[421]&m[423]&m[424])|(m[404]&m[420]&m[421]&m[423]&m[424]))):InitCond[359];
    m[426] = run?((((m[301]&~m[425]&~m[427]&~m[428]&~m[429])|(~m[301]&~m[425]&~m[427]&m[428]&~m[429])|(m[301]&m[425]&~m[427]&m[428]&~m[429])|(m[301]&~m[425]&m[427]&m[428]&~m[429])|(~m[301]&m[425]&~m[427]&~m[428]&m[429])|(~m[301]&~m[425]&m[427]&~m[428]&m[429])|(m[301]&m[425]&m[427]&~m[428]&m[429])|(~m[301]&m[425]&m[427]&m[428]&m[429]))&UnbiasedRNG[121])|((m[301]&~m[425]&~m[427]&m[428]&~m[429])|(~m[301]&~m[425]&~m[427]&~m[428]&m[429])|(m[301]&~m[425]&~m[427]&~m[428]&m[429])|(m[301]&m[425]&~m[427]&~m[428]&m[429])|(m[301]&~m[425]&m[427]&~m[428]&m[429])|(~m[301]&~m[425]&~m[427]&m[428]&m[429])|(m[301]&~m[425]&~m[427]&m[428]&m[429])|(~m[301]&m[425]&~m[427]&m[428]&m[429])|(m[301]&m[425]&~m[427]&m[428]&m[429])|(~m[301]&~m[425]&m[427]&m[428]&m[429])|(m[301]&~m[425]&m[427]&m[428]&m[429])|(m[301]&m[425]&m[427]&m[428]&m[429]))):InitCond[360];
    m[431] = run?((((m[310]&~m[430]&~m[432]&~m[433]&~m[434])|(~m[310]&~m[430]&~m[432]&m[433]&~m[434])|(m[310]&m[430]&~m[432]&m[433]&~m[434])|(m[310]&~m[430]&m[432]&m[433]&~m[434])|(~m[310]&m[430]&~m[432]&~m[433]&m[434])|(~m[310]&~m[430]&m[432]&~m[433]&m[434])|(m[310]&m[430]&m[432]&~m[433]&m[434])|(~m[310]&m[430]&m[432]&m[433]&m[434]))&UnbiasedRNG[122])|((m[310]&~m[430]&~m[432]&m[433]&~m[434])|(~m[310]&~m[430]&~m[432]&~m[433]&m[434])|(m[310]&~m[430]&~m[432]&~m[433]&m[434])|(m[310]&m[430]&~m[432]&~m[433]&m[434])|(m[310]&~m[430]&m[432]&~m[433]&m[434])|(~m[310]&~m[430]&~m[432]&m[433]&m[434])|(m[310]&~m[430]&~m[432]&m[433]&m[434])|(~m[310]&m[430]&~m[432]&m[433]&m[434])|(m[310]&m[430]&~m[432]&m[433]&m[434])|(~m[310]&~m[430]&m[432]&m[433]&m[434])|(m[310]&~m[430]&m[432]&m[433]&m[434])|(m[310]&m[430]&m[432]&m[433]&m[434]))):InitCond[361];
    m[436] = run?((((m[275]&~m[435]&~m[437]&~m[438]&~m[439])|(~m[275]&~m[435]&~m[437]&m[438]&~m[439])|(m[275]&m[435]&~m[437]&m[438]&~m[439])|(m[275]&~m[435]&m[437]&m[438]&~m[439])|(~m[275]&m[435]&~m[437]&~m[438]&m[439])|(~m[275]&~m[435]&m[437]&~m[438]&m[439])|(m[275]&m[435]&m[437]&~m[438]&m[439])|(~m[275]&m[435]&m[437]&m[438]&m[439]))&UnbiasedRNG[123])|((m[275]&~m[435]&~m[437]&m[438]&~m[439])|(~m[275]&~m[435]&~m[437]&~m[438]&m[439])|(m[275]&~m[435]&~m[437]&~m[438]&m[439])|(m[275]&m[435]&~m[437]&~m[438]&m[439])|(m[275]&~m[435]&m[437]&~m[438]&m[439])|(~m[275]&~m[435]&~m[437]&m[438]&m[439])|(m[275]&~m[435]&~m[437]&m[438]&m[439])|(~m[275]&m[435]&~m[437]&m[438]&m[439])|(m[275]&m[435]&~m[437]&m[438]&m[439])|(~m[275]&~m[435]&m[437]&m[438]&m[439])|(m[275]&~m[435]&m[437]&m[438]&m[439])|(m[275]&m[435]&m[437]&m[438]&m[439]))):InitCond[362];
    m[442] = run?((((m[419]&~m[440]&~m[441]&~m[443]&~m[444])|(~m[419]&~m[440]&~m[441]&m[443]&~m[444])|(m[419]&m[440]&~m[441]&m[443]&~m[444])|(m[419]&~m[440]&m[441]&m[443]&~m[444])|(~m[419]&m[440]&~m[441]&~m[443]&m[444])|(~m[419]&~m[440]&m[441]&~m[443]&m[444])|(m[419]&m[440]&m[441]&~m[443]&m[444])|(~m[419]&m[440]&m[441]&m[443]&m[444]))&UnbiasedRNG[124])|((m[419]&~m[440]&~m[441]&m[443]&~m[444])|(~m[419]&~m[440]&~m[441]&~m[443]&m[444])|(m[419]&~m[440]&~m[441]&~m[443]&m[444])|(m[419]&m[440]&~m[441]&~m[443]&m[444])|(m[419]&~m[440]&m[441]&~m[443]&m[444])|(~m[419]&~m[440]&~m[441]&m[443]&m[444])|(m[419]&~m[440]&~m[441]&m[443]&m[444])|(~m[419]&m[440]&~m[441]&m[443]&m[444])|(m[419]&m[440]&~m[441]&m[443]&m[444])|(~m[419]&~m[440]&m[441]&m[443]&m[444])|(m[419]&~m[440]&m[441]&m[443]&m[444])|(m[419]&m[440]&m[441]&m[443]&m[444]))):InitCond[363];
    m[447] = run?((((m[424]&~m[445]&~m[446]&~m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&m[448]&~m[449])|(m[424]&m[445]&~m[446]&m[448]&~m[449])|(m[424]&~m[445]&m[446]&m[448]&~m[449])|(~m[424]&m[445]&~m[446]&~m[448]&m[449])|(~m[424]&~m[445]&m[446]&~m[448]&m[449])|(m[424]&m[445]&m[446]&~m[448]&m[449])|(~m[424]&m[445]&m[446]&m[448]&m[449]))&UnbiasedRNG[125])|((m[424]&~m[445]&~m[446]&m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&m[446]&~m[448]&m[449])|(~m[424]&~m[445]&~m[446]&m[448]&m[449])|(m[424]&~m[445]&~m[446]&m[448]&m[449])|(~m[424]&m[445]&~m[446]&m[448]&m[449])|(m[424]&m[445]&~m[446]&m[448]&m[449])|(~m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&m[445]&m[446]&m[448]&m[449]))):InitCond[364];
    m[452] = run?((((m[429]&~m[450]&~m[451]&~m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&m[453]&~m[454])|(m[429]&m[450]&~m[451]&m[453]&~m[454])|(m[429]&~m[450]&m[451]&m[453]&~m[454])|(~m[429]&m[450]&~m[451]&~m[453]&m[454])|(~m[429]&~m[450]&m[451]&~m[453]&m[454])|(m[429]&m[450]&m[451]&~m[453]&m[454])|(~m[429]&m[450]&m[451]&m[453]&m[454]))&UnbiasedRNG[126])|((m[429]&~m[450]&~m[451]&m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&m[451]&~m[453]&m[454])|(~m[429]&~m[450]&~m[451]&m[453]&m[454])|(m[429]&~m[450]&~m[451]&m[453]&m[454])|(~m[429]&m[450]&~m[451]&m[453]&m[454])|(m[429]&m[450]&~m[451]&m[453]&m[454])|(~m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&m[450]&m[451]&m[453]&m[454]))):InitCond[365];
    m[456] = run?((((m[311]&~m[455]&~m[457]&~m[458]&~m[459])|(~m[311]&~m[455]&~m[457]&m[458]&~m[459])|(m[311]&m[455]&~m[457]&m[458]&~m[459])|(m[311]&~m[455]&m[457]&m[458]&~m[459])|(~m[311]&m[455]&~m[457]&~m[458]&m[459])|(~m[311]&~m[455]&m[457]&~m[458]&m[459])|(m[311]&m[455]&m[457]&~m[458]&m[459])|(~m[311]&m[455]&m[457]&m[458]&m[459]))&UnbiasedRNG[127])|((m[311]&~m[455]&~m[457]&m[458]&~m[459])|(~m[311]&~m[455]&~m[457]&~m[458]&m[459])|(m[311]&~m[455]&~m[457]&~m[458]&m[459])|(m[311]&m[455]&~m[457]&~m[458]&m[459])|(m[311]&~m[455]&m[457]&~m[458]&m[459])|(~m[311]&~m[455]&~m[457]&m[458]&m[459])|(m[311]&~m[455]&~m[457]&m[458]&m[459])|(~m[311]&m[455]&~m[457]&m[458]&m[459])|(m[311]&m[455]&~m[457]&m[458]&m[459])|(~m[311]&~m[455]&m[457]&m[458]&m[459])|(m[311]&~m[455]&m[457]&m[458]&m[459])|(m[311]&m[455]&m[457]&m[458]&m[459]))):InitCond[366];
    m[461] = run?((((m[320]&~m[460]&~m[462]&~m[463]&~m[464])|(~m[320]&~m[460]&~m[462]&m[463]&~m[464])|(m[320]&m[460]&~m[462]&m[463]&~m[464])|(m[320]&~m[460]&m[462]&m[463]&~m[464])|(~m[320]&m[460]&~m[462]&~m[463]&m[464])|(~m[320]&~m[460]&m[462]&~m[463]&m[464])|(m[320]&m[460]&m[462]&~m[463]&m[464])|(~m[320]&m[460]&m[462]&m[463]&m[464]))&UnbiasedRNG[128])|((m[320]&~m[460]&~m[462]&m[463]&~m[464])|(~m[320]&~m[460]&~m[462]&~m[463]&m[464])|(m[320]&~m[460]&~m[462]&~m[463]&m[464])|(m[320]&m[460]&~m[462]&~m[463]&m[464])|(m[320]&~m[460]&m[462]&~m[463]&m[464])|(~m[320]&~m[460]&~m[462]&m[463]&m[464])|(m[320]&~m[460]&~m[462]&m[463]&m[464])|(~m[320]&m[460]&~m[462]&m[463]&m[464])|(m[320]&m[460]&~m[462]&m[463]&m[464])|(~m[320]&~m[460]&m[462]&m[463]&m[464])|(m[320]&~m[460]&m[462]&m[463]&m[464])|(m[320]&m[460]&m[462]&m[463]&m[464]))):InitCond[367];
    m[466] = run?((((m[276]&~m[465]&~m[467]&~m[468]&~m[469])|(~m[276]&~m[465]&~m[467]&m[468]&~m[469])|(m[276]&m[465]&~m[467]&m[468]&~m[469])|(m[276]&~m[465]&m[467]&m[468]&~m[469])|(~m[276]&m[465]&~m[467]&~m[468]&m[469])|(~m[276]&~m[465]&m[467]&~m[468]&m[469])|(m[276]&m[465]&m[467]&~m[468]&m[469])|(~m[276]&m[465]&m[467]&m[468]&m[469]))&UnbiasedRNG[129])|((m[276]&~m[465]&~m[467]&m[468]&~m[469])|(~m[276]&~m[465]&~m[467]&~m[468]&m[469])|(m[276]&~m[465]&~m[467]&~m[468]&m[469])|(m[276]&m[465]&~m[467]&~m[468]&m[469])|(m[276]&~m[465]&m[467]&~m[468]&m[469])|(~m[276]&~m[465]&~m[467]&m[468]&m[469])|(m[276]&~m[465]&~m[467]&m[468]&m[469])|(~m[276]&m[465]&~m[467]&m[468]&m[469])|(m[276]&m[465]&~m[467]&m[468]&m[469])|(~m[276]&~m[465]&m[467]&m[468]&m[469])|(m[276]&~m[465]&m[467]&m[468]&m[469])|(m[276]&m[465]&m[467]&m[468]&m[469]))):InitCond[368];
    m[472] = run?((((m[444]&~m[470]&~m[471]&~m[473]&~m[474])|(~m[444]&~m[470]&~m[471]&m[473]&~m[474])|(m[444]&m[470]&~m[471]&m[473]&~m[474])|(m[444]&~m[470]&m[471]&m[473]&~m[474])|(~m[444]&m[470]&~m[471]&~m[473]&m[474])|(~m[444]&~m[470]&m[471]&~m[473]&m[474])|(m[444]&m[470]&m[471]&~m[473]&m[474])|(~m[444]&m[470]&m[471]&m[473]&m[474]))&UnbiasedRNG[130])|((m[444]&~m[470]&~m[471]&m[473]&~m[474])|(~m[444]&~m[470]&~m[471]&~m[473]&m[474])|(m[444]&~m[470]&~m[471]&~m[473]&m[474])|(m[444]&m[470]&~m[471]&~m[473]&m[474])|(m[444]&~m[470]&m[471]&~m[473]&m[474])|(~m[444]&~m[470]&~m[471]&m[473]&m[474])|(m[444]&~m[470]&~m[471]&m[473]&m[474])|(~m[444]&m[470]&~m[471]&m[473]&m[474])|(m[444]&m[470]&~m[471]&m[473]&m[474])|(~m[444]&~m[470]&m[471]&m[473]&m[474])|(m[444]&~m[470]&m[471]&m[473]&m[474])|(m[444]&m[470]&m[471]&m[473]&m[474]))):InitCond[369];
    m[477] = run?((((m[449]&~m[475]&~m[476]&~m[478]&~m[479])|(~m[449]&~m[475]&~m[476]&m[478]&~m[479])|(m[449]&m[475]&~m[476]&m[478]&~m[479])|(m[449]&~m[475]&m[476]&m[478]&~m[479])|(~m[449]&m[475]&~m[476]&~m[478]&m[479])|(~m[449]&~m[475]&m[476]&~m[478]&m[479])|(m[449]&m[475]&m[476]&~m[478]&m[479])|(~m[449]&m[475]&m[476]&m[478]&m[479]))&UnbiasedRNG[131])|((m[449]&~m[475]&~m[476]&m[478]&~m[479])|(~m[449]&~m[475]&~m[476]&~m[478]&m[479])|(m[449]&~m[475]&~m[476]&~m[478]&m[479])|(m[449]&m[475]&~m[476]&~m[478]&m[479])|(m[449]&~m[475]&m[476]&~m[478]&m[479])|(~m[449]&~m[475]&~m[476]&m[478]&m[479])|(m[449]&~m[475]&~m[476]&m[478]&m[479])|(~m[449]&m[475]&~m[476]&m[478]&m[479])|(m[449]&m[475]&~m[476]&m[478]&m[479])|(~m[449]&~m[475]&m[476]&m[478]&m[479])|(m[449]&~m[475]&m[476]&m[478]&m[479])|(m[449]&m[475]&m[476]&m[478]&m[479]))):InitCond[370];
    m[482] = run?((((m[454]&~m[480]&~m[481]&~m[483]&~m[484])|(~m[454]&~m[480]&~m[481]&m[483]&~m[484])|(m[454]&m[480]&~m[481]&m[483]&~m[484])|(m[454]&~m[480]&m[481]&m[483]&~m[484])|(~m[454]&m[480]&~m[481]&~m[483]&m[484])|(~m[454]&~m[480]&m[481]&~m[483]&m[484])|(m[454]&m[480]&m[481]&~m[483]&m[484])|(~m[454]&m[480]&m[481]&m[483]&m[484]))&UnbiasedRNG[132])|((m[454]&~m[480]&~m[481]&m[483]&~m[484])|(~m[454]&~m[480]&~m[481]&~m[483]&m[484])|(m[454]&~m[480]&~m[481]&~m[483]&m[484])|(m[454]&m[480]&~m[481]&~m[483]&m[484])|(m[454]&~m[480]&m[481]&~m[483]&m[484])|(~m[454]&~m[480]&~m[481]&m[483]&m[484])|(m[454]&~m[480]&~m[481]&m[483]&m[484])|(~m[454]&m[480]&~m[481]&m[483]&m[484])|(m[454]&m[480]&~m[481]&m[483]&m[484])|(~m[454]&~m[480]&m[481]&m[483]&m[484])|(m[454]&~m[480]&m[481]&m[483]&m[484])|(m[454]&m[480]&m[481]&m[483]&m[484]))):InitCond[371];
    m[487] = run?((((m[459]&~m[485]&~m[486]&~m[488]&~m[489])|(~m[459]&~m[485]&~m[486]&m[488]&~m[489])|(m[459]&m[485]&~m[486]&m[488]&~m[489])|(m[459]&~m[485]&m[486]&m[488]&~m[489])|(~m[459]&m[485]&~m[486]&~m[488]&m[489])|(~m[459]&~m[485]&m[486]&~m[488]&m[489])|(m[459]&m[485]&m[486]&~m[488]&m[489])|(~m[459]&m[485]&m[486]&m[488]&m[489]))&UnbiasedRNG[133])|((m[459]&~m[485]&~m[486]&m[488]&~m[489])|(~m[459]&~m[485]&~m[486]&~m[488]&m[489])|(m[459]&~m[485]&~m[486]&~m[488]&m[489])|(m[459]&m[485]&~m[486]&~m[488]&m[489])|(m[459]&~m[485]&m[486]&~m[488]&m[489])|(~m[459]&~m[485]&~m[486]&m[488]&m[489])|(m[459]&~m[485]&~m[486]&m[488]&m[489])|(~m[459]&m[485]&~m[486]&m[488]&m[489])|(m[459]&m[485]&~m[486]&m[488]&m[489])|(~m[459]&~m[485]&m[486]&m[488]&m[489])|(m[459]&~m[485]&m[486]&m[488]&m[489])|(m[459]&m[485]&m[486]&m[488]&m[489]))):InitCond[372];
    m[491] = run?((((m[321]&~m[490]&~m[492]&~m[493]&~m[494])|(~m[321]&~m[490]&~m[492]&m[493]&~m[494])|(m[321]&m[490]&~m[492]&m[493]&~m[494])|(m[321]&~m[490]&m[492]&m[493]&~m[494])|(~m[321]&m[490]&~m[492]&~m[493]&m[494])|(~m[321]&~m[490]&m[492]&~m[493]&m[494])|(m[321]&m[490]&m[492]&~m[493]&m[494])|(~m[321]&m[490]&m[492]&m[493]&m[494]))&UnbiasedRNG[134])|((m[321]&~m[490]&~m[492]&m[493]&~m[494])|(~m[321]&~m[490]&~m[492]&~m[493]&m[494])|(m[321]&~m[490]&~m[492]&~m[493]&m[494])|(m[321]&m[490]&~m[492]&~m[493]&m[494])|(m[321]&~m[490]&m[492]&~m[493]&m[494])|(~m[321]&~m[490]&~m[492]&m[493]&m[494])|(m[321]&~m[490]&~m[492]&m[493]&m[494])|(~m[321]&m[490]&~m[492]&m[493]&m[494])|(m[321]&m[490]&~m[492]&m[493]&m[494])|(~m[321]&~m[490]&m[492]&m[493]&m[494])|(m[321]&~m[490]&m[492]&m[493]&m[494])|(m[321]&m[490]&m[492]&m[493]&m[494]))):InitCond[373];
    m[496] = run?((((m[330]&~m[495]&~m[497]&~m[498]&~m[499])|(~m[330]&~m[495]&~m[497]&m[498]&~m[499])|(m[330]&m[495]&~m[497]&m[498]&~m[499])|(m[330]&~m[495]&m[497]&m[498]&~m[499])|(~m[330]&m[495]&~m[497]&~m[498]&m[499])|(~m[330]&~m[495]&m[497]&~m[498]&m[499])|(m[330]&m[495]&m[497]&~m[498]&m[499])|(~m[330]&m[495]&m[497]&m[498]&m[499]))&UnbiasedRNG[135])|((m[330]&~m[495]&~m[497]&m[498]&~m[499])|(~m[330]&~m[495]&~m[497]&~m[498]&m[499])|(m[330]&~m[495]&~m[497]&~m[498]&m[499])|(m[330]&m[495]&~m[497]&~m[498]&m[499])|(m[330]&~m[495]&m[497]&~m[498]&m[499])|(~m[330]&~m[495]&~m[497]&m[498]&m[499])|(m[330]&~m[495]&~m[497]&m[498]&m[499])|(~m[330]&m[495]&~m[497]&m[498]&m[499])|(m[330]&m[495]&~m[497]&m[498]&m[499])|(~m[330]&~m[495]&m[497]&m[498]&m[499])|(m[330]&~m[495]&m[497]&m[498]&m[499])|(m[330]&m[495]&m[497]&m[498]&m[499]))):InitCond[374];
    m[501] = run?((((m[277]&~m[500]&~m[502]&~m[503]&~m[504])|(~m[277]&~m[500]&~m[502]&m[503]&~m[504])|(m[277]&m[500]&~m[502]&m[503]&~m[504])|(m[277]&~m[500]&m[502]&m[503]&~m[504])|(~m[277]&m[500]&~m[502]&~m[503]&m[504])|(~m[277]&~m[500]&m[502]&~m[503]&m[504])|(m[277]&m[500]&m[502]&~m[503]&m[504])|(~m[277]&m[500]&m[502]&m[503]&m[504]))&UnbiasedRNG[136])|((m[277]&~m[500]&~m[502]&m[503]&~m[504])|(~m[277]&~m[500]&~m[502]&~m[503]&m[504])|(m[277]&~m[500]&~m[502]&~m[503]&m[504])|(m[277]&m[500]&~m[502]&~m[503]&m[504])|(m[277]&~m[500]&m[502]&~m[503]&m[504])|(~m[277]&~m[500]&~m[502]&m[503]&m[504])|(m[277]&~m[500]&~m[502]&m[503]&m[504])|(~m[277]&m[500]&~m[502]&m[503]&m[504])|(m[277]&m[500]&~m[502]&m[503]&m[504])|(~m[277]&~m[500]&m[502]&m[503]&m[504])|(m[277]&~m[500]&m[502]&m[503]&m[504])|(m[277]&m[500]&m[502]&m[503]&m[504]))):InitCond[375];
    m[507] = run?((((m[474]&~m[505]&~m[506]&~m[508]&~m[509])|(~m[474]&~m[505]&~m[506]&m[508]&~m[509])|(m[474]&m[505]&~m[506]&m[508]&~m[509])|(m[474]&~m[505]&m[506]&m[508]&~m[509])|(~m[474]&m[505]&~m[506]&~m[508]&m[509])|(~m[474]&~m[505]&m[506]&~m[508]&m[509])|(m[474]&m[505]&m[506]&~m[508]&m[509])|(~m[474]&m[505]&m[506]&m[508]&m[509]))&UnbiasedRNG[137])|((m[474]&~m[505]&~m[506]&m[508]&~m[509])|(~m[474]&~m[505]&~m[506]&~m[508]&m[509])|(m[474]&~m[505]&~m[506]&~m[508]&m[509])|(m[474]&m[505]&~m[506]&~m[508]&m[509])|(m[474]&~m[505]&m[506]&~m[508]&m[509])|(~m[474]&~m[505]&~m[506]&m[508]&m[509])|(m[474]&~m[505]&~m[506]&m[508]&m[509])|(~m[474]&m[505]&~m[506]&m[508]&m[509])|(m[474]&m[505]&~m[506]&m[508]&m[509])|(~m[474]&~m[505]&m[506]&m[508]&m[509])|(m[474]&~m[505]&m[506]&m[508]&m[509])|(m[474]&m[505]&m[506]&m[508]&m[509]))):InitCond[376];
    m[512] = run?((((m[479]&~m[510]&~m[511]&~m[513]&~m[514])|(~m[479]&~m[510]&~m[511]&m[513]&~m[514])|(m[479]&m[510]&~m[511]&m[513]&~m[514])|(m[479]&~m[510]&m[511]&m[513]&~m[514])|(~m[479]&m[510]&~m[511]&~m[513]&m[514])|(~m[479]&~m[510]&m[511]&~m[513]&m[514])|(m[479]&m[510]&m[511]&~m[513]&m[514])|(~m[479]&m[510]&m[511]&m[513]&m[514]))&UnbiasedRNG[138])|((m[479]&~m[510]&~m[511]&m[513]&~m[514])|(~m[479]&~m[510]&~m[511]&~m[513]&m[514])|(m[479]&~m[510]&~m[511]&~m[513]&m[514])|(m[479]&m[510]&~m[511]&~m[513]&m[514])|(m[479]&~m[510]&m[511]&~m[513]&m[514])|(~m[479]&~m[510]&~m[511]&m[513]&m[514])|(m[479]&~m[510]&~m[511]&m[513]&m[514])|(~m[479]&m[510]&~m[511]&m[513]&m[514])|(m[479]&m[510]&~m[511]&m[513]&m[514])|(~m[479]&~m[510]&m[511]&m[513]&m[514])|(m[479]&~m[510]&m[511]&m[513]&m[514])|(m[479]&m[510]&m[511]&m[513]&m[514]))):InitCond[377];
    m[517] = run?((((m[484]&~m[515]&~m[516]&~m[518]&~m[519])|(~m[484]&~m[515]&~m[516]&m[518]&~m[519])|(m[484]&m[515]&~m[516]&m[518]&~m[519])|(m[484]&~m[515]&m[516]&m[518]&~m[519])|(~m[484]&m[515]&~m[516]&~m[518]&m[519])|(~m[484]&~m[515]&m[516]&~m[518]&m[519])|(m[484]&m[515]&m[516]&~m[518]&m[519])|(~m[484]&m[515]&m[516]&m[518]&m[519]))&UnbiasedRNG[139])|((m[484]&~m[515]&~m[516]&m[518]&~m[519])|(~m[484]&~m[515]&~m[516]&~m[518]&m[519])|(m[484]&~m[515]&~m[516]&~m[518]&m[519])|(m[484]&m[515]&~m[516]&~m[518]&m[519])|(m[484]&~m[515]&m[516]&~m[518]&m[519])|(~m[484]&~m[515]&~m[516]&m[518]&m[519])|(m[484]&~m[515]&~m[516]&m[518]&m[519])|(~m[484]&m[515]&~m[516]&m[518]&m[519])|(m[484]&m[515]&~m[516]&m[518]&m[519])|(~m[484]&~m[515]&m[516]&m[518]&m[519])|(m[484]&~m[515]&m[516]&m[518]&m[519])|(m[484]&m[515]&m[516]&m[518]&m[519]))):InitCond[378];
    m[522] = run?((((m[489]&~m[520]&~m[521]&~m[523]&~m[524])|(~m[489]&~m[520]&~m[521]&m[523]&~m[524])|(m[489]&m[520]&~m[521]&m[523]&~m[524])|(m[489]&~m[520]&m[521]&m[523]&~m[524])|(~m[489]&m[520]&~m[521]&~m[523]&m[524])|(~m[489]&~m[520]&m[521]&~m[523]&m[524])|(m[489]&m[520]&m[521]&~m[523]&m[524])|(~m[489]&m[520]&m[521]&m[523]&m[524]))&UnbiasedRNG[140])|((m[489]&~m[520]&~m[521]&m[523]&~m[524])|(~m[489]&~m[520]&~m[521]&~m[523]&m[524])|(m[489]&~m[520]&~m[521]&~m[523]&m[524])|(m[489]&m[520]&~m[521]&~m[523]&m[524])|(m[489]&~m[520]&m[521]&~m[523]&m[524])|(~m[489]&~m[520]&~m[521]&m[523]&m[524])|(m[489]&~m[520]&~m[521]&m[523]&m[524])|(~m[489]&m[520]&~m[521]&m[523]&m[524])|(m[489]&m[520]&~m[521]&m[523]&m[524])|(~m[489]&~m[520]&m[521]&m[523]&m[524])|(m[489]&~m[520]&m[521]&m[523]&m[524])|(m[489]&m[520]&m[521]&m[523]&m[524]))):InitCond[379];
    m[527] = run?((((m[494]&~m[525]&~m[526]&~m[528]&~m[529])|(~m[494]&~m[525]&~m[526]&m[528]&~m[529])|(m[494]&m[525]&~m[526]&m[528]&~m[529])|(m[494]&~m[525]&m[526]&m[528]&~m[529])|(~m[494]&m[525]&~m[526]&~m[528]&m[529])|(~m[494]&~m[525]&m[526]&~m[528]&m[529])|(m[494]&m[525]&m[526]&~m[528]&m[529])|(~m[494]&m[525]&m[526]&m[528]&m[529]))&UnbiasedRNG[141])|((m[494]&~m[525]&~m[526]&m[528]&~m[529])|(~m[494]&~m[525]&~m[526]&~m[528]&m[529])|(m[494]&~m[525]&~m[526]&~m[528]&m[529])|(m[494]&m[525]&~m[526]&~m[528]&m[529])|(m[494]&~m[525]&m[526]&~m[528]&m[529])|(~m[494]&~m[525]&~m[526]&m[528]&m[529])|(m[494]&~m[525]&~m[526]&m[528]&m[529])|(~m[494]&m[525]&~m[526]&m[528]&m[529])|(m[494]&m[525]&~m[526]&m[528]&m[529])|(~m[494]&~m[525]&m[526]&m[528]&m[529])|(m[494]&~m[525]&m[526]&m[528]&m[529])|(m[494]&m[525]&m[526]&m[528]&m[529]))):InitCond[380];
    m[531] = run?((((m[331]&~m[530]&~m[532]&~m[533]&~m[534])|(~m[331]&~m[530]&~m[532]&m[533]&~m[534])|(m[331]&m[530]&~m[532]&m[533]&~m[534])|(m[331]&~m[530]&m[532]&m[533]&~m[534])|(~m[331]&m[530]&~m[532]&~m[533]&m[534])|(~m[331]&~m[530]&m[532]&~m[533]&m[534])|(m[331]&m[530]&m[532]&~m[533]&m[534])|(~m[331]&m[530]&m[532]&m[533]&m[534]))&UnbiasedRNG[142])|((m[331]&~m[530]&~m[532]&m[533]&~m[534])|(~m[331]&~m[530]&~m[532]&~m[533]&m[534])|(m[331]&~m[530]&~m[532]&~m[533]&m[534])|(m[331]&m[530]&~m[532]&~m[533]&m[534])|(m[331]&~m[530]&m[532]&~m[533]&m[534])|(~m[331]&~m[530]&~m[532]&m[533]&m[534])|(m[331]&~m[530]&~m[532]&m[533]&m[534])|(~m[331]&m[530]&~m[532]&m[533]&m[534])|(m[331]&m[530]&~m[532]&m[533]&m[534])|(~m[331]&~m[530]&m[532]&m[533]&m[534])|(m[331]&~m[530]&m[532]&m[533]&m[534])|(m[331]&m[530]&m[532]&m[533]&m[534]))):InitCond[381];
    m[536] = run?((((m[340]&~m[535]&~m[537]&~m[538]&~m[539])|(~m[340]&~m[535]&~m[537]&m[538]&~m[539])|(m[340]&m[535]&~m[537]&m[538]&~m[539])|(m[340]&~m[535]&m[537]&m[538]&~m[539])|(~m[340]&m[535]&~m[537]&~m[538]&m[539])|(~m[340]&~m[535]&m[537]&~m[538]&m[539])|(m[340]&m[535]&m[537]&~m[538]&m[539])|(~m[340]&m[535]&m[537]&m[538]&m[539]))&UnbiasedRNG[143])|((m[340]&~m[535]&~m[537]&m[538]&~m[539])|(~m[340]&~m[535]&~m[537]&~m[538]&m[539])|(m[340]&~m[535]&~m[537]&~m[538]&m[539])|(m[340]&m[535]&~m[537]&~m[538]&m[539])|(m[340]&~m[535]&m[537]&~m[538]&m[539])|(~m[340]&~m[535]&~m[537]&m[538]&m[539])|(m[340]&~m[535]&~m[537]&m[538]&m[539])|(~m[340]&m[535]&~m[537]&m[538]&m[539])|(m[340]&m[535]&~m[537]&m[538]&m[539])|(~m[340]&~m[535]&m[537]&m[538]&m[539])|(m[340]&~m[535]&m[537]&m[538]&m[539])|(m[340]&m[535]&m[537]&m[538]&m[539]))):InitCond[382];
    m[541] = run?((((m[278]&~m[540]&~m[542]&~m[543]&~m[544])|(~m[278]&~m[540]&~m[542]&m[543]&~m[544])|(m[278]&m[540]&~m[542]&m[543]&~m[544])|(m[278]&~m[540]&m[542]&m[543]&~m[544])|(~m[278]&m[540]&~m[542]&~m[543]&m[544])|(~m[278]&~m[540]&m[542]&~m[543]&m[544])|(m[278]&m[540]&m[542]&~m[543]&m[544])|(~m[278]&m[540]&m[542]&m[543]&m[544]))&UnbiasedRNG[144])|((m[278]&~m[540]&~m[542]&m[543]&~m[544])|(~m[278]&~m[540]&~m[542]&~m[543]&m[544])|(m[278]&~m[540]&~m[542]&~m[543]&m[544])|(m[278]&m[540]&~m[542]&~m[543]&m[544])|(m[278]&~m[540]&m[542]&~m[543]&m[544])|(~m[278]&~m[540]&~m[542]&m[543]&m[544])|(m[278]&~m[540]&~m[542]&m[543]&m[544])|(~m[278]&m[540]&~m[542]&m[543]&m[544])|(m[278]&m[540]&~m[542]&m[543]&m[544])|(~m[278]&~m[540]&m[542]&m[543]&m[544])|(m[278]&~m[540]&m[542]&m[543]&m[544])|(m[278]&m[540]&m[542]&m[543]&m[544]))):InitCond[383];
    m[547] = run?((((m[509]&~m[545]&~m[546]&~m[548]&~m[549])|(~m[509]&~m[545]&~m[546]&m[548]&~m[549])|(m[509]&m[545]&~m[546]&m[548]&~m[549])|(m[509]&~m[545]&m[546]&m[548]&~m[549])|(~m[509]&m[545]&~m[546]&~m[548]&m[549])|(~m[509]&~m[545]&m[546]&~m[548]&m[549])|(m[509]&m[545]&m[546]&~m[548]&m[549])|(~m[509]&m[545]&m[546]&m[548]&m[549]))&UnbiasedRNG[145])|((m[509]&~m[545]&~m[546]&m[548]&~m[549])|(~m[509]&~m[545]&~m[546]&~m[548]&m[549])|(m[509]&~m[545]&~m[546]&~m[548]&m[549])|(m[509]&m[545]&~m[546]&~m[548]&m[549])|(m[509]&~m[545]&m[546]&~m[548]&m[549])|(~m[509]&~m[545]&~m[546]&m[548]&m[549])|(m[509]&~m[545]&~m[546]&m[548]&m[549])|(~m[509]&m[545]&~m[546]&m[548]&m[549])|(m[509]&m[545]&~m[546]&m[548]&m[549])|(~m[509]&~m[545]&m[546]&m[548]&m[549])|(m[509]&~m[545]&m[546]&m[548]&m[549])|(m[509]&m[545]&m[546]&m[548]&m[549]))):InitCond[384];
    m[552] = run?((((m[514]&~m[550]&~m[551]&~m[553]&~m[554])|(~m[514]&~m[550]&~m[551]&m[553]&~m[554])|(m[514]&m[550]&~m[551]&m[553]&~m[554])|(m[514]&~m[550]&m[551]&m[553]&~m[554])|(~m[514]&m[550]&~m[551]&~m[553]&m[554])|(~m[514]&~m[550]&m[551]&~m[553]&m[554])|(m[514]&m[550]&m[551]&~m[553]&m[554])|(~m[514]&m[550]&m[551]&m[553]&m[554]))&UnbiasedRNG[146])|((m[514]&~m[550]&~m[551]&m[553]&~m[554])|(~m[514]&~m[550]&~m[551]&~m[553]&m[554])|(m[514]&~m[550]&~m[551]&~m[553]&m[554])|(m[514]&m[550]&~m[551]&~m[553]&m[554])|(m[514]&~m[550]&m[551]&~m[553]&m[554])|(~m[514]&~m[550]&~m[551]&m[553]&m[554])|(m[514]&~m[550]&~m[551]&m[553]&m[554])|(~m[514]&m[550]&~m[551]&m[553]&m[554])|(m[514]&m[550]&~m[551]&m[553]&m[554])|(~m[514]&~m[550]&m[551]&m[553]&m[554])|(m[514]&~m[550]&m[551]&m[553]&m[554])|(m[514]&m[550]&m[551]&m[553]&m[554]))):InitCond[385];
    m[557] = run?((((m[519]&~m[555]&~m[556]&~m[558]&~m[559])|(~m[519]&~m[555]&~m[556]&m[558]&~m[559])|(m[519]&m[555]&~m[556]&m[558]&~m[559])|(m[519]&~m[555]&m[556]&m[558]&~m[559])|(~m[519]&m[555]&~m[556]&~m[558]&m[559])|(~m[519]&~m[555]&m[556]&~m[558]&m[559])|(m[519]&m[555]&m[556]&~m[558]&m[559])|(~m[519]&m[555]&m[556]&m[558]&m[559]))&UnbiasedRNG[147])|((m[519]&~m[555]&~m[556]&m[558]&~m[559])|(~m[519]&~m[555]&~m[556]&~m[558]&m[559])|(m[519]&~m[555]&~m[556]&~m[558]&m[559])|(m[519]&m[555]&~m[556]&~m[558]&m[559])|(m[519]&~m[555]&m[556]&~m[558]&m[559])|(~m[519]&~m[555]&~m[556]&m[558]&m[559])|(m[519]&~m[555]&~m[556]&m[558]&m[559])|(~m[519]&m[555]&~m[556]&m[558]&m[559])|(m[519]&m[555]&~m[556]&m[558]&m[559])|(~m[519]&~m[555]&m[556]&m[558]&m[559])|(m[519]&~m[555]&m[556]&m[558]&m[559])|(m[519]&m[555]&m[556]&m[558]&m[559]))):InitCond[386];
    m[562] = run?((((m[524]&~m[560]&~m[561]&~m[563]&~m[564])|(~m[524]&~m[560]&~m[561]&m[563]&~m[564])|(m[524]&m[560]&~m[561]&m[563]&~m[564])|(m[524]&~m[560]&m[561]&m[563]&~m[564])|(~m[524]&m[560]&~m[561]&~m[563]&m[564])|(~m[524]&~m[560]&m[561]&~m[563]&m[564])|(m[524]&m[560]&m[561]&~m[563]&m[564])|(~m[524]&m[560]&m[561]&m[563]&m[564]))&UnbiasedRNG[148])|((m[524]&~m[560]&~m[561]&m[563]&~m[564])|(~m[524]&~m[560]&~m[561]&~m[563]&m[564])|(m[524]&~m[560]&~m[561]&~m[563]&m[564])|(m[524]&m[560]&~m[561]&~m[563]&m[564])|(m[524]&~m[560]&m[561]&~m[563]&m[564])|(~m[524]&~m[560]&~m[561]&m[563]&m[564])|(m[524]&~m[560]&~m[561]&m[563]&m[564])|(~m[524]&m[560]&~m[561]&m[563]&m[564])|(m[524]&m[560]&~m[561]&m[563]&m[564])|(~m[524]&~m[560]&m[561]&m[563]&m[564])|(m[524]&~m[560]&m[561]&m[563]&m[564])|(m[524]&m[560]&m[561]&m[563]&m[564]))):InitCond[387];
    m[567] = run?((((m[529]&~m[565]&~m[566]&~m[568]&~m[569])|(~m[529]&~m[565]&~m[566]&m[568]&~m[569])|(m[529]&m[565]&~m[566]&m[568]&~m[569])|(m[529]&~m[565]&m[566]&m[568]&~m[569])|(~m[529]&m[565]&~m[566]&~m[568]&m[569])|(~m[529]&~m[565]&m[566]&~m[568]&m[569])|(m[529]&m[565]&m[566]&~m[568]&m[569])|(~m[529]&m[565]&m[566]&m[568]&m[569]))&UnbiasedRNG[149])|((m[529]&~m[565]&~m[566]&m[568]&~m[569])|(~m[529]&~m[565]&~m[566]&~m[568]&m[569])|(m[529]&~m[565]&~m[566]&~m[568]&m[569])|(m[529]&m[565]&~m[566]&~m[568]&m[569])|(m[529]&~m[565]&m[566]&~m[568]&m[569])|(~m[529]&~m[565]&~m[566]&m[568]&m[569])|(m[529]&~m[565]&~m[566]&m[568]&m[569])|(~m[529]&m[565]&~m[566]&m[568]&m[569])|(m[529]&m[565]&~m[566]&m[568]&m[569])|(~m[529]&~m[565]&m[566]&m[568]&m[569])|(m[529]&~m[565]&m[566]&m[568]&m[569])|(m[529]&m[565]&m[566]&m[568]&m[569]))):InitCond[388];
    m[572] = run?((((m[534]&~m[570]&~m[571]&~m[573]&~m[574])|(~m[534]&~m[570]&~m[571]&m[573]&~m[574])|(m[534]&m[570]&~m[571]&m[573]&~m[574])|(m[534]&~m[570]&m[571]&m[573]&~m[574])|(~m[534]&m[570]&~m[571]&~m[573]&m[574])|(~m[534]&~m[570]&m[571]&~m[573]&m[574])|(m[534]&m[570]&m[571]&~m[573]&m[574])|(~m[534]&m[570]&m[571]&m[573]&m[574]))&UnbiasedRNG[150])|((m[534]&~m[570]&~m[571]&m[573]&~m[574])|(~m[534]&~m[570]&~m[571]&~m[573]&m[574])|(m[534]&~m[570]&~m[571]&~m[573]&m[574])|(m[534]&m[570]&~m[571]&~m[573]&m[574])|(m[534]&~m[570]&m[571]&~m[573]&m[574])|(~m[534]&~m[570]&~m[571]&m[573]&m[574])|(m[534]&~m[570]&~m[571]&m[573]&m[574])|(~m[534]&m[570]&~m[571]&m[573]&m[574])|(m[534]&m[570]&~m[571]&m[573]&m[574])|(~m[534]&~m[570]&m[571]&m[573]&m[574])|(m[534]&~m[570]&m[571]&m[573]&m[574])|(m[534]&m[570]&m[571]&m[573]&m[574]))):InitCond[389];
    m[576] = run?((((m[341]&~m[575]&~m[577]&~m[578]&~m[579])|(~m[341]&~m[575]&~m[577]&m[578]&~m[579])|(m[341]&m[575]&~m[577]&m[578]&~m[579])|(m[341]&~m[575]&m[577]&m[578]&~m[579])|(~m[341]&m[575]&~m[577]&~m[578]&m[579])|(~m[341]&~m[575]&m[577]&~m[578]&m[579])|(m[341]&m[575]&m[577]&~m[578]&m[579])|(~m[341]&m[575]&m[577]&m[578]&m[579]))&UnbiasedRNG[151])|((m[341]&~m[575]&~m[577]&m[578]&~m[579])|(~m[341]&~m[575]&~m[577]&~m[578]&m[579])|(m[341]&~m[575]&~m[577]&~m[578]&m[579])|(m[341]&m[575]&~m[577]&~m[578]&m[579])|(m[341]&~m[575]&m[577]&~m[578]&m[579])|(~m[341]&~m[575]&~m[577]&m[578]&m[579])|(m[341]&~m[575]&~m[577]&m[578]&m[579])|(~m[341]&m[575]&~m[577]&m[578]&m[579])|(m[341]&m[575]&~m[577]&m[578]&m[579])|(~m[341]&~m[575]&m[577]&m[578]&m[579])|(m[341]&~m[575]&m[577]&m[578]&m[579])|(m[341]&m[575]&m[577]&m[578]&m[579]))):InitCond[390];
    m[581] = run?((((m[350]&~m[580]&~m[582]&~m[583]&~m[584])|(~m[350]&~m[580]&~m[582]&m[583]&~m[584])|(m[350]&m[580]&~m[582]&m[583]&~m[584])|(m[350]&~m[580]&m[582]&m[583]&~m[584])|(~m[350]&m[580]&~m[582]&~m[583]&m[584])|(~m[350]&~m[580]&m[582]&~m[583]&m[584])|(m[350]&m[580]&m[582]&~m[583]&m[584])|(~m[350]&m[580]&m[582]&m[583]&m[584]))&UnbiasedRNG[152])|((m[350]&~m[580]&~m[582]&m[583]&~m[584])|(~m[350]&~m[580]&~m[582]&~m[583]&m[584])|(m[350]&~m[580]&~m[582]&~m[583]&m[584])|(m[350]&m[580]&~m[582]&~m[583]&m[584])|(m[350]&~m[580]&m[582]&~m[583]&m[584])|(~m[350]&~m[580]&~m[582]&m[583]&m[584])|(m[350]&~m[580]&~m[582]&m[583]&m[584])|(~m[350]&m[580]&~m[582]&m[583]&m[584])|(m[350]&m[580]&~m[582]&m[583]&m[584])|(~m[350]&~m[580]&m[582]&m[583]&m[584])|(m[350]&~m[580]&m[582]&m[583]&m[584])|(m[350]&m[580]&m[582]&m[583]&m[584]))):InitCond[391];
    m[586] = run?((((m[279]&~m[585]&~m[587]&~m[588]&~m[589])|(~m[279]&~m[585]&~m[587]&m[588]&~m[589])|(m[279]&m[585]&~m[587]&m[588]&~m[589])|(m[279]&~m[585]&m[587]&m[588]&~m[589])|(~m[279]&m[585]&~m[587]&~m[588]&m[589])|(~m[279]&~m[585]&m[587]&~m[588]&m[589])|(m[279]&m[585]&m[587]&~m[588]&m[589])|(~m[279]&m[585]&m[587]&m[588]&m[589]))&UnbiasedRNG[153])|((m[279]&~m[585]&~m[587]&m[588]&~m[589])|(~m[279]&~m[585]&~m[587]&~m[588]&m[589])|(m[279]&~m[585]&~m[587]&~m[588]&m[589])|(m[279]&m[585]&~m[587]&~m[588]&m[589])|(m[279]&~m[585]&m[587]&~m[588]&m[589])|(~m[279]&~m[585]&~m[587]&m[588]&m[589])|(m[279]&~m[585]&~m[587]&m[588]&m[589])|(~m[279]&m[585]&~m[587]&m[588]&m[589])|(m[279]&m[585]&~m[587]&m[588]&m[589])|(~m[279]&~m[585]&m[587]&m[588]&m[589])|(m[279]&~m[585]&m[587]&m[588]&m[589])|(m[279]&m[585]&m[587]&m[588]&m[589]))):InitCond[392];
    m[592] = run?((((m[549]&~m[590]&~m[591]&~m[593]&~m[594])|(~m[549]&~m[590]&~m[591]&m[593]&~m[594])|(m[549]&m[590]&~m[591]&m[593]&~m[594])|(m[549]&~m[590]&m[591]&m[593]&~m[594])|(~m[549]&m[590]&~m[591]&~m[593]&m[594])|(~m[549]&~m[590]&m[591]&~m[593]&m[594])|(m[549]&m[590]&m[591]&~m[593]&m[594])|(~m[549]&m[590]&m[591]&m[593]&m[594]))&UnbiasedRNG[154])|((m[549]&~m[590]&~m[591]&m[593]&~m[594])|(~m[549]&~m[590]&~m[591]&~m[593]&m[594])|(m[549]&~m[590]&~m[591]&~m[593]&m[594])|(m[549]&m[590]&~m[591]&~m[593]&m[594])|(m[549]&~m[590]&m[591]&~m[593]&m[594])|(~m[549]&~m[590]&~m[591]&m[593]&m[594])|(m[549]&~m[590]&~m[591]&m[593]&m[594])|(~m[549]&m[590]&~m[591]&m[593]&m[594])|(m[549]&m[590]&~m[591]&m[593]&m[594])|(~m[549]&~m[590]&m[591]&m[593]&m[594])|(m[549]&~m[590]&m[591]&m[593]&m[594])|(m[549]&m[590]&m[591]&m[593]&m[594]))):InitCond[393];
    m[597] = run?((((m[554]&~m[595]&~m[596]&~m[598]&~m[599])|(~m[554]&~m[595]&~m[596]&m[598]&~m[599])|(m[554]&m[595]&~m[596]&m[598]&~m[599])|(m[554]&~m[595]&m[596]&m[598]&~m[599])|(~m[554]&m[595]&~m[596]&~m[598]&m[599])|(~m[554]&~m[595]&m[596]&~m[598]&m[599])|(m[554]&m[595]&m[596]&~m[598]&m[599])|(~m[554]&m[595]&m[596]&m[598]&m[599]))&UnbiasedRNG[155])|((m[554]&~m[595]&~m[596]&m[598]&~m[599])|(~m[554]&~m[595]&~m[596]&~m[598]&m[599])|(m[554]&~m[595]&~m[596]&~m[598]&m[599])|(m[554]&m[595]&~m[596]&~m[598]&m[599])|(m[554]&~m[595]&m[596]&~m[598]&m[599])|(~m[554]&~m[595]&~m[596]&m[598]&m[599])|(m[554]&~m[595]&~m[596]&m[598]&m[599])|(~m[554]&m[595]&~m[596]&m[598]&m[599])|(m[554]&m[595]&~m[596]&m[598]&m[599])|(~m[554]&~m[595]&m[596]&m[598]&m[599])|(m[554]&~m[595]&m[596]&m[598]&m[599])|(m[554]&m[595]&m[596]&m[598]&m[599]))):InitCond[394];
    m[602] = run?((((m[559]&~m[600]&~m[601]&~m[603]&~m[604])|(~m[559]&~m[600]&~m[601]&m[603]&~m[604])|(m[559]&m[600]&~m[601]&m[603]&~m[604])|(m[559]&~m[600]&m[601]&m[603]&~m[604])|(~m[559]&m[600]&~m[601]&~m[603]&m[604])|(~m[559]&~m[600]&m[601]&~m[603]&m[604])|(m[559]&m[600]&m[601]&~m[603]&m[604])|(~m[559]&m[600]&m[601]&m[603]&m[604]))&UnbiasedRNG[156])|((m[559]&~m[600]&~m[601]&m[603]&~m[604])|(~m[559]&~m[600]&~m[601]&~m[603]&m[604])|(m[559]&~m[600]&~m[601]&~m[603]&m[604])|(m[559]&m[600]&~m[601]&~m[603]&m[604])|(m[559]&~m[600]&m[601]&~m[603]&m[604])|(~m[559]&~m[600]&~m[601]&m[603]&m[604])|(m[559]&~m[600]&~m[601]&m[603]&m[604])|(~m[559]&m[600]&~m[601]&m[603]&m[604])|(m[559]&m[600]&~m[601]&m[603]&m[604])|(~m[559]&~m[600]&m[601]&m[603]&m[604])|(m[559]&~m[600]&m[601]&m[603]&m[604])|(m[559]&m[600]&m[601]&m[603]&m[604]))):InitCond[395];
    m[607] = run?((((m[564]&~m[605]&~m[606]&~m[608]&~m[609])|(~m[564]&~m[605]&~m[606]&m[608]&~m[609])|(m[564]&m[605]&~m[606]&m[608]&~m[609])|(m[564]&~m[605]&m[606]&m[608]&~m[609])|(~m[564]&m[605]&~m[606]&~m[608]&m[609])|(~m[564]&~m[605]&m[606]&~m[608]&m[609])|(m[564]&m[605]&m[606]&~m[608]&m[609])|(~m[564]&m[605]&m[606]&m[608]&m[609]))&UnbiasedRNG[157])|((m[564]&~m[605]&~m[606]&m[608]&~m[609])|(~m[564]&~m[605]&~m[606]&~m[608]&m[609])|(m[564]&~m[605]&~m[606]&~m[608]&m[609])|(m[564]&m[605]&~m[606]&~m[608]&m[609])|(m[564]&~m[605]&m[606]&~m[608]&m[609])|(~m[564]&~m[605]&~m[606]&m[608]&m[609])|(m[564]&~m[605]&~m[606]&m[608]&m[609])|(~m[564]&m[605]&~m[606]&m[608]&m[609])|(m[564]&m[605]&~m[606]&m[608]&m[609])|(~m[564]&~m[605]&m[606]&m[608]&m[609])|(m[564]&~m[605]&m[606]&m[608]&m[609])|(m[564]&m[605]&m[606]&m[608]&m[609]))):InitCond[396];
    m[612] = run?((((m[569]&~m[610]&~m[611]&~m[613]&~m[614])|(~m[569]&~m[610]&~m[611]&m[613]&~m[614])|(m[569]&m[610]&~m[611]&m[613]&~m[614])|(m[569]&~m[610]&m[611]&m[613]&~m[614])|(~m[569]&m[610]&~m[611]&~m[613]&m[614])|(~m[569]&~m[610]&m[611]&~m[613]&m[614])|(m[569]&m[610]&m[611]&~m[613]&m[614])|(~m[569]&m[610]&m[611]&m[613]&m[614]))&UnbiasedRNG[158])|((m[569]&~m[610]&~m[611]&m[613]&~m[614])|(~m[569]&~m[610]&~m[611]&~m[613]&m[614])|(m[569]&~m[610]&~m[611]&~m[613]&m[614])|(m[569]&m[610]&~m[611]&~m[613]&m[614])|(m[569]&~m[610]&m[611]&~m[613]&m[614])|(~m[569]&~m[610]&~m[611]&m[613]&m[614])|(m[569]&~m[610]&~m[611]&m[613]&m[614])|(~m[569]&m[610]&~m[611]&m[613]&m[614])|(m[569]&m[610]&~m[611]&m[613]&m[614])|(~m[569]&~m[610]&m[611]&m[613]&m[614])|(m[569]&~m[610]&m[611]&m[613]&m[614])|(m[569]&m[610]&m[611]&m[613]&m[614]))):InitCond[397];
    m[617] = run?((((m[574]&~m[615]&~m[616]&~m[618]&~m[619])|(~m[574]&~m[615]&~m[616]&m[618]&~m[619])|(m[574]&m[615]&~m[616]&m[618]&~m[619])|(m[574]&~m[615]&m[616]&m[618]&~m[619])|(~m[574]&m[615]&~m[616]&~m[618]&m[619])|(~m[574]&~m[615]&m[616]&~m[618]&m[619])|(m[574]&m[615]&m[616]&~m[618]&m[619])|(~m[574]&m[615]&m[616]&m[618]&m[619]))&UnbiasedRNG[159])|((m[574]&~m[615]&~m[616]&m[618]&~m[619])|(~m[574]&~m[615]&~m[616]&~m[618]&m[619])|(m[574]&~m[615]&~m[616]&~m[618]&m[619])|(m[574]&m[615]&~m[616]&~m[618]&m[619])|(m[574]&~m[615]&m[616]&~m[618]&m[619])|(~m[574]&~m[615]&~m[616]&m[618]&m[619])|(m[574]&~m[615]&~m[616]&m[618]&m[619])|(~m[574]&m[615]&~m[616]&m[618]&m[619])|(m[574]&m[615]&~m[616]&m[618]&m[619])|(~m[574]&~m[615]&m[616]&m[618]&m[619])|(m[574]&~m[615]&m[616]&m[618]&m[619])|(m[574]&m[615]&m[616]&m[618]&m[619]))):InitCond[398];
    m[622] = run?((((m[579]&~m[620]&~m[621]&~m[623]&~m[624])|(~m[579]&~m[620]&~m[621]&m[623]&~m[624])|(m[579]&m[620]&~m[621]&m[623]&~m[624])|(m[579]&~m[620]&m[621]&m[623]&~m[624])|(~m[579]&m[620]&~m[621]&~m[623]&m[624])|(~m[579]&~m[620]&m[621]&~m[623]&m[624])|(m[579]&m[620]&m[621]&~m[623]&m[624])|(~m[579]&m[620]&m[621]&m[623]&m[624]))&UnbiasedRNG[160])|((m[579]&~m[620]&~m[621]&m[623]&~m[624])|(~m[579]&~m[620]&~m[621]&~m[623]&m[624])|(m[579]&~m[620]&~m[621]&~m[623]&m[624])|(m[579]&m[620]&~m[621]&~m[623]&m[624])|(m[579]&~m[620]&m[621]&~m[623]&m[624])|(~m[579]&~m[620]&~m[621]&m[623]&m[624])|(m[579]&~m[620]&~m[621]&m[623]&m[624])|(~m[579]&m[620]&~m[621]&m[623]&m[624])|(m[579]&m[620]&~m[621]&m[623]&m[624])|(~m[579]&~m[620]&m[621]&m[623]&m[624])|(m[579]&~m[620]&m[621]&m[623]&m[624])|(m[579]&m[620]&m[621]&m[623]&m[624]))):InitCond[399];
    m[626] = run?((((m[351]&~m[625]&~m[627]&~m[628]&~m[629])|(~m[351]&~m[625]&~m[627]&m[628]&~m[629])|(m[351]&m[625]&~m[627]&m[628]&~m[629])|(m[351]&~m[625]&m[627]&m[628]&~m[629])|(~m[351]&m[625]&~m[627]&~m[628]&m[629])|(~m[351]&~m[625]&m[627]&~m[628]&m[629])|(m[351]&m[625]&m[627]&~m[628]&m[629])|(~m[351]&m[625]&m[627]&m[628]&m[629]))&UnbiasedRNG[161])|((m[351]&~m[625]&~m[627]&m[628]&~m[629])|(~m[351]&~m[625]&~m[627]&~m[628]&m[629])|(m[351]&~m[625]&~m[627]&~m[628]&m[629])|(m[351]&m[625]&~m[627]&~m[628]&m[629])|(m[351]&~m[625]&m[627]&~m[628]&m[629])|(~m[351]&~m[625]&~m[627]&m[628]&m[629])|(m[351]&~m[625]&~m[627]&m[628]&m[629])|(~m[351]&m[625]&~m[627]&m[628]&m[629])|(m[351]&m[625]&~m[627]&m[628]&m[629])|(~m[351]&~m[625]&m[627]&m[628]&m[629])|(m[351]&~m[625]&m[627]&m[628]&m[629])|(m[351]&m[625]&m[627]&m[628]&m[629]))):InitCond[400];
    m[632] = run?((((m[594]&~m[630]&~m[631]&~m[633]&~m[634])|(~m[594]&~m[630]&~m[631]&m[633]&~m[634])|(m[594]&m[630]&~m[631]&m[633]&~m[634])|(m[594]&~m[630]&m[631]&m[633]&~m[634])|(~m[594]&m[630]&~m[631]&~m[633]&m[634])|(~m[594]&~m[630]&m[631]&~m[633]&m[634])|(m[594]&m[630]&m[631]&~m[633]&m[634])|(~m[594]&m[630]&m[631]&m[633]&m[634]))&UnbiasedRNG[162])|((m[594]&~m[630]&~m[631]&m[633]&~m[634])|(~m[594]&~m[630]&~m[631]&~m[633]&m[634])|(m[594]&~m[630]&~m[631]&~m[633]&m[634])|(m[594]&m[630]&~m[631]&~m[633]&m[634])|(m[594]&~m[630]&m[631]&~m[633]&m[634])|(~m[594]&~m[630]&~m[631]&m[633]&m[634])|(m[594]&~m[630]&~m[631]&m[633]&m[634])|(~m[594]&m[630]&~m[631]&m[633]&m[634])|(m[594]&m[630]&~m[631]&m[633]&m[634])|(~m[594]&~m[630]&m[631]&m[633]&m[634])|(m[594]&~m[630]&m[631]&m[633]&m[634])|(m[594]&m[630]&m[631]&m[633]&m[634]))):InitCond[401];
    m[637] = run?((((m[599]&~m[635]&~m[636]&~m[638]&~m[639])|(~m[599]&~m[635]&~m[636]&m[638]&~m[639])|(m[599]&m[635]&~m[636]&m[638]&~m[639])|(m[599]&~m[635]&m[636]&m[638]&~m[639])|(~m[599]&m[635]&~m[636]&~m[638]&m[639])|(~m[599]&~m[635]&m[636]&~m[638]&m[639])|(m[599]&m[635]&m[636]&~m[638]&m[639])|(~m[599]&m[635]&m[636]&m[638]&m[639]))&UnbiasedRNG[163])|((m[599]&~m[635]&~m[636]&m[638]&~m[639])|(~m[599]&~m[635]&~m[636]&~m[638]&m[639])|(m[599]&~m[635]&~m[636]&~m[638]&m[639])|(m[599]&m[635]&~m[636]&~m[638]&m[639])|(m[599]&~m[635]&m[636]&~m[638]&m[639])|(~m[599]&~m[635]&~m[636]&m[638]&m[639])|(m[599]&~m[635]&~m[636]&m[638]&m[639])|(~m[599]&m[635]&~m[636]&m[638]&m[639])|(m[599]&m[635]&~m[636]&m[638]&m[639])|(~m[599]&~m[635]&m[636]&m[638]&m[639])|(m[599]&~m[635]&m[636]&m[638]&m[639])|(m[599]&m[635]&m[636]&m[638]&m[639]))):InitCond[402];
    m[642] = run?((((m[604]&~m[640]&~m[641]&~m[643]&~m[644])|(~m[604]&~m[640]&~m[641]&m[643]&~m[644])|(m[604]&m[640]&~m[641]&m[643]&~m[644])|(m[604]&~m[640]&m[641]&m[643]&~m[644])|(~m[604]&m[640]&~m[641]&~m[643]&m[644])|(~m[604]&~m[640]&m[641]&~m[643]&m[644])|(m[604]&m[640]&m[641]&~m[643]&m[644])|(~m[604]&m[640]&m[641]&m[643]&m[644]))&UnbiasedRNG[164])|((m[604]&~m[640]&~m[641]&m[643]&~m[644])|(~m[604]&~m[640]&~m[641]&~m[643]&m[644])|(m[604]&~m[640]&~m[641]&~m[643]&m[644])|(m[604]&m[640]&~m[641]&~m[643]&m[644])|(m[604]&~m[640]&m[641]&~m[643]&m[644])|(~m[604]&~m[640]&~m[641]&m[643]&m[644])|(m[604]&~m[640]&~m[641]&m[643]&m[644])|(~m[604]&m[640]&~m[641]&m[643]&m[644])|(m[604]&m[640]&~m[641]&m[643]&m[644])|(~m[604]&~m[640]&m[641]&m[643]&m[644])|(m[604]&~m[640]&m[641]&m[643]&m[644])|(m[604]&m[640]&m[641]&m[643]&m[644]))):InitCond[403];
    m[647] = run?((((m[609]&~m[645]&~m[646]&~m[648]&~m[649])|(~m[609]&~m[645]&~m[646]&m[648]&~m[649])|(m[609]&m[645]&~m[646]&m[648]&~m[649])|(m[609]&~m[645]&m[646]&m[648]&~m[649])|(~m[609]&m[645]&~m[646]&~m[648]&m[649])|(~m[609]&~m[645]&m[646]&~m[648]&m[649])|(m[609]&m[645]&m[646]&~m[648]&m[649])|(~m[609]&m[645]&m[646]&m[648]&m[649]))&UnbiasedRNG[165])|((m[609]&~m[645]&~m[646]&m[648]&~m[649])|(~m[609]&~m[645]&~m[646]&~m[648]&m[649])|(m[609]&~m[645]&~m[646]&~m[648]&m[649])|(m[609]&m[645]&~m[646]&~m[648]&m[649])|(m[609]&~m[645]&m[646]&~m[648]&m[649])|(~m[609]&~m[645]&~m[646]&m[648]&m[649])|(m[609]&~m[645]&~m[646]&m[648]&m[649])|(~m[609]&m[645]&~m[646]&m[648]&m[649])|(m[609]&m[645]&~m[646]&m[648]&m[649])|(~m[609]&~m[645]&m[646]&m[648]&m[649])|(m[609]&~m[645]&m[646]&m[648]&m[649])|(m[609]&m[645]&m[646]&m[648]&m[649]))):InitCond[404];
    m[652] = run?((((m[614]&~m[650]&~m[651]&~m[653]&~m[654])|(~m[614]&~m[650]&~m[651]&m[653]&~m[654])|(m[614]&m[650]&~m[651]&m[653]&~m[654])|(m[614]&~m[650]&m[651]&m[653]&~m[654])|(~m[614]&m[650]&~m[651]&~m[653]&m[654])|(~m[614]&~m[650]&m[651]&~m[653]&m[654])|(m[614]&m[650]&m[651]&~m[653]&m[654])|(~m[614]&m[650]&m[651]&m[653]&m[654]))&UnbiasedRNG[166])|((m[614]&~m[650]&~m[651]&m[653]&~m[654])|(~m[614]&~m[650]&~m[651]&~m[653]&m[654])|(m[614]&~m[650]&~m[651]&~m[653]&m[654])|(m[614]&m[650]&~m[651]&~m[653]&m[654])|(m[614]&~m[650]&m[651]&~m[653]&m[654])|(~m[614]&~m[650]&~m[651]&m[653]&m[654])|(m[614]&~m[650]&~m[651]&m[653]&m[654])|(~m[614]&m[650]&~m[651]&m[653]&m[654])|(m[614]&m[650]&~m[651]&m[653]&m[654])|(~m[614]&~m[650]&m[651]&m[653]&m[654])|(m[614]&~m[650]&m[651]&m[653]&m[654])|(m[614]&m[650]&m[651]&m[653]&m[654]))):InitCond[405];
    m[657] = run?((((m[619]&~m[655]&~m[656]&~m[658]&~m[659])|(~m[619]&~m[655]&~m[656]&m[658]&~m[659])|(m[619]&m[655]&~m[656]&m[658]&~m[659])|(m[619]&~m[655]&m[656]&m[658]&~m[659])|(~m[619]&m[655]&~m[656]&~m[658]&m[659])|(~m[619]&~m[655]&m[656]&~m[658]&m[659])|(m[619]&m[655]&m[656]&~m[658]&m[659])|(~m[619]&m[655]&m[656]&m[658]&m[659]))&UnbiasedRNG[167])|((m[619]&~m[655]&~m[656]&m[658]&~m[659])|(~m[619]&~m[655]&~m[656]&~m[658]&m[659])|(m[619]&~m[655]&~m[656]&~m[658]&m[659])|(m[619]&m[655]&~m[656]&~m[658]&m[659])|(m[619]&~m[655]&m[656]&~m[658]&m[659])|(~m[619]&~m[655]&~m[656]&m[658]&m[659])|(m[619]&~m[655]&~m[656]&m[658]&m[659])|(~m[619]&m[655]&~m[656]&m[658]&m[659])|(m[619]&m[655]&~m[656]&m[658]&m[659])|(~m[619]&~m[655]&m[656]&m[658]&m[659])|(m[619]&~m[655]&m[656]&m[658]&m[659])|(m[619]&m[655]&m[656]&m[658]&m[659]))):InitCond[406];
    m[662] = run?((((m[624]&~m[660]&~m[661]&~m[663]&~m[664])|(~m[624]&~m[660]&~m[661]&m[663]&~m[664])|(m[624]&m[660]&~m[661]&m[663]&~m[664])|(m[624]&~m[660]&m[661]&m[663]&~m[664])|(~m[624]&m[660]&~m[661]&~m[663]&m[664])|(~m[624]&~m[660]&m[661]&~m[663]&m[664])|(m[624]&m[660]&m[661]&~m[663]&m[664])|(~m[624]&m[660]&m[661]&m[663]&m[664]))&UnbiasedRNG[168])|((m[624]&~m[660]&~m[661]&m[663]&~m[664])|(~m[624]&~m[660]&~m[661]&~m[663]&m[664])|(m[624]&~m[660]&~m[661]&~m[663]&m[664])|(m[624]&m[660]&~m[661]&~m[663]&m[664])|(m[624]&~m[660]&m[661]&~m[663]&m[664])|(~m[624]&~m[660]&~m[661]&m[663]&m[664])|(m[624]&~m[660]&~m[661]&m[663]&m[664])|(~m[624]&m[660]&~m[661]&m[663]&m[664])|(m[624]&m[660]&~m[661]&m[663]&m[664])|(~m[624]&~m[660]&m[661]&m[663]&m[664])|(m[624]&~m[660]&m[661]&m[663]&m[664])|(m[624]&m[660]&m[661]&m[663]&m[664]))):InitCond[407];
    m[667] = run?((((m[629]&~m[665]&~m[666]&~m[668]&~m[669])|(~m[629]&~m[665]&~m[666]&m[668]&~m[669])|(m[629]&m[665]&~m[666]&m[668]&~m[669])|(m[629]&~m[665]&m[666]&m[668]&~m[669])|(~m[629]&m[665]&~m[666]&~m[668]&m[669])|(~m[629]&~m[665]&m[666]&~m[668]&m[669])|(m[629]&m[665]&m[666]&~m[668]&m[669])|(~m[629]&m[665]&m[666]&m[668]&m[669]))&UnbiasedRNG[169])|((m[629]&~m[665]&~m[666]&m[668]&~m[669])|(~m[629]&~m[665]&~m[666]&~m[668]&m[669])|(m[629]&~m[665]&~m[666]&~m[668]&m[669])|(m[629]&m[665]&~m[666]&~m[668]&m[669])|(m[629]&~m[665]&m[666]&~m[668]&m[669])|(~m[629]&~m[665]&~m[666]&m[668]&m[669])|(m[629]&~m[665]&~m[666]&m[668]&m[669])|(~m[629]&m[665]&~m[666]&m[668]&m[669])|(m[629]&m[665]&~m[666]&m[668]&m[669])|(~m[629]&~m[665]&m[666]&m[668]&m[669])|(m[629]&~m[665]&m[666]&m[668]&m[669])|(m[629]&m[665]&m[666]&m[668]&m[669]))):InitCond[408];
    m[672] = run?((((m[639]&~m[670]&~m[671]&~m[673]&~m[674])|(~m[639]&~m[670]&~m[671]&m[673]&~m[674])|(m[639]&m[670]&~m[671]&m[673]&~m[674])|(m[639]&~m[670]&m[671]&m[673]&~m[674])|(~m[639]&m[670]&~m[671]&~m[673]&m[674])|(~m[639]&~m[670]&m[671]&~m[673]&m[674])|(m[639]&m[670]&m[671]&~m[673]&m[674])|(~m[639]&m[670]&m[671]&m[673]&m[674]))&UnbiasedRNG[170])|((m[639]&~m[670]&~m[671]&m[673]&~m[674])|(~m[639]&~m[670]&~m[671]&~m[673]&m[674])|(m[639]&~m[670]&~m[671]&~m[673]&m[674])|(m[639]&m[670]&~m[671]&~m[673]&m[674])|(m[639]&~m[670]&m[671]&~m[673]&m[674])|(~m[639]&~m[670]&~m[671]&m[673]&m[674])|(m[639]&~m[670]&~m[671]&m[673]&m[674])|(~m[639]&m[670]&~m[671]&m[673]&m[674])|(m[639]&m[670]&~m[671]&m[673]&m[674])|(~m[639]&~m[670]&m[671]&m[673]&m[674])|(m[639]&~m[670]&m[671]&m[673]&m[674])|(m[639]&m[670]&m[671]&m[673]&m[674]))):InitCond[409];
    m[677] = run?((((m[644]&~m[675]&~m[676]&~m[678]&~m[679])|(~m[644]&~m[675]&~m[676]&m[678]&~m[679])|(m[644]&m[675]&~m[676]&m[678]&~m[679])|(m[644]&~m[675]&m[676]&m[678]&~m[679])|(~m[644]&m[675]&~m[676]&~m[678]&m[679])|(~m[644]&~m[675]&m[676]&~m[678]&m[679])|(m[644]&m[675]&m[676]&~m[678]&m[679])|(~m[644]&m[675]&m[676]&m[678]&m[679]))&UnbiasedRNG[171])|((m[644]&~m[675]&~m[676]&m[678]&~m[679])|(~m[644]&~m[675]&~m[676]&~m[678]&m[679])|(m[644]&~m[675]&~m[676]&~m[678]&m[679])|(m[644]&m[675]&~m[676]&~m[678]&m[679])|(m[644]&~m[675]&m[676]&~m[678]&m[679])|(~m[644]&~m[675]&~m[676]&m[678]&m[679])|(m[644]&~m[675]&~m[676]&m[678]&m[679])|(~m[644]&m[675]&~m[676]&m[678]&m[679])|(m[644]&m[675]&~m[676]&m[678]&m[679])|(~m[644]&~m[675]&m[676]&m[678]&m[679])|(m[644]&~m[675]&m[676]&m[678]&m[679])|(m[644]&m[675]&m[676]&m[678]&m[679]))):InitCond[410];
    m[682] = run?((((m[649]&~m[680]&~m[681]&~m[683]&~m[684])|(~m[649]&~m[680]&~m[681]&m[683]&~m[684])|(m[649]&m[680]&~m[681]&m[683]&~m[684])|(m[649]&~m[680]&m[681]&m[683]&~m[684])|(~m[649]&m[680]&~m[681]&~m[683]&m[684])|(~m[649]&~m[680]&m[681]&~m[683]&m[684])|(m[649]&m[680]&m[681]&~m[683]&m[684])|(~m[649]&m[680]&m[681]&m[683]&m[684]))&UnbiasedRNG[172])|((m[649]&~m[680]&~m[681]&m[683]&~m[684])|(~m[649]&~m[680]&~m[681]&~m[683]&m[684])|(m[649]&~m[680]&~m[681]&~m[683]&m[684])|(m[649]&m[680]&~m[681]&~m[683]&m[684])|(m[649]&~m[680]&m[681]&~m[683]&m[684])|(~m[649]&~m[680]&~m[681]&m[683]&m[684])|(m[649]&~m[680]&~m[681]&m[683]&m[684])|(~m[649]&m[680]&~m[681]&m[683]&m[684])|(m[649]&m[680]&~m[681]&m[683]&m[684])|(~m[649]&~m[680]&m[681]&m[683]&m[684])|(m[649]&~m[680]&m[681]&m[683]&m[684])|(m[649]&m[680]&m[681]&m[683]&m[684]))):InitCond[411];
    m[687] = run?((((m[654]&~m[685]&~m[686]&~m[688]&~m[689])|(~m[654]&~m[685]&~m[686]&m[688]&~m[689])|(m[654]&m[685]&~m[686]&m[688]&~m[689])|(m[654]&~m[685]&m[686]&m[688]&~m[689])|(~m[654]&m[685]&~m[686]&~m[688]&m[689])|(~m[654]&~m[685]&m[686]&~m[688]&m[689])|(m[654]&m[685]&m[686]&~m[688]&m[689])|(~m[654]&m[685]&m[686]&m[688]&m[689]))&UnbiasedRNG[173])|((m[654]&~m[685]&~m[686]&m[688]&~m[689])|(~m[654]&~m[685]&~m[686]&~m[688]&m[689])|(m[654]&~m[685]&~m[686]&~m[688]&m[689])|(m[654]&m[685]&~m[686]&~m[688]&m[689])|(m[654]&~m[685]&m[686]&~m[688]&m[689])|(~m[654]&~m[685]&~m[686]&m[688]&m[689])|(m[654]&~m[685]&~m[686]&m[688]&m[689])|(~m[654]&m[685]&~m[686]&m[688]&m[689])|(m[654]&m[685]&~m[686]&m[688]&m[689])|(~m[654]&~m[685]&m[686]&m[688]&m[689])|(m[654]&~m[685]&m[686]&m[688]&m[689])|(m[654]&m[685]&m[686]&m[688]&m[689]))):InitCond[412];
    m[692] = run?((((m[659]&~m[690]&~m[691]&~m[693]&~m[694])|(~m[659]&~m[690]&~m[691]&m[693]&~m[694])|(m[659]&m[690]&~m[691]&m[693]&~m[694])|(m[659]&~m[690]&m[691]&m[693]&~m[694])|(~m[659]&m[690]&~m[691]&~m[693]&m[694])|(~m[659]&~m[690]&m[691]&~m[693]&m[694])|(m[659]&m[690]&m[691]&~m[693]&m[694])|(~m[659]&m[690]&m[691]&m[693]&m[694]))&UnbiasedRNG[174])|((m[659]&~m[690]&~m[691]&m[693]&~m[694])|(~m[659]&~m[690]&~m[691]&~m[693]&m[694])|(m[659]&~m[690]&~m[691]&~m[693]&m[694])|(m[659]&m[690]&~m[691]&~m[693]&m[694])|(m[659]&~m[690]&m[691]&~m[693]&m[694])|(~m[659]&~m[690]&~m[691]&m[693]&m[694])|(m[659]&~m[690]&~m[691]&m[693]&m[694])|(~m[659]&m[690]&~m[691]&m[693]&m[694])|(m[659]&m[690]&~m[691]&m[693]&m[694])|(~m[659]&~m[690]&m[691]&m[693]&m[694])|(m[659]&~m[690]&m[691]&m[693]&m[694])|(m[659]&m[690]&m[691]&m[693]&m[694]))):InitCond[413];
    m[697] = run?((((m[664]&~m[695]&~m[696]&~m[698]&~m[699])|(~m[664]&~m[695]&~m[696]&m[698]&~m[699])|(m[664]&m[695]&~m[696]&m[698]&~m[699])|(m[664]&~m[695]&m[696]&m[698]&~m[699])|(~m[664]&m[695]&~m[696]&~m[698]&m[699])|(~m[664]&~m[695]&m[696]&~m[698]&m[699])|(m[664]&m[695]&m[696]&~m[698]&m[699])|(~m[664]&m[695]&m[696]&m[698]&m[699]))&UnbiasedRNG[175])|((m[664]&~m[695]&~m[696]&m[698]&~m[699])|(~m[664]&~m[695]&~m[696]&~m[698]&m[699])|(m[664]&~m[695]&~m[696]&~m[698]&m[699])|(m[664]&m[695]&~m[696]&~m[698]&m[699])|(m[664]&~m[695]&m[696]&~m[698]&m[699])|(~m[664]&~m[695]&~m[696]&m[698]&m[699])|(m[664]&~m[695]&~m[696]&m[698]&m[699])|(~m[664]&m[695]&~m[696]&m[698]&m[699])|(m[664]&m[695]&~m[696]&m[698]&m[699])|(~m[664]&~m[695]&m[696]&m[698]&m[699])|(m[664]&~m[695]&m[696]&m[698]&m[699])|(m[664]&m[695]&m[696]&m[698]&m[699]))):InitCond[414];
    m[702] = run?((((m[669]&~m[700]&~m[701]&~m[703]&~m[704])|(~m[669]&~m[700]&~m[701]&m[703]&~m[704])|(m[669]&m[700]&~m[701]&m[703]&~m[704])|(m[669]&~m[700]&m[701]&m[703]&~m[704])|(~m[669]&m[700]&~m[701]&~m[703]&m[704])|(~m[669]&~m[700]&m[701]&~m[703]&m[704])|(m[669]&m[700]&m[701]&~m[703]&m[704])|(~m[669]&m[700]&m[701]&m[703]&m[704]))&UnbiasedRNG[176])|((m[669]&~m[700]&~m[701]&m[703]&~m[704])|(~m[669]&~m[700]&~m[701]&~m[703]&m[704])|(m[669]&~m[700]&~m[701]&~m[703]&m[704])|(m[669]&m[700]&~m[701]&~m[703]&m[704])|(m[669]&~m[700]&m[701]&~m[703]&m[704])|(~m[669]&~m[700]&~m[701]&m[703]&m[704])|(m[669]&~m[700]&~m[701]&m[703]&m[704])|(~m[669]&m[700]&~m[701]&m[703]&m[704])|(m[669]&m[700]&~m[701]&m[703]&m[704])|(~m[669]&~m[700]&m[701]&m[703]&m[704])|(m[669]&~m[700]&m[701]&m[703]&m[704])|(m[669]&m[700]&m[701]&m[703]&m[704]))):InitCond[415];
    m[707] = run?((((m[679]&~m[705]&~m[706]&~m[708]&~m[709])|(~m[679]&~m[705]&~m[706]&m[708]&~m[709])|(m[679]&m[705]&~m[706]&m[708]&~m[709])|(m[679]&~m[705]&m[706]&m[708]&~m[709])|(~m[679]&m[705]&~m[706]&~m[708]&m[709])|(~m[679]&~m[705]&m[706]&~m[708]&m[709])|(m[679]&m[705]&m[706]&~m[708]&m[709])|(~m[679]&m[705]&m[706]&m[708]&m[709]))&UnbiasedRNG[177])|((m[679]&~m[705]&~m[706]&m[708]&~m[709])|(~m[679]&~m[705]&~m[706]&~m[708]&m[709])|(m[679]&~m[705]&~m[706]&~m[708]&m[709])|(m[679]&m[705]&~m[706]&~m[708]&m[709])|(m[679]&~m[705]&m[706]&~m[708]&m[709])|(~m[679]&~m[705]&~m[706]&m[708]&m[709])|(m[679]&~m[705]&~m[706]&m[708]&m[709])|(~m[679]&m[705]&~m[706]&m[708]&m[709])|(m[679]&m[705]&~m[706]&m[708]&m[709])|(~m[679]&~m[705]&m[706]&m[708]&m[709])|(m[679]&~m[705]&m[706]&m[708]&m[709])|(m[679]&m[705]&m[706]&m[708]&m[709]))):InitCond[416];
    m[712] = run?((((m[684]&~m[710]&~m[711]&~m[713]&~m[714])|(~m[684]&~m[710]&~m[711]&m[713]&~m[714])|(m[684]&m[710]&~m[711]&m[713]&~m[714])|(m[684]&~m[710]&m[711]&m[713]&~m[714])|(~m[684]&m[710]&~m[711]&~m[713]&m[714])|(~m[684]&~m[710]&m[711]&~m[713]&m[714])|(m[684]&m[710]&m[711]&~m[713]&m[714])|(~m[684]&m[710]&m[711]&m[713]&m[714]))&UnbiasedRNG[178])|((m[684]&~m[710]&~m[711]&m[713]&~m[714])|(~m[684]&~m[710]&~m[711]&~m[713]&m[714])|(m[684]&~m[710]&~m[711]&~m[713]&m[714])|(m[684]&m[710]&~m[711]&~m[713]&m[714])|(m[684]&~m[710]&m[711]&~m[713]&m[714])|(~m[684]&~m[710]&~m[711]&m[713]&m[714])|(m[684]&~m[710]&~m[711]&m[713]&m[714])|(~m[684]&m[710]&~m[711]&m[713]&m[714])|(m[684]&m[710]&~m[711]&m[713]&m[714])|(~m[684]&~m[710]&m[711]&m[713]&m[714])|(m[684]&~m[710]&m[711]&m[713]&m[714])|(m[684]&m[710]&m[711]&m[713]&m[714]))):InitCond[417];
    m[717] = run?((((m[689]&~m[715]&~m[716]&~m[718]&~m[719])|(~m[689]&~m[715]&~m[716]&m[718]&~m[719])|(m[689]&m[715]&~m[716]&m[718]&~m[719])|(m[689]&~m[715]&m[716]&m[718]&~m[719])|(~m[689]&m[715]&~m[716]&~m[718]&m[719])|(~m[689]&~m[715]&m[716]&~m[718]&m[719])|(m[689]&m[715]&m[716]&~m[718]&m[719])|(~m[689]&m[715]&m[716]&m[718]&m[719]))&UnbiasedRNG[179])|((m[689]&~m[715]&~m[716]&m[718]&~m[719])|(~m[689]&~m[715]&~m[716]&~m[718]&m[719])|(m[689]&~m[715]&~m[716]&~m[718]&m[719])|(m[689]&m[715]&~m[716]&~m[718]&m[719])|(m[689]&~m[715]&m[716]&~m[718]&m[719])|(~m[689]&~m[715]&~m[716]&m[718]&m[719])|(m[689]&~m[715]&~m[716]&m[718]&m[719])|(~m[689]&m[715]&~m[716]&m[718]&m[719])|(m[689]&m[715]&~m[716]&m[718]&m[719])|(~m[689]&~m[715]&m[716]&m[718]&m[719])|(m[689]&~m[715]&m[716]&m[718]&m[719])|(m[689]&m[715]&m[716]&m[718]&m[719]))):InitCond[418];
    m[722] = run?((((m[694]&~m[720]&~m[721]&~m[723]&~m[724])|(~m[694]&~m[720]&~m[721]&m[723]&~m[724])|(m[694]&m[720]&~m[721]&m[723]&~m[724])|(m[694]&~m[720]&m[721]&m[723]&~m[724])|(~m[694]&m[720]&~m[721]&~m[723]&m[724])|(~m[694]&~m[720]&m[721]&~m[723]&m[724])|(m[694]&m[720]&m[721]&~m[723]&m[724])|(~m[694]&m[720]&m[721]&m[723]&m[724]))&UnbiasedRNG[180])|((m[694]&~m[720]&~m[721]&m[723]&~m[724])|(~m[694]&~m[720]&~m[721]&~m[723]&m[724])|(m[694]&~m[720]&~m[721]&~m[723]&m[724])|(m[694]&m[720]&~m[721]&~m[723]&m[724])|(m[694]&~m[720]&m[721]&~m[723]&m[724])|(~m[694]&~m[720]&~m[721]&m[723]&m[724])|(m[694]&~m[720]&~m[721]&m[723]&m[724])|(~m[694]&m[720]&~m[721]&m[723]&m[724])|(m[694]&m[720]&~m[721]&m[723]&m[724])|(~m[694]&~m[720]&m[721]&m[723]&m[724])|(m[694]&~m[720]&m[721]&m[723]&m[724])|(m[694]&m[720]&m[721]&m[723]&m[724]))):InitCond[419];
    m[727] = run?((((m[699]&~m[725]&~m[726]&~m[728]&~m[729])|(~m[699]&~m[725]&~m[726]&m[728]&~m[729])|(m[699]&m[725]&~m[726]&m[728]&~m[729])|(m[699]&~m[725]&m[726]&m[728]&~m[729])|(~m[699]&m[725]&~m[726]&~m[728]&m[729])|(~m[699]&~m[725]&m[726]&~m[728]&m[729])|(m[699]&m[725]&m[726]&~m[728]&m[729])|(~m[699]&m[725]&m[726]&m[728]&m[729]))&UnbiasedRNG[181])|((m[699]&~m[725]&~m[726]&m[728]&~m[729])|(~m[699]&~m[725]&~m[726]&~m[728]&m[729])|(m[699]&~m[725]&~m[726]&~m[728]&m[729])|(m[699]&m[725]&~m[726]&~m[728]&m[729])|(m[699]&~m[725]&m[726]&~m[728]&m[729])|(~m[699]&~m[725]&~m[726]&m[728]&m[729])|(m[699]&~m[725]&~m[726]&m[728]&m[729])|(~m[699]&m[725]&~m[726]&m[728]&m[729])|(m[699]&m[725]&~m[726]&m[728]&m[729])|(~m[699]&~m[725]&m[726]&m[728]&m[729])|(m[699]&~m[725]&m[726]&m[728]&m[729])|(m[699]&m[725]&m[726]&m[728]&m[729]))):InitCond[420];
    m[732] = run?((((m[704]&~m[730]&~m[731]&~m[733]&~m[734])|(~m[704]&~m[730]&~m[731]&m[733]&~m[734])|(m[704]&m[730]&~m[731]&m[733]&~m[734])|(m[704]&~m[730]&m[731]&m[733]&~m[734])|(~m[704]&m[730]&~m[731]&~m[733]&m[734])|(~m[704]&~m[730]&m[731]&~m[733]&m[734])|(m[704]&m[730]&m[731]&~m[733]&m[734])|(~m[704]&m[730]&m[731]&m[733]&m[734]))&UnbiasedRNG[182])|((m[704]&~m[730]&~m[731]&m[733]&~m[734])|(~m[704]&~m[730]&~m[731]&~m[733]&m[734])|(m[704]&~m[730]&~m[731]&~m[733]&m[734])|(m[704]&m[730]&~m[731]&~m[733]&m[734])|(m[704]&~m[730]&m[731]&~m[733]&m[734])|(~m[704]&~m[730]&~m[731]&m[733]&m[734])|(m[704]&~m[730]&~m[731]&m[733]&m[734])|(~m[704]&m[730]&~m[731]&m[733]&m[734])|(m[704]&m[730]&~m[731]&m[733]&m[734])|(~m[704]&~m[730]&m[731]&m[733]&m[734])|(m[704]&~m[730]&m[731]&m[733]&m[734])|(m[704]&m[730]&m[731]&m[733]&m[734]))):InitCond[421];
    m[737] = run?((((m[714]&~m[735]&~m[736]&~m[738]&~m[739])|(~m[714]&~m[735]&~m[736]&m[738]&~m[739])|(m[714]&m[735]&~m[736]&m[738]&~m[739])|(m[714]&~m[735]&m[736]&m[738]&~m[739])|(~m[714]&m[735]&~m[736]&~m[738]&m[739])|(~m[714]&~m[735]&m[736]&~m[738]&m[739])|(m[714]&m[735]&m[736]&~m[738]&m[739])|(~m[714]&m[735]&m[736]&m[738]&m[739]))&UnbiasedRNG[183])|((m[714]&~m[735]&~m[736]&m[738]&~m[739])|(~m[714]&~m[735]&~m[736]&~m[738]&m[739])|(m[714]&~m[735]&~m[736]&~m[738]&m[739])|(m[714]&m[735]&~m[736]&~m[738]&m[739])|(m[714]&~m[735]&m[736]&~m[738]&m[739])|(~m[714]&~m[735]&~m[736]&m[738]&m[739])|(m[714]&~m[735]&~m[736]&m[738]&m[739])|(~m[714]&m[735]&~m[736]&m[738]&m[739])|(m[714]&m[735]&~m[736]&m[738]&m[739])|(~m[714]&~m[735]&m[736]&m[738]&m[739])|(m[714]&~m[735]&m[736]&m[738]&m[739])|(m[714]&m[735]&m[736]&m[738]&m[739]))):InitCond[422];
    m[742] = run?((((m[719]&~m[740]&~m[741]&~m[743]&~m[744])|(~m[719]&~m[740]&~m[741]&m[743]&~m[744])|(m[719]&m[740]&~m[741]&m[743]&~m[744])|(m[719]&~m[740]&m[741]&m[743]&~m[744])|(~m[719]&m[740]&~m[741]&~m[743]&m[744])|(~m[719]&~m[740]&m[741]&~m[743]&m[744])|(m[719]&m[740]&m[741]&~m[743]&m[744])|(~m[719]&m[740]&m[741]&m[743]&m[744]))&UnbiasedRNG[184])|((m[719]&~m[740]&~m[741]&m[743]&~m[744])|(~m[719]&~m[740]&~m[741]&~m[743]&m[744])|(m[719]&~m[740]&~m[741]&~m[743]&m[744])|(m[719]&m[740]&~m[741]&~m[743]&m[744])|(m[719]&~m[740]&m[741]&~m[743]&m[744])|(~m[719]&~m[740]&~m[741]&m[743]&m[744])|(m[719]&~m[740]&~m[741]&m[743]&m[744])|(~m[719]&m[740]&~m[741]&m[743]&m[744])|(m[719]&m[740]&~m[741]&m[743]&m[744])|(~m[719]&~m[740]&m[741]&m[743]&m[744])|(m[719]&~m[740]&m[741]&m[743]&m[744])|(m[719]&m[740]&m[741]&m[743]&m[744]))):InitCond[423];
    m[747] = run?((((m[724]&~m[745]&~m[746]&~m[748]&~m[749])|(~m[724]&~m[745]&~m[746]&m[748]&~m[749])|(m[724]&m[745]&~m[746]&m[748]&~m[749])|(m[724]&~m[745]&m[746]&m[748]&~m[749])|(~m[724]&m[745]&~m[746]&~m[748]&m[749])|(~m[724]&~m[745]&m[746]&~m[748]&m[749])|(m[724]&m[745]&m[746]&~m[748]&m[749])|(~m[724]&m[745]&m[746]&m[748]&m[749]))&UnbiasedRNG[185])|((m[724]&~m[745]&~m[746]&m[748]&~m[749])|(~m[724]&~m[745]&~m[746]&~m[748]&m[749])|(m[724]&~m[745]&~m[746]&~m[748]&m[749])|(m[724]&m[745]&~m[746]&~m[748]&m[749])|(m[724]&~m[745]&m[746]&~m[748]&m[749])|(~m[724]&~m[745]&~m[746]&m[748]&m[749])|(m[724]&~m[745]&~m[746]&m[748]&m[749])|(~m[724]&m[745]&~m[746]&m[748]&m[749])|(m[724]&m[745]&~m[746]&m[748]&m[749])|(~m[724]&~m[745]&m[746]&m[748]&m[749])|(m[724]&~m[745]&m[746]&m[748]&m[749])|(m[724]&m[745]&m[746]&m[748]&m[749]))):InitCond[424];
    m[752] = run?((((m[729]&~m[750]&~m[751]&~m[753]&~m[754])|(~m[729]&~m[750]&~m[751]&m[753]&~m[754])|(m[729]&m[750]&~m[751]&m[753]&~m[754])|(m[729]&~m[750]&m[751]&m[753]&~m[754])|(~m[729]&m[750]&~m[751]&~m[753]&m[754])|(~m[729]&~m[750]&m[751]&~m[753]&m[754])|(m[729]&m[750]&m[751]&~m[753]&m[754])|(~m[729]&m[750]&m[751]&m[753]&m[754]))&UnbiasedRNG[186])|((m[729]&~m[750]&~m[751]&m[753]&~m[754])|(~m[729]&~m[750]&~m[751]&~m[753]&m[754])|(m[729]&~m[750]&~m[751]&~m[753]&m[754])|(m[729]&m[750]&~m[751]&~m[753]&m[754])|(m[729]&~m[750]&m[751]&~m[753]&m[754])|(~m[729]&~m[750]&~m[751]&m[753]&m[754])|(m[729]&~m[750]&~m[751]&m[753]&m[754])|(~m[729]&m[750]&~m[751]&m[753]&m[754])|(m[729]&m[750]&~m[751]&m[753]&m[754])|(~m[729]&~m[750]&m[751]&m[753]&m[754])|(m[729]&~m[750]&m[751]&m[753]&m[754])|(m[729]&m[750]&m[751]&m[753]&m[754]))):InitCond[425];
    m[757] = run?((((m[734]&~m[755]&~m[756]&~m[758]&~m[759])|(~m[734]&~m[755]&~m[756]&m[758]&~m[759])|(m[734]&m[755]&~m[756]&m[758]&~m[759])|(m[734]&~m[755]&m[756]&m[758]&~m[759])|(~m[734]&m[755]&~m[756]&~m[758]&m[759])|(~m[734]&~m[755]&m[756]&~m[758]&m[759])|(m[734]&m[755]&m[756]&~m[758]&m[759])|(~m[734]&m[755]&m[756]&m[758]&m[759]))&UnbiasedRNG[187])|((m[734]&~m[755]&~m[756]&m[758]&~m[759])|(~m[734]&~m[755]&~m[756]&~m[758]&m[759])|(m[734]&~m[755]&~m[756]&~m[758]&m[759])|(m[734]&m[755]&~m[756]&~m[758]&m[759])|(m[734]&~m[755]&m[756]&~m[758]&m[759])|(~m[734]&~m[755]&~m[756]&m[758]&m[759])|(m[734]&~m[755]&~m[756]&m[758]&m[759])|(~m[734]&m[755]&~m[756]&m[758]&m[759])|(m[734]&m[755]&~m[756]&m[758]&m[759])|(~m[734]&~m[755]&m[756]&m[758]&m[759])|(m[734]&~m[755]&m[756]&m[758]&m[759])|(m[734]&m[755]&m[756]&m[758]&m[759]))):InitCond[426];
    m[762] = run?((((m[744]&~m[760]&~m[761]&~m[763]&~m[764])|(~m[744]&~m[760]&~m[761]&m[763]&~m[764])|(m[744]&m[760]&~m[761]&m[763]&~m[764])|(m[744]&~m[760]&m[761]&m[763]&~m[764])|(~m[744]&m[760]&~m[761]&~m[763]&m[764])|(~m[744]&~m[760]&m[761]&~m[763]&m[764])|(m[744]&m[760]&m[761]&~m[763]&m[764])|(~m[744]&m[760]&m[761]&m[763]&m[764]))&UnbiasedRNG[188])|((m[744]&~m[760]&~m[761]&m[763]&~m[764])|(~m[744]&~m[760]&~m[761]&~m[763]&m[764])|(m[744]&~m[760]&~m[761]&~m[763]&m[764])|(m[744]&m[760]&~m[761]&~m[763]&m[764])|(m[744]&~m[760]&m[761]&~m[763]&m[764])|(~m[744]&~m[760]&~m[761]&m[763]&m[764])|(m[744]&~m[760]&~m[761]&m[763]&m[764])|(~m[744]&m[760]&~m[761]&m[763]&m[764])|(m[744]&m[760]&~m[761]&m[763]&m[764])|(~m[744]&~m[760]&m[761]&m[763]&m[764])|(m[744]&~m[760]&m[761]&m[763]&m[764])|(m[744]&m[760]&m[761]&m[763]&m[764]))):InitCond[427];
    m[767] = run?((((m[749]&~m[765]&~m[766]&~m[768]&~m[769])|(~m[749]&~m[765]&~m[766]&m[768]&~m[769])|(m[749]&m[765]&~m[766]&m[768]&~m[769])|(m[749]&~m[765]&m[766]&m[768]&~m[769])|(~m[749]&m[765]&~m[766]&~m[768]&m[769])|(~m[749]&~m[765]&m[766]&~m[768]&m[769])|(m[749]&m[765]&m[766]&~m[768]&m[769])|(~m[749]&m[765]&m[766]&m[768]&m[769]))&UnbiasedRNG[189])|((m[749]&~m[765]&~m[766]&m[768]&~m[769])|(~m[749]&~m[765]&~m[766]&~m[768]&m[769])|(m[749]&~m[765]&~m[766]&~m[768]&m[769])|(m[749]&m[765]&~m[766]&~m[768]&m[769])|(m[749]&~m[765]&m[766]&~m[768]&m[769])|(~m[749]&~m[765]&~m[766]&m[768]&m[769])|(m[749]&~m[765]&~m[766]&m[768]&m[769])|(~m[749]&m[765]&~m[766]&m[768]&m[769])|(m[749]&m[765]&~m[766]&m[768]&m[769])|(~m[749]&~m[765]&m[766]&m[768]&m[769])|(m[749]&~m[765]&m[766]&m[768]&m[769])|(m[749]&m[765]&m[766]&m[768]&m[769]))):InitCond[428];
    m[772] = run?((((m[754]&~m[770]&~m[771]&~m[773]&~m[774])|(~m[754]&~m[770]&~m[771]&m[773]&~m[774])|(m[754]&m[770]&~m[771]&m[773]&~m[774])|(m[754]&~m[770]&m[771]&m[773]&~m[774])|(~m[754]&m[770]&~m[771]&~m[773]&m[774])|(~m[754]&~m[770]&m[771]&~m[773]&m[774])|(m[754]&m[770]&m[771]&~m[773]&m[774])|(~m[754]&m[770]&m[771]&m[773]&m[774]))&UnbiasedRNG[190])|((m[754]&~m[770]&~m[771]&m[773]&~m[774])|(~m[754]&~m[770]&~m[771]&~m[773]&m[774])|(m[754]&~m[770]&~m[771]&~m[773]&m[774])|(m[754]&m[770]&~m[771]&~m[773]&m[774])|(m[754]&~m[770]&m[771]&~m[773]&m[774])|(~m[754]&~m[770]&~m[771]&m[773]&m[774])|(m[754]&~m[770]&~m[771]&m[773]&m[774])|(~m[754]&m[770]&~m[771]&m[773]&m[774])|(m[754]&m[770]&~m[771]&m[773]&m[774])|(~m[754]&~m[770]&m[771]&m[773]&m[774])|(m[754]&~m[770]&m[771]&m[773]&m[774])|(m[754]&m[770]&m[771]&m[773]&m[774]))):InitCond[429];
    m[777] = run?((((m[759]&~m[775]&~m[776]&~m[778]&~m[779])|(~m[759]&~m[775]&~m[776]&m[778]&~m[779])|(m[759]&m[775]&~m[776]&m[778]&~m[779])|(m[759]&~m[775]&m[776]&m[778]&~m[779])|(~m[759]&m[775]&~m[776]&~m[778]&m[779])|(~m[759]&~m[775]&m[776]&~m[778]&m[779])|(m[759]&m[775]&m[776]&~m[778]&m[779])|(~m[759]&m[775]&m[776]&m[778]&m[779]))&UnbiasedRNG[191])|((m[759]&~m[775]&~m[776]&m[778]&~m[779])|(~m[759]&~m[775]&~m[776]&~m[778]&m[779])|(m[759]&~m[775]&~m[776]&~m[778]&m[779])|(m[759]&m[775]&~m[776]&~m[778]&m[779])|(m[759]&~m[775]&m[776]&~m[778]&m[779])|(~m[759]&~m[775]&~m[776]&m[778]&m[779])|(m[759]&~m[775]&~m[776]&m[778]&m[779])|(~m[759]&m[775]&~m[776]&m[778]&m[779])|(m[759]&m[775]&~m[776]&m[778]&m[779])|(~m[759]&~m[775]&m[776]&m[778]&m[779])|(m[759]&~m[775]&m[776]&m[778]&m[779])|(m[759]&m[775]&m[776]&m[778]&m[779]))):InitCond[430];
    m[782] = run?((((m[769]&~m[780]&~m[781]&~m[783]&~m[784])|(~m[769]&~m[780]&~m[781]&m[783]&~m[784])|(m[769]&m[780]&~m[781]&m[783]&~m[784])|(m[769]&~m[780]&m[781]&m[783]&~m[784])|(~m[769]&m[780]&~m[781]&~m[783]&m[784])|(~m[769]&~m[780]&m[781]&~m[783]&m[784])|(m[769]&m[780]&m[781]&~m[783]&m[784])|(~m[769]&m[780]&m[781]&m[783]&m[784]))&UnbiasedRNG[192])|((m[769]&~m[780]&~m[781]&m[783]&~m[784])|(~m[769]&~m[780]&~m[781]&~m[783]&m[784])|(m[769]&~m[780]&~m[781]&~m[783]&m[784])|(m[769]&m[780]&~m[781]&~m[783]&m[784])|(m[769]&~m[780]&m[781]&~m[783]&m[784])|(~m[769]&~m[780]&~m[781]&m[783]&m[784])|(m[769]&~m[780]&~m[781]&m[783]&m[784])|(~m[769]&m[780]&~m[781]&m[783]&m[784])|(m[769]&m[780]&~m[781]&m[783]&m[784])|(~m[769]&~m[780]&m[781]&m[783]&m[784])|(m[769]&~m[780]&m[781]&m[783]&m[784])|(m[769]&m[780]&m[781]&m[783]&m[784]))):InitCond[431];
    m[787] = run?((((m[774]&~m[785]&~m[786]&~m[788]&~m[789])|(~m[774]&~m[785]&~m[786]&m[788]&~m[789])|(m[774]&m[785]&~m[786]&m[788]&~m[789])|(m[774]&~m[785]&m[786]&m[788]&~m[789])|(~m[774]&m[785]&~m[786]&~m[788]&m[789])|(~m[774]&~m[785]&m[786]&~m[788]&m[789])|(m[774]&m[785]&m[786]&~m[788]&m[789])|(~m[774]&m[785]&m[786]&m[788]&m[789]))&UnbiasedRNG[193])|((m[774]&~m[785]&~m[786]&m[788]&~m[789])|(~m[774]&~m[785]&~m[786]&~m[788]&m[789])|(m[774]&~m[785]&~m[786]&~m[788]&m[789])|(m[774]&m[785]&~m[786]&~m[788]&m[789])|(m[774]&~m[785]&m[786]&~m[788]&m[789])|(~m[774]&~m[785]&~m[786]&m[788]&m[789])|(m[774]&~m[785]&~m[786]&m[788]&m[789])|(~m[774]&m[785]&~m[786]&m[788]&m[789])|(m[774]&m[785]&~m[786]&m[788]&m[789])|(~m[774]&~m[785]&m[786]&m[788]&m[789])|(m[774]&~m[785]&m[786]&m[788]&m[789])|(m[774]&m[785]&m[786]&m[788]&m[789]))):InitCond[432];
    m[792] = run?((((m[779]&~m[790]&~m[791]&~m[793]&~m[794])|(~m[779]&~m[790]&~m[791]&m[793]&~m[794])|(m[779]&m[790]&~m[791]&m[793]&~m[794])|(m[779]&~m[790]&m[791]&m[793]&~m[794])|(~m[779]&m[790]&~m[791]&~m[793]&m[794])|(~m[779]&~m[790]&m[791]&~m[793]&m[794])|(m[779]&m[790]&m[791]&~m[793]&m[794])|(~m[779]&m[790]&m[791]&m[793]&m[794]))&UnbiasedRNG[194])|((m[779]&~m[790]&~m[791]&m[793]&~m[794])|(~m[779]&~m[790]&~m[791]&~m[793]&m[794])|(m[779]&~m[790]&~m[791]&~m[793]&m[794])|(m[779]&m[790]&~m[791]&~m[793]&m[794])|(m[779]&~m[790]&m[791]&~m[793]&m[794])|(~m[779]&~m[790]&~m[791]&m[793]&m[794])|(m[779]&~m[790]&~m[791]&m[793]&m[794])|(~m[779]&m[790]&~m[791]&m[793]&m[794])|(m[779]&m[790]&~m[791]&m[793]&m[794])|(~m[779]&~m[790]&m[791]&m[793]&m[794])|(m[779]&~m[790]&m[791]&m[793]&m[794])|(m[779]&m[790]&m[791]&m[793]&m[794]))):InitCond[433];
    m[797] = run?((((m[789]&~m[795]&~m[796]&~m[798]&~m[799])|(~m[789]&~m[795]&~m[796]&m[798]&~m[799])|(m[789]&m[795]&~m[796]&m[798]&~m[799])|(m[789]&~m[795]&m[796]&m[798]&~m[799])|(~m[789]&m[795]&~m[796]&~m[798]&m[799])|(~m[789]&~m[795]&m[796]&~m[798]&m[799])|(m[789]&m[795]&m[796]&~m[798]&m[799])|(~m[789]&m[795]&m[796]&m[798]&m[799]))&UnbiasedRNG[195])|((m[789]&~m[795]&~m[796]&m[798]&~m[799])|(~m[789]&~m[795]&~m[796]&~m[798]&m[799])|(m[789]&~m[795]&~m[796]&~m[798]&m[799])|(m[789]&m[795]&~m[796]&~m[798]&m[799])|(m[789]&~m[795]&m[796]&~m[798]&m[799])|(~m[789]&~m[795]&~m[796]&m[798]&m[799])|(m[789]&~m[795]&~m[796]&m[798]&m[799])|(~m[789]&m[795]&~m[796]&m[798]&m[799])|(m[789]&m[795]&~m[796]&m[798]&m[799])|(~m[789]&~m[795]&m[796]&m[798]&m[799])|(m[789]&~m[795]&m[796]&m[798]&m[799])|(m[789]&m[795]&m[796]&m[798]&m[799]))):InitCond[434];
    m[802] = run?((((m[794]&~m[800]&~m[801]&~m[803]&~m[804])|(~m[794]&~m[800]&~m[801]&m[803]&~m[804])|(m[794]&m[800]&~m[801]&m[803]&~m[804])|(m[794]&~m[800]&m[801]&m[803]&~m[804])|(~m[794]&m[800]&~m[801]&~m[803]&m[804])|(~m[794]&~m[800]&m[801]&~m[803]&m[804])|(m[794]&m[800]&m[801]&~m[803]&m[804])|(~m[794]&m[800]&m[801]&m[803]&m[804]))&UnbiasedRNG[196])|((m[794]&~m[800]&~m[801]&m[803]&~m[804])|(~m[794]&~m[800]&~m[801]&~m[803]&m[804])|(m[794]&~m[800]&~m[801]&~m[803]&m[804])|(m[794]&m[800]&~m[801]&~m[803]&m[804])|(m[794]&~m[800]&m[801]&~m[803]&m[804])|(~m[794]&~m[800]&~m[801]&m[803]&m[804])|(m[794]&~m[800]&~m[801]&m[803]&m[804])|(~m[794]&m[800]&~m[801]&m[803]&m[804])|(m[794]&m[800]&~m[801]&m[803]&m[804])|(~m[794]&~m[800]&m[801]&m[803]&m[804])|(m[794]&~m[800]&m[801]&m[803]&m[804])|(m[794]&m[800]&m[801]&m[803]&m[804]))):InitCond[435];
    m[807] = run?((((m[804]&~m[805]&~m[806]&~m[808]&~m[809])|(~m[804]&~m[805]&~m[806]&m[808]&~m[809])|(m[804]&m[805]&~m[806]&m[808]&~m[809])|(m[804]&~m[805]&m[806]&m[808]&~m[809])|(~m[804]&m[805]&~m[806]&~m[808]&m[809])|(~m[804]&~m[805]&m[806]&~m[808]&m[809])|(m[804]&m[805]&m[806]&~m[808]&m[809])|(~m[804]&m[805]&m[806]&m[808]&m[809]))&UnbiasedRNG[197])|((m[804]&~m[805]&~m[806]&m[808]&~m[809])|(~m[804]&~m[805]&~m[806]&~m[808]&m[809])|(m[804]&~m[805]&~m[806]&~m[808]&m[809])|(m[804]&m[805]&~m[806]&~m[808]&m[809])|(m[804]&~m[805]&m[806]&~m[808]&m[809])|(~m[804]&~m[805]&~m[806]&m[808]&m[809])|(m[804]&~m[805]&~m[806]&m[808]&m[809])|(~m[804]&m[805]&~m[806]&m[808]&m[809])|(m[804]&m[805]&~m[806]&m[808]&m[809])|(~m[804]&~m[805]&m[806]&m[808]&m[809])|(m[804]&~m[805]&m[806]&m[808]&m[809])|(m[804]&m[805]&m[806]&m[808]&m[809]))):InitCond[436];
end

always @(posedge color2_clk) begin
    m[160] = run?((((~m[10]&~m[60]&~m[260])|(m[10]&m[60]&~m[260]))&BiasedRNG[239])|(((m[10]&~m[60]&~m[260])|(~m[10]&m[60]&m[260]))&~BiasedRNG[239])|((~m[10]&~m[60]&m[260])|(m[10]&~m[60]&m[260])|(m[10]&m[60]&m[260]))):InitCond[437];
    m[161] = run?((((~m[10]&~m[70]&~m[261])|(m[10]&m[70]&~m[261]))&BiasedRNG[240])|(((m[10]&~m[70]&~m[261])|(~m[10]&m[70]&m[261]))&~BiasedRNG[240])|((~m[10]&~m[70]&m[261])|(m[10]&~m[70]&m[261])|(m[10]&m[70]&m[261]))):InitCond[438];
    m[170] = run?((((~m[11]&~m[61]&~m[270])|(m[11]&m[61]&~m[270]))&BiasedRNG[241])|(((m[11]&~m[61]&~m[270])|(~m[11]&m[61]&m[270]))&~BiasedRNG[241])|((~m[11]&~m[61]&m[270])|(m[11]&~m[61]&m[270])|(m[11]&m[61]&m[270]))):InitCond[439];
    m[171] = run?((((~m[11]&~m[71]&~m[271])|(m[11]&m[71]&~m[271]))&BiasedRNG[242])|(((m[11]&~m[71]&~m[271])|(~m[11]&m[71]&m[271]))&~BiasedRNG[242])|((~m[11]&~m[71]&m[271])|(m[11]&~m[71]&m[271])|(m[11]&m[71]&m[271]))):InitCond[440];
    m[182] = run?((((~m[44]&~m[82]&~m[282])|(m[44]&m[82]&~m[282]))&BiasedRNG[243])|(((m[44]&~m[82]&~m[282])|(~m[44]&m[82]&m[282]))&~BiasedRNG[243])|((~m[44]&~m[82]&m[282])|(m[44]&~m[82]&m[282])|(m[44]&m[82]&m[282]))):InitCond[441];
    m[183] = run?((((~m[44]&~m[92]&~m[283])|(m[44]&m[92]&~m[283]))&BiasedRNG[244])|(((m[44]&~m[92]&~m[283])|(~m[44]&m[92]&m[283]))&~BiasedRNG[244])|((~m[44]&~m[92]&m[283])|(m[44]&~m[92]&m[283])|(m[44]&m[92]&m[283]))):InitCond[442];
    m[184] = run?((((~m[44]&~m[102]&~m[284])|(m[44]&m[102]&~m[284]))&BiasedRNG[245])|(((m[44]&~m[102]&~m[284])|(~m[44]&m[102]&m[284]))&~BiasedRNG[245])|((~m[44]&~m[102]&m[284])|(m[44]&~m[102]&m[284])|(m[44]&m[102]&m[284]))):InitCond[443];
    m[185] = run?((((~m[44]&~m[112]&~m[285])|(m[44]&m[112]&~m[285]))&BiasedRNG[246])|(((m[44]&~m[112]&~m[285])|(~m[44]&m[112]&m[285]))&~BiasedRNG[246])|((~m[44]&~m[112]&m[285])|(m[44]&~m[112]&m[285])|(m[44]&m[112]&m[285]))):InitCond[444];
    m[186] = run?((((~m[45]&~m[122]&~m[286])|(m[45]&m[122]&~m[286]))&BiasedRNG[247])|(((m[45]&~m[122]&~m[286])|(~m[45]&m[122]&m[286]))&~BiasedRNG[247])|((~m[45]&~m[122]&m[286])|(m[45]&~m[122]&m[286])|(m[45]&m[122]&m[286]))):InitCond[445];
    m[187] = run?((((~m[45]&~m[132]&~m[287])|(m[45]&m[132]&~m[287]))&BiasedRNG[248])|(((m[45]&~m[132]&~m[287])|(~m[45]&m[132]&m[287]))&~BiasedRNG[248])|((~m[45]&~m[132]&m[287])|(m[45]&~m[132]&m[287])|(m[45]&m[132]&m[287]))):InitCond[446];
    m[188] = run?((((~m[45]&~m[142]&~m[288])|(m[45]&m[142]&~m[288]))&BiasedRNG[249])|(((m[45]&~m[142]&~m[288])|(~m[45]&m[142]&m[288]))&~BiasedRNG[249])|((~m[45]&~m[142]&m[288])|(m[45]&~m[142]&m[288])|(m[45]&m[142]&m[288]))):InitCond[447];
    m[189] = run?((((~m[45]&~m[152]&~m[289])|(m[45]&m[152]&~m[289]))&BiasedRNG[250])|(((m[45]&~m[152]&~m[289])|(~m[45]&m[152]&m[289]))&~BiasedRNG[250])|((~m[45]&~m[152]&m[289])|(m[45]&~m[152]&m[289])|(m[45]&m[152]&m[289]))):InitCond[448];
    m[192] = run?((((~m[46]&~m[83]&~m[292])|(m[46]&m[83]&~m[292]))&BiasedRNG[251])|(((m[46]&~m[83]&~m[292])|(~m[46]&m[83]&m[292]))&~BiasedRNG[251])|((~m[46]&~m[83]&m[292])|(m[46]&~m[83]&m[292])|(m[46]&m[83]&m[292]))):InitCond[449];
    m[193] = run?((((~m[46]&~m[93]&~m[293])|(m[46]&m[93]&~m[293]))&BiasedRNG[252])|(((m[46]&~m[93]&~m[293])|(~m[46]&m[93]&m[293]))&~BiasedRNG[252])|((~m[46]&~m[93]&m[293])|(m[46]&~m[93]&m[293])|(m[46]&m[93]&m[293]))):InitCond[450];
    m[194] = run?((((~m[46]&~m[103]&~m[294])|(m[46]&m[103]&~m[294]))&BiasedRNG[253])|(((m[46]&~m[103]&~m[294])|(~m[46]&m[103]&m[294]))&~BiasedRNG[253])|((~m[46]&~m[103]&m[294])|(m[46]&~m[103]&m[294])|(m[46]&m[103]&m[294]))):InitCond[451];
    m[195] = run?((((~m[46]&~m[113]&~m[295])|(m[46]&m[113]&~m[295]))&BiasedRNG[254])|(((m[46]&~m[113]&~m[295])|(~m[46]&m[113]&m[295]))&~BiasedRNG[254])|((~m[46]&~m[113]&m[295])|(m[46]&~m[113]&m[295])|(m[46]&m[113]&m[295]))):InitCond[452];
    m[196] = run?((((~m[47]&~m[123]&~m[296])|(m[47]&m[123]&~m[296]))&BiasedRNG[255])|(((m[47]&~m[123]&~m[296])|(~m[47]&m[123]&m[296]))&~BiasedRNG[255])|((~m[47]&~m[123]&m[296])|(m[47]&~m[123]&m[296])|(m[47]&m[123]&m[296]))):InitCond[453];
    m[197] = run?((((~m[47]&~m[133]&~m[297])|(m[47]&m[133]&~m[297]))&BiasedRNG[256])|(((m[47]&~m[133]&~m[297])|(~m[47]&m[133]&m[297]))&~BiasedRNG[256])|((~m[47]&~m[133]&m[297])|(m[47]&~m[133]&m[297])|(m[47]&m[133]&m[297]))):InitCond[454];
    m[198] = run?((((~m[47]&~m[143]&~m[298])|(m[47]&m[143]&~m[298]))&BiasedRNG[257])|(((m[47]&~m[143]&~m[298])|(~m[47]&m[143]&m[298]))&~BiasedRNG[257])|((~m[47]&~m[143]&m[298])|(m[47]&~m[143]&m[298])|(m[47]&m[143]&m[298]))):InitCond[455];
    m[199] = run?((((~m[47]&~m[153]&~m[299])|(m[47]&m[153]&~m[299]))&BiasedRNG[258])|(((m[47]&~m[153]&~m[299])|(~m[47]&m[153]&m[299]))&~BiasedRNG[258])|((~m[47]&~m[153]&m[299])|(m[47]&~m[153]&m[299])|(m[47]&m[153]&m[299]))):InitCond[456];
    m[202] = run?((((~m[48]&~m[84]&~m[302])|(m[48]&m[84]&~m[302]))&BiasedRNG[259])|(((m[48]&~m[84]&~m[302])|(~m[48]&m[84]&m[302]))&~BiasedRNG[259])|((~m[48]&~m[84]&m[302])|(m[48]&~m[84]&m[302])|(m[48]&m[84]&m[302]))):InitCond[457];
    m[203] = run?((((~m[48]&~m[94]&~m[303])|(m[48]&m[94]&~m[303]))&BiasedRNG[260])|(((m[48]&~m[94]&~m[303])|(~m[48]&m[94]&m[303]))&~BiasedRNG[260])|((~m[48]&~m[94]&m[303])|(m[48]&~m[94]&m[303])|(m[48]&m[94]&m[303]))):InitCond[458];
    m[204] = run?((((~m[48]&~m[104]&~m[304])|(m[48]&m[104]&~m[304]))&BiasedRNG[261])|(((m[48]&~m[104]&~m[304])|(~m[48]&m[104]&m[304]))&~BiasedRNG[261])|((~m[48]&~m[104]&m[304])|(m[48]&~m[104]&m[304])|(m[48]&m[104]&m[304]))):InitCond[459];
    m[205] = run?((((~m[48]&~m[114]&~m[305])|(m[48]&m[114]&~m[305]))&BiasedRNG[262])|(((m[48]&~m[114]&~m[305])|(~m[48]&m[114]&m[305]))&~BiasedRNG[262])|((~m[48]&~m[114]&m[305])|(m[48]&~m[114]&m[305])|(m[48]&m[114]&m[305]))):InitCond[460];
    m[206] = run?((((~m[49]&~m[124]&~m[306])|(m[49]&m[124]&~m[306]))&BiasedRNG[263])|(((m[49]&~m[124]&~m[306])|(~m[49]&m[124]&m[306]))&~BiasedRNG[263])|((~m[49]&~m[124]&m[306])|(m[49]&~m[124]&m[306])|(m[49]&m[124]&m[306]))):InitCond[461];
    m[207] = run?((((~m[49]&~m[134]&~m[307])|(m[49]&m[134]&~m[307]))&BiasedRNG[264])|(((m[49]&~m[134]&~m[307])|(~m[49]&m[134]&m[307]))&~BiasedRNG[264])|((~m[49]&~m[134]&m[307])|(m[49]&~m[134]&m[307])|(m[49]&m[134]&m[307]))):InitCond[462];
    m[208] = run?((((~m[49]&~m[144]&~m[308])|(m[49]&m[144]&~m[308]))&BiasedRNG[265])|(((m[49]&~m[144]&~m[308])|(~m[49]&m[144]&m[308]))&~BiasedRNG[265])|((~m[49]&~m[144]&m[308])|(m[49]&~m[144]&m[308])|(m[49]&m[144]&m[308]))):InitCond[463];
    m[209] = run?((((~m[49]&~m[154]&~m[309])|(m[49]&m[154]&~m[309]))&BiasedRNG[266])|(((m[49]&~m[154]&~m[309])|(~m[49]&m[154]&m[309]))&~BiasedRNG[266])|((~m[49]&~m[154]&m[309])|(m[49]&~m[154]&m[309])|(m[49]&m[154]&m[309]))):InitCond[464];
    m[212] = run?((((~m[50]&~m[85]&~m[312])|(m[50]&m[85]&~m[312]))&BiasedRNG[267])|(((m[50]&~m[85]&~m[312])|(~m[50]&m[85]&m[312]))&~BiasedRNG[267])|((~m[50]&~m[85]&m[312])|(m[50]&~m[85]&m[312])|(m[50]&m[85]&m[312]))):InitCond[465];
    m[213] = run?((((~m[50]&~m[95]&~m[313])|(m[50]&m[95]&~m[313]))&BiasedRNG[268])|(((m[50]&~m[95]&~m[313])|(~m[50]&m[95]&m[313]))&~BiasedRNG[268])|((~m[50]&~m[95]&m[313])|(m[50]&~m[95]&m[313])|(m[50]&m[95]&m[313]))):InitCond[466];
    m[214] = run?((((~m[50]&~m[105]&~m[314])|(m[50]&m[105]&~m[314]))&BiasedRNG[269])|(((m[50]&~m[105]&~m[314])|(~m[50]&m[105]&m[314]))&~BiasedRNG[269])|((~m[50]&~m[105]&m[314])|(m[50]&~m[105]&m[314])|(m[50]&m[105]&m[314]))):InitCond[467];
    m[215] = run?((((~m[50]&~m[115]&~m[315])|(m[50]&m[115]&~m[315]))&BiasedRNG[270])|(((m[50]&~m[115]&~m[315])|(~m[50]&m[115]&m[315]))&~BiasedRNG[270])|((~m[50]&~m[115]&m[315])|(m[50]&~m[115]&m[315])|(m[50]&m[115]&m[315]))):InitCond[468];
    m[216] = run?((((~m[51]&~m[125]&~m[316])|(m[51]&m[125]&~m[316]))&BiasedRNG[271])|(((m[51]&~m[125]&~m[316])|(~m[51]&m[125]&m[316]))&~BiasedRNG[271])|((~m[51]&~m[125]&m[316])|(m[51]&~m[125]&m[316])|(m[51]&m[125]&m[316]))):InitCond[469];
    m[217] = run?((((~m[51]&~m[135]&~m[317])|(m[51]&m[135]&~m[317]))&BiasedRNG[272])|(((m[51]&~m[135]&~m[317])|(~m[51]&m[135]&m[317]))&~BiasedRNG[272])|((~m[51]&~m[135]&m[317])|(m[51]&~m[135]&m[317])|(m[51]&m[135]&m[317]))):InitCond[470];
    m[218] = run?((((~m[51]&~m[145]&~m[318])|(m[51]&m[145]&~m[318]))&BiasedRNG[273])|(((m[51]&~m[145]&~m[318])|(~m[51]&m[145]&m[318]))&~BiasedRNG[273])|((~m[51]&~m[145]&m[318])|(m[51]&~m[145]&m[318])|(m[51]&m[145]&m[318]))):InitCond[471];
    m[219] = run?((((~m[51]&~m[155]&~m[319])|(m[51]&m[155]&~m[319]))&BiasedRNG[274])|(((m[51]&~m[155]&~m[319])|(~m[51]&m[155]&m[319]))&~BiasedRNG[274])|((~m[51]&~m[155]&m[319])|(m[51]&~m[155]&m[319])|(m[51]&m[155]&m[319]))):InitCond[472];
    m[222] = run?((((~m[52]&~m[86]&~m[322])|(m[52]&m[86]&~m[322]))&BiasedRNG[275])|(((m[52]&~m[86]&~m[322])|(~m[52]&m[86]&m[322]))&~BiasedRNG[275])|((~m[52]&~m[86]&m[322])|(m[52]&~m[86]&m[322])|(m[52]&m[86]&m[322]))):InitCond[473];
    m[223] = run?((((~m[52]&~m[96]&~m[323])|(m[52]&m[96]&~m[323]))&BiasedRNG[276])|(((m[52]&~m[96]&~m[323])|(~m[52]&m[96]&m[323]))&~BiasedRNG[276])|((~m[52]&~m[96]&m[323])|(m[52]&~m[96]&m[323])|(m[52]&m[96]&m[323]))):InitCond[474];
    m[224] = run?((((~m[52]&~m[106]&~m[324])|(m[52]&m[106]&~m[324]))&BiasedRNG[277])|(((m[52]&~m[106]&~m[324])|(~m[52]&m[106]&m[324]))&~BiasedRNG[277])|((~m[52]&~m[106]&m[324])|(m[52]&~m[106]&m[324])|(m[52]&m[106]&m[324]))):InitCond[475];
    m[225] = run?((((~m[52]&~m[116]&~m[325])|(m[52]&m[116]&~m[325]))&BiasedRNG[278])|(((m[52]&~m[116]&~m[325])|(~m[52]&m[116]&m[325]))&~BiasedRNG[278])|((~m[52]&~m[116]&m[325])|(m[52]&~m[116]&m[325])|(m[52]&m[116]&m[325]))):InitCond[476];
    m[226] = run?((((~m[53]&~m[126]&~m[326])|(m[53]&m[126]&~m[326]))&BiasedRNG[279])|(((m[53]&~m[126]&~m[326])|(~m[53]&m[126]&m[326]))&~BiasedRNG[279])|((~m[53]&~m[126]&m[326])|(m[53]&~m[126]&m[326])|(m[53]&m[126]&m[326]))):InitCond[477];
    m[227] = run?((((~m[53]&~m[136]&~m[327])|(m[53]&m[136]&~m[327]))&BiasedRNG[280])|(((m[53]&~m[136]&~m[327])|(~m[53]&m[136]&m[327]))&~BiasedRNG[280])|((~m[53]&~m[136]&m[327])|(m[53]&~m[136]&m[327])|(m[53]&m[136]&m[327]))):InitCond[478];
    m[228] = run?((((~m[53]&~m[146]&~m[328])|(m[53]&m[146]&~m[328]))&BiasedRNG[281])|(((m[53]&~m[146]&~m[328])|(~m[53]&m[146]&m[328]))&~BiasedRNG[281])|((~m[53]&~m[146]&m[328])|(m[53]&~m[146]&m[328])|(m[53]&m[146]&m[328]))):InitCond[479];
    m[229] = run?((((~m[53]&~m[156]&~m[329])|(m[53]&m[156]&~m[329]))&BiasedRNG[282])|(((m[53]&~m[156]&~m[329])|(~m[53]&m[156]&m[329]))&~BiasedRNG[282])|((~m[53]&~m[156]&m[329])|(m[53]&~m[156]&m[329])|(m[53]&m[156]&m[329]))):InitCond[480];
    m[232] = run?((((~m[54]&~m[87]&~m[332])|(m[54]&m[87]&~m[332]))&BiasedRNG[283])|(((m[54]&~m[87]&~m[332])|(~m[54]&m[87]&m[332]))&~BiasedRNG[283])|((~m[54]&~m[87]&m[332])|(m[54]&~m[87]&m[332])|(m[54]&m[87]&m[332]))):InitCond[481];
    m[233] = run?((((~m[54]&~m[97]&~m[333])|(m[54]&m[97]&~m[333]))&BiasedRNG[284])|(((m[54]&~m[97]&~m[333])|(~m[54]&m[97]&m[333]))&~BiasedRNG[284])|((~m[54]&~m[97]&m[333])|(m[54]&~m[97]&m[333])|(m[54]&m[97]&m[333]))):InitCond[482];
    m[234] = run?((((~m[54]&~m[107]&~m[334])|(m[54]&m[107]&~m[334]))&BiasedRNG[285])|(((m[54]&~m[107]&~m[334])|(~m[54]&m[107]&m[334]))&~BiasedRNG[285])|((~m[54]&~m[107]&m[334])|(m[54]&~m[107]&m[334])|(m[54]&m[107]&m[334]))):InitCond[483];
    m[235] = run?((((~m[54]&~m[117]&~m[335])|(m[54]&m[117]&~m[335]))&BiasedRNG[286])|(((m[54]&~m[117]&~m[335])|(~m[54]&m[117]&m[335]))&~BiasedRNG[286])|((~m[54]&~m[117]&m[335])|(m[54]&~m[117]&m[335])|(m[54]&m[117]&m[335]))):InitCond[484];
    m[236] = run?((((~m[55]&~m[127]&~m[336])|(m[55]&m[127]&~m[336]))&BiasedRNG[287])|(((m[55]&~m[127]&~m[336])|(~m[55]&m[127]&m[336]))&~BiasedRNG[287])|((~m[55]&~m[127]&m[336])|(m[55]&~m[127]&m[336])|(m[55]&m[127]&m[336]))):InitCond[485];
    m[237] = run?((((~m[55]&~m[137]&~m[337])|(m[55]&m[137]&~m[337]))&BiasedRNG[288])|(((m[55]&~m[137]&~m[337])|(~m[55]&m[137]&m[337]))&~BiasedRNG[288])|((~m[55]&~m[137]&m[337])|(m[55]&~m[137]&m[337])|(m[55]&m[137]&m[337]))):InitCond[486];
    m[238] = run?((((~m[55]&~m[147]&~m[338])|(m[55]&m[147]&~m[338]))&BiasedRNG[289])|(((m[55]&~m[147]&~m[338])|(~m[55]&m[147]&m[338]))&~BiasedRNG[289])|((~m[55]&~m[147]&m[338])|(m[55]&~m[147]&m[338])|(m[55]&m[147]&m[338]))):InitCond[487];
    m[239] = run?((((~m[55]&~m[157]&~m[339])|(m[55]&m[157]&~m[339]))&BiasedRNG[290])|(((m[55]&~m[157]&~m[339])|(~m[55]&m[157]&m[339]))&~BiasedRNG[290])|((~m[55]&~m[157]&m[339])|(m[55]&~m[157]&m[339])|(m[55]&m[157]&m[339]))):InitCond[488];
    m[242] = run?((((~m[56]&~m[88]&~m[342])|(m[56]&m[88]&~m[342]))&BiasedRNG[291])|(((m[56]&~m[88]&~m[342])|(~m[56]&m[88]&m[342]))&~BiasedRNG[291])|((~m[56]&~m[88]&m[342])|(m[56]&~m[88]&m[342])|(m[56]&m[88]&m[342]))):InitCond[489];
    m[243] = run?((((~m[56]&~m[98]&~m[343])|(m[56]&m[98]&~m[343]))&BiasedRNG[292])|(((m[56]&~m[98]&~m[343])|(~m[56]&m[98]&m[343]))&~BiasedRNG[292])|((~m[56]&~m[98]&m[343])|(m[56]&~m[98]&m[343])|(m[56]&m[98]&m[343]))):InitCond[490];
    m[244] = run?((((~m[56]&~m[108]&~m[344])|(m[56]&m[108]&~m[344]))&BiasedRNG[293])|(((m[56]&~m[108]&~m[344])|(~m[56]&m[108]&m[344]))&~BiasedRNG[293])|((~m[56]&~m[108]&m[344])|(m[56]&~m[108]&m[344])|(m[56]&m[108]&m[344]))):InitCond[491];
    m[245] = run?((((~m[56]&~m[118]&~m[345])|(m[56]&m[118]&~m[345]))&BiasedRNG[294])|(((m[56]&~m[118]&~m[345])|(~m[56]&m[118]&m[345]))&~BiasedRNG[294])|((~m[56]&~m[118]&m[345])|(m[56]&~m[118]&m[345])|(m[56]&m[118]&m[345]))):InitCond[492];
    m[246] = run?((((~m[57]&~m[128]&~m[346])|(m[57]&m[128]&~m[346]))&BiasedRNG[295])|(((m[57]&~m[128]&~m[346])|(~m[57]&m[128]&m[346]))&~BiasedRNG[295])|((~m[57]&~m[128]&m[346])|(m[57]&~m[128]&m[346])|(m[57]&m[128]&m[346]))):InitCond[493];
    m[247] = run?((((~m[57]&~m[138]&~m[347])|(m[57]&m[138]&~m[347]))&BiasedRNG[296])|(((m[57]&~m[138]&~m[347])|(~m[57]&m[138]&m[347]))&~BiasedRNG[296])|((~m[57]&~m[138]&m[347])|(m[57]&~m[138]&m[347])|(m[57]&m[138]&m[347]))):InitCond[494];
    m[248] = run?((((~m[57]&~m[148]&~m[348])|(m[57]&m[148]&~m[348]))&BiasedRNG[297])|(((m[57]&~m[148]&~m[348])|(~m[57]&m[148]&m[348]))&~BiasedRNG[297])|((~m[57]&~m[148]&m[348])|(m[57]&~m[148]&m[348])|(m[57]&m[148]&m[348]))):InitCond[495];
    m[249] = run?((((~m[57]&~m[158]&~m[349])|(m[57]&m[158]&~m[349]))&BiasedRNG[298])|(((m[57]&~m[158]&~m[349])|(~m[57]&m[158]&m[349]))&~BiasedRNG[298])|((~m[57]&~m[158]&m[349])|(m[57]&~m[158]&m[349])|(m[57]&m[158]&m[349]))):InitCond[496];
    m[252] = run?((((~m[58]&~m[89]&~m[352])|(m[58]&m[89]&~m[352]))&BiasedRNG[299])|(((m[58]&~m[89]&~m[352])|(~m[58]&m[89]&m[352]))&~BiasedRNG[299])|((~m[58]&~m[89]&m[352])|(m[58]&~m[89]&m[352])|(m[58]&m[89]&m[352]))):InitCond[497];
    m[253] = run?((((~m[58]&~m[99]&~m[353])|(m[58]&m[99]&~m[353]))&BiasedRNG[300])|(((m[58]&~m[99]&~m[353])|(~m[58]&m[99]&m[353]))&~BiasedRNG[300])|((~m[58]&~m[99]&m[353])|(m[58]&~m[99]&m[353])|(m[58]&m[99]&m[353]))):InitCond[498];
    m[254] = run?((((~m[58]&~m[109]&~m[354])|(m[58]&m[109]&~m[354]))&BiasedRNG[301])|(((m[58]&~m[109]&~m[354])|(~m[58]&m[109]&m[354]))&~BiasedRNG[301])|((~m[58]&~m[109]&m[354])|(m[58]&~m[109]&m[354])|(m[58]&m[109]&m[354]))):InitCond[499];
    m[255] = run?((((~m[58]&~m[119]&~m[355])|(m[58]&m[119]&~m[355]))&BiasedRNG[302])|(((m[58]&~m[119]&~m[355])|(~m[58]&m[119]&m[355]))&~BiasedRNG[302])|((~m[58]&~m[119]&m[355])|(m[58]&~m[119]&m[355])|(m[58]&m[119]&m[355]))):InitCond[500];
    m[256] = run?((((~m[59]&~m[129]&~m[356])|(m[59]&m[129]&~m[356]))&BiasedRNG[303])|(((m[59]&~m[129]&~m[356])|(~m[59]&m[129]&m[356]))&~BiasedRNG[303])|((~m[59]&~m[129]&m[356])|(m[59]&~m[129]&m[356])|(m[59]&m[129]&m[356]))):InitCond[501];
    m[257] = run?((((~m[59]&~m[139]&~m[357])|(m[59]&m[139]&~m[357]))&BiasedRNG[304])|(((m[59]&~m[139]&~m[357])|(~m[59]&m[139]&m[357]))&~BiasedRNG[304])|((~m[59]&~m[139]&m[357])|(m[59]&~m[139]&m[357])|(m[59]&m[139]&m[357]))):InitCond[502];
    m[258] = run?((((~m[59]&~m[149]&~m[358])|(m[59]&m[149]&~m[358]))&BiasedRNG[305])|(((m[59]&~m[149]&~m[358])|(~m[59]&m[149]&m[358]))&~BiasedRNG[305])|((~m[59]&~m[149]&m[358])|(m[59]&~m[149]&m[358])|(m[59]&m[149]&m[358]))):InitCond[503];
    m[259] = run?((((~m[59]&~m[159]&~m[359])|(m[59]&m[159]&~m[359]))&BiasedRNG[306])|(((m[59]&~m[159]&~m[359])|(~m[59]&m[159]&m[359]))&~BiasedRNG[306])|((~m[59]&~m[159]&m[359])|(m[59]&~m[159]&m[359])|(m[59]&m[159]&m[359]))):InitCond[504];
    m[262] = run?((((m[80]&~m[162]&m[365])|(~m[80]&m[162]&m[365]))&BiasedRNG[307])|(((m[80]&m[162]&~m[365]))&~BiasedRNG[307])|((m[80]&m[162]&m[365]))):InitCond[505];
    m[263] = run?((((m[90]&~m[163]&m[375])|(~m[90]&m[163]&m[375]))&BiasedRNG[308])|(((m[90]&m[163]&~m[375]))&~BiasedRNG[308])|((m[90]&m[163]&m[375]))):InitCond[506];
    m[264] = run?((((m[100]&~m[164]&m[390])|(~m[100]&m[164]&m[390]))&BiasedRNG[309])|(((m[100]&m[164]&~m[390]))&~BiasedRNG[309])|((m[100]&m[164]&m[390]))):InitCond[507];
    m[265] = run?((((m[110]&~m[165]&m[410])|(~m[110]&m[165]&m[410]))&BiasedRNG[310])|(((m[110]&m[165]&~m[410]))&~BiasedRNG[310])|((m[110]&m[165]&m[410]))):InitCond[508];
    m[266] = run?((((m[120]&~m[166]&m[435])|(~m[120]&m[166]&m[435]))&BiasedRNG[311])|(((m[120]&m[166]&~m[435]))&~BiasedRNG[311])|((m[120]&m[166]&m[435]))):InitCond[509];
    m[267] = run?((((m[130]&~m[167]&m[465])|(~m[130]&m[167]&m[465]))&BiasedRNG[312])|(((m[130]&m[167]&~m[465]))&~BiasedRNG[312])|((m[130]&m[167]&m[465]))):InitCond[510];
    m[268] = run?((((m[140]&~m[168]&m[500])|(~m[140]&m[168]&m[500]))&BiasedRNG[313])|(((m[140]&m[168]&~m[500]))&~BiasedRNG[313])|((m[140]&m[168]&m[500]))):InitCond[511];
    m[269] = run?((((m[150]&~m[169]&m[540])|(~m[150]&m[169]&m[540]))&BiasedRNG[314])|(((m[150]&m[169]&~m[540]))&~BiasedRNG[314])|((m[150]&m[169]&m[540]))):InitCond[512];
    m[272] = run?((((m[81]&~m[172]&m[376])|(~m[81]&m[172]&m[376]))&BiasedRNG[315])|(((m[81]&m[172]&~m[376]))&~BiasedRNG[315])|((m[81]&m[172]&m[376]))):InitCond[513];
    m[273] = run?((((m[91]&~m[173]&m[391])|(~m[91]&m[173]&m[391]))&BiasedRNG[316])|(((m[91]&m[173]&~m[391]))&~BiasedRNG[316])|((m[91]&m[173]&m[391]))):InitCond[514];
    m[274] = run?((((m[101]&~m[174]&m[411])|(~m[101]&m[174]&m[411]))&BiasedRNG[317])|(((m[101]&m[174]&~m[411]))&~BiasedRNG[317])|((m[101]&m[174]&m[411]))):InitCond[515];
    m[275] = run?((((m[111]&~m[175]&m[436])|(~m[111]&m[175]&m[436]))&BiasedRNG[318])|(((m[111]&m[175]&~m[436]))&~BiasedRNG[318])|((m[111]&m[175]&m[436]))):InitCond[516];
    m[276] = run?((((m[121]&~m[176]&m[466])|(~m[121]&m[176]&m[466]))&BiasedRNG[319])|(((m[121]&m[176]&~m[466]))&~BiasedRNG[319])|((m[121]&m[176]&m[466]))):InitCond[517];
    m[277] = run?((((m[131]&~m[177]&m[501])|(~m[131]&m[177]&m[501]))&BiasedRNG[320])|(((m[131]&m[177]&~m[501]))&~BiasedRNG[320])|((m[131]&m[177]&m[501]))):InitCond[518];
    m[278] = run?((((m[141]&~m[178]&m[541])|(~m[141]&m[178]&m[541]))&BiasedRNG[321])|(((m[141]&m[178]&~m[541]))&~BiasedRNG[321])|((m[141]&m[178]&m[541]))):InitCond[519];
    m[279] = run?((((m[151]&~m[179]&m[586])|(~m[151]&m[179]&m[586]))&BiasedRNG[322])|(((m[151]&m[179]&~m[586]))&~BiasedRNG[322])|((m[151]&m[179]&m[586]))):InitCond[520];
    m[280] = run?((((m[62]&~m[180]&m[371])|(~m[62]&m[180]&m[371]))&BiasedRNG[323])|(((m[62]&m[180]&~m[371]))&~BiasedRNG[323])|((m[62]&m[180]&m[371]))):InitCond[521];
    m[281] = run?((((m[72]&~m[181]&m[381])|(~m[72]&m[181]&m[381]))&BiasedRNG[324])|(((m[72]&m[181]&~m[381]))&~BiasedRNG[324])|((m[72]&m[181]&m[381]))):InitCond[522];
    m[290] = run?((((m[63]&~m[190]&m[386])|(~m[63]&m[190]&m[386]))&BiasedRNG[325])|(((m[63]&m[190]&~m[386]))&~BiasedRNG[325])|((m[63]&m[190]&m[386]))):InitCond[523];
    m[291] = run?((((m[73]&~m[191]&m[401])|(~m[73]&m[191]&m[401]))&BiasedRNG[326])|(((m[73]&m[191]&~m[401]))&~BiasedRNG[326])|((m[73]&m[191]&m[401]))):InitCond[524];
    m[300] = run?((((m[64]&~m[200]&m[406])|(~m[64]&m[200]&m[406]))&BiasedRNG[327])|(((m[64]&m[200]&~m[406]))&~BiasedRNG[327])|((m[64]&m[200]&m[406]))):InitCond[525];
    m[301] = run?((((m[74]&~m[201]&m[426])|(~m[74]&m[201]&m[426]))&BiasedRNG[328])|(((m[74]&m[201]&~m[426]))&~BiasedRNG[328])|((m[74]&m[201]&m[426]))):InitCond[526];
    m[310] = run?((((m[65]&~m[210]&m[431])|(~m[65]&m[210]&m[431]))&BiasedRNG[329])|(((m[65]&m[210]&~m[431]))&~BiasedRNG[329])|((m[65]&m[210]&m[431]))):InitCond[527];
    m[311] = run?((((m[75]&~m[211]&m[456])|(~m[75]&m[211]&m[456]))&BiasedRNG[330])|(((m[75]&m[211]&~m[456]))&~BiasedRNG[330])|((m[75]&m[211]&m[456]))):InitCond[528];
    m[320] = run?((((m[66]&~m[220]&m[461])|(~m[66]&m[220]&m[461]))&BiasedRNG[331])|(((m[66]&m[220]&~m[461]))&~BiasedRNG[331])|((m[66]&m[220]&m[461]))):InitCond[529];
    m[321] = run?((((m[76]&~m[221]&m[491])|(~m[76]&m[221]&m[491]))&BiasedRNG[332])|(((m[76]&m[221]&~m[491]))&~BiasedRNG[332])|((m[76]&m[221]&m[491]))):InitCond[530];
    m[330] = run?((((m[67]&~m[230]&m[496])|(~m[67]&m[230]&m[496]))&BiasedRNG[333])|(((m[67]&m[230]&~m[496]))&~BiasedRNG[333])|((m[67]&m[230]&m[496]))):InitCond[531];
    m[331] = run?((((m[77]&~m[231]&m[531])|(~m[77]&m[231]&m[531]))&BiasedRNG[334])|(((m[77]&m[231]&~m[531]))&~BiasedRNG[334])|((m[77]&m[231]&m[531]))):InitCond[532];
    m[340] = run?((((m[68]&~m[240]&m[536])|(~m[68]&m[240]&m[536]))&BiasedRNG[335])|(((m[68]&m[240]&~m[536]))&~BiasedRNG[335])|((m[68]&m[240]&m[536]))):InitCond[533];
    m[341] = run?((((m[78]&~m[241]&m[576])|(~m[78]&m[241]&m[576]))&BiasedRNG[336])|(((m[78]&m[241]&~m[576]))&~BiasedRNG[336])|((m[78]&m[241]&m[576]))):InitCond[534];
    m[350] = run?((((m[69]&~m[250]&m[581])|(~m[69]&m[250]&m[581]))&BiasedRNG[337])|(((m[69]&m[250]&~m[581]))&~BiasedRNG[337])|((m[69]&m[250]&m[581]))):InitCond[535];
    m[351] = run?((((m[79]&~m[251]&m[626])|(~m[79]&m[251]&m[626]))&BiasedRNG[338])|(((m[79]&m[251]&~m[626]))&~BiasedRNG[338])|((m[79]&m[251]&m[626]))):InitCond[536];
    m[361] = run?((((m[270]&~m[360]&~m[362]&~m[363]&~m[364])|(~m[270]&~m[360]&~m[362]&m[363]&~m[364])|(m[270]&m[360]&~m[362]&m[363]&~m[364])|(m[270]&~m[360]&m[362]&m[363]&~m[364])|(~m[270]&m[360]&~m[362]&~m[363]&m[364])|(~m[270]&~m[360]&m[362]&~m[363]&m[364])|(m[270]&m[360]&m[362]&~m[363]&m[364])|(~m[270]&m[360]&m[362]&m[363]&m[364]))&UnbiasedRNG[198])|((m[270]&~m[360]&~m[362]&m[363]&~m[364])|(~m[270]&~m[360]&~m[362]&~m[363]&m[364])|(m[270]&~m[360]&~m[362]&~m[363]&m[364])|(m[270]&m[360]&~m[362]&~m[363]&m[364])|(m[270]&~m[360]&m[362]&~m[363]&m[364])|(~m[270]&~m[360]&~m[362]&m[363]&m[364])|(m[270]&~m[360]&~m[362]&m[363]&m[364])|(~m[270]&m[360]&~m[362]&m[363]&m[364])|(m[270]&m[360]&~m[362]&m[363]&m[364])|(~m[270]&~m[360]&m[362]&m[363]&m[364])|(m[270]&~m[360]&m[362]&m[363]&m[364])|(m[270]&m[360]&m[362]&m[363]&m[364]))):InitCond[537];
    m[367] = run?((((m[364]&~m[365]&~m[366]&~m[368]&~m[369])|(~m[364]&~m[365]&~m[366]&m[368]&~m[369])|(m[364]&m[365]&~m[366]&m[368]&~m[369])|(m[364]&~m[365]&m[366]&m[368]&~m[369])|(~m[364]&m[365]&~m[366]&~m[368]&m[369])|(~m[364]&~m[365]&m[366]&~m[368]&m[369])|(m[364]&m[365]&m[366]&~m[368]&m[369])|(~m[364]&m[365]&m[366]&m[368]&m[369]))&UnbiasedRNG[199])|((m[364]&~m[365]&~m[366]&m[368]&~m[369])|(~m[364]&~m[365]&~m[366]&~m[368]&m[369])|(m[364]&~m[365]&~m[366]&~m[368]&m[369])|(m[364]&m[365]&~m[366]&~m[368]&m[369])|(m[364]&~m[365]&m[366]&~m[368]&m[369])|(~m[364]&~m[365]&~m[366]&m[368]&m[369])|(m[364]&~m[365]&~m[366]&m[368]&m[369])|(~m[364]&m[365]&~m[366]&m[368]&m[369])|(m[364]&m[365]&~m[366]&m[368]&m[369])|(~m[364]&~m[365]&m[366]&m[368]&m[369])|(m[364]&~m[365]&m[366]&m[368]&m[369])|(m[364]&m[365]&m[366]&m[368]&m[369]))):InitCond[538];
    m[377] = run?((((m[369]&~m[375]&~m[376]&~m[378]&~m[379])|(~m[369]&~m[375]&~m[376]&m[378]&~m[379])|(m[369]&m[375]&~m[376]&m[378]&~m[379])|(m[369]&~m[375]&m[376]&m[378]&~m[379])|(~m[369]&m[375]&~m[376]&~m[378]&m[379])|(~m[369]&~m[375]&m[376]&~m[378]&m[379])|(m[369]&m[375]&m[376]&~m[378]&m[379])|(~m[369]&m[375]&m[376]&m[378]&m[379]))&UnbiasedRNG[200])|((m[369]&~m[375]&~m[376]&m[378]&~m[379])|(~m[369]&~m[375]&~m[376]&~m[378]&m[379])|(m[369]&~m[375]&~m[376]&~m[378]&m[379])|(m[369]&m[375]&~m[376]&~m[378]&m[379])|(m[369]&~m[375]&m[376]&~m[378]&m[379])|(~m[369]&~m[375]&~m[376]&m[378]&m[379])|(m[369]&~m[375]&~m[376]&m[378]&m[379])|(~m[369]&m[375]&~m[376]&m[378]&m[379])|(m[369]&m[375]&~m[376]&m[378]&m[379])|(~m[369]&~m[375]&m[376]&m[378]&m[379])|(m[369]&~m[375]&m[376]&m[378]&m[379])|(m[369]&m[375]&m[376]&m[378]&m[379]))):InitCond[539];
    m[382] = run?((((m[374]&~m[380]&~m[381]&~m[383]&~m[384])|(~m[374]&~m[380]&~m[381]&m[383]&~m[384])|(m[374]&m[380]&~m[381]&m[383]&~m[384])|(m[374]&~m[380]&m[381]&m[383]&~m[384])|(~m[374]&m[380]&~m[381]&~m[383]&m[384])|(~m[374]&~m[380]&m[381]&~m[383]&m[384])|(m[374]&m[380]&m[381]&~m[383]&m[384])|(~m[374]&m[380]&m[381]&m[383]&m[384]))&UnbiasedRNG[201])|((m[374]&~m[380]&~m[381]&m[383]&~m[384])|(~m[374]&~m[380]&~m[381]&~m[383]&m[384])|(m[374]&~m[380]&~m[381]&~m[383]&m[384])|(m[374]&m[380]&~m[381]&~m[383]&m[384])|(m[374]&~m[380]&m[381]&~m[383]&m[384])|(~m[374]&~m[380]&~m[381]&m[383]&m[384])|(m[374]&~m[380]&~m[381]&m[383]&m[384])|(~m[374]&m[380]&~m[381]&m[383]&m[384])|(m[374]&m[380]&~m[381]&m[383]&m[384])|(~m[374]&~m[380]&m[381]&m[383]&m[384])|(m[374]&~m[380]&m[381]&m[383]&m[384])|(m[374]&m[380]&m[381]&m[383]&m[384]))):InitCond[540];
    m[392] = run?((((m[379]&~m[390]&~m[391]&~m[393]&~m[394])|(~m[379]&~m[390]&~m[391]&m[393]&~m[394])|(m[379]&m[390]&~m[391]&m[393]&~m[394])|(m[379]&~m[390]&m[391]&m[393]&~m[394])|(~m[379]&m[390]&~m[391]&~m[393]&m[394])|(~m[379]&~m[390]&m[391]&~m[393]&m[394])|(m[379]&m[390]&m[391]&~m[393]&m[394])|(~m[379]&m[390]&m[391]&m[393]&m[394]))&UnbiasedRNG[202])|((m[379]&~m[390]&~m[391]&m[393]&~m[394])|(~m[379]&~m[390]&~m[391]&~m[393]&m[394])|(m[379]&~m[390]&~m[391]&~m[393]&m[394])|(m[379]&m[390]&~m[391]&~m[393]&m[394])|(m[379]&~m[390]&m[391]&~m[393]&m[394])|(~m[379]&~m[390]&~m[391]&m[393]&m[394])|(m[379]&~m[390]&~m[391]&m[393]&m[394])|(~m[379]&m[390]&~m[391]&m[393]&m[394])|(m[379]&m[390]&~m[391]&m[393]&m[394])|(~m[379]&~m[390]&m[391]&m[393]&m[394])|(m[379]&~m[390]&m[391]&m[393]&m[394])|(m[379]&m[390]&m[391]&m[393]&m[394]))):InitCond[541];
    m[396] = run?((((m[282]&~m[395]&~m[397]&~m[398]&~m[399])|(~m[282]&~m[395]&~m[397]&m[398]&~m[399])|(m[282]&m[395]&~m[397]&m[398]&~m[399])|(m[282]&~m[395]&m[397]&m[398]&~m[399])|(~m[282]&m[395]&~m[397]&~m[398]&m[399])|(~m[282]&~m[395]&m[397]&~m[398]&m[399])|(m[282]&m[395]&m[397]&~m[398]&m[399])|(~m[282]&m[395]&m[397]&m[398]&m[399]))&UnbiasedRNG[203])|((m[282]&~m[395]&~m[397]&m[398]&~m[399])|(~m[282]&~m[395]&~m[397]&~m[398]&m[399])|(m[282]&~m[395]&~m[397]&~m[398]&m[399])|(m[282]&m[395]&~m[397]&~m[398]&m[399])|(m[282]&~m[395]&m[397]&~m[398]&m[399])|(~m[282]&~m[395]&~m[397]&m[398]&m[399])|(m[282]&~m[395]&~m[397]&m[398]&m[399])|(~m[282]&m[395]&~m[397]&m[398]&m[399])|(m[282]&m[395]&~m[397]&m[398]&m[399])|(~m[282]&~m[395]&m[397]&m[398]&m[399])|(m[282]&~m[395]&m[397]&m[398]&m[399])|(m[282]&m[395]&m[397]&m[398]&m[399]))):InitCond[542];
    m[402] = run?((((m[389]&~m[400]&~m[401]&~m[403]&~m[404])|(~m[389]&~m[400]&~m[401]&m[403]&~m[404])|(m[389]&m[400]&~m[401]&m[403]&~m[404])|(m[389]&~m[400]&m[401]&m[403]&~m[404])|(~m[389]&m[400]&~m[401]&~m[403]&m[404])|(~m[389]&~m[400]&m[401]&~m[403]&m[404])|(m[389]&m[400]&m[401]&~m[403]&m[404])|(~m[389]&m[400]&m[401]&m[403]&m[404]))&UnbiasedRNG[204])|((m[389]&~m[400]&~m[401]&m[403]&~m[404])|(~m[389]&~m[400]&~m[401]&~m[403]&m[404])|(m[389]&~m[400]&~m[401]&~m[403]&m[404])|(m[389]&m[400]&~m[401]&~m[403]&m[404])|(m[389]&~m[400]&m[401]&~m[403]&m[404])|(~m[389]&~m[400]&~m[401]&m[403]&m[404])|(m[389]&~m[400]&~m[401]&m[403]&m[404])|(~m[389]&m[400]&~m[401]&m[403]&m[404])|(m[389]&m[400]&~m[401]&m[403]&m[404])|(~m[389]&~m[400]&m[401]&m[403]&m[404])|(m[389]&~m[400]&m[401]&m[403]&m[404])|(m[389]&m[400]&m[401]&m[403]&m[404]))):InitCond[543];
    m[412] = run?((((m[394]&~m[410]&~m[411]&~m[413]&~m[414])|(~m[394]&~m[410]&~m[411]&m[413]&~m[414])|(m[394]&m[410]&~m[411]&m[413]&~m[414])|(m[394]&~m[410]&m[411]&m[413]&~m[414])|(~m[394]&m[410]&~m[411]&~m[413]&m[414])|(~m[394]&~m[410]&m[411]&~m[413]&m[414])|(m[394]&m[410]&m[411]&~m[413]&m[414])|(~m[394]&m[410]&m[411]&m[413]&m[414]))&UnbiasedRNG[205])|((m[394]&~m[410]&~m[411]&m[413]&~m[414])|(~m[394]&~m[410]&~m[411]&~m[413]&m[414])|(m[394]&~m[410]&~m[411]&~m[413]&m[414])|(m[394]&m[410]&~m[411]&~m[413]&m[414])|(m[394]&~m[410]&m[411]&~m[413]&m[414])|(~m[394]&~m[410]&~m[411]&m[413]&m[414])|(m[394]&~m[410]&~m[411]&m[413]&m[414])|(~m[394]&m[410]&~m[411]&m[413]&m[414])|(m[394]&m[410]&~m[411]&m[413]&m[414])|(~m[394]&~m[410]&m[411]&m[413]&m[414])|(m[394]&~m[410]&m[411]&m[413]&m[414])|(m[394]&m[410]&m[411]&m[413]&m[414]))):InitCond[544];
    m[416] = run?((((m[283]&~m[415]&~m[417]&~m[418]&~m[419])|(~m[283]&~m[415]&~m[417]&m[418]&~m[419])|(m[283]&m[415]&~m[417]&m[418]&~m[419])|(m[283]&~m[415]&m[417]&m[418]&~m[419])|(~m[283]&m[415]&~m[417]&~m[418]&m[419])|(~m[283]&~m[415]&m[417]&~m[418]&m[419])|(m[283]&m[415]&m[417]&~m[418]&m[419])|(~m[283]&m[415]&m[417]&m[418]&m[419]))&UnbiasedRNG[206])|((m[283]&~m[415]&~m[417]&m[418]&~m[419])|(~m[283]&~m[415]&~m[417]&~m[418]&m[419])|(m[283]&~m[415]&~m[417]&~m[418]&m[419])|(m[283]&m[415]&~m[417]&~m[418]&m[419])|(m[283]&~m[415]&m[417]&~m[418]&m[419])|(~m[283]&~m[415]&~m[417]&m[418]&m[419])|(m[283]&~m[415]&~m[417]&m[418]&m[419])|(~m[283]&m[415]&~m[417]&m[418]&m[419])|(m[283]&m[415]&~m[417]&m[418]&m[419])|(~m[283]&~m[415]&m[417]&m[418]&m[419])|(m[283]&~m[415]&m[417]&m[418]&m[419])|(m[283]&m[415]&m[417]&m[418]&m[419]))):InitCond[545];
    m[421] = run?((((m[292]&~m[420]&~m[422]&~m[423]&~m[424])|(~m[292]&~m[420]&~m[422]&m[423]&~m[424])|(m[292]&m[420]&~m[422]&m[423]&~m[424])|(m[292]&~m[420]&m[422]&m[423]&~m[424])|(~m[292]&m[420]&~m[422]&~m[423]&m[424])|(~m[292]&~m[420]&m[422]&~m[423]&m[424])|(m[292]&m[420]&m[422]&~m[423]&m[424])|(~m[292]&m[420]&m[422]&m[423]&m[424]))&UnbiasedRNG[207])|((m[292]&~m[420]&~m[422]&m[423]&~m[424])|(~m[292]&~m[420]&~m[422]&~m[423]&m[424])|(m[292]&~m[420]&~m[422]&~m[423]&m[424])|(m[292]&m[420]&~m[422]&~m[423]&m[424])|(m[292]&~m[420]&m[422]&~m[423]&m[424])|(~m[292]&~m[420]&~m[422]&m[423]&m[424])|(m[292]&~m[420]&~m[422]&m[423]&m[424])|(~m[292]&m[420]&~m[422]&m[423]&m[424])|(m[292]&m[420]&~m[422]&m[423]&m[424])|(~m[292]&~m[420]&m[422]&m[423]&m[424])|(m[292]&~m[420]&m[422]&m[423]&m[424])|(m[292]&m[420]&m[422]&m[423]&m[424]))):InitCond[546];
    m[427] = run?((((m[409]&~m[425]&~m[426]&~m[428]&~m[429])|(~m[409]&~m[425]&~m[426]&m[428]&~m[429])|(m[409]&m[425]&~m[426]&m[428]&~m[429])|(m[409]&~m[425]&m[426]&m[428]&~m[429])|(~m[409]&m[425]&~m[426]&~m[428]&m[429])|(~m[409]&~m[425]&m[426]&~m[428]&m[429])|(m[409]&m[425]&m[426]&~m[428]&m[429])|(~m[409]&m[425]&m[426]&m[428]&m[429]))&UnbiasedRNG[208])|((m[409]&~m[425]&~m[426]&m[428]&~m[429])|(~m[409]&~m[425]&~m[426]&~m[428]&m[429])|(m[409]&~m[425]&~m[426]&~m[428]&m[429])|(m[409]&m[425]&~m[426]&~m[428]&m[429])|(m[409]&~m[425]&m[426]&~m[428]&m[429])|(~m[409]&~m[425]&~m[426]&m[428]&m[429])|(m[409]&~m[425]&~m[426]&m[428]&m[429])|(~m[409]&m[425]&~m[426]&m[428]&m[429])|(m[409]&m[425]&~m[426]&m[428]&m[429])|(~m[409]&~m[425]&m[426]&m[428]&m[429])|(m[409]&~m[425]&m[426]&m[428]&m[429])|(m[409]&m[425]&m[426]&m[428]&m[429]))):InitCond[547];
    m[437] = run?((((m[414]&~m[435]&~m[436]&~m[438]&~m[439])|(~m[414]&~m[435]&~m[436]&m[438]&~m[439])|(m[414]&m[435]&~m[436]&m[438]&~m[439])|(m[414]&~m[435]&m[436]&m[438]&~m[439])|(~m[414]&m[435]&~m[436]&~m[438]&m[439])|(~m[414]&~m[435]&m[436]&~m[438]&m[439])|(m[414]&m[435]&m[436]&~m[438]&m[439])|(~m[414]&m[435]&m[436]&m[438]&m[439]))&UnbiasedRNG[209])|((m[414]&~m[435]&~m[436]&m[438]&~m[439])|(~m[414]&~m[435]&~m[436]&~m[438]&m[439])|(m[414]&~m[435]&~m[436]&~m[438]&m[439])|(m[414]&m[435]&~m[436]&~m[438]&m[439])|(m[414]&~m[435]&m[436]&~m[438]&m[439])|(~m[414]&~m[435]&~m[436]&m[438]&m[439])|(m[414]&~m[435]&~m[436]&m[438]&m[439])|(~m[414]&m[435]&~m[436]&m[438]&m[439])|(m[414]&m[435]&~m[436]&m[438]&m[439])|(~m[414]&~m[435]&m[436]&m[438]&m[439])|(m[414]&~m[435]&m[436]&m[438]&m[439])|(m[414]&m[435]&m[436]&m[438]&m[439]))):InitCond[548];
    m[441] = run?((((m[284]&~m[440]&~m[442]&~m[443]&~m[444])|(~m[284]&~m[440]&~m[442]&m[443]&~m[444])|(m[284]&m[440]&~m[442]&m[443]&~m[444])|(m[284]&~m[440]&m[442]&m[443]&~m[444])|(~m[284]&m[440]&~m[442]&~m[443]&m[444])|(~m[284]&~m[440]&m[442]&~m[443]&m[444])|(m[284]&m[440]&m[442]&~m[443]&m[444])|(~m[284]&m[440]&m[442]&m[443]&m[444]))&UnbiasedRNG[210])|((m[284]&~m[440]&~m[442]&m[443]&~m[444])|(~m[284]&~m[440]&~m[442]&~m[443]&m[444])|(m[284]&~m[440]&~m[442]&~m[443]&m[444])|(m[284]&m[440]&~m[442]&~m[443]&m[444])|(m[284]&~m[440]&m[442]&~m[443]&m[444])|(~m[284]&~m[440]&~m[442]&m[443]&m[444])|(m[284]&~m[440]&~m[442]&m[443]&m[444])|(~m[284]&m[440]&~m[442]&m[443]&m[444])|(m[284]&m[440]&~m[442]&m[443]&m[444])|(~m[284]&~m[440]&m[442]&m[443]&m[444])|(m[284]&~m[440]&m[442]&m[443]&m[444])|(m[284]&m[440]&m[442]&m[443]&m[444]))):InitCond[549];
    m[446] = run?((((m[293]&~m[445]&~m[447]&~m[448]&~m[449])|(~m[293]&~m[445]&~m[447]&m[448]&~m[449])|(m[293]&m[445]&~m[447]&m[448]&~m[449])|(m[293]&~m[445]&m[447]&m[448]&~m[449])|(~m[293]&m[445]&~m[447]&~m[448]&m[449])|(~m[293]&~m[445]&m[447]&~m[448]&m[449])|(m[293]&m[445]&m[447]&~m[448]&m[449])|(~m[293]&m[445]&m[447]&m[448]&m[449]))&UnbiasedRNG[211])|((m[293]&~m[445]&~m[447]&m[448]&~m[449])|(~m[293]&~m[445]&~m[447]&~m[448]&m[449])|(m[293]&~m[445]&~m[447]&~m[448]&m[449])|(m[293]&m[445]&~m[447]&~m[448]&m[449])|(m[293]&~m[445]&m[447]&~m[448]&m[449])|(~m[293]&~m[445]&~m[447]&m[448]&m[449])|(m[293]&~m[445]&~m[447]&m[448]&m[449])|(~m[293]&m[445]&~m[447]&m[448]&m[449])|(m[293]&m[445]&~m[447]&m[448]&m[449])|(~m[293]&~m[445]&m[447]&m[448]&m[449])|(m[293]&~m[445]&m[447]&m[448]&m[449])|(m[293]&m[445]&m[447]&m[448]&m[449]))):InitCond[550];
    m[451] = run?((((m[302]&~m[450]&~m[452]&~m[453]&~m[454])|(~m[302]&~m[450]&~m[452]&m[453]&~m[454])|(m[302]&m[450]&~m[452]&m[453]&~m[454])|(m[302]&~m[450]&m[452]&m[453]&~m[454])|(~m[302]&m[450]&~m[452]&~m[453]&m[454])|(~m[302]&~m[450]&m[452]&~m[453]&m[454])|(m[302]&m[450]&m[452]&~m[453]&m[454])|(~m[302]&m[450]&m[452]&m[453]&m[454]))&UnbiasedRNG[212])|((m[302]&~m[450]&~m[452]&m[453]&~m[454])|(~m[302]&~m[450]&~m[452]&~m[453]&m[454])|(m[302]&~m[450]&~m[452]&~m[453]&m[454])|(m[302]&m[450]&~m[452]&~m[453]&m[454])|(m[302]&~m[450]&m[452]&~m[453]&m[454])|(~m[302]&~m[450]&~m[452]&m[453]&m[454])|(m[302]&~m[450]&~m[452]&m[453]&m[454])|(~m[302]&m[450]&~m[452]&m[453]&m[454])|(m[302]&m[450]&~m[452]&m[453]&m[454])|(~m[302]&~m[450]&m[452]&m[453]&m[454])|(m[302]&~m[450]&m[452]&m[453]&m[454])|(m[302]&m[450]&m[452]&m[453]&m[454]))):InitCond[551];
    m[457] = run?((((m[434]&~m[455]&~m[456]&~m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&m[458]&~m[459])|(m[434]&m[455]&~m[456]&m[458]&~m[459])|(m[434]&~m[455]&m[456]&m[458]&~m[459])|(~m[434]&m[455]&~m[456]&~m[458]&m[459])|(~m[434]&~m[455]&m[456]&~m[458]&m[459])|(m[434]&m[455]&m[456]&~m[458]&m[459])|(~m[434]&m[455]&m[456]&m[458]&m[459]))&UnbiasedRNG[213])|((m[434]&~m[455]&~m[456]&m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&m[456]&~m[458]&m[459])|(~m[434]&~m[455]&~m[456]&m[458]&m[459])|(m[434]&~m[455]&~m[456]&m[458]&m[459])|(~m[434]&m[455]&~m[456]&m[458]&m[459])|(m[434]&m[455]&~m[456]&m[458]&m[459])|(~m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&m[455]&m[456]&m[458]&m[459]))):InitCond[552];
    m[467] = run?((((m[439]&~m[465]&~m[466]&~m[468]&~m[469])|(~m[439]&~m[465]&~m[466]&m[468]&~m[469])|(m[439]&m[465]&~m[466]&m[468]&~m[469])|(m[439]&~m[465]&m[466]&m[468]&~m[469])|(~m[439]&m[465]&~m[466]&~m[468]&m[469])|(~m[439]&~m[465]&m[466]&~m[468]&m[469])|(m[439]&m[465]&m[466]&~m[468]&m[469])|(~m[439]&m[465]&m[466]&m[468]&m[469]))&UnbiasedRNG[214])|((m[439]&~m[465]&~m[466]&m[468]&~m[469])|(~m[439]&~m[465]&~m[466]&~m[468]&m[469])|(m[439]&~m[465]&~m[466]&~m[468]&m[469])|(m[439]&m[465]&~m[466]&~m[468]&m[469])|(m[439]&~m[465]&m[466]&~m[468]&m[469])|(~m[439]&~m[465]&~m[466]&m[468]&m[469])|(m[439]&~m[465]&~m[466]&m[468]&m[469])|(~m[439]&m[465]&~m[466]&m[468]&m[469])|(m[439]&m[465]&~m[466]&m[468]&m[469])|(~m[439]&~m[465]&m[466]&m[468]&m[469])|(m[439]&~m[465]&m[466]&m[468]&m[469])|(m[439]&m[465]&m[466]&m[468]&m[469]))):InitCond[553];
    m[471] = run?((((m[285]&~m[470]&~m[472]&~m[473]&~m[474])|(~m[285]&~m[470]&~m[472]&m[473]&~m[474])|(m[285]&m[470]&~m[472]&m[473]&~m[474])|(m[285]&~m[470]&m[472]&m[473]&~m[474])|(~m[285]&m[470]&~m[472]&~m[473]&m[474])|(~m[285]&~m[470]&m[472]&~m[473]&m[474])|(m[285]&m[470]&m[472]&~m[473]&m[474])|(~m[285]&m[470]&m[472]&m[473]&m[474]))&UnbiasedRNG[215])|((m[285]&~m[470]&~m[472]&m[473]&~m[474])|(~m[285]&~m[470]&~m[472]&~m[473]&m[474])|(m[285]&~m[470]&~m[472]&~m[473]&m[474])|(m[285]&m[470]&~m[472]&~m[473]&m[474])|(m[285]&~m[470]&m[472]&~m[473]&m[474])|(~m[285]&~m[470]&~m[472]&m[473]&m[474])|(m[285]&~m[470]&~m[472]&m[473]&m[474])|(~m[285]&m[470]&~m[472]&m[473]&m[474])|(m[285]&m[470]&~m[472]&m[473]&m[474])|(~m[285]&~m[470]&m[472]&m[473]&m[474])|(m[285]&~m[470]&m[472]&m[473]&m[474])|(m[285]&m[470]&m[472]&m[473]&m[474]))):InitCond[554];
    m[476] = run?((((m[294]&~m[475]&~m[477]&~m[478]&~m[479])|(~m[294]&~m[475]&~m[477]&m[478]&~m[479])|(m[294]&m[475]&~m[477]&m[478]&~m[479])|(m[294]&~m[475]&m[477]&m[478]&~m[479])|(~m[294]&m[475]&~m[477]&~m[478]&m[479])|(~m[294]&~m[475]&m[477]&~m[478]&m[479])|(m[294]&m[475]&m[477]&~m[478]&m[479])|(~m[294]&m[475]&m[477]&m[478]&m[479]))&UnbiasedRNG[216])|((m[294]&~m[475]&~m[477]&m[478]&~m[479])|(~m[294]&~m[475]&~m[477]&~m[478]&m[479])|(m[294]&~m[475]&~m[477]&~m[478]&m[479])|(m[294]&m[475]&~m[477]&~m[478]&m[479])|(m[294]&~m[475]&m[477]&~m[478]&m[479])|(~m[294]&~m[475]&~m[477]&m[478]&m[479])|(m[294]&~m[475]&~m[477]&m[478]&m[479])|(~m[294]&m[475]&~m[477]&m[478]&m[479])|(m[294]&m[475]&~m[477]&m[478]&m[479])|(~m[294]&~m[475]&m[477]&m[478]&m[479])|(m[294]&~m[475]&m[477]&m[478]&m[479])|(m[294]&m[475]&m[477]&m[478]&m[479]))):InitCond[555];
    m[481] = run?((((m[303]&~m[480]&~m[482]&~m[483]&~m[484])|(~m[303]&~m[480]&~m[482]&m[483]&~m[484])|(m[303]&m[480]&~m[482]&m[483]&~m[484])|(m[303]&~m[480]&m[482]&m[483]&~m[484])|(~m[303]&m[480]&~m[482]&~m[483]&m[484])|(~m[303]&~m[480]&m[482]&~m[483]&m[484])|(m[303]&m[480]&m[482]&~m[483]&m[484])|(~m[303]&m[480]&m[482]&m[483]&m[484]))&UnbiasedRNG[217])|((m[303]&~m[480]&~m[482]&m[483]&~m[484])|(~m[303]&~m[480]&~m[482]&~m[483]&m[484])|(m[303]&~m[480]&~m[482]&~m[483]&m[484])|(m[303]&m[480]&~m[482]&~m[483]&m[484])|(m[303]&~m[480]&m[482]&~m[483]&m[484])|(~m[303]&~m[480]&~m[482]&m[483]&m[484])|(m[303]&~m[480]&~m[482]&m[483]&m[484])|(~m[303]&m[480]&~m[482]&m[483]&m[484])|(m[303]&m[480]&~m[482]&m[483]&m[484])|(~m[303]&~m[480]&m[482]&m[483]&m[484])|(m[303]&~m[480]&m[482]&m[483]&m[484])|(m[303]&m[480]&m[482]&m[483]&m[484]))):InitCond[556];
    m[486] = run?((((m[312]&~m[485]&~m[487]&~m[488]&~m[489])|(~m[312]&~m[485]&~m[487]&m[488]&~m[489])|(m[312]&m[485]&~m[487]&m[488]&~m[489])|(m[312]&~m[485]&m[487]&m[488]&~m[489])|(~m[312]&m[485]&~m[487]&~m[488]&m[489])|(~m[312]&~m[485]&m[487]&~m[488]&m[489])|(m[312]&m[485]&m[487]&~m[488]&m[489])|(~m[312]&m[485]&m[487]&m[488]&m[489]))&UnbiasedRNG[218])|((m[312]&~m[485]&~m[487]&m[488]&~m[489])|(~m[312]&~m[485]&~m[487]&~m[488]&m[489])|(m[312]&~m[485]&~m[487]&~m[488]&m[489])|(m[312]&m[485]&~m[487]&~m[488]&m[489])|(m[312]&~m[485]&m[487]&~m[488]&m[489])|(~m[312]&~m[485]&~m[487]&m[488]&m[489])|(m[312]&~m[485]&~m[487]&m[488]&m[489])|(~m[312]&m[485]&~m[487]&m[488]&m[489])|(m[312]&m[485]&~m[487]&m[488]&m[489])|(~m[312]&~m[485]&m[487]&m[488]&m[489])|(m[312]&~m[485]&m[487]&m[488]&m[489])|(m[312]&m[485]&m[487]&m[488]&m[489]))):InitCond[557];
    m[492] = run?((((m[464]&~m[490]&~m[491]&~m[493]&~m[494])|(~m[464]&~m[490]&~m[491]&m[493]&~m[494])|(m[464]&m[490]&~m[491]&m[493]&~m[494])|(m[464]&~m[490]&m[491]&m[493]&~m[494])|(~m[464]&m[490]&~m[491]&~m[493]&m[494])|(~m[464]&~m[490]&m[491]&~m[493]&m[494])|(m[464]&m[490]&m[491]&~m[493]&m[494])|(~m[464]&m[490]&m[491]&m[493]&m[494]))&UnbiasedRNG[219])|((m[464]&~m[490]&~m[491]&m[493]&~m[494])|(~m[464]&~m[490]&~m[491]&~m[493]&m[494])|(m[464]&~m[490]&~m[491]&~m[493]&m[494])|(m[464]&m[490]&~m[491]&~m[493]&m[494])|(m[464]&~m[490]&m[491]&~m[493]&m[494])|(~m[464]&~m[490]&~m[491]&m[493]&m[494])|(m[464]&~m[490]&~m[491]&m[493]&m[494])|(~m[464]&m[490]&~m[491]&m[493]&m[494])|(m[464]&m[490]&~m[491]&m[493]&m[494])|(~m[464]&~m[490]&m[491]&m[493]&m[494])|(m[464]&~m[490]&m[491]&m[493]&m[494])|(m[464]&m[490]&m[491]&m[493]&m[494]))):InitCond[558];
    m[502] = run?((((m[469]&~m[500]&~m[501]&~m[503]&~m[504])|(~m[469]&~m[500]&~m[501]&m[503]&~m[504])|(m[469]&m[500]&~m[501]&m[503]&~m[504])|(m[469]&~m[500]&m[501]&m[503]&~m[504])|(~m[469]&m[500]&~m[501]&~m[503]&m[504])|(~m[469]&~m[500]&m[501]&~m[503]&m[504])|(m[469]&m[500]&m[501]&~m[503]&m[504])|(~m[469]&m[500]&m[501]&m[503]&m[504]))&UnbiasedRNG[220])|((m[469]&~m[500]&~m[501]&m[503]&~m[504])|(~m[469]&~m[500]&~m[501]&~m[503]&m[504])|(m[469]&~m[500]&~m[501]&~m[503]&m[504])|(m[469]&m[500]&~m[501]&~m[503]&m[504])|(m[469]&~m[500]&m[501]&~m[503]&m[504])|(~m[469]&~m[500]&~m[501]&m[503]&m[504])|(m[469]&~m[500]&~m[501]&m[503]&m[504])|(~m[469]&m[500]&~m[501]&m[503]&m[504])|(m[469]&m[500]&~m[501]&m[503]&m[504])|(~m[469]&~m[500]&m[501]&m[503]&m[504])|(m[469]&~m[500]&m[501]&m[503]&m[504])|(m[469]&m[500]&m[501]&m[503]&m[504]))):InitCond[559];
    m[506] = run?((((m[286]&~m[505]&~m[507]&~m[508]&~m[509])|(~m[286]&~m[505]&~m[507]&m[508]&~m[509])|(m[286]&m[505]&~m[507]&m[508]&~m[509])|(m[286]&~m[505]&m[507]&m[508]&~m[509])|(~m[286]&m[505]&~m[507]&~m[508]&m[509])|(~m[286]&~m[505]&m[507]&~m[508]&m[509])|(m[286]&m[505]&m[507]&~m[508]&m[509])|(~m[286]&m[505]&m[507]&m[508]&m[509]))&UnbiasedRNG[221])|((m[286]&~m[505]&~m[507]&m[508]&~m[509])|(~m[286]&~m[505]&~m[507]&~m[508]&m[509])|(m[286]&~m[505]&~m[507]&~m[508]&m[509])|(m[286]&m[505]&~m[507]&~m[508]&m[509])|(m[286]&~m[505]&m[507]&~m[508]&m[509])|(~m[286]&~m[505]&~m[507]&m[508]&m[509])|(m[286]&~m[505]&~m[507]&m[508]&m[509])|(~m[286]&m[505]&~m[507]&m[508]&m[509])|(m[286]&m[505]&~m[507]&m[508]&m[509])|(~m[286]&~m[505]&m[507]&m[508]&m[509])|(m[286]&~m[505]&m[507]&m[508]&m[509])|(m[286]&m[505]&m[507]&m[508]&m[509]))):InitCond[560];
    m[511] = run?((((m[295]&~m[510]&~m[512]&~m[513]&~m[514])|(~m[295]&~m[510]&~m[512]&m[513]&~m[514])|(m[295]&m[510]&~m[512]&m[513]&~m[514])|(m[295]&~m[510]&m[512]&m[513]&~m[514])|(~m[295]&m[510]&~m[512]&~m[513]&m[514])|(~m[295]&~m[510]&m[512]&~m[513]&m[514])|(m[295]&m[510]&m[512]&~m[513]&m[514])|(~m[295]&m[510]&m[512]&m[513]&m[514]))&UnbiasedRNG[222])|((m[295]&~m[510]&~m[512]&m[513]&~m[514])|(~m[295]&~m[510]&~m[512]&~m[513]&m[514])|(m[295]&~m[510]&~m[512]&~m[513]&m[514])|(m[295]&m[510]&~m[512]&~m[513]&m[514])|(m[295]&~m[510]&m[512]&~m[513]&m[514])|(~m[295]&~m[510]&~m[512]&m[513]&m[514])|(m[295]&~m[510]&~m[512]&m[513]&m[514])|(~m[295]&m[510]&~m[512]&m[513]&m[514])|(m[295]&m[510]&~m[512]&m[513]&m[514])|(~m[295]&~m[510]&m[512]&m[513]&m[514])|(m[295]&~m[510]&m[512]&m[513]&m[514])|(m[295]&m[510]&m[512]&m[513]&m[514]))):InitCond[561];
    m[516] = run?((((m[304]&~m[515]&~m[517]&~m[518]&~m[519])|(~m[304]&~m[515]&~m[517]&m[518]&~m[519])|(m[304]&m[515]&~m[517]&m[518]&~m[519])|(m[304]&~m[515]&m[517]&m[518]&~m[519])|(~m[304]&m[515]&~m[517]&~m[518]&m[519])|(~m[304]&~m[515]&m[517]&~m[518]&m[519])|(m[304]&m[515]&m[517]&~m[518]&m[519])|(~m[304]&m[515]&m[517]&m[518]&m[519]))&UnbiasedRNG[223])|((m[304]&~m[515]&~m[517]&m[518]&~m[519])|(~m[304]&~m[515]&~m[517]&~m[518]&m[519])|(m[304]&~m[515]&~m[517]&~m[518]&m[519])|(m[304]&m[515]&~m[517]&~m[518]&m[519])|(m[304]&~m[515]&m[517]&~m[518]&m[519])|(~m[304]&~m[515]&~m[517]&m[518]&m[519])|(m[304]&~m[515]&~m[517]&m[518]&m[519])|(~m[304]&m[515]&~m[517]&m[518]&m[519])|(m[304]&m[515]&~m[517]&m[518]&m[519])|(~m[304]&~m[515]&m[517]&m[518]&m[519])|(m[304]&~m[515]&m[517]&m[518]&m[519])|(m[304]&m[515]&m[517]&m[518]&m[519]))):InitCond[562];
    m[521] = run?((((m[313]&~m[520]&~m[522]&~m[523]&~m[524])|(~m[313]&~m[520]&~m[522]&m[523]&~m[524])|(m[313]&m[520]&~m[522]&m[523]&~m[524])|(m[313]&~m[520]&m[522]&m[523]&~m[524])|(~m[313]&m[520]&~m[522]&~m[523]&m[524])|(~m[313]&~m[520]&m[522]&~m[523]&m[524])|(m[313]&m[520]&m[522]&~m[523]&m[524])|(~m[313]&m[520]&m[522]&m[523]&m[524]))&UnbiasedRNG[224])|((m[313]&~m[520]&~m[522]&m[523]&~m[524])|(~m[313]&~m[520]&~m[522]&~m[523]&m[524])|(m[313]&~m[520]&~m[522]&~m[523]&m[524])|(m[313]&m[520]&~m[522]&~m[523]&m[524])|(m[313]&~m[520]&m[522]&~m[523]&m[524])|(~m[313]&~m[520]&~m[522]&m[523]&m[524])|(m[313]&~m[520]&~m[522]&m[523]&m[524])|(~m[313]&m[520]&~m[522]&m[523]&m[524])|(m[313]&m[520]&~m[522]&m[523]&m[524])|(~m[313]&~m[520]&m[522]&m[523]&m[524])|(m[313]&~m[520]&m[522]&m[523]&m[524])|(m[313]&m[520]&m[522]&m[523]&m[524]))):InitCond[563];
    m[526] = run?((((m[322]&~m[525]&~m[527]&~m[528]&~m[529])|(~m[322]&~m[525]&~m[527]&m[528]&~m[529])|(m[322]&m[525]&~m[527]&m[528]&~m[529])|(m[322]&~m[525]&m[527]&m[528]&~m[529])|(~m[322]&m[525]&~m[527]&~m[528]&m[529])|(~m[322]&~m[525]&m[527]&~m[528]&m[529])|(m[322]&m[525]&m[527]&~m[528]&m[529])|(~m[322]&m[525]&m[527]&m[528]&m[529]))&UnbiasedRNG[225])|((m[322]&~m[525]&~m[527]&m[528]&~m[529])|(~m[322]&~m[525]&~m[527]&~m[528]&m[529])|(m[322]&~m[525]&~m[527]&~m[528]&m[529])|(m[322]&m[525]&~m[527]&~m[528]&m[529])|(m[322]&~m[525]&m[527]&~m[528]&m[529])|(~m[322]&~m[525]&~m[527]&m[528]&m[529])|(m[322]&~m[525]&~m[527]&m[528]&m[529])|(~m[322]&m[525]&~m[527]&m[528]&m[529])|(m[322]&m[525]&~m[527]&m[528]&m[529])|(~m[322]&~m[525]&m[527]&m[528]&m[529])|(m[322]&~m[525]&m[527]&m[528]&m[529])|(m[322]&m[525]&m[527]&m[528]&m[529]))):InitCond[564];
    m[532] = run?((((m[499]&~m[530]&~m[531]&~m[533]&~m[534])|(~m[499]&~m[530]&~m[531]&m[533]&~m[534])|(m[499]&m[530]&~m[531]&m[533]&~m[534])|(m[499]&~m[530]&m[531]&m[533]&~m[534])|(~m[499]&m[530]&~m[531]&~m[533]&m[534])|(~m[499]&~m[530]&m[531]&~m[533]&m[534])|(m[499]&m[530]&m[531]&~m[533]&m[534])|(~m[499]&m[530]&m[531]&m[533]&m[534]))&UnbiasedRNG[226])|((m[499]&~m[530]&~m[531]&m[533]&~m[534])|(~m[499]&~m[530]&~m[531]&~m[533]&m[534])|(m[499]&~m[530]&~m[531]&~m[533]&m[534])|(m[499]&m[530]&~m[531]&~m[533]&m[534])|(m[499]&~m[530]&m[531]&~m[533]&m[534])|(~m[499]&~m[530]&~m[531]&m[533]&m[534])|(m[499]&~m[530]&~m[531]&m[533]&m[534])|(~m[499]&m[530]&~m[531]&m[533]&m[534])|(m[499]&m[530]&~m[531]&m[533]&m[534])|(~m[499]&~m[530]&m[531]&m[533]&m[534])|(m[499]&~m[530]&m[531]&m[533]&m[534])|(m[499]&m[530]&m[531]&m[533]&m[534]))):InitCond[565];
    m[542] = run?((((m[504]&~m[540]&~m[541]&~m[543]&~m[544])|(~m[504]&~m[540]&~m[541]&m[543]&~m[544])|(m[504]&m[540]&~m[541]&m[543]&~m[544])|(m[504]&~m[540]&m[541]&m[543]&~m[544])|(~m[504]&m[540]&~m[541]&~m[543]&m[544])|(~m[504]&~m[540]&m[541]&~m[543]&m[544])|(m[504]&m[540]&m[541]&~m[543]&m[544])|(~m[504]&m[540]&m[541]&m[543]&m[544]))&UnbiasedRNG[227])|((m[504]&~m[540]&~m[541]&m[543]&~m[544])|(~m[504]&~m[540]&~m[541]&~m[543]&m[544])|(m[504]&~m[540]&~m[541]&~m[543]&m[544])|(m[504]&m[540]&~m[541]&~m[543]&m[544])|(m[504]&~m[540]&m[541]&~m[543]&m[544])|(~m[504]&~m[540]&~m[541]&m[543]&m[544])|(m[504]&~m[540]&~m[541]&m[543]&m[544])|(~m[504]&m[540]&~m[541]&m[543]&m[544])|(m[504]&m[540]&~m[541]&m[543]&m[544])|(~m[504]&~m[540]&m[541]&m[543]&m[544])|(m[504]&~m[540]&m[541]&m[543]&m[544])|(m[504]&m[540]&m[541]&m[543]&m[544]))):InitCond[566];
    m[546] = run?((((m[287]&~m[545]&~m[547]&~m[548]&~m[549])|(~m[287]&~m[545]&~m[547]&m[548]&~m[549])|(m[287]&m[545]&~m[547]&m[548]&~m[549])|(m[287]&~m[545]&m[547]&m[548]&~m[549])|(~m[287]&m[545]&~m[547]&~m[548]&m[549])|(~m[287]&~m[545]&m[547]&~m[548]&m[549])|(m[287]&m[545]&m[547]&~m[548]&m[549])|(~m[287]&m[545]&m[547]&m[548]&m[549]))&UnbiasedRNG[228])|((m[287]&~m[545]&~m[547]&m[548]&~m[549])|(~m[287]&~m[545]&~m[547]&~m[548]&m[549])|(m[287]&~m[545]&~m[547]&~m[548]&m[549])|(m[287]&m[545]&~m[547]&~m[548]&m[549])|(m[287]&~m[545]&m[547]&~m[548]&m[549])|(~m[287]&~m[545]&~m[547]&m[548]&m[549])|(m[287]&~m[545]&~m[547]&m[548]&m[549])|(~m[287]&m[545]&~m[547]&m[548]&m[549])|(m[287]&m[545]&~m[547]&m[548]&m[549])|(~m[287]&~m[545]&m[547]&m[548]&m[549])|(m[287]&~m[545]&m[547]&m[548]&m[549])|(m[287]&m[545]&m[547]&m[548]&m[549]))):InitCond[567];
    m[551] = run?((((m[296]&~m[550]&~m[552]&~m[553]&~m[554])|(~m[296]&~m[550]&~m[552]&m[553]&~m[554])|(m[296]&m[550]&~m[552]&m[553]&~m[554])|(m[296]&~m[550]&m[552]&m[553]&~m[554])|(~m[296]&m[550]&~m[552]&~m[553]&m[554])|(~m[296]&~m[550]&m[552]&~m[553]&m[554])|(m[296]&m[550]&m[552]&~m[553]&m[554])|(~m[296]&m[550]&m[552]&m[553]&m[554]))&UnbiasedRNG[229])|((m[296]&~m[550]&~m[552]&m[553]&~m[554])|(~m[296]&~m[550]&~m[552]&~m[553]&m[554])|(m[296]&~m[550]&~m[552]&~m[553]&m[554])|(m[296]&m[550]&~m[552]&~m[553]&m[554])|(m[296]&~m[550]&m[552]&~m[553]&m[554])|(~m[296]&~m[550]&~m[552]&m[553]&m[554])|(m[296]&~m[550]&~m[552]&m[553]&m[554])|(~m[296]&m[550]&~m[552]&m[553]&m[554])|(m[296]&m[550]&~m[552]&m[553]&m[554])|(~m[296]&~m[550]&m[552]&m[553]&m[554])|(m[296]&~m[550]&m[552]&m[553]&m[554])|(m[296]&m[550]&m[552]&m[553]&m[554]))):InitCond[568];
    m[556] = run?((((m[305]&~m[555]&~m[557]&~m[558]&~m[559])|(~m[305]&~m[555]&~m[557]&m[558]&~m[559])|(m[305]&m[555]&~m[557]&m[558]&~m[559])|(m[305]&~m[555]&m[557]&m[558]&~m[559])|(~m[305]&m[555]&~m[557]&~m[558]&m[559])|(~m[305]&~m[555]&m[557]&~m[558]&m[559])|(m[305]&m[555]&m[557]&~m[558]&m[559])|(~m[305]&m[555]&m[557]&m[558]&m[559]))&UnbiasedRNG[230])|((m[305]&~m[555]&~m[557]&m[558]&~m[559])|(~m[305]&~m[555]&~m[557]&~m[558]&m[559])|(m[305]&~m[555]&~m[557]&~m[558]&m[559])|(m[305]&m[555]&~m[557]&~m[558]&m[559])|(m[305]&~m[555]&m[557]&~m[558]&m[559])|(~m[305]&~m[555]&~m[557]&m[558]&m[559])|(m[305]&~m[555]&~m[557]&m[558]&m[559])|(~m[305]&m[555]&~m[557]&m[558]&m[559])|(m[305]&m[555]&~m[557]&m[558]&m[559])|(~m[305]&~m[555]&m[557]&m[558]&m[559])|(m[305]&~m[555]&m[557]&m[558]&m[559])|(m[305]&m[555]&m[557]&m[558]&m[559]))):InitCond[569];
    m[561] = run?((((m[314]&~m[560]&~m[562]&~m[563]&~m[564])|(~m[314]&~m[560]&~m[562]&m[563]&~m[564])|(m[314]&m[560]&~m[562]&m[563]&~m[564])|(m[314]&~m[560]&m[562]&m[563]&~m[564])|(~m[314]&m[560]&~m[562]&~m[563]&m[564])|(~m[314]&~m[560]&m[562]&~m[563]&m[564])|(m[314]&m[560]&m[562]&~m[563]&m[564])|(~m[314]&m[560]&m[562]&m[563]&m[564]))&UnbiasedRNG[231])|((m[314]&~m[560]&~m[562]&m[563]&~m[564])|(~m[314]&~m[560]&~m[562]&~m[563]&m[564])|(m[314]&~m[560]&~m[562]&~m[563]&m[564])|(m[314]&m[560]&~m[562]&~m[563]&m[564])|(m[314]&~m[560]&m[562]&~m[563]&m[564])|(~m[314]&~m[560]&~m[562]&m[563]&m[564])|(m[314]&~m[560]&~m[562]&m[563]&m[564])|(~m[314]&m[560]&~m[562]&m[563]&m[564])|(m[314]&m[560]&~m[562]&m[563]&m[564])|(~m[314]&~m[560]&m[562]&m[563]&m[564])|(m[314]&~m[560]&m[562]&m[563]&m[564])|(m[314]&m[560]&m[562]&m[563]&m[564]))):InitCond[570];
    m[566] = run?((((m[323]&~m[565]&~m[567]&~m[568]&~m[569])|(~m[323]&~m[565]&~m[567]&m[568]&~m[569])|(m[323]&m[565]&~m[567]&m[568]&~m[569])|(m[323]&~m[565]&m[567]&m[568]&~m[569])|(~m[323]&m[565]&~m[567]&~m[568]&m[569])|(~m[323]&~m[565]&m[567]&~m[568]&m[569])|(m[323]&m[565]&m[567]&~m[568]&m[569])|(~m[323]&m[565]&m[567]&m[568]&m[569]))&UnbiasedRNG[232])|((m[323]&~m[565]&~m[567]&m[568]&~m[569])|(~m[323]&~m[565]&~m[567]&~m[568]&m[569])|(m[323]&~m[565]&~m[567]&~m[568]&m[569])|(m[323]&m[565]&~m[567]&~m[568]&m[569])|(m[323]&~m[565]&m[567]&~m[568]&m[569])|(~m[323]&~m[565]&~m[567]&m[568]&m[569])|(m[323]&~m[565]&~m[567]&m[568]&m[569])|(~m[323]&m[565]&~m[567]&m[568]&m[569])|(m[323]&m[565]&~m[567]&m[568]&m[569])|(~m[323]&~m[565]&m[567]&m[568]&m[569])|(m[323]&~m[565]&m[567]&m[568]&m[569])|(m[323]&m[565]&m[567]&m[568]&m[569]))):InitCond[571];
    m[571] = run?((((m[332]&~m[570]&~m[572]&~m[573]&~m[574])|(~m[332]&~m[570]&~m[572]&m[573]&~m[574])|(m[332]&m[570]&~m[572]&m[573]&~m[574])|(m[332]&~m[570]&m[572]&m[573]&~m[574])|(~m[332]&m[570]&~m[572]&~m[573]&m[574])|(~m[332]&~m[570]&m[572]&~m[573]&m[574])|(m[332]&m[570]&m[572]&~m[573]&m[574])|(~m[332]&m[570]&m[572]&m[573]&m[574]))&UnbiasedRNG[233])|((m[332]&~m[570]&~m[572]&m[573]&~m[574])|(~m[332]&~m[570]&~m[572]&~m[573]&m[574])|(m[332]&~m[570]&~m[572]&~m[573]&m[574])|(m[332]&m[570]&~m[572]&~m[573]&m[574])|(m[332]&~m[570]&m[572]&~m[573]&m[574])|(~m[332]&~m[570]&~m[572]&m[573]&m[574])|(m[332]&~m[570]&~m[572]&m[573]&m[574])|(~m[332]&m[570]&~m[572]&m[573]&m[574])|(m[332]&m[570]&~m[572]&m[573]&m[574])|(~m[332]&~m[570]&m[572]&m[573]&m[574])|(m[332]&~m[570]&m[572]&m[573]&m[574])|(m[332]&m[570]&m[572]&m[573]&m[574]))):InitCond[572];
    m[577] = run?((((m[539]&~m[575]&~m[576]&~m[578]&~m[579])|(~m[539]&~m[575]&~m[576]&m[578]&~m[579])|(m[539]&m[575]&~m[576]&m[578]&~m[579])|(m[539]&~m[575]&m[576]&m[578]&~m[579])|(~m[539]&m[575]&~m[576]&~m[578]&m[579])|(~m[539]&~m[575]&m[576]&~m[578]&m[579])|(m[539]&m[575]&m[576]&~m[578]&m[579])|(~m[539]&m[575]&m[576]&m[578]&m[579]))&UnbiasedRNG[234])|((m[539]&~m[575]&~m[576]&m[578]&~m[579])|(~m[539]&~m[575]&~m[576]&~m[578]&m[579])|(m[539]&~m[575]&~m[576]&~m[578]&m[579])|(m[539]&m[575]&~m[576]&~m[578]&m[579])|(m[539]&~m[575]&m[576]&~m[578]&m[579])|(~m[539]&~m[575]&~m[576]&m[578]&m[579])|(m[539]&~m[575]&~m[576]&m[578]&m[579])|(~m[539]&m[575]&~m[576]&m[578]&m[579])|(m[539]&m[575]&~m[576]&m[578]&m[579])|(~m[539]&~m[575]&m[576]&m[578]&m[579])|(m[539]&~m[575]&m[576]&m[578]&m[579])|(m[539]&m[575]&m[576]&m[578]&m[579]))):InitCond[573];
    m[587] = run?((((m[544]&~m[585]&~m[586]&~m[588]&~m[589])|(~m[544]&~m[585]&~m[586]&m[588]&~m[589])|(m[544]&m[585]&~m[586]&m[588]&~m[589])|(m[544]&~m[585]&m[586]&m[588]&~m[589])|(~m[544]&m[585]&~m[586]&~m[588]&m[589])|(~m[544]&~m[585]&m[586]&~m[588]&m[589])|(m[544]&m[585]&m[586]&~m[588]&m[589])|(~m[544]&m[585]&m[586]&m[588]&m[589]))&UnbiasedRNG[235])|((m[544]&~m[585]&~m[586]&m[588]&~m[589])|(~m[544]&~m[585]&~m[586]&~m[588]&m[589])|(m[544]&~m[585]&~m[586]&~m[588]&m[589])|(m[544]&m[585]&~m[586]&~m[588]&m[589])|(m[544]&~m[585]&m[586]&~m[588]&m[589])|(~m[544]&~m[585]&~m[586]&m[588]&m[589])|(m[544]&~m[585]&~m[586]&m[588]&m[589])|(~m[544]&m[585]&~m[586]&m[588]&m[589])|(m[544]&m[585]&~m[586]&m[588]&m[589])|(~m[544]&~m[585]&m[586]&m[588]&m[589])|(m[544]&~m[585]&m[586]&m[588]&m[589])|(m[544]&m[585]&m[586]&m[588]&m[589]))):InitCond[574];
    m[591] = run?((((m[288]&~m[590]&~m[592]&~m[593]&~m[594])|(~m[288]&~m[590]&~m[592]&m[593]&~m[594])|(m[288]&m[590]&~m[592]&m[593]&~m[594])|(m[288]&~m[590]&m[592]&m[593]&~m[594])|(~m[288]&m[590]&~m[592]&~m[593]&m[594])|(~m[288]&~m[590]&m[592]&~m[593]&m[594])|(m[288]&m[590]&m[592]&~m[593]&m[594])|(~m[288]&m[590]&m[592]&m[593]&m[594]))&UnbiasedRNG[236])|((m[288]&~m[590]&~m[592]&m[593]&~m[594])|(~m[288]&~m[590]&~m[592]&~m[593]&m[594])|(m[288]&~m[590]&~m[592]&~m[593]&m[594])|(m[288]&m[590]&~m[592]&~m[593]&m[594])|(m[288]&~m[590]&m[592]&~m[593]&m[594])|(~m[288]&~m[590]&~m[592]&m[593]&m[594])|(m[288]&~m[590]&~m[592]&m[593]&m[594])|(~m[288]&m[590]&~m[592]&m[593]&m[594])|(m[288]&m[590]&~m[592]&m[593]&m[594])|(~m[288]&~m[590]&m[592]&m[593]&m[594])|(m[288]&~m[590]&m[592]&m[593]&m[594])|(m[288]&m[590]&m[592]&m[593]&m[594]))):InitCond[575];
    m[596] = run?((((m[297]&~m[595]&~m[597]&~m[598]&~m[599])|(~m[297]&~m[595]&~m[597]&m[598]&~m[599])|(m[297]&m[595]&~m[597]&m[598]&~m[599])|(m[297]&~m[595]&m[597]&m[598]&~m[599])|(~m[297]&m[595]&~m[597]&~m[598]&m[599])|(~m[297]&~m[595]&m[597]&~m[598]&m[599])|(m[297]&m[595]&m[597]&~m[598]&m[599])|(~m[297]&m[595]&m[597]&m[598]&m[599]))&UnbiasedRNG[237])|((m[297]&~m[595]&~m[597]&m[598]&~m[599])|(~m[297]&~m[595]&~m[597]&~m[598]&m[599])|(m[297]&~m[595]&~m[597]&~m[598]&m[599])|(m[297]&m[595]&~m[597]&~m[598]&m[599])|(m[297]&~m[595]&m[597]&~m[598]&m[599])|(~m[297]&~m[595]&~m[597]&m[598]&m[599])|(m[297]&~m[595]&~m[597]&m[598]&m[599])|(~m[297]&m[595]&~m[597]&m[598]&m[599])|(m[297]&m[595]&~m[597]&m[598]&m[599])|(~m[297]&~m[595]&m[597]&m[598]&m[599])|(m[297]&~m[595]&m[597]&m[598]&m[599])|(m[297]&m[595]&m[597]&m[598]&m[599]))):InitCond[576];
    m[601] = run?((((m[306]&~m[600]&~m[602]&~m[603]&~m[604])|(~m[306]&~m[600]&~m[602]&m[603]&~m[604])|(m[306]&m[600]&~m[602]&m[603]&~m[604])|(m[306]&~m[600]&m[602]&m[603]&~m[604])|(~m[306]&m[600]&~m[602]&~m[603]&m[604])|(~m[306]&~m[600]&m[602]&~m[603]&m[604])|(m[306]&m[600]&m[602]&~m[603]&m[604])|(~m[306]&m[600]&m[602]&m[603]&m[604]))&UnbiasedRNG[238])|((m[306]&~m[600]&~m[602]&m[603]&~m[604])|(~m[306]&~m[600]&~m[602]&~m[603]&m[604])|(m[306]&~m[600]&~m[602]&~m[603]&m[604])|(m[306]&m[600]&~m[602]&~m[603]&m[604])|(m[306]&~m[600]&m[602]&~m[603]&m[604])|(~m[306]&~m[600]&~m[602]&m[603]&m[604])|(m[306]&~m[600]&~m[602]&m[603]&m[604])|(~m[306]&m[600]&~m[602]&m[603]&m[604])|(m[306]&m[600]&~m[602]&m[603]&m[604])|(~m[306]&~m[600]&m[602]&m[603]&m[604])|(m[306]&~m[600]&m[602]&m[603]&m[604])|(m[306]&m[600]&m[602]&m[603]&m[604]))):InitCond[577];
    m[606] = run?((((m[315]&~m[605]&~m[607]&~m[608]&~m[609])|(~m[315]&~m[605]&~m[607]&m[608]&~m[609])|(m[315]&m[605]&~m[607]&m[608]&~m[609])|(m[315]&~m[605]&m[607]&m[608]&~m[609])|(~m[315]&m[605]&~m[607]&~m[608]&m[609])|(~m[315]&~m[605]&m[607]&~m[608]&m[609])|(m[315]&m[605]&m[607]&~m[608]&m[609])|(~m[315]&m[605]&m[607]&m[608]&m[609]))&UnbiasedRNG[239])|((m[315]&~m[605]&~m[607]&m[608]&~m[609])|(~m[315]&~m[605]&~m[607]&~m[608]&m[609])|(m[315]&~m[605]&~m[607]&~m[608]&m[609])|(m[315]&m[605]&~m[607]&~m[608]&m[609])|(m[315]&~m[605]&m[607]&~m[608]&m[609])|(~m[315]&~m[605]&~m[607]&m[608]&m[609])|(m[315]&~m[605]&~m[607]&m[608]&m[609])|(~m[315]&m[605]&~m[607]&m[608]&m[609])|(m[315]&m[605]&~m[607]&m[608]&m[609])|(~m[315]&~m[605]&m[607]&m[608]&m[609])|(m[315]&~m[605]&m[607]&m[608]&m[609])|(m[315]&m[605]&m[607]&m[608]&m[609]))):InitCond[578];
    m[611] = run?((((m[324]&~m[610]&~m[612]&~m[613]&~m[614])|(~m[324]&~m[610]&~m[612]&m[613]&~m[614])|(m[324]&m[610]&~m[612]&m[613]&~m[614])|(m[324]&~m[610]&m[612]&m[613]&~m[614])|(~m[324]&m[610]&~m[612]&~m[613]&m[614])|(~m[324]&~m[610]&m[612]&~m[613]&m[614])|(m[324]&m[610]&m[612]&~m[613]&m[614])|(~m[324]&m[610]&m[612]&m[613]&m[614]))&UnbiasedRNG[240])|((m[324]&~m[610]&~m[612]&m[613]&~m[614])|(~m[324]&~m[610]&~m[612]&~m[613]&m[614])|(m[324]&~m[610]&~m[612]&~m[613]&m[614])|(m[324]&m[610]&~m[612]&~m[613]&m[614])|(m[324]&~m[610]&m[612]&~m[613]&m[614])|(~m[324]&~m[610]&~m[612]&m[613]&m[614])|(m[324]&~m[610]&~m[612]&m[613]&m[614])|(~m[324]&m[610]&~m[612]&m[613]&m[614])|(m[324]&m[610]&~m[612]&m[613]&m[614])|(~m[324]&~m[610]&m[612]&m[613]&m[614])|(m[324]&~m[610]&m[612]&m[613]&m[614])|(m[324]&m[610]&m[612]&m[613]&m[614]))):InitCond[579];
    m[616] = run?((((m[333]&~m[615]&~m[617]&~m[618]&~m[619])|(~m[333]&~m[615]&~m[617]&m[618]&~m[619])|(m[333]&m[615]&~m[617]&m[618]&~m[619])|(m[333]&~m[615]&m[617]&m[618]&~m[619])|(~m[333]&m[615]&~m[617]&~m[618]&m[619])|(~m[333]&~m[615]&m[617]&~m[618]&m[619])|(m[333]&m[615]&m[617]&~m[618]&m[619])|(~m[333]&m[615]&m[617]&m[618]&m[619]))&UnbiasedRNG[241])|((m[333]&~m[615]&~m[617]&m[618]&~m[619])|(~m[333]&~m[615]&~m[617]&~m[618]&m[619])|(m[333]&~m[615]&~m[617]&~m[618]&m[619])|(m[333]&m[615]&~m[617]&~m[618]&m[619])|(m[333]&~m[615]&m[617]&~m[618]&m[619])|(~m[333]&~m[615]&~m[617]&m[618]&m[619])|(m[333]&~m[615]&~m[617]&m[618]&m[619])|(~m[333]&m[615]&~m[617]&m[618]&m[619])|(m[333]&m[615]&~m[617]&m[618]&m[619])|(~m[333]&~m[615]&m[617]&m[618]&m[619])|(m[333]&~m[615]&m[617]&m[618]&m[619])|(m[333]&m[615]&m[617]&m[618]&m[619]))):InitCond[580];
    m[621] = run?((((m[342]&~m[620]&~m[622]&~m[623]&~m[624])|(~m[342]&~m[620]&~m[622]&m[623]&~m[624])|(m[342]&m[620]&~m[622]&m[623]&~m[624])|(m[342]&~m[620]&m[622]&m[623]&~m[624])|(~m[342]&m[620]&~m[622]&~m[623]&m[624])|(~m[342]&~m[620]&m[622]&~m[623]&m[624])|(m[342]&m[620]&m[622]&~m[623]&m[624])|(~m[342]&m[620]&m[622]&m[623]&m[624]))&UnbiasedRNG[242])|((m[342]&~m[620]&~m[622]&m[623]&~m[624])|(~m[342]&~m[620]&~m[622]&~m[623]&m[624])|(m[342]&~m[620]&~m[622]&~m[623]&m[624])|(m[342]&m[620]&~m[622]&~m[623]&m[624])|(m[342]&~m[620]&m[622]&~m[623]&m[624])|(~m[342]&~m[620]&~m[622]&m[623]&m[624])|(m[342]&~m[620]&~m[622]&m[623]&m[624])|(~m[342]&m[620]&~m[622]&m[623]&m[624])|(m[342]&m[620]&~m[622]&m[623]&m[624])|(~m[342]&~m[620]&m[622]&m[623]&m[624])|(m[342]&~m[620]&m[622]&m[623]&m[624])|(m[342]&m[620]&m[622]&m[623]&m[624]))):InitCond[581];
    m[627] = run?((((m[584]&~m[625]&~m[626]&~m[628]&~m[629])|(~m[584]&~m[625]&~m[626]&m[628]&~m[629])|(m[584]&m[625]&~m[626]&m[628]&~m[629])|(m[584]&~m[625]&m[626]&m[628]&~m[629])|(~m[584]&m[625]&~m[626]&~m[628]&m[629])|(~m[584]&~m[625]&m[626]&~m[628]&m[629])|(m[584]&m[625]&m[626]&~m[628]&m[629])|(~m[584]&m[625]&m[626]&m[628]&m[629]))&UnbiasedRNG[243])|((m[584]&~m[625]&~m[626]&m[628]&~m[629])|(~m[584]&~m[625]&~m[626]&~m[628]&m[629])|(m[584]&~m[625]&~m[626]&~m[628]&m[629])|(m[584]&m[625]&~m[626]&~m[628]&m[629])|(m[584]&~m[625]&m[626]&~m[628]&m[629])|(~m[584]&~m[625]&~m[626]&m[628]&m[629])|(m[584]&~m[625]&~m[626]&m[628]&m[629])|(~m[584]&m[625]&~m[626]&m[628]&m[629])|(m[584]&m[625]&~m[626]&m[628]&m[629])|(~m[584]&~m[625]&m[626]&m[628]&m[629])|(m[584]&~m[625]&m[626]&m[628]&m[629])|(m[584]&m[625]&m[626]&m[628]&m[629]))):InitCond[582];
    m[631] = run?((((m[289]&~m[630]&~m[632]&~m[633]&~m[634])|(~m[289]&~m[630]&~m[632]&m[633]&~m[634])|(m[289]&m[630]&~m[632]&m[633]&~m[634])|(m[289]&~m[630]&m[632]&m[633]&~m[634])|(~m[289]&m[630]&~m[632]&~m[633]&m[634])|(~m[289]&~m[630]&m[632]&~m[633]&m[634])|(m[289]&m[630]&m[632]&~m[633]&m[634])|(~m[289]&m[630]&m[632]&m[633]&m[634]))&UnbiasedRNG[244])|((m[289]&~m[630]&~m[632]&m[633]&~m[634])|(~m[289]&~m[630]&~m[632]&~m[633]&m[634])|(m[289]&~m[630]&~m[632]&~m[633]&m[634])|(m[289]&m[630]&~m[632]&~m[633]&m[634])|(m[289]&~m[630]&m[632]&~m[633]&m[634])|(~m[289]&~m[630]&~m[632]&m[633]&m[634])|(m[289]&~m[630]&~m[632]&m[633]&m[634])|(~m[289]&m[630]&~m[632]&m[633]&m[634])|(m[289]&m[630]&~m[632]&m[633]&m[634])|(~m[289]&~m[630]&m[632]&m[633]&m[634])|(m[289]&~m[630]&m[632]&m[633]&m[634])|(m[289]&m[630]&m[632]&m[633]&m[634]))):InitCond[583];
    m[636] = run?((((m[298]&~m[635]&~m[637]&~m[638]&~m[639])|(~m[298]&~m[635]&~m[637]&m[638]&~m[639])|(m[298]&m[635]&~m[637]&m[638]&~m[639])|(m[298]&~m[635]&m[637]&m[638]&~m[639])|(~m[298]&m[635]&~m[637]&~m[638]&m[639])|(~m[298]&~m[635]&m[637]&~m[638]&m[639])|(m[298]&m[635]&m[637]&~m[638]&m[639])|(~m[298]&m[635]&m[637]&m[638]&m[639]))&UnbiasedRNG[245])|((m[298]&~m[635]&~m[637]&m[638]&~m[639])|(~m[298]&~m[635]&~m[637]&~m[638]&m[639])|(m[298]&~m[635]&~m[637]&~m[638]&m[639])|(m[298]&m[635]&~m[637]&~m[638]&m[639])|(m[298]&~m[635]&m[637]&~m[638]&m[639])|(~m[298]&~m[635]&~m[637]&m[638]&m[639])|(m[298]&~m[635]&~m[637]&m[638]&m[639])|(~m[298]&m[635]&~m[637]&m[638]&m[639])|(m[298]&m[635]&~m[637]&m[638]&m[639])|(~m[298]&~m[635]&m[637]&m[638]&m[639])|(m[298]&~m[635]&m[637]&m[638]&m[639])|(m[298]&m[635]&m[637]&m[638]&m[639]))):InitCond[584];
    m[641] = run?((((m[307]&~m[640]&~m[642]&~m[643]&~m[644])|(~m[307]&~m[640]&~m[642]&m[643]&~m[644])|(m[307]&m[640]&~m[642]&m[643]&~m[644])|(m[307]&~m[640]&m[642]&m[643]&~m[644])|(~m[307]&m[640]&~m[642]&~m[643]&m[644])|(~m[307]&~m[640]&m[642]&~m[643]&m[644])|(m[307]&m[640]&m[642]&~m[643]&m[644])|(~m[307]&m[640]&m[642]&m[643]&m[644]))&UnbiasedRNG[246])|((m[307]&~m[640]&~m[642]&m[643]&~m[644])|(~m[307]&~m[640]&~m[642]&~m[643]&m[644])|(m[307]&~m[640]&~m[642]&~m[643]&m[644])|(m[307]&m[640]&~m[642]&~m[643]&m[644])|(m[307]&~m[640]&m[642]&~m[643]&m[644])|(~m[307]&~m[640]&~m[642]&m[643]&m[644])|(m[307]&~m[640]&~m[642]&m[643]&m[644])|(~m[307]&m[640]&~m[642]&m[643]&m[644])|(m[307]&m[640]&~m[642]&m[643]&m[644])|(~m[307]&~m[640]&m[642]&m[643]&m[644])|(m[307]&~m[640]&m[642]&m[643]&m[644])|(m[307]&m[640]&m[642]&m[643]&m[644]))):InitCond[585];
    m[646] = run?((((m[316]&~m[645]&~m[647]&~m[648]&~m[649])|(~m[316]&~m[645]&~m[647]&m[648]&~m[649])|(m[316]&m[645]&~m[647]&m[648]&~m[649])|(m[316]&~m[645]&m[647]&m[648]&~m[649])|(~m[316]&m[645]&~m[647]&~m[648]&m[649])|(~m[316]&~m[645]&m[647]&~m[648]&m[649])|(m[316]&m[645]&m[647]&~m[648]&m[649])|(~m[316]&m[645]&m[647]&m[648]&m[649]))&UnbiasedRNG[247])|((m[316]&~m[645]&~m[647]&m[648]&~m[649])|(~m[316]&~m[645]&~m[647]&~m[648]&m[649])|(m[316]&~m[645]&~m[647]&~m[648]&m[649])|(m[316]&m[645]&~m[647]&~m[648]&m[649])|(m[316]&~m[645]&m[647]&~m[648]&m[649])|(~m[316]&~m[645]&~m[647]&m[648]&m[649])|(m[316]&~m[645]&~m[647]&m[648]&m[649])|(~m[316]&m[645]&~m[647]&m[648]&m[649])|(m[316]&m[645]&~m[647]&m[648]&m[649])|(~m[316]&~m[645]&m[647]&m[648]&m[649])|(m[316]&~m[645]&m[647]&m[648]&m[649])|(m[316]&m[645]&m[647]&m[648]&m[649]))):InitCond[586];
    m[651] = run?((((m[325]&~m[650]&~m[652]&~m[653]&~m[654])|(~m[325]&~m[650]&~m[652]&m[653]&~m[654])|(m[325]&m[650]&~m[652]&m[653]&~m[654])|(m[325]&~m[650]&m[652]&m[653]&~m[654])|(~m[325]&m[650]&~m[652]&~m[653]&m[654])|(~m[325]&~m[650]&m[652]&~m[653]&m[654])|(m[325]&m[650]&m[652]&~m[653]&m[654])|(~m[325]&m[650]&m[652]&m[653]&m[654]))&UnbiasedRNG[248])|((m[325]&~m[650]&~m[652]&m[653]&~m[654])|(~m[325]&~m[650]&~m[652]&~m[653]&m[654])|(m[325]&~m[650]&~m[652]&~m[653]&m[654])|(m[325]&m[650]&~m[652]&~m[653]&m[654])|(m[325]&~m[650]&m[652]&~m[653]&m[654])|(~m[325]&~m[650]&~m[652]&m[653]&m[654])|(m[325]&~m[650]&~m[652]&m[653]&m[654])|(~m[325]&m[650]&~m[652]&m[653]&m[654])|(m[325]&m[650]&~m[652]&m[653]&m[654])|(~m[325]&~m[650]&m[652]&m[653]&m[654])|(m[325]&~m[650]&m[652]&m[653]&m[654])|(m[325]&m[650]&m[652]&m[653]&m[654]))):InitCond[587];
    m[656] = run?((((m[334]&~m[655]&~m[657]&~m[658]&~m[659])|(~m[334]&~m[655]&~m[657]&m[658]&~m[659])|(m[334]&m[655]&~m[657]&m[658]&~m[659])|(m[334]&~m[655]&m[657]&m[658]&~m[659])|(~m[334]&m[655]&~m[657]&~m[658]&m[659])|(~m[334]&~m[655]&m[657]&~m[658]&m[659])|(m[334]&m[655]&m[657]&~m[658]&m[659])|(~m[334]&m[655]&m[657]&m[658]&m[659]))&UnbiasedRNG[249])|((m[334]&~m[655]&~m[657]&m[658]&~m[659])|(~m[334]&~m[655]&~m[657]&~m[658]&m[659])|(m[334]&~m[655]&~m[657]&~m[658]&m[659])|(m[334]&m[655]&~m[657]&~m[658]&m[659])|(m[334]&~m[655]&m[657]&~m[658]&m[659])|(~m[334]&~m[655]&~m[657]&m[658]&m[659])|(m[334]&~m[655]&~m[657]&m[658]&m[659])|(~m[334]&m[655]&~m[657]&m[658]&m[659])|(m[334]&m[655]&~m[657]&m[658]&m[659])|(~m[334]&~m[655]&m[657]&m[658]&m[659])|(m[334]&~m[655]&m[657]&m[658]&m[659])|(m[334]&m[655]&m[657]&m[658]&m[659]))):InitCond[588];
    m[661] = run?((((m[343]&~m[660]&~m[662]&~m[663]&~m[664])|(~m[343]&~m[660]&~m[662]&m[663]&~m[664])|(m[343]&m[660]&~m[662]&m[663]&~m[664])|(m[343]&~m[660]&m[662]&m[663]&~m[664])|(~m[343]&m[660]&~m[662]&~m[663]&m[664])|(~m[343]&~m[660]&m[662]&~m[663]&m[664])|(m[343]&m[660]&m[662]&~m[663]&m[664])|(~m[343]&m[660]&m[662]&m[663]&m[664]))&UnbiasedRNG[250])|((m[343]&~m[660]&~m[662]&m[663]&~m[664])|(~m[343]&~m[660]&~m[662]&~m[663]&m[664])|(m[343]&~m[660]&~m[662]&~m[663]&m[664])|(m[343]&m[660]&~m[662]&~m[663]&m[664])|(m[343]&~m[660]&m[662]&~m[663]&m[664])|(~m[343]&~m[660]&~m[662]&m[663]&m[664])|(m[343]&~m[660]&~m[662]&m[663]&m[664])|(~m[343]&m[660]&~m[662]&m[663]&m[664])|(m[343]&m[660]&~m[662]&m[663]&m[664])|(~m[343]&~m[660]&m[662]&m[663]&m[664])|(m[343]&~m[660]&m[662]&m[663]&m[664])|(m[343]&m[660]&m[662]&m[663]&m[664]))):InitCond[589];
    m[666] = run?((((m[352]&~m[665]&~m[667]&~m[668]&~m[669])|(~m[352]&~m[665]&~m[667]&m[668]&~m[669])|(m[352]&m[665]&~m[667]&m[668]&~m[669])|(m[352]&~m[665]&m[667]&m[668]&~m[669])|(~m[352]&m[665]&~m[667]&~m[668]&m[669])|(~m[352]&~m[665]&m[667]&~m[668]&m[669])|(m[352]&m[665]&m[667]&~m[668]&m[669])|(~m[352]&m[665]&m[667]&m[668]&m[669]))&UnbiasedRNG[251])|((m[352]&~m[665]&~m[667]&m[668]&~m[669])|(~m[352]&~m[665]&~m[667]&~m[668]&m[669])|(m[352]&~m[665]&~m[667]&~m[668]&m[669])|(m[352]&m[665]&~m[667]&~m[668]&m[669])|(m[352]&~m[665]&m[667]&~m[668]&m[669])|(~m[352]&~m[665]&~m[667]&m[668]&m[669])|(m[352]&~m[665]&~m[667]&m[668]&m[669])|(~m[352]&m[665]&~m[667]&m[668]&m[669])|(m[352]&m[665]&~m[667]&m[668]&m[669])|(~m[352]&~m[665]&m[667]&m[668]&m[669])|(m[352]&~m[665]&m[667]&m[668]&m[669])|(m[352]&m[665]&m[667]&m[668]&m[669]))):InitCond[590];
    m[671] = run?((((m[299]&~m[670]&~m[672]&~m[673]&~m[674])|(~m[299]&~m[670]&~m[672]&m[673]&~m[674])|(m[299]&m[670]&~m[672]&m[673]&~m[674])|(m[299]&~m[670]&m[672]&m[673]&~m[674])|(~m[299]&m[670]&~m[672]&~m[673]&m[674])|(~m[299]&~m[670]&m[672]&~m[673]&m[674])|(m[299]&m[670]&m[672]&~m[673]&m[674])|(~m[299]&m[670]&m[672]&m[673]&m[674]))&UnbiasedRNG[252])|((m[299]&~m[670]&~m[672]&m[673]&~m[674])|(~m[299]&~m[670]&~m[672]&~m[673]&m[674])|(m[299]&~m[670]&~m[672]&~m[673]&m[674])|(m[299]&m[670]&~m[672]&~m[673]&m[674])|(m[299]&~m[670]&m[672]&~m[673]&m[674])|(~m[299]&~m[670]&~m[672]&m[673]&m[674])|(m[299]&~m[670]&~m[672]&m[673]&m[674])|(~m[299]&m[670]&~m[672]&m[673]&m[674])|(m[299]&m[670]&~m[672]&m[673]&m[674])|(~m[299]&~m[670]&m[672]&m[673]&m[674])|(m[299]&~m[670]&m[672]&m[673]&m[674])|(m[299]&m[670]&m[672]&m[673]&m[674]))):InitCond[591];
    m[676] = run?((((m[308]&~m[675]&~m[677]&~m[678]&~m[679])|(~m[308]&~m[675]&~m[677]&m[678]&~m[679])|(m[308]&m[675]&~m[677]&m[678]&~m[679])|(m[308]&~m[675]&m[677]&m[678]&~m[679])|(~m[308]&m[675]&~m[677]&~m[678]&m[679])|(~m[308]&~m[675]&m[677]&~m[678]&m[679])|(m[308]&m[675]&m[677]&~m[678]&m[679])|(~m[308]&m[675]&m[677]&m[678]&m[679]))&UnbiasedRNG[253])|((m[308]&~m[675]&~m[677]&m[678]&~m[679])|(~m[308]&~m[675]&~m[677]&~m[678]&m[679])|(m[308]&~m[675]&~m[677]&~m[678]&m[679])|(m[308]&m[675]&~m[677]&~m[678]&m[679])|(m[308]&~m[675]&m[677]&~m[678]&m[679])|(~m[308]&~m[675]&~m[677]&m[678]&m[679])|(m[308]&~m[675]&~m[677]&m[678]&m[679])|(~m[308]&m[675]&~m[677]&m[678]&m[679])|(m[308]&m[675]&~m[677]&m[678]&m[679])|(~m[308]&~m[675]&m[677]&m[678]&m[679])|(m[308]&~m[675]&m[677]&m[678]&m[679])|(m[308]&m[675]&m[677]&m[678]&m[679]))):InitCond[592];
    m[681] = run?((((m[317]&~m[680]&~m[682]&~m[683]&~m[684])|(~m[317]&~m[680]&~m[682]&m[683]&~m[684])|(m[317]&m[680]&~m[682]&m[683]&~m[684])|(m[317]&~m[680]&m[682]&m[683]&~m[684])|(~m[317]&m[680]&~m[682]&~m[683]&m[684])|(~m[317]&~m[680]&m[682]&~m[683]&m[684])|(m[317]&m[680]&m[682]&~m[683]&m[684])|(~m[317]&m[680]&m[682]&m[683]&m[684]))&UnbiasedRNG[254])|((m[317]&~m[680]&~m[682]&m[683]&~m[684])|(~m[317]&~m[680]&~m[682]&~m[683]&m[684])|(m[317]&~m[680]&~m[682]&~m[683]&m[684])|(m[317]&m[680]&~m[682]&~m[683]&m[684])|(m[317]&~m[680]&m[682]&~m[683]&m[684])|(~m[317]&~m[680]&~m[682]&m[683]&m[684])|(m[317]&~m[680]&~m[682]&m[683]&m[684])|(~m[317]&m[680]&~m[682]&m[683]&m[684])|(m[317]&m[680]&~m[682]&m[683]&m[684])|(~m[317]&~m[680]&m[682]&m[683]&m[684])|(m[317]&~m[680]&m[682]&m[683]&m[684])|(m[317]&m[680]&m[682]&m[683]&m[684]))):InitCond[593];
    m[686] = run?((((m[326]&~m[685]&~m[687]&~m[688]&~m[689])|(~m[326]&~m[685]&~m[687]&m[688]&~m[689])|(m[326]&m[685]&~m[687]&m[688]&~m[689])|(m[326]&~m[685]&m[687]&m[688]&~m[689])|(~m[326]&m[685]&~m[687]&~m[688]&m[689])|(~m[326]&~m[685]&m[687]&~m[688]&m[689])|(m[326]&m[685]&m[687]&~m[688]&m[689])|(~m[326]&m[685]&m[687]&m[688]&m[689]))&UnbiasedRNG[255])|((m[326]&~m[685]&~m[687]&m[688]&~m[689])|(~m[326]&~m[685]&~m[687]&~m[688]&m[689])|(m[326]&~m[685]&~m[687]&~m[688]&m[689])|(m[326]&m[685]&~m[687]&~m[688]&m[689])|(m[326]&~m[685]&m[687]&~m[688]&m[689])|(~m[326]&~m[685]&~m[687]&m[688]&m[689])|(m[326]&~m[685]&~m[687]&m[688]&m[689])|(~m[326]&m[685]&~m[687]&m[688]&m[689])|(m[326]&m[685]&~m[687]&m[688]&m[689])|(~m[326]&~m[685]&m[687]&m[688]&m[689])|(m[326]&~m[685]&m[687]&m[688]&m[689])|(m[326]&m[685]&m[687]&m[688]&m[689]))):InitCond[594];
    m[691] = run?((((m[335]&~m[690]&~m[692]&~m[693]&~m[694])|(~m[335]&~m[690]&~m[692]&m[693]&~m[694])|(m[335]&m[690]&~m[692]&m[693]&~m[694])|(m[335]&~m[690]&m[692]&m[693]&~m[694])|(~m[335]&m[690]&~m[692]&~m[693]&m[694])|(~m[335]&~m[690]&m[692]&~m[693]&m[694])|(m[335]&m[690]&m[692]&~m[693]&m[694])|(~m[335]&m[690]&m[692]&m[693]&m[694]))&UnbiasedRNG[256])|((m[335]&~m[690]&~m[692]&m[693]&~m[694])|(~m[335]&~m[690]&~m[692]&~m[693]&m[694])|(m[335]&~m[690]&~m[692]&~m[693]&m[694])|(m[335]&m[690]&~m[692]&~m[693]&m[694])|(m[335]&~m[690]&m[692]&~m[693]&m[694])|(~m[335]&~m[690]&~m[692]&m[693]&m[694])|(m[335]&~m[690]&~m[692]&m[693]&m[694])|(~m[335]&m[690]&~m[692]&m[693]&m[694])|(m[335]&m[690]&~m[692]&m[693]&m[694])|(~m[335]&~m[690]&m[692]&m[693]&m[694])|(m[335]&~m[690]&m[692]&m[693]&m[694])|(m[335]&m[690]&m[692]&m[693]&m[694]))):InitCond[595];
    m[696] = run?((((m[344]&~m[695]&~m[697]&~m[698]&~m[699])|(~m[344]&~m[695]&~m[697]&m[698]&~m[699])|(m[344]&m[695]&~m[697]&m[698]&~m[699])|(m[344]&~m[695]&m[697]&m[698]&~m[699])|(~m[344]&m[695]&~m[697]&~m[698]&m[699])|(~m[344]&~m[695]&m[697]&~m[698]&m[699])|(m[344]&m[695]&m[697]&~m[698]&m[699])|(~m[344]&m[695]&m[697]&m[698]&m[699]))&UnbiasedRNG[257])|((m[344]&~m[695]&~m[697]&m[698]&~m[699])|(~m[344]&~m[695]&~m[697]&~m[698]&m[699])|(m[344]&~m[695]&~m[697]&~m[698]&m[699])|(m[344]&m[695]&~m[697]&~m[698]&m[699])|(m[344]&~m[695]&m[697]&~m[698]&m[699])|(~m[344]&~m[695]&~m[697]&m[698]&m[699])|(m[344]&~m[695]&~m[697]&m[698]&m[699])|(~m[344]&m[695]&~m[697]&m[698]&m[699])|(m[344]&m[695]&~m[697]&m[698]&m[699])|(~m[344]&~m[695]&m[697]&m[698]&m[699])|(m[344]&~m[695]&m[697]&m[698]&m[699])|(m[344]&m[695]&m[697]&m[698]&m[699]))):InitCond[596];
    m[701] = run?((((m[353]&~m[700]&~m[702]&~m[703]&~m[704])|(~m[353]&~m[700]&~m[702]&m[703]&~m[704])|(m[353]&m[700]&~m[702]&m[703]&~m[704])|(m[353]&~m[700]&m[702]&m[703]&~m[704])|(~m[353]&m[700]&~m[702]&~m[703]&m[704])|(~m[353]&~m[700]&m[702]&~m[703]&m[704])|(m[353]&m[700]&m[702]&~m[703]&m[704])|(~m[353]&m[700]&m[702]&m[703]&m[704]))&UnbiasedRNG[258])|((m[353]&~m[700]&~m[702]&m[703]&~m[704])|(~m[353]&~m[700]&~m[702]&~m[703]&m[704])|(m[353]&~m[700]&~m[702]&~m[703]&m[704])|(m[353]&m[700]&~m[702]&~m[703]&m[704])|(m[353]&~m[700]&m[702]&~m[703]&m[704])|(~m[353]&~m[700]&~m[702]&m[703]&m[704])|(m[353]&~m[700]&~m[702]&m[703]&m[704])|(~m[353]&m[700]&~m[702]&m[703]&m[704])|(m[353]&m[700]&~m[702]&m[703]&m[704])|(~m[353]&~m[700]&m[702]&m[703]&m[704])|(m[353]&~m[700]&m[702]&m[703]&m[704])|(m[353]&m[700]&m[702]&m[703]&m[704]))):InitCond[597];
    m[706] = run?((((m[309]&~m[705]&~m[707]&~m[708]&~m[709])|(~m[309]&~m[705]&~m[707]&m[708]&~m[709])|(m[309]&m[705]&~m[707]&m[708]&~m[709])|(m[309]&~m[705]&m[707]&m[708]&~m[709])|(~m[309]&m[705]&~m[707]&~m[708]&m[709])|(~m[309]&~m[705]&m[707]&~m[708]&m[709])|(m[309]&m[705]&m[707]&~m[708]&m[709])|(~m[309]&m[705]&m[707]&m[708]&m[709]))&UnbiasedRNG[259])|((m[309]&~m[705]&~m[707]&m[708]&~m[709])|(~m[309]&~m[705]&~m[707]&~m[708]&m[709])|(m[309]&~m[705]&~m[707]&~m[708]&m[709])|(m[309]&m[705]&~m[707]&~m[708]&m[709])|(m[309]&~m[705]&m[707]&~m[708]&m[709])|(~m[309]&~m[705]&~m[707]&m[708]&m[709])|(m[309]&~m[705]&~m[707]&m[708]&m[709])|(~m[309]&m[705]&~m[707]&m[708]&m[709])|(m[309]&m[705]&~m[707]&m[708]&m[709])|(~m[309]&~m[705]&m[707]&m[708]&m[709])|(m[309]&~m[705]&m[707]&m[708]&m[709])|(m[309]&m[705]&m[707]&m[708]&m[709]))):InitCond[598];
    m[711] = run?((((m[318]&~m[710]&~m[712]&~m[713]&~m[714])|(~m[318]&~m[710]&~m[712]&m[713]&~m[714])|(m[318]&m[710]&~m[712]&m[713]&~m[714])|(m[318]&~m[710]&m[712]&m[713]&~m[714])|(~m[318]&m[710]&~m[712]&~m[713]&m[714])|(~m[318]&~m[710]&m[712]&~m[713]&m[714])|(m[318]&m[710]&m[712]&~m[713]&m[714])|(~m[318]&m[710]&m[712]&m[713]&m[714]))&UnbiasedRNG[260])|((m[318]&~m[710]&~m[712]&m[713]&~m[714])|(~m[318]&~m[710]&~m[712]&~m[713]&m[714])|(m[318]&~m[710]&~m[712]&~m[713]&m[714])|(m[318]&m[710]&~m[712]&~m[713]&m[714])|(m[318]&~m[710]&m[712]&~m[713]&m[714])|(~m[318]&~m[710]&~m[712]&m[713]&m[714])|(m[318]&~m[710]&~m[712]&m[713]&m[714])|(~m[318]&m[710]&~m[712]&m[713]&m[714])|(m[318]&m[710]&~m[712]&m[713]&m[714])|(~m[318]&~m[710]&m[712]&m[713]&m[714])|(m[318]&~m[710]&m[712]&m[713]&m[714])|(m[318]&m[710]&m[712]&m[713]&m[714]))):InitCond[599];
    m[716] = run?((((m[327]&~m[715]&~m[717]&~m[718]&~m[719])|(~m[327]&~m[715]&~m[717]&m[718]&~m[719])|(m[327]&m[715]&~m[717]&m[718]&~m[719])|(m[327]&~m[715]&m[717]&m[718]&~m[719])|(~m[327]&m[715]&~m[717]&~m[718]&m[719])|(~m[327]&~m[715]&m[717]&~m[718]&m[719])|(m[327]&m[715]&m[717]&~m[718]&m[719])|(~m[327]&m[715]&m[717]&m[718]&m[719]))&UnbiasedRNG[261])|((m[327]&~m[715]&~m[717]&m[718]&~m[719])|(~m[327]&~m[715]&~m[717]&~m[718]&m[719])|(m[327]&~m[715]&~m[717]&~m[718]&m[719])|(m[327]&m[715]&~m[717]&~m[718]&m[719])|(m[327]&~m[715]&m[717]&~m[718]&m[719])|(~m[327]&~m[715]&~m[717]&m[718]&m[719])|(m[327]&~m[715]&~m[717]&m[718]&m[719])|(~m[327]&m[715]&~m[717]&m[718]&m[719])|(m[327]&m[715]&~m[717]&m[718]&m[719])|(~m[327]&~m[715]&m[717]&m[718]&m[719])|(m[327]&~m[715]&m[717]&m[718]&m[719])|(m[327]&m[715]&m[717]&m[718]&m[719]))):InitCond[600];
    m[721] = run?((((m[336]&~m[720]&~m[722]&~m[723]&~m[724])|(~m[336]&~m[720]&~m[722]&m[723]&~m[724])|(m[336]&m[720]&~m[722]&m[723]&~m[724])|(m[336]&~m[720]&m[722]&m[723]&~m[724])|(~m[336]&m[720]&~m[722]&~m[723]&m[724])|(~m[336]&~m[720]&m[722]&~m[723]&m[724])|(m[336]&m[720]&m[722]&~m[723]&m[724])|(~m[336]&m[720]&m[722]&m[723]&m[724]))&UnbiasedRNG[262])|((m[336]&~m[720]&~m[722]&m[723]&~m[724])|(~m[336]&~m[720]&~m[722]&~m[723]&m[724])|(m[336]&~m[720]&~m[722]&~m[723]&m[724])|(m[336]&m[720]&~m[722]&~m[723]&m[724])|(m[336]&~m[720]&m[722]&~m[723]&m[724])|(~m[336]&~m[720]&~m[722]&m[723]&m[724])|(m[336]&~m[720]&~m[722]&m[723]&m[724])|(~m[336]&m[720]&~m[722]&m[723]&m[724])|(m[336]&m[720]&~m[722]&m[723]&m[724])|(~m[336]&~m[720]&m[722]&m[723]&m[724])|(m[336]&~m[720]&m[722]&m[723]&m[724])|(m[336]&m[720]&m[722]&m[723]&m[724]))):InitCond[601];
    m[726] = run?((((m[345]&~m[725]&~m[727]&~m[728]&~m[729])|(~m[345]&~m[725]&~m[727]&m[728]&~m[729])|(m[345]&m[725]&~m[727]&m[728]&~m[729])|(m[345]&~m[725]&m[727]&m[728]&~m[729])|(~m[345]&m[725]&~m[727]&~m[728]&m[729])|(~m[345]&~m[725]&m[727]&~m[728]&m[729])|(m[345]&m[725]&m[727]&~m[728]&m[729])|(~m[345]&m[725]&m[727]&m[728]&m[729]))&UnbiasedRNG[263])|((m[345]&~m[725]&~m[727]&m[728]&~m[729])|(~m[345]&~m[725]&~m[727]&~m[728]&m[729])|(m[345]&~m[725]&~m[727]&~m[728]&m[729])|(m[345]&m[725]&~m[727]&~m[728]&m[729])|(m[345]&~m[725]&m[727]&~m[728]&m[729])|(~m[345]&~m[725]&~m[727]&m[728]&m[729])|(m[345]&~m[725]&~m[727]&m[728]&m[729])|(~m[345]&m[725]&~m[727]&m[728]&m[729])|(m[345]&m[725]&~m[727]&m[728]&m[729])|(~m[345]&~m[725]&m[727]&m[728]&m[729])|(m[345]&~m[725]&m[727]&m[728]&m[729])|(m[345]&m[725]&m[727]&m[728]&m[729]))):InitCond[602];
    m[731] = run?((((m[354]&~m[730]&~m[732]&~m[733]&~m[734])|(~m[354]&~m[730]&~m[732]&m[733]&~m[734])|(m[354]&m[730]&~m[732]&m[733]&~m[734])|(m[354]&~m[730]&m[732]&m[733]&~m[734])|(~m[354]&m[730]&~m[732]&~m[733]&m[734])|(~m[354]&~m[730]&m[732]&~m[733]&m[734])|(m[354]&m[730]&m[732]&~m[733]&m[734])|(~m[354]&m[730]&m[732]&m[733]&m[734]))&UnbiasedRNG[264])|((m[354]&~m[730]&~m[732]&m[733]&~m[734])|(~m[354]&~m[730]&~m[732]&~m[733]&m[734])|(m[354]&~m[730]&~m[732]&~m[733]&m[734])|(m[354]&m[730]&~m[732]&~m[733]&m[734])|(m[354]&~m[730]&m[732]&~m[733]&m[734])|(~m[354]&~m[730]&~m[732]&m[733]&m[734])|(m[354]&~m[730]&~m[732]&m[733]&m[734])|(~m[354]&m[730]&~m[732]&m[733]&m[734])|(m[354]&m[730]&~m[732]&m[733]&m[734])|(~m[354]&~m[730]&m[732]&m[733]&m[734])|(m[354]&~m[730]&m[732]&m[733]&m[734])|(m[354]&m[730]&m[732]&m[733]&m[734]))):InitCond[603];
    m[736] = run?((((m[319]&~m[735]&~m[737]&~m[738]&~m[739])|(~m[319]&~m[735]&~m[737]&m[738]&~m[739])|(m[319]&m[735]&~m[737]&m[738]&~m[739])|(m[319]&~m[735]&m[737]&m[738]&~m[739])|(~m[319]&m[735]&~m[737]&~m[738]&m[739])|(~m[319]&~m[735]&m[737]&~m[738]&m[739])|(m[319]&m[735]&m[737]&~m[738]&m[739])|(~m[319]&m[735]&m[737]&m[738]&m[739]))&UnbiasedRNG[265])|((m[319]&~m[735]&~m[737]&m[738]&~m[739])|(~m[319]&~m[735]&~m[737]&~m[738]&m[739])|(m[319]&~m[735]&~m[737]&~m[738]&m[739])|(m[319]&m[735]&~m[737]&~m[738]&m[739])|(m[319]&~m[735]&m[737]&~m[738]&m[739])|(~m[319]&~m[735]&~m[737]&m[738]&m[739])|(m[319]&~m[735]&~m[737]&m[738]&m[739])|(~m[319]&m[735]&~m[737]&m[738]&m[739])|(m[319]&m[735]&~m[737]&m[738]&m[739])|(~m[319]&~m[735]&m[737]&m[738]&m[739])|(m[319]&~m[735]&m[737]&m[738]&m[739])|(m[319]&m[735]&m[737]&m[738]&m[739]))):InitCond[604];
    m[741] = run?((((m[328]&~m[740]&~m[742]&~m[743]&~m[744])|(~m[328]&~m[740]&~m[742]&m[743]&~m[744])|(m[328]&m[740]&~m[742]&m[743]&~m[744])|(m[328]&~m[740]&m[742]&m[743]&~m[744])|(~m[328]&m[740]&~m[742]&~m[743]&m[744])|(~m[328]&~m[740]&m[742]&~m[743]&m[744])|(m[328]&m[740]&m[742]&~m[743]&m[744])|(~m[328]&m[740]&m[742]&m[743]&m[744]))&UnbiasedRNG[266])|((m[328]&~m[740]&~m[742]&m[743]&~m[744])|(~m[328]&~m[740]&~m[742]&~m[743]&m[744])|(m[328]&~m[740]&~m[742]&~m[743]&m[744])|(m[328]&m[740]&~m[742]&~m[743]&m[744])|(m[328]&~m[740]&m[742]&~m[743]&m[744])|(~m[328]&~m[740]&~m[742]&m[743]&m[744])|(m[328]&~m[740]&~m[742]&m[743]&m[744])|(~m[328]&m[740]&~m[742]&m[743]&m[744])|(m[328]&m[740]&~m[742]&m[743]&m[744])|(~m[328]&~m[740]&m[742]&m[743]&m[744])|(m[328]&~m[740]&m[742]&m[743]&m[744])|(m[328]&m[740]&m[742]&m[743]&m[744]))):InitCond[605];
    m[746] = run?((((m[337]&~m[745]&~m[747]&~m[748]&~m[749])|(~m[337]&~m[745]&~m[747]&m[748]&~m[749])|(m[337]&m[745]&~m[747]&m[748]&~m[749])|(m[337]&~m[745]&m[747]&m[748]&~m[749])|(~m[337]&m[745]&~m[747]&~m[748]&m[749])|(~m[337]&~m[745]&m[747]&~m[748]&m[749])|(m[337]&m[745]&m[747]&~m[748]&m[749])|(~m[337]&m[745]&m[747]&m[748]&m[749]))&UnbiasedRNG[267])|((m[337]&~m[745]&~m[747]&m[748]&~m[749])|(~m[337]&~m[745]&~m[747]&~m[748]&m[749])|(m[337]&~m[745]&~m[747]&~m[748]&m[749])|(m[337]&m[745]&~m[747]&~m[748]&m[749])|(m[337]&~m[745]&m[747]&~m[748]&m[749])|(~m[337]&~m[745]&~m[747]&m[748]&m[749])|(m[337]&~m[745]&~m[747]&m[748]&m[749])|(~m[337]&m[745]&~m[747]&m[748]&m[749])|(m[337]&m[745]&~m[747]&m[748]&m[749])|(~m[337]&~m[745]&m[747]&m[748]&m[749])|(m[337]&~m[745]&m[747]&m[748]&m[749])|(m[337]&m[745]&m[747]&m[748]&m[749]))):InitCond[606];
    m[751] = run?((((m[346]&~m[750]&~m[752]&~m[753]&~m[754])|(~m[346]&~m[750]&~m[752]&m[753]&~m[754])|(m[346]&m[750]&~m[752]&m[753]&~m[754])|(m[346]&~m[750]&m[752]&m[753]&~m[754])|(~m[346]&m[750]&~m[752]&~m[753]&m[754])|(~m[346]&~m[750]&m[752]&~m[753]&m[754])|(m[346]&m[750]&m[752]&~m[753]&m[754])|(~m[346]&m[750]&m[752]&m[753]&m[754]))&UnbiasedRNG[268])|((m[346]&~m[750]&~m[752]&m[753]&~m[754])|(~m[346]&~m[750]&~m[752]&~m[753]&m[754])|(m[346]&~m[750]&~m[752]&~m[753]&m[754])|(m[346]&m[750]&~m[752]&~m[753]&m[754])|(m[346]&~m[750]&m[752]&~m[753]&m[754])|(~m[346]&~m[750]&~m[752]&m[753]&m[754])|(m[346]&~m[750]&~m[752]&m[753]&m[754])|(~m[346]&m[750]&~m[752]&m[753]&m[754])|(m[346]&m[750]&~m[752]&m[753]&m[754])|(~m[346]&~m[750]&m[752]&m[753]&m[754])|(m[346]&~m[750]&m[752]&m[753]&m[754])|(m[346]&m[750]&m[752]&m[753]&m[754]))):InitCond[607];
    m[756] = run?((((m[355]&~m[755]&~m[757]&~m[758]&~m[759])|(~m[355]&~m[755]&~m[757]&m[758]&~m[759])|(m[355]&m[755]&~m[757]&m[758]&~m[759])|(m[355]&~m[755]&m[757]&m[758]&~m[759])|(~m[355]&m[755]&~m[757]&~m[758]&m[759])|(~m[355]&~m[755]&m[757]&~m[758]&m[759])|(m[355]&m[755]&m[757]&~m[758]&m[759])|(~m[355]&m[755]&m[757]&m[758]&m[759]))&UnbiasedRNG[269])|((m[355]&~m[755]&~m[757]&m[758]&~m[759])|(~m[355]&~m[755]&~m[757]&~m[758]&m[759])|(m[355]&~m[755]&~m[757]&~m[758]&m[759])|(m[355]&m[755]&~m[757]&~m[758]&m[759])|(m[355]&~m[755]&m[757]&~m[758]&m[759])|(~m[355]&~m[755]&~m[757]&m[758]&m[759])|(m[355]&~m[755]&~m[757]&m[758]&m[759])|(~m[355]&m[755]&~m[757]&m[758]&m[759])|(m[355]&m[755]&~m[757]&m[758]&m[759])|(~m[355]&~m[755]&m[757]&m[758]&m[759])|(m[355]&~m[755]&m[757]&m[758]&m[759])|(m[355]&m[755]&m[757]&m[758]&m[759]))):InitCond[608];
    m[761] = run?((((m[329]&~m[760]&~m[762]&~m[763]&~m[764])|(~m[329]&~m[760]&~m[762]&m[763]&~m[764])|(m[329]&m[760]&~m[762]&m[763]&~m[764])|(m[329]&~m[760]&m[762]&m[763]&~m[764])|(~m[329]&m[760]&~m[762]&~m[763]&m[764])|(~m[329]&~m[760]&m[762]&~m[763]&m[764])|(m[329]&m[760]&m[762]&~m[763]&m[764])|(~m[329]&m[760]&m[762]&m[763]&m[764]))&UnbiasedRNG[270])|((m[329]&~m[760]&~m[762]&m[763]&~m[764])|(~m[329]&~m[760]&~m[762]&~m[763]&m[764])|(m[329]&~m[760]&~m[762]&~m[763]&m[764])|(m[329]&m[760]&~m[762]&~m[763]&m[764])|(m[329]&~m[760]&m[762]&~m[763]&m[764])|(~m[329]&~m[760]&~m[762]&m[763]&m[764])|(m[329]&~m[760]&~m[762]&m[763]&m[764])|(~m[329]&m[760]&~m[762]&m[763]&m[764])|(m[329]&m[760]&~m[762]&m[763]&m[764])|(~m[329]&~m[760]&m[762]&m[763]&m[764])|(m[329]&~m[760]&m[762]&m[763]&m[764])|(m[329]&m[760]&m[762]&m[763]&m[764]))):InitCond[609];
    m[766] = run?((((m[338]&~m[765]&~m[767]&~m[768]&~m[769])|(~m[338]&~m[765]&~m[767]&m[768]&~m[769])|(m[338]&m[765]&~m[767]&m[768]&~m[769])|(m[338]&~m[765]&m[767]&m[768]&~m[769])|(~m[338]&m[765]&~m[767]&~m[768]&m[769])|(~m[338]&~m[765]&m[767]&~m[768]&m[769])|(m[338]&m[765]&m[767]&~m[768]&m[769])|(~m[338]&m[765]&m[767]&m[768]&m[769]))&UnbiasedRNG[271])|((m[338]&~m[765]&~m[767]&m[768]&~m[769])|(~m[338]&~m[765]&~m[767]&~m[768]&m[769])|(m[338]&~m[765]&~m[767]&~m[768]&m[769])|(m[338]&m[765]&~m[767]&~m[768]&m[769])|(m[338]&~m[765]&m[767]&~m[768]&m[769])|(~m[338]&~m[765]&~m[767]&m[768]&m[769])|(m[338]&~m[765]&~m[767]&m[768]&m[769])|(~m[338]&m[765]&~m[767]&m[768]&m[769])|(m[338]&m[765]&~m[767]&m[768]&m[769])|(~m[338]&~m[765]&m[767]&m[768]&m[769])|(m[338]&~m[765]&m[767]&m[768]&m[769])|(m[338]&m[765]&m[767]&m[768]&m[769]))):InitCond[610];
    m[771] = run?((((m[347]&~m[770]&~m[772]&~m[773]&~m[774])|(~m[347]&~m[770]&~m[772]&m[773]&~m[774])|(m[347]&m[770]&~m[772]&m[773]&~m[774])|(m[347]&~m[770]&m[772]&m[773]&~m[774])|(~m[347]&m[770]&~m[772]&~m[773]&m[774])|(~m[347]&~m[770]&m[772]&~m[773]&m[774])|(m[347]&m[770]&m[772]&~m[773]&m[774])|(~m[347]&m[770]&m[772]&m[773]&m[774]))&UnbiasedRNG[272])|((m[347]&~m[770]&~m[772]&m[773]&~m[774])|(~m[347]&~m[770]&~m[772]&~m[773]&m[774])|(m[347]&~m[770]&~m[772]&~m[773]&m[774])|(m[347]&m[770]&~m[772]&~m[773]&m[774])|(m[347]&~m[770]&m[772]&~m[773]&m[774])|(~m[347]&~m[770]&~m[772]&m[773]&m[774])|(m[347]&~m[770]&~m[772]&m[773]&m[774])|(~m[347]&m[770]&~m[772]&m[773]&m[774])|(m[347]&m[770]&~m[772]&m[773]&m[774])|(~m[347]&~m[770]&m[772]&m[773]&m[774])|(m[347]&~m[770]&m[772]&m[773]&m[774])|(m[347]&m[770]&m[772]&m[773]&m[774]))):InitCond[611];
    m[776] = run?((((m[356]&~m[775]&~m[777]&~m[778]&~m[779])|(~m[356]&~m[775]&~m[777]&m[778]&~m[779])|(m[356]&m[775]&~m[777]&m[778]&~m[779])|(m[356]&~m[775]&m[777]&m[778]&~m[779])|(~m[356]&m[775]&~m[777]&~m[778]&m[779])|(~m[356]&~m[775]&m[777]&~m[778]&m[779])|(m[356]&m[775]&m[777]&~m[778]&m[779])|(~m[356]&m[775]&m[777]&m[778]&m[779]))&UnbiasedRNG[273])|((m[356]&~m[775]&~m[777]&m[778]&~m[779])|(~m[356]&~m[775]&~m[777]&~m[778]&m[779])|(m[356]&~m[775]&~m[777]&~m[778]&m[779])|(m[356]&m[775]&~m[777]&~m[778]&m[779])|(m[356]&~m[775]&m[777]&~m[778]&m[779])|(~m[356]&~m[775]&~m[777]&m[778]&m[779])|(m[356]&~m[775]&~m[777]&m[778]&m[779])|(~m[356]&m[775]&~m[777]&m[778]&m[779])|(m[356]&m[775]&~m[777]&m[778]&m[779])|(~m[356]&~m[775]&m[777]&m[778]&m[779])|(m[356]&~m[775]&m[777]&m[778]&m[779])|(m[356]&m[775]&m[777]&m[778]&m[779]))):InitCond[612];
    m[781] = run?((((m[339]&~m[780]&~m[782]&~m[783]&~m[784])|(~m[339]&~m[780]&~m[782]&m[783]&~m[784])|(m[339]&m[780]&~m[782]&m[783]&~m[784])|(m[339]&~m[780]&m[782]&m[783]&~m[784])|(~m[339]&m[780]&~m[782]&~m[783]&m[784])|(~m[339]&~m[780]&m[782]&~m[783]&m[784])|(m[339]&m[780]&m[782]&~m[783]&m[784])|(~m[339]&m[780]&m[782]&m[783]&m[784]))&UnbiasedRNG[274])|((m[339]&~m[780]&~m[782]&m[783]&~m[784])|(~m[339]&~m[780]&~m[782]&~m[783]&m[784])|(m[339]&~m[780]&~m[782]&~m[783]&m[784])|(m[339]&m[780]&~m[782]&~m[783]&m[784])|(m[339]&~m[780]&m[782]&~m[783]&m[784])|(~m[339]&~m[780]&~m[782]&m[783]&m[784])|(m[339]&~m[780]&~m[782]&m[783]&m[784])|(~m[339]&m[780]&~m[782]&m[783]&m[784])|(m[339]&m[780]&~m[782]&m[783]&m[784])|(~m[339]&~m[780]&m[782]&m[783]&m[784])|(m[339]&~m[780]&m[782]&m[783]&m[784])|(m[339]&m[780]&m[782]&m[783]&m[784]))):InitCond[613];
    m[786] = run?((((m[348]&~m[785]&~m[787]&~m[788]&~m[789])|(~m[348]&~m[785]&~m[787]&m[788]&~m[789])|(m[348]&m[785]&~m[787]&m[788]&~m[789])|(m[348]&~m[785]&m[787]&m[788]&~m[789])|(~m[348]&m[785]&~m[787]&~m[788]&m[789])|(~m[348]&~m[785]&m[787]&~m[788]&m[789])|(m[348]&m[785]&m[787]&~m[788]&m[789])|(~m[348]&m[785]&m[787]&m[788]&m[789]))&UnbiasedRNG[275])|((m[348]&~m[785]&~m[787]&m[788]&~m[789])|(~m[348]&~m[785]&~m[787]&~m[788]&m[789])|(m[348]&~m[785]&~m[787]&~m[788]&m[789])|(m[348]&m[785]&~m[787]&~m[788]&m[789])|(m[348]&~m[785]&m[787]&~m[788]&m[789])|(~m[348]&~m[785]&~m[787]&m[788]&m[789])|(m[348]&~m[785]&~m[787]&m[788]&m[789])|(~m[348]&m[785]&~m[787]&m[788]&m[789])|(m[348]&m[785]&~m[787]&m[788]&m[789])|(~m[348]&~m[785]&m[787]&m[788]&m[789])|(m[348]&~m[785]&m[787]&m[788]&m[789])|(m[348]&m[785]&m[787]&m[788]&m[789]))):InitCond[614];
    m[791] = run?((((m[357]&~m[790]&~m[792]&~m[793]&~m[794])|(~m[357]&~m[790]&~m[792]&m[793]&~m[794])|(m[357]&m[790]&~m[792]&m[793]&~m[794])|(m[357]&~m[790]&m[792]&m[793]&~m[794])|(~m[357]&m[790]&~m[792]&~m[793]&m[794])|(~m[357]&~m[790]&m[792]&~m[793]&m[794])|(m[357]&m[790]&m[792]&~m[793]&m[794])|(~m[357]&m[790]&m[792]&m[793]&m[794]))&UnbiasedRNG[276])|((m[357]&~m[790]&~m[792]&m[793]&~m[794])|(~m[357]&~m[790]&~m[792]&~m[793]&m[794])|(m[357]&~m[790]&~m[792]&~m[793]&m[794])|(m[357]&m[790]&~m[792]&~m[793]&m[794])|(m[357]&~m[790]&m[792]&~m[793]&m[794])|(~m[357]&~m[790]&~m[792]&m[793]&m[794])|(m[357]&~m[790]&~m[792]&m[793]&m[794])|(~m[357]&m[790]&~m[792]&m[793]&m[794])|(m[357]&m[790]&~m[792]&m[793]&m[794])|(~m[357]&~m[790]&m[792]&m[793]&m[794])|(m[357]&~m[790]&m[792]&m[793]&m[794])|(m[357]&m[790]&m[792]&m[793]&m[794]))):InitCond[615];
    m[796] = run?((((m[349]&~m[795]&~m[797]&~m[798]&~m[799])|(~m[349]&~m[795]&~m[797]&m[798]&~m[799])|(m[349]&m[795]&~m[797]&m[798]&~m[799])|(m[349]&~m[795]&m[797]&m[798]&~m[799])|(~m[349]&m[795]&~m[797]&~m[798]&m[799])|(~m[349]&~m[795]&m[797]&~m[798]&m[799])|(m[349]&m[795]&m[797]&~m[798]&m[799])|(~m[349]&m[795]&m[797]&m[798]&m[799]))&UnbiasedRNG[277])|((m[349]&~m[795]&~m[797]&m[798]&~m[799])|(~m[349]&~m[795]&~m[797]&~m[798]&m[799])|(m[349]&~m[795]&~m[797]&~m[798]&m[799])|(m[349]&m[795]&~m[797]&~m[798]&m[799])|(m[349]&~m[795]&m[797]&~m[798]&m[799])|(~m[349]&~m[795]&~m[797]&m[798]&m[799])|(m[349]&~m[795]&~m[797]&m[798]&m[799])|(~m[349]&m[795]&~m[797]&m[798]&m[799])|(m[349]&m[795]&~m[797]&m[798]&m[799])|(~m[349]&~m[795]&m[797]&m[798]&m[799])|(m[349]&~m[795]&m[797]&m[798]&m[799])|(m[349]&m[795]&m[797]&m[798]&m[799]))):InitCond[616];
    m[801] = run?((((m[358]&~m[800]&~m[802]&~m[803]&~m[804])|(~m[358]&~m[800]&~m[802]&m[803]&~m[804])|(m[358]&m[800]&~m[802]&m[803]&~m[804])|(m[358]&~m[800]&m[802]&m[803]&~m[804])|(~m[358]&m[800]&~m[802]&~m[803]&m[804])|(~m[358]&~m[800]&m[802]&~m[803]&m[804])|(m[358]&m[800]&m[802]&~m[803]&m[804])|(~m[358]&m[800]&m[802]&m[803]&m[804]))&UnbiasedRNG[278])|((m[358]&~m[800]&~m[802]&m[803]&~m[804])|(~m[358]&~m[800]&~m[802]&~m[803]&m[804])|(m[358]&~m[800]&~m[802]&~m[803]&m[804])|(m[358]&m[800]&~m[802]&~m[803]&m[804])|(m[358]&~m[800]&m[802]&~m[803]&m[804])|(~m[358]&~m[800]&~m[802]&m[803]&m[804])|(m[358]&~m[800]&~m[802]&m[803]&m[804])|(~m[358]&m[800]&~m[802]&m[803]&m[804])|(m[358]&m[800]&~m[802]&m[803]&m[804])|(~m[358]&~m[800]&m[802]&m[803]&m[804])|(m[358]&~m[800]&m[802]&m[803]&m[804])|(m[358]&m[800]&m[802]&m[803]&m[804]))):InitCond[617];
    m[806] = run?((((m[359]&~m[805]&~m[807]&~m[808]&~m[809])|(~m[359]&~m[805]&~m[807]&m[808]&~m[809])|(m[359]&m[805]&~m[807]&m[808]&~m[809])|(m[359]&~m[805]&m[807]&m[808]&~m[809])|(~m[359]&m[805]&~m[807]&~m[808]&m[809])|(~m[359]&~m[805]&m[807]&~m[808]&m[809])|(m[359]&m[805]&m[807]&~m[808]&m[809])|(~m[359]&m[805]&m[807]&m[808]&m[809]))&UnbiasedRNG[279])|((m[359]&~m[805]&~m[807]&m[808]&~m[809])|(~m[359]&~m[805]&~m[807]&~m[808]&m[809])|(m[359]&~m[805]&~m[807]&~m[808]&m[809])|(m[359]&m[805]&~m[807]&~m[808]&m[809])|(m[359]&~m[805]&m[807]&~m[808]&m[809])|(~m[359]&~m[805]&~m[807]&m[808]&m[809])|(m[359]&~m[805]&~m[807]&m[808]&m[809])|(~m[359]&m[805]&~m[807]&m[808]&m[809])|(m[359]&m[805]&~m[807]&m[808]&m[809])|(~m[359]&~m[805]&m[807]&m[808]&m[809])|(m[359]&~m[805]&m[807]&m[808]&m[809])|(m[359]&m[805]&m[807]&m[808]&m[809]))):InitCond[618];
end

always @(posedge color3_clk) begin
    m[368] = run?((((m[365]&~m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&~m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&m[369]&~m[370])|(~m[365]&~m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&m[369]&m[370])|(m[365]&~m[366]&m[367]&m[369]&m[370])|(~m[365]&m[366]&m[367]&m[369]&m[370]))&UnbiasedRNG[280])|((m[365]&m[366]&~m[367]&~m[369]&~m[370])|(m[365]&~m[366]&m[367]&~m[369]&~m[370])|(~m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&~m[366]&~m[367]&~m[369]&m[370])|(~m[365]&m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&~m[369]&m[370])|(~m[365]&~m[366]&m[367]&~m[369]&m[370])|(m[365]&~m[366]&m[367]&~m[369]&m[370])|(~m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&m[369]&m[370]))):InitCond[619];
    m[378] = run?((((m[375]&~m[376]&~m[377]&~m[379]&~m[380])|(~m[375]&m[376]&~m[377]&~m[379]&~m[380])|(~m[375]&~m[376]&m[377]&~m[379]&~m[380])|(m[375]&m[376]&m[377]&m[379]&~m[380])|(~m[375]&~m[376]&~m[377]&~m[379]&m[380])|(m[375]&m[376]&~m[377]&m[379]&m[380])|(m[375]&~m[376]&m[377]&m[379]&m[380])|(~m[375]&m[376]&m[377]&m[379]&m[380]))&UnbiasedRNG[281])|((m[375]&m[376]&~m[377]&~m[379]&~m[380])|(m[375]&~m[376]&m[377]&~m[379]&~m[380])|(~m[375]&m[376]&m[377]&~m[379]&~m[380])|(m[375]&m[376]&m[377]&~m[379]&~m[380])|(m[375]&~m[376]&~m[377]&~m[379]&m[380])|(~m[375]&m[376]&~m[377]&~m[379]&m[380])|(m[375]&m[376]&~m[377]&~m[379]&m[380])|(~m[375]&~m[376]&m[377]&~m[379]&m[380])|(m[375]&~m[376]&m[377]&~m[379]&m[380])|(~m[375]&m[376]&m[377]&~m[379]&m[380])|(m[375]&m[376]&m[377]&~m[379]&m[380])|(m[375]&m[376]&m[377]&m[379]&m[380]))):InitCond[620];
    m[383] = run?((((m[380]&~m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&~m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&m[384]&~m[385])|(~m[380]&~m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&m[384]&m[385])|(m[380]&~m[381]&m[382]&m[384]&m[385])|(~m[380]&m[381]&m[382]&m[384]&m[385]))&UnbiasedRNG[282])|((m[380]&m[381]&~m[382]&~m[384]&~m[385])|(m[380]&~m[381]&m[382]&~m[384]&~m[385])|(~m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&~m[381]&~m[382]&~m[384]&m[385])|(~m[380]&m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&~m[384]&m[385])|(~m[380]&~m[381]&m[382]&~m[384]&m[385])|(m[380]&~m[381]&m[382]&~m[384]&m[385])|(~m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&m[384]&m[385]))):InitCond[621];
    m[393] = run?((((m[390]&~m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&~m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&m[394]&~m[395])|(~m[390]&~m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&m[394]&m[395])|(m[390]&~m[391]&m[392]&m[394]&m[395])|(~m[390]&m[391]&m[392]&m[394]&m[395]))&UnbiasedRNG[283])|((m[390]&m[391]&~m[392]&~m[394]&~m[395])|(m[390]&~m[391]&m[392]&~m[394]&~m[395])|(~m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&~m[391]&~m[392]&~m[394]&m[395])|(~m[390]&m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&~m[394]&m[395])|(~m[390]&~m[391]&m[392]&~m[394]&m[395])|(m[390]&~m[391]&m[392]&~m[394]&m[395])|(~m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&m[394]&m[395]))):InitCond[622];
    m[398] = run?((((m[395]&~m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&~m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&m[399]&~m[400])|(~m[395]&~m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&m[399]&m[400])|(m[395]&~m[396]&m[397]&m[399]&m[400])|(~m[395]&m[396]&m[397]&m[399]&m[400]))&UnbiasedRNG[284])|((m[395]&m[396]&~m[397]&~m[399]&~m[400])|(m[395]&~m[396]&m[397]&~m[399]&~m[400])|(~m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&~m[396]&~m[397]&~m[399]&m[400])|(~m[395]&m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&~m[399]&m[400])|(~m[395]&~m[396]&m[397]&~m[399]&m[400])|(m[395]&~m[396]&m[397]&~m[399]&m[400])|(~m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&m[399]&m[400]))):InitCond[623];
    m[403] = run?((((m[400]&~m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&~m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&m[404]&~m[405])|(~m[400]&~m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&m[404]&m[405])|(m[400]&~m[401]&m[402]&m[404]&m[405])|(~m[400]&m[401]&m[402]&m[404]&m[405]))&UnbiasedRNG[285])|((m[400]&m[401]&~m[402]&~m[404]&~m[405])|(m[400]&~m[401]&m[402]&~m[404]&~m[405])|(~m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&~m[401]&~m[402]&~m[404]&m[405])|(~m[400]&m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&~m[404]&m[405])|(~m[400]&~m[401]&m[402]&~m[404]&m[405])|(m[400]&~m[401]&m[402]&~m[404]&m[405])|(~m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&m[404]&m[405]))):InitCond[624];
    m[413] = run?((((m[410]&~m[411]&~m[412]&~m[414]&~m[415])|(~m[410]&m[411]&~m[412]&~m[414]&~m[415])|(~m[410]&~m[411]&m[412]&~m[414]&~m[415])|(m[410]&m[411]&m[412]&m[414]&~m[415])|(~m[410]&~m[411]&~m[412]&~m[414]&m[415])|(m[410]&m[411]&~m[412]&m[414]&m[415])|(m[410]&~m[411]&m[412]&m[414]&m[415])|(~m[410]&m[411]&m[412]&m[414]&m[415]))&UnbiasedRNG[286])|((m[410]&m[411]&~m[412]&~m[414]&~m[415])|(m[410]&~m[411]&m[412]&~m[414]&~m[415])|(~m[410]&m[411]&m[412]&~m[414]&~m[415])|(m[410]&m[411]&m[412]&~m[414]&~m[415])|(m[410]&~m[411]&~m[412]&~m[414]&m[415])|(~m[410]&m[411]&~m[412]&~m[414]&m[415])|(m[410]&m[411]&~m[412]&~m[414]&m[415])|(~m[410]&~m[411]&m[412]&~m[414]&m[415])|(m[410]&~m[411]&m[412]&~m[414]&m[415])|(~m[410]&m[411]&m[412]&~m[414]&m[415])|(m[410]&m[411]&m[412]&~m[414]&m[415])|(m[410]&m[411]&m[412]&m[414]&m[415]))):InitCond[625];
    m[418] = run?((((m[415]&~m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&~m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&m[419]&~m[420])|(~m[415]&~m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&m[419]&m[420])|(m[415]&~m[416]&m[417]&m[419]&m[420])|(~m[415]&m[416]&m[417]&m[419]&m[420]))&UnbiasedRNG[287])|((m[415]&m[416]&~m[417]&~m[419]&~m[420])|(m[415]&~m[416]&m[417]&~m[419]&~m[420])|(~m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&~m[416]&~m[417]&~m[419]&m[420])|(~m[415]&m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&~m[419]&m[420])|(~m[415]&~m[416]&m[417]&~m[419]&m[420])|(m[415]&~m[416]&m[417]&~m[419]&m[420])|(~m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&m[419]&m[420]))):InitCond[626];
    m[423] = run?((((m[420]&~m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&~m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&m[424]&~m[425])|(~m[420]&~m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&m[424]&m[425])|(m[420]&~m[421]&m[422]&m[424]&m[425])|(~m[420]&m[421]&m[422]&m[424]&m[425]))&UnbiasedRNG[288])|((m[420]&m[421]&~m[422]&~m[424]&~m[425])|(m[420]&~m[421]&m[422]&~m[424]&~m[425])|(~m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&~m[421]&~m[422]&~m[424]&m[425])|(~m[420]&m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&~m[424]&m[425])|(~m[420]&~m[421]&m[422]&~m[424]&m[425])|(m[420]&~m[421]&m[422]&~m[424]&m[425])|(~m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&m[424]&m[425]))):InitCond[627];
    m[428] = run?((((m[425]&~m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&~m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&m[429]&~m[430])|(~m[425]&~m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&m[429]&m[430])|(m[425]&~m[426]&m[427]&m[429]&m[430])|(~m[425]&m[426]&m[427]&m[429]&m[430]))&UnbiasedRNG[289])|((m[425]&m[426]&~m[427]&~m[429]&~m[430])|(m[425]&~m[426]&m[427]&~m[429]&~m[430])|(~m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&~m[426]&~m[427]&~m[429]&m[430])|(~m[425]&m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&~m[429]&m[430])|(~m[425]&~m[426]&m[427]&~m[429]&m[430])|(m[425]&~m[426]&m[427]&~m[429]&m[430])|(~m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&m[429]&m[430]))):InitCond[628];
    m[438] = run?((((m[435]&~m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&~m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&m[439]&~m[440])|(~m[435]&~m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&m[439]&m[440])|(m[435]&~m[436]&m[437]&m[439]&m[440])|(~m[435]&m[436]&m[437]&m[439]&m[440]))&UnbiasedRNG[290])|((m[435]&m[436]&~m[437]&~m[439]&~m[440])|(m[435]&~m[436]&m[437]&~m[439]&~m[440])|(~m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&~m[436]&~m[437]&~m[439]&m[440])|(~m[435]&m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&~m[439]&m[440])|(~m[435]&~m[436]&m[437]&~m[439]&m[440])|(m[435]&~m[436]&m[437]&~m[439]&m[440])|(~m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&m[439]&m[440]))):InitCond[629];
    m[443] = run?((((m[440]&~m[441]&~m[442]&~m[444]&~m[445])|(~m[440]&m[441]&~m[442]&~m[444]&~m[445])|(~m[440]&~m[441]&m[442]&~m[444]&~m[445])|(m[440]&m[441]&m[442]&m[444]&~m[445])|(~m[440]&~m[441]&~m[442]&~m[444]&m[445])|(m[440]&m[441]&~m[442]&m[444]&m[445])|(m[440]&~m[441]&m[442]&m[444]&m[445])|(~m[440]&m[441]&m[442]&m[444]&m[445]))&UnbiasedRNG[291])|((m[440]&m[441]&~m[442]&~m[444]&~m[445])|(m[440]&~m[441]&m[442]&~m[444]&~m[445])|(~m[440]&m[441]&m[442]&~m[444]&~m[445])|(m[440]&m[441]&m[442]&~m[444]&~m[445])|(m[440]&~m[441]&~m[442]&~m[444]&m[445])|(~m[440]&m[441]&~m[442]&~m[444]&m[445])|(m[440]&m[441]&~m[442]&~m[444]&m[445])|(~m[440]&~m[441]&m[442]&~m[444]&m[445])|(m[440]&~m[441]&m[442]&~m[444]&m[445])|(~m[440]&m[441]&m[442]&~m[444]&m[445])|(m[440]&m[441]&m[442]&~m[444]&m[445])|(m[440]&m[441]&m[442]&m[444]&m[445]))):InitCond[630];
    m[448] = run?((((m[445]&~m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&~m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&m[449]&~m[450])|(~m[445]&~m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&m[449]&m[450])|(m[445]&~m[446]&m[447]&m[449]&m[450])|(~m[445]&m[446]&m[447]&m[449]&m[450]))&UnbiasedRNG[292])|((m[445]&m[446]&~m[447]&~m[449]&~m[450])|(m[445]&~m[446]&m[447]&~m[449]&~m[450])|(~m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&~m[446]&~m[447]&~m[449]&m[450])|(~m[445]&m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&~m[449]&m[450])|(~m[445]&~m[446]&m[447]&~m[449]&m[450])|(m[445]&~m[446]&m[447]&~m[449]&m[450])|(~m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&m[449]&m[450]))):InitCond[631];
    m[453] = run?((((m[450]&~m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&~m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&m[454]&~m[455])|(~m[450]&~m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&m[454]&m[455])|(m[450]&~m[451]&m[452]&m[454]&m[455])|(~m[450]&m[451]&m[452]&m[454]&m[455]))&UnbiasedRNG[293])|((m[450]&m[451]&~m[452]&~m[454]&~m[455])|(m[450]&~m[451]&m[452]&~m[454]&~m[455])|(~m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&~m[451]&~m[452]&~m[454]&m[455])|(~m[450]&m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&~m[454]&m[455])|(~m[450]&~m[451]&m[452]&~m[454]&m[455])|(m[450]&~m[451]&m[452]&~m[454]&m[455])|(~m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&m[454]&m[455]))):InitCond[632];
    m[458] = run?((((m[455]&~m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&~m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&m[459]&~m[460])|(~m[455]&~m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&m[459]&m[460])|(m[455]&~m[456]&m[457]&m[459]&m[460])|(~m[455]&m[456]&m[457]&m[459]&m[460]))&UnbiasedRNG[294])|((m[455]&m[456]&~m[457]&~m[459]&~m[460])|(m[455]&~m[456]&m[457]&~m[459]&~m[460])|(~m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&~m[456]&~m[457]&~m[459]&m[460])|(~m[455]&m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&~m[459]&m[460])|(~m[455]&~m[456]&m[457]&~m[459]&m[460])|(m[455]&~m[456]&m[457]&~m[459]&m[460])|(~m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&m[459]&m[460]))):InitCond[633];
    m[468] = run?((((m[465]&~m[466]&~m[467]&~m[469]&~m[470])|(~m[465]&m[466]&~m[467]&~m[469]&~m[470])|(~m[465]&~m[466]&m[467]&~m[469]&~m[470])|(m[465]&m[466]&m[467]&m[469]&~m[470])|(~m[465]&~m[466]&~m[467]&~m[469]&m[470])|(m[465]&m[466]&~m[467]&m[469]&m[470])|(m[465]&~m[466]&m[467]&m[469]&m[470])|(~m[465]&m[466]&m[467]&m[469]&m[470]))&UnbiasedRNG[295])|((m[465]&m[466]&~m[467]&~m[469]&~m[470])|(m[465]&~m[466]&m[467]&~m[469]&~m[470])|(~m[465]&m[466]&m[467]&~m[469]&~m[470])|(m[465]&m[466]&m[467]&~m[469]&~m[470])|(m[465]&~m[466]&~m[467]&~m[469]&m[470])|(~m[465]&m[466]&~m[467]&~m[469]&m[470])|(m[465]&m[466]&~m[467]&~m[469]&m[470])|(~m[465]&~m[466]&m[467]&~m[469]&m[470])|(m[465]&~m[466]&m[467]&~m[469]&m[470])|(~m[465]&m[466]&m[467]&~m[469]&m[470])|(m[465]&m[466]&m[467]&~m[469]&m[470])|(m[465]&m[466]&m[467]&m[469]&m[470]))):InitCond[634];
    m[473] = run?((((m[470]&~m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&~m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&m[474]&~m[475])|(~m[470]&~m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&m[474]&m[475])|(m[470]&~m[471]&m[472]&m[474]&m[475])|(~m[470]&m[471]&m[472]&m[474]&m[475]))&UnbiasedRNG[296])|((m[470]&m[471]&~m[472]&~m[474]&~m[475])|(m[470]&~m[471]&m[472]&~m[474]&~m[475])|(~m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&~m[471]&~m[472]&~m[474]&m[475])|(~m[470]&m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&~m[474]&m[475])|(~m[470]&~m[471]&m[472]&~m[474]&m[475])|(m[470]&~m[471]&m[472]&~m[474]&m[475])|(~m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&m[474]&m[475]))):InitCond[635];
    m[478] = run?((((m[475]&~m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&~m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&m[479]&~m[480])|(~m[475]&~m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&m[479]&m[480])|(m[475]&~m[476]&m[477]&m[479]&m[480])|(~m[475]&m[476]&m[477]&m[479]&m[480]))&UnbiasedRNG[297])|((m[475]&m[476]&~m[477]&~m[479]&~m[480])|(m[475]&~m[476]&m[477]&~m[479]&~m[480])|(~m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&~m[476]&~m[477]&~m[479]&m[480])|(~m[475]&m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&~m[479]&m[480])|(~m[475]&~m[476]&m[477]&~m[479]&m[480])|(m[475]&~m[476]&m[477]&~m[479]&m[480])|(~m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&m[479]&m[480]))):InitCond[636];
    m[483] = run?((((m[480]&~m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&~m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&m[484]&~m[485])|(~m[480]&~m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&m[484]&m[485])|(m[480]&~m[481]&m[482]&m[484]&m[485])|(~m[480]&m[481]&m[482]&m[484]&m[485]))&UnbiasedRNG[298])|((m[480]&m[481]&~m[482]&~m[484]&~m[485])|(m[480]&~m[481]&m[482]&~m[484]&~m[485])|(~m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&~m[481]&~m[482]&~m[484]&m[485])|(~m[480]&m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&~m[484]&m[485])|(~m[480]&~m[481]&m[482]&~m[484]&m[485])|(m[480]&~m[481]&m[482]&~m[484]&m[485])|(~m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&m[484]&m[485]))):InitCond[637];
    m[488] = run?((((m[485]&~m[486]&~m[487]&~m[489]&~m[490])|(~m[485]&m[486]&~m[487]&~m[489]&~m[490])|(~m[485]&~m[486]&m[487]&~m[489]&~m[490])|(m[485]&m[486]&m[487]&m[489]&~m[490])|(~m[485]&~m[486]&~m[487]&~m[489]&m[490])|(m[485]&m[486]&~m[487]&m[489]&m[490])|(m[485]&~m[486]&m[487]&m[489]&m[490])|(~m[485]&m[486]&m[487]&m[489]&m[490]))&UnbiasedRNG[299])|((m[485]&m[486]&~m[487]&~m[489]&~m[490])|(m[485]&~m[486]&m[487]&~m[489]&~m[490])|(~m[485]&m[486]&m[487]&~m[489]&~m[490])|(m[485]&m[486]&m[487]&~m[489]&~m[490])|(m[485]&~m[486]&~m[487]&~m[489]&m[490])|(~m[485]&m[486]&~m[487]&~m[489]&m[490])|(m[485]&m[486]&~m[487]&~m[489]&m[490])|(~m[485]&~m[486]&m[487]&~m[489]&m[490])|(m[485]&~m[486]&m[487]&~m[489]&m[490])|(~m[485]&m[486]&m[487]&~m[489]&m[490])|(m[485]&m[486]&m[487]&~m[489]&m[490])|(m[485]&m[486]&m[487]&m[489]&m[490]))):InitCond[638];
    m[493] = run?((((m[490]&~m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&~m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&m[494]&~m[495])|(~m[490]&~m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&m[494]&m[495])|(m[490]&~m[491]&m[492]&m[494]&m[495])|(~m[490]&m[491]&m[492]&m[494]&m[495]))&UnbiasedRNG[300])|((m[490]&m[491]&~m[492]&~m[494]&~m[495])|(m[490]&~m[491]&m[492]&~m[494]&~m[495])|(~m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&~m[491]&~m[492]&~m[494]&m[495])|(~m[490]&m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&~m[494]&m[495])|(~m[490]&~m[491]&m[492]&~m[494]&m[495])|(m[490]&~m[491]&m[492]&~m[494]&m[495])|(~m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&m[494]&m[495]))):InitCond[639];
    m[503] = run?((((m[500]&~m[501]&~m[502]&~m[504]&~m[505])|(~m[500]&m[501]&~m[502]&~m[504]&~m[505])|(~m[500]&~m[501]&m[502]&~m[504]&~m[505])|(m[500]&m[501]&m[502]&m[504]&~m[505])|(~m[500]&~m[501]&~m[502]&~m[504]&m[505])|(m[500]&m[501]&~m[502]&m[504]&m[505])|(m[500]&~m[501]&m[502]&m[504]&m[505])|(~m[500]&m[501]&m[502]&m[504]&m[505]))&UnbiasedRNG[301])|((m[500]&m[501]&~m[502]&~m[504]&~m[505])|(m[500]&~m[501]&m[502]&~m[504]&~m[505])|(~m[500]&m[501]&m[502]&~m[504]&~m[505])|(m[500]&m[501]&m[502]&~m[504]&~m[505])|(m[500]&~m[501]&~m[502]&~m[504]&m[505])|(~m[500]&m[501]&~m[502]&~m[504]&m[505])|(m[500]&m[501]&~m[502]&~m[504]&m[505])|(~m[500]&~m[501]&m[502]&~m[504]&m[505])|(m[500]&~m[501]&m[502]&~m[504]&m[505])|(~m[500]&m[501]&m[502]&~m[504]&m[505])|(m[500]&m[501]&m[502]&~m[504]&m[505])|(m[500]&m[501]&m[502]&m[504]&m[505]))):InitCond[640];
    m[508] = run?((((m[505]&~m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&~m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&m[509]&~m[510])|(~m[505]&~m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&m[509]&m[510])|(m[505]&~m[506]&m[507]&m[509]&m[510])|(~m[505]&m[506]&m[507]&m[509]&m[510]))&UnbiasedRNG[302])|((m[505]&m[506]&~m[507]&~m[509]&~m[510])|(m[505]&~m[506]&m[507]&~m[509]&~m[510])|(~m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&~m[506]&~m[507]&~m[509]&m[510])|(~m[505]&m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&~m[509]&m[510])|(~m[505]&~m[506]&m[507]&~m[509]&m[510])|(m[505]&~m[506]&m[507]&~m[509]&m[510])|(~m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&m[509]&m[510]))):InitCond[641];
    m[513] = run?((((m[510]&~m[511]&~m[512]&~m[514]&~m[515])|(~m[510]&m[511]&~m[512]&~m[514]&~m[515])|(~m[510]&~m[511]&m[512]&~m[514]&~m[515])|(m[510]&m[511]&m[512]&m[514]&~m[515])|(~m[510]&~m[511]&~m[512]&~m[514]&m[515])|(m[510]&m[511]&~m[512]&m[514]&m[515])|(m[510]&~m[511]&m[512]&m[514]&m[515])|(~m[510]&m[511]&m[512]&m[514]&m[515]))&UnbiasedRNG[303])|((m[510]&m[511]&~m[512]&~m[514]&~m[515])|(m[510]&~m[511]&m[512]&~m[514]&~m[515])|(~m[510]&m[511]&m[512]&~m[514]&~m[515])|(m[510]&m[511]&m[512]&~m[514]&~m[515])|(m[510]&~m[511]&~m[512]&~m[514]&m[515])|(~m[510]&m[511]&~m[512]&~m[514]&m[515])|(m[510]&m[511]&~m[512]&~m[514]&m[515])|(~m[510]&~m[511]&m[512]&~m[514]&m[515])|(m[510]&~m[511]&m[512]&~m[514]&m[515])|(~m[510]&m[511]&m[512]&~m[514]&m[515])|(m[510]&m[511]&m[512]&~m[514]&m[515])|(m[510]&m[511]&m[512]&m[514]&m[515]))):InitCond[642];
    m[518] = run?((((m[515]&~m[516]&~m[517]&~m[519]&~m[520])|(~m[515]&m[516]&~m[517]&~m[519]&~m[520])|(~m[515]&~m[516]&m[517]&~m[519]&~m[520])|(m[515]&m[516]&m[517]&m[519]&~m[520])|(~m[515]&~m[516]&~m[517]&~m[519]&m[520])|(m[515]&m[516]&~m[517]&m[519]&m[520])|(m[515]&~m[516]&m[517]&m[519]&m[520])|(~m[515]&m[516]&m[517]&m[519]&m[520]))&UnbiasedRNG[304])|((m[515]&m[516]&~m[517]&~m[519]&~m[520])|(m[515]&~m[516]&m[517]&~m[519]&~m[520])|(~m[515]&m[516]&m[517]&~m[519]&~m[520])|(m[515]&m[516]&m[517]&~m[519]&~m[520])|(m[515]&~m[516]&~m[517]&~m[519]&m[520])|(~m[515]&m[516]&~m[517]&~m[519]&m[520])|(m[515]&m[516]&~m[517]&~m[519]&m[520])|(~m[515]&~m[516]&m[517]&~m[519]&m[520])|(m[515]&~m[516]&m[517]&~m[519]&m[520])|(~m[515]&m[516]&m[517]&~m[519]&m[520])|(m[515]&m[516]&m[517]&~m[519]&m[520])|(m[515]&m[516]&m[517]&m[519]&m[520]))):InitCond[643];
    m[523] = run?((((m[520]&~m[521]&~m[522]&~m[524]&~m[525])|(~m[520]&m[521]&~m[522]&~m[524]&~m[525])|(~m[520]&~m[521]&m[522]&~m[524]&~m[525])|(m[520]&m[521]&m[522]&m[524]&~m[525])|(~m[520]&~m[521]&~m[522]&~m[524]&m[525])|(m[520]&m[521]&~m[522]&m[524]&m[525])|(m[520]&~m[521]&m[522]&m[524]&m[525])|(~m[520]&m[521]&m[522]&m[524]&m[525]))&UnbiasedRNG[305])|((m[520]&m[521]&~m[522]&~m[524]&~m[525])|(m[520]&~m[521]&m[522]&~m[524]&~m[525])|(~m[520]&m[521]&m[522]&~m[524]&~m[525])|(m[520]&m[521]&m[522]&~m[524]&~m[525])|(m[520]&~m[521]&~m[522]&~m[524]&m[525])|(~m[520]&m[521]&~m[522]&~m[524]&m[525])|(m[520]&m[521]&~m[522]&~m[524]&m[525])|(~m[520]&~m[521]&m[522]&~m[524]&m[525])|(m[520]&~m[521]&m[522]&~m[524]&m[525])|(~m[520]&m[521]&m[522]&~m[524]&m[525])|(m[520]&m[521]&m[522]&~m[524]&m[525])|(m[520]&m[521]&m[522]&m[524]&m[525]))):InitCond[644];
    m[528] = run?((((m[525]&~m[526]&~m[527]&~m[529]&~m[530])|(~m[525]&m[526]&~m[527]&~m[529]&~m[530])|(~m[525]&~m[526]&m[527]&~m[529]&~m[530])|(m[525]&m[526]&m[527]&m[529]&~m[530])|(~m[525]&~m[526]&~m[527]&~m[529]&m[530])|(m[525]&m[526]&~m[527]&m[529]&m[530])|(m[525]&~m[526]&m[527]&m[529]&m[530])|(~m[525]&m[526]&m[527]&m[529]&m[530]))&UnbiasedRNG[306])|((m[525]&m[526]&~m[527]&~m[529]&~m[530])|(m[525]&~m[526]&m[527]&~m[529]&~m[530])|(~m[525]&m[526]&m[527]&~m[529]&~m[530])|(m[525]&m[526]&m[527]&~m[529]&~m[530])|(m[525]&~m[526]&~m[527]&~m[529]&m[530])|(~m[525]&m[526]&~m[527]&~m[529]&m[530])|(m[525]&m[526]&~m[527]&~m[529]&m[530])|(~m[525]&~m[526]&m[527]&~m[529]&m[530])|(m[525]&~m[526]&m[527]&~m[529]&m[530])|(~m[525]&m[526]&m[527]&~m[529]&m[530])|(m[525]&m[526]&m[527]&~m[529]&m[530])|(m[525]&m[526]&m[527]&m[529]&m[530]))):InitCond[645];
    m[533] = run?((((m[530]&~m[531]&~m[532]&~m[534]&~m[535])|(~m[530]&m[531]&~m[532]&~m[534]&~m[535])|(~m[530]&~m[531]&m[532]&~m[534]&~m[535])|(m[530]&m[531]&m[532]&m[534]&~m[535])|(~m[530]&~m[531]&~m[532]&~m[534]&m[535])|(m[530]&m[531]&~m[532]&m[534]&m[535])|(m[530]&~m[531]&m[532]&m[534]&m[535])|(~m[530]&m[531]&m[532]&m[534]&m[535]))&UnbiasedRNG[307])|((m[530]&m[531]&~m[532]&~m[534]&~m[535])|(m[530]&~m[531]&m[532]&~m[534]&~m[535])|(~m[530]&m[531]&m[532]&~m[534]&~m[535])|(m[530]&m[531]&m[532]&~m[534]&~m[535])|(m[530]&~m[531]&~m[532]&~m[534]&m[535])|(~m[530]&m[531]&~m[532]&~m[534]&m[535])|(m[530]&m[531]&~m[532]&~m[534]&m[535])|(~m[530]&~m[531]&m[532]&~m[534]&m[535])|(m[530]&~m[531]&m[532]&~m[534]&m[535])|(~m[530]&m[531]&m[532]&~m[534]&m[535])|(m[530]&m[531]&m[532]&~m[534]&m[535])|(m[530]&m[531]&m[532]&m[534]&m[535]))):InitCond[646];
    m[543] = run?((((m[540]&~m[541]&~m[542]&~m[544]&~m[545])|(~m[540]&m[541]&~m[542]&~m[544]&~m[545])|(~m[540]&~m[541]&m[542]&~m[544]&~m[545])|(m[540]&m[541]&m[542]&m[544]&~m[545])|(~m[540]&~m[541]&~m[542]&~m[544]&m[545])|(m[540]&m[541]&~m[542]&m[544]&m[545])|(m[540]&~m[541]&m[542]&m[544]&m[545])|(~m[540]&m[541]&m[542]&m[544]&m[545]))&UnbiasedRNG[308])|((m[540]&m[541]&~m[542]&~m[544]&~m[545])|(m[540]&~m[541]&m[542]&~m[544]&~m[545])|(~m[540]&m[541]&m[542]&~m[544]&~m[545])|(m[540]&m[541]&m[542]&~m[544]&~m[545])|(m[540]&~m[541]&~m[542]&~m[544]&m[545])|(~m[540]&m[541]&~m[542]&~m[544]&m[545])|(m[540]&m[541]&~m[542]&~m[544]&m[545])|(~m[540]&~m[541]&m[542]&~m[544]&m[545])|(m[540]&~m[541]&m[542]&~m[544]&m[545])|(~m[540]&m[541]&m[542]&~m[544]&m[545])|(m[540]&m[541]&m[542]&~m[544]&m[545])|(m[540]&m[541]&m[542]&m[544]&m[545]))):InitCond[647];
    m[548] = run?((((m[545]&~m[546]&~m[547]&~m[549]&~m[550])|(~m[545]&m[546]&~m[547]&~m[549]&~m[550])|(~m[545]&~m[546]&m[547]&~m[549]&~m[550])|(m[545]&m[546]&m[547]&m[549]&~m[550])|(~m[545]&~m[546]&~m[547]&~m[549]&m[550])|(m[545]&m[546]&~m[547]&m[549]&m[550])|(m[545]&~m[546]&m[547]&m[549]&m[550])|(~m[545]&m[546]&m[547]&m[549]&m[550]))&UnbiasedRNG[309])|((m[545]&m[546]&~m[547]&~m[549]&~m[550])|(m[545]&~m[546]&m[547]&~m[549]&~m[550])|(~m[545]&m[546]&m[547]&~m[549]&~m[550])|(m[545]&m[546]&m[547]&~m[549]&~m[550])|(m[545]&~m[546]&~m[547]&~m[549]&m[550])|(~m[545]&m[546]&~m[547]&~m[549]&m[550])|(m[545]&m[546]&~m[547]&~m[549]&m[550])|(~m[545]&~m[546]&m[547]&~m[549]&m[550])|(m[545]&~m[546]&m[547]&~m[549]&m[550])|(~m[545]&m[546]&m[547]&~m[549]&m[550])|(m[545]&m[546]&m[547]&~m[549]&m[550])|(m[545]&m[546]&m[547]&m[549]&m[550]))):InitCond[648];
    m[553] = run?((((m[550]&~m[551]&~m[552]&~m[554]&~m[555])|(~m[550]&m[551]&~m[552]&~m[554]&~m[555])|(~m[550]&~m[551]&m[552]&~m[554]&~m[555])|(m[550]&m[551]&m[552]&m[554]&~m[555])|(~m[550]&~m[551]&~m[552]&~m[554]&m[555])|(m[550]&m[551]&~m[552]&m[554]&m[555])|(m[550]&~m[551]&m[552]&m[554]&m[555])|(~m[550]&m[551]&m[552]&m[554]&m[555]))&UnbiasedRNG[310])|((m[550]&m[551]&~m[552]&~m[554]&~m[555])|(m[550]&~m[551]&m[552]&~m[554]&~m[555])|(~m[550]&m[551]&m[552]&~m[554]&~m[555])|(m[550]&m[551]&m[552]&~m[554]&~m[555])|(m[550]&~m[551]&~m[552]&~m[554]&m[555])|(~m[550]&m[551]&~m[552]&~m[554]&m[555])|(m[550]&m[551]&~m[552]&~m[554]&m[555])|(~m[550]&~m[551]&m[552]&~m[554]&m[555])|(m[550]&~m[551]&m[552]&~m[554]&m[555])|(~m[550]&m[551]&m[552]&~m[554]&m[555])|(m[550]&m[551]&m[552]&~m[554]&m[555])|(m[550]&m[551]&m[552]&m[554]&m[555]))):InitCond[649];
    m[558] = run?((((m[555]&~m[556]&~m[557]&~m[559]&~m[560])|(~m[555]&m[556]&~m[557]&~m[559]&~m[560])|(~m[555]&~m[556]&m[557]&~m[559]&~m[560])|(m[555]&m[556]&m[557]&m[559]&~m[560])|(~m[555]&~m[556]&~m[557]&~m[559]&m[560])|(m[555]&m[556]&~m[557]&m[559]&m[560])|(m[555]&~m[556]&m[557]&m[559]&m[560])|(~m[555]&m[556]&m[557]&m[559]&m[560]))&UnbiasedRNG[311])|((m[555]&m[556]&~m[557]&~m[559]&~m[560])|(m[555]&~m[556]&m[557]&~m[559]&~m[560])|(~m[555]&m[556]&m[557]&~m[559]&~m[560])|(m[555]&m[556]&m[557]&~m[559]&~m[560])|(m[555]&~m[556]&~m[557]&~m[559]&m[560])|(~m[555]&m[556]&~m[557]&~m[559]&m[560])|(m[555]&m[556]&~m[557]&~m[559]&m[560])|(~m[555]&~m[556]&m[557]&~m[559]&m[560])|(m[555]&~m[556]&m[557]&~m[559]&m[560])|(~m[555]&m[556]&m[557]&~m[559]&m[560])|(m[555]&m[556]&m[557]&~m[559]&m[560])|(m[555]&m[556]&m[557]&m[559]&m[560]))):InitCond[650];
    m[563] = run?((((m[560]&~m[561]&~m[562]&~m[564]&~m[565])|(~m[560]&m[561]&~m[562]&~m[564]&~m[565])|(~m[560]&~m[561]&m[562]&~m[564]&~m[565])|(m[560]&m[561]&m[562]&m[564]&~m[565])|(~m[560]&~m[561]&~m[562]&~m[564]&m[565])|(m[560]&m[561]&~m[562]&m[564]&m[565])|(m[560]&~m[561]&m[562]&m[564]&m[565])|(~m[560]&m[561]&m[562]&m[564]&m[565]))&UnbiasedRNG[312])|((m[560]&m[561]&~m[562]&~m[564]&~m[565])|(m[560]&~m[561]&m[562]&~m[564]&~m[565])|(~m[560]&m[561]&m[562]&~m[564]&~m[565])|(m[560]&m[561]&m[562]&~m[564]&~m[565])|(m[560]&~m[561]&~m[562]&~m[564]&m[565])|(~m[560]&m[561]&~m[562]&~m[564]&m[565])|(m[560]&m[561]&~m[562]&~m[564]&m[565])|(~m[560]&~m[561]&m[562]&~m[564]&m[565])|(m[560]&~m[561]&m[562]&~m[564]&m[565])|(~m[560]&m[561]&m[562]&~m[564]&m[565])|(m[560]&m[561]&m[562]&~m[564]&m[565])|(m[560]&m[561]&m[562]&m[564]&m[565]))):InitCond[651];
    m[568] = run?((((m[565]&~m[566]&~m[567]&~m[569]&~m[570])|(~m[565]&m[566]&~m[567]&~m[569]&~m[570])|(~m[565]&~m[566]&m[567]&~m[569]&~m[570])|(m[565]&m[566]&m[567]&m[569]&~m[570])|(~m[565]&~m[566]&~m[567]&~m[569]&m[570])|(m[565]&m[566]&~m[567]&m[569]&m[570])|(m[565]&~m[566]&m[567]&m[569]&m[570])|(~m[565]&m[566]&m[567]&m[569]&m[570]))&UnbiasedRNG[313])|((m[565]&m[566]&~m[567]&~m[569]&~m[570])|(m[565]&~m[566]&m[567]&~m[569]&~m[570])|(~m[565]&m[566]&m[567]&~m[569]&~m[570])|(m[565]&m[566]&m[567]&~m[569]&~m[570])|(m[565]&~m[566]&~m[567]&~m[569]&m[570])|(~m[565]&m[566]&~m[567]&~m[569]&m[570])|(m[565]&m[566]&~m[567]&~m[569]&m[570])|(~m[565]&~m[566]&m[567]&~m[569]&m[570])|(m[565]&~m[566]&m[567]&~m[569]&m[570])|(~m[565]&m[566]&m[567]&~m[569]&m[570])|(m[565]&m[566]&m[567]&~m[569]&m[570])|(m[565]&m[566]&m[567]&m[569]&m[570]))):InitCond[652];
    m[573] = run?((((m[570]&~m[571]&~m[572]&~m[574]&~m[575])|(~m[570]&m[571]&~m[572]&~m[574]&~m[575])|(~m[570]&~m[571]&m[572]&~m[574]&~m[575])|(m[570]&m[571]&m[572]&m[574]&~m[575])|(~m[570]&~m[571]&~m[572]&~m[574]&m[575])|(m[570]&m[571]&~m[572]&m[574]&m[575])|(m[570]&~m[571]&m[572]&m[574]&m[575])|(~m[570]&m[571]&m[572]&m[574]&m[575]))&UnbiasedRNG[314])|((m[570]&m[571]&~m[572]&~m[574]&~m[575])|(m[570]&~m[571]&m[572]&~m[574]&~m[575])|(~m[570]&m[571]&m[572]&~m[574]&~m[575])|(m[570]&m[571]&m[572]&~m[574]&~m[575])|(m[570]&~m[571]&~m[572]&~m[574]&m[575])|(~m[570]&m[571]&~m[572]&~m[574]&m[575])|(m[570]&m[571]&~m[572]&~m[574]&m[575])|(~m[570]&~m[571]&m[572]&~m[574]&m[575])|(m[570]&~m[571]&m[572]&~m[574]&m[575])|(~m[570]&m[571]&m[572]&~m[574]&m[575])|(m[570]&m[571]&m[572]&~m[574]&m[575])|(m[570]&m[571]&m[572]&m[574]&m[575]))):InitCond[653];
    m[578] = run?((((m[575]&~m[576]&~m[577]&~m[579]&~m[580])|(~m[575]&m[576]&~m[577]&~m[579]&~m[580])|(~m[575]&~m[576]&m[577]&~m[579]&~m[580])|(m[575]&m[576]&m[577]&m[579]&~m[580])|(~m[575]&~m[576]&~m[577]&~m[579]&m[580])|(m[575]&m[576]&~m[577]&m[579]&m[580])|(m[575]&~m[576]&m[577]&m[579]&m[580])|(~m[575]&m[576]&m[577]&m[579]&m[580]))&UnbiasedRNG[315])|((m[575]&m[576]&~m[577]&~m[579]&~m[580])|(m[575]&~m[576]&m[577]&~m[579]&~m[580])|(~m[575]&m[576]&m[577]&~m[579]&~m[580])|(m[575]&m[576]&m[577]&~m[579]&~m[580])|(m[575]&~m[576]&~m[577]&~m[579]&m[580])|(~m[575]&m[576]&~m[577]&~m[579]&m[580])|(m[575]&m[576]&~m[577]&~m[579]&m[580])|(~m[575]&~m[576]&m[577]&~m[579]&m[580])|(m[575]&~m[576]&m[577]&~m[579]&m[580])|(~m[575]&m[576]&m[577]&~m[579]&m[580])|(m[575]&m[576]&m[577]&~m[579]&m[580])|(m[575]&m[576]&m[577]&m[579]&m[580]))):InitCond[654];
    m[588] = run?((((m[585]&~m[586]&~m[587]&~m[589]&~m[590])|(~m[585]&m[586]&~m[587]&~m[589]&~m[590])|(~m[585]&~m[586]&m[587]&~m[589]&~m[590])|(m[585]&m[586]&m[587]&m[589]&~m[590])|(~m[585]&~m[586]&~m[587]&~m[589]&m[590])|(m[585]&m[586]&~m[587]&m[589]&m[590])|(m[585]&~m[586]&m[587]&m[589]&m[590])|(~m[585]&m[586]&m[587]&m[589]&m[590]))&UnbiasedRNG[316])|((m[585]&m[586]&~m[587]&~m[589]&~m[590])|(m[585]&~m[586]&m[587]&~m[589]&~m[590])|(~m[585]&m[586]&m[587]&~m[589]&~m[590])|(m[585]&m[586]&m[587]&~m[589]&~m[590])|(m[585]&~m[586]&~m[587]&~m[589]&m[590])|(~m[585]&m[586]&~m[587]&~m[589]&m[590])|(m[585]&m[586]&~m[587]&~m[589]&m[590])|(~m[585]&~m[586]&m[587]&~m[589]&m[590])|(m[585]&~m[586]&m[587]&~m[589]&m[590])|(~m[585]&m[586]&m[587]&~m[589]&m[590])|(m[585]&m[586]&m[587]&~m[589]&m[590])|(m[585]&m[586]&m[587]&m[589]&m[590]))):InitCond[655];
    m[593] = run?((((m[590]&~m[591]&~m[592]&~m[594]&~m[595])|(~m[590]&m[591]&~m[592]&~m[594]&~m[595])|(~m[590]&~m[591]&m[592]&~m[594]&~m[595])|(m[590]&m[591]&m[592]&m[594]&~m[595])|(~m[590]&~m[591]&~m[592]&~m[594]&m[595])|(m[590]&m[591]&~m[592]&m[594]&m[595])|(m[590]&~m[591]&m[592]&m[594]&m[595])|(~m[590]&m[591]&m[592]&m[594]&m[595]))&UnbiasedRNG[317])|((m[590]&m[591]&~m[592]&~m[594]&~m[595])|(m[590]&~m[591]&m[592]&~m[594]&~m[595])|(~m[590]&m[591]&m[592]&~m[594]&~m[595])|(m[590]&m[591]&m[592]&~m[594]&~m[595])|(m[590]&~m[591]&~m[592]&~m[594]&m[595])|(~m[590]&m[591]&~m[592]&~m[594]&m[595])|(m[590]&m[591]&~m[592]&~m[594]&m[595])|(~m[590]&~m[591]&m[592]&~m[594]&m[595])|(m[590]&~m[591]&m[592]&~m[594]&m[595])|(~m[590]&m[591]&m[592]&~m[594]&m[595])|(m[590]&m[591]&m[592]&~m[594]&m[595])|(m[590]&m[591]&m[592]&m[594]&m[595]))):InitCond[656];
    m[598] = run?((((m[595]&~m[596]&~m[597]&~m[599]&~m[600])|(~m[595]&m[596]&~m[597]&~m[599]&~m[600])|(~m[595]&~m[596]&m[597]&~m[599]&~m[600])|(m[595]&m[596]&m[597]&m[599]&~m[600])|(~m[595]&~m[596]&~m[597]&~m[599]&m[600])|(m[595]&m[596]&~m[597]&m[599]&m[600])|(m[595]&~m[596]&m[597]&m[599]&m[600])|(~m[595]&m[596]&m[597]&m[599]&m[600]))&UnbiasedRNG[318])|((m[595]&m[596]&~m[597]&~m[599]&~m[600])|(m[595]&~m[596]&m[597]&~m[599]&~m[600])|(~m[595]&m[596]&m[597]&~m[599]&~m[600])|(m[595]&m[596]&m[597]&~m[599]&~m[600])|(m[595]&~m[596]&~m[597]&~m[599]&m[600])|(~m[595]&m[596]&~m[597]&~m[599]&m[600])|(m[595]&m[596]&~m[597]&~m[599]&m[600])|(~m[595]&~m[596]&m[597]&~m[599]&m[600])|(m[595]&~m[596]&m[597]&~m[599]&m[600])|(~m[595]&m[596]&m[597]&~m[599]&m[600])|(m[595]&m[596]&m[597]&~m[599]&m[600])|(m[595]&m[596]&m[597]&m[599]&m[600]))):InitCond[657];
    m[603] = run?((((m[600]&~m[601]&~m[602]&~m[604]&~m[605])|(~m[600]&m[601]&~m[602]&~m[604]&~m[605])|(~m[600]&~m[601]&m[602]&~m[604]&~m[605])|(m[600]&m[601]&m[602]&m[604]&~m[605])|(~m[600]&~m[601]&~m[602]&~m[604]&m[605])|(m[600]&m[601]&~m[602]&m[604]&m[605])|(m[600]&~m[601]&m[602]&m[604]&m[605])|(~m[600]&m[601]&m[602]&m[604]&m[605]))&UnbiasedRNG[319])|((m[600]&m[601]&~m[602]&~m[604]&~m[605])|(m[600]&~m[601]&m[602]&~m[604]&~m[605])|(~m[600]&m[601]&m[602]&~m[604]&~m[605])|(m[600]&m[601]&m[602]&~m[604]&~m[605])|(m[600]&~m[601]&~m[602]&~m[604]&m[605])|(~m[600]&m[601]&~m[602]&~m[604]&m[605])|(m[600]&m[601]&~m[602]&~m[604]&m[605])|(~m[600]&~m[601]&m[602]&~m[604]&m[605])|(m[600]&~m[601]&m[602]&~m[604]&m[605])|(~m[600]&m[601]&m[602]&~m[604]&m[605])|(m[600]&m[601]&m[602]&~m[604]&m[605])|(m[600]&m[601]&m[602]&m[604]&m[605]))):InitCond[658];
    m[608] = run?((((m[605]&~m[606]&~m[607]&~m[609]&~m[610])|(~m[605]&m[606]&~m[607]&~m[609]&~m[610])|(~m[605]&~m[606]&m[607]&~m[609]&~m[610])|(m[605]&m[606]&m[607]&m[609]&~m[610])|(~m[605]&~m[606]&~m[607]&~m[609]&m[610])|(m[605]&m[606]&~m[607]&m[609]&m[610])|(m[605]&~m[606]&m[607]&m[609]&m[610])|(~m[605]&m[606]&m[607]&m[609]&m[610]))&UnbiasedRNG[320])|((m[605]&m[606]&~m[607]&~m[609]&~m[610])|(m[605]&~m[606]&m[607]&~m[609]&~m[610])|(~m[605]&m[606]&m[607]&~m[609]&~m[610])|(m[605]&m[606]&m[607]&~m[609]&~m[610])|(m[605]&~m[606]&~m[607]&~m[609]&m[610])|(~m[605]&m[606]&~m[607]&~m[609]&m[610])|(m[605]&m[606]&~m[607]&~m[609]&m[610])|(~m[605]&~m[606]&m[607]&~m[609]&m[610])|(m[605]&~m[606]&m[607]&~m[609]&m[610])|(~m[605]&m[606]&m[607]&~m[609]&m[610])|(m[605]&m[606]&m[607]&~m[609]&m[610])|(m[605]&m[606]&m[607]&m[609]&m[610]))):InitCond[659];
    m[613] = run?((((m[610]&~m[611]&~m[612]&~m[614]&~m[615])|(~m[610]&m[611]&~m[612]&~m[614]&~m[615])|(~m[610]&~m[611]&m[612]&~m[614]&~m[615])|(m[610]&m[611]&m[612]&m[614]&~m[615])|(~m[610]&~m[611]&~m[612]&~m[614]&m[615])|(m[610]&m[611]&~m[612]&m[614]&m[615])|(m[610]&~m[611]&m[612]&m[614]&m[615])|(~m[610]&m[611]&m[612]&m[614]&m[615]))&UnbiasedRNG[321])|((m[610]&m[611]&~m[612]&~m[614]&~m[615])|(m[610]&~m[611]&m[612]&~m[614]&~m[615])|(~m[610]&m[611]&m[612]&~m[614]&~m[615])|(m[610]&m[611]&m[612]&~m[614]&~m[615])|(m[610]&~m[611]&~m[612]&~m[614]&m[615])|(~m[610]&m[611]&~m[612]&~m[614]&m[615])|(m[610]&m[611]&~m[612]&~m[614]&m[615])|(~m[610]&~m[611]&m[612]&~m[614]&m[615])|(m[610]&~m[611]&m[612]&~m[614]&m[615])|(~m[610]&m[611]&m[612]&~m[614]&m[615])|(m[610]&m[611]&m[612]&~m[614]&m[615])|(m[610]&m[611]&m[612]&m[614]&m[615]))):InitCond[660];
    m[618] = run?((((m[615]&~m[616]&~m[617]&~m[619]&~m[620])|(~m[615]&m[616]&~m[617]&~m[619]&~m[620])|(~m[615]&~m[616]&m[617]&~m[619]&~m[620])|(m[615]&m[616]&m[617]&m[619]&~m[620])|(~m[615]&~m[616]&~m[617]&~m[619]&m[620])|(m[615]&m[616]&~m[617]&m[619]&m[620])|(m[615]&~m[616]&m[617]&m[619]&m[620])|(~m[615]&m[616]&m[617]&m[619]&m[620]))&UnbiasedRNG[322])|((m[615]&m[616]&~m[617]&~m[619]&~m[620])|(m[615]&~m[616]&m[617]&~m[619]&~m[620])|(~m[615]&m[616]&m[617]&~m[619]&~m[620])|(m[615]&m[616]&m[617]&~m[619]&~m[620])|(m[615]&~m[616]&~m[617]&~m[619]&m[620])|(~m[615]&m[616]&~m[617]&~m[619]&m[620])|(m[615]&m[616]&~m[617]&~m[619]&m[620])|(~m[615]&~m[616]&m[617]&~m[619]&m[620])|(m[615]&~m[616]&m[617]&~m[619]&m[620])|(~m[615]&m[616]&m[617]&~m[619]&m[620])|(m[615]&m[616]&m[617]&~m[619]&m[620])|(m[615]&m[616]&m[617]&m[619]&m[620]))):InitCond[661];
    m[623] = run?((((m[620]&~m[621]&~m[622]&~m[624]&~m[625])|(~m[620]&m[621]&~m[622]&~m[624]&~m[625])|(~m[620]&~m[621]&m[622]&~m[624]&~m[625])|(m[620]&m[621]&m[622]&m[624]&~m[625])|(~m[620]&~m[621]&~m[622]&~m[624]&m[625])|(m[620]&m[621]&~m[622]&m[624]&m[625])|(m[620]&~m[621]&m[622]&m[624]&m[625])|(~m[620]&m[621]&m[622]&m[624]&m[625]))&UnbiasedRNG[323])|((m[620]&m[621]&~m[622]&~m[624]&~m[625])|(m[620]&~m[621]&m[622]&~m[624]&~m[625])|(~m[620]&m[621]&m[622]&~m[624]&~m[625])|(m[620]&m[621]&m[622]&~m[624]&~m[625])|(m[620]&~m[621]&~m[622]&~m[624]&m[625])|(~m[620]&m[621]&~m[622]&~m[624]&m[625])|(m[620]&m[621]&~m[622]&~m[624]&m[625])|(~m[620]&~m[621]&m[622]&~m[624]&m[625])|(m[620]&~m[621]&m[622]&~m[624]&m[625])|(~m[620]&m[621]&m[622]&~m[624]&m[625])|(m[620]&m[621]&m[622]&~m[624]&m[625])|(m[620]&m[621]&m[622]&m[624]&m[625]))):InitCond[662];
    m[633] = run?((((m[630]&~m[631]&~m[632]&~m[634]&~m[635])|(~m[630]&m[631]&~m[632]&~m[634]&~m[635])|(~m[630]&~m[631]&m[632]&~m[634]&~m[635])|(m[630]&m[631]&m[632]&m[634]&~m[635])|(~m[630]&~m[631]&~m[632]&~m[634]&m[635])|(m[630]&m[631]&~m[632]&m[634]&m[635])|(m[630]&~m[631]&m[632]&m[634]&m[635])|(~m[630]&m[631]&m[632]&m[634]&m[635]))&UnbiasedRNG[324])|((m[630]&m[631]&~m[632]&~m[634]&~m[635])|(m[630]&~m[631]&m[632]&~m[634]&~m[635])|(~m[630]&m[631]&m[632]&~m[634]&~m[635])|(m[630]&m[631]&m[632]&~m[634]&~m[635])|(m[630]&~m[631]&~m[632]&~m[634]&m[635])|(~m[630]&m[631]&~m[632]&~m[634]&m[635])|(m[630]&m[631]&~m[632]&~m[634]&m[635])|(~m[630]&~m[631]&m[632]&~m[634]&m[635])|(m[630]&~m[631]&m[632]&~m[634]&m[635])|(~m[630]&m[631]&m[632]&~m[634]&m[635])|(m[630]&m[631]&m[632]&~m[634]&m[635])|(m[630]&m[631]&m[632]&m[634]&m[635]))):InitCond[663];
    m[638] = run?((((m[635]&~m[636]&~m[637]&~m[639]&~m[640])|(~m[635]&m[636]&~m[637]&~m[639]&~m[640])|(~m[635]&~m[636]&m[637]&~m[639]&~m[640])|(m[635]&m[636]&m[637]&m[639]&~m[640])|(~m[635]&~m[636]&~m[637]&~m[639]&m[640])|(m[635]&m[636]&~m[637]&m[639]&m[640])|(m[635]&~m[636]&m[637]&m[639]&m[640])|(~m[635]&m[636]&m[637]&m[639]&m[640]))&UnbiasedRNG[325])|((m[635]&m[636]&~m[637]&~m[639]&~m[640])|(m[635]&~m[636]&m[637]&~m[639]&~m[640])|(~m[635]&m[636]&m[637]&~m[639]&~m[640])|(m[635]&m[636]&m[637]&~m[639]&~m[640])|(m[635]&~m[636]&~m[637]&~m[639]&m[640])|(~m[635]&m[636]&~m[637]&~m[639]&m[640])|(m[635]&m[636]&~m[637]&~m[639]&m[640])|(~m[635]&~m[636]&m[637]&~m[639]&m[640])|(m[635]&~m[636]&m[637]&~m[639]&m[640])|(~m[635]&m[636]&m[637]&~m[639]&m[640])|(m[635]&m[636]&m[637]&~m[639]&m[640])|(m[635]&m[636]&m[637]&m[639]&m[640]))):InitCond[664];
    m[643] = run?((((m[640]&~m[641]&~m[642]&~m[644]&~m[645])|(~m[640]&m[641]&~m[642]&~m[644]&~m[645])|(~m[640]&~m[641]&m[642]&~m[644]&~m[645])|(m[640]&m[641]&m[642]&m[644]&~m[645])|(~m[640]&~m[641]&~m[642]&~m[644]&m[645])|(m[640]&m[641]&~m[642]&m[644]&m[645])|(m[640]&~m[641]&m[642]&m[644]&m[645])|(~m[640]&m[641]&m[642]&m[644]&m[645]))&UnbiasedRNG[326])|((m[640]&m[641]&~m[642]&~m[644]&~m[645])|(m[640]&~m[641]&m[642]&~m[644]&~m[645])|(~m[640]&m[641]&m[642]&~m[644]&~m[645])|(m[640]&m[641]&m[642]&~m[644]&~m[645])|(m[640]&~m[641]&~m[642]&~m[644]&m[645])|(~m[640]&m[641]&~m[642]&~m[644]&m[645])|(m[640]&m[641]&~m[642]&~m[644]&m[645])|(~m[640]&~m[641]&m[642]&~m[644]&m[645])|(m[640]&~m[641]&m[642]&~m[644]&m[645])|(~m[640]&m[641]&m[642]&~m[644]&m[645])|(m[640]&m[641]&m[642]&~m[644]&m[645])|(m[640]&m[641]&m[642]&m[644]&m[645]))):InitCond[665];
    m[648] = run?((((m[645]&~m[646]&~m[647]&~m[649]&~m[650])|(~m[645]&m[646]&~m[647]&~m[649]&~m[650])|(~m[645]&~m[646]&m[647]&~m[649]&~m[650])|(m[645]&m[646]&m[647]&m[649]&~m[650])|(~m[645]&~m[646]&~m[647]&~m[649]&m[650])|(m[645]&m[646]&~m[647]&m[649]&m[650])|(m[645]&~m[646]&m[647]&m[649]&m[650])|(~m[645]&m[646]&m[647]&m[649]&m[650]))&UnbiasedRNG[327])|((m[645]&m[646]&~m[647]&~m[649]&~m[650])|(m[645]&~m[646]&m[647]&~m[649]&~m[650])|(~m[645]&m[646]&m[647]&~m[649]&~m[650])|(m[645]&m[646]&m[647]&~m[649]&~m[650])|(m[645]&~m[646]&~m[647]&~m[649]&m[650])|(~m[645]&m[646]&~m[647]&~m[649]&m[650])|(m[645]&m[646]&~m[647]&~m[649]&m[650])|(~m[645]&~m[646]&m[647]&~m[649]&m[650])|(m[645]&~m[646]&m[647]&~m[649]&m[650])|(~m[645]&m[646]&m[647]&~m[649]&m[650])|(m[645]&m[646]&m[647]&~m[649]&m[650])|(m[645]&m[646]&m[647]&m[649]&m[650]))):InitCond[666];
    m[653] = run?((((m[650]&~m[651]&~m[652]&~m[654]&~m[655])|(~m[650]&m[651]&~m[652]&~m[654]&~m[655])|(~m[650]&~m[651]&m[652]&~m[654]&~m[655])|(m[650]&m[651]&m[652]&m[654]&~m[655])|(~m[650]&~m[651]&~m[652]&~m[654]&m[655])|(m[650]&m[651]&~m[652]&m[654]&m[655])|(m[650]&~m[651]&m[652]&m[654]&m[655])|(~m[650]&m[651]&m[652]&m[654]&m[655]))&UnbiasedRNG[328])|((m[650]&m[651]&~m[652]&~m[654]&~m[655])|(m[650]&~m[651]&m[652]&~m[654]&~m[655])|(~m[650]&m[651]&m[652]&~m[654]&~m[655])|(m[650]&m[651]&m[652]&~m[654]&~m[655])|(m[650]&~m[651]&~m[652]&~m[654]&m[655])|(~m[650]&m[651]&~m[652]&~m[654]&m[655])|(m[650]&m[651]&~m[652]&~m[654]&m[655])|(~m[650]&~m[651]&m[652]&~m[654]&m[655])|(m[650]&~m[651]&m[652]&~m[654]&m[655])|(~m[650]&m[651]&m[652]&~m[654]&m[655])|(m[650]&m[651]&m[652]&~m[654]&m[655])|(m[650]&m[651]&m[652]&m[654]&m[655]))):InitCond[667];
    m[658] = run?((((m[655]&~m[656]&~m[657]&~m[659]&~m[660])|(~m[655]&m[656]&~m[657]&~m[659]&~m[660])|(~m[655]&~m[656]&m[657]&~m[659]&~m[660])|(m[655]&m[656]&m[657]&m[659]&~m[660])|(~m[655]&~m[656]&~m[657]&~m[659]&m[660])|(m[655]&m[656]&~m[657]&m[659]&m[660])|(m[655]&~m[656]&m[657]&m[659]&m[660])|(~m[655]&m[656]&m[657]&m[659]&m[660]))&UnbiasedRNG[329])|((m[655]&m[656]&~m[657]&~m[659]&~m[660])|(m[655]&~m[656]&m[657]&~m[659]&~m[660])|(~m[655]&m[656]&m[657]&~m[659]&~m[660])|(m[655]&m[656]&m[657]&~m[659]&~m[660])|(m[655]&~m[656]&~m[657]&~m[659]&m[660])|(~m[655]&m[656]&~m[657]&~m[659]&m[660])|(m[655]&m[656]&~m[657]&~m[659]&m[660])|(~m[655]&~m[656]&m[657]&~m[659]&m[660])|(m[655]&~m[656]&m[657]&~m[659]&m[660])|(~m[655]&m[656]&m[657]&~m[659]&m[660])|(m[655]&m[656]&m[657]&~m[659]&m[660])|(m[655]&m[656]&m[657]&m[659]&m[660]))):InitCond[668];
    m[663] = run?((((m[660]&~m[661]&~m[662]&~m[664]&~m[665])|(~m[660]&m[661]&~m[662]&~m[664]&~m[665])|(~m[660]&~m[661]&m[662]&~m[664]&~m[665])|(m[660]&m[661]&m[662]&m[664]&~m[665])|(~m[660]&~m[661]&~m[662]&~m[664]&m[665])|(m[660]&m[661]&~m[662]&m[664]&m[665])|(m[660]&~m[661]&m[662]&m[664]&m[665])|(~m[660]&m[661]&m[662]&m[664]&m[665]))&UnbiasedRNG[330])|((m[660]&m[661]&~m[662]&~m[664]&~m[665])|(m[660]&~m[661]&m[662]&~m[664]&~m[665])|(~m[660]&m[661]&m[662]&~m[664]&~m[665])|(m[660]&m[661]&m[662]&~m[664]&~m[665])|(m[660]&~m[661]&~m[662]&~m[664]&m[665])|(~m[660]&m[661]&~m[662]&~m[664]&m[665])|(m[660]&m[661]&~m[662]&~m[664]&m[665])|(~m[660]&~m[661]&m[662]&~m[664]&m[665])|(m[660]&~m[661]&m[662]&~m[664]&m[665])|(~m[660]&m[661]&m[662]&~m[664]&m[665])|(m[660]&m[661]&m[662]&~m[664]&m[665])|(m[660]&m[661]&m[662]&m[664]&m[665]))):InitCond[669];
    m[673] = run?((((m[670]&~m[671]&~m[672]&~m[674]&~m[675])|(~m[670]&m[671]&~m[672]&~m[674]&~m[675])|(~m[670]&~m[671]&m[672]&~m[674]&~m[675])|(m[670]&m[671]&m[672]&m[674]&~m[675])|(~m[670]&~m[671]&~m[672]&~m[674]&m[675])|(m[670]&m[671]&~m[672]&m[674]&m[675])|(m[670]&~m[671]&m[672]&m[674]&m[675])|(~m[670]&m[671]&m[672]&m[674]&m[675]))&UnbiasedRNG[331])|((m[670]&m[671]&~m[672]&~m[674]&~m[675])|(m[670]&~m[671]&m[672]&~m[674]&~m[675])|(~m[670]&m[671]&m[672]&~m[674]&~m[675])|(m[670]&m[671]&m[672]&~m[674]&~m[675])|(m[670]&~m[671]&~m[672]&~m[674]&m[675])|(~m[670]&m[671]&~m[672]&~m[674]&m[675])|(m[670]&m[671]&~m[672]&~m[674]&m[675])|(~m[670]&~m[671]&m[672]&~m[674]&m[675])|(m[670]&~m[671]&m[672]&~m[674]&m[675])|(~m[670]&m[671]&m[672]&~m[674]&m[675])|(m[670]&m[671]&m[672]&~m[674]&m[675])|(m[670]&m[671]&m[672]&m[674]&m[675]))):InitCond[670];
    m[678] = run?((((m[675]&~m[676]&~m[677]&~m[679]&~m[680])|(~m[675]&m[676]&~m[677]&~m[679]&~m[680])|(~m[675]&~m[676]&m[677]&~m[679]&~m[680])|(m[675]&m[676]&m[677]&m[679]&~m[680])|(~m[675]&~m[676]&~m[677]&~m[679]&m[680])|(m[675]&m[676]&~m[677]&m[679]&m[680])|(m[675]&~m[676]&m[677]&m[679]&m[680])|(~m[675]&m[676]&m[677]&m[679]&m[680]))&UnbiasedRNG[332])|((m[675]&m[676]&~m[677]&~m[679]&~m[680])|(m[675]&~m[676]&m[677]&~m[679]&~m[680])|(~m[675]&m[676]&m[677]&~m[679]&~m[680])|(m[675]&m[676]&m[677]&~m[679]&~m[680])|(m[675]&~m[676]&~m[677]&~m[679]&m[680])|(~m[675]&m[676]&~m[677]&~m[679]&m[680])|(m[675]&m[676]&~m[677]&~m[679]&m[680])|(~m[675]&~m[676]&m[677]&~m[679]&m[680])|(m[675]&~m[676]&m[677]&~m[679]&m[680])|(~m[675]&m[676]&m[677]&~m[679]&m[680])|(m[675]&m[676]&m[677]&~m[679]&m[680])|(m[675]&m[676]&m[677]&m[679]&m[680]))):InitCond[671];
    m[683] = run?((((m[680]&~m[681]&~m[682]&~m[684]&~m[685])|(~m[680]&m[681]&~m[682]&~m[684]&~m[685])|(~m[680]&~m[681]&m[682]&~m[684]&~m[685])|(m[680]&m[681]&m[682]&m[684]&~m[685])|(~m[680]&~m[681]&~m[682]&~m[684]&m[685])|(m[680]&m[681]&~m[682]&m[684]&m[685])|(m[680]&~m[681]&m[682]&m[684]&m[685])|(~m[680]&m[681]&m[682]&m[684]&m[685]))&UnbiasedRNG[333])|((m[680]&m[681]&~m[682]&~m[684]&~m[685])|(m[680]&~m[681]&m[682]&~m[684]&~m[685])|(~m[680]&m[681]&m[682]&~m[684]&~m[685])|(m[680]&m[681]&m[682]&~m[684]&~m[685])|(m[680]&~m[681]&~m[682]&~m[684]&m[685])|(~m[680]&m[681]&~m[682]&~m[684]&m[685])|(m[680]&m[681]&~m[682]&~m[684]&m[685])|(~m[680]&~m[681]&m[682]&~m[684]&m[685])|(m[680]&~m[681]&m[682]&~m[684]&m[685])|(~m[680]&m[681]&m[682]&~m[684]&m[685])|(m[680]&m[681]&m[682]&~m[684]&m[685])|(m[680]&m[681]&m[682]&m[684]&m[685]))):InitCond[672];
    m[688] = run?((((m[685]&~m[686]&~m[687]&~m[689]&~m[690])|(~m[685]&m[686]&~m[687]&~m[689]&~m[690])|(~m[685]&~m[686]&m[687]&~m[689]&~m[690])|(m[685]&m[686]&m[687]&m[689]&~m[690])|(~m[685]&~m[686]&~m[687]&~m[689]&m[690])|(m[685]&m[686]&~m[687]&m[689]&m[690])|(m[685]&~m[686]&m[687]&m[689]&m[690])|(~m[685]&m[686]&m[687]&m[689]&m[690]))&UnbiasedRNG[334])|((m[685]&m[686]&~m[687]&~m[689]&~m[690])|(m[685]&~m[686]&m[687]&~m[689]&~m[690])|(~m[685]&m[686]&m[687]&~m[689]&~m[690])|(m[685]&m[686]&m[687]&~m[689]&~m[690])|(m[685]&~m[686]&~m[687]&~m[689]&m[690])|(~m[685]&m[686]&~m[687]&~m[689]&m[690])|(m[685]&m[686]&~m[687]&~m[689]&m[690])|(~m[685]&~m[686]&m[687]&~m[689]&m[690])|(m[685]&~m[686]&m[687]&~m[689]&m[690])|(~m[685]&m[686]&m[687]&~m[689]&m[690])|(m[685]&m[686]&m[687]&~m[689]&m[690])|(m[685]&m[686]&m[687]&m[689]&m[690]))):InitCond[673];
    m[693] = run?((((m[690]&~m[691]&~m[692]&~m[694]&~m[695])|(~m[690]&m[691]&~m[692]&~m[694]&~m[695])|(~m[690]&~m[691]&m[692]&~m[694]&~m[695])|(m[690]&m[691]&m[692]&m[694]&~m[695])|(~m[690]&~m[691]&~m[692]&~m[694]&m[695])|(m[690]&m[691]&~m[692]&m[694]&m[695])|(m[690]&~m[691]&m[692]&m[694]&m[695])|(~m[690]&m[691]&m[692]&m[694]&m[695]))&UnbiasedRNG[335])|((m[690]&m[691]&~m[692]&~m[694]&~m[695])|(m[690]&~m[691]&m[692]&~m[694]&~m[695])|(~m[690]&m[691]&m[692]&~m[694]&~m[695])|(m[690]&m[691]&m[692]&~m[694]&~m[695])|(m[690]&~m[691]&~m[692]&~m[694]&m[695])|(~m[690]&m[691]&~m[692]&~m[694]&m[695])|(m[690]&m[691]&~m[692]&~m[694]&m[695])|(~m[690]&~m[691]&m[692]&~m[694]&m[695])|(m[690]&~m[691]&m[692]&~m[694]&m[695])|(~m[690]&m[691]&m[692]&~m[694]&m[695])|(m[690]&m[691]&m[692]&~m[694]&m[695])|(m[690]&m[691]&m[692]&m[694]&m[695]))):InitCond[674];
    m[698] = run?((((m[695]&~m[696]&~m[697]&~m[699]&~m[700])|(~m[695]&m[696]&~m[697]&~m[699]&~m[700])|(~m[695]&~m[696]&m[697]&~m[699]&~m[700])|(m[695]&m[696]&m[697]&m[699]&~m[700])|(~m[695]&~m[696]&~m[697]&~m[699]&m[700])|(m[695]&m[696]&~m[697]&m[699]&m[700])|(m[695]&~m[696]&m[697]&m[699]&m[700])|(~m[695]&m[696]&m[697]&m[699]&m[700]))&UnbiasedRNG[336])|((m[695]&m[696]&~m[697]&~m[699]&~m[700])|(m[695]&~m[696]&m[697]&~m[699]&~m[700])|(~m[695]&m[696]&m[697]&~m[699]&~m[700])|(m[695]&m[696]&m[697]&~m[699]&~m[700])|(m[695]&~m[696]&~m[697]&~m[699]&m[700])|(~m[695]&m[696]&~m[697]&~m[699]&m[700])|(m[695]&m[696]&~m[697]&~m[699]&m[700])|(~m[695]&~m[696]&m[697]&~m[699]&m[700])|(m[695]&~m[696]&m[697]&~m[699]&m[700])|(~m[695]&m[696]&m[697]&~m[699]&m[700])|(m[695]&m[696]&m[697]&~m[699]&m[700])|(m[695]&m[696]&m[697]&m[699]&m[700]))):InitCond[675];
    m[708] = run?((((m[705]&~m[706]&~m[707]&~m[709]&~m[710])|(~m[705]&m[706]&~m[707]&~m[709]&~m[710])|(~m[705]&~m[706]&m[707]&~m[709]&~m[710])|(m[705]&m[706]&m[707]&m[709]&~m[710])|(~m[705]&~m[706]&~m[707]&~m[709]&m[710])|(m[705]&m[706]&~m[707]&m[709]&m[710])|(m[705]&~m[706]&m[707]&m[709]&m[710])|(~m[705]&m[706]&m[707]&m[709]&m[710]))&UnbiasedRNG[337])|((m[705]&m[706]&~m[707]&~m[709]&~m[710])|(m[705]&~m[706]&m[707]&~m[709]&~m[710])|(~m[705]&m[706]&m[707]&~m[709]&~m[710])|(m[705]&m[706]&m[707]&~m[709]&~m[710])|(m[705]&~m[706]&~m[707]&~m[709]&m[710])|(~m[705]&m[706]&~m[707]&~m[709]&m[710])|(m[705]&m[706]&~m[707]&~m[709]&m[710])|(~m[705]&~m[706]&m[707]&~m[709]&m[710])|(m[705]&~m[706]&m[707]&~m[709]&m[710])|(~m[705]&m[706]&m[707]&~m[709]&m[710])|(m[705]&m[706]&m[707]&~m[709]&m[710])|(m[705]&m[706]&m[707]&m[709]&m[710]))):InitCond[676];
    m[713] = run?((((m[710]&~m[711]&~m[712]&~m[714]&~m[715])|(~m[710]&m[711]&~m[712]&~m[714]&~m[715])|(~m[710]&~m[711]&m[712]&~m[714]&~m[715])|(m[710]&m[711]&m[712]&m[714]&~m[715])|(~m[710]&~m[711]&~m[712]&~m[714]&m[715])|(m[710]&m[711]&~m[712]&m[714]&m[715])|(m[710]&~m[711]&m[712]&m[714]&m[715])|(~m[710]&m[711]&m[712]&m[714]&m[715]))&UnbiasedRNG[338])|((m[710]&m[711]&~m[712]&~m[714]&~m[715])|(m[710]&~m[711]&m[712]&~m[714]&~m[715])|(~m[710]&m[711]&m[712]&~m[714]&~m[715])|(m[710]&m[711]&m[712]&~m[714]&~m[715])|(m[710]&~m[711]&~m[712]&~m[714]&m[715])|(~m[710]&m[711]&~m[712]&~m[714]&m[715])|(m[710]&m[711]&~m[712]&~m[714]&m[715])|(~m[710]&~m[711]&m[712]&~m[714]&m[715])|(m[710]&~m[711]&m[712]&~m[714]&m[715])|(~m[710]&m[711]&m[712]&~m[714]&m[715])|(m[710]&m[711]&m[712]&~m[714]&m[715])|(m[710]&m[711]&m[712]&m[714]&m[715]))):InitCond[677];
    m[718] = run?((((m[715]&~m[716]&~m[717]&~m[719]&~m[720])|(~m[715]&m[716]&~m[717]&~m[719]&~m[720])|(~m[715]&~m[716]&m[717]&~m[719]&~m[720])|(m[715]&m[716]&m[717]&m[719]&~m[720])|(~m[715]&~m[716]&~m[717]&~m[719]&m[720])|(m[715]&m[716]&~m[717]&m[719]&m[720])|(m[715]&~m[716]&m[717]&m[719]&m[720])|(~m[715]&m[716]&m[717]&m[719]&m[720]))&UnbiasedRNG[339])|((m[715]&m[716]&~m[717]&~m[719]&~m[720])|(m[715]&~m[716]&m[717]&~m[719]&~m[720])|(~m[715]&m[716]&m[717]&~m[719]&~m[720])|(m[715]&m[716]&m[717]&~m[719]&~m[720])|(m[715]&~m[716]&~m[717]&~m[719]&m[720])|(~m[715]&m[716]&~m[717]&~m[719]&m[720])|(m[715]&m[716]&~m[717]&~m[719]&m[720])|(~m[715]&~m[716]&m[717]&~m[719]&m[720])|(m[715]&~m[716]&m[717]&~m[719]&m[720])|(~m[715]&m[716]&m[717]&~m[719]&m[720])|(m[715]&m[716]&m[717]&~m[719]&m[720])|(m[715]&m[716]&m[717]&m[719]&m[720]))):InitCond[678];
    m[723] = run?((((m[720]&~m[721]&~m[722]&~m[724]&~m[725])|(~m[720]&m[721]&~m[722]&~m[724]&~m[725])|(~m[720]&~m[721]&m[722]&~m[724]&~m[725])|(m[720]&m[721]&m[722]&m[724]&~m[725])|(~m[720]&~m[721]&~m[722]&~m[724]&m[725])|(m[720]&m[721]&~m[722]&m[724]&m[725])|(m[720]&~m[721]&m[722]&m[724]&m[725])|(~m[720]&m[721]&m[722]&m[724]&m[725]))&UnbiasedRNG[340])|((m[720]&m[721]&~m[722]&~m[724]&~m[725])|(m[720]&~m[721]&m[722]&~m[724]&~m[725])|(~m[720]&m[721]&m[722]&~m[724]&~m[725])|(m[720]&m[721]&m[722]&~m[724]&~m[725])|(m[720]&~m[721]&~m[722]&~m[724]&m[725])|(~m[720]&m[721]&~m[722]&~m[724]&m[725])|(m[720]&m[721]&~m[722]&~m[724]&m[725])|(~m[720]&~m[721]&m[722]&~m[724]&m[725])|(m[720]&~m[721]&m[722]&~m[724]&m[725])|(~m[720]&m[721]&m[722]&~m[724]&m[725])|(m[720]&m[721]&m[722]&~m[724]&m[725])|(m[720]&m[721]&m[722]&m[724]&m[725]))):InitCond[679];
    m[728] = run?((((m[725]&~m[726]&~m[727]&~m[729]&~m[730])|(~m[725]&m[726]&~m[727]&~m[729]&~m[730])|(~m[725]&~m[726]&m[727]&~m[729]&~m[730])|(m[725]&m[726]&m[727]&m[729]&~m[730])|(~m[725]&~m[726]&~m[727]&~m[729]&m[730])|(m[725]&m[726]&~m[727]&m[729]&m[730])|(m[725]&~m[726]&m[727]&m[729]&m[730])|(~m[725]&m[726]&m[727]&m[729]&m[730]))&UnbiasedRNG[341])|((m[725]&m[726]&~m[727]&~m[729]&~m[730])|(m[725]&~m[726]&m[727]&~m[729]&~m[730])|(~m[725]&m[726]&m[727]&~m[729]&~m[730])|(m[725]&m[726]&m[727]&~m[729]&~m[730])|(m[725]&~m[726]&~m[727]&~m[729]&m[730])|(~m[725]&m[726]&~m[727]&~m[729]&m[730])|(m[725]&m[726]&~m[727]&~m[729]&m[730])|(~m[725]&~m[726]&m[727]&~m[729]&m[730])|(m[725]&~m[726]&m[727]&~m[729]&m[730])|(~m[725]&m[726]&m[727]&~m[729]&m[730])|(m[725]&m[726]&m[727]&~m[729]&m[730])|(m[725]&m[726]&m[727]&m[729]&m[730]))):InitCond[680];
    m[738] = run?((((m[735]&~m[736]&~m[737]&~m[739]&~m[740])|(~m[735]&m[736]&~m[737]&~m[739]&~m[740])|(~m[735]&~m[736]&m[737]&~m[739]&~m[740])|(m[735]&m[736]&m[737]&m[739]&~m[740])|(~m[735]&~m[736]&~m[737]&~m[739]&m[740])|(m[735]&m[736]&~m[737]&m[739]&m[740])|(m[735]&~m[736]&m[737]&m[739]&m[740])|(~m[735]&m[736]&m[737]&m[739]&m[740]))&UnbiasedRNG[342])|((m[735]&m[736]&~m[737]&~m[739]&~m[740])|(m[735]&~m[736]&m[737]&~m[739]&~m[740])|(~m[735]&m[736]&m[737]&~m[739]&~m[740])|(m[735]&m[736]&m[737]&~m[739]&~m[740])|(m[735]&~m[736]&~m[737]&~m[739]&m[740])|(~m[735]&m[736]&~m[737]&~m[739]&m[740])|(m[735]&m[736]&~m[737]&~m[739]&m[740])|(~m[735]&~m[736]&m[737]&~m[739]&m[740])|(m[735]&~m[736]&m[737]&~m[739]&m[740])|(~m[735]&m[736]&m[737]&~m[739]&m[740])|(m[735]&m[736]&m[737]&~m[739]&m[740])|(m[735]&m[736]&m[737]&m[739]&m[740]))):InitCond[681];
    m[743] = run?((((m[740]&~m[741]&~m[742]&~m[744]&~m[745])|(~m[740]&m[741]&~m[742]&~m[744]&~m[745])|(~m[740]&~m[741]&m[742]&~m[744]&~m[745])|(m[740]&m[741]&m[742]&m[744]&~m[745])|(~m[740]&~m[741]&~m[742]&~m[744]&m[745])|(m[740]&m[741]&~m[742]&m[744]&m[745])|(m[740]&~m[741]&m[742]&m[744]&m[745])|(~m[740]&m[741]&m[742]&m[744]&m[745]))&UnbiasedRNG[343])|((m[740]&m[741]&~m[742]&~m[744]&~m[745])|(m[740]&~m[741]&m[742]&~m[744]&~m[745])|(~m[740]&m[741]&m[742]&~m[744]&~m[745])|(m[740]&m[741]&m[742]&~m[744]&~m[745])|(m[740]&~m[741]&~m[742]&~m[744]&m[745])|(~m[740]&m[741]&~m[742]&~m[744]&m[745])|(m[740]&m[741]&~m[742]&~m[744]&m[745])|(~m[740]&~m[741]&m[742]&~m[744]&m[745])|(m[740]&~m[741]&m[742]&~m[744]&m[745])|(~m[740]&m[741]&m[742]&~m[744]&m[745])|(m[740]&m[741]&m[742]&~m[744]&m[745])|(m[740]&m[741]&m[742]&m[744]&m[745]))):InitCond[682];
    m[748] = run?((((m[745]&~m[746]&~m[747]&~m[749]&~m[750])|(~m[745]&m[746]&~m[747]&~m[749]&~m[750])|(~m[745]&~m[746]&m[747]&~m[749]&~m[750])|(m[745]&m[746]&m[747]&m[749]&~m[750])|(~m[745]&~m[746]&~m[747]&~m[749]&m[750])|(m[745]&m[746]&~m[747]&m[749]&m[750])|(m[745]&~m[746]&m[747]&m[749]&m[750])|(~m[745]&m[746]&m[747]&m[749]&m[750]))&UnbiasedRNG[344])|((m[745]&m[746]&~m[747]&~m[749]&~m[750])|(m[745]&~m[746]&m[747]&~m[749]&~m[750])|(~m[745]&m[746]&m[747]&~m[749]&~m[750])|(m[745]&m[746]&m[747]&~m[749]&~m[750])|(m[745]&~m[746]&~m[747]&~m[749]&m[750])|(~m[745]&m[746]&~m[747]&~m[749]&m[750])|(m[745]&m[746]&~m[747]&~m[749]&m[750])|(~m[745]&~m[746]&m[747]&~m[749]&m[750])|(m[745]&~m[746]&m[747]&~m[749]&m[750])|(~m[745]&m[746]&m[747]&~m[749]&m[750])|(m[745]&m[746]&m[747]&~m[749]&m[750])|(m[745]&m[746]&m[747]&m[749]&m[750]))):InitCond[683];
    m[753] = run?((((m[750]&~m[751]&~m[752]&~m[754]&~m[755])|(~m[750]&m[751]&~m[752]&~m[754]&~m[755])|(~m[750]&~m[751]&m[752]&~m[754]&~m[755])|(m[750]&m[751]&m[752]&m[754]&~m[755])|(~m[750]&~m[751]&~m[752]&~m[754]&m[755])|(m[750]&m[751]&~m[752]&m[754]&m[755])|(m[750]&~m[751]&m[752]&m[754]&m[755])|(~m[750]&m[751]&m[752]&m[754]&m[755]))&UnbiasedRNG[345])|((m[750]&m[751]&~m[752]&~m[754]&~m[755])|(m[750]&~m[751]&m[752]&~m[754]&~m[755])|(~m[750]&m[751]&m[752]&~m[754]&~m[755])|(m[750]&m[751]&m[752]&~m[754]&~m[755])|(m[750]&~m[751]&~m[752]&~m[754]&m[755])|(~m[750]&m[751]&~m[752]&~m[754]&m[755])|(m[750]&m[751]&~m[752]&~m[754]&m[755])|(~m[750]&~m[751]&m[752]&~m[754]&m[755])|(m[750]&~m[751]&m[752]&~m[754]&m[755])|(~m[750]&m[751]&m[752]&~m[754]&m[755])|(m[750]&m[751]&m[752]&~m[754]&m[755])|(m[750]&m[751]&m[752]&m[754]&m[755]))):InitCond[684];
    m[763] = run?((((m[760]&~m[761]&~m[762]&~m[764]&~m[765])|(~m[760]&m[761]&~m[762]&~m[764]&~m[765])|(~m[760]&~m[761]&m[762]&~m[764]&~m[765])|(m[760]&m[761]&m[762]&m[764]&~m[765])|(~m[760]&~m[761]&~m[762]&~m[764]&m[765])|(m[760]&m[761]&~m[762]&m[764]&m[765])|(m[760]&~m[761]&m[762]&m[764]&m[765])|(~m[760]&m[761]&m[762]&m[764]&m[765]))&UnbiasedRNG[346])|((m[760]&m[761]&~m[762]&~m[764]&~m[765])|(m[760]&~m[761]&m[762]&~m[764]&~m[765])|(~m[760]&m[761]&m[762]&~m[764]&~m[765])|(m[760]&m[761]&m[762]&~m[764]&~m[765])|(m[760]&~m[761]&~m[762]&~m[764]&m[765])|(~m[760]&m[761]&~m[762]&~m[764]&m[765])|(m[760]&m[761]&~m[762]&~m[764]&m[765])|(~m[760]&~m[761]&m[762]&~m[764]&m[765])|(m[760]&~m[761]&m[762]&~m[764]&m[765])|(~m[760]&m[761]&m[762]&~m[764]&m[765])|(m[760]&m[761]&m[762]&~m[764]&m[765])|(m[760]&m[761]&m[762]&m[764]&m[765]))):InitCond[685];
    m[768] = run?((((m[765]&~m[766]&~m[767]&~m[769]&~m[770])|(~m[765]&m[766]&~m[767]&~m[769]&~m[770])|(~m[765]&~m[766]&m[767]&~m[769]&~m[770])|(m[765]&m[766]&m[767]&m[769]&~m[770])|(~m[765]&~m[766]&~m[767]&~m[769]&m[770])|(m[765]&m[766]&~m[767]&m[769]&m[770])|(m[765]&~m[766]&m[767]&m[769]&m[770])|(~m[765]&m[766]&m[767]&m[769]&m[770]))&UnbiasedRNG[347])|((m[765]&m[766]&~m[767]&~m[769]&~m[770])|(m[765]&~m[766]&m[767]&~m[769]&~m[770])|(~m[765]&m[766]&m[767]&~m[769]&~m[770])|(m[765]&m[766]&m[767]&~m[769]&~m[770])|(m[765]&~m[766]&~m[767]&~m[769]&m[770])|(~m[765]&m[766]&~m[767]&~m[769]&m[770])|(m[765]&m[766]&~m[767]&~m[769]&m[770])|(~m[765]&~m[766]&m[767]&~m[769]&m[770])|(m[765]&~m[766]&m[767]&~m[769]&m[770])|(~m[765]&m[766]&m[767]&~m[769]&m[770])|(m[765]&m[766]&m[767]&~m[769]&m[770])|(m[765]&m[766]&m[767]&m[769]&m[770]))):InitCond[686];
    m[773] = run?((((m[770]&~m[771]&~m[772]&~m[774]&~m[775])|(~m[770]&m[771]&~m[772]&~m[774]&~m[775])|(~m[770]&~m[771]&m[772]&~m[774]&~m[775])|(m[770]&m[771]&m[772]&m[774]&~m[775])|(~m[770]&~m[771]&~m[772]&~m[774]&m[775])|(m[770]&m[771]&~m[772]&m[774]&m[775])|(m[770]&~m[771]&m[772]&m[774]&m[775])|(~m[770]&m[771]&m[772]&m[774]&m[775]))&UnbiasedRNG[348])|((m[770]&m[771]&~m[772]&~m[774]&~m[775])|(m[770]&~m[771]&m[772]&~m[774]&~m[775])|(~m[770]&m[771]&m[772]&~m[774]&~m[775])|(m[770]&m[771]&m[772]&~m[774]&~m[775])|(m[770]&~m[771]&~m[772]&~m[774]&m[775])|(~m[770]&m[771]&~m[772]&~m[774]&m[775])|(m[770]&m[771]&~m[772]&~m[774]&m[775])|(~m[770]&~m[771]&m[772]&~m[774]&m[775])|(m[770]&~m[771]&m[772]&~m[774]&m[775])|(~m[770]&m[771]&m[772]&~m[774]&m[775])|(m[770]&m[771]&m[772]&~m[774]&m[775])|(m[770]&m[771]&m[772]&m[774]&m[775]))):InitCond[687];
    m[783] = run?((((m[780]&~m[781]&~m[782]&~m[784]&~m[785])|(~m[780]&m[781]&~m[782]&~m[784]&~m[785])|(~m[780]&~m[781]&m[782]&~m[784]&~m[785])|(m[780]&m[781]&m[782]&m[784]&~m[785])|(~m[780]&~m[781]&~m[782]&~m[784]&m[785])|(m[780]&m[781]&~m[782]&m[784]&m[785])|(m[780]&~m[781]&m[782]&m[784]&m[785])|(~m[780]&m[781]&m[782]&m[784]&m[785]))&UnbiasedRNG[349])|((m[780]&m[781]&~m[782]&~m[784]&~m[785])|(m[780]&~m[781]&m[782]&~m[784]&~m[785])|(~m[780]&m[781]&m[782]&~m[784]&~m[785])|(m[780]&m[781]&m[782]&~m[784]&~m[785])|(m[780]&~m[781]&~m[782]&~m[784]&m[785])|(~m[780]&m[781]&~m[782]&~m[784]&m[785])|(m[780]&m[781]&~m[782]&~m[784]&m[785])|(~m[780]&~m[781]&m[782]&~m[784]&m[785])|(m[780]&~m[781]&m[782]&~m[784]&m[785])|(~m[780]&m[781]&m[782]&~m[784]&m[785])|(m[780]&m[781]&m[782]&~m[784]&m[785])|(m[780]&m[781]&m[782]&m[784]&m[785]))):InitCond[688];
    m[788] = run?((((m[785]&~m[786]&~m[787]&~m[789]&~m[790])|(~m[785]&m[786]&~m[787]&~m[789]&~m[790])|(~m[785]&~m[786]&m[787]&~m[789]&~m[790])|(m[785]&m[786]&m[787]&m[789]&~m[790])|(~m[785]&~m[786]&~m[787]&~m[789]&m[790])|(m[785]&m[786]&~m[787]&m[789]&m[790])|(m[785]&~m[786]&m[787]&m[789]&m[790])|(~m[785]&m[786]&m[787]&m[789]&m[790]))&UnbiasedRNG[350])|((m[785]&m[786]&~m[787]&~m[789]&~m[790])|(m[785]&~m[786]&m[787]&~m[789]&~m[790])|(~m[785]&m[786]&m[787]&~m[789]&~m[790])|(m[785]&m[786]&m[787]&~m[789]&~m[790])|(m[785]&~m[786]&~m[787]&~m[789]&m[790])|(~m[785]&m[786]&~m[787]&~m[789]&m[790])|(m[785]&m[786]&~m[787]&~m[789]&m[790])|(~m[785]&~m[786]&m[787]&~m[789]&m[790])|(m[785]&~m[786]&m[787]&~m[789]&m[790])|(~m[785]&m[786]&m[787]&~m[789]&m[790])|(m[785]&m[786]&m[787]&~m[789]&m[790])|(m[785]&m[786]&m[787]&m[789]&m[790]))):InitCond[689];
    m[798] = run?((((m[795]&~m[796]&~m[797]&~m[799]&~m[800])|(~m[795]&m[796]&~m[797]&~m[799]&~m[800])|(~m[795]&~m[796]&m[797]&~m[799]&~m[800])|(m[795]&m[796]&m[797]&m[799]&~m[800])|(~m[795]&~m[796]&~m[797]&~m[799]&m[800])|(m[795]&m[796]&~m[797]&m[799]&m[800])|(m[795]&~m[796]&m[797]&m[799]&m[800])|(~m[795]&m[796]&m[797]&m[799]&m[800]))&UnbiasedRNG[351])|((m[795]&m[796]&~m[797]&~m[799]&~m[800])|(m[795]&~m[796]&m[797]&~m[799]&~m[800])|(~m[795]&m[796]&m[797]&~m[799]&~m[800])|(m[795]&m[796]&m[797]&~m[799]&~m[800])|(m[795]&~m[796]&~m[797]&~m[799]&m[800])|(~m[795]&m[796]&~m[797]&~m[799]&m[800])|(m[795]&m[796]&~m[797]&~m[799]&m[800])|(~m[795]&~m[796]&m[797]&~m[799]&m[800])|(m[795]&~m[796]&m[797]&~m[799]&m[800])|(~m[795]&m[796]&m[797]&~m[799]&m[800])|(m[795]&m[796]&m[797]&~m[799]&m[800])|(m[795]&m[796]&m[797]&m[799]&m[800]))):InitCond[690];
end

always @(posedge color4_clk) begin
    m[364] = run?((((m[360]&~m[361]&~m[362]&~m[363]&~m[367])|(~m[360]&m[361]&~m[362]&~m[363]&~m[367])|(~m[360]&~m[361]&m[362]&~m[363]&~m[367])|(m[360]&m[361]&~m[362]&m[363]&~m[367])|(m[360]&~m[361]&m[362]&m[363]&~m[367])|(~m[360]&m[361]&m[362]&m[363]&~m[367]))&BiasedRNG[339])|(((m[360]&~m[361]&~m[362]&~m[363]&m[367])|(~m[360]&m[361]&~m[362]&~m[363]&m[367])|(~m[360]&~m[361]&m[362]&~m[363]&m[367])|(m[360]&m[361]&~m[362]&m[363]&m[367])|(m[360]&~m[361]&m[362]&m[363]&m[367])|(~m[360]&m[361]&m[362]&m[363]&m[367]))&~BiasedRNG[339])|((m[360]&m[361]&~m[362]&~m[363]&~m[367])|(m[360]&~m[361]&m[362]&~m[363]&~m[367])|(~m[360]&m[361]&m[362]&~m[363]&~m[367])|(m[360]&m[361]&m[362]&~m[363]&~m[367])|(m[360]&m[361]&m[362]&m[363]&~m[367])|(m[360]&m[361]&~m[362]&~m[363]&m[367])|(m[360]&~m[361]&m[362]&~m[363]&m[367])|(~m[360]&m[361]&m[362]&~m[363]&m[367])|(m[360]&m[361]&m[362]&~m[363]&m[367])|(m[360]&m[361]&m[362]&m[363]&m[367]))):InitCond[691];
    m[369] = run?((((m[365]&~m[366]&~m[367]&~m[368]&~m[377])|(~m[365]&m[366]&~m[367]&~m[368]&~m[377])|(~m[365]&~m[366]&m[367]&~m[368]&~m[377])|(m[365]&m[366]&~m[367]&m[368]&~m[377])|(m[365]&~m[366]&m[367]&m[368]&~m[377])|(~m[365]&m[366]&m[367]&m[368]&~m[377]))&BiasedRNG[340])|(((m[365]&~m[366]&~m[367]&~m[368]&m[377])|(~m[365]&m[366]&~m[367]&~m[368]&m[377])|(~m[365]&~m[366]&m[367]&~m[368]&m[377])|(m[365]&m[366]&~m[367]&m[368]&m[377])|(m[365]&~m[366]&m[367]&m[368]&m[377])|(~m[365]&m[366]&m[367]&m[368]&m[377]))&~BiasedRNG[340])|((m[365]&m[366]&~m[367]&~m[368]&~m[377])|(m[365]&~m[366]&m[367]&~m[368]&~m[377])|(~m[365]&m[366]&m[367]&~m[368]&~m[377])|(m[365]&m[366]&m[367]&~m[368]&~m[377])|(m[365]&m[366]&m[367]&m[368]&~m[377])|(m[365]&m[366]&~m[367]&~m[368]&m[377])|(m[365]&~m[366]&m[367]&~m[368]&m[377])|(~m[365]&m[366]&m[367]&~m[368]&m[377])|(m[365]&m[366]&m[367]&~m[368]&m[377])|(m[365]&m[366]&m[367]&m[368]&m[377]))):InitCond[692];
    m[374] = run?((((m[370]&~m[371]&~m[372]&~m[373]&~m[382])|(~m[370]&m[371]&~m[372]&~m[373]&~m[382])|(~m[370]&~m[371]&m[372]&~m[373]&~m[382])|(m[370]&m[371]&~m[372]&m[373]&~m[382])|(m[370]&~m[371]&m[372]&m[373]&~m[382])|(~m[370]&m[371]&m[372]&m[373]&~m[382]))&BiasedRNG[341])|(((m[370]&~m[371]&~m[372]&~m[373]&m[382])|(~m[370]&m[371]&~m[372]&~m[373]&m[382])|(~m[370]&~m[371]&m[372]&~m[373]&m[382])|(m[370]&m[371]&~m[372]&m[373]&m[382])|(m[370]&~m[371]&m[372]&m[373]&m[382])|(~m[370]&m[371]&m[372]&m[373]&m[382]))&~BiasedRNG[341])|((m[370]&m[371]&~m[372]&~m[373]&~m[382])|(m[370]&~m[371]&m[372]&~m[373]&~m[382])|(~m[370]&m[371]&m[372]&~m[373]&~m[382])|(m[370]&m[371]&m[372]&~m[373]&~m[382])|(m[370]&m[371]&m[372]&m[373]&~m[382])|(m[370]&m[371]&~m[372]&~m[373]&m[382])|(m[370]&~m[371]&m[372]&~m[373]&m[382])|(~m[370]&m[371]&m[372]&~m[373]&m[382])|(m[370]&m[371]&m[372]&~m[373]&m[382])|(m[370]&m[371]&m[372]&m[373]&m[382]))):InitCond[693];
    m[379] = run?((((m[375]&~m[376]&~m[377]&~m[378]&~m[392])|(~m[375]&m[376]&~m[377]&~m[378]&~m[392])|(~m[375]&~m[376]&m[377]&~m[378]&~m[392])|(m[375]&m[376]&~m[377]&m[378]&~m[392])|(m[375]&~m[376]&m[377]&m[378]&~m[392])|(~m[375]&m[376]&m[377]&m[378]&~m[392]))&BiasedRNG[342])|(((m[375]&~m[376]&~m[377]&~m[378]&m[392])|(~m[375]&m[376]&~m[377]&~m[378]&m[392])|(~m[375]&~m[376]&m[377]&~m[378]&m[392])|(m[375]&m[376]&~m[377]&m[378]&m[392])|(m[375]&~m[376]&m[377]&m[378]&m[392])|(~m[375]&m[376]&m[377]&m[378]&m[392]))&~BiasedRNG[342])|((m[375]&m[376]&~m[377]&~m[378]&~m[392])|(m[375]&~m[376]&m[377]&~m[378]&~m[392])|(~m[375]&m[376]&m[377]&~m[378]&~m[392])|(m[375]&m[376]&m[377]&~m[378]&~m[392])|(m[375]&m[376]&m[377]&m[378]&~m[392])|(m[375]&m[376]&~m[377]&~m[378]&m[392])|(m[375]&~m[376]&m[377]&~m[378]&m[392])|(~m[375]&m[376]&m[377]&~m[378]&m[392])|(m[375]&m[376]&m[377]&~m[378]&m[392])|(m[375]&m[376]&m[377]&m[378]&m[392]))):InitCond[694];
    m[384] = run?((((m[380]&~m[381]&~m[382]&~m[383]&~m[397])|(~m[380]&m[381]&~m[382]&~m[383]&~m[397])|(~m[380]&~m[381]&m[382]&~m[383]&~m[397])|(m[380]&m[381]&~m[382]&m[383]&~m[397])|(m[380]&~m[381]&m[382]&m[383]&~m[397])|(~m[380]&m[381]&m[382]&m[383]&~m[397]))&BiasedRNG[343])|(((m[380]&~m[381]&~m[382]&~m[383]&m[397])|(~m[380]&m[381]&~m[382]&~m[383]&m[397])|(~m[380]&~m[381]&m[382]&~m[383]&m[397])|(m[380]&m[381]&~m[382]&m[383]&m[397])|(m[380]&~m[381]&m[382]&m[383]&m[397])|(~m[380]&m[381]&m[382]&m[383]&m[397]))&~BiasedRNG[343])|((m[380]&m[381]&~m[382]&~m[383]&~m[397])|(m[380]&~m[381]&m[382]&~m[383]&~m[397])|(~m[380]&m[381]&m[382]&~m[383]&~m[397])|(m[380]&m[381]&m[382]&~m[383]&~m[397])|(m[380]&m[381]&m[382]&m[383]&~m[397])|(m[380]&m[381]&~m[382]&~m[383]&m[397])|(m[380]&~m[381]&m[382]&~m[383]&m[397])|(~m[380]&m[381]&m[382]&~m[383]&m[397])|(m[380]&m[381]&m[382]&~m[383]&m[397])|(m[380]&m[381]&m[382]&m[383]&m[397]))):InitCond[695];
    m[389] = run?((((m[385]&~m[386]&~m[387]&~m[388]&~m[402])|(~m[385]&m[386]&~m[387]&~m[388]&~m[402])|(~m[385]&~m[386]&m[387]&~m[388]&~m[402])|(m[385]&m[386]&~m[387]&m[388]&~m[402])|(m[385]&~m[386]&m[387]&m[388]&~m[402])|(~m[385]&m[386]&m[387]&m[388]&~m[402]))&BiasedRNG[344])|(((m[385]&~m[386]&~m[387]&~m[388]&m[402])|(~m[385]&m[386]&~m[387]&~m[388]&m[402])|(~m[385]&~m[386]&m[387]&~m[388]&m[402])|(m[385]&m[386]&~m[387]&m[388]&m[402])|(m[385]&~m[386]&m[387]&m[388]&m[402])|(~m[385]&m[386]&m[387]&m[388]&m[402]))&~BiasedRNG[344])|((m[385]&m[386]&~m[387]&~m[388]&~m[402])|(m[385]&~m[386]&m[387]&~m[388]&~m[402])|(~m[385]&m[386]&m[387]&~m[388]&~m[402])|(m[385]&m[386]&m[387]&~m[388]&~m[402])|(m[385]&m[386]&m[387]&m[388]&~m[402])|(m[385]&m[386]&~m[387]&~m[388]&m[402])|(m[385]&~m[386]&m[387]&~m[388]&m[402])|(~m[385]&m[386]&m[387]&~m[388]&m[402])|(m[385]&m[386]&m[387]&~m[388]&m[402])|(m[385]&m[386]&m[387]&m[388]&m[402]))):InitCond[696];
    m[394] = run?((((m[390]&~m[391]&~m[392]&~m[393]&~m[412])|(~m[390]&m[391]&~m[392]&~m[393]&~m[412])|(~m[390]&~m[391]&m[392]&~m[393]&~m[412])|(m[390]&m[391]&~m[392]&m[393]&~m[412])|(m[390]&~m[391]&m[392]&m[393]&~m[412])|(~m[390]&m[391]&m[392]&m[393]&~m[412]))&BiasedRNG[345])|(((m[390]&~m[391]&~m[392]&~m[393]&m[412])|(~m[390]&m[391]&~m[392]&~m[393]&m[412])|(~m[390]&~m[391]&m[392]&~m[393]&m[412])|(m[390]&m[391]&~m[392]&m[393]&m[412])|(m[390]&~m[391]&m[392]&m[393]&m[412])|(~m[390]&m[391]&m[392]&m[393]&m[412]))&~BiasedRNG[345])|((m[390]&m[391]&~m[392]&~m[393]&~m[412])|(m[390]&~m[391]&m[392]&~m[393]&~m[412])|(~m[390]&m[391]&m[392]&~m[393]&~m[412])|(m[390]&m[391]&m[392]&~m[393]&~m[412])|(m[390]&m[391]&m[392]&m[393]&~m[412])|(m[390]&m[391]&~m[392]&~m[393]&m[412])|(m[390]&~m[391]&m[392]&~m[393]&m[412])|(~m[390]&m[391]&m[392]&~m[393]&m[412])|(m[390]&m[391]&m[392]&~m[393]&m[412])|(m[390]&m[391]&m[392]&m[393]&m[412]))):InitCond[697];
    m[399] = run?((((m[395]&~m[396]&~m[397]&~m[398]&~m[417])|(~m[395]&m[396]&~m[397]&~m[398]&~m[417])|(~m[395]&~m[396]&m[397]&~m[398]&~m[417])|(m[395]&m[396]&~m[397]&m[398]&~m[417])|(m[395]&~m[396]&m[397]&m[398]&~m[417])|(~m[395]&m[396]&m[397]&m[398]&~m[417]))&BiasedRNG[346])|(((m[395]&~m[396]&~m[397]&~m[398]&m[417])|(~m[395]&m[396]&~m[397]&~m[398]&m[417])|(~m[395]&~m[396]&m[397]&~m[398]&m[417])|(m[395]&m[396]&~m[397]&m[398]&m[417])|(m[395]&~m[396]&m[397]&m[398]&m[417])|(~m[395]&m[396]&m[397]&m[398]&m[417]))&~BiasedRNG[346])|((m[395]&m[396]&~m[397]&~m[398]&~m[417])|(m[395]&~m[396]&m[397]&~m[398]&~m[417])|(~m[395]&m[396]&m[397]&~m[398]&~m[417])|(m[395]&m[396]&m[397]&~m[398]&~m[417])|(m[395]&m[396]&m[397]&m[398]&~m[417])|(m[395]&m[396]&~m[397]&~m[398]&m[417])|(m[395]&~m[396]&m[397]&~m[398]&m[417])|(~m[395]&m[396]&m[397]&~m[398]&m[417])|(m[395]&m[396]&m[397]&~m[398]&m[417])|(m[395]&m[396]&m[397]&m[398]&m[417]))):InitCond[698];
    m[404] = run?((((m[400]&~m[401]&~m[402]&~m[403]&~m[422])|(~m[400]&m[401]&~m[402]&~m[403]&~m[422])|(~m[400]&~m[401]&m[402]&~m[403]&~m[422])|(m[400]&m[401]&~m[402]&m[403]&~m[422])|(m[400]&~m[401]&m[402]&m[403]&~m[422])|(~m[400]&m[401]&m[402]&m[403]&~m[422]))&BiasedRNG[347])|(((m[400]&~m[401]&~m[402]&~m[403]&m[422])|(~m[400]&m[401]&~m[402]&~m[403]&m[422])|(~m[400]&~m[401]&m[402]&~m[403]&m[422])|(m[400]&m[401]&~m[402]&m[403]&m[422])|(m[400]&~m[401]&m[402]&m[403]&m[422])|(~m[400]&m[401]&m[402]&m[403]&m[422]))&~BiasedRNG[347])|((m[400]&m[401]&~m[402]&~m[403]&~m[422])|(m[400]&~m[401]&m[402]&~m[403]&~m[422])|(~m[400]&m[401]&m[402]&~m[403]&~m[422])|(m[400]&m[401]&m[402]&~m[403]&~m[422])|(m[400]&m[401]&m[402]&m[403]&~m[422])|(m[400]&m[401]&~m[402]&~m[403]&m[422])|(m[400]&~m[401]&m[402]&~m[403]&m[422])|(~m[400]&m[401]&m[402]&~m[403]&m[422])|(m[400]&m[401]&m[402]&~m[403]&m[422])|(m[400]&m[401]&m[402]&m[403]&m[422]))):InitCond[699];
    m[409] = run?((((m[405]&~m[406]&~m[407]&~m[408]&~m[427])|(~m[405]&m[406]&~m[407]&~m[408]&~m[427])|(~m[405]&~m[406]&m[407]&~m[408]&~m[427])|(m[405]&m[406]&~m[407]&m[408]&~m[427])|(m[405]&~m[406]&m[407]&m[408]&~m[427])|(~m[405]&m[406]&m[407]&m[408]&~m[427]))&BiasedRNG[348])|(((m[405]&~m[406]&~m[407]&~m[408]&m[427])|(~m[405]&m[406]&~m[407]&~m[408]&m[427])|(~m[405]&~m[406]&m[407]&~m[408]&m[427])|(m[405]&m[406]&~m[407]&m[408]&m[427])|(m[405]&~m[406]&m[407]&m[408]&m[427])|(~m[405]&m[406]&m[407]&m[408]&m[427]))&~BiasedRNG[348])|((m[405]&m[406]&~m[407]&~m[408]&~m[427])|(m[405]&~m[406]&m[407]&~m[408]&~m[427])|(~m[405]&m[406]&m[407]&~m[408]&~m[427])|(m[405]&m[406]&m[407]&~m[408]&~m[427])|(m[405]&m[406]&m[407]&m[408]&~m[427])|(m[405]&m[406]&~m[407]&~m[408]&m[427])|(m[405]&~m[406]&m[407]&~m[408]&m[427])|(~m[405]&m[406]&m[407]&~m[408]&m[427])|(m[405]&m[406]&m[407]&~m[408]&m[427])|(m[405]&m[406]&m[407]&m[408]&m[427]))):InitCond[700];
    m[414] = run?((((m[410]&~m[411]&~m[412]&~m[413]&~m[437])|(~m[410]&m[411]&~m[412]&~m[413]&~m[437])|(~m[410]&~m[411]&m[412]&~m[413]&~m[437])|(m[410]&m[411]&~m[412]&m[413]&~m[437])|(m[410]&~m[411]&m[412]&m[413]&~m[437])|(~m[410]&m[411]&m[412]&m[413]&~m[437]))&BiasedRNG[349])|(((m[410]&~m[411]&~m[412]&~m[413]&m[437])|(~m[410]&m[411]&~m[412]&~m[413]&m[437])|(~m[410]&~m[411]&m[412]&~m[413]&m[437])|(m[410]&m[411]&~m[412]&m[413]&m[437])|(m[410]&~m[411]&m[412]&m[413]&m[437])|(~m[410]&m[411]&m[412]&m[413]&m[437]))&~BiasedRNG[349])|((m[410]&m[411]&~m[412]&~m[413]&~m[437])|(m[410]&~m[411]&m[412]&~m[413]&~m[437])|(~m[410]&m[411]&m[412]&~m[413]&~m[437])|(m[410]&m[411]&m[412]&~m[413]&~m[437])|(m[410]&m[411]&m[412]&m[413]&~m[437])|(m[410]&m[411]&~m[412]&~m[413]&m[437])|(m[410]&~m[411]&m[412]&~m[413]&m[437])|(~m[410]&m[411]&m[412]&~m[413]&m[437])|(m[410]&m[411]&m[412]&~m[413]&m[437])|(m[410]&m[411]&m[412]&m[413]&m[437]))):InitCond[701];
    m[419] = run?((((m[415]&~m[416]&~m[417]&~m[418]&~m[442])|(~m[415]&m[416]&~m[417]&~m[418]&~m[442])|(~m[415]&~m[416]&m[417]&~m[418]&~m[442])|(m[415]&m[416]&~m[417]&m[418]&~m[442])|(m[415]&~m[416]&m[417]&m[418]&~m[442])|(~m[415]&m[416]&m[417]&m[418]&~m[442]))&BiasedRNG[350])|(((m[415]&~m[416]&~m[417]&~m[418]&m[442])|(~m[415]&m[416]&~m[417]&~m[418]&m[442])|(~m[415]&~m[416]&m[417]&~m[418]&m[442])|(m[415]&m[416]&~m[417]&m[418]&m[442])|(m[415]&~m[416]&m[417]&m[418]&m[442])|(~m[415]&m[416]&m[417]&m[418]&m[442]))&~BiasedRNG[350])|((m[415]&m[416]&~m[417]&~m[418]&~m[442])|(m[415]&~m[416]&m[417]&~m[418]&~m[442])|(~m[415]&m[416]&m[417]&~m[418]&~m[442])|(m[415]&m[416]&m[417]&~m[418]&~m[442])|(m[415]&m[416]&m[417]&m[418]&~m[442])|(m[415]&m[416]&~m[417]&~m[418]&m[442])|(m[415]&~m[416]&m[417]&~m[418]&m[442])|(~m[415]&m[416]&m[417]&~m[418]&m[442])|(m[415]&m[416]&m[417]&~m[418]&m[442])|(m[415]&m[416]&m[417]&m[418]&m[442]))):InitCond[702];
    m[424] = run?((((m[420]&~m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&~m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&~m[422]&m[423]&~m[447])|(m[420]&~m[421]&m[422]&m[423]&~m[447])|(~m[420]&m[421]&m[422]&m[423]&~m[447]))&BiasedRNG[351])|(((m[420]&~m[421]&~m[422]&~m[423]&m[447])|(~m[420]&m[421]&~m[422]&~m[423]&m[447])|(~m[420]&~m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&~m[422]&m[423]&m[447])|(m[420]&~m[421]&m[422]&m[423]&m[447])|(~m[420]&m[421]&m[422]&m[423]&m[447]))&~BiasedRNG[351])|((m[420]&m[421]&~m[422]&~m[423]&~m[447])|(m[420]&~m[421]&m[422]&~m[423]&~m[447])|(~m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&m[423]&~m[447])|(m[420]&m[421]&~m[422]&~m[423]&m[447])|(m[420]&~m[421]&m[422]&~m[423]&m[447])|(~m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&m[423]&m[447]))):InitCond[703];
    m[429] = run?((((m[425]&~m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&~m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&~m[427]&m[428]&~m[452])|(m[425]&~m[426]&m[427]&m[428]&~m[452])|(~m[425]&m[426]&m[427]&m[428]&~m[452]))&BiasedRNG[352])|(((m[425]&~m[426]&~m[427]&~m[428]&m[452])|(~m[425]&m[426]&~m[427]&~m[428]&m[452])|(~m[425]&~m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&~m[427]&m[428]&m[452])|(m[425]&~m[426]&m[427]&m[428]&m[452])|(~m[425]&m[426]&m[427]&m[428]&m[452]))&~BiasedRNG[352])|((m[425]&m[426]&~m[427]&~m[428]&~m[452])|(m[425]&~m[426]&m[427]&~m[428]&~m[452])|(~m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&m[428]&~m[452])|(m[425]&m[426]&~m[427]&~m[428]&m[452])|(m[425]&~m[426]&m[427]&~m[428]&m[452])|(~m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&m[428]&m[452]))):InitCond[704];
    m[434] = run?((((m[430]&~m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&~m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&~m[432]&m[433]&~m[457])|(m[430]&~m[431]&m[432]&m[433]&~m[457])|(~m[430]&m[431]&m[432]&m[433]&~m[457]))&BiasedRNG[353])|(((m[430]&~m[431]&~m[432]&~m[433]&m[457])|(~m[430]&m[431]&~m[432]&~m[433]&m[457])|(~m[430]&~m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&~m[432]&m[433]&m[457])|(m[430]&~m[431]&m[432]&m[433]&m[457])|(~m[430]&m[431]&m[432]&m[433]&m[457]))&~BiasedRNG[353])|((m[430]&m[431]&~m[432]&~m[433]&~m[457])|(m[430]&~m[431]&m[432]&~m[433]&~m[457])|(~m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&m[433]&~m[457])|(m[430]&m[431]&~m[432]&~m[433]&m[457])|(m[430]&~m[431]&m[432]&~m[433]&m[457])|(~m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&m[433]&m[457]))):InitCond[705];
    m[439] = run?((((m[435]&~m[436]&~m[437]&~m[438]&~m[467])|(~m[435]&m[436]&~m[437]&~m[438]&~m[467])|(~m[435]&~m[436]&m[437]&~m[438]&~m[467])|(m[435]&m[436]&~m[437]&m[438]&~m[467])|(m[435]&~m[436]&m[437]&m[438]&~m[467])|(~m[435]&m[436]&m[437]&m[438]&~m[467]))&BiasedRNG[354])|(((m[435]&~m[436]&~m[437]&~m[438]&m[467])|(~m[435]&m[436]&~m[437]&~m[438]&m[467])|(~m[435]&~m[436]&m[437]&~m[438]&m[467])|(m[435]&m[436]&~m[437]&m[438]&m[467])|(m[435]&~m[436]&m[437]&m[438]&m[467])|(~m[435]&m[436]&m[437]&m[438]&m[467]))&~BiasedRNG[354])|((m[435]&m[436]&~m[437]&~m[438]&~m[467])|(m[435]&~m[436]&m[437]&~m[438]&~m[467])|(~m[435]&m[436]&m[437]&~m[438]&~m[467])|(m[435]&m[436]&m[437]&~m[438]&~m[467])|(m[435]&m[436]&m[437]&m[438]&~m[467])|(m[435]&m[436]&~m[437]&~m[438]&m[467])|(m[435]&~m[436]&m[437]&~m[438]&m[467])|(~m[435]&m[436]&m[437]&~m[438]&m[467])|(m[435]&m[436]&m[437]&~m[438]&m[467])|(m[435]&m[436]&m[437]&m[438]&m[467]))):InitCond[706];
    m[444] = run?((((m[440]&~m[441]&~m[442]&~m[443]&~m[472])|(~m[440]&m[441]&~m[442]&~m[443]&~m[472])|(~m[440]&~m[441]&m[442]&~m[443]&~m[472])|(m[440]&m[441]&~m[442]&m[443]&~m[472])|(m[440]&~m[441]&m[442]&m[443]&~m[472])|(~m[440]&m[441]&m[442]&m[443]&~m[472]))&BiasedRNG[355])|(((m[440]&~m[441]&~m[442]&~m[443]&m[472])|(~m[440]&m[441]&~m[442]&~m[443]&m[472])|(~m[440]&~m[441]&m[442]&~m[443]&m[472])|(m[440]&m[441]&~m[442]&m[443]&m[472])|(m[440]&~m[441]&m[442]&m[443]&m[472])|(~m[440]&m[441]&m[442]&m[443]&m[472]))&~BiasedRNG[355])|((m[440]&m[441]&~m[442]&~m[443]&~m[472])|(m[440]&~m[441]&m[442]&~m[443]&~m[472])|(~m[440]&m[441]&m[442]&~m[443]&~m[472])|(m[440]&m[441]&m[442]&~m[443]&~m[472])|(m[440]&m[441]&m[442]&m[443]&~m[472])|(m[440]&m[441]&~m[442]&~m[443]&m[472])|(m[440]&~m[441]&m[442]&~m[443]&m[472])|(~m[440]&m[441]&m[442]&~m[443]&m[472])|(m[440]&m[441]&m[442]&~m[443]&m[472])|(m[440]&m[441]&m[442]&m[443]&m[472]))):InitCond[707];
    m[449] = run?((((m[445]&~m[446]&~m[447]&~m[448]&~m[477])|(~m[445]&m[446]&~m[447]&~m[448]&~m[477])|(~m[445]&~m[446]&m[447]&~m[448]&~m[477])|(m[445]&m[446]&~m[447]&m[448]&~m[477])|(m[445]&~m[446]&m[447]&m[448]&~m[477])|(~m[445]&m[446]&m[447]&m[448]&~m[477]))&BiasedRNG[356])|(((m[445]&~m[446]&~m[447]&~m[448]&m[477])|(~m[445]&m[446]&~m[447]&~m[448]&m[477])|(~m[445]&~m[446]&m[447]&~m[448]&m[477])|(m[445]&m[446]&~m[447]&m[448]&m[477])|(m[445]&~m[446]&m[447]&m[448]&m[477])|(~m[445]&m[446]&m[447]&m[448]&m[477]))&~BiasedRNG[356])|((m[445]&m[446]&~m[447]&~m[448]&~m[477])|(m[445]&~m[446]&m[447]&~m[448]&~m[477])|(~m[445]&m[446]&m[447]&~m[448]&~m[477])|(m[445]&m[446]&m[447]&~m[448]&~m[477])|(m[445]&m[446]&m[447]&m[448]&~m[477])|(m[445]&m[446]&~m[447]&~m[448]&m[477])|(m[445]&~m[446]&m[447]&~m[448]&m[477])|(~m[445]&m[446]&m[447]&~m[448]&m[477])|(m[445]&m[446]&m[447]&~m[448]&m[477])|(m[445]&m[446]&m[447]&m[448]&m[477]))):InitCond[708];
    m[454] = run?((((m[450]&~m[451]&~m[452]&~m[453]&~m[482])|(~m[450]&m[451]&~m[452]&~m[453]&~m[482])|(~m[450]&~m[451]&m[452]&~m[453]&~m[482])|(m[450]&m[451]&~m[452]&m[453]&~m[482])|(m[450]&~m[451]&m[452]&m[453]&~m[482])|(~m[450]&m[451]&m[452]&m[453]&~m[482]))&BiasedRNG[357])|(((m[450]&~m[451]&~m[452]&~m[453]&m[482])|(~m[450]&m[451]&~m[452]&~m[453]&m[482])|(~m[450]&~m[451]&m[452]&~m[453]&m[482])|(m[450]&m[451]&~m[452]&m[453]&m[482])|(m[450]&~m[451]&m[452]&m[453]&m[482])|(~m[450]&m[451]&m[452]&m[453]&m[482]))&~BiasedRNG[357])|((m[450]&m[451]&~m[452]&~m[453]&~m[482])|(m[450]&~m[451]&m[452]&~m[453]&~m[482])|(~m[450]&m[451]&m[452]&~m[453]&~m[482])|(m[450]&m[451]&m[452]&~m[453]&~m[482])|(m[450]&m[451]&m[452]&m[453]&~m[482])|(m[450]&m[451]&~m[452]&~m[453]&m[482])|(m[450]&~m[451]&m[452]&~m[453]&m[482])|(~m[450]&m[451]&m[452]&~m[453]&m[482])|(m[450]&m[451]&m[452]&~m[453]&m[482])|(m[450]&m[451]&m[452]&m[453]&m[482]))):InitCond[709];
    m[459] = run?((((m[455]&~m[456]&~m[457]&~m[458]&~m[487])|(~m[455]&m[456]&~m[457]&~m[458]&~m[487])|(~m[455]&~m[456]&m[457]&~m[458]&~m[487])|(m[455]&m[456]&~m[457]&m[458]&~m[487])|(m[455]&~m[456]&m[457]&m[458]&~m[487])|(~m[455]&m[456]&m[457]&m[458]&~m[487]))&BiasedRNG[358])|(((m[455]&~m[456]&~m[457]&~m[458]&m[487])|(~m[455]&m[456]&~m[457]&~m[458]&m[487])|(~m[455]&~m[456]&m[457]&~m[458]&m[487])|(m[455]&m[456]&~m[457]&m[458]&m[487])|(m[455]&~m[456]&m[457]&m[458]&m[487])|(~m[455]&m[456]&m[457]&m[458]&m[487]))&~BiasedRNG[358])|((m[455]&m[456]&~m[457]&~m[458]&~m[487])|(m[455]&~m[456]&m[457]&~m[458]&~m[487])|(~m[455]&m[456]&m[457]&~m[458]&~m[487])|(m[455]&m[456]&m[457]&~m[458]&~m[487])|(m[455]&m[456]&m[457]&m[458]&~m[487])|(m[455]&m[456]&~m[457]&~m[458]&m[487])|(m[455]&~m[456]&m[457]&~m[458]&m[487])|(~m[455]&m[456]&m[457]&~m[458]&m[487])|(m[455]&m[456]&m[457]&~m[458]&m[487])|(m[455]&m[456]&m[457]&m[458]&m[487]))):InitCond[710];
    m[464] = run?((((m[460]&~m[461]&~m[462]&~m[463]&~m[492])|(~m[460]&m[461]&~m[462]&~m[463]&~m[492])|(~m[460]&~m[461]&m[462]&~m[463]&~m[492])|(m[460]&m[461]&~m[462]&m[463]&~m[492])|(m[460]&~m[461]&m[462]&m[463]&~m[492])|(~m[460]&m[461]&m[462]&m[463]&~m[492]))&BiasedRNG[359])|(((m[460]&~m[461]&~m[462]&~m[463]&m[492])|(~m[460]&m[461]&~m[462]&~m[463]&m[492])|(~m[460]&~m[461]&m[462]&~m[463]&m[492])|(m[460]&m[461]&~m[462]&m[463]&m[492])|(m[460]&~m[461]&m[462]&m[463]&m[492])|(~m[460]&m[461]&m[462]&m[463]&m[492]))&~BiasedRNG[359])|((m[460]&m[461]&~m[462]&~m[463]&~m[492])|(m[460]&~m[461]&m[462]&~m[463]&~m[492])|(~m[460]&m[461]&m[462]&~m[463]&~m[492])|(m[460]&m[461]&m[462]&~m[463]&~m[492])|(m[460]&m[461]&m[462]&m[463]&~m[492])|(m[460]&m[461]&~m[462]&~m[463]&m[492])|(m[460]&~m[461]&m[462]&~m[463]&m[492])|(~m[460]&m[461]&m[462]&~m[463]&m[492])|(m[460]&m[461]&m[462]&~m[463]&m[492])|(m[460]&m[461]&m[462]&m[463]&m[492]))):InitCond[711];
    m[469] = run?((((m[465]&~m[466]&~m[467]&~m[468]&~m[502])|(~m[465]&m[466]&~m[467]&~m[468]&~m[502])|(~m[465]&~m[466]&m[467]&~m[468]&~m[502])|(m[465]&m[466]&~m[467]&m[468]&~m[502])|(m[465]&~m[466]&m[467]&m[468]&~m[502])|(~m[465]&m[466]&m[467]&m[468]&~m[502]))&BiasedRNG[360])|(((m[465]&~m[466]&~m[467]&~m[468]&m[502])|(~m[465]&m[466]&~m[467]&~m[468]&m[502])|(~m[465]&~m[466]&m[467]&~m[468]&m[502])|(m[465]&m[466]&~m[467]&m[468]&m[502])|(m[465]&~m[466]&m[467]&m[468]&m[502])|(~m[465]&m[466]&m[467]&m[468]&m[502]))&~BiasedRNG[360])|((m[465]&m[466]&~m[467]&~m[468]&~m[502])|(m[465]&~m[466]&m[467]&~m[468]&~m[502])|(~m[465]&m[466]&m[467]&~m[468]&~m[502])|(m[465]&m[466]&m[467]&~m[468]&~m[502])|(m[465]&m[466]&m[467]&m[468]&~m[502])|(m[465]&m[466]&~m[467]&~m[468]&m[502])|(m[465]&~m[466]&m[467]&~m[468]&m[502])|(~m[465]&m[466]&m[467]&~m[468]&m[502])|(m[465]&m[466]&m[467]&~m[468]&m[502])|(m[465]&m[466]&m[467]&m[468]&m[502]))):InitCond[712];
    m[474] = run?((((m[470]&~m[471]&~m[472]&~m[473]&~m[507])|(~m[470]&m[471]&~m[472]&~m[473]&~m[507])|(~m[470]&~m[471]&m[472]&~m[473]&~m[507])|(m[470]&m[471]&~m[472]&m[473]&~m[507])|(m[470]&~m[471]&m[472]&m[473]&~m[507])|(~m[470]&m[471]&m[472]&m[473]&~m[507]))&BiasedRNG[361])|(((m[470]&~m[471]&~m[472]&~m[473]&m[507])|(~m[470]&m[471]&~m[472]&~m[473]&m[507])|(~m[470]&~m[471]&m[472]&~m[473]&m[507])|(m[470]&m[471]&~m[472]&m[473]&m[507])|(m[470]&~m[471]&m[472]&m[473]&m[507])|(~m[470]&m[471]&m[472]&m[473]&m[507]))&~BiasedRNG[361])|((m[470]&m[471]&~m[472]&~m[473]&~m[507])|(m[470]&~m[471]&m[472]&~m[473]&~m[507])|(~m[470]&m[471]&m[472]&~m[473]&~m[507])|(m[470]&m[471]&m[472]&~m[473]&~m[507])|(m[470]&m[471]&m[472]&m[473]&~m[507])|(m[470]&m[471]&~m[472]&~m[473]&m[507])|(m[470]&~m[471]&m[472]&~m[473]&m[507])|(~m[470]&m[471]&m[472]&~m[473]&m[507])|(m[470]&m[471]&m[472]&~m[473]&m[507])|(m[470]&m[471]&m[472]&m[473]&m[507]))):InitCond[713];
    m[479] = run?((((m[475]&~m[476]&~m[477]&~m[478]&~m[512])|(~m[475]&m[476]&~m[477]&~m[478]&~m[512])|(~m[475]&~m[476]&m[477]&~m[478]&~m[512])|(m[475]&m[476]&~m[477]&m[478]&~m[512])|(m[475]&~m[476]&m[477]&m[478]&~m[512])|(~m[475]&m[476]&m[477]&m[478]&~m[512]))&BiasedRNG[362])|(((m[475]&~m[476]&~m[477]&~m[478]&m[512])|(~m[475]&m[476]&~m[477]&~m[478]&m[512])|(~m[475]&~m[476]&m[477]&~m[478]&m[512])|(m[475]&m[476]&~m[477]&m[478]&m[512])|(m[475]&~m[476]&m[477]&m[478]&m[512])|(~m[475]&m[476]&m[477]&m[478]&m[512]))&~BiasedRNG[362])|((m[475]&m[476]&~m[477]&~m[478]&~m[512])|(m[475]&~m[476]&m[477]&~m[478]&~m[512])|(~m[475]&m[476]&m[477]&~m[478]&~m[512])|(m[475]&m[476]&m[477]&~m[478]&~m[512])|(m[475]&m[476]&m[477]&m[478]&~m[512])|(m[475]&m[476]&~m[477]&~m[478]&m[512])|(m[475]&~m[476]&m[477]&~m[478]&m[512])|(~m[475]&m[476]&m[477]&~m[478]&m[512])|(m[475]&m[476]&m[477]&~m[478]&m[512])|(m[475]&m[476]&m[477]&m[478]&m[512]))):InitCond[714];
    m[484] = run?((((m[480]&~m[481]&~m[482]&~m[483]&~m[517])|(~m[480]&m[481]&~m[482]&~m[483]&~m[517])|(~m[480]&~m[481]&m[482]&~m[483]&~m[517])|(m[480]&m[481]&~m[482]&m[483]&~m[517])|(m[480]&~m[481]&m[482]&m[483]&~m[517])|(~m[480]&m[481]&m[482]&m[483]&~m[517]))&BiasedRNG[363])|(((m[480]&~m[481]&~m[482]&~m[483]&m[517])|(~m[480]&m[481]&~m[482]&~m[483]&m[517])|(~m[480]&~m[481]&m[482]&~m[483]&m[517])|(m[480]&m[481]&~m[482]&m[483]&m[517])|(m[480]&~m[481]&m[482]&m[483]&m[517])|(~m[480]&m[481]&m[482]&m[483]&m[517]))&~BiasedRNG[363])|((m[480]&m[481]&~m[482]&~m[483]&~m[517])|(m[480]&~m[481]&m[482]&~m[483]&~m[517])|(~m[480]&m[481]&m[482]&~m[483]&~m[517])|(m[480]&m[481]&m[482]&~m[483]&~m[517])|(m[480]&m[481]&m[482]&m[483]&~m[517])|(m[480]&m[481]&~m[482]&~m[483]&m[517])|(m[480]&~m[481]&m[482]&~m[483]&m[517])|(~m[480]&m[481]&m[482]&~m[483]&m[517])|(m[480]&m[481]&m[482]&~m[483]&m[517])|(m[480]&m[481]&m[482]&m[483]&m[517]))):InitCond[715];
    m[489] = run?((((m[485]&~m[486]&~m[487]&~m[488]&~m[522])|(~m[485]&m[486]&~m[487]&~m[488]&~m[522])|(~m[485]&~m[486]&m[487]&~m[488]&~m[522])|(m[485]&m[486]&~m[487]&m[488]&~m[522])|(m[485]&~m[486]&m[487]&m[488]&~m[522])|(~m[485]&m[486]&m[487]&m[488]&~m[522]))&BiasedRNG[364])|(((m[485]&~m[486]&~m[487]&~m[488]&m[522])|(~m[485]&m[486]&~m[487]&~m[488]&m[522])|(~m[485]&~m[486]&m[487]&~m[488]&m[522])|(m[485]&m[486]&~m[487]&m[488]&m[522])|(m[485]&~m[486]&m[487]&m[488]&m[522])|(~m[485]&m[486]&m[487]&m[488]&m[522]))&~BiasedRNG[364])|((m[485]&m[486]&~m[487]&~m[488]&~m[522])|(m[485]&~m[486]&m[487]&~m[488]&~m[522])|(~m[485]&m[486]&m[487]&~m[488]&~m[522])|(m[485]&m[486]&m[487]&~m[488]&~m[522])|(m[485]&m[486]&m[487]&m[488]&~m[522])|(m[485]&m[486]&~m[487]&~m[488]&m[522])|(m[485]&~m[486]&m[487]&~m[488]&m[522])|(~m[485]&m[486]&m[487]&~m[488]&m[522])|(m[485]&m[486]&m[487]&~m[488]&m[522])|(m[485]&m[486]&m[487]&m[488]&m[522]))):InitCond[716];
    m[494] = run?((((m[490]&~m[491]&~m[492]&~m[493]&~m[527])|(~m[490]&m[491]&~m[492]&~m[493]&~m[527])|(~m[490]&~m[491]&m[492]&~m[493]&~m[527])|(m[490]&m[491]&~m[492]&m[493]&~m[527])|(m[490]&~m[491]&m[492]&m[493]&~m[527])|(~m[490]&m[491]&m[492]&m[493]&~m[527]))&BiasedRNG[365])|(((m[490]&~m[491]&~m[492]&~m[493]&m[527])|(~m[490]&m[491]&~m[492]&~m[493]&m[527])|(~m[490]&~m[491]&m[492]&~m[493]&m[527])|(m[490]&m[491]&~m[492]&m[493]&m[527])|(m[490]&~m[491]&m[492]&m[493]&m[527])|(~m[490]&m[491]&m[492]&m[493]&m[527]))&~BiasedRNG[365])|((m[490]&m[491]&~m[492]&~m[493]&~m[527])|(m[490]&~m[491]&m[492]&~m[493]&~m[527])|(~m[490]&m[491]&m[492]&~m[493]&~m[527])|(m[490]&m[491]&m[492]&~m[493]&~m[527])|(m[490]&m[491]&m[492]&m[493]&~m[527])|(m[490]&m[491]&~m[492]&~m[493]&m[527])|(m[490]&~m[491]&m[492]&~m[493]&m[527])|(~m[490]&m[491]&m[492]&~m[493]&m[527])|(m[490]&m[491]&m[492]&~m[493]&m[527])|(m[490]&m[491]&m[492]&m[493]&m[527]))):InitCond[717];
    m[499] = run?((((m[495]&~m[496]&~m[497]&~m[498]&~m[532])|(~m[495]&m[496]&~m[497]&~m[498]&~m[532])|(~m[495]&~m[496]&m[497]&~m[498]&~m[532])|(m[495]&m[496]&~m[497]&m[498]&~m[532])|(m[495]&~m[496]&m[497]&m[498]&~m[532])|(~m[495]&m[496]&m[497]&m[498]&~m[532]))&BiasedRNG[366])|(((m[495]&~m[496]&~m[497]&~m[498]&m[532])|(~m[495]&m[496]&~m[497]&~m[498]&m[532])|(~m[495]&~m[496]&m[497]&~m[498]&m[532])|(m[495]&m[496]&~m[497]&m[498]&m[532])|(m[495]&~m[496]&m[497]&m[498]&m[532])|(~m[495]&m[496]&m[497]&m[498]&m[532]))&~BiasedRNG[366])|((m[495]&m[496]&~m[497]&~m[498]&~m[532])|(m[495]&~m[496]&m[497]&~m[498]&~m[532])|(~m[495]&m[496]&m[497]&~m[498]&~m[532])|(m[495]&m[496]&m[497]&~m[498]&~m[532])|(m[495]&m[496]&m[497]&m[498]&~m[532])|(m[495]&m[496]&~m[497]&~m[498]&m[532])|(m[495]&~m[496]&m[497]&~m[498]&m[532])|(~m[495]&m[496]&m[497]&~m[498]&m[532])|(m[495]&m[496]&m[497]&~m[498]&m[532])|(m[495]&m[496]&m[497]&m[498]&m[532]))):InitCond[718];
    m[504] = run?((((m[500]&~m[501]&~m[502]&~m[503]&~m[542])|(~m[500]&m[501]&~m[502]&~m[503]&~m[542])|(~m[500]&~m[501]&m[502]&~m[503]&~m[542])|(m[500]&m[501]&~m[502]&m[503]&~m[542])|(m[500]&~m[501]&m[502]&m[503]&~m[542])|(~m[500]&m[501]&m[502]&m[503]&~m[542]))&BiasedRNG[367])|(((m[500]&~m[501]&~m[502]&~m[503]&m[542])|(~m[500]&m[501]&~m[502]&~m[503]&m[542])|(~m[500]&~m[501]&m[502]&~m[503]&m[542])|(m[500]&m[501]&~m[502]&m[503]&m[542])|(m[500]&~m[501]&m[502]&m[503]&m[542])|(~m[500]&m[501]&m[502]&m[503]&m[542]))&~BiasedRNG[367])|((m[500]&m[501]&~m[502]&~m[503]&~m[542])|(m[500]&~m[501]&m[502]&~m[503]&~m[542])|(~m[500]&m[501]&m[502]&~m[503]&~m[542])|(m[500]&m[501]&m[502]&~m[503]&~m[542])|(m[500]&m[501]&m[502]&m[503]&~m[542])|(m[500]&m[501]&~m[502]&~m[503]&m[542])|(m[500]&~m[501]&m[502]&~m[503]&m[542])|(~m[500]&m[501]&m[502]&~m[503]&m[542])|(m[500]&m[501]&m[502]&~m[503]&m[542])|(m[500]&m[501]&m[502]&m[503]&m[542]))):InitCond[719];
    m[509] = run?((((m[505]&~m[506]&~m[507]&~m[508]&~m[547])|(~m[505]&m[506]&~m[507]&~m[508]&~m[547])|(~m[505]&~m[506]&m[507]&~m[508]&~m[547])|(m[505]&m[506]&~m[507]&m[508]&~m[547])|(m[505]&~m[506]&m[507]&m[508]&~m[547])|(~m[505]&m[506]&m[507]&m[508]&~m[547]))&BiasedRNG[368])|(((m[505]&~m[506]&~m[507]&~m[508]&m[547])|(~m[505]&m[506]&~m[507]&~m[508]&m[547])|(~m[505]&~m[506]&m[507]&~m[508]&m[547])|(m[505]&m[506]&~m[507]&m[508]&m[547])|(m[505]&~m[506]&m[507]&m[508]&m[547])|(~m[505]&m[506]&m[507]&m[508]&m[547]))&~BiasedRNG[368])|((m[505]&m[506]&~m[507]&~m[508]&~m[547])|(m[505]&~m[506]&m[507]&~m[508]&~m[547])|(~m[505]&m[506]&m[507]&~m[508]&~m[547])|(m[505]&m[506]&m[507]&~m[508]&~m[547])|(m[505]&m[506]&m[507]&m[508]&~m[547])|(m[505]&m[506]&~m[507]&~m[508]&m[547])|(m[505]&~m[506]&m[507]&~m[508]&m[547])|(~m[505]&m[506]&m[507]&~m[508]&m[547])|(m[505]&m[506]&m[507]&~m[508]&m[547])|(m[505]&m[506]&m[507]&m[508]&m[547]))):InitCond[720];
    m[514] = run?((((m[510]&~m[511]&~m[512]&~m[513]&~m[552])|(~m[510]&m[511]&~m[512]&~m[513]&~m[552])|(~m[510]&~m[511]&m[512]&~m[513]&~m[552])|(m[510]&m[511]&~m[512]&m[513]&~m[552])|(m[510]&~m[511]&m[512]&m[513]&~m[552])|(~m[510]&m[511]&m[512]&m[513]&~m[552]))&BiasedRNG[369])|(((m[510]&~m[511]&~m[512]&~m[513]&m[552])|(~m[510]&m[511]&~m[512]&~m[513]&m[552])|(~m[510]&~m[511]&m[512]&~m[513]&m[552])|(m[510]&m[511]&~m[512]&m[513]&m[552])|(m[510]&~m[511]&m[512]&m[513]&m[552])|(~m[510]&m[511]&m[512]&m[513]&m[552]))&~BiasedRNG[369])|((m[510]&m[511]&~m[512]&~m[513]&~m[552])|(m[510]&~m[511]&m[512]&~m[513]&~m[552])|(~m[510]&m[511]&m[512]&~m[513]&~m[552])|(m[510]&m[511]&m[512]&~m[513]&~m[552])|(m[510]&m[511]&m[512]&m[513]&~m[552])|(m[510]&m[511]&~m[512]&~m[513]&m[552])|(m[510]&~m[511]&m[512]&~m[513]&m[552])|(~m[510]&m[511]&m[512]&~m[513]&m[552])|(m[510]&m[511]&m[512]&~m[513]&m[552])|(m[510]&m[511]&m[512]&m[513]&m[552]))):InitCond[721];
    m[519] = run?((((m[515]&~m[516]&~m[517]&~m[518]&~m[557])|(~m[515]&m[516]&~m[517]&~m[518]&~m[557])|(~m[515]&~m[516]&m[517]&~m[518]&~m[557])|(m[515]&m[516]&~m[517]&m[518]&~m[557])|(m[515]&~m[516]&m[517]&m[518]&~m[557])|(~m[515]&m[516]&m[517]&m[518]&~m[557]))&BiasedRNG[370])|(((m[515]&~m[516]&~m[517]&~m[518]&m[557])|(~m[515]&m[516]&~m[517]&~m[518]&m[557])|(~m[515]&~m[516]&m[517]&~m[518]&m[557])|(m[515]&m[516]&~m[517]&m[518]&m[557])|(m[515]&~m[516]&m[517]&m[518]&m[557])|(~m[515]&m[516]&m[517]&m[518]&m[557]))&~BiasedRNG[370])|((m[515]&m[516]&~m[517]&~m[518]&~m[557])|(m[515]&~m[516]&m[517]&~m[518]&~m[557])|(~m[515]&m[516]&m[517]&~m[518]&~m[557])|(m[515]&m[516]&m[517]&~m[518]&~m[557])|(m[515]&m[516]&m[517]&m[518]&~m[557])|(m[515]&m[516]&~m[517]&~m[518]&m[557])|(m[515]&~m[516]&m[517]&~m[518]&m[557])|(~m[515]&m[516]&m[517]&~m[518]&m[557])|(m[515]&m[516]&m[517]&~m[518]&m[557])|(m[515]&m[516]&m[517]&m[518]&m[557]))):InitCond[722];
    m[524] = run?((((m[520]&~m[521]&~m[522]&~m[523]&~m[562])|(~m[520]&m[521]&~m[522]&~m[523]&~m[562])|(~m[520]&~m[521]&m[522]&~m[523]&~m[562])|(m[520]&m[521]&~m[522]&m[523]&~m[562])|(m[520]&~m[521]&m[522]&m[523]&~m[562])|(~m[520]&m[521]&m[522]&m[523]&~m[562]))&BiasedRNG[371])|(((m[520]&~m[521]&~m[522]&~m[523]&m[562])|(~m[520]&m[521]&~m[522]&~m[523]&m[562])|(~m[520]&~m[521]&m[522]&~m[523]&m[562])|(m[520]&m[521]&~m[522]&m[523]&m[562])|(m[520]&~m[521]&m[522]&m[523]&m[562])|(~m[520]&m[521]&m[522]&m[523]&m[562]))&~BiasedRNG[371])|((m[520]&m[521]&~m[522]&~m[523]&~m[562])|(m[520]&~m[521]&m[522]&~m[523]&~m[562])|(~m[520]&m[521]&m[522]&~m[523]&~m[562])|(m[520]&m[521]&m[522]&~m[523]&~m[562])|(m[520]&m[521]&m[522]&m[523]&~m[562])|(m[520]&m[521]&~m[522]&~m[523]&m[562])|(m[520]&~m[521]&m[522]&~m[523]&m[562])|(~m[520]&m[521]&m[522]&~m[523]&m[562])|(m[520]&m[521]&m[522]&~m[523]&m[562])|(m[520]&m[521]&m[522]&m[523]&m[562]))):InitCond[723];
    m[529] = run?((((m[525]&~m[526]&~m[527]&~m[528]&~m[567])|(~m[525]&m[526]&~m[527]&~m[528]&~m[567])|(~m[525]&~m[526]&m[527]&~m[528]&~m[567])|(m[525]&m[526]&~m[527]&m[528]&~m[567])|(m[525]&~m[526]&m[527]&m[528]&~m[567])|(~m[525]&m[526]&m[527]&m[528]&~m[567]))&BiasedRNG[372])|(((m[525]&~m[526]&~m[527]&~m[528]&m[567])|(~m[525]&m[526]&~m[527]&~m[528]&m[567])|(~m[525]&~m[526]&m[527]&~m[528]&m[567])|(m[525]&m[526]&~m[527]&m[528]&m[567])|(m[525]&~m[526]&m[527]&m[528]&m[567])|(~m[525]&m[526]&m[527]&m[528]&m[567]))&~BiasedRNG[372])|((m[525]&m[526]&~m[527]&~m[528]&~m[567])|(m[525]&~m[526]&m[527]&~m[528]&~m[567])|(~m[525]&m[526]&m[527]&~m[528]&~m[567])|(m[525]&m[526]&m[527]&~m[528]&~m[567])|(m[525]&m[526]&m[527]&m[528]&~m[567])|(m[525]&m[526]&~m[527]&~m[528]&m[567])|(m[525]&~m[526]&m[527]&~m[528]&m[567])|(~m[525]&m[526]&m[527]&~m[528]&m[567])|(m[525]&m[526]&m[527]&~m[528]&m[567])|(m[525]&m[526]&m[527]&m[528]&m[567]))):InitCond[724];
    m[534] = run?((((m[530]&~m[531]&~m[532]&~m[533]&~m[572])|(~m[530]&m[531]&~m[532]&~m[533]&~m[572])|(~m[530]&~m[531]&m[532]&~m[533]&~m[572])|(m[530]&m[531]&~m[532]&m[533]&~m[572])|(m[530]&~m[531]&m[532]&m[533]&~m[572])|(~m[530]&m[531]&m[532]&m[533]&~m[572]))&BiasedRNG[373])|(((m[530]&~m[531]&~m[532]&~m[533]&m[572])|(~m[530]&m[531]&~m[532]&~m[533]&m[572])|(~m[530]&~m[531]&m[532]&~m[533]&m[572])|(m[530]&m[531]&~m[532]&m[533]&m[572])|(m[530]&~m[531]&m[532]&m[533]&m[572])|(~m[530]&m[531]&m[532]&m[533]&m[572]))&~BiasedRNG[373])|((m[530]&m[531]&~m[532]&~m[533]&~m[572])|(m[530]&~m[531]&m[532]&~m[533]&~m[572])|(~m[530]&m[531]&m[532]&~m[533]&~m[572])|(m[530]&m[531]&m[532]&~m[533]&~m[572])|(m[530]&m[531]&m[532]&m[533]&~m[572])|(m[530]&m[531]&~m[532]&~m[533]&m[572])|(m[530]&~m[531]&m[532]&~m[533]&m[572])|(~m[530]&m[531]&m[532]&~m[533]&m[572])|(m[530]&m[531]&m[532]&~m[533]&m[572])|(m[530]&m[531]&m[532]&m[533]&m[572]))):InitCond[725];
    m[539] = run?((((m[535]&~m[536]&~m[537]&~m[538]&~m[577])|(~m[535]&m[536]&~m[537]&~m[538]&~m[577])|(~m[535]&~m[536]&m[537]&~m[538]&~m[577])|(m[535]&m[536]&~m[537]&m[538]&~m[577])|(m[535]&~m[536]&m[537]&m[538]&~m[577])|(~m[535]&m[536]&m[537]&m[538]&~m[577]))&BiasedRNG[374])|(((m[535]&~m[536]&~m[537]&~m[538]&m[577])|(~m[535]&m[536]&~m[537]&~m[538]&m[577])|(~m[535]&~m[536]&m[537]&~m[538]&m[577])|(m[535]&m[536]&~m[537]&m[538]&m[577])|(m[535]&~m[536]&m[537]&m[538]&m[577])|(~m[535]&m[536]&m[537]&m[538]&m[577]))&~BiasedRNG[374])|((m[535]&m[536]&~m[537]&~m[538]&~m[577])|(m[535]&~m[536]&m[537]&~m[538]&~m[577])|(~m[535]&m[536]&m[537]&~m[538]&~m[577])|(m[535]&m[536]&m[537]&~m[538]&~m[577])|(m[535]&m[536]&m[537]&m[538]&~m[577])|(m[535]&m[536]&~m[537]&~m[538]&m[577])|(m[535]&~m[536]&m[537]&~m[538]&m[577])|(~m[535]&m[536]&m[537]&~m[538]&m[577])|(m[535]&m[536]&m[537]&~m[538]&m[577])|(m[535]&m[536]&m[537]&m[538]&m[577]))):InitCond[726];
    m[544] = run?((((m[540]&~m[541]&~m[542]&~m[543]&~m[587])|(~m[540]&m[541]&~m[542]&~m[543]&~m[587])|(~m[540]&~m[541]&m[542]&~m[543]&~m[587])|(m[540]&m[541]&~m[542]&m[543]&~m[587])|(m[540]&~m[541]&m[542]&m[543]&~m[587])|(~m[540]&m[541]&m[542]&m[543]&~m[587]))&BiasedRNG[375])|(((m[540]&~m[541]&~m[542]&~m[543]&m[587])|(~m[540]&m[541]&~m[542]&~m[543]&m[587])|(~m[540]&~m[541]&m[542]&~m[543]&m[587])|(m[540]&m[541]&~m[542]&m[543]&m[587])|(m[540]&~m[541]&m[542]&m[543]&m[587])|(~m[540]&m[541]&m[542]&m[543]&m[587]))&~BiasedRNG[375])|((m[540]&m[541]&~m[542]&~m[543]&~m[587])|(m[540]&~m[541]&m[542]&~m[543]&~m[587])|(~m[540]&m[541]&m[542]&~m[543]&~m[587])|(m[540]&m[541]&m[542]&~m[543]&~m[587])|(m[540]&m[541]&m[542]&m[543]&~m[587])|(m[540]&m[541]&~m[542]&~m[543]&m[587])|(m[540]&~m[541]&m[542]&~m[543]&m[587])|(~m[540]&m[541]&m[542]&~m[543]&m[587])|(m[540]&m[541]&m[542]&~m[543]&m[587])|(m[540]&m[541]&m[542]&m[543]&m[587]))):InitCond[727];
    m[549] = run?((((m[545]&~m[546]&~m[547]&~m[548]&~m[592])|(~m[545]&m[546]&~m[547]&~m[548]&~m[592])|(~m[545]&~m[546]&m[547]&~m[548]&~m[592])|(m[545]&m[546]&~m[547]&m[548]&~m[592])|(m[545]&~m[546]&m[547]&m[548]&~m[592])|(~m[545]&m[546]&m[547]&m[548]&~m[592]))&BiasedRNG[376])|(((m[545]&~m[546]&~m[547]&~m[548]&m[592])|(~m[545]&m[546]&~m[547]&~m[548]&m[592])|(~m[545]&~m[546]&m[547]&~m[548]&m[592])|(m[545]&m[546]&~m[547]&m[548]&m[592])|(m[545]&~m[546]&m[547]&m[548]&m[592])|(~m[545]&m[546]&m[547]&m[548]&m[592]))&~BiasedRNG[376])|((m[545]&m[546]&~m[547]&~m[548]&~m[592])|(m[545]&~m[546]&m[547]&~m[548]&~m[592])|(~m[545]&m[546]&m[547]&~m[548]&~m[592])|(m[545]&m[546]&m[547]&~m[548]&~m[592])|(m[545]&m[546]&m[547]&m[548]&~m[592])|(m[545]&m[546]&~m[547]&~m[548]&m[592])|(m[545]&~m[546]&m[547]&~m[548]&m[592])|(~m[545]&m[546]&m[547]&~m[548]&m[592])|(m[545]&m[546]&m[547]&~m[548]&m[592])|(m[545]&m[546]&m[547]&m[548]&m[592]))):InitCond[728];
    m[554] = run?((((m[550]&~m[551]&~m[552]&~m[553]&~m[597])|(~m[550]&m[551]&~m[552]&~m[553]&~m[597])|(~m[550]&~m[551]&m[552]&~m[553]&~m[597])|(m[550]&m[551]&~m[552]&m[553]&~m[597])|(m[550]&~m[551]&m[552]&m[553]&~m[597])|(~m[550]&m[551]&m[552]&m[553]&~m[597]))&BiasedRNG[377])|(((m[550]&~m[551]&~m[552]&~m[553]&m[597])|(~m[550]&m[551]&~m[552]&~m[553]&m[597])|(~m[550]&~m[551]&m[552]&~m[553]&m[597])|(m[550]&m[551]&~m[552]&m[553]&m[597])|(m[550]&~m[551]&m[552]&m[553]&m[597])|(~m[550]&m[551]&m[552]&m[553]&m[597]))&~BiasedRNG[377])|((m[550]&m[551]&~m[552]&~m[553]&~m[597])|(m[550]&~m[551]&m[552]&~m[553]&~m[597])|(~m[550]&m[551]&m[552]&~m[553]&~m[597])|(m[550]&m[551]&m[552]&~m[553]&~m[597])|(m[550]&m[551]&m[552]&m[553]&~m[597])|(m[550]&m[551]&~m[552]&~m[553]&m[597])|(m[550]&~m[551]&m[552]&~m[553]&m[597])|(~m[550]&m[551]&m[552]&~m[553]&m[597])|(m[550]&m[551]&m[552]&~m[553]&m[597])|(m[550]&m[551]&m[552]&m[553]&m[597]))):InitCond[729];
    m[559] = run?((((m[555]&~m[556]&~m[557]&~m[558]&~m[602])|(~m[555]&m[556]&~m[557]&~m[558]&~m[602])|(~m[555]&~m[556]&m[557]&~m[558]&~m[602])|(m[555]&m[556]&~m[557]&m[558]&~m[602])|(m[555]&~m[556]&m[557]&m[558]&~m[602])|(~m[555]&m[556]&m[557]&m[558]&~m[602]))&BiasedRNG[378])|(((m[555]&~m[556]&~m[557]&~m[558]&m[602])|(~m[555]&m[556]&~m[557]&~m[558]&m[602])|(~m[555]&~m[556]&m[557]&~m[558]&m[602])|(m[555]&m[556]&~m[557]&m[558]&m[602])|(m[555]&~m[556]&m[557]&m[558]&m[602])|(~m[555]&m[556]&m[557]&m[558]&m[602]))&~BiasedRNG[378])|((m[555]&m[556]&~m[557]&~m[558]&~m[602])|(m[555]&~m[556]&m[557]&~m[558]&~m[602])|(~m[555]&m[556]&m[557]&~m[558]&~m[602])|(m[555]&m[556]&m[557]&~m[558]&~m[602])|(m[555]&m[556]&m[557]&m[558]&~m[602])|(m[555]&m[556]&~m[557]&~m[558]&m[602])|(m[555]&~m[556]&m[557]&~m[558]&m[602])|(~m[555]&m[556]&m[557]&~m[558]&m[602])|(m[555]&m[556]&m[557]&~m[558]&m[602])|(m[555]&m[556]&m[557]&m[558]&m[602]))):InitCond[730];
    m[564] = run?((((m[560]&~m[561]&~m[562]&~m[563]&~m[607])|(~m[560]&m[561]&~m[562]&~m[563]&~m[607])|(~m[560]&~m[561]&m[562]&~m[563]&~m[607])|(m[560]&m[561]&~m[562]&m[563]&~m[607])|(m[560]&~m[561]&m[562]&m[563]&~m[607])|(~m[560]&m[561]&m[562]&m[563]&~m[607]))&BiasedRNG[379])|(((m[560]&~m[561]&~m[562]&~m[563]&m[607])|(~m[560]&m[561]&~m[562]&~m[563]&m[607])|(~m[560]&~m[561]&m[562]&~m[563]&m[607])|(m[560]&m[561]&~m[562]&m[563]&m[607])|(m[560]&~m[561]&m[562]&m[563]&m[607])|(~m[560]&m[561]&m[562]&m[563]&m[607]))&~BiasedRNG[379])|((m[560]&m[561]&~m[562]&~m[563]&~m[607])|(m[560]&~m[561]&m[562]&~m[563]&~m[607])|(~m[560]&m[561]&m[562]&~m[563]&~m[607])|(m[560]&m[561]&m[562]&~m[563]&~m[607])|(m[560]&m[561]&m[562]&m[563]&~m[607])|(m[560]&m[561]&~m[562]&~m[563]&m[607])|(m[560]&~m[561]&m[562]&~m[563]&m[607])|(~m[560]&m[561]&m[562]&~m[563]&m[607])|(m[560]&m[561]&m[562]&~m[563]&m[607])|(m[560]&m[561]&m[562]&m[563]&m[607]))):InitCond[731];
    m[569] = run?((((m[565]&~m[566]&~m[567]&~m[568]&~m[612])|(~m[565]&m[566]&~m[567]&~m[568]&~m[612])|(~m[565]&~m[566]&m[567]&~m[568]&~m[612])|(m[565]&m[566]&~m[567]&m[568]&~m[612])|(m[565]&~m[566]&m[567]&m[568]&~m[612])|(~m[565]&m[566]&m[567]&m[568]&~m[612]))&BiasedRNG[380])|(((m[565]&~m[566]&~m[567]&~m[568]&m[612])|(~m[565]&m[566]&~m[567]&~m[568]&m[612])|(~m[565]&~m[566]&m[567]&~m[568]&m[612])|(m[565]&m[566]&~m[567]&m[568]&m[612])|(m[565]&~m[566]&m[567]&m[568]&m[612])|(~m[565]&m[566]&m[567]&m[568]&m[612]))&~BiasedRNG[380])|((m[565]&m[566]&~m[567]&~m[568]&~m[612])|(m[565]&~m[566]&m[567]&~m[568]&~m[612])|(~m[565]&m[566]&m[567]&~m[568]&~m[612])|(m[565]&m[566]&m[567]&~m[568]&~m[612])|(m[565]&m[566]&m[567]&m[568]&~m[612])|(m[565]&m[566]&~m[567]&~m[568]&m[612])|(m[565]&~m[566]&m[567]&~m[568]&m[612])|(~m[565]&m[566]&m[567]&~m[568]&m[612])|(m[565]&m[566]&m[567]&~m[568]&m[612])|(m[565]&m[566]&m[567]&m[568]&m[612]))):InitCond[732];
    m[574] = run?((((m[570]&~m[571]&~m[572]&~m[573]&~m[617])|(~m[570]&m[571]&~m[572]&~m[573]&~m[617])|(~m[570]&~m[571]&m[572]&~m[573]&~m[617])|(m[570]&m[571]&~m[572]&m[573]&~m[617])|(m[570]&~m[571]&m[572]&m[573]&~m[617])|(~m[570]&m[571]&m[572]&m[573]&~m[617]))&BiasedRNG[381])|(((m[570]&~m[571]&~m[572]&~m[573]&m[617])|(~m[570]&m[571]&~m[572]&~m[573]&m[617])|(~m[570]&~m[571]&m[572]&~m[573]&m[617])|(m[570]&m[571]&~m[572]&m[573]&m[617])|(m[570]&~m[571]&m[572]&m[573]&m[617])|(~m[570]&m[571]&m[572]&m[573]&m[617]))&~BiasedRNG[381])|((m[570]&m[571]&~m[572]&~m[573]&~m[617])|(m[570]&~m[571]&m[572]&~m[573]&~m[617])|(~m[570]&m[571]&m[572]&~m[573]&~m[617])|(m[570]&m[571]&m[572]&~m[573]&~m[617])|(m[570]&m[571]&m[572]&m[573]&~m[617])|(m[570]&m[571]&~m[572]&~m[573]&m[617])|(m[570]&~m[571]&m[572]&~m[573]&m[617])|(~m[570]&m[571]&m[572]&~m[573]&m[617])|(m[570]&m[571]&m[572]&~m[573]&m[617])|(m[570]&m[571]&m[572]&m[573]&m[617]))):InitCond[733];
    m[579] = run?((((m[575]&~m[576]&~m[577]&~m[578]&~m[622])|(~m[575]&m[576]&~m[577]&~m[578]&~m[622])|(~m[575]&~m[576]&m[577]&~m[578]&~m[622])|(m[575]&m[576]&~m[577]&m[578]&~m[622])|(m[575]&~m[576]&m[577]&m[578]&~m[622])|(~m[575]&m[576]&m[577]&m[578]&~m[622]))&BiasedRNG[382])|(((m[575]&~m[576]&~m[577]&~m[578]&m[622])|(~m[575]&m[576]&~m[577]&~m[578]&m[622])|(~m[575]&~m[576]&m[577]&~m[578]&m[622])|(m[575]&m[576]&~m[577]&m[578]&m[622])|(m[575]&~m[576]&m[577]&m[578]&m[622])|(~m[575]&m[576]&m[577]&m[578]&m[622]))&~BiasedRNG[382])|((m[575]&m[576]&~m[577]&~m[578]&~m[622])|(m[575]&~m[576]&m[577]&~m[578]&~m[622])|(~m[575]&m[576]&m[577]&~m[578]&~m[622])|(m[575]&m[576]&m[577]&~m[578]&~m[622])|(m[575]&m[576]&m[577]&m[578]&~m[622])|(m[575]&m[576]&~m[577]&~m[578]&m[622])|(m[575]&~m[576]&m[577]&~m[578]&m[622])|(~m[575]&m[576]&m[577]&~m[578]&m[622])|(m[575]&m[576]&m[577]&~m[578]&m[622])|(m[575]&m[576]&m[577]&m[578]&m[622]))):InitCond[734];
    m[584] = run?((((m[580]&~m[581]&~m[582]&~m[583]&~m[627])|(~m[580]&m[581]&~m[582]&~m[583]&~m[627])|(~m[580]&~m[581]&m[582]&~m[583]&~m[627])|(m[580]&m[581]&~m[582]&m[583]&~m[627])|(m[580]&~m[581]&m[582]&m[583]&~m[627])|(~m[580]&m[581]&m[582]&m[583]&~m[627]))&BiasedRNG[383])|(((m[580]&~m[581]&~m[582]&~m[583]&m[627])|(~m[580]&m[581]&~m[582]&~m[583]&m[627])|(~m[580]&~m[581]&m[582]&~m[583]&m[627])|(m[580]&m[581]&~m[582]&m[583]&m[627])|(m[580]&~m[581]&m[582]&m[583]&m[627])|(~m[580]&m[581]&m[582]&m[583]&m[627]))&~BiasedRNG[383])|((m[580]&m[581]&~m[582]&~m[583]&~m[627])|(m[580]&~m[581]&m[582]&~m[583]&~m[627])|(~m[580]&m[581]&m[582]&~m[583]&~m[627])|(m[580]&m[581]&m[582]&~m[583]&~m[627])|(m[580]&m[581]&m[582]&m[583]&~m[627])|(m[580]&m[581]&~m[582]&~m[583]&m[627])|(m[580]&~m[581]&m[582]&~m[583]&m[627])|(~m[580]&m[581]&m[582]&~m[583]&m[627])|(m[580]&m[581]&m[582]&~m[583]&m[627])|(m[580]&m[581]&m[582]&m[583]&m[627]))):InitCond[735];
    m[589] = run?((((m[585]&~m[586]&~m[587]&~m[588]&~m[630])|(~m[585]&m[586]&~m[587]&~m[588]&~m[630])|(~m[585]&~m[586]&m[587]&~m[588]&~m[630])|(m[585]&m[586]&~m[587]&m[588]&~m[630])|(m[585]&~m[586]&m[587]&m[588]&~m[630])|(~m[585]&m[586]&m[587]&m[588]&~m[630]))&BiasedRNG[384])|(((m[585]&~m[586]&~m[587]&~m[588]&m[630])|(~m[585]&m[586]&~m[587]&~m[588]&m[630])|(~m[585]&~m[586]&m[587]&~m[588]&m[630])|(m[585]&m[586]&~m[587]&m[588]&m[630])|(m[585]&~m[586]&m[587]&m[588]&m[630])|(~m[585]&m[586]&m[587]&m[588]&m[630]))&~BiasedRNG[384])|((m[585]&m[586]&~m[587]&~m[588]&~m[630])|(m[585]&~m[586]&m[587]&~m[588]&~m[630])|(~m[585]&m[586]&m[587]&~m[588]&~m[630])|(m[585]&m[586]&m[587]&~m[588]&~m[630])|(m[585]&m[586]&m[587]&m[588]&~m[630])|(m[585]&m[586]&~m[587]&~m[588]&m[630])|(m[585]&~m[586]&m[587]&~m[588]&m[630])|(~m[585]&m[586]&m[587]&~m[588]&m[630])|(m[585]&m[586]&m[587]&~m[588]&m[630])|(m[585]&m[586]&m[587]&m[588]&m[630]))):InitCond[736];
    m[594] = run?((((m[590]&~m[591]&~m[592]&~m[593]&~m[632])|(~m[590]&m[591]&~m[592]&~m[593]&~m[632])|(~m[590]&~m[591]&m[592]&~m[593]&~m[632])|(m[590]&m[591]&~m[592]&m[593]&~m[632])|(m[590]&~m[591]&m[592]&m[593]&~m[632])|(~m[590]&m[591]&m[592]&m[593]&~m[632]))&BiasedRNG[385])|(((m[590]&~m[591]&~m[592]&~m[593]&m[632])|(~m[590]&m[591]&~m[592]&~m[593]&m[632])|(~m[590]&~m[591]&m[592]&~m[593]&m[632])|(m[590]&m[591]&~m[592]&m[593]&m[632])|(m[590]&~m[591]&m[592]&m[593]&m[632])|(~m[590]&m[591]&m[592]&m[593]&m[632]))&~BiasedRNG[385])|((m[590]&m[591]&~m[592]&~m[593]&~m[632])|(m[590]&~m[591]&m[592]&~m[593]&~m[632])|(~m[590]&m[591]&m[592]&~m[593]&~m[632])|(m[590]&m[591]&m[592]&~m[593]&~m[632])|(m[590]&m[591]&m[592]&m[593]&~m[632])|(m[590]&m[591]&~m[592]&~m[593]&m[632])|(m[590]&~m[591]&m[592]&~m[593]&m[632])|(~m[590]&m[591]&m[592]&~m[593]&m[632])|(m[590]&m[591]&m[592]&~m[593]&m[632])|(m[590]&m[591]&m[592]&m[593]&m[632]))):InitCond[737];
    m[599] = run?((((m[595]&~m[596]&~m[597]&~m[598]&~m[637])|(~m[595]&m[596]&~m[597]&~m[598]&~m[637])|(~m[595]&~m[596]&m[597]&~m[598]&~m[637])|(m[595]&m[596]&~m[597]&m[598]&~m[637])|(m[595]&~m[596]&m[597]&m[598]&~m[637])|(~m[595]&m[596]&m[597]&m[598]&~m[637]))&BiasedRNG[386])|(((m[595]&~m[596]&~m[597]&~m[598]&m[637])|(~m[595]&m[596]&~m[597]&~m[598]&m[637])|(~m[595]&~m[596]&m[597]&~m[598]&m[637])|(m[595]&m[596]&~m[597]&m[598]&m[637])|(m[595]&~m[596]&m[597]&m[598]&m[637])|(~m[595]&m[596]&m[597]&m[598]&m[637]))&~BiasedRNG[386])|((m[595]&m[596]&~m[597]&~m[598]&~m[637])|(m[595]&~m[596]&m[597]&~m[598]&~m[637])|(~m[595]&m[596]&m[597]&~m[598]&~m[637])|(m[595]&m[596]&m[597]&~m[598]&~m[637])|(m[595]&m[596]&m[597]&m[598]&~m[637])|(m[595]&m[596]&~m[597]&~m[598]&m[637])|(m[595]&~m[596]&m[597]&~m[598]&m[637])|(~m[595]&m[596]&m[597]&~m[598]&m[637])|(m[595]&m[596]&m[597]&~m[598]&m[637])|(m[595]&m[596]&m[597]&m[598]&m[637]))):InitCond[738];
    m[604] = run?((((m[600]&~m[601]&~m[602]&~m[603]&~m[642])|(~m[600]&m[601]&~m[602]&~m[603]&~m[642])|(~m[600]&~m[601]&m[602]&~m[603]&~m[642])|(m[600]&m[601]&~m[602]&m[603]&~m[642])|(m[600]&~m[601]&m[602]&m[603]&~m[642])|(~m[600]&m[601]&m[602]&m[603]&~m[642]))&BiasedRNG[387])|(((m[600]&~m[601]&~m[602]&~m[603]&m[642])|(~m[600]&m[601]&~m[602]&~m[603]&m[642])|(~m[600]&~m[601]&m[602]&~m[603]&m[642])|(m[600]&m[601]&~m[602]&m[603]&m[642])|(m[600]&~m[601]&m[602]&m[603]&m[642])|(~m[600]&m[601]&m[602]&m[603]&m[642]))&~BiasedRNG[387])|((m[600]&m[601]&~m[602]&~m[603]&~m[642])|(m[600]&~m[601]&m[602]&~m[603]&~m[642])|(~m[600]&m[601]&m[602]&~m[603]&~m[642])|(m[600]&m[601]&m[602]&~m[603]&~m[642])|(m[600]&m[601]&m[602]&m[603]&~m[642])|(m[600]&m[601]&~m[602]&~m[603]&m[642])|(m[600]&~m[601]&m[602]&~m[603]&m[642])|(~m[600]&m[601]&m[602]&~m[603]&m[642])|(m[600]&m[601]&m[602]&~m[603]&m[642])|(m[600]&m[601]&m[602]&m[603]&m[642]))):InitCond[739];
    m[609] = run?((((m[605]&~m[606]&~m[607]&~m[608]&~m[647])|(~m[605]&m[606]&~m[607]&~m[608]&~m[647])|(~m[605]&~m[606]&m[607]&~m[608]&~m[647])|(m[605]&m[606]&~m[607]&m[608]&~m[647])|(m[605]&~m[606]&m[607]&m[608]&~m[647])|(~m[605]&m[606]&m[607]&m[608]&~m[647]))&BiasedRNG[388])|(((m[605]&~m[606]&~m[607]&~m[608]&m[647])|(~m[605]&m[606]&~m[607]&~m[608]&m[647])|(~m[605]&~m[606]&m[607]&~m[608]&m[647])|(m[605]&m[606]&~m[607]&m[608]&m[647])|(m[605]&~m[606]&m[607]&m[608]&m[647])|(~m[605]&m[606]&m[607]&m[608]&m[647]))&~BiasedRNG[388])|((m[605]&m[606]&~m[607]&~m[608]&~m[647])|(m[605]&~m[606]&m[607]&~m[608]&~m[647])|(~m[605]&m[606]&m[607]&~m[608]&~m[647])|(m[605]&m[606]&m[607]&~m[608]&~m[647])|(m[605]&m[606]&m[607]&m[608]&~m[647])|(m[605]&m[606]&~m[607]&~m[608]&m[647])|(m[605]&~m[606]&m[607]&~m[608]&m[647])|(~m[605]&m[606]&m[607]&~m[608]&m[647])|(m[605]&m[606]&m[607]&~m[608]&m[647])|(m[605]&m[606]&m[607]&m[608]&m[647]))):InitCond[740];
    m[614] = run?((((m[610]&~m[611]&~m[612]&~m[613]&~m[652])|(~m[610]&m[611]&~m[612]&~m[613]&~m[652])|(~m[610]&~m[611]&m[612]&~m[613]&~m[652])|(m[610]&m[611]&~m[612]&m[613]&~m[652])|(m[610]&~m[611]&m[612]&m[613]&~m[652])|(~m[610]&m[611]&m[612]&m[613]&~m[652]))&BiasedRNG[389])|(((m[610]&~m[611]&~m[612]&~m[613]&m[652])|(~m[610]&m[611]&~m[612]&~m[613]&m[652])|(~m[610]&~m[611]&m[612]&~m[613]&m[652])|(m[610]&m[611]&~m[612]&m[613]&m[652])|(m[610]&~m[611]&m[612]&m[613]&m[652])|(~m[610]&m[611]&m[612]&m[613]&m[652]))&~BiasedRNG[389])|((m[610]&m[611]&~m[612]&~m[613]&~m[652])|(m[610]&~m[611]&m[612]&~m[613]&~m[652])|(~m[610]&m[611]&m[612]&~m[613]&~m[652])|(m[610]&m[611]&m[612]&~m[613]&~m[652])|(m[610]&m[611]&m[612]&m[613]&~m[652])|(m[610]&m[611]&~m[612]&~m[613]&m[652])|(m[610]&~m[611]&m[612]&~m[613]&m[652])|(~m[610]&m[611]&m[612]&~m[613]&m[652])|(m[610]&m[611]&m[612]&~m[613]&m[652])|(m[610]&m[611]&m[612]&m[613]&m[652]))):InitCond[741];
    m[619] = run?((((m[615]&~m[616]&~m[617]&~m[618]&~m[657])|(~m[615]&m[616]&~m[617]&~m[618]&~m[657])|(~m[615]&~m[616]&m[617]&~m[618]&~m[657])|(m[615]&m[616]&~m[617]&m[618]&~m[657])|(m[615]&~m[616]&m[617]&m[618]&~m[657])|(~m[615]&m[616]&m[617]&m[618]&~m[657]))&BiasedRNG[390])|(((m[615]&~m[616]&~m[617]&~m[618]&m[657])|(~m[615]&m[616]&~m[617]&~m[618]&m[657])|(~m[615]&~m[616]&m[617]&~m[618]&m[657])|(m[615]&m[616]&~m[617]&m[618]&m[657])|(m[615]&~m[616]&m[617]&m[618]&m[657])|(~m[615]&m[616]&m[617]&m[618]&m[657]))&~BiasedRNG[390])|((m[615]&m[616]&~m[617]&~m[618]&~m[657])|(m[615]&~m[616]&m[617]&~m[618]&~m[657])|(~m[615]&m[616]&m[617]&~m[618]&~m[657])|(m[615]&m[616]&m[617]&~m[618]&~m[657])|(m[615]&m[616]&m[617]&m[618]&~m[657])|(m[615]&m[616]&~m[617]&~m[618]&m[657])|(m[615]&~m[616]&m[617]&~m[618]&m[657])|(~m[615]&m[616]&m[617]&~m[618]&m[657])|(m[615]&m[616]&m[617]&~m[618]&m[657])|(m[615]&m[616]&m[617]&m[618]&m[657]))):InitCond[742];
    m[624] = run?((((m[620]&~m[621]&~m[622]&~m[623]&~m[662])|(~m[620]&m[621]&~m[622]&~m[623]&~m[662])|(~m[620]&~m[621]&m[622]&~m[623]&~m[662])|(m[620]&m[621]&~m[622]&m[623]&~m[662])|(m[620]&~m[621]&m[622]&m[623]&~m[662])|(~m[620]&m[621]&m[622]&m[623]&~m[662]))&BiasedRNG[391])|(((m[620]&~m[621]&~m[622]&~m[623]&m[662])|(~m[620]&m[621]&~m[622]&~m[623]&m[662])|(~m[620]&~m[621]&m[622]&~m[623]&m[662])|(m[620]&m[621]&~m[622]&m[623]&m[662])|(m[620]&~m[621]&m[622]&m[623]&m[662])|(~m[620]&m[621]&m[622]&m[623]&m[662]))&~BiasedRNG[391])|((m[620]&m[621]&~m[622]&~m[623]&~m[662])|(m[620]&~m[621]&m[622]&~m[623]&~m[662])|(~m[620]&m[621]&m[622]&~m[623]&~m[662])|(m[620]&m[621]&m[622]&~m[623]&~m[662])|(m[620]&m[621]&m[622]&m[623]&~m[662])|(m[620]&m[621]&~m[622]&~m[623]&m[662])|(m[620]&~m[621]&m[622]&~m[623]&m[662])|(~m[620]&m[621]&m[622]&~m[623]&m[662])|(m[620]&m[621]&m[622]&~m[623]&m[662])|(m[620]&m[621]&m[622]&m[623]&m[662]))):InitCond[743];
    m[629] = run?((((m[625]&~m[626]&~m[627]&~m[628]&~m[667])|(~m[625]&m[626]&~m[627]&~m[628]&~m[667])|(~m[625]&~m[626]&m[627]&~m[628]&~m[667])|(m[625]&m[626]&~m[627]&m[628]&~m[667])|(m[625]&~m[626]&m[627]&m[628]&~m[667])|(~m[625]&m[626]&m[627]&m[628]&~m[667]))&BiasedRNG[392])|(((m[625]&~m[626]&~m[627]&~m[628]&m[667])|(~m[625]&m[626]&~m[627]&~m[628]&m[667])|(~m[625]&~m[626]&m[627]&~m[628]&m[667])|(m[625]&m[626]&~m[627]&m[628]&m[667])|(m[625]&~m[626]&m[627]&m[628]&m[667])|(~m[625]&m[626]&m[627]&m[628]&m[667]))&~BiasedRNG[392])|((m[625]&m[626]&~m[627]&~m[628]&~m[667])|(m[625]&~m[626]&m[627]&~m[628]&~m[667])|(~m[625]&m[626]&m[627]&~m[628]&~m[667])|(m[625]&m[626]&m[627]&~m[628]&~m[667])|(m[625]&m[626]&m[627]&m[628]&~m[667])|(m[625]&m[626]&~m[627]&~m[628]&m[667])|(m[625]&~m[626]&m[627]&~m[628]&m[667])|(~m[625]&m[626]&m[627]&~m[628]&m[667])|(m[625]&m[626]&m[627]&~m[628]&m[667])|(m[625]&m[626]&m[627]&m[628]&m[667]))):InitCond[744];
    m[634] = run?((((m[630]&~m[631]&~m[632]&~m[633]&~m[670])|(~m[630]&m[631]&~m[632]&~m[633]&~m[670])|(~m[630]&~m[631]&m[632]&~m[633]&~m[670])|(m[630]&m[631]&~m[632]&m[633]&~m[670])|(m[630]&~m[631]&m[632]&m[633]&~m[670])|(~m[630]&m[631]&m[632]&m[633]&~m[670]))&BiasedRNG[393])|(((m[630]&~m[631]&~m[632]&~m[633]&m[670])|(~m[630]&m[631]&~m[632]&~m[633]&m[670])|(~m[630]&~m[631]&m[632]&~m[633]&m[670])|(m[630]&m[631]&~m[632]&m[633]&m[670])|(m[630]&~m[631]&m[632]&m[633]&m[670])|(~m[630]&m[631]&m[632]&m[633]&m[670]))&~BiasedRNG[393])|((m[630]&m[631]&~m[632]&~m[633]&~m[670])|(m[630]&~m[631]&m[632]&~m[633]&~m[670])|(~m[630]&m[631]&m[632]&~m[633]&~m[670])|(m[630]&m[631]&m[632]&~m[633]&~m[670])|(m[630]&m[631]&m[632]&m[633]&~m[670])|(m[630]&m[631]&~m[632]&~m[633]&m[670])|(m[630]&~m[631]&m[632]&~m[633]&m[670])|(~m[630]&m[631]&m[632]&~m[633]&m[670])|(m[630]&m[631]&m[632]&~m[633]&m[670])|(m[630]&m[631]&m[632]&m[633]&m[670]))):InitCond[745];
    m[639] = run?((((m[635]&~m[636]&~m[637]&~m[638]&~m[672])|(~m[635]&m[636]&~m[637]&~m[638]&~m[672])|(~m[635]&~m[636]&m[637]&~m[638]&~m[672])|(m[635]&m[636]&~m[637]&m[638]&~m[672])|(m[635]&~m[636]&m[637]&m[638]&~m[672])|(~m[635]&m[636]&m[637]&m[638]&~m[672]))&BiasedRNG[394])|(((m[635]&~m[636]&~m[637]&~m[638]&m[672])|(~m[635]&m[636]&~m[637]&~m[638]&m[672])|(~m[635]&~m[636]&m[637]&~m[638]&m[672])|(m[635]&m[636]&~m[637]&m[638]&m[672])|(m[635]&~m[636]&m[637]&m[638]&m[672])|(~m[635]&m[636]&m[637]&m[638]&m[672]))&~BiasedRNG[394])|((m[635]&m[636]&~m[637]&~m[638]&~m[672])|(m[635]&~m[636]&m[637]&~m[638]&~m[672])|(~m[635]&m[636]&m[637]&~m[638]&~m[672])|(m[635]&m[636]&m[637]&~m[638]&~m[672])|(m[635]&m[636]&m[637]&m[638]&~m[672])|(m[635]&m[636]&~m[637]&~m[638]&m[672])|(m[635]&~m[636]&m[637]&~m[638]&m[672])|(~m[635]&m[636]&m[637]&~m[638]&m[672])|(m[635]&m[636]&m[637]&~m[638]&m[672])|(m[635]&m[636]&m[637]&m[638]&m[672]))):InitCond[746];
    m[644] = run?((((m[640]&~m[641]&~m[642]&~m[643]&~m[677])|(~m[640]&m[641]&~m[642]&~m[643]&~m[677])|(~m[640]&~m[641]&m[642]&~m[643]&~m[677])|(m[640]&m[641]&~m[642]&m[643]&~m[677])|(m[640]&~m[641]&m[642]&m[643]&~m[677])|(~m[640]&m[641]&m[642]&m[643]&~m[677]))&BiasedRNG[395])|(((m[640]&~m[641]&~m[642]&~m[643]&m[677])|(~m[640]&m[641]&~m[642]&~m[643]&m[677])|(~m[640]&~m[641]&m[642]&~m[643]&m[677])|(m[640]&m[641]&~m[642]&m[643]&m[677])|(m[640]&~m[641]&m[642]&m[643]&m[677])|(~m[640]&m[641]&m[642]&m[643]&m[677]))&~BiasedRNG[395])|((m[640]&m[641]&~m[642]&~m[643]&~m[677])|(m[640]&~m[641]&m[642]&~m[643]&~m[677])|(~m[640]&m[641]&m[642]&~m[643]&~m[677])|(m[640]&m[641]&m[642]&~m[643]&~m[677])|(m[640]&m[641]&m[642]&m[643]&~m[677])|(m[640]&m[641]&~m[642]&~m[643]&m[677])|(m[640]&~m[641]&m[642]&~m[643]&m[677])|(~m[640]&m[641]&m[642]&~m[643]&m[677])|(m[640]&m[641]&m[642]&~m[643]&m[677])|(m[640]&m[641]&m[642]&m[643]&m[677]))):InitCond[747];
    m[649] = run?((((m[645]&~m[646]&~m[647]&~m[648]&~m[682])|(~m[645]&m[646]&~m[647]&~m[648]&~m[682])|(~m[645]&~m[646]&m[647]&~m[648]&~m[682])|(m[645]&m[646]&~m[647]&m[648]&~m[682])|(m[645]&~m[646]&m[647]&m[648]&~m[682])|(~m[645]&m[646]&m[647]&m[648]&~m[682]))&BiasedRNG[396])|(((m[645]&~m[646]&~m[647]&~m[648]&m[682])|(~m[645]&m[646]&~m[647]&~m[648]&m[682])|(~m[645]&~m[646]&m[647]&~m[648]&m[682])|(m[645]&m[646]&~m[647]&m[648]&m[682])|(m[645]&~m[646]&m[647]&m[648]&m[682])|(~m[645]&m[646]&m[647]&m[648]&m[682]))&~BiasedRNG[396])|((m[645]&m[646]&~m[647]&~m[648]&~m[682])|(m[645]&~m[646]&m[647]&~m[648]&~m[682])|(~m[645]&m[646]&m[647]&~m[648]&~m[682])|(m[645]&m[646]&m[647]&~m[648]&~m[682])|(m[645]&m[646]&m[647]&m[648]&~m[682])|(m[645]&m[646]&~m[647]&~m[648]&m[682])|(m[645]&~m[646]&m[647]&~m[648]&m[682])|(~m[645]&m[646]&m[647]&~m[648]&m[682])|(m[645]&m[646]&m[647]&~m[648]&m[682])|(m[645]&m[646]&m[647]&m[648]&m[682]))):InitCond[748];
    m[654] = run?((((m[650]&~m[651]&~m[652]&~m[653]&~m[687])|(~m[650]&m[651]&~m[652]&~m[653]&~m[687])|(~m[650]&~m[651]&m[652]&~m[653]&~m[687])|(m[650]&m[651]&~m[652]&m[653]&~m[687])|(m[650]&~m[651]&m[652]&m[653]&~m[687])|(~m[650]&m[651]&m[652]&m[653]&~m[687]))&BiasedRNG[397])|(((m[650]&~m[651]&~m[652]&~m[653]&m[687])|(~m[650]&m[651]&~m[652]&~m[653]&m[687])|(~m[650]&~m[651]&m[652]&~m[653]&m[687])|(m[650]&m[651]&~m[652]&m[653]&m[687])|(m[650]&~m[651]&m[652]&m[653]&m[687])|(~m[650]&m[651]&m[652]&m[653]&m[687]))&~BiasedRNG[397])|((m[650]&m[651]&~m[652]&~m[653]&~m[687])|(m[650]&~m[651]&m[652]&~m[653]&~m[687])|(~m[650]&m[651]&m[652]&~m[653]&~m[687])|(m[650]&m[651]&m[652]&~m[653]&~m[687])|(m[650]&m[651]&m[652]&m[653]&~m[687])|(m[650]&m[651]&~m[652]&~m[653]&m[687])|(m[650]&~m[651]&m[652]&~m[653]&m[687])|(~m[650]&m[651]&m[652]&~m[653]&m[687])|(m[650]&m[651]&m[652]&~m[653]&m[687])|(m[650]&m[651]&m[652]&m[653]&m[687]))):InitCond[749];
    m[659] = run?((((m[655]&~m[656]&~m[657]&~m[658]&~m[692])|(~m[655]&m[656]&~m[657]&~m[658]&~m[692])|(~m[655]&~m[656]&m[657]&~m[658]&~m[692])|(m[655]&m[656]&~m[657]&m[658]&~m[692])|(m[655]&~m[656]&m[657]&m[658]&~m[692])|(~m[655]&m[656]&m[657]&m[658]&~m[692]))&BiasedRNG[398])|(((m[655]&~m[656]&~m[657]&~m[658]&m[692])|(~m[655]&m[656]&~m[657]&~m[658]&m[692])|(~m[655]&~m[656]&m[657]&~m[658]&m[692])|(m[655]&m[656]&~m[657]&m[658]&m[692])|(m[655]&~m[656]&m[657]&m[658]&m[692])|(~m[655]&m[656]&m[657]&m[658]&m[692]))&~BiasedRNG[398])|((m[655]&m[656]&~m[657]&~m[658]&~m[692])|(m[655]&~m[656]&m[657]&~m[658]&~m[692])|(~m[655]&m[656]&m[657]&~m[658]&~m[692])|(m[655]&m[656]&m[657]&~m[658]&~m[692])|(m[655]&m[656]&m[657]&m[658]&~m[692])|(m[655]&m[656]&~m[657]&~m[658]&m[692])|(m[655]&~m[656]&m[657]&~m[658]&m[692])|(~m[655]&m[656]&m[657]&~m[658]&m[692])|(m[655]&m[656]&m[657]&~m[658]&m[692])|(m[655]&m[656]&m[657]&m[658]&m[692]))):InitCond[750];
    m[664] = run?((((m[660]&~m[661]&~m[662]&~m[663]&~m[697])|(~m[660]&m[661]&~m[662]&~m[663]&~m[697])|(~m[660]&~m[661]&m[662]&~m[663]&~m[697])|(m[660]&m[661]&~m[662]&m[663]&~m[697])|(m[660]&~m[661]&m[662]&m[663]&~m[697])|(~m[660]&m[661]&m[662]&m[663]&~m[697]))&BiasedRNG[399])|(((m[660]&~m[661]&~m[662]&~m[663]&m[697])|(~m[660]&m[661]&~m[662]&~m[663]&m[697])|(~m[660]&~m[661]&m[662]&~m[663]&m[697])|(m[660]&m[661]&~m[662]&m[663]&m[697])|(m[660]&~m[661]&m[662]&m[663]&m[697])|(~m[660]&m[661]&m[662]&m[663]&m[697]))&~BiasedRNG[399])|((m[660]&m[661]&~m[662]&~m[663]&~m[697])|(m[660]&~m[661]&m[662]&~m[663]&~m[697])|(~m[660]&m[661]&m[662]&~m[663]&~m[697])|(m[660]&m[661]&m[662]&~m[663]&~m[697])|(m[660]&m[661]&m[662]&m[663]&~m[697])|(m[660]&m[661]&~m[662]&~m[663]&m[697])|(m[660]&~m[661]&m[662]&~m[663]&m[697])|(~m[660]&m[661]&m[662]&~m[663]&m[697])|(m[660]&m[661]&m[662]&~m[663]&m[697])|(m[660]&m[661]&m[662]&m[663]&m[697]))):InitCond[751];
    m[669] = run?((((m[665]&~m[666]&~m[667]&~m[668]&~m[702])|(~m[665]&m[666]&~m[667]&~m[668]&~m[702])|(~m[665]&~m[666]&m[667]&~m[668]&~m[702])|(m[665]&m[666]&~m[667]&m[668]&~m[702])|(m[665]&~m[666]&m[667]&m[668]&~m[702])|(~m[665]&m[666]&m[667]&m[668]&~m[702]))&BiasedRNG[400])|(((m[665]&~m[666]&~m[667]&~m[668]&m[702])|(~m[665]&m[666]&~m[667]&~m[668]&m[702])|(~m[665]&~m[666]&m[667]&~m[668]&m[702])|(m[665]&m[666]&~m[667]&m[668]&m[702])|(m[665]&~m[666]&m[667]&m[668]&m[702])|(~m[665]&m[666]&m[667]&m[668]&m[702]))&~BiasedRNG[400])|((m[665]&m[666]&~m[667]&~m[668]&~m[702])|(m[665]&~m[666]&m[667]&~m[668]&~m[702])|(~m[665]&m[666]&m[667]&~m[668]&~m[702])|(m[665]&m[666]&m[667]&~m[668]&~m[702])|(m[665]&m[666]&m[667]&m[668]&~m[702])|(m[665]&m[666]&~m[667]&~m[668]&m[702])|(m[665]&~m[666]&m[667]&~m[668]&m[702])|(~m[665]&m[666]&m[667]&~m[668]&m[702])|(m[665]&m[666]&m[667]&~m[668]&m[702])|(m[665]&m[666]&m[667]&m[668]&m[702]))):InitCond[752];
    m[674] = run?((((m[670]&~m[671]&~m[672]&~m[673]&~m[705])|(~m[670]&m[671]&~m[672]&~m[673]&~m[705])|(~m[670]&~m[671]&m[672]&~m[673]&~m[705])|(m[670]&m[671]&~m[672]&m[673]&~m[705])|(m[670]&~m[671]&m[672]&m[673]&~m[705])|(~m[670]&m[671]&m[672]&m[673]&~m[705]))&BiasedRNG[401])|(((m[670]&~m[671]&~m[672]&~m[673]&m[705])|(~m[670]&m[671]&~m[672]&~m[673]&m[705])|(~m[670]&~m[671]&m[672]&~m[673]&m[705])|(m[670]&m[671]&~m[672]&m[673]&m[705])|(m[670]&~m[671]&m[672]&m[673]&m[705])|(~m[670]&m[671]&m[672]&m[673]&m[705]))&~BiasedRNG[401])|((m[670]&m[671]&~m[672]&~m[673]&~m[705])|(m[670]&~m[671]&m[672]&~m[673]&~m[705])|(~m[670]&m[671]&m[672]&~m[673]&~m[705])|(m[670]&m[671]&m[672]&~m[673]&~m[705])|(m[670]&m[671]&m[672]&m[673]&~m[705])|(m[670]&m[671]&~m[672]&~m[673]&m[705])|(m[670]&~m[671]&m[672]&~m[673]&m[705])|(~m[670]&m[671]&m[672]&~m[673]&m[705])|(m[670]&m[671]&m[672]&~m[673]&m[705])|(m[670]&m[671]&m[672]&m[673]&m[705]))):InitCond[753];
    m[679] = run?((((m[675]&~m[676]&~m[677]&~m[678]&~m[707])|(~m[675]&m[676]&~m[677]&~m[678]&~m[707])|(~m[675]&~m[676]&m[677]&~m[678]&~m[707])|(m[675]&m[676]&~m[677]&m[678]&~m[707])|(m[675]&~m[676]&m[677]&m[678]&~m[707])|(~m[675]&m[676]&m[677]&m[678]&~m[707]))&BiasedRNG[402])|(((m[675]&~m[676]&~m[677]&~m[678]&m[707])|(~m[675]&m[676]&~m[677]&~m[678]&m[707])|(~m[675]&~m[676]&m[677]&~m[678]&m[707])|(m[675]&m[676]&~m[677]&m[678]&m[707])|(m[675]&~m[676]&m[677]&m[678]&m[707])|(~m[675]&m[676]&m[677]&m[678]&m[707]))&~BiasedRNG[402])|((m[675]&m[676]&~m[677]&~m[678]&~m[707])|(m[675]&~m[676]&m[677]&~m[678]&~m[707])|(~m[675]&m[676]&m[677]&~m[678]&~m[707])|(m[675]&m[676]&m[677]&~m[678]&~m[707])|(m[675]&m[676]&m[677]&m[678]&~m[707])|(m[675]&m[676]&~m[677]&~m[678]&m[707])|(m[675]&~m[676]&m[677]&~m[678]&m[707])|(~m[675]&m[676]&m[677]&~m[678]&m[707])|(m[675]&m[676]&m[677]&~m[678]&m[707])|(m[675]&m[676]&m[677]&m[678]&m[707]))):InitCond[754];
    m[684] = run?((((m[680]&~m[681]&~m[682]&~m[683]&~m[712])|(~m[680]&m[681]&~m[682]&~m[683]&~m[712])|(~m[680]&~m[681]&m[682]&~m[683]&~m[712])|(m[680]&m[681]&~m[682]&m[683]&~m[712])|(m[680]&~m[681]&m[682]&m[683]&~m[712])|(~m[680]&m[681]&m[682]&m[683]&~m[712]))&BiasedRNG[403])|(((m[680]&~m[681]&~m[682]&~m[683]&m[712])|(~m[680]&m[681]&~m[682]&~m[683]&m[712])|(~m[680]&~m[681]&m[682]&~m[683]&m[712])|(m[680]&m[681]&~m[682]&m[683]&m[712])|(m[680]&~m[681]&m[682]&m[683]&m[712])|(~m[680]&m[681]&m[682]&m[683]&m[712]))&~BiasedRNG[403])|((m[680]&m[681]&~m[682]&~m[683]&~m[712])|(m[680]&~m[681]&m[682]&~m[683]&~m[712])|(~m[680]&m[681]&m[682]&~m[683]&~m[712])|(m[680]&m[681]&m[682]&~m[683]&~m[712])|(m[680]&m[681]&m[682]&m[683]&~m[712])|(m[680]&m[681]&~m[682]&~m[683]&m[712])|(m[680]&~m[681]&m[682]&~m[683]&m[712])|(~m[680]&m[681]&m[682]&~m[683]&m[712])|(m[680]&m[681]&m[682]&~m[683]&m[712])|(m[680]&m[681]&m[682]&m[683]&m[712]))):InitCond[755];
    m[689] = run?((((m[685]&~m[686]&~m[687]&~m[688]&~m[717])|(~m[685]&m[686]&~m[687]&~m[688]&~m[717])|(~m[685]&~m[686]&m[687]&~m[688]&~m[717])|(m[685]&m[686]&~m[687]&m[688]&~m[717])|(m[685]&~m[686]&m[687]&m[688]&~m[717])|(~m[685]&m[686]&m[687]&m[688]&~m[717]))&BiasedRNG[404])|(((m[685]&~m[686]&~m[687]&~m[688]&m[717])|(~m[685]&m[686]&~m[687]&~m[688]&m[717])|(~m[685]&~m[686]&m[687]&~m[688]&m[717])|(m[685]&m[686]&~m[687]&m[688]&m[717])|(m[685]&~m[686]&m[687]&m[688]&m[717])|(~m[685]&m[686]&m[687]&m[688]&m[717]))&~BiasedRNG[404])|((m[685]&m[686]&~m[687]&~m[688]&~m[717])|(m[685]&~m[686]&m[687]&~m[688]&~m[717])|(~m[685]&m[686]&m[687]&~m[688]&~m[717])|(m[685]&m[686]&m[687]&~m[688]&~m[717])|(m[685]&m[686]&m[687]&m[688]&~m[717])|(m[685]&m[686]&~m[687]&~m[688]&m[717])|(m[685]&~m[686]&m[687]&~m[688]&m[717])|(~m[685]&m[686]&m[687]&~m[688]&m[717])|(m[685]&m[686]&m[687]&~m[688]&m[717])|(m[685]&m[686]&m[687]&m[688]&m[717]))):InitCond[756];
    m[694] = run?((((m[690]&~m[691]&~m[692]&~m[693]&~m[722])|(~m[690]&m[691]&~m[692]&~m[693]&~m[722])|(~m[690]&~m[691]&m[692]&~m[693]&~m[722])|(m[690]&m[691]&~m[692]&m[693]&~m[722])|(m[690]&~m[691]&m[692]&m[693]&~m[722])|(~m[690]&m[691]&m[692]&m[693]&~m[722]))&BiasedRNG[405])|(((m[690]&~m[691]&~m[692]&~m[693]&m[722])|(~m[690]&m[691]&~m[692]&~m[693]&m[722])|(~m[690]&~m[691]&m[692]&~m[693]&m[722])|(m[690]&m[691]&~m[692]&m[693]&m[722])|(m[690]&~m[691]&m[692]&m[693]&m[722])|(~m[690]&m[691]&m[692]&m[693]&m[722]))&~BiasedRNG[405])|((m[690]&m[691]&~m[692]&~m[693]&~m[722])|(m[690]&~m[691]&m[692]&~m[693]&~m[722])|(~m[690]&m[691]&m[692]&~m[693]&~m[722])|(m[690]&m[691]&m[692]&~m[693]&~m[722])|(m[690]&m[691]&m[692]&m[693]&~m[722])|(m[690]&m[691]&~m[692]&~m[693]&m[722])|(m[690]&~m[691]&m[692]&~m[693]&m[722])|(~m[690]&m[691]&m[692]&~m[693]&m[722])|(m[690]&m[691]&m[692]&~m[693]&m[722])|(m[690]&m[691]&m[692]&m[693]&m[722]))):InitCond[757];
    m[699] = run?((((m[695]&~m[696]&~m[697]&~m[698]&~m[727])|(~m[695]&m[696]&~m[697]&~m[698]&~m[727])|(~m[695]&~m[696]&m[697]&~m[698]&~m[727])|(m[695]&m[696]&~m[697]&m[698]&~m[727])|(m[695]&~m[696]&m[697]&m[698]&~m[727])|(~m[695]&m[696]&m[697]&m[698]&~m[727]))&BiasedRNG[406])|(((m[695]&~m[696]&~m[697]&~m[698]&m[727])|(~m[695]&m[696]&~m[697]&~m[698]&m[727])|(~m[695]&~m[696]&m[697]&~m[698]&m[727])|(m[695]&m[696]&~m[697]&m[698]&m[727])|(m[695]&~m[696]&m[697]&m[698]&m[727])|(~m[695]&m[696]&m[697]&m[698]&m[727]))&~BiasedRNG[406])|((m[695]&m[696]&~m[697]&~m[698]&~m[727])|(m[695]&~m[696]&m[697]&~m[698]&~m[727])|(~m[695]&m[696]&m[697]&~m[698]&~m[727])|(m[695]&m[696]&m[697]&~m[698]&~m[727])|(m[695]&m[696]&m[697]&m[698]&~m[727])|(m[695]&m[696]&~m[697]&~m[698]&m[727])|(m[695]&~m[696]&m[697]&~m[698]&m[727])|(~m[695]&m[696]&m[697]&~m[698]&m[727])|(m[695]&m[696]&m[697]&~m[698]&m[727])|(m[695]&m[696]&m[697]&m[698]&m[727]))):InitCond[758];
    m[704] = run?((((m[700]&~m[701]&~m[702]&~m[703]&~m[732])|(~m[700]&m[701]&~m[702]&~m[703]&~m[732])|(~m[700]&~m[701]&m[702]&~m[703]&~m[732])|(m[700]&m[701]&~m[702]&m[703]&~m[732])|(m[700]&~m[701]&m[702]&m[703]&~m[732])|(~m[700]&m[701]&m[702]&m[703]&~m[732]))&BiasedRNG[407])|(((m[700]&~m[701]&~m[702]&~m[703]&m[732])|(~m[700]&m[701]&~m[702]&~m[703]&m[732])|(~m[700]&~m[701]&m[702]&~m[703]&m[732])|(m[700]&m[701]&~m[702]&m[703]&m[732])|(m[700]&~m[701]&m[702]&m[703]&m[732])|(~m[700]&m[701]&m[702]&m[703]&m[732]))&~BiasedRNG[407])|((m[700]&m[701]&~m[702]&~m[703]&~m[732])|(m[700]&~m[701]&m[702]&~m[703]&~m[732])|(~m[700]&m[701]&m[702]&~m[703]&~m[732])|(m[700]&m[701]&m[702]&~m[703]&~m[732])|(m[700]&m[701]&m[702]&m[703]&~m[732])|(m[700]&m[701]&~m[702]&~m[703]&m[732])|(m[700]&~m[701]&m[702]&~m[703]&m[732])|(~m[700]&m[701]&m[702]&~m[703]&m[732])|(m[700]&m[701]&m[702]&~m[703]&m[732])|(m[700]&m[701]&m[702]&m[703]&m[732]))):InitCond[759];
    m[709] = run?((((m[705]&~m[706]&~m[707]&~m[708]&~m[735])|(~m[705]&m[706]&~m[707]&~m[708]&~m[735])|(~m[705]&~m[706]&m[707]&~m[708]&~m[735])|(m[705]&m[706]&~m[707]&m[708]&~m[735])|(m[705]&~m[706]&m[707]&m[708]&~m[735])|(~m[705]&m[706]&m[707]&m[708]&~m[735]))&BiasedRNG[408])|(((m[705]&~m[706]&~m[707]&~m[708]&m[735])|(~m[705]&m[706]&~m[707]&~m[708]&m[735])|(~m[705]&~m[706]&m[707]&~m[708]&m[735])|(m[705]&m[706]&~m[707]&m[708]&m[735])|(m[705]&~m[706]&m[707]&m[708]&m[735])|(~m[705]&m[706]&m[707]&m[708]&m[735]))&~BiasedRNG[408])|((m[705]&m[706]&~m[707]&~m[708]&~m[735])|(m[705]&~m[706]&m[707]&~m[708]&~m[735])|(~m[705]&m[706]&m[707]&~m[708]&~m[735])|(m[705]&m[706]&m[707]&~m[708]&~m[735])|(m[705]&m[706]&m[707]&m[708]&~m[735])|(m[705]&m[706]&~m[707]&~m[708]&m[735])|(m[705]&~m[706]&m[707]&~m[708]&m[735])|(~m[705]&m[706]&m[707]&~m[708]&m[735])|(m[705]&m[706]&m[707]&~m[708]&m[735])|(m[705]&m[706]&m[707]&m[708]&m[735]))):InitCond[760];
    m[714] = run?((((m[710]&~m[711]&~m[712]&~m[713]&~m[737])|(~m[710]&m[711]&~m[712]&~m[713]&~m[737])|(~m[710]&~m[711]&m[712]&~m[713]&~m[737])|(m[710]&m[711]&~m[712]&m[713]&~m[737])|(m[710]&~m[711]&m[712]&m[713]&~m[737])|(~m[710]&m[711]&m[712]&m[713]&~m[737]))&BiasedRNG[409])|(((m[710]&~m[711]&~m[712]&~m[713]&m[737])|(~m[710]&m[711]&~m[712]&~m[713]&m[737])|(~m[710]&~m[711]&m[712]&~m[713]&m[737])|(m[710]&m[711]&~m[712]&m[713]&m[737])|(m[710]&~m[711]&m[712]&m[713]&m[737])|(~m[710]&m[711]&m[712]&m[713]&m[737]))&~BiasedRNG[409])|((m[710]&m[711]&~m[712]&~m[713]&~m[737])|(m[710]&~m[711]&m[712]&~m[713]&~m[737])|(~m[710]&m[711]&m[712]&~m[713]&~m[737])|(m[710]&m[711]&m[712]&~m[713]&~m[737])|(m[710]&m[711]&m[712]&m[713]&~m[737])|(m[710]&m[711]&~m[712]&~m[713]&m[737])|(m[710]&~m[711]&m[712]&~m[713]&m[737])|(~m[710]&m[711]&m[712]&~m[713]&m[737])|(m[710]&m[711]&m[712]&~m[713]&m[737])|(m[710]&m[711]&m[712]&m[713]&m[737]))):InitCond[761];
    m[719] = run?((((m[715]&~m[716]&~m[717]&~m[718]&~m[742])|(~m[715]&m[716]&~m[717]&~m[718]&~m[742])|(~m[715]&~m[716]&m[717]&~m[718]&~m[742])|(m[715]&m[716]&~m[717]&m[718]&~m[742])|(m[715]&~m[716]&m[717]&m[718]&~m[742])|(~m[715]&m[716]&m[717]&m[718]&~m[742]))&BiasedRNG[410])|(((m[715]&~m[716]&~m[717]&~m[718]&m[742])|(~m[715]&m[716]&~m[717]&~m[718]&m[742])|(~m[715]&~m[716]&m[717]&~m[718]&m[742])|(m[715]&m[716]&~m[717]&m[718]&m[742])|(m[715]&~m[716]&m[717]&m[718]&m[742])|(~m[715]&m[716]&m[717]&m[718]&m[742]))&~BiasedRNG[410])|((m[715]&m[716]&~m[717]&~m[718]&~m[742])|(m[715]&~m[716]&m[717]&~m[718]&~m[742])|(~m[715]&m[716]&m[717]&~m[718]&~m[742])|(m[715]&m[716]&m[717]&~m[718]&~m[742])|(m[715]&m[716]&m[717]&m[718]&~m[742])|(m[715]&m[716]&~m[717]&~m[718]&m[742])|(m[715]&~m[716]&m[717]&~m[718]&m[742])|(~m[715]&m[716]&m[717]&~m[718]&m[742])|(m[715]&m[716]&m[717]&~m[718]&m[742])|(m[715]&m[716]&m[717]&m[718]&m[742]))):InitCond[762];
    m[724] = run?((((m[720]&~m[721]&~m[722]&~m[723]&~m[747])|(~m[720]&m[721]&~m[722]&~m[723]&~m[747])|(~m[720]&~m[721]&m[722]&~m[723]&~m[747])|(m[720]&m[721]&~m[722]&m[723]&~m[747])|(m[720]&~m[721]&m[722]&m[723]&~m[747])|(~m[720]&m[721]&m[722]&m[723]&~m[747]))&BiasedRNG[411])|(((m[720]&~m[721]&~m[722]&~m[723]&m[747])|(~m[720]&m[721]&~m[722]&~m[723]&m[747])|(~m[720]&~m[721]&m[722]&~m[723]&m[747])|(m[720]&m[721]&~m[722]&m[723]&m[747])|(m[720]&~m[721]&m[722]&m[723]&m[747])|(~m[720]&m[721]&m[722]&m[723]&m[747]))&~BiasedRNG[411])|((m[720]&m[721]&~m[722]&~m[723]&~m[747])|(m[720]&~m[721]&m[722]&~m[723]&~m[747])|(~m[720]&m[721]&m[722]&~m[723]&~m[747])|(m[720]&m[721]&m[722]&~m[723]&~m[747])|(m[720]&m[721]&m[722]&m[723]&~m[747])|(m[720]&m[721]&~m[722]&~m[723]&m[747])|(m[720]&~m[721]&m[722]&~m[723]&m[747])|(~m[720]&m[721]&m[722]&~m[723]&m[747])|(m[720]&m[721]&m[722]&~m[723]&m[747])|(m[720]&m[721]&m[722]&m[723]&m[747]))):InitCond[763];
    m[729] = run?((((m[725]&~m[726]&~m[727]&~m[728]&~m[752])|(~m[725]&m[726]&~m[727]&~m[728]&~m[752])|(~m[725]&~m[726]&m[727]&~m[728]&~m[752])|(m[725]&m[726]&~m[727]&m[728]&~m[752])|(m[725]&~m[726]&m[727]&m[728]&~m[752])|(~m[725]&m[726]&m[727]&m[728]&~m[752]))&BiasedRNG[412])|(((m[725]&~m[726]&~m[727]&~m[728]&m[752])|(~m[725]&m[726]&~m[727]&~m[728]&m[752])|(~m[725]&~m[726]&m[727]&~m[728]&m[752])|(m[725]&m[726]&~m[727]&m[728]&m[752])|(m[725]&~m[726]&m[727]&m[728]&m[752])|(~m[725]&m[726]&m[727]&m[728]&m[752]))&~BiasedRNG[412])|((m[725]&m[726]&~m[727]&~m[728]&~m[752])|(m[725]&~m[726]&m[727]&~m[728]&~m[752])|(~m[725]&m[726]&m[727]&~m[728]&~m[752])|(m[725]&m[726]&m[727]&~m[728]&~m[752])|(m[725]&m[726]&m[727]&m[728]&~m[752])|(m[725]&m[726]&~m[727]&~m[728]&m[752])|(m[725]&~m[726]&m[727]&~m[728]&m[752])|(~m[725]&m[726]&m[727]&~m[728]&m[752])|(m[725]&m[726]&m[727]&~m[728]&m[752])|(m[725]&m[726]&m[727]&m[728]&m[752]))):InitCond[764];
    m[734] = run?((((m[730]&~m[731]&~m[732]&~m[733]&~m[757])|(~m[730]&m[731]&~m[732]&~m[733]&~m[757])|(~m[730]&~m[731]&m[732]&~m[733]&~m[757])|(m[730]&m[731]&~m[732]&m[733]&~m[757])|(m[730]&~m[731]&m[732]&m[733]&~m[757])|(~m[730]&m[731]&m[732]&m[733]&~m[757]))&BiasedRNG[413])|(((m[730]&~m[731]&~m[732]&~m[733]&m[757])|(~m[730]&m[731]&~m[732]&~m[733]&m[757])|(~m[730]&~m[731]&m[732]&~m[733]&m[757])|(m[730]&m[731]&~m[732]&m[733]&m[757])|(m[730]&~m[731]&m[732]&m[733]&m[757])|(~m[730]&m[731]&m[732]&m[733]&m[757]))&~BiasedRNG[413])|((m[730]&m[731]&~m[732]&~m[733]&~m[757])|(m[730]&~m[731]&m[732]&~m[733]&~m[757])|(~m[730]&m[731]&m[732]&~m[733]&~m[757])|(m[730]&m[731]&m[732]&~m[733]&~m[757])|(m[730]&m[731]&m[732]&m[733]&~m[757])|(m[730]&m[731]&~m[732]&~m[733]&m[757])|(m[730]&~m[731]&m[732]&~m[733]&m[757])|(~m[730]&m[731]&m[732]&~m[733]&m[757])|(m[730]&m[731]&m[732]&~m[733]&m[757])|(m[730]&m[731]&m[732]&m[733]&m[757]))):InitCond[765];
    m[739] = run?((((m[735]&~m[736]&~m[737]&~m[738]&~m[760])|(~m[735]&m[736]&~m[737]&~m[738]&~m[760])|(~m[735]&~m[736]&m[737]&~m[738]&~m[760])|(m[735]&m[736]&~m[737]&m[738]&~m[760])|(m[735]&~m[736]&m[737]&m[738]&~m[760])|(~m[735]&m[736]&m[737]&m[738]&~m[760]))&BiasedRNG[414])|(((m[735]&~m[736]&~m[737]&~m[738]&m[760])|(~m[735]&m[736]&~m[737]&~m[738]&m[760])|(~m[735]&~m[736]&m[737]&~m[738]&m[760])|(m[735]&m[736]&~m[737]&m[738]&m[760])|(m[735]&~m[736]&m[737]&m[738]&m[760])|(~m[735]&m[736]&m[737]&m[738]&m[760]))&~BiasedRNG[414])|((m[735]&m[736]&~m[737]&~m[738]&~m[760])|(m[735]&~m[736]&m[737]&~m[738]&~m[760])|(~m[735]&m[736]&m[737]&~m[738]&~m[760])|(m[735]&m[736]&m[737]&~m[738]&~m[760])|(m[735]&m[736]&m[737]&m[738]&~m[760])|(m[735]&m[736]&~m[737]&~m[738]&m[760])|(m[735]&~m[736]&m[737]&~m[738]&m[760])|(~m[735]&m[736]&m[737]&~m[738]&m[760])|(m[735]&m[736]&m[737]&~m[738]&m[760])|(m[735]&m[736]&m[737]&m[738]&m[760]))):InitCond[766];
    m[744] = run?((((m[740]&~m[741]&~m[742]&~m[743]&~m[762])|(~m[740]&m[741]&~m[742]&~m[743]&~m[762])|(~m[740]&~m[741]&m[742]&~m[743]&~m[762])|(m[740]&m[741]&~m[742]&m[743]&~m[762])|(m[740]&~m[741]&m[742]&m[743]&~m[762])|(~m[740]&m[741]&m[742]&m[743]&~m[762]))&BiasedRNG[415])|(((m[740]&~m[741]&~m[742]&~m[743]&m[762])|(~m[740]&m[741]&~m[742]&~m[743]&m[762])|(~m[740]&~m[741]&m[742]&~m[743]&m[762])|(m[740]&m[741]&~m[742]&m[743]&m[762])|(m[740]&~m[741]&m[742]&m[743]&m[762])|(~m[740]&m[741]&m[742]&m[743]&m[762]))&~BiasedRNG[415])|((m[740]&m[741]&~m[742]&~m[743]&~m[762])|(m[740]&~m[741]&m[742]&~m[743]&~m[762])|(~m[740]&m[741]&m[742]&~m[743]&~m[762])|(m[740]&m[741]&m[742]&~m[743]&~m[762])|(m[740]&m[741]&m[742]&m[743]&~m[762])|(m[740]&m[741]&~m[742]&~m[743]&m[762])|(m[740]&~m[741]&m[742]&~m[743]&m[762])|(~m[740]&m[741]&m[742]&~m[743]&m[762])|(m[740]&m[741]&m[742]&~m[743]&m[762])|(m[740]&m[741]&m[742]&m[743]&m[762]))):InitCond[767];
    m[749] = run?((((m[745]&~m[746]&~m[747]&~m[748]&~m[767])|(~m[745]&m[746]&~m[747]&~m[748]&~m[767])|(~m[745]&~m[746]&m[747]&~m[748]&~m[767])|(m[745]&m[746]&~m[747]&m[748]&~m[767])|(m[745]&~m[746]&m[747]&m[748]&~m[767])|(~m[745]&m[746]&m[747]&m[748]&~m[767]))&BiasedRNG[416])|(((m[745]&~m[746]&~m[747]&~m[748]&m[767])|(~m[745]&m[746]&~m[747]&~m[748]&m[767])|(~m[745]&~m[746]&m[747]&~m[748]&m[767])|(m[745]&m[746]&~m[747]&m[748]&m[767])|(m[745]&~m[746]&m[747]&m[748]&m[767])|(~m[745]&m[746]&m[747]&m[748]&m[767]))&~BiasedRNG[416])|((m[745]&m[746]&~m[747]&~m[748]&~m[767])|(m[745]&~m[746]&m[747]&~m[748]&~m[767])|(~m[745]&m[746]&m[747]&~m[748]&~m[767])|(m[745]&m[746]&m[747]&~m[748]&~m[767])|(m[745]&m[746]&m[747]&m[748]&~m[767])|(m[745]&m[746]&~m[747]&~m[748]&m[767])|(m[745]&~m[746]&m[747]&~m[748]&m[767])|(~m[745]&m[746]&m[747]&~m[748]&m[767])|(m[745]&m[746]&m[747]&~m[748]&m[767])|(m[745]&m[746]&m[747]&m[748]&m[767]))):InitCond[768];
    m[754] = run?((((m[750]&~m[751]&~m[752]&~m[753]&~m[772])|(~m[750]&m[751]&~m[752]&~m[753]&~m[772])|(~m[750]&~m[751]&m[752]&~m[753]&~m[772])|(m[750]&m[751]&~m[752]&m[753]&~m[772])|(m[750]&~m[751]&m[752]&m[753]&~m[772])|(~m[750]&m[751]&m[752]&m[753]&~m[772]))&BiasedRNG[417])|(((m[750]&~m[751]&~m[752]&~m[753]&m[772])|(~m[750]&m[751]&~m[752]&~m[753]&m[772])|(~m[750]&~m[751]&m[752]&~m[753]&m[772])|(m[750]&m[751]&~m[752]&m[753]&m[772])|(m[750]&~m[751]&m[752]&m[753]&m[772])|(~m[750]&m[751]&m[752]&m[753]&m[772]))&~BiasedRNG[417])|((m[750]&m[751]&~m[752]&~m[753]&~m[772])|(m[750]&~m[751]&m[752]&~m[753]&~m[772])|(~m[750]&m[751]&m[752]&~m[753]&~m[772])|(m[750]&m[751]&m[752]&~m[753]&~m[772])|(m[750]&m[751]&m[752]&m[753]&~m[772])|(m[750]&m[751]&~m[752]&~m[753]&m[772])|(m[750]&~m[751]&m[752]&~m[753]&m[772])|(~m[750]&m[751]&m[752]&~m[753]&m[772])|(m[750]&m[751]&m[752]&~m[753]&m[772])|(m[750]&m[751]&m[752]&m[753]&m[772]))):InitCond[769];
    m[759] = run?((((m[755]&~m[756]&~m[757]&~m[758]&~m[777])|(~m[755]&m[756]&~m[757]&~m[758]&~m[777])|(~m[755]&~m[756]&m[757]&~m[758]&~m[777])|(m[755]&m[756]&~m[757]&m[758]&~m[777])|(m[755]&~m[756]&m[757]&m[758]&~m[777])|(~m[755]&m[756]&m[757]&m[758]&~m[777]))&BiasedRNG[418])|(((m[755]&~m[756]&~m[757]&~m[758]&m[777])|(~m[755]&m[756]&~m[757]&~m[758]&m[777])|(~m[755]&~m[756]&m[757]&~m[758]&m[777])|(m[755]&m[756]&~m[757]&m[758]&m[777])|(m[755]&~m[756]&m[757]&m[758]&m[777])|(~m[755]&m[756]&m[757]&m[758]&m[777]))&~BiasedRNG[418])|((m[755]&m[756]&~m[757]&~m[758]&~m[777])|(m[755]&~m[756]&m[757]&~m[758]&~m[777])|(~m[755]&m[756]&m[757]&~m[758]&~m[777])|(m[755]&m[756]&m[757]&~m[758]&~m[777])|(m[755]&m[756]&m[757]&m[758]&~m[777])|(m[755]&m[756]&~m[757]&~m[758]&m[777])|(m[755]&~m[756]&m[757]&~m[758]&m[777])|(~m[755]&m[756]&m[757]&~m[758]&m[777])|(m[755]&m[756]&m[757]&~m[758]&m[777])|(m[755]&m[756]&m[757]&m[758]&m[777]))):InitCond[770];
    m[764] = run?((((m[760]&~m[761]&~m[762]&~m[763]&~m[780])|(~m[760]&m[761]&~m[762]&~m[763]&~m[780])|(~m[760]&~m[761]&m[762]&~m[763]&~m[780])|(m[760]&m[761]&~m[762]&m[763]&~m[780])|(m[760]&~m[761]&m[762]&m[763]&~m[780])|(~m[760]&m[761]&m[762]&m[763]&~m[780]))&BiasedRNG[419])|(((m[760]&~m[761]&~m[762]&~m[763]&m[780])|(~m[760]&m[761]&~m[762]&~m[763]&m[780])|(~m[760]&~m[761]&m[762]&~m[763]&m[780])|(m[760]&m[761]&~m[762]&m[763]&m[780])|(m[760]&~m[761]&m[762]&m[763]&m[780])|(~m[760]&m[761]&m[762]&m[763]&m[780]))&~BiasedRNG[419])|((m[760]&m[761]&~m[762]&~m[763]&~m[780])|(m[760]&~m[761]&m[762]&~m[763]&~m[780])|(~m[760]&m[761]&m[762]&~m[763]&~m[780])|(m[760]&m[761]&m[762]&~m[763]&~m[780])|(m[760]&m[761]&m[762]&m[763]&~m[780])|(m[760]&m[761]&~m[762]&~m[763]&m[780])|(m[760]&~m[761]&m[762]&~m[763]&m[780])|(~m[760]&m[761]&m[762]&~m[763]&m[780])|(m[760]&m[761]&m[762]&~m[763]&m[780])|(m[760]&m[761]&m[762]&m[763]&m[780]))):InitCond[771];
    m[769] = run?((((m[765]&~m[766]&~m[767]&~m[768]&~m[782])|(~m[765]&m[766]&~m[767]&~m[768]&~m[782])|(~m[765]&~m[766]&m[767]&~m[768]&~m[782])|(m[765]&m[766]&~m[767]&m[768]&~m[782])|(m[765]&~m[766]&m[767]&m[768]&~m[782])|(~m[765]&m[766]&m[767]&m[768]&~m[782]))&BiasedRNG[420])|(((m[765]&~m[766]&~m[767]&~m[768]&m[782])|(~m[765]&m[766]&~m[767]&~m[768]&m[782])|(~m[765]&~m[766]&m[767]&~m[768]&m[782])|(m[765]&m[766]&~m[767]&m[768]&m[782])|(m[765]&~m[766]&m[767]&m[768]&m[782])|(~m[765]&m[766]&m[767]&m[768]&m[782]))&~BiasedRNG[420])|((m[765]&m[766]&~m[767]&~m[768]&~m[782])|(m[765]&~m[766]&m[767]&~m[768]&~m[782])|(~m[765]&m[766]&m[767]&~m[768]&~m[782])|(m[765]&m[766]&m[767]&~m[768]&~m[782])|(m[765]&m[766]&m[767]&m[768]&~m[782])|(m[765]&m[766]&~m[767]&~m[768]&m[782])|(m[765]&~m[766]&m[767]&~m[768]&m[782])|(~m[765]&m[766]&m[767]&~m[768]&m[782])|(m[765]&m[766]&m[767]&~m[768]&m[782])|(m[765]&m[766]&m[767]&m[768]&m[782]))):InitCond[772];
    m[774] = run?((((m[770]&~m[771]&~m[772]&~m[773]&~m[787])|(~m[770]&m[771]&~m[772]&~m[773]&~m[787])|(~m[770]&~m[771]&m[772]&~m[773]&~m[787])|(m[770]&m[771]&~m[772]&m[773]&~m[787])|(m[770]&~m[771]&m[772]&m[773]&~m[787])|(~m[770]&m[771]&m[772]&m[773]&~m[787]))&BiasedRNG[421])|(((m[770]&~m[771]&~m[772]&~m[773]&m[787])|(~m[770]&m[771]&~m[772]&~m[773]&m[787])|(~m[770]&~m[771]&m[772]&~m[773]&m[787])|(m[770]&m[771]&~m[772]&m[773]&m[787])|(m[770]&~m[771]&m[772]&m[773]&m[787])|(~m[770]&m[771]&m[772]&m[773]&m[787]))&~BiasedRNG[421])|((m[770]&m[771]&~m[772]&~m[773]&~m[787])|(m[770]&~m[771]&m[772]&~m[773]&~m[787])|(~m[770]&m[771]&m[772]&~m[773]&~m[787])|(m[770]&m[771]&m[772]&~m[773]&~m[787])|(m[770]&m[771]&m[772]&m[773]&~m[787])|(m[770]&m[771]&~m[772]&~m[773]&m[787])|(m[770]&~m[771]&m[772]&~m[773]&m[787])|(~m[770]&m[771]&m[772]&~m[773]&m[787])|(m[770]&m[771]&m[772]&~m[773]&m[787])|(m[770]&m[771]&m[772]&m[773]&m[787]))):InitCond[773];
    m[779] = run?((((m[775]&~m[776]&~m[777]&~m[778]&~m[792])|(~m[775]&m[776]&~m[777]&~m[778]&~m[792])|(~m[775]&~m[776]&m[777]&~m[778]&~m[792])|(m[775]&m[776]&~m[777]&m[778]&~m[792])|(m[775]&~m[776]&m[777]&m[778]&~m[792])|(~m[775]&m[776]&m[777]&m[778]&~m[792]))&BiasedRNG[422])|(((m[775]&~m[776]&~m[777]&~m[778]&m[792])|(~m[775]&m[776]&~m[777]&~m[778]&m[792])|(~m[775]&~m[776]&m[777]&~m[778]&m[792])|(m[775]&m[776]&~m[777]&m[778]&m[792])|(m[775]&~m[776]&m[777]&m[778]&m[792])|(~m[775]&m[776]&m[777]&m[778]&m[792]))&~BiasedRNG[422])|((m[775]&m[776]&~m[777]&~m[778]&~m[792])|(m[775]&~m[776]&m[777]&~m[778]&~m[792])|(~m[775]&m[776]&m[777]&~m[778]&~m[792])|(m[775]&m[776]&m[777]&~m[778]&~m[792])|(m[775]&m[776]&m[777]&m[778]&~m[792])|(m[775]&m[776]&~m[777]&~m[778]&m[792])|(m[775]&~m[776]&m[777]&~m[778]&m[792])|(~m[775]&m[776]&m[777]&~m[778]&m[792])|(m[775]&m[776]&m[777]&~m[778]&m[792])|(m[775]&m[776]&m[777]&m[778]&m[792]))):InitCond[774];
    m[784] = run?((((m[780]&~m[781]&~m[782]&~m[783]&~m[795])|(~m[780]&m[781]&~m[782]&~m[783]&~m[795])|(~m[780]&~m[781]&m[782]&~m[783]&~m[795])|(m[780]&m[781]&~m[782]&m[783]&~m[795])|(m[780]&~m[781]&m[782]&m[783]&~m[795])|(~m[780]&m[781]&m[782]&m[783]&~m[795]))&BiasedRNG[423])|(((m[780]&~m[781]&~m[782]&~m[783]&m[795])|(~m[780]&m[781]&~m[782]&~m[783]&m[795])|(~m[780]&~m[781]&m[782]&~m[783]&m[795])|(m[780]&m[781]&~m[782]&m[783]&m[795])|(m[780]&~m[781]&m[782]&m[783]&m[795])|(~m[780]&m[781]&m[782]&m[783]&m[795]))&~BiasedRNG[423])|((m[780]&m[781]&~m[782]&~m[783]&~m[795])|(m[780]&~m[781]&m[782]&~m[783]&~m[795])|(~m[780]&m[781]&m[782]&~m[783]&~m[795])|(m[780]&m[781]&m[782]&~m[783]&~m[795])|(m[780]&m[781]&m[782]&m[783]&~m[795])|(m[780]&m[781]&~m[782]&~m[783]&m[795])|(m[780]&~m[781]&m[782]&~m[783]&m[795])|(~m[780]&m[781]&m[782]&~m[783]&m[795])|(m[780]&m[781]&m[782]&~m[783]&m[795])|(m[780]&m[781]&m[782]&m[783]&m[795]))):InitCond[775];
    m[789] = run?((((m[785]&~m[786]&~m[787]&~m[788]&~m[797])|(~m[785]&m[786]&~m[787]&~m[788]&~m[797])|(~m[785]&~m[786]&m[787]&~m[788]&~m[797])|(m[785]&m[786]&~m[787]&m[788]&~m[797])|(m[785]&~m[786]&m[787]&m[788]&~m[797])|(~m[785]&m[786]&m[787]&m[788]&~m[797]))&BiasedRNG[424])|(((m[785]&~m[786]&~m[787]&~m[788]&m[797])|(~m[785]&m[786]&~m[787]&~m[788]&m[797])|(~m[785]&~m[786]&m[787]&~m[788]&m[797])|(m[785]&m[786]&~m[787]&m[788]&m[797])|(m[785]&~m[786]&m[787]&m[788]&m[797])|(~m[785]&m[786]&m[787]&m[788]&m[797]))&~BiasedRNG[424])|((m[785]&m[786]&~m[787]&~m[788]&~m[797])|(m[785]&~m[786]&m[787]&~m[788]&~m[797])|(~m[785]&m[786]&m[787]&~m[788]&~m[797])|(m[785]&m[786]&m[787]&~m[788]&~m[797])|(m[785]&m[786]&m[787]&m[788]&~m[797])|(m[785]&m[786]&~m[787]&~m[788]&m[797])|(m[785]&~m[786]&m[787]&~m[788]&m[797])|(~m[785]&m[786]&m[787]&~m[788]&m[797])|(m[785]&m[786]&m[787]&~m[788]&m[797])|(m[785]&m[786]&m[787]&m[788]&m[797]))):InitCond[776];
    m[794] = run?((((m[790]&~m[791]&~m[792]&~m[793]&~m[802])|(~m[790]&m[791]&~m[792]&~m[793]&~m[802])|(~m[790]&~m[791]&m[792]&~m[793]&~m[802])|(m[790]&m[791]&~m[792]&m[793]&~m[802])|(m[790]&~m[791]&m[792]&m[793]&~m[802])|(~m[790]&m[791]&m[792]&m[793]&~m[802]))&BiasedRNG[425])|(((m[790]&~m[791]&~m[792]&~m[793]&m[802])|(~m[790]&m[791]&~m[792]&~m[793]&m[802])|(~m[790]&~m[791]&m[792]&~m[793]&m[802])|(m[790]&m[791]&~m[792]&m[793]&m[802])|(m[790]&~m[791]&m[792]&m[793]&m[802])|(~m[790]&m[791]&m[792]&m[793]&m[802]))&~BiasedRNG[425])|((m[790]&m[791]&~m[792]&~m[793]&~m[802])|(m[790]&~m[791]&m[792]&~m[793]&~m[802])|(~m[790]&m[791]&m[792]&~m[793]&~m[802])|(m[790]&m[791]&m[792]&~m[793]&~m[802])|(m[790]&m[791]&m[792]&m[793]&~m[802])|(m[790]&m[791]&~m[792]&~m[793]&m[802])|(m[790]&~m[791]&m[792]&~m[793]&m[802])|(~m[790]&m[791]&m[792]&~m[793]&m[802])|(m[790]&m[791]&m[792]&~m[793]&m[802])|(m[790]&m[791]&m[792]&m[793]&m[802]))):InitCond[777];
    m[799] = run?((((m[795]&~m[796]&~m[797]&~m[798]&~m[805])|(~m[795]&m[796]&~m[797]&~m[798]&~m[805])|(~m[795]&~m[796]&m[797]&~m[798]&~m[805])|(m[795]&m[796]&~m[797]&m[798]&~m[805])|(m[795]&~m[796]&m[797]&m[798]&~m[805])|(~m[795]&m[796]&m[797]&m[798]&~m[805]))&BiasedRNG[426])|(((m[795]&~m[796]&~m[797]&~m[798]&m[805])|(~m[795]&m[796]&~m[797]&~m[798]&m[805])|(~m[795]&~m[796]&m[797]&~m[798]&m[805])|(m[795]&m[796]&~m[797]&m[798]&m[805])|(m[795]&~m[796]&m[797]&m[798]&m[805])|(~m[795]&m[796]&m[797]&m[798]&m[805]))&~BiasedRNG[426])|((m[795]&m[796]&~m[797]&~m[798]&~m[805])|(m[795]&~m[796]&m[797]&~m[798]&~m[805])|(~m[795]&m[796]&m[797]&~m[798]&~m[805])|(m[795]&m[796]&m[797]&~m[798]&~m[805])|(m[795]&m[796]&m[797]&m[798]&~m[805])|(m[795]&m[796]&~m[797]&~m[798]&m[805])|(m[795]&~m[796]&m[797]&~m[798]&m[805])|(~m[795]&m[796]&m[797]&~m[798]&m[805])|(m[795]&m[796]&m[797]&~m[798]&m[805])|(m[795]&m[796]&m[797]&m[798]&m[805]))):InitCond[778];
    m[804] = run?((((m[800]&~m[801]&~m[802]&~m[803]&~m[807])|(~m[800]&m[801]&~m[802]&~m[803]&~m[807])|(~m[800]&~m[801]&m[802]&~m[803]&~m[807])|(m[800]&m[801]&~m[802]&m[803]&~m[807])|(m[800]&~m[801]&m[802]&m[803]&~m[807])|(~m[800]&m[801]&m[802]&m[803]&~m[807]))&BiasedRNG[427])|(((m[800]&~m[801]&~m[802]&~m[803]&m[807])|(~m[800]&m[801]&~m[802]&~m[803]&m[807])|(~m[800]&~m[801]&m[802]&~m[803]&m[807])|(m[800]&m[801]&~m[802]&m[803]&m[807])|(m[800]&~m[801]&m[802]&m[803]&m[807])|(~m[800]&m[801]&m[802]&m[803]&m[807]))&~BiasedRNG[427])|((m[800]&m[801]&~m[802]&~m[803]&~m[807])|(m[800]&~m[801]&m[802]&~m[803]&~m[807])|(~m[800]&m[801]&m[802]&~m[803]&~m[807])|(m[800]&m[801]&m[802]&~m[803]&~m[807])|(m[800]&m[801]&m[802]&m[803]&~m[807])|(m[800]&m[801]&~m[802]&~m[803]&m[807])|(m[800]&~m[801]&m[802]&~m[803]&m[807])|(~m[800]&m[801]&m[802]&~m[803]&m[807])|(m[800]&m[801]&m[802]&~m[803]&m[807])|(m[800]&m[801]&m[802]&m[803]&m[807]))):InitCond[779];
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[159]&LFSRcolor0[54]&LFSRcolor0[378]);
    BiasedRNG[1] = (LFSRcolor0[208]&LFSRcolor0[340]&LFSRcolor0[403]);
    BiasedRNG[2] = (LFSRcolor0[350]&LFSRcolor0[274]&LFSRcolor0[71]);
    BiasedRNG[3] = (LFSRcolor0[371]&LFSRcolor0[74]&LFSRcolor0[36]);
    BiasedRNG[4] = (LFSRcolor0[389]&LFSRcolor0[413]&LFSRcolor0[409]);
    BiasedRNG[5] = (LFSRcolor0[211]&LFSRcolor0[174]&LFSRcolor0[412]);
    BiasedRNG[6] = (LFSRcolor0[384]&LFSRcolor0[92]&LFSRcolor0[112]);
    BiasedRNG[7] = (LFSRcolor0[76]&LFSRcolor0[163]&LFSRcolor0[227]);
    BiasedRNG[8] = (LFSRcolor0[268]&LFSRcolor0[301]&LFSRcolor0[372]);
    BiasedRNG[9] = (LFSRcolor0[387]&LFSRcolor0[400]&LFSRcolor0[207]);
    BiasedRNG[10] = (LFSRcolor0[243]&LFSRcolor0[186]&LFSRcolor0[158]);
    BiasedRNG[11] = (LFSRcolor0[72]&LFSRcolor0[183]&LFSRcolor0[261]);
    BiasedRNG[12] = (LFSRcolor0[317]&LFSRcolor0[16]&LFSRcolor0[290]);
    BiasedRNG[13] = (LFSRcolor0[266]&LFSRcolor0[334]&LFSRcolor0[385]);
    BiasedRNG[14] = (LFSRcolor0[50]&LFSRcolor0[122]&LFSRcolor0[256]);
    BiasedRNG[15] = (LFSRcolor0[131]&LFSRcolor0[226]&LFSRcolor0[199]);
    BiasedRNG[16] = (LFSRcolor0[352]&LFSRcolor0[172]&LFSRcolor0[347]);
    BiasedRNG[17] = (LFSRcolor0[322]&LFSRcolor0[5]&LFSRcolor0[333]);
    BiasedRNG[18] = (LFSRcolor0[98]&LFSRcolor0[286]&LFSRcolor0[304]);
    BiasedRNG[19] = (LFSRcolor0[7]&LFSRcolor0[282]&LFSRcolor0[130]);
    BiasedRNG[20] = (LFSRcolor0[306]&LFSRcolor0[37]&LFSRcolor0[359]);
    BiasedRNG[21] = (LFSRcolor0[156]&LFSRcolor0[49]&LFSRcolor0[247]);
    BiasedRNG[22] = (LFSRcolor0[355]&LFSRcolor0[21]&LFSRcolor0[214]);
    BiasedRNG[23] = (LFSRcolor0[60]&LFSRcolor0[265]&LFSRcolor0[251]);
    BiasedRNG[24] = (LFSRcolor0[198]&LFSRcolor0[179]&LFSRcolor0[160]);
    BiasedRNG[25] = (LFSRcolor0[59]&LFSRcolor0[277]&LFSRcolor0[390]);
    BiasedRNG[26] = (LFSRcolor0[296]&LFSRcolor0[281]&LFSRcolor0[48]);
    BiasedRNG[27] = (LFSRcolor0[55]&LFSRcolor0[3]&LFSRcolor0[275]);
    BiasedRNG[28] = (LFSRcolor0[1]&LFSRcolor0[376]&LFSRcolor0[396]);
    BiasedRNG[29] = (LFSRcolor0[13]&LFSRcolor0[346]&LFSRcolor0[377]);
    BiasedRNG[30] = (LFSRcolor0[242]&LFSRcolor0[106]&LFSRcolor0[177]);
    BiasedRNG[31] = (LFSRcolor0[43]&LFSRcolor0[65]&LFSRcolor0[231]);
    BiasedRNG[32] = (LFSRcolor0[284]&LFSRcolor0[254]&LFSRcolor0[197]);
    BiasedRNG[33] = (LFSRcolor0[285]&LFSRcolor0[234]&LFSRcolor0[116]);
    BiasedRNG[34] = (LFSRcolor0[383]&LFSRcolor0[224]&LFSRcolor0[341]);
    BiasedRNG[35] = (LFSRcolor0[259]&LFSRcolor0[178]&LFSRcolor0[365]);
    BiasedRNG[36] = (LFSRcolor0[288]&LFSRcolor0[107]&LFSRcolor0[212]);
    BiasedRNG[37] = (LFSRcolor0[165]&LFSRcolor0[23]&LFSRcolor0[364]);
    BiasedRNG[38] = (LFSRcolor0[176]&LFSRcolor0[185]&LFSRcolor0[102]);
    BiasedRNG[39] = (LFSRcolor0[219]&LFSRcolor0[129]&LFSRcolor0[260]);
    BiasedRNG[40] = (LFSRcolor0[311]&LFSRcolor0[338]&LFSRcolor0[133]);
    BiasedRNG[41] = (LFSRcolor0[332]&LFSRcolor0[68]&LFSRcolor0[111]);
    BiasedRNG[42] = (LFSRcolor0[117]&LFSRcolor0[132]&LFSRcolor0[119]);
    BiasedRNG[43] = (LFSRcolor0[41]&LFSRcolor0[305]&LFSRcolor0[169]);
    BiasedRNG[44] = (LFSRcolor0[34]&LFSRcolor0[123]&LFSRcolor0[10]);
    BiasedRNG[45] = (LFSRcolor0[15]&LFSRcolor0[331]&LFSRcolor0[135]);
    BiasedRNG[46] = (LFSRcolor0[95]&LFSRcolor0[295]&LFSRcolor0[166]);
    BiasedRNG[47] = (LFSRcolor0[366]&LFSRcolor0[392]&LFSRcolor0[382]);
    BiasedRNG[48] = (LFSRcolor0[250]&LFSRcolor0[147]&LFSRcolor0[302]);
    BiasedRNG[49] = (LFSRcolor0[374]&LFSRcolor0[221]&LFSRcolor0[363]);
    BiasedRNG[50] = (LFSRcolor0[56]&LFSRcolor0[6]&LFSRcolor0[40]);
    BiasedRNG[51] = (LFSRcolor0[157]&LFSRcolor0[171]&LFSRcolor0[38]);
    BiasedRNG[52] = (LFSRcolor0[86]&LFSRcolor0[233]&LFSRcolor0[127]);
    BiasedRNG[53] = (LFSRcolor0[272]&LFSRcolor0[100]&LFSRcolor0[18]);
    BiasedRNG[54] = (LFSRcolor0[61]&LFSRcolor0[120]&LFSRcolor0[58]);
    BiasedRNG[55] = (LFSRcolor0[181]&LFSRcolor0[379]&LFSRcolor0[252]);
    BiasedRNG[56] = (LFSRcolor0[57]&LFSRcolor0[2]&LFSRcolor0[90]);
    BiasedRNG[57] = (LFSRcolor0[25]&LFSRcolor0[328]&LFSRcolor0[175]);
    BiasedRNG[58] = (LFSRcolor0[375]&LFSRcolor0[337]&LFSRcolor0[373]);
    BiasedRNG[59] = (LFSRcolor0[206]&LFSRcolor0[293]&LFSRcolor0[73]);
    BiasedRNG[60] = (LFSRcolor0[279]&LFSRcolor0[238]&LFSRcolor0[29]);
    BiasedRNG[61] = (LFSRcolor0[24]&LFSRcolor0[210]&LFSRcolor0[248]);
    BiasedRNG[62] = (LFSRcolor0[356]&LFSRcolor0[182]&LFSRcolor0[351]);
    BiasedRNG[63] = (LFSRcolor0[52]&LFSRcolor0[358]&LFSRcolor0[343]);
    BiasedRNG[64] = (LFSRcolor0[381]&LFSRcolor0[110]&LFSRcolor0[369]);
    BiasedRNG[65] = (LFSRcolor0[321]&LFSRcolor0[168]&LFSRcolor0[209]);
    BiasedRNG[66] = (LFSRcolor0[138]&LFSRcolor0[83]&LFSRcolor0[4]);
    BiasedRNG[67] = (LFSRcolor0[314]&LFSRcolor0[89]&LFSRcolor0[407]);
    BiasedRNG[68] = (LFSRcolor0[287]&LFSRcolor0[357]&LFSRcolor0[146]);
    BiasedRNG[69] = (LFSRcolor0[294]&LFSRcolor0[398]&LFSRcolor0[399]);
    BiasedRNG[70] = (LFSRcolor0[367]&LFSRcolor0[270]&LFSRcolor0[342]);
    BiasedRNG[71] = (LFSRcolor0[35]&LFSRcolor0[31]&LFSRcolor0[237]);
    BiasedRNG[72] = (LFSRcolor0[152]&LFSRcolor0[81]&LFSRcolor0[101]);
    BiasedRNG[73] = (LFSRcolor0[94]&LFSRcolor0[222]&LFSRcolor0[195]);
    BiasedRNG[74] = (LFSRcolor0[269]&LFSRcolor0[386]&LFSRcolor0[298]);
    BiasedRNG[75] = (LFSRcolor0[406]&LFSRcolor0[244]&LFSRcolor0[28]);
    BiasedRNG[76] = (LFSRcolor0[401]&LFSRcolor0[19]&LFSRcolor0[124]);
    BiasedRNG[77] = (LFSRcolor0[194]&LFSRcolor0[325]&LFSRcolor0[391]);
    BiasedRNG[78] = (LFSRcolor0[404]&LFSRcolor0[75]&LFSRcolor0[109]);
    BiasedRNG[79] = (LFSRcolor0[253]&LFSRcolor0[153]&LFSRcolor0[303]);
    BiasedRNG[80] = (LFSRcolor0[154]&LFSRcolor0[215]&LFSRcolor0[137]);
    BiasedRNG[81] = (LFSRcolor0[11]&LFSRcolor0[45]&LFSRcolor0[114]);
    BiasedRNG[82] = (LFSRcolor0[258]&LFSRcolor0[91]&LFSRcolor0[307]);
    BiasedRNG[83] = (LFSRcolor0[330]&LFSRcolor0[82]&LFSRcolor0[319]);
    BiasedRNG[84] = (LFSRcolor0[229]&LFSRcolor0[62]&LFSRcolor0[410]);
    BiasedRNG[85] = (LFSRcolor0[262]&LFSRcolor0[145]&LFSRcolor0[315]);
    BiasedRNG[86] = (LFSRcolor0[236]&LFSRcolor0[84]&LFSRcolor0[218]);
    BiasedRNG[87] = (LFSRcolor0[397]&LFSRcolor0[323]&LFSRcolor0[280]);
    BiasedRNG[88] = (LFSRcolor0[170]&LFSRcolor0[180]&LFSRcolor0[292]);
    BiasedRNG[89] = (LFSRcolor0[136]&LFSRcolor0[139]&LFSRcolor0[118]);
    BiasedRNG[90] = (LFSRcolor0[273]&LFSRcolor0[380]&LFSRcolor0[318]);
    BiasedRNG[91] = (LFSRcolor0[149]&LFSRcolor0[14]&LFSRcolor0[257]);
    BiasedRNG[92] = (LFSRcolor0[249]&LFSRcolor0[27]&LFSRcolor0[291]);
    BiasedRNG[93] = (LFSRcolor0[22]&LFSRcolor0[161]&LFSRcolor0[77]);
    BiasedRNG[94] = (LFSRcolor0[167]&LFSRcolor0[125]&LFSRcolor0[121]);
    BiasedRNG[95] = (LFSRcolor0[30]&LFSRcolor0[349]&LFSRcolor0[164]);
    BiasedRNG[96] = (LFSRcolor0[143]&LFSRcolor0[205]&LFSRcolor0[370]);
    BiasedRNG[97] = (LFSRcolor0[20]&LFSRcolor0[326]&LFSRcolor0[99]);
    BiasedRNG[98] = (LFSRcolor0[329]&LFSRcolor0[8]&LFSRcolor0[64]);
    UnbiasedRNG[0] = LFSRcolor0[239];
    UnbiasedRNG[1] = LFSRcolor0[32];
    UnbiasedRNG[2] = LFSRcolor0[193];
    UnbiasedRNG[3] = LFSRcolor0[232];
    UnbiasedRNG[4] = LFSRcolor0[402];
    UnbiasedRNG[5] = LFSRcolor0[312];
    UnbiasedRNG[6] = LFSRcolor0[267];
    UnbiasedRNG[7] = LFSRcolor0[47];
    UnbiasedRNG[8] = LFSRcolor0[200];
    UnbiasedRNG[9] = LFSRcolor0[204];
    UnbiasedRNG[10] = LFSRcolor0[213];
    UnbiasedRNG[11] = LFSRcolor0[53];
    UnbiasedRNG[12] = LFSRcolor0[241];
    UnbiasedRNG[13] = LFSRcolor0[228];
    UnbiasedRNG[14] = LFSRcolor0[162];
    UnbiasedRNG[15] = LFSRcolor0[246];
    UnbiasedRNG[16] = LFSRcolor0[151];
    UnbiasedRNG[17] = LFSRcolor0[128];
    UnbiasedRNG[18] = LFSRcolor0[344];
    UnbiasedRNG[19] = LFSRcolor0[276];
    UnbiasedRNG[20] = LFSRcolor0[33];
    UnbiasedRNG[21] = LFSRcolor0[66];
    UnbiasedRNG[22] = LFSRcolor0[235];
    UnbiasedRNG[23] = LFSRcolor0[278];
    UnbiasedRNG[24] = LFSRcolor0[196];
    UnbiasedRNG[25] = LFSRcolor0[217];
    UnbiasedRNG[26] = LFSRcolor0[271];
    UnbiasedRNG[27] = LFSRcolor0[96];
    UnbiasedRNG[28] = LFSRcolor0[202];
    UnbiasedRNG[29] = LFSRcolor0[230];
    UnbiasedRNG[30] = LFSRcolor0[316];
    UnbiasedRNG[31] = LFSRcolor0[140];
    UnbiasedRNG[32] = LFSRcolor0[192];
    UnbiasedRNG[33] = LFSRcolor0[148];
    UnbiasedRNG[34] = LFSRcolor0[190];
    UnbiasedRNG[35] = LFSRcolor0[191];
    UnbiasedRNG[36] = LFSRcolor0[360];
    UnbiasedRNG[37] = LFSRcolor0[104];
    UnbiasedRNG[38] = LFSRcolor0[335];
    UnbiasedRNG[39] = LFSRcolor0[184];
    UnbiasedRNG[40] = LFSRcolor0[85];
    UnbiasedRNG[41] = LFSRcolor0[17];
    UnbiasedRNG[42] = LFSRcolor0[105];
    UnbiasedRNG[43] = LFSRcolor0[299];
    UnbiasedRNG[44] = LFSRcolor0[216];
    UnbiasedRNG[45] = LFSRcolor0[327];
    UnbiasedRNG[46] = LFSRcolor0[297];
    UnbiasedRNG[47] = LFSRcolor0[240];
    UnbiasedRNG[48] = LFSRcolor0[126];
    UnbiasedRNG[49] = LFSRcolor0[368];
    UnbiasedRNG[50] = LFSRcolor0[187];
    UnbiasedRNG[51] = LFSRcolor0[308];
    UnbiasedRNG[52] = LFSRcolor0[223];
    UnbiasedRNG[53] = LFSRcolor0[245];
    UnbiasedRNG[54] = LFSRcolor0[39];
    UnbiasedRNG[55] = LFSRcolor0[353];
    UnbiasedRNG[56] = LFSRcolor0[313];
    UnbiasedRNG[57] = LFSRcolor0[9];
    UnbiasedRNG[58] = LFSRcolor0[26];
    UnbiasedRNG[59] = LFSRcolor0[393];
    UnbiasedRNG[60] = LFSRcolor0[51];
    UnbiasedRNG[61] = LFSRcolor0[220];
    UnbiasedRNG[62] = LFSRcolor0[97];
    UnbiasedRNG[63] = LFSRcolor0[78];
    UnbiasedRNG[64] = LFSRcolor0[144];
    UnbiasedRNG[65] = LFSRcolor0[88];
    UnbiasedRNG[66] = LFSRcolor0[80];
    UnbiasedRNG[67] = LFSRcolor0[300];
    UnbiasedRNG[68] = LFSRcolor0[263];
    UnbiasedRNG[69] = LFSRcolor0[0];
    UnbiasedRNG[70] = LFSRcolor0[225];
    UnbiasedRNG[71] = LFSRcolor0[67];
    UnbiasedRNG[72] = LFSRcolor0[320];
    UnbiasedRNG[73] = LFSRcolor0[134];
    UnbiasedRNG[74] = LFSRcolor0[188];
    UnbiasedRNG[75] = LFSRcolor0[289];
    UnbiasedRNG[76] = LFSRcolor0[103];
    UnbiasedRNG[77] = LFSRcolor0[150];
    UnbiasedRNG[78] = LFSRcolor0[189];
    UnbiasedRNG[79] = LFSRcolor0[394];
    UnbiasedRNG[80] = LFSRcolor0[93];
    UnbiasedRNG[81] = LFSRcolor0[141];
    UnbiasedRNG[82] = LFSRcolor0[339];
    UnbiasedRNG[83] = LFSRcolor0[336];
    UnbiasedRNG[84] = LFSRcolor0[411];
    UnbiasedRNG[85] = LFSRcolor0[309];
    UnbiasedRNG[86] = LFSRcolor0[79];
    UnbiasedRNG[87] = LFSRcolor0[70];
    UnbiasedRNG[88] = LFSRcolor0[87];
    UnbiasedRNG[89] = LFSRcolor0[408];
    UnbiasedRNG[90] = LFSRcolor0[324];
    UnbiasedRNG[91] = LFSRcolor0[46];
    UnbiasedRNG[92] = LFSRcolor0[113];
    UnbiasedRNG[93] = LFSRcolor0[115];
    UnbiasedRNG[94] = LFSRcolor0[362];
    UnbiasedRNG[95] = LFSRcolor0[405];
    UnbiasedRNG[96] = LFSRcolor0[173];
    UnbiasedRNG[97] = LFSRcolor0[201];
    UnbiasedRNG[98] = LFSRcolor0[361];
    UnbiasedRNG[99] = LFSRcolor0[42];
    UnbiasedRNG[100] = LFSRcolor0[255];
    UnbiasedRNG[101] = LFSRcolor0[348];
    UnbiasedRNG[102] = LFSRcolor0[108];
    UnbiasedRNG[103] = LFSRcolor0[345];
    UnbiasedRNG[104] = LFSRcolor0[283];
    UnbiasedRNG[105] = LFSRcolor0[310];
    UnbiasedRNG[106] = LFSRcolor0[142];
    UnbiasedRNG[107] = LFSRcolor0[63];
end

always @(posedge color0_clk) begin
    BiasedRNG[99] = (LFSRcolor1[331]&LFSRcolor1[67]&LFSRcolor1[69]);
    BiasedRNG[100] = (LFSRcolor1[89]&LFSRcolor1[282]&LFSRcolor1[19]);
    BiasedRNG[101] = (LFSRcolor1[470]&LFSRcolor1[166]&LFSRcolor1[531]);
    BiasedRNG[102] = (LFSRcolor1[246]&LFSRcolor1[494]&LFSRcolor1[493]);
    BiasedRNG[103] = (LFSRcolor1[262]&LFSRcolor1[290]&LFSRcolor1[130]);
    BiasedRNG[104] = (LFSRcolor1[103]&LFSRcolor1[272]&LFSRcolor1[491]);
    BiasedRNG[105] = (LFSRcolor1[17]&LFSRcolor1[462]&LFSRcolor1[160]);
    BiasedRNG[106] = (LFSRcolor1[530]&LFSRcolor1[525]&LFSRcolor1[140]);
    BiasedRNG[107] = (LFSRcolor1[203]&LFSRcolor1[253]&LFSRcolor1[116]);
    BiasedRNG[108] = (LFSRcolor1[247]&LFSRcolor1[469]&LFSRcolor1[52]);
    BiasedRNG[109] = (LFSRcolor1[128]&LFSRcolor1[409]&LFSRcolor1[218]);
    BiasedRNG[110] = (LFSRcolor1[417]&LFSRcolor1[327]&LFSRcolor1[308]);
    BiasedRNG[111] = (LFSRcolor1[162]&LFSRcolor1[446]&LFSRcolor1[47]);
    BiasedRNG[112] = (LFSRcolor1[480]&LFSRcolor1[392]&LFSRcolor1[377]);
    BiasedRNG[113] = (LFSRcolor1[447]&LFSRcolor1[520]&LFSRcolor1[92]);
    BiasedRNG[114] = (LFSRcolor1[210]&LFSRcolor1[68]&LFSRcolor1[81]);
    BiasedRNG[115] = (LFSRcolor1[232]&LFSRcolor1[418]&LFSRcolor1[41]);
    BiasedRNG[116] = (LFSRcolor1[535]&LFSRcolor1[234]&LFSRcolor1[400]);
    BiasedRNG[117] = (LFSRcolor1[289]&LFSRcolor1[74]&LFSRcolor1[291]);
    BiasedRNG[118] = (LFSRcolor1[102]&LFSRcolor1[159]&LFSRcolor1[33]);
    BiasedRNG[119] = (LFSRcolor1[224]&LFSRcolor1[50]&LFSRcolor1[178]);
    BiasedRNG[120] = (LFSRcolor1[57]&LFSRcolor1[550]&LFSRcolor1[292]);
    BiasedRNG[121] = (LFSRcolor1[135]&LFSRcolor1[302]&LFSRcolor1[396]);
    BiasedRNG[122] = (LFSRcolor1[547]&LFSRcolor1[346]&LFSRcolor1[222]);
    BiasedRNG[123] = (LFSRcolor1[402]&LFSRcolor1[53]&LFSRcolor1[95]);
    BiasedRNG[124] = (LFSRcolor1[112]&LFSRcolor1[245]&LFSRcolor1[212]);
    BiasedRNG[125] = (LFSRcolor1[24]&LFSRcolor1[342]&LFSRcolor1[411]);
    BiasedRNG[126] = (LFSRcolor1[169]&LFSRcolor1[269]&LFSRcolor1[475]);
    BiasedRNG[127] = (LFSRcolor1[482]&LFSRcolor1[181]&LFSRcolor1[223]);
    BiasedRNG[128] = (LFSRcolor1[157]&LFSRcolor1[455]&LFSRcolor1[215]);
    BiasedRNG[129] = (LFSRcolor1[254]&LFSRcolor1[349]&LFSRcolor1[478]);
    BiasedRNG[130] = (LFSRcolor1[229]&LFSRcolor1[288]&LFSRcolor1[388]);
    BiasedRNG[131] = (LFSRcolor1[529]&LFSRcolor1[179]&LFSRcolor1[412]);
    BiasedRNG[132] = (LFSRcolor1[73]&LFSRcolor1[184]&LFSRcolor1[295]);
    BiasedRNG[133] = (LFSRcolor1[176]&LFSRcolor1[216]&LFSRcolor1[136]);
    BiasedRNG[134] = (LFSRcolor1[158]&LFSRcolor1[40]&LFSRcolor1[523]);
    BiasedRNG[135] = (LFSRcolor1[370]&LFSRcolor1[72]&LFSRcolor1[512]);
    BiasedRNG[136] = (LFSRcolor1[114]&LFSRcolor1[153]&LFSRcolor1[382]);
    BiasedRNG[137] = (LFSRcolor1[268]&LFSRcolor1[543]&LFSRcolor1[318]);
    BiasedRNG[138] = (LFSRcolor1[167]&LFSRcolor1[298]&LFSRcolor1[362]);
    BiasedRNG[139] = (LFSRcolor1[98]&LFSRcolor1[301]&LFSRcolor1[275]);
    BiasedRNG[140] = (LFSRcolor1[249]&LFSRcolor1[326]&LFSRcolor1[197]);
    BiasedRNG[141] = (LFSRcolor1[123]&LFSRcolor1[80]&LFSRcolor1[427]);
    BiasedRNG[142] = (LFSRcolor1[26]&LFSRcolor1[406]&LFSRcolor1[479]);
    BiasedRNG[143] = (LFSRcolor1[42]&LFSRcolor1[451]&LFSRcolor1[338]);
    BiasedRNG[144] = (LFSRcolor1[363]&LFSRcolor1[536]&LFSRcolor1[97]);
    BiasedRNG[145] = (LFSRcolor1[38]&LFSRcolor1[294]&LFSRcolor1[344]);
    BiasedRNG[146] = (LFSRcolor1[329]&LFSRcolor1[60]&LFSRcolor1[271]);
    BiasedRNG[147] = (LFSRcolor1[231]&LFSRcolor1[424]&LFSRcolor1[0]);
    BiasedRNG[148] = (LFSRcolor1[23]&LFSRcolor1[433]&LFSRcolor1[214]);
    BiasedRNG[149] = (LFSRcolor1[78]&LFSRcolor1[273]&LFSRcolor1[30]);
    BiasedRNG[150] = (LFSRcolor1[460]&LFSRcolor1[445]&LFSRcolor1[332]);
    BiasedRNG[151] = (LFSRcolor1[325]&LFSRcolor1[55]&LFSRcolor1[172]);
    BiasedRNG[152] = (LFSRcolor1[175]&LFSRcolor1[339]&LFSRcolor1[449]);
    BiasedRNG[153] = (LFSRcolor1[351]&LFSRcolor1[39]&LFSRcolor1[439]);
    BiasedRNG[154] = (LFSRcolor1[414]&LFSRcolor1[526]&LFSRcolor1[532]);
    BiasedRNG[155] = (LFSRcolor1[36]&LFSRcolor1[313]&LFSRcolor1[322]);
    BiasedRNG[156] = (LFSRcolor1[452]&LFSRcolor1[152]&LFSRcolor1[101]);
    BiasedRNG[157] = (LFSRcolor1[94]&LFSRcolor1[147]&LFSRcolor1[538]);
    BiasedRNG[158] = (LFSRcolor1[328]&LFSRcolor1[28]&LFSRcolor1[261]);
    BiasedRNG[159] = (LFSRcolor1[236]&LFSRcolor1[255]&LFSRcolor1[546]);
    BiasedRNG[160] = (LFSRcolor1[1]&LFSRcolor1[539]&LFSRcolor1[165]);
    BiasedRNG[161] = (LFSRcolor1[353]&LFSRcolor1[537]&LFSRcolor1[3]);
    BiasedRNG[162] = (LFSRcolor1[155]&LFSRcolor1[58]&LFSRcolor1[144]);
    BiasedRNG[163] = (LFSRcolor1[143]&LFSRcolor1[134]&LFSRcolor1[62]);
    BiasedRNG[164] = (LFSRcolor1[117]&LFSRcolor1[173]&LFSRcolor1[208]);
    BiasedRNG[165] = (LFSRcolor1[228]&LFSRcolor1[148]&LFSRcolor1[122]);
    BiasedRNG[166] = (LFSRcolor1[35]&LFSRcolor1[337]&LFSRcolor1[335]);
    BiasedRNG[167] = (LFSRcolor1[336]&LFSRcolor1[201]&LFSRcolor1[518]);
    BiasedRNG[168] = (LFSRcolor1[86]&LFSRcolor1[421]&LFSRcolor1[473]);
    BiasedRNG[169] = (LFSRcolor1[507]&LFSRcolor1[321]&LFSRcolor1[474]);
    BiasedRNG[170] = (LFSRcolor1[503]&LFSRcolor1[263]&LFSRcolor1[260]);
    BiasedRNG[171] = (LFSRcolor1[368]&LFSRcolor1[186]&LFSRcolor1[476]);
    BiasedRNG[172] = (LFSRcolor1[391]&LFSRcolor1[459]&LFSRcolor1[2]);
    BiasedRNG[173] = (LFSRcolor1[293]&LFSRcolor1[506]&LFSRcolor1[516]);
    BiasedRNG[174] = (LFSRcolor1[49]&LFSRcolor1[59]&LFSRcolor1[65]);
    BiasedRNG[175] = (LFSRcolor1[513]&LFSRcolor1[180]&LFSRcolor1[366]);
    BiasedRNG[176] = (LFSRcolor1[450]&LFSRcolor1[32]&LFSRcolor1[468]);
    BiasedRNG[177] = (LFSRcolor1[367]&LFSRcolor1[490]&LFSRcolor1[204]);
    BiasedRNG[178] = (LFSRcolor1[248]&LFSRcolor1[185]&LFSRcolor1[299]);
    BiasedRNG[179] = (LFSRcolor1[434]&LFSRcolor1[287]&LFSRcolor1[238]);
    BiasedRNG[180] = (LFSRcolor1[357]&LFSRcolor1[22]&LFSRcolor1[227]);
    BiasedRNG[181] = (LFSRcolor1[82]&LFSRcolor1[10]&LFSRcolor1[296]);
    BiasedRNG[182] = (LFSRcolor1[405]&LFSRcolor1[14]&LFSRcolor1[124]);
    BiasedRNG[183] = (LFSRcolor1[315]&LFSRcolor1[458]&LFSRcolor1[241]);
    BiasedRNG[184] = (LFSRcolor1[12]&LFSRcolor1[316]&LFSRcolor1[190]);
    BiasedRNG[185] = (LFSRcolor1[499]&LFSRcolor1[4]&LFSRcolor1[483]);
    BiasedRNG[186] = (LFSRcolor1[11]&LFSRcolor1[467]&LFSRcolor1[8]);
    BiasedRNG[187] = (LFSRcolor1[384]&LFSRcolor1[425]&LFSRcolor1[211]);
    BiasedRNG[188] = (LFSRcolor1[380]&LFSRcolor1[435]&LFSRcolor1[266]);
    BiasedRNG[189] = (LFSRcolor1[311]&LFSRcolor1[375]&LFSRcolor1[386]);
    BiasedRNG[190] = (LFSRcolor1[436]&LFSRcolor1[70]&LFSRcolor1[286]);
    BiasedRNG[191] = (LFSRcolor1[171]&LFSRcolor1[240]&LFSRcolor1[151]);
    BiasedRNG[192] = (LFSRcolor1[132]&LFSRcolor1[456]&LFSRcolor1[355]);
    BiasedRNG[193] = (LFSRcolor1[205]&LFSRcolor1[361]&LFSRcolor1[256]);
    BiasedRNG[194] = (LFSRcolor1[509]&LFSRcolor1[358]&LFSRcolor1[438]);
    BiasedRNG[195] = (LFSRcolor1[527]&LFSRcolor1[235]&LFSRcolor1[258]);
    BiasedRNG[196] = (LFSRcolor1[200]&LFSRcolor1[484]&LFSRcolor1[113]);
    BiasedRNG[197] = (LFSRcolor1[463]&LFSRcolor1[374]&LFSRcolor1[45]);
    BiasedRNG[198] = (LFSRcolor1[317]&LFSRcolor1[307]&LFSRcolor1[549]);
    BiasedRNG[199] = (LFSRcolor1[407]&LFSRcolor1[27]&LFSRcolor1[192]);
    BiasedRNG[200] = (LFSRcolor1[304]&LFSRcolor1[133]&LFSRcolor1[161]);
    BiasedRNG[201] = (LFSRcolor1[76]&LFSRcolor1[533]&LFSRcolor1[330]);
    BiasedRNG[202] = (LFSRcolor1[466]&LFSRcolor1[220]&LFSRcolor1[515]);
    BiasedRNG[203] = (LFSRcolor1[381]&LFSRcolor1[429]&LFSRcolor1[371]);
    BiasedRNG[204] = (LFSRcolor1[394]&LFSRcolor1[163]&LFSRcolor1[442]);
    BiasedRNG[205] = (LFSRcolor1[504]&LFSRcolor1[309]&LFSRcolor1[149]);
    BiasedRNG[206] = (LFSRcolor1[448]&LFSRcolor1[511]&LFSRcolor1[221]);
    BiasedRNG[207] = (LFSRcolor1[109]&LFSRcolor1[115]&LFSRcolor1[63]);
    BiasedRNG[208] = (LFSRcolor1[489]&LFSRcolor1[43]&LFSRcolor1[419]);
    BiasedRNG[209] = (LFSRcolor1[372]&LFSRcolor1[306]&LFSRcolor1[267]);
    BiasedRNG[210] = (LFSRcolor1[90]&LFSRcolor1[541]&LFSRcolor1[111]);
    BiasedRNG[211] = (LFSRcolor1[120]&LFSRcolor1[343]&LFSRcolor1[110]);
    BiasedRNG[212] = (LFSRcolor1[281]&LFSRcolor1[194]&LFSRcolor1[347]);
    BiasedRNG[213] = (LFSRcolor1[233]&LFSRcolor1[310]&LFSRcolor1[18]);
    BiasedRNG[214] = (LFSRcolor1[395]&LFSRcolor1[303]&LFSRcolor1[5]);
    BiasedRNG[215] = (LFSRcolor1[426]&LFSRcolor1[79]&LFSRcolor1[164]);
    BiasedRNG[216] = (LFSRcolor1[100]&LFSRcolor1[487]&LFSRcolor1[9]);
    BiasedRNG[217] = (LFSRcolor1[219]&LFSRcolor1[283]&LFSRcolor1[510]);
    BiasedRNG[218] = (LFSRcolor1[84]&LFSRcolor1[237]&LFSRcolor1[142]);
    BiasedRNG[219] = (LFSRcolor1[521]&LFSRcolor1[416]&LFSRcolor1[244]);
    BiasedRNG[220] = (LFSRcolor1[46]&LFSRcolor1[48]&LFSRcolor1[437]);
    BiasedRNG[221] = (LFSRcolor1[56]&LFSRcolor1[334]&LFSRcolor1[430]);
    BiasedRNG[222] = (LFSRcolor1[385]&LFSRcolor1[202]&LFSRcolor1[420]);
    BiasedRNG[223] = (LFSRcolor1[51]&LFSRcolor1[193]&LFSRcolor1[492]);
    BiasedRNG[224] = (LFSRcolor1[548]&LFSRcolor1[187]&LFSRcolor1[376]);
    BiasedRNG[225] = (LFSRcolor1[383]&LFSRcolor1[323]&LFSRcolor1[496]);
    BiasedRNG[226] = (LFSRcolor1[64]&LFSRcolor1[191]&LFSRcolor1[314]);
    BiasedRNG[227] = (LFSRcolor1[551]&LFSRcolor1[119]&LFSRcolor1[410]);
    BiasedRNG[228] = (LFSRcolor1[196]&LFSRcolor1[213]&LFSRcolor1[230]);
    BiasedRNG[229] = (LFSRcolor1[251]&LFSRcolor1[514]&LFSRcolor1[156]);
    BiasedRNG[230] = (LFSRcolor1[183]&LFSRcolor1[545]&LFSRcolor1[305]);
    BiasedRNG[231] = (LFSRcolor1[542]&LFSRcolor1[486]&LFSRcolor1[390]);
    BiasedRNG[232] = (LFSRcolor1[508]&LFSRcolor1[472]&LFSRcolor1[501]);
    BiasedRNG[233] = (LFSRcolor1[397]&LFSRcolor1[239]&LFSRcolor1[198]);
    BiasedRNG[234] = (LFSRcolor1[127]&LFSRcolor1[279]&LFSRcolor1[29]);
    BiasedRNG[235] = (LFSRcolor1[519]&LFSRcolor1[398]&LFSRcolor1[243]);
    BiasedRNG[236] = (LFSRcolor1[195]&LFSRcolor1[77]&LFSRcolor1[96]);
    BiasedRNG[237] = (LFSRcolor1[71]&LFSRcolor1[422]&LFSRcolor1[502]);
    BiasedRNG[238] = (LFSRcolor1[131]&LFSRcolor1[145]&LFSRcolor1[93]);
    UnbiasedRNG[108] = LFSRcolor1[121];
    UnbiasedRNG[109] = LFSRcolor1[454];
    UnbiasedRNG[110] = LFSRcolor1[284];
    UnbiasedRNG[111] = LFSRcolor1[364];
    UnbiasedRNG[112] = LFSRcolor1[108];
    UnbiasedRNG[113] = LFSRcolor1[83];
    UnbiasedRNG[114] = LFSRcolor1[21];
    UnbiasedRNG[115] = LFSRcolor1[365];
    UnbiasedRNG[116] = LFSRcolor1[403];
    UnbiasedRNG[117] = LFSRcolor1[415];
    UnbiasedRNG[118] = LFSRcolor1[280];
    UnbiasedRNG[119] = LFSRcolor1[276];
    UnbiasedRNG[120] = LFSRcolor1[354];
    UnbiasedRNG[121] = LFSRcolor1[528];
    UnbiasedRNG[122] = LFSRcolor1[373];
    UnbiasedRNG[123] = LFSRcolor1[524];
    UnbiasedRNG[124] = LFSRcolor1[413];
    UnbiasedRNG[125] = LFSRcolor1[440];
    UnbiasedRNG[126] = LFSRcolor1[319];
    UnbiasedRNG[127] = LFSRcolor1[500];
    UnbiasedRNG[128] = LFSRcolor1[350];
    UnbiasedRNG[129] = LFSRcolor1[300];
    UnbiasedRNG[130] = LFSRcolor1[252];
    UnbiasedRNG[131] = LFSRcolor1[259];
    UnbiasedRNG[132] = LFSRcolor1[150];
    UnbiasedRNG[133] = LFSRcolor1[225];
    UnbiasedRNG[134] = LFSRcolor1[278];
    UnbiasedRNG[135] = LFSRcolor1[444];
    UnbiasedRNG[136] = LFSRcolor1[188];
    UnbiasedRNG[137] = LFSRcolor1[360];
    UnbiasedRNG[138] = LFSRcolor1[477];
    UnbiasedRNG[139] = LFSRcolor1[189];
    UnbiasedRNG[140] = LFSRcolor1[387];
    UnbiasedRNG[141] = LFSRcolor1[379];
    UnbiasedRNG[142] = LFSRcolor1[107];
    UnbiasedRNG[143] = LFSRcolor1[378];
    UnbiasedRNG[144] = LFSRcolor1[498];
    UnbiasedRNG[145] = LFSRcolor1[320];
    UnbiasedRNG[146] = LFSRcolor1[404];
    UnbiasedRNG[147] = LFSRcolor1[105];
    UnbiasedRNG[148] = LFSRcolor1[401];
    UnbiasedRNG[149] = LFSRcolor1[348];
    UnbiasedRNG[150] = LFSRcolor1[88];
    UnbiasedRNG[151] = LFSRcolor1[250];
    UnbiasedRNG[152] = LFSRcolor1[226];
    UnbiasedRNG[153] = LFSRcolor1[138];
    UnbiasedRNG[154] = LFSRcolor1[125];
    UnbiasedRNG[155] = LFSRcolor1[505];
    UnbiasedRNG[156] = LFSRcolor1[129];
    UnbiasedRNG[157] = LFSRcolor1[497];
    UnbiasedRNG[158] = LFSRcolor1[146];
    UnbiasedRNG[159] = LFSRcolor1[168];
    UnbiasedRNG[160] = LFSRcolor1[517];
    UnbiasedRNG[161] = LFSRcolor1[182];
    UnbiasedRNG[162] = LFSRcolor1[91];
    UnbiasedRNG[163] = LFSRcolor1[432];
    UnbiasedRNG[164] = LFSRcolor1[481];
    UnbiasedRNG[165] = LFSRcolor1[356];
    UnbiasedRNG[166] = LFSRcolor1[441];
    UnbiasedRNG[167] = LFSRcolor1[461];
    UnbiasedRNG[168] = LFSRcolor1[20];
    UnbiasedRNG[169] = LFSRcolor1[126];
    UnbiasedRNG[170] = LFSRcolor1[177];
    UnbiasedRNG[171] = LFSRcolor1[137];
    UnbiasedRNG[172] = LFSRcolor1[522];
    UnbiasedRNG[173] = LFSRcolor1[37];
    UnbiasedRNG[174] = LFSRcolor1[485];
    UnbiasedRNG[175] = LFSRcolor1[393];
    UnbiasedRNG[176] = LFSRcolor1[139];
    UnbiasedRNG[177] = LFSRcolor1[25];
    UnbiasedRNG[178] = LFSRcolor1[217];
    UnbiasedRNG[179] = LFSRcolor1[31];
    UnbiasedRNG[180] = LFSRcolor1[341];
    UnbiasedRNG[181] = LFSRcolor1[408];
    UnbiasedRNG[182] = LFSRcolor1[285];
    UnbiasedRNG[183] = LFSRcolor1[352];
    UnbiasedRNG[184] = LFSRcolor1[274];
    UnbiasedRNG[185] = LFSRcolor1[443];
    UnbiasedRNG[186] = LFSRcolor1[141];
    UnbiasedRNG[187] = LFSRcolor1[333];
    UnbiasedRNG[188] = LFSRcolor1[465];
    UnbiasedRNG[189] = LFSRcolor1[431];
    UnbiasedRNG[190] = LFSRcolor1[265];
    UnbiasedRNG[191] = LFSRcolor1[16];
    UnbiasedRNG[192] = LFSRcolor1[54];
    UnbiasedRNG[193] = LFSRcolor1[340];
    UnbiasedRNG[194] = LFSRcolor1[15];
    UnbiasedRNG[195] = LFSRcolor1[389];
    UnbiasedRNG[196] = LFSRcolor1[534];
    UnbiasedRNG[197] = LFSRcolor1[104];
end

always @(posedge color1_clk) begin
    BiasedRNG[239] = (LFSRcolor2[239]&LFSRcolor2[295]&LFSRcolor2[341]);
    BiasedRNG[240] = (LFSRcolor2[135]&LFSRcolor2[219]&LFSRcolor2[331]);
    BiasedRNG[241] = (LFSRcolor2[45]&LFSRcolor2[62]&LFSRcolor2[247]);
    BiasedRNG[242] = (LFSRcolor2[388]&LFSRcolor2[71]&LFSRcolor2[406]);
    BiasedRNG[243] = (LFSRcolor2[90]&LFSRcolor2[41]&LFSRcolor2[187]);
    BiasedRNG[244] = (LFSRcolor2[377]&LFSRcolor2[384]&LFSRcolor2[292]);
    BiasedRNG[245] = (LFSRcolor2[407]&LFSRcolor2[28]&LFSRcolor2[191]);
    BiasedRNG[246] = (LFSRcolor2[117]&LFSRcolor2[33]&LFSRcolor2[404]);
    BiasedRNG[247] = (LFSRcolor2[189]&LFSRcolor2[397]&LFSRcolor2[125]);
    BiasedRNG[248] = (LFSRcolor2[25]&LFSRcolor2[227]&LFSRcolor2[196]);
    BiasedRNG[249] = (LFSRcolor2[112]&LFSRcolor2[48]&LFSRcolor2[380]);
    BiasedRNG[250] = (LFSRcolor2[336]&LFSRcolor2[305]&LFSRcolor2[365]);
    BiasedRNG[251] = (LFSRcolor2[356]&LFSRcolor2[87]&LFSRcolor2[316]);
    BiasedRNG[252] = (LFSRcolor2[11]&LFSRcolor2[127]&LFSRcolor2[378]);
    BiasedRNG[253] = (LFSRcolor2[96]&LFSRcolor2[287]&LFSRcolor2[166]);
    BiasedRNG[254] = (LFSRcolor2[75]&LFSRcolor2[134]&LFSRcolor2[6]);
    BiasedRNG[255] = (LFSRcolor2[374]&LFSRcolor2[333]&LFSRcolor2[172]);
    BiasedRNG[256] = (LFSRcolor2[73]&LFSRcolor2[88]&LFSRcolor2[58]);
    BiasedRNG[257] = (LFSRcolor2[398]&LFSRcolor2[355]&LFSRcolor2[139]);
    BiasedRNG[258] = (LFSRcolor2[201]&LFSRcolor2[138]&LFSRcolor2[146]);
    BiasedRNG[259] = (LFSRcolor2[206]&LFSRcolor2[129]&LFSRcolor2[349]);
    BiasedRNG[260] = (LFSRcolor2[133]&LFSRcolor2[317]&LFSRcolor2[268]);
    BiasedRNG[261] = (LFSRcolor2[325]&LFSRcolor2[154]&LFSRcolor2[213]);
    BiasedRNG[262] = (LFSRcolor2[385]&LFSRcolor2[106]&LFSRcolor2[392]);
    BiasedRNG[263] = (LFSRcolor2[221]&LFSRcolor2[65]&LFSRcolor2[362]);
    BiasedRNG[264] = (LFSRcolor2[38]&LFSRcolor2[400]&LFSRcolor2[181]);
    BiasedRNG[265] = (LFSRcolor2[144]&LFSRcolor2[83]&LFSRcolor2[2]);
    BiasedRNG[266] = (LFSRcolor2[202]&LFSRcolor2[303]&LFSRcolor2[238]);
    BiasedRNG[267] = (LFSRcolor2[97]&LFSRcolor2[311]&LFSRcolor2[59]);
    BiasedRNG[268] = (LFSRcolor2[32]&LFSRcolor2[399]&LFSRcolor2[160]);
    BiasedRNG[269] = (LFSRcolor2[282]&LFSRcolor2[80]&LFSRcolor2[12]);
    BiasedRNG[270] = (LFSRcolor2[225]&LFSRcolor2[35]&LFSRcolor2[193]);
    BiasedRNG[271] = (LFSRcolor2[366]&LFSRcolor2[405]&LFSRcolor2[68]);
    BiasedRNG[272] = (LFSRcolor2[164]&LFSRcolor2[148]&LFSRcolor2[61]);
    BiasedRNG[273] = (LFSRcolor2[15]&LFSRcolor2[115]&LFSRcolor2[122]);
    BiasedRNG[274] = (LFSRcolor2[288]&LFSRcolor2[168]&LFSRcolor2[77]);
    BiasedRNG[275] = (LFSRcolor2[343]&LFSRcolor2[232]&LFSRcolor2[159]);
    BiasedRNG[276] = (LFSRcolor2[389]&LFSRcolor2[260]&LFSRcolor2[315]);
    BiasedRNG[277] = (LFSRcolor2[264]&LFSRcolor2[228]&LFSRcolor2[137]);
    BiasedRNG[278] = (LFSRcolor2[4]&LFSRcolor2[103]&LFSRcolor2[81]);
    BiasedRNG[279] = (LFSRcolor2[214]&LFSRcolor2[396]&LFSRcolor2[40]);
    BiasedRNG[280] = (LFSRcolor2[391]&LFSRcolor2[205]&LFSRcolor2[57]);
    BiasedRNG[281] = (LFSRcolor2[373]&LFSRcolor2[308]&LFSRcolor2[177]);
    BiasedRNG[282] = (LFSRcolor2[158]&LFSRcolor2[310]&LFSRcolor2[116]);
    BiasedRNG[283] = (LFSRcolor2[153]&LFSRcolor2[169]&LFSRcolor2[176]);
    BiasedRNG[284] = (LFSRcolor2[14]&LFSRcolor2[155]&LFSRcolor2[229]);
    BiasedRNG[285] = (LFSRcolor2[285]&LFSRcolor2[7]&LFSRcolor2[344]);
    BiasedRNG[286] = (LFSRcolor2[5]&LFSRcolor2[387]&LFSRcolor2[237]);
    BiasedRNG[287] = (LFSRcolor2[203]&LFSRcolor2[222]&LFSRcolor2[171]);
    BiasedRNG[288] = (LFSRcolor2[283]&LFSRcolor2[314]&LFSRcolor2[18]);
    BiasedRNG[289] = (LFSRcolor2[353]&LFSRcolor2[321]&LFSRcolor2[174]);
    BiasedRNG[290] = (LFSRcolor2[246]&LFSRcolor2[132]&LFSRcolor2[242]);
    BiasedRNG[291] = (LFSRcolor2[141]&LFSRcolor2[34]&LFSRcolor2[270]);
    BiasedRNG[292] = (LFSRcolor2[263]&LFSRcolor2[412]&LFSRcolor2[276]);
    BiasedRNG[293] = (LFSRcolor2[383]&LFSRcolor2[324]&LFSRcolor2[3]);
    BiasedRNG[294] = (LFSRcolor2[121]&LFSRcolor2[79]&LFSRcolor2[267]);
    BiasedRNG[295] = (LFSRcolor2[1]&LFSRcolor2[379]&LFSRcolor2[386]);
    BiasedRNG[296] = (LFSRcolor2[30]&LFSRcolor2[199]&LFSRcolor2[175]);
    BiasedRNG[297] = (LFSRcolor2[51]&LFSRcolor2[302]&LFSRcolor2[275]);
    BiasedRNG[298] = (LFSRcolor2[266]&LFSRcolor2[29]&LFSRcolor2[210]);
    BiasedRNG[299] = (LFSRcolor2[367]&LFSRcolor2[256]&LFSRcolor2[52]);
    BiasedRNG[300] = (LFSRcolor2[351]&LFSRcolor2[329]&LFSRcolor2[277]);
    BiasedRNG[301] = (LFSRcolor2[198]&LFSRcolor2[190]&LFSRcolor2[332]);
    BiasedRNG[302] = (LFSRcolor2[364]&LFSRcolor2[274]&LFSRcolor2[265]);
    BiasedRNG[303] = (LFSRcolor2[179]&LFSRcolor2[13]&LFSRcolor2[24]);
    BiasedRNG[304] = (LFSRcolor2[212]&LFSRcolor2[31]&LFSRcolor2[352]);
    BiasedRNG[305] = (LFSRcolor2[124]&LFSRcolor2[224]&LFSRcolor2[255]);
    BiasedRNG[306] = (LFSRcolor2[244]&LFSRcolor2[233]&LFSRcolor2[312]);
    BiasedRNG[307] = (LFSRcolor2[330]&LFSRcolor2[78]&LFSRcolor2[100]);
    BiasedRNG[308] = (LFSRcolor2[16]&LFSRcolor2[252]&LFSRcolor2[180]);
    BiasedRNG[309] = (LFSRcolor2[163]&LFSRcolor2[50]&LFSRcolor2[408]);
    BiasedRNG[310] = (LFSRcolor2[131]&LFSRcolor2[394]&LFSRcolor2[149]);
    BiasedRNG[311] = (LFSRcolor2[220]&LFSRcolor2[74]&LFSRcolor2[85]);
    BiasedRNG[312] = (LFSRcolor2[216]&LFSRcolor2[147]&LFSRcolor2[371]);
    BiasedRNG[313] = (LFSRcolor2[358]&LFSRcolor2[271]&LFSRcolor2[409]);
    BiasedRNG[314] = (LFSRcolor2[84]&LFSRcolor2[92]&LFSRcolor2[248]);
    BiasedRNG[315] = (LFSRcolor2[64]&LFSRcolor2[357]&LFSRcolor2[323]);
    BiasedRNG[316] = (LFSRcolor2[300]&LFSRcolor2[347]&LFSRcolor2[91]);
    BiasedRNG[317] = (LFSRcolor2[338]&LFSRcolor2[286]&LFSRcolor2[261]);
    BiasedRNG[318] = (LFSRcolor2[37]&LFSRcolor2[207]&LFSRcolor2[150]);
    BiasedRNG[319] = (LFSRcolor2[294]&LFSRcolor2[200]&LFSRcolor2[395]);
    BiasedRNG[320] = (LFSRcolor2[241]&LFSRcolor2[9]&LFSRcolor2[184]);
    BiasedRNG[321] = (LFSRcolor2[208]&LFSRcolor2[236]&LFSRcolor2[279]);
    BiasedRNG[322] = (LFSRcolor2[162]&LFSRcolor2[413]&LFSRcolor2[151]);
    BiasedRNG[323] = (LFSRcolor2[123]&LFSRcolor2[313]&LFSRcolor2[393]);
    BiasedRNG[324] = (LFSRcolor2[319]&LFSRcolor2[309]&LFSRcolor2[250]);
    BiasedRNG[325] = (LFSRcolor2[70]&LFSRcolor2[249]&LFSRcolor2[43]);
    BiasedRNG[326] = (LFSRcolor2[289]&LFSRcolor2[76]&LFSRcolor2[56]);
    BiasedRNG[327] = (LFSRcolor2[156]&LFSRcolor2[107]&LFSRcolor2[126]);
    BiasedRNG[328] = (LFSRcolor2[182]&LFSRcolor2[111]&LFSRcolor2[381]);
    BiasedRNG[329] = (LFSRcolor2[258]&LFSRcolor2[188]&LFSRcolor2[350]);
    BiasedRNG[330] = (LFSRcolor2[186]&LFSRcolor2[297]&LFSRcolor2[167]);
    BiasedRNG[331] = (LFSRcolor2[17]&LFSRcolor2[94]&LFSRcolor2[299]);
    BiasedRNG[332] = (LFSRcolor2[82]&LFSRcolor2[340]&LFSRcolor2[93]);
    BiasedRNG[333] = (LFSRcolor2[185]&LFSRcolor2[259]&LFSRcolor2[337]);
    BiasedRNG[334] = (LFSRcolor2[231]&LFSRcolor2[195]&LFSRcolor2[363]);
    BiasedRNG[335] = (LFSRcolor2[240]&LFSRcolor2[269]&LFSRcolor2[217]);
    BiasedRNG[336] = (LFSRcolor2[20]&LFSRcolor2[328]&LFSRcolor2[140]);
    BiasedRNG[337] = (LFSRcolor2[226]&LFSRcolor2[342]&LFSRcolor2[69]);
    BiasedRNG[338] = (LFSRcolor2[192]&LFSRcolor2[262]&LFSRcolor2[290]);
    UnbiasedRNG[198] = LFSRcolor2[101];
    UnbiasedRNG[199] = LFSRcolor2[44];
    UnbiasedRNG[200] = LFSRcolor2[253];
    UnbiasedRNG[201] = LFSRcolor2[327];
    UnbiasedRNG[202] = LFSRcolor2[145];
    UnbiasedRNG[203] = LFSRcolor2[390];
    UnbiasedRNG[204] = LFSRcolor2[376];
    UnbiasedRNG[205] = LFSRcolor2[27];
    UnbiasedRNG[206] = LFSRcolor2[243];
    UnbiasedRNG[207] = LFSRcolor2[53];
    UnbiasedRNG[208] = LFSRcolor2[143];
    UnbiasedRNG[209] = LFSRcolor2[194];
    UnbiasedRNG[210] = LFSRcolor2[307];
    UnbiasedRNG[211] = LFSRcolor2[136];
    UnbiasedRNG[212] = LFSRcolor2[142];
    UnbiasedRNG[213] = LFSRcolor2[60];
    UnbiasedRNG[214] = LFSRcolor2[354];
    UnbiasedRNG[215] = LFSRcolor2[67];
    UnbiasedRNG[216] = LFSRcolor2[234];
    UnbiasedRNG[217] = LFSRcolor2[301];
    UnbiasedRNG[218] = LFSRcolor2[215];
    UnbiasedRNG[219] = LFSRcolor2[55];
    UnbiasedRNG[220] = LFSRcolor2[36];
    UnbiasedRNG[221] = LFSRcolor2[348];
    UnbiasedRNG[222] = LFSRcolor2[8];
    UnbiasedRNG[223] = LFSRcolor2[46];
    UnbiasedRNG[224] = LFSRcolor2[165];
    UnbiasedRNG[225] = LFSRcolor2[257];
    UnbiasedRNG[226] = LFSRcolor2[318];
    UnbiasedRNG[227] = LFSRcolor2[293];
    UnbiasedRNG[228] = LFSRcolor2[335];
    UnbiasedRNG[229] = LFSRcolor2[218];
    UnbiasedRNG[230] = LFSRcolor2[211];
    UnbiasedRNG[231] = LFSRcolor2[47];
    UnbiasedRNG[232] = LFSRcolor2[298];
    UnbiasedRNG[233] = LFSRcolor2[339];
    UnbiasedRNG[234] = LFSRcolor2[304];
    UnbiasedRNG[235] = LFSRcolor2[368];
    UnbiasedRNG[236] = LFSRcolor2[152];
    UnbiasedRNG[237] = LFSRcolor2[99];
    UnbiasedRNG[238] = LFSRcolor2[346];
    UnbiasedRNG[239] = LFSRcolor2[369];
    UnbiasedRNG[240] = LFSRcolor2[119];
    UnbiasedRNG[241] = LFSRcolor2[281];
    UnbiasedRNG[242] = LFSRcolor2[10];
    UnbiasedRNG[243] = LFSRcolor2[113];
    UnbiasedRNG[244] = LFSRcolor2[370];
    UnbiasedRNG[245] = LFSRcolor2[120];
    UnbiasedRNG[246] = LFSRcolor2[72];
    UnbiasedRNG[247] = LFSRcolor2[22];
    UnbiasedRNG[248] = LFSRcolor2[410];
    UnbiasedRNG[249] = LFSRcolor2[110];
    UnbiasedRNG[250] = LFSRcolor2[157];
    UnbiasedRNG[251] = LFSRcolor2[235];
    UnbiasedRNG[252] = LFSRcolor2[102];
    UnbiasedRNG[253] = LFSRcolor2[66];
    UnbiasedRNG[254] = LFSRcolor2[98];
    UnbiasedRNG[255] = LFSRcolor2[245];
    UnbiasedRNG[256] = LFSRcolor2[306];
    UnbiasedRNG[257] = LFSRcolor2[254];
    UnbiasedRNG[258] = LFSRcolor2[284];
    UnbiasedRNG[259] = LFSRcolor2[326];
    UnbiasedRNG[260] = LFSRcolor2[104];
    UnbiasedRNG[261] = LFSRcolor2[39];
    UnbiasedRNG[262] = LFSRcolor2[345];
    UnbiasedRNG[263] = LFSRcolor2[375];
    UnbiasedRNG[264] = LFSRcolor2[401];
    UnbiasedRNG[265] = LFSRcolor2[382];
    UnbiasedRNG[266] = LFSRcolor2[26];
    UnbiasedRNG[267] = LFSRcolor2[278];
    UnbiasedRNG[268] = LFSRcolor2[334];
    UnbiasedRNG[269] = LFSRcolor2[320];
    UnbiasedRNG[270] = LFSRcolor2[63];
    UnbiasedRNG[271] = LFSRcolor2[21];
    UnbiasedRNG[272] = LFSRcolor2[114];
    UnbiasedRNG[273] = LFSRcolor2[296];
    UnbiasedRNG[274] = LFSRcolor2[360];
    UnbiasedRNG[275] = LFSRcolor2[170];
    UnbiasedRNG[276] = LFSRcolor2[230];
    UnbiasedRNG[277] = LFSRcolor2[372];
    UnbiasedRNG[278] = LFSRcolor2[161];
    UnbiasedRNG[279] = LFSRcolor2[273];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[280] = LFSRcolor3[23];
    UnbiasedRNG[281] = LFSRcolor3[81];
    UnbiasedRNG[282] = LFSRcolor3[48];
    UnbiasedRNG[283] = LFSRcolor3[64];
    UnbiasedRNG[284] = LFSRcolor3[0];
    UnbiasedRNG[285] = LFSRcolor3[38];
    UnbiasedRNG[286] = LFSRcolor3[72];
    UnbiasedRNG[287] = LFSRcolor3[33];
    UnbiasedRNG[288] = LFSRcolor3[78];
    UnbiasedRNG[289] = LFSRcolor3[21];
    UnbiasedRNG[290] = LFSRcolor3[86];
    UnbiasedRNG[291] = LFSRcolor3[44];
    UnbiasedRNG[292] = LFSRcolor3[4];
    UnbiasedRNG[293] = LFSRcolor3[67];
    UnbiasedRNG[294] = LFSRcolor3[47];
    UnbiasedRNG[295] = LFSRcolor3[11];
    UnbiasedRNG[296] = LFSRcolor3[15];
    UnbiasedRNG[297] = LFSRcolor3[2];
    UnbiasedRNG[298] = LFSRcolor3[25];
    UnbiasedRNG[299] = LFSRcolor3[69];
    UnbiasedRNG[300] = LFSRcolor3[32];
    UnbiasedRNG[301] = LFSRcolor3[52];
    UnbiasedRNG[302] = LFSRcolor3[75];
    UnbiasedRNG[303] = LFSRcolor3[24];
    UnbiasedRNG[304] = LFSRcolor3[43];
    UnbiasedRNG[305] = LFSRcolor3[45];
    UnbiasedRNG[306] = LFSRcolor3[20];
    UnbiasedRNG[307] = LFSRcolor3[6];
    UnbiasedRNG[308] = LFSRcolor3[7];
    UnbiasedRNG[309] = LFSRcolor3[68];
    UnbiasedRNG[310] = LFSRcolor3[61];
    UnbiasedRNG[311] = LFSRcolor3[62];
    UnbiasedRNG[312] = LFSRcolor3[90];
    UnbiasedRNG[313] = LFSRcolor3[60];
    UnbiasedRNG[314] = LFSRcolor3[88];
    UnbiasedRNG[315] = LFSRcolor3[42];
    UnbiasedRNG[316] = LFSRcolor3[18];
    UnbiasedRNG[317] = LFSRcolor3[13];
    UnbiasedRNG[318] = LFSRcolor3[79];
    UnbiasedRNG[319] = LFSRcolor3[30];
    UnbiasedRNG[320] = LFSRcolor3[10];
    UnbiasedRNG[321] = LFSRcolor3[91];
    UnbiasedRNG[322] = LFSRcolor3[51];
    UnbiasedRNG[323] = LFSRcolor3[26];
    UnbiasedRNG[324] = LFSRcolor3[49];
    UnbiasedRNG[325] = LFSRcolor3[19];
    UnbiasedRNG[326] = LFSRcolor3[77];
    UnbiasedRNG[327] = LFSRcolor3[71];
    UnbiasedRNG[328] = LFSRcolor3[70];
    UnbiasedRNG[329] = LFSRcolor3[57];
    UnbiasedRNG[330] = LFSRcolor3[37];
    UnbiasedRNG[331] = LFSRcolor3[55];
    UnbiasedRNG[332] = LFSRcolor3[3];
    UnbiasedRNG[333] = LFSRcolor3[1];
    UnbiasedRNG[334] = LFSRcolor3[58];
    UnbiasedRNG[335] = LFSRcolor3[41];
    UnbiasedRNG[336] = LFSRcolor3[89];
    UnbiasedRNG[337] = LFSRcolor3[84];
    UnbiasedRNG[338] = LFSRcolor3[66];
    UnbiasedRNG[339] = LFSRcolor3[9];
    UnbiasedRNG[340] = LFSRcolor3[73];
    UnbiasedRNG[341] = LFSRcolor3[28];
    UnbiasedRNG[342] = LFSRcolor3[16];
    UnbiasedRNG[343] = LFSRcolor3[27];
    UnbiasedRNG[344] = LFSRcolor3[5];
    UnbiasedRNG[345] = LFSRcolor3[40];
    UnbiasedRNG[346] = LFSRcolor3[12];
    UnbiasedRNG[347] = LFSRcolor3[74];
    UnbiasedRNG[348] = LFSRcolor3[8];
    UnbiasedRNG[349] = LFSRcolor3[46];
    UnbiasedRNG[350] = LFSRcolor3[50];
    UnbiasedRNG[351] = LFSRcolor3[39];
end

always @(posedge color3_clk) begin
    BiasedRNG[339] = (LFSRcolor4[85]&LFSRcolor4[249]&LFSRcolor4[112]);
    BiasedRNG[340] = (LFSRcolor4[262]&LFSRcolor4[143]&LFSRcolor4[50]);
    BiasedRNG[341] = (LFSRcolor4[20]&LFSRcolor4[55]&LFSRcolor4[164]);
    BiasedRNG[342] = (LFSRcolor4[5]&LFSRcolor4[82]&LFSRcolor4[225]);
    BiasedRNG[343] = (LFSRcolor4[37]&LFSRcolor4[0]&LFSRcolor4[9]);
    BiasedRNG[344] = (LFSRcolor4[13]&LFSRcolor4[71]&LFSRcolor4[30]);
    BiasedRNG[345] = (LFSRcolor4[116]&LFSRcolor4[270]&LFSRcolor4[107]);
    BiasedRNG[346] = (LFSRcolor4[29]&LFSRcolor4[25]&LFSRcolor4[66]);
    BiasedRNG[347] = (LFSRcolor4[130]&LFSRcolor4[39]&LFSRcolor4[131]);
    BiasedRNG[348] = (LFSRcolor4[192]&LFSRcolor4[264]&LFSRcolor4[90]);
    BiasedRNG[349] = (LFSRcolor4[146]&LFSRcolor4[75]&LFSRcolor4[35]);
    BiasedRNG[350] = (LFSRcolor4[21]&LFSRcolor4[123]&LFSRcolor4[258]);
    BiasedRNG[351] = (LFSRcolor4[149]&LFSRcolor4[6]&LFSRcolor4[273]);
    BiasedRNG[352] = (LFSRcolor4[232]&LFSRcolor4[255]&LFSRcolor4[64]);
    BiasedRNG[353] = (LFSRcolor4[221]&LFSRcolor4[137]&LFSRcolor4[250]);
    BiasedRNG[354] = (LFSRcolor4[34]&LFSRcolor4[119]&LFSRcolor4[22]);
    BiasedRNG[355] = (LFSRcolor4[102]&LFSRcolor4[60]&LFSRcolor4[170]);
    BiasedRNG[356] = (LFSRcolor4[108]&LFSRcolor4[187]&LFSRcolor4[10]);
    BiasedRNG[357] = (LFSRcolor4[172]&LFSRcolor4[125]&LFSRcolor4[114]);
    BiasedRNG[358] = (LFSRcolor4[220]&LFSRcolor4[218]&LFSRcolor4[103]);
    BiasedRNG[359] = (LFSRcolor4[217]&LFSRcolor4[97]&LFSRcolor4[191]);
    BiasedRNG[360] = (LFSRcolor4[152]&LFSRcolor4[62]&LFSRcolor4[223]);
    BiasedRNG[361] = (LFSRcolor4[77]&LFSRcolor4[127]&LFSRcolor4[267]);
    BiasedRNG[362] = (LFSRcolor4[8]&LFSRcolor4[245]&LFSRcolor4[128]);
    BiasedRNG[363] = (LFSRcolor4[28]&LFSRcolor4[42]&LFSRcolor4[195]);
    BiasedRNG[364] = (LFSRcolor4[109]&LFSRcolor4[205]&LFSRcolor4[260]);
    BiasedRNG[365] = (LFSRcolor4[58]&LFSRcolor4[256]&LFSRcolor4[48]);
    BiasedRNG[366] = (LFSRcolor4[158]&LFSRcolor4[185]&LFSRcolor4[84]);
    BiasedRNG[367] = (LFSRcolor4[43]&LFSRcolor4[265]&LFSRcolor4[199]);
    BiasedRNG[368] = (LFSRcolor4[202]&LFSRcolor4[157]&LFSRcolor4[198]);
    BiasedRNG[369] = (LFSRcolor4[165]&LFSRcolor4[117]&LFSRcolor4[38]);
    BiasedRNG[370] = (LFSRcolor4[115]&LFSRcolor4[244]&LFSRcolor4[4]);
    BiasedRNG[371] = (LFSRcolor4[68]&LFSRcolor4[259]&LFSRcolor4[138]);
    BiasedRNG[372] = (LFSRcolor4[175]&LFSRcolor4[161]&LFSRcolor4[257]);
    BiasedRNG[373] = (LFSRcolor4[132]&LFSRcolor4[83]&LFSRcolor4[88]);
    BiasedRNG[374] = (LFSRcolor4[224]&LFSRcolor4[26]&LFSRcolor4[181]);
    BiasedRNG[375] = (LFSRcolor4[200]&LFSRcolor4[144]&LFSRcolor4[126]);
    BiasedRNG[376] = (LFSRcolor4[150]&LFSRcolor4[247]&LFSRcolor4[18]);
    BiasedRNG[377] = (LFSRcolor4[261]&LFSRcolor4[211]&LFSRcolor4[70]);
    BiasedRNG[378] = (LFSRcolor4[275]&LFSRcolor4[141]&LFSRcolor4[101]);
    BiasedRNG[379] = (LFSRcolor4[274]&LFSRcolor4[222]&LFSRcolor4[76]);
    BiasedRNG[380] = (LFSRcolor4[78]&LFSRcolor4[243]&LFSRcolor4[52]);
    BiasedRNG[381] = (LFSRcolor4[167]&LFSRcolor4[7]&LFSRcolor4[73]);
    BiasedRNG[382] = (LFSRcolor4[86]&LFSRcolor4[253]&LFSRcolor4[234]);
    BiasedRNG[383] = (LFSRcolor4[235]&LFSRcolor4[2]&LFSRcolor4[56]);
    BiasedRNG[384] = (LFSRcolor4[136]&LFSRcolor4[227]&LFSRcolor4[230]);
    BiasedRNG[385] = (LFSRcolor4[19]&LFSRcolor4[12]&LFSRcolor4[41]);
    BiasedRNG[386] = (LFSRcolor4[120]&LFSRcolor4[14]&LFSRcolor4[197]);
    BiasedRNG[387] = (LFSRcolor4[184]&LFSRcolor4[155]&LFSRcolor4[129]);
    BiasedRNG[388] = (LFSRcolor4[251]&LFSRcolor4[239]&LFSRcolor4[240]);
    BiasedRNG[389] = (LFSRcolor4[151]&LFSRcolor4[242]&LFSRcolor4[174]);
    BiasedRNG[390] = (LFSRcolor4[163]&LFSRcolor4[148]&LFSRcolor4[254]);
    BiasedRNG[391] = (LFSRcolor4[91]&LFSRcolor4[142]&LFSRcolor4[1]);
    BiasedRNG[392] = (LFSRcolor4[216]&LFSRcolor4[67]&LFSRcolor4[162]);
    BiasedRNG[393] = (LFSRcolor4[237]&LFSRcolor4[15]&LFSRcolor4[47]);
    BiasedRNG[394] = (LFSRcolor4[171]&LFSRcolor4[36]&LFSRcolor4[104]);
    BiasedRNG[395] = (LFSRcolor4[153]&LFSRcolor4[177]&LFSRcolor4[238]);
    BiasedRNG[396] = (LFSRcolor4[229]&LFSRcolor4[210]&LFSRcolor4[252]);
    BiasedRNG[397] = (LFSRcolor4[179]&LFSRcolor4[166]&LFSRcolor4[80]);
    BiasedRNG[398] = (LFSRcolor4[40]&LFSRcolor4[92]&LFSRcolor4[61]);
    BiasedRNG[399] = (LFSRcolor4[140]&LFSRcolor4[215]&LFSRcolor4[32]);
    BiasedRNG[400] = (LFSRcolor4[178]&LFSRcolor4[203]&LFSRcolor4[241]);
    BiasedRNG[401] = (LFSRcolor4[231]&LFSRcolor4[124]&LFSRcolor4[159]);
    BiasedRNG[402] = (LFSRcolor4[113]&LFSRcolor4[118]&LFSRcolor4[269]);
    BiasedRNG[403] = (LFSRcolor4[133]&LFSRcolor4[121]&LFSRcolor4[183]);
    BiasedRNG[404] = (LFSRcolor4[201]&LFSRcolor4[213]&LFSRcolor4[59]);
    BiasedRNG[405] = (LFSRcolor4[111]&LFSRcolor4[79]&LFSRcolor4[95]);
    BiasedRNG[406] = (LFSRcolor4[94]&LFSRcolor4[145]&LFSRcolor4[23]);
    BiasedRNG[407] = (LFSRcolor4[233]&LFSRcolor4[74]&LFSRcolor4[87]);
    BiasedRNG[408] = (LFSRcolor4[147]&LFSRcolor4[173]&LFSRcolor4[176]);
    BiasedRNG[409] = (LFSRcolor4[236]&LFSRcolor4[263]&LFSRcolor4[31]);
    BiasedRNG[410] = (LFSRcolor4[89]&LFSRcolor4[98]&LFSRcolor4[122]);
    BiasedRNG[411] = (LFSRcolor4[196]&LFSRcolor4[190]&LFSRcolor4[63]);
    BiasedRNG[412] = (LFSRcolor4[134]&LFSRcolor4[180]&LFSRcolor4[44]);
    BiasedRNG[413] = (LFSRcolor4[105]&LFSRcolor4[160]&LFSRcolor4[51]);
    BiasedRNG[414] = (LFSRcolor4[188]&LFSRcolor4[106]&LFSRcolor4[208]);
    BiasedRNG[415] = (LFSRcolor4[72]&LFSRcolor4[54]&LFSRcolor4[204]);
    BiasedRNG[416] = (LFSRcolor4[100]&LFSRcolor4[168]&LFSRcolor4[194]);
    BiasedRNG[417] = (LFSRcolor4[65]&LFSRcolor4[182]&LFSRcolor4[214]);
    BiasedRNG[418] = (LFSRcolor4[186]&LFSRcolor4[57]&LFSRcolor4[16]);
    BiasedRNG[419] = (LFSRcolor4[110]&LFSRcolor4[169]&LFSRcolor4[266]);
    BiasedRNG[420] = (LFSRcolor4[11]&LFSRcolor4[156]&LFSRcolor4[268]);
    BiasedRNG[421] = (LFSRcolor4[154]&LFSRcolor4[81]&LFSRcolor4[209]);
    BiasedRNG[422] = (LFSRcolor4[53]&LFSRcolor4[219]&LFSRcolor4[99]);
    BiasedRNG[423] = (LFSRcolor4[139]&LFSRcolor4[33]&LFSRcolor4[135]);
    BiasedRNG[424] = (LFSRcolor4[206]&LFSRcolor4[96]&LFSRcolor4[27]);
    BiasedRNG[425] = (LFSRcolor4[248]&LFSRcolor4[69]&LFSRcolor4[93]);
    BiasedRNG[426] = (LFSRcolor4[212]&LFSRcolor4[17]&LFSRcolor4[228]);
    BiasedRNG[427] = (LFSRcolor4[3]&LFSRcolor4[189]&LFSRcolor4[272]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

//Generate the ILA for data collection:
ila_0 ILAinst(.clk(sample_clk),.probe0(run),.probe1(solution_flag),.probe2(failure),.probe3(counter[37:0]));

//Instantiate VIO:
vio_0 VIOinst (.clk(sample_clk),.probe_out0(reset),.probe_out1(solution_set[19:0]));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule