//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [27:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [1241:0] LFSRcolor0;
wire [1195:0] LFSRcolor1;
wire [965:0] LFSRcolor2;
wire [183:0] LFSRcolor3;
wire [735:0] LFSRcolor4;
reg [879:0] BiasedRNG;       //For I=+/-1 cases
reg [715:0] UnbiasedRNG;   //For I=0 cases
reg [0:1637] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[532] = 1'b1;
initial m[731] = 1'b1;
initial m[741] = 1'b1;
initial m[756] = 1'b0;
initial m[776] = 1'b0;
initial m[801] = 1'b0;
initial m[831] = 1'b1;
initial m[866] = 1'b0;
initial m[906] = 1'b0;
initial m[951] = 1'b1;
initial m[1001] = 1'b0;
initial m[1056] = 1'b0;
initial m[1116] = 1'b0;
initial m[1181] = 1'b1;
initial m[1246] = 1'b0;
initial m[1306] = 1'b0;
initial m[1361] = 1'b0;
initial m[1411] = 1'b1;
initial m[1456] = 1'b1;
initial m[1496] = 1'b1;
initial m[1531] = 1'b0;
initial m[1561] = 1'b0;
initial m[1586] = 1'b1;
initial m[1606] = 1'b1;
initial m[1621] = 1'b1;
initial m[1631] = 1'b1;
initial m[1636] = 1'b1;
initial m[1637] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[730] = 1'b0;
initial m[740] = 1'b0;
initial m[755] = 1'b0;
initial m[775] = 1'b0;
initial m[800] = 1'b0;
initial m[830] = 1'b0;
initial m[865] = 1'b0;
initial m[905] = 1'b0;
initial m[950] = 1'b0;
initial m[1000] = 1'b0;
initial m[1055] = 1'b0;
initial m[1115] = 1'b0;
initial m[1180] = 1'b0;
initial m[1183] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR0_8(.LFSRregister(LFSRcolor0[413:368]),.clk(sample_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR0_9(.LFSRregister(LFSRcolor0[459:414]),.clk(sample_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR0_10(.LFSRregister(LFSRcolor0[505:460]),.clk(sample_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR0_11(.LFSRregister(LFSRcolor0[551:506]),.clk(sample_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR0_12(.LFSRregister(LFSRcolor0[597:552]),.clk(sample_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR0_13(.LFSRregister(LFSRcolor0[643:598]),.clk(sample_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR0_14(.LFSRregister(LFSRcolor0[689:644]),.clk(sample_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR0_15(.LFSRregister(LFSRcolor0[735:690]),.clk(sample_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR0_16(.LFSRregister(LFSRcolor0[781:736]),.clk(sample_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR0_17(.LFSRregister(LFSRcolor0[827:782]),.clk(sample_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR0_18(.LFSRregister(LFSRcolor0[873:828]),.clk(sample_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR0_19(.LFSRregister(LFSRcolor0[919:874]),.clk(sample_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR0_20(.LFSRregister(LFSRcolor0[965:920]),.clk(sample_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR0_21(.LFSRregister(LFSRcolor0[1011:966]),.clk(sample_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR0_22(.LFSRregister(LFSRcolor0[1057:1012]),.clk(sample_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR0_23(.LFSRregister(LFSRcolor0[1103:1058]),.clk(sample_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR0_24(.LFSRregister(LFSRcolor0[1149:1104]),.clk(sample_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR0_25(.LFSRregister(LFSRcolor0[1195:1150]),.clk(sample_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR0_26(.LFSRregister(LFSRcolor0[1241:1196]),.clk(sample_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b0100011100010000010101011001010001111101000000)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b1000101110000100010101010111001111101101001001)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b1100100101010011101001000011100111000000101011)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b1010101011010011100001001101101100110011110011)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0110111001001001100111011011011101101100001101)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b0111010100000100101111101111001010100011110111)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b1010111000011111000010100110001011101010111110)) LFSR1_10(.LFSRregister(LFSRcolor1[505:460]),.clk(color0_clk));
lfsr #(.seed(46'b0111001111101001110000011010001101011011101111)) LFSR1_11(.LFSRregister(LFSRcolor1[551:506]),.clk(color0_clk));
lfsr #(.seed(46'b1001001111101100101100100000101100111110011010)) LFSR1_12(.LFSRregister(LFSRcolor1[597:552]),.clk(color0_clk));
lfsr #(.seed(46'b1001111111100011100000010111111101110010011110)) LFSR1_13(.LFSRregister(LFSRcolor1[643:598]),.clk(color0_clk));
lfsr #(.seed(46'b0000000111011001111111000111110100110000111101)) LFSR1_14(.LFSRregister(LFSRcolor1[689:644]),.clk(color0_clk));
lfsr #(.seed(46'b0100000011011100110101110101010010111001010000)) LFSR1_15(.LFSRregister(LFSRcolor1[735:690]),.clk(color0_clk));
lfsr #(.seed(46'b1010010111011000101010101111011000010011001010)) LFSR1_16(.LFSRregister(LFSRcolor1[781:736]),.clk(color0_clk));
lfsr #(.seed(46'b1011010100011001010110010011101110100011101010)) LFSR1_17(.LFSRregister(LFSRcolor1[827:782]),.clk(color0_clk));
lfsr #(.seed(46'b0111011011101111010101001100011100100100110000)) LFSR1_18(.LFSRregister(LFSRcolor1[873:828]),.clk(color0_clk));
lfsr #(.seed(46'b1110110011110011000100010100111110011101010011)) LFSR1_19(.LFSRregister(LFSRcolor1[919:874]),.clk(color0_clk));
lfsr #(.seed(46'b0011001000010001001111001110101111011111000110)) LFSR1_20(.LFSRregister(LFSRcolor1[965:920]),.clk(color0_clk));
lfsr #(.seed(46'b0101000110100000010101001000010000101101100110)) LFSR1_21(.LFSRregister(LFSRcolor1[1011:966]),.clk(color0_clk));
lfsr #(.seed(46'b1110011010010011001010111010100101111111100000)) LFSR1_22(.LFSRregister(LFSRcolor1[1057:1012]),.clk(color0_clk));
lfsr #(.seed(46'b1001111000010100100001100010110000001111101011)) LFSR1_23(.LFSRregister(LFSRcolor1[1103:1058]),.clk(color0_clk));
lfsr #(.seed(46'b0011101001111100110111000000010000101100111110)) LFSR1_24(.LFSRregister(LFSRcolor1[1149:1104]),.clk(color0_clk));
lfsr #(.seed(46'b1010111010001100001100010110010011100100101100)) LFSR1_25(.LFSRregister(LFSRcolor1[1195:1150]),.clk(color0_clk));
lfsr #(.seed(46'b1101010000110001000001011010110100010000110101)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0111111000001001010001100011001110110101101001)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b0111011110101100100001111000001001111001010010)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b0110010001011011111100000000110011011110000100)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b1100101101001001110010011101110000001110111111)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b1110010100000011100111110011000001001000000101)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b1100111110111110000101110101010111111010101000)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b1101101000110111001110111111011011100011111101)) LFSR2_7(.LFSRregister(LFSRcolor2[367:322]),.clk(color1_clk));
lfsr #(.seed(46'b1011100111101011110000001101111100001111100011)) LFSR2_8(.LFSRregister(LFSRcolor2[413:368]),.clk(color1_clk));
lfsr #(.seed(46'b1000011101010100110111010000000111000111010111)) LFSR2_9(.LFSRregister(LFSRcolor2[459:414]),.clk(color1_clk));
lfsr #(.seed(46'b0011001001101100101110110001011100100100110000)) LFSR2_10(.LFSRregister(LFSRcolor2[505:460]),.clk(color1_clk));
lfsr #(.seed(46'b0011110010011101000111111110100110110100101000)) LFSR2_11(.LFSRregister(LFSRcolor2[551:506]),.clk(color1_clk));
lfsr #(.seed(46'b1100000100011100010111001011000000101100110100)) LFSR2_12(.LFSRregister(LFSRcolor2[597:552]),.clk(color1_clk));
lfsr #(.seed(46'b1001101001101101001001111001110100110001100010)) LFSR2_13(.LFSRregister(LFSRcolor2[643:598]),.clk(color1_clk));
lfsr #(.seed(46'b1000000000001101011011010100000001101001001111)) LFSR2_14(.LFSRregister(LFSRcolor2[689:644]),.clk(color1_clk));
lfsr #(.seed(46'b1000011000100000010011100100110100001010000001)) LFSR2_15(.LFSRregister(LFSRcolor2[735:690]),.clk(color1_clk));
lfsr #(.seed(46'b0101000011110010010110011011111101010101011010)) LFSR2_16(.LFSRregister(LFSRcolor2[781:736]),.clk(color1_clk));
lfsr #(.seed(46'b0011111001110010110000110100101000000000100010)) LFSR2_17(.LFSRregister(LFSRcolor2[827:782]),.clk(color1_clk));
lfsr #(.seed(46'b0011101001110100101101111100101010101100110000)) LFSR2_18(.LFSRregister(LFSRcolor2[873:828]),.clk(color1_clk));
lfsr #(.seed(46'b1100111100001111010111011100011110001010110011)) LFSR2_19(.LFSRregister(LFSRcolor2[919:874]),.clk(color1_clk));
lfsr #(.seed(46'b0101101111111000101111101010111101100011110011)) LFSR2_20(.LFSRregister(LFSRcolor2[965:920]),.clk(color1_clk));
lfsr #(.seed(46'b1100101101101111100100111011110111010010100100)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b0110001110010011010100101010010010100100011000)) LFSR3_1(.LFSRregister(LFSRcolor3[91:46]),.clk(color2_clk));
lfsr #(.seed(46'b0010101111101011001110100001110011000100001001)) LFSR3_2(.LFSRregister(LFSRcolor3[137:92]),.clk(color2_clk));
lfsr #(.seed(46'b0100110100101000110001000110101010001110100101)) LFSR3_3(.LFSRregister(LFSRcolor3[183:138]),.clk(color2_clk));
lfsr #(.seed(46'b1111010011010001011111110011011111011111011010)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b0011000010001101011100101011111101010001010111)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b0011010011011000100111011100010000001110001110)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0010110000011111111111101000111101111100101000)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b1110000110010010100110000110010000011111100110)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));
lfsr #(.seed(46'b0011101100010010111110000100001011000110001101)) LFSR4_5(.LFSRregister(LFSRcolor4[275:230]),.clk(color3_clk));
lfsr #(.seed(46'b0010001010111001000011110110110110100001001011)) LFSR4_6(.LFSRregister(LFSRcolor4[321:276]),.clk(color3_clk));
lfsr #(.seed(46'b1010111110010100100000100111111111101010101011)) LFSR4_7(.LFSRregister(LFSRcolor4[367:322]),.clk(color3_clk));
lfsr #(.seed(46'b0000001101010010101110010000001110111100000000)) LFSR4_8(.LFSRregister(LFSRcolor4[413:368]),.clk(color3_clk));
lfsr #(.seed(46'b0001101011110001101001101001111111011101001010)) LFSR4_9(.LFSRregister(LFSRcolor4[459:414]),.clk(color3_clk));
lfsr #(.seed(46'b1010111010011010101000111010001000010011110111)) LFSR4_10(.LFSRregister(LFSRcolor4[505:460]),.clk(color3_clk));
lfsr #(.seed(46'b0001100101111110101010111111100101111000000011)) LFSR4_11(.LFSRregister(LFSRcolor4[551:506]),.clk(color3_clk));
lfsr #(.seed(46'b1110110011101111100000001011100011010010100101)) LFSR4_12(.LFSRregister(LFSRcolor4[597:552]),.clk(color3_clk));
lfsr #(.seed(46'b1110101011011010101011001110110110100100110110)) LFSR4_13(.LFSRregister(LFSRcolor4[643:598]),.clk(color3_clk));
lfsr #(.seed(46'b0011111111100000000000011101001000101110111011)) LFSR4_14(.LFSRregister(LFSRcolor4[689:644]),.clk(color3_clk));
lfsr #(.seed(46'b0111111111000000001010100101100111000000010111)) LFSR4_15(.LFSRregister(LFSRcolor4[735:690]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 0;
initial m[1] = 0;
initial m[2] = 1;
initial m[3] = 0;
initial m[4] = 1;
initial m[5] = 1;
initial m[6] = 1;
initial m[7] = 0;
initial m[8] = 0;
initial m[9] = 0;
initial m[10] = 1;
initial m[11] = 1;
initial m[12] = 0;
initial m[13] = 0;
initial m[14] = 1;
initial m[15] = 0;
initial m[16] = 0;
initial m[17] = 0;
initial m[18] = 0;
initial m[19] = 0;
initial m[20] = 0;
initial m[21] = 0;
initial m[22] = 1;
initial m[23] = 1;
initial m[24] = 0;
initial m[25] = 1;
initial m[26] = 0;
initial m[27] = 0;
initial m[28] = 0;
initial m[29] = 1;
initial m[30] = 1;
initial m[31] = 0;
initial m[32] = 1;
initial m[33] = 1;
initial m[34] = 0;
initial m[35] = 0;
initial m[36] = 1;
initial m[37] = 1;
initial m[38] = 0;
initial m[39] = 1;
initial m[40] = 0;
initial m[41] = 0;
initial m[42] = 0;
initial m[43] = 0;
initial m[44] = 0;
initial m[45] = 0;
initial m[46] = 1;
initial m[47] = 1;
initial m[48] = 0;
initial m[49] = 1;
initial m[50] = 1;
initial m[51] = 0;
initial m[52] = 1;
initial m[53] = 0;
initial m[54] = 1;
initial m[55] = 1;
initial m[56] = 0;
initial m[57] = 0;
initial m[58] = 0;
initial m[59] = 1;
initial m[60] = 1;
initial m[61] = 0;
initial m[62] = 1;
initial m[63] = 1;
initial m[64] = 1;
initial m[65] = 1;
initial m[66] = 0;
initial m[67] = 0;
initial m[68] = 1;
initial m[69] = 0;
initial m[70] = 1;
initial m[71] = 0;
initial m[72] = 0;
initial m[73] = 1;
initial m[74] = 1;
initial m[75] = 0;
initial m[76] = 0;
initial m[77] = 0;
initial m[78] = 1;
initial m[79] = 1;
initial m[80] = 0;
initial m[81] = 1;
initial m[82] = 0;
initial m[83] = 1;
initial m[84] = 0;
initial m[85] = 0;
initial m[86] = 1;
initial m[87] = 1;
initial m[88] = 1;
initial m[89] = 0;
initial m[90] = 0;
initial m[91] = 1;
initial m[92] = 1;
initial m[93] = 1;
initial m[94] = 1;
initial m[95] = 1;
initial m[96] = 0;
initial m[97] = 1;
initial m[98] = 1;
initial m[99] = 1;
initial m[100] = 1;
initial m[101] = 1;
initial m[102] = 0;
initial m[103] = 1;
initial m[104] = 0;
initial m[105] = 0;
initial m[106] = 0;
initial m[107] = 0;
initial m[108] = 0;
initial m[109] = 1;
initial m[110] = 1;
initial m[111] = 0;
initial m[112] = 1;
initial m[113] = 1;
initial m[114] = 0;
initial m[115] = 1;
initial m[116] = 0;
initial m[117] = 1;
initial m[118] = 1;
initial m[119] = 0;
initial m[120] = 1;
initial m[121] = 1;
initial m[122] = 0;
initial m[123] = 0;
initial m[124] = 0;
initial m[125] = 0;
initial m[126] = 0;
initial m[127] = 1;
initial m[128] = 1;
initial m[129] = 1;
initial m[130] = 0;
initial m[131] = 0;
initial m[132] = 0;
initial m[133] = 0;
initial m[134] = 1;
initial m[135] = 0;
initial m[136] = 0;
initial m[137] = 1;
initial m[138] = 1;
initial m[139] = 1;
initial m[140] = 1;
initial m[141] = 1;
initial m[142] = 1;
initial m[143] = 0;
initial m[144] = 1;
initial m[145] = 0;
initial m[146] = 1;
initial m[147] = 1;
initial m[148] = 0;
initial m[149] = 0;
initial m[150] = 0;
initial m[151] = 0;
initial m[152] = 0;
initial m[153] = 1;
initial m[154] = 0;
initial m[155] = 1;
initial m[156] = 0;
initial m[157] = 1;
initial m[158] = 0;
initial m[159] = 1;
initial m[160] = 1;
initial m[161] = 1;
initial m[162] = 1;
initial m[163] = 1;
initial m[164] = 0;
initial m[165] = 1;
initial m[166] = 1;
initial m[167] = 1;
initial m[168] = 1;
initial m[169] = 1;
initial m[170] = 0;
initial m[171] = 0;
initial m[172] = 0;
initial m[173] = 1;
initial m[174] = 0;
initial m[175] = 0;
initial m[176] = 1;
initial m[177] = 0;
initial m[178] = 1;
initial m[179] = 1;
initial m[180] = 0;
initial m[181] = 0;
initial m[182] = 1;
initial m[183] = 1;
initial m[184] = 0;
initial m[185] = 1;
initial m[186] = 0;
initial m[187] = 1;
initial m[188] = 1;
initial m[189] = 0;
initial m[190] = 0;
initial m[191] = 1;
initial m[192] = 0;
initial m[193] = 1;
initial m[194] = 1;
initial m[195] = 1;
initial m[196] = 0;
initial m[197] = 0;
initial m[198] = 0;
initial m[199] = 1;
initial m[200] = 0;
initial m[201] = 0;
initial m[202] = 1;
initial m[203] = 0;
initial m[204] = 0;
initial m[205] = 1;
initial m[206] = 0;
initial m[207] = 0;
initial m[208] = 1;
initial m[209] = 1;
initial m[210] = 0;
initial m[211] = 1;
initial m[212] = 0;
initial m[213] = 1;
initial m[214] = 1;
initial m[215] = 1;
initial m[216] = 1;
initial m[217] = 0;
initial m[218] = 1;
initial m[219] = 1;
initial m[220] = 1;
initial m[221] = 0;
initial m[222] = 0;
initial m[223] = 1;
initial m[224] = 0;
initial m[225] = 1;
initial m[226] = 0;
initial m[227] = 0;
initial m[228] = 1;
initial m[229] = 0;
initial m[230] = 1;
initial m[231] = 1;
initial m[232] = 0;
initial m[233] = 1;
initial m[234] = 1;
initial m[235] = 0;
initial m[236] = 1;
initial m[237] = 0;
initial m[238] = 0;
initial m[239] = 1;
initial m[240] = 1;
initial m[241] = 1;
initial m[242] = 1;
initial m[243] = 0;
initial m[244] = 1;
initial m[245] = 0;
initial m[246] = 0;
initial m[247] = 0;
initial m[248] = 0;
initial m[249] = 0;
initial m[250] = 1;
initial m[251] = 0;
initial m[252] = 0;
initial m[253] = 1;
initial m[254] = 0;
initial m[255] = 0;
initial m[256] = 1;
initial m[257] = 0;
initial m[258] = 0;
initial m[259] = 0;
initial m[260] = 0;
initial m[261] = 1;
initial m[262] = 0;
initial m[263] = 0;
initial m[264] = 1;
initial m[265] = 1;
initial m[266] = 1;
initial m[267] = 1;
initial m[268] = 1;
initial m[269] = 0;
initial m[270] = 0;
initial m[271] = 1;
initial m[272] = 0;
initial m[273] = 0;
initial m[274] = 0;
initial m[275] = 1;
initial m[276] = 1;
initial m[277] = 1;
initial m[278] = 1;
initial m[279] = 1;
initial m[280] = 0;
initial m[281] = 0;
initial m[282] = 0;
initial m[283] = 0;
initial m[284] = 0;
initial m[285] = 0;
initial m[286] = 1;
initial m[287] = 0;
initial m[288] = 1;
initial m[289] = 1;
initial m[290] = 0;
initial m[291] = 0;
initial m[292] = 1;
initial m[293] = 0;
initial m[294] = 1;
initial m[295] = 1;
initial m[296] = 0;
initial m[297] = 1;
initial m[298] = 0;
initial m[299] = 1;
initial m[300] = 1;
initial m[301] = 0;
initial m[302] = 1;
initial m[303] = 0;
initial m[304] = 0;
initial m[305] = 1;
initial m[306] = 1;
initial m[307] = 1;
initial m[308] = 1;
initial m[309] = 0;
initial m[310] = 0;
initial m[311] = 0;
initial m[312] = 0;
initial m[313] = 1;
initial m[314] = 0;
initial m[315] = 0;
initial m[316] = 1;
initial m[317] = 1;
initial m[318] = 0;
initial m[319] = 0;
initial m[320] = 1;
initial m[321] = 1;
initial m[322] = 1;
initial m[323] = 1;
initial m[324] = 0;
initial m[325] = 1;
initial m[326] = 0;
initial m[327] = 1;
initial m[328] = 0;
initial m[329] = 1;
initial m[330] = 0;
initial m[331] = 1;
initial m[332] = 1;
initial m[333] = 1;
initial m[334] = 1;
initial m[335] = 1;
initial m[336] = 1;
initial m[337] = 1;
initial m[338] = 0;
initial m[339] = 1;
initial m[340] = 1;
initial m[341] = 1;
initial m[342] = 0;
initial m[343] = 0;
initial m[344] = 0;
initial m[345] = 1;
initial m[346] = 1;
initial m[347] = 0;
initial m[348] = 0;
initial m[349] = 1;
initial m[350] = 1;
initial m[351] = 1;
initial m[352] = 0;
initial m[353] = 1;
initial m[354] = 0;
initial m[355] = 1;
initial m[356] = 1;
initial m[357] = 0;
initial m[358] = 0;
initial m[359] = 1;
initial m[360] = 1;
initial m[361] = 0;
initial m[362] = 1;
initial m[363] = 1;
initial m[364] = 1;
initial m[365] = 0;
initial m[366] = 0;
initial m[367] = 1;
initial m[368] = 1;
initial m[369] = 0;
initial m[370] = 0;
initial m[371] = 0;
initial m[372] = 0;
initial m[373] = 1;
initial m[374] = 1;
initial m[375] = 1;
initial m[376] = 1;
initial m[377] = 1;
initial m[378] = 1;
initial m[379] = 0;
initial m[380] = 0;
initial m[381] = 1;
initial m[382] = 0;
initial m[383] = 0;
initial m[384] = 1;
initial m[385] = 0;
initial m[386] = 1;
initial m[387] = 0;
initial m[388] = 1;
initial m[389] = 1;
initial m[390] = 0;
initial m[391] = 1;
initial m[392] = 1;
initial m[393] = 0;
initial m[394] = 1;
initial m[395] = 1;
initial m[396] = 1;
initial m[397] = 1;
initial m[398] = 1;
initial m[399] = 0;
initial m[400] = 0;
initial m[401] = 0;
initial m[402] = 0;
initial m[403] = 0;
initial m[404] = 1;
initial m[405] = 1;
initial m[406] = 0;
initial m[407] = 0;
initial m[408] = 0;
initial m[409] = 0;
initial m[410] = 0;
initial m[411] = 0;
initial m[412] = 1;
initial m[413] = 1;
initial m[414] = 1;
initial m[415] = 0;
initial m[416] = 1;
initial m[417] = 1;
initial m[418] = 0;
initial m[419] = 0;
initial m[420] = 1;
initial m[421] = 1;
initial m[422] = 0;
initial m[423] = 0;
initial m[424] = 0;
initial m[425] = 1;
initial m[426] = 0;
initial m[427] = 1;
initial m[428] = 1;
initial m[429] = 0;
initial m[430] = 1;
initial m[431] = 0;
initial m[432] = 1;
initial m[433] = 1;
initial m[434] = 0;
initial m[435] = 0;
initial m[436] = 0;
initial m[437] = 0;
initial m[438] = 0;
initial m[439] = 1;
initial m[440] = 1;
initial m[441] = 1;
initial m[442] = 0;
initial m[443] = 1;
initial m[444] = 1;
initial m[445] = 1;
initial m[446] = 1;
initial m[447] = 1;
initial m[448] = 1;
initial m[449] = 0;
initial m[450] = 1;
initial m[451] = 0;
initial m[452] = 0;
initial m[453] = 0;
initial m[454] = 0;
initial m[455] = 1;
initial m[456] = 0;
initial m[457] = 1;
initial m[458] = 0;
initial m[459] = 0;
initial m[460] = 0;
initial m[461] = 1;
initial m[462] = 0;
initial m[463] = 0;
initial m[464] = 1;
initial m[465] = 1;
initial m[466] = 1;
initial m[467] = 1;
initial m[468] = 1;
initial m[469] = 1;
initial m[470] = 0;
initial m[471] = 0;
initial m[472] = 0;
initial m[473] = 1;
initial m[474] = 0;
initial m[475] = 1;
initial m[476] = 0;
initial m[477] = 1;
initial m[478] = 1;
initial m[479] = 0;
initial m[480] = 1;
initial m[481] = 1;
initial m[482] = 1;
initial m[483] = 1;
initial m[484] = 1;
initial m[485] = 1;
initial m[486] = 0;
initial m[487] = 0;
initial m[488] = 1;
initial m[489] = 0;
initial m[490] = 0;
initial m[491] = 1;
initial m[492] = 1;
initial m[493] = 0;
initial m[494] = 1;
initial m[495] = 0;
initial m[496] = 0;
initial m[497] = 0;
initial m[498] = 0;
initial m[499] = 1;
initial m[500] = 0;
initial m[501] = 1;
initial m[502] = 0;
initial m[503] = 0;
initial m[504] = 1;
initial m[505] = 0;
initial m[506] = 1;
initial m[507] = 0;
initial m[508] = 0;
initial m[509] = 0;
initial m[510] = 1;
initial m[511] = 1;
initial m[512] = 1;
initial m[513] = 0;
initial m[514] = 1;
initial m[515] = 0;
initial m[516] = 0;
initial m[517] = 0;
initial m[518] = 1;
initial m[519] = 0;
initial m[520] = 1;
initial m[521] = 0;
initial m[522] = 0;
initial m[523] = 0;
initial m[524] = 0;
initial m[525] = 0;
initial m[526] = 1;
initial m[527] = 1;
initial m[528] = 1;
initial m[529] = 1;
initial m[530] = 0;
initial m[531] = 0;
initial m[533] = 0;
initial m[534] = 1;
initial m[535] = 1;
initial m[536] = 0;
initial m[537] = 0;
initial m[538] = 1;
initial m[539] = 1;
initial m[540] = 1;
initial m[541] = 1;
initial m[542] = 1;
initial m[543] = 0;
initial m[544] = 1;
initial m[545] = 0;
initial m[546] = 0;
initial m[547] = 1;
initial m[548] = 1;
initial m[549] = 0;
initial m[550] = 1;
initial m[551] = 1;
initial m[552] = 0;
initial m[553] = 1;
initial m[554] = 1;
initial m[555] = 0;
initial m[556] = 0;
initial m[557] = 0;
initial m[558] = 0;
initial m[559] = 0;
initial m[560] = 1;
initial m[561] = 0;
initial m[562] = 0;
initial m[563] = 1;
initial m[564] = 1;
initial m[565] = 1;
initial m[566] = 0;
initial m[567] = 1;
initial m[568] = 1;
initial m[569] = 0;
initial m[570] = 1;
initial m[571] = 0;
initial m[572] = 1;
initial m[573] = 0;
initial m[574] = 1;
initial m[575] = 0;
initial m[576] = 1;
initial m[577] = 0;
initial m[578] = 1;
initial m[579] = 0;
initial m[580] = 0;
initial m[581] = 0;
initial m[582] = 1;
initial m[583] = 1;
initial m[584] = 0;
initial m[585] = 1;
initial m[586] = 0;
initial m[587] = 0;
initial m[588] = 1;
initial m[589] = 0;
initial m[590] = 0;
initial m[591] = 1;
initial m[592] = 1;
initial m[593] = 0;
initial m[594] = 1;
initial m[595] = 0;
initial m[596] = 0;
initial m[597] = 0;
initial m[598] = 0;
initial m[599] = 0;
initial m[600] = 1;
initial m[601] = 0;
initial m[602] = 1;
initial m[603] = 0;
initial m[604] = 1;
initial m[605] = 0;
initial m[606] = 1;
initial m[607] = 1;
initial m[608] = 0;
initial m[609] = 0;
initial m[610] = 0;
initial m[611] = 1;
initial m[612] = 0;
initial m[613] = 1;
initial m[614] = 1;
initial m[615] = 1;
initial m[616] = 1;
initial m[617] = 0;
initial m[618] = 1;
initial m[619] = 0;
initial m[620] = 0;
initial m[621] = 0;
initial m[622] = 0;
initial m[623] = 1;
initial m[624] = 0;
initial m[625] = 1;
initial m[626] = 0;
initial m[627] = 1;
initial m[628] = 1;
initial m[629] = 0;
initial m[630] = 1;
initial m[631] = 1;
initial m[632] = 1;
initial m[633] = 0;
initial m[634] = 0;
initial m[635] = 0;
initial m[636] = 0;
initial m[637] = 1;
initial m[638] = 1;
initial m[639] = 0;
initial m[640] = 0;
initial m[641] = 0;
initial m[642] = 1;
initial m[643] = 1;
initial m[644] = 0;
initial m[645] = 0;
initial m[646] = 1;
initial m[647] = 1;
initial m[648] = 0;
initial m[649] = 1;
initial m[650] = 0;
initial m[651] = 0;
initial m[652] = 1;
initial m[653] = 1;
initial m[654] = 0;
initial m[655] = 1;
initial m[656] = 0;
initial m[657] = 0;
initial m[658] = 0;
initial m[659] = 1;
initial m[660] = 0;
initial m[661] = 1;
initial m[662] = 1;
initial m[663] = 1;
initial m[664] = 0;
initial m[665] = 0;
initial m[666] = 0;
initial m[667] = 1;
initial m[668] = 0;
initial m[669] = 1;
initial m[670] = 0;
initial m[671] = 0;
initial m[672] = 0;
initial m[673] = 1;
initial m[674] = 0;
initial m[675] = 0;
initial m[676] = 0;
initial m[677] = 1;
initial m[678] = 0;
initial m[679] = 1;
initial m[680] = 1;
initial m[681] = 0;
initial m[682] = 0;
initial m[683] = 1;
initial m[684] = 1;
initial m[685] = 0;
initial m[686] = 0;
initial m[687] = 1;
initial m[688] = 0;
initial m[689] = 1;
initial m[690] = 0;
initial m[691] = 1;
initial m[692] = 1;
initial m[693] = 0;
initial m[694] = 1;
initial m[695] = 1;
initial m[696] = 0;
initial m[697] = 1;
initial m[698] = 0;
initial m[699] = 1;
initial m[700] = 1;
initial m[701] = 0;
initial m[702] = 0;
initial m[703] = 0;
initial m[704] = 1;
initial m[705] = 1;
initial m[706] = 1;
initial m[707] = 1;
initial m[708] = 1;
initial m[709] = 0;
initial m[710] = 1;
initial m[711] = 1;
initial m[712] = 1;
initial m[713] = 1;
initial m[714] = 0;
initial m[715] = 0;
initial m[716] = 1;
initial m[717] = 0;
initial m[718] = 0;
initial m[719] = 1;
initial m[720] = 0;
initial m[721] = 1;
initial m[722] = 0;
initial m[723] = 0;
initial m[724] = 1;
initial m[725] = 0;
initial m[726] = 0;
initial m[727] = 1;
initial m[728] = 0;
initial m[729] = 0;
initial m[732] = 0;
initial m[733] = 0;
initial m[734] = 0;
initial m[735] = 1;
initial m[736] = 0;
initial m[737] = 0;
initial m[738] = 0;
initial m[739] = 0;
initial m[742] = 1;
initial m[743] = 0;
initial m[744] = 0;
initial m[745] = 1;
initial m[746] = 0;
initial m[747] = 1;
initial m[748] = 0;
initial m[749] = 1;
initial m[750] = 0;
initial m[751] = 1;
initial m[752] = 0;
initial m[753] = 1;
initial m[754] = 1;
initial m[757] = 1;
initial m[758] = 1;
initial m[759] = 1;
initial m[760] = 1;
initial m[761] = 1;
initial m[762] = 1;
initial m[763] = 1;
initial m[764] = 0;
initial m[765] = 0;
initial m[766] = 0;
initial m[767] = 1;
initial m[768] = 1;
initial m[769] = 1;
initial m[770] = 1;
initial m[771] = 1;
initial m[772] = 0;
initial m[773] = 0;
initial m[774] = 1;
initial m[777] = 0;
initial m[778] = 0;
initial m[779] = 1;
initial m[780] = 0;
initial m[781] = 0;
initial m[782] = 1;
initial m[783] = 0;
initial m[784] = 0;
initial m[785] = 0;
initial m[786] = 0;
initial m[787] = 0;
initial m[788] = 0;
initial m[789] = 1;
initial m[790] = 0;
initial m[791] = 0;
initial m[792] = 0;
initial m[793] = 0;
initial m[794] = 0;
initial m[795] = 0;
initial m[796] = 0;
initial m[797] = 1;
initial m[798] = 0;
initial m[799] = 1;
initial m[802] = 1;
initial m[803] = 0;
initial m[804] = 0;
initial m[805] = 1;
initial m[806] = 1;
initial m[807] = 1;
initial m[808] = 1;
initial m[809] = 1;
initial m[810] = 0;
initial m[811] = 0;
initial m[812] = 0;
initial m[813] = 1;
initial m[814] = 1;
initial m[815] = 1;
initial m[816] = 0;
initial m[817] = 0;
initial m[818] = 1;
initial m[819] = 0;
initial m[820] = 1;
initial m[821] = 1;
initial m[822] = 1;
initial m[823] = 1;
initial m[824] = 1;
initial m[825] = 1;
initial m[826] = 0;
initial m[827] = 0;
initial m[828] = 1;
initial m[829] = 1;
initial m[832] = 1;
initial m[833] = 1;
initial m[834] = 1;
initial m[835] = 1;
initial m[836] = 1;
initial m[837] = 0;
initial m[838] = 0;
initial m[839] = 1;
initial m[840] = 1;
initial m[841] = 0;
initial m[842] = 0;
initial m[843] = 0;
initial m[844] = 0;
initial m[845] = 0;
initial m[846] = 1;
initial m[847] = 1;
initial m[848] = 0;
initial m[849] = 0;
initial m[850] = 1;
initial m[851] = 0;
initial m[852] = 1;
initial m[853] = 1;
initial m[854] = 0;
initial m[855] = 0;
initial m[856] = 0;
initial m[857] = 0;
initial m[858] = 0;
initial m[859] = 1;
initial m[860] = 1;
initial m[861] = 0;
initial m[862] = 0;
initial m[863] = 0;
initial m[864] = 0;
initial m[867] = 1;
initial m[868] = 0;
initial m[869] = 1;
initial m[870] = 1;
initial m[871] = 0;
initial m[872] = 0;
initial m[873] = 1;
initial m[874] = 1;
initial m[875] = 1;
initial m[876] = 1;
initial m[877] = 0;
initial m[878] = 1;
initial m[879] = 1;
initial m[880] = 0;
initial m[881] = 1;
initial m[882] = 0;
initial m[883] = 1;
initial m[884] = 1;
initial m[885] = 0;
initial m[886] = 0;
initial m[887] = 0;
initial m[888] = 0;
initial m[889] = 0;
initial m[890] = 0;
initial m[891] = 1;
initial m[892] = 1;
initial m[893] = 0;
initial m[894] = 1;
initial m[895] = 0;
initial m[896] = 0;
initial m[897] = 0;
initial m[898] = 1;
initial m[899] = 1;
initial m[900] = 0;
initial m[901] = 1;
initial m[902] = 0;
initial m[903] = 0;
initial m[904] = 0;
initial m[907] = 0;
initial m[908] = 1;
initial m[909] = 1;
initial m[910] = 0;
initial m[911] = 1;
initial m[912] = 1;
initial m[913] = 1;
initial m[914] = 0;
initial m[915] = 1;
initial m[916] = 1;
initial m[917] = 0;
initial m[918] = 1;
initial m[919] = 0;
initial m[920] = 0;
initial m[921] = 1;
initial m[922] = 1;
initial m[923] = 0;
initial m[924] = 0;
initial m[925] = 0;
initial m[926] = 0;
initial m[927] = 0;
initial m[928] = 1;
initial m[929] = 1;
initial m[930] = 1;
initial m[931] = 1;
initial m[932] = 1;
initial m[933] = 0;
initial m[934] = 0;
initial m[935] = 0;
initial m[936] = 1;
initial m[937] = 1;
initial m[938] = 1;
initial m[939] = 1;
initial m[940] = 0;
initial m[941] = 1;
initial m[942] = 0;
initial m[943] = 1;
initial m[944] = 0;
initial m[945] = 1;
initial m[946] = 0;
initial m[947] = 0;
initial m[948] = 1;
initial m[949] = 0;
initial m[952] = 0;
initial m[953] = 0;
initial m[954] = 1;
initial m[955] = 0;
initial m[956] = 1;
initial m[957] = 0;
initial m[958] = 1;
initial m[959] = 1;
initial m[960] = 1;
initial m[961] = 1;
initial m[962] = 0;
initial m[963] = 0;
initial m[964] = 1;
initial m[965] = 0;
initial m[966] = 0;
initial m[967] = 1;
initial m[968] = 0;
initial m[969] = 0;
initial m[970] = 0;
initial m[971] = 1;
initial m[972] = 1;
initial m[973] = 1;
initial m[974] = 1;
initial m[975] = 0;
initial m[976] = 0;
initial m[977] = 0;
initial m[978] = 1;
initial m[979] = 1;
initial m[980] = 1;
initial m[981] = 0;
initial m[982] = 1;
initial m[983] = 1;
initial m[984] = 1;
initial m[985] = 0;
initial m[986] = 0;
initial m[987] = 0;
initial m[988] = 0;
initial m[989] = 1;
initial m[990] = 0;
initial m[991] = 1;
initial m[992] = 0;
initial m[993] = 0;
initial m[994] = 1;
initial m[995] = 0;
initial m[996] = 1;
initial m[997] = 0;
initial m[998] = 1;
initial m[999] = 1;
initial m[1002] = 1;
initial m[1003] = 1;
initial m[1004] = 1;
initial m[1005] = 0;
initial m[1006] = 0;
initial m[1007] = 0;
initial m[1008] = 0;
initial m[1009] = 0;
initial m[1010] = 1;
initial m[1011] = 0;
initial m[1012] = 0;
initial m[1013] = 1;
initial m[1014] = 1;
initial m[1015] = 1;
initial m[1016] = 1;
initial m[1017] = 0;
initial m[1018] = 0;
initial m[1019] = 0;
initial m[1020] = 0;
initial m[1021] = 1;
initial m[1022] = 1;
initial m[1023] = 0;
initial m[1024] = 1;
initial m[1025] = 1;
initial m[1026] = 1;
initial m[1027] = 1;
initial m[1028] = 0;
initial m[1029] = 1;
initial m[1030] = 0;
initial m[1031] = 1;
initial m[1032] = 1;
initial m[1033] = 0;
initial m[1034] = 0;
initial m[1035] = 0;
initial m[1036] = 0;
initial m[1037] = 0;
initial m[1038] = 1;
initial m[1039] = 1;
initial m[1040] = 1;
initial m[1041] = 1;
initial m[1042] = 0;
initial m[1043] = 0;
initial m[1044] = 0;
initial m[1045] = 1;
initial m[1046] = 0;
initial m[1047] = 1;
initial m[1048] = 1;
initial m[1049] = 0;
initial m[1050] = 1;
initial m[1051] = 1;
initial m[1052] = 0;
initial m[1053] = 0;
initial m[1054] = 0;
initial m[1057] = 0;
initial m[1058] = 1;
initial m[1059] = 0;
initial m[1060] = 0;
initial m[1061] = 1;
initial m[1062] = 0;
initial m[1063] = 1;
initial m[1064] = 0;
initial m[1065] = 1;
initial m[1066] = 1;
initial m[1067] = 0;
initial m[1068] = 1;
initial m[1069] = 1;
initial m[1070] = 0;
initial m[1071] = 1;
initial m[1072] = 0;
initial m[1073] = 0;
initial m[1074] = 1;
initial m[1075] = 1;
initial m[1076] = 0;
initial m[1077] = 0;
initial m[1078] = 1;
initial m[1079] = 0;
initial m[1080] = 0;
initial m[1081] = 0;
initial m[1082] = 0;
initial m[1083] = 1;
initial m[1084] = 1;
initial m[1085] = 1;
initial m[1086] = 1;
initial m[1087] = 0;
initial m[1088] = 0;
initial m[1089] = 1;
initial m[1090] = 0;
initial m[1091] = 1;
initial m[1092] = 0;
initial m[1093] = 1;
initial m[1094] = 1;
initial m[1095] = 0;
initial m[1096] = 1;
initial m[1097] = 1;
initial m[1098] = 1;
initial m[1099] = 1;
initial m[1100] = 0;
initial m[1101] = 0;
initial m[1102] = 1;
initial m[1103] = 0;
initial m[1104] = 0;
initial m[1105] = 0;
initial m[1106] = 0;
initial m[1107] = 0;
initial m[1108] = 0;
initial m[1109] = 0;
initial m[1110] = 1;
initial m[1111] = 1;
initial m[1112] = 1;
initial m[1113] = 1;
initial m[1114] = 0;
initial m[1117] = 0;
initial m[1118] = 0;
initial m[1119] = 0;
initial m[1120] = 1;
initial m[1121] = 1;
initial m[1122] = 1;
initial m[1123] = 1;
initial m[1124] = 1;
initial m[1125] = 0;
initial m[1126] = 1;
initial m[1127] = 1;
initial m[1128] = 0;
initial m[1129] = 0;
initial m[1130] = 0;
initial m[1131] = 0;
initial m[1132] = 1;
initial m[1133] = 0;
initial m[1134] = 1;
initial m[1135] = 1;
initial m[1136] = 1;
initial m[1137] = 1;
initial m[1138] = 0;
initial m[1139] = 0;
initial m[1140] = 0;
initial m[1141] = 1;
initial m[1142] = 0;
initial m[1143] = 1;
initial m[1144] = 0;
initial m[1145] = 0;
initial m[1146] = 1;
initial m[1147] = 1;
initial m[1148] = 0;
initial m[1149] = 1;
initial m[1150] = 1;
initial m[1151] = 0;
initial m[1152] = 1;
initial m[1153] = 0;
initial m[1154] = 0;
initial m[1155] = 0;
initial m[1156] = 1;
initial m[1157] = 0;
initial m[1158] = 1;
initial m[1159] = 0;
initial m[1160] = 0;
initial m[1161] = 1;
initial m[1162] = 1;
initial m[1163] = 1;
initial m[1164] = 0;
initial m[1165] = 0;
initial m[1166] = 0;
initial m[1167] = 0;
initial m[1168] = 1;
initial m[1169] = 1;
initial m[1170] = 0;
initial m[1171] = 0;
initial m[1172] = 1;
initial m[1173] = 1;
initial m[1174] = 1;
initial m[1175] = 0;
initial m[1176] = 0;
initial m[1177] = 1;
initial m[1178] = 0;
initial m[1179] = 0;
initial m[1182] = 1;
initial m[1184] = 1;
initial m[1185] = 0;
initial m[1186] = 0;
initial m[1187] = 1;
initial m[1188] = 1;
initial m[1189] = 0;
initial m[1190] = 1;
initial m[1191] = 0;
initial m[1192] = 1;
initial m[1193] = 0;
initial m[1194] = 0;
initial m[1195] = 0;
initial m[1196] = 1;
initial m[1197] = 0;
initial m[1198] = 0;
initial m[1199] = 0;
initial m[1200] = 1;
initial m[1201] = 0;
initial m[1202] = 1;
initial m[1203] = 0;
initial m[1204] = 0;
initial m[1205] = 1;
initial m[1206] = 0;
initial m[1207] = 0;
initial m[1208] = 1;
initial m[1209] = 0;
initial m[1210] = 1;
initial m[1211] = 0;
initial m[1212] = 1;
initial m[1213] = 0;
initial m[1214] = 1;
initial m[1215] = 0;
initial m[1216] = 1;
initial m[1217] = 0;
initial m[1218] = 1;
initial m[1219] = 1;
initial m[1220] = 0;
initial m[1221] = 0;
initial m[1222] = 0;
initial m[1223] = 0;
initial m[1224] = 1;
initial m[1225] = 0;
initial m[1226] = 1;
initial m[1227] = 0;
initial m[1228] = 0;
initial m[1229] = 0;
initial m[1230] = 1;
initial m[1231] = 0;
initial m[1232] = 1;
initial m[1233] = 1;
initial m[1234] = 0;
initial m[1235] = 0;
initial m[1236] = 1;
initial m[1237] = 1;
initial m[1238] = 1;
initial m[1239] = 0;
initial m[1240] = 0;
initial m[1241] = 0;
initial m[1242] = 1;
initial m[1243] = 1;
initial m[1244] = 1;
initial m[1245] = 0;
initial m[1247] = 1;
initial m[1248] = 1;
initial m[1249] = 0;
initial m[1250] = 0;
initial m[1251] = 1;
initial m[1252] = 0;
initial m[1253] = 0;
initial m[1254] = 0;
initial m[1255] = 0;
initial m[1256] = 0;
initial m[1257] = 1;
initial m[1258] = 0;
initial m[1259] = 1;
initial m[1260] = 0;
initial m[1261] = 0;
initial m[1262] = 0;
initial m[1263] = 1;
initial m[1264] = 1;
initial m[1265] = 0;
initial m[1266] = 1;
initial m[1267] = 1;
initial m[1268] = 0;
initial m[1269] = 0;
initial m[1270] = 0;
initial m[1271] = 1;
initial m[1272] = 0;
initial m[1273] = 0;
initial m[1274] = 1;
initial m[1275] = 1;
initial m[1276] = 0;
initial m[1277] = 1;
initial m[1278] = 0;
initial m[1279] = 1;
initial m[1280] = 0;
initial m[1281] = 0;
initial m[1282] = 1;
initial m[1283] = 1;
initial m[1284] = 1;
initial m[1285] = 1;
initial m[1286] = 0;
initial m[1287] = 1;
initial m[1288] = 0;
initial m[1289] = 0;
initial m[1290] = 0;
initial m[1291] = 1;
initial m[1292] = 1;
initial m[1293] = 1;
initial m[1294] = 1;
initial m[1295] = 0;
initial m[1296] = 1;
initial m[1297] = 0;
initial m[1298] = 0;
initial m[1299] = 0;
initial m[1300] = 1;
initial m[1301] = 0;
initial m[1302] = 1;
initial m[1303] = 1;
initial m[1304] = 0;
initial m[1305] = 0;
initial m[1307] = 1;
initial m[1308] = 1;
initial m[1309] = 0;
initial m[1310] = 0;
initial m[1311] = 1;
initial m[1312] = 1;
initial m[1313] = 1;
initial m[1314] = 0;
initial m[1315] = 0;
initial m[1316] = 0;
initial m[1317] = 1;
initial m[1318] = 1;
initial m[1319] = 1;
initial m[1320] = 1;
initial m[1321] = 0;
initial m[1322] = 0;
initial m[1323] = 0;
initial m[1324] = 0;
initial m[1325] = 0;
initial m[1326] = 0;
initial m[1327] = 1;
initial m[1328] = 0;
initial m[1329] = 1;
initial m[1330] = 1;
initial m[1331] = 0;
initial m[1332] = 0;
initial m[1333] = 0;
initial m[1334] = 1;
initial m[1335] = 0;
initial m[1336] = 1;
initial m[1337] = 1;
initial m[1338] = 1;
initial m[1339] = 1;
initial m[1340] = 1;
initial m[1341] = 1;
initial m[1342] = 1;
initial m[1343] = 1;
initial m[1344] = 0;
initial m[1345] = 0;
initial m[1346] = 1;
initial m[1347] = 0;
initial m[1348] = 1;
initial m[1349] = 1;
initial m[1350] = 1;
initial m[1351] = 1;
initial m[1352] = 1;
initial m[1353] = 1;
initial m[1354] = 1;
initial m[1355] = 1;
initial m[1356] = 0;
initial m[1357] = 1;
initial m[1358] = 0;
initial m[1359] = 1;
initial m[1360] = 1;
initial m[1362] = 1;
initial m[1363] = 1;
initial m[1364] = 0;
initial m[1365] = 1;
initial m[1366] = 1;
initial m[1367] = 0;
initial m[1368] = 1;
initial m[1369] = 0;
initial m[1370] = 0;
initial m[1371] = 0;
initial m[1372] = 0;
initial m[1373] = 1;
initial m[1374] = 1;
initial m[1375] = 1;
initial m[1376] = 1;
initial m[1377] = 1;
initial m[1378] = 0;
initial m[1379] = 1;
initial m[1380] = 1;
initial m[1381] = 1;
initial m[1382] = 1;
initial m[1383] = 1;
initial m[1384] = 1;
initial m[1385] = 1;
initial m[1386] = 1;
initial m[1387] = 1;
initial m[1388] = 0;
initial m[1389] = 1;
initial m[1390] = 0;
initial m[1391] = 1;
initial m[1392] = 1;
initial m[1393] = 1;
initial m[1394] = 0;
initial m[1395] = 0;
initial m[1396] = 0;
initial m[1397] = 0;
initial m[1398] = 1;
initial m[1399] = 1;
initial m[1400] = 1;
initial m[1401] = 1;
initial m[1402] = 0;
initial m[1403] = 0;
initial m[1404] = 0;
initial m[1405] = 1;
initial m[1406] = 1;
initial m[1407] = 0;
initial m[1408] = 0;
initial m[1409] = 1;
initial m[1410] = 0;
initial m[1412] = 1;
initial m[1413] = 1;
initial m[1414] = 1;
initial m[1415] = 0;
initial m[1416] = 0;
initial m[1417] = 1;
initial m[1418] = 0;
initial m[1419] = 1;
initial m[1420] = 0;
initial m[1421] = 1;
initial m[1422] = 0;
initial m[1423] = 1;
initial m[1424] = 1;
initial m[1425] = 1;
initial m[1426] = 0;
initial m[1427] = 0;
initial m[1428] = 1;
initial m[1429] = 0;
initial m[1430] = 0;
initial m[1431] = 0;
initial m[1432] = 1;
initial m[1433] = 1;
initial m[1434] = 0;
initial m[1435] = 1;
initial m[1436] = 1;
initial m[1437] = 1;
initial m[1438] = 0;
initial m[1439] = 1;
initial m[1440] = 0;
initial m[1441] = 1;
initial m[1442] = 1;
initial m[1443] = 1;
initial m[1444] = 0;
initial m[1445] = 0;
initial m[1446] = 0;
initial m[1447] = 0;
initial m[1448] = 0;
initial m[1449] = 1;
initial m[1450] = 1;
initial m[1451] = 1;
initial m[1452] = 0;
initial m[1453] = 0;
initial m[1454] = 1;
initial m[1455] = 0;
initial m[1457] = 1;
initial m[1458] = 0;
initial m[1459] = 1;
initial m[1460] = 1;
initial m[1461] = 0;
initial m[1462] = 1;
initial m[1463] = 1;
initial m[1464] = 1;
initial m[1465] = 0;
initial m[1466] = 1;
initial m[1467] = 1;
initial m[1468] = 1;
initial m[1469] = 1;
initial m[1470] = 1;
initial m[1471] = 0;
initial m[1472] = 0;
initial m[1473] = 0;
initial m[1474] = 0;
initial m[1475] = 0;
initial m[1476] = 1;
initial m[1477] = 0;
initial m[1478] = 0;
initial m[1479] = 1;
initial m[1480] = 1;
initial m[1481] = 0;
initial m[1482] = 1;
initial m[1483] = 0;
initial m[1484] = 1;
initial m[1485] = 0;
initial m[1486] = 1;
initial m[1487] = 1;
initial m[1488] = 1;
initial m[1489] = 0;
initial m[1490] = 0;
initial m[1491] = 0;
initial m[1492] = 1;
initial m[1493] = 0;
initial m[1494] = 0;
initial m[1495] = 1;
initial m[1497] = 1;
initial m[1498] = 1;
initial m[1499] = 1;
initial m[1500] = 0;
initial m[1501] = 1;
initial m[1502] = 0;
initial m[1503] = 1;
initial m[1504] = 0;
initial m[1505] = 1;
initial m[1506] = 1;
initial m[1507] = 0;
initial m[1508] = 1;
initial m[1509] = 1;
initial m[1510] = 0;
initial m[1511] = 0;
initial m[1512] = 1;
initial m[1513] = 1;
initial m[1514] = 1;
initial m[1515] = 1;
initial m[1516] = 1;
initial m[1517] = 0;
initial m[1518] = 0;
initial m[1519] = 0;
initial m[1520] = 1;
initial m[1521] = 1;
initial m[1522] = 1;
initial m[1523] = 1;
initial m[1524] = 0;
initial m[1525] = 0;
initial m[1526] = 0;
initial m[1527] = 1;
initial m[1528] = 1;
initial m[1529] = 1;
initial m[1530] = 1;
initial m[1532] = 0;
initial m[1533] = 1;
initial m[1534] = 0;
initial m[1535] = 1;
initial m[1536] = 0;
initial m[1537] = 0;
initial m[1538] = 0;
initial m[1539] = 1;
initial m[1540] = 1;
initial m[1541] = 1;
initial m[1542] = 1;
initial m[1543] = 1;
initial m[1544] = 1;
initial m[1545] = 0;
initial m[1546] = 0;
initial m[1547] = 1;
initial m[1548] = 1;
initial m[1549] = 0;
initial m[1550] = 0;
initial m[1551] = 1;
initial m[1552] = 1;
initial m[1553] = 1;
initial m[1554] = 0;
initial m[1555] = 0;
initial m[1556] = 0;
initial m[1557] = 1;
initial m[1558] = 1;
initial m[1559] = 1;
initial m[1560] = 1;
initial m[1562] = 0;
initial m[1563] = 1;
initial m[1564] = 1;
initial m[1565] = 0;
initial m[1566] = 1;
initial m[1567] = 0;
initial m[1568] = 1;
initial m[1569] = 1;
initial m[1570] = 1;
initial m[1571] = 0;
initial m[1572] = 1;
initial m[1573] = 1;
initial m[1574] = 0;
initial m[1575] = 1;
initial m[1576] = 1;
initial m[1577] = 0;
initial m[1578] = 0;
initial m[1579] = 1;
initial m[1580] = 1;
initial m[1581] = 0;
initial m[1582] = 1;
initial m[1583] = 0;
initial m[1584] = 1;
initial m[1585] = 1;
initial m[1587] = 0;
initial m[1588] = 0;
initial m[1589] = 1;
initial m[1590] = 1;
initial m[1591] = 0;
initial m[1592] = 1;
initial m[1593] = 1;
initial m[1594] = 1;
initial m[1595] = 0;
initial m[1596] = 1;
initial m[1597] = 0;
initial m[1598] = 0;
initial m[1599] = 0;
initial m[1600] = 0;
initial m[1601] = 1;
initial m[1602] = 0;
initial m[1603] = 0;
initial m[1604] = 0;
initial m[1605] = 0;
initial m[1607] = 0;
initial m[1608] = 1;
initial m[1609] = 0;
initial m[1610] = 0;
initial m[1611] = 0;
initial m[1612] = 0;
initial m[1613] = 0;
initial m[1614] = 1;
initial m[1615] = 0;
initial m[1616] = 0;
initial m[1617] = 1;
initial m[1618] = 0;
initial m[1619] = 1;
initial m[1620] = 0;
initial m[1622] = 1;
initial m[1623] = 0;
initial m[1624] = 0;
initial m[1625] = 1;
initial m[1626] = 1;
initial m[1627] = 1;
initial m[1628] = 0;
initial m[1629] = 1;
initial m[1630] = 0;
initial m[1632] = 1;
initial m[1633] = 1;
initial m[1634] = 1;
initial m[1635] = 0;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[13],m[12],m[11],m[10],m[9],m[8],m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[27],m[26],m[25],m[24],m[23],m[22],m[21],m[20],m[19],m[18],m[17],m[16],m[15],m[14]};
end

always @(negedge sample_clk) begin
    if (solution == 28'b1111110011100010001001000111)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[28]&~m[56])|(~m[28]&m[56]))&UnbiasedRNG[0])|((m[28]&m[56]));
    m[1] = (((m[29]&~m[59])|(~m[29]&m[59]))&UnbiasedRNG[1])|((m[29]&m[59]));
    m[2] = (((m[30]&~m[62])|(~m[30]&m[62]))&UnbiasedRNG[2])|((m[30]&m[62]));
    m[3] = (((m[31]&~m[65])|(~m[31]&m[65]))&UnbiasedRNG[3])|((m[31]&m[65]));
    m[4] = (((m[32]&~m[68])|(~m[32]&m[68]))&UnbiasedRNG[4])|((m[32]&m[68]));
    m[5] = (((m[33]&~m[71])|(~m[33]&m[71]))&UnbiasedRNG[5])|((m[33]&m[71]));
    m[6] = (((m[34]&~m[74])|(~m[34]&m[74]))&UnbiasedRNG[6])|((m[34]&m[74]));
    m[7] = (((m[35]&~m[77])|(~m[35]&m[77]))&UnbiasedRNG[7])|((m[35]&m[77]));
    m[8] = (((m[36]&~m[80])|(~m[36]&m[80]))&UnbiasedRNG[8])|((m[36]&m[80]));
    m[9] = (((m[37]&~m[83])|(~m[37]&m[83]))&UnbiasedRNG[9])|((m[37]&m[83]));
    m[10] = (((m[38]&~m[86])|(~m[38]&m[86]))&UnbiasedRNG[10])|((m[38]&m[86]));
    m[11] = (((m[39]&~m[89])|(~m[39]&m[89]))&UnbiasedRNG[11])|((m[39]&m[89]));
    m[12] = (((m[40]&~m[92])|(~m[40]&m[92]))&UnbiasedRNG[12])|((m[40]&m[92]));
    m[13] = (((m[41]&~m[95])|(~m[41]&m[95]))&UnbiasedRNG[13])|((m[41]&m[95]));
    m[14] = (((m[42]&~m[98])|(~m[42]&m[98]))&UnbiasedRNG[14])|((m[42]&m[98]));
    m[15] = (((m[43]&~m[101])|(~m[43]&m[101]))&UnbiasedRNG[15])|((m[43]&m[101]));
    m[16] = (((m[44]&~m[104])|(~m[44]&m[104]))&UnbiasedRNG[16])|((m[44]&m[104]));
    m[17] = (((m[45]&~m[107])|(~m[45]&m[107]))&UnbiasedRNG[17])|((m[45]&m[107]));
    m[18] = (((m[46]&~m[110])|(~m[46]&m[110]))&UnbiasedRNG[18])|((m[46]&m[110]));
    m[19] = (((m[47]&~m[113])|(~m[47]&m[113]))&UnbiasedRNG[19])|((m[47]&m[113]));
    m[20] = (((m[48]&~m[116])|(~m[48]&m[116]))&UnbiasedRNG[20])|((m[48]&m[116]));
    m[21] = (((m[49]&~m[119])|(~m[49]&m[119]))&UnbiasedRNG[21])|((m[49]&m[119]));
    m[22] = (((m[50]&~m[122])|(~m[50]&m[122]))&UnbiasedRNG[22])|((m[50]&m[122]));
    m[23] = (((m[51]&~m[125])|(~m[51]&m[125]))&UnbiasedRNG[23])|((m[51]&m[125]));
    m[24] = (((m[52]&~m[128])|(~m[52]&m[128]))&UnbiasedRNG[24])|((m[52]&m[128]));
    m[25] = (((m[53]&~m[131])|(~m[53]&m[131]))&UnbiasedRNG[25])|((m[53]&m[131]));
    m[26] = (((m[54]&~m[134])|(~m[54]&m[134]))&UnbiasedRNG[26])|((m[54]&m[134]));
    m[27] = (((m[55]&~m[137])|(~m[55]&m[137]))&UnbiasedRNG[27])|((m[55]&m[137]));
    m[57] = (((m[28]&m[146]&~m[147]&~m[148]&~m[149])|(m[28]&~m[146]&m[147]&~m[148]&~m[149])|(~m[28]&m[146]&m[147]&~m[148]&~m[149])|(m[28]&~m[146]&~m[147]&m[148]&~m[149])|(~m[28]&m[146]&~m[147]&m[148]&~m[149])|(~m[28]&~m[146]&m[147]&m[148]&~m[149])|(m[28]&~m[146]&~m[147]&~m[148]&m[149])|(~m[28]&m[146]&~m[147]&~m[148]&m[149])|(~m[28]&~m[146]&m[147]&~m[148]&m[149])|(~m[28]&~m[146]&~m[147]&m[148]&m[149]))&BiasedRNG[0])|(((m[28]&m[146]&m[147]&~m[148]&~m[149])|(m[28]&m[146]&~m[147]&m[148]&~m[149])|(m[28]&~m[146]&m[147]&m[148]&~m[149])|(~m[28]&m[146]&m[147]&m[148]&~m[149])|(m[28]&m[146]&~m[147]&~m[148]&m[149])|(m[28]&~m[146]&m[147]&~m[148]&m[149])|(~m[28]&m[146]&m[147]&~m[148]&m[149])|(m[28]&~m[146]&~m[147]&m[148]&m[149])|(~m[28]&m[146]&~m[147]&m[148]&m[149])|(~m[28]&~m[146]&m[147]&m[148]&m[149]))&~BiasedRNG[0])|((m[28]&m[146]&m[147]&m[148]&~m[149])|(m[28]&m[146]&m[147]&~m[148]&m[149])|(m[28]&m[146]&~m[147]&m[148]&m[149])|(m[28]&~m[146]&m[147]&m[148]&m[149])|(~m[28]&m[146]&m[147]&m[148]&m[149])|(m[28]&m[146]&m[147]&m[148]&m[149]));
    m[58] = (((m[28]&m[150]&~m[151]&~m[152]&~m[153])|(m[28]&~m[150]&m[151]&~m[152]&~m[153])|(~m[28]&m[150]&m[151]&~m[152]&~m[153])|(m[28]&~m[150]&~m[151]&m[152]&~m[153])|(~m[28]&m[150]&~m[151]&m[152]&~m[153])|(~m[28]&~m[150]&m[151]&m[152]&~m[153])|(m[28]&~m[150]&~m[151]&~m[152]&m[153])|(~m[28]&m[150]&~m[151]&~m[152]&m[153])|(~m[28]&~m[150]&m[151]&~m[152]&m[153])|(~m[28]&~m[150]&~m[151]&m[152]&m[153]))&BiasedRNG[1])|(((m[28]&m[150]&m[151]&~m[152]&~m[153])|(m[28]&m[150]&~m[151]&m[152]&~m[153])|(m[28]&~m[150]&m[151]&m[152]&~m[153])|(~m[28]&m[150]&m[151]&m[152]&~m[153])|(m[28]&m[150]&~m[151]&~m[152]&m[153])|(m[28]&~m[150]&m[151]&~m[152]&m[153])|(~m[28]&m[150]&m[151]&~m[152]&m[153])|(m[28]&~m[150]&~m[151]&m[152]&m[153])|(~m[28]&m[150]&~m[151]&m[152]&m[153])|(~m[28]&~m[150]&m[151]&m[152]&m[153]))&~BiasedRNG[1])|((m[28]&m[150]&m[151]&m[152]&~m[153])|(m[28]&m[150]&m[151]&~m[152]&m[153])|(m[28]&m[150]&~m[151]&m[152]&m[153])|(m[28]&~m[150]&m[151]&m[152]&m[153])|(~m[28]&m[150]&m[151]&m[152]&m[153])|(m[28]&m[150]&m[151]&m[152]&m[153]));
    m[60] = (((m[29]&m[160]&~m[161]&~m[162]&~m[163])|(m[29]&~m[160]&m[161]&~m[162]&~m[163])|(~m[29]&m[160]&m[161]&~m[162]&~m[163])|(m[29]&~m[160]&~m[161]&m[162]&~m[163])|(~m[29]&m[160]&~m[161]&m[162]&~m[163])|(~m[29]&~m[160]&m[161]&m[162]&~m[163])|(m[29]&~m[160]&~m[161]&~m[162]&m[163])|(~m[29]&m[160]&~m[161]&~m[162]&m[163])|(~m[29]&~m[160]&m[161]&~m[162]&m[163])|(~m[29]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[2])|(((m[29]&m[160]&m[161]&~m[162]&~m[163])|(m[29]&m[160]&~m[161]&m[162]&~m[163])|(m[29]&~m[160]&m[161]&m[162]&~m[163])|(~m[29]&m[160]&m[161]&m[162]&~m[163])|(m[29]&m[160]&~m[161]&~m[162]&m[163])|(m[29]&~m[160]&m[161]&~m[162]&m[163])|(~m[29]&m[160]&m[161]&~m[162]&m[163])|(m[29]&~m[160]&~m[161]&m[162]&m[163])|(~m[29]&m[160]&~m[161]&m[162]&m[163])|(~m[29]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[2])|((m[29]&m[160]&m[161]&m[162]&~m[163])|(m[29]&m[160]&m[161]&~m[162]&m[163])|(m[29]&m[160]&~m[161]&m[162]&m[163])|(m[29]&~m[160]&m[161]&m[162]&m[163])|(~m[29]&m[160]&m[161]&m[162]&m[163])|(m[29]&m[160]&m[161]&m[162]&m[163]));
    m[61] = (((m[29]&m[164]&~m[165]&~m[166]&~m[167])|(m[29]&~m[164]&m[165]&~m[166]&~m[167])|(~m[29]&m[164]&m[165]&~m[166]&~m[167])|(m[29]&~m[164]&~m[165]&m[166]&~m[167])|(~m[29]&m[164]&~m[165]&m[166]&~m[167])|(~m[29]&~m[164]&m[165]&m[166]&~m[167])|(m[29]&~m[164]&~m[165]&~m[166]&m[167])|(~m[29]&m[164]&~m[165]&~m[166]&m[167])|(~m[29]&~m[164]&m[165]&~m[166]&m[167])|(~m[29]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[3])|(((m[29]&m[164]&m[165]&~m[166]&~m[167])|(m[29]&m[164]&~m[165]&m[166]&~m[167])|(m[29]&~m[164]&m[165]&m[166]&~m[167])|(~m[29]&m[164]&m[165]&m[166]&~m[167])|(m[29]&m[164]&~m[165]&~m[166]&m[167])|(m[29]&~m[164]&m[165]&~m[166]&m[167])|(~m[29]&m[164]&m[165]&~m[166]&m[167])|(m[29]&~m[164]&~m[165]&m[166]&m[167])|(~m[29]&m[164]&~m[165]&m[166]&m[167])|(~m[29]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[3])|((m[29]&m[164]&m[165]&m[166]&~m[167])|(m[29]&m[164]&m[165]&~m[166]&m[167])|(m[29]&m[164]&~m[165]&m[166]&m[167])|(m[29]&~m[164]&m[165]&m[166]&m[167])|(~m[29]&m[164]&m[165]&m[166]&m[167])|(m[29]&m[164]&m[165]&m[166]&m[167]));
    m[63] = (((m[30]&m[174]&~m[175]&~m[176]&~m[177])|(m[30]&~m[174]&m[175]&~m[176]&~m[177])|(~m[30]&m[174]&m[175]&~m[176]&~m[177])|(m[30]&~m[174]&~m[175]&m[176]&~m[177])|(~m[30]&m[174]&~m[175]&m[176]&~m[177])|(~m[30]&~m[174]&m[175]&m[176]&~m[177])|(m[30]&~m[174]&~m[175]&~m[176]&m[177])|(~m[30]&m[174]&~m[175]&~m[176]&m[177])|(~m[30]&~m[174]&m[175]&~m[176]&m[177])|(~m[30]&~m[174]&~m[175]&m[176]&m[177]))&BiasedRNG[4])|(((m[30]&m[174]&m[175]&~m[176]&~m[177])|(m[30]&m[174]&~m[175]&m[176]&~m[177])|(m[30]&~m[174]&m[175]&m[176]&~m[177])|(~m[30]&m[174]&m[175]&m[176]&~m[177])|(m[30]&m[174]&~m[175]&~m[176]&m[177])|(m[30]&~m[174]&m[175]&~m[176]&m[177])|(~m[30]&m[174]&m[175]&~m[176]&m[177])|(m[30]&~m[174]&~m[175]&m[176]&m[177])|(~m[30]&m[174]&~m[175]&m[176]&m[177])|(~m[30]&~m[174]&m[175]&m[176]&m[177]))&~BiasedRNG[4])|((m[30]&m[174]&m[175]&m[176]&~m[177])|(m[30]&m[174]&m[175]&~m[176]&m[177])|(m[30]&m[174]&~m[175]&m[176]&m[177])|(m[30]&~m[174]&m[175]&m[176]&m[177])|(~m[30]&m[174]&m[175]&m[176]&m[177])|(m[30]&m[174]&m[175]&m[176]&m[177]));
    m[64] = (((m[30]&m[178]&~m[179]&~m[180]&~m[181])|(m[30]&~m[178]&m[179]&~m[180]&~m[181])|(~m[30]&m[178]&m[179]&~m[180]&~m[181])|(m[30]&~m[178]&~m[179]&m[180]&~m[181])|(~m[30]&m[178]&~m[179]&m[180]&~m[181])|(~m[30]&~m[178]&m[179]&m[180]&~m[181])|(m[30]&~m[178]&~m[179]&~m[180]&m[181])|(~m[30]&m[178]&~m[179]&~m[180]&m[181])|(~m[30]&~m[178]&m[179]&~m[180]&m[181])|(~m[30]&~m[178]&~m[179]&m[180]&m[181]))&BiasedRNG[5])|(((m[30]&m[178]&m[179]&~m[180]&~m[181])|(m[30]&m[178]&~m[179]&m[180]&~m[181])|(m[30]&~m[178]&m[179]&m[180]&~m[181])|(~m[30]&m[178]&m[179]&m[180]&~m[181])|(m[30]&m[178]&~m[179]&~m[180]&m[181])|(m[30]&~m[178]&m[179]&~m[180]&m[181])|(~m[30]&m[178]&m[179]&~m[180]&m[181])|(m[30]&~m[178]&~m[179]&m[180]&m[181])|(~m[30]&m[178]&~m[179]&m[180]&m[181])|(~m[30]&~m[178]&m[179]&m[180]&m[181]))&~BiasedRNG[5])|((m[30]&m[178]&m[179]&m[180]&~m[181])|(m[30]&m[178]&m[179]&~m[180]&m[181])|(m[30]&m[178]&~m[179]&m[180]&m[181])|(m[30]&~m[178]&m[179]&m[180]&m[181])|(~m[30]&m[178]&m[179]&m[180]&m[181])|(m[30]&m[178]&m[179]&m[180]&m[181]));
    m[66] = (((m[31]&m[188]&~m[189]&~m[190]&~m[191])|(m[31]&~m[188]&m[189]&~m[190]&~m[191])|(~m[31]&m[188]&m[189]&~m[190]&~m[191])|(m[31]&~m[188]&~m[189]&m[190]&~m[191])|(~m[31]&m[188]&~m[189]&m[190]&~m[191])|(~m[31]&~m[188]&m[189]&m[190]&~m[191])|(m[31]&~m[188]&~m[189]&~m[190]&m[191])|(~m[31]&m[188]&~m[189]&~m[190]&m[191])|(~m[31]&~m[188]&m[189]&~m[190]&m[191])|(~m[31]&~m[188]&~m[189]&m[190]&m[191]))&BiasedRNG[6])|(((m[31]&m[188]&m[189]&~m[190]&~m[191])|(m[31]&m[188]&~m[189]&m[190]&~m[191])|(m[31]&~m[188]&m[189]&m[190]&~m[191])|(~m[31]&m[188]&m[189]&m[190]&~m[191])|(m[31]&m[188]&~m[189]&~m[190]&m[191])|(m[31]&~m[188]&m[189]&~m[190]&m[191])|(~m[31]&m[188]&m[189]&~m[190]&m[191])|(m[31]&~m[188]&~m[189]&m[190]&m[191])|(~m[31]&m[188]&~m[189]&m[190]&m[191])|(~m[31]&~m[188]&m[189]&m[190]&m[191]))&~BiasedRNG[6])|((m[31]&m[188]&m[189]&m[190]&~m[191])|(m[31]&m[188]&m[189]&~m[190]&m[191])|(m[31]&m[188]&~m[189]&m[190]&m[191])|(m[31]&~m[188]&m[189]&m[190]&m[191])|(~m[31]&m[188]&m[189]&m[190]&m[191])|(m[31]&m[188]&m[189]&m[190]&m[191]));
    m[67] = (((m[31]&m[192]&~m[193]&~m[194]&~m[195])|(m[31]&~m[192]&m[193]&~m[194]&~m[195])|(~m[31]&m[192]&m[193]&~m[194]&~m[195])|(m[31]&~m[192]&~m[193]&m[194]&~m[195])|(~m[31]&m[192]&~m[193]&m[194]&~m[195])|(~m[31]&~m[192]&m[193]&m[194]&~m[195])|(m[31]&~m[192]&~m[193]&~m[194]&m[195])|(~m[31]&m[192]&~m[193]&~m[194]&m[195])|(~m[31]&~m[192]&m[193]&~m[194]&m[195])|(~m[31]&~m[192]&~m[193]&m[194]&m[195]))&BiasedRNG[7])|(((m[31]&m[192]&m[193]&~m[194]&~m[195])|(m[31]&m[192]&~m[193]&m[194]&~m[195])|(m[31]&~m[192]&m[193]&m[194]&~m[195])|(~m[31]&m[192]&m[193]&m[194]&~m[195])|(m[31]&m[192]&~m[193]&~m[194]&m[195])|(m[31]&~m[192]&m[193]&~m[194]&m[195])|(~m[31]&m[192]&m[193]&~m[194]&m[195])|(m[31]&~m[192]&~m[193]&m[194]&m[195])|(~m[31]&m[192]&~m[193]&m[194]&m[195])|(~m[31]&~m[192]&m[193]&m[194]&m[195]))&~BiasedRNG[7])|((m[31]&m[192]&m[193]&m[194]&~m[195])|(m[31]&m[192]&m[193]&~m[194]&m[195])|(m[31]&m[192]&~m[193]&m[194]&m[195])|(m[31]&~m[192]&m[193]&m[194]&m[195])|(~m[31]&m[192]&m[193]&m[194]&m[195])|(m[31]&m[192]&m[193]&m[194]&m[195]));
    m[69] = (((m[32]&m[202]&~m[203]&~m[204]&~m[205])|(m[32]&~m[202]&m[203]&~m[204]&~m[205])|(~m[32]&m[202]&m[203]&~m[204]&~m[205])|(m[32]&~m[202]&~m[203]&m[204]&~m[205])|(~m[32]&m[202]&~m[203]&m[204]&~m[205])|(~m[32]&~m[202]&m[203]&m[204]&~m[205])|(m[32]&~m[202]&~m[203]&~m[204]&m[205])|(~m[32]&m[202]&~m[203]&~m[204]&m[205])|(~m[32]&~m[202]&m[203]&~m[204]&m[205])|(~m[32]&~m[202]&~m[203]&m[204]&m[205]))&BiasedRNG[8])|(((m[32]&m[202]&m[203]&~m[204]&~m[205])|(m[32]&m[202]&~m[203]&m[204]&~m[205])|(m[32]&~m[202]&m[203]&m[204]&~m[205])|(~m[32]&m[202]&m[203]&m[204]&~m[205])|(m[32]&m[202]&~m[203]&~m[204]&m[205])|(m[32]&~m[202]&m[203]&~m[204]&m[205])|(~m[32]&m[202]&m[203]&~m[204]&m[205])|(m[32]&~m[202]&~m[203]&m[204]&m[205])|(~m[32]&m[202]&~m[203]&m[204]&m[205])|(~m[32]&~m[202]&m[203]&m[204]&m[205]))&~BiasedRNG[8])|((m[32]&m[202]&m[203]&m[204]&~m[205])|(m[32]&m[202]&m[203]&~m[204]&m[205])|(m[32]&m[202]&~m[203]&m[204]&m[205])|(m[32]&~m[202]&m[203]&m[204]&m[205])|(~m[32]&m[202]&m[203]&m[204]&m[205])|(m[32]&m[202]&m[203]&m[204]&m[205]));
    m[70] = (((m[32]&m[206]&~m[207]&~m[208]&~m[209])|(m[32]&~m[206]&m[207]&~m[208]&~m[209])|(~m[32]&m[206]&m[207]&~m[208]&~m[209])|(m[32]&~m[206]&~m[207]&m[208]&~m[209])|(~m[32]&m[206]&~m[207]&m[208]&~m[209])|(~m[32]&~m[206]&m[207]&m[208]&~m[209])|(m[32]&~m[206]&~m[207]&~m[208]&m[209])|(~m[32]&m[206]&~m[207]&~m[208]&m[209])|(~m[32]&~m[206]&m[207]&~m[208]&m[209])|(~m[32]&~m[206]&~m[207]&m[208]&m[209]))&BiasedRNG[9])|(((m[32]&m[206]&m[207]&~m[208]&~m[209])|(m[32]&m[206]&~m[207]&m[208]&~m[209])|(m[32]&~m[206]&m[207]&m[208]&~m[209])|(~m[32]&m[206]&m[207]&m[208]&~m[209])|(m[32]&m[206]&~m[207]&~m[208]&m[209])|(m[32]&~m[206]&m[207]&~m[208]&m[209])|(~m[32]&m[206]&m[207]&~m[208]&m[209])|(m[32]&~m[206]&~m[207]&m[208]&m[209])|(~m[32]&m[206]&~m[207]&m[208]&m[209])|(~m[32]&~m[206]&m[207]&m[208]&m[209]))&~BiasedRNG[9])|((m[32]&m[206]&m[207]&m[208]&~m[209])|(m[32]&m[206]&m[207]&~m[208]&m[209])|(m[32]&m[206]&~m[207]&m[208]&m[209])|(m[32]&~m[206]&m[207]&m[208]&m[209])|(~m[32]&m[206]&m[207]&m[208]&m[209])|(m[32]&m[206]&m[207]&m[208]&m[209]));
    m[72] = (((m[33]&m[216]&~m[217]&~m[218]&~m[219])|(m[33]&~m[216]&m[217]&~m[218]&~m[219])|(~m[33]&m[216]&m[217]&~m[218]&~m[219])|(m[33]&~m[216]&~m[217]&m[218]&~m[219])|(~m[33]&m[216]&~m[217]&m[218]&~m[219])|(~m[33]&~m[216]&m[217]&m[218]&~m[219])|(m[33]&~m[216]&~m[217]&~m[218]&m[219])|(~m[33]&m[216]&~m[217]&~m[218]&m[219])|(~m[33]&~m[216]&m[217]&~m[218]&m[219])|(~m[33]&~m[216]&~m[217]&m[218]&m[219]))&BiasedRNG[10])|(((m[33]&m[216]&m[217]&~m[218]&~m[219])|(m[33]&m[216]&~m[217]&m[218]&~m[219])|(m[33]&~m[216]&m[217]&m[218]&~m[219])|(~m[33]&m[216]&m[217]&m[218]&~m[219])|(m[33]&m[216]&~m[217]&~m[218]&m[219])|(m[33]&~m[216]&m[217]&~m[218]&m[219])|(~m[33]&m[216]&m[217]&~m[218]&m[219])|(m[33]&~m[216]&~m[217]&m[218]&m[219])|(~m[33]&m[216]&~m[217]&m[218]&m[219])|(~m[33]&~m[216]&m[217]&m[218]&m[219]))&~BiasedRNG[10])|((m[33]&m[216]&m[217]&m[218]&~m[219])|(m[33]&m[216]&m[217]&~m[218]&m[219])|(m[33]&m[216]&~m[217]&m[218]&m[219])|(m[33]&~m[216]&m[217]&m[218]&m[219])|(~m[33]&m[216]&m[217]&m[218]&m[219])|(m[33]&m[216]&m[217]&m[218]&m[219]));
    m[73] = (((m[33]&m[220]&~m[221]&~m[222]&~m[223])|(m[33]&~m[220]&m[221]&~m[222]&~m[223])|(~m[33]&m[220]&m[221]&~m[222]&~m[223])|(m[33]&~m[220]&~m[221]&m[222]&~m[223])|(~m[33]&m[220]&~m[221]&m[222]&~m[223])|(~m[33]&~m[220]&m[221]&m[222]&~m[223])|(m[33]&~m[220]&~m[221]&~m[222]&m[223])|(~m[33]&m[220]&~m[221]&~m[222]&m[223])|(~m[33]&~m[220]&m[221]&~m[222]&m[223])|(~m[33]&~m[220]&~m[221]&m[222]&m[223]))&BiasedRNG[11])|(((m[33]&m[220]&m[221]&~m[222]&~m[223])|(m[33]&m[220]&~m[221]&m[222]&~m[223])|(m[33]&~m[220]&m[221]&m[222]&~m[223])|(~m[33]&m[220]&m[221]&m[222]&~m[223])|(m[33]&m[220]&~m[221]&~m[222]&m[223])|(m[33]&~m[220]&m[221]&~m[222]&m[223])|(~m[33]&m[220]&m[221]&~m[222]&m[223])|(m[33]&~m[220]&~m[221]&m[222]&m[223])|(~m[33]&m[220]&~m[221]&m[222]&m[223])|(~m[33]&~m[220]&m[221]&m[222]&m[223]))&~BiasedRNG[11])|((m[33]&m[220]&m[221]&m[222]&~m[223])|(m[33]&m[220]&m[221]&~m[222]&m[223])|(m[33]&m[220]&~m[221]&m[222]&m[223])|(m[33]&~m[220]&m[221]&m[222]&m[223])|(~m[33]&m[220]&m[221]&m[222]&m[223])|(m[33]&m[220]&m[221]&m[222]&m[223]));
    m[75] = (((m[34]&m[230]&~m[231]&~m[232]&~m[233])|(m[34]&~m[230]&m[231]&~m[232]&~m[233])|(~m[34]&m[230]&m[231]&~m[232]&~m[233])|(m[34]&~m[230]&~m[231]&m[232]&~m[233])|(~m[34]&m[230]&~m[231]&m[232]&~m[233])|(~m[34]&~m[230]&m[231]&m[232]&~m[233])|(m[34]&~m[230]&~m[231]&~m[232]&m[233])|(~m[34]&m[230]&~m[231]&~m[232]&m[233])|(~m[34]&~m[230]&m[231]&~m[232]&m[233])|(~m[34]&~m[230]&~m[231]&m[232]&m[233]))&BiasedRNG[12])|(((m[34]&m[230]&m[231]&~m[232]&~m[233])|(m[34]&m[230]&~m[231]&m[232]&~m[233])|(m[34]&~m[230]&m[231]&m[232]&~m[233])|(~m[34]&m[230]&m[231]&m[232]&~m[233])|(m[34]&m[230]&~m[231]&~m[232]&m[233])|(m[34]&~m[230]&m[231]&~m[232]&m[233])|(~m[34]&m[230]&m[231]&~m[232]&m[233])|(m[34]&~m[230]&~m[231]&m[232]&m[233])|(~m[34]&m[230]&~m[231]&m[232]&m[233])|(~m[34]&~m[230]&m[231]&m[232]&m[233]))&~BiasedRNG[12])|((m[34]&m[230]&m[231]&m[232]&~m[233])|(m[34]&m[230]&m[231]&~m[232]&m[233])|(m[34]&m[230]&~m[231]&m[232]&m[233])|(m[34]&~m[230]&m[231]&m[232]&m[233])|(~m[34]&m[230]&m[231]&m[232]&m[233])|(m[34]&m[230]&m[231]&m[232]&m[233]));
    m[76] = (((m[34]&m[234]&~m[235]&~m[236]&~m[237])|(m[34]&~m[234]&m[235]&~m[236]&~m[237])|(~m[34]&m[234]&m[235]&~m[236]&~m[237])|(m[34]&~m[234]&~m[235]&m[236]&~m[237])|(~m[34]&m[234]&~m[235]&m[236]&~m[237])|(~m[34]&~m[234]&m[235]&m[236]&~m[237])|(m[34]&~m[234]&~m[235]&~m[236]&m[237])|(~m[34]&m[234]&~m[235]&~m[236]&m[237])|(~m[34]&~m[234]&m[235]&~m[236]&m[237])|(~m[34]&~m[234]&~m[235]&m[236]&m[237]))&BiasedRNG[13])|(((m[34]&m[234]&m[235]&~m[236]&~m[237])|(m[34]&m[234]&~m[235]&m[236]&~m[237])|(m[34]&~m[234]&m[235]&m[236]&~m[237])|(~m[34]&m[234]&m[235]&m[236]&~m[237])|(m[34]&m[234]&~m[235]&~m[236]&m[237])|(m[34]&~m[234]&m[235]&~m[236]&m[237])|(~m[34]&m[234]&m[235]&~m[236]&m[237])|(m[34]&~m[234]&~m[235]&m[236]&m[237])|(~m[34]&m[234]&~m[235]&m[236]&m[237])|(~m[34]&~m[234]&m[235]&m[236]&m[237]))&~BiasedRNG[13])|((m[34]&m[234]&m[235]&m[236]&~m[237])|(m[34]&m[234]&m[235]&~m[236]&m[237])|(m[34]&m[234]&~m[235]&m[236]&m[237])|(m[34]&~m[234]&m[235]&m[236]&m[237])|(~m[34]&m[234]&m[235]&m[236]&m[237])|(m[34]&m[234]&m[235]&m[236]&m[237]));
    m[78] = (((m[35]&m[244]&~m[245]&~m[246]&~m[247])|(m[35]&~m[244]&m[245]&~m[246]&~m[247])|(~m[35]&m[244]&m[245]&~m[246]&~m[247])|(m[35]&~m[244]&~m[245]&m[246]&~m[247])|(~m[35]&m[244]&~m[245]&m[246]&~m[247])|(~m[35]&~m[244]&m[245]&m[246]&~m[247])|(m[35]&~m[244]&~m[245]&~m[246]&m[247])|(~m[35]&m[244]&~m[245]&~m[246]&m[247])|(~m[35]&~m[244]&m[245]&~m[246]&m[247])|(~m[35]&~m[244]&~m[245]&m[246]&m[247]))&BiasedRNG[14])|(((m[35]&m[244]&m[245]&~m[246]&~m[247])|(m[35]&m[244]&~m[245]&m[246]&~m[247])|(m[35]&~m[244]&m[245]&m[246]&~m[247])|(~m[35]&m[244]&m[245]&m[246]&~m[247])|(m[35]&m[244]&~m[245]&~m[246]&m[247])|(m[35]&~m[244]&m[245]&~m[246]&m[247])|(~m[35]&m[244]&m[245]&~m[246]&m[247])|(m[35]&~m[244]&~m[245]&m[246]&m[247])|(~m[35]&m[244]&~m[245]&m[246]&m[247])|(~m[35]&~m[244]&m[245]&m[246]&m[247]))&~BiasedRNG[14])|((m[35]&m[244]&m[245]&m[246]&~m[247])|(m[35]&m[244]&m[245]&~m[246]&m[247])|(m[35]&m[244]&~m[245]&m[246]&m[247])|(m[35]&~m[244]&m[245]&m[246]&m[247])|(~m[35]&m[244]&m[245]&m[246]&m[247])|(m[35]&m[244]&m[245]&m[246]&m[247]));
    m[79] = (((m[35]&m[248]&~m[249]&~m[250]&~m[251])|(m[35]&~m[248]&m[249]&~m[250]&~m[251])|(~m[35]&m[248]&m[249]&~m[250]&~m[251])|(m[35]&~m[248]&~m[249]&m[250]&~m[251])|(~m[35]&m[248]&~m[249]&m[250]&~m[251])|(~m[35]&~m[248]&m[249]&m[250]&~m[251])|(m[35]&~m[248]&~m[249]&~m[250]&m[251])|(~m[35]&m[248]&~m[249]&~m[250]&m[251])|(~m[35]&~m[248]&m[249]&~m[250]&m[251])|(~m[35]&~m[248]&~m[249]&m[250]&m[251]))&BiasedRNG[15])|(((m[35]&m[248]&m[249]&~m[250]&~m[251])|(m[35]&m[248]&~m[249]&m[250]&~m[251])|(m[35]&~m[248]&m[249]&m[250]&~m[251])|(~m[35]&m[248]&m[249]&m[250]&~m[251])|(m[35]&m[248]&~m[249]&~m[250]&m[251])|(m[35]&~m[248]&m[249]&~m[250]&m[251])|(~m[35]&m[248]&m[249]&~m[250]&m[251])|(m[35]&~m[248]&~m[249]&m[250]&m[251])|(~m[35]&m[248]&~m[249]&m[250]&m[251])|(~m[35]&~m[248]&m[249]&m[250]&m[251]))&~BiasedRNG[15])|((m[35]&m[248]&m[249]&m[250]&~m[251])|(m[35]&m[248]&m[249]&~m[250]&m[251])|(m[35]&m[248]&~m[249]&m[250]&m[251])|(m[35]&~m[248]&m[249]&m[250]&m[251])|(~m[35]&m[248]&m[249]&m[250]&m[251])|(m[35]&m[248]&m[249]&m[250]&m[251]));
    m[81] = (((m[36]&m[258]&~m[259]&~m[260]&~m[261])|(m[36]&~m[258]&m[259]&~m[260]&~m[261])|(~m[36]&m[258]&m[259]&~m[260]&~m[261])|(m[36]&~m[258]&~m[259]&m[260]&~m[261])|(~m[36]&m[258]&~m[259]&m[260]&~m[261])|(~m[36]&~m[258]&m[259]&m[260]&~m[261])|(m[36]&~m[258]&~m[259]&~m[260]&m[261])|(~m[36]&m[258]&~m[259]&~m[260]&m[261])|(~m[36]&~m[258]&m[259]&~m[260]&m[261])|(~m[36]&~m[258]&~m[259]&m[260]&m[261]))&BiasedRNG[16])|(((m[36]&m[258]&m[259]&~m[260]&~m[261])|(m[36]&m[258]&~m[259]&m[260]&~m[261])|(m[36]&~m[258]&m[259]&m[260]&~m[261])|(~m[36]&m[258]&m[259]&m[260]&~m[261])|(m[36]&m[258]&~m[259]&~m[260]&m[261])|(m[36]&~m[258]&m[259]&~m[260]&m[261])|(~m[36]&m[258]&m[259]&~m[260]&m[261])|(m[36]&~m[258]&~m[259]&m[260]&m[261])|(~m[36]&m[258]&~m[259]&m[260]&m[261])|(~m[36]&~m[258]&m[259]&m[260]&m[261]))&~BiasedRNG[16])|((m[36]&m[258]&m[259]&m[260]&~m[261])|(m[36]&m[258]&m[259]&~m[260]&m[261])|(m[36]&m[258]&~m[259]&m[260]&m[261])|(m[36]&~m[258]&m[259]&m[260]&m[261])|(~m[36]&m[258]&m[259]&m[260]&m[261])|(m[36]&m[258]&m[259]&m[260]&m[261]));
    m[82] = (((m[36]&m[262]&~m[263]&~m[264]&~m[265])|(m[36]&~m[262]&m[263]&~m[264]&~m[265])|(~m[36]&m[262]&m[263]&~m[264]&~m[265])|(m[36]&~m[262]&~m[263]&m[264]&~m[265])|(~m[36]&m[262]&~m[263]&m[264]&~m[265])|(~m[36]&~m[262]&m[263]&m[264]&~m[265])|(m[36]&~m[262]&~m[263]&~m[264]&m[265])|(~m[36]&m[262]&~m[263]&~m[264]&m[265])|(~m[36]&~m[262]&m[263]&~m[264]&m[265])|(~m[36]&~m[262]&~m[263]&m[264]&m[265]))&BiasedRNG[17])|(((m[36]&m[262]&m[263]&~m[264]&~m[265])|(m[36]&m[262]&~m[263]&m[264]&~m[265])|(m[36]&~m[262]&m[263]&m[264]&~m[265])|(~m[36]&m[262]&m[263]&m[264]&~m[265])|(m[36]&m[262]&~m[263]&~m[264]&m[265])|(m[36]&~m[262]&m[263]&~m[264]&m[265])|(~m[36]&m[262]&m[263]&~m[264]&m[265])|(m[36]&~m[262]&~m[263]&m[264]&m[265])|(~m[36]&m[262]&~m[263]&m[264]&m[265])|(~m[36]&~m[262]&m[263]&m[264]&m[265]))&~BiasedRNG[17])|((m[36]&m[262]&m[263]&m[264]&~m[265])|(m[36]&m[262]&m[263]&~m[264]&m[265])|(m[36]&m[262]&~m[263]&m[264]&m[265])|(m[36]&~m[262]&m[263]&m[264]&m[265])|(~m[36]&m[262]&m[263]&m[264]&m[265])|(m[36]&m[262]&m[263]&m[264]&m[265]));
    m[84] = (((m[37]&m[272]&~m[273]&~m[274]&~m[275])|(m[37]&~m[272]&m[273]&~m[274]&~m[275])|(~m[37]&m[272]&m[273]&~m[274]&~m[275])|(m[37]&~m[272]&~m[273]&m[274]&~m[275])|(~m[37]&m[272]&~m[273]&m[274]&~m[275])|(~m[37]&~m[272]&m[273]&m[274]&~m[275])|(m[37]&~m[272]&~m[273]&~m[274]&m[275])|(~m[37]&m[272]&~m[273]&~m[274]&m[275])|(~m[37]&~m[272]&m[273]&~m[274]&m[275])|(~m[37]&~m[272]&~m[273]&m[274]&m[275]))&BiasedRNG[18])|(((m[37]&m[272]&m[273]&~m[274]&~m[275])|(m[37]&m[272]&~m[273]&m[274]&~m[275])|(m[37]&~m[272]&m[273]&m[274]&~m[275])|(~m[37]&m[272]&m[273]&m[274]&~m[275])|(m[37]&m[272]&~m[273]&~m[274]&m[275])|(m[37]&~m[272]&m[273]&~m[274]&m[275])|(~m[37]&m[272]&m[273]&~m[274]&m[275])|(m[37]&~m[272]&~m[273]&m[274]&m[275])|(~m[37]&m[272]&~m[273]&m[274]&m[275])|(~m[37]&~m[272]&m[273]&m[274]&m[275]))&~BiasedRNG[18])|((m[37]&m[272]&m[273]&m[274]&~m[275])|(m[37]&m[272]&m[273]&~m[274]&m[275])|(m[37]&m[272]&~m[273]&m[274]&m[275])|(m[37]&~m[272]&m[273]&m[274]&m[275])|(~m[37]&m[272]&m[273]&m[274]&m[275])|(m[37]&m[272]&m[273]&m[274]&m[275]));
    m[85] = (((m[37]&m[276]&~m[277]&~m[278]&~m[279])|(m[37]&~m[276]&m[277]&~m[278]&~m[279])|(~m[37]&m[276]&m[277]&~m[278]&~m[279])|(m[37]&~m[276]&~m[277]&m[278]&~m[279])|(~m[37]&m[276]&~m[277]&m[278]&~m[279])|(~m[37]&~m[276]&m[277]&m[278]&~m[279])|(m[37]&~m[276]&~m[277]&~m[278]&m[279])|(~m[37]&m[276]&~m[277]&~m[278]&m[279])|(~m[37]&~m[276]&m[277]&~m[278]&m[279])|(~m[37]&~m[276]&~m[277]&m[278]&m[279]))&BiasedRNG[19])|(((m[37]&m[276]&m[277]&~m[278]&~m[279])|(m[37]&m[276]&~m[277]&m[278]&~m[279])|(m[37]&~m[276]&m[277]&m[278]&~m[279])|(~m[37]&m[276]&m[277]&m[278]&~m[279])|(m[37]&m[276]&~m[277]&~m[278]&m[279])|(m[37]&~m[276]&m[277]&~m[278]&m[279])|(~m[37]&m[276]&m[277]&~m[278]&m[279])|(m[37]&~m[276]&~m[277]&m[278]&m[279])|(~m[37]&m[276]&~m[277]&m[278]&m[279])|(~m[37]&~m[276]&m[277]&m[278]&m[279]))&~BiasedRNG[19])|((m[37]&m[276]&m[277]&m[278]&~m[279])|(m[37]&m[276]&m[277]&~m[278]&m[279])|(m[37]&m[276]&~m[277]&m[278]&m[279])|(m[37]&~m[276]&m[277]&m[278]&m[279])|(~m[37]&m[276]&m[277]&m[278]&m[279])|(m[37]&m[276]&m[277]&m[278]&m[279]));
    m[87] = (((m[38]&m[286]&~m[287]&~m[288]&~m[289])|(m[38]&~m[286]&m[287]&~m[288]&~m[289])|(~m[38]&m[286]&m[287]&~m[288]&~m[289])|(m[38]&~m[286]&~m[287]&m[288]&~m[289])|(~m[38]&m[286]&~m[287]&m[288]&~m[289])|(~m[38]&~m[286]&m[287]&m[288]&~m[289])|(m[38]&~m[286]&~m[287]&~m[288]&m[289])|(~m[38]&m[286]&~m[287]&~m[288]&m[289])|(~m[38]&~m[286]&m[287]&~m[288]&m[289])|(~m[38]&~m[286]&~m[287]&m[288]&m[289]))&BiasedRNG[20])|(((m[38]&m[286]&m[287]&~m[288]&~m[289])|(m[38]&m[286]&~m[287]&m[288]&~m[289])|(m[38]&~m[286]&m[287]&m[288]&~m[289])|(~m[38]&m[286]&m[287]&m[288]&~m[289])|(m[38]&m[286]&~m[287]&~m[288]&m[289])|(m[38]&~m[286]&m[287]&~m[288]&m[289])|(~m[38]&m[286]&m[287]&~m[288]&m[289])|(m[38]&~m[286]&~m[287]&m[288]&m[289])|(~m[38]&m[286]&~m[287]&m[288]&m[289])|(~m[38]&~m[286]&m[287]&m[288]&m[289]))&~BiasedRNG[20])|((m[38]&m[286]&m[287]&m[288]&~m[289])|(m[38]&m[286]&m[287]&~m[288]&m[289])|(m[38]&m[286]&~m[287]&m[288]&m[289])|(m[38]&~m[286]&m[287]&m[288]&m[289])|(~m[38]&m[286]&m[287]&m[288]&m[289])|(m[38]&m[286]&m[287]&m[288]&m[289]));
    m[88] = (((m[38]&m[290]&~m[291]&~m[292]&~m[293])|(m[38]&~m[290]&m[291]&~m[292]&~m[293])|(~m[38]&m[290]&m[291]&~m[292]&~m[293])|(m[38]&~m[290]&~m[291]&m[292]&~m[293])|(~m[38]&m[290]&~m[291]&m[292]&~m[293])|(~m[38]&~m[290]&m[291]&m[292]&~m[293])|(m[38]&~m[290]&~m[291]&~m[292]&m[293])|(~m[38]&m[290]&~m[291]&~m[292]&m[293])|(~m[38]&~m[290]&m[291]&~m[292]&m[293])|(~m[38]&~m[290]&~m[291]&m[292]&m[293]))&BiasedRNG[21])|(((m[38]&m[290]&m[291]&~m[292]&~m[293])|(m[38]&m[290]&~m[291]&m[292]&~m[293])|(m[38]&~m[290]&m[291]&m[292]&~m[293])|(~m[38]&m[290]&m[291]&m[292]&~m[293])|(m[38]&m[290]&~m[291]&~m[292]&m[293])|(m[38]&~m[290]&m[291]&~m[292]&m[293])|(~m[38]&m[290]&m[291]&~m[292]&m[293])|(m[38]&~m[290]&~m[291]&m[292]&m[293])|(~m[38]&m[290]&~m[291]&m[292]&m[293])|(~m[38]&~m[290]&m[291]&m[292]&m[293]))&~BiasedRNG[21])|((m[38]&m[290]&m[291]&m[292]&~m[293])|(m[38]&m[290]&m[291]&~m[292]&m[293])|(m[38]&m[290]&~m[291]&m[292]&m[293])|(m[38]&~m[290]&m[291]&m[292]&m[293])|(~m[38]&m[290]&m[291]&m[292]&m[293])|(m[38]&m[290]&m[291]&m[292]&m[293]));
    m[90] = (((m[39]&m[300]&~m[301]&~m[302]&~m[303])|(m[39]&~m[300]&m[301]&~m[302]&~m[303])|(~m[39]&m[300]&m[301]&~m[302]&~m[303])|(m[39]&~m[300]&~m[301]&m[302]&~m[303])|(~m[39]&m[300]&~m[301]&m[302]&~m[303])|(~m[39]&~m[300]&m[301]&m[302]&~m[303])|(m[39]&~m[300]&~m[301]&~m[302]&m[303])|(~m[39]&m[300]&~m[301]&~m[302]&m[303])|(~m[39]&~m[300]&m[301]&~m[302]&m[303])|(~m[39]&~m[300]&~m[301]&m[302]&m[303]))&BiasedRNG[22])|(((m[39]&m[300]&m[301]&~m[302]&~m[303])|(m[39]&m[300]&~m[301]&m[302]&~m[303])|(m[39]&~m[300]&m[301]&m[302]&~m[303])|(~m[39]&m[300]&m[301]&m[302]&~m[303])|(m[39]&m[300]&~m[301]&~m[302]&m[303])|(m[39]&~m[300]&m[301]&~m[302]&m[303])|(~m[39]&m[300]&m[301]&~m[302]&m[303])|(m[39]&~m[300]&~m[301]&m[302]&m[303])|(~m[39]&m[300]&~m[301]&m[302]&m[303])|(~m[39]&~m[300]&m[301]&m[302]&m[303]))&~BiasedRNG[22])|((m[39]&m[300]&m[301]&m[302]&~m[303])|(m[39]&m[300]&m[301]&~m[302]&m[303])|(m[39]&m[300]&~m[301]&m[302]&m[303])|(m[39]&~m[300]&m[301]&m[302]&m[303])|(~m[39]&m[300]&m[301]&m[302]&m[303])|(m[39]&m[300]&m[301]&m[302]&m[303]));
    m[91] = (((m[39]&m[304]&~m[305]&~m[306]&~m[307])|(m[39]&~m[304]&m[305]&~m[306]&~m[307])|(~m[39]&m[304]&m[305]&~m[306]&~m[307])|(m[39]&~m[304]&~m[305]&m[306]&~m[307])|(~m[39]&m[304]&~m[305]&m[306]&~m[307])|(~m[39]&~m[304]&m[305]&m[306]&~m[307])|(m[39]&~m[304]&~m[305]&~m[306]&m[307])|(~m[39]&m[304]&~m[305]&~m[306]&m[307])|(~m[39]&~m[304]&m[305]&~m[306]&m[307])|(~m[39]&~m[304]&~m[305]&m[306]&m[307]))&BiasedRNG[23])|(((m[39]&m[304]&m[305]&~m[306]&~m[307])|(m[39]&m[304]&~m[305]&m[306]&~m[307])|(m[39]&~m[304]&m[305]&m[306]&~m[307])|(~m[39]&m[304]&m[305]&m[306]&~m[307])|(m[39]&m[304]&~m[305]&~m[306]&m[307])|(m[39]&~m[304]&m[305]&~m[306]&m[307])|(~m[39]&m[304]&m[305]&~m[306]&m[307])|(m[39]&~m[304]&~m[305]&m[306]&m[307])|(~m[39]&m[304]&~m[305]&m[306]&m[307])|(~m[39]&~m[304]&m[305]&m[306]&m[307]))&~BiasedRNG[23])|((m[39]&m[304]&m[305]&m[306]&~m[307])|(m[39]&m[304]&m[305]&~m[306]&m[307])|(m[39]&m[304]&~m[305]&m[306]&m[307])|(m[39]&~m[304]&m[305]&m[306]&m[307])|(~m[39]&m[304]&m[305]&m[306]&m[307])|(m[39]&m[304]&m[305]&m[306]&m[307]));
    m[93] = (((m[40]&m[314]&~m[315]&~m[316]&~m[317])|(m[40]&~m[314]&m[315]&~m[316]&~m[317])|(~m[40]&m[314]&m[315]&~m[316]&~m[317])|(m[40]&~m[314]&~m[315]&m[316]&~m[317])|(~m[40]&m[314]&~m[315]&m[316]&~m[317])|(~m[40]&~m[314]&m[315]&m[316]&~m[317])|(m[40]&~m[314]&~m[315]&~m[316]&m[317])|(~m[40]&m[314]&~m[315]&~m[316]&m[317])|(~m[40]&~m[314]&m[315]&~m[316]&m[317])|(~m[40]&~m[314]&~m[315]&m[316]&m[317]))&BiasedRNG[24])|(((m[40]&m[314]&m[315]&~m[316]&~m[317])|(m[40]&m[314]&~m[315]&m[316]&~m[317])|(m[40]&~m[314]&m[315]&m[316]&~m[317])|(~m[40]&m[314]&m[315]&m[316]&~m[317])|(m[40]&m[314]&~m[315]&~m[316]&m[317])|(m[40]&~m[314]&m[315]&~m[316]&m[317])|(~m[40]&m[314]&m[315]&~m[316]&m[317])|(m[40]&~m[314]&~m[315]&m[316]&m[317])|(~m[40]&m[314]&~m[315]&m[316]&m[317])|(~m[40]&~m[314]&m[315]&m[316]&m[317]))&~BiasedRNG[24])|((m[40]&m[314]&m[315]&m[316]&~m[317])|(m[40]&m[314]&m[315]&~m[316]&m[317])|(m[40]&m[314]&~m[315]&m[316]&m[317])|(m[40]&~m[314]&m[315]&m[316]&m[317])|(~m[40]&m[314]&m[315]&m[316]&m[317])|(m[40]&m[314]&m[315]&m[316]&m[317]));
    m[94] = (((m[40]&m[318]&~m[319]&~m[320]&~m[321])|(m[40]&~m[318]&m[319]&~m[320]&~m[321])|(~m[40]&m[318]&m[319]&~m[320]&~m[321])|(m[40]&~m[318]&~m[319]&m[320]&~m[321])|(~m[40]&m[318]&~m[319]&m[320]&~m[321])|(~m[40]&~m[318]&m[319]&m[320]&~m[321])|(m[40]&~m[318]&~m[319]&~m[320]&m[321])|(~m[40]&m[318]&~m[319]&~m[320]&m[321])|(~m[40]&~m[318]&m[319]&~m[320]&m[321])|(~m[40]&~m[318]&~m[319]&m[320]&m[321]))&BiasedRNG[25])|(((m[40]&m[318]&m[319]&~m[320]&~m[321])|(m[40]&m[318]&~m[319]&m[320]&~m[321])|(m[40]&~m[318]&m[319]&m[320]&~m[321])|(~m[40]&m[318]&m[319]&m[320]&~m[321])|(m[40]&m[318]&~m[319]&~m[320]&m[321])|(m[40]&~m[318]&m[319]&~m[320]&m[321])|(~m[40]&m[318]&m[319]&~m[320]&m[321])|(m[40]&~m[318]&~m[319]&m[320]&m[321])|(~m[40]&m[318]&~m[319]&m[320]&m[321])|(~m[40]&~m[318]&m[319]&m[320]&m[321]))&~BiasedRNG[25])|((m[40]&m[318]&m[319]&m[320]&~m[321])|(m[40]&m[318]&m[319]&~m[320]&m[321])|(m[40]&m[318]&~m[319]&m[320]&m[321])|(m[40]&~m[318]&m[319]&m[320]&m[321])|(~m[40]&m[318]&m[319]&m[320]&m[321])|(m[40]&m[318]&m[319]&m[320]&m[321]));
    m[96] = (((m[41]&m[328]&~m[329]&~m[330]&~m[331])|(m[41]&~m[328]&m[329]&~m[330]&~m[331])|(~m[41]&m[328]&m[329]&~m[330]&~m[331])|(m[41]&~m[328]&~m[329]&m[330]&~m[331])|(~m[41]&m[328]&~m[329]&m[330]&~m[331])|(~m[41]&~m[328]&m[329]&m[330]&~m[331])|(m[41]&~m[328]&~m[329]&~m[330]&m[331])|(~m[41]&m[328]&~m[329]&~m[330]&m[331])|(~m[41]&~m[328]&m[329]&~m[330]&m[331])|(~m[41]&~m[328]&~m[329]&m[330]&m[331]))&BiasedRNG[26])|(((m[41]&m[328]&m[329]&~m[330]&~m[331])|(m[41]&m[328]&~m[329]&m[330]&~m[331])|(m[41]&~m[328]&m[329]&m[330]&~m[331])|(~m[41]&m[328]&m[329]&m[330]&~m[331])|(m[41]&m[328]&~m[329]&~m[330]&m[331])|(m[41]&~m[328]&m[329]&~m[330]&m[331])|(~m[41]&m[328]&m[329]&~m[330]&m[331])|(m[41]&~m[328]&~m[329]&m[330]&m[331])|(~m[41]&m[328]&~m[329]&m[330]&m[331])|(~m[41]&~m[328]&m[329]&m[330]&m[331]))&~BiasedRNG[26])|((m[41]&m[328]&m[329]&m[330]&~m[331])|(m[41]&m[328]&m[329]&~m[330]&m[331])|(m[41]&m[328]&~m[329]&m[330]&m[331])|(m[41]&~m[328]&m[329]&m[330]&m[331])|(~m[41]&m[328]&m[329]&m[330]&m[331])|(m[41]&m[328]&m[329]&m[330]&m[331]));
    m[97] = (((m[41]&m[332]&~m[333]&~m[334]&~m[335])|(m[41]&~m[332]&m[333]&~m[334]&~m[335])|(~m[41]&m[332]&m[333]&~m[334]&~m[335])|(m[41]&~m[332]&~m[333]&m[334]&~m[335])|(~m[41]&m[332]&~m[333]&m[334]&~m[335])|(~m[41]&~m[332]&m[333]&m[334]&~m[335])|(m[41]&~m[332]&~m[333]&~m[334]&m[335])|(~m[41]&m[332]&~m[333]&~m[334]&m[335])|(~m[41]&~m[332]&m[333]&~m[334]&m[335])|(~m[41]&~m[332]&~m[333]&m[334]&m[335]))&BiasedRNG[27])|(((m[41]&m[332]&m[333]&~m[334]&~m[335])|(m[41]&m[332]&~m[333]&m[334]&~m[335])|(m[41]&~m[332]&m[333]&m[334]&~m[335])|(~m[41]&m[332]&m[333]&m[334]&~m[335])|(m[41]&m[332]&~m[333]&~m[334]&m[335])|(m[41]&~m[332]&m[333]&~m[334]&m[335])|(~m[41]&m[332]&m[333]&~m[334]&m[335])|(m[41]&~m[332]&~m[333]&m[334]&m[335])|(~m[41]&m[332]&~m[333]&m[334]&m[335])|(~m[41]&~m[332]&m[333]&m[334]&m[335]))&~BiasedRNG[27])|((m[41]&m[332]&m[333]&m[334]&~m[335])|(m[41]&m[332]&m[333]&~m[334]&m[335])|(m[41]&m[332]&~m[333]&m[334]&m[335])|(m[41]&~m[332]&m[333]&m[334]&m[335])|(~m[41]&m[332]&m[333]&m[334]&m[335])|(m[41]&m[332]&m[333]&m[334]&m[335]));
    m[99] = (((m[42]&m[342]&~m[343]&~m[344]&~m[345])|(m[42]&~m[342]&m[343]&~m[344]&~m[345])|(~m[42]&m[342]&m[343]&~m[344]&~m[345])|(m[42]&~m[342]&~m[343]&m[344]&~m[345])|(~m[42]&m[342]&~m[343]&m[344]&~m[345])|(~m[42]&~m[342]&m[343]&m[344]&~m[345])|(m[42]&~m[342]&~m[343]&~m[344]&m[345])|(~m[42]&m[342]&~m[343]&~m[344]&m[345])|(~m[42]&~m[342]&m[343]&~m[344]&m[345])|(~m[42]&~m[342]&~m[343]&m[344]&m[345]))&BiasedRNG[28])|(((m[42]&m[342]&m[343]&~m[344]&~m[345])|(m[42]&m[342]&~m[343]&m[344]&~m[345])|(m[42]&~m[342]&m[343]&m[344]&~m[345])|(~m[42]&m[342]&m[343]&m[344]&~m[345])|(m[42]&m[342]&~m[343]&~m[344]&m[345])|(m[42]&~m[342]&m[343]&~m[344]&m[345])|(~m[42]&m[342]&m[343]&~m[344]&m[345])|(m[42]&~m[342]&~m[343]&m[344]&m[345])|(~m[42]&m[342]&~m[343]&m[344]&m[345])|(~m[42]&~m[342]&m[343]&m[344]&m[345]))&~BiasedRNG[28])|((m[42]&m[342]&m[343]&m[344]&~m[345])|(m[42]&m[342]&m[343]&~m[344]&m[345])|(m[42]&m[342]&~m[343]&m[344]&m[345])|(m[42]&~m[342]&m[343]&m[344]&m[345])|(~m[42]&m[342]&m[343]&m[344]&m[345])|(m[42]&m[342]&m[343]&m[344]&m[345]));
    m[100] = (((m[42]&m[346]&~m[347]&~m[348]&~m[349])|(m[42]&~m[346]&m[347]&~m[348]&~m[349])|(~m[42]&m[346]&m[347]&~m[348]&~m[349])|(m[42]&~m[346]&~m[347]&m[348]&~m[349])|(~m[42]&m[346]&~m[347]&m[348]&~m[349])|(~m[42]&~m[346]&m[347]&m[348]&~m[349])|(m[42]&~m[346]&~m[347]&~m[348]&m[349])|(~m[42]&m[346]&~m[347]&~m[348]&m[349])|(~m[42]&~m[346]&m[347]&~m[348]&m[349])|(~m[42]&~m[346]&~m[347]&m[348]&m[349]))&BiasedRNG[29])|(((m[42]&m[346]&m[347]&~m[348]&~m[349])|(m[42]&m[346]&~m[347]&m[348]&~m[349])|(m[42]&~m[346]&m[347]&m[348]&~m[349])|(~m[42]&m[346]&m[347]&m[348]&~m[349])|(m[42]&m[346]&~m[347]&~m[348]&m[349])|(m[42]&~m[346]&m[347]&~m[348]&m[349])|(~m[42]&m[346]&m[347]&~m[348]&m[349])|(m[42]&~m[346]&~m[347]&m[348]&m[349])|(~m[42]&m[346]&~m[347]&m[348]&m[349])|(~m[42]&~m[346]&m[347]&m[348]&m[349]))&~BiasedRNG[29])|((m[42]&m[346]&m[347]&m[348]&~m[349])|(m[42]&m[346]&m[347]&~m[348]&m[349])|(m[42]&m[346]&~m[347]&m[348]&m[349])|(m[42]&~m[346]&m[347]&m[348]&m[349])|(~m[42]&m[346]&m[347]&m[348]&m[349])|(m[42]&m[346]&m[347]&m[348]&m[349]));
    m[102] = (((m[43]&m[356]&~m[357]&~m[358]&~m[359])|(m[43]&~m[356]&m[357]&~m[358]&~m[359])|(~m[43]&m[356]&m[357]&~m[358]&~m[359])|(m[43]&~m[356]&~m[357]&m[358]&~m[359])|(~m[43]&m[356]&~m[357]&m[358]&~m[359])|(~m[43]&~m[356]&m[357]&m[358]&~m[359])|(m[43]&~m[356]&~m[357]&~m[358]&m[359])|(~m[43]&m[356]&~m[357]&~m[358]&m[359])|(~m[43]&~m[356]&m[357]&~m[358]&m[359])|(~m[43]&~m[356]&~m[357]&m[358]&m[359]))&BiasedRNG[30])|(((m[43]&m[356]&m[357]&~m[358]&~m[359])|(m[43]&m[356]&~m[357]&m[358]&~m[359])|(m[43]&~m[356]&m[357]&m[358]&~m[359])|(~m[43]&m[356]&m[357]&m[358]&~m[359])|(m[43]&m[356]&~m[357]&~m[358]&m[359])|(m[43]&~m[356]&m[357]&~m[358]&m[359])|(~m[43]&m[356]&m[357]&~m[358]&m[359])|(m[43]&~m[356]&~m[357]&m[358]&m[359])|(~m[43]&m[356]&~m[357]&m[358]&m[359])|(~m[43]&~m[356]&m[357]&m[358]&m[359]))&~BiasedRNG[30])|((m[43]&m[356]&m[357]&m[358]&~m[359])|(m[43]&m[356]&m[357]&~m[358]&m[359])|(m[43]&m[356]&~m[357]&m[358]&m[359])|(m[43]&~m[356]&m[357]&m[358]&m[359])|(~m[43]&m[356]&m[357]&m[358]&m[359])|(m[43]&m[356]&m[357]&m[358]&m[359]));
    m[103] = (((m[43]&m[360]&~m[361]&~m[362]&~m[363])|(m[43]&~m[360]&m[361]&~m[362]&~m[363])|(~m[43]&m[360]&m[361]&~m[362]&~m[363])|(m[43]&~m[360]&~m[361]&m[362]&~m[363])|(~m[43]&m[360]&~m[361]&m[362]&~m[363])|(~m[43]&~m[360]&m[361]&m[362]&~m[363])|(m[43]&~m[360]&~m[361]&~m[362]&m[363])|(~m[43]&m[360]&~m[361]&~m[362]&m[363])|(~m[43]&~m[360]&m[361]&~m[362]&m[363])|(~m[43]&~m[360]&~m[361]&m[362]&m[363]))&BiasedRNG[31])|(((m[43]&m[360]&m[361]&~m[362]&~m[363])|(m[43]&m[360]&~m[361]&m[362]&~m[363])|(m[43]&~m[360]&m[361]&m[362]&~m[363])|(~m[43]&m[360]&m[361]&m[362]&~m[363])|(m[43]&m[360]&~m[361]&~m[362]&m[363])|(m[43]&~m[360]&m[361]&~m[362]&m[363])|(~m[43]&m[360]&m[361]&~m[362]&m[363])|(m[43]&~m[360]&~m[361]&m[362]&m[363])|(~m[43]&m[360]&~m[361]&m[362]&m[363])|(~m[43]&~m[360]&m[361]&m[362]&m[363]))&~BiasedRNG[31])|((m[43]&m[360]&m[361]&m[362]&~m[363])|(m[43]&m[360]&m[361]&~m[362]&m[363])|(m[43]&m[360]&~m[361]&m[362]&m[363])|(m[43]&~m[360]&m[361]&m[362]&m[363])|(~m[43]&m[360]&m[361]&m[362]&m[363])|(m[43]&m[360]&m[361]&m[362]&m[363]));
    m[105] = (((m[44]&m[370]&~m[371]&~m[372]&~m[373])|(m[44]&~m[370]&m[371]&~m[372]&~m[373])|(~m[44]&m[370]&m[371]&~m[372]&~m[373])|(m[44]&~m[370]&~m[371]&m[372]&~m[373])|(~m[44]&m[370]&~m[371]&m[372]&~m[373])|(~m[44]&~m[370]&m[371]&m[372]&~m[373])|(m[44]&~m[370]&~m[371]&~m[372]&m[373])|(~m[44]&m[370]&~m[371]&~m[372]&m[373])|(~m[44]&~m[370]&m[371]&~m[372]&m[373])|(~m[44]&~m[370]&~m[371]&m[372]&m[373]))&BiasedRNG[32])|(((m[44]&m[370]&m[371]&~m[372]&~m[373])|(m[44]&m[370]&~m[371]&m[372]&~m[373])|(m[44]&~m[370]&m[371]&m[372]&~m[373])|(~m[44]&m[370]&m[371]&m[372]&~m[373])|(m[44]&m[370]&~m[371]&~m[372]&m[373])|(m[44]&~m[370]&m[371]&~m[372]&m[373])|(~m[44]&m[370]&m[371]&~m[372]&m[373])|(m[44]&~m[370]&~m[371]&m[372]&m[373])|(~m[44]&m[370]&~m[371]&m[372]&m[373])|(~m[44]&~m[370]&m[371]&m[372]&m[373]))&~BiasedRNG[32])|((m[44]&m[370]&m[371]&m[372]&~m[373])|(m[44]&m[370]&m[371]&~m[372]&m[373])|(m[44]&m[370]&~m[371]&m[372]&m[373])|(m[44]&~m[370]&m[371]&m[372]&m[373])|(~m[44]&m[370]&m[371]&m[372]&m[373])|(m[44]&m[370]&m[371]&m[372]&m[373]));
    m[106] = (((m[44]&m[374]&~m[375]&~m[376]&~m[377])|(m[44]&~m[374]&m[375]&~m[376]&~m[377])|(~m[44]&m[374]&m[375]&~m[376]&~m[377])|(m[44]&~m[374]&~m[375]&m[376]&~m[377])|(~m[44]&m[374]&~m[375]&m[376]&~m[377])|(~m[44]&~m[374]&m[375]&m[376]&~m[377])|(m[44]&~m[374]&~m[375]&~m[376]&m[377])|(~m[44]&m[374]&~m[375]&~m[376]&m[377])|(~m[44]&~m[374]&m[375]&~m[376]&m[377])|(~m[44]&~m[374]&~m[375]&m[376]&m[377]))&BiasedRNG[33])|(((m[44]&m[374]&m[375]&~m[376]&~m[377])|(m[44]&m[374]&~m[375]&m[376]&~m[377])|(m[44]&~m[374]&m[375]&m[376]&~m[377])|(~m[44]&m[374]&m[375]&m[376]&~m[377])|(m[44]&m[374]&~m[375]&~m[376]&m[377])|(m[44]&~m[374]&m[375]&~m[376]&m[377])|(~m[44]&m[374]&m[375]&~m[376]&m[377])|(m[44]&~m[374]&~m[375]&m[376]&m[377])|(~m[44]&m[374]&~m[375]&m[376]&m[377])|(~m[44]&~m[374]&m[375]&m[376]&m[377]))&~BiasedRNG[33])|((m[44]&m[374]&m[375]&m[376]&~m[377])|(m[44]&m[374]&m[375]&~m[376]&m[377])|(m[44]&m[374]&~m[375]&m[376]&m[377])|(m[44]&~m[374]&m[375]&m[376]&m[377])|(~m[44]&m[374]&m[375]&m[376]&m[377])|(m[44]&m[374]&m[375]&m[376]&m[377]));
    m[108] = (((m[45]&m[384]&~m[385]&~m[386]&~m[387])|(m[45]&~m[384]&m[385]&~m[386]&~m[387])|(~m[45]&m[384]&m[385]&~m[386]&~m[387])|(m[45]&~m[384]&~m[385]&m[386]&~m[387])|(~m[45]&m[384]&~m[385]&m[386]&~m[387])|(~m[45]&~m[384]&m[385]&m[386]&~m[387])|(m[45]&~m[384]&~m[385]&~m[386]&m[387])|(~m[45]&m[384]&~m[385]&~m[386]&m[387])|(~m[45]&~m[384]&m[385]&~m[386]&m[387])|(~m[45]&~m[384]&~m[385]&m[386]&m[387]))&BiasedRNG[34])|(((m[45]&m[384]&m[385]&~m[386]&~m[387])|(m[45]&m[384]&~m[385]&m[386]&~m[387])|(m[45]&~m[384]&m[385]&m[386]&~m[387])|(~m[45]&m[384]&m[385]&m[386]&~m[387])|(m[45]&m[384]&~m[385]&~m[386]&m[387])|(m[45]&~m[384]&m[385]&~m[386]&m[387])|(~m[45]&m[384]&m[385]&~m[386]&m[387])|(m[45]&~m[384]&~m[385]&m[386]&m[387])|(~m[45]&m[384]&~m[385]&m[386]&m[387])|(~m[45]&~m[384]&m[385]&m[386]&m[387]))&~BiasedRNG[34])|((m[45]&m[384]&m[385]&m[386]&~m[387])|(m[45]&m[384]&m[385]&~m[386]&m[387])|(m[45]&m[384]&~m[385]&m[386]&m[387])|(m[45]&~m[384]&m[385]&m[386]&m[387])|(~m[45]&m[384]&m[385]&m[386]&m[387])|(m[45]&m[384]&m[385]&m[386]&m[387]));
    m[109] = (((m[45]&m[388]&~m[389]&~m[390]&~m[391])|(m[45]&~m[388]&m[389]&~m[390]&~m[391])|(~m[45]&m[388]&m[389]&~m[390]&~m[391])|(m[45]&~m[388]&~m[389]&m[390]&~m[391])|(~m[45]&m[388]&~m[389]&m[390]&~m[391])|(~m[45]&~m[388]&m[389]&m[390]&~m[391])|(m[45]&~m[388]&~m[389]&~m[390]&m[391])|(~m[45]&m[388]&~m[389]&~m[390]&m[391])|(~m[45]&~m[388]&m[389]&~m[390]&m[391])|(~m[45]&~m[388]&~m[389]&m[390]&m[391]))&BiasedRNG[35])|(((m[45]&m[388]&m[389]&~m[390]&~m[391])|(m[45]&m[388]&~m[389]&m[390]&~m[391])|(m[45]&~m[388]&m[389]&m[390]&~m[391])|(~m[45]&m[388]&m[389]&m[390]&~m[391])|(m[45]&m[388]&~m[389]&~m[390]&m[391])|(m[45]&~m[388]&m[389]&~m[390]&m[391])|(~m[45]&m[388]&m[389]&~m[390]&m[391])|(m[45]&~m[388]&~m[389]&m[390]&m[391])|(~m[45]&m[388]&~m[389]&m[390]&m[391])|(~m[45]&~m[388]&m[389]&m[390]&m[391]))&~BiasedRNG[35])|((m[45]&m[388]&m[389]&m[390]&~m[391])|(m[45]&m[388]&m[389]&~m[390]&m[391])|(m[45]&m[388]&~m[389]&m[390]&m[391])|(m[45]&~m[388]&m[389]&m[390]&m[391])|(~m[45]&m[388]&m[389]&m[390]&m[391])|(m[45]&m[388]&m[389]&m[390]&m[391]));
    m[111] = (((m[46]&m[398]&~m[399]&~m[400]&~m[401])|(m[46]&~m[398]&m[399]&~m[400]&~m[401])|(~m[46]&m[398]&m[399]&~m[400]&~m[401])|(m[46]&~m[398]&~m[399]&m[400]&~m[401])|(~m[46]&m[398]&~m[399]&m[400]&~m[401])|(~m[46]&~m[398]&m[399]&m[400]&~m[401])|(m[46]&~m[398]&~m[399]&~m[400]&m[401])|(~m[46]&m[398]&~m[399]&~m[400]&m[401])|(~m[46]&~m[398]&m[399]&~m[400]&m[401])|(~m[46]&~m[398]&~m[399]&m[400]&m[401]))&BiasedRNG[36])|(((m[46]&m[398]&m[399]&~m[400]&~m[401])|(m[46]&m[398]&~m[399]&m[400]&~m[401])|(m[46]&~m[398]&m[399]&m[400]&~m[401])|(~m[46]&m[398]&m[399]&m[400]&~m[401])|(m[46]&m[398]&~m[399]&~m[400]&m[401])|(m[46]&~m[398]&m[399]&~m[400]&m[401])|(~m[46]&m[398]&m[399]&~m[400]&m[401])|(m[46]&~m[398]&~m[399]&m[400]&m[401])|(~m[46]&m[398]&~m[399]&m[400]&m[401])|(~m[46]&~m[398]&m[399]&m[400]&m[401]))&~BiasedRNG[36])|((m[46]&m[398]&m[399]&m[400]&~m[401])|(m[46]&m[398]&m[399]&~m[400]&m[401])|(m[46]&m[398]&~m[399]&m[400]&m[401])|(m[46]&~m[398]&m[399]&m[400]&m[401])|(~m[46]&m[398]&m[399]&m[400]&m[401])|(m[46]&m[398]&m[399]&m[400]&m[401]));
    m[112] = (((m[46]&m[402]&~m[403]&~m[404]&~m[405])|(m[46]&~m[402]&m[403]&~m[404]&~m[405])|(~m[46]&m[402]&m[403]&~m[404]&~m[405])|(m[46]&~m[402]&~m[403]&m[404]&~m[405])|(~m[46]&m[402]&~m[403]&m[404]&~m[405])|(~m[46]&~m[402]&m[403]&m[404]&~m[405])|(m[46]&~m[402]&~m[403]&~m[404]&m[405])|(~m[46]&m[402]&~m[403]&~m[404]&m[405])|(~m[46]&~m[402]&m[403]&~m[404]&m[405])|(~m[46]&~m[402]&~m[403]&m[404]&m[405]))&BiasedRNG[37])|(((m[46]&m[402]&m[403]&~m[404]&~m[405])|(m[46]&m[402]&~m[403]&m[404]&~m[405])|(m[46]&~m[402]&m[403]&m[404]&~m[405])|(~m[46]&m[402]&m[403]&m[404]&~m[405])|(m[46]&m[402]&~m[403]&~m[404]&m[405])|(m[46]&~m[402]&m[403]&~m[404]&m[405])|(~m[46]&m[402]&m[403]&~m[404]&m[405])|(m[46]&~m[402]&~m[403]&m[404]&m[405])|(~m[46]&m[402]&~m[403]&m[404]&m[405])|(~m[46]&~m[402]&m[403]&m[404]&m[405]))&~BiasedRNG[37])|((m[46]&m[402]&m[403]&m[404]&~m[405])|(m[46]&m[402]&m[403]&~m[404]&m[405])|(m[46]&m[402]&~m[403]&m[404]&m[405])|(m[46]&~m[402]&m[403]&m[404]&m[405])|(~m[46]&m[402]&m[403]&m[404]&m[405])|(m[46]&m[402]&m[403]&m[404]&m[405]));
    m[114] = (((m[47]&m[412]&~m[413]&~m[414]&~m[415])|(m[47]&~m[412]&m[413]&~m[414]&~m[415])|(~m[47]&m[412]&m[413]&~m[414]&~m[415])|(m[47]&~m[412]&~m[413]&m[414]&~m[415])|(~m[47]&m[412]&~m[413]&m[414]&~m[415])|(~m[47]&~m[412]&m[413]&m[414]&~m[415])|(m[47]&~m[412]&~m[413]&~m[414]&m[415])|(~m[47]&m[412]&~m[413]&~m[414]&m[415])|(~m[47]&~m[412]&m[413]&~m[414]&m[415])|(~m[47]&~m[412]&~m[413]&m[414]&m[415]))&BiasedRNG[38])|(((m[47]&m[412]&m[413]&~m[414]&~m[415])|(m[47]&m[412]&~m[413]&m[414]&~m[415])|(m[47]&~m[412]&m[413]&m[414]&~m[415])|(~m[47]&m[412]&m[413]&m[414]&~m[415])|(m[47]&m[412]&~m[413]&~m[414]&m[415])|(m[47]&~m[412]&m[413]&~m[414]&m[415])|(~m[47]&m[412]&m[413]&~m[414]&m[415])|(m[47]&~m[412]&~m[413]&m[414]&m[415])|(~m[47]&m[412]&~m[413]&m[414]&m[415])|(~m[47]&~m[412]&m[413]&m[414]&m[415]))&~BiasedRNG[38])|((m[47]&m[412]&m[413]&m[414]&~m[415])|(m[47]&m[412]&m[413]&~m[414]&m[415])|(m[47]&m[412]&~m[413]&m[414]&m[415])|(m[47]&~m[412]&m[413]&m[414]&m[415])|(~m[47]&m[412]&m[413]&m[414]&m[415])|(m[47]&m[412]&m[413]&m[414]&m[415]));
    m[115] = (((m[47]&m[416]&~m[417]&~m[418]&~m[419])|(m[47]&~m[416]&m[417]&~m[418]&~m[419])|(~m[47]&m[416]&m[417]&~m[418]&~m[419])|(m[47]&~m[416]&~m[417]&m[418]&~m[419])|(~m[47]&m[416]&~m[417]&m[418]&~m[419])|(~m[47]&~m[416]&m[417]&m[418]&~m[419])|(m[47]&~m[416]&~m[417]&~m[418]&m[419])|(~m[47]&m[416]&~m[417]&~m[418]&m[419])|(~m[47]&~m[416]&m[417]&~m[418]&m[419])|(~m[47]&~m[416]&~m[417]&m[418]&m[419]))&BiasedRNG[39])|(((m[47]&m[416]&m[417]&~m[418]&~m[419])|(m[47]&m[416]&~m[417]&m[418]&~m[419])|(m[47]&~m[416]&m[417]&m[418]&~m[419])|(~m[47]&m[416]&m[417]&m[418]&~m[419])|(m[47]&m[416]&~m[417]&~m[418]&m[419])|(m[47]&~m[416]&m[417]&~m[418]&m[419])|(~m[47]&m[416]&m[417]&~m[418]&m[419])|(m[47]&~m[416]&~m[417]&m[418]&m[419])|(~m[47]&m[416]&~m[417]&m[418]&m[419])|(~m[47]&~m[416]&m[417]&m[418]&m[419]))&~BiasedRNG[39])|((m[47]&m[416]&m[417]&m[418]&~m[419])|(m[47]&m[416]&m[417]&~m[418]&m[419])|(m[47]&m[416]&~m[417]&m[418]&m[419])|(m[47]&~m[416]&m[417]&m[418]&m[419])|(~m[47]&m[416]&m[417]&m[418]&m[419])|(m[47]&m[416]&m[417]&m[418]&m[419]));
    m[117] = (((m[48]&m[426]&~m[427]&~m[428]&~m[429])|(m[48]&~m[426]&m[427]&~m[428]&~m[429])|(~m[48]&m[426]&m[427]&~m[428]&~m[429])|(m[48]&~m[426]&~m[427]&m[428]&~m[429])|(~m[48]&m[426]&~m[427]&m[428]&~m[429])|(~m[48]&~m[426]&m[427]&m[428]&~m[429])|(m[48]&~m[426]&~m[427]&~m[428]&m[429])|(~m[48]&m[426]&~m[427]&~m[428]&m[429])|(~m[48]&~m[426]&m[427]&~m[428]&m[429])|(~m[48]&~m[426]&~m[427]&m[428]&m[429]))&BiasedRNG[40])|(((m[48]&m[426]&m[427]&~m[428]&~m[429])|(m[48]&m[426]&~m[427]&m[428]&~m[429])|(m[48]&~m[426]&m[427]&m[428]&~m[429])|(~m[48]&m[426]&m[427]&m[428]&~m[429])|(m[48]&m[426]&~m[427]&~m[428]&m[429])|(m[48]&~m[426]&m[427]&~m[428]&m[429])|(~m[48]&m[426]&m[427]&~m[428]&m[429])|(m[48]&~m[426]&~m[427]&m[428]&m[429])|(~m[48]&m[426]&~m[427]&m[428]&m[429])|(~m[48]&~m[426]&m[427]&m[428]&m[429]))&~BiasedRNG[40])|((m[48]&m[426]&m[427]&m[428]&~m[429])|(m[48]&m[426]&m[427]&~m[428]&m[429])|(m[48]&m[426]&~m[427]&m[428]&m[429])|(m[48]&~m[426]&m[427]&m[428]&m[429])|(~m[48]&m[426]&m[427]&m[428]&m[429])|(m[48]&m[426]&m[427]&m[428]&m[429]));
    m[118] = (((m[48]&m[430]&~m[431]&~m[432]&~m[433])|(m[48]&~m[430]&m[431]&~m[432]&~m[433])|(~m[48]&m[430]&m[431]&~m[432]&~m[433])|(m[48]&~m[430]&~m[431]&m[432]&~m[433])|(~m[48]&m[430]&~m[431]&m[432]&~m[433])|(~m[48]&~m[430]&m[431]&m[432]&~m[433])|(m[48]&~m[430]&~m[431]&~m[432]&m[433])|(~m[48]&m[430]&~m[431]&~m[432]&m[433])|(~m[48]&~m[430]&m[431]&~m[432]&m[433])|(~m[48]&~m[430]&~m[431]&m[432]&m[433]))&BiasedRNG[41])|(((m[48]&m[430]&m[431]&~m[432]&~m[433])|(m[48]&m[430]&~m[431]&m[432]&~m[433])|(m[48]&~m[430]&m[431]&m[432]&~m[433])|(~m[48]&m[430]&m[431]&m[432]&~m[433])|(m[48]&m[430]&~m[431]&~m[432]&m[433])|(m[48]&~m[430]&m[431]&~m[432]&m[433])|(~m[48]&m[430]&m[431]&~m[432]&m[433])|(m[48]&~m[430]&~m[431]&m[432]&m[433])|(~m[48]&m[430]&~m[431]&m[432]&m[433])|(~m[48]&~m[430]&m[431]&m[432]&m[433]))&~BiasedRNG[41])|((m[48]&m[430]&m[431]&m[432]&~m[433])|(m[48]&m[430]&m[431]&~m[432]&m[433])|(m[48]&m[430]&~m[431]&m[432]&m[433])|(m[48]&~m[430]&m[431]&m[432]&m[433])|(~m[48]&m[430]&m[431]&m[432]&m[433])|(m[48]&m[430]&m[431]&m[432]&m[433]));
    m[120] = (((m[49]&m[440]&~m[441]&~m[442]&~m[443])|(m[49]&~m[440]&m[441]&~m[442]&~m[443])|(~m[49]&m[440]&m[441]&~m[442]&~m[443])|(m[49]&~m[440]&~m[441]&m[442]&~m[443])|(~m[49]&m[440]&~m[441]&m[442]&~m[443])|(~m[49]&~m[440]&m[441]&m[442]&~m[443])|(m[49]&~m[440]&~m[441]&~m[442]&m[443])|(~m[49]&m[440]&~m[441]&~m[442]&m[443])|(~m[49]&~m[440]&m[441]&~m[442]&m[443])|(~m[49]&~m[440]&~m[441]&m[442]&m[443]))&BiasedRNG[42])|(((m[49]&m[440]&m[441]&~m[442]&~m[443])|(m[49]&m[440]&~m[441]&m[442]&~m[443])|(m[49]&~m[440]&m[441]&m[442]&~m[443])|(~m[49]&m[440]&m[441]&m[442]&~m[443])|(m[49]&m[440]&~m[441]&~m[442]&m[443])|(m[49]&~m[440]&m[441]&~m[442]&m[443])|(~m[49]&m[440]&m[441]&~m[442]&m[443])|(m[49]&~m[440]&~m[441]&m[442]&m[443])|(~m[49]&m[440]&~m[441]&m[442]&m[443])|(~m[49]&~m[440]&m[441]&m[442]&m[443]))&~BiasedRNG[42])|((m[49]&m[440]&m[441]&m[442]&~m[443])|(m[49]&m[440]&m[441]&~m[442]&m[443])|(m[49]&m[440]&~m[441]&m[442]&m[443])|(m[49]&~m[440]&m[441]&m[442]&m[443])|(~m[49]&m[440]&m[441]&m[442]&m[443])|(m[49]&m[440]&m[441]&m[442]&m[443]));
    m[121] = (((m[49]&m[444]&~m[445]&~m[446]&~m[447])|(m[49]&~m[444]&m[445]&~m[446]&~m[447])|(~m[49]&m[444]&m[445]&~m[446]&~m[447])|(m[49]&~m[444]&~m[445]&m[446]&~m[447])|(~m[49]&m[444]&~m[445]&m[446]&~m[447])|(~m[49]&~m[444]&m[445]&m[446]&~m[447])|(m[49]&~m[444]&~m[445]&~m[446]&m[447])|(~m[49]&m[444]&~m[445]&~m[446]&m[447])|(~m[49]&~m[444]&m[445]&~m[446]&m[447])|(~m[49]&~m[444]&~m[445]&m[446]&m[447]))&BiasedRNG[43])|(((m[49]&m[444]&m[445]&~m[446]&~m[447])|(m[49]&m[444]&~m[445]&m[446]&~m[447])|(m[49]&~m[444]&m[445]&m[446]&~m[447])|(~m[49]&m[444]&m[445]&m[446]&~m[447])|(m[49]&m[444]&~m[445]&~m[446]&m[447])|(m[49]&~m[444]&m[445]&~m[446]&m[447])|(~m[49]&m[444]&m[445]&~m[446]&m[447])|(m[49]&~m[444]&~m[445]&m[446]&m[447])|(~m[49]&m[444]&~m[445]&m[446]&m[447])|(~m[49]&~m[444]&m[445]&m[446]&m[447]))&~BiasedRNG[43])|((m[49]&m[444]&m[445]&m[446]&~m[447])|(m[49]&m[444]&m[445]&~m[446]&m[447])|(m[49]&m[444]&~m[445]&m[446]&m[447])|(m[49]&~m[444]&m[445]&m[446]&m[447])|(~m[49]&m[444]&m[445]&m[446]&m[447])|(m[49]&m[444]&m[445]&m[446]&m[447]));
    m[123] = (((m[50]&m[454]&~m[455]&~m[456]&~m[457])|(m[50]&~m[454]&m[455]&~m[456]&~m[457])|(~m[50]&m[454]&m[455]&~m[456]&~m[457])|(m[50]&~m[454]&~m[455]&m[456]&~m[457])|(~m[50]&m[454]&~m[455]&m[456]&~m[457])|(~m[50]&~m[454]&m[455]&m[456]&~m[457])|(m[50]&~m[454]&~m[455]&~m[456]&m[457])|(~m[50]&m[454]&~m[455]&~m[456]&m[457])|(~m[50]&~m[454]&m[455]&~m[456]&m[457])|(~m[50]&~m[454]&~m[455]&m[456]&m[457]))&BiasedRNG[44])|(((m[50]&m[454]&m[455]&~m[456]&~m[457])|(m[50]&m[454]&~m[455]&m[456]&~m[457])|(m[50]&~m[454]&m[455]&m[456]&~m[457])|(~m[50]&m[454]&m[455]&m[456]&~m[457])|(m[50]&m[454]&~m[455]&~m[456]&m[457])|(m[50]&~m[454]&m[455]&~m[456]&m[457])|(~m[50]&m[454]&m[455]&~m[456]&m[457])|(m[50]&~m[454]&~m[455]&m[456]&m[457])|(~m[50]&m[454]&~m[455]&m[456]&m[457])|(~m[50]&~m[454]&m[455]&m[456]&m[457]))&~BiasedRNG[44])|((m[50]&m[454]&m[455]&m[456]&~m[457])|(m[50]&m[454]&m[455]&~m[456]&m[457])|(m[50]&m[454]&~m[455]&m[456]&m[457])|(m[50]&~m[454]&m[455]&m[456]&m[457])|(~m[50]&m[454]&m[455]&m[456]&m[457])|(m[50]&m[454]&m[455]&m[456]&m[457]));
    m[124] = (((m[50]&m[458]&~m[459]&~m[460]&~m[461])|(m[50]&~m[458]&m[459]&~m[460]&~m[461])|(~m[50]&m[458]&m[459]&~m[460]&~m[461])|(m[50]&~m[458]&~m[459]&m[460]&~m[461])|(~m[50]&m[458]&~m[459]&m[460]&~m[461])|(~m[50]&~m[458]&m[459]&m[460]&~m[461])|(m[50]&~m[458]&~m[459]&~m[460]&m[461])|(~m[50]&m[458]&~m[459]&~m[460]&m[461])|(~m[50]&~m[458]&m[459]&~m[460]&m[461])|(~m[50]&~m[458]&~m[459]&m[460]&m[461]))&BiasedRNG[45])|(((m[50]&m[458]&m[459]&~m[460]&~m[461])|(m[50]&m[458]&~m[459]&m[460]&~m[461])|(m[50]&~m[458]&m[459]&m[460]&~m[461])|(~m[50]&m[458]&m[459]&m[460]&~m[461])|(m[50]&m[458]&~m[459]&~m[460]&m[461])|(m[50]&~m[458]&m[459]&~m[460]&m[461])|(~m[50]&m[458]&m[459]&~m[460]&m[461])|(m[50]&~m[458]&~m[459]&m[460]&m[461])|(~m[50]&m[458]&~m[459]&m[460]&m[461])|(~m[50]&~m[458]&m[459]&m[460]&m[461]))&~BiasedRNG[45])|((m[50]&m[458]&m[459]&m[460]&~m[461])|(m[50]&m[458]&m[459]&~m[460]&m[461])|(m[50]&m[458]&~m[459]&m[460]&m[461])|(m[50]&~m[458]&m[459]&m[460]&m[461])|(~m[50]&m[458]&m[459]&m[460]&m[461])|(m[50]&m[458]&m[459]&m[460]&m[461]));
    m[126] = (((m[51]&m[468]&~m[469]&~m[470]&~m[471])|(m[51]&~m[468]&m[469]&~m[470]&~m[471])|(~m[51]&m[468]&m[469]&~m[470]&~m[471])|(m[51]&~m[468]&~m[469]&m[470]&~m[471])|(~m[51]&m[468]&~m[469]&m[470]&~m[471])|(~m[51]&~m[468]&m[469]&m[470]&~m[471])|(m[51]&~m[468]&~m[469]&~m[470]&m[471])|(~m[51]&m[468]&~m[469]&~m[470]&m[471])|(~m[51]&~m[468]&m[469]&~m[470]&m[471])|(~m[51]&~m[468]&~m[469]&m[470]&m[471]))&BiasedRNG[46])|(((m[51]&m[468]&m[469]&~m[470]&~m[471])|(m[51]&m[468]&~m[469]&m[470]&~m[471])|(m[51]&~m[468]&m[469]&m[470]&~m[471])|(~m[51]&m[468]&m[469]&m[470]&~m[471])|(m[51]&m[468]&~m[469]&~m[470]&m[471])|(m[51]&~m[468]&m[469]&~m[470]&m[471])|(~m[51]&m[468]&m[469]&~m[470]&m[471])|(m[51]&~m[468]&~m[469]&m[470]&m[471])|(~m[51]&m[468]&~m[469]&m[470]&m[471])|(~m[51]&~m[468]&m[469]&m[470]&m[471]))&~BiasedRNG[46])|((m[51]&m[468]&m[469]&m[470]&~m[471])|(m[51]&m[468]&m[469]&~m[470]&m[471])|(m[51]&m[468]&~m[469]&m[470]&m[471])|(m[51]&~m[468]&m[469]&m[470]&m[471])|(~m[51]&m[468]&m[469]&m[470]&m[471])|(m[51]&m[468]&m[469]&m[470]&m[471]));
    m[127] = (((m[51]&m[472]&~m[473]&~m[474]&~m[475])|(m[51]&~m[472]&m[473]&~m[474]&~m[475])|(~m[51]&m[472]&m[473]&~m[474]&~m[475])|(m[51]&~m[472]&~m[473]&m[474]&~m[475])|(~m[51]&m[472]&~m[473]&m[474]&~m[475])|(~m[51]&~m[472]&m[473]&m[474]&~m[475])|(m[51]&~m[472]&~m[473]&~m[474]&m[475])|(~m[51]&m[472]&~m[473]&~m[474]&m[475])|(~m[51]&~m[472]&m[473]&~m[474]&m[475])|(~m[51]&~m[472]&~m[473]&m[474]&m[475]))&BiasedRNG[47])|(((m[51]&m[472]&m[473]&~m[474]&~m[475])|(m[51]&m[472]&~m[473]&m[474]&~m[475])|(m[51]&~m[472]&m[473]&m[474]&~m[475])|(~m[51]&m[472]&m[473]&m[474]&~m[475])|(m[51]&m[472]&~m[473]&~m[474]&m[475])|(m[51]&~m[472]&m[473]&~m[474]&m[475])|(~m[51]&m[472]&m[473]&~m[474]&m[475])|(m[51]&~m[472]&~m[473]&m[474]&m[475])|(~m[51]&m[472]&~m[473]&m[474]&m[475])|(~m[51]&~m[472]&m[473]&m[474]&m[475]))&~BiasedRNG[47])|((m[51]&m[472]&m[473]&m[474]&~m[475])|(m[51]&m[472]&m[473]&~m[474]&m[475])|(m[51]&m[472]&~m[473]&m[474]&m[475])|(m[51]&~m[472]&m[473]&m[474]&m[475])|(~m[51]&m[472]&m[473]&m[474]&m[475])|(m[51]&m[472]&m[473]&m[474]&m[475]));
    m[129] = (((m[52]&m[482]&~m[483]&~m[484]&~m[485])|(m[52]&~m[482]&m[483]&~m[484]&~m[485])|(~m[52]&m[482]&m[483]&~m[484]&~m[485])|(m[52]&~m[482]&~m[483]&m[484]&~m[485])|(~m[52]&m[482]&~m[483]&m[484]&~m[485])|(~m[52]&~m[482]&m[483]&m[484]&~m[485])|(m[52]&~m[482]&~m[483]&~m[484]&m[485])|(~m[52]&m[482]&~m[483]&~m[484]&m[485])|(~m[52]&~m[482]&m[483]&~m[484]&m[485])|(~m[52]&~m[482]&~m[483]&m[484]&m[485]))&BiasedRNG[48])|(((m[52]&m[482]&m[483]&~m[484]&~m[485])|(m[52]&m[482]&~m[483]&m[484]&~m[485])|(m[52]&~m[482]&m[483]&m[484]&~m[485])|(~m[52]&m[482]&m[483]&m[484]&~m[485])|(m[52]&m[482]&~m[483]&~m[484]&m[485])|(m[52]&~m[482]&m[483]&~m[484]&m[485])|(~m[52]&m[482]&m[483]&~m[484]&m[485])|(m[52]&~m[482]&~m[483]&m[484]&m[485])|(~m[52]&m[482]&~m[483]&m[484]&m[485])|(~m[52]&~m[482]&m[483]&m[484]&m[485]))&~BiasedRNG[48])|((m[52]&m[482]&m[483]&m[484]&~m[485])|(m[52]&m[482]&m[483]&~m[484]&m[485])|(m[52]&m[482]&~m[483]&m[484]&m[485])|(m[52]&~m[482]&m[483]&m[484]&m[485])|(~m[52]&m[482]&m[483]&m[484]&m[485])|(m[52]&m[482]&m[483]&m[484]&m[485]));
    m[130] = (((m[52]&m[486]&~m[487]&~m[488]&~m[489])|(m[52]&~m[486]&m[487]&~m[488]&~m[489])|(~m[52]&m[486]&m[487]&~m[488]&~m[489])|(m[52]&~m[486]&~m[487]&m[488]&~m[489])|(~m[52]&m[486]&~m[487]&m[488]&~m[489])|(~m[52]&~m[486]&m[487]&m[488]&~m[489])|(m[52]&~m[486]&~m[487]&~m[488]&m[489])|(~m[52]&m[486]&~m[487]&~m[488]&m[489])|(~m[52]&~m[486]&m[487]&~m[488]&m[489])|(~m[52]&~m[486]&~m[487]&m[488]&m[489]))&BiasedRNG[49])|(((m[52]&m[486]&m[487]&~m[488]&~m[489])|(m[52]&m[486]&~m[487]&m[488]&~m[489])|(m[52]&~m[486]&m[487]&m[488]&~m[489])|(~m[52]&m[486]&m[487]&m[488]&~m[489])|(m[52]&m[486]&~m[487]&~m[488]&m[489])|(m[52]&~m[486]&m[487]&~m[488]&m[489])|(~m[52]&m[486]&m[487]&~m[488]&m[489])|(m[52]&~m[486]&~m[487]&m[488]&m[489])|(~m[52]&m[486]&~m[487]&m[488]&m[489])|(~m[52]&~m[486]&m[487]&m[488]&m[489]))&~BiasedRNG[49])|((m[52]&m[486]&m[487]&m[488]&~m[489])|(m[52]&m[486]&m[487]&~m[488]&m[489])|(m[52]&m[486]&~m[487]&m[488]&m[489])|(m[52]&~m[486]&m[487]&m[488]&m[489])|(~m[52]&m[486]&m[487]&m[488]&m[489])|(m[52]&m[486]&m[487]&m[488]&m[489]));
    m[132] = (((m[53]&m[496]&~m[497]&~m[498]&~m[499])|(m[53]&~m[496]&m[497]&~m[498]&~m[499])|(~m[53]&m[496]&m[497]&~m[498]&~m[499])|(m[53]&~m[496]&~m[497]&m[498]&~m[499])|(~m[53]&m[496]&~m[497]&m[498]&~m[499])|(~m[53]&~m[496]&m[497]&m[498]&~m[499])|(m[53]&~m[496]&~m[497]&~m[498]&m[499])|(~m[53]&m[496]&~m[497]&~m[498]&m[499])|(~m[53]&~m[496]&m[497]&~m[498]&m[499])|(~m[53]&~m[496]&~m[497]&m[498]&m[499]))&BiasedRNG[50])|(((m[53]&m[496]&m[497]&~m[498]&~m[499])|(m[53]&m[496]&~m[497]&m[498]&~m[499])|(m[53]&~m[496]&m[497]&m[498]&~m[499])|(~m[53]&m[496]&m[497]&m[498]&~m[499])|(m[53]&m[496]&~m[497]&~m[498]&m[499])|(m[53]&~m[496]&m[497]&~m[498]&m[499])|(~m[53]&m[496]&m[497]&~m[498]&m[499])|(m[53]&~m[496]&~m[497]&m[498]&m[499])|(~m[53]&m[496]&~m[497]&m[498]&m[499])|(~m[53]&~m[496]&m[497]&m[498]&m[499]))&~BiasedRNG[50])|((m[53]&m[496]&m[497]&m[498]&~m[499])|(m[53]&m[496]&m[497]&~m[498]&m[499])|(m[53]&m[496]&~m[497]&m[498]&m[499])|(m[53]&~m[496]&m[497]&m[498]&m[499])|(~m[53]&m[496]&m[497]&m[498]&m[499])|(m[53]&m[496]&m[497]&m[498]&m[499]));
    m[133] = (((m[53]&m[500]&~m[501]&~m[502]&~m[503])|(m[53]&~m[500]&m[501]&~m[502]&~m[503])|(~m[53]&m[500]&m[501]&~m[502]&~m[503])|(m[53]&~m[500]&~m[501]&m[502]&~m[503])|(~m[53]&m[500]&~m[501]&m[502]&~m[503])|(~m[53]&~m[500]&m[501]&m[502]&~m[503])|(m[53]&~m[500]&~m[501]&~m[502]&m[503])|(~m[53]&m[500]&~m[501]&~m[502]&m[503])|(~m[53]&~m[500]&m[501]&~m[502]&m[503])|(~m[53]&~m[500]&~m[501]&m[502]&m[503]))&BiasedRNG[51])|(((m[53]&m[500]&m[501]&~m[502]&~m[503])|(m[53]&m[500]&~m[501]&m[502]&~m[503])|(m[53]&~m[500]&m[501]&m[502]&~m[503])|(~m[53]&m[500]&m[501]&m[502]&~m[503])|(m[53]&m[500]&~m[501]&~m[502]&m[503])|(m[53]&~m[500]&m[501]&~m[502]&m[503])|(~m[53]&m[500]&m[501]&~m[502]&m[503])|(m[53]&~m[500]&~m[501]&m[502]&m[503])|(~m[53]&m[500]&~m[501]&m[502]&m[503])|(~m[53]&~m[500]&m[501]&m[502]&m[503]))&~BiasedRNG[51])|((m[53]&m[500]&m[501]&m[502]&~m[503])|(m[53]&m[500]&m[501]&~m[502]&m[503])|(m[53]&m[500]&~m[501]&m[502]&m[503])|(m[53]&~m[500]&m[501]&m[502]&m[503])|(~m[53]&m[500]&m[501]&m[502]&m[503])|(m[53]&m[500]&m[501]&m[502]&m[503]));
    m[135] = (((m[54]&m[510]&~m[511]&~m[512]&~m[513])|(m[54]&~m[510]&m[511]&~m[512]&~m[513])|(~m[54]&m[510]&m[511]&~m[512]&~m[513])|(m[54]&~m[510]&~m[511]&m[512]&~m[513])|(~m[54]&m[510]&~m[511]&m[512]&~m[513])|(~m[54]&~m[510]&m[511]&m[512]&~m[513])|(m[54]&~m[510]&~m[511]&~m[512]&m[513])|(~m[54]&m[510]&~m[511]&~m[512]&m[513])|(~m[54]&~m[510]&m[511]&~m[512]&m[513])|(~m[54]&~m[510]&~m[511]&m[512]&m[513]))&BiasedRNG[52])|(((m[54]&m[510]&m[511]&~m[512]&~m[513])|(m[54]&m[510]&~m[511]&m[512]&~m[513])|(m[54]&~m[510]&m[511]&m[512]&~m[513])|(~m[54]&m[510]&m[511]&m[512]&~m[513])|(m[54]&m[510]&~m[511]&~m[512]&m[513])|(m[54]&~m[510]&m[511]&~m[512]&m[513])|(~m[54]&m[510]&m[511]&~m[512]&m[513])|(m[54]&~m[510]&~m[511]&m[512]&m[513])|(~m[54]&m[510]&~m[511]&m[512]&m[513])|(~m[54]&~m[510]&m[511]&m[512]&m[513]))&~BiasedRNG[52])|((m[54]&m[510]&m[511]&m[512]&~m[513])|(m[54]&m[510]&m[511]&~m[512]&m[513])|(m[54]&m[510]&~m[511]&m[512]&m[513])|(m[54]&~m[510]&m[511]&m[512]&m[513])|(~m[54]&m[510]&m[511]&m[512]&m[513])|(m[54]&m[510]&m[511]&m[512]&m[513]));
    m[136] = (((m[54]&m[514]&~m[515]&~m[516]&~m[517])|(m[54]&~m[514]&m[515]&~m[516]&~m[517])|(~m[54]&m[514]&m[515]&~m[516]&~m[517])|(m[54]&~m[514]&~m[515]&m[516]&~m[517])|(~m[54]&m[514]&~m[515]&m[516]&~m[517])|(~m[54]&~m[514]&m[515]&m[516]&~m[517])|(m[54]&~m[514]&~m[515]&~m[516]&m[517])|(~m[54]&m[514]&~m[515]&~m[516]&m[517])|(~m[54]&~m[514]&m[515]&~m[516]&m[517])|(~m[54]&~m[514]&~m[515]&m[516]&m[517]))&BiasedRNG[53])|(((m[54]&m[514]&m[515]&~m[516]&~m[517])|(m[54]&m[514]&~m[515]&m[516]&~m[517])|(m[54]&~m[514]&m[515]&m[516]&~m[517])|(~m[54]&m[514]&m[515]&m[516]&~m[517])|(m[54]&m[514]&~m[515]&~m[516]&m[517])|(m[54]&~m[514]&m[515]&~m[516]&m[517])|(~m[54]&m[514]&m[515]&~m[516]&m[517])|(m[54]&~m[514]&~m[515]&m[516]&m[517])|(~m[54]&m[514]&~m[515]&m[516]&m[517])|(~m[54]&~m[514]&m[515]&m[516]&m[517]))&~BiasedRNG[53])|((m[54]&m[514]&m[515]&m[516]&~m[517])|(m[54]&m[514]&m[515]&~m[516]&m[517])|(m[54]&m[514]&~m[515]&m[516]&m[517])|(m[54]&~m[514]&m[515]&m[516]&m[517])|(~m[54]&m[514]&m[515]&m[516]&m[517])|(m[54]&m[514]&m[515]&m[516]&m[517]));
    m[138] = (((m[55]&m[524]&~m[525]&~m[526]&~m[527])|(m[55]&~m[524]&m[525]&~m[526]&~m[527])|(~m[55]&m[524]&m[525]&~m[526]&~m[527])|(m[55]&~m[524]&~m[525]&m[526]&~m[527])|(~m[55]&m[524]&~m[525]&m[526]&~m[527])|(~m[55]&~m[524]&m[525]&m[526]&~m[527])|(m[55]&~m[524]&~m[525]&~m[526]&m[527])|(~m[55]&m[524]&~m[525]&~m[526]&m[527])|(~m[55]&~m[524]&m[525]&~m[526]&m[527])|(~m[55]&~m[524]&~m[525]&m[526]&m[527]))&BiasedRNG[54])|(((m[55]&m[524]&m[525]&~m[526]&~m[527])|(m[55]&m[524]&~m[525]&m[526]&~m[527])|(m[55]&~m[524]&m[525]&m[526]&~m[527])|(~m[55]&m[524]&m[525]&m[526]&~m[527])|(m[55]&m[524]&~m[525]&~m[526]&m[527])|(m[55]&~m[524]&m[525]&~m[526]&m[527])|(~m[55]&m[524]&m[525]&~m[526]&m[527])|(m[55]&~m[524]&~m[525]&m[526]&m[527])|(~m[55]&m[524]&~m[525]&m[526]&m[527])|(~m[55]&~m[524]&m[525]&m[526]&m[527]))&~BiasedRNG[54])|((m[55]&m[524]&m[525]&m[526]&~m[527])|(m[55]&m[524]&m[525]&~m[526]&m[527])|(m[55]&m[524]&~m[525]&m[526]&m[527])|(m[55]&~m[524]&m[525]&m[526]&m[527])|(~m[55]&m[524]&m[525]&m[526]&m[527])|(m[55]&m[524]&m[525]&m[526]&m[527]));
    m[139] = (((m[55]&m[528]&~m[529]&~m[530]&~m[531])|(m[55]&~m[528]&m[529]&~m[530]&~m[531])|(~m[55]&m[528]&m[529]&~m[530]&~m[531])|(m[55]&~m[528]&~m[529]&m[530]&~m[531])|(~m[55]&m[528]&~m[529]&m[530]&~m[531])|(~m[55]&~m[528]&m[529]&m[530]&~m[531])|(m[55]&~m[528]&~m[529]&~m[530]&m[531])|(~m[55]&m[528]&~m[529]&~m[530]&m[531])|(~m[55]&~m[528]&m[529]&~m[530]&m[531])|(~m[55]&~m[528]&~m[529]&m[530]&m[531]))&BiasedRNG[55])|(((m[55]&m[528]&m[529]&~m[530]&~m[531])|(m[55]&m[528]&~m[529]&m[530]&~m[531])|(m[55]&~m[528]&m[529]&m[530]&~m[531])|(~m[55]&m[528]&m[529]&m[530]&~m[531])|(m[55]&m[528]&~m[529]&~m[530]&m[531])|(m[55]&~m[528]&m[529]&~m[530]&m[531])|(~m[55]&m[528]&m[529]&~m[530]&m[531])|(m[55]&~m[528]&~m[529]&m[530]&m[531])|(~m[55]&m[528]&~m[529]&m[530]&m[531])|(~m[55]&~m[528]&m[529]&m[530]&m[531]))&~BiasedRNG[55])|((m[55]&m[528]&m[529]&m[530]&~m[531])|(m[55]&m[528]&m[529]&~m[530]&m[531])|(m[55]&m[528]&~m[529]&m[530]&m[531])|(m[55]&~m[528]&m[529]&m[530]&m[531])|(~m[55]&m[528]&m[529]&m[530]&m[531])|(m[55]&m[528]&m[529]&m[530]&m[531]));
    m[140] = (((~m[28]&~m[336]&~m[532])|(m[28]&m[336]&~m[532]))&BiasedRNG[56])|(((m[28]&~m[336]&~m[532])|(~m[28]&m[336]&m[532]))&~BiasedRNG[56])|((~m[28]&~m[336]&m[532])|(m[28]&~m[336]&m[532])|(m[28]&m[336]&m[532]));
    m[141] = (((~m[28]&~m[350]&~m[546])|(m[28]&m[350]&~m[546]))&BiasedRNG[57])|(((m[28]&~m[350]&~m[546])|(~m[28]&m[350]&m[546]))&~BiasedRNG[57])|((~m[28]&~m[350]&m[546])|(m[28]&~m[350]&m[546])|(m[28]&m[350]&m[546]));
    m[142] = (((~m[56]&~m[364]&~m[560])|(m[56]&m[364]&~m[560]))&BiasedRNG[58])|(((m[56]&~m[364]&~m[560])|(~m[56]&m[364]&m[560]))&~BiasedRNG[58])|((~m[56]&~m[364]&m[560])|(m[56]&~m[364]&m[560])|(m[56]&m[364]&m[560]));
    m[143] = (((~m[56]&~m[378]&~m[574])|(m[56]&m[378]&~m[574]))&BiasedRNG[59])|(((m[56]&~m[378]&~m[574])|(~m[56]&m[378]&m[574]))&~BiasedRNG[59])|((~m[56]&~m[378]&m[574])|(m[56]&~m[378]&m[574])|(m[56]&m[378]&m[574]));
    m[144] = (((~m[56]&~m[392]&~m[588])|(m[56]&m[392]&~m[588]))&BiasedRNG[60])|(((m[56]&~m[392]&~m[588])|(~m[56]&m[392]&m[588]))&~BiasedRNG[60])|((~m[56]&~m[392]&m[588])|(m[56]&~m[392]&m[588])|(m[56]&m[392]&m[588]));
    m[145] = (((~m[56]&~m[406]&~m[602])|(m[56]&m[406]&~m[602]))&BiasedRNG[61])|(((m[56]&~m[406]&~m[602])|(~m[56]&m[406]&m[602]))&~BiasedRNG[61])|((~m[56]&~m[406]&m[602])|(m[56]&~m[406]&m[602])|(m[56]&m[406]&m[602]));
    m[154] = (((~m[29]&~m[337]&~m[533])|(m[29]&m[337]&~m[533]))&BiasedRNG[62])|(((m[29]&~m[337]&~m[533])|(~m[29]&m[337]&m[533]))&~BiasedRNG[62])|((~m[29]&~m[337]&m[533])|(m[29]&~m[337]&m[533])|(m[29]&m[337]&m[533]));
    m[155] = (((~m[29]&~m[351]&~m[547])|(m[29]&m[351]&~m[547]))&BiasedRNG[63])|(((m[29]&~m[351]&~m[547])|(~m[29]&m[351]&m[547]))&~BiasedRNG[63])|((~m[29]&~m[351]&m[547])|(m[29]&~m[351]&m[547])|(m[29]&m[351]&m[547]));
    m[156] = (((~m[59]&~m[365]&~m[561])|(m[59]&m[365]&~m[561]))&BiasedRNG[64])|(((m[59]&~m[365]&~m[561])|(~m[59]&m[365]&m[561]))&~BiasedRNG[64])|((~m[59]&~m[365]&m[561])|(m[59]&~m[365]&m[561])|(m[59]&m[365]&m[561]));
    m[157] = (((~m[59]&~m[379]&~m[575])|(m[59]&m[379]&~m[575]))&BiasedRNG[65])|(((m[59]&~m[379]&~m[575])|(~m[59]&m[379]&m[575]))&~BiasedRNG[65])|((~m[59]&~m[379]&m[575])|(m[59]&~m[379]&m[575])|(m[59]&m[379]&m[575]));
    m[158] = (((~m[59]&~m[393]&~m[589])|(m[59]&m[393]&~m[589]))&BiasedRNG[66])|(((m[59]&~m[393]&~m[589])|(~m[59]&m[393]&m[589]))&~BiasedRNG[66])|((~m[59]&~m[393]&m[589])|(m[59]&~m[393]&m[589])|(m[59]&m[393]&m[589]));
    m[159] = (((~m[59]&~m[407]&~m[603])|(m[59]&m[407]&~m[603]))&BiasedRNG[67])|(((m[59]&~m[407]&~m[603])|(~m[59]&m[407]&m[603]))&~BiasedRNG[67])|((~m[59]&~m[407]&m[603])|(m[59]&~m[407]&m[603])|(m[59]&m[407]&m[603]));
    m[168] = (((~m[30]&~m[338]&~m[534])|(m[30]&m[338]&~m[534]))&BiasedRNG[68])|(((m[30]&~m[338]&~m[534])|(~m[30]&m[338]&m[534]))&~BiasedRNG[68])|((~m[30]&~m[338]&m[534])|(m[30]&~m[338]&m[534])|(m[30]&m[338]&m[534]));
    m[169] = (((~m[30]&~m[352]&~m[548])|(m[30]&m[352]&~m[548]))&BiasedRNG[69])|(((m[30]&~m[352]&~m[548])|(~m[30]&m[352]&m[548]))&~BiasedRNG[69])|((~m[30]&~m[352]&m[548])|(m[30]&~m[352]&m[548])|(m[30]&m[352]&m[548]));
    m[170] = (((~m[62]&~m[366]&~m[562])|(m[62]&m[366]&~m[562]))&BiasedRNG[70])|(((m[62]&~m[366]&~m[562])|(~m[62]&m[366]&m[562]))&~BiasedRNG[70])|((~m[62]&~m[366]&m[562])|(m[62]&~m[366]&m[562])|(m[62]&m[366]&m[562]));
    m[171] = (((~m[62]&~m[380]&~m[576])|(m[62]&m[380]&~m[576]))&BiasedRNG[71])|(((m[62]&~m[380]&~m[576])|(~m[62]&m[380]&m[576]))&~BiasedRNG[71])|((~m[62]&~m[380]&m[576])|(m[62]&~m[380]&m[576])|(m[62]&m[380]&m[576]));
    m[172] = (((~m[62]&~m[394]&~m[590])|(m[62]&m[394]&~m[590]))&BiasedRNG[72])|(((m[62]&~m[394]&~m[590])|(~m[62]&m[394]&m[590]))&~BiasedRNG[72])|((~m[62]&~m[394]&m[590])|(m[62]&~m[394]&m[590])|(m[62]&m[394]&m[590]));
    m[173] = (((~m[62]&~m[408]&~m[604])|(m[62]&m[408]&~m[604]))&BiasedRNG[73])|(((m[62]&~m[408]&~m[604])|(~m[62]&m[408]&m[604]))&~BiasedRNG[73])|((~m[62]&~m[408]&m[604])|(m[62]&~m[408]&m[604])|(m[62]&m[408]&m[604]));
    m[182] = (((~m[31]&~m[339]&~m[535])|(m[31]&m[339]&~m[535]))&BiasedRNG[74])|(((m[31]&~m[339]&~m[535])|(~m[31]&m[339]&m[535]))&~BiasedRNG[74])|((~m[31]&~m[339]&m[535])|(m[31]&~m[339]&m[535])|(m[31]&m[339]&m[535]));
    m[183] = (((~m[31]&~m[353]&~m[549])|(m[31]&m[353]&~m[549]))&BiasedRNG[75])|(((m[31]&~m[353]&~m[549])|(~m[31]&m[353]&m[549]))&~BiasedRNG[75])|((~m[31]&~m[353]&m[549])|(m[31]&~m[353]&m[549])|(m[31]&m[353]&m[549]));
    m[184] = (((~m[65]&~m[367]&~m[563])|(m[65]&m[367]&~m[563]))&BiasedRNG[76])|(((m[65]&~m[367]&~m[563])|(~m[65]&m[367]&m[563]))&~BiasedRNG[76])|((~m[65]&~m[367]&m[563])|(m[65]&~m[367]&m[563])|(m[65]&m[367]&m[563]));
    m[185] = (((~m[65]&~m[381]&~m[577])|(m[65]&m[381]&~m[577]))&BiasedRNG[77])|(((m[65]&~m[381]&~m[577])|(~m[65]&m[381]&m[577]))&~BiasedRNG[77])|((~m[65]&~m[381]&m[577])|(m[65]&~m[381]&m[577])|(m[65]&m[381]&m[577]));
    m[186] = (((~m[65]&~m[395]&~m[591])|(m[65]&m[395]&~m[591]))&BiasedRNG[78])|(((m[65]&~m[395]&~m[591])|(~m[65]&m[395]&m[591]))&~BiasedRNG[78])|((~m[65]&~m[395]&m[591])|(m[65]&~m[395]&m[591])|(m[65]&m[395]&m[591]));
    m[187] = (((~m[65]&~m[409]&~m[605])|(m[65]&m[409]&~m[605]))&BiasedRNG[79])|(((m[65]&~m[409]&~m[605])|(~m[65]&m[409]&m[605]))&~BiasedRNG[79])|((~m[65]&~m[409]&m[605])|(m[65]&~m[409]&m[605])|(m[65]&m[409]&m[605]));
    m[196] = (((~m[32]&~m[340]&~m[536])|(m[32]&m[340]&~m[536]))&BiasedRNG[80])|(((m[32]&~m[340]&~m[536])|(~m[32]&m[340]&m[536]))&~BiasedRNG[80])|((~m[32]&~m[340]&m[536])|(m[32]&~m[340]&m[536])|(m[32]&m[340]&m[536]));
    m[197] = (((~m[32]&~m[354]&~m[550])|(m[32]&m[354]&~m[550]))&BiasedRNG[81])|(((m[32]&~m[354]&~m[550])|(~m[32]&m[354]&m[550]))&~BiasedRNG[81])|((~m[32]&~m[354]&m[550])|(m[32]&~m[354]&m[550])|(m[32]&m[354]&m[550]));
    m[198] = (((~m[68]&~m[368]&~m[564])|(m[68]&m[368]&~m[564]))&BiasedRNG[82])|(((m[68]&~m[368]&~m[564])|(~m[68]&m[368]&m[564]))&~BiasedRNG[82])|((~m[68]&~m[368]&m[564])|(m[68]&~m[368]&m[564])|(m[68]&m[368]&m[564]));
    m[199] = (((~m[68]&~m[382]&~m[578])|(m[68]&m[382]&~m[578]))&BiasedRNG[83])|(((m[68]&~m[382]&~m[578])|(~m[68]&m[382]&m[578]))&~BiasedRNG[83])|((~m[68]&~m[382]&m[578])|(m[68]&~m[382]&m[578])|(m[68]&m[382]&m[578]));
    m[200] = (((~m[68]&~m[396]&~m[592])|(m[68]&m[396]&~m[592]))&BiasedRNG[84])|(((m[68]&~m[396]&~m[592])|(~m[68]&m[396]&m[592]))&~BiasedRNG[84])|((~m[68]&~m[396]&m[592])|(m[68]&~m[396]&m[592])|(m[68]&m[396]&m[592]));
    m[201] = (((~m[68]&~m[410]&~m[606])|(m[68]&m[410]&~m[606]))&BiasedRNG[85])|(((m[68]&~m[410]&~m[606])|(~m[68]&m[410]&m[606]))&~BiasedRNG[85])|((~m[68]&~m[410]&m[606])|(m[68]&~m[410]&m[606])|(m[68]&m[410]&m[606]));
    m[210] = (((~m[33]&~m[341]&~m[537])|(m[33]&m[341]&~m[537]))&BiasedRNG[86])|(((m[33]&~m[341]&~m[537])|(~m[33]&m[341]&m[537]))&~BiasedRNG[86])|((~m[33]&~m[341]&m[537])|(m[33]&~m[341]&m[537])|(m[33]&m[341]&m[537]));
    m[211] = (((~m[33]&~m[355]&~m[551])|(m[33]&m[355]&~m[551]))&BiasedRNG[87])|(((m[33]&~m[355]&~m[551])|(~m[33]&m[355]&m[551]))&~BiasedRNG[87])|((~m[33]&~m[355]&m[551])|(m[33]&~m[355]&m[551])|(m[33]&m[355]&m[551]));
    m[212] = (((~m[71]&~m[369]&~m[565])|(m[71]&m[369]&~m[565]))&BiasedRNG[88])|(((m[71]&~m[369]&~m[565])|(~m[71]&m[369]&m[565]))&~BiasedRNG[88])|((~m[71]&~m[369]&m[565])|(m[71]&~m[369]&m[565])|(m[71]&m[369]&m[565]));
    m[213] = (((~m[71]&~m[383]&~m[579])|(m[71]&m[383]&~m[579]))&BiasedRNG[89])|(((m[71]&~m[383]&~m[579])|(~m[71]&m[383]&m[579]))&~BiasedRNG[89])|((~m[71]&~m[383]&m[579])|(m[71]&~m[383]&m[579])|(m[71]&m[383]&m[579]));
    m[214] = (((~m[71]&~m[397]&~m[593])|(m[71]&m[397]&~m[593]))&BiasedRNG[90])|(((m[71]&~m[397]&~m[593])|(~m[71]&m[397]&m[593]))&~BiasedRNG[90])|((~m[71]&~m[397]&m[593])|(m[71]&~m[397]&m[593])|(m[71]&m[397]&m[593]));
    m[215] = (((~m[71]&~m[411]&~m[607])|(m[71]&m[411]&~m[607]))&BiasedRNG[91])|(((m[71]&~m[411]&~m[607])|(~m[71]&m[411]&m[607]))&~BiasedRNG[91])|((~m[71]&~m[411]&m[607])|(m[71]&~m[411]&m[607])|(m[71]&m[411]&m[607]));
    m[224] = (((~m[34]&~m[342]&~m[538])|(m[34]&m[342]&~m[538]))&BiasedRNG[92])|(((m[34]&~m[342]&~m[538])|(~m[34]&m[342]&m[538]))&~BiasedRNG[92])|((~m[34]&~m[342]&m[538])|(m[34]&~m[342]&m[538])|(m[34]&m[342]&m[538]));
    m[225] = (((~m[34]&~m[356]&~m[552])|(m[34]&m[356]&~m[552]))&BiasedRNG[93])|(((m[34]&~m[356]&~m[552])|(~m[34]&m[356]&m[552]))&~BiasedRNG[93])|((~m[34]&~m[356]&m[552])|(m[34]&~m[356]&m[552])|(m[34]&m[356]&m[552]));
    m[226] = (((~m[74]&~m[370]&~m[566])|(m[74]&m[370]&~m[566]))&BiasedRNG[94])|(((m[74]&~m[370]&~m[566])|(~m[74]&m[370]&m[566]))&~BiasedRNG[94])|((~m[74]&~m[370]&m[566])|(m[74]&~m[370]&m[566])|(m[74]&m[370]&m[566]));
    m[227] = (((~m[74]&~m[384]&~m[580])|(m[74]&m[384]&~m[580]))&BiasedRNG[95])|(((m[74]&~m[384]&~m[580])|(~m[74]&m[384]&m[580]))&~BiasedRNG[95])|((~m[74]&~m[384]&m[580])|(m[74]&~m[384]&m[580])|(m[74]&m[384]&m[580]));
    m[228] = (((~m[74]&~m[398]&~m[594])|(m[74]&m[398]&~m[594]))&BiasedRNG[96])|(((m[74]&~m[398]&~m[594])|(~m[74]&m[398]&m[594]))&~BiasedRNG[96])|((~m[74]&~m[398]&m[594])|(m[74]&~m[398]&m[594])|(m[74]&m[398]&m[594]));
    m[229] = (((~m[74]&~m[412]&~m[608])|(m[74]&m[412]&~m[608]))&BiasedRNG[97])|(((m[74]&~m[412]&~m[608])|(~m[74]&m[412]&m[608]))&~BiasedRNG[97])|((~m[74]&~m[412]&m[608])|(m[74]&~m[412]&m[608])|(m[74]&m[412]&m[608]));
    m[238] = (((~m[35]&~m[343]&~m[539])|(m[35]&m[343]&~m[539]))&BiasedRNG[98])|(((m[35]&~m[343]&~m[539])|(~m[35]&m[343]&m[539]))&~BiasedRNG[98])|((~m[35]&~m[343]&m[539])|(m[35]&~m[343]&m[539])|(m[35]&m[343]&m[539]));
    m[239] = (((~m[35]&~m[357]&~m[553])|(m[35]&m[357]&~m[553]))&BiasedRNG[99])|(((m[35]&~m[357]&~m[553])|(~m[35]&m[357]&m[553]))&~BiasedRNG[99])|((~m[35]&~m[357]&m[553])|(m[35]&~m[357]&m[553])|(m[35]&m[357]&m[553]));
    m[240] = (((~m[77]&~m[371]&~m[567])|(m[77]&m[371]&~m[567]))&BiasedRNG[100])|(((m[77]&~m[371]&~m[567])|(~m[77]&m[371]&m[567]))&~BiasedRNG[100])|((~m[77]&~m[371]&m[567])|(m[77]&~m[371]&m[567])|(m[77]&m[371]&m[567]));
    m[241] = (((~m[77]&~m[385]&~m[581])|(m[77]&m[385]&~m[581]))&BiasedRNG[101])|(((m[77]&~m[385]&~m[581])|(~m[77]&m[385]&m[581]))&~BiasedRNG[101])|((~m[77]&~m[385]&m[581])|(m[77]&~m[385]&m[581])|(m[77]&m[385]&m[581]));
    m[242] = (((~m[77]&~m[399]&~m[595])|(m[77]&m[399]&~m[595]))&BiasedRNG[102])|(((m[77]&~m[399]&~m[595])|(~m[77]&m[399]&m[595]))&~BiasedRNG[102])|((~m[77]&~m[399]&m[595])|(m[77]&~m[399]&m[595])|(m[77]&m[399]&m[595]));
    m[243] = (((~m[77]&~m[413]&~m[609])|(m[77]&m[413]&~m[609]))&BiasedRNG[103])|(((m[77]&~m[413]&~m[609])|(~m[77]&m[413]&m[609]))&~BiasedRNG[103])|((~m[77]&~m[413]&m[609])|(m[77]&~m[413]&m[609])|(m[77]&m[413]&m[609]));
    m[252] = (((~m[36]&~m[344]&~m[540])|(m[36]&m[344]&~m[540]))&BiasedRNG[104])|(((m[36]&~m[344]&~m[540])|(~m[36]&m[344]&m[540]))&~BiasedRNG[104])|((~m[36]&~m[344]&m[540])|(m[36]&~m[344]&m[540])|(m[36]&m[344]&m[540]));
    m[253] = (((~m[36]&~m[358]&~m[554])|(m[36]&m[358]&~m[554]))&BiasedRNG[105])|(((m[36]&~m[358]&~m[554])|(~m[36]&m[358]&m[554]))&~BiasedRNG[105])|((~m[36]&~m[358]&m[554])|(m[36]&~m[358]&m[554])|(m[36]&m[358]&m[554]));
    m[254] = (((~m[80]&~m[372]&~m[568])|(m[80]&m[372]&~m[568]))&BiasedRNG[106])|(((m[80]&~m[372]&~m[568])|(~m[80]&m[372]&m[568]))&~BiasedRNG[106])|((~m[80]&~m[372]&m[568])|(m[80]&~m[372]&m[568])|(m[80]&m[372]&m[568]));
    m[255] = (((~m[80]&~m[386]&~m[582])|(m[80]&m[386]&~m[582]))&BiasedRNG[107])|(((m[80]&~m[386]&~m[582])|(~m[80]&m[386]&m[582]))&~BiasedRNG[107])|((~m[80]&~m[386]&m[582])|(m[80]&~m[386]&m[582])|(m[80]&m[386]&m[582]));
    m[256] = (((~m[80]&~m[400]&~m[596])|(m[80]&m[400]&~m[596]))&BiasedRNG[108])|(((m[80]&~m[400]&~m[596])|(~m[80]&m[400]&m[596]))&~BiasedRNG[108])|((~m[80]&~m[400]&m[596])|(m[80]&~m[400]&m[596])|(m[80]&m[400]&m[596]));
    m[257] = (((~m[80]&~m[414]&~m[610])|(m[80]&m[414]&~m[610]))&BiasedRNG[109])|(((m[80]&~m[414]&~m[610])|(~m[80]&m[414]&m[610]))&~BiasedRNG[109])|((~m[80]&~m[414]&m[610])|(m[80]&~m[414]&m[610])|(m[80]&m[414]&m[610]));
    m[266] = (((~m[37]&~m[345]&~m[541])|(m[37]&m[345]&~m[541]))&BiasedRNG[110])|(((m[37]&~m[345]&~m[541])|(~m[37]&m[345]&m[541]))&~BiasedRNG[110])|((~m[37]&~m[345]&m[541])|(m[37]&~m[345]&m[541])|(m[37]&m[345]&m[541]));
    m[267] = (((~m[37]&~m[359]&~m[555])|(m[37]&m[359]&~m[555]))&BiasedRNG[111])|(((m[37]&~m[359]&~m[555])|(~m[37]&m[359]&m[555]))&~BiasedRNG[111])|((~m[37]&~m[359]&m[555])|(m[37]&~m[359]&m[555])|(m[37]&m[359]&m[555]));
    m[268] = (((~m[83]&~m[373]&~m[569])|(m[83]&m[373]&~m[569]))&BiasedRNG[112])|(((m[83]&~m[373]&~m[569])|(~m[83]&m[373]&m[569]))&~BiasedRNG[112])|((~m[83]&~m[373]&m[569])|(m[83]&~m[373]&m[569])|(m[83]&m[373]&m[569]));
    m[269] = (((~m[83]&~m[387]&~m[583])|(m[83]&m[387]&~m[583]))&BiasedRNG[113])|(((m[83]&~m[387]&~m[583])|(~m[83]&m[387]&m[583]))&~BiasedRNG[113])|((~m[83]&~m[387]&m[583])|(m[83]&~m[387]&m[583])|(m[83]&m[387]&m[583]));
    m[270] = (((~m[83]&~m[401]&~m[597])|(m[83]&m[401]&~m[597]))&BiasedRNG[114])|(((m[83]&~m[401]&~m[597])|(~m[83]&m[401]&m[597]))&~BiasedRNG[114])|((~m[83]&~m[401]&m[597])|(m[83]&~m[401]&m[597])|(m[83]&m[401]&m[597]));
    m[271] = (((~m[83]&~m[415]&~m[611])|(m[83]&m[415]&~m[611]))&BiasedRNG[115])|(((m[83]&~m[415]&~m[611])|(~m[83]&m[415]&m[611]))&~BiasedRNG[115])|((~m[83]&~m[415]&m[611])|(m[83]&~m[415]&m[611])|(m[83]&m[415]&m[611]));
    m[280] = (((~m[38]&~m[346]&~m[542])|(m[38]&m[346]&~m[542]))&BiasedRNG[116])|(((m[38]&~m[346]&~m[542])|(~m[38]&m[346]&m[542]))&~BiasedRNG[116])|((~m[38]&~m[346]&m[542])|(m[38]&~m[346]&m[542])|(m[38]&m[346]&m[542]));
    m[281] = (((~m[38]&~m[360]&~m[556])|(m[38]&m[360]&~m[556]))&BiasedRNG[117])|(((m[38]&~m[360]&~m[556])|(~m[38]&m[360]&m[556]))&~BiasedRNG[117])|((~m[38]&~m[360]&m[556])|(m[38]&~m[360]&m[556])|(m[38]&m[360]&m[556]));
    m[282] = (((~m[86]&~m[374]&~m[570])|(m[86]&m[374]&~m[570]))&BiasedRNG[118])|(((m[86]&~m[374]&~m[570])|(~m[86]&m[374]&m[570]))&~BiasedRNG[118])|((~m[86]&~m[374]&m[570])|(m[86]&~m[374]&m[570])|(m[86]&m[374]&m[570]));
    m[283] = (((~m[86]&~m[388]&~m[584])|(m[86]&m[388]&~m[584]))&BiasedRNG[119])|(((m[86]&~m[388]&~m[584])|(~m[86]&m[388]&m[584]))&~BiasedRNG[119])|((~m[86]&~m[388]&m[584])|(m[86]&~m[388]&m[584])|(m[86]&m[388]&m[584]));
    m[284] = (((~m[86]&~m[402]&~m[598])|(m[86]&m[402]&~m[598]))&BiasedRNG[120])|(((m[86]&~m[402]&~m[598])|(~m[86]&m[402]&m[598]))&~BiasedRNG[120])|((~m[86]&~m[402]&m[598])|(m[86]&~m[402]&m[598])|(m[86]&m[402]&m[598]));
    m[285] = (((~m[86]&~m[416]&~m[612])|(m[86]&m[416]&~m[612]))&BiasedRNG[121])|(((m[86]&~m[416]&~m[612])|(~m[86]&m[416]&m[612]))&~BiasedRNG[121])|((~m[86]&~m[416]&m[612])|(m[86]&~m[416]&m[612])|(m[86]&m[416]&m[612]));
    m[294] = (((~m[39]&~m[347]&~m[543])|(m[39]&m[347]&~m[543]))&BiasedRNG[122])|(((m[39]&~m[347]&~m[543])|(~m[39]&m[347]&m[543]))&~BiasedRNG[122])|((~m[39]&~m[347]&m[543])|(m[39]&~m[347]&m[543])|(m[39]&m[347]&m[543]));
    m[295] = (((~m[39]&~m[361]&~m[557])|(m[39]&m[361]&~m[557]))&BiasedRNG[123])|(((m[39]&~m[361]&~m[557])|(~m[39]&m[361]&m[557]))&~BiasedRNG[123])|((~m[39]&~m[361]&m[557])|(m[39]&~m[361]&m[557])|(m[39]&m[361]&m[557]));
    m[296] = (((~m[89]&~m[375]&~m[571])|(m[89]&m[375]&~m[571]))&BiasedRNG[124])|(((m[89]&~m[375]&~m[571])|(~m[89]&m[375]&m[571]))&~BiasedRNG[124])|((~m[89]&~m[375]&m[571])|(m[89]&~m[375]&m[571])|(m[89]&m[375]&m[571]));
    m[297] = (((~m[89]&~m[389]&~m[585])|(m[89]&m[389]&~m[585]))&BiasedRNG[125])|(((m[89]&~m[389]&~m[585])|(~m[89]&m[389]&m[585]))&~BiasedRNG[125])|((~m[89]&~m[389]&m[585])|(m[89]&~m[389]&m[585])|(m[89]&m[389]&m[585]));
    m[298] = (((~m[89]&~m[403]&~m[599])|(m[89]&m[403]&~m[599]))&BiasedRNG[126])|(((m[89]&~m[403]&~m[599])|(~m[89]&m[403]&m[599]))&~BiasedRNG[126])|((~m[89]&~m[403]&m[599])|(m[89]&~m[403]&m[599])|(m[89]&m[403]&m[599]));
    m[299] = (((~m[89]&~m[417]&~m[613])|(m[89]&m[417]&~m[613]))&BiasedRNG[127])|(((m[89]&~m[417]&~m[613])|(~m[89]&m[417]&m[613]))&~BiasedRNG[127])|((~m[89]&~m[417]&m[613])|(m[89]&~m[417]&m[613])|(m[89]&m[417]&m[613]));
    m[308] = (((~m[40]&~m[348]&~m[544])|(m[40]&m[348]&~m[544]))&BiasedRNG[128])|(((m[40]&~m[348]&~m[544])|(~m[40]&m[348]&m[544]))&~BiasedRNG[128])|((~m[40]&~m[348]&m[544])|(m[40]&~m[348]&m[544])|(m[40]&m[348]&m[544]));
    m[309] = (((~m[40]&~m[362]&~m[558])|(m[40]&m[362]&~m[558]))&BiasedRNG[129])|(((m[40]&~m[362]&~m[558])|(~m[40]&m[362]&m[558]))&~BiasedRNG[129])|((~m[40]&~m[362]&m[558])|(m[40]&~m[362]&m[558])|(m[40]&m[362]&m[558]));
    m[310] = (((~m[92]&~m[376]&~m[572])|(m[92]&m[376]&~m[572]))&BiasedRNG[130])|(((m[92]&~m[376]&~m[572])|(~m[92]&m[376]&m[572]))&~BiasedRNG[130])|((~m[92]&~m[376]&m[572])|(m[92]&~m[376]&m[572])|(m[92]&m[376]&m[572]));
    m[311] = (((~m[92]&~m[390]&~m[586])|(m[92]&m[390]&~m[586]))&BiasedRNG[131])|(((m[92]&~m[390]&~m[586])|(~m[92]&m[390]&m[586]))&~BiasedRNG[131])|((~m[92]&~m[390]&m[586])|(m[92]&~m[390]&m[586])|(m[92]&m[390]&m[586]));
    m[312] = (((~m[92]&~m[404]&~m[600])|(m[92]&m[404]&~m[600]))&BiasedRNG[132])|(((m[92]&~m[404]&~m[600])|(~m[92]&m[404]&m[600]))&~BiasedRNG[132])|((~m[92]&~m[404]&m[600])|(m[92]&~m[404]&m[600])|(m[92]&m[404]&m[600]));
    m[313] = (((~m[92]&~m[418]&~m[614])|(m[92]&m[418]&~m[614]))&BiasedRNG[133])|(((m[92]&~m[418]&~m[614])|(~m[92]&m[418]&m[614]))&~BiasedRNG[133])|((~m[92]&~m[418]&m[614])|(m[92]&~m[418]&m[614])|(m[92]&m[418]&m[614]));
    m[322] = (((~m[41]&~m[349]&~m[545])|(m[41]&m[349]&~m[545]))&BiasedRNG[134])|(((m[41]&~m[349]&~m[545])|(~m[41]&m[349]&m[545]))&~BiasedRNG[134])|((~m[41]&~m[349]&m[545])|(m[41]&~m[349]&m[545])|(m[41]&m[349]&m[545]));
    m[323] = (((~m[41]&~m[363]&~m[559])|(m[41]&m[363]&~m[559]))&BiasedRNG[135])|(((m[41]&~m[363]&~m[559])|(~m[41]&m[363]&m[559]))&~BiasedRNG[135])|((~m[41]&~m[363]&m[559])|(m[41]&~m[363]&m[559])|(m[41]&m[363]&m[559]));
    m[324] = (((~m[95]&~m[377]&~m[573])|(m[95]&m[377]&~m[573]))&BiasedRNG[136])|(((m[95]&~m[377]&~m[573])|(~m[95]&m[377]&m[573]))&~BiasedRNG[136])|((~m[95]&~m[377]&m[573])|(m[95]&~m[377]&m[573])|(m[95]&m[377]&m[573]));
    m[325] = (((~m[95]&~m[391]&~m[587])|(m[95]&m[391]&~m[587]))&BiasedRNG[137])|(((m[95]&~m[391]&~m[587])|(~m[95]&m[391]&m[587]))&~BiasedRNG[137])|((~m[95]&~m[391]&m[587])|(m[95]&~m[391]&m[587])|(m[95]&m[391]&m[587]));
    m[326] = (((~m[95]&~m[405]&~m[601])|(m[95]&m[405]&~m[601]))&BiasedRNG[138])|(((m[95]&~m[405]&~m[601])|(~m[95]&m[405]&m[601]))&~BiasedRNG[138])|((~m[95]&~m[405]&m[601])|(m[95]&~m[405]&m[601])|(m[95]&m[405]&m[601]));
    m[327] = (((~m[95]&~m[419]&~m[615])|(m[95]&m[419]&~m[615]))&BiasedRNG[139])|(((m[95]&~m[419]&~m[615])|(~m[95]&m[419]&m[615]))&~BiasedRNG[139])|((~m[95]&~m[419]&m[615])|(m[95]&~m[419]&m[615])|(m[95]&m[419]&m[615]));
    m[420] = (((~m[48]&~m[146]&~m[616])|(m[48]&m[146]&~m[616]))&BiasedRNG[140])|(((m[48]&~m[146]&~m[616])|(~m[48]&m[146]&m[616]))&~BiasedRNG[140])|((~m[48]&~m[146]&m[616])|(m[48]&~m[146]&m[616])|(m[48]&m[146]&m[616]));
    m[421] = (((~m[48]&~m[160]&~m[617])|(m[48]&m[160]&~m[617]))&BiasedRNG[141])|(((m[48]&~m[160]&~m[617])|(~m[48]&m[160]&m[617]))&~BiasedRNG[141])|((~m[48]&~m[160]&m[617])|(m[48]&~m[160]&m[617])|(m[48]&m[160]&m[617]));
    m[422] = (((~m[116]&~m[174]&~m[618])|(m[116]&m[174]&~m[618]))&BiasedRNG[142])|(((m[116]&~m[174]&~m[618])|(~m[116]&m[174]&m[618]))&~BiasedRNG[142])|((~m[116]&~m[174]&m[618])|(m[116]&~m[174]&m[618])|(m[116]&m[174]&m[618]));
    m[423] = (((~m[116]&~m[188]&~m[619])|(m[116]&m[188]&~m[619]))&BiasedRNG[143])|(((m[116]&~m[188]&~m[619])|(~m[116]&m[188]&m[619]))&~BiasedRNG[143])|((~m[116]&~m[188]&m[619])|(m[116]&~m[188]&m[619])|(m[116]&m[188]&m[619]));
    m[424] = (((~m[116]&~m[202]&~m[620])|(m[116]&m[202]&~m[620]))&BiasedRNG[144])|(((m[116]&~m[202]&~m[620])|(~m[116]&m[202]&m[620]))&~BiasedRNG[144])|((~m[116]&~m[202]&m[620])|(m[116]&~m[202]&m[620])|(m[116]&m[202]&m[620]));
    m[425] = (((~m[116]&~m[216]&~m[621])|(m[116]&m[216]&~m[621]))&BiasedRNG[145])|(((m[116]&~m[216]&~m[621])|(~m[116]&m[216]&m[621]))&~BiasedRNG[145])|((~m[116]&~m[216]&m[621])|(m[116]&~m[216]&m[621])|(m[116]&m[216]&m[621]));
    m[434] = (((~m[49]&~m[147]&~m[630])|(m[49]&m[147]&~m[630]))&BiasedRNG[146])|(((m[49]&~m[147]&~m[630])|(~m[49]&m[147]&m[630]))&~BiasedRNG[146])|((~m[49]&~m[147]&m[630])|(m[49]&~m[147]&m[630])|(m[49]&m[147]&m[630]));
    m[435] = (((~m[49]&~m[161]&~m[631])|(m[49]&m[161]&~m[631]))&BiasedRNG[147])|(((m[49]&~m[161]&~m[631])|(~m[49]&m[161]&m[631]))&~BiasedRNG[147])|((~m[49]&~m[161]&m[631])|(m[49]&~m[161]&m[631])|(m[49]&m[161]&m[631]));
    m[436] = (((~m[119]&~m[175]&~m[632])|(m[119]&m[175]&~m[632]))&BiasedRNG[148])|(((m[119]&~m[175]&~m[632])|(~m[119]&m[175]&m[632]))&~BiasedRNG[148])|((~m[119]&~m[175]&m[632])|(m[119]&~m[175]&m[632])|(m[119]&m[175]&m[632]));
    m[437] = (((~m[119]&~m[189]&~m[633])|(m[119]&m[189]&~m[633]))&BiasedRNG[149])|(((m[119]&~m[189]&~m[633])|(~m[119]&m[189]&m[633]))&~BiasedRNG[149])|((~m[119]&~m[189]&m[633])|(m[119]&~m[189]&m[633])|(m[119]&m[189]&m[633]));
    m[438] = (((~m[119]&~m[203]&~m[634])|(m[119]&m[203]&~m[634]))&BiasedRNG[150])|(((m[119]&~m[203]&~m[634])|(~m[119]&m[203]&m[634]))&~BiasedRNG[150])|((~m[119]&~m[203]&m[634])|(m[119]&~m[203]&m[634])|(m[119]&m[203]&m[634]));
    m[439] = (((~m[119]&~m[217]&~m[635])|(m[119]&m[217]&~m[635]))&BiasedRNG[151])|(((m[119]&~m[217]&~m[635])|(~m[119]&m[217]&m[635]))&~BiasedRNG[151])|((~m[119]&~m[217]&m[635])|(m[119]&~m[217]&m[635])|(m[119]&m[217]&m[635]));
    m[448] = (((~m[50]&~m[148]&~m[644])|(m[50]&m[148]&~m[644]))&BiasedRNG[152])|(((m[50]&~m[148]&~m[644])|(~m[50]&m[148]&m[644]))&~BiasedRNG[152])|((~m[50]&~m[148]&m[644])|(m[50]&~m[148]&m[644])|(m[50]&m[148]&m[644]));
    m[449] = (((~m[50]&~m[162]&~m[645])|(m[50]&m[162]&~m[645]))&BiasedRNG[153])|(((m[50]&~m[162]&~m[645])|(~m[50]&m[162]&m[645]))&~BiasedRNG[153])|((~m[50]&~m[162]&m[645])|(m[50]&~m[162]&m[645])|(m[50]&m[162]&m[645]));
    m[450] = (((~m[122]&~m[176]&~m[646])|(m[122]&m[176]&~m[646]))&BiasedRNG[154])|(((m[122]&~m[176]&~m[646])|(~m[122]&m[176]&m[646]))&~BiasedRNG[154])|((~m[122]&~m[176]&m[646])|(m[122]&~m[176]&m[646])|(m[122]&m[176]&m[646]));
    m[451] = (((~m[122]&~m[190]&~m[647])|(m[122]&m[190]&~m[647]))&BiasedRNG[155])|(((m[122]&~m[190]&~m[647])|(~m[122]&m[190]&m[647]))&~BiasedRNG[155])|((~m[122]&~m[190]&m[647])|(m[122]&~m[190]&m[647])|(m[122]&m[190]&m[647]));
    m[452] = (((~m[122]&~m[204]&~m[648])|(m[122]&m[204]&~m[648]))&BiasedRNG[156])|(((m[122]&~m[204]&~m[648])|(~m[122]&m[204]&m[648]))&~BiasedRNG[156])|((~m[122]&~m[204]&m[648])|(m[122]&~m[204]&m[648])|(m[122]&m[204]&m[648]));
    m[453] = (((~m[122]&~m[218]&~m[649])|(m[122]&m[218]&~m[649]))&BiasedRNG[157])|(((m[122]&~m[218]&~m[649])|(~m[122]&m[218]&m[649]))&~BiasedRNG[157])|((~m[122]&~m[218]&m[649])|(m[122]&~m[218]&m[649])|(m[122]&m[218]&m[649]));
    m[462] = (((~m[51]&~m[149]&~m[658])|(m[51]&m[149]&~m[658]))&BiasedRNG[158])|(((m[51]&~m[149]&~m[658])|(~m[51]&m[149]&m[658]))&~BiasedRNG[158])|((~m[51]&~m[149]&m[658])|(m[51]&~m[149]&m[658])|(m[51]&m[149]&m[658]));
    m[463] = (((~m[51]&~m[163]&~m[659])|(m[51]&m[163]&~m[659]))&BiasedRNG[159])|(((m[51]&~m[163]&~m[659])|(~m[51]&m[163]&m[659]))&~BiasedRNG[159])|((~m[51]&~m[163]&m[659])|(m[51]&~m[163]&m[659])|(m[51]&m[163]&m[659]));
    m[464] = (((~m[125]&~m[177]&~m[660])|(m[125]&m[177]&~m[660]))&BiasedRNG[160])|(((m[125]&~m[177]&~m[660])|(~m[125]&m[177]&m[660]))&~BiasedRNG[160])|((~m[125]&~m[177]&m[660])|(m[125]&~m[177]&m[660])|(m[125]&m[177]&m[660]));
    m[465] = (((~m[125]&~m[191]&~m[661])|(m[125]&m[191]&~m[661]))&BiasedRNG[161])|(((m[125]&~m[191]&~m[661])|(~m[125]&m[191]&m[661]))&~BiasedRNG[161])|((~m[125]&~m[191]&m[661])|(m[125]&~m[191]&m[661])|(m[125]&m[191]&m[661]));
    m[466] = (((~m[125]&~m[205]&~m[662])|(m[125]&m[205]&~m[662]))&BiasedRNG[162])|(((m[125]&~m[205]&~m[662])|(~m[125]&m[205]&m[662]))&~BiasedRNG[162])|((~m[125]&~m[205]&m[662])|(m[125]&~m[205]&m[662])|(m[125]&m[205]&m[662]));
    m[467] = (((~m[125]&~m[219]&~m[663])|(m[125]&m[219]&~m[663]))&BiasedRNG[163])|(((m[125]&~m[219]&~m[663])|(~m[125]&m[219]&m[663]))&~BiasedRNG[163])|((~m[125]&~m[219]&m[663])|(m[125]&~m[219]&m[663])|(m[125]&m[219]&m[663]));
    m[476] = (((~m[52]&~m[150]&~m[672])|(m[52]&m[150]&~m[672]))&BiasedRNG[164])|(((m[52]&~m[150]&~m[672])|(~m[52]&m[150]&m[672]))&~BiasedRNG[164])|((~m[52]&~m[150]&m[672])|(m[52]&~m[150]&m[672])|(m[52]&m[150]&m[672]));
    m[477] = (((~m[52]&~m[164]&~m[673])|(m[52]&m[164]&~m[673]))&BiasedRNG[165])|(((m[52]&~m[164]&~m[673])|(~m[52]&m[164]&m[673]))&~BiasedRNG[165])|((~m[52]&~m[164]&m[673])|(m[52]&~m[164]&m[673])|(m[52]&m[164]&m[673]));
    m[478] = (((~m[128]&~m[178]&~m[674])|(m[128]&m[178]&~m[674]))&BiasedRNG[166])|(((m[128]&~m[178]&~m[674])|(~m[128]&m[178]&m[674]))&~BiasedRNG[166])|((~m[128]&~m[178]&m[674])|(m[128]&~m[178]&m[674])|(m[128]&m[178]&m[674]));
    m[479] = (((~m[128]&~m[192]&~m[675])|(m[128]&m[192]&~m[675]))&BiasedRNG[167])|(((m[128]&~m[192]&~m[675])|(~m[128]&m[192]&m[675]))&~BiasedRNG[167])|((~m[128]&~m[192]&m[675])|(m[128]&~m[192]&m[675])|(m[128]&m[192]&m[675]));
    m[480] = (((~m[128]&~m[206]&~m[676])|(m[128]&m[206]&~m[676]))&BiasedRNG[168])|(((m[128]&~m[206]&~m[676])|(~m[128]&m[206]&m[676]))&~BiasedRNG[168])|((~m[128]&~m[206]&m[676])|(m[128]&~m[206]&m[676])|(m[128]&m[206]&m[676]));
    m[481] = (((~m[128]&~m[220]&~m[677])|(m[128]&m[220]&~m[677]))&BiasedRNG[169])|(((m[128]&~m[220]&~m[677])|(~m[128]&m[220]&m[677]))&~BiasedRNG[169])|((~m[128]&~m[220]&m[677])|(m[128]&~m[220]&m[677])|(m[128]&m[220]&m[677]));
    m[490] = (((~m[53]&~m[151]&~m[686])|(m[53]&m[151]&~m[686]))&BiasedRNG[170])|(((m[53]&~m[151]&~m[686])|(~m[53]&m[151]&m[686]))&~BiasedRNG[170])|((~m[53]&~m[151]&m[686])|(m[53]&~m[151]&m[686])|(m[53]&m[151]&m[686]));
    m[491] = (((~m[53]&~m[165]&~m[687])|(m[53]&m[165]&~m[687]))&BiasedRNG[171])|(((m[53]&~m[165]&~m[687])|(~m[53]&m[165]&m[687]))&~BiasedRNG[171])|((~m[53]&~m[165]&m[687])|(m[53]&~m[165]&m[687])|(m[53]&m[165]&m[687]));
    m[492] = (((~m[131]&~m[179]&~m[688])|(m[131]&m[179]&~m[688]))&BiasedRNG[172])|(((m[131]&~m[179]&~m[688])|(~m[131]&m[179]&m[688]))&~BiasedRNG[172])|((~m[131]&~m[179]&m[688])|(m[131]&~m[179]&m[688])|(m[131]&m[179]&m[688]));
    m[493] = (((~m[131]&~m[193]&~m[689])|(m[131]&m[193]&~m[689]))&BiasedRNG[173])|(((m[131]&~m[193]&~m[689])|(~m[131]&m[193]&m[689]))&~BiasedRNG[173])|((~m[131]&~m[193]&m[689])|(m[131]&~m[193]&m[689])|(m[131]&m[193]&m[689]));
    m[494] = (((~m[131]&~m[207]&~m[690])|(m[131]&m[207]&~m[690]))&BiasedRNG[174])|(((m[131]&~m[207]&~m[690])|(~m[131]&m[207]&m[690]))&~BiasedRNG[174])|((~m[131]&~m[207]&m[690])|(m[131]&~m[207]&m[690])|(m[131]&m[207]&m[690]));
    m[495] = (((~m[131]&~m[221]&~m[691])|(m[131]&m[221]&~m[691]))&BiasedRNG[175])|(((m[131]&~m[221]&~m[691])|(~m[131]&m[221]&m[691]))&~BiasedRNG[175])|((~m[131]&~m[221]&m[691])|(m[131]&~m[221]&m[691])|(m[131]&m[221]&m[691]));
    m[504] = (((~m[54]&~m[152]&~m[700])|(m[54]&m[152]&~m[700]))&BiasedRNG[176])|(((m[54]&~m[152]&~m[700])|(~m[54]&m[152]&m[700]))&~BiasedRNG[176])|((~m[54]&~m[152]&m[700])|(m[54]&~m[152]&m[700])|(m[54]&m[152]&m[700]));
    m[505] = (((~m[54]&~m[166]&~m[701])|(m[54]&m[166]&~m[701]))&BiasedRNG[177])|(((m[54]&~m[166]&~m[701])|(~m[54]&m[166]&m[701]))&~BiasedRNG[177])|((~m[54]&~m[166]&m[701])|(m[54]&~m[166]&m[701])|(m[54]&m[166]&m[701]));
    m[506] = (((~m[134]&~m[180]&~m[702])|(m[134]&m[180]&~m[702]))&BiasedRNG[178])|(((m[134]&~m[180]&~m[702])|(~m[134]&m[180]&m[702]))&~BiasedRNG[178])|((~m[134]&~m[180]&m[702])|(m[134]&~m[180]&m[702])|(m[134]&m[180]&m[702]));
    m[507] = (((~m[134]&~m[194]&~m[703])|(m[134]&m[194]&~m[703]))&BiasedRNG[179])|(((m[134]&~m[194]&~m[703])|(~m[134]&m[194]&m[703]))&~BiasedRNG[179])|((~m[134]&~m[194]&m[703])|(m[134]&~m[194]&m[703])|(m[134]&m[194]&m[703]));
    m[508] = (((~m[134]&~m[208]&~m[704])|(m[134]&m[208]&~m[704]))&BiasedRNG[180])|(((m[134]&~m[208]&~m[704])|(~m[134]&m[208]&m[704]))&~BiasedRNG[180])|((~m[134]&~m[208]&m[704])|(m[134]&~m[208]&m[704])|(m[134]&m[208]&m[704]));
    m[509] = (((~m[134]&~m[222]&~m[705])|(m[134]&m[222]&~m[705]))&BiasedRNG[181])|(((m[134]&~m[222]&~m[705])|(~m[134]&m[222]&m[705]))&~BiasedRNG[181])|((~m[134]&~m[222]&m[705])|(m[134]&~m[222]&m[705])|(m[134]&m[222]&m[705]));
    m[518] = (((~m[55]&~m[153]&~m[714])|(m[55]&m[153]&~m[714]))&BiasedRNG[182])|(((m[55]&~m[153]&~m[714])|(~m[55]&m[153]&m[714]))&~BiasedRNG[182])|((~m[55]&~m[153]&m[714])|(m[55]&~m[153]&m[714])|(m[55]&m[153]&m[714]));
    m[519] = (((~m[55]&~m[167]&~m[715])|(m[55]&m[167]&~m[715]))&BiasedRNG[183])|(((m[55]&~m[167]&~m[715])|(~m[55]&m[167]&m[715]))&~BiasedRNG[183])|((~m[55]&~m[167]&m[715])|(m[55]&~m[167]&m[715])|(m[55]&m[167]&m[715]));
    m[520] = (((~m[137]&~m[181]&~m[716])|(m[137]&m[181]&~m[716]))&BiasedRNG[184])|(((m[137]&~m[181]&~m[716])|(~m[137]&m[181]&m[716]))&~BiasedRNG[184])|((~m[137]&~m[181]&m[716])|(m[137]&~m[181]&m[716])|(m[137]&m[181]&m[716]));
    m[521] = (((~m[137]&~m[195]&~m[717])|(m[137]&m[195]&~m[717]))&BiasedRNG[185])|(((m[137]&~m[195]&~m[717])|(~m[137]&m[195]&m[717]))&~BiasedRNG[185])|((~m[137]&~m[195]&m[717])|(m[137]&~m[195]&m[717])|(m[137]&m[195]&m[717]));
    m[522] = (((~m[137]&~m[209]&~m[718])|(m[137]&m[209]&~m[718]))&BiasedRNG[186])|(((m[137]&~m[209]&~m[718])|(~m[137]&m[209]&m[718]))&~BiasedRNG[186])|((~m[137]&~m[209]&m[718])|(m[137]&~m[209]&m[718])|(m[137]&m[209]&m[718]));
    m[523] = (((~m[137]&~m[223]&~m[719])|(m[137]&m[223]&~m[719]))&BiasedRNG[187])|(((m[137]&~m[223]&~m[719])|(~m[137]&m[223]&m[719]))&~BiasedRNG[187])|((~m[137]&~m[223]&m[719])|(m[137]&~m[223]&m[719])|(m[137]&m[223]&m[719]));
    m[622] = (((m[230]&~m[426]&m[1084])|(~m[230]&m[426]&m[1084]))&BiasedRNG[188])|(((m[230]&m[426]&~m[1084]))&~BiasedRNG[188])|((m[230]&m[426]&m[1084]));
    m[623] = (((m[244]&~m[427]&m[1144])|(~m[244]&m[427]&m[1144]))&BiasedRNG[189])|(((m[244]&m[427]&~m[1144]))&~BiasedRNG[189])|((m[244]&m[427]&m[1144]));
    m[624] = (((m[258]&~m[428]&m[1209])|(~m[258]&m[428]&m[1209]))&BiasedRNG[190])|(((m[258]&m[428]&~m[1209]))&~BiasedRNG[190])|((m[258]&m[428]&m[1209]));
    m[625] = (((m[272]&~m[429]&m[1269])|(~m[272]&m[429]&m[1269]))&BiasedRNG[191])|(((m[272]&m[429]&~m[1269]))&~BiasedRNG[191])|((m[272]&m[429]&m[1269]));
    m[626] = (((m[286]&~m[430]&m[1324])|(~m[286]&m[430]&m[1324]))&BiasedRNG[192])|(((m[286]&m[430]&~m[1324]))&~BiasedRNG[192])|((m[286]&m[430]&m[1324]));
    m[627] = (((m[300]&~m[431]&m[1374])|(~m[300]&m[431]&m[1374]))&BiasedRNG[193])|(((m[300]&m[431]&~m[1374]))&~BiasedRNG[193])|((m[300]&m[431]&m[1374]));
    m[628] = (((m[314]&~m[432]&m[1419])|(~m[314]&m[432]&m[1419]))&BiasedRNG[194])|(((m[314]&m[432]&~m[1419]))&~BiasedRNG[194])|((m[314]&m[432]&m[1419]));
    m[629] = (((m[328]&~m[433]&m[1459])|(~m[328]&m[433]&m[1459]))&BiasedRNG[195])|(((m[328]&m[433]&~m[1459]))&~BiasedRNG[195])|((m[328]&m[433]&m[1459]));
    m[636] = (((m[231]&~m[440]&m[1149])|(~m[231]&m[440]&m[1149]))&BiasedRNG[196])|(((m[231]&m[440]&~m[1149]))&~BiasedRNG[196])|((m[231]&m[440]&m[1149]));
    m[637] = (((m[245]&~m[441]&m[1214])|(~m[245]&m[441]&m[1214]))&BiasedRNG[197])|(((m[245]&m[441]&~m[1214]))&~BiasedRNG[197])|((m[245]&m[441]&m[1214]));
    m[638] = (((m[259]&~m[442]&m[1274])|(~m[259]&m[442]&m[1274]))&BiasedRNG[198])|(((m[259]&m[442]&~m[1274]))&~BiasedRNG[198])|((m[259]&m[442]&m[1274]));
    m[639] = (((m[273]&~m[443]&m[1329])|(~m[273]&m[443]&m[1329]))&BiasedRNG[199])|(((m[273]&m[443]&~m[1329]))&~BiasedRNG[199])|((m[273]&m[443]&m[1329]));
    m[640] = (((m[287]&~m[444]&m[1379])|(~m[287]&m[444]&m[1379]))&BiasedRNG[200])|(((m[287]&m[444]&~m[1379]))&~BiasedRNG[200])|((m[287]&m[444]&m[1379]));
    m[641] = (((m[301]&~m[445]&m[1424])|(~m[301]&m[445]&m[1424]))&BiasedRNG[201])|(((m[301]&m[445]&~m[1424]))&~BiasedRNG[201])|((m[301]&m[445]&m[1424]));
    m[642] = (((m[315]&~m[446]&m[1464])|(~m[315]&m[446]&m[1464]))&BiasedRNG[202])|(((m[315]&m[446]&~m[1464]))&~BiasedRNG[202])|((m[315]&m[446]&m[1464]));
    m[643] = (((m[329]&~m[447]&m[1499])|(~m[329]&m[447]&m[1499]))&BiasedRNG[203])|(((m[329]&m[447]&~m[1499]))&~BiasedRNG[203])|((m[329]&m[447]&m[1499]));
    m[650] = (((m[232]&~m[454]&m[1219])|(~m[232]&m[454]&m[1219]))&BiasedRNG[204])|(((m[232]&m[454]&~m[1219]))&~BiasedRNG[204])|((m[232]&m[454]&m[1219]));
    m[651] = (((m[246]&~m[455]&m[1279])|(~m[246]&m[455]&m[1279]))&BiasedRNG[205])|(((m[246]&m[455]&~m[1279]))&~BiasedRNG[205])|((m[246]&m[455]&m[1279]));
    m[652] = (((m[260]&~m[456]&m[1334])|(~m[260]&m[456]&m[1334]))&BiasedRNG[206])|(((m[260]&m[456]&~m[1334]))&~BiasedRNG[206])|((m[260]&m[456]&m[1334]));
    m[653] = (((m[274]&~m[457]&m[1384])|(~m[274]&m[457]&m[1384]))&BiasedRNG[207])|(((m[274]&m[457]&~m[1384]))&~BiasedRNG[207])|((m[274]&m[457]&m[1384]));
    m[654] = (((m[288]&~m[458]&m[1429])|(~m[288]&m[458]&m[1429]))&BiasedRNG[208])|(((m[288]&m[458]&~m[1429]))&~BiasedRNG[208])|((m[288]&m[458]&m[1429]));
    m[655] = (((m[302]&~m[459]&m[1469])|(~m[302]&m[459]&m[1469]))&BiasedRNG[209])|(((m[302]&m[459]&~m[1469]))&~BiasedRNG[209])|((m[302]&m[459]&m[1469]));
    m[656] = (((m[316]&~m[460]&m[1504])|(~m[316]&m[460]&m[1504]))&BiasedRNG[210])|(((m[316]&m[460]&~m[1504]))&~BiasedRNG[210])|((m[316]&m[460]&m[1504]));
    m[657] = (((m[330]&~m[461]&m[1534])|(~m[330]&m[461]&m[1534]))&BiasedRNG[211])|(((m[330]&m[461]&~m[1534]))&~BiasedRNG[211])|((m[330]&m[461]&m[1534]));
    m[664] = (((m[233]&~m[468]&m[1284])|(~m[233]&m[468]&m[1284]))&BiasedRNG[212])|(((m[233]&m[468]&~m[1284]))&~BiasedRNG[212])|((m[233]&m[468]&m[1284]));
    m[665] = (((m[247]&~m[469]&m[1339])|(~m[247]&m[469]&m[1339]))&BiasedRNG[213])|(((m[247]&m[469]&~m[1339]))&~BiasedRNG[213])|((m[247]&m[469]&m[1339]));
    m[666] = (((m[261]&~m[470]&m[1389])|(~m[261]&m[470]&m[1389]))&BiasedRNG[214])|(((m[261]&m[470]&~m[1389]))&~BiasedRNG[214])|((m[261]&m[470]&m[1389]));
    m[667] = (((m[275]&~m[471]&m[1434])|(~m[275]&m[471]&m[1434]))&BiasedRNG[215])|(((m[275]&m[471]&~m[1434]))&~BiasedRNG[215])|((m[275]&m[471]&m[1434]));
    m[668] = (((m[289]&~m[472]&m[1474])|(~m[289]&m[472]&m[1474]))&BiasedRNG[216])|(((m[289]&m[472]&~m[1474]))&~BiasedRNG[216])|((m[289]&m[472]&m[1474]));
    m[669] = (((m[303]&~m[473]&m[1509])|(~m[303]&m[473]&m[1509]))&BiasedRNG[217])|(((m[303]&m[473]&~m[1509]))&~BiasedRNG[217])|((m[303]&m[473]&m[1509]));
    m[670] = (((m[317]&~m[474]&m[1539])|(~m[317]&m[474]&m[1539]))&BiasedRNG[218])|(((m[317]&m[474]&~m[1539]))&~BiasedRNG[218])|((m[317]&m[474]&m[1539]));
    m[671] = (((m[331]&~m[475]&m[1564])|(~m[331]&m[475]&m[1564]))&BiasedRNG[219])|(((m[331]&m[475]&~m[1564]))&~BiasedRNG[219])|((m[331]&m[475]&m[1564]));
    m[678] = (((m[234]&~m[482]&m[1344])|(~m[234]&m[482]&m[1344]))&BiasedRNG[220])|(((m[234]&m[482]&~m[1344]))&~BiasedRNG[220])|((m[234]&m[482]&m[1344]));
    m[679] = (((m[248]&~m[483]&m[1394])|(~m[248]&m[483]&m[1394]))&BiasedRNG[221])|(((m[248]&m[483]&~m[1394]))&~BiasedRNG[221])|((m[248]&m[483]&m[1394]));
    m[680] = (((m[262]&~m[484]&m[1439])|(~m[262]&m[484]&m[1439]))&BiasedRNG[222])|(((m[262]&m[484]&~m[1439]))&~BiasedRNG[222])|((m[262]&m[484]&m[1439]));
    m[681] = (((m[276]&~m[485]&m[1479])|(~m[276]&m[485]&m[1479]))&BiasedRNG[223])|(((m[276]&m[485]&~m[1479]))&~BiasedRNG[223])|((m[276]&m[485]&m[1479]));
    m[682] = (((m[290]&~m[486]&m[1514])|(~m[290]&m[486]&m[1514]))&BiasedRNG[224])|(((m[290]&m[486]&~m[1514]))&~BiasedRNG[224])|((m[290]&m[486]&m[1514]));
    m[683] = (((m[304]&~m[487]&m[1544])|(~m[304]&m[487]&m[1544]))&BiasedRNG[225])|(((m[304]&m[487]&~m[1544]))&~BiasedRNG[225])|((m[304]&m[487]&m[1544]));
    m[684] = (((m[318]&~m[488]&m[1569])|(~m[318]&m[488]&m[1569]))&BiasedRNG[226])|(((m[318]&m[488]&~m[1569]))&~BiasedRNG[226])|((m[318]&m[488]&m[1569]));
    m[685] = (((m[332]&~m[489]&m[1589])|(~m[332]&m[489]&m[1589]))&BiasedRNG[227])|(((m[332]&m[489]&~m[1589]))&~BiasedRNG[227])|((m[332]&m[489]&m[1589]));
    m[692] = (((m[235]&~m[496]&m[1399])|(~m[235]&m[496]&m[1399]))&BiasedRNG[228])|(((m[235]&m[496]&~m[1399]))&~BiasedRNG[228])|((m[235]&m[496]&m[1399]));
    m[693] = (((m[249]&~m[497]&m[1444])|(~m[249]&m[497]&m[1444]))&BiasedRNG[229])|(((m[249]&m[497]&~m[1444]))&~BiasedRNG[229])|((m[249]&m[497]&m[1444]));
    m[694] = (((m[263]&~m[498]&m[1484])|(~m[263]&m[498]&m[1484]))&BiasedRNG[230])|(((m[263]&m[498]&~m[1484]))&~BiasedRNG[230])|((m[263]&m[498]&m[1484]));
    m[695] = (((m[277]&~m[499]&m[1519])|(~m[277]&m[499]&m[1519]))&BiasedRNG[231])|(((m[277]&m[499]&~m[1519]))&~BiasedRNG[231])|((m[277]&m[499]&m[1519]));
    m[696] = (((m[291]&~m[500]&m[1549])|(~m[291]&m[500]&m[1549]))&BiasedRNG[232])|(((m[291]&m[500]&~m[1549]))&~BiasedRNG[232])|((m[291]&m[500]&m[1549]));
    m[697] = (((m[305]&~m[501]&m[1574])|(~m[305]&m[501]&m[1574]))&BiasedRNG[233])|(((m[305]&m[501]&~m[1574]))&~BiasedRNG[233])|((m[305]&m[501]&m[1574]));
    m[698] = (((m[319]&~m[502]&m[1594])|(~m[319]&m[502]&m[1594]))&BiasedRNG[234])|(((m[319]&m[502]&~m[1594]))&~BiasedRNG[234])|((m[319]&m[502]&m[1594]));
    m[699] = (((m[333]&~m[503]&m[1609])|(~m[333]&m[503]&m[1609]))&BiasedRNG[235])|(((m[333]&m[503]&~m[1609]))&~BiasedRNG[235])|((m[333]&m[503]&m[1609]));
    m[706] = (((m[236]&~m[510]&m[1449])|(~m[236]&m[510]&m[1449]))&BiasedRNG[236])|(((m[236]&m[510]&~m[1449]))&~BiasedRNG[236])|((m[236]&m[510]&m[1449]));
    m[707] = (((m[250]&~m[511]&m[1489])|(~m[250]&m[511]&m[1489]))&BiasedRNG[237])|(((m[250]&m[511]&~m[1489]))&~BiasedRNG[237])|((m[250]&m[511]&m[1489]));
    m[708] = (((m[264]&~m[512]&m[1524])|(~m[264]&m[512]&m[1524]))&BiasedRNG[238])|(((m[264]&m[512]&~m[1524]))&~BiasedRNG[238])|((m[264]&m[512]&m[1524]));
    m[709] = (((m[278]&~m[513]&m[1554])|(~m[278]&m[513]&m[1554]))&BiasedRNG[239])|(((m[278]&m[513]&~m[1554]))&~BiasedRNG[239])|((m[278]&m[513]&m[1554]));
    m[710] = (((m[292]&~m[514]&m[1579])|(~m[292]&m[514]&m[1579]))&BiasedRNG[240])|(((m[292]&m[514]&~m[1579]))&~BiasedRNG[240])|((m[292]&m[514]&m[1579]));
    m[711] = (((m[306]&~m[515]&m[1599])|(~m[306]&m[515]&m[1599]))&BiasedRNG[241])|(((m[306]&m[515]&~m[1599]))&~BiasedRNG[241])|((m[306]&m[515]&m[1599]));
    m[712] = (((m[320]&~m[516]&m[1614])|(~m[320]&m[516]&m[1614]))&BiasedRNG[242])|(((m[320]&m[516]&~m[1614]))&~BiasedRNG[242])|((m[320]&m[516]&m[1614]));
    m[713] = (((m[334]&~m[517]&m[1624])|(~m[334]&m[517]&m[1624]))&BiasedRNG[243])|(((m[334]&m[517]&~m[1624]))&~BiasedRNG[243])|((m[334]&m[517]&m[1624]));
    m[720] = (((m[237]&~m[524]&m[1494])|(~m[237]&m[524]&m[1494]))&BiasedRNG[244])|(((m[237]&m[524]&~m[1494]))&~BiasedRNG[244])|((m[237]&m[524]&m[1494]));
    m[721] = (((m[251]&~m[525]&m[1529])|(~m[251]&m[525]&m[1529]))&BiasedRNG[245])|(((m[251]&m[525]&~m[1529]))&~BiasedRNG[245])|((m[251]&m[525]&m[1529]));
    m[722] = (((m[265]&~m[526]&m[1559])|(~m[265]&m[526]&m[1559]))&BiasedRNG[246])|(((m[265]&m[526]&~m[1559]))&~BiasedRNG[246])|((m[265]&m[526]&m[1559]));
    m[723] = (((m[279]&~m[527]&m[1584])|(~m[279]&m[527]&m[1584]))&BiasedRNG[247])|(((m[279]&m[527]&~m[1584]))&~BiasedRNG[247])|((m[279]&m[527]&m[1584]));
    m[724] = (((m[293]&~m[528]&m[1604])|(~m[293]&m[528]&m[1604]))&BiasedRNG[248])|(((m[293]&m[528]&~m[1604]))&~BiasedRNG[248])|((m[293]&m[528]&m[1604]));
    m[725] = (((m[307]&~m[529]&m[1619])|(~m[307]&m[529]&m[1619]))&BiasedRNG[249])|(((m[307]&m[529]&~m[1619]))&~BiasedRNG[249])|((m[307]&m[529]&m[1619]));
    m[726] = (((m[321]&~m[530]&m[1629])|(~m[321]&m[530]&m[1629]))&BiasedRNG[250])|(((m[321]&m[530]&~m[1629]))&~BiasedRNG[250])|((m[321]&m[530]&m[1629]));
    m[727] = (((m[335]&~m[531]&m[1634])|(~m[335]&m[531]&m[1634]))&BiasedRNG[251])|(((m[335]&m[531]&~m[1634]))&~BiasedRNG[251])|((m[335]&m[531]&m[1634]));
    m[728] = (((m[533]&~m[729]&~m[730]&~m[731]&~m[732])|(~m[533]&~m[729]&~m[730]&m[731]&~m[732])|(m[533]&m[729]&~m[730]&m[731]&~m[732])|(m[533]&~m[729]&m[730]&m[731]&~m[732])|(~m[533]&m[729]&~m[730]&~m[731]&m[732])|(~m[533]&~m[729]&m[730]&~m[731]&m[732])|(m[533]&m[729]&m[730]&~m[731]&m[732])|(~m[533]&m[729]&m[730]&m[731]&m[732]))&UnbiasedRNG[28])|((m[533]&~m[729]&~m[730]&m[731]&~m[732])|(~m[533]&~m[729]&~m[730]&~m[731]&m[732])|(m[533]&~m[729]&~m[730]&~m[731]&m[732])|(m[533]&m[729]&~m[730]&~m[731]&m[732])|(m[533]&~m[729]&m[730]&~m[731]&m[732])|(~m[533]&~m[729]&~m[730]&m[731]&m[732])|(m[533]&~m[729]&~m[730]&m[731]&m[732])|(~m[533]&m[729]&~m[730]&m[731]&m[732])|(m[533]&m[729]&~m[730]&m[731]&m[732])|(~m[533]&~m[729]&m[730]&m[731]&m[732])|(m[533]&~m[729]&m[730]&m[731]&m[732])|(m[533]&m[729]&m[730]&m[731]&m[732]));
    m[733] = (((m[534]&~m[734]&~m[735]&~m[736]&~m[737])|(~m[534]&~m[734]&~m[735]&m[736]&~m[737])|(m[534]&m[734]&~m[735]&m[736]&~m[737])|(m[534]&~m[734]&m[735]&m[736]&~m[737])|(~m[534]&m[734]&~m[735]&~m[736]&m[737])|(~m[534]&~m[734]&m[735]&~m[736]&m[737])|(m[534]&m[734]&m[735]&~m[736]&m[737])|(~m[534]&m[734]&m[735]&m[736]&m[737]))&UnbiasedRNG[29])|((m[534]&~m[734]&~m[735]&m[736]&~m[737])|(~m[534]&~m[734]&~m[735]&~m[736]&m[737])|(m[534]&~m[734]&~m[735]&~m[736]&m[737])|(m[534]&m[734]&~m[735]&~m[736]&m[737])|(m[534]&~m[734]&m[735]&~m[736]&m[737])|(~m[534]&~m[734]&~m[735]&m[736]&m[737])|(m[534]&~m[734]&~m[735]&m[736]&m[737])|(~m[534]&m[734]&~m[735]&m[736]&m[737])|(m[534]&m[734]&~m[735]&m[736]&m[737])|(~m[534]&~m[734]&m[735]&m[736]&m[737])|(m[534]&~m[734]&m[735]&m[736]&m[737])|(m[534]&m[734]&m[735]&m[736]&m[737]));
    m[738] = (((m[736]&~m[739]&~m[740]&~m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&m[741]&~m[742])|(m[736]&m[739]&~m[740]&m[741]&~m[742])|(m[736]&~m[739]&m[740]&m[741]&~m[742])|(~m[736]&m[739]&~m[740]&~m[741]&m[742])|(~m[736]&~m[739]&m[740]&~m[741]&m[742])|(m[736]&m[739]&m[740]&~m[741]&m[742])|(~m[736]&m[739]&m[740]&m[741]&m[742]))&UnbiasedRNG[30])|((m[736]&~m[739]&~m[740]&m[741]&~m[742])|(~m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&~m[740]&~m[741]&m[742])|(m[736]&m[739]&~m[740]&~m[741]&m[742])|(m[736]&~m[739]&m[740]&~m[741]&m[742])|(~m[736]&~m[739]&~m[740]&m[741]&m[742])|(m[736]&~m[739]&~m[740]&m[741]&m[742])|(~m[736]&m[739]&~m[740]&m[741]&m[742])|(m[736]&m[739]&~m[740]&m[741]&m[742])|(~m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&~m[739]&m[740]&m[741]&m[742])|(m[736]&m[739]&m[740]&m[741]&m[742]));
    m[743] = (((m[535]&~m[744]&~m[745]&~m[746]&~m[747])|(~m[535]&~m[744]&~m[745]&m[746]&~m[747])|(m[535]&m[744]&~m[745]&m[746]&~m[747])|(m[535]&~m[744]&m[745]&m[746]&~m[747])|(~m[535]&m[744]&~m[745]&~m[746]&m[747])|(~m[535]&~m[744]&m[745]&~m[746]&m[747])|(m[535]&m[744]&m[745]&~m[746]&m[747])|(~m[535]&m[744]&m[745]&m[746]&m[747]))&UnbiasedRNG[31])|((m[535]&~m[744]&~m[745]&m[746]&~m[747])|(~m[535]&~m[744]&~m[745]&~m[746]&m[747])|(m[535]&~m[744]&~m[745]&~m[746]&m[747])|(m[535]&m[744]&~m[745]&~m[746]&m[747])|(m[535]&~m[744]&m[745]&~m[746]&m[747])|(~m[535]&~m[744]&~m[745]&m[746]&m[747])|(m[535]&~m[744]&~m[745]&m[746]&m[747])|(~m[535]&m[744]&~m[745]&m[746]&m[747])|(m[535]&m[744]&~m[745]&m[746]&m[747])|(~m[535]&~m[744]&m[745]&m[746]&m[747])|(m[535]&~m[744]&m[745]&m[746]&m[747])|(m[535]&m[744]&m[745]&m[746]&m[747]));
    m[748] = (((m[746]&~m[749]&~m[750]&~m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&m[751]&~m[752])|(m[746]&m[749]&~m[750]&m[751]&~m[752])|(m[746]&~m[749]&m[750]&m[751]&~m[752])|(~m[746]&m[749]&~m[750]&~m[751]&m[752])|(~m[746]&~m[749]&m[750]&~m[751]&m[752])|(m[746]&m[749]&m[750]&~m[751]&m[752])|(~m[746]&m[749]&m[750]&m[751]&m[752]))&UnbiasedRNG[32])|((m[746]&~m[749]&~m[750]&m[751]&~m[752])|(~m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&~m[750]&~m[751]&m[752])|(m[746]&m[749]&~m[750]&~m[751]&m[752])|(m[746]&~m[749]&m[750]&~m[751]&m[752])|(~m[746]&~m[749]&~m[750]&m[751]&m[752])|(m[746]&~m[749]&~m[750]&m[751]&m[752])|(~m[746]&m[749]&~m[750]&m[751]&m[752])|(m[746]&m[749]&~m[750]&m[751]&m[752])|(~m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&~m[749]&m[750]&m[751]&m[752])|(m[746]&m[749]&m[750]&m[751]&m[752]));
    m[753] = (((m[751]&~m[754]&~m[755]&~m[756]&~m[757])|(~m[751]&~m[754]&~m[755]&m[756]&~m[757])|(m[751]&m[754]&~m[755]&m[756]&~m[757])|(m[751]&~m[754]&m[755]&m[756]&~m[757])|(~m[751]&m[754]&~m[755]&~m[756]&m[757])|(~m[751]&~m[754]&m[755]&~m[756]&m[757])|(m[751]&m[754]&m[755]&~m[756]&m[757])|(~m[751]&m[754]&m[755]&m[756]&m[757]))&UnbiasedRNG[33])|((m[751]&~m[754]&~m[755]&m[756]&~m[757])|(~m[751]&~m[754]&~m[755]&~m[756]&m[757])|(m[751]&~m[754]&~m[755]&~m[756]&m[757])|(m[751]&m[754]&~m[755]&~m[756]&m[757])|(m[751]&~m[754]&m[755]&~m[756]&m[757])|(~m[751]&~m[754]&~m[755]&m[756]&m[757])|(m[751]&~m[754]&~m[755]&m[756]&m[757])|(~m[751]&m[754]&~m[755]&m[756]&m[757])|(m[751]&m[754]&~m[755]&m[756]&m[757])|(~m[751]&~m[754]&m[755]&m[756]&m[757])|(m[751]&~m[754]&m[755]&m[756]&m[757])|(m[751]&m[754]&m[755]&m[756]&m[757]));
    m[758] = (((m[536]&~m[759]&~m[760]&~m[761]&~m[762])|(~m[536]&~m[759]&~m[760]&m[761]&~m[762])|(m[536]&m[759]&~m[760]&m[761]&~m[762])|(m[536]&~m[759]&m[760]&m[761]&~m[762])|(~m[536]&m[759]&~m[760]&~m[761]&m[762])|(~m[536]&~m[759]&m[760]&~m[761]&m[762])|(m[536]&m[759]&m[760]&~m[761]&m[762])|(~m[536]&m[759]&m[760]&m[761]&m[762]))&UnbiasedRNG[34])|((m[536]&~m[759]&~m[760]&m[761]&~m[762])|(~m[536]&~m[759]&~m[760]&~m[761]&m[762])|(m[536]&~m[759]&~m[760]&~m[761]&m[762])|(m[536]&m[759]&~m[760]&~m[761]&m[762])|(m[536]&~m[759]&m[760]&~m[761]&m[762])|(~m[536]&~m[759]&~m[760]&m[761]&m[762])|(m[536]&~m[759]&~m[760]&m[761]&m[762])|(~m[536]&m[759]&~m[760]&m[761]&m[762])|(m[536]&m[759]&~m[760]&m[761]&m[762])|(~m[536]&~m[759]&m[760]&m[761]&m[762])|(m[536]&~m[759]&m[760]&m[761]&m[762])|(m[536]&m[759]&m[760]&m[761]&m[762]));
    m[763] = (((m[761]&~m[764]&~m[765]&~m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&m[766]&~m[767])|(m[761]&m[764]&~m[765]&m[766]&~m[767])|(m[761]&~m[764]&m[765]&m[766]&~m[767])|(~m[761]&m[764]&~m[765]&~m[766]&m[767])|(~m[761]&~m[764]&m[765]&~m[766]&m[767])|(m[761]&m[764]&m[765]&~m[766]&m[767])|(~m[761]&m[764]&m[765]&m[766]&m[767]))&UnbiasedRNG[35])|((m[761]&~m[764]&~m[765]&m[766]&~m[767])|(~m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&~m[765]&~m[766]&m[767])|(m[761]&m[764]&~m[765]&~m[766]&m[767])|(m[761]&~m[764]&m[765]&~m[766]&m[767])|(~m[761]&~m[764]&~m[765]&m[766]&m[767])|(m[761]&~m[764]&~m[765]&m[766]&m[767])|(~m[761]&m[764]&~m[765]&m[766]&m[767])|(m[761]&m[764]&~m[765]&m[766]&m[767])|(~m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&~m[764]&m[765]&m[766]&m[767])|(m[761]&m[764]&m[765]&m[766]&m[767]));
    m[768] = (((m[766]&~m[769]&~m[770]&~m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&m[771]&~m[772])|(m[766]&m[769]&~m[770]&m[771]&~m[772])|(m[766]&~m[769]&m[770]&m[771]&~m[772])|(~m[766]&m[769]&~m[770]&~m[771]&m[772])|(~m[766]&~m[769]&m[770]&~m[771]&m[772])|(m[766]&m[769]&m[770]&~m[771]&m[772])|(~m[766]&m[769]&m[770]&m[771]&m[772]))&UnbiasedRNG[36])|((m[766]&~m[769]&~m[770]&m[771]&~m[772])|(~m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&~m[770]&~m[771]&m[772])|(m[766]&m[769]&~m[770]&~m[771]&m[772])|(m[766]&~m[769]&m[770]&~m[771]&m[772])|(~m[766]&~m[769]&~m[770]&m[771]&m[772])|(m[766]&~m[769]&~m[770]&m[771]&m[772])|(~m[766]&m[769]&~m[770]&m[771]&m[772])|(m[766]&m[769]&~m[770]&m[771]&m[772])|(~m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&~m[769]&m[770]&m[771]&m[772])|(m[766]&m[769]&m[770]&m[771]&m[772]));
    m[773] = (((m[771]&~m[774]&~m[775]&~m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&m[776]&~m[777])|(m[771]&m[774]&~m[775]&m[776]&~m[777])|(m[771]&~m[774]&m[775]&m[776]&~m[777])|(~m[771]&m[774]&~m[775]&~m[776]&m[777])|(~m[771]&~m[774]&m[775]&~m[776]&m[777])|(m[771]&m[774]&m[775]&~m[776]&m[777])|(~m[771]&m[774]&m[775]&m[776]&m[777]))&UnbiasedRNG[37])|((m[771]&~m[774]&~m[775]&m[776]&~m[777])|(~m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&~m[775]&~m[776]&m[777])|(m[771]&m[774]&~m[775]&~m[776]&m[777])|(m[771]&~m[774]&m[775]&~m[776]&m[777])|(~m[771]&~m[774]&~m[775]&m[776]&m[777])|(m[771]&~m[774]&~m[775]&m[776]&m[777])|(~m[771]&m[774]&~m[775]&m[776]&m[777])|(m[771]&m[774]&~m[775]&m[776]&m[777])|(~m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&~m[774]&m[775]&m[776]&m[777])|(m[771]&m[774]&m[775]&m[776]&m[777]));
    m[778] = (((m[537]&~m[779]&~m[780]&~m[781]&~m[782])|(~m[537]&~m[779]&~m[780]&m[781]&~m[782])|(m[537]&m[779]&~m[780]&m[781]&~m[782])|(m[537]&~m[779]&m[780]&m[781]&~m[782])|(~m[537]&m[779]&~m[780]&~m[781]&m[782])|(~m[537]&~m[779]&m[780]&~m[781]&m[782])|(m[537]&m[779]&m[780]&~m[781]&m[782])|(~m[537]&m[779]&m[780]&m[781]&m[782]))&UnbiasedRNG[38])|((m[537]&~m[779]&~m[780]&m[781]&~m[782])|(~m[537]&~m[779]&~m[780]&~m[781]&m[782])|(m[537]&~m[779]&~m[780]&~m[781]&m[782])|(m[537]&m[779]&~m[780]&~m[781]&m[782])|(m[537]&~m[779]&m[780]&~m[781]&m[782])|(~m[537]&~m[779]&~m[780]&m[781]&m[782])|(m[537]&~m[779]&~m[780]&m[781]&m[782])|(~m[537]&m[779]&~m[780]&m[781]&m[782])|(m[537]&m[779]&~m[780]&m[781]&m[782])|(~m[537]&~m[779]&m[780]&m[781]&m[782])|(m[537]&~m[779]&m[780]&m[781]&m[782])|(m[537]&m[779]&m[780]&m[781]&m[782]));
    m[783] = (((m[781]&~m[784]&~m[785]&~m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&m[786]&~m[787])|(m[781]&m[784]&~m[785]&m[786]&~m[787])|(m[781]&~m[784]&m[785]&m[786]&~m[787])|(~m[781]&m[784]&~m[785]&~m[786]&m[787])|(~m[781]&~m[784]&m[785]&~m[786]&m[787])|(m[781]&m[784]&m[785]&~m[786]&m[787])|(~m[781]&m[784]&m[785]&m[786]&m[787]))&UnbiasedRNG[39])|((m[781]&~m[784]&~m[785]&m[786]&~m[787])|(~m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&~m[785]&~m[786]&m[787])|(m[781]&m[784]&~m[785]&~m[786]&m[787])|(m[781]&~m[784]&m[785]&~m[786]&m[787])|(~m[781]&~m[784]&~m[785]&m[786]&m[787])|(m[781]&~m[784]&~m[785]&m[786]&m[787])|(~m[781]&m[784]&~m[785]&m[786]&m[787])|(m[781]&m[784]&~m[785]&m[786]&m[787])|(~m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&~m[784]&m[785]&m[786]&m[787])|(m[781]&m[784]&m[785]&m[786]&m[787]));
    m[788] = (((m[786]&~m[789]&~m[790]&~m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&m[791]&~m[792])|(m[786]&m[789]&~m[790]&m[791]&~m[792])|(m[786]&~m[789]&m[790]&m[791]&~m[792])|(~m[786]&m[789]&~m[790]&~m[791]&m[792])|(~m[786]&~m[789]&m[790]&~m[791]&m[792])|(m[786]&m[789]&m[790]&~m[791]&m[792])|(~m[786]&m[789]&m[790]&m[791]&m[792]))&UnbiasedRNG[40])|((m[786]&~m[789]&~m[790]&m[791]&~m[792])|(~m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&~m[790]&~m[791]&m[792])|(m[786]&m[789]&~m[790]&~m[791]&m[792])|(m[786]&~m[789]&m[790]&~m[791]&m[792])|(~m[786]&~m[789]&~m[790]&m[791]&m[792])|(m[786]&~m[789]&~m[790]&m[791]&m[792])|(~m[786]&m[789]&~m[790]&m[791]&m[792])|(m[786]&m[789]&~m[790]&m[791]&m[792])|(~m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&~m[789]&m[790]&m[791]&m[792])|(m[786]&m[789]&m[790]&m[791]&m[792]));
    m[793] = (((m[791]&~m[794]&~m[795]&~m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&m[796]&~m[797])|(m[791]&m[794]&~m[795]&m[796]&~m[797])|(m[791]&~m[794]&m[795]&m[796]&~m[797])|(~m[791]&m[794]&~m[795]&~m[796]&m[797])|(~m[791]&~m[794]&m[795]&~m[796]&m[797])|(m[791]&m[794]&m[795]&~m[796]&m[797])|(~m[791]&m[794]&m[795]&m[796]&m[797]))&UnbiasedRNG[41])|((m[791]&~m[794]&~m[795]&m[796]&~m[797])|(~m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&~m[795]&~m[796]&m[797])|(m[791]&m[794]&~m[795]&~m[796]&m[797])|(m[791]&~m[794]&m[795]&~m[796]&m[797])|(~m[791]&~m[794]&~m[795]&m[796]&m[797])|(m[791]&~m[794]&~m[795]&m[796]&m[797])|(~m[791]&m[794]&~m[795]&m[796]&m[797])|(m[791]&m[794]&~m[795]&m[796]&m[797])|(~m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&~m[794]&m[795]&m[796]&m[797])|(m[791]&m[794]&m[795]&m[796]&m[797]));
    m[798] = (((m[796]&~m[799]&~m[800]&~m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&m[801]&~m[802])|(m[796]&m[799]&~m[800]&m[801]&~m[802])|(m[796]&~m[799]&m[800]&m[801]&~m[802])|(~m[796]&m[799]&~m[800]&~m[801]&m[802])|(~m[796]&~m[799]&m[800]&~m[801]&m[802])|(m[796]&m[799]&m[800]&~m[801]&m[802])|(~m[796]&m[799]&m[800]&m[801]&m[802]))&UnbiasedRNG[42])|((m[796]&~m[799]&~m[800]&m[801]&~m[802])|(~m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&~m[800]&~m[801]&m[802])|(m[796]&m[799]&~m[800]&~m[801]&m[802])|(m[796]&~m[799]&m[800]&~m[801]&m[802])|(~m[796]&~m[799]&~m[800]&m[801]&m[802])|(m[796]&~m[799]&~m[800]&m[801]&m[802])|(~m[796]&m[799]&~m[800]&m[801]&m[802])|(m[796]&m[799]&~m[800]&m[801]&m[802])|(~m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&~m[799]&m[800]&m[801]&m[802])|(m[796]&m[799]&m[800]&m[801]&m[802]));
    m[803] = (((m[538]&~m[804]&~m[805]&~m[806]&~m[807])|(~m[538]&~m[804]&~m[805]&m[806]&~m[807])|(m[538]&m[804]&~m[805]&m[806]&~m[807])|(m[538]&~m[804]&m[805]&m[806]&~m[807])|(~m[538]&m[804]&~m[805]&~m[806]&m[807])|(~m[538]&~m[804]&m[805]&~m[806]&m[807])|(m[538]&m[804]&m[805]&~m[806]&m[807])|(~m[538]&m[804]&m[805]&m[806]&m[807]))&UnbiasedRNG[43])|((m[538]&~m[804]&~m[805]&m[806]&~m[807])|(~m[538]&~m[804]&~m[805]&~m[806]&m[807])|(m[538]&~m[804]&~m[805]&~m[806]&m[807])|(m[538]&m[804]&~m[805]&~m[806]&m[807])|(m[538]&~m[804]&m[805]&~m[806]&m[807])|(~m[538]&~m[804]&~m[805]&m[806]&m[807])|(m[538]&~m[804]&~m[805]&m[806]&m[807])|(~m[538]&m[804]&~m[805]&m[806]&m[807])|(m[538]&m[804]&~m[805]&m[806]&m[807])|(~m[538]&~m[804]&m[805]&m[806]&m[807])|(m[538]&~m[804]&m[805]&m[806]&m[807])|(m[538]&m[804]&m[805]&m[806]&m[807]));
    m[808] = (((m[806]&~m[809]&~m[810]&~m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&m[811]&~m[812])|(m[806]&m[809]&~m[810]&m[811]&~m[812])|(m[806]&~m[809]&m[810]&m[811]&~m[812])|(~m[806]&m[809]&~m[810]&~m[811]&m[812])|(~m[806]&~m[809]&m[810]&~m[811]&m[812])|(m[806]&m[809]&m[810]&~m[811]&m[812])|(~m[806]&m[809]&m[810]&m[811]&m[812]))&UnbiasedRNG[44])|((m[806]&~m[809]&~m[810]&m[811]&~m[812])|(~m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&~m[810]&~m[811]&m[812])|(m[806]&m[809]&~m[810]&~m[811]&m[812])|(m[806]&~m[809]&m[810]&~m[811]&m[812])|(~m[806]&~m[809]&~m[810]&m[811]&m[812])|(m[806]&~m[809]&~m[810]&m[811]&m[812])|(~m[806]&m[809]&~m[810]&m[811]&m[812])|(m[806]&m[809]&~m[810]&m[811]&m[812])|(~m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&~m[809]&m[810]&m[811]&m[812])|(m[806]&m[809]&m[810]&m[811]&m[812]));
    m[813] = (((m[811]&~m[814]&~m[815]&~m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&m[816]&~m[817])|(m[811]&m[814]&~m[815]&m[816]&~m[817])|(m[811]&~m[814]&m[815]&m[816]&~m[817])|(~m[811]&m[814]&~m[815]&~m[816]&m[817])|(~m[811]&~m[814]&m[815]&~m[816]&m[817])|(m[811]&m[814]&m[815]&~m[816]&m[817])|(~m[811]&m[814]&m[815]&m[816]&m[817]))&UnbiasedRNG[45])|((m[811]&~m[814]&~m[815]&m[816]&~m[817])|(~m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&~m[815]&~m[816]&m[817])|(m[811]&m[814]&~m[815]&~m[816]&m[817])|(m[811]&~m[814]&m[815]&~m[816]&m[817])|(~m[811]&~m[814]&~m[815]&m[816]&m[817])|(m[811]&~m[814]&~m[815]&m[816]&m[817])|(~m[811]&m[814]&~m[815]&m[816]&m[817])|(m[811]&m[814]&~m[815]&m[816]&m[817])|(~m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&~m[814]&m[815]&m[816]&m[817])|(m[811]&m[814]&m[815]&m[816]&m[817]));
    m[818] = (((m[816]&~m[819]&~m[820]&~m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&m[821]&~m[822])|(m[816]&m[819]&~m[820]&m[821]&~m[822])|(m[816]&~m[819]&m[820]&m[821]&~m[822])|(~m[816]&m[819]&~m[820]&~m[821]&m[822])|(~m[816]&~m[819]&m[820]&~m[821]&m[822])|(m[816]&m[819]&m[820]&~m[821]&m[822])|(~m[816]&m[819]&m[820]&m[821]&m[822]))&UnbiasedRNG[46])|((m[816]&~m[819]&~m[820]&m[821]&~m[822])|(~m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&~m[820]&~m[821]&m[822])|(m[816]&m[819]&~m[820]&~m[821]&m[822])|(m[816]&~m[819]&m[820]&~m[821]&m[822])|(~m[816]&~m[819]&~m[820]&m[821]&m[822])|(m[816]&~m[819]&~m[820]&m[821]&m[822])|(~m[816]&m[819]&~m[820]&m[821]&m[822])|(m[816]&m[819]&~m[820]&m[821]&m[822])|(~m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&~m[819]&m[820]&m[821]&m[822])|(m[816]&m[819]&m[820]&m[821]&m[822]));
    m[823] = (((m[821]&~m[824]&~m[825]&~m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&m[826]&~m[827])|(m[821]&m[824]&~m[825]&m[826]&~m[827])|(m[821]&~m[824]&m[825]&m[826]&~m[827])|(~m[821]&m[824]&~m[825]&~m[826]&m[827])|(~m[821]&~m[824]&m[825]&~m[826]&m[827])|(m[821]&m[824]&m[825]&~m[826]&m[827])|(~m[821]&m[824]&m[825]&m[826]&m[827]))&UnbiasedRNG[47])|((m[821]&~m[824]&~m[825]&m[826]&~m[827])|(~m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&~m[825]&~m[826]&m[827])|(m[821]&m[824]&~m[825]&~m[826]&m[827])|(m[821]&~m[824]&m[825]&~m[826]&m[827])|(~m[821]&~m[824]&~m[825]&m[826]&m[827])|(m[821]&~m[824]&~m[825]&m[826]&m[827])|(~m[821]&m[824]&~m[825]&m[826]&m[827])|(m[821]&m[824]&~m[825]&m[826]&m[827])|(~m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&~m[824]&m[825]&m[826]&m[827])|(m[821]&m[824]&m[825]&m[826]&m[827]));
    m[828] = (((m[826]&~m[829]&~m[830]&~m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&m[831]&~m[832])|(m[826]&m[829]&~m[830]&m[831]&~m[832])|(m[826]&~m[829]&m[830]&m[831]&~m[832])|(~m[826]&m[829]&~m[830]&~m[831]&m[832])|(~m[826]&~m[829]&m[830]&~m[831]&m[832])|(m[826]&m[829]&m[830]&~m[831]&m[832])|(~m[826]&m[829]&m[830]&m[831]&m[832]))&UnbiasedRNG[48])|((m[826]&~m[829]&~m[830]&m[831]&~m[832])|(~m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&~m[830]&~m[831]&m[832])|(m[826]&m[829]&~m[830]&~m[831]&m[832])|(m[826]&~m[829]&m[830]&~m[831]&m[832])|(~m[826]&~m[829]&~m[830]&m[831]&m[832])|(m[826]&~m[829]&~m[830]&m[831]&m[832])|(~m[826]&m[829]&~m[830]&m[831]&m[832])|(m[826]&m[829]&~m[830]&m[831]&m[832])|(~m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&~m[829]&m[830]&m[831]&m[832])|(m[826]&m[829]&m[830]&m[831]&m[832]));
    m[833] = (((m[539]&~m[834]&~m[835]&~m[836]&~m[837])|(~m[539]&~m[834]&~m[835]&m[836]&~m[837])|(m[539]&m[834]&~m[835]&m[836]&~m[837])|(m[539]&~m[834]&m[835]&m[836]&~m[837])|(~m[539]&m[834]&~m[835]&~m[836]&m[837])|(~m[539]&~m[834]&m[835]&~m[836]&m[837])|(m[539]&m[834]&m[835]&~m[836]&m[837])|(~m[539]&m[834]&m[835]&m[836]&m[837]))&UnbiasedRNG[49])|((m[539]&~m[834]&~m[835]&m[836]&~m[837])|(~m[539]&~m[834]&~m[835]&~m[836]&m[837])|(m[539]&~m[834]&~m[835]&~m[836]&m[837])|(m[539]&m[834]&~m[835]&~m[836]&m[837])|(m[539]&~m[834]&m[835]&~m[836]&m[837])|(~m[539]&~m[834]&~m[835]&m[836]&m[837])|(m[539]&~m[834]&~m[835]&m[836]&m[837])|(~m[539]&m[834]&~m[835]&m[836]&m[837])|(m[539]&m[834]&~m[835]&m[836]&m[837])|(~m[539]&~m[834]&m[835]&m[836]&m[837])|(m[539]&~m[834]&m[835]&m[836]&m[837])|(m[539]&m[834]&m[835]&m[836]&m[837]));
    m[838] = (((m[836]&~m[839]&~m[840]&~m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&m[841]&~m[842])|(m[836]&m[839]&~m[840]&m[841]&~m[842])|(m[836]&~m[839]&m[840]&m[841]&~m[842])|(~m[836]&m[839]&~m[840]&~m[841]&m[842])|(~m[836]&~m[839]&m[840]&~m[841]&m[842])|(m[836]&m[839]&m[840]&~m[841]&m[842])|(~m[836]&m[839]&m[840]&m[841]&m[842]))&UnbiasedRNG[50])|((m[836]&~m[839]&~m[840]&m[841]&~m[842])|(~m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&~m[840]&~m[841]&m[842])|(m[836]&m[839]&~m[840]&~m[841]&m[842])|(m[836]&~m[839]&m[840]&~m[841]&m[842])|(~m[836]&~m[839]&~m[840]&m[841]&m[842])|(m[836]&~m[839]&~m[840]&m[841]&m[842])|(~m[836]&m[839]&~m[840]&m[841]&m[842])|(m[836]&m[839]&~m[840]&m[841]&m[842])|(~m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&~m[839]&m[840]&m[841]&m[842])|(m[836]&m[839]&m[840]&m[841]&m[842]));
    m[843] = (((m[841]&~m[844]&~m[845]&~m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&m[846]&~m[847])|(m[841]&m[844]&~m[845]&m[846]&~m[847])|(m[841]&~m[844]&m[845]&m[846]&~m[847])|(~m[841]&m[844]&~m[845]&~m[846]&m[847])|(~m[841]&~m[844]&m[845]&~m[846]&m[847])|(m[841]&m[844]&m[845]&~m[846]&m[847])|(~m[841]&m[844]&m[845]&m[846]&m[847]))&UnbiasedRNG[51])|((m[841]&~m[844]&~m[845]&m[846]&~m[847])|(~m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&~m[845]&~m[846]&m[847])|(m[841]&m[844]&~m[845]&~m[846]&m[847])|(m[841]&~m[844]&m[845]&~m[846]&m[847])|(~m[841]&~m[844]&~m[845]&m[846]&m[847])|(m[841]&~m[844]&~m[845]&m[846]&m[847])|(~m[841]&m[844]&~m[845]&m[846]&m[847])|(m[841]&m[844]&~m[845]&m[846]&m[847])|(~m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&~m[844]&m[845]&m[846]&m[847])|(m[841]&m[844]&m[845]&m[846]&m[847]));
    m[848] = (((m[846]&~m[849]&~m[850]&~m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&m[851]&~m[852])|(m[846]&m[849]&~m[850]&m[851]&~m[852])|(m[846]&~m[849]&m[850]&m[851]&~m[852])|(~m[846]&m[849]&~m[850]&~m[851]&m[852])|(~m[846]&~m[849]&m[850]&~m[851]&m[852])|(m[846]&m[849]&m[850]&~m[851]&m[852])|(~m[846]&m[849]&m[850]&m[851]&m[852]))&UnbiasedRNG[52])|((m[846]&~m[849]&~m[850]&m[851]&~m[852])|(~m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&~m[850]&~m[851]&m[852])|(m[846]&m[849]&~m[850]&~m[851]&m[852])|(m[846]&~m[849]&m[850]&~m[851]&m[852])|(~m[846]&~m[849]&~m[850]&m[851]&m[852])|(m[846]&~m[849]&~m[850]&m[851]&m[852])|(~m[846]&m[849]&~m[850]&m[851]&m[852])|(m[846]&m[849]&~m[850]&m[851]&m[852])|(~m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&~m[849]&m[850]&m[851]&m[852])|(m[846]&m[849]&m[850]&m[851]&m[852]));
    m[853] = (((m[851]&~m[854]&~m[855]&~m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&m[856]&~m[857])|(m[851]&m[854]&~m[855]&m[856]&~m[857])|(m[851]&~m[854]&m[855]&m[856]&~m[857])|(~m[851]&m[854]&~m[855]&~m[856]&m[857])|(~m[851]&~m[854]&m[855]&~m[856]&m[857])|(m[851]&m[854]&m[855]&~m[856]&m[857])|(~m[851]&m[854]&m[855]&m[856]&m[857]))&UnbiasedRNG[53])|((m[851]&~m[854]&~m[855]&m[856]&~m[857])|(~m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&~m[855]&~m[856]&m[857])|(m[851]&m[854]&~m[855]&~m[856]&m[857])|(m[851]&~m[854]&m[855]&~m[856]&m[857])|(~m[851]&~m[854]&~m[855]&m[856]&m[857])|(m[851]&~m[854]&~m[855]&m[856]&m[857])|(~m[851]&m[854]&~m[855]&m[856]&m[857])|(m[851]&m[854]&~m[855]&m[856]&m[857])|(~m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&~m[854]&m[855]&m[856]&m[857])|(m[851]&m[854]&m[855]&m[856]&m[857]));
    m[858] = (((m[856]&~m[859]&~m[860]&~m[861]&~m[862])|(~m[856]&~m[859]&~m[860]&m[861]&~m[862])|(m[856]&m[859]&~m[860]&m[861]&~m[862])|(m[856]&~m[859]&m[860]&m[861]&~m[862])|(~m[856]&m[859]&~m[860]&~m[861]&m[862])|(~m[856]&~m[859]&m[860]&~m[861]&m[862])|(m[856]&m[859]&m[860]&~m[861]&m[862])|(~m[856]&m[859]&m[860]&m[861]&m[862]))&UnbiasedRNG[54])|((m[856]&~m[859]&~m[860]&m[861]&~m[862])|(~m[856]&~m[859]&~m[860]&~m[861]&m[862])|(m[856]&~m[859]&~m[860]&~m[861]&m[862])|(m[856]&m[859]&~m[860]&~m[861]&m[862])|(m[856]&~m[859]&m[860]&~m[861]&m[862])|(~m[856]&~m[859]&~m[860]&m[861]&m[862])|(m[856]&~m[859]&~m[860]&m[861]&m[862])|(~m[856]&m[859]&~m[860]&m[861]&m[862])|(m[856]&m[859]&~m[860]&m[861]&m[862])|(~m[856]&~m[859]&m[860]&m[861]&m[862])|(m[856]&~m[859]&m[860]&m[861]&m[862])|(m[856]&m[859]&m[860]&m[861]&m[862]));
    m[863] = (((m[861]&~m[864]&~m[865]&~m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&m[866]&~m[867])|(m[861]&m[864]&~m[865]&m[866]&~m[867])|(m[861]&~m[864]&m[865]&m[866]&~m[867])|(~m[861]&m[864]&~m[865]&~m[866]&m[867])|(~m[861]&~m[864]&m[865]&~m[866]&m[867])|(m[861]&m[864]&m[865]&~m[866]&m[867])|(~m[861]&m[864]&m[865]&m[866]&m[867]))&UnbiasedRNG[55])|((m[861]&~m[864]&~m[865]&m[866]&~m[867])|(~m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&~m[865]&~m[866]&m[867])|(m[861]&m[864]&~m[865]&~m[866]&m[867])|(m[861]&~m[864]&m[865]&~m[866]&m[867])|(~m[861]&~m[864]&~m[865]&m[866]&m[867])|(m[861]&~m[864]&~m[865]&m[866]&m[867])|(~m[861]&m[864]&~m[865]&m[866]&m[867])|(m[861]&m[864]&~m[865]&m[866]&m[867])|(~m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&~m[864]&m[865]&m[866]&m[867])|(m[861]&m[864]&m[865]&m[866]&m[867]));
    m[868] = (((m[540]&~m[869]&~m[870]&~m[871]&~m[872])|(~m[540]&~m[869]&~m[870]&m[871]&~m[872])|(m[540]&m[869]&~m[870]&m[871]&~m[872])|(m[540]&~m[869]&m[870]&m[871]&~m[872])|(~m[540]&m[869]&~m[870]&~m[871]&m[872])|(~m[540]&~m[869]&m[870]&~m[871]&m[872])|(m[540]&m[869]&m[870]&~m[871]&m[872])|(~m[540]&m[869]&m[870]&m[871]&m[872]))&UnbiasedRNG[56])|((m[540]&~m[869]&~m[870]&m[871]&~m[872])|(~m[540]&~m[869]&~m[870]&~m[871]&m[872])|(m[540]&~m[869]&~m[870]&~m[871]&m[872])|(m[540]&m[869]&~m[870]&~m[871]&m[872])|(m[540]&~m[869]&m[870]&~m[871]&m[872])|(~m[540]&~m[869]&~m[870]&m[871]&m[872])|(m[540]&~m[869]&~m[870]&m[871]&m[872])|(~m[540]&m[869]&~m[870]&m[871]&m[872])|(m[540]&m[869]&~m[870]&m[871]&m[872])|(~m[540]&~m[869]&m[870]&m[871]&m[872])|(m[540]&~m[869]&m[870]&m[871]&m[872])|(m[540]&m[869]&m[870]&m[871]&m[872]));
    m[873] = (((m[871]&~m[874]&~m[875]&~m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&m[876]&~m[877])|(m[871]&m[874]&~m[875]&m[876]&~m[877])|(m[871]&~m[874]&m[875]&m[876]&~m[877])|(~m[871]&m[874]&~m[875]&~m[876]&m[877])|(~m[871]&~m[874]&m[875]&~m[876]&m[877])|(m[871]&m[874]&m[875]&~m[876]&m[877])|(~m[871]&m[874]&m[875]&m[876]&m[877]))&UnbiasedRNG[57])|((m[871]&~m[874]&~m[875]&m[876]&~m[877])|(~m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&~m[875]&~m[876]&m[877])|(m[871]&m[874]&~m[875]&~m[876]&m[877])|(m[871]&~m[874]&m[875]&~m[876]&m[877])|(~m[871]&~m[874]&~m[875]&m[876]&m[877])|(m[871]&~m[874]&~m[875]&m[876]&m[877])|(~m[871]&m[874]&~m[875]&m[876]&m[877])|(m[871]&m[874]&~m[875]&m[876]&m[877])|(~m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&~m[874]&m[875]&m[876]&m[877])|(m[871]&m[874]&m[875]&m[876]&m[877]));
    m[878] = (((m[876]&~m[879]&~m[880]&~m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&m[881]&~m[882])|(m[876]&m[879]&~m[880]&m[881]&~m[882])|(m[876]&~m[879]&m[880]&m[881]&~m[882])|(~m[876]&m[879]&~m[880]&~m[881]&m[882])|(~m[876]&~m[879]&m[880]&~m[881]&m[882])|(m[876]&m[879]&m[880]&~m[881]&m[882])|(~m[876]&m[879]&m[880]&m[881]&m[882]))&UnbiasedRNG[58])|((m[876]&~m[879]&~m[880]&m[881]&~m[882])|(~m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&~m[880]&~m[881]&m[882])|(m[876]&m[879]&~m[880]&~m[881]&m[882])|(m[876]&~m[879]&m[880]&~m[881]&m[882])|(~m[876]&~m[879]&~m[880]&m[881]&m[882])|(m[876]&~m[879]&~m[880]&m[881]&m[882])|(~m[876]&m[879]&~m[880]&m[881]&m[882])|(m[876]&m[879]&~m[880]&m[881]&m[882])|(~m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&~m[879]&m[880]&m[881]&m[882])|(m[876]&m[879]&m[880]&m[881]&m[882]));
    m[883] = (((m[881]&~m[884]&~m[885]&~m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&m[886]&~m[887])|(m[881]&m[884]&~m[885]&m[886]&~m[887])|(m[881]&~m[884]&m[885]&m[886]&~m[887])|(~m[881]&m[884]&~m[885]&~m[886]&m[887])|(~m[881]&~m[884]&m[885]&~m[886]&m[887])|(m[881]&m[884]&m[885]&~m[886]&m[887])|(~m[881]&m[884]&m[885]&m[886]&m[887]))&UnbiasedRNG[59])|((m[881]&~m[884]&~m[885]&m[886]&~m[887])|(~m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&~m[885]&~m[886]&m[887])|(m[881]&m[884]&~m[885]&~m[886]&m[887])|(m[881]&~m[884]&m[885]&~m[886]&m[887])|(~m[881]&~m[884]&~m[885]&m[886]&m[887])|(m[881]&~m[884]&~m[885]&m[886]&m[887])|(~m[881]&m[884]&~m[885]&m[886]&m[887])|(m[881]&m[884]&~m[885]&m[886]&m[887])|(~m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&~m[884]&m[885]&m[886]&m[887])|(m[881]&m[884]&m[885]&m[886]&m[887]));
    m[888] = (((m[886]&~m[889]&~m[890]&~m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&m[891]&~m[892])|(m[886]&m[889]&~m[890]&m[891]&~m[892])|(m[886]&~m[889]&m[890]&m[891]&~m[892])|(~m[886]&m[889]&~m[890]&~m[891]&m[892])|(~m[886]&~m[889]&m[890]&~m[891]&m[892])|(m[886]&m[889]&m[890]&~m[891]&m[892])|(~m[886]&m[889]&m[890]&m[891]&m[892]))&UnbiasedRNG[60])|((m[886]&~m[889]&~m[890]&m[891]&~m[892])|(~m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&~m[890]&~m[891]&m[892])|(m[886]&m[889]&~m[890]&~m[891]&m[892])|(m[886]&~m[889]&m[890]&~m[891]&m[892])|(~m[886]&~m[889]&~m[890]&m[891]&m[892])|(m[886]&~m[889]&~m[890]&m[891]&m[892])|(~m[886]&m[889]&~m[890]&m[891]&m[892])|(m[886]&m[889]&~m[890]&m[891]&m[892])|(~m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&~m[889]&m[890]&m[891]&m[892])|(m[886]&m[889]&m[890]&m[891]&m[892]));
    m[893] = (((m[891]&~m[894]&~m[895]&~m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&m[896]&~m[897])|(m[891]&m[894]&~m[895]&m[896]&~m[897])|(m[891]&~m[894]&m[895]&m[896]&~m[897])|(~m[891]&m[894]&~m[895]&~m[896]&m[897])|(~m[891]&~m[894]&m[895]&~m[896]&m[897])|(m[891]&m[894]&m[895]&~m[896]&m[897])|(~m[891]&m[894]&m[895]&m[896]&m[897]))&UnbiasedRNG[61])|((m[891]&~m[894]&~m[895]&m[896]&~m[897])|(~m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&~m[895]&~m[896]&m[897])|(m[891]&m[894]&~m[895]&~m[896]&m[897])|(m[891]&~m[894]&m[895]&~m[896]&m[897])|(~m[891]&~m[894]&~m[895]&m[896]&m[897])|(m[891]&~m[894]&~m[895]&m[896]&m[897])|(~m[891]&m[894]&~m[895]&m[896]&m[897])|(m[891]&m[894]&~m[895]&m[896]&m[897])|(~m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&~m[894]&m[895]&m[896]&m[897])|(m[891]&m[894]&m[895]&m[896]&m[897]));
    m[898] = (((m[896]&~m[899]&~m[900]&~m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&m[901]&~m[902])|(m[896]&m[899]&~m[900]&m[901]&~m[902])|(m[896]&~m[899]&m[900]&m[901]&~m[902])|(~m[896]&m[899]&~m[900]&~m[901]&m[902])|(~m[896]&~m[899]&m[900]&~m[901]&m[902])|(m[896]&m[899]&m[900]&~m[901]&m[902])|(~m[896]&m[899]&m[900]&m[901]&m[902]))&UnbiasedRNG[62])|((m[896]&~m[899]&~m[900]&m[901]&~m[902])|(~m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&~m[900]&~m[901]&m[902])|(m[896]&m[899]&~m[900]&~m[901]&m[902])|(m[896]&~m[899]&m[900]&~m[901]&m[902])|(~m[896]&~m[899]&~m[900]&m[901]&m[902])|(m[896]&~m[899]&~m[900]&m[901]&m[902])|(~m[896]&m[899]&~m[900]&m[901]&m[902])|(m[896]&m[899]&~m[900]&m[901]&m[902])|(~m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&~m[899]&m[900]&m[901]&m[902])|(m[896]&m[899]&m[900]&m[901]&m[902]));
    m[903] = (((m[901]&~m[904]&~m[905]&~m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&m[906]&~m[907])|(m[901]&m[904]&~m[905]&m[906]&~m[907])|(m[901]&~m[904]&m[905]&m[906]&~m[907])|(~m[901]&m[904]&~m[905]&~m[906]&m[907])|(~m[901]&~m[904]&m[905]&~m[906]&m[907])|(m[901]&m[904]&m[905]&~m[906]&m[907])|(~m[901]&m[904]&m[905]&m[906]&m[907]))&UnbiasedRNG[63])|((m[901]&~m[904]&~m[905]&m[906]&~m[907])|(~m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&~m[905]&~m[906]&m[907])|(m[901]&m[904]&~m[905]&~m[906]&m[907])|(m[901]&~m[904]&m[905]&~m[906]&m[907])|(~m[901]&~m[904]&~m[905]&m[906]&m[907])|(m[901]&~m[904]&~m[905]&m[906]&m[907])|(~m[901]&m[904]&~m[905]&m[906]&m[907])|(m[901]&m[904]&~m[905]&m[906]&m[907])|(~m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&~m[904]&m[905]&m[906]&m[907])|(m[901]&m[904]&m[905]&m[906]&m[907]));
    m[908] = (((m[541]&~m[909]&~m[910]&~m[911]&~m[912])|(~m[541]&~m[909]&~m[910]&m[911]&~m[912])|(m[541]&m[909]&~m[910]&m[911]&~m[912])|(m[541]&~m[909]&m[910]&m[911]&~m[912])|(~m[541]&m[909]&~m[910]&~m[911]&m[912])|(~m[541]&~m[909]&m[910]&~m[911]&m[912])|(m[541]&m[909]&m[910]&~m[911]&m[912])|(~m[541]&m[909]&m[910]&m[911]&m[912]))&UnbiasedRNG[64])|((m[541]&~m[909]&~m[910]&m[911]&~m[912])|(~m[541]&~m[909]&~m[910]&~m[911]&m[912])|(m[541]&~m[909]&~m[910]&~m[911]&m[912])|(m[541]&m[909]&~m[910]&~m[911]&m[912])|(m[541]&~m[909]&m[910]&~m[911]&m[912])|(~m[541]&~m[909]&~m[910]&m[911]&m[912])|(m[541]&~m[909]&~m[910]&m[911]&m[912])|(~m[541]&m[909]&~m[910]&m[911]&m[912])|(m[541]&m[909]&~m[910]&m[911]&m[912])|(~m[541]&~m[909]&m[910]&m[911]&m[912])|(m[541]&~m[909]&m[910]&m[911]&m[912])|(m[541]&m[909]&m[910]&m[911]&m[912]));
    m[913] = (((m[911]&~m[914]&~m[915]&~m[916]&~m[917])|(~m[911]&~m[914]&~m[915]&m[916]&~m[917])|(m[911]&m[914]&~m[915]&m[916]&~m[917])|(m[911]&~m[914]&m[915]&m[916]&~m[917])|(~m[911]&m[914]&~m[915]&~m[916]&m[917])|(~m[911]&~m[914]&m[915]&~m[916]&m[917])|(m[911]&m[914]&m[915]&~m[916]&m[917])|(~m[911]&m[914]&m[915]&m[916]&m[917]))&UnbiasedRNG[65])|((m[911]&~m[914]&~m[915]&m[916]&~m[917])|(~m[911]&~m[914]&~m[915]&~m[916]&m[917])|(m[911]&~m[914]&~m[915]&~m[916]&m[917])|(m[911]&m[914]&~m[915]&~m[916]&m[917])|(m[911]&~m[914]&m[915]&~m[916]&m[917])|(~m[911]&~m[914]&~m[915]&m[916]&m[917])|(m[911]&~m[914]&~m[915]&m[916]&m[917])|(~m[911]&m[914]&~m[915]&m[916]&m[917])|(m[911]&m[914]&~m[915]&m[916]&m[917])|(~m[911]&~m[914]&m[915]&m[916]&m[917])|(m[911]&~m[914]&m[915]&m[916]&m[917])|(m[911]&m[914]&m[915]&m[916]&m[917]));
    m[918] = (((m[916]&~m[919]&~m[920]&~m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&m[921]&~m[922])|(m[916]&m[919]&~m[920]&m[921]&~m[922])|(m[916]&~m[919]&m[920]&m[921]&~m[922])|(~m[916]&m[919]&~m[920]&~m[921]&m[922])|(~m[916]&~m[919]&m[920]&~m[921]&m[922])|(m[916]&m[919]&m[920]&~m[921]&m[922])|(~m[916]&m[919]&m[920]&m[921]&m[922]))&UnbiasedRNG[66])|((m[916]&~m[919]&~m[920]&m[921]&~m[922])|(~m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&~m[920]&~m[921]&m[922])|(m[916]&m[919]&~m[920]&~m[921]&m[922])|(m[916]&~m[919]&m[920]&~m[921]&m[922])|(~m[916]&~m[919]&~m[920]&m[921]&m[922])|(m[916]&~m[919]&~m[920]&m[921]&m[922])|(~m[916]&m[919]&~m[920]&m[921]&m[922])|(m[916]&m[919]&~m[920]&m[921]&m[922])|(~m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&~m[919]&m[920]&m[921]&m[922])|(m[916]&m[919]&m[920]&m[921]&m[922]));
    m[923] = (((m[921]&~m[924]&~m[925]&~m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&m[926]&~m[927])|(m[921]&m[924]&~m[925]&m[926]&~m[927])|(m[921]&~m[924]&m[925]&m[926]&~m[927])|(~m[921]&m[924]&~m[925]&~m[926]&m[927])|(~m[921]&~m[924]&m[925]&~m[926]&m[927])|(m[921]&m[924]&m[925]&~m[926]&m[927])|(~m[921]&m[924]&m[925]&m[926]&m[927]))&UnbiasedRNG[67])|((m[921]&~m[924]&~m[925]&m[926]&~m[927])|(~m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&~m[925]&~m[926]&m[927])|(m[921]&m[924]&~m[925]&~m[926]&m[927])|(m[921]&~m[924]&m[925]&~m[926]&m[927])|(~m[921]&~m[924]&~m[925]&m[926]&m[927])|(m[921]&~m[924]&~m[925]&m[926]&m[927])|(~m[921]&m[924]&~m[925]&m[926]&m[927])|(m[921]&m[924]&~m[925]&m[926]&m[927])|(~m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&~m[924]&m[925]&m[926]&m[927])|(m[921]&m[924]&m[925]&m[926]&m[927]));
    m[928] = (((m[926]&~m[929]&~m[930]&~m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&m[931]&~m[932])|(m[926]&m[929]&~m[930]&m[931]&~m[932])|(m[926]&~m[929]&m[930]&m[931]&~m[932])|(~m[926]&m[929]&~m[930]&~m[931]&m[932])|(~m[926]&~m[929]&m[930]&~m[931]&m[932])|(m[926]&m[929]&m[930]&~m[931]&m[932])|(~m[926]&m[929]&m[930]&m[931]&m[932]))&UnbiasedRNG[68])|((m[926]&~m[929]&~m[930]&m[931]&~m[932])|(~m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&~m[930]&~m[931]&m[932])|(m[926]&m[929]&~m[930]&~m[931]&m[932])|(m[926]&~m[929]&m[930]&~m[931]&m[932])|(~m[926]&~m[929]&~m[930]&m[931]&m[932])|(m[926]&~m[929]&~m[930]&m[931]&m[932])|(~m[926]&m[929]&~m[930]&m[931]&m[932])|(m[926]&m[929]&~m[930]&m[931]&m[932])|(~m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&~m[929]&m[930]&m[931]&m[932])|(m[926]&m[929]&m[930]&m[931]&m[932]));
    m[933] = (((m[931]&~m[934]&~m[935]&~m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&m[936]&~m[937])|(m[931]&m[934]&~m[935]&m[936]&~m[937])|(m[931]&~m[934]&m[935]&m[936]&~m[937])|(~m[931]&m[934]&~m[935]&~m[936]&m[937])|(~m[931]&~m[934]&m[935]&~m[936]&m[937])|(m[931]&m[934]&m[935]&~m[936]&m[937])|(~m[931]&m[934]&m[935]&m[936]&m[937]))&UnbiasedRNG[69])|((m[931]&~m[934]&~m[935]&m[936]&~m[937])|(~m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&~m[935]&~m[936]&m[937])|(m[931]&m[934]&~m[935]&~m[936]&m[937])|(m[931]&~m[934]&m[935]&~m[936]&m[937])|(~m[931]&~m[934]&~m[935]&m[936]&m[937])|(m[931]&~m[934]&~m[935]&m[936]&m[937])|(~m[931]&m[934]&~m[935]&m[936]&m[937])|(m[931]&m[934]&~m[935]&m[936]&m[937])|(~m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&~m[934]&m[935]&m[936]&m[937])|(m[931]&m[934]&m[935]&m[936]&m[937]));
    m[938] = (((m[936]&~m[939]&~m[940]&~m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&m[941]&~m[942])|(m[936]&m[939]&~m[940]&m[941]&~m[942])|(m[936]&~m[939]&m[940]&m[941]&~m[942])|(~m[936]&m[939]&~m[940]&~m[941]&m[942])|(~m[936]&~m[939]&m[940]&~m[941]&m[942])|(m[936]&m[939]&m[940]&~m[941]&m[942])|(~m[936]&m[939]&m[940]&m[941]&m[942]))&UnbiasedRNG[70])|((m[936]&~m[939]&~m[940]&m[941]&~m[942])|(~m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&~m[940]&~m[941]&m[942])|(m[936]&m[939]&~m[940]&~m[941]&m[942])|(m[936]&~m[939]&m[940]&~m[941]&m[942])|(~m[936]&~m[939]&~m[940]&m[941]&m[942])|(m[936]&~m[939]&~m[940]&m[941]&m[942])|(~m[936]&m[939]&~m[940]&m[941]&m[942])|(m[936]&m[939]&~m[940]&m[941]&m[942])|(~m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&~m[939]&m[940]&m[941]&m[942])|(m[936]&m[939]&m[940]&m[941]&m[942]));
    m[943] = (((m[941]&~m[944]&~m[945]&~m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&m[946]&~m[947])|(m[941]&m[944]&~m[945]&m[946]&~m[947])|(m[941]&~m[944]&m[945]&m[946]&~m[947])|(~m[941]&m[944]&~m[945]&~m[946]&m[947])|(~m[941]&~m[944]&m[945]&~m[946]&m[947])|(m[941]&m[944]&m[945]&~m[946]&m[947])|(~m[941]&m[944]&m[945]&m[946]&m[947]))&UnbiasedRNG[71])|((m[941]&~m[944]&~m[945]&m[946]&~m[947])|(~m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&~m[945]&~m[946]&m[947])|(m[941]&m[944]&~m[945]&~m[946]&m[947])|(m[941]&~m[944]&m[945]&~m[946]&m[947])|(~m[941]&~m[944]&~m[945]&m[946]&m[947])|(m[941]&~m[944]&~m[945]&m[946]&m[947])|(~m[941]&m[944]&~m[945]&m[946]&m[947])|(m[941]&m[944]&~m[945]&m[946]&m[947])|(~m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&~m[944]&m[945]&m[946]&m[947])|(m[941]&m[944]&m[945]&m[946]&m[947]));
    m[948] = (((m[946]&~m[949]&~m[950]&~m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&m[951]&~m[952])|(m[946]&m[949]&~m[950]&m[951]&~m[952])|(m[946]&~m[949]&m[950]&m[951]&~m[952])|(~m[946]&m[949]&~m[950]&~m[951]&m[952])|(~m[946]&~m[949]&m[950]&~m[951]&m[952])|(m[946]&m[949]&m[950]&~m[951]&m[952])|(~m[946]&m[949]&m[950]&m[951]&m[952]))&UnbiasedRNG[72])|((m[946]&~m[949]&~m[950]&m[951]&~m[952])|(~m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&~m[950]&~m[951]&m[952])|(m[946]&m[949]&~m[950]&~m[951]&m[952])|(m[946]&~m[949]&m[950]&~m[951]&m[952])|(~m[946]&~m[949]&~m[950]&m[951]&m[952])|(m[946]&~m[949]&~m[950]&m[951]&m[952])|(~m[946]&m[949]&~m[950]&m[951]&m[952])|(m[946]&m[949]&~m[950]&m[951]&m[952])|(~m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&~m[949]&m[950]&m[951]&m[952])|(m[946]&m[949]&m[950]&m[951]&m[952]));
    m[953] = (((m[542]&~m[954]&~m[955]&~m[956]&~m[957])|(~m[542]&~m[954]&~m[955]&m[956]&~m[957])|(m[542]&m[954]&~m[955]&m[956]&~m[957])|(m[542]&~m[954]&m[955]&m[956]&~m[957])|(~m[542]&m[954]&~m[955]&~m[956]&m[957])|(~m[542]&~m[954]&m[955]&~m[956]&m[957])|(m[542]&m[954]&m[955]&~m[956]&m[957])|(~m[542]&m[954]&m[955]&m[956]&m[957]))&UnbiasedRNG[73])|((m[542]&~m[954]&~m[955]&m[956]&~m[957])|(~m[542]&~m[954]&~m[955]&~m[956]&m[957])|(m[542]&~m[954]&~m[955]&~m[956]&m[957])|(m[542]&m[954]&~m[955]&~m[956]&m[957])|(m[542]&~m[954]&m[955]&~m[956]&m[957])|(~m[542]&~m[954]&~m[955]&m[956]&m[957])|(m[542]&~m[954]&~m[955]&m[956]&m[957])|(~m[542]&m[954]&~m[955]&m[956]&m[957])|(m[542]&m[954]&~m[955]&m[956]&m[957])|(~m[542]&~m[954]&m[955]&m[956]&m[957])|(m[542]&~m[954]&m[955]&m[956]&m[957])|(m[542]&m[954]&m[955]&m[956]&m[957]));
    m[958] = (((m[956]&~m[959]&~m[960]&~m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&m[961]&~m[962])|(m[956]&m[959]&~m[960]&m[961]&~m[962])|(m[956]&~m[959]&m[960]&m[961]&~m[962])|(~m[956]&m[959]&~m[960]&~m[961]&m[962])|(~m[956]&~m[959]&m[960]&~m[961]&m[962])|(m[956]&m[959]&m[960]&~m[961]&m[962])|(~m[956]&m[959]&m[960]&m[961]&m[962]))&UnbiasedRNG[74])|((m[956]&~m[959]&~m[960]&m[961]&~m[962])|(~m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&~m[960]&~m[961]&m[962])|(m[956]&m[959]&~m[960]&~m[961]&m[962])|(m[956]&~m[959]&m[960]&~m[961]&m[962])|(~m[956]&~m[959]&~m[960]&m[961]&m[962])|(m[956]&~m[959]&~m[960]&m[961]&m[962])|(~m[956]&m[959]&~m[960]&m[961]&m[962])|(m[956]&m[959]&~m[960]&m[961]&m[962])|(~m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&~m[959]&m[960]&m[961]&m[962])|(m[956]&m[959]&m[960]&m[961]&m[962]));
    m[963] = (((m[961]&~m[964]&~m[965]&~m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&m[966]&~m[967])|(m[961]&m[964]&~m[965]&m[966]&~m[967])|(m[961]&~m[964]&m[965]&m[966]&~m[967])|(~m[961]&m[964]&~m[965]&~m[966]&m[967])|(~m[961]&~m[964]&m[965]&~m[966]&m[967])|(m[961]&m[964]&m[965]&~m[966]&m[967])|(~m[961]&m[964]&m[965]&m[966]&m[967]))&UnbiasedRNG[75])|((m[961]&~m[964]&~m[965]&m[966]&~m[967])|(~m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&~m[965]&~m[966]&m[967])|(m[961]&m[964]&~m[965]&~m[966]&m[967])|(m[961]&~m[964]&m[965]&~m[966]&m[967])|(~m[961]&~m[964]&~m[965]&m[966]&m[967])|(m[961]&~m[964]&~m[965]&m[966]&m[967])|(~m[961]&m[964]&~m[965]&m[966]&m[967])|(m[961]&m[964]&~m[965]&m[966]&m[967])|(~m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&~m[964]&m[965]&m[966]&m[967])|(m[961]&m[964]&m[965]&m[966]&m[967]));
    m[968] = (((m[966]&~m[969]&~m[970]&~m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&m[971]&~m[972])|(m[966]&m[969]&~m[970]&m[971]&~m[972])|(m[966]&~m[969]&m[970]&m[971]&~m[972])|(~m[966]&m[969]&~m[970]&~m[971]&m[972])|(~m[966]&~m[969]&m[970]&~m[971]&m[972])|(m[966]&m[969]&m[970]&~m[971]&m[972])|(~m[966]&m[969]&m[970]&m[971]&m[972]))&UnbiasedRNG[76])|((m[966]&~m[969]&~m[970]&m[971]&~m[972])|(~m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&~m[970]&~m[971]&m[972])|(m[966]&m[969]&~m[970]&~m[971]&m[972])|(m[966]&~m[969]&m[970]&~m[971]&m[972])|(~m[966]&~m[969]&~m[970]&m[971]&m[972])|(m[966]&~m[969]&~m[970]&m[971]&m[972])|(~m[966]&m[969]&~m[970]&m[971]&m[972])|(m[966]&m[969]&~m[970]&m[971]&m[972])|(~m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&~m[969]&m[970]&m[971]&m[972])|(m[966]&m[969]&m[970]&m[971]&m[972]));
    m[973] = (((m[971]&~m[974]&~m[975]&~m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&m[976]&~m[977])|(m[971]&m[974]&~m[975]&m[976]&~m[977])|(m[971]&~m[974]&m[975]&m[976]&~m[977])|(~m[971]&m[974]&~m[975]&~m[976]&m[977])|(~m[971]&~m[974]&m[975]&~m[976]&m[977])|(m[971]&m[974]&m[975]&~m[976]&m[977])|(~m[971]&m[974]&m[975]&m[976]&m[977]))&UnbiasedRNG[77])|((m[971]&~m[974]&~m[975]&m[976]&~m[977])|(~m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&~m[975]&~m[976]&m[977])|(m[971]&m[974]&~m[975]&~m[976]&m[977])|(m[971]&~m[974]&m[975]&~m[976]&m[977])|(~m[971]&~m[974]&~m[975]&m[976]&m[977])|(m[971]&~m[974]&~m[975]&m[976]&m[977])|(~m[971]&m[974]&~m[975]&m[976]&m[977])|(m[971]&m[974]&~m[975]&m[976]&m[977])|(~m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&~m[974]&m[975]&m[976]&m[977])|(m[971]&m[974]&m[975]&m[976]&m[977]));
    m[978] = (((m[976]&~m[979]&~m[980]&~m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&m[981]&~m[982])|(m[976]&m[979]&~m[980]&m[981]&~m[982])|(m[976]&~m[979]&m[980]&m[981]&~m[982])|(~m[976]&m[979]&~m[980]&~m[981]&m[982])|(~m[976]&~m[979]&m[980]&~m[981]&m[982])|(m[976]&m[979]&m[980]&~m[981]&m[982])|(~m[976]&m[979]&m[980]&m[981]&m[982]))&UnbiasedRNG[78])|((m[976]&~m[979]&~m[980]&m[981]&~m[982])|(~m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&~m[980]&~m[981]&m[982])|(m[976]&m[979]&~m[980]&~m[981]&m[982])|(m[976]&~m[979]&m[980]&~m[981]&m[982])|(~m[976]&~m[979]&~m[980]&m[981]&m[982])|(m[976]&~m[979]&~m[980]&m[981]&m[982])|(~m[976]&m[979]&~m[980]&m[981]&m[982])|(m[976]&m[979]&~m[980]&m[981]&m[982])|(~m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&~m[979]&m[980]&m[981]&m[982])|(m[976]&m[979]&m[980]&m[981]&m[982]));
    m[983] = (((m[981]&~m[984]&~m[985]&~m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&m[986]&~m[987])|(m[981]&m[984]&~m[985]&m[986]&~m[987])|(m[981]&~m[984]&m[985]&m[986]&~m[987])|(~m[981]&m[984]&~m[985]&~m[986]&m[987])|(~m[981]&~m[984]&m[985]&~m[986]&m[987])|(m[981]&m[984]&m[985]&~m[986]&m[987])|(~m[981]&m[984]&m[985]&m[986]&m[987]))&UnbiasedRNG[79])|((m[981]&~m[984]&~m[985]&m[986]&~m[987])|(~m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&~m[985]&~m[986]&m[987])|(m[981]&m[984]&~m[985]&~m[986]&m[987])|(m[981]&~m[984]&m[985]&~m[986]&m[987])|(~m[981]&~m[984]&~m[985]&m[986]&m[987])|(m[981]&~m[984]&~m[985]&m[986]&m[987])|(~m[981]&m[984]&~m[985]&m[986]&m[987])|(m[981]&m[984]&~m[985]&m[986]&m[987])|(~m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&~m[984]&m[985]&m[986]&m[987])|(m[981]&m[984]&m[985]&m[986]&m[987]));
    m[988] = (((m[986]&~m[989]&~m[990]&~m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&m[991]&~m[992])|(m[986]&m[989]&~m[990]&m[991]&~m[992])|(m[986]&~m[989]&m[990]&m[991]&~m[992])|(~m[986]&m[989]&~m[990]&~m[991]&m[992])|(~m[986]&~m[989]&m[990]&~m[991]&m[992])|(m[986]&m[989]&m[990]&~m[991]&m[992])|(~m[986]&m[989]&m[990]&m[991]&m[992]))&UnbiasedRNG[80])|((m[986]&~m[989]&~m[990]&m[991]&~m[992])|(~m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&~m[990]&~m[991]&m[992])|(m[986]&m[989]&~m[990]&~m[991]&m[992])|(m[986]&~m[989]&m[990]&~m[991]&m[992])|(~m[986]&~m[989]&~m[990]&m[991]&m[992])|(m[986]&~m[989]&~m[990]&m[991]&m[992])|(~m[986]&m[989]&~m[990]&m[991]&m[992])|(m[986]&m[989]&~m[990]&m[991]&m[992])|(~m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&~m[989]&m[990]&m[991]&m[992])|(m[986]&m[989]&m[990]&m[991]&m[992]));
    m[993] = (((m[991]&~m[994]&~m[995]&~m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&m[996]&~m[997])|(m[991]&m[994]&~m[995]&m[996]&~m[997])|(m[991]&~m[994]&m[995]&m[996]&~m[997])|(~m[991]&m[994]&~m[995]&~m[996]&m[997])|(~m[991]&~m[994]&m[995]&~m[996]&m[997])|(m[991]&m[994]&m[995]&~m[996]&m[997])|(~m[991]&m[994]&m[995]&m[996]&m[997]))&UnbiasedRNG[81])|((m[991]&~m[994]&~m[995]&m[996]&~m[997])|(~m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&~m[995]&~m[996]&m[997])|(m[991]&m[994]&~m[995]&~m[996]&m[997])|(m[991]&~m[994]&m[995]&~m[996]&m[997])|(~m[991]&~m[994]&~m[995]&m[996]&m[997])|(m[991]&~m[994]&~m[995]&m[996]&m[997])|(~m[991]&m[994]&~m[995]&m[996]&m[997])|(m[991]&m[994]&~m[995]&m[996]&m[997])|(~m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&~m[994]&m[995]&m[996]&m[997])|(m[991]&m[994]&m[995]&m[996]&m[997]));
    m[998] = (((m[996]&~m[999]&~m[1000]&~m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&~m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&~m[1002])|(~m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&m[999]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[82])|((m[996]&~m[999]&~m[1000]&m[1001]&~m[1002])|(~m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&~m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&~m[1001]&m[1002])|(~m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(m[996]&m[999]&~m[1000]&m[1001]&m[1002])|(~m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&~m[999]&m[1000]&m[1001]&m[1002])|(m[996]&m[999]&m[1000]&m[1001]&m[1002]));
    m[1003] = (((m[543]&~m[1004]&~m[1005]&~m[1006]&~m[1007])|(~m[543]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(m[543]&m[1004]&~m[1005]&m[1006]&~m[1007])|(m[543]&~m[1004]&m[1005]&m[1006]&~m[1007])|(~m[543]&m[1004]&~m[1005]&~m[1006]&m[1007])|(~m[543]&~m[1004]&m[1005]&~m[1006]&m[1007])|(m[543]&m[1004]&m[1005]&~m[1006]&m[1007])|(~m[543]&m[1004]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[83])|((m[543]&~m[1004]&~m[1005]&m[1006]&~m[1007])|(~m[543]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[543]&~m[1004]&~m[1005]&~m[1006]&m[1007])|(m[543]&m[1004]&~m[1005]&~m[1006]&m[1007])|(m[543]&~m[1004]&m[1005]&~m[1006]&m[1007])|(~m[543]&~m[1004]&~m[1005]&m[1006]&m[1007])|(m[543]&~m[1004]&~m[1005]&m[1006]&m[1007])|(~m[543]&m[1004]&~m[1005]&m[1006]&m[1007])|(m[543]&m[1004]&~m[1005]&m[1006]&m[1007])|(~m[543]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[543]&~m[1004]&m[1005]&m[1006]&m[1007])|(m[543]&m[1004]&m[1005]&m[1006]&m[1007]));
    m[1008] = (((m[1006]&~m[1009]&~m[1010]&~m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&~m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&~m[1012])|(~m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&m[1009]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[84])|((m[1006]&~m[1009]&~m[1010]&m[1011]&~m[1012])|(~m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&~m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&~m[1011]&m[1012])|(~m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&~m[1010]&m[1011]&m[1012])|(~m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&~m[1009]&m[1010]&m[1011]&m[1012])|(m[1006]&m[1009]&m[1010]&m[1011]&m[1012]));
    m[1013] = (((m[1011]&~m[1014]&~m[1015]&~m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&~m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&~m[1017])|(~m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&m[1014]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[85])|((m[1011]&~m[1014]&~m[1015]&m[1016]&~m[1017])|(~m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&~m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&~m[1016]&m[1017])|(~m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&~m[1015]&m[1016]&m[1017])|(~m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&~m[1014]&m[1015]&m[1016]&m[1017])|(m[1011]&m[1014]&m[1015]&m[1016]&m[1017]));
    m[1018] = (((m[1016]&~m[1019]&~m[1020]&~m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&~m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&~m[1022])|(~m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&m[1019]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[86])|((m[1016]&~m[1019]&~m[1020]&m[1021]&~m[1022])|(~m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&~m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&~m[1021]&m[1022])|(~m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&~m[1020]&m[1021]&m[1022])|(~m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&~m[1019]&m[1020]&m[1021]&m[1022])|(m[1016]&m[1019]&m[1020]&m[1021]&m[1022]));
    m[1023] = (((m[1021]&~m[1024]&~m[1025]&~m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&~m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&~m[1027])|(~m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&m[1024]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[87])|((m[1021]&~m[1024]&~m[1025]&m[1026]&~m[1027])|(~m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&~m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&~m[1026]&m[1027])|(~m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&~m[1025]&m[1026]&m[1027])|(~m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&~m[1024]&m[1025]&m[1026]&m[1027])|(m[1021]&m[1024]&m[1025]&m[1026]&m[1027]));
    m[1028] = (((m[1026]&~m[1029]&~m[1030]&~m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&~m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&~m[1032])|(~m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&m[1029]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[88])|((m[1026]&~m[1029]&~m[1030]&m[1031]&~m[1032])|(~m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&~m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&~m[1031]&m[1032])|(~m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&~m[1030]&m[1031]&m[1032])|(~m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&~m[1029]&m[1030]&m[1031]&m[1032])|(m[1026]&m[1029]&m[1030]&m[1031]&m[1032]));
    m[1033] = (((m[1031]&~m[1034]&~m[1035]&~m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&~m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&~m[1037])|(~m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&m[1034]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[89])|((m[1031]&~m[1034]&~m[1035]&m[1036]&~m[1037])|(~m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&~m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&~m[1036]&m[1037])|(~m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&~m[1035]&m[1036]&m[1037])|(~m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&~m[1034]&m[1035]&m[1036]&m[1037])|(m[1031]&m[1034]&m[1035]&m[1036]&m[1037]));
    m[1038] = (((m[1036]&~m[1039]&~m[1040]&~m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&~m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&~m[1042])|(~m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&m[1039]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[90])|((m[1036]&~m[1039]&~m[1040]&m[1041]&~m[1042])|(~m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&~m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&~m[1041]&m[1042])|(~m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&~m[1040]&m[1041]&m[1042])|(~m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&~m[1039]&m[1040]&m[1041]&m[1042])|(m[1036]&m[1039]&m[1040]&m[1041]&m[1042]));
    m[1043] = (((m[1041]&~m[1044]&~m[1045]&~m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&~m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&~m[1047])|(~m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&m[1044]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[91])|((m[1041]&~m[1044]&~m[1045]&m[1046]&~m[1047])|(~m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&~m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&~m[1046]&m[1047])|(~m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&~m[1045]&m[1046]&m[1047])|(~m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&~m[1044]&m[1045]&m[1046]&m[1047])|(m[1041]&m[1044]&m[1045]&m[1046]&m[1047]));
    m[1048] = (((m[1046]&~m[1049]&~m[1050]&~m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&~m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&~m[1052])|(~m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&m[1049]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[92])|((m[1046]&~m[1049]&~m[1050]&m[1051]&~m[1052])|(~m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&~m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&~m[1051]&m[1052])|(~m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&~m[1050]&m[1051]&m[1052])|(~m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&~m[1049]&m[1050]&m[1051]&m[1052])|(m[1046]&m[1049]&m[1050]&m[1051]&m[1052]));
    m[1053] = (((m[1051]&~m[1054]&~m[1055]&~m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&~m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&~m[1057])|(~m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&m[1054]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[93])|((m[1051]&~m[1054]&~m[1055]&m[1056]&~m[1057])|(~m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&~m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&~m[1056]&m[1057])|(~m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&~m[1055]&m[1056]&m[1057])|(~m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&~m[1054]&m[1055]&m[1056]&m[1057])|(m[1051]&m[1054]&m[1055]&m[1056]&m[1057]));
    m[1058] = (((m[544]&~m[1059]&~m[1060]&~m[1061]&~m[1062])|(~m[544]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(m[544]&m[1059]&~m[1060]&m[1061]&~m[1062])|(m[544]&~m[1059]&m[1060]&m[1061]&~m[1062])|(~m[544]&m[1059]&~m[1060]&~m[1061]&m[1062])|(~m[544]&~m[1059]&m[1060]&~m[1061]&m[1062])|(m[544]&m[1059]&m[1060]&~m[1061]&m[1062])|(~m[544]&m[1059]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[94])|((m[544]&~m[1059]&~m[1060]&m[1061]&~m[1062])|(~m[544]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[544]&~m[1059]&~m[1060]&~m[1061]&m[1062])|(m[544]&m[1059]&~m[1060]&~m[1061]&m[1062])|(m[544]&~m[1059]&m[1060]&~m[1061]&m[1062])|(~m[544]&~m[1059]&~m[1060]&m[1061]&m[1062])|(m[544]&~m[1059]&~m[1060]&m[1061]&m[1062])|(~m[544]&m[1059]&~m[1060]&m[1061]&m[1062])|(m[544]&m[1059]&~m[1060]&m[1061]&m[1062])|(~m[544]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[544]&~m[1059]&m[1060]&m[1061]&m[1062])|(m[544]&m[1059]&m[1060]&m[1061]&m[1062]));
    m[1063] = (((m[1061]&~m[1064]&~m[1065]&~m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&~m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&~m[1067])|(~m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&m[1064]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[95])|((m[1061]&~m[1064]&~m[1065]&m[1066]&~m[1067])|(~m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&~m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&~m[1066]&m[1067])|(~m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&~m[1065]&m[1066]&m[1067])|(~m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&~m[1064]&m[1065]&m[1066]&m[1067])|(m[1061]&m[1064]&m[1065]&m[1066]&m[1067]));
    m[1068] = (((m[1066]&~m[1069]&~m[1070]&~m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&~m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&~m[1072])|(~m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&m[1069]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[96])|((m[1066]&~m[1069]&~m[1070]&m[1071]&~m[1072])|(~m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&~m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&~m[1071]&m[1072])|(~m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&~m[1070]&m[1071]&m[1072])|(~m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&~m[1069]&m[1070]&m[1071]&m[1072])|(m[1066]&m[1069]&m[1070]&m[1071]&m[1072]));
    m[1073] = (((m[1071]&~m[1074]&~m[1075]&~m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&~m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&~m[1077])|(~m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&m[1074]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[97])|((m[1071]&~m[1074]&~m[1075]&m[1076]&~m[1077])|(~m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&~m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&~m[1076]&m[1077])|(~m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&~m[1075]&m[1076]&m[1077])|(~m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&~m[1074]&m[1075]&m[1076]&m[1077])|(m[1071]&m[1074]&m[1075]&m[1076]&m[1077]));
    m[1078] = (((m[1076]&~m[1079]&~m[1080]&~m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&~m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&~m[1082])|(~m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&m[1079]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[98])|((m[1076]&~m[1079]&~m[1080]&m[1081]&~m[1082])|(~m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&~m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&~m[1081]&m[1082])|(~m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&~m[1080]&m[1081]&m[1082])|(~m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&~m[1079]&m[1080]&m[1081]&m[1082])|(m[1076]&m[1079]&m[1080]&m[1081]&m[1082]));
    m[1083] = (((m[1081]&~m[1084]&~m[1085]&~m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&~m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&~m[1087])|(~m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&m[1084]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[99])|((m[1081]&~m[1084]&~m[1085]&m[1086]&~m[1087])|(~m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&~m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&~m[1086]&m[1087])|(~m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&~m[1085]&m[1086]&m[1087])|(~m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&~m[1084]&m[1085]&m[1086]&m[1087])|(m[1081]&m[1084]&m[1085]&m[1086]&m[1087]));
    m[1088] = (((m[1086]&~m[1089]&~m[1090]&~m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&~m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&~m[1092])|(~m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&m[1089]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[100])|((m[1086]&~m[1089]&~m[1090]&m[1091]&~m[1092])|(~m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&~m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&~m[1091]&m[1092])|(~m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&~m[1090]&m[1091]&m[1092])|(~m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&~m[1089]&m[1090]&m[1091]&m[1092])|(m[1086]&m[1089]&m[1090]&m[1091]&m[1092]));
    m[1093] = (((m[1091]&~m[1094]&~m[1095]&~m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&~m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&~m[1097])|(~m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&m[1094]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[101])|((m[1091]&~m[1094]&~m[1095]&m[1096]&~m[1097])|(~m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&~m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&~m[1096]&m[1097])|(~m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&~m[1095]&m[1096]&m[1097])|(~m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&~m[1094]&m[1095]&m[1096]&m[1097])|(m[1091]&m[1094]&m[1095]&m[1096]&m[1097]));
    m[1098] = (((m[1096]&~m[1099]&~m[1100]&~m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&~m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&~m[1102])|(~m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&m[1099]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[102])|((m[1096]&~m[1099]&~m[1100]&m[1101]&~m[1102])|(~m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&~m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&~m[1101]&m[1102])|(~m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&~m[1100]&m[1101]&m[1102])|(~m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&~m[1099]&m[1100]&m[1101]&m[1102])|(m[1096]&m[1099]&m[1100]&m[1101]&m[1102]));
    m[1103] = (((m[1101]&~m[1104]&~m[1105]&~m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&~m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&~m[1107])|(~m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&m[1104]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[103])|((m[1101]&~m[1104]&~m[1105]&m[1106]&~m[1107])|(~m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&~m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&~m[1106]&m[1107])|(~m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&~m[1105]&m[1106]&m[1107])|(~m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&~m[1104]&m[1105]&m[1106]&m[1107])|(m[1101]&m[1104]&m[1105]&m[1106]&m[1107]));
    m[1108] = (((m[1106]&~m[1109]&~m[1110]&~m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&~m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&~m[1112])|(~m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&m[1109]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[104])|((m[1106]&~m[1109]&~m[1110]&m[1111]&~m[1112])|(~m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&~m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&~m[1111]&m[1112])|(~m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&~m[1110]&m[1111]&m[1112])|(~m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&~m[1109]&m[1110]&m[1111]&m[1112])|(m[1106]&m[1109]&m[1110]&m[1111]&m[1112]));
    m[1113] = (((m[1111]&~m[1114]&~m[1115]&~m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&~m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&~m[1117])|(~m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&m[1114]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[105])|((m[1111]&~m[1114]&~m[1115]&m[1116]&~m[1117])|(~m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&~m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&~m[1116]&m[1117])|(~m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&~m[1115]&m[1116]&m[1117])|(~m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&~m[1114]&m[1115]&m[1116]&m[1117])|(m[1111]&m[1114]&m[1115]&m[1116]&m[1117]));
    m[1118] = (((m[545]&~m[1119]&~m[1120]&~m[1121]&~m[1122])|(~m[545]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(m[545]&m[1119]&~m[1120]&m[1121]&~m[1122])|(m[545]&~m[1119]&m[1120]&m[1121]&~m[1122])|(~m[545]&m[1119]&~m[1120]&~m[1121]&m[1122])|(~m[545]&~m[1119]&m[1120]&~m[1121]&m[1122])|(m[545]&m[1119]&m[1120]&~m[1121]&m[1122])|(~m[545]&m[1119]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[106])|((m[545]&~m[1119]&~m[1120]&m[1121]&~m[1122])|(~m[545]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[545]&~m[1119]&~m[1120]&~m[1121]&m[1122])|(m[545]&m[1119]&~m[1120]&~m[1121]&m[1122])|(m[545]&~m[1119]&m[1120]&~m[1121]&m[1122])|(~m[545]&~m[1119]&~m[1120]&m[1121]&m[1122])|(m[545]&~m[1119]&~m[1120]&m[1121]&m[1122])|(~m[545]&m[1119]&~m[1120]&m[1121]&m[1122])|(m[545]&m[1119]&~m[1120]&m[1121]&m[1122])|(~m[545]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[545]&~m[1119]&m[1120]&m[1121]&m[1122])|(m[545]&m[1119]&m[1120]&m[1121]&m[1122]));
    m[1123] = (((m[1121]&~m[1124]&~m[1125]&~m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&~m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&~m[1127])|(~m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&m[1124]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[107])|((m[1121]&~m[1124]&~m[1125]&m[1126]&~m[1127])|(~m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&~m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&~m[1126]&m[1127])|(~m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&~m[1125]&m[1126]&m[1127])|(~m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&~m[1124]&m[1125]&m[1126]&m[1127])|(m[1121]&m[1124]&m[1125]&m[1126]&m[1127]));
    m[1128] = (((m[1126]&~m[1129]&~m[1130]&~m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&~m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&~m[1132])|(~m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&m[1129]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[108])|((m[1126]&~m[1129]&~m[1130]&m[1131]&~m[1132])|(~m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&~m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&~m[1131]&m[1132])|(~m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&~m[1130]&m[1131]&m[1132])|(~m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&~m[1129]&m[1130]&m[1131]&m[1132])|(m[1126]&m[1129]&m[1130]&m[1131]&m[1132]));
    m[1133] = (((m[1131]&~m[1134]&~m[1135]&~m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&~m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&~m[1137])|(~m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&m[1134]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[109])|((m[1131]&~m[1134]&~m[1135]&m[1136]&~m[1137])|(~m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&~m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&~m[1136]&m[1137])|(~m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&~m[1135]&m[1136]&m[1137])|(~m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&~m[1134]&m[1135]&m[1136]&m[1137])|(m[1131]&m[1134]&m[1135]&m[1136]&m[1137]));
    m[1138] = (((m[1136]&~m[1139]&~m[1140]&~m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&~m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&~m[1142])|(~m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&m[1139]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[110])|((m[1136]&~m[1139]&~m[1140]&m[1141]&~m[1142])|(~m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&~m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&~m[1141]&m[1142])|(~m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&~m[1140]&m[1141]&m[1142])|(~m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&~m[1139]&m[1140]&m[1141]&m[1142])|(m[1136]&m[1139]&m[1140]&m[1141]&m[1142]));
    m[1143] = (((m[1141]&~m[1144]&~m[1145]&~m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&~m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&~m[1147])|(~m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&m[1144]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[111])|((m[1141]&~m[1144]&~m[1145]&m[1146]&~m[1147])|(~m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&~m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&~m[1146]&m[1147])|(~m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&~m[1145]&m[1146]&m[1147])|(~m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&~m[1144]&m[1145]&m[1146]&m[1147])|(m[1141]&m[1144]&m[1145]&m[1146]&m[1147]));
    m[1148] = (((m[1146]&~m[1149]&~m[1150]&~m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&~m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&~m[1152])|(~m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&m[1149]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[112])|((m[1146]&~m[1149]&~m[1150]&m[1151]&~m[1152])|(~m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&~m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&~m[1151]&m[1152])|(~m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&~m[1150]&m[1151]&m[1152])|(~m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&~m[1149]&m[1150]&m[1151]&m[1152])|(m[1146]&m[1149]&m[1150]&m[1151]&m[1152]));
    m[1153] = (((m[1151]&~m[1154]&~m[1155]&~m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&~m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&~m[1157])|(~m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&m[1154]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[113])|((m[1151]&~m[1154]&~m[1155]&m[1156]&~m[1157])|(~m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&~m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&~m[1156]&m[1157])|(~m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&~m[1155]&m[1156]&m[1157])|(~m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&~m[1154]&m[1155]&m[1156]&m[1157])|(m[1151]&m[1154]&m[1155]&m[1156]&m[1157]));
    m[1158] = (((m[1156]&~m[1159]&~m[1160]&~m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&~m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&~m[1162])|(~m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&m[1159]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[114])|((m[1156]&~m[1159]&~m[1160]&m[1161]&~m[1162])|(~m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&~m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&~m[1161]&m[1162])|(~m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&~m[1160]&m[1161]&m[1162])|(~m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&~m[1159]&m[1160]&m[1161]&m[1162])|(m[1156]&m[1159]&m[1160]&m[1161]&m[1162]));
    m[1163] = (((m[1161]&~m[1164]&~m[1165]&~m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&~m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&~m[1167])|(~m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&m[1164]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[115])|((m[1161]&~m[1164]&~m[1165]&m[1166]&~m[1167])|(~m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&~m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&~m[1166]&m[1167])|(~m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&~m[1165]&m[1166]&m[1167])|(~m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&~m[1164]&m[1165]&m[1166]&m[1167])|(m[1161]&m[1164]&m[1165]&m[1166]&m[1167]));
    m[1168] = (((m[1166]&~m[1169]&~m[1170]&~m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&~m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&~m[1172])|(~m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&m[1169]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[116])|((m[1166]&~m[1169]&~m[1170]&m[1171]&~m[1172])|(~m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&~m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&~m[1171]&m[1172])|(~m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&~m[1170]&m[1171]&m[1172])|(~m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&~m[1169]&m[1170]&m[1171]&m[1172])|(m[1166]&m[1169]&m[1170]&m[1171]&m[1172]));
    m[1173] = (((m[1171]&~m[1174]&~m[1175]&~m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&~m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&~m[1177])|(~m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&m[1174]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[117])|((m[1171]&~m[1174]&~m[1175]&m[1176]&~m[1177])|(~m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&~m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&~m[1176]&m[1177])|(~m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&~m[1175]&m[1176]&m[1177])|(~m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&~m[1174]&m[1175]&m[1176]&m[1177])|(m[1171]&m[1174]&m[1175]&m[1176]&m[1177]));
    m[1178] = (((m[1176]&~m[1179]&~m[1180]&~m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&~m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&~m[1182])|(~m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&m[1179]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[118])|((m[1176]&~m[1179]&~m[1180]&m[1181]&~m[1182])|(~m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&~m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&~m[1181]&m[1182])|(~m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&~m[1180]&m[1181]&m[1182])|(~m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&~m[1179]&m[1180]&m[1181]&m[1182])|(m[1176]&m[1179]&m[1180]&m[1181]&m[1182]));
    m[1188] = (((m[1186]&~m[1189]&~m[1190]&~m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&~m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&~m[1192])|(~m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&m[1189]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[119])|((m[1186]&~m[1189]&~m[1190]&m[1191]&~m[1192])|(~m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&~m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&~m[1191]&m[1192])|(~m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&~m[1190]&m[1191]&m[1192])|(~m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&~m[1189]&m[1190]&m[1191]&m[1192])|(m[1186]&m[1189]&m[1190]&m[1191]&m[1192]));
    m[1193] = (((m[1191]&~m[1194]&~m[1195]&~m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&~m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&~m[1197])|(~m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&m[1194]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[120])|((m[1191]&~m[1194]&~m[1195]&m[1196]&~m[1197])|(~m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&~m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&~m[1196]&m[1197])|(~m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&~m[1195]&m[1196]&m[1197])|(~m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&~m[1194]&m[1195]&m[1196]&m[1197])|(m[1191]&m[1194]&m[1195]&m[1196]&m[1197]));
    m[1198] = (((m[1196]&~m[1199]&~m[1200]&~m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&~m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&~m[1202])|(~m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&m[1199]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[121])|((m[1196]&~m[1199]&~m[1200]&m[1201]&~m[1202])|(~m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&~m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&~m[1201]&m[1202])|(~m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&~m[1200]&m[1201]&m[1202])|(~m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&~m[1199]&m[1200]&m[1201]&m[1202])|(m[1196]&m[1199]&m[1200]&m[1201]&m[1202]));
    m[1203] = (((m[1201]&~m[1204]&~m[1205]&~m[1206]&~m[1207])|(~m[1201]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(m[1201]&m[1204]&~m[1205]&m[1206]&~m[1207])|(m[1201]&~m[1204]&m[1205]&m[1206]&~m[1207])|(~m[1201]&m[1204]&~m[1205]&~m[1206]&m[1207])|(~m[1201]&~m[1204]&m[1205]&~m[1206]&m[1207])|(m[1201]&m[1204]&m[1205]&~m[1206]&m[1207])|(~m[1201]&m[1204]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[122])|((m[1201]&~m[1204]&~m[1205]&m[1206]&~m[1207])|(~m[1201]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[1201]&~m[1204]&~m[1205]&~m[1206]&m[1207])|(m[1201]&m[1204]&~m[1205]&~m[1206]&m[1207])|(m[1201]&~m[1204]&m[1205]&~m[1206]&m[1207])|(~m[1201]&~m[1204]&~m[1205]&m[1206]&m[1207])|(m[1201]&~m[1204]&~m[1205]&m[1206]&m[1207])|(~m[1201]&m[1204]&~m[1205]&m[1206]&m[1207])|(m[1201]&m[1204]&~m[1205]&m[1206]&m[1207])|(~m[1201]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[1201]&~m[1204]&m[1205]&m[1206]&m[1207])|(m[1201]&m[1204]&m[1205]&m[1206]&m[1207]));
    m[1208] = (((m[1206]&~m[1209]&~m[1210]&~m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&~m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&~m[1212])|(~m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&m[1209]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[123])|((m[1206]&~m[1209]&~m[1210]&m[1211]&~m[1212])|(~m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&~m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&~m[1211]&m[1212])|(~m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&~m[1210]&m[1211]&m[1212])|(~m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&~m[1209]&m[1210]&m[1211]&m[1212])|(m[1206]&m[1209]&m[1210]&m[1211]&m[1212]));
    m[1213] = (((m[1211]&~m[1214]&~m[1215]&~m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&~m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&~m[1217])|(~m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&m[1214]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[124])|((m[1211]&~m[1214]&~m[1215]&m[1216]&~m[1217])|(~m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&~m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&~m[1216]&m[1217])|(~m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&~m[1215]&m[1216]&m[1217])|(~m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&~m[1214]&m[1215]&m[1216]&m[1217])|(m[1211]&m[1214]&m[1215]&m[1216]&m[1217]));
    m[1218] = (((m[1216]&~m[1219]&~m[1220]&~m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&~m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&~m[1222])|(~m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&m[1219]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[125])|((m[1216]&~m[1219]&~m[1220]&m[1221]&~m[1222])|(~m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&~m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&~m[1221]&m[1222])|(~m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&~m[1220]&m[1221]&m[1222])|(~m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&~m[1219]&m[1220]&m[1221]&m[1222])|(m[1216]&m[1219]&m[1220]&m[1221]&m[1222]));
    m[1223] = (((m[1221]&~m[1224]&~m[1225]&~m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&~m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&~m[1227])|(~m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&m[1224]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[126])|((m[1221]&~m[1224]&~m[1225]&m[1226]&~m[1227])|(~m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&~m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&~m[1226]&m[1227])|(~m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&~m[1225]&m[1226]&m[1227])|(~m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&~m[1224]&m[1225]&m[1226]&m[1227])|(m[1221]&m[1224]&m[1225]&m[1226]&m[1227]));
    m[1228] = (((m[1226]&~m[1229]&~m[1230]&~m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&~m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&~m[1232])|(~m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&m[1229]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[127])|((m[1226]&~m[1229]&~m[1230]&m[1231]&~m[1232])|(~m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&~m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&~m[1231]&m[1232])|(~m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&~m[1230]&m[1231]&m[1232])|(~m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&~m[1229]&m[1230]&m[1231]&m[1232])|(m[1226]&m[1229]&m[1230]&m[1231]&m[1232]));
    m[1233] = (((m[1231]&~m[1234]&~m[1235]&~m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&~m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&~m[1237])|(~m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&m[1234]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[128])|((m[1231]&~m[1234]&~m[1235]&m[1236]&~m[1237])|(~m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&~m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&~m[1236]&m[1237])|(~m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&~m[1235]&m[1236]&m[1237])|(~m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&~m[1234]&m[1235]&m[1236]&m[1237])|(m[1231]&m[1234]&m[1235]&m[1236]&m[1237]));
    m[1238] = (((m[1236]&~m[1239]&~m[1240]&~m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&~m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&~m[1242])|(~m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&m[1239]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[129])|((m[1236]&~m[1239]&~m[1240]&m[1241]&~m[1242])|(~m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&~m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&~m[1241]&m[1242])|(~m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&~m[1240]&m[1241]&m[1242])|(~m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&~m[1239]&m[1240]&m[1241]&m[1242])|(m[1236]&m[1239]&m[1240]&m[1241]&m[1242]));
    m[1243] = (((m[1241]&~m[1244]&~m[1245]&~m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&~m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&~m[1247])|(~m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&m[1244]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[130])|((m[1241]&~m[1244]&~m[1245]&m[1246]&~m[1247])|(~m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&~m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&~m[1246]&m[1247])|(~m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&~m[1245]&m[1246]&m[1247])|(~m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&~m[1244]&m[1245]&m[1246]&m[1247])|(m[1241]&m[1244]&m[1245]&m[1246]&m[1247]));
    m[1248] = (((m[1187]&~m[1249]&~m[1250]&~m[1251]&~m[1252])|(~m[1187]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1187]&m[1249]&~m[1250]&m[1251]&~m[1252])|(m[1187]&~m[1249]&m[1250]&m[1251]&~m[1252])|(~m[1187]&m[1249]&~m[1250]&~m[1251]&m[1252])|(~m[1187]&~m[1249]&m[1250]&~m[1251]&m[1252])|(m[1187]&m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1187]&m[1249]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[131])|((m[1187]&~m[1249]&~m[1250]&m[1251]&~m[1252])|(~m[1187]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1187]&~m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1187]&m[1249]&~m[1250]&~m[1251]&m[1252])|(m[1187]&~m[1249]&m[1250]&~m[1251]&m[1252])|(~m[1187]&~m[1249]&~m[1250]&m[1251]&m[1252])|(m[1187]&~m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1187]&m[1249]&~m[1250]&m[1251]&m[1252])|(m[1187]&m[1249]&~m[1250]&m[1251]&m[1252])|(~m[1187]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1187]&~m[1249]&m[1250]&m[1251]&m[1252])|(m[1187]&m[1249]&m[1250]&m[1251]&m[1252]));
    m[1253] = (((m[1251]&~m[1254]&~m[1255]&~m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&~m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&~m[1257])|(~m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&m[1254]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[132])|((m[1251]&~m[1254]&~m[1255]&m[1256]&~m[1257])|(~m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&~m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&~m[1256]&m[1257])|(~m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&~m[1255]&m[1256]&m[1257])|(~m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&~m[1254]&m[1255]&m[1256]&m[1257])|(m[1251]&m[1254]&m[1255]&m[1256]&m[1257]));
    m[1258] = (((m[1256]&~m[1259]&~m[1260]&~m[1261]&~m[1262])|(~m[1256]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(m[1256]&m[1259]&~m[1260]&m[1261]&~m[1262])|(m[1256]&~m[1259]&m[1260]&m[1261]&~m[1262])|(~m[1256]&m[1259]&~m[1260]&~m[1261]&m[1262])|(~m[1256]&~m[1259]&m[1260]&~m[1261]&m[1262])|(m[1256]&m[1259]&m[1260]&~m[1261]&m[1262])|(~m[1256]&m[1259]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[133])|((m[1256]&~m[1259]&~m[1260]&m[1261]&~m[1262])|(~m[1256]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[1256]&~m[1259]&~m[1260]&~m[1261]&m[1262])|(m[1256]&m[1259]&~m[1260]&~m[1261]&m[1262])|(m[1256]&~m[1259]&m[1260]&~m[1261]&m[1262])|(~m[1256]&~m[1259]&~m[1260]&m[1261]&m[1262])|(m[1256]&~m[1259]&~m[1260]&m[1261]&m[1262])|(~m[1256]&m[1259]&~m[1260]&m[1261]&m[1262])|(m[1256]&m[1259]&~m[1260]&m[1261]&m[1262])|(~m[1256]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[1256]&~m[1259]&m[1260]&m[1261]&m[1262])|(m[1256]&m[1259]&m[1260]&m[1261]&m[1262]));
    m[1263] = (((m[1261]&~m[1264]&~m[1265]&~m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&~m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&~m[1267])|(~m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&m[1264]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[134])|((m[1261]&~m[1264]&~m[1265]&m[1266]&~m[1267])|(~m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&~m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&~m[1266]&m[1267])|(~m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&~m[1265]&m[1266]&m[1267])|(~m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&~m[1264]&m[1265]&m[1266]&m[1267])|(m[1261]&m[1264]&m[1265]&m[1266]&m[1267]));
    m[1268] = (((m[1266]&~m[1269]&~m[1270]&~m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&~m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&~m[1272])|(~m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&m[1269]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[135])|((m[1266]&~m[1269]&~m[1270]&m[1271]&~m[1272])|(~m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&~m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&~m[1271]&m[1272])|(~m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&~m[1270]&m[1271]&m[1272])|(~m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&~m[1269]&m[1270]&m[1271]&m[1272])|(m[1266]&m[1269]&m[1270]&m[1271]&m[1272]));
    m[1273] = (((m[1271]&~m[1274]&~m[1275]&~m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&~m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&~m[1277])|(~m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&m[1274]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[136])|((m[1271]&~m[1274]&~m[1275]&m[1276]&~m[1277])|(~m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&~m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&~m[1276]&m[1277])|(~m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&~m[1275]&m[1276]&m[1277])|(~m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&~m[1274]&m[1275]&m[1276]&m[1277])|(m[1271]&m[1274]&m[1275]&m[1276]&m[1277]));
    m[1278] = (((m[1276]&~m[1279]&~m[1280]&~m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&~m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&~m[1282])|(~m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&m[1279]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[137])|((m[1276]&~m[1279]&~m[1280]&m[1281]&~m[1282])|(~m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&~m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&~m[1281]&m[1282])|(~m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&~m[1280]&m[1281]&m[1282])|(~m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&~m[1279]&m[1280]&m[1281]&m[1282])|(m[1276]&m[1279]&m[1280]&m[1281]&m[1282]));
    m[1283] = (((m[1281]&~m[1284]&~m[1285]&~m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&~m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&~m[1287])|(~m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&m[1284]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[138])|((m[1281]&~m[1284]&~m[1285]&m[1286]&~m[1287])|(~m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&~m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&~m[1286]&m[1287])|(~m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&~m[1285]&m[1286]&m[1287])|(~m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&~m[1284]&m[1285]&m[1286]&m[1287])|(m[1281]&m[1284]&m[1285]&m[1286]&m[1287]));
    m[1288] = (((m[1286]&~m[1289]&~m[1290]&~m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&~m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&~m[1292])|(~m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&m[1289]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[139])|((m[1286]&~m[1289]&~m[1290]&m[1291]&~m[1292])|(~m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&~m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&~m[1291]&m[1292])|(~m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&~m[1290]&m[1291]&m[1292])|(~m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&~m[1289]&m[1290]&m[1291]&m[1292])|(m[1286]&m[1289]&m[1290]&m[1291]&m[1292]));
    m[1293] = (((m[1291]&~m[1294]&~m[1295]&~m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&~m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&~m[1297])|(~m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&m[1294]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[140])|((m[1291]&~m[1294]&~m[1295]&m[1296]&~m[1297])|(~m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&~m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&~m[1296]&m[1297])|(~m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&~m[1295]&m[1296]&m[1297])|(~m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&~m[1294]&m[1295]&m[1296]&m[1297])|(m[1291]&m[1294]&m[1295]&m[1296]&m[1297]));
    m[1298] = (((m[1296]&~m[1299]&~m[1300]&~m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&~m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&~m[1302])|(~m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&m[1299]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[141])|((m[1296]&~m[1299]&~m[1300]&m[1301]&~m[1302])|(~m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&~m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&~m[1301]&m[1302])|(~m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&~m[1300]&m[1301]&m[1302])|(~m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&~m[1299]&m[1300]&m[1301]&m[1302])|(m[1296]&m[1299]&m[1300]&m[1301]&m[1302]));
    m[1303] = (((m[1301]&~m[1304]&~m[1305]&~m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&~m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&~m[1307])|(~m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&m[1304]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[142])|((m[1301]&~m[1304]&~m[1305]&m[1306]&~m[1307])|(~m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&~m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&~m[1306]&m[1307])|(~m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&~m[1305]&m[1306]&m[1307])|(~m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&~m[1304]&m[1305]&m[1306]&m[1307])|(m[1301]&m[1304]&m[1305]&m[1306]&m[1307]));
    m[1308] = (((m[1252]&~m[1309]&~m[1310]&~m[1311]&~m[1312])|(~m[1252]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1252]&m[1309]&~m[1310]&m[1311]&~m[1312])|(m[1252]&~m[1309]&m[1310]&m[1311]&~m[1312])|(~m[1252]&m[1309]&~m[1310]&~m[1311]&m[1312])|(~m[1252]&~m[1309]&m[1310]&~m[1311]&m[1312])|(m[1252]&m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1252]&m[1309]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[143])|((m[1252]&~m[1309]&~m[1310]&m[1311]&~m[1312])|(~m[1252]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1252]&~m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1252]&m[1309]&~m[1310]&~m[1311]&m[1312])|(m[1252]&~m[1309]&m[1310]&~m[1311]&m[1312])|(~m[1252]&~m[1309]&~m[1310]&m[1311]&m[1312])|(m[1252]&~m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1252]&m[1309]&~m[1310]&m[1311]&m[1312])|(m[1252]&m[1309]&~m[1310]&m[1311]&m[1312])|(~m[1252]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1252]&~m[1309]&m[1310]&m[1311]&m[1312])|(m[1252]&m[1309]&m[1310]&m[1311]&m[1312]));
    m[1313] = (((m[1311]&~m[1314]&~m[1315]&~m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&~m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&~m[1317])|(~m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&m[1314]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[144])|((m[1311]&~m[1314]&~m[1315]&m[1316]&~m[1317])|(~m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&~m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&~m[1316]&m[1317])|(~m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&~m[1315]&m[1316]&m[1317])|(~m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&~m[1314]&m[1315]&m[1316]&m[1317])|(m[1311]&m[1314]&m[1315]&m[1316]&m[1317]));
    m[1318] = (((m[1316]&~m[1319]&~m[1320]&~m[1321]&~m[1322])|(~m[1316]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(m[1316]&m[1319]&~m[1320]&m[1321]&~m[1322])|(m[1316]&~m[1319]&m[1320]&m[1321]&~m[1322])|(~m[1316]&m[1319]&~m[1320]&~m[1321]&m[1322])|(~m[1316]&~m[1319]&m[1320]&~m[1321]&m[1322])|(m[1316]&m[1319]&m[1320]&~m[1321]&m[1322])|(~m[1316]&m[1319]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[145])|((m[1316]&~m[1319]&~m[1320]&m[1321]&~m[1322])|(~m[1316]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[1316]&~m[1319]&~m[1320]&~m[1321]&m[1322])|(m[1316]&m[1319]&~m[1320]&~m[1321]&m[1322])|(m[1316]&~m[1319]&m[1320]&~m[1321]&m[1322])|(~m[1316]&~m[1319]&~m[1320]&m[1321]&m[1322])|(m[1316]&~m[1319]&~m[1320]&m[1321]&m[1322])|(~m[1316]&m[1319]&~m[1320]&m[1321]&m[1322])|(m[1316]&m[1319]&~m[1320]&m[1321]&m[1322])|(~m[1316]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[1316]&~m[1319]&m[1320]&m[1321]&m[1322])|(m[1316]&m[1319]&m[1320]&m[1321]&m[1322]));
    m[1323] = (((m[1321]&~m[1324]&~m[1325]&~m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&~m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&~m[1327])|(~m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&m[1324]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[146])|((m[1321]&~m[1324]&~m[1325]&m[1326]&~m[1327])|(~m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&~m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&~m[1326]&m[1327])|(~m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&~m[1325]&m[1326]&m[1327])|(~m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&~m[1324]&m[1325]&m[1326]&m[1327])|(m[1321]&m[1324]&m[1325]&m[1326]&m[1327]));
    m[1328] = (((m[1326]&~m[1329]&~m[1330]&~m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&~m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&~m[1332])|(~m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&m[1329]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[147])|((m[1326]&~m[1329]&~m[1330]&m[1331]&~m[1332])|(~m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&~m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&~m[1331]&m[1332])|(~m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&~m[1330]&m[1331]&m[1332])|(~m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&~m[1329]&m[1330]&m[1331]&m[1332])|(m[1326]&m[1329]&m[1330]&m[1331]&m[1332]));
    m[1333] = (((m[1331]&~m[1334]&~m[1335]&~m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&~m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&~m[1337])|(~m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&m[1334]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[148])|((m[1331]&~m[1334]&~m[1335]&m[1336]&~m[1337])|(~m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&~m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&~m[1336]&m[1337])|(~m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&~m[1335]&m[1336]&m[1337])|(~m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&~m[1334]&m[1335]&m[1336]&m[1337])|(m[1331]&m[1334]&m[1335]&m[1336]&m[1337]));
    m[1338] = (((m[1336]&~m[1339]&~m[1340]&~m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&~m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&~m[1342])|(~m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&m[1339]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[149])|((m[1336]&~m[1339]&~m[1340]&m[1341]&~m[1342])|(~m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&~m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&~m[1341]&m[1342])|(~m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&~m[1340]&m[1341]&m[1342])|(~m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&~m[1339]&m[1340]&m[1341]&m[1342])|(m[1336]&m[1339]&m[1340]&m[1341]&m[1342]));
    m[1343] = (((m[1341]&~m[1344]&~m[1345]&~m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&~m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&~m[1347])|(~m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&m[1344]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[150])|((m[1341]&~m[1344]&~m[1345]&m[1346]&~m[1347])|(~m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&~m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&~m[1346]&m[1347])|(~m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&~m[1345]&m[1346]&m[1347])|(~m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&~m[1344]&m[1345]&m[1346]&m[1347])|(m[1341]&m[1344]&m[1345]&m[1346]&m[1347]));
    m[1348] = (((m[1346]&~m[1349]&~m[1350]&~m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&~m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&~m[1352])|(~m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&m[1349]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[151])|((m[1346]&~m[1349]&~m[1350]&m[1351]&~m[1352])|(~m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&~m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&~m[1351]&m[1352])|(~m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&~m[1350]&m[1351]&m[1352])|(~m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&~m[1349]&m[1350]&m[1351]&m[1352])|(m[1346]&m[1349]&m[1350]&m[1351]&m[1352]));
    m[1353] = (((m[1351]&~m[1354]&~m[1355]&~m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&~m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&~m[1357])|(~m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&m[1354]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[152])|((m[1351]&~m[1354]&~m[1355]&m[1356]&~m[1357])|(~m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&~m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&~m[1356]&m[1357])|(~m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&~m[1355]&m[1356]&m[1357])|(~m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&~m[1354]&m[1355]&m[1356]&m[1357])|(m[1351]&m[1354]&m[1355]&m[1356]&m[1357]));
    m[1358] = (((m[1356]&~m[1359]&~m[1360]&~m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&~m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&~m[1362])|(~m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&m[1359]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[153])|((m[1356]&~m[1359]&~m[1360]&m[1361]&~m[1362])|(~m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&~m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&~m[1361]&m[1362])|(~m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&~m[1360]&m[1361]&m[1362])|(~m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&~m[1359]&m[1360]&m[1361]&m[1362])|(m[1356]&m[1359]&m[1360]&m[1361]&m[1362]));
    m[1363] = (((m[1312]&~m[1364]&~m[1365]&~m[1366]&~m[1367])|(~m[1312]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1312]&m[1364]&~m[1365]&m[1366]&~m[1367])|(m[1312]&~m[1364]&m[1365]&m[1366]&~m[1367])|(~m[1312]&m[1364]&~m[1365]&~m[1366]&m[1367])|(~m[1312]&~m[1364]&m[1365]&~m[1366]&m[1367])|(m[1312]&m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1312]&m[1364]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[154])|((m[1312]&~m[1364]&~m[1365]&m[1366]&~m[1367])|(~m[1312]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1312]&~m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1312]&m[1364]&~m[1365]&~m[1366]&m[1367])|(m[1312]&~m[1364]&m[1365]&~m[1366]&m[1367])|(~m[1312]&~m[1364]&~m[1365]&m[1366]&m[1367])|(m[1312]&~m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1312]&m[1364]&~m[1365]&m[1366]&m[1367])|(m[1312]&m[1364]&~m[1365]&m[1366]&m[1367])|(~m[1312]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1312]&~m[1364]&m[1365]&m[1366]&m[1367])|(m[1312]&m[1364]&m[1365]&m[1366]&m[1367]));
    m[1368] = (((m[1366]&~m[1369]&~m[1370]&~m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&~m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&~m[1372])|(~m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&m[1369]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[155])|((m[1366]&~m[1369]&~m[1370]&m[1371]&~m[1372])|(~m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&~m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&~m[1371]&m[1372])|(~m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&~m[1370]&m[1371]&m[1372])|(~m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&~m[1369]&m[1370]&m[1371]&m[1372])|(m[1366]&m[1369]&m[1370]&m[1371]&m[1372]));
    m[1373] = (((m[1371]&~m[1374]&~m[1375]&~m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&~m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&~m[1377])|(~m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&m[1374]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[156])|((m[1371]&~m[1374]&~m[1375]&m[1376]&~m[1377])|(~m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&~m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&~m[1376]&m[1377])|(~m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&~m[1375]&m[1376]&m[1377])|(~m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&~m[1374]&m[1375]&m[1376]&m[1377])|(m[1371]&m[1374]&m[1375]&m[1376]&m[1377]));
    m[1378] = (((m[1376]&~m[1379]&~m[1380]&~m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&~m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&~m[1382])|(~m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&m[1379]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[157])|((m[1376]&~m[1379]&~m[1380]&m[1381]&~m[1382])|(~m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&~m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&~m[1381]&m[1382])|(~m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&~m[1380]&m[1381]&m[1382])|(~m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&~m[1379]&m[1380]&m[1381]&m[1382])|(m[1376]&m[1379]&m[1380]&m[1381]&m[1382]));
    m[1383] = (((m[1381]&~m[1384]&~m[1385]&~m[1386]&~m[1387])|(~m[1381]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(m[1381]&m[1384]&~m[1385]&m[1386]&~m[1387])|(m[1381]&~m[1384]&m[1385]&m[1386]&~m[1387])|(~m[1381]&m[1384]&~m[1385]&~m[1386]&m[1387])|(~m[1381]&~m[1384]&m[1385]&~m[1386]&m[1387])|(m[1381]&m[1384]&m[1385]&~m[1386]&m[1387])|(~m[1381]&m[1384]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[158])|((m[1381]&~m[1384]&~m[1385]&m[1386]&~m[1387])|(~m[1381]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[1381]&~m[1384]&~m[1385]&~m[1386]&m[1387])|(m[1381]&m[1384]&~m[1385]&~m[1386]&m[1387])|(m[1381]&~m[1384]&m[1385]&~m[1386]&m[1387])|(~m[1381]&~m[1384]&~m[1385]&m[1386]&m[1387])|(m[1381]&~m[1384]&~m[1385]&m[1386]&m[1387])|(~m[1381]&m[1384]&~m[1385]&m[1386]&m[1387])|(m[1381]&m[1384]&~m[1385]&m[1386]&m[1387])|(~m[1381]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[1381]&~m[1384]&m[1385]&m[1386]&m[1387])|(m[1381]&m[1384]&m[1385]&m[1386]&m[1387]));
    m[1388] = (((m[1386]&~m[1389]&~m[1390]&~m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&~m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&~m[1392])|(~m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&m[1389]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[159])|((m[1386]&~m[1389]&~m[1390]&m[1391]&~m[1392])|(~m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&~m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&~m[1391]&m[1392])|(~m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&~m[1390]&m[1391]&m[1392])|(~m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&~m[1389]&m[1390]&m[1391]&m[1392])|(m[1386]&m[1389]&m[1390]&m[1391]&m[1392]));
    m[1393] = (((m[1391]&~m[1394]&~m[1395]&~m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&~m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&~m[1397])|(~m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&m[1394]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[160])|((m[1391]&~m[1394]&~m[1395]&m[1396]&~m[1397])|(~m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&~m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&~m[1396]&m[1397])|(~m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&~m[1395]&m[1396]&m[1397])|(~m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&~m[1394]&m[1395]&m[1396]&m[1397])|(m[1391]&m[1394]&m[1395]&m[1396]&m[1397]));
    m[1398] = (((m[1396]&~m[1399]&~m[1400]&~m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&~m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&~m[1402])|(~m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&m[1399]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[161])|((m[1396]&~m[1399]&~m[1400]&m[1401]&~m[1402])|(~m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&~m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&~m[1401]&m[1402])|(~m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&~m[1400]&m[1401]&m[1402])|(~m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&~m[1399]&m[1400]&m[1401]&m[1402])|(m[1396]&m[1399]&m[1400]&m[1401]&m[1402]));
    m[1403] = (((m[1401]&~m[1404]&~m[1405]&~m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&~m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&~m[1407])|(~m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&m[1404]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[162])|((m[1401]&~m[1404]&~m[1405]&m[1406]&~m[1407])|(~m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&~m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&~m[1406]&m[1407])|(~m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&~m[1405]&m[1406]&m[1407])|(~m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&~m[1404]&m[1405]&m[1406]&m[1407])|(m[1401]&m[1404]&m[1405]&m[1406]&m[1407]));
    m[1408] = (((m[1406]&~m[1409]&~m[1410]&~m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&~m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&~m[1412])|(~m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&m[1409]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[163])|((m[1406]&~m[1409]&~m[1410]&m[1411]&~m[1412])|(~m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&~m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&~m[1411]&m[1412])|(~m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&~m[1410]&m[1411]&m[1412])|(~m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&~m[1409]&m[1410]&m[1411]&m[1412])|(m[1406]&m[1409]&m[1410]&m[1411]&m[1412]));
    m[1413] = (((m[1367]&~m[1414]&~m[1415]&~m[1416]&~m[1417])|(~m[1367]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1367]&m[1414]&~m[1415]&m[1416]&~m[1417])|(m[1367]&~m[1414]&m[1415]&m[1416]&~m[1417])|(~m[1367]&m[1414]&~m[1415]&~m[1416]&m[1417])|(~m[1367]&~m[1414]&m[1415]&~m[1416]&m[1417])|(m[1367]&m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1367]&m[1414]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[164])|((m[1367]&~m[1414]&~m[1415]&m[1416]&~m[1417])|(~m[1367]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1367]&~m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1367]&m[1414]&~m[1415]&~m[1416]&m[1417])|(m[1367]&~m[1414]&m[1415]&~m[1416]&m[1417])|(~m[1367]&~m[1414]&~m[1415]&m[1416]&m[1417])|(m[1367]&~m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1367]&m[1414]&~m[1415]&m[1416]&m[1417])|(m[1367]&m[1414]&~m[1415]&m[1416]&m[1417])|(~m[1367]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1367]&~m[1414]&m[1415]&m[1416]&m[1417])|(m[1367]&m[1414]&m[1415]&m[1416]&m[1417]));
    m[1418] = (((m[1416]&~m[1419]&~m[1420]&~m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&~m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&~m[1422])|(~m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&m[1419]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[165])|((m[1416]&~m[1419]&~m[1420]&m[1421]&~m[1422])|(~m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&~m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&~m[1421]&m[1422])|(~m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&~m[1420]&m[1421]&m[1422])|(~m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&~m[1419]&m[1420]&m[1421]&m[1422])|(m[1416]&m[1419]&m[1420]&m[1421]&m[1422]));
    m[1423] = (((m[1421]&~m[1424]&~m[1425]&~m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&~m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&~m[1427])|(~m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&m[1424]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[166])|((m[1421]&~m[1424]&~m[1425]&m[1426]&~m[1427])|(~m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&~m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&~m[1426]&m[1427])|(~m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&~m[1425]&m[1426]&m[1427])|(~m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&~m[1424]&m[1425]&m[1426]&m[1427])|(m[1421]&m[1424]&m[1425]&m[1426]&m[1427]));
    m[1428] = (((m[1426]&~m[1429]&~m[1430]&~m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&~m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&~m[1432])|(~m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&m[1429]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[167])|((m[1426]&~m[1429]&~m[1430]&m[1431]&~m[1432])|(~m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&~m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&~m[1431]&m[1432])|(~m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&~m[1430]&m[1431]&m[1432])|(~m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&~m[1429]&m[1430]&m[1431]&m[1432])|(m[1426]&m[1429]&m[1430]&m[1431]&m[1432]));
    m[1433] = (((m[1431]&~m[1434]&~m[1435]&~m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&~m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&~m[1437])|(~m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&m[1434]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[168])|((m[1431]&~m[1434]&~m[1435]&m[1436]&~m[1437])|(~m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&~m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&~m[1436]&m[1437])|(~m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&~m[1435]&m[1436]&m[1437])|(~m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&~m[1434]&m[1435]&m[1436]&m[1437])|(m[1431]&m[1434]&m[1435]&m[1436]&m[1437]));
    m[1438] = (((m[1436]&~m[1439]&~m[1440]&~m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&~m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&~m[1442])|(~m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&m[1439]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[169])|((m[1436]&~m[1439]&~m[1440]&m[1441]&~m[1442])|(~m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&~m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&~m[1441]&m[1442])|(~m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&~m[1440]&m[1441]&m[1442])|(~m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&~m[1439]&m[1440]&m[1441]&m[1442])|(m[1436]&m[1439]&m[1440]&m[1441]&m[1442]));
    m[1443] = (((m[1441]&~m[1444]&~m[1445]&~m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&~m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&~m[1447])|(~m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&m[1444]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[170])|((m[1441]&~m[1444]&~m[1445]&m[1446]&~m[1447])|(~m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&~m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&~m[1446]&m[1447])|(~m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&~m[1445]&m[1446]&m[1447])|(~m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&~m[1444]&m[1445]&m[1446]&m[1447])|(m[1441]&m[1444]&m[1445]&m[1446]&m[1447]));
    m[1448] = (((m[1446]&~m[1449]&~m[1450]&~m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&~m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&~m[1452])|(~m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&m[1449]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[171])|((m[1446]&~m[1449]&~m[1450]&m[1451]&~m[1452])|(~m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&~m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&~m[1451]&m[1452])|(~m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&~m[1450]&m[1451]&m[1452])|(~m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&~m[1449]&m[1450]&m[1451]&m[1452])|(m[1446]&m[1449]&m[1450]&m[1451]&m[1452]));
    m[1453] = (((m[1451]&~m[1454]&~m[1455]&~m[1456]&~m[1457])|(~m[1451]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(m[1451]&m[1454]&~m[1455]&m[1456]&~m[1457])|(m[1451]&~m[1454]&m[1455]&m[1456]&~m[1457])|(~m[1451]&m[1454]&~m[1455]&~m[1456]&m[1457])|(~m[1451]&~m[1454]&m[1455]&~m[1456]&m[1457])|(m[1451]&m[1454]&m[1455]&~m[1456]&m[1457])|(~m[1451]&m[1454]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[172])|((m[1451]&~m[1454]&~m[1455]&m[1456]&~m[1457])|(~m[1451]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[1451]&~m[1454]&~m[1455]&~m[1456]&m[1457])|(m[1451]&m[1454]&~m[1455]&~m[1456]&m[1457])|(m[1451]&~m[1454]&m[1455]&~m[1456]&m[1457])|(~m[1451]&~m[1454]&~m[1455]&m[1456]&m[1457])|(m[1451]&~m[1454]&~m[1455]&m[1456]&m[1457])|(~m[1451]&m[1454]&~m[1455]&m[1456]&m[1457])|(m[1451]&m[1454]&~m[1455]&m[1456]&m[1457])|(~m[1451]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[1451]&~m[1454]&m[1455]&m[1456]&m[1457])|(m[1451]&m[1454]&m[1455]&m[1456]&m[1457]));
    m[1458] = (((m[1417]&~m[1459]&~m[1460]&~m[1461]&~m[1462])|(~m[1417]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1417]&m[1459]&~m[1460]&m[1461]&~m[1462])|(m[1417]&~m[1459]&m[1460]&m[1461]&~m[1462])|(~m[1417]&m[1459]&~m[1460]&~m[1461]&m[1462])|(~m[1417]&~m[1459]&m[1460]&~m[1461]&m[1462])|(m[1417]&m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1417]&m[1459]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[173])|((m[1417]&~m[1459]&~m[1460]&m[1461]&~m[1462])|(~m[1417]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1417]&~m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1417]&m[1459]&~m[1460]&~m[1461]&m[1462])|(m[1417]&~m[1459]&m[1460]&~m[1461]&m[1462])|(~m[1417]&~m[1459]&~m[1460]&m[1461]&m[1462])|(m[1417]&~m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1417]&m[1459]&~m[1460]&m[1461]&m[1462])|(m[1417]&m[1459]&~m[1460]&m[1461]&m[1462])|(~m[1417]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1417]&~m[1459]&m[1460]&m[1461]&m[1462])|(m[1417]&m[1459]&m[1460]&m[1461]&m[1462]));
    m[1463] = (((m[1461]&~m[1464]&~m[1465]&~m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&~m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&~m[1467])|(~m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&m[1464]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[174])|((m[1461]&~m[1464]&~m[1465]&m[1466]&~m[1467])|(~m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&~m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&~m[1466]&m[1467])|(~m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&~m[1465]&m[1466]&m[1467])|(~m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&~m[1464]&m[1465]&m[1466]&m[1467])|(m[1461]&m[1464]&m[1465]&m[1466]&m[1467]));
    m[1468] = (((m[1466]&~m[1469]&~m[1470]&~m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&~m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&~m[1472])|(~m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&m[1469]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[175])|((m[1466]&~m[1469]&~m[1470]&m[1471]&~m[1472])|(~m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&~m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&~m[1471]&m[1472])|(~m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&~m[1470]&m[1471]&m[1472])|(~m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&~m[1469]&m[1470]&m[1471]&m[1472])|(m[1466]&m[1469]&m[1470]&m[1471]&m[1472]));
    m[1473] = (((m[1471]&~m[1474]&~m[1475]&~m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&~m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&~m[1477])|(~m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&m[1474]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[176])|((m[1471]&~m[1474]&~m[1475]&m[1476]&~m[1477])|(~m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&~m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&~m[1476]&m[1477])|(~m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&~m[1475]&m[1476]&m[1477])|(~m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&~m[1474]&m[1475]&m[1476]&m[1477])|(m[1471]&m[1474]&m[1475]&m[1476]&m[1477]));
    m[1478] = (((m[1476]&~m[1479]&~m[1480]&~m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&~m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&~m[1482])|(~m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&m[1479]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[177])|((m[1476]&~m[1479]&~m[1480]&m[1481]&~m[1482])|(~m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&~m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&~m[1481]&m[1482])|(~m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&~m[1480]&m[1481]&m[1482])|(~m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&~m[1479]&m[1480]&m[1481]&m[1482])|(m[1476]&m[1479]&m[1480]&m[1481]&m[1482]));
    m[1483] = (((m[1481]&~m[1484]&~m[1485]&~m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&~m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&~m[1487])|(~m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&m[1484]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[178])|((m[1481]&~m[1484]&~m[1485]&m[1486]&~m[1487])|(~m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&~m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&~m[1486]&m[1487])|(~m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&~m[1485]&m[1486]&m[1487])|(~m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&~m[1484]&m[1485]&m[1486]&m[1487])|(m[1481]&m[1484]&m[1485]&m[1486]&m[1487]));
    m[1488] = (((m[1486]&~m[1489]&~m[1490]&~m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&~m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&~m[1492])|(~m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&m[1489]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[179])|((m[1486]&~m[1489]&~m[1490]&m[1491]&~m[1492])|(~m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&~m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&~m[1491]&m[1492])|(~m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&~m[1490]&m[1491]&m[1492])|(~m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&~m[1489]&m[1490]&m[1491]&m[1492])|(m[1486]&m[1489]&m[1490]&m[1491]&m[1492]));
    m[1493] = (((m[1491]&~m[1494]&~m[1495]&~m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&~m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&~m[1497])|(~m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&m[1494]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[180])|((m[1491]&~m[1494]&~m[1495]&m[1496]&~m[1497])|(~m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&~m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&~m[1496]&m[1497])|(~m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&~m[1495]&m[1496]&m[1497])|(~m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&~m[1494]&m[1495]&m[1496]&m[1497])|(m[1491]&m[1494]&m[1495]&m[1496]&m[1497]));
    m[1498] = (((m[1462]&~m[1499]&~m[1500]&~m[1501]&~m[1502])|(~m[1462]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1462]&m[1499]&~m[1500]&m[1501]&~m[1502])|(m[1462]&~m[1499]&m[1500]&m[1501]&~m[1502])|(~m[1462]&m[1499]&~m[1500]&~m[1501]&m[1502])|(~m[1462]&~m[1499]&m[1500]&~m[1501]&m[1502])|(m[1462]&m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1462]&m[1499]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[181])|((m[1462]&~m[1499]&~m[1500]&m[1501]&~m[1502])|(~m[1462]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1462]&~m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1462]&m[1499]&~m[1500]&~m[1501]&m[1502])|(m[1462]&~m[1499]&m[1500]&~m[1501]&m[1502])|(~m[1462]&~m[1499]&~m[1500]&m[1501]&m[1502])|(m[1462]&~m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1462]&m[1499]&~m[1500]&m[1501]&m[1502])|(m[1462]&m[1499]&~m[1500]&m[1501]&m[1502])|(~m[1462]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1462]&~m[1499]&m[1500]&m[1501]&m[1502])|(m[1462]&m[1499]&m[1500]&m[1501]&m[1502]));
    m[1503] = (((m[1501]&~m[1504]&~m[1505]&~m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&~m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&~m[1507])|(~m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&m[1504]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[182])|((m[1501]&~m[1504]&~m[1505]&m[1506]&~m[1507])|(~m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&~m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&~m[1506]&m[1507])|(~m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&~m[1505]&m[1506]&m[1507])|(~m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&~m[1504]&m[1505]&m[1506]&m[1507])|(m[1501]&m[1504]&m[1505]&m[1506]&m[1507]));
    m[1508] = (((m[1506]&~m[1509]&~m[1510]&~m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&~m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&~m[1512])|(~m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&m[1509]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[183])|((m[1506]&~m[1509]&~m[1510]&m[1511]&~m[1512])|(~m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&~m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&~m[1511]&m[1512])|(~m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&~m[1510]&m[1511]&m[1512])|(~m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&~m[1509]&m[1510]&m[1511]&m[1512])|(m[1506]&m[1509]&m[1510]&m[1511]&m[1512]));
    m[1513] = (((m[1511]&~m[1514]&~m[1515]&~m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&~m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&~m[1517])|(~m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&m[1514]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[184])|((m[1511]&~m[1514]&~m[1515]&m[1516]&~m[1517])|(~m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&~m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&~m[1516]&m[1517])|(~m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&~m[1515]&m[1516]&m[1517])|(~m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&~m[1514]&m[1515]&m[1516]&m[1517])|(m[1511]&m[1514]&m[1515]&m[1516]&m[1517]));
    m[1518] = (((m[1516]&~m[1519]&~m[1520]&~m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&~m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&~m[1522])|(~m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&m[1519]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[185])|((m[1516]&~m[1519]&~m[1520]&m[1521]&~m[1522])|(~m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&~m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&~m[1521]&m[1522])|(~m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&~m[1520]&m[1521]&m[1522])|(~m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&~m[1519]&m[1520]&m[1521]&m[1522])|(m[1516]&m[1519]&m[1520]&m[1521]&m[1522]));
    m[1523] = (((m[1521]&~m[1524]&~m[1525]&~m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&~m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&~m[1527])|(~m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&m[1524]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[186])|((m[1521]&~m[1524]&~m[1525]&m[1526]&~m[1527])|(~m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&~m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&~m[1526]&m[1527])|(~m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&~m[1525]&m[1526]&m[1527])|(~m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&~m[1524]&m[1525]&m[1526]&m[1527])|(m[1521]&m[1524]&m[1525]&m[1526]&m[1527]));
    m[1528] = (((m[1526]&~m[1529]&~m[1530]&~m[1531]&~m[1532])|(~m[1526]&~m[1529]&~m[1530]&m[1531]&~m[1532])|(m[1526]&m[1529]&~m[1530]&m[1531]&~m[1532])|(m[1526]&~m[1529]&m[1530]&m[1531]&~m[1532])|(~m[1526]&m[1529]&~m[1530]&~m[1531]&m[1532])|(~m[1526]&~m[1529]&m[1530]&~m[1531]&m[1532])|(m[1526]&m[1529]&m[1530]&~m[1531]&m[1532])|(~m[1526]&m[1529]&m[1530]&m[1531]&m[1532]))&UnbiasedRNG[187])|((m[1526]&~m[1529]&~m[1530]&m[1531]&~m[1532])|(~m[1526]&~m[1529]&~m[1530]&~m[1531]&m[1532])|(m[1526]&~m[1529]&~m[1530]&~m[1531]&m[1532])|(m[1526]&m[1529]&~m[1530]&~m[1531]&m[1532])|(m[1526]&~m[1529]&m[1530]&~m[1531]&m[1532])|(~m[1526]&~m[1529]&~m[1530]&m[1531]&m[1532])|(m[1526]&~m[1529]&~m[1530]&m[1531]&m[1532])|(~m[1526]&m[1529]&~m[1530]&m[1531]&m[1532])|(m[1526]&m[1529]&~m[1530]&m[1531]&m[1532])|(~m[1526]&~m[1529]&m[1530]&m[1531]&m[1532])|(m[1526]&~m[1529]&m[1530]&m[1531]&m[1532])|(m[1526]&m[1529]&m[1530]&m[1531]&m[1532]));
    m[1533] = (((m[1502]&~m[1534]&~m[1535]&~m[1536]&~m[1537])|(~m[1502]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1502]&m[1534]&~m[1535]&m[1536]&~m[1537])|(m[1502]&~m[1534]&m[1535]&m[1536]&~m[1537])|(~m[1502]&m[1534]&~m[1535]&~m[1536]&m[1537])|(~m[1502]&~m[1534]&m[1535]&~m[1536]&m[1537])|(m[1502]&m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1502]&m[1534]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[188])|((m[1502]&~m[1534]&~m[1535]&m[1536]&~m[1537])|(~m[1502]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1502]&~m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1502]&m[1534]&~m[1535]&~m[1536]&m[1537])|(m[1502]&~m[1534]&m[1535]&~m[1536]&m[1537])|(~m[1502]&~m[1534]&~m[1535]&m[1536]&m[1537])|(m[1502]&~m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1502]&m[1534]&~m[1535]&m[1536]&m[1537])|(m[1502]&m[1534]&~m[1535]&m[1536]&m[1537])|(~m[1502]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1502]&~m[1534]&m[1535]&m[1536]&m[1537])|(m[1502]&m[1534]&m[1535]&m[1536]&m[1537]));
    m[1538] = (((m[1536]&~m[1539]&~m[1540]&~m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&~m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&~m[1542])|(~m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&m[1539]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[189])|((m[1536]&~m[1539]&~m[1540]&m[1541]&~m[1542])|(~m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&~m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&~m[1541]&m[1542])|(~m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&~m[1540]&m[1541]&m[1542])|(~m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&~m[1539]&m[1540]&m[1541]&m[1542])|(m[1536]&m[1539]&m[1540]&m[1541]&m[1542]));
    m[1543] = (((m[1541]&~m[1544]&~m[1545]&~m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&~m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&~m[1547])|(~m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&m[1544]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[190])|((m[1541]&~m[1544]&~m[1545]&m[1546]&~m[1547])|(~m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&~m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&~m[1546]&m[1547])|(~m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&~m[1545]&m[1546]&m[1547])|(~m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&~m[1544]&m[1545]&m[1546]&m[1547])|(m[1541]&m[1544]&m[1545]&m[1546]&m[1547]));
    m[1548] = (((m[1546]&~m[1549]&~m[1550]&~m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&~m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&~m[1552])|(~m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&m[1549]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[191])|((m[1546]&~m[1549]&~m[1550]&m[1551]&~m[1552])|(~m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&~m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&~m[1551]&m[1552])|(~m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&~m[1550]&m[1551]&m[1552])|(~m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&~m[1549]&m[1550]&m[1551]&m[1552])|(m[1546]&m[1549]&m[1550]&m[1551]&m[1552]));
    m[1553] = (((m[1551]&~m[1554]&~m[1555]&~m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&~m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&~m[1557])|(~m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&m[1554]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[192])|((m[1551]&~m[1554]&~m[1555]&m[1556]&~m[1557])|(~m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&~m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&~m[1556]&m[1557])|(~m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&~m[1555]&m[1556]&m[1557])|(~m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&~m[1554]&m[1555]&m[1556]&m[1557])|(m[1551]&m[1554]&m[1555]&m[1556]&m[1557]));
    m[1558] = (((m[1556]&~m[1559]&~m[1560]&~m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&~m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&~m[1562])|(~m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&m[1559]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[193])|((m[1556]&~m[1559]&~m[1560]&m[1561]&~m[1562])|(~m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&~m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&~m[1561]&m[1562])|(~m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&~m[1560]&m[1561]&m[1562])|(~m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&~m[1559]&m[1560]&m[1561]&m[1562])|(m[1556]&m[1559]&m[1560]&m[1561]&m[1562]));
    m[1563] = (((m[1537]&~m[1564]&~m[1565]&~m[1566]&~m[1567])|(~m[1537]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1537]&m[1564]&~m[1565]&m[1566]&~m[1567])|(m[1537]&~m[1564]&m[1565]&m[1566]&~m[1567])|(~m[1537]&m[1564]&~m[1565]&~m[1566]&m[1567])|(~m[1537]&~m[1564]&m[1565]&~m[1566]&m[1567])|(m[1537]&m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1537]&m[1564]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[194])|((m[1537]&~m[1564]&~m[1565]&m[1566]&~m[1567])|(~m[1537]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1537]&~m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1537]&m[1564]&~m[1565]&~m[1566]&m[1567])|(m[1537]&~m[1564]&m[1565]&~m[1566]&m[1567])|(~m[1537]&~m[1564]&~m[1565]&m[1566]&m[1567])|(m[1537]&~m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1537]&m[1564]&~m[1565]&m[1566]&m[1567])|(m[1537]&m[1564]&~m[1565]&m[1566]&m[1567])|(~m[1537]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1537]&~m[1564]&m[1565]&m[1566]&m[1567])|(m[1537]&m[1564]&m[1565]&m[1566]&m[1567]));
    m[1568] = (((m[1566]&~m[1569]&~m[1570]&~m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&~m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&~m[1572])|(~m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&m[1569]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[195])|((m[1566]&~m[1569]&~m[1570]&m[1571]&~m[1572])|(~m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&~m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&~m[1571]&m[1572])|(~m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&~m[1570]&m[1571]&m[1572])|(~m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&~m[1569]&m[1570]&m[1571]&m[1572])|(m[1566]&m[1569]&m[1570]&m[1571]&m[1572]));
    m[1573] = (((m[1571]&~m[1574]&~m[1575]&~m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&~m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&~m[1577])|(~m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&m[1574]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[196])|((m[1571]&~m[1574]&~m[1575]&m[1576]&~m[1577])|(~m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&~m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&~m[1576]&m[1577])|(~m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&~m[1575]&m[1576]&m[1577])|(~m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&~m[1574]&m[1575]&m[1576]&m[1577])|(m[1571]&m[1574]&m[1575]&m[1576]&m[1577]));
    m[1578] = (((m[1576]&~m[1579]&~m[1580]&~m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&~m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&~m[1582])|(~m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&m[1579]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[197])|((m[1576]&~m[1579]&~m[1580]&m[1581]&~m[1582])|(~m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&~m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&~m[1581]&m[1582])|(~m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&~m[1580]&m[1581]&m[1582])|(~m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&~m[1579]&m[1580]&m[1581]&m[1582])|(m[1576]&m[1579]&m[1580]&m[1581]&m[1582]));
    m[1583] = (((m[1581]&~m[1584]&~m[1585]&~m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&~m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&~m[1587])|(~m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&m[1584]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[198])|((m[1581]&~m[1584]&~m[1585]&m[1586]&~m[1587])|(~m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&~m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&~m[1586]&m[1587])|(~m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&~m[1585]&m[1586]&m[1587])|(~m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&~m[1584]&m[1585]&m[1586]&m[1587])|(m[1581]&m[1584]&m[1585]&m[1586]&m[1587]));
    m[1588] = (((m[1567]&~m[1589]&~m[1590]&~m[1591]&~m[1592])|(~m[1567]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1567]&m[1589]&~m[1590]&m[1591]&~m[1592])|(m[1567]&~m[1589]&m[1590]&m[1591]&~m[1592])|(~m[1567]&m[1589]&~m[1590]&~m[1591]&m[1592])|(~m[1567]&~m[1589]&m[1590]&~m[1591]&m[1592])|(m[1567]&m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1567]&m[1589]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[199])|((m[1567]&~m[1589]&~m[1590]&m[1591]&~m[1592])|(~m[1567]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1567]&~m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1567]&m[1589]&~m[1590]&~m[1591]&m[1592])|(m[1567]&~m[1589]&m[1590]&~m[1591]&m[1592])|(~m[1567]&~m[1589]&~m[1590]&m[1591]&m[1592])|(m[1567]&~m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1567]&m[1589]&~m[1590]&m[1591]&m[1592])|(m[1567]&m[1589]&~m[1590]&m[1591]&m[1592])|(~m[1567]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1567]&~m[1589]&m[1590]&m[1591]&m[1592])|(m[1567]&m[1589]&m[1590]&m[1591]&m[1592]));
    m[1593] = (((m[1591]&~m[1594]&~m[1595]&~m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&~m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&~m[1597])|(~m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&m[1594]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[200])|((m[1591]&~m[1594]&~m[1595]&m[1596]&~m[1597])|(~m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&~m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&~m[1596]&m[1597])|(~m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&~m[1595]&m[1596]&m[1597])|(~m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&~m[1594]&m[1595]&m[1596]&m[1597])|(m[1591]&m[1594]&m[1595]&m[1596]&m[1597]));
    m[1598] = (((m[1596]&~m[1599]&~m[1600]&~m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&~m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&~m[1602])|(~m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&m[1599]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[201])|((m[1596]&~m[1599]&~m[1600]&m[1601]&~m[1602])|(~m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&~m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&~m[1601]&m[1602])|(~m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&~m[1600]&m[1601]&m[1602])|(~m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&~m[1599]&m[1600]&m[1601]&m[1602])|(m[1596]&m[1599]&m[1600]&m[1601]&m[1602]));
    m[1603] = (((m[1601]&~m[1604]&~m[1605]&~m[1606]&~m[1607])|(~m[1601]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1601]&m[1604]&~m[1605]&m[1606]&~m[1607])|(m[1601]&~m[1604]&m[1605]&m[1606]&~m[1607])|(~m[1601]&m[1604]&~m[1605]&~m[1606]&m[1607])|(~m[1601]&~m[1604]&m[1605]&~m[1606]&m[1607])|(m[1601]&m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1601]&m[1604]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[202])|((m[1601]&~m[1604]&~m[1605]&m[1606]&~m[1607])|(~m[1601]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1601]&~m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1601]&m[1604]&~m[1605]&~m[1606]&m[1607])|(m[1601]&~m[1604]&m[1605]&~m[1606]&m[1607])|(~m[1601]&~m[1604]&~m[1605]&m[1606]&m[1607])|(m[1601]&~m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1601]&m[1604]&~m[1605]&m[1606]&m[1607])|(m[1601]&m[1604]&~m[1605]&m[1606]&m[1607])|(~m[1601]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1601]&~m[1604]&m[1605]&m[1606]&m[1607])|(m[1601]&m[1604]&m[1605]&m[1606]&m[1607]));
    m[1608] = (((m[1592]&~m[1609]&~m[1610]&~m[1611]&~m[1612])|(~m[1592]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1592]&m[1609]&~m[1610]&m[1611]&~m[1612])|(m[1592]&~m[1609]&m[1610]&m[1611]&~m[1612])|(~m[1592]&m[1609]&~m[1610]&~m[1611]&m[1612])|(~m[1592]&~m[1609]&m[1610]&~m[1611]&m[1612])|(m[1592]&m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1592]&m[1609]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[203])|((m[1592]&~m[1609]&~m[1610]&m[1611]&~m[1612])|(~m[1592]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1592]&~m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1592]&m[1609]&~m[1610]&~m[1611]&m[1612])|(m[1592]&~m[1609]&m[1610]&~m[1611]&m[1612])|(~m[1592]&~m[1609]&~m[1610]&m[1611]&m[1612])|(m[1592]&~m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1592]&m[1609]&~m[1610]&m[1611]&m[1612])|(m[1592]&m[1609]&~m[1610]&m[1611]&m[1612])|(~m[1592]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1592]&~m[1609]&m[1610]&m[1611]&m[1612])|(m[1592]&m[1609]&m[1610]&m[1611]&m[1612]));
    m[1613] = (((m[1611]&~m[1614]&~m[1615]&~m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&~m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&~m[1617])|(~m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&m[1614]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[204])|((m[1611]&~m[1614]&~m[1615]&m[1616]&~m[1617])|(~m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&~m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&~m[1616]&m[1617])|(~m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&~m[1615]&m[1616]&m[1617])|(~m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&~m[1614]&m[1615]&m[1616]&m[1617])|(m[1611]&m[1614]&m[1615]&m[1616]&m[1617]));
    m[1618] = (((m[1616]&~m[1619]&~m[1620]&~m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&~m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&~m[1622])|(~m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&m[1619]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[205])|((m[1616]&~m[1619]&~m[1620]&m[1621]&~m[1622])|(~m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&~m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&~m[1621]&m[1622])|(~m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&~m[1620]&m[1621]&m[1622])|(~m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&~m[1619]&m[1620]&m[1621]&m[1622])|(m[1616]&m[1619]&m[1620]&m[1621]&m[1622]));
    m[1623] = (((m[1612]&~m[1624]&~m[1625]&~m[1626]&~m[1627])|(~m[1612]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1612]&m[1624]&~m[1625]&m[1626]&~m[1627])|(m[1612]&~m[1624]&m[1625]&m[1626]&~m[1627])|(~m[1612]&m[1624]&~m[1625]&~m[1626]&m[1627])|(~m[1612]&~m[1624]&m[1625]&~m[1626]&m[1627])|(m[1612]&m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1612]&m[1624]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[206])|((m[1612]&~m[1624]&~m[1625]&m[1626]&~m[1627])|(~m[1612]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1612]&~m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1612]&m[1624]&~m[1625]&~m[1626]&m[1627])|(m[1612]&~m[1624]&m[1625]&~m[1626]&m[1627])|(~m[1612]&~m[1624]&~m[1625]&m[1626]&m[1627])|(m[1612]&~m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1612]&m[1624]&~m[1625]&m[1626]&m[1627])|(m[1612]&m[1624]&~m[1625]&m[1626]&m[1627])|(~m[1612]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1612]&~m[1624]&m[1625]&m[1626]&m[1627])|(m[1612]&m[1624]&m[1625]&m[1626]&m[1627]));
    m[1628] = (((m[1626]&~m[1629]&~m[1630]&~m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&~m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&~m[1632])|(~m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&m[1629]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[207])|((m[1626]&~m[1629]&~m[1630]&m[1631]&~m[1632])|(~m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&~m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&~m[1631]&m[1632])|(~m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&~m[1630]&m[1631]&m[1632])|(~m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&~m[1629]&m[1630]&m[1631]&m[1632])|(m[1626]&m[1629]&m[1630]&m[1631]&m[1632]));
    m[1633] = (((m[1627]&~m[1634]&~m[1635]&~m[1636]&~m[1637])|(~m[1627]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1627]&m[1634]&~m[1635]&m[1636]&~m[1637])|(m[1627]&~m[1634]&m[1635]&m[1636]&~m[1637])|(~m[1627]&m[1634]&~m[1635]&~m[1636]&m[1637])|(~m[1627]&~m[1634]&m[1635]&~m[1636]&m[1637])|(m[1627]&m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1627]&m[1634]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[208])|((m[1627]&~m[1634]&~m[1635]&m[1636]&~m[1637])|(~m[1627]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1627]&~m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1627]&m[1634]&~m[1635]&~m[1636]&m[1637])|(m[1627]&~m[1634]&m[1635]&~m[1636]&m[1637])|(~m[1627]&~m[1634]&~m[1635]&m[1636]&m[1637])|(m[1627]&~m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1627]&m[1634]&~m[1635]&m[1636]&m[1637])|(m[1627]&m[1634]&~m[1635]&m[1636]&m[1637])|(~m[1627]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1627]&~m[1634]&m[1635]&m[1636]&m[1637])|(m[1627]&m[1634]&m[1635]&m[1636]&m[1637]));
end

always @(posedge color1_clk) begin
    m[28] = (((m[0]&m[57]&~m[58]&~m[140]&~m[141])|(m[0]&~m[57]&m[58]&~m[140]&~m[141])|(~m[0]&m[57]&m[58]&~m[140]&~m[141])|(m[0]&~m[57]&~m[58]&m[140]&~m[141])|(~m[0]&m[57]&~m[58]&m[140]&~m[141])|(~m[0]&~m[57]&m[58]&m[140]&~m[141])|(m[0]&~m[57]&~m[58]&~m[140]&m[141])|(~m[0]&m[57]&~m[58]&~m[140]&m[141])|(~m[0]&~m[57]&m[58]&~m[140]&m[141])|(~m[0]&~m[57]&~m[58]&m[140]&m[141]))&BiasedRNG[252])|(((m[0]&m[57]&m[58]&~m[140]&~m[141])|(m[0]&m[57]&~m[58]&m[140]&~m[141])|(m[0]&~m[57]&m[58]&m[140]&~m[141])|(~m[0]&m[57]&m[58]&m[140]&~m[141])|(m[0]&m[57]&~m[58]&~m[140]&m[141])|(m[0]&~m[57]&m[58]&~m[140]&m[141])|(~m[0]&m[57]&m[58]&~m[140]&m[141])|(m[0]&~m[57]&~m[58]&m[140]&m[141])|(~m[0]&m[57]&~m[58]&m[140]&m[141])|(~m[0]&~m[57]&m[58]&m[140]&m[141]))&~BiasedRNG[252])|((m[0]&m[57]&m[58]&m[140]&~m[141])|(m[0]&m[57]&m[58]&~m[140]&m[141])|(m[0]&m[57]&~m[58]&m[140]&m[141])|(m[0]&~m[57]&m[58]&m[140]&m[141])|(~m[0]&m[57]&m[58]&m[140]&m[141])|(m[0]&m[57]&m[58]&m[140]&m[141]));
    m[29] = (((m[1]&m[60]&~m[61]&~m[154]&~m[155])|(m[1]&~m[60]&m[61]&~m[154]&~m[155])|(~m[1]&m[60]&m[61]&~m[154]&~m[155])|(m[1]&~m[60]&~m[61]&m[154]&~m[155])|(~m[1]&m[60]&~m[61]&m[154]&~m[155])|(~m[1]&~m[60]&m[61]&m[154]&~m[155])|(m[1]&~m[60]&~m[61]&~m[154]&m[155])|(~m[1]&m[60]&~m[61]&~m[154]&m[155])|(~m[1]&~m[60]&m[61]&~m[154]&m[155])|(~m[1]&~m[60]&~m[61]&m[154]&m[155]))&BiasedRNG[253])|(((m[1]&m[60]&m[61]&~m[154]&~m[155])|(m[1]&m[60]&~m[61]&m[154]&~m[155])|(m[1]&~m[60]&m[61]&m[154]&~m[155])|(~m[1]&m[60]&m[61]&m[154]&~m[155])|(m[1]&m[60]&~m[61]&~m[154]&m[155])|(m[1]&~m[60]&m[61]&~m[154]&m[155])|(~m[1]&m[60]&m[61]&~m[154]&m[155])|(m[1]&~m[60]&~m[61]&m[154]&m[155])|(~m[1]&m[60]&~m[61]&m[154]&m[155])|(~m[1]&~m[60]&m[61]&m[154]&m[155]))&~BiasedRNG[253])|((m[1]&m[60]&m[61]&m[154]&~m[155])|(m[1]&m[60]&m[61]&~m[154]&m[155])|(m[1]&m[60]&~m[61]&m[154]&m[155])|(m[1]&~m[60]&m[61]&m[154]&m[155])|(~m[1]&m[60]&m[61]&m[154]&m[155])|(m[1]&m[60]&m[61]&m[154]&m[155]));
    m[30] = (((m[2]&m[63]&~m[64]&~m[168]&~m[169])|(m[2]&~m[63]&m[64]&~m[168]&~m[169])|(~m[2]&m[63]&m[64]&~m[168]&~m[169])|(m[2]&~m[63]&~m[64]&m[168]&~m[169])|(~m[2]&m[63]&~m[64]&m[168]&~m[169])|(~m[2]&~m[63]&m[64]&m[168]&~m[169])|(m[2]&~m[63]&~m[64]&~m[168]&m[169])|(~m[2]&m[63]&~m[64]&~m[168]&m[169])|(~m[2]&~m[63]&m[64]&~m[168]&m[169])|(~m[2]&~m[63]&~m[64]&m[168]&m[169]))&BiasedRNG[254])|(((m[2]&m[63]&m[64]&~m[168]&~m[169])|(m[2]&m[63]&~m[64]&m[168]&~m[169])|(m[2]&~m[63]&m[64]&m[168]&~m[169])|(~m[2]&m[63]&m[64]&m[168]&~m[169])|(m[2]&m[63]&~m[64]&~m[168]&m[169])|(m[2]&~m[63]&m[64]&~m[168]&m[169])|(~m[2]&m[63]&m[64]&~m[168]&m[169])|(m[2]&~m[63]&~m[64]&m[168]&m[169])|(~m[2]&m[63]&~m[64]&m[168]&m[169])|(~m[2]&~m[63]&m[64]&m[168]&m[169]))&~BiasedRNG[254])|((m[2]&m[63]&m[64]&m[168]&~m[169])|(m[2]&m[63]&m[64]&~m[168]&m[169])|(m[2]&m[63]&~m[64]&m[168]&m[169])|(m[2]&~m[63]&m[64]&m[168]&m[169])|(~m[2]&m[63]&m[64]&m[168]&m[169])|(m[2]&m[63]&m[64]&m[168]&m[169]));
    m[31] = (((m[3]&m[66]&~m[67]&~m[182]&~m[183])|(m[3]&~m[66]&m[67]&~m[182]&~m[183])|(~m[3]&m[66]&m[67]&~m[182]&~m[183])|(m[3]&~m[66]&~m[67]&m[182]&~m[183])|(~m[3]&m[66]&~m[67]&m[182]&~m[183])|(~m[3]&~m[66]&m[67]&m[182]&~m[183])|(m[3]&~m[66]&~m[67]&~m[182]&m[183])|(~m[3]&m[66]&~m[67]&~m[182]&m[183])|(~m[3]&~m[66]&m[67]&~m[182]&m[183])|(~m[3]&~m[66]&~m[67]&m[182]&m[183]))&BiasedRNG[255])|(((m[3]&m[66]&m[67]&~m[182]&~m[183])|(m[3]&m[66]&~m[67]&m[182]&~m[183])|(m[3]&~m[66]&m[67]&m[182]&~m[183])|(~m[3]&m[66]&m[67]&m[182]&~m[183])|(m[3]&m[66]&~m[67]&~m[182]&m[183])|(m[3]&~m[66]&m[67]&~m[182]&m[183])|(~m[3]&m[66]&m[67]&~m[182]&m[183])|(m[3]&~m[66]&~m[67]&m[182]&m[183])|(~m[3]&m[66]&~m[67]&m[182]&m[183])|(~m[3]&~m[66]&m[67]&m[182]&m[183]))&~BiasedRNG[255])|((m[3]&m[66]&m[67]&m[182]&~m[183])|(m[3]&m[66]&m[67]&~m[182]&m[183])|(m[3]&m[66]&~m[67]&m[182]&m[183])|(m[3]&~m[66]&m[67]&m[182]&m[183])|(~m[3]&m[66]&m[67]&m[182]&m[183])|(m[3]&m[66]&m[67]&m[182]&m[183]));
    m[32] = (((m[4]&m[69]&~m[70]&~m[196]&~m[197])|(m[4]&~m[69]&m[70]&~m[196]&~m[197])|(~m[4]&m[69]&m[70]&~m[196]&~m[197])|(m[4]&~m[69]&~m[70]&m[196]&~m[197])|(~m[4]&m[69]&~m[70]&m[196]&~m[197])|(~m[4]&~m[69]&m[70]&m[196]&~m[197])|(m[4]&~m[69]&~m[70]&~m[196]&m[197])|(~m[4]&m[69]&~m[70]&~m[196]&m[197])|(~m[4]&~m[69]&m[70]&~m[196]&m[197])|(~m[4]&~m[69]&~m[70]&m[196]&m[197]))&BiasedRNG[256])|(((m[4]&m[69]&m[70]&~m[196]&~m[197])|(m[4]&m[69]&~m[70]&m[196]&~m[197])|(m[4]&~m[69]&m[70]&m[196]&~m[197])|(~m[4]&m[69]&m[70]&m[196]&~m[197])|(m[4]&m[69]&~m[70]&~m[196]&m[197])|(m[4]&~m[69]&m[70]&~m[196]&m[197])|(~m[4]&m[69]&m[70]&~m[196]&m[197])|(m[4]&~m[69]&~m[70]&m[196]&m[197])|(~m[4]&m[69]&~m[70]&m[196]&m[197])|(~m[4]&~m[69]&m[70]&m[196]&m[197]))&~BiasedRNG[256])|((m[4]&m[69]&m[70]&m[196]&~m[197])|(m[4]&m[69]&m[70]&~m[196]&m[197])|(m[4]&m[69]&~m[70]&m[196]&m[197])|(m[4]&~m[69]&m[70]&m[196]&m[197])|(~m[4]&m[69]&m[70]&m[196]&m[197])|(m[4]&m[69]&m[70]&m[196]&m[197]));
    m[33] = (((m[5]&m[72]&~m[73]&~m[210]&~m[211])|(m[5]&~m[72]&m[73]&~m[210]&~m[211])|(~m[5]&m[72]&m[73]&~m[210]&~m[211])|(m[5]&~m[72]&~m[73]&m[210]&~m[211])|(~m[5]&m[72]&~m[73]&m[210]&~m[211])|(~m[5]&~m[72]&m[73]&m[210]&~m[211])|(m[5]&~m[72]&~m[73]&~m[210]&m[211])|(~m[5]&m[72]&~m[73]&~m[210]&m[211])|(~m[5]&~m[72]&m[73]&~m[210]&m[211])|(~m[5]&~m[72]&~m[73]&m[210]&m[211]))&BiasedRNG[257])|(((m[5]&m[72]&m[73]&~m[210]&~m[211])|(m[5]&m[72]&~m[73]&m[210]&~m[211])|(m[5]&~m[72]&m[73]&m[210]&~m[211])|(~m[5]&m[72]&m[73]&m[210]&~m[211])|(m[5]&m[72]&~m[73]&~m[210]&m[211])|(m[5]&~m[72]&m[73]&~m[210]&m[211])|(~m[5]&m[72]&m[73]&~m[210]&m[211])|(m[5]&~m[72]&~m[73]&m[210]&m[211])|(~m[5]&m[72]&~m[73]&m[210]&m[211])|(~m[5]&~m[72]&m[73]&m[210]&m[211]))&~BiasedRNG[257])|((m[5]&m[72]&m[73]&m[210]&~m[211])|(m[5]&m[72]&m[73]&~m[210]&m[211])|(m[5]&m[72]&~m[73]&m[210]&m[211])|(m[5]&~m[72]&m[73]&m[210]&m[211])|(~m[5]&m[72]&m[73]&m[210]&m[211])|(m[5]&m[72]&m[73]&m[210]&m[211]));
    m[34] = (((m[6]&m[75]&~m[76]&~m[224]&~m[225])|(m[6]&~m[75]&m[76]&~m[224]&~m[225])|(~m[6]&m[75]&m[76]&~m[224]&~m[225])|(m[6]&~m[75]&~m[76]&m[224]&~m[225])|(~m[6]&m[75]&~m[76]&m[224]&~m[225])|(~m[6]&~m[75]&m[76]&m[224]&~m[225])|(m[6]&~m[75]&~m[76]&~m[224]&m[225])|(~m[6]&m[75]&~m[76]&~m[224]&m[225])|(~m[6]&~m[75]&m[76]&~m[224]&m[225])|(~m[6]&~m[75]&~m[76]&m[224]&m[225]))&BiasedRNG[258])|(((m[6]&m[75]&m[76]&~m[224]&~m[225])|(m[6]&m[75]&~m[76]&m[224]&~m[225])|(m[6]&~m[75]&m[76]&m[224]&~m[225])|(~m[6]&m[75]&m[76]&m[224]&~m[225])|(m[6]&m[75]&~m[76]&~m[224]&m[225])|(m[6]&~m[75]&m[76]&~m[224]&m[225])|(~m[6]&m[75]&m[76]&~m[224]&m[225])|(m[6]&~m[75]&~m[76]&m[224]&m[225])|(~m[6]&m[75]&~m[76]&m[224]&m[225])|(~m[6]&~m[75]&m[76]&m[224]&m[225]))&~BiasedRNG[258])|((m[6]&m[75]&m[76]&m[224]&~m[225])|(m[6]&m[75]&m[76]&~m[224]&m[225])|(m[6]&m[75]&~m[76]&m[224]&m[225])|(m[6]&~m[75]&m[76]&m[224]&m[225])|(~m[6]&m[75]&m[76]&m[224]&m[225])|(m[6]&m[75]&m[76]&m[224]&m[225]));
    m[35] = (((m[7]&m[78]&~m[79]&~m[238]&~m[239])|(m[7]&~m[78]&m[79]&~m[238]&~m[239])|(~m[7]&m[78]&m[79]&~m[238]&~m[239])|(m[7]&~m[78]&~m[79]&m[238]&~m[239])|(~m[7]&m[78]&~m[79]&m[238]&~m[239])|(~m[7]&~m[78]&m[79]&m[238]&~m[239])|(m[7]&~m[78]&~m[79]&~m[238]&m[239])|(~m[7]&m[78]&~m[79]&~m[238]&m[239])|(~m[7]&~m[78]&m[79]&~m[238]&m[239])|(~m[7]&~m[78]&~m[79]&m[238]&m[239]))&BiasedRNG[259])|(((m[7]&m[78]&m[79]&~m[238]&~m[239])|(m[7]&m[78]&~m[79]&m[238]&~m[239])|(m[7]&~m[78]&m[79]&m[238]&~m[239])|(~m[7]&m[78]&m[79]&m[238]&~m[239])|(m[7]&m[78]&~m[79]&~m[238]&m[239])|(m[7]&~m[78]&m[79]&~m[238]&m[239])|(~m[7]&m[78]&m[79]&~m[238]&m[239])|(m[7]&~m[78]&~m[79]&m[238]&m[239])|(~m[7]&m[78]&~m[79]&m[238]&m[239])|(~m[7]&~m[78]&m[79]&m[238]&m[239]))&~BiasedRNG[259])|((m[7]&m[78]&m[79]&m[238]&~m[239])|(m[7]&m[78]&m[79]&~m[238]&m[239])|(m[7]&m[78]&~m[79]&m[238]&m[239])|(m[7]&~m[78]&m[79]&m[238]&m[239])|(~m[7]&m[78]&m[79]&m[238]&m[239])|(m[7]&m[78]&m[79]&m[238]&m[239]));
    m[36] = (((m[8]&m[81]&~m[82]&~m[252]&~m[253])|(m[8]&~m[81]&m[82]&~m[252]&~m[253])|(~m[8]&m[81]&m[82]&~m[252]&~m[253])|(m[8]&~m[81]&~m[82]&m[252]&~m[253])|(~m[8]&m[81]&~m[82]&m[252]&~m[253])|(~m[8]&~m[81]&m[82]&m[252]&~m[253])|(m[8]&~m[81]&~m[82]&~m[252]&m[253])|(~m[8]&m[81]&~m[82]&~m[252]&m[253])|(~m[8]&~m[81]&m[82]&~m[252]&m[253])|(~m[8]&~m[81]&~m[82]&m[252]&m[253]))&BiasedRNG[260])|(((m[8]&m[81]&m[82]&~m[252]&~m[253])|(m[8]&m[81]&~m[82]&m[252]&~m[253])|(m[8]&~m[81]&m[82]&m[252]&~m[253])|(~m[8]&m[81]&m[82]&m[252]&~m[253])|(m[8]&m[81]&~m[82]&~m[252]&m[253])|(m[8]&~m[81]&m[82]&~m[252]&m[253])|(~m[8]&m[81]&m[82]&~m[252]&m[253])|(m[8]&~m[81]&~m[82]&m[252]&m[253])|(~m[8]&m[81]&~m[82]&m[252]&m[253])|(~m[8]&~m[81]&m[82]&m[252]&m[253]))&~BiasedRNG[260])|((m[8]&m[81]&m[82]&m[252]&~m[253])|(m[8]&m[81]&m[82]&~m[252]&m[253])|(m[8]&m[81]&~m[82]&m[252]&m[253])|(m[8]&~m[81]&m[82]&m[252]&m[253])|(~m[8]&m[81]&m[82]&m[252]&m[253])|(m[8]&m[81]&m[82]&m[252]&m[253]));
    m[37] = (((m[9]&m[84]&~m[85]&~m[266]&~m[267])|(m[9]&~m[84]&m[85]&~m[266]&~m[267])|(~m[9]&m[84]&m[85]&~m[266]&~m[267])|(m[9]&~m[84]&~m[85]&m[266]&~m[267])|(~m[9]&m[84]&~m[85]&m[266]&~m[267])|(~m[9]&~m[84]&m[85]&m[266]&~m[267])|(m[9]&~m[84]&~m[85]&~m[266]&m[267])|(~m[9]&m[84]&~m[85]&~m[266]&m[267])|(~m[9]&~m[84]&m[85]&~m[266]&m[267])|(~m[9]&~m[84]&~m[85]&m[266]&m[267]))&BiasedRNG[261])|(((m[9]&m[84]&m[85]&~m[266]&~m[267])|(m[9]&m[84]&~m[85]&m[266]&~m[267])|(m[9]&~m[84]&m[85]&m[266]&~m[267])|(~m[9]&m[84]&m[85]&m[266]&~m[267])|(m[9]&m[84]&~m[85]&~m[266]&m[267])|(m[9]&~m[84]&m[85]&~m[266]&m[267])|(~m[9]&m[84]&m[85]&~m[266]&m[267])|(m[9]&~m[84]&~m[85]&m[266]&m[267])|(~m[9]&m[84]&~m[85]&m[266]&m[267])|(~m[9]&~m[84]&m[85]&m[266]&m[267]))&~BiasedRNG[261])|((m[9]&m[84]&m[85]&m[266]&~m[267])|(m[9]&m[84]&m[85]&~m[266]&m[267])|(m[9]&m[84]&~m[85]&m[266]&m[267])|(m[9]&~m[84]&m[85]&m[266]&m[267])|(~m[9]&m[84]&m[85]&m[266]&m[267])|(m[9]&m[84]&m[85]&m[266]&m[267]));
    m[38] = (((m[10]&m[87]&~m[88]&~m[280]&~m[281])|(m[10]&~m[87]&m[88]&~m[280]&~m[281])|(~m[10]&m[87]&m[88]&~m[280]&~m[281])|(m[10]&~m[87]&~m[88]&m[280]&~m[281])|(~m[10]&m[87]&~m[88]&m[280]&~m[281])|(~m[10]&~m[87]&m[88]&m[280]&~m[281])|(m[10]&~m[87]&~m[88]&~m[280]&m[281])|(~m[10]&m[87]&~m[88]&~m[280]&m[281])|(~m[10]&~m[87]&m[88]&~m[280]&m[281])|(~m[10]&~m[87]&~m[88]&m[280]&m[281]))&BiasedRNG[262])|(((m[10]&m[87]&m[88]&~m[280]&~m[281])|(m[10]&m[87]&~m[88]&m[280]&~m[281])|(m[10]&~m[87]&m[88]&m[280]&~m[281])|(~m[10]&m[87]&m[88]&m[280]&~m[281])|(m[10]&m[87]&~m[88]&~m[280]&m[281])|(m[10]&~m[87]&m[88]&~m[280]&m[281])|(~m[10]&m[87]&m[88]&~m[280]&m[281])|(m[10]&~m[87]&~m[88]&m[280]&m[281])|(~m[10]&m[87]&~m[88]&m[280]&m[281])|(~m[10]&~m[87]&m[88]&m[280]&m[281]))&~BiasedRNG[262])|((m[10]&m[87]&m[88]&m[280]&~m[281])|(m[10]&m[87]&m[88]&~m[280]&m[281])|(m[10]&m[87]&~m[88]&m[280]&m[281])|(m[10]&~m[87]&m[88]&m[280]&m[281])|(~m[10]&m[87]&m[88]&m[280]&m[281])|(m[10]&m[87]&m[88]&m[280]&m[281]));
    m[39] = (((m[11]&m[90]&~m[91]&~m[294]&~m[295])|(m[11]&~m[90]&m[91]&~m[294]&~m[295])|(~m[11]&m[90]&m[91]&~m[294]&~m[295])|(m[11]&~m[90]&~m[91]&m[294]&~m[295])|(~m[11]&m[90]&~m[91]&m[294]&~m[295])|(~m[11]&~m[90]&m[91]&m[294]&~m[295])|(m[11]&~m[90]&~m[91]&~m[294]&m[295])|(~m[11]&m[90]&~m[91]&~m[294]&m[295])|(~m[11]&~m[90]&m[91]&~m[294]&m[295])|(~m[11]&~m[90]&~m[91]&m[294]&m[295]))&BiasedRNG[263])|(((m[11]&m[90]&m[91]&~m[294]&~m[295])|(m[11]&m[90]&~m[91]&m[294]&~m[295])|(m[11]&~m[90]&m[91]&m[294]&~m[295])|(~m[11]&m[90]&m[91]&m[294]&~m[295])|(m[11]&m[90]&~m[91]&~m[294]&m[295])|(m[11]&~m[90]&m[91]&~m[294]&m[295])|(~m[11]&m[90]&m[91]&~m[294]&m[295])|(m[11]&~m[90]&~m[91]&m[294]&m[295])|(~m[11]&m[90]&~m[91]&m[294]&m[295])|(~m[11]&~m[90]&m[91]&m[294]&m[295]))&~BiasedRNG[263])|((m[11]&m[90]&m[91]&m[294]&~m[295])|(m[11]&m[90]&m[91]&~m[294]&m[295])|(m[11]&m[90]&~m[91]&m[294]&m[295])|(m[11]&~m[90]&m[91]&m[294]&m[295])|(~m[11]&m[90]&m[91]&m[294]&m[295])|(m[11]&m[90]&m[91]&m[294]&m[295]));
    m[40] = (((m[12]&m[93]&~m[94]&~m[308]&~m[309])|(m[12]&~m[93]&m[94]&~m[308]&~m[309])|(~m[12]&m[93]&m[94]&~m[308]&~m[309])|(m[12]&~m[93]&~m[94]&m[308]&~m[309])|(~m[12]&m[93]&~m[94]&m[308]&~m[309])|(~m[12]&~m[93]&m[94]&m[308]&~m[309])|(m[12]&~m[93]&~m[94]&~m[308]&m[309])|(~m[12]&m[93]&~m[94]&~m[308]&m[309])|(~m[12]&~m[93]&m[94]&~m[308]&m[309])|(~m[12]&~m[93]&~m[94]&m[308]&m[309]))&BiasedRNG[264])|(((m[12]&m[93]&m[94]&~m[308]&~m[309])|(m[12]&m[93]&~m[94]&m[308]&~m[309])|(m[12]&~m[93]&m[94]&m[308]&~m[309])|(~m[12]&m[93]&m[94]&m[308]&~m[309])|(m[12]&m[93]&~m[94]&~m[308]&m[309])|(m[12]&~m[93]&m[94]&~m[308]&m[309])|(~m[12]&m[93]&m[94]&~m[308]&m[309])|(m[12]&~m[93]&~m[94]&m[308]&m[309])|(~m[12]&m[93]&~m[94]&m[308]&m[309])|(~m[12]&~m[93]&m[94]&m[308]&m[309]))&~BiasedRNG[264])|((m[12]&m[93]&m[94]&m[308]&~m[309])|(m[12]&m[93]&m[94]&~m[308]&m[309])|(m[12]&m[93]&~m[94]&m[308]&m[309])|(m[12]&~m[93]&m[94]&m[308]&m[309])|(~m[12]&m[93]&m[94]&m[308]&m[309])|(m[12]&m[93]&m[94]&m[308]&m[309]));
    m[41] = (((m[13]&m[96]&~m[97]&~m[322]&~m[323])|(m[13]&~m[96]&m[97]&~m[322]&~m[323])|(~m[13]&m[96]&m[97]&~m[322]&~m[323])|(m[13]&~m[96]&~m[97]&m[322]&~m[323])|(~m[13]&m[96]&~m[97]&m[322]&~m[323])|(~m[13]&~m[96]&m[97]&m[322]&~m[323])|(m[13]&~m[96]&~m[97]&~m[322]&m[323])|(~m[13]&m[96]&~m[97]&~m[322]&m[323])|(~m[13]&~m[96]&m[97]&~m[322]&m[323])|(~m[13]&~m[96]&~m[97]&m[322]&m[323]))&BiasedRNG[265])|(((m[13]&m[96]&m[97]&~m[322]&~m[323])|(m[13]&m[96]&~m[97]&m[322]&~m[323])|(m[13]&~m[96]&m[97]&m[322]&~m[323])|(~m[13]&m[96]&m[97]&m[322]&~m[323])|(m[13]&m[96]&~m[97]&~m[322]&m[323])|(m[13]&~m[96]&m[97]&~m[322]&m[323])|(~m[13]&m[96]&m[97]&~m[322]&m[323])|(m[13]&~m[96]&~m[97]&m[322]&m[323])|(~m[13]&m[96]&~m[97]&m[322]&m[323])|(~m[13]&~m[96]&m[97]&m[322]&m[323]))&~BiasedRNG[265])|((m[13]&m[96]&m[97]&m[322]&~m[323])|(m[13]&m[96]&m[97]&~m[322]&m[323])|(m[13]&m[96]&~m[97]&m[322]&m[323])|(m[13]&~m[96]&m[97]&m[322]&m[323])|(~m[13]&m[96]&m[97]&m[322]&m[323])|(m[13]&m[96]&m[97]&m[322]&m[323]));
    m[42] = (((m[14]&m[99]&~m[100]&~m[336]&~m[337])|(m[14]&~m[99]&m[100]&~m[336]&~m[337])|(~m[14]&m[99]&m[100]&~m[336]&~m[337])|(m[14]&~m[99]&~m[100]&m[336]&~m[337])|(~m[14]&m[99]&~m[100]&m[336]&~m[337])|(~m[14]&~m[99]&m[100]&m[336]&~m[337])|(m[14]&~m[99]&~m[100]&~m[336]&m[337])|(~m[14]&m[99]&~m[100]&~m[336]&m[337])|(~m[14]&~m[99]&m[100]&~m[336]&m[337])|(~m[14]&~m[99]&~m[100]&m[336]&m[337]))&BiasedRNG[266])|(((m[14]&m[99]&m[100]&~m[336]&~m[337])|(m[14]&m[99]&~m[100]&m[336]&~m[337])|(m[14]&~m[99]&m[100]&m[336]&~m[337])|(~m[14]&m[99]&m[100]&m[336]&~m[337])|(m[14]&m[99]&~m[100]&~m[336]&m[337])|(m[14]&~m[99]&m[100]&~m[336]&m[337])|(~m[14]&m[99]&m[100]&~m[336]&m[337])|(m[14]&~m[99]&~m[100]&m[336]&m[337])|(~m[14]&m[99]&~m[100]&m[336]&m[337])|(~m[14]&~m[99]&m[100]&m[336]&m[337]))&~BiasedRNG[266])|((m[14]&m[99]&m[100]&m[336]&~m[337])|(m[14]&m[99]&m[100]&~m[336]&m[337])|(m[14]&m[99]&~m[100]&m[336]&m[337])|(m[14]&~m[99]&m[100]&m[336]&m[337])|(~m[14]&m[99]&m[100]&m[336]&m[337])|(m[14]&m[99]&m[100]&m[336]&m[337]));
    m[43] = (((m[15]&m[102]&~m[103]&~m[350]&~m[351])|(m[15]&~m[102]&m[103]&~m[350]&~m[351])|(~m[15]&m[102]&m[103]&~m[350]&~m[351])|(m[15]&~m[102]&~m[103]&m[350]&~m[351])|(~m[15]&m[102]&~m[103]&m[350]&~m[351])|(~m[15]&~m[102]&m[103]&m[350]&~m[351])|(m[15]&~m[102]&~m[103]&~m[350]&m[351])|(~m[15]&m[102]&~m[103]&~m[350]&m[351])|(~m[15]&~m[102]&m[103]&~m[350]&m[351])|(~m[15]&~m[102]&~m[103]&m[350]&m[351]))&BiasedRNG[267])|(((m[15]&m[102]&m[103]&~m[350]&~m[351])|(m[15]&m[102]&~m[103]&m[350]&~m[351])|(m[15]&~m[102]&m[103]&m[350]&~m[351])|(~m[15]&m[102]&m[103]&m[350]&~m[351])|(m[15]&m[102]&~m[103]&~m[350]&m[351])|(m[15]&~m[102]&m[103]&~m[350]&m[351])|(~m[15]&m[102]&m[103]&~m[350]&m[351])|(m[15]&~m[102]&~m[103]&m[350]&m[351])|(~m[15]&m[102]&~m[103]&m[350]&m[351])|(~m[15]&~m[102]&m[103]&m[350]&m[351]))&~BiasedRNG[267])|((m[15]&m[102]&m[103]&m[350]&~m[351])|(m[15]&m[102]&m[103]&~m[350]&m[351])|(m[15]&m[102]&~m[103]&m[350]&m[351])|(m[15]&~m[102]&m[103]&m[350]&m[351])|(~m[15]&m[102]&m[103]&m[350]&m[351])|(m[15]&m[102]&m[103]&m[350]&m[351]));
    m[44] = (((m[16]&m[105]&~m[106]&~m[364]&~m[365])|(m[16]&~m[105]&m[106]&~m[364]&~m[365])|(~m[16]&m[105]&m[106]&~m[364]&~m[365])|(m[16]&~m[105]&~m[106]&m[364]&~m[365])|(~m[16]&m[105]&~m[106]&m[364]&~m[365])|(~m[16]&~m[105]&m[106]&m[364]&~m[365])|(m[16]&~m[105]&~m[106]&~m[364]&m[365])|(~m[16]&m[105]&~m[106]&~m[364]&m[365])|(~m[16]&~m[105]&m[106]&~m[364]&m[365])|(~m[16]&~m[105]&~m[106]&m[364]&m[365]))&BiasedRNG[268])|(((m[16]&m[105]&m[106]&~m[364]&~m[365])|(m[16]&m[105]&~m[106]&m[364]&~m[365])|(m[16]&~m[105]&m[106]&m[364]&~m[365])|(~m[16]&m[105]&m[106]&m[364]&~m[365])|(m[16]&m[105]&~m[106]&~m[364]&m[365])|(m[16]&~m[105]&m[106]&~m[364]&m[365])|(~m[16]&m[105]&m[106]&~m[364]&m[365])|(m[16]&~m[105]&~m[106]&m[364]&m[365])|(~m[16]&m[105]&~m[106]&m[364]&m[365])|(~m[16]&~m[105]&m[106]&m[364]&m[365]))&~BiasedRNG[268])|((m[16]&m[105]&m[106]&m[364]&~m[365])|(m[16]&m[105]&m[106]&~m[364]&m[365])|(m[16]&m[105]&~m[106]&m[364]&m[365])|(m[16]&~m[105]&m[106]&m[364]&m[365])|(~m[16]&m[105]&m[106]&m[364]&m[365])|(m[16]&m[105]&m[106]&m[364]&m[365]));
    m[45] = (((m[17]&m[108]&~m[109]&~m[378]&~m[379])|(m[17]&~m[108]&m[109]&~m[378]&~m[379])|(~m[17]&m[108]&m[109]&~m[378]&~m[379])|(m[17]&~m[108]&~m[109]&m[378]&~m[379])|(~m[17]&m[108]&~m[109]&m[378]&~m[379])|(~m[17]&~m[108]&m[109]&m[378]&~m[379])|(m[17]&~m[108]&~m[109]&~m[378]&m[379])|(~m[17]&m[108]&~m[109]&~m[378]&m[379])|(~m[17]&~m[108]&m[109]&~m[378]&m[379])|(~m[17]&~m[108]&~m[109]&m[378]&m[379]))&BiasedRNG[269])|(((m[17]&m[108]&m[109]&~m[378]&~m[379])|(m[17]&m[108]&~m[109]&m[378]&~m[379])|(m[17]&~m[108]&m[109]&m[378]&~m[379])|(~m[17]&m[108]&m[109]&m[378]&~m[379])|(m[17]&m[108]&~m[109]&~m[378]&m[379])|(m[17]&~m[108]&m[109]&~m[378]&m[379])|(~m[17]&m[108]&m[109]&~m[378]&m[379])|(m[17]&~m[108]&~m[109]&m[378]&m[379])|(~m[17]&m[108]&~m[109]&m[378]&m[379])|(~m[17]&~m[108]&m[109]&m[378]&m[379]))&~BiasedRNG[269])|((m[17]&m[108]&m[109]&m[378]&~m[379])|(m[17]&m[108]&m[109]&~m[378]&m[379])|(m[17]&m[108]&~m[109]&m[378]&m[379])|(m[17]&~m[108]&m[109]&m[378]&m[379])|(~m[17]&m[108]&m[109]&m[378]&m[379])|(m[17]&m[108]&m[109]&m[378]&m[379]));
    m[46] = (((m[18]&m[111]&~m[112]&~m[392]&~m[393])|(m[18]&~m[111]&m[112]&~m[392]&~m[393])|(~m[18]&m[111]&m[112]&~m[392]&~m[393])|(m[18]&~m[111]&~m[112]&m[392]&~m[393])|(~m[18]&m[111]&~m[112]&m[392]&~m[393])|(~m[18]&~m[111]&m[112]&m[392]&~m[393])|(m[18]&~m[111]&~m[112]&~m[392]&m[393])|(~m[18]&m[111]&~m[112]&~m[392]&m[393])|(~m[18]&~m[111]&m[112]&~m[392]&m[393])|(~m[18]&~m[111]&~m[112]&m[392]&m[393]))&BiasedRNG[270])|(((m[18]&m[111]&m[112]&~m[392]&~m[393])|(m[18]&m[111]&~m[112]&m[392]&~m[393])|(m[18]&~m[111]&m[112]&m[392]&~m[393])|(~m[18]&m[111]&m[112]&m[392]&~m[393])|(m[18]&m[111]&~m[112]&~m[392]&m[393])|(m[18]&~m[111]&m[112]&~m[392]&m[393])|(~m[18]&m[111]&m[112]&~m[392]&m[393])|(m[18]&~m[111]&~m[112]&m[392]&m[393])|(~m[18]&m[111]&~m[112]&m[392]&m[393])|(~m[18]&~m[111]&m[112]&m[392]&m[393]))&~BiasedRNG[270])|((m[18]&m[111]&m[112]&m[392]&~m[393])|(m[18]&m[111]&m[112]&~m[392]&m[393])|(m[18]&m[111]&~m[112]&m[392]&m[393])|(m[18]&~m[111]&m[112]&m[392]&m[393])|(~m[18]&m[111]&m[112]&m[392]&m[393])|(m[18]&m[111]&m[112]&m[392]&m[393]));
    m[47] = (((m[19]&m[114]&~m[115]&~m[406]&~m[407])|(m[19]&~m[114]&m[115]&~m[406]&~m[407])|(~m[19]&m[114]&m[115]&~m[406]&~m[407])|(m[19]&~m[114]&~m[115]&m[406]&~m[407])|(~m[19]&m[114]&~m[115]&m[406]&~m[407])|(~m[19]&~m[114]&m[115]&m[406]&~m[407])|(m[19]&~m[114]&~m[115]&~m[406]&m[407])|(~m[19]&m[114]&~m[115]&~m[406]&m[407])|(~m[19]&~m[114]&m[115]&~m[406]&m[407])|(~m[19]&~m[114]&~m[115]&m[406]&m[407]))&BiasedRNG[271])|(((m[19]&m[114]&m[115]&~m[406]&~m[407])|(m[19]&m[114]&~m[115]&m[406]&~m[407])|(m[19]&~m[114]&m[115]&m[406]&~m[407])|(~m[19]&m[114]&m[115]&m[406]&~m[407])|(m[19]&m[114]&~m[115]&~m[406]&m[407])|(m[19]&~m[114]&m[115]&~m[406]&m[407])|(~m[19]&m[114]&m[115]&~m[406]&m[407])|(m[19]&~m[114]&~m[115]&m[406]&m[407])|(~m[19]&m[114]&~m[115]&m[406]&m[407])|(~m[19]&~m[114]&m[115]&m[406]&m[407]))&~BiasedRNG[271])|((m[19]&m[114]&m[115]&m[406]&~m[407])|(m[19]&m[114]&m[115]&~m[406]&m[407])|(m[19]&m[114]&~m[115]&m[406]&m[407])|(m[19]&~m[114]&m[115]&m[406]&m[407])|(~m[19]&m[114]&m[115]&m[406]&m[407])|(m[19]&m[114]&m[115]&m[406]&m[407]));
    m[48] = (((m[20]&m[117]&~m[118]&~m[420]&~m[421])|(m[20]&~m[117]&m[118]&~m[420]&~m[421])|(~m[20]&m[117]&m[118]&~m[420]&~m[421])|(m[20]&~m[117]&~m[118]&m[420]&~m[421])|(~m[20]&m[117]&~m[118]&m[420]&~m[421])|(~m[20]&~m[117]&m[118]&m[420]&~m[421])|(m[20]&~m[117]&~m[118]&~m[420]&m[421])|(~m[20]&m[117]&~m[118]&~m[420]&m[421])|(~m[20]&~m[117]&m[118]&~m[420]&m[421])|(~m[20]&~m[117]&~m[118]&m[420]&m[421]))&BiasedRNG[272])|(((m[20]&m[117]&m[118]&~m[420]&~m[421])|(m[20]&m[117]&~m[118]&m[420]&~m[421])|(m[20]&~m[117]&m[118]&m[420]&~m[421])|(~m[20]&m[117]&m[118]&m[420]&~m[421])|(m[20]&m[117]&~m[118]&~m[420]&m[421])|(m[20]&~m[117]&m[118]&~m[420]&m[421])|(~m[20]&m[117]&m[118]&~m[420]&m[421])|(m[20]&~m[117]&~m[118]&m[420]&m[421])|(~m[20]&m[117]&~m[118]&m[420]&m[421])|(~m[20]&~m[117]&m[118]&m[420]&m[421]))&~BiasedRNG[272])|((m[20]&m[117]&m[118]&m[420]&~m[421])|(m[20]&m[117]&m[118]&~m[420]&m[421])|(m[20]&m[117]&~m[118]&m[420]&m[421])|(m[20]&~m[117]&m[118]&m[420]&m[421])|(~m[20]&m[117]&m[118]&m[420]&m[421])|(m[20]&m[117]&m[118]&m[420]&m[421]));
    m[49] = (((m[21]&m[120]&~m[121]&~m[434]&~m[435])|(m[21]&~m[120]&m[121]&~m[434]&~m[435])|(~m[21]&m[120]&m[121]&~m[434]&~m[435])|(m[21]&~m[120]&~m[121]&m[434]&~m[435])|(~m[21]&m[120]&~m[121]&m[434]&~m[435])|(~m[21]&~m[120]&m[121]&m[434]&~m[435])|(m[21]&~m[120]&~m[121]&~m[434]&m[435])|(~m[21]&m[120]&~m[121]&~m[434]&m[435])|(~m[21]&~m[120]&m[121]&~m[434]&m[435])|(~m[21]&~m[120]&~m[121]&m[434]&m[435]))&BiasedRNG[273])|(((m[21]&m[120]&m[121]&~m[434]&~m[435])|(m[21]&m[120]&~m[121]&m[434]&~m[435])|(m[21]&~m[120]&m[121]&m[434]&~m[435])|(~m[21]&m[120]&m[121]&m[434]&~m[435])|(m[21]&m[120]&~m[121]&~m[434]&m[435])|(m[21]&~m[120]&m[121]&~m[434]&m[435])|(~m[21]&m[120]&m[121]&~m[434]&m[435])|(m[21]&~m[120]&~m[121]&m[434]&m[435])|(~m[21]&m[120]&~m[121]&m[434]&m[435])|(~m[21]&~m[120]&m[121]&m[434]&m[435]))&~BiasedRNG[273])|((m[21]&m[120]&m[121]&m[434]&~m[435])|(m[21]&m[120]&m[121]&~m[434]&m[435])|(m[21]&m[120]&~m[121]&m[434]&m[435])|(m[21]&~m[120]&m[121]&m[434]&m[435])|(~m[21]&m[120]&m[121]&m[434]&m[435])|(m[21]&m[120]&m[121]&m[434]&m[435]));
    m[50] = (((m[22]&m[123]&~m[124]&~m[448]&~m[449])|(m[22]&~m[123]&m[124]&~m[448]&~m[449])|(~m[22]&m[123]&m[124]&~m[448]&~m[449])|(m[22]&~m[123]&~m[124]&m[448]&~m[449])|(~m[22]&m[123]&~m[124]&m[448]&~m[449])|(~m[22]&~m[123]&m[124]&m[448]&~m[449])|(m[22]&~m[123]&~m[124]&~m[448]&m[449])|(~m[22]&m[123]&~m[124]&~m[448]&m[449])|(~m[22]&~m[123]&m[124]&~m[448]&m[449])|(~m[22]&~m[123]&~m[124]&m[448]&m[449]))&BiasedRNG[274])|(((m[22]&m[123]&m[124]&~m[448]&~m[449])|(m[22]&m[123]&~m[124]&m[448]&~m[449])|(m[22]&~m[123]&m[124]&m[448]&~m[449])|(~m[22]&m[123]&m[124]&m[448]&~m[449])|(m[22]&m[123]&~m[124]&~m[448]&m[449])|(m[22]&~m[123]&m[124]&~m[448]&m[449])|(~m[22]&m[123]&m[124]&~m[448]&m[449])|(m[22]&~m[123]&~m[124]&m[448]&m[449])|(~m[22]&m[123]&~m[124]&m[448]&m[449])|(~m[22]&~m[123]&m[124]&m[448]&m[449]))&~BiasedRNG[274])|((m[22]&m[123]&m[124]&m[448]&~m[449])|(m[22]&m[123]&m[124]&~m[448]&m[449])|(m[22]&m[123]&~m[124]&m[448]&m[449])|(m[22]&~m[123]&m[124]&m[448]&m[449])|(~m[22]&m[123]&m[124]&m[448]&m[449])|(m[22]&m[123]&m[124]&m[448]&m[449]));
    m[51] = (((m[23]&m[126]&~m[127]&~m[462]&~m[463])|(m[23]&~m[126]&m[127]&~m[462]&~m[463])|(~m[23]&m[126]&m[127]&~m[462]&~m[463])|(m[23]&~m[126]&~m[127]&m[462]&~m[463])|(~m[23]&m[126]&~m[127]&m[462]&~m[463])|(~m[23]&~m[126]&m[127]&m[462]&~m[463])|(m[23]&~m[126]&~m[127]&~m[462]&m[463])|(~m[23]&m[126]&~m[127]&~m[462]&m[463])|(~m[23]&~m[126]&m[127]&~m[462]&m[463])|(~m[23]&~m[126]&~m[127]&m[462]&m[463]))&BiasedRNG[275])|(((m[23]&m[126]&m[127]&~m[462]&~m[463])|(m[23]&m[126]&~m[127]&m[462]&~m[463])|(m[23]&~m[126]&m[127]&m[462]&~m[463])|(~m[23]&m[126]&m[127]&m[462]&~m[463])|(m[23]&m[126]&~m[127]&~m[462]&m[463])|(m[23]&~m[126]&m[127]&~m[462]&m[463])|(~m[23]&m[126]&m[127]&~m[462]&m[463])|(m[23]&~m[126]&~m[127]&m[462]&m[463])|(~m[23]&m[126]&~m[127]&m[462]&m[463])|(~m[23]&~m[126]&m[127]&m[462]&m[463]))&~BiasedRNG[275])|((m[23]&m[126]&m[127]&m[462]&~m[463])|(m[23]&m[126]&m[127]&~m[462]&m[463])|(m[23]&m[126]&~m[127]&m[462]&m[463])|(m[23]&~m[126]&m[127]&m[462]&m[463])|(~m[23]&m[126]&m[127]&m[462]&m[463])|(m[23]&m[126]&m[127]&m[462]&m[463]));
    m[52] = (((m[24]&m[129]&~m[130]&~m[476]&~m[477])|(m[24]&~m[129]&m[130]&~m[476]&~m[477])|(~m[24]&m[129]&m[130]&~m[476]&~m[477])|(m[24]&~m[129]&~m[130]&m[476]&~m[477])|(~m[24]&m[129]&~m[130]&m[476]&~m[477])|(~m[24]&~m[129]&m[130]&m[476]&~m[477])|(m[24]&~m[129]&~m[130]&~m[476]&m[477])|(~m[24]&m[129]&~m[130]&~m[476]&m[477])|(~m[24]&~m[129]&m[130]&~m[476]&m[477])|(~m[24]&~m[129]&~m[130]&m[476]&m[477]))&BiasedRNG[276])|(((m[24]&m[129]&m[130]&~m[476]&~m[477])|(m[24]&m[129]&~m[130]&m[476]&~m[477])|(m[24]&~m[129]&m[130]&m[476]&~m[477])|(~m[24]&m[129]&m[130]&m[476]&~m[477])|(m[24]&m[129]&~m[130]&~m[476]&m[477])|(m[24]&~m[129]&m[130]&~m[476]&m[477])|(~m[24]&m[129]&m[130]&~m[476]&m[477])|(m[24]&~m[129]&~m[130]&m[476]&m[477])|(~m[24]&m[129]&~m[130]&m[476]&m[477])|(~m[24]&~m[129]&m[130]&m[476]&m[477]))&~BiasedRNG[276])|((m[24]&m[129]&m[130]&m[476]&~m[477])|(m[24]&m[129]&m[130]&~m[476]&m[477])|(m[24]&m[129]&~m[130]&m[476]&m[477])|(m[24]&~m[129]&m[130]&m[476]&m[477])|(~m[24]&m[129]&m[130]&m[476]&m[477])|(m[24]&m[129]&m[130]&m[476]&m[477]));
    m[53] = (((m[25]&m[132]&~m[133]&~m[490]&~m[491])|(m[25]&~m[132]&m[133]&~m[490]&~m[491])|(~m[25]&m[132]&m[133]&~m[490]&~m[491])|(m[25]&~m[132]&~m[133]&m[490]&~m[491])|(~m[25]&m[132]&~m[133]&m[490]&~m[491])|(~m[25]&~m[132]&m[133]&m[490]&~m[491])|(m[25]&~m[132]&~m[133]&~m[490]&m[491])|(~m[25]&m[132]&~m[133]&~m[490]&m[491])|(~m[25]&~m[132]&m[133]&~m[490]&m[491])|(~m[25]&~m[132]&~m[133]&m[490]&m[491]))&BiasedRNG[277])|(((m[25]&m[132]&m[133]&~m[490]&~m[491])|(m[25]&m[132]&~m[133]&m[490]&~m[491])|(m[25]&~m[132]&m[133]&m[490]&~m[491])|(~m[25]&m[132]&m[133]&m[490]&~m[491])|(m[25]&m[132]&~m[133]&~m[490]&m[491])|(m[25]&~m[132]&m[133]&~m[490]&m[491])|(~m[25]&m[132]&m[133]&~m[490]&m[491])|(m[25]&~m[132]&~m[133]&m[490]&m[491])|(~m[25]&m[132]&~m[133]&m[490]&m[491])|(~m[25]&~m[132]&m[133]&m[490]&m[491]))&~BiasedRNG[277])|((m[25]&m[132]&m[133]&m[490]&~m[491])|(m[25]&m[132]&m[133]&~m[490]&m[491])|(m[25]&m[132]&~m[133]&m[490]&m[491])|(m[25]&~m[132]&m[133]&m[490]&m[491])|(~m[25]&m[132]&m[133]&m[490]&m[491])|(m[25]&m[132]&m[133]&m[490]&m[491]));
    m[54] = (((m[26]&m[135]&~m[136]&~m[504]&~m[505])|(m[26]&~m[135]&m[136]&~m[504]&~m[505])|(~m[26]&m[135]&m[136]&~m[504]&~m[505])|(m[26]&~m[135]&~m[136]&m[504]&~m[505])|(~m[26]&m[135]&~m[136]&m[504]&~m[505])|(~m[26]&~m[135]&m[136]&m[504]&~m[505])|(m[26]&~m[135]&~m[136]&~m[504]&m[505])|(~m[26]&m[135]&~m[136]&~m[504]&m[505])|(~m[26]&~m[135]&m[136]&~m[504]&m[505])|(~m[26]&~m[135]&~m[136]&m[504]&m[505]))&BiasedRNG[278])|(((m[26]&m[135]&m[136]&~m[504]&~m[505])|(m[26]&m[135]&~m[136]&m[504]&~m[505])|(m[26]&~m[135]&m[136]&m[504]&~m[505])|(~m[26]&m[135]&m[136]&m[504]&~m[505])|(m[26]&m[135]&~m[136]&~m[504]&m[505])|(m[26]&~m[135]&m[136]&~m[504]&m[505])|(~m[26]&m[135]&m[136]&~m[504]&m[505])|(m[26]&~m[135]&~m[136]&m[504]&m[505])|(~m[26]&m[135]&~m[136]&m[504]&m[505])|(~m[26]&~m[135]&m[136]&m[504]&m[505]))&~BiasedRNG[278])|((m[26]&m[135]&m[136]&m[504]&~m[505])|(m[26]&m[135]&m[136]&~m[504]&m[505])|(m[26]&m[135]&~m[136]&m[504]&m[505])|(m[26]&~m[135]&m[136]&m[504]&m[505])|(~m[26]&m[135]&m[136]&m[504]&m[505])|(m[26]&m[135]&m[136]&m[504]&m[505]));
    m[55] = (((m[27]&m[138]&~m[139]&~m[518]&~m[519])|(m[27]&~m[138]&m[139]&~m[518]&~m[519])|(~m[27]&m[138]&m[139]&~m[518]&~m[519])|(m[27]&~m[138]&~m[139]&m[518]&~m[519])|(~m[27]&m[138]&~m[139]&m[518]&~m[519])|(~m[27]&~m[138]&m[139]&m[518]&~m[519])|(m[27]&~m[138]&~m[139]&~m[518]&m[519])|(~m[27]&m[138]&~m[139]&~m[518]&m[519])|(~m[27]&~m[138]&m[139]&~m[518]&m[519])|(~m[27]&~m[138]&~m[139]&m[518]&m[519]))&BiasedRNG[279])|(((m[27]&m[138]&m[139]&~m[518]&~m[519])|(m[27]&m[138]&~m[139]&m[518]&~m[519])|(m[27]&~m[138]&m[139]&m[518]&~m[519])|(~m[27]&m[138]&m[139]&m[518]&~m[519])|(m[27]&m[138]&~m[139]&~m[518]&m[519])|(m[27]&~m[138]&m[139]&~m[518]&m[519])|(~m[27]&m[138]&m[139]&~m[518]&m[519])|(m[27]&~m[138]&~m[139]&m[518]&m[519])|(~m[27]&m[138]&~m[139]&m[518]&m[519])|(~m[27]&~m[138]&m[139]&m[518]&m[519]))&~BiasedRNG[279])|((m[27]&m[138]&m[139]&m[518]&~m[519])|(m[27]&m[138]&m[139]&~m[518]&m[519])|(m[27]&m[138]&~m[139]&m[518]&m[519])|(m[27]&~m[138]&m[139]&m[518]&m[519])|(~m[27]&m[138]&m[139]&m[518]&m[519])|(m[27]&m[138]&m[139]&m[518]&m[519]));
    m[56] = (((m[0]&m[142]&~m[143]&~m[144]&~m[145])|(m[0]&~m[142]&m[143]&~m[144]&~m[145])|(~m[0]&m[142]&m[143]&~m[144]&~m[145])|(m[0]&~m[142]&~m[143]&m[144]&~m[145])|(~m[0]&m[142]&~m[143]&m[144]&~m[145])|(~m[0]&~m[142]&m[143]&m[144]&~m[145])|(m[0]&~m[142]&~m[143]&~m[144]&m[145])|(~m[0]&m[142]&~m[143]&~m[144]&m[145])|(~m[0]&~m[142]&m[143]&~m[144]&m[145])|(~m[0]&~m[142]&~m[143]&m[144]&m[145]))&BiasedRNG[280])|(((m[0]&m[142]&m[143]&~m[144]&~m[145])|(m[0]&m[142]&~m[143]&m[144]&~m[145])|(m[0]&~m[142]&m[143]&m[144]&~m[145])|(~m[0]&m[142]&m[143]&m[144]&~m[145])|(m[0]&m[142]&~m[143]&~m[144]&m[145])|(m[0]&~m[142]&m[143]&~m[144]&m[145])|(~m[0]&m[142]&m[143]&~m[144]&m[145])|(m[0]&~m[142]&~m[143]&m[144]&m[145])|(~m[0]&m[142]&~m[143]&m[144]&m[145])|(~m[0]&~m[142]&m[143]&m[144]&m[145]))&~BiasedRNG[280])|((m[0]&m[142]&m[143]&m[144]&~m[145])|(m[0]&m[142]&m[143]&~m[144]&m[145])|(m[0]&m[142]&~m[143]&m[144]&m[145])|(m[0]&~m[142]&m[143]&m[144]&m[145])|(~m[0]&m[142]&m[143]&m[144]&m[145])|(m[0]&m[142]&m[143]&m[144]&m[145]));
    m[59] = (((m[1]&m[156]&~m[157]&~m[158]&~m[159])|(m[1]&~m[156]&m[157]&~m[158]&~m[159])|(~m[1]&m[156]&m[157]&~m[158]&~m[159])|(m[1]&~m[156]&~m[157]&m[158]&~m[159])|(~m[1]&m[156]&~m[157]&m[158]&~m[159])|(~m[1]&~m[156]&m[157]&m[158]&~m[159])|(m[1]&~m[156]&~m[157]&~m[158]&m[159])|(~m[1]&m[156]&~m[157]&~m[158]&m[159])|(~m[1]&~m[156]&m[157]&~m[158]&m[159])|(~m[1]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[281])|(((m[1]&m[156]&m[157]&~m[158]&~m[159])|(m[1]&m[156]&~m[157]&m[158]&~m[159])|(m[1]&~m[156]&m[157]&m[158]&~m[159])|(~m[1]&m[156]&m[157]&m[158]&~m[159])|(m[1]&m[156]&~m[157]&~m[158]&m[159])|(m[1]&~m[156]&m[157]&~m[158]&m[159])|(~m[1]&m[156]&m[157]&~m[158]&m[159])|(m[1]&~m[156]&~m[157]&m[158]&m[159])|(~m[1]&m[156]&~m[157]&m[158]&m[159])|(~m[1]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[281])|((m[1]&m[156]&m[157]&m[158]&~m[159])|(m[1]&m[156]&m[157]&~m[158]&m[159])|(m[1]&m[156]&~m[157]&m[158]&m[159])|(m[1]&~m[156]&m[157]&m[158]&m[159])|(~m[1]&m[156]&m[157]&m[158]&m[159])|(m[1]&m[156]&m[157]&m[158]&m[159]));
    m[62] = (((m[2]&m[170]&~m[171]&~m[172]&~m[173])|(m[2]&~m[170]&m[171]&~m[172]&~m[173])|(~m[2]&m[170]&m[171]&~m[172]&~m[173])|(m[2]&~m[170]&~m[171]&m[172]&~m[173])|(~m[2]&m[170]&~m[171]&m[172]&~m[173])|(~m[2]&~m[170]&m[171]&m[172]&~m[173])|(m[2]&~m[170]&~m[171]&~m[172]&m[173])|(~m[2]&m[170]&~m[171]&~m[172]&m[173])|(~m[2]&~m[170]&m[171]&~m[172]&m[173])|(~m[2]&~m[170]&~m[171]&m[172]&m[173]))&BiasedRNG[282])|(((m[2]&m[170]&m[171]&~m[172]&~m[173])|(m[2]&m[170]&~m[171]&m[172]&~m[173])|(m[2]&~m[170]&m[171]&m[172]&~m[173])|(~m[2]&m[170]&m[171]&m[172]&~m[173])|(m[2]&m[170]&~m[171]&~m[172]&m[173])|(m[2]&~m[170]&m[171]&~m[172]&m[173])|(~m[2]&m[170]&m[171]&~m[172]&m[173])|(m[2]&~m[170]&~m[171]&m[172]&m[173])|(~m[2]&m[170]&~m[171]&m[172]&m[173])|(~m[2]&~m[170]&m[171]&m[172]&m[173]))&~BiasedRNG[282])|((m[2]&m[170]&m[171]&m[172]&~m[173])|(m[2]&m[170]&m[171]&~m[172]&m[173])|(m[2]&m[170]&~m[171]&m[172]&m[173])|(m[2]&~m[170]&m[171]&m[172]&m[173])|(~m[2]&m[170]&m[171]&m[172]&m[173])|(m[2]&m[170]&m[171]&m[172]&m[173]));
    m[65] = (((m[3]&m[184]&~m[185]&~m[186]&~m[187])|(m[3]&~m[184]&m[185]&~m[186]&~m[187])|(~m[3]&m[184]&m[185]&~m[186]&~m[187])|(m[3]&~m[184]&~m[185]&m[186]&~m[187])|(~m[3]&m[184]&~m[185]&m[186]&~m[187])|(~m[3]&~m[184]&m[185]&m[186]&~m[187])|(m[3]&~m[184]&~m[185]&~m[186]&m[187])|(~m[3]&m[184]&~m[185]&~m[186]&m[187])|(~m[3]&~m[184]&m[185]&~m[186]&m[187])|(~m[3]&~m[184]&~m[185]&m[186]&m[187]))&BiasedRNG[283])|(((m[3]&m[184]&m[185]&~m[186]&~m[187])|(m[3]&m[184]&~m[185]&m[186]&~m[187])|(m[3]&~m[184]&m[185]&m[186]&~m[187])|(~m[3]&m[184]&m[185]&m[186]&~m[187])|(m[3]&m[184]&~m[185]&~m[186]&m[187])|(m[3]&~m[184]&m[185]&~m[186]&m[187])|(~m[3]&m[184]&m[185]&~m[186]&m[187])|(m[3]&~m[184]&~m[185]&m[186]&m[187])|(~m[3]&m[184]&~m[185]&m[186]&m[187])|(~m[3]&~m[184]&m[185]&m[186]&m[187]))&~BiasedRNG[283])|((m[3]&m[184]&m[185]&m[186]&~m[187])|(m[3]&m[184]&m[185]&~m[186]&m[187])|(m[3]&m[184]&~m[185]&m[186]&m[187])|(m[3]&~m[184]&m[185]&m[186]&m[187])|(~m[3]&m[184]&m[185]&m[186]&m[187])|(m[3]&m[184]&m[185]&m[186]&m[187]));
    m[68] = (((m[4]&m[198]&~m[199]&~m[200]&~m[201])|(m[4]&~m[198]&m[199]&~m[200]&~m[201])|(~m[4]&m[198]&m[199]&~m[200]&~m[201])|(m[4]&~m[198]&~m[199]&m[200]&~m[201])|(~m[4]&m[198]&~m[199]&m[200]&~m[201])|(~m[4]&~m[198]&m[199]&m[200]&~m[201])|(m[4]&~m[198]&~m[199]&~m[200]&m[201])|(~m[4]&m[198]&~m[199]&~m[200]&m[201])|(~m[4]&~m[198]&m[199]&~m[200]&m[201])|(~m[4]&~m[198]&~m[199]&m[200]&m[201]))&BiasedRNG[284])|(((m[4]&m[198]&m[199]&~m[200]&~m[201])|(m[4]&m[198]&~m[199]&m[200]&~m[201])|(m[4]&~m[198]&m[199]&m[200]&~m[201])|(~m[4]&m[198]&m[199]&m[200]&~m[201])|(m[4]&m[198]&~m[199]&~m[200]&m[201])|(m[4]&~m[198]&m[199]&~m[200]&m[201])|(~m[4]&m[198]&m[199]&~m[200]&m[201])|(m[4]&~m[198]&~m[199]&m[200]&m[201])|(~m[4]&m[198]&~m[199]&m[200]&m[201])|(~m[4]&~m[198]&m[199]&m[200]&m[201]))&~BiasedRNG[284])|((m[4]&m[198]&m[199]&m[200]&~m[201])|(m[4]&m[198]&m[199]&~m[200]&m[201])|(m[4]&m[198]&~m[199]&m[200]&m[201])|(m[4]&~m[198]&m[199]&m[200]&m[201])|(~m[4]&m[198]&m[199]&m[200]&m[201])|(m[4]&m[198]&m[199]&m[200]&m[201]));
    m[71] = (((m[5]&m[212]&~m[213]&~m[214]&~m[215])|(m[5]&~m[212]&m[213]&~m[214]&~m[215])|(~m[5]&m[212]&m[213]&~m[214]&~m[215])|(m[5]&~m[212]&~m[213]&m[214]&~m[215])|(~m[5]&m[212]&~m[213]&m[214]&~m[215])|(~m[5]&~m[212]&m[213]&m[214]&~m[215])|(m[5]&~m[212]&~m[213]&~m[214]&m[215])|(~m[5]&m[212]&~m[213]&~m[214]&m[215])|(~m[5]&~m[212]&m[213]&~m[214]&m[215])|(~m[5]&~m[212]&~m[213]&m[214]&m[215]))&BiasedRNG[285])|(((m[5]&m[212]&m[213]&~m[214]&~m[215])|(m[5]&m[212]&~m[213]&m[214]&~m[215])|(m[5]&~m[212]&m[213]&m[214]&~m[215])|(~m[5]&m[212]&m[213]&m[214]&~m[215])|(m[5]&m[212]&~m[213]&~m[214]&m[215])|(m[5]&~m[212]&m[213]&~m[214]&m[215])|(~m[5]&m[212]&m[213]&~m[214]&m[215])|(m[5]&~m[212]&~m[213]&m[214]&m[215])|(~m[5]&m[212]&~m[213]&m[214]&m[215])|(~m[5]&~m[212]&m[213]&m[214]&m[215]))&~BiasedRNG[285])|((m[5]&m[212]&m[213]&m[214]&~m[215])|(m[5]&m[212]&m[213]&~m[214]&m[215])|(m[5]&m[212]&~m[213]&m[214]&m[215])|(m[5]&~m[212]&m[213]&m[214]&m[215])|(~m[5]&m[212]&m[213]&m[214]&m[215])|(m[5]&m[212]&m[213]&m[214]&m[215]));
    m[74] = (((m[6]&m[226]&~m[227]&~m[228]&~m[229])|(m[6]&~m[226]&m[227]&~m[228]&~m[229])|(~m[6]&m[226]&m[227]&~m[228]&~m[229])|(m[6]&~m[226]&~m[227]&m[228]&~m[229])|(~m[6]&m[226]&~m[227]&m[228]&~m[229])|(~m[6]&~m[226]&m[227]&m[228]&~m[229])|(m[6]&~m[226]&~m[227]&~m[228]&m[229])|(~m[6]&m[226]&~m[227]&~m[228]&m[229])|(~m[6]&~m[226]&m[227]&~m[228]&m[229])|(~m[6]&~m[226]&~m[227]&m[228]&m[229]))&BiasedRNG[286])|(((m[6]&m[226]&m[227]&~m[228]&~m[229])|(m[6]&m[226]&~m[227]&m[228]&~m[229])|(m[6]&~m[226]&m[227]&m[228]&~m[229])|(~m[6]&m[226]&m[227]&m[228]&~m[229])|(m[6]&m[226]&~m[227]&~m[228]&m[229])|(m[6]&~m[226]&m[227]&~m[228]&m[229])|(~m[6]&m[226]&m[227]&~m[228]&m[229])|(m[6]&~m[226]&~m[227]&m[228]&m[229])|(~m[6]&m[226]&~m[227]&m[228]&m[229])|(~m[6]&~m[226]&m[227]&m[228]&m[229]))&~BiasedRNG[286])|((m[6]&m[226]&m[227]&m[228]&~m[229])|(m[6]&m[226]&m[227]&~m[228]&m[229])|(m[6]&m[226]&~m[227]&m[228]&m[229])|(m[6]&~m[226]&m[227]&m[228]&m[229])|(~m[6]&m[226]&m[227]&m[228]&m[229])|(m[6]&m[226]&m[227]&m[228]&m[229]));
    m[77] = (((m[7]&m[240]&~m[241]&~m[242]&~m[243])|(m[7]&~m[240]&m[241]&~m[242]&~m[243])|(~m[7]&m[240]&m[241]&~m[242]&~m[243])|(m[7]&~m[240]&~m[241]&m[242]&~m[243])|(~m[7]&m[240]&~m[241]&m[242]&~m[243])|(~m[7]&~m[240]&m[241]&m[242]&~m[243])|(m[7]&~m[240]&~m[241]&~m[242]&m[243])|(~m[7]&m[240]&~m[241]&~m[242]&m[243])|(~m[7]&~m[240]&m[241]&~m[242]&m[243])|(~m[7]&~m[240]&~m[241]&m[242]&m[243]))&BiasedRNG[287])|(((m[7]&m[240]&m[241]&~m[242]&~m[243])|(m[7]&m[240]&~m[241]&m[242]&~m[243])|(m[7]&~m[240]&m[241]&m[242]&~m[243])|(~m[7]&m[240]&m[241]&m[242]&~m[243])|(m[7]&m[240]&~m[241]&~m[242]&m[243])|(m[7]&~m[240]&m[241]&~m[242]&m[243])|(~m[7]&m[240]&m[241]&~m[242]&m[243])|(m[7]&~m[240]&~m[241]&m[242]&m[243])|(~m[7]&m[240]&~m[241]&m[242]&m[243])|(~m[7]&~m[240]&m[241]&m[242]&m[243]))&~BiasedRNG[287])|((m[7]&m[240]&m[241]&m[242]&~m[243])|(m[7]&m[240]&m[241]&~m[242]&m[243])|(m[7]&m[240]&~m[241]&m[242]&m[243])|(m[7]&~m[240]&m[241]&m[242]&m[243])|(~m[7]&m[240]&m[241]&m[242]&m[243])|(m[7]&m[240]&m[241]&m[242]&m[243]));
    m[80] = (((m[8]&m[254]&~m[255]&~m[256]&~m[257])|(m[8]&~m[254]&m[255]&~m[256]&~m[257])|(~m[8]&m[254]&m[255]&~m[256]&~m[257])|(m[8]&~m[254]&~m[255]&m[256]&~m[257])|(~m[8]&m[254]&~m[255]&m[256]&~m[257])|(~m[8]&~m[254]&m[255]&m[256]&~m[257])|(m[8]&~m[254]&~m[255]&~m[256]&m[257])|(~m[8]&m[254]&~m[255]&~m[256]&m[257])|(~m[8]&~m[254]&m[255]&~m[256]&m[257])|(~m[8]&~m[254]&~m[255]&m[256]&m[257]))&BiasedRNG[288])|(((m[8]&m[254]&m[255]&~m[256]&~m[257])|(m[8]&m[254]&~m[255]&m[256]&~m[257])|(m[8]&~m[254]&m[255]&m[256]&~m[257])|(~m[8]&m[254]&m[255]&m[256]&~m[257])|(m[8]&m[254]&~m[255]&~m[256]&m[257])|(m[8]&~m[254]&m[255]&~m[256]&m[257])|(~m[8]&m[254]&m[255]&~m[256]&m[257])|(m[8]&~m[254]&~m[255]&m[256]&m[257])|(~m[8]&m[254]&~m[255]&m[256]&m[257])|(~m[8]&~m[254]&m[255]&m[256]&m[257]))&~BiasedRNG[288])|((m[8]&m[254]&m[255]&m[256]&~m[257])|(m[8]&m[254]&m[255]&~m[256]&m[257])|(m[8]&m[254]&~m[255]&m[256]&m[257])|(m[8]&~m[254]&m[255]&m[256]&m[257])|(~m[8]&m[254]&m[255]&m[256]&m[257])|(m[8]&m[254]&m[255]&m[256]&m[257]));
    m[83] = (((m[9]&m[268]&~m[269]&~m[270]&~m[271])|(m[9]&~m[268]&m[269]&~m[270]&~m[271])|(~m[9]&m[268]&m[269]&~m[270]&~m[271])|(m[9]&~m[268]&~m[269]&m[270]&~m[271])|(~m[9]&m[268]&~m[269]&m[270]&~m[271])|(~m[9]&~m[268]&m[269]&m[270]&~m[271])|(m[9]&~m[268]&~m[269]&~m[270]&m[271])|(~m[9]&m[268]&~m[269]&~m[270]&m[271])|(~m[9]&~m[268]&m[269]&~m[270]&m[271])|(~m[9]&~m[268]&~m[269]&m[270]&m[271]))&BiasedRNG[289])|(((m[9]&m[268]&m[269]&~m[270]&~m[271])|(m[9]&m[268]&~m[269]&m[270]&~m[271])|(m[9]&~m[268]&m[269]&m[270]&~m[271])|(~m[9]&m[268]&m[269]&m[270]&~m[271])|(m[9]&m[268]&~m[269]&~m[270]&m[271])|(m[9]&~m[268]&m[269]&~m[270]&m[271])|(~m[9]&m[268]&m[269]&~m[270]&m[271])|(m[9]&~m[268]&~m[269]&m[270]&m[271])|(~m[9]&m[268]&~m[269]&m[270]&m[271])|(~m[9]&~m[268]&m[269]&m[270]&m[271]))&~BiasedRNG[289])|((m[9]&m[268]&m[269]&m[270]&~m[271])|(m[9]&m[268]&m[269]&~m[270]&m[271])|(m[9]&m[268]&~m[269]&m[270]&m[271])|(m[9]&~m[268]&m[269]&m[270]&m[271])|(~m[9]&m[268]&m[269]&m[270]&m[271])|(m[9]&m[268]&m[269]&m[270]&m[271]));
    m[86] = (((m[10]&m[282]&~m[283]&~m[284]&~m[285])|(m[10]&~m[282]&m[283]&~m[284]&~m[285])|(~m[10]&m[282]&m[283]&~m[284]&~m[285])|(m[10]&~m[282]&~m[283]&m[284]&~m[285])|(~m[10]&m[282]&~m[283]&m[284]&~m[285])|(~m[10]&~m[282]&m[283]&m[284]&~m[285])|(m[10]&~m[282]&~m[283]&~m[284]&m[285])|(~m[10]&m[282]&~m[283]&~m[284]&m[285])|(~m[10]&~m[282]&m[283]&~m[284]&m[285])|(~m[10]&~m[282]&~m[283]&m[284]&m[285]))&BiasedRNG[290])|(((m[10]&m[282]&m[283]&~m[284]&~m[285])|(m[10]&m[282]&~m[283]&m[284]&~m[285])|(m[10]&~m[282]&m[283]&m[284]&~m[285])|(~m[10]&m[282]&m[283]&m[284]&~m[285])|(m[10]&m[282]&~m[283]&~m[284]&m[285])|(m[10]&~m[282]&m[283]&~m[284]&m[285])|(~m[10]&m[282]&m[283]&~m[284]&m[285])|(m[10]&~m[282]&~m[283]&m[284]&m[285])|(~m[10]&m[282]&~m[283]&m[284]&m[285])|(~m[10]&~m[282]&m[283]&m[284]&m[285]))&~BiasedRNG[290])|((m[10]&m[282]&m[283]&m[284]&~m[285])|(m[10]&m[282]&m[283]&~m[284]&m[285])|(m[10]&m[282]&~m[283]&m[284]&m[285])|(m[10]&~m[282]&m[283]&m[284]&m[285])|(~m[10]&m[282]&m[283]&m[284]&m[285])|(m[10]&m[282]&m[283]&m[284]&m[285]));
    m[89] = (((m[11]&m[296]&~m[297]&~m[298]&~m[299])|(m[11]&~m[296]&m[297]&~m[298]&~m[299])|(~m[11]&m[296]&m[297]&~m[298]&~m[299])|(m[11]&~m[296]&~m[297]&m[298]&~m[299])|(~m[11]&m[296]&~m[297]&m[298]&~m[299])|(~m[11]&~m[296]&m[297]&m[298]&~m[299])|(m[11]&~m[296]&~m[297]&~m[298]&m[299])|(~m[11]&m[296]&~m[297]&~m[298]&m[299])|(~m[11]&~m[296]&m[297]&~m[298]&m[299])|(~m[11]&~m[296]&~m[297]&m[298]&m[299]))&BiasedRNG[291])|(((m[11]&m[296]&m[297]&~m[298]&~m[299])|(m[11]&m[296]&~m[297]&m[298]&~m[299])|(m[11]&~m[296]&m[297]&m[298]&~m[299])|(~m[11]&m[296]&m[297]&m[298]&~m[299])|(m[11]&m[296]&~m[297]&~m[298]&m[299])|(m[11]&~m[296]&m[297]&~m[298]&m[299])|(~m[11]&m[296]&m[297]&~m[298]&m[299])|(m[11]&~m[296]&~m[297]&m[298]&m[299])|(~m[11]&m[296]&~m[297]&m[298]&m[299])|(~m[11]&~m[296]&m[297]&m[298]&m[299]))&~BiasedRNG[291])|((m[11]&m[296]&m[297]&m[298]&~m[299])|(m[11]&m[296]&m[297]&~m[298]&m[299])|(m[11]&m[296]&~m[297]&m[298]&m[299])|(m[11]&~m[296]&m[297]&m[298]&m[299])|(~m[11]&m[296]&m[297]&m[298]&m[299])|(m[11]&m[296]&m[297]&m[298]&m[299]));
    m[92] = (((m[12]&m[310]&~m[311]&~m[312]&~m[313])|(m[12]&~m[310]&m[311]&~m[312]&~m[313])|(~m[12]&m[310]&m[311]&~m[312]&~m[313])|(m[12]&~m[310]&~m[311]&m[312]&~m[313])|(~m[12]&m[310]&~m[311]&m[312]&~m[313])|(~m[12]&~m[310]&m[311]&m[312]&~m[313])|(m[12]&~m[310]&~m[311]&~m[312]&m[313])|(~m[12]&m[310]&~m[311]&~m[312]&m[313])|(~m[12]&~m[310]&m[311]&~m[312]&m[313])|(~m[12]&~m[310]&~m[311]&m[312]&m[313]))&BiasedRNG[292])|(((m[12]&m[310]&m[311]&~m[312]&~m[313])|(m[12]&m[310]&~m[311]&m[312]&~m[313])|(m[12]&~m[310]&m[311]&m[312]&~m[313])|(~m[12]&m[310]&m[311]&m[312]&~m[313])|(m[12]&m[310]&~m[311]&~m[312]&m[313])|(m[12]&~m[310]&m[311]&~m[312]&m[313])|(~m[12]&m[310]&m[311]&~m[312]&m[313])|(m[12]&~m[310]&~m[311]&m[312]&m[313])|(~m[12]&m[310]&~m[311]&m[312]&m[313])|(~m[12]&~m[310]&m[311]&m[312]&m[313]))&~BiasedRNG[292])|((m[12]&m[310]&m[311]&m[312]&~m[313])|(m[12]&m[310]&m[311]&~m[312]&m[313])|(m[12]&m[310]&~m[311]&m[312]&m[313])|(m[12]&~m[310]&m[311]&m[312]&m[313])|(~m[12]&m[310]&m[311]&m[312]&m[313])|(m[12]&m[310]&m[311]&m[312]&m[313]));
    m[95] = (((m[13]&m[324]&~m[325]&~m[326]&~m[327])|(m[13]&~m[324]&m[325]&~m[326]&~m[327])|(~m[13]&m[324]&m[325]&~m[326]&~m[327])|(m[13]&~m[324]&~m[325]&m[326]&~m[327])|(~m[13]&m[324]&~m[325]&m[326]&~m[327])|(~m[13]&~m[324]&m[325]&m[326]&~m[327])|(m[13]&~m[324]&~m[325]&~m[326]&m[327])|(~m[13]&m[324]&~m[325]&~m[326]&m[327])|(~m[13]&~m[324]&m[325]&~m[326]&m[327])|(~m[13]&~m[324]&~m[325]&m[326]&m[327]))&BiasedRNG[293])|(((m[13]&m[324]&m[325]&~m[326]&~m[327])|(m[13]&m[324]&~m[325]&m[326]&~m[327])|(m[13]&~m[324]&m[325]&m[326]&~m[327])|(~m[13]&m[324]&m[325]&m[326]&~m[327])|(m[13]&m[324]&~m[325]&~m[326]&m[327])|(m[13]&~m[324]&m[325]&~m[326]&m[327])|(~m[13]&m[324]&m[325]&~m[326]&m[327])|(m[13]&~m[324]&~m[325]&m[326]&m[327])|(~m[13]&m[324]&~m[325]&m[326]&m[327])|(~m[13]&~m[324]&m[325]&m[326]&m[327]))&~BiasedRNG[293])|((m[13]&m[324]&m[325]&m[326]&~m[327])|(m[13]&m[324]&m[325]&~m[326]&m[327])|(m[13]&m[324]&~m[325]&m[326]&m[327])|(m[13]&~m[324]&m[325]&m[326]&m[327])|(~m[13]&m[324]&m[325]&m[326]&m[327])|(m[13]&m[324]&m[325]&m[326]&m[327]));
    m[98] = (((m[14]&m[338]&~m[339]&~m[340]&~m[341])|(m[14]&~m[338]&m[339]&~m[340]&~m[341])|(~m[14]&m[338]&m[339]&~m[340]&~m[341])|(m[14]&~m[338]&~m[339]&m[340]&~m[341])|(~m[14]&m[338]&~m[339]&m[340]&~m[341])|(~m[14]&~m[338]&m[339]&m[340]&~m[341])|(m[14]&~m[338]&~m[339]&~m[340]&m[341])|(~m[14]&m[338]&~m[339]&~m[340]&m[341])|(~m[14]&~m[338]&m[339]&~m[340]&m[341])|(~m[14]&~m[338]&~m[339]&m[340]&m[341]))&BiasedRNG[294])|(((m[14]&m[338]&m[339]&~m[340]&~m[341])|(m[14]&m[338]&~m[339]&m[340]&~m[341])|(m[14]&~m[338]&m[339]&m[340]&~m[341])|(~m[14]&m[338]&m[339]&m[340]&~m[341])|(m[14]&m[338]&~m[339]&~m[340]&m[341])|(m[14]&~m[338]&m[339]&~m[340]&m[341])|(~m[14]&m[338]&m[339]&~m[340]&m[341])|(m[14]&~m[338]&~m[339]&m[340]&m[341])|(~m[14]&m[338]&~m[339]&m[340]&m[341])|(~m[14]&~m[338]&m[339]&m[340]&m[341]))&~BiasedRNG[294])|((m[14]&m[338]&m[339]&m[340]&~m[341])|(m[14]&m[338]&m[339]&~m[340]&m[341])|(m[14]&m[338]&~m[339]&m[340]&m[341])|(m[14]&~m[338]&m[339]&m[340]&m[341])|(~m[14]&m[338]&m[339]&m[340]&m[341])|(m[14]&m[338]&m[339]&m[340]&m[341]));
    m[101] = (((m[15]&m[352]&~m[353]&~m[354]&~m[355])|(m[15]&~m[352]&m[353]&~m[354]&~m[355])|(~m[15]&m[352]&m[353]&~m[354]&~m[355])|(m[15]&~m[352]&~m[353]&m[354]&~m[355])|(~m[15]&m[352]&~m[353]&m[354]&~m[355])|(~m[15]&~m[352]&m[353]&m[354]&~m[355])|(m[15]&~m[352]&~m[353]&~m[354]&m[355])|(~m[15]&m[352]&~m[353]&~m[354]&m[355])|(~m[15]&~m[352]&m[353]&~m[354]&m[355])|(~m[15]&~m[352]&~m[353]&m[354]&m[355]))&BiasedRNG[295])|(((m[15]&m[352]&m[353]&~m[354]&~m[355])|(m[15]&m[352]&~m[353]&m[354]&~m[355])|(m[15]&~m[352]&m[353]&m[354]&~m[355])|(~m[15]&m[352]&m[353]&m[354]&~m[355])|(m[15]&m[352]&~m[353]&~m[354]&m[355])|(m[15]&~m[352]&m[353]&~m[354]&m[355])|(~m[15]&m[352]&m[353]&~m[354]&m[355])|(m[15]&~m[352]&~m[353]&m[354]&m[355])|(~m[15]&m[352]&~m[353]&m[354]&m[355])|(~m[15]&~m[352]&m[353]&m[354]&m[355]))&~BiasedRNG[295])|((m[15]&m[352]&m[353]&m[354]&~m[355])|(m[15]&m[352]&m[353]&~m[354]&m[355])|(m[15]&m[352]&~m[353]&m[354]&m[355])|(m[15]&~m[352]&m[353]&m[354]&m[355])|(~m[15]&m[352]&m[353]&m[354]&m[355])|(m[15]&m[352]&m[353]&m[354]&m[355]));
    m[104] = (((m[16]&m[366]&~m[367]&~m[368]&~m[369])|(m[16]&~m[366]&m[367]&~m[368]&~m[369])|(~m[16]&m[366]&m[367]&~m[368]&~m[369])|(m[16]&~m[366]&~m[367]&m[368]&~m[369])|(~m[16]&m[366]&~m[367]&m[368]&~m[369])|(~m[16]&~m[366]&m[367]&m[368]&~m[369])|(m[16]&~m[366]&~m[367]&~m[368]&m[369])|(~m[16]&m[366]&~m[367]&~m[368]&m[369])|(~m[16]&~m[366]&m[367]&~m[368]&m[369])|(~m[16]&~m[366]&~m[367]&m[368]&m[369]))&BiasedRNG[296])|(((m[16]&m[366]&m[367]&~m[368]&~m[369])|(m[16]&m[366]&~m[367]&m[368]&~m[369])|(m[16]&~m[366]&m[367]&m[368]&~m[369])|(~m[16]&m[366]&m[367]&m[368]&~m[369])|(m[16]&m[366]&~m[367]&~m[368]&m[369])|(m[16]&~m[366]&m[367]&~m[368]&m[369])|(~m[16]&m[366]&m[367]&~m[368]&m[369])|(m[16]&~m[366]&~m[367]&m[368]&m[369])|(~m[16]&m[366]&~m[367]&m[368]&m[369])|(~m[16]&~m[366]&m[367]&m[368]&m[369]))&~BiasedRNG[296])|((m[16]&m[366]&m[367]&m[368]&~m[369])|(m[16]&m[366]&m[367]&~m[368]&m[369])|(m[16]&m[366]&~m[367]&m[368]&m[369])|(m[16]&~m[366]&m[367]&m[368]&m[369])|(~m[16]&m[366]&m[367]&m[368]&m[369])|(m[16]&m[366]&m[367]&m[368]&m[369]));
    m[107] = (((m[17]&m[380]&~m[381]&~m[382]&~m[383])|(m[17]&~m[380]&m[381]&~m[382]&~m[383])|(~m[17]&m[380]&m[381]&~m[382]&~m[383])|(m[17]&~m[380]&~m[381]&m[382]&~m[383])|(~m[17]&m[380]&~m[381]&m[382]&~m[383])|(~m[17]&~m[380]&m[381]&m[382]&~m[383])|(m[17]&~m[380]&~m[381]&~m[382]&m[383])|(~m[17]&m[380]&~m[381]&~m[382]&m[383])|(~m[17]&~m[380]&m[381]&~m[382]&m[383])|(~m[17]&~m[380]&~m[381]&m[382]&m[383]))&BiasedRNG[297])|(((m[17]&m[380]&m[381]&~m[382]&~m[383])|(m[17]&m[380]&~m[381]&m[382]&~m[383])|(m[17]&~m[380]&m[381]&m[382]&~m[383])|(~m[17]&m[380]&m[381]&m[382]&~m[383])|(m[17]&m[380]&~m[381]&~m[382]&m[383])|(m[17]&~m[380]&m[381]&~m[382]&m[383])|(~m[17]&m[380]&m[381]&~m[382]&m[383])|(m[17]&~m[380]&~m[381]&m[382]&m[383])|(~m[17]&m[380]&~m[381]&m[382]&m[383])|(~m[17]&~m[380]&m[381]&m[382]&m[383]))&~BiasedRNG[297])|((m[17]&m[380]&m[381]&m[382]&~m[383])|(m[17]&m[380]&m[381]&~m[382]&m[383])|(m[17]&m[380]&~m[381]&m[382]&m[383])|(m[17]&~m[380]&m[381]&m[382]&m[383])|(~m[17]&m[380]&m[381]&m[382]&m[383])|(m[17]&m[380]&m[381]&m[382]&m[383]));
    m[110] = (((m[18]&m[394]&~m[395]&~m[396]&~m[397])|(m[18]&~m[394]&m[395]&~m[396]&~m[397])|(~m[18]&m[394]&m[395]&~m[396]&~m[397])|(m[18]&~m[394]&~m[395]&m[396]&~m[397])|(~m[18]&m[394]&~m[395]&m[396]&~m[397])|(~m[18]&~m[394]&m[395]&m[396]&~m[397])|(m[18]&~m[394]&~m[395]&~m[396]&m[397])|(~m[18]&m[394]&~m[395]&~m[396]&m[397])|(~m[18]&~m[394]&m[395]&~m[396]&m[397])|(~m[18]&~m[394]&~m[395]&m[396]&m[397]))&BiasedRNG[298])|(((m[18]&m[394]&m[395]&~m[396]&~m[397])|(m[18]&m[394]&~m[395]&m[396]&~m[397])|(m[18]&~m[394]&m[395]&m[396]&~m[397])|(~m[18]&m[394]&m[395]&m[396]&~m[397])|(m[18]&m[394]&~m[395]&~m[396]&m[397])|(m[18]&~m[394]&m[395]&~m[396]&m[397])|(~m[18]&m[394]&m[395]&~m[396]&m[397])|(m[18]&~m[394]&~m[395]&m[396]&m[397])|(~m[18]&m[394]&~m[395]&m[396]&m[397])|(~m[18]&~m[394]&m[395]&m[396]&m[397]))&~BiasedRNG[298])|((m[18]&m[394]&m[395]&m[396]&~m[397])|(m[18]&m[394]&m[395]&~m[396]&m[397])|(m[18]&m[394]&~m[395]&m[396]&m[397])|(m[18]&~m[394]&m[395]&m[396]&m[397])|(~m[18]&m[394]&m[395]&m[396]&m[397])|(m[18]&m[394]&m[395]&m[396]&m[397]));
    m[113] = (((m[19]&m[408]&~m[409]&~m[410]&~m[411])|(m[19]&~m[408]&m[409]&~m[410]&~m[411])|(~m[19]&m[408]&m[409]&~m[410]&~m[411])|(m[19]&~m[408]&~m[409]&m[410]&~m[411])|(~m[19]&m[408]&~m[409]&m[410]&~m[411])|(~m[19]&~m[408]&m[409]&m[410]&~m[411])|(m[19]&~m[408]&~m[409]&~m[410]&m[411])|(~m[19]&m[408]&~m[409]&~m[410]&m[411])|(~m[19]&~m[408]&m[409]&~m[410]&m[411])|(~m[19]&~m[408]&~m[409]&m[410]&m[411]))&BiasedRNG[299])|(((m[19]&m[408]&m[409]&~m[410]&~m[411])|(m[19]&m[408]&~m[409]&m[410]&~m[411])|(m[19]&~m[408]&m[409]&m[410]&~m[411])|(~m[19]&m[408]&m[409]&m[410]&~m[411])|(m[19]&m[408]&~m[409]&~m[410]&m[411])|(m[19]&~m[408]&m[409]&~m[410]&m[411])|(~m[19]&m[408]&m[409]&~m[410]&m[411])|(m[19]&~m[408]&~m[409]&m[410]&m[411])|(~m[19]&m[408]&~m[409]&m[410]&m[411])|(~m[19]&~m[408]&m[409]&m[410]&m[411]))&~BiasedRNG[299])|((m[19]&m[408]&m[409]&m[410]&~m[411])|(m[19]&m[408]&m[409]&~m[410]&m[411])|(m[19]&m[408]&~m[409]&m[410]&m[411])|(m[19]&~m[408]&m[409]&m[410]&m[411])|(~m[19]&m[408]&m[409]&m[410]&m[411])|(m[19]&m[408]&m[409]&m[410]&m[411]));
    m[116] = (((m[20]&m[422]&~m[423]&~m[424]&~m[425])|(m[20]&~m[422]&m[423]&~m[424]&~m[425])|(~m[20]&m[422]&m[423]&~m[424]&~m[425])|(m[20]&~m[422]&~m[423]&m[424]&~m[425])|(~m[20]&m[422]&~m[423]&m[424]&~m[425])|(~m[20]&~m[422]&m[423]&m[424]&~m[425])|(m[20]&~m[422]&~m[423]&~m[424]&m[425])|(~m[20]&m[422]&~m[423]&~m[424]&m[425])|(~m[20]&~m[422]&m[423]&~m[424]&m[425])|(~m[20]&~m[422]&~m[423]&m[424]&m[425]))&BiasedRNG[300])|(((m[20]&m[422]&m[423]&~m[424]&~m[425])|(m[20]&m[422]&~m[423]&m[424]&~m[425])|(m[20]&~m[422]&m[423]&m[424]&~m[425])|(~m[20]&m[422]&m[423]&m[424]&~m[425])|(m[20]&m[422]&~m[423]&~m[424]&m[425])|(m[20]&~m[422]&m[423]&~m[424]&m[425])|(~m[20]&m[422]&m[423]&~m[424]&m[425])|(m[20]&~m[422]&~m[423]&m[424]&m[425])|(~m[20]&m[422]&~m[423]&m[424]&m[425])|(~m[20]&~m[422]&m[423]&m[424]&m[425]))&~BiasedRNG[300])|((m[20]&m[422]&m[423]&m[424]&~m[425])|(m[20]&m[422]&m[423]&~m[424]&m[425])|(m[20]&m[422]&~m[423]&m[424]&m[425])|(m[20]&~m[422]&m[423]&m[424]&m[425])|(~m[20]&m[422]&m[423]&m[424]&m[425])|(m[20]&m[422]&m[423]&m[424]&m[425]));
    m[119] = (((m[21]&m[436]&~m[437]&~m[438]&~m[439])|(m[21]&~m[436]&m[437]&~m[438]&~m[439])|(~m[21]&m[436]&m[437]&~m[438]&~m[439])|(m[21]&~m[436]&~m[437]&m[438]&~m[439])|(~m[21]&m[436]&~m[437]&m[438]&~m[439])|(~m[21]&~m[436]&m[437]&m[438]&~m[439])|(m[21]&~m[436]&~m[437]&~m[438]&m[439])|(~m[21]&m[436]&~m[437]&~m[438]&m[439])|(~m[21]&~m[436]&m[437]&~m[438]&m[439])|(~m[21]&~m[436]&~m[437]&m[438]&m[439]))&BiasedRNG[301])|(((m[21]&m[436]&m[437]&~m[438]&~m[439])|(m[21]&m[436]&~m[437]&m[438]&~m[439])|(m[21]&~m[436]&m[437]&m[438]&~m[439])|(~m[21]&m[436]&m[437]&m[438]&~m[439])|(m[21]&m[436]&~m[437]&~m[438]&m[439])|(m[21]&~m[436]&m[437]&~m[438]&m[439])|(~m[21]&m[436]&m[437]&~m[438]&m[439])|(m[21]&~m[436]&~m[437]&m[438]&m[439])|(~m[21]&m[436]&~m[437]&m[438]&m[439])|(~m[21]&~m[436]&m[437]&m[438]&m[439]))&~BiasedRNG[301])|((m[21]&m[436]&m[437]&m[438]&~m[439])|(m[21]&m[436]&m[437]&~m[438]&m[439])|(m[21]&m[436]&~m[437]&m[438]&m[439])|(m[21]&~m[436]&m[437]&m[438]&m[439])|(~m[21]&m[436]&m[437]&m[438]&m[439])|(m[21]&m[436]&m[437]&m[438]&m[439]));
    m[122] = (((m[22]&m[450]&~m[451]&~m[452]&~m[453])|(m[22]&~m[450]&m[451]&~m[452]&~m[453])|(~m[22]&m[450]&m[451]&~m[452]&~m[453])|(m[22]&~m[450]&~m[451]&m[452]&~m[453])|(~m[22]&m[450]&~m[451]&m[452]&~m[453])|(~m[22]&~m[450]&m[451]&m[452]&~m[453])|(m[22]&~m[450]&~m[451]&~m[452]&m[453])|(~m[22]&m[450]&~m[451]&~m[452]&m[453])|(~m[22]&~m[450]&m[451]&~m[452]&m[453])|(~m[22]&~m[450]&~m[451]&m[452]&m[453]))&BiasedRNG[302])|(((m[22]&m[450]&m[451]&~m[452]&~m[453])|(m[22]&m[450]&~m[451]&m[452]&~m[453])|(m[22]&~m[450]&m[451]&m[452]&~m[453])|(~m[22]&m[450]&m[451]&m[452]&~m[453])|(m[22]&m[450]&~m[451]&~m[452]&m[453])|(m[22]&~m[450]&m[451]&~m[452]&m[453])|(~m[22]&m[450]&m[451]&~m[452]&m[453])|(m[22]&~m[450]&~m[451]&m[452]&m[453])|(~m[22]&m[450]&~m[451]&m[452]&m[453])|(~m[22]&~m[450]&m[451]&m[452]&m[453]))&~BiasedRNG[302])|((m[22]&m[450]&m[451]&m[452]&~m[453])|(m[22]&m[450]&m[451]&~m[452]&m[453])|(m[22]&m[450]&~m[451]&m[452]&m[453])|(m[22]&~m[450]&m[451]&m[452]&m[453])|(~m[22]&m[450]&m[451]&m[452]&m[453])|(m[22]&m[450]&m[451]&m[452]&m[453]));
    m[125] = (((m[23]&m[464]&~m[465]&~m[466]&~m[467])|(m[23]&~m[464]&m[465]&~m[466]&~m[467])|(~m[23]&m[464]&m[465]&~m[466]&~m[467])|(m[23]&~m[464]&~m[465]&m[466]&~m[467])|(~m[23]&m[464]&~m[465]&m[466]&~m[467])|(~m[23]&~m[464]&m[465]&m[466]&~m[467])|(m[23]&~m[464]&~m[465]&~m[466]&m[467])|(~m[23]&m[464]&~m[465]&~m[466]&m[467])|(~m[23]&~m[464]&m[465]&~m[466]&m[467])|(~m[23]&~m[464]&~m[465]&m[466]&m[467]))&BiasedRNG[303])|(((m[23]&m[464]&m[465]&~m[466]&~m[467])|(m[23]&m[464]&~m[465]&m[466]&~m[467])|(m[23]&~m[464]&m[465]&m[466]&~m[467])|(~m[23]&m[464]&m[465]&m[466]&~m[467])|(m[23]&m[464]&~m[465]&~m[466]&m[467])|(m[23]&~m[464]&m[465]&~m[466]&m[467])|(~m[23]&m[464]&m[465]&~m[466]&m[467])|(m[23]&~m[464]&~m[465]&m[466]&m[467])|(~m[23]&m[464]&~m[465]&m[466]&m[467])|(~m[23]&~m[464]&m[465]&m[466]&m[467]))&~BiasedRNG[303])|((m[23]&m[464]&m[465]&m[466]&~m[467])|(m[23]&m[464]&m[465]&~m[466]&m[467])|(m[23]&m[464]&~m[465]&m[466]&m[467])|(m[23]&~m[464]&m[465]&m[466]&m[467])|(~m[23]&m[464]&m[465]&m[466]&m[467])|(m[23]&m[464]&m[465]&m[466]&m[467]));
    m[128] = (((m[24]&m[478]&~m[479]&~m[480]&~m[481])|(m[24]&~m[478]&m[479]&~m[480]&~m[481])|(~m[24]&m[478]&m[479]&~m[480]&~m[481])|(m[24]&~m[478]&~m[479]&m[480]&~m[481])|(~m[24]&m[478]&~m[479]&m[480]&~m[481])|(~m[24]&~m[478]&m[479]&m[480]&~m[481])|(m[24]&~m[478]&~m[479]&~m[480]&m[481])|(~m[24]&m[478]&~m[479]&~m[480]&m[481])|(~m[24]&~m[478]&m[479]&~m[480]&m[481])|(~m[24]&~m[478]&~m[479]&m[480]&m[481]))&BiasedRNG[304])|(((m[24]&m[478]&m[479]&~m[480]&~m[481])|(m[24]&m[478]&~m[479]&m[480]&~m[481])|(m[24]&~m[478]&m[479]&m[480]&~m[481])|(~m[24]&m[478]&m[479]&m[480]&~m[481])|(m[24]&m[478]&~m[479]&~m[480]&m[481])|(m[24]&~m[478]&m[479]&~m[480]&m[481])|(~m[24]&m[478]&m[479]&~m[480]&m[481])|(m[24]&~m[478]&~m[479]&m[480]&m[481])|(~m[24]&m[478]&~m[479]&m[480]&m[481])|(~m[24]&~m[478]&m[479]&m[480]&m[481]))&~BiasedRNG[304])|((m[24]&m[478]&m[479]&m[480]&~m[481])|(m[24]&m[478]&m[479]&~m[480]&m[481])|(m[24]&m[478]&~m[479]&m[480]&m[481])|(m[24]&~m[478]&m[479]&m[480]&m[481])|(~m[24]&m[478]&m[479]&m[480]&m[481])|(m[24]&m[478]&m[479]&m[480]&m[481]));
    m[131] = (((m[25]&m[492]&~m[493]&~m[494]&~m[495])|(m[25]&~m[492]&m[493]&~m[494]&~m[495])|(~m[25]&m[492]&m[493]&~m[494]&~m[495])|(m[25]&~m[492]&~m[493]&m[494]&~m[495])|(~m[25]&m[492]&~m[493]&m[494]&~m[495])|(~m[25]&~m[492]&m[493]&m[494]&~m[495])|(m[25]&~m[492]&~m[493]&~m[494]&m[495])|(~m[25]&m[492]&~m[493]&~m[494]&m[495])|(~m[25]&~m[492]&m[493]&~m[494]&m[495])|(~m[25]&~m[492]&~m[493]&m[494]&m[495]))&BiasedRNG[305])|(((m[25]&m[492]&m[493]&~m[494]&~m[495])|(m[25]&m[492]&~m[493]&m[494]&~m[495])|(m[25]&~m[492]&m[493]&m[494]&~m[495])|(~m[25]&m[492]&m[493]&m[494]&~m[495])|(m[25]&m[492]&~m[493]&~m[494]&m[495])|(m[25]&~m[492]&m[493]&~m[494]&m[495])|(~m[25]&m[492]&m[493]&~m[494]&m[495])|(m[25]&~m[492]&~m[493]&m[494]&m[495])|(~m[25]&m[492]&~m[493]&m[494]&m[495])|(~m[25]&~m[492]&m[493]&m[494]&m[495]))&~BiasedRNG[305])|((m[25]&m[492]&m[493]&m[494]&~m[495])|(m[25]&m[492]&m[493]&~m[494]&m[495])|(m[25]&m[492]&~m[493]&m[494]&m[495])|(m[25]&~m[492]&m[493]&m[494]&m[495])|(~m[25]&m[492]&m[493]&m[494]&m[495])|(m[25]&m[492]&m[493]&m[494]&m[495]));
    m[134] = (((m[26]&m[506]&~m[507]&~m[508]&~m[509])|(m[26]&~m[506]&m[507]&~m[508]&~m[509])|(~m[26]&m[506]&m[507]&~m[508]&~m[509])|(m[26]&~m[506]&~m[507]&m[508]&~m[509])|(~m[26]&m[506]&~m[507]&m[508]&~m[509])|(~m[26]&~m[506]&m[507]&m[508]&~m[509])|(m[26]&~m[506]&~m[507]&~m[508]&m[509])|(~m[26]&m[506]&~m[507]&~m[508]&m[509])|(~m[26]&~m[506]&m[507]&~m[508]&m[509])|(~m[26]&~m[506]&~m[507]&m[508]&m[509]))&BiasedRNG[306])|(((m[26]&m[506]&m[507]&~m[508]&~m[509])|(m[26]&m[506]&~m[507]&m[508]&~m[509])|(m[26]&~m[506]&m[507]&m[508]&~m[509])|(~m[26]&m[506]&m[507]&m[508]&~m[509])|(m[26]&m[506]&~m[507]&~m[508]&m[509])|(m[26]&~m[506]&m[507]&~m[508]&m[509])|(~m[26]&m[506]&m[507]&~m[508]&m[509])|(m[26]&~m[506]&~m[507]&m[508]&m[509])|(~m[26]&m[506]&~m[507]&m[508]&m[509])|(~m[26]&~m[506]&m[507]&m[508]&m[509]))&~BiasedRNG[306])|((m[26]&m[506]&m[507]&m[508]&~m[509])|(m[26]&m[506]&m[507]&~m[508]&m[509])|(m[26]&m[506]&~m[507]&m[508]&m[509])|(m[26]&~m[506]&m[507]&m[508]&m[509])|(~m[26]&m[506]&m[507]&m[508]&m[509])|(m[26]&m[506]&m[507]&m[508]&m[509]));
    m[137] = (((m[27]&m[520]&~m[521]&~m[522]&~m[523])|(m[27]&~m[520]&m[521]&~m[522]&~m[523])|(~m[27]&m[520]&m[521]&~m[522]&~m[523])|(m[27]&~m[520]&~m[521]&m[522]&~m[523])|(~m[27]&m[520]&~m[521]&m[522]&~m[523])|(~m[27]&~m[520]&m[521]&m[522]&~m[523])|(m[27]&~m[520]&~m[521]&~m[522]&m[523])|(~m[27]&m[520]&~m[521]&~m[522]&m[523])|(~m[27]&~m[520]&m[521]&~m[522]&m[523])|(~m[27]&~m[520]&~m[521]&m[522]&m[523]))&BiasedRNG[307])|(((m[27]&m[520]&m[521]&~m[522]&~m[523])|(m[27]&m[520]&~m[521]&m[522]&~m[523])|(m[27]&~m[520]&m[521]&m[522]&~m[523])|(~m[27]&m[520]&m[521]&m[522]&~m[523])|(m[27]&m[520]&~m[521]&~m[522]&m[523])|(m[27]&~m[520]&m[521]&~m[522]&m[523])|(~m[27]&m[520]&m[521]&~m[522]&m[523])|(m[27]&~m[520]&~m[521]&m[522]&m[523])|(~m[27]&m[520]&~m[521]&m[522]&m[523])|(~m[27]&~m[520]&m[521]&m[522]&m[523]))&~BiasedRNG[307])|((m[27]&m[520]&m[521]&m[522]&~m[523])|(m[27]&m[520]&m[521]&~m[522]&m[523])|(m[27]&m[520]&~m[521]&m[522]&m[523])|(m[27]&~m[520]&m[521]&m[522]&m[523])|(~m[27]&m[520]&m[521]&m[522]&m[523])|(m[27]&m[520]&m[521]&m[522]&m[523]));
    m[146] = (((~m[57]&~m[420]&~m[616])|(m[57]&m[420]&~m[616]))&BiasedRNG[308])|(((m[57]&~m[420]&~m[616])|(~m[57]&m[420]&m[616]))&~BiasedRNG[308])|((~m[57]&~m[420]&m[616])|(m[57]&~m[420]&m[616])|(m[57]&m[420]&m[616]));
    m[147] = (((~m[57]&~m[434]&~m[630])|(m[57]&m[434]&~m[630]))&BiasedRNG[309])|(((m[57]&~m[434]&~m[630])|(~m[57]&m[434]&m[630]))&~BiasedRNG[309])|((~m[57]&~m[434]&m[630])|(m[57]&~m[434]&m[630])|(m[57]&m[434]&m[630]));
    m[148] = (((~m[57]&~m[448]&~m[644])|(m[57]&m[448]&~m[644]))&BiasedRNG[310])|(((m[57]&~m[448]&~m[644])|(~m[57]&m[448]&m[644]))&~BiasedRNG[310])|((~m[57]&~m[448]&m[644])|(m[57]&~m[448]&m[644])|(m[57]&m[448]&m[644]));
    m[149] = (((~m[57]&~m[462]&~m[658])|(m[57]&m[462]&~m[658]))&BiasedRNG[311])|(((m[57]&~m[462]&~m[658])|(~m[57]&m[462]&m[658]))&~BiasedRNG[311])|((~m[57]&~m[462]&m[658])|(m[57]&~m[462]&m[658])|(m[57]&m[462]&m[658]));
    m[150] = (((~m[58]&~m[476]&~m[672])|(m[58]&m[476]&~m[672]))&BiasedRNG[312])|(((m[58]&~m[476]&~m[672])|(~m[58]&m[476]&m[672]))&~BiasedRNG[312])|((~m[58]&~m[476]&m[672])|(m[58]&~m[476]&m[672])|(m[58]&m[476]&m[672]));
    m[151] = (((~m[58]&~m[490]&~m[686])|(m[58]&m[490]&~m[686]))&BiasedRNG[313])|(((m[58]&~m[490]&~m[686])|(~m[58]&m[490]&m[686]))&~BiasedRNG[313])|((~m[58]&~m[490]&m[686])|(m[58]&~m[490]&m[686])|(m[58]&m[490]&m[686]));
    m[152] = (((~m[58]&~m[504]&~m[700])|(m[58]&m[504]&~m[700]))&BiasedRNG[314])|(((m[58]&~m[504]&~m[700])|(~m[58]&m[504]&m[700]))&~BiasedRNG[314])|((~m[58]&~m[504]&m[700])|(m[58]&~m[504]&m[700])|(m[58]&m[504]&m[700]));
    m[153] = (((~m[58]&~m[518]&~m[714])|(m[58]&m[518]&~m[714]))&BiasedRNG[315])|(((m[58]&~m[518]&~m[714])|(~m[58]&m[518]&m[714]))&~BiasedRNG[315])|((~m[58]&~m[518]&m[714])|(m[58]&~m[518]&m[714])|(m[58]&m[518]&m[714]));
    m[160] = (((~m[60]&~m[421]&~m[617])|(m[60]&m[421]&~m[617]))&BiasedRNG[316])|(((m[60]&~m[421]&~m[617])|(~m[60]&m[421]&m[617]))&~BiasedRNG[316])|((~m[60]&~m[421]&m[617])|(m[60]&~m[421]&m[617])|(m[60]&m[421]&m[617]));
    m[161] = (((~m[60]&~m[435]&~m[631])|(m[60]&m[435]&~m[631]))&BiasedRNG[317])|(((m[60]&~m[435]&~m[631])|(~m[60]&m[435]&m[631]))&~BiasedRNG[317])|((~m[60]&~m[435]&m[631])|(m[60]&~m[435]&m[631])|(m[60]&m[435]&m[631]));
    m[162] = (((~m[60]&~m[449]&~m[645])|(m[60]&m[449]&~m[645]))&BiasedRNG[318])|(((m[60]&~m[449]&~m[645])|(~m[60]&m[449]&m[645]))&~BiasedRNG[318])|((~m[60]&~m[449]&m[645])|(m[60]&~m[449]&m[645])|(m[60]&m[449]&m[645]));
    m[163] = (((~m[60]&~m[463]&~m[659])|(m[60]&m[463]&~m[659]))&BiasedRNG[319])|(((m[60]&~m[463]&~m[659])|(~m[60]&m[463]&m[659]))&~BiasedRNG[319])|((~m[60]&~m[463]&m[659])|(m[60]&~m[463]&m[659])|(m[60]&m[463]&m[659]));
    m[164] = (((~m[61]&~m[477]&~m[673])|(m[61]&m[477]&~m[673]))&BiasedRNG[320])|(((m[61]&~m[477]&~m[673])|(~m[61]&m[477]&m[673]))&~BiasedRNG[320])|((~m[61]&~m[477]&m[673])|(m[61]&~m[477]&m[673])|(m[61]&m[477]&m[673]));
    m[165] = (((~m[61]&~m[491]&~m[687])|(m[61]&m[491]&~m[687]))&BiasedRNG[321])|(((m[61]&~m[491]&~m[687])|(~m[61]&m[491]&m[687]))&~BiasedRNG[321])|((~m[61]&~m[491]&m[687])|(m[61]&~m[491]&m[687])|(m[61]&m[491]&m[687]));
    m[166] = (((~m[61]&~m[505]&~m[701])|(m[61]&m[505]&~m[701]))&BiasedRNG[322])|(((m[61]&~m[505]&~m[701])|(~m[61]&m[505]&m[701]))&~BiasedRNG[322])|((~m[61]&~m[505]&m[701])|(m[61]&~m[505]&m[701])|(m[61]&m[505]&m[701]));
    m[167] = (((~m[61]&~m[519]&~m[715])|(m[61]&m[519]&~m[715]))&BiasedRNG[323])|(((m[61]&~m[519]&~m[715])|(~m[61]&m[519]&m[715]))&~BiasedRNG[323])|((~m[61]&~m[519]&m[715])|(m[61]&~m[519]&m[715])|(m[61]&m[519]&m[715]));
    m[174] = (((~m[63]&~m[422]&~m[618])|(m[63]&m[422]&~m[618]))&BiasedRNG[324])|(((m[63]&~m[422]&~m[618])|(~m[63]&m[422]&m[618]))&~BiasedRNG[324])|((~m[63]&~m[422]&m[618])|(m[63]&~m[422]&m[618])|(m[63]&m[422]&m[618]));
    m[175] = (((~m[63]&~m[436]&~m[632])|(m[63]&m[436]&~m[632]))&BiasedRNG[325])|(((m[63]&~m[436]&~m[632])|(~m[63]&m[436]&m[632]))&~BiasedRNG[325])|((~m[63]&~m[436]&m[632])|(m[63]&~m[436]&m[632])|(m[63]&m[436]&m[632]));
    m[176] = (((~m[63]&~m[450]&~m[646])|(m[63]&m[450]&~m[646]))&BiasedRNG[326])|(((m[63]&~m[450]&~m[646])|(~m[63]&m[450]&m[646]))&~BiasedRNG[326])|((~m[63]&~m[450]&m[646])|(m[63]&~m[450]&m[646])|(m[63]&m[450]&m[646]));
    m[177] = (((~m[63]&~m[464]&~m[660])|(m[63]&m[464]&~m[660]))&BiasedRNG[327])|(((m[63]&~m[464]&~m[660])|(~m[63]&m[464]&m[660]))&~BiasedRNG[327])|((~m[63]&~m[464]&m[660])|(m[63]&~m[464]&m[660])|(m[63]&m[464]&m[660]));
    m[178] = (((~m[64]&~m[478]&~m[674])|(m[64]&m[478]&~m[674]))&BiasedRNG[328])|(((m[64]&~m[478]&~m[674])|(~m[64]&m[478]&m[674]))&~BiasedRNG[328])|((~m[64]&~m[478]&m[674])|(m[64]&~m[478]&m[674])|(m[64]&m[478]&m[674]));
    m[179] = (((~m[64]&~m[492]&~m[688])|(m[64]&m[492]&~m[688]))&BiasedRNG[329])|(((m[64]&~m[492]&~m[688])|(~m[64]&m[492]&m[688]))&~BiasedRNG[329])|((~m[64]&~m[492]&m[688])|(m[64]&~m[492]&m[688])|(m[64]&m[492]&m[688]));
    m[180] = (((~m[64]&~m[506]&~m[702])|(m[64]&m[506]&~m[702]))&BiasedRNG[330])|(((m[64]&~m[506]&~m[702])|(~m[64]&m[506]&m[702]))&~BiasedRNG[330])|((~m[64]&~m[506]&m[702])|(m[64]&~m[506]&m[702])|(m[64]&m[506]&m[702]));
    m[181] = (((~m[64]&~m[520]&~m[716])|(m[64]&m[520]&~m[716]))&BiasedRNG[331])|(((m[64]&~m[520]&~m[716])|(~m[64]&m[520]&m[716]))&~BiasedRNG[331])|((~m[64]&~m[520]&m[716])|(m[64]&~m[520]&m[716])|(m[64]&m[520]&m[716]));
    m[188] = (((~m[66]&~m[423]&~m[619])|(m[66]&m[423]&~m[619]))&BiasedRNG[332])|(((m[66]&~m[423]&~m[619])|(~m[66]&m[423]&m[619]))&~BiasedRNG[332])|((~m[66]&~m[423]&m[619])|(m[66]&~m[423]&m[619])|(m[66]&m[423]&m[619]));
    m[189] = (((~m[66]&~m[437]&~m[633])|(m[66]&m[437]&~m[633]))&BiasedRNG[333])|(((m[66]&~m[437]&~m[633])|(~m[66]&m[437]&m[633]))&~BiasedRNG[333])|((~m[66]&~m[437]&m[633])|(m[66]&~m[437]&m[633])|(m[66]&m[437]&m[633]));
    m[190] = (((~m[66]&~m[451]&~m[647])|(m[66]&m[451]&~m[647]))&BiasedRNG[334])|(((m[66]&~m[451]&~m[647])|(~m[66]&m[451]&m[647]))&~BiasedRNG[334])|((~m[66]&~m[451]&m[647])|(m[66]&~m[451]&m[647])|(m[66]&m[451]&m[647]));
    m[191] = (((~m[66]&~m[465]&~m[661])|(m[66]&m[465]&~m[661]))&BiasedRNG[335])|(((m[66]&~m[465]&~m[661])|(~m[66]&m[465]&m[661]))&~BiasedRNG[335])|((~m[66]&~m[465]&m[661])|(m[66]&~m[465]&m[661])|(m[66]&m[465]&m[661]));
    m[192] = (((~m[67]&~m[479]&~m[675])|(m[67]&m[479]&~m[675]))&BiasedRNG[336])|(((m[67]&~m[479]&~m[675])|(~m[67]&m[479]&m[675]))&~BiasedRNG[336])|((~m[67]&~m[479]&m[675])|(m[67]&~m[479]&m[675])|(m[67]&m[479]&m[675]));
    m[193] = (((~m[67]&~m[493]&~m[689])|(m[67]&m[493]&~m[689]))&BiasedRNG[337])|(((m[67]&~m[493]&~m[689])|(~m[67]&m[493]&m[689]))&~BiasedRNG[337])|((~m[67]&~m[493]&m[689])|(m[67]&~m[493]&m[689])|(m[67]&m[493]&m[689]));
    m[194] = (((~m[67]&~m[507]&~m[703])|(m[67]&m[507]&~m[703]))&BiasedRNG[338])|(((m[67]&~m[507]&~m[703])|(~m[67]&m[507]&m[703]))&~BiasedRNG[338])|((~m[67]&~m[507]&m[703])|(m[67]&~m[507]&m[703])|(m[67]&m[507]&m[703]));
    m[195] = (((~m[67]&~m[521]&~m[717])|(m[67]&m[521]&~m[717]))&BiasedRNG[339])|(((m[67]&~m[521]&~m[717])|(~m[67]&m[521]&m[717]))&~BiasedRNG[339])|((~m[67]&~m[521]&m[717])|(m[67]&~m[521]&m[717])|(m[67]&m[521]&m[717]));
    m[202] = (((~m[69]&~m[424]&~m[620])|(m[69]&m[424]&~m[620]))&BiasedRNG[340])|(((m[69]&~m[424]&~m[620])|(~m[69]&m[424]&m[620]))&~BiasedRNG[340])|((~m[69]&~m[424]&m[620])|(m[69]&~m[424]&m[620])|(m[69]&m[424]&m[620]));
    m[203] = (((~m[69]&~m[438]&~m[634])|(m[69]&m[438]&~m[634]))&BiasedRNG[341])|(((m[69]&~m[438]&~m[634])|(~m[69]&m[438]&m[634]))&~BiasedRNG[341])|((~m[69]&~m[438]&m[634])|(m[69]&~m[438]&m[634])|(m[69]&m[438]&m[634]));
    m[204] = (((~m[69]&~m[452]&~m[648])|(m[69]&m[452]&~m[648]))&BiasedRNG[342])|(((m[69]&~m[452]&~m[648])|(~m[69]&m[452]&m[648]))&~BiasedRNG[342])|((~m[69]&~m[452]&m[648])|(m[69]&~m[452]&m[648])|(m[69]&m[452]&m[648]));
    m[205] = (((~m[69]&~m[466]&~m[662])|(m[69]&m[466]&~m[662]))&BiasedRNG[343])|(((m[69]&~m[466]&~m[662])|(~m[69]&m[466]&m[662]))&~BiasedRNG[343])|((~m[69]&~m[466]&m[662])|(m[69]&~m[466]&m[662])|(m[69]&m[466]&m[662]));
    m[206] = (((~m[70]&~m[480]&~m[676])|(m[70]&m[480]&~m[676]))&BiasedRNG[344])|(((m[70]&~m[480]&~m[676])|(~m[70]&m[480]&m[676]))&~BiasedRNG[344])|((~m[70]&~m[480]&m[676])|(m[70]&~m[480]&m[676])|(m[70]&m[480]&m[676]));
    m[207] = (((~m[70]&~m[494]&~m[690])|(m[70]&m[494]&~m[690]))&BiasedRNG[345])|(((m[70]&~m[494]&~m[690])|(~m[70]&m[494]&m[690]))&~BiasedRNG[345])|((~m[70]&~m[494]&m[690])|(m[70]&~m[494]&m[690])|(m[70]&m[494]&m[690]));
    m[208] = (((~m[70]&~m[508]&~m[704])|(m[70]&m[508]&~m[704]))&BiasedRNG[346])|(((m[70]&~m[508]&~m[704])|(~m[70]&m[508]&m[704]))&~BiasedRNG[346])|((~m[70]&~m[508]&m[704])|(m[70]&~m[508]&m[704])|(m[70]&m[508]&m[704]));
    m[209] = (((~m[70]&~m[522]&~m[718])|(m[70]&m[522]&~m[718]))&BiasedRNG[347])|(((m[70]&~m[522]&~m[718])|(~m[70]&m[522]&m[718]))&~BiasedRNG[347])|((~m[70]&~m[522]&m[718])|(m[70]&~m[522]&m[718])|(m[70]&m[522]&m[718]));
    m[216] = (((~m[72]&~m[425]&~m[621])|(m[72]&m[425]&~m[621]))&BiasedRNG[348])|(((m[72]&~m[425]&~m[621])|(~m[72]&m[425]&m[621]))&~BiasedRNG[348])|((~m[72]&~m[425]&m[621])|(m[72]&~m[425]&m[621])|(m[72]&m[425]&m[621]));
    m[217] = (((~m[72]&~m[439]&~m[635])|(m[72]&m[439]&~m[635]))&BiasedRNG[349])|(((m[72]&~m[439]&~m[635])|(~m[72]&m[439]&m[635]))&~BiasedRNG[349])|((~m[72]&~m[439]&m[635])|(m[72]&~m[439]&m[635])|(m[72]&m[439]&m[635]));
    m[218] = (((~m[72]&~m[453]&~m[649])|(m[72]&m[453]&~m[649]))&BiasedRNG[350])|(((m[72]&~m[453]&~m[649])|(~m[72]&m[453]&m[649]))&~BiasedRNG[350])|((~m[72]&~m[453]&m[649])|(m[72]&~m[453]&m[649])|(m[72]&m[453]&m[649]));
    m[219] = (((~m[72]&~m[467]&~m[663])|(m[72]&m[467]&~m[663]))&BiasedRNG[351])|(((m[72]&~m[467]&~m[663])|(~m[72]&m[467]&m[663]))&~BiasedRNG[351])|((~m[72]&~m[467]&m[663])|(m[72]&~m[467]&m[663])|(m[72]&m[467]&m[663]));
    m[220] = (((~m[73]&~m[481]&~m[677])|(m[73]&m[481]&~m[677]))&BiasedRNG[352])|(((m[73]&~m[481]&~m[677])|(~m[73]&m[481]&m[677]))&~BiasedRNG[352])|((~m[73]&~m[481]&m[677])|(m[73]&~m[481]&m[677])|(m[73]&m[481]&m[677]));
    m[221] = (((~m[73]&~m[495]&~m[691])|(m[73]&m[495]&~m[691]))&BiasedRNG[353])|(((m[73]&~m[495]&~m[691])|(~m[73]&m[495]&m[691]))&~BiasedRNG[353])|((~m[73]&~m[495]&m[691])|(m[73]&~m[495]&m[691])|(m[73]&m[495]&m[691]));
    m[222] = (((~m[73]&~m[509]&~m[705])|(m[73]&m[509]&~m[705]))&BiasedRNG[354])|(((m[73]&~m[509]&~m[705])|(~m[73]&m[509]&m[705]))&~BiasedRNG[354])|((~m[73]&~m[509]&m[705])|(m[73]&~m[509]&m[705])|(m[73]&m[509]&m[705]));
    m[223] = (((~m[73]&~m[523]&~m[719])|(m[73]&m[523]&~m[719]))&BiasedRNG[355])|(((m[73]&~m[523]&~m[719])|(~m[73]&m[523]&m[719]))&~BiasedRNG[355])|((~m[73]&~m[523]&m[719])|(m[73]&~m[523]&m[719])|(m[73]&m[523]&m[719]));
    m[230] = (((~m[75]&~m[426]&~m[622])|(m[75]&m[426]&~m[622]))&BiasedRNG[356])|(((m[75]&~m[426]&~m[622])|(~m[75]&m[426]&m[622]))&~BiasedRNG[356])|((~m[75]&~m[426]&m[622])|(m[75]&~m[426]&m[622])|(m[75]&m[426]&m[622]));
    m[231] = (((~m[75]&~m[440]&~m[636])|(m[75]&m[440]&~m[636]))&BiasedRNG[357])|(((m[75]&~m[440]&~m[636])|(~m[75]&m[440]&m[636]))&~BiasedRNG[357])|((~m[75]&~m[440]&m[636])|(m[75]&~m[440]&m[636])|(m[75]&m[440]&m[636]));
    m[232] = (((~m[75]&~m[454]&~m[650])|(m[75]&m[454]&~m[650]))&BiasedRNG[358])|(((m[75]&~m[454]&~m[650])|(~m[75]&m[454]&m[650]))&~BiasedRNG[358])|((~m[75]&~m[454]&m[650])|(m[75]&~m[454]&m[650])|(m[75]&m[454]&m[650]));
    m[233] = (((~m[75]&~m[468]&~m[664])|(m[75]&m[468]&~m[664]))&BiasedRNG[359])|(((m[75]&~m[468]&~m[664])|(~m[75]&m[468]&m[664]))&~BiasedRNG[359])|((~m[75]&~m[468]&m[664])|(m[75]&~m[468]&m[664])|(m[75]&m[468]&m[664]));
    m[234] = (((~m[76]&~m[482]&~m[678])|(m[76]&m[482]&~m[678]))&BiasedRNG[360])|(((m[76]&~m[482]&~m[678])|(~m[76]&m[482]&m[678]))&~BiasedRNG[360])|((~m[76]&~m[482]&m[678])|(m[76]&~m[482]&m[678])|(m[76]&m[482]&m[678]));
    m[235] = (((~m[76]&~m[496]&~m[692])|(m[76]&m[496]&~m[692]))&BiasedRNG[361])|(((m[76]&~m[496]&~m[692])|(~m[76]&m[496]&m[692]))&~BiasedRNG[361])|((~m[76]&~m[496]&m[692])|(m[76]&~m[496]&m[692])|(m[76]&m[496]&m[692]));
    m[236] = (((~m[76]&~m[510]&~m[706])|(m[76]&m[510]&~m[706]))&BiasedRNG[362])|(((m[76]&~m[510]&~m[706])|(~m[76]&m[510]&m[706]))&~BiasedRNG[362])|((~m[76]&~m[510]&m[706])|(m[76]&~m[510]&m[706])|(m[76]&m[510]&m[706]));
    m[237] = (((~m[76]&~m[524]&~m[720])|(m[76]&m[524]&~m[720]))&BiasedRNG[363])|(((m[76]&~m[524]&~m[720])|(~m[76]&m[524]&m[720]))&~BiasedRNG[363])|((~m[76]&~m[524]&m[720])|(m[76]&~m[524]&m[720])|(m[76]&m[524]&m[720]));
    m[244] = (((~m[78]&~m[427]&~m[623])|(m[78]&m[427]&~m[623]))&BiasedRNG[364])|(((m[78]&~m[427]&~m[623])|(~m[78]&m[427]&m[623]))&~BiasedRNG[364])|((~m[78]&~m[427]&m[623])|(m[78]&~m[427]&m[623])|(m[78]&m[427]&m[623]));
    m[245] = (((~m[78]&~m[441]&~m[637])|(m[78]&m[441]&~m[637]))&BiasedRNG[365])|(((m[78]&~m[441]&~m[637])|(~m[78]&m[441]&m[637]))&~BiasedRNG[365])|((~m[78]&~m[441]&m[637])|(m[78]&~m[441]&m[637])|(m[78]&m[441]&m[637]));
    m[246] = (((~m[78]&~m[455]&~m[651])|(m[78]&m[455]&~m[651]))&BiasedRNG[366])|(((m[78]&~m[455]&~m[651])|(~m[78]&m[455]&m[651]))&~BiasedRNG[366])|((~m[78]&~m[455]&m[651])|(m[78]&~m[455]&m[651])|(m[78]&m[455]&m[651]));
    m[247] = (((~m[78]&~m[469]&~m[665])|(m[78]&m[469]&~m[665]))&BiasedRNG[367])|(((m[78]&~m[469]&~m[665])|(~m[78]&m[469]&m[665]))&~BiasedRNG[367])|((~m[78]&~m[469]&m[665])|(m[78]&~m[469]&m[665])|(m[78]&m[469]&m[665]));
    m[248] = (((~m[79]&~m[483]&~m[679])|(m[79]&m[483]&~m[679]))&BiasedRNG[368])|(((m[79]&~m[483]&~m[679])|(~m[79]&m[483]&m[679]))&~BiasedRNG[368])|((~m[79]&~m[483]&m[679])|(m[79]&~m[483]&m[679])|(m[79]&m[483]&m[679]));
    m[249] = (((~m[79]&~m[497]&~m[693])|(m[79]&m[497]&~m[693]))&BiasedRNG[369])|(((m[79]&~m[497]&~m[693])|(~m[79]&m[497]&m[693]))&~BiasedRNG[369])|((~m[79]&~m[497]&m[693])|(m[79]&~m[497]&m[693])|(m[79]&m[497]&m[693]));
    m[250] = (((~m[79]&~m[511]&~m[707])|(m[79]&m[511]&~m[707]))&BiasedRNG[370])|(((m[79]&~m[511]&~m[707])|(~m[79]&m[511]&m[707]))&~BiasedRNG[370])|((~m[79]&~m[511]&m[707])|(m[79]&~m[511]&m[707])|(m[79]&m[511]&m[707]));
    m[251] = (((~m[79]&~m[525]&~m[721])|(m[79]&m[525]&~m[721]))&BiasedRNG[371])|(((m[79]&~m[525]&~m[721])|(~m[79]&m[525]&m[721]))&~BiasedRNG[371])|((~m[79]&~m[525]&m[721])|(m[79]&~m[525]&m[721])|(m[79]&m[525]&m[721]));
    m[258] = (((~m[81]&~m[428]&~m[624])|(m[81]&m[428]&~m[624]))&BiasedRNG[372])|(((m[81]&~m[428]&~m[624])|(~m[81]&m[428]&m[624]))&~BiasedRNG[372])|((~m[81]&~m[428]&m[624])|(m[81]&~m[428]&m[624])|(m[81]&m[428]&m[624]));
    m[259] = (((~m[81]&~m[442]&~m[638])|(m[81]&m[442]&~m[638]))&BiasedRNG[373])|(((m[81]&~m[442]&~m[638])|(~m[81]&m[442]&m[638]))&~BiasedRNG[373])|((~m[81]&~m[442]&m[638])|(m[81]&~m[442]&m[638])|(m[81]&m[442]&m[638]));
    m[260] = (((~m[81]&~m[456]&~m[652])|(m[81]&m[456]&~m[652]))&BiasedRNG[374])|(((m[81]&~m[456]&~m[652])|(~m[81]&m[456]&m[652]))&~BiasedRNG[374])|((~m[81]&~m[456]&m[652])|(m[81]&~m[456]&m[652])|(m[81]&m[456]&m[652]));
    m[261] = (((~m[81]&~m[470]&~m[666])|(m[81]&m[470]&~m[666]))&BiasedRNG[375])|(((m[81]&~m[470]&~m[666])|(~m[81]&m[470]&m[666]))&~BiasedRNG[375])|((~m[81]&~m[470]&m[666])|(m[81]&~m[470]&m[666])|(m[81]&m[470]&m[666]));
    m[262] = (((~m[82]&~m[484]&~m[680])|(m[82]&m[484]&~m[680]))&BiasedRNG[376])|(((m[82]&~m[484]&~m[680])|(~m[82]&m[484]&m[680]))&~BiasedRNG[376])|((~m[82]&~m[484]&m[680])|(m[82]&~m[484]&m[680])|(m[82]&m[484]&m[680]));
    m[263] = (((~m[82]&~m[498]&~m[694])|(m[82]&m[498]&~m[694]))&BiasedRNG[377])|(((m[82]&~m[498]&~m[694])|(~m[82]&m[498]&m[694]))&~BiasedRNG[377])|((~m[82]&~m[498]&m[694])|(m[82]&~m[498]&m[694])|(m[82]&m[498]&m[694]));
    m[264] = (((~m[82]&~m[512]&~m[708])|(m[82]&m[512]&~m[708]))&BiasedRNG[378])|(((m[82]&~m[512]&~m[708])|(~m[82]&m[512]&m[708]))&~BiasedRNG[378])|((~m[82]&~m[512]&m[708])|(m[82]&~m[512]&m[708])|(m[82]&m[512]&m[708]));
    m[265] = (((~m[82]&~m[526]&~m[722])|(m[82]&m[526]&~m[722]))&BiasedRNG[379])|(((m[82]&~m[526]&~m[722])|(~m[82]&m[526]&m[722]))&~BiasedRNG[379])|((~m[82]&~m[526]&m[722])|(m[82]&~m[526]&m[722])|(m[82]&m[526]&m[722]));
    m[272] = (((~m[84]&~m[429]&~m[625])|(m[84]&m[429]&~m[625]))&BiasedRNG[380])|(((m[84]&~m[429]&~m[625])|(~m[84]&m[429]&m[625]))&~BiasedRNG[380])|((~m[84]&~m[429]&m[625])|(m[84]&~m[429]&m[625])|(m[84]&m[429]&m[625]));
    m[273] = (((~m[84]&~m[443]&~m[639])|(m[84]&m[443]&~m[639]))&BiasedRNG[381])|(((m[84]&~m[443]&~m[639])|(~m[84]&m[443]&m[639]))&~BiasedRNG[381])|((~m[84]&~m[443]&m[639])|(m[84]&~m[443]&m[639])|(m[84]&m[443]&m[639]));
    m[274] = (((~m[84]&~m[457]&~m[653])|(m[84]&m[457]&~m[653]))&BiasedRNG[382])|(((m[84]&~m[457]&~m[653])|(~m[84]&m[457]&m[653]))&~BiasedRNG[382])|((~m[84]&~m[457]&m[653])|(m[84]&~m[457]&m[653])|(m[84]&m[457]&m[653]));
    m[275] = (((~m[84]&~m[471]&~m[667])|(m[84]&m[471]&~m[667]))&BiasedRNG[383])|(((m[84]&~m[471]&~m[667])|(~m[84]&m[471]&m[667]))&~BiasedRNG[383])|((~m[84]&~m[471]&m[667])|(m[84]&~m[471]&m[667])|(m[84]&m[471]&m[667]));
    m[276] = (((~m[85]&~m[485]&~m[681])|(m[85]&m[485]&~m[681]))&BiasedRNG[384])|(((m[85]&~m[485]&~m[681])|(~m[85]&m[485]&m[681]))&~BiasedRNG[384])|((~m[85]&~m[485]&m[681])|(m[85]&~m[485]&m[681])|(m[85]&m[485]&m[681]));
    m[277] = (((~m[85]&~m[499]&~m[695])|(m[85]&m[499]&~m[695]))&BiasedRNG[385])|(((m[85]&~m[499]&~m[695])|(~m[85]&m[499]&m[695]))&~BiasedRNG[385])|((~m[85]&~m[499]&m[695])|(m[85]&~m[499]&m[695])|(m[85]&m[499]&m[695]));
    m[278] = (((~m[85]&~m[513]&~m[709])|(m[85]&m[513]&~m[709]))&BiasedRNG[386])|(((m[85]&~m[513]&~m[709])|(~m[85]&m[513]&m[709]))&~BiasedRNG[386])|((~m[85]&~m[513]&m[709])|(m[85]&~m[513]&m[709])|(m[85]&m[513]&m[709]));
    m[279] = (((~m[85]&~m[527]&~m[723])|(m[85]&m[527]&~m[723]))&BiasedRNG[387])|(((m[85]&~m[527]&~m[723])|(~m[85]&m[527]&m[723]))&~BiasedRNG[387])|((~m[85]&~m[527]&m[723])|(m[85]&~m[527]&m[723])|(m[85]&m[527]&m[723]));
    m[286] = (((~m[87]&~m[430]&~m[626])|(m[87]&m[430]&~m[626]))&BiasedRNG[388])|(((m[87]&~m[430]&~m[626])|(~m[87]&m[430]&m[626]))&~BiasedRNG[388])|((~m[87]&~m[430]&m[626])|(m[87]&~m[430]&m[626])|(m[87]&m[430]&m[626]));
    m[287] = (((~m[87]&~m[444]&~m[640])|(m[87]&m[444]&~m[640]))&BiasedRNG[389])|(((m[87]&~m[444]&~m[640])|(~m[87]&m[444]&m[640]))&~BiasedRNG[389])|((~m[87]&~m[444]&m[640])|(m[87]&~m[444]&m[640])|(m[87]&m[444]&m[640]));
    m[288] = (((~m[87]&~m[458]&~m[654])|(m[87]&m[458]&~m[654]))&BiasedRNG[390])|(((m[87]&~m[458]&~m[654])|(~m[87]&m[458]&m[654]))&~BiasedRNG[390])|((~m[87]&~m[458]&m[654])|(m[87]&~m[458]&m[654])|(m[87]&m[458]&m[654]));
    m[289] = (((~m[87]&~m[472]&~m[668])|(m[87]&m[472]&~m[668]))&BiasedRNG[391])|(((m[87]&~m[472]&~m[668])|(~m[87]&m[472]&m[668]))&~BiasedRNG[391])|((~m[87]&~m[472]&m[668])|(m[87]&~m[472]&m[668])|(m[87]&m[472]&m[668]));
    m[290] = (((~m[88]&~m[486]&~m[682])|(m[88]&m[486]&~m[682]))&BiasedRNG[392])|(((m[88]&~m[486]&~m[682])|(~m[88]&m[486]&m[682]))&~BiasedRNG[392])|((~m[88]&~m[486]&m[682])|(m[88]&~m[486]&m[682])|(m[88]&m[486]&m[682]));
    m[291] = (((~m[88]&~m[500]&~m[696])|(m[88]&m[500]&~m[696]))&BiasedRNG[393])|(((m[88]&~m[500]&~m[696])|(~m[88]&m[500]&m[696]))&~BiasedRNG[393])|((~m[88]&~m[500]&m[696])|(m[88]&~m[500]&m[696])|(m[88]&m[500]&m[696]));
    m[292] = (((~m[88]&~m[514]&~m[710])|(m[88]&m[514]&~m[710]))&BiasedRNG[394])|(((m[88]&~m[514]&~m[710])|(~m[88]&m[514]&m[710]))&~BiasedRNG[394])|((~m[88]&~m[514]&m[710])|(m[88]&~m[514]&m[710])|(m[88]&m[514]&m[710]));
    m[293] = (((~m[88]&~m[528]&~m[724])|(m[88]&m[528]&~m[724]))&BiasedRNG[395])|(((m[88]&~m[528]&~m[724])|(~m[88]&m[528]&m[724]))&~BiasedRNG[395])|((~m[88]&~m[528]&m[724])|(m[88]&~m[528]&m[724])|(m[88]&m[528]&m[724]));
    m[300] = (((~m[90]&~m[431]&~m[627])|(m[90]&m[431]&~m[627]))&BiasedRNG[396])|(((m[90]&~m[431]&~m[627])|(~m[90]&m[431]&m[627]))&~BiasedRNG[396])|((~m[90]&~m[431]&m[627])|(m[90]&~m[431]&m[627])|(m[90]&m[431]&m[627]));
    m[301] = (((~m[90]&~m[445]&~m[641])|(m[90]&m[445]&~m[641]))&BiasedRNG[397])|(((m[90]&~m[445]&~m[641])|(~m[90]&m[445]&m[641]))&~BiasedRNG[397])|((~m[90]&~m[445]&m[641])|(m[90]&~m[445]&m[641])|(m[90]&m[445]&m[641]));
    m[302] = (((~m[90]&~m[459]&~m[655])|(m[90]&m[459]&~m[655]))&BiasedRNG[398])|(((m[90]&~m[459]&~m[655])|(~m[90]&m[459]&m[655]))&~BiasedRNG[398])|((~m[90]&~m[459]&m[655])|(m[90]&~m[459]&m[655])|(m[90]&m[459]&m[655]));
    m[303] = (((~m[90]&~m[473]&~m[669])|(m[90]&m[473]&~m[669]))&BiasedRNG[399])|(((m[90]&~m[473]&~m[669])|(~m[90]&m[473]&m[669]))&~BiasedRNG[399])|((~m[90]&~m[473]&m[669])|(m[90]&~m[473]&m[669])|(m[90]&m[473]&m[669]));
    m[304] = (((~m[91]&~m[487]&~m[683])|(m[91]&m[487]&~m[683]))&BiasedRNG[400])|(((m[91]&~m[487]&~m[683])|(~m[91]&m[487]&m[683]))&~BiasedRNG[400])|((~m[91]&~m[487]&m[683])|(m[91]&~m[487]&m[683])|(m[91]&m[487]&m[683]));
    m[305] = (((~m[91]&~m[501]&~m[697])|(m[91]&m[501]&~m[697]))&BiasedRNG[401])|(((m[91]&~m[501]&~m[697])|(~m[91]&m[501]&m[697]))&~BiasedRNG[401])|((~m[91]&~m[501]&m[697])|(m[91]&~m[501]&m[697])|(m[91]&m[501]&m[697]));
    m[306] = (((~m[91]&~m[515]&~m[711])|(m[91]&m[515]&~m[711]))&BiasedRNG[402])|(((m[91]&~m[515]&~m[711])|(~m[91]&m[515]&m[711]))&~BiasedRNG[402])|((~m[91]&~m[515]&m[711])|(m[91]&~m[515]&m[711])|(m[91]&m[515]&m[711]));
    m[307] = (((~m[91]&~m[529]&~m[725])|(m[91]&m[529]&~m[725]))&BiasedRNG[403])|(((m[91]&~m[529]&~m[725])|(~m[91]&m[529]&m[725]))&~BiasedRNG[403])|((~m[91]&~m[529]&m[725])|(m[91]&~m[529]&m[725])|(m[91]&m[529]&m[725]));
    m[314] = (((~m[93]&~m[432]&~m[628])|(m[93]&m[432]&~m[628]))&BiasedRNG[404])|(((m[93]&~m[432]&~m[628])|(~m[93]&m[432]&m[628]))&~BiasedRNG[404])|((~m[93]&~m[432]&m[628])|(m[93]&~m[432]&m[628])|(m[93]&m[432]&m[628]));
    m[315] = (((~m[93]&~m[446]&~m[642])|(m[93]&m[446]&~m[642]))&BiasedRNG[405])|(((m[93]&~m[446]&~m[642])|(~m[93]&m[446]&m[642]))&~BiasedRNG[405])|((~m[93]&~m[446]&m[642])|(m[93]&~m[446]&m[642])|(m[93]&m[446]&m[642]));
    m[316] = (((~m[93]&~m[460]&~m[656])|(m[93]&m[460]&~m[656]))&BiasedRNG[406])|(((m[93]&~m[460]&~m[656])|(~m[93]&m[460]&m[656]))&~BiasedRNG[406])|((~m[93]&~m[460]&m[656])|(m[93]&~m[460]&m[656])|(m[93]&m[460]&m[656]));
    m[317] = (((~m[93]&~m[474]&~m[670])|(m[93]&m[474]&~m[670]))&BiasedRNG[407])|(((m[93]&~m[474]&~m[670])|(~m[93]&m[474]&m[670]))&~BiasedRNG[407])|((~m[93]&~m[474]&m[670])|(m[93]&~m[474]&m[670])|(m[93]&m[474]&m[670]));
    m[318] = (((~m[94]&~m[488]&~m[684])|(m[94]&m[488]&~m[684]))&BiasedRNG[408])|(((m[94]&~m[488]&~m[684])|(~m[94]&m[488]&m[684]))&~BiasedRNG[408])|((~m[94]&~m[488]&m[684])|(m[94]&~m[488]&m[684])|(m[94]&m[488]&m[684]));
    m[319] = (((~m[94]&~m[502]&~m[698])|(m[94]&m[502]&~m[698]))&BiasedRNG[409])|(((m[94]&~m[502]&~m[698])|(~m[94]&m[502]&m[698]))&~BiasedRNG[409])|((~m[94]&~m[502]&m[698])|(m[94]&~m[502]&m[698])|(m[94]&m[502]&m[698]));
    m[320] = (((~m[94]&~m[516]&~m[712])|(m[94]&m[516]&~m[712]))&BiasedRNG[410])|(((m[94]&~m[516]&~m[712])|(~m[94]&m[516]&m[712]))&~BiasedRNG[410])|((~m[94]&~m[516]&m[712])|(m[94]&~m[516]&m[712])|(m[94]&m[516]&m[712]));
    m[321] = (((~m[94]&~m[530]&~m[726])|(m[94]&m[530]&~m[726]))&BiasedRNG[411])|(((m[94]&~m[530]&~m[726])|(~m[94]&m[530]&m[726]))&~BiasedRNG[411])|((~m[94]&~m[530]&m[726])|(m[94]&~m[530]&m[726])|(m[94]&m[530]&m[726]));
    m[328] = (((~m[96]&~m[433]&~m[629])|(m[96]&m[433]&~m[629]))&BiasedRNG[412])|(((m[96]&~m[433]&~m[629])|(~m[96]&m[433]&m[629]))&~BiasedRNG[412])|((~m[96]&~m[433]&m[629])|(m[96]&~m[433]&m[629])|(m[96]&m[433]&m[629]));
    m[329] = (((~m[96]&~m[447]&~m[643])|(m[96]&m[447]&~m[643]))&BiasedRNG[413])|(((m[96]&~m[447]&~m[643])|(~m[96]&m[447]&m[643]))&~BiasedRNG[413])|((~m[96]&~m[447]&m[643])|(m[96]&~m[447]&m[643])|(m[96]&m[447]&m[643]));
    m[330] = (((~m[96]&~m[461]&~m[657])|(m[96]&m[461]&~m[657]))&BiasedRNG[414])|(((m[96]&~m[461]&~m[657])|(~m[96]&m[461]&m[657]))&~BiasedRNG[414])|((~m[96]&~m[461]&m[657])|(m[96]&~m[461]&m[657])|(m[96]&m[461]&m[657]));
    m[331] = (((~m[96]&~m[475]&~m[671])|(m[96]&m[475]&~m[671]))&BiasedRNG[415])|(((m[96]&~m[475]&~m[671])|(~m[96]&m[475]&m[671]))&~BiasedRNG[415])|((~m[96]&~m[475]&m[671])|(m[96]&~m[475]&m[671])|(m[96]&m[475]&m[671]));
    m[332] = (((~m[97]&~m[489]&~m[685])|(m[97]&m[489]&~m[685]))&BiasedRNG[416])|(((m[97]&~m[489]&~m[685])|(~m[97]&m[489]&m[685]))&~BiasedRNG[416])|((~m[97]&~m[489]&m[685])|(m[97]&~m[489]&m[685])|(m[97]&m[489]&m[685]));
    m[333] = (((~m[97]&~m[503]&~m[699])|(m[97]&m[503]&~m[699]))&BiasedRNG[417])|(((m[97]&~m[503]&~m[699])|(~m[97]&m[503]&m[699]))&~BiasedRNG[417])|((~m[97]&~m[503]&m[699])|(m[97]&~m[503]&m[699])|(m[97]&m[503]&m[699]));
    m[334] = (((~m[97]&~m[517]&~m[713])|(m[97]&m[517]&~m[713]))&BiasedRNG[418])|(((m[97]&~m[517]&~m[713])|(~m[97]&m[517]&m[713]))&~BiasedRNG[418])|((~m[97]&~m[517]&m[713])|(m[97]&~m[517]&m[713])|(m[97]&m[517]&m[713]));
    m[335] = (((~m[97]&~m[531]&~m[727])|(m[97]&m[531]&~m[727]))&BiasedRNG[419])|(((m[97]&~m[531]&~m[727])|(~m[97]&m[531]&m[727]))&~BiasedRNG[419])|((~m[97]&~m[531]&m[727])|(m[97]&~m[531]&m[727])|(m[97]&m[531]&m[727]));
    m[342] = (((~m[99]&~m[224]&~m[538])|(m[99]&m[224]&~m[538]))&BiasedRNG[420])|(((m[99]&~m[224]&~m[538])|(~m[99]&m[224]&m[538]))&~BiasedRNG[420])|((~m[99]&~m[224]&m[538])|(m[99]&~m[224]&m[538])|(m[99]&m[224]&m[538]));
    m[343] = (((~m[99]&~m[238]&~m[539])|(m[99]&m[238]&~m[539]))&BiasedRNG[421])|(((m[99]&~m[238]&~m[539])|(~m[99]&m[238]&m[539]))&~BiasedRNG[421])|((~m[99]&~m[238]&m[539])|(m[99]&~m[238]&m[539])|(m[99]&m[238]&m[539]));
    m[344] = (((~m[99]&~m[252]&~m[540])|(m[99]&m[252]&~m[540]))&BiasedRNG[422])|(((m[99]&~m[252]&~m[540])|(~m[99]&m[252]&m[540]))&~BiasedRNG[422])|((~m[99]&~m[252]&m[540])|(m[99]&~m[252]&m[540])|(m[99]&m[252]&m[540]));
    m[345] = (((~m[99]&~m[266]&~m[541])|(m[99]&m[266]&~m[541]))&BiasedRNG[423])|(((m[99]&~m[266]&~m[541])|(~m[99]&m[266]&m[541]))&~BiasedRNG[423])|((~m[99]&~m[266]&m[541])|(m[99]&~m[266]&m[541])|(m[99]&m[266]&m[541]));
    m[346] = (((~m[100]&~m[280]&~m[542])|(m[100]&m[280]&~m[542]))&BiasedRNG[424])|(((m[100]&~m[280]&~m[542])|(~m[100]&m[280]&m[542]))&~BiasedRNG[424])|((~m[100]&~m[280]&m[542])|(m[100]&~m[280]&m[542])|(m[100]&m[280]&m[542]));
    m[347] = (((~m[100]&~m[294]&~m[543])|(m[100]&m[294]&~m[543]))&BiasedRNG[425])|(((m[100]&~m[294]&~m[543])|(~m[100]&m[294]&m[543]))&~BiasedRNG[425])|((~m[100]&~m[294]&m[543])|(m[100]&~m[294]&m[543])|(m[100]&m[294]&m[543]));
    m[348] = (((~m[100]&~m[308]&~m[544])|(m[100]&m[308]&~m[544]))&BiasedRNG[426])|(((m[100]&~m[308]&~m[544])|(~m[100]&m[308]&m[544]))&~BiasedRNG[426])|((~m[100]&~m[308]&m[544])|(m[100]&~m[308]&m[544])|(m[100]&m[308]&m[544]));
    m[349] = (((~m[100]&~m[322]&~m[545])|(m[100]&m[322]&~m[545]))&BiasedRNG[427])|(((m[100]&~m[322]&~m[545])|(~m[100]&m[322]&m[545]))&~BiasedRNG[427])|((~m[100]&~m[322]&m[545])|(m[100]&~m[322]&m[545])|(m[100]&m[322]&m[545]));
    m[356] = (((~m[102]&~m[225]&~m[552])|(m[102]&m[225]&~m[552]))&BiasedRNG[428])|(((m[102]&~m[225]&~m[552])|(~m[102]&m[225]&m[552]))&~BiasedRNG[428])|((~m[102]&~m[225]&m[552])|(m[102]&~m[225]&m[552])|(m[102]&m[225]&m[552]));
    m[357] = (((~m[102]&~m[239]&~m[553])|(m[102]&m[239]&~m[553]))&BiasedRNG[429])|(((m[102]&~m[239]&~m[553])|(~m[102]&m[239]&m[553]))&~BiasedRNG[429])|((~m[102]&~m[239]&m[553])|(m[102]&~m[239]&m[553])|(m[102]&m[239]&m[553]));
    m[358] = (((~m[102]&~m[253]&~m[554])|(m[102]&m[253]&~m[554]))&BiasedRNG[430])|(((m[102]&~m[253]&~m[554])|(~m[102]&m[253]&m[554]))&~BiasedRNG[430])|((~m[102]&~m[253]&m[554])|(m[102]&~m[253]&m[554])|(m[102]&m[253]&m[554]));
    m[359] = (((~m[102]&~m[267]&~m[555])|(m[102]&m[267]&~m[555]))&BiasedRNG[431])|(((m[102]&~m[267]&~m[555])|(~m[102]&m[267]&m[555]))&~BiasedRNG[431])|((~m[102]&~m[267]&m[555])|(m[102]&~m[267]&m[555])|(m[102]&m[267]&m[555]));
    m[360] = (((~m[103]&~m[281]&~m[556])|(m[103]&m[281]&~m[556]))&BiasedRNG[432])|(((m[103]&~m[281]&~m[556])|(~m[103]&m[281]&m[556]))&~BiasedRNG[432])|((~m[103]&~m[281]&m[556])|(m[103]&~m[281]&m[556])|(m[103]&m[281]&m[556]));
    m[361] = (((~m[103]&~m[295]&~m[557])|(m[103]&m[295]&~m[557]))&BiasedRNG[433])|(((m[103]&~m[295]&~m[557])|(~m[103]&m[295]&m[557]))&~BiasedRNG[433])|((~m[103]&~m[295]&m[557])|(m[103]&~m[295]&m[557])|(m[103]&m[295]&m[557]));
    m[362] = (((~m[103]&~m[309]&~m[558])|(m[103]&m[309]&~m[558]))&BiasedRNG[434])|(((m[103]&~m[309]&~m[558])|(~m[103]&m[309]&m[558]))&~BiasedRNG[434])|((~m[103]&~m[309]&m[558])|(m[103]&~m[309]&m[558])|(m[103]&m[309]&m[558]));
    m[363] = (((~m[103]&~m[323]&~m[559])|(m[103]&m[323]&~m[559]))&BiasedRNG[435])|(((m[103]&~m[323]&~m[559])|(~m[103]&m[323]&m[559]))&~BiasedRNG[435])|((~m[103]&~m[323]&m[559])|(m[103]&~m[323]&m[559])|(m[103]&m[323]&m[559]));
    m[370] = (((~m[105]&~m[226]&~m[566])|(m[105]&m[226]&~m[566]))&BiasedRNG[436])|(((m[105]&~m[226]&~m[566])|(~m[105]&m[226]&m[566]))&~BiasedRNG[436])|((~m[105]&~m[226]&m[566])|(m[105]&~m[226]&m[566])|(m[105]&m[226]&m[566]));
    m[371] = (((~m[105]&~m[240]&~m[567])|(m[105]&m[240]&~m[567]))&BiasedRNG[437])|(((m[105]&~m[240]&~m[567])|(~m[105]&m[240]&m[567]))&~BiasedRNG[437])|((~m[105]&~m[240]&m[567])|(m[105]&~m[240]&m[567])|(m[105]&m[240]&m[567]));
    m[372] = (((~m[105]&~m[254]&~m[568])|(m[105]&m[254]&~m[568]))&BiasedRNG[438])|(((m[105]&~m[254]&~m[568])|(~m[105]&m[254]&m[568]))&~BiasedRNG[438])|((~m[105]&~m[254]&m[568])|(m[105]&~m[254]&m[568])|(m[105]&m[254]&m[568]));
    m[373] = (((~m[105]&~m[268]&~m[569])|(m[105]&m[268]&~m[569]))&BiasedRNG[439])|(((m[105]&~m[268]&~m[569])|(~m[105]&m[268]&m[569]))&~BiasedRNG[439])|((~m[105]&~m[268]&m[569])|(m[105]&~m[268]&m[569])|(m[105]&m[268]&m[569]));
    m[374] = (((~m[106]&~m[282]&~m[570])|(m[106]&m[282]&~m[570]))&BiasedRNG[440])|(((m[106]&~m[282]&~m[570])|(~m[106]&m[282]&m[570]))&~BiasedRNG[440])|((~m[106]&~m[282]&m[570])|(m[106]&~m[282]&m[570])|(m[106]&m[282]&m[570]));
    m[375] = (((~m[106]&~m[296]&~m[571])|(m[106]&m[296]&~m[571]))&BiasedRNG[441])|(((m[106]&~m[296]&~m[571])|(~m[106]&m[296]&m[571]))&~BiasedRNG[441])|((~m[106]&~m[296]&m[571])|(m[106]&~m[296]&m[571])|(m[106]&m[296]&m[571]));
    m[376] = (((~m[106]&~m[310]&~m[572])|(m[106]&m[310]&~m[572]))&BiasedRNG[442])|(((m[106]&~m[310]&~m[572])|(~m[106]&m[310]&m[572]))&~BiasedRNG[442])|((~m[106]&~m[310]&m[572])|(m[106]&~m[310]&m[572])|(m[106]&m[310]&m[572]));
    m[377] = (((~m[106]&~m[324]&~m[573])|(m[106]&m[324]&~m[573]))&BiasedRNG[443])|(((m[106]&~m[324]&~m[573])|(~m[106]&m[324]&m[573]))&~BiasedRNG[443])|((~m[106]&~m[324]&m[573])|(m[106]&~m[324]&m[573])|(m[106]&m[324]&m[573]));
    m[384] = (((~m[108]&~m[227]&~m[580])|(m[108]&m[227]&~m[580]))&BiasedRNG[444])|(((m[108]&~m[227]&~m[580])|(~m[108]&m[227]&m[580]))&~BiasedRNG[444])|((~m[108]&~m[227]&m[580])|(m[108]&~m[227]&m[580])|(m[108]&m[227]&m[580]));
    m[385] = (((~m[108]&~m[241]&~m[581])|(m[108]&m[241]&~m[581]))&BiasedRNG[445])|(((m[108]&~m[241]&~m[581])|(~m[108]&m[241]&m[581]))&~BiasedRNG[445])|((~m[108]&~m[241]&m[581])|(m[108]&~m[241]&m[581])|(m[108]&m[241]&m[581]));
    m[386] = (((~m[108]&~m[255]&~m[582])|(m[108]&m[255]&~m[582]))&BiasedRNG[446])|(((m[108]&~m[255]&~m[582])|(~m[108]&m[255]&m[582]))&~BiasedRNG[446])|((~m[108]&~m[255]&m[582])|(m[108]&~m[255]&m[582])|(m[108]&m[255]&m[582]));
    m[387] = (((~m[108]&~m[269]&~m[583])|(m[108]&m[269]&~m[583]))&BiasedRNG[447])|(((m[108]&~m[269]&~m[583])|(~m[108]&m[269]&m[583]))&~BiasedRNG[447])|((~m[108]&~m[269]&m[583])|(m[108]&~m[269]&m[583])|(m[108]&m[269]&m[583]));
    m[388] = (((~m[109]&~m[283]&~m[584])|(m[109]&m[283]&~m[584]))&BiasedRNG[448])|(((m[109]&~m[283]&~m[584])|(~m[109]&m[283]&m[584]))&~BiasedRNG[448])|((~m[109]&~m[283]&m[584])|(m[109]&~m[283]&m[584])|(m[109]&m[283]&m[584]));
    m[389] = (((~m[109]&~m[297]&~m[585])|(m[109]&m[297]&~m[585]))&BiasedRNG[449])|(((m[109]&~m[297]&~m[585])|(~m[109]&m[297]&m[585]))&~BiasedRNG[449])|((~m[109]&~m[297]&m[585])|(m[109]&~m[297]&m[585])|(m[109]&m[297]&m[585]));
    m[390] = (((~m[109]&~m[311]&~m[586])|(m[109]&m[311]&~m[586]))&BiasedRNG[450])|(((m[109]&~m[311]&~m[586])|(~m[109]&m[311]&m[586]))&~BiasedRNG[450])|((~m[109]&~m[311]&m[586])|(m[109]&~m[311]&m[586])|(m[109]&m[311]&m[586]));
    m[391] = (((~m[109]&~m[325]&~m[587])|(m[109]&m[325]&~m[587]))&BiasedRNG[451])|(((m[109]&~m[325]&~m[587])|(~m[109]&m[325]&m[587]))&~BiasedRNG[451])|((~m[109]&~m[325]&m[587])|(m[109]&~m[325]&m[587])|(m[109]&m[325]&m[587]));
    m[398] = (((~m[111]&~m[228]&~m[594])|(m[111]&m[228]&~m[594]))&BiasedRNG[452])|(((m[111]&~m[228]&~m[594])|(~m[111]&m[228]&m[594]))&~BiasedRNG[452])|((~m[111]&~m[228]&m[594])|(m[111]&~m[228]&m[594])|(m[111]&m[228]&m[594]));
    m[399] = (((~m[111]&~m[242]&~m[595])|(m[111]&m[242]&~m[595]))&BiasedRNG[453])|(((m[111]&~m[242]&~m[595])|(~m[111]&m[242]&m[595]))&~BiasedRNG[453])|((~m[111]&~m[242]&m[595])|(m[111]&~m[242]&m[595])|(m[111]&m[242]&m[595]));
    m[400] = (((~m[111]&~m[256]&~m[596])|(m[111]&m[256]&~m[596]))&BiasedRNG[454])|(((m[111]&~m[256]&~m[596])|(~m[111]&m[256]&m[596]))&~BiasedRNG[454])|((~m[111]&~m[256]&m[596])|(m[111]&~m[256]&m[596])|(m[111]&m[256]&m[596]));
    m[401] = (((~m[111]&~m[270]&~m[597])|(m[111]&m[270]&~m[597]))&BiasedRNG[455])|(((m[111]&~m[270]&~m[597])|(~m[111]&m[270]&m[597]))&~BiasedRNG[455])|((~m[111]&~m[270]&m[597])|(m[111]&~m[270]&m[597])|(m[111]&m[270]&m[597]));
    m[402] = (((~m[112]&~m[284]&~m[598])|(m[112]&m[284]&~m[598]))&BiasedRNG[456])|(((m[112]&~m[284]&~m[598])|(~m[112]&m[284]&m[598]))&~BiasedRNG[456])|((~m[112]&~m[284]&m[598])|(m[112]&~m[284]&m[598])|(m[112]&m[284]&m[598]));
    m[403] = (((~m[112]&~m[298]&~m[599])|(m[112]&m[298]&~m[599]))&BiasedRNG[457])|(((m[112]&~m[298]&~m[599])|(~m[112]&m[298]&m[599]))&~BiasedRNG[457])|((~m[112]&~m[298]&m[599])|(m[112]&~m[298]&m[599])|(m[112]&m[298]&m[599]));
    m[404] = (((~m[112]&~m[312]&~m[600])|(m[112]&m[312]&~m[600]))&BiasedRNG[458])|(((m[112]&~m[312]&~m[600])|(~m[112]&m[312]&m[600]))&~BiasedRNG[458])|((~m[112]&~m[312]&m[600])|(m[112]&~m[312]&m[600])|(m[112]&m[312]&m[600]));
    m[405] = (((~m[112]&~m[326]&~m[601])|(m[112]&m[326]&~m[601]))&BiasedRNG[459])|(((m[112]&~m[326]&~m[601])|(~m[112]&m[326]&m[601]))&~BiasedRNG[459])|((~m[112]&~m[326]&m[601])|(m[112]&~m[326]&m[601])|(m[112]&m[326]&m[601]));
    m[412] = (((~m[114]&~m[229]&~m[608])|(m[114]&m[229]&~m[608]))&BiasedRNG[460])|(((m[114]&~m[229]&~m[608])|(~m[114]&m[229]&m[608]))&~BiasedRNG[460])|((~m[114]&~m[229]&m[608])|(m[114]&~m[229]&m[608])|(m[114]&m[229]&m[608]));
    m[413] = (((~m[114]&~m[243]&~m[609])|(m[114]&m[243]&~m[609]))&BiasedRNG[461])|(((m[114]&~m[243]&~m[609])|(~m[114]&m[243]&m[609]))&~BiasedRNG[461])|((~m[114]&~m[243]&m[609])|(m[114]&~m[243]&m[609])|(m[114]&m[243]&m[609]));
    m[414] = (((~m[114]&~m[257]&~m[610])|(m[114]&m[257]&~m[610]))&BiasedRNG[462])|(((m[114]&~m[257]&~m[610])|(~m[114]&m[257]&m[610]))&~BiasedRNG[462])|((~m[114]&~m[257]&m[610])|(m[114]&~m[257]&m[610])|(m[114]&m[257]&m[610]));
    m[415] = (((~m[114]&~m[271]&~m[611])|(m[114]&m[271]&~m[611]))&BiasedRNG[463])|(((m[114]&~m[271]&~m[611])|(~m[114]&m[271]&m[611]))&~BiasedRNG[463])|((~m[114]&~m[271]&m[611])|(m[114]&~m[271]&m[611])|(m[114]&m[271]&m[611]));
    m[416] = (((~m[115]&~m[285]&~m[612])|(m[115]&m[285]&~m[612]))&BiasedRNG[464])|(((m[115]&~m[285]&~m[612])|(~m[115]&m[285]&m[612]))&~BiasedRNG[464])|((~m[115]&~m[285]&m[612])|(m[115]&~m[285]&m[612])|(m[115]&m[285]&m[612]));
    m[417] = (((~m[115]&~m[299]&~m[613])|(m[115]&m[299]&~m[613]))&BiasedRNG[465])|(((m[115]&~m[299]&~m[613])|(~m[115]&m[299]&m[613]))&~BiasedRNG[465])|((~m[115]&~m[299]&m[613])|(m[115]&~m[299]&m[613])|(m[115]&m[299]&m[613]));
    m[418] = (((~m[115]&~m[313]&~m[614])|(m[115]&m[313]&~m[614]))&BiasedRNG[466])|(((m[115]&~m[313]&~m[614])|(~m[115]&m[313]&m[614]))&~BiasedRNG[466])|((~m[115]&~m[313]&m[614])|(m[115]&~m[313]&m[614])|(m[115]&m[313]&m[614]));
    m[419] = (((~m[115]&~m[327]&~m[615])|(m[115]&m[327]&~m[615]))&BiasedRNG[467])|(((m[115]&~m[327]&~m[615])|(~m[115]&m[327]&m[615]))&~BiasedRNG[467])|((~m[115]&~m[327]&m[615])|(m[115]&~m[327]&m[615])|(m[115]&m[327]&m[615]));
    m[533] = (((m[154]&~m[337]&m[728])|(~m[154]&m[337]&m[728]))&BiasedRNG[468])|(((m[154]&m[337]&~m[728]))&~BiasedRNG[468])|((m[154]&m[337]&m[728]));
    m[534] = (((m[168]&~m[338]&m[733])|(~m[168]&m[338]&m[733]))&BiasedRNG[469])|(((m[168]&m[338]&~m[733]))&~BiasedRNG[469])|((m[168]&m[338]&m[733]));
    m[535] = (((m[182]&~m[339]&m[743])|(~m[182]&m[339]&m[743]))&BiasedRNG[470])|(((m[182]&m[339]&~m[743]))&~BiasedRNG[470])|((m[182]&m[339]&m[743]));
    m[536] = (((m[196]&~m[340]&m[758])|(~m[196]&m[340]&m[758]))&BiasedRNG[471])|(((m[196]&m[340]&~m[758]))&~BiasedRNG[471])|((m[196]&m[340]&m[758]));
    m[537] = (((m[210]&~m[341]&m[778])|(~m[210]&m[341]&m[778]))&BiasedRNG[472])|(((m[210]&m[341]&~m[778]))&~BiasedRNG[472])|((m[210]&m[341]&m[778]));
    m[546] = (((m[141]&~m[350]&m[729])|(~m[141]&m[350]&m[729]))&BiasedRNG[473])|(((m[141]&m[350]&~m[729]))&~BiasedRNG[473])|((m[141]&m[350]&m[729]));
    m[547] = (((m[155]&~m[351]&m[734])|(~m[155]&m[351]&m[734]))&BiasedRNG[474])|(((m[155]&m[351]&~m[734]))&~BiasedRNG[474])|((m[155]&m[351]&m[734]));
    m[548] = (((m[169]&~m[352]&m[744])|(~m[169]&m[352]&m[744]))&BiasedRNG[475])|(((m[169]&m[352]&~m[744]))&~BiasedRNG[475])|((m[169]&m[352]&m[744]));
    m[549] = (((m[183]&~m[353]&m[759])|(~m[183]&m[353]&m[759]))&BiasedRNG[476])|(((m[183]&m[353]&~m[759]))&~BiasedRNG[476])|((m[183]&m[353]&m[759]));
    m[550] = (((m[197]&~m[354]&m[779])|(~m[197]&m[354]&m[779]))&BiasedRNG[477])|(((m[197]&m[354]&~m[779]))&~BiasedRNG[477])|((m[197]&m[354]&m[779]));
    m[551] = (((m[211]&~m[355]&m[804])|(~m[211]&m[355]&m[804]))&BiasedRNG[478])|(((m[211]&m[355]&~m[804]))&~BiasedRNG[478])|((m[211]&m[355]&m[804]));
    m[560] = (((m[142]&~m[364]&m[739])|(~m[142]&m[364]&m[739]))&BiasedRNG[479])|(((m[142]&m[364]&~m[739]))&~BiasedRNG[479])|((m[142]&m[364]&m[739]));
    m[561] = (((m[156]&~m[365]&m[749])|(~m[156]&m[365]&m[749]))&BiasedRNG[480])|(((m[156]&m[365]&~m[749]))&~BiasedRNG[480])|((m[156]&m[365]&m[749]));
    m[562] = (((m[170]&~m[366]&m[764])|(~m[170]&m[366]&m[764]))&BiasedRNG[481])|(((m[170]&m[366]&~m[764]))&~BiasedRNG[481])|((m[170]&m[366]&m[764]));
    m[563] = (((m[184]&~m[367]&m[784])|(~m[184]&m[367]&m[784]))&BiasedRNG[482])|(((m[184]&m[367]&~m[784]))&~BiasedRNG[482])|((m[184]&m[367]&m[784]));
    m[564] = (((m[198]&~m[368]&m[809])|(~m[198]&m[368]&m[809]))&BiasedRNG[483])|(((m[198]&m[368]&~m[809]))&~BiasedRNG[483])|((m[198]&m[368]&m[809]));
    m[565] = (((m[212]&~m[369]&m[839])|(~m[212]&m[369]&m[839]))&BiasedRNG[484])|(((m[212]&m[369]&~m[839]))&~BiasedRNG[484])|((m[212]&m[369]&m[839]));
    m[574] = (((m[143]&~m[378]&m[754])|(~m[143]&m[378]&m[754]))&BiasedRNG[485])|(((m[143]&m[378]&~m[754]))&~BiasedRNG[485])|((m[143]&m[378]&m[754]));
    m[575] = (((m[157]&~m[379]&m[769])|(~m[157]&m[379]&m[769]))&BiasedRNG[486])|(((m[157]&m[379]&~m[769]))&~BiasedRNG[486])|((m[157]&m[379]&m[769]));
    m[576] = (((m[171]&~m[380]&m[789])|(~m[171]&m[380]&m[789]))&BiasedRNG[487])|(((m[171]&m[380]&~m[789]))&~BiasedRNG[487])|((m[171]&m[380]&m[789]));
    m[577] = (((m[185]&~m[381]&m[814])|(~m[185]&m[381]&m[814]))&BiasedRNG[488])|(((m[185]&m[381]&~m[814]))&~BiasedRNG[488])|((m[185]&m[381]&m[814]));
    m[578] = (((m[199]&~m[382]&m[844])|(~m[199]&m[382]&m[844]))&BiasedRNG[489])|(((m[199]&m[382]&~m[844]))&~BiasedRNG[489])|((m[199]&m[382]&m[844]));
    m[579] = (((m[213]&~m[383]&m[879])|(~m[213]&m[383]&m[879]))&BiasedRNG[490])|(((m[213]&m[383]&~m[879]))&~BiasedRNG[490])|((m[213]&m[383]&m[879]));
    m[588] = (((m[144]&~m[392]&m[774])|(~m[144]&m[392]&m[774]))&BiasedRNG[491])|(((m[144]&m[392]&~m[774]))&~BiasedRNG[491])|((m[144]&m[392]&m[774]));
    m[589] = (((m[158]&~m[393]&m[794])|(~m[158]&m[393]&m[794]))&BiasedRNG[492])|(((m[158]&m[393]&~m[794]))&~BiasedRNG[492])|((m[158]&m[393]&m[794]));
    m[590] = (((m[172]&~m[394]&m[819])|(~m[172]&m[394]&m[819]))&BiasedRNG[493])|(((m[172]&m[394]&~m[819]))&~BiasedRNG[493])|((m[172]&m[394]&m[819]));
    m[591] = (((m[186]&~m[395]&m[849])|(~m[186]&m[395]&m[849]))&BiasedRNG[494])|(((m[186]&m[395]&~m[849]))&~BiasedRNG[494])|((m[186]&m[395]&m[849]));
    m[592] = (((m[200]&~m[396]&m[884])|(~m[200]&m[396]&m[884]))&BiasedRNG[495])|(((m[200]&m[396]&~m[884]))&~BiasedRNG[495])|((m[200]&m[396]&m[884]));
    m[593] = (((m[214]&~m[397]&m[924])|(~m[214]&m[397]&m[924]))&BiasedRNG[496])|(((m[214]&m[397]&~m[924]))&~BiasedRNG[496])|((m[214]&m[397]&m[924]));
    m[602] = (((m[145]&~m[406]&m[799])|(~m[145]&m[406]&m[799]))&BiasedRNG[497])|(((m[145]&m[406]&~m[799]))&~BiasedRNG[497])|((m[145]&m[406]&m[799]));
    m[603] = (((m[159]&~m[407]&m[824])|(~m[159]&m[407]&m[824]))&BiasedRNG[498])|(((m[159]&m[407]&~m[824]))&~BiasedRNG[498])|((m[159]&m[407]&m[824]));
    m[604] = (((m[173]&~m[408]&m[854])|(~m[173]&m[408]&m[854]))&BiasedRNG[499])|(((m[173]&m[408]&~m[854]))&~BiasedRNG[499])|((m[173]&m[408]&m[854]));
    m[605] = (((m[187]&~m[409]&m[889])|(~m[187]&m[409]&m[889]))&BiasedRNG[500])|(((m[187]&m[409]&~m[889]))&~BiasedRNG[500])|((m[187]&m[409]&m[889]));
    m[606] = (((m[201]&~m[410]&m[929])|(~m[201]&m[410]&m[929]))&BiasedRNG[501])|(((m[201]&m[410]&~m[929]))&~BiasedRNG[501])|((m[201]&m[410]&m[929]));
    m[607] = (((m[215]&~m[411]&m[974])|(~m[215]&m[411]&m[974]))&BiasedRNG[502])|(((m[215]&m[411]&~m[974]))&~BiasedRNG[502])|((m[215]&m[411]&m[974]));
    m[735] = (((m[732]&~m[733]&~m[734]&~m[736]&~m[737])|(~m[732]&~m[733]&~m[734]&m[736]&~m[737])|(m[732]&m[733]&~m[734]&m[736]&~m[737])|(m[732]&~m[733]&m[734]&m[736]&~m[737])|(~m[732]&m[733]&~m[734]&~m[736]&m[737])|(~m[732]&~m[733]&m[734]&~m[736]&m[737])|(m[732]&m[733]&m[734]&~m[736]&m[737])|(~m[732]&m[733]&m[734]&m[736]&m[737]))&UnbiasedRNG[209])|((m[732]&~m[733]&~m[734]&m[736]&~m[737])|(~m[732]&~m[733]&~m[734]&~m[736]&m[737])|(m[732]&~m[733]&~m[734]&~m[736]&m[737])|(m[732]&m[733]&~m[734]&~m[736]&m[737])|(m[732]&~m[733]&m[734]&~m[736]&m[737])|(~m[732]&~m[733]&~m[734]&m[736]&m[737])|(m[732]&~m[733]&~m[734]&m[736]&m[737])|(~m[732]&m[733]&~m[734]&m[736]&m[737])|(m[732]&m[733]&~m[734]&m[736]&m[737])|(~m[732]&~m[733]&m[734]&m[736]&m[737])|(m[732]&~m[733]&m[734]&m[736]&m[737])|(m[732]&m[733]&m[734]&m[736]&m[737]));
    m[745] = (((m[737]&~m[743]&~m[744]&~m[746]&~m[747])|(~m[737]&~m[743]&~m[744]&m[746]&~m[747])|(m[737]&m[743]&~m[744]&m[746]&~m[747])|(m[737]&~m[743]&m[744]&m[746]&~m[747])|(~m[737]&m[743]&~m[744]&~m[746]&m[747])|(~m[737]&~m[743]&m[744]&~m[746]&m[747])|(m[737]&m[743]&m[744]&~m[746]&m[747])|(~m[737]&m[743]&m[744]&m[746]&m[747]))&UnbiasedRNG[210])|((m[737]&~m[743]&~m[744]&m[746]&~m[747])|(~m[737]&~m[743]&~m[744]&~m[746]&m[747])|(m[737]&~m[743]&~m[744]&~m[746]&m[747])|(m[737]&m[743]&~m[744]&~m[746]&m[747])|(m[737]&~m[743]&m[744]&~m[746]&m[747])|(~m[737]&~m[743]&~m[744]&m[746]&m[747])|(m[737]&~m[743]&~m[744]&m[746]&m[747])|(~m[737]&m[743]&~m[744]&m[746]&m[747])|(m[737]&m[743]&~m[744]&m[746]&m[747])|(~m[737]&~m[743]&m[744]&m[746]&m[747])|(m[737]&~m[743]&m[744]&m[746]&m[747])|(m[737]&m[743]&m[744]&m[746]&m[747]));
    m[750] = (((m[742]&~m[748]&~m[749]&~m[751]&~m[752])|(~m[742]&~m[748]&~m[749]&m[751]&~m[752])|(m[742]&m[748]&~m[749]&m[751]&~m[752])|(m[742]&~m[748]&m[749]&m[751]&~m[752])|(~m[742]&m[748]&~m[749]&~m[751]&m[752])|(~m[742]&~m[748]&m[749]&~m[751]&m[752])|(m[742]&m[748]&m[749]&~m[751]&m[752])|(~m[742]&m[748]&m[749]&m[751]&m[752]))&UnbiasedRNG[211])|((m[742]&~m[748]&~m[749]&m[751]&~m[752])|(~m[742]&~m[748]&~m[749]&~m[751]&m[752])|(m[742]&~m[748]&~m[749]&~m[751]&m[752])|(m[742]&m[748]&~m[749]&~m[751]&m[752])|(m[742]&~m[748]&m[749]&~m[751]&m[752])|(~m[742]&~m[748]&~m[749]&m[751]&m[752])|(m[742]&~m[748]&~m[749]&m[751]&m[752])|(~m[742]&m[748]&~m[749]&m[751]&m[752])|(m[742]&m[748]&~m[749]&m[751]&m[752])|(~m[742]&~m[748]&m[749]&m[751]&m[752])|(m[742]&~m[748]&m[749]&m[751]&m[752])|(m[742]&m[748]&m[749]&m[751]&m[752]));
    m[760] = (((m[747]&~m[758]&~m[759]&~m[761]&~m[762])|(~m[747]&~m[758]&~m[759]&m[761]&~m[762])|(m[747]&m[758]&~m[759]&m[761]&~m[762])|(m[747]&~m[758]&m[759]&m[761]&~m[762])|(~m[747]&m[758]&~m[759]&~m[761]&m[762])|(~m[747]&~m[758]&m[759]&~m[761]&m[762])|(m[747]&m[758]&m[759]&~m[761]&m[762])|(~m[747]&m[758]&m[759]&m[761]&m[762]))&UnbiasedRNG[212])|((m[747]&~m[758]&~m[759]&m[761]&~m[762])|(~m[747]&~m[758]&~m[759]&~m[761]&m[762])|(m[747]&~m[758]&~m[759]&~m[761]&m[762])|(m[747]&m[758]&~m[759]&~m[761]&m[762])|(m[747]&~m[758]&m[759]&~m[761]&m[762])|(~m[747]&~m[758]&~m[759]&m[761]&m[762])|(m[747]&~m[758]&~m[759]&m[761]&m[762])|(~m[747]&m[758]&~m[759]&m[761]&m[762])|(m[747]&m[758]&~m[759]&m[761]&m[762])|(~m[747]&~m[758]&m[759]&m[761]&m[762])|(m[747]&~m[758]&m[759]&m[761]&m[762])|(m[747]&m[758]&m[759]&m[761]&m[762]));
    m[765] = (((m[752]&~m[763]&~m[764]&~m[766]&~m[767])|(~m[752]&~m[763]&~m[764]&m[766]&~m[767])|(m[752]&m[763]&~m[764]&m[766]&~m[767])|(m[752]&~m[763]&m[764]&m[766]&~m[767])|(~m[752]&m[763]&~m[764]&~m[766]&m[767])|(~m[752]&~m[763]&m[764]&~m[766]&m[767])|(m[752]&m[763]&m[764]&~m[766]&m[767])|(~m[752]&m[763]&m[764]&m[766]&m[767]))&UnbiasedRNG[213])|((m[752]&~m[763]&~m[764]&m[766]&~m[767])|(~m[752]&~m[763]&~m[764]&~m[766]&m[767])|(m[752]&~m[763]&~m[764]&~m[766]&m[767])|(m[752]&m[763]&~m[764]&~m[766]&m[767])|(m[752]&~m[763]&m[764]&~m[766]&m[767])|(~m[752]&~m[763]&~m[764]&m[766]&m[767])|(m[752]&~m[763]&~m[764]&m[766]&m[767])|(~m[752]&m[763]&~m[764]&m[766]&m[767])|(m[752]&m[763]&~m[764]&m[766]&m[767])|(~m[752]&~m[763]&m[764]&m[766]&m[767])|(m[752]&~m[763]&m[764]&m[766]&m[767])|(m[752]&m[763]&m[764]&m[766]&m[767]));
    m[770] = (((m[757]&~m[768]&~m[769]&~m[771]&~m[772])|(~m[757]&~m[768]&~m[769]&m[771]&~m[772])|(m[757]&m[768]&~m[769]&m[771]&~m[772])|(m[757]&~m[768]&m[769]&m[771]&~m[772])|(~m[757]&m[768]&~m[769]&~m[771]&m[772])|(~m[757]&~m[768]&m[769]&~m[771]&m[772])|(m[757]&m[768]&m[769]&~m[771]&m[772])|(~m[757]&m[768]&m[769]&m[771]&m[772]))&UnbiasedRNG[214])|((m[757]&~m[768]&~m[769]&m[771]&~m[772])|(~m[757]&~m[768]&~m[769]&~m[771]&m[772])|(m[757]&~m[768]&~m[769]&~m[771]&m[772])|(m[757]&m[768]&~m[769]&~m[771]&m[772])|(m[757]&~m[768]&m[769]&~m[771]&m[772])|(~m[757]&~m[768]&~m[769]&m[771]&m[772])|(m[757]&~m[768]&~m[769]&m[771]&m[772])|(~m[757]&m[768]&~m[769]&m[771]&m[772])|(m[757]&m[768]&~m[769]&m[771]&m[772])|(~m[757]&~m[768]&m[769]&m[771]&m[772])|(m[757]&~m[768]&m[769]&m[771]&m[772])|(m[757]&m[768]&m[769]&m[771]&m[772]));
    m[780] = (((m[762]&~m[778]&~m[779]&~m[781]&~m[782])|(~m[762]&~m[778]&~m[779]&m[781]&~m[782])|(m[762]&m[778]&~m[779]&m[781]&~m[782])|(m[762]&~m[778]&m[779]&m[781]&~m[782])|(~m[762]&m[778]&~m[779]&~m[781]&m[782])|(~m[762]&~m[778]&m[779]&~m[781]&m[782])|(m[762]&m[778]&m[779]&~m[781]&m[782])|(~m[762]&m[778]&m[779]&m[781]&m[782]))&UnbiasedRNG[215])|((m[762]&~m[778]&~m[779]&m[781]&~m[782])|(~m[762]&~m[778]&~m[779]&~m[781]&m[782])|(m[762]&~m[778]&~m[779]&~m[781]&m[782])|(m[762]&m[778]&~m[779]&~m[781]&m[782])|(m[762]&~m[778]&m[779]&~m[781]&m[782])|(~m[762]&~m[778]&~m[779]&m[781]&m[782])|(m[762]&~m[778]&~m[779]&m[781]&m[782])|(~m[762]&m[778]&~m[779]&m[781]&m[782])|(m[762]&m[778]&~m[779]&m[781]&m[782])|(~m[762]&~m[778]&m[779]&m[781]&m[782])|(m[762]&~m[778]&m[779]&m[781]&m[782])|(m[762]&m[778]&m[779]&m[781]&m[782]));
    m[785] = (((m[767]&~m[783]&~m[784]&~m[786]&~m[787])|(~m[767]&~m[783]&~m[784]&m[786]&~m[787])|(m[767]&m[783]&~m[784]&m[786]&~m[787])|(m[767]&~m[783]&m[784]&m[786]&~m[787])|(~m[767]&m[783]&~m[784]&~m[786]&m[787])|(~m[767]&~m[783]&m[784]&~m[786]&m[787])|(m[767]&m[783]&m[784]&~m[786]&m[787])|(~m[767]&m[783]&m[784]&m[786]&m[787]))&UnbiasedRNG[216])|((m[767]&~m[783]&~m[784]&m[786]&~m[787])|(~m[767]&~m[783]&~m[784]&~m[786]&m[787])|(m[767]&~m[783]&~m[784]&~m[786]&m[787])|(m[767]&m[783]&~m[784]&~m[786]&m[787])|(m[767]&~m[783]&m[784]&~m[786]&m[787])|(~m[767]&~m[783]&~m[784]&m[786]&m[787])|(m[767]&~m[783]&~m[784]&m[786]&m[787])|(~m[767]&m[783]&~m[784]&m[786]&m[787])|(m[767]&m[783]&~m[784]&m[786]&m[787])|(~m[767]&~m[783]&m[784]&m[786]&m[787])|(m[767]&~m[783]&m[784]&m[786]&m[787])|(m[767]&m[783]&m[784]&m[786]&m[787]));
    m[790] = (((m[772]&~m[788]&~m[789]&~m[791]&~m[792])|(~m[772]&~m[788]&~m[789]&m[791]&~m[792])|(m[772]&m[788]&~m[789]&m[791]&~m[792])|(m[772]&~m[788]&m[789]&m[791]&~m[792])|(~m[772]&m[788]&~m[789]&~m[791]&m[792])|(~m[772]&~m[788]&m[789]&~m[791]&m[792])|(m[772]&m[788]&m[789]&~m[791]&m[792])|(~m[772]&m[788]&m[789]&m[791]&m[792]))&UnbiasedRNG[217])|((m[772]&~m[788]&~m[789]&m[791]&~m[792])|(~m[772]&~m[788]&~m[789]&~m[791]&m[792])|(m[772]&~m[788]&~m[789]&~m[791]&m[792])|(m[772]&m[788]&~m[789]&~m[791]&m[792])|(m[772]&~m[788]&m[789]&~m[791]&m[792])|(~m[772]&~m[788]&~m[789]&m[791]&m[792])|(m[772]&~m[788]&~m[789]&m[791]&m[792])|(~m[772]&m[788]&~m[789]&m[791]&m[792])|(m[772]&m[788]&~m[789]&m[791]&m[792])|(~m[772]&~m[788]&m[789]&m[791]&m[792])|(m[772]&~m[788]&m[789]&m[791]&m[792])|(m[772]&m[788]&m[789]&m[791]&m[792]));
    m[795] = (((m[777]&~m[793]&~m[794]&~m[796]&~m[797])|(~m[777]&~m[793]&~m[794]&m[796]&~m[797])|(m[777]&m[793]&~m[794]&m[796]&~m[797])|(m[777]&~m[793]&m[794]&m[796]&~m[797])|(~m[777]&m[793]&~m[794]&~m[796]&m[797])|(~m[777]&~m[793]&m[794]&~m[796]&m[797])|(m[777]&m[793]&m[794]&~m[796]&m[797])|(~m[777]&m[793]&m[794]&m[796]&m[797]))&UnbiasedRNG[218])|((m[777]&~m[793]&~m[794]&m[796]&~m[797])|(~m[777]&~m[793]&~m[794]&~m[796]&m[797])|(m[777]&~m[793]&~m[794]&~m[796]&m[797])|(m[777]&m[793]&~m[794]&~m[796]&m[797])|(m[777]&~m[793]&m[794]&~m[796]&m[797])|(~m[777]&~m[793]&~m[794]&m[796]&m[797])|(m[777]&~m[793]&~m[794]&m[796]&m[797])|(~m[777]&m[793]&~m[794]&m[796]&m[797])|(m[777]&m[793]&~m[794]&m[796]&m[797])|(~m[777]&~m[793]&m[794]&m[796]&m[797])|(m[777]&~m[793]&m[794]&m[796]&m[797])|(m[777]&m[793]&m[794]&m[796]&m[797]));
    m[805] = (((m[782]&~m[803]&~m[804]&~m[806]&~m[807])|(~m[782]&~m[803]&~m[804]&m[806]&~m[807])|(m[782]&m[803]&~m[804]&m[806]&~m[807])|(m[782]&~m[803]&m[804]&m[806]&~m[807])|(~m[782]&m[803]&~m[804]&~m[806]&m[807])|(~m[782]&~m[803]&m[804]&~m[806]&m[807])|(m[782]&m[803]&m[804]&~m[806]&m[807])|(~m[782]&m[803]&m[804]&m[806]&m[807]))&UnbiasedRNG[219])|((m[782]&~m[803]&~m[804]&m[806]&~m[807])|(~m[782]&~m[803]&~m[804]&~m[806]&m[807])|(m[782]&~m[803]&~m[804]&~m[806]&m[807])|(m[782]&m[803]&~m[804]&~m[806]&m[807])|(m[782]&~m[803]&m[804]&~m[806]&m[807])|(~m[782]&~m[803]&~m[804]&m[806]&m[807])|(m[782]&~m[803]&~m[804]&m[806]&m[807])|(~m[782]&m[803]&~m[804]&m[806]&m[807])|(m[782]&m[803]&~m[804]&m[806]&m[807])|(~m[782]&~m[803]&m[804]&m[806]&m[807])|(m[782]&~m[803]&m[804]&m[806]&m[807])|(m[782]&m[803]&m[804]&m[806]&m[807]));
    m[810] = (((m[787]&~m[808]&~m[809]&~m[811]&~m[812])|(~m[787]&~m[808]&~m[809]&m[811]&~m[812])|(m[787]&m[808]&~m[809]&m[811]&~m[812])|(m[787]&~m[808]&m[809]&m[811]&~m[812])|(~m[787]&m[808]&~m[809]&~m[811]&m[812])|(~m[787]&~m[808]&m[809]&~m[811]&m[812])|(m[787]&m[808]&m[809]&~m[811]&m[812])|(~m[787]&m[808]&m[809]&m[811]&m[812]))&UnbiasedRNG[220])|((m[787]&~m[808]&~m[809]&m[811]&~m[812])|(~m[787]&~m[808]&~m[809]&~m[811]&m[812])|(m[787]&~m[808]&~m[809]&~m[811]&m[812])|(m[787]&m[808]&~m[809]&~m[811]&m[812])|(m[787]&~m[808]&m[809]&~m[811]&m[812])|(~m[787]&~m[808]&~m[809]&m[811]&m[812])|(m[787]&~m[808]&~m[809]&m[811]&m[812])|(~m[787]&m[808]&~m[809]&m[811]&m[812])|(m[787]&m[808]&~m[809]&m[811]&m[812])|(~m[787]&~m[808]&m[809]&m[811]&m[812])|(m[787]&~m[808]&m[809]&m[811]&m[812])|(m[787]&m[808]&m[809]&m[811]&m[812]));
    m[815] = (((m[792]&~m[813]&~m[814]&~m[816]&~m[817])|(~m[792]&~m[813]&~m[814]&m[816]&~m[817])|(m[792]&m[813]&~m[814]&m[816]&~m[817])|(m[792]&~m[813]&m[814]&m[816]&~m[817])|(~m[792]&m[813]&~m[814]&~m[816]&m[817])|(~m[792]&~m[813]&m[814]&~m[816]&m[817])|(m[792]&m[813]&m[814]&~m[816]&m[817])|(~m[792]&m[813]&m[814]&m[816]&m[817]))&UnbiasedRNG[221])|((m[792]&~m[813]&~m[814]&m[816]&~m[817])|(~m[792]&~m[813]&~m[814]&~m[816]&m[817])|(m[792]&~m[813]&~m[814]&~m[816]&m[817])|(m[792]&m[813]&~m[814]&~m[816]&m[817])|(m[792]&~m[813]&m[814]&~m[816]&m[817])|(~m[792]&~m[813]&~m[814]&m[816]&m[817])|(m[792]&~m[813]&~m[814]&m[816]&m[817])|(~m[792]&m[813]&~m[814]&m[816]&m[817])|(m[792]&m[813]&~m[814]&m[816]&m[817])|(~m[792]&~m[813]&m[814]&m[816]&m[817])|(m[792]&~m[813]&m[814]&m[816]&m[817])|(m[792]&m[813]&m[814]&m[816]&m[817]));
    m[820] = (((m[797]&~m[818]&~m[819]&~m[821]&~m[822])|(~m[797]&~m[818]&~m[819]&m[821]&~m[822])|(m[797]&m[818]&~m[819]&m[821]&~m[822])|(m[797]&~m[818]&m[819]&m[821]&~m[822])|(~m[797]&m[818]&~m[819]&~m[821]&m[822])|(~m[797]&~m[818]&m[819]&~m[821]&m[822])|(m[797]&m[818]&m[819]&~m[821]&m[822])|(~m[797]&m[818]&m[819]&m[821]&m[822]))&UnbiasedRNG[222])|((m[797]&~m[818]&~m[819]&m[821]&~m[822])|(~m[797]&~m[818]&~m[819]&~m[821]&m[822])|(m[797]&~m[818]&~m[819]&~m[821]&m[822])|(m[797]&m[818]&~m[819]&~m[821]&m[822])|(m[797]&~m[818]&m[819]&~m[821]&m[822])|(~m[797]&~m[818]&~m[819]&m[821]&m[822])|(m[797]&~m[818]&~m[819]&m[821]&m[822])|(~m[797]&m[818]&~m[819]&m[821]&m[822])|(m[797]&m[818]&~m[819]&m[821]&m[822])|(~m[797]&~m[818]&m[819]&m[821]&m[822])|(m[797]&~m[818]&m[819]&m[821]&m[822])|(m[797]&m[818]&m[819]&m[821]&m[822]));
    m[825] = (((m[802]&~m[823]&~m[824]&~m[826]&~m[827])|(~m[802]&~m[823]&~m[824]&m[826]&~m[827])|(m[802]&m[823]&~m[824]&m[826]&~m[827])|(m[802]&~m[823]&m[824]&m[826]&~m[827])|(~m[802]&m[823]&~m[824]&~m[826]&m[827])|(~m[802]&~m[823]&m[824]&~m[826]&m[827])|(m[802]&m[823]&m[824]&~m[826]&m[827])|(~m[802]&m[823]&m[824]&m[826]&m[827]))&UnbiasedRNG[223])|((m[802]&~m[823]&~m[824]&m[826]&~m[827])|(~m[802]&~m[823]&~m[824]&~m[826]&m[827])|(m[802]&~m[823]&~m[824]&~m[826]&m[827])|(m[802]&m[823]&~m[824]&~m[826]&m[827])|(m[802]&~m[823]&m[824]&~m[826]&m[827])|(~m[802]&~m[823]&~m[824]&m[826]&m[827])|(m[802]&~m[823]&~m[824]&m[826]&m[827])|(~m[802]&m[823]&~m[824]&m[826]&m[827])|(m[802]&m[823]&~m[824]&m[826]&m[827])|(~m[802]&~m[823]&m[824]&m[826]&m[827])|(m[802]&~m[823]&m[824]&m[826]&m[827])|(m[802]&m[823]&m[824]&m[826]&m[827]));
    m[829] = (((m[616]&~m[828]&~m[830]&~m[831]&~m[832])|(~m[616]&~m[828]&~m[830]&m[831]&~m[832])|(m[616]&m[828]&~m[830]&m[831]&~m[832])|(m[616]&~m[828]&m[830]&m[831]&~m[832])|(~m[616]&m[828]&~m[830]&~m[831]&m[832])|(~m[616]&~m[828]&m[830]&~m[831]&m[832])|(m[616]&m[828]&m[830]&~m[831]&m[832])|(~m[616]&m[828]&m[830]&m[831]&m[832]))&UnbiasedRNG[224])|((m[616]&~m[828]&~m[830]&m[831]&~m[832])|(~m[616]&~m[828]&~m[830]&~m[831]&m[832])|(m[616]&~m[828]&~m[830]&~m[831]&m[832])|(m[616]&m[828]&~m[830]&~m[831]&m[832])|(m[616]&~m[828]&m[830]&~m[831]&m[832])|(~m[616]&~m[828]&~m[830]&m[831]&m[832])|(m[616]&~m[828]&~m[830]&m[831]&m[832])|(~m[616]&m[828]&~m[830]&m[831]&m[832])|(m[616]&m[828]&~m[830]&m[831]&m[832])|(~m[616]&~m[828]&m[830]&m[831]&m[832])|(m[616]&~m[828]&m[830]&m[831]&m[832])|(m[616]&m[828]&m[830]&m[831]&m[832]));
    m[834] = (((m[552]&~m[833]&~m[835]&~m[836]&~m[837])|(~m[552]&~m[833]&~m[835]&m[836]&~m[837])|(m[552]&m[833]&~m[835]&m[836]&~m[837])|(m[552]&~m[833]&m[835]&m[836]&~m[837])|(~m[552]&m[833]&~m[835]&~m[836]&m[837])|(~m[552]&~m[833]&m[835]&~m[836]&m[837])|(m[552]&m[833]&m[835]&~m[836]&m[837])|(~m[552]&m[833]&m[835]&m[836]&m[837]))&UnbiasedRNG[225])|((m[552]&~m[833]&~m[835]&m[836]&~m[837])|(~m[552]&~m[833]&~m[835]&~m[836]&m[837])|(m[552]&~m[833]&~m[835]&~m[836]&m[837])|(m[552]&m[833]&~m[835]&~m[836]&m[837])|(m[552]&~m[833]&m[835]&~m[836]&m[837])|(~m[552]&~m[833]&~m[835]&m[836]&m[837])|(m[552]&~m[833]&~m[835]&m[836]&m[837])|(~m[552]&m[833]&~m[835]&m[836]&m[837])|(m[552]&m[833]&~m[835]&m[836]&m[837])|(~m[552]&~m[833]&m[835]&m[836]&m[837])|(m[552]&~m[833]&m[835]&m[836]&m[837])|(m[552]&m[833]&m[835]&m[836]&m[837]));
    m[840] = (((m[812]&~m[838]&~m[839]&~m[841]&~m[842])|(~m[812]&~m[838]&~m[839]&m[841]&~m[842])|(m[812]&m[838]&~m[839]&m[841]&~m[842])|(m[812]&~m[838]&m[839]&m[841]&~m[842])|(~m[812]&m[838]&~m[839]&~m[841]&m[842])|(~m[812]&~m[838]&m[839]&~m[841]&m[842])|(m[812]&m[838]&m[839]&~m[841]&m[842])|(~m[812]&m[838]&m[839]&m[841]&m[842]))&UnbiasedRNG[226])|((m[812]&~m[838]&~m[839]&m[841]&~m[842])|(~m[812]&~m[838]&~m[839]&~m[841]&m[842])|(m[812]&~m[838]&~m[839]&~m[841]&m[842])|(m[812]&m[838]&~m[839]&~m[841]&m[842])|(m[812]&~m[838]&m[839]&~m[841]&m[842])|(~m[812]&~m[838]&~m[839]&m[841]&m[842])|(m[812]&~m[838]&~m[839]&m[841]&m[842])|(~m[812]&m[838]&~m[839]&m[841]&m[842])|(m[812]&m[838]&~m[839]&m[841]&m[842])|(~m[812]&~m[838]&m[839]&m[841]&m[842])|(m[812]&~m[838]&m[839]&m[841]&m[842])|(m[812]&m[838]&m[839]&m[841]&m[842]));
    m[845] = (((m[817]&~m[843]&~m[844]&~m[846]&~m[847])|(~m[817]&~m[843]&~m[844]&m[846]&~m[847])|(m[817]&m[843]&~m[844]&m[846]&~m[847])|(m[817]&~m[843]&m[844]&m[846]&~m[847])|(~m[817]&m[843]&~m[844]&~m[846]&m[847])|(~m[817]&~m[843]&m[844]&~m[846]&m[847])|(m[817]&m[843]&m[844]&~m[846]&m[847])|(~m[817]&m[843]&m[844]&m[846]&m[847]))&UnbiasedRNG[227])|((m[817]&~m[843]&~m[844]&m[846]&~m[847])|(~m[817]&~m[843]&~m[844]&~m[846]&m[847])|(m[817]&~m[843]&~m[844]&~m[846]&m[847])|(m[817]&m[843]&~m[844]&~m[846]&m[847])|(m[817]&~m[843]&m[844]&~m[846]&m[847])|(~m[817]&~m[843]&~m[844]&m[846]&m[847])|(m[817]&~m[843]&~m[844]&m[846]&m[847])|(~m[817]&m[843]&~m[844]&m[846]&m[847])|(m[817]&m[843]&~m[844]&m[846]&m[847])|(~m[817]&~m[843]&m[844]&m[846]&m[847])|(m[817]&~m[843]&m[844]&m[846]&m[847])|(m[817]&m[843]&m[844]&m[846]&m[847]));
    m[850] = (((m[822]&~m[848]&~m[849]&~m[851]&~m[852])|(~m[822]&~m[848]&~m[849]&m[851]&~m[852])|(m[822]&m[848]&~m[849]&m[851]&~m[852])|(m[822]&~m[848]&m[849]&m[851]&~m[852])|(~m[822]&m[848]&~m[849]&~m[851]&m[852])|(~m[822]&~m[848]&m[849]&~m[851]&m[852])|(m[822]&m[848]&m[849]&~m[851]&m[852])|(~m[822]&m[848]&m[849]&m[851]&m[852]))&UnbiasedRNG[228])|((m[822]&~m[848]&~m[849]&m[851]&~m[852])|(~m[822]&~m[848]&~m[849]&~m[851]&m[852])|(m[822]&~m[848]&~m[849]&~m[851]&m[852])|(m[822]&m[848]&~m[849]&~m[851]&m[852])|(m[822]&~m[848]&m[849]&~m[851]&m[852])|(~m[822]&~m[848]&~m[849]&m[851]&m[852])|(m[822]&~m[848]&~m[849]&m[851]&m[852])|(~m[822]&m[848]&~m[849]&m[851]&m[852])|(m[822]&m[848]&~m[849]&m[851]&m[852])|(~m[822]&~m[848]&m[849]&m[851]&m[852])|(m[822]&~m[848]&m[849]&m[851]&m[852])|(m[822]&m[848]&m[849]&m[851]&m[852]));
    m[855] = (((m[827]&~m[853]&~m[854]&~m[856]&~m[857])|(~m[827]&~m[853]&~m[854]&m[856]&~m[857])|(m[827]&m[853]&~m[854]&m[856]&~m[857])|(m[827]&~m[853]&m[854]&m[856]&~m[857])|(~m[827]&m[853]&~m[854]&~m[856]&m[857])|(~m[827]&~m[853]&m[854]&~m[856]&m[857])|(m[827]&m[853]&m[854]&~m[856]&m[857])|(~m[827]&m[853]&m[854]&m[856]&m[857]))&UnbiasedRNG[229])|((m[827]&~m[853]&~m[854]&m[856]&~m[857])|(~m[827]&~m[853]&~m[854]&~m[856]&m[857])|(m[827]&~m[853]&~m[854]&~m[856]&m[857])|(m[827]&m[853]&~m[854]&~m[856]&m[857])|(m[827]&~m[853]&m[854]&~m[856]&m[857])|(~m[827]&~m[853]&~m[854]&m[856]&m[857])|(m[827]&~m[853]&~m[854]&m[856]&m[857])|(~m[827]&m[853]&~m[854]&m[856]&m[857])|(m[827]&m[853]&~m[854]&m[856]&m[857])|(~m[827]&~m[853]&m[854]&m[856]&m[857])|(m[827]&~m[853]&m[854]&m[856]&m[857])|(m[827]&m[853]&m[854]&m[856]&m[857]));
    m[859] = (((m[617]&~m[858]&~m[860]&~m[861]&~m[862])|(~m[617]&~m[858]&~m[860]&m[861]&~m[862])|(m[617]&m[858]&~m[860]&m[861]&~m[862])|(m[617]&~m[858]&m[860]&m[861]&~m[862])|(~m[617]&m[858]&~m[860]&~m[861]&m[862])|(~m[617]&~m[858]&m[860]&~m[861]&m[862])|(m[617]&m[858]&m[860]&~m[861]&m[862])|(~m[617]&m[858]&m[860]&m[861]&m[862]))&UnbiasedRNG[230])|((m[617]&~m[858]&~m[860]&m[861]&~m[862])|(~m[617]&~m[858]&~m[860]&~m[861]&m[862])|(m[617]&~m[858]&~m[860]&~m[861]&m[862])|(m[617]&m[858]&~m[860]&~m[861]&m[862])|(m[617]&~m[858]&m[860]&~m[861]&m[862])|(~m[617]&~m[858]&~m[860]&m[861]&m[862])|(m[617]&~m[858]&~m[860]&m[861]&m[862])|(~m[617]&m[858]&~m[860]&m[861]&m[862])|(m[617]&m[858]&~m[860]&m[861]&m[862])|(~m[617]&~m[858]&m[860]&m[861]&m[862])|(m[617]&~m[858]&m[860]&m[861]&m[862])|(m[617]&m[858]&m[860]&m[861]&m[862]));
    m[864] = (((m[630]&~m[863]&~m[865]&~m[866]&~m[867])|(~m[630]&~m[863]&~m[865]&m[866]&~m[867])|(m[630]&m[863]&~m[865]&m[866]&~m[867])|(m[630]&~m[863]&m[865]&m[866]&~m[867])|(~m[630]&m[863]&~m[865]&~m[866]&m[867])|(~m[630]&~m[863]&m[865]&~m[866]&m[867])|(m[630]&m[863]&m[865]&~m[866]&m[867])|(~m[630]&m[863]&m[865]&m[866]&m[867]))&UnbiasedRNG[231])|((m[630]&~m[863]&~m[865]&m[866]&~m[867])|(~m[630]&~m[863]&~m[865]&~m[866]&m[867])|(m[630]&~m[863]&~m[865]&~m[866]&m[867])|(m[630]&m[863]&~m[865]&~m[866]&m[867])|(m[630]&~m[863]&m[865]&~m[866]&m[867])|(~m[630]&~m[863]&~m[865]&m[866]&m[867])|(m[630]&~m[863]&~m[865]&m[866]&m[867])|(~m[630]&m[863]&~m[865]&m[866]&m[867])|(m[630]&m[863]&~m[865]&m[866]&m[867])|(~m[630]&~m[863]&m[865]&m[866]&m[867])|(m[630]&~m[863]&m[865]&m[866]&m[867])|(m[630]&m[863]&m[865]&m[866]&m[867]));
    m[869] = (((m[553]&~m[868]&~m[870]&~m[871]&~m[872])|(~m[553]&~m[868]&~m[870]&m[871]&~m[872])|(m[553]&m[868]&~m[870]&m[871]&~m[872])|(m[553]&~m[868]&m[870]&m[871]&~m[872])|(~m[553]&m[868]&~m[870]&~m[871]&m[872])|(~m[553]&~m[868]&m[870]&~m[871]&m[872])|(m[553]&m[868]&m[870]&~m[871]&m[872])|(~m[553]&m[868]&m[870]&m[871]&m[872]))&UnbiasedRNG[232])|((m[553]&~m[868]&~m[870]&m[871]&~m[872])|(~m[553]&~m[868]&~m[870]&~m[871]&m[872])|(m[553]&~m[868]&~m[870]&~m[871]&m[872])|(m[553]&m[868]&~m[870]&~m[871]&m[872])|(m[553]&~m[868]&m[870]&~m[871]&m[872])|(~m[553]&~m[868]&~m[870]&m[871]&m[872])|(m[553]&~m[868]&~m[870]&m[871]&m[872])|(~m[553]&m[868]&~m[870]&m[871]&m[872])|(m[553]&m[868]&~m[870]&m[871]&m[872])|(~m[553]&~m[868]&m[870]&m[871]&m[872])|(m[553]&~m[868]&m[870]&m[871]&m[872])|(m[553]&m[868]&m[870]&m[871]&m[872]));
    m[874] = (((m[566]&~m[873]&~m[875]&~m[876]&~m[877])|(~m[566]&~m[873]&~m[875]&m[876]&~m[877])|(m[566]&m[873]&~m[875]&m[876]&~m[877])|(m[566]&~m[873]&m[875]&m[876]&~m[877])|(~m[566]&m[873]&~m[875]&~m[876]&m[877])|(~m[566]&~m[873]&m[875]&~m[876]&m[877])|(m[566]&m[873]&m[875]&~m[876]&m[877])|(~m[566]&m[873]&m[875]&m[876]&m[877]))&UnbiasedRNG[233])|((m[566]&~m[873]&~m[875]&m[876]&~m[877])|(~m[566]&~m[873]&~m[875]&~m[876]&m[877])|(m[566]&~m[873]&~m[875]&~m[876]&m[877])|(m[566]&m[873]&~m[875]&~m[876]&m[877])|(m[566]&~m[873]&m[875]&~m[876]&m[877])|(~m[566]&~m[873]&~m[875]&m[876]&m[877])|(m[566]&~m[873]&~m[875]&m[876]&m[877])|(~m[566]&m[873]&~m[875]&m[876]&m[877])|(m[566]&m[873]&~m[875]&m[876]&m[877])|(~m[566]&~m[873]&m[875]&m[876]&m[877])|(m[566]&~m[873]&m[875]&m[876]&m[877])|(m[566]&m[873]&m[875]&m[876]&m[877]));
    m[880] = (((m[847]&~m[878]&~m[879]&~m[881]&~m[882])|(~m[847]&~m[878]&~m[879]&m[881]&~m[882])|(m[847]&m[878]&~m[879]&m[881]&~m[882])|(m[847]&~m[878]&m[879]&m[881]&~m[882])|(~m[847]&m[878]&~m[879]&~m[881]&m[882])|(~m[847]&~m[878]&m[879]&~m[881]&m[882])|(m[847]&m[878]&m[879]&~m[881]&m[882])|(~m[847]&m[878]&m[879]&m[881]&m[882]))&UnbiasedRNG[234])|((m[847]&~m[878]&~m[879]&m[881]&~m[882])|(~m[847]&~m[878]&~m[879]&~m[881]&m[882])|(m[847]&~m[878]&~m[879]&~m[881]&m[882])|(m[847]&m[878]&~m[879]&~m[881]&m[882])|(m[847]&~m[878]&m[879]&~m[881]&m[882])|(~m[847]&~m[878]&~m[879]&m[881]&m[882])|(m[847]&~m[878]&~m[879]&m[881]&m[882])|(~m[847]&m[878]&~m[879]&m[881]&m[882])|(m[847]&m[878]&~m[879]&m[881]&m[882])|(~m[847]&~m[878]&m[879]&m[881]&m[882])|(m[847]&~m[878]&m[879]&m[881]&m[882])|(m[847]&m[878]&m[879]&m[881]&m[882]));
    m[885] = (((m[852]&~m[883]&~m[884]&~m[886]&~m[887])|(~m[852]&~m[883]&~m[884]&m[886]&~m[887])|(m[852]&m[883]&~m[884]&m[886]&~m[887])|(m[852]&~m[883]&m[884]&m[886]&~m[887])|(~m[852]&m[883]&~m[884]&~m[886]&m[887])|(~m[852]&~m[883]&m[884]&~m[886]&m[887])|(m[852]&m[883]&m[884]&~m[886]&m[887])|(~m[852]&m[883]&m[884]&m[886]&m[887]))&UnbiasedRNG[235])|((m[852]&~m[883]&~m[884]&m[886]&~m[887])|(~m[852]&~m[883]&~m[884]&~m[886]&m[887])|(m[852]&~m[883]&~m[884]&~m[886]&m[887])|(m[852]&m[883]&~m[884]&~m[886]&m[887])|(m[852]&~m[883]&m[884]&~m[886]&m[887])|(~m[852]&~m[883]&~m[884]&m[886]&m[887])|(m[852]&~m[883]&~m[884]&m[886]&m[887])|(~m[852]&m[883]&~m[884]&m[886]&m[887])|(m[852]&m[883]&~m[884]&m[886]&m[887])|(~m[852]&~m[883]&m[884]&m[886]&m[887])|(m[852]&~m[883]&m[884]&m[886]&m[887])|(m[852]&m[883]&m[884]&m[886]&m[887]));
    m[890] = (((m[857]&~m[888]&~m[889]&~m[891]&~m[892])|(~m[857]&~m[888]&~m[889]&m[891]&~m[892])|(m[857]&m[888]&~m[889]&m[891]&~m[892])|(m[857]&~m[888]&m[889]&m[891]&~m[892])|(~m[857]&m[888]&~m[889]&~m[891]&m[892])|(~m[857]&~m[888]&m[889]&~m[891]&m[892])|(m[857]&m[888]&m[889]&~m[891]&m[892])|(~m[857]&m[888]&m[889]&m[891]&m[892]))&UnbiasedRNG[236])|((m[857]&~m[888]&~m[889]&m[891]&~m[892])|(~m[857]&~m[888]&~m[889]&~m[891]&m[892])|(m[857]&~m[888]&~m[889]&~m[891]&m[892])|(m[857]&m[888]&~m[889]&~m[891]&m[892])|(m[857]&~m[888]&m[889]&~m[891]&m[892])|(~m[857]&~m[888]&~m[889]&m[891]&m[892])|(m[857]&~m[888]&~m[889]&m[891]&m[892])|(~m[857]&m[888]&~m[889]&m[891]&m[892])|(m[857]&m[888]&~m[889]&m[891]&m[892])|(~m[857]&~m[888]&m[889]&m[891]&m[892])|(m[857]&~m[888]&m[889]&m[891]&m[892])|(m[857]&m[888]&m[889]&m[891]&m[892]));
    m[894] = (((m[618]&~m[893]&~m[895]&~m[896]&~m[897])|(~m[618]&~m[893]&~m[895]&m[896]&~m[897])|(m[618]&m[893]&~m[895]&m[896]&~m[897])|(m[618]&~m[893]&m[895]&m[896]&~m[897])|(~m[618]&m[893]&~m[895]&~m[896]&m[897])|(~m[618]&~m[893]&m[895]&~m[896]&m[897])|(m[618]&m[893]&m[895]&~m[896]&m[897])|(~m[618]&m[893]&m[895]&m[896]&m[897]))&UnbiasedRNG[237])|((m[618]&~m[893]&~m[895]&m[896]&~m[897])|(~m[618]&~m[893]&~m[895]&~m[896]&m[897])|(m[618]&~m[893]&~m[895]&~m[896]&m[897])|(m[618]&m[893]&~m[895]&~m[896]&m[897])|(m[618]&~m[893]&m[895]&~m[896]&m[897])|(~m[618]&~m[893]&~m[895]&m[896]&m[897])|(m[618]&~m[893]&~m[895]&m[896]&m[897])|(~m[618]&m[893]&~m[895]&m[896]&m[897])|(m[618]&m[893]&~m[895]&m[896]&m[897])|(~m[618]&~m[893]&m[895]&m[896]&m[897])|(m[618]&~m[893]&m[895]&m[896]&m[897])|(m[618]&m[893]&m[895]&m[896]&m[897]));
    m[899] = (((m[631]&~m[898]&~m[900]&~m[901]&~m[902])|(~m[631]&~m[898]&~m[900]&m[901]&~m[902])|(m[631]&m[898]&~m[900]&m[901]&~m[902])|(m[631]&~m[898]&m[900]&m[901]&~m[902])|(~m[631]&m[898]&~m[900]&~m[901]&m[902])|(~m[631]&~m[898]&m[900]&~m[901]&m[902])|(m[631]&m[898]&m[900]&~m[901]&m[902])|(~m[631]&m[898]&m[900]&m[901]&m[902]))&UnbiasedRNG[238])|((m[631]&~m[898]&~m[900]&m[901]&~m[902])|(~m[631]&~m[898]&~m[900]&~m[901]&m[902])|(m[631]&~m[898]&~m[900]&~m[901]&m[902])|(m[631]&m[898]&~m[900]&~m[901]&m[902])|(m[631]&~m[898]&m[900]&~m[901]&m[902])|(~m[631]&~m[898]&~m[900]&m[901]&m[902])|(m[631]&~m[898]&~m[900]&m[901]&m[902])|(~m[631]&m[898]&~m[900]&m[901]&m[902])|(m[631]&m[898]&~m[900]&m[901]&m[902])|(~m[631]&~m[898]&m[900]&m[901]&m[902])|(m[631]&~m[898]&m[900]&m[901]&m[902])|(m[631]&m[898]&m[900]&m[901]&m[902]));
    m[904] = (((m[644]&~m[903]&~m[905]&~m[906]&~m[907])|(~m[644]&~m[903]&~m[905]&m[906]&~m[907])|(m[644]&m[903]&~m[905]&m[906]&~m[907])|(m[644]&~m[903]&m[905]&m[906]&~m[907])|(~m[644]&m[903]&~m[905]&~m[906]&m[907])|(~m[644]&~m[903]&m[905]&~m[906]&m[907])|(m[644]&m[903]&m[905]&~m[906]&m[907])|(~m[644]&m[903]&m[905]&m[906]&m[907]))&UnbiasedRNG[239])|((m[644]&~m[903]&~m[905]&m[906]&~m[907])|(~m[644]&~m[903]&~m[905]&~m[906]&m[907])|(m[644]&~m[903]&~m[905]&~m[906]&m[907])|(m[644]&m[903]&~m[905]&~m[906]&m[907])|(m[644]&~m[903]&m[905]&~m[906]&m[907])|(~m[644]&~m[903]&~m[905]&m[906]&m[907])|(m[644]&~m[903]&~m[905]&m[906]&m[907])|(~m[644]&m[903]&~m[905]&m[906]&m[907])|(m[644]&m[903]&~m[905]&m[906]&m[907])|(~m[644]&~m[903]&m[905]&m[906]&m[907])|(m[644]&~m[903]&m[905]&m[906]&m[907])|(m[644]&m[903]&m[905]&m[906]&m[907]));
    m[909] = (((m[554]&~m[908]&~m[910]&~m[911]&~m[912])|(~m[554]&~m[908]&~m[910]&m[911]&~m[912])|(m[554]&m[908]&~m[910]&m[911]&~m[912])|(m[554]&~m[908]&m[910]&m[911]&~m[912])|(~m[554]&m[908]&~m[910]&~m[911]&m[912])|(~m[554]&~m[908]&m[910]&~m[911]&m[912])|(m[554]&m[908]&m[910]&~m[911]&m[912])|(~m[554]&m[908]&m[910]&m[911]&m[912]))&UnbiasedRNG[240])|((m[554]&~m[908]&~m[910]&m[911]&~m[912])|(~m[554]&~m[908]&~m[910]&~m[911]&m[912])|(m[554]&~m[908]&~m[910]&~m[911]&m[912])|(m[554]&m[908]&~m[910]&~m[911]&m[912])|(m[554]&~m[908]&m[910]&~m[911]&m[912])|(~m[554]&~m[908]&~m[910]&m[911]&m[912])|(m[554]&~m[908]&~m[910]&m[911]&m[912])|(~m[554]&m[908]&~m[910]&m[911]&m[912])|(m[554]&m[908]&~m[910]&m[911]&m[912])|(~m[554]&~m[908]&m[910]&m[911]&m[912])|(m[554]&~m[908]&m[910]&m[911]&m[912])|(m[554]&m[908]&m[910]&m[911]&m[912]));
    m[914] = (((m[567]&~m[913]&~m[915]&~m[916]&~m[917])|(~m[567]&~m[913]&~m[915]&m[916]&~m[917])|(m[567]&m[913]&~m[915]&m[916]&~m[917])|(m[567]&~m[913]&m[915]&m[916]&~m[917])|(~m[567]&m[913]&~m[915]&~m[916]&m[917])|(~m[567]&~m[913]&m[915]&~m[916]&m[917])|(m[567]&m[913]&m[915]&~m[916]&m[917])|(~m[567]&m[913]&m[915]&m[916]&m[917]))&UnbiasedRNG[241])|((m[567]&~m[913]&~m[915]&m[916]&~m[917])|(~m[567]&~m[913]&~m[915]&~m[916]&m[917])|(m[567]&~m[913]&~m[915]&~m[916]&m[917])|(m[567]&m[913]&~m[915]&~m[916]&m[917])|(m[567]&~m[913]&m[915]&~m[916]&m[917])|(~m[567]&~m[913]&~m[915]&m[916]&m[917])|(m[567]&~m[913]&~m[915]&m[916]&m[917])|(~m[567]&m[913]&~m[915]&m[916]&m[917])|(m[567]&m[913]&~m[915]&m[916]&m[917])|(~m[567]&~m[913]&m[915]&m[916]&m[917])|(m[567]&~m[913]&m[915]&m[916]&m[917])|(m[567]&m[913]&m[915]&m[916]&m[917]));
    m[919] = (((m[580]&~m[918]&~m[920]&~m[921]&~m[922])|(~m[580]&~m[918]&~m[920]&m[921]&~m[922])|(m[580]&m[918]&~m[920]&m[921]&~m[922])|(m[580]&~m[918]&m[920]&m[921]&~m[922])|(~m[580]&m[918]&~m[920]&~m[921]&m[922])|(~m[580]&~m[918]&m[920]&~m[921]&m[922])|(m[580]&m[918]&m[920]&~m[921]&m[922])|(~m[580]&m[918]&m[920]&m[921]&m[922]))&UnbiasedRNG[242])|((m[580]&~m[918]&~m[920]&m[921]&~m[922])|(~m[580]&~m[918]&~m[920]&~m[921]&m[922])|(m[580]&~m[918]&~m[920]&~m[921]&m[922])|(m[580]&m[918]&~m[920]&~m[921]&m[922])|(m[580]&~m[918]&m[920]&~m[921]&m[922])|(~m[580]&~m[918]&~m[920]&m[921]&m[922])|(m[580]&~m[918]&~m[920]&m[921]&m[922])|(~m[580]&m[918]&~m[920]&m[921]&m[922])|(m[580]&m[918]&~m[920]&m[921]&m[922])|(~m[580]&~m[918]&m[920]&m[921]&m[922])|(m[580]&~m[918]&m[920]&m[921]&m[922])|(m[580]&m[918]&m[920]&m[921]&m[922]));
    m[925] = (((m[887]&~m[923]&~m[924]&~m[926]&~m[927])|(~m[887]&~m[923]&~m[924]&m[926]&~m[927])|(m[887]&m[923]&~m[924]&m[926]&~m[927])|(m[887]&~m[923]&m[924]&m[926]&~m[927])|(~m[887]&m[923]&~m[924]&~m[926]&m[927])|(~m[887]&~m[923]&m[924]&~m[926]&m[927])|(m[887]&m[923]&m[924]&~m[926]&m[927])|(~m[887]&m[923]&m[924]&m[926]&m[927]))&UnbiasedRNG[243])|((m[887]&~m[923]&~m[924]&m[926]&~m[927])|(~m[887]&~m[923]&~m[924]&~m[926]&m[927])|(m[887]&~m[923]&~m[924]&~m[926]&m[927])|(m[887]&m[923]&~m[924]&~m[926]&m[927])|(m[887]&~m[923]&m[924]&~m[926]&m[927])|(~m[887]&~m[923]&~m[924]&m[926]&m[927])|(m[887]&~m[923]&~m[924]&m[926]&m[927])|(~m[887]&m[923]&~m[924]&m[926]&m[927])|(m[887]&m[923]&~m[924]&m[926]&m[927])|(~m[887]&~m[923]&m[924]&m[926]&m[927])|(m[887]&~m[923]&m[924]&m[926]&m[927])|(m[887]&m[923]&m[924]&m[926]&m[927]));
    m[930] = (((m[892]&~m[928]&~m[929]&~m[931]&~m[932])|(~m[892]&~m[928]&~m[929]&m[931]&~m[932])|(m[892]&m[928]&~m[929]&m[931]&~m[932])|(m[892]&~m[928]&m[929]&m[931]&~m[932])|(~m[892]&m[928]&~m[929]&~m[931]&m[932])|(~m[892]&~m[928]&m[929]&~m[931]&m[932])|(m[892]&m[928]&m[929]&~m[931]&m[932])|(~m[892]&m[928]&m[929]&m[931]&m[932]))&UnbiasedRNG[244])|((m[892]&~m[928]&~m[929]&m[931]&~m[932])|(~m[892]&~m[928]&~m[929]&~m[931]&m[932])|(m[892]&~m[928]&~m[929]&~m[931]&m[932])|(m[892]&m[928]&~m[929]&~m[931]&m[932])|(m[892]&~m[928]&m[929]&~m[931]&m[932])|(~m[892]&~m[928]&~m[929]&m[931]&m[932])|(m[892]&~m[928]&~m[929]&m[931]&m[932])|(~m[892]&m[928]&~m[929]&m[931]&m[932])|(m[892]&m[928]&~m[929]&m[931]&m[932])|(~m[892]&~m[928]&m[929]&m[931]&m[932])|(m[892]&~m[928]&m[929]&m[931]&m[932])|(m[892]&m[928]&m[929]&m[931]&m[932]));
    m[934] = (((m[619]&~m[933]&~m[935]&~m[936]&~m[937])|(~m[619]&~m[933]&~m[935]&m[936]&~m[937])|(m[619]&m[933]&~m[935]&m[936]&~m[937])|(m[619]&~m[933]&m[935]&m[936]&~m[937])|(~m[619]&m[933]&~m[935]&~m[936]&m[937])|(~m[619]&~m[933]&m[935]&~m[936]&m[937])|(m[619]&m[933]&m[935]&~m[936]&m[937])|(~m[619]&m[933]&m[935]&m[936]&m[937]))&UnbiasedRNG[245])|((m[619]&~m[933]&~m[935]&m[936]&~m[937])|(~m[619]&~m[933]&~m[935]&~m[936]&m[937])|(m[619]&~m[933]&~m[935]&~m[936]&m[937])|(m[619]&m[933]&~m[935]&~m[936]&m[937])|(m[619]&~m[933]&m[935]&~m[936]&m[937])|(~m[619]&~m[933]&~m[935]&m[936]&m[937])|(m[619]&~m[933]&~m[935]&m[936]&m[937])|(~m[619]&m[933]&~m[935]&m[936]&m[937])|(m[619]&m[933]&~m[935]&m[936]&m[937])|(~m[619]&~m[933]&m[935]&m[936]&m[937])|(m[619]&~m[933]&m[935]&m[936]&m[937])|(m[619]&m[933]&m[935]&m[936]&m[937]));
    m[939] = (((m[632]&~m[938]&~m[940]&~m[941]&~m[942])|(~m[632]&~m[938]&~m[940]&m[941]&~m[942])|(m[632]&m[938]&~m[940]&m[941]&~m[942])|(m[632]&~m[938]&m[940]&m[941]&~m[942])|(~m[632]&m[938]&~m[940]&~m[941]&m[942])|(~m[632]&~m[938]&m[940]&~m[941]&m[942])|(m[632]&m[938]&m[940]&~m[941]&m[942])|(~m[632]&m[938]&m[940]&m[941]&m[942]))&UnbiasedRNG[246])|((m[632]&~m[938]&~m[940]&m[941]&~m[942])|(~m[632]&~m[938]&~m[940]&~m[941]&m[942])|(m[632]&~m[938]&~m[940]&~m[941]&m[942])|(m[632]&m[938]&~m[940]&~m[941]&m[942])|(m[632]&~m[938]&m[940]&~m[941]&m[942])|(~m[632]&~m[938]&~m[940]&m[941]&m[942])|(m[632]&~m[938]&~m[940]&m[941]&m[942])|(~m[632]&m[938]&~m[940]&m[941]&m[942])|(m[632]&m[938]&~m[940]&m[941]&m[942])|(~m[632]&~m[938]&m[940]&m[941]&m[942])|(m[632]&~m[938]&m[940]&m[941]&m[942])|(m[632]&m[938]&m[940]&m[941]&m[942]));
    m[944] = (((m[645]&~m[943]&~m[945]&~m[946]&~m[947])|(~m[645]&~m[943]&~m[945]&m[946]&~m[947])|(m[645]&m[943]&~m[945]&m[946]&~m[947])|(m[645]&~m[943]&m[945]&m[946]&~m[947])|(~m[645]&m[943]&~m[945]&~m[946]&m[947])|(~m[645]&~m[943]&m[945]&~m[946]&m[947])|(m[645]&m[943]&m[945]&~m[946]&m[947])|(~m[645]&m[943]&m[945]&m[946]&m[947]))&UnbiasedRNG[247])|((m[645]&~m[943]&~m[945]&m[946]&~m[947])|(~m[645]&~m[943]&~m[945]&~m[946]&m[947])|(m[645]&~m[943]&~m[945]&~m[946]&m[947])|(m[645]&m[943]&~m[945]&~m[946]&m[947])|(m[645]&~m[943]&m[945]&~m[946]&m[947])|(~m[645]&~m[943]&~m[945]&m[946]&m[947])|(m[645]&~m[943]&~m[945]&m[946]&m[947])|(~m[645]&m[943]&~m[945]&m[946]&m[947])|(m[645]&m[943]&~m[945]&m[946]&m[947])|(~m[645]&~m[943]&m[945]&m[946]&m[947])|(m[645]&~m[943]&m[945]&m[946]&m[947])|(m[645]&m[943]&m[945]&m[946]&m[947]));
    m[949] = (((m[658]&~m[948]&~m[950]&~m[951]&~m[952])|(~m[658]&~m[948]&~m[950]&m[951]&~m[952])|(m[658]&m[948]&~m[950]&m[951]&~m[952])|(m[658]&~m[948]&m[950]&m[951]&~m[952])|(~m[658]&m[948]&~m[950]&~m[951]&m[952])|(~m[658]&~m[948]&m[950]&~m[951]&m[952])|(m[658]&m[948]&m[950]&~m[951]&m[952])|(~m[658]&m[948]&m[950]&m[951]&m[952]))&UnbiasedRNG[248])|((m[658]&~m[948]&~m[950]&m[951]&~m[952])|(~m[658]&~m[948]&~m[950]&~m[951]&m[952])|(m[658]&~m[948]&~m[950]&~m[951]&m[952])|(m[658]&m[948]&~m[950]&~m[951]&m[952])|(m[658]&~m[948]&m[950]&~m[951]&m[952])|(~m[658]&~m[948]&~m[950]&m[951]&m[952])|(m[658]&~m[948]&~m[950]&m[951]&m[952])|(~m[658]&m[948]&~m[950]&m[951]&m[952])|(m[658]&m[948]&~m[950]&m[951]&m[952])|(~m[658]&~m[948]&m[950]&m[951]&m[952])|(m[658]&~m[948]&m[950]&m[951]&m[952])|(m[658]&m[948]&m[950]&m[951]&m[952]));
    m[954] = (((m[555]&~m[953]&~m[955]&~m[956]&~m[957])|(~m[555]&~m[953]&~m[955]&m[956]&~m[957])|(m[555]&m[953]&~m[955]&m[956]&~m[957])|(m[555]&~m[953]&m[955]&m[956]&~m[957])|(~m[555]&m[953]&~m[955]&~m[956]&m[957])|(~m[555]&~m[953]&m[955]&~m[956]&m[957])|(m[555]&m[953]&m[955]&~m[956]&m[957])|(~m[555]&m[953]&m[955]&m[956]&m[957]))&UnbiasedRNG[249])|((m[555]&~m[953]&~m[955]&m[956]&~m[957])|(~m[555]&~m[953]&~m[955]&~m[956]&m[957])|(m[555]&~m[953]&~m[955]&~m[956]&m[957])|(m[555]&m[953]&~m[955]&~m[956]&m[957])|(m[555]&~m[953]&m[955]&~m[956]&m[957])|(~m[555]&~m[953]&~m[955]&m[956]&m[957])|(m[555]&~m[953]&~m[955]&m[956]&m[957])|(~m[555]&m[953]&~m[955]&m[956]&m[957])|(m[555]&m[953]&~m[955]&m[956]&m[957])|(~m[555]&~m[953]&m[955]&m[956]&m[957])|(m[555]&~m[953]&m[955]&m[956]&m[957])|(m[555]&m[953]&m[955]&m[956]&m[957]));
    m[959] = (((m[568]&~m[958]&~m[960]&~m[961]&~m[962])|(~m[568]&~m[958]&~m[960]&m[961]&~m[962])|(m[568]&m[958]&~m[960]&m[961]&~m[962])|(m[568]&~m[958]&m[960]&m[961]&~m[962])|(~m[568]&m[958]&~m[960]&~m[961]&m[962])|(~m[568]&~m[958]&m[960]&~m[961]&m[962])|(m[568]&m[958]&m[960]&~m[961]&m[962])|(~m[568]&m[958]&m[960]&m[961]&m[962]))&UnbiasedRNG[250])|((m[568]&~m[958]&~m[960]&m[961]&~m[962])|(~m[568]&~m[958]&~m[960]&~m[961]&m[962])|(m[568]&~m[958]&~m[960]&~m[961]&m[962])|(m[568]&m[958]&~m[960]&~m[961]&m[962])|(m[568]&~m[958]&m[960]&~m[961]&m[962])|(~m[568]&~m[958]&~m[960]&m[961]&m[962])|(m[568]&~m[958]&~m[960]&m[961]&m[962])|(~m[568]&m[958]&~m[960]&m[961]&m[962])|(m[568]&m[958]&~m[960]&m[961]&m[962])|(~m[568]&~m[958]&m[960]&m[961]&m[962])|(m[568]&~m[958]&m[960]&m[961]&m[962])|(m[568]&m[958]&m[960]&m[961]&m[962]));
    m[964] = (((m[581]&~m[963]&~m[965]&~m[966]&~m[967])|(~m[581]&~m[963]&~m[965]&m[966]&~m[967])|(m[581]&m[963]&~m[965]&m[966]&~m[967])|(m[581]&~m[963]&m[965]&m[966]&~m[967])|(~m[581]&m[963]&~m[965]&~m[966]&m[967])|(~m[581]&~m[963]&m[965]&~m[966]&m[967])|(m[581]&m[963]&m[965]&~m[966]&m[967])|(~m[581]&m[963]&m[965]&m[966]&m[967]))&UnbiasedRNG[251])|((m[581]&~m[963]&~m[965]&m[966]&~m[967])|(~m[581]&~m[963]&~m[965]&~m[966]&m[967])|(m[581]&~m[963]&~m[965]&~m[966]&m[967])|(m[581]&m[963]&~m[965]&~m[966]&m[967])|(m[581]&~m[963]&m[965]&~m[966]&m[967])|(~m[581]&~m[963]&~m[965]&m[966]&m[967])|(m[581]&~m[963]&~m[965]&m[966]&m[967])|(~m[581]&m[963]&~m[965]&m[966]&m[967])|(m[581]&m[963]&~m[965]&m[966]&m[967])|(~m[581]&~m[963]&m[965]&m[966]&m[967])|(m[581]&~m[963]&m[965]&m[966]&m[967])|(m[581]&m[963]&m[965]&m[966]&m[967]));
    m[969] = (((m[594]&~m[968]&~m[970]&~m[971]&~m[972])|(~m[594]&~m[968]&~m[970]&m[971]&~m[972])|(m[594]&m[968]&~m[970]&m[971]&~m[972])|(m[594]&~m[968]&m[970]&m[971]&~m[972])|(~m[594]&m[968]&~m[970]&~m[971]&m[972])|(~m[594]&~m[968]&m[970]&~m[971]&m[972])|(m[594]&m[968]&m[970]&~m[971]&m[972])|(~m[594]&m[968]&m[970]&m[971]&m[972]))&UnbiasedRNG[252])|((m[594]&~m[968]&~m[970]&m[971]&~m[972])|(~m[594]&~m[968]&~m[970]&~m[971]&m[972])|(m[594]&~m[968]&~m[970]&~m[971]&m[972])|(m[594]&m[968]&~m[970]&~m[971]&m[972])|(m[594]&~m[968]&m[970]&~m[971]&m[972])|(~m[594]&~m[968]&~m[970]&m[971]&m[972])|(m[594]&~m[968]&~m[970]&m[971]&m[972])|(~m[594]&m[968]&~m[970]&m[971]&m[972])|(m[594]&m[968]&~m[970]&m[971]&m[972])|(~m[594]&~m[968]&m[970]&m[971]&m[972])|(m[594]&~m[968]&m[970]&m[971]&m[972])|(m[594]&m[968]&m[970]&m[971]&m[972]));
    m[975] = (((m[932]&~m[973]&~m[974]&~m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&m[976]&~m[977])|(m[932]&m[973]&~m[974]&m[976]&~m[977])|(m[932]&~m[973]&m[974]&m[976]&~m[977])|(~m[932]&m[973]&~m[974]&~m[976]&m[977])|(~m[932]&~m[973]&m[974]&~m[976]&m[977])|(m[932]&m[973]&m[974]&~m[976]&m[977])|(~m[932]&m[973]&m[974]&m[976]&m[977]))&UnbiasedRNG[253])|((m[932]&~m[973]&~m[974]&m[976]&~m[977])|(~m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&~m[974]&~m[976]&m[977])|(m[932]&m[973]&~m[974]&~m[976]&m[977])|(m[932]&~m[973]&m[974]&~m[976]&m[977])|(~m[932]&~m[973]&~m[974]&m[976]&m[977])|(m[932]&~m[973]&~m[974]&m[976]&m[977])|(~m[932]&m[973]&~m[974]&m[976]&m[977])|(m[932]&m[973]&~m[974]&m[976]&m[977])|(~m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&~m[973]&m[974]&m[976]&m[977])|(m[932]&m[973]&m[974]&m[976]&m[977]));
    m[979] = (((m[620]&~m[978]&~m[980]&~m[981]&~m[982])|(~m[620]&~m[978]&~m[980]&m[981]&~m[982])|(m[620]&m[978]&~m[980]&m[981]&~m[982])|(m[620]&~m[978]&m[980]&m[981]&~m[982])|(~m[620]&m[978]&~m[980]&~m[981]&m[982])|(~m[620]&~m[978]&m[980]&~m[981]&m[982])|(m[620]&m[978]&m[980]&~m[981]&m[982])|(~m[620]&m[978]&m[980]&m[981]&m[982]))&UnbiasedRNG[254])|((m[620]&~m[978]&~m[980]&m[981]&~m[982])|(~m[620]&~m[978]&~m[980]&~m[981]&m[982])|(m[620]&~m[978]&~m[980]&~m[981]&m[982])|(m[620]&m[978]&~m[980]&~m[981]&m[982])|(m[620]&~m[978]&m[980]&~m[981]&m[982])|(~m[620]&~m[978]&~m[980]&m[981]&m[982])|(m[620]&~m[978]&~m[980]&m[981]&m[982])|(~m[620]&m[978]&~m[980]&m[981]&m[982])|(m[620]&m[978]&~m[980]&m[981]&m[982])|(~m[620]&~m[978]&m[980]&m[981]&m[982])|(m[620]&~m[978]&m[980]&m[981]&m[982])|(m[620]&m[978]&m[980]&m[981]&m[982]));
    m[984] = (((m[633]&~m[983]&~m[985]&~m[986]&~m[987])|(~m[633]&~m[983]&~m[985]&m[986]&~m[987])|(m[633]&m[983]&~m[985]&m[986]&~m[987])|(m[633]&~m[983]&m[985]&m[986]&~m[987])|(~m[633]&m[983]&~m[985]&~m[986]&m[987])|(~m[633]&~m[983]&m[985]&~m[986]&m[987])|(m[633]&m[983]&m[985]&~m[986]&m[987])|(~m[633]&m[983]&m[985]&m[986]&m[987]))&UnbiasedRNG[255])|((m[633]&~m[983]&~m[985]&m[986]&~m[987])|(~m[633]&~m[983]&~m[985]&~m[986]&m[987])|(m[633]&~m[983]&~m[985]&~m[986]&m[987])|(m[633]&m[983]&~m[985]&~m[986]&m[987])|(m[633]&~m[983]&m[985]&~m[986]&m[987])|(~m[633]&~m[983]&~m[985]&m[986]&m[987])|(m[633]&~m[983]&~m[985]&m[986]&m[987])|(~m[633]&m[983]&~m[985]&m[986]&m[987])|(m[633]&m[983]&~m[985]&m[986]&m[987])|(~m[633]&~m[983]&m[985]&m[986]&m[987])|(m[633]&~m[983]&m[985]&m[986]&m[987])|(m[633]&m[983]&m[985]&m[986]&m[987]));
    m[989] = (((m[646]&~m[988]&~m[990]&~m[991]&~m[992])|(~m[646]&~m[988]&~m[990]&m[991]&~m[992])|(m[646]&m[988]&~m[990]&m[991]&~m[992])|(m[646]&~m[988]&m[990]&m[991]&~m[992])|(~m[646]&m[988]&~m[990]&~m[991]&m[992])|(~m[646]&~m[988]&m[990]&~m[991]&m[992])|(m[646]&m[988]&m[990]&~m[991]&m[992])|(~m[646]&m[988]&m[990]&m[991]&m[992]))&UnbiasedRNG[256])|((m[646]&~m[988]&~m[990]&m[991]&~m[992])|(~m[646]&~m[988]&~m[990]&~m[991]&m[992])|(m[646]&~m[988]&~m[990]&~m[991]&m[992])|(m[646]&m[988]&~m[990]&~m[991]&m[992])|(m[646]&~m[988]&m[990]&~m[991]&m[992])|(~m[646]&~m[988]&~m[990]&m[991]&m[992])|(m[646]&~m[988]&~m[990]&m[991]&m[992])|(~m[646]&m[988]&~m[990]&m[991]&m[992])|(m[646]&m[988]&~m[990]&m[991]&m[992])|(~m[646]&~m[988]&m[990]&m[991]&m[992])|(m[646]&~m[988]&m[990]&m[991]&m[992])|(m[646]&m[988]&m[990]&m[991]&m[992]));
    m[994] = (((m[659]&~m[993]&~m[995]&~m[996]&~m[997])|(~m[659]&~m[993]&~m[995]&m[996]&~m[997])|(m[659]&m[993]&~m[995]&m[996]&~m[997])|(m[659]&~m[993]&m[995]&m[996]&~m[997])|(~m[659]&m[993]&~m[995]&~m[996]&m[997])|(~m[659]&~m[993]&m[995]&~m[996]&m[997])|(m[659]&m[993]&m[995]&~m[996]&m[997])|(~m[659]&m[993]&m[995]&m[996]&m[997]))&UnbiasedRNG[257])|((m[659]&~m[993]&~m[995]&m[996]&~m[997])|(~m[659]&~m[993]&~m[995]&~m[996]&m[997])|(m[659]&~m[993]&~m[995]&~m[996]&m[997])|(m[659]&m[993]&~m[995]&~m[996]&m[997])|(m[659]&~m[993]&m[995]&~m[996]&m[997])|(~m[659]&~m[993]&~m[995]&m[996]&m[997])|(m[659]&~m[993]&~m[995]&m[996]&m[997])|(~m[659]&m[993]&~m[995]&m[996]&m[997])|(m[659]&m[993]&~m[995]&m[996]&m[997])|(~m[659]&~m[993]&m[995]&m[996]&m[997])|(m[659]&~m[993]&m[995]&m[996]&m[997])|(m[659]&m[993]&m[995]&m[996]&m[997]));
    m[999] = (((m[672]&~m[998]&~m[1000]&~m[1001]&~m[1002])|(~m[672]&~m[998]&~m[1000]&m[1001]&~m[1002])|(m[672]&m[998]&~m[1000]&m[1001]&~m[1002])|(m[672]&~m[998]&m[1000]&m[1001]&~m[1002])|(~m[672]&m[998]&~m[1000]&~m[1001]&m[1002])|(~m[672]&~m[998]&m[1000]&~m[1001]&m[1002])|(m[672]&m[998]&m[1000]&~m[1001]&m[1002])|(~m[672]&m[998]&m[1000]&m[1001]&m[1002]))&UnbiasedRNG[258])|((m[672]&~m[998]&~m[1000]&m[1001]&~m[1002])|(~m[672]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[672]&~m[998]&~m[1000]&~m[1001]&m[1002])|(m[672]&m[998]&~m[1000]&~m[1001]&m[1002])|(m[672]&~m[998]&m[1000]&~m[1001]&m[1002])|(~m[672]&~m[998]&~m[1000]&m[1001]&m[1002])|(m[672]&~m[998]&~m[1000]&m[1001]&m[1002])|(~m[672]&m[998]&~m[1000]&m[1001]&m[1002])|(m[672]&m[998]&~m[1000]&m[1001]&m[1002])|(~m[672]&~m[998]&m[1000]&m[1001]&m[1002])|(m[672]&~m[998]&m[1000]&m[1001]&m[1002])|(m[672]&m[998]&m[1000]&m[1001]&m[1002]));
    m[1004] = (((m[556]&~m[1003]&~m[1005]&~m[1006]&~m[1007])|(~m[556]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(m[556]&m[1003]&~m[1005]&m[1006]&~m[1007])|(m[556]&~m[1003]&m[1005]&m[1006]&~m[1007])|(~m[556]&m[1003]&~m[1005]&~m[1006]&m[1007])|(~m[556]&~m[1003]&m[1005]&~m[1006]&m[1007])|(m[556]&m[1003]&m[1005]&~m[1006]&m[1007])|(~m[556]&m[1003]&m[1005]&m[1006]&m[1007]))&UnbiasedRNG[259])|((m[556]&~m[1003]&~m[1005]&m[1006]&~m[1007])|(~m[556]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[556]&~m[1003]&~m[1005]&~m[1006]&m[1007])|(m[556]&m[1003]&~m[1005]&~m[1006]&m[1007])|(m[556]&~m[1003]&m[1005]&~m[1006]&m[1007])|(~m[556]&~m[1003]&~m[1005]&m[1006]&m[1007])|(m[556]&~m[1003]&~m[1005]&m[1006]&m[1007])|(~m[556]&m[1003]&~m[1005]&m[1006]&m[1007])|(m[556]&m[1003]&~m[1005]&m[1006]&m[1007])|(~m[556]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[556]&~m[1003]&m[1005]&m[1006]&m[1007])|(m[556]&m[1003]&m[1005]&m[1006]&m[1007]));
    m[1009] = (((m[569]&~m[1008]&~m[1010]&~m[1011]&~m[1012])|(~m[569]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(m[569]&m[1008]&~m[1010]&m[1011]&~m[1012])|(m[569]&~m[1008]&m[1010]&m[1011]&~m[1012])|(~m[569]&m[1008]&~m[1010]&~m[1011]&m[1012])|(~m[569]&~m[1008]&m[1010]&~m[1011]&m[1012])|(m[569]&m[1008]&m[1010]&~m[1011]&m[1012])|(~m[569]&m[1008]&m[1010]&m[1011]&m[1012]))&UnbiasedRNG[260])|((m[569]&~m[1008]&~m[1010]&m[1011]&~m[1012])|(~m[569]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[569]&~m[1008]&~m[1010]&~m[1011]&m[1012])|(m[569]&m[1008]&~m[1010]&~m[1011]&m[1012])|(m[569]&~m[1008]&m[1010]&~m[1011]&m[1012])|(~m[569]&~m[1008]&~m[1010]&m[1011]&m[1012])|(m[569]&~m[1008]&~m[1010]&m[1011]&m[1012])|(~m[569]&m[1008]&~m[1010]&m[1011]&m[1012])|(m[569]&m[1008]&~m[1010]&m[1011]&m[1012])|(~m[569]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[569]&~m[1008]&m[1010]&m[1011]&m[1012])|(m[569]&m[1008]&m[1010]&m[1011]&m[1012]));
    m[1014] = (((m[582]&~m[1013]&~m[1015]&~m[1016]&~m[1017])|(~m[582]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(m[582]&m[1013]&~m[1015]&m[1016]&~m[1017])|(m[582]&~m[1013]&m[1015]&m[1016]&~m[1017])|(~m[582]&m[1013]&~m[1015]&~m[1016]&m[1017])|(~m[582]&~m[1013]&m[1015]&~m[1016]&m[1017])|(m[582]&m[1013]&m[1015]&~m[1016]&m[1017])|(~m[582]&m[1013]&m[1015]&m[1016]&m[1017]))&UnbiasedRNG[261])|((m[582]&~m[1013]&~m[1015]&m[1016]&~m[1017])|(~m[582]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[582]&~m[1013]&~m[1015]&~m[1016]&m[1017])|(m[582]&m[1013]&~m[1015]&~m[1016]&m[1017])|(m[582]&~m[1013]&m[1015]&~m[1016]&m[1017])|(~m[582]&~m[1013]&~m[1015]&m[1016]&m[1017])|(m[582]&~m[1013]&~m[1015]&m[1016]&m[1017])|(~m[582]&m[1013]&~m[1015]&m[1016]&m[1017])|(m[582]&m[1013]&~m[1015]&m[1016]&m[1017])|(~m[582]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[582]&~m[1013]&m[1015]&m[1016]&m[1017])|(m[582]&m[1013]&m[1015]&m[1016]&m[1017]));
    m[1019] = (((m[595]&~m[1018]&~m[1020]&~m[1021]&~m[1022])|(~m[595]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(m[595]&m[1018]&~m[1020]&m[1021]&~m[1022])|(m[595]&~m[1018]&m[1020]&m[1021]&~m[1022])|(~m[595]&m[1018]&~m[1020]&~m[1021]&m[1022])|(~m[595]&~m[1018]&m[1020]&~m[1021]&m[1022])|(m[595]&m[1018]&m[1020]&~m[1021]&m[1022])|(~m[595]&m[1018]&m[1020]&m[1021]&m[1022]))&UnbiasedRNG[262])|((m[595]&~m[1018]&~m[1020]&m[1021]&~m[1022])|(~m[595]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[595]&~m[1018]&~m[1020]&~m[1021]&m[1022])|(m[595]&m[1018]&~m[1020]&~m[1021]&m[1022])|(m[595]&~m[1018]&m[1020]&~m[1021]&m[1022])|(~m[595]&~m[1018]&~m[1020]&m[1021]&m[1022])|(m[595]&~m[1018]&~m[1020]&m[1021]&m[1022])|(~m[595]&m[1018]&~m[1020]&m[1021]&m[1022])|(m[595]&m[1018]&~m[1020]&m[1021]&m[1022])|(~m[595]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[595]&~m[1018]&m[1020]&m[1021]&m[1022])|(m[595]&m[1018]&m[1020]&m[1021]&m[1022]));
    m[1024] = (((m[608]&~m[1023]&~m[1025]&~m[1026]&~m[1027])|(~m[608]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(m[608]&m[1023]&~m[1025]&m[1026]&~m[1027])|(m[608]&~m[1023]&m[1025]&m[1026]&~m[1027])|(~m[608]&m[1023]&~m[1025]&~m[1026]&m[1027])|(~m[608]&~m[1023]&m[1025]&~m[1026]&m[1027])|(m[608]&m[1023]&m[1025]&~m[1026]&m[1027])|(~m[608]&m[1023]&m[1025]&m[1026]&m[1027]))&UnbiasedRNG[263])|((m[608]&~m[1023]&~m[1025]&m[1026]&~m[1027])|(~m[608]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[608]&~m[1023]&~m[1025]&~m[1026]&m[1027])|(m[608]&m[1023]&~m[1025]&~m[1026]&m[1027])|(m[608]&~m[1023]&m[1025]&~m[1026]&m[1027])|(~m[608]&~m[1023]&~m[1025]&m[1026]&m[1027])|(m[608]&~m[1023]&~m[1025]&m[1026]&m[1027])|(~m[608]&m[1023]&~m[1025]&m[1026]&m[1027])|(m[608]&m[1023]&~m[1025]&m[1026]&m[1027])|(~m[608]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[608]&~m[1023]&m[1025]&m[1026]&m[1027])|(m[608]&m[1023]&m[1025]&m[1026]&m[1027]));
    m[1029] = (((m[621]&~m[1028]&~m[1030]&~m[1031]&~m[1032])|(~m[621]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(m[621]&m[1028]&~m[1030]&m[1031]&~m[1032])|(m[621]&~m[1028]&m[1030]&m[1031]&~m[1032])|(~m[621]&m[1028]&~m[1030]&~m[1031]&m[1032])|(~m[621]&~m[1028]&m[1030]&~m[1031]&m[1032])|(m[621]&m[1028]&m[1030]&~m[1031]&m[1032])|(~m[621]&m[1028]&m[1030]&m[1031]&m[1032]))&UnbiasedRNG[264])|((m[621]&~m[1028]&~m[1030]&m[1031]&~m[1032])|(~m[621]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[621]&~m[1028]&~m[1030]&~m[1031]&m[1032])|(m[621]&m[1028]&~m[1030]&~m[1031]&m[1032])|(m[621]&~m[1028]&m[1030]&~m[1031]&m[1032])|(~m[621]&~m[1028]&~m[1030]&m[1031]&m[1032])|(m[621]&~m[1028]&~m[1030]&m[1031]&m[1032])|(~m[621]&m[1028]&~m[1030]&m[1031]&m[1032])|(m[621]&m[1028]&~m[1030]&m[1031]&m[1032])|(~m[621]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[621]&~m[1028]&m[1030]&m[1031]&m[1032])|(m[621]&m[1028]&m[1030]&m[1031]&m[1032]));
    m[1034] = (((m[634]&~m[1033]&~m[1035]&~m[1036]&~m[1037])|(~m[634]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(m[634]&m[1033]&~m[1035]&m[1036]&~m[1037])|(m[634]&~m[1033]&m[1035]&m[1036]&~m[1037])|(~m[634]&m[1033]&~m[1035]&~m[1036]&m[1037])|(~m[634]&~m[1033]&m[1035]&~m[1036]&m[1037])|(m[634]&m[1033]&m[1035]&~m[1036]&m[1037])|(~m[634]&m[1033]&m[1035]&m[1036]&m[1037]))&UnbiasedRNG[265])|((m[634]&~m[1033]&~m[1035]&m[1036]&~m[1037])|(~m[634]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[634]&~m[1033]&~m[1035]&~m[1036]&m[1037])|(m[634]&m[1033]&~m[1035]&~m[1036]&m[1037])|(m[634]&~m[1033]&m[1035]&~m[1036]&m[1037])|(~m[634]&~m[1033]&~m[1035]&m[1036]&m[1037])|(m[634]&~m[1033]&~m[1035]&m[1036]&m[1037])|(~m[634]&m[1033]&~m[1035]&m[1036]&m[1037])|(m[634]&m[1033]&~m[1035]&m[1036]&m[1037])|(~m[634]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[634]&~m[1033]&m[1035]&m[1036]&m[1037])|(m[634]&m[1033]&m[1035]&m[1036]&m[1037]));
    m[1039] = (((m[647]&~m[1038]&~m[1040]&~m[1041]&~m[1042])|(~m[647]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(m[647]&m[1038]&~m[1040]&m[1041]&~m[1042])|(m[647]&~m[1038]&m[1040]&m[1041]&~m[1042])|(~m[647]&m[1038]&~m[1040]&~m[1041]&m[1042])|(~m[647]&~m[1038]&m[1040]&~m[1041]&m[1042])|(m[647]&m[1038]&m[1040]&~m[1041]&m[1042])|(~m[647]&m[1038]&m[1040]&m[1041]&m[1042]))&UnbiasedRNG[266])|((m[647]&~m[1038]&~m[1040]&m[1041]&~m[1042])|(~m[647]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[647]&~m[1038]&~m[1040]&~m[1041]&m[1042])|(m[647]&m[1038]&~m[1040]&~m[1041]&m[1042])|(m[647]&~m[1038]&m[1040]&~m[1041]&m[1042])|(~m[647]&~m[1038]&~m[1040]&m[1041]&m[1042])|(m[647]&~m[1038]&~m[1040]&m[1041]&m[1042])|(~m[647]&m[1038]&~m[1040]&m[1041]&m[1042])|(m[647]&m[1038]&~m[1040]&m[1041]&m[1042])|(~m[647]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[647]&~m[1038]&m[1040]&m[1041]&m[1042])|(m[647]&m[1038]&m[1040]&m[1041]&m[1042]));
    m[1044] = (((m[660]&~m[1043]&~m[1045]&~m[1046]&~m[1047])|(~m[660]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(m[660]&m[1043]&~m[1045]&m[1046]&~m[1047])|(m[660]&~m[1043]&m[1045]&m[1046]&~m[1047])|(~m[660]&m[1043]&~m[1045]&~m[1046]&m[1047])|(~m[660]&~m[1043]&m[1045]&~m[1046]&m[1047])|(m[660]&m[1043]&m[1045]&~m[1046]&m[1047])|(~m[660]&m[1043]&m[1045]&m[1046]&m[1047]))&UnbiasedRNG[267])|((m[660]&~m[1043]&~m[1045]&m[1046]&~m[1047])|(~m[660]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[660]&~m[1043]&~m[1045]&~m[1046]&m[1047])|(m[660]&m[1043]&~m[1045]&~m[1046]&m[1047])|(m[660]&~m[1043]&m[1045]&~m[1046]&m[1047])|(~m[660]&~m[1043]&~m[1045]&m[1046]&m[1047])|(m[660]&~m[1043]&~m[1045]&m[1046]&m[1047])|(~m[660]&m[1043]&~m[1045]&m[1046]&m[1047])|(m[660]&m[1043]&~m[1045]&m[1046]&m[1047])|(~m[660]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[660]&~m[1043]&m[1045]&m[1046]&m[1047])|(m[660]&m[1043]&m[1045]&m[1046]&m[1047]));
    m[1049] = (((m[673]&~m[1048]&~m[1050]&~m[1051]&~m[1052])|(~m[673]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(m[673]&m[1048]&~m[1050]&m[1051]&~m[1052])|(m[673]&~m[1048]&m[1050]&m[1051]&~m[1052])|(~m[673]&m[1048]&~m[1050]&~m[1051]&m[1052])|(~m[673]&~m[1048]&m[1050]&~m[1051]&m[1052])|(m[673]&m[1048]&m[1050]&~m[1051]&m[1052])|(~m[673]&m[1048]&m[1050]&m[1051]&m[1052]))&UnbiasedRNG[268])|((m[673]&~m[1048]&~m[1050]&m[1051]&~m[1052])|(~m[673]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[673]&~m[1048]&~m[1050]&~m[1051]&m[1052])|(m[673]&m[1048]&~m[1050]&~m[1051]&m[1052])|(m[673]&~m[1048]&m[1050]&~m[1051]&m[1052])|(~m[673]&~m[1048]&~m[1050]&m[1051]&m[1052])|(m[673]&~m[1048]&~m[1050]&m[1051]&m[1052])|(~m[673]&m[1048]&~m[1050]&m[1051]&m[1052])|(m[673]&m[1048]&~m[1050]&m[1051]&m[1052])|(~m[673]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[673]&~m[1048]&m[1050]&m[1051]&m[1052])|(m[673]&m[1048]&m[1050]&m[1051]&m[1052]));
    m[1054] = (((m[686]&~m[1053]&~m[1055]&~m[1056]&~m[1057])|(~m[686]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(m[686]&m[1053]&~m[1055]&m[1056]&~m[1057])|(m[686]&~m[1053]&m[1055]&m[1056]&~m[1057])|(~m[686]&m[1053]&~m[1055]&~m[1056]&m[1057])|(~m[686]&~m[1053]&m[1055]&~m[1056]&m[1057])|(m[686]&m[1053]&m[1055]&~m[1056]&m[1057])|(~m[686]&m[1053]&m[1055]&m[1056]&m[1057]))&UnbiasedRNG[269])|((m[686]&~m[1053]&~m[1055]&m[1056]&~m[1057])|(~m[686]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[686]&~m[1053]&~m[1055]&~m[1056]&m[1057])|(m[686]&m[1053]&~m[1055]&~m[1056]&m[1057])|(m[686]&~m[1053]&m[1055]&~m[1056]&m[1057])|(~m[686]&~m[1053]&~m[1055]&m[1056]&m[1057])|(m[686]&~m[1053]&~m[1055]&m[1056]&m[1057])|(~m[686]&m[1053]&~m[1055]&m[1056]&m[1057])|(m[686]&m[1053]&~m[1055]&m[1056]&m[1057])|(~m[686]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[686]&~m[1053]&m[1055]&m[1056]&m[1057])|(m[686]&m[1053]&m[1055]&m[1056]&m[1057]));
    m[1059] = (((m[557]&~m[1058]&~m[1060]&~m[1061]&~m[1062])|(~m[557]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(m[557]&m[1058]&~m[1060]&m[1061]&~m[1062])|(m[557]&~m[1058]&m[1060]&m[1061]&~m[1062])|(~m[557]&m[1058]&~m[1060]&~m[1061]&m[1062])|(~m[557]&~m[1058]&m[1060]&~m[1061]&m[1062])|(m[557]&m[1058]&m[1060]&~m[1061]&m[1062])|(~m[557]&m[1058]&m[1060]&m[1061]&m[1062]))&UnbiasedRNG[270])|((m[557]&~m[1058]&~m[1060]&m[1061]&~m[1062])|(~m[557]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[557]&~m[1058]&~m[1060]&~m[1061]&m[1062])|(m[557]&m[1058]&~m[1060]&~m[1061]&m[1062])|(m[557]&~m[1058]&m[1060]&~m[1061]&m[1062])|(~m[557]&~m[1058]&~m[1060]&m[1061]&m[1062])|(m[557]&~m[1058]&~m[1060]&m[1061]&m[1062])|(~m[557]&m[1058]&~m[1060]&m[1061]&m[1062])|(m[557]&m[1058]&~m[1060]&m[1061]&m[1062])|(~m[557]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[557]&~m[1058]&m[1060]&m[1061]&m[1062])|(m[557]&m[1058]&m[1060]&m[1061]&m[1062]));
    m[1064] = (((m[570]&~m[1063]&~m[1065]&~m[1066]&~m[1067])|(~m[570]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(m[570]&m[1063]&~m[1065]&m[1066]&~m[1067])|(m[570]&~m[1063]&m[1065]&m[1066]&~m[1067])|(~m[570]&m[1063]&~m[1065]&~m[1066]&m[1067])|(~m[570]&~m[1063]&m[1065]&~m[1066]&m[1067])|(m[570]&m[1063]&m[1065]&~m[1066]&m[1067])|(~m[570]&m[1063]&m[1065]&m[1066]&m[1067]))&UnbiasedRNG[271])|((m[570]&~m[1063]&~m[1065]&m[1066]&~m[1067])|(~m[570]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[570]&~m[1063]&~m[1065]&~m[1066]&m[1067])|(m[570]&m[1063]&~m[1065]&~m[1066]&m[1067])|(m[570]&~m[1063]&m[1065]&~m[1066]&m[1067])|(~m[570]&~m[1063]&~m[1065]&m[1066]&m[1067])|(m[570]&~m[1063]&~m[1065]&m[1066]&m[1067])|(~m[570]&m[1063]&~m[1065]&m[1066]&m[1067])|(m[570]&m[1063]&~m[1065]&m[1066]&m[1067])|(~m[570]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[570]&~m[1063]&m[1065]&m[1066]&m[1067])|(m[570]&m[1063]&m[1065]&m[1066]&m[1067]));
    m[1069] = (((m[583]&~m[1068]&~m[1070]&~m[1071]&~m[1072])|(~m[583]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(m[583]&m[1068]&~m[1070]&m[1071]&~m[1072])|(m[583]&~m[1068]&m[1070]&m[1071]&~m[1072])|(~m[583]&m[1068]&~m[1070]&~m[1071]&m[1072])|(~m[583]&~m[1068]&m[1070]&~m[1071]&m[1072])|(m[583]&m[1068]&m[1070]&~m[1071]&m[1072])|(~m[583]&m[1068]&m[1070]&m[1071]&m[1072]))&UnbiasedRNG[272])|((m[583]&~m[1068]&~m[1070]&m[1071]&~m[1072])|(~m[583]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[583]&~m[1068]&~m[1070]&~m[1071]&m[1072])|(m[583]&m[1068]&~m[1070]&~m[1071]&m[1072])|(m[583]&~m[1068]&m[1070]&~m[1071]&m[1072])|(~m[583]&~m[1068]&~m[1070]&m[1071]&m[1072])|(m[583]&~m[1068]&~m[1070]&m[1071]&m[1072])|(~m[583]&m[1068]&~m[1070]&m[1071]&m[1072])|(m[583]&m[1068]&~m[1070]&m[1071]&m[1072])|(~m[583]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[583]&~m[1068]&m[1070]&m[1071]&m[1072])|(m[583]&m[1068]&m[1070]&m[1071]&m[1072]));
    m[1074] = (((m[596]&~m[1073]&~m[1075]&~m[1076]&~m[1077])|(~m[596]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(m[596]&m[1073]&~m[1075]&m[1076]&~m[1077])|(m[596]&~m[1073]&m[1075]&m[1076]&~m[1077])|(~m[596]&m[1073]&~m[1075]&~m[1076]&m[1077])|(~m[596]&~m[1073]&m[1075]&~m[1076]&m[1077])|(m[596]&m[1073]&m[1075]&~m[1076]&m[1077])|(~m[596]&m[1073]&m[1075]&m[1076]&m[1077]))&UnbiasedRNG[273])|((m[596]&~m[1073]&~m[1075]&m[1076]&~m[1077])|(~m[596]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[596]&~m[1073]&~m[1075]&~m[1076]&m[1077])|(m[596]&m[1073]&~m[1075]&~m[1076]&m[1077])|(m[596]&~m[1073]&m[1075]&~m[1076]&m[1077])|(~m[596]&~m[1073]&~m[1075]&m[1076]&m[1077])|(m[596]&~m[1073]&~m[1075]&m[1076]&m[1077])|(~m[596]&m[1073]&~m[1075]&m[1076]&m[1077])|(m[596]&m[1073]&~m[1075]&m[1076]&m[1077])|(~m[596]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[596]&~m[1073]&m[1075]&m[1076]&m[1077])|(m[596]&m[1073]&m[1075]&m[1076]&m[1077]));
    m[1079] = (((m[609]&~m[1078]&~m[1080]&~m[1081]&~m[1082])|(~m[609]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(m[609]&m[1078]&~m[1080]&m[1081]&~m[1082])|(m[609]&~m[1078]&m[1080]&m[1081]&~m[1082])|(~m[609]&m[1078]&~m[1080]&~m[1081]&m[1082])|(~m[609]&~m[1078]&m[1080]&~m[1081]&m[1082])|(m[609]&m[1078]&m[1080]&~m[1081]&m[1082])|(~m[609]&m[1078]&m[1080]&m[1081]&m[1082]))&UnbiasedRNG[274])|((m[609]&~m[1078]&~m[1080]&m[1081]&~m[1082])|(~m[609]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[609]&~m[1078]&~m[1080]&~m[1081]&m[1082])|(m[609]&m[1078]&~m[1080]&~m[1081]&m[1082])|(m[609]&~m[1078]&m[1080]&~m[1081]&m[1082])|(~m[609]&~m[1078]&~m[1080]&m[1081]&m[1082])|(m[609]&~m[1078]&~m[1080]&m[1081]&m[1082])|(~m[609]&m[1078]&~m[1080]&m[1081]&m[1082])|(m[609]&m[1078]&~m[1080]&m[1081]&m[1082])|(~m[609]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[609]&~m[1078]&m[1080]&m[1081]&m[1082])|(m[609]&m[1078]&m[1080]&m[1081]&m[1082]));
    m[1084] = (((m[622]&~m[1083]&~m[1085]&~m[1086]&~m[1087])|(~m[622]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(m[622]&m[1083]&~m[1085]&m[1086]&~m[1087])|(m[622]&~m[1083]&m[1085]&m[1086]&~m[1087])|(~m[622]&m[1083]&~m[1085]&~m[1086]&m[1087])|(~m[622]&~m[1083]&m[1085]&~m[1086]&m[1087])|(m[622]&m[1083]&m[1085]&~m[1086]&m[1087])|(~m[622]&m[1083]&m[1085]&m[1086]&m[1087]))&UnbiasedRNG[275])|((m[622]&~m[1083]&~m[1085]&m[1086]&~m[1087])|(~m[622]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[622]&~m[1083]&~m[1085]&~m[1086]&m[1087])|(m[622]&m[1083]&~m[1085]&~m[1086]&m[1087])|(m[622]&~m[1083]&m[1085]&~m[1086]&m[1087])|(~m[622]&~m[1083]&~m[1085]&m[1086]&m[1087])|(m[622]&~m[1083]&~m[1085]&m[1086]&m[1087])|(~m[622]&m[1083]&~m[1085]&m[1086]&m[1087])|(m[622]&m[1083]&~m[1085]&m[1086]&m[1087])|(~m[622]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[622]&~m[1083]&m[1085]&m[1086]&m[1087])|(m[622]&m[1083]&m[1085]&m[1086]&m[1087]));
    m[1089] = (((m[635]&~m[1088]&~m[1090]&~m[1091]&~m[1092])|(~m[635]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(m[635]&m[1088]&~m[1090]&m[1091]&~m[1092])|(m[635]&~m[1088]&m[1090]&m[1091]&~m[1092])|(~m[635]&m[1088]&~m[1090]&~m[1091]&m[1092])|(~m[635]&~m[1088]&m[1090]&~m[1091]&m[1092])|(m[635]&m[1088]&m[1090]&~m[1091]&m[1092])|(~m[635]&m[1088]&m[1090]&m[1091]&m[1092]))&UnbiasedRNG[276])|((m[635]&~m[1088]&~m[1090]&m[1091]&~m[1092])|(~m[635]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[635]&~m[1088]&~m[1090]&~m[1091]&m[1092])|(m[635]&m[1088]&~m[1090]&~m[1091]&m[1092])|(m[635]&~m[1088]&m[1090]&~m[1091]&m[1092])|(~m[635]&~m[1088]&~m[1090]&m[1091]&m[1092])|(m[635]&~m[1088]&~m[1090]&m[1091]&m[1092])|(~m[635]&m[1088]&~m[1090]&m[1091]&m[1092])|(m[635]&m[1088]&~m[1090]&m[1091]&m[1092])|(~m[635]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[635]&~m[1088]&m[1090]&m[1091]&m[1092])|(m[635]&m[1088]&m[1090]&m[1091]&m[1092]));
    m[1094] = (((m[648]&~m[1093]&~m[1095]&~m[1096]&~m[1097])|(~m[648]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(m[648]&m[1093]&~m[1095]&m[1096]&~m[1097])|(m[648]&~m[1093]&m[1095]&m[1096]&~m[1097])|(~m[648]&m[1093]&~m[1095]&~m[1096]&m[1097])|(~m[648]&~m[1093]&m[1095]&~m[1096]&m[1097])|(m[648]&m[1093]&m[1095]&~m[1096]&m[1097])|(~m[648]&m[1093]&m[1095]&m[1096]&m[1097]))&UnbiasedRNG[277])|((m[648]&~m[1093]&~m[1095]&m[1096]&~m[1097])|(~m[648]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[648]&~m[1093]&~m[1095]&~m[1096]&m[1097])|(m[648]&m[1093]&~m[1095]&~m[1096]&m[1097])|(m[648]&~m[1093]&m[1095]&~m[1096]&m[1097])|(~m[648]&~m[1093]&~m[1095]&m[1096]&m[1097])|(m[648]&~m[1093]&~m[1095]&m[1096]&m[1097])|(~m[648]&m[1093]&~m[1095]&m[1096]&m[1097])|(m[648]&m[1093]&~m[1095]&m[1096]&m[1097])|(~m[648]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[648]&~m[1093]&m[1095]&m[1096]&m[1097])|(m[648]&m[1093]&m[1095]&m[1096]&m[1097]));
    m[1099] = (((m[661]&~m[1098]&~m[1100]&~m[1101]&~m[1102])|(~m[661]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(m[661]&m[1098]&~m[1100]&m[1101]&~m[1102])|(m[661]&~m[1098]&m[1100]&m[1101]&~m[1102])|(~m[661]&m[1098]&~m[1100]&~m[1101]&m[1102])|(~m[661]&~m[1098]&m[1100]&~m[1101]&m[1102])|(m[661]&m[1098]&m[1100]&~m[1101]&m[1102])|(~m[661]&m[1098]&m[1100]&m[1101]&m[1102]))&UnbiasedRNG[278])|((m[661]&~m[1098]&~m[1100]&m[1101]&~m[1102])|(~m[661]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[661]&~m[1098]&~m[1100]&~m[1101]&m[1102])|(m[661]&m[1098]&~m[1100]&~m[1101]&m[1102])|(m[661]&~m[1098]&m[1100]&~m[1101]&m[1102])|(~m[661]&~m[1098]&~m[1100]&m[1101]&m[1102])|(m[661]&~m[1098]&~m[1100]&m[1101]&m[1102])|(~m[661]&m[1098]&~m[1100]&m[1101]&m[1102])|(m[661]&m[1098]&~m[1100]&m[1101]&m[1102])|(~m[661]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[661]&~m[1098]&m[1100]&m[1101]&m[1102])|(m[661]&m[1098]&m[1100]&m[1101]&m[1102]));
    m[1104] = (((m[674]&~m[1103]&~m[1105]&~m[1106]&~m[1107])|(~m[674]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(m[674]&m[1103]&~m[1105]&m[1106]&~m[1107])|(m[674]&~m[1103]&m[1105]&m[1106]&~m[1107])|(~m[674]&m[1103]&~m[1105]&~m[1106]&m[1107])|(~m[674]&~m[1103]&m[1105]&~m[1106]&m[1107])|(m[674]&m[1103]&m[1105]&~m[1106]&m[1107])|(~m[674]&m[1103]&m[1105]&m[1106]&m[1107]))&UnbiasedRNG[279])|((m[674]&~m[1103]&~m[1105]&m[1106]&~m[1107])|(~m[674]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[674]&~m[1103]&~m[1105]&~m[1106]&m[1107])|(m[674]&m[1103]&~m[1105]&~m[1106]&m[1107])|(m[674]&~m[1103]&m[1105]&~m[1106]&m[1107])|(~m[674]&~m[1103]&~m[1105]&m[1106]&m[1107])|(m[674]&~m[1103]&~m[1105]&m[1106]&m[1107])|(~m[674]&m[1103]&~m[1105]&m[1106]&m[1107])|(m[674]&m[1103]&~m[1105]&m[1106]&m[1107])|(~m[674]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[674]&~m[1103]&m[1105]&m[1106]&m[1107])|(m[674]&m[1103]&m[1105]&m[1106]&m[1107]));
    m[1109] = (((m[687]&~m[1108]&~m[1110]&~m[1111]&~m[1112])|(~m[687]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(m[687]&m[1108]&~m[1110]&m[1111]&~m[1112])|(m[687]&~m[1108]&m[1110]&m[1111]&~m[1112])|(~m[687]&m[1108]&~m[1110]&~m[1111]&m[1112])|(~m[687]&~m[1108]&m[1110]&~m[1111]&m[1112])|(m[687]&m[1108]&m[1110]&~m[1111]&m[1112])|(~m[687]&m[1108]&m[1110]&m[1111]&m[1112]))&UnbiasedRNG[280])|((m[687]&~m[1108]&~m[1110]&m[1111]&~m[1112])|(~m[687]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[687]&~m[1108]&~m[1110]&~m[1111]&m[1112])|(m[687]&m[1108]&~m[1110]&~m[1111]&m[1112])|(m[687]&~m[1108]&m[1110]&~m[1111]&m[1112])|(~m[687]&~m[1108]&~m[1110]&m[1111]&m[1112])|(m[687]&~m[1108]&~m[1110]&m[1111]&m[1112])|(~m[687]&m[1108]&~m[1110]&m[1111]&m[1112])|(m[687]&m[1108]&~m[1110]&m[1111]&m[1112])|(~m[687]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[687]&~m[1108]&m[1110]&m[1111]&m[1112])|(m[687]&m[1108]&m[1110]&m[1111]&m[1112]));
    m[1114] = (((m[700]&~m[1113]&~m[1115]&~m[1116]&~m[1117])|(~m[700]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(m[700]&m[1113]&~m[1115]&m[1116]&~m[1117])|(m[700]&~m[1113]&m[1115]&m[1116]&~m[1117])|(~m[700]&m[1113]&~m[1115]&~m[1116]&m[1117])|(~m[700]&~m[1113]&m[1115]&~m[1116]&m[1117])|(m[700]&m[1113]&m[1115]&~m[1116]&m[1117])|(~m[700]&m[1113]&m[1115]&m[1116]&m[1117]))&UnbiasedRNG[281])|((m[700]&~m[1113]&~m[1115]&m[1116]&~m[1117])|(~m[700]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[700]&~m[1113]&~m[1115]&~m[1116]&m[1117])|(m[700]&m[1113]&~m[1115]&~m[1116]&m[1117])|(m[700]&~m[1113]&m[1115]&~m[1116]&m[1117])|(~m[700]&~m[1113]&~m[1115]&m[1116]&m[1117])|(m[700]&~m[1113]&~m[1115]&m[1116]&m[1117])|(~m[700]&m[1113]&~m[1115]&m[1116]&m[1117])|(m[700]&m[1113]&~m[1115]&m[1116]&m[1117])|(~m[700]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[700]&~m[1113]&m[1115]&m[1116]&m[1117])|(m[700]&m[1113]&m[1115]&m[1116]&m[1117]));
    m[1119] = (((m[558]&~m[1118]&~m[1120]&~m[1121]&~m[1122])|(~m[558]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(m[558]&m[1118]&~m[1120]&m[1121]&~m[1122])|(m[558]&~m[1118]&m[1120]&m[1121]&~m[1122])|(~m[558]&m[1118]&~m[1120]&~m[1121]&m[1122])|(~m[558]&~m[1118]&m[1120]&~m[1121]&m[1122])|(m[558]&m[1118]&m[1120]&~m[1121]&m[1122])|(~m[558]&m[1118]&m[1120]&m[1121]&m[1122]))&UnbiasedRNG[282])|((m[558]&~m[1118]&~m[1120]&m[1121]&~m[1122])|(~m[558]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[558]&~m[1118]&~m[1120]&~m[1121]&m[1122])|(m[558]&m[1118]&~m[1120]&~m[1121]&m[1122])|(m[558]&~m[1118]&m[1120]&~m[1121]&m[1122])|(~m[558]&~m[1118]&~m[1120]&m[1121]&m[1122])|(m[558]&~m[1118]&~m[1120]&m[1121]&m[1122])|(~m[558]&m[1118]&~m[1120]&m[1121]&m[1122])|(m[558]&m[1118]&~m[1120]&m[1121]&m[1122])|(~m[558]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[558]&~m[1118]&m[1120]&m[1121]&m[1122])|(m[558]&m[1118]&m[1120]&m[1121]&m[1122]));
    m[1124] = (((m[571]&~m[1123]&~m[1125]&~m[1126]&~m[1127])|(~m[571]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(m[571]&m[1123]&~m[1125]&m[1126]&~m[1127])|(m[571]&~m[1123]&m[1125]&m[1126]&~m[1127])|(~m[571]&m[1123]&~m[1125]&~m[1126]&m[1127])|(~m[571]&~m[1123]&m[1125]&~m[1126]&m[1127])|(m[571]&m[1123]&m[1125]&~m[1126]&m[1127])|(~m[571]&m[1123]&m[1125]&m[1126]&m[1127]))&UnbiasedRNG[283])|((m[571]&~m[1123]&~m[1125]&m[1126]&~m[1127])|(~m[571]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[571]&~m[1123]&~m[1125]&~m[1126]&m[1127])|(m[571]&m[1123]&~m[1125]&~m[1126]&m[1127])|(m[571]&~m[1123]&m[1125]&~m[1126]&m[1127])|(~m[571]&~m[1123]&~m[1125]&m[1126]&m[1127])|(m[571]&~m[1123]&~m[1125]&m[1126]&m[1127])|(~m[571]&m[1123]&~m[1125]&m[1126]&m[1127])|(m[571]&m[1123]&~m[1125]&m[1126]&m[1127])|(~m[571]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[571]&~m[1123]&m[1125]&m[1126]&m[1127])|(m[571]&m[1123]&m[1125]&m[1126]&m[1127]));
    m[1129] = (((m[584]&~m[1128]&~m[1130]&~m[1131]&~m[1132])|(~m[584]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(m[584]&m[1128]&~m[1130]&m[1131]&~m[1132])|(m[584]&~m[1128]&m[1130]&m[1131]&~m[1132])|(~m[584]&m[1128]&~m[1130]&~m[1131]&m[1132])|(~m[584]&~m[1128]&m[1130]&~m[1131]&m[1132])|(m[584]&m[1128]&m[1130]&~m[1131]&m[1132])|(~m[584]&m[1128]&m[1130]&m[1131]&m[1132]))&UnbiasedRNG[284])|((m[584]&~m[1128]&~m[1130]&m[1131]&~m[1132])|(~m[584]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[584]&~m[1128]&~m[1130]&~m[1131]&m[1132])|(m[584]&m[1128]&~m[1130]&~m[1131]&m[1132])|(m[584]&~m[1128]&m[1130]&~m[1131]&m[1132])|(~m[584]&~m[1128]&~m[1130]&m[1131]&m[1132])|(m[584]&~m[1128]&~m[1130]&m[1131]&m[1132])|(~m[584]&m[1128]&~m[1130]&m[1131]&m[1132])|(m[584]&m[1128]&~m[1130]&m[1131]&m[1132])|(~m[584]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[584]&~m[1128]&m[1130]&m[1131]&m[1132])|(m[584]&m[1128]&m[1130]&m[1131]&m[1132]));
    m[1134] = (((m[597]&~m[1133]&~m[1135]&~m[1136]&~m[1137])|(~m[597]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(m[597]&m[1133]&~m[1135]&m[1136]&~m[1137])|(m[597]&~m[1133]&m[1135]&m[1136]&~m[1137])|(~m[597]&m[1133]&~m[1135]&~m[1136]&m[1137])|(~m[597]&~m[1133]&m[1135]&~m[1136]&m[1137])|(m[597]&m[1133]&m[1135]&~m[1136]&m[1137])|(~m[597]&m[1133]&m[1135]&m[1136]&m[1137]))&UnbiasedRNG[285])|((m[597]&~m[1133]&~m[1135]&m[1136]&~m[1137])|(~m[597]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[597]&~m[1133]&~m[1135]&~m[1136]&m[1137])|(m[597]&m[1133]&~m[1135]&~m[1136]&m[1137])|(m[597]&~m[1133]&m[1135]&~m[1136]&m[1137])|(~m[597]&~m[1133]&~m[1135]&m[1136]&m[1137])|(m[597]&~m[1133]&~m[1135]&m[1136]&m[1137])|(~m[597]&m[1133]&~m[1135]&m[1136]&m[1137])|(m[597]&m[1133]&~m[1135]&m[1136]&m[1137])|(~m[597]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[597]&~m[1133]&m[1135]&m[1136]&m[1137])|(m[597]&m[1133]&m[1135]&m[1136]&m[1137]));
    m[1139] = (((m[610]&~m[1138]&~m[1140]&~m[1141]&~m[1142])|(~m[610]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(m[610]&m[1138]&~m[1140]&m[1141]&~m[1142])|(m[610]&~m[1138]&m[1140]&m[1141]&~m[1142])|(~m[610]&m[1138]&~m[1140]&~m[1141]&m[1142])|(~m[610]&~m[1138]&m[1140]&~m[1141]&m[1142])|(m[610]&m[1138]&m[1140]&~m[1141]&m[1142])|(~m[610]&m[1138]&m[1140]&m[1141]&m[1142]))&UnbiasedRNG[286])|((m[610]&~m[1138]&~m[1140]&m[1141]&~m[1142])|(~m[610]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[610]&~m[1138]&~m[1140]&~m[1141]&m[1142])|(m[610]&m[1138]&~m[1140]&~m[1141]&m[1142])|(m[610]&~m[1138]&m[1140]&~m[1141]&m[1142])|(~m[610]&~m[1138]&~m[1140]&m[1141]&m[1142])|(m[610]&~m[1138]&~m[1140]&m[1141]&m[1142])|(~m[610]&m[1138]&~m[1140]&m[1141]&m[1142])|(m[610]&m[1138]&~m[1140]&m[1141]&m[1142])|(~m[610]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[610]&~m[1138]&m[1140]&m[1141]&m[1142])|(m[610]&m[1138]&m[1140]&m[1141]&m[1142]));
    m[1144] = (((m[623]&~m[1143]&~m[1145]&~m[1146]&~m[1147])|(~m[623]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(m[623]&m[1143]&~m[1145]&m[1146]&~m[1147])|(m[623]&~m[1143]&m[1145]&m[1146]&~m[1147])|(~m[623]&m[1143]&~m[1145]&~m[1146]&m[1147])|(~m[623]&~m[1143]&m[1145]&~m[1146]&m[1147])|(m[623]&m[1143]&m[1145]&~m[1146]&m[1147])|(~m[623]&m[1143]&m[1145]&m[1146]&m[1147]))&UnbiasedRNG[287])|((m[623]&~m[1143]&~m[1145]&m[1146]&~m[1147])|(~m[623]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[623]&~m[1143]&~m[1145]&~m[1146]&m[1147])|(m[623]&m[1143]&~m[1145]&~m[1146]&m[1147])|(m[623]&~m[1143]&m[1145]&~m[1146]&m[1147])|(~m[623]&~m[1143]&~m[1145]&m[1146]&m[1147])|(m[623]&~m[1143]&~m[1145]&m[1146]&m[1147])|(~m[623]&m[1143]&~m[1145]&m[1146]&m[1147])|(m[623]&m[1143]&~m[1145]&m[1146]&m[1147])|(~m[623]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[623]&~m[1143]&m[1145]&m[1146]&m[1147])|(m[623]&m[1143]&m[1145]&m[1146]&m[1147]));
    m[1149] = (((m[636]&~m[1148]&~m[1150]&~m[1151]&~m[1152])|(~m[636]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(m[636]&m[1148]&~m[1150]&m[1151]&~m[1152])|(m[636]&~m[1148]&m[1150]&m[1151]&~m[1152])|(~m[636]&m[1148]&~m[1150]&~m[1151]&m[1152])|(~m[636]&~m[1148]&m[1150]&~m[1151]&m[1152])|(m[636]&m[1148]&m[1150]&~m[1151]&m[1152])|(~m[636]&m[1148]&m[1150]&m[1151]&m[1152]))&UnbiasedRNG[288])|((m[636]&~m[1148]&~m[1150]&m[1151]&~m[1152])|(~m[636]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[636]&~m[1148]&~m[1150]&~m[1151]&m[1152])|(m[636]&m[1148]&~m[1150]&~m[1151]&m[1152])|(m[636]&~m[1148]&m[1150]&~m[1151]&m[1152])|(~m[636]&~m[1148]&~m[1150]&m[1151]&m[1152])|(m[636]&~m[1148]&~m[1150]&m[1151]&m[1152])|(~m[636]&m[1148]&~m[1150]&m[1151]&m[1152])|(m[636]&m[1148]&~m[1150]&m[1151]&m[1152])|(~m[636]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[636]&~m[1148]&m[1150]&m[1151]&m[1152])|(m[636]&m[1148]&m[1150]&m[1151]&m[1152]));
    m[1154] = (((m[649]&~m[1153]&~m[1155]&~m[1156]&~m[1157])|(~m[649]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(m[649]&m[1153]&~m[1155]&m[1156]&~m[1157])|(m[649]&~m[1153]&m[1155]&m[1156]&~m[1157])|(~m[649]&m[1153]&~m[1155]&~m[1156]&m[1157])|(~m[649]&~m[1153]&m[1155]&~m[1156]&m[1157])|(m[649]&m[1153]&m[1155]&~m[1156]&m[1157])|(~m[649]&m[1153]&m[1155]&m[1156]&m[1157]))&UnbiasedRNG[289])|((m[649]&~m[1153]&~m[1155]&m[1156]&~m[1157])|(~m[649]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[649]&~m[1153]&~m[1155]&~m[1156]&m[1157])|(m[649]&m[1153]&~m[1155]&~m[1156]&m[1157])|(m[649]&~m[1153]&m[1155]&~m[1156]&m[1157])|(~m[649]&~m[1153]&~m[1155]&m[1156]&m[1157])|(m[649]&~m[1153]&~m[1155]&m[1156]&m[1157])|(~m[649]&m[1153]&~m[1155]&m[1156]&m[1157])|(m[649]&m[1153]&~m[1155]&m[1156]&m[1157])|(~m[649]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[649]&~m[1153]&m[1155]&m[1156]&m[1157])|(m[649]&m[1153]&m[1155]&m[1156]&m[1157]));
    m[1159] = (((m[662]&~m[1158]&~m[1160]&~m[1161]&~m[1162])|(~m[662]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(m[662]&m[1158]&~m[1160]&m[1161]&~m[1162])|(m[662]&~m[1158]&m[1160]&m[1161]&~m[1162])|(~m[662]&m[1158]&~m[1160]&~m[1161]&m[1162])|(~m[662]&~m[1158]&m[1160]&~m[1161]&m[1162])|(m[662]&m[1158]&m[1160]&~m[1161]&m[1162])|(~m[662]&m[1158]&m[1160]&m[1161]&m[1162]))&UnbiasedRNG[290])|((m[662]&~m[1158]&~m[1160]&m[1161]&~m[1162])|(~m[662]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[662]&~m[1158]&~m[1160]&~m[1161]&m[1162])|(m[662]&m[1158]&~m[1160]&~m[1161]&m[1162])|(m[662]&~m[1158]&m[1160]&~m[1161]&m[1162])|(~m[662]&~m[1158]&~m[1160]&m[1161]&m[1162])|(m[662]&~m[1158]&~m[1160]&m[1161]&m[1162])|(~m[662]&m[1158]&~m[1160]&m[1161]&m[1162])|(m[662]&m[1158]&~m[1160]&m[1161]&m[1162])|(~m[662]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[662]&~m[1158]&m[1160]&m[1161]&m[1162])|(m[662]&m[1158]&m[1160]&m[1161]&m[1162]));
    m[1164] = (((m[675]&~m[1163]&~m[1165]&~m[1166]&~m[1167])|(~m[675]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(m[675]&m[1163]&~m[1165]&m[1166]&~m[1167])|(m[675]&~m[1163]&m[1165]&m[1166]&~m[1167])|(~m[675]&m[1163]&~m[1165]&~m[1166]&m[1167])|(~m[675]&~m[1163]&m[1165]&~m[1166]&m[1167])|(m[675]&m[1163]&m[1165]&~m[1166]&m[1167])|(~m[675]&m[1163]&m[1165]&m[1166]&m[1167]))&UnbiasedRNG[291])|((m[675]&~m[1163]&~m[1165]&m[1166]&~m[1167])|(~m[675]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[675]&~m[1163]&~m[1165]&~m[1166]&m[1167])|(m[675]&m[1163]&~m[1165]&~m[1166]&m[1167])|(m[675]&~m[1163]&m[1165]&~m[1166]&m[1167])|(~m[675]&~m[1163]&~m[1165]&m[1166]&m[1167])|(m[675]&~m[1163]&~m[1165]&m[1166]&m[1167])|(~m[675]&m[1163]&~m[1165]&m[1166]&m[1167])|(m[675]&m[1163]&~m[1165]&m[1166]&m[1167])|(~m[675]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[675]&~m[1163]&m[1165]&m[1166]&m[1167])|(m[675]&m[1163]&m[1165]&m[1166]&m[1167]));
    m[1169] = (((m[688]&~m[1168]&~m[1170]&~m[1171]&~m[1172])|(~m[688]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(m[688]&m[1168]&~m[1170]&m[1171]&~m[1172])|(m[688]&~m[1168]&m[1170]&m[1171]&~m[1172])|(~m[688]&m[1168]&~m[1170]&~m[1171]&m[1172])|(~m[688]&~m[1168]&m[1170]&~m[1171]&m[1172])|(m[688]&m[1168]&m[1170]&~m[1171]&m[1172])|(~m[688]&m[1168]&m[1170]&m[1171]&m[1172]))&UnbiasedRNG[292])|((m[688]&~m[1168]&~m[1170]&m[1171]&~m[1172])|(~m[688]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[688]&~m[1168]&~m[1170]&~m[1171]&m[1172])|(m[688]&m[1168]&~m[1170]&~m[1171]&m[1172])|(m[688]&~m[1168]&m[1170]&~m[1171]&m[1172])|(~m[688]&~m[1168]&~m[1170]&m[1171]&m[1172])|(m[688]&~m[1168]&~m[1170]&m[1171]&m[1172])|(~m[688]&m[1168]&~m[1170]&m[1171]&m[1172])|(m[688]&m[1168]&~m[1170]&m[1171]&m[1172])|(~m[688]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[688]&~m[1168]&m[1170]&m[1171]&m[1172])|(m[688]&m[1168]&m[1170]&m[1171]&m[1172]));
    m[1174] = (((m[701]&~m[1173]&~m[1175]&~m[1176]&~m[1177])|(~m[701]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(m[701]&m[1173]&~m[1175]&m[1176]&~m[1177])|(m[701]&~m[1173]&m[1175]&m[1176]&~m[1177])|(~m[701]&m[1173]&~m[1175]&~m[1176]&m[1177])|(~m[701]&~m[1173]&m[1175]&~m[1176]&m[1177])|(m[701]&m[1173]&m[1175]&~m[1176]&m[1177])|(~m[701]&m[1173]&m[1175]&m[1176]&m[1177]))&UnbiasedRNG[293])|((m[701]&~m[1173]&~m[1175]&m[1176]&~m[1177])|(~m[701]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[701]&~m[1173]&~m[1175]&~m[1176]&m[1177])|(m[701]&m[1173]&~m[1175]&~m[1176]&m[1177])|(m[701]&~m[1173]&m[1175]&~m[1176]&m[1177])|(~m[701]&~m[1173]&~m[1175]&m[1176]&m[1177])|(m[701]&~m[1173]&~m[1175]&m[1176]&m[1177])|(~m[701]&m[1173]&~m[1175]&m[1176]&m[1177])|(m[701]&m[1173]&~m[1175]&m[1176]&m[1177])|(~m[701]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[701]&~m[1173]&m[1175]&m[1176]&m[1177])|(m[701]&m[1173]&m[1175]&m[1176]&m[1177]));
    m[1179] = (((m[714]&~m[1178]&~m[1180]&~m[1181]&~m[1182])|(~m[714]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(m[714]&m[1178]&~m[1180]&m[1181]&~m[1182])|(m[714]&~m[1178]&m[1180]&m[1181]&~m[1182])|(~m[714]&m[1178]&~m[1180]&~m[1181]&m[1182])|(~m[714]&~m[1178]&m[1180]&~m[1181]&m[1182])|(m[714]&m[1178]&m[1180]&~m[1181]&m[1182])|(~m[714]&m[1178]&m[1180]&m[1181]&m[1182]))&UnbiasedRNG[294])|((m[714]&~m[1178]&~m[1180]&m[1181]&~m[1182])|(~m[714]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[714]&~m[1178]&~m[1180]&~m[1181]&m[1182])|(m[714]&m[1178]&~m[1180]&~m[1181]&m[1182])|(m[714]&~m[1178]&m[1180]&~m[1181]&m[1182])|(~m[714]&~m[1178]&~m[1180]&m[1181]&m[1182])|(m[714]&~m[1178]&~m[1180]&m[1181]&m[1182])|(~m[714]&m[1178]&~m[1180]&m[1181]&m[1182])|(m[714]&m[1178]&~m[1180]&m[1181]&m[1182])|(~m[714]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[714]&~m[1178]&m[1180]&m[1181]&m[1182])|(m[714]&m[1178]&m[1180]&m[1181]&m[1182]));
    m[1184] = (((m[559]&~m[1183]&~m[1185]&~m[1186]&~m[1187])|(~m[559]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(m[559]&m[1183]&~m[1185]&m[1186]&~m[1187])|(m[559]&~m[1183]&m[1185]&m[1186]&~m[1187])|(~m[559]&m[1183]&~m[1185]&~m[1186]&m[1187])|(~m[559]&~m[1183]&m[1185]&~m[1186]&m[1187])|(m[559]&m[1183]&m[1185]&~m[1186]&m[1187])|(~m[559]&m[1183]&m[1185]&m[1186]&m[1187]))&UnbiasedRNG[295])|((m[559]&~m[1183]&~m[1185]&m[1186]&~m[1187])|(~m[559]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[559]&~m[1183]&~m[1185]&~m[1186]&m[1187])|(m[559]&m[1183]&~m[1185]&~m[1186]&m[1187])|(m[559]&~m[1183]&m[1185]&~m[1186]&m[1187])|(~m[559]&~m[1183]&~m[1185]&m[1186]&m[1187])|(m[559]&~m[1183]&~m[1185]&m[1186]&m[1187])|(~m[559]&m[1183]&~m[1185]&m[1186]&m[1187])|(m[559]&m[1183]&~m[1185]&m[1186]&m[1187])|(~m[559]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[559]&~m[1183]&m[1185]&m[1186]&m[1187])|(m[559]&m[1183]&m[1185]&m[1186]&m[1187]));
    m[1189] = (((m[572]&~m[1188]&~m[1190]&~m[1191]&~m[1192])|(~m[572]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(m[572]&m[1188]&~m[1190]&m[1191]&~m[1192])|(m[572]&~m[1188]&m[1190]&m[1191]&~m[1192])|(~m[572]&m[1188]&~m[1190]&~m[1191]&m[1192])|(~m[572]&~m[1188]&m[1190]&~m[1191]&m[1192])|(m[572]&m[1188]&m[1190]&~m[1191]&m[1192])|(~m[572]&m[1188]&m[1190]&m[1191]&m[1192]))&UnbiasedRNG[296])|((m[572]&~m[1188]&~m[1190]&m[1191]&~m[1192])|(~m[572]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[572]&~m[1188]&~m[1190]&~m[1191]&m[1192])|(m[572]&m[1188]&~m[1190]&~m[1191]&m[1192])|(m[572]&~m[1188]&m[1190]&~m[1191]&m[1192])|(~m[572]&~m[1188]&~m[1190]&m[1191]&m[1192])|(m[572]&~m[1188]&~m[1190]&m[1191]&m[1192])|(~m[572]&m[1188]&~m[1190]&m[1191]&m[1192])|(m[572]&m[1188]&~m[1190]&m[1191]&m[1192])|(~m[572]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[572]&~m[1188]&m[1190]&m[1191]&m[1192])|(m[572]&m[1188]&m[1190]&m[1191]&m[1192]));
    m[1194] = (((m[585]&~m[1193]&~m[1195]&~m[1196]&~m[1197])|(~m[585]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(m[585]&m[1193]&~m[1195]&m[1196]&~m[1197])|(m[585]&~m[1193]&m[1195]&m[1196]&~m[1197])|(~m[585]&m[1193]&~m[1195]&~m[1196]&m[1197])|(~m[585]&~m[1193]&m[1195]&~m[1196]&m[1197])|(m[585]&m[1193]&m[1195]&~m[1196]&m[1197])|(~m[585]&m[1193]&m[1195]&m[1196]&m[1197]))&UnbiasedRNG[297])|((m[585]&~m[1193]&~m[1195]&m[1196]&~m[1197])|(~m[585]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[585]&~m[1193]&~m[1195]&~m[1196]&m[1197])|(m[585]&m[1193]&~m[1195]&~m[1196]&m[1197])|(m[585]&~m[1193]&m[1195]&~m[1196]&m[1197])|(~m[585]&~m[1193]&~m[1195]&m[1196]&m[1197])|(m[585]&~m[1193]&~m[1195]&m[1196]&m[1197])|(~m[585]&m[1193]&~m[1195]&m[1196]&m[1197])|(m[585]&m[1193]&~m[1195]&m[1196]&m[1197])|(~m[585]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[585]&~m[1193]&m[1195]&m[1196]&m[1197])|(m[585]&m[1193]&m[1195]&m[1196]&m[1197]));
    m[1199] = (((m[598]&~m[1198]&~m[1200]&~m[1201]&~m[1202])|(~m[598]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(m[598]&m[1198]&~m[1200]&m[1201]&~m[1202])|(m[598]&~m[1198]&m[1200]&m[1201]&~m[1202])|(~m[598]&m[1198]&~m[1200]&~m[1201]&m[1202])|(~m[598]&~m[1198]&m[1200]&~m[1201]&m[1202])|(m[598]&m[1198]&m[1200]&~m[1201]&m[1202])|(~m[598]&m[1198]&m[1200]&m[1201]&m[1202]))&UnbiasedRNG[298])|((m[598]&~m[1198]&~m[1200]&m[1201]&~m[1202])|(~m[598]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[598]&~m[1198]&~m[1200]&~m[1201]&m[1202])|(m[598]&m[1198]&~m[1200]&~m[1201]&m[1202])|(m[598]&~m[1198]&m[1200]&~m[1201]&m[1202])|(~m[598]&~m[1198]&~m[1200]&m[1201]&m[1202])|(m[598]&~m[1198]&~m[1200]&m[1201]&m[1202])|(~m[598]&m[1198]&~m[1200]&m[1201]&m[1202])|(m[598]&m[1198]&~m[1200]&m[1201]&m[1202])|(~m[598]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[598]&~m[1198]&m[1200]&m[1201]&m[1202])|(m[598]&m[1198]&m[1200]&m[1201]&m[1202]));
    m[1204] = (((m[611]&~m[1203]&~m[1205]&~m[1206]&~m[1207])|(~m[611]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(m[611]&m[1203]&~m[1205]&m[1206]&~m[1207])|(m[611]&~m[1203]&m[1205]&m[1206]&~m[1207])|(~m[611]&m[1203]&~m[1205]&~m[1206]&m[1207])|(~m[611]&~m[1203]&m[1205]&~m[1206]&m[1207])|(m[611]&m[1203]&m[1205]&~m[1206]&m[1207])|(~m[611]&m[1203]&m[1205]&m[1206]&m[1207]))&UnbiasedRNG[299])|((m[611]&~m[1203]&~m[1205]&m[1206]&~m[1207])|(~m[611]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[611]&~m[1203]&~m[1205]&~m[1206]&m[1207])|(m[611]&m[1203]&~m[1205]&~m[1206]&m[1207])|(m[611]&~m[1203]&m[1205]&~m[1206]&m[1207])|(~m[611]&~m[1203]&~m[1205]&m[1206]&m[1207])|(m[611]&~m[1203]&~m[1205]&m[1206]&m[1207])|(~m[611]&m[1203]&~m[1205]&m[1206]&m[1207])|(m[611]&m[1203]&~m[1205]&m[1206]&m[1207])|(~m[611]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[611]&~m[1203]&m[1205]&m[1206]&m[1207])|(m[611]&m[1203]&m[1205]&m[1206]&m[1207]));
    m[1209] = (((m[624]&~m[1208]&~m[1210]&~m[1211]&~m[1212])|(~m[624]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(m[624]&m[1208]&~m[1210]&m[1211]&~m[1212])|(m[624]&~m[1208]&m[1210]&m[1211]&~m[1212])|(~m[624]&m[1208]&~m[1210]&~m[1211]&m[1212])|(~m[624]&~m[1208]&m[1210]&~m[1211]&m[1212])|(m[624]&m[1208]&m[1210]&~m[1211]&m[1212])|(~m[624]&m[1208]&m[1210]&m[1211]&m[1212]))&UnbiasedRNG[300])|((m[624]&~m[1208]&~m[1210]&m[1211]&~m[1212])|(~m[624]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[624]&~m[1208]&~m[1210]&~m[1211]&m[1212])|(m[624]&m[1208]&~m[1210]&~m[1211]&m[1212])|(m[624]&~m[1208]&m[1210]&~m[1211]&m[1212])|(~m[624]&~m[1208]&~m[1210]&m[1211]&m[1212])|(m[624]&~m[1208]&~m[1210]&m[1211]&m[1212])|(~m[624]&m[1208]&~m[1210]&m[1211]&m[1212])|(m[624]&m[1208]&~m[1210]&m[1211]&m[1212])|(~m[624]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[624]&~m[1208]&m[1210]&m[1211]&m[1212])|(m[624]&m[1208]&m[1210]&m[1211]&m[1212]));
    m[1214] = (((m[637]&~m[1213]&~m[1215]&~m[1216]&~m[1217])|(~m[637]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(m[637]&m[1213]&~m[1215]&m[1216]&~m[1217])|(m[637]&~m[1213]&m[1215]&m[1216]&~m[1217])|(~m[637]&m[1213]&~m[1215]&~m[1216]&m[1217])|(~m[637]&~m[1213]&m[1215]&~m[1216]&m[1217])|(m[637]&m[1213]&m[1215]&~m[1216]&m[1217])|(~m[637]&m[1213]&m[1215]&m[1216]&m[1217]))&UnbiasedRNG[301])|((m[637]&~m[1213]&~m[1215]&m[1216]&~m[1217])|(~m[637]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[637]&~m[1213]&~m[1215]&~m[1216]&m[1217])|(m[637]&m[1213]&~m[1215]&~m[1216]&m[1217])|(m[637]&~m[1213]&m[1215]&~m[1216]&m[1217])|(~m[637]&~m[1213]&~m[1215]&m[1216]&m[1217])|(m[637]&~m[1213]&~m[1215]&m[1216]&m[1217])|(~m[637]&m[1213]&~m[1215]&m[1216]&m[1217])|(m[637]&m[1213]&~m[1215]&m[1216]&m[1217])|(~m[637]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[637]&~m[1213]&m[1215]&m[1216]&m[1217])|(m[637]&m[1213]&m[1215]&m[1216]&m[1217]));
    m[1219] = (((m[650]&~m[1218]&~m[1220]&~m[1221]&~m[1222])|(~m[650]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(m[650]&m[1218]&~m[1220]&m[1221]&~m[1222])|(m[650]&~m[1218]&m[1220]&m[1221]&~m[1222])|(~m[650]&m[1218]&~m[1220]&~m[1221]&m[1222])|(~m[650]&~m[1218]&m[1220]&~m[1221]&m[1222])|(m[650]&m[1218]&m[1220]&~m[1221]&m[1222])|(~m[650]&m[1218]&m[1220]&m[1221]&m[1222]))&UnbiasedRNG[302])|((m[650]&~m[1218]&~m[1220]&m[1221]&~m[1222])|(~m[650]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[650]&~m[1218]&~m[1220]&~m[1221]&m[1222])|(m[650]&m[1218]&~m[1220]&~m[1221]&m[1222])|(m[650]&~m[1218]&m[1220]&~m[1221]&m[1222])|(~m[650]&~m[1218]&~m[1220]&m[1221]&m[1222])|(m[650]&~m[1218]&~m[1220]&m[1221]&m[1222])|(~m[650]&m[1218]&~m[1220]&m[1221]&m[1222])|(m[650]&m[1218]&~m[1220]&m[1221]&m[1222])|(~m[650]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[650]&~m[1218]&m[1220]&m[1221]&m[1222])|(m[650]&m[1218]&m[1220]&m[1221]&m[1222]));
    m[1224] = (((m[663]&~m[1223]&~m[1225]&~m[1226]&~m[1227])|(~m[663]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(m[663]&m[1223]&~m[1225]&m[1226]&~m[1227])|(m[663]&~m[1223]&m[1225]&m[1226]&~m[1227])|(~m[663]&m[1223]&~m[1225]&~m[1226]&m[1227])|(~m[663]&~m[1223]&m[1225]&~m[1226]&m[1227])|(m[663]&m[1223]&m[1225]&~m[1226]&m[1227])|(~m[663]&m[1223]&m[1225]&m[1226]&m[1227]))&UnbiasedRNG[303])|((m[663]&~m[1223]&~m[1225]&m[1226]&~m[1227])|(~m[663]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[663]&~m[1223]&~m[1225]&~m[1226]&m[1227])|(m[663]&m[1223]&~m[1225]&~m[1226]&m[1227])|(m[663]&~m[1223]&m[1225]&~m[1226]&m[1227])|(~m[663]&~m[1223]&~m[1225]&m[1226]&m[1227])|(m[663]&~m[1223]&~m[1225]&m[1226]&m[1227])|(~m[663]&m[1223]&~m[1225]&m[1226]&m[1227])|(m[663]&m[1223]&~m[1225]&m[1226]&m[1227])|(~m[663]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[663]&~m[1223]&m[1225]&m[1226]&m[1227])|(m[663]&m[1223]&m[1225]&m[1226]&m[1227]));
    m[1229] = (((m[676]&~m[1228]&~m[1230]&~m[1231]&~m[1232])|(~m[676]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(m[676]&m[1228]&~m[1230]&m[1231]&~m[1232])|(m[676]&~m[1228]&m[1230]&m[1231]&~m[1232])|(~m[676]&m[1228]&~m[1230]&~m[1231]&m[1232])|(~m[676]&~m[1228]&m[1230]&~m[1231]&m[1232])|(m[676]&m[1228]&m[1230]&~m[1231]&m[1232])|(~m[676]&m[1228]&m[1230]&m[1231]&m[1232]))&UnbiasedRNG[304])|((m[676]&~m[1228]&~m[1230]&m[1231]&~m[1232])|(~m[676]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[676]&~m[1228]&~m[1230]&~m[1231]&m[1232])|(m[676]&m[1228]&~m[1230]&~m[1231]&m[1232])|(m[676]&~m[1228]&m[1230]&~m[1231]&m[1232])|(~m[676]&~m[1228]&~m[1230]&m[1231]&m[1232])|(m[676]&~m[1228]&~m[1230]&m[1231]&m[1232])|(~m[676]&m[1228]&~m[1230]&m[1231]&m[1232])|(m[676]&m[1228]&~m[1230]&m[1231]&m[1232])|(~m[676]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[676]&~m[1228]&m[1230]&m[1231]&m[1232])|(m[676]&m[1228]&m[1230]&m[1231]&m[1232]));
    m[1234] = (((m[689]&~m[1233]&~m[1235]&~m[1236]&~m[1237])|(~m[689]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(m[689]&m[1233]&~m[1235]&m[1236]&~m[1237])|(m[689]&~m[1233]&m[1235]&m[1236]&~m[1237])|(~m[689]&m[1233]&~m[1235]&~m[1236]&m[1237])|(~m[689]&~m[1233]&m[1235]&~m[1236]&m[1237])|(m[689]&m[1233]&m[1235]&~m[1236]&m[1237])|(~m[689]&m[1233]&m[1235]&m[1236]&m[1237]))&UnbiasedRNG[305])|((m[689]&~m[1233]&~m[1235]&m[1236]&~m[1237])|(~m[689]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[689]&~m[1233]&~m[1235]&~m[1236]&m[1237])|(m[689]&m[1233]&~m[1235]&~m[1236]&m[1237])|(m[689]&~m[1233]&m[1235]&~m[1236]&m[1237])|(~m[689]&~m[1233]&~m[1235]&m[1236]&m[1237])|(m[689]&~m[1233]&~m[1235]&m[1236]&m[1237])|(~m[689]&m[1233]&~m[1235]&m[1236]&m[1237])|(m[689]&m[1233]&~m[1235]&m[1236]&m[1237])|(~m[689]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[689]&~m[1233]&m[1235]&m[1236]&m[1237])|(m[689]&m[1233]&m[1235]&m[1236]&m[1237]));
    m[1239] = (((m[702]&~m[1238]&~m[1240]&~m[1241]&~m[1242])|(~m[702]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(m[702]&m[1238]&~m[1240]&m[1241]&~m[1242])|(m[702]&~m[1238]&m[1240]&m[1241]&~m[1242])|(~m[702]&m[1238]&~m[1240]&~m[1241]&m[1242])|(~m[702]&~m[1238]&m[1240]&~m[1241]&m[1242])|(m[702]&m[1238]&m[1240]&~m[1241]&m[1242])|(~m[702]&m[1238]&m[1240]&m[1241]&m[1242]))&UnbiasedRNG[306])|((m[702]&~m[1238]&~m[1240]&m[1241]&~m[1242])|(~m[702]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[702]&~m[1238]&~m[1240]&~m[1241]&m[1242])|(m[702]&m[1238]&~m[1240]&~m[1241]&m[1242])|(m[702]&~m[1238]&m[1240]&~m[1241]&m[1242])|(~m[702]&~m[1238]&~m[1240]&m[1241]&m[1242])|(m[702]&~m[1238]&~m[1240]&m[1241]&m[1242])|(~m[702]&m[1238]&~m[1240]&m[1241]&m[1242])|(m[702]&m[1238]&~m[1240]&m[1241]&m[1242])|(~m[702]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[702]&~m[1238]&m[1240]&m[1241]&m[1242])|(m[702]&m[1238]&m[1240]&m[1241]&m[1242]));
    m[1244] = (((m[715]&~m[1243]&~m[1245]&~m[1246]&~m[1247])|(~m[715]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(m[715]&m[1243]&~m[1245]&m[1246]&~m[1247])|(m[715]&~m[1243]&m[1245]&m[1246]&~m[1247])|(~m[715]&m[1243]&~m[1245]&~m[1246]&m[1247])|(~m[715]&~m[1243]&m[1245]&~m[1246]&m[1247])|(m[715]&m[1243]&m[1245]&~m[1246]&m[1247])|(~m[715]&m[1243]&m[1245]&m[1246]&m[1247]))&UnbiasedRNG[307])|((m[715]&~m[1243]&~m[1245]&m[1246]&~m[1247])|(~m[715]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[715]&~m[1243]&~m[1245]&~m[1246]&m[1247])|(m[715]&m[1243]&~m[1245]&~m[1246]&m[1247])|(m[715]&~m[1243]&m[1245]&~m[1246]&m[1247])|(~m[715]&~m[1243]&~m[1245]&m[1246]&m[1247])|(m[715]&~m[1243]&~m[1245]&m[1246]&m[1247])|(~m[715]&m[1243]&~m[1245]&m[1246]&m[1247])|(m[715]&m[1243]&~m[1245]&m[1246]&m[1247])|(~m[715]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[715]&~m[1243]&m[1245]&m[1246]&m[1247])|(m[715]&m[1243]&m[1245]&m[1246]&m[1247]));
    m[1249] = (((m[573]&~m[1248]&~m[1250]&~m[1251]&~m[1252])|(~m[573]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(m[573]&m[1248]&~m[1250]&m[1251]&~m[1252])|(m[573]&~m[1248]&m[1250]&m[1251]&~m[1252])|(~m[573]&m[1248]&~m[1250]&~m[1251]&m[1252])|(~m[573]&~m[1248]&m[1250]&~m[1251]&m[1252])|(m[573]&m[1248]&m[1250]&~m[1251]&m[1252])|(~m[573]&m[1248]&m[1250]&m[1251]&m[1252]))&UnbiasedRNG[308])|((m[573]&~m[1248]&~m[1250]&m[1251]&~m[1252])|(~m[573]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[573]&~m[1248]&~m[1250]&~m[1251]&m[1252])|(m[573]&m[1248]&~m[1250]&~m[1251]&m[1252])|(m[573]&~m[1248]&m[1250]&~m[1251]&m[1252])|(~m[573]&~m[1248]&~m[1250]&m[1251]&m[1252])|(m[573]&~m[1248]&~m[1250]&m[1251]&m[1252])|(~m[573]&m[1248]&~m[1250]&m[1251]&m[1252])|(m[573]&m[1248]&~m[1250]&m[1251]&m[1252])|(~m[573]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[573]&~m[1248]&m[1250]&m[1251]&m[1252])|(m[573]&m[1248]&m[1250]&m[1251]&m[1252]));
    m[1254] = (((m[586]&~m[1253]&~m[1255]&~m[1256]&~m[1257])|(~m[586]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(m[586]&m[1253]&~m[1255]&m[1256]&~m[1257])|(m[586]&~m[1253]&m[1255]&m[1256]&~m[1257])|(~m[586]&m[1253]&~m[1255]&~m[1256]&m[1257])|(~m[586]&~m[1253]&m[1255]&~m[1256]&m[1257])|(m[586]&m[1253]&m[1255]&~m[1256]&m[1257])|(~m[586]&m[1253]&m[1255]&m[1256]&m[1257]))&UnbiasedRNG[309])|((m[586]&~m[1253]&~m[1255]&m[1256]&~m[1257])|(~m[586]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[586]&~m[1253]&~m[1255]&~m[1256]&m[1257])|(m[586]&m[1253]&~m[1255]&~m[1256]&m[1257])|(m[586]&~m[1253]&m[1255]&~m[1256]&m[1257])|(~m[586]&~m[1253]&~m[1255]&m[1256]&m[1257])|(m[586]&~m[1253]&~m[1255]&m[1256]&m[1257])|(~m[586]&m[1253]&~m[1255]&m[1256]&m[1257])|(m[586]&m[1253]&~m[1255]&m[1256]&m[1257])|(~m[586]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[586]&~m[1253]&m[1255]&m[1256]&m[1257])|(m[586]&m[1253]&m[1255]&m[1256]&m[1257]));
    m[1259] = (((m[599]&~m[1258]&~m[1260]&~m[1261]&~m[1262])|(~m[599]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(m[599]&m[1258]&~m[1260]&m[1261]&~m[1262])|(m[599]&~m[1258]&m[1260]&m[1261]&~m[1262])|(~m[599]&m[1258]&~m[1260]&~m[1261]&m[1262])|(~m[599]&~m[1258]&m[1260]&~m[1261]&m[1262])|(m[599]&m[1258]&m[1260]&~m[1261]&m[1262])|(~m[599]&m[1258]&m[1260]&m[1261]&m[1262]))&UnbiasedRNG[310])|((m[599]&~m[1258]&~m[1260]&m[1261]&~m[1262])|(~m[599]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[599]&~m[1258]&~m[1260]&~m[1261]&m[1262])|(m[599]&m[1258]&~m[1260]&~m[1261]&m[1262])|(m[599]&~m[1258]&m[1260]&~m[1261]&m[1262])|(~m[599]&~m[1258]&~m[1260]&m[1261]&m[1262])|(m[599]&~m[1258]&~m[1260]&m[1261]&m[1262])|(~m[599]&m[1258]&~m[1260]&m[1261]&m[1262])|(m[599]&m[1258]&~m[1260]&m[1261]&m[1262])|(~m[599]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[599]&~m[1258]&m[1260]&m[1261]&m[1262])|(m[599]&m[1258]&m[1260]&m[1261]&m[1262]));
    m[1264] = (((m[612]&~m[1263]&~m[1265]&~m[1266]&~m[1267])|(~m[612]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(m[612]&m[1263]&~m[1265]&m[1266]&~m[1267])|(m[612]&~m[1263]&m[1265]&m[1266]&~m[1267])|(~m[612]&m[1263]&~m[1265]&~m[1266]&m[1267])|(~m[612]&~m[1263]&m[1265]&~m[1266]&m[1267])|(m[612]&m[1263]&m[1265]&~m[1266]&m[1267])|(~m[612]&m[1263]&m[1265]&m[1266]&m[1267]))&UnbiasedRNG[311])|((m[612]&~m[1263]&~m[1265]&m[1266]&~m[1267])|(~m[612]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[612]&~m[1263]&~m[1265]&~m[1266]&m[1267])|(m[612]&m[1263]&~m[1265]&~m[1266]&m[1267])|(m[612]&~m[1263]&m[1265]&~m[1266]&m[1267])|(~m[612]&~m[1263]&~m[1265]&m[1266]&m[1267])|(m[612]&~m[1263]&~m[1265]&m[1266]&m[1267])|(~m[612]&m[1263]&~m[1265]&m[1266]&m[1267])|(m[612]&m[1263]&~m[1265]&m[1266]&m[1267])|(~m[612]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[612]&~m[1263]&m[1265]&m[1266]&m[1267])|(m[612]&m[1263]&m[1265]&m[1266]&m[1267]));
    m[1269] = (((m[625]&~m[1268]&~m[1270]&~m[1271]&~m[1272])|(~m[625]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(m[625]&m[1268]&~m[1270]&m[1271]&~m[1272])|(m[625]&~m[1268]&m[1270]&m[1271]&~m[1272])|(~m[625]&m[1268]&~m[1270]&~m[1271]&m[1272])|(~m[625]&~m[1268]&m[1270]&~m[1271]&m[1272])|(m[625]&m[1268]&m[1270]&~m[1271]&m[1272])|(~m[625]&m[1268]&m[1270]&m[1271]&m[1272]))&UnbiasedRNG[312])|((m[625]&~m[1268]&~m[1270]&m[1271]&~m[1272])|(~m[625]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[625]&~m[1268]&~m[1270]&~m[1271]&m[1272])|(m[625]&m[1268]&~m[1270]&~m[1271]&m[1272])|(m[625]&~m[1268]&m[1270]&~m[1271]&m[1272])|(~m[625]&~m[1268]&~m[1270]&m[1271]&m[1272])|(m[625]&~m[1268]&~m[1270]&m[1271]&m[1272])|(~m[625]&m[1268]&~m[1270]&m[1271]&m[1272])|(m[625]&m[1268]&~m[1270]&m[1271]&m[1272])|(~m[625]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[625]&~m[1268]&m[1270]&m[1271]&m[1272])|(m[625]&m[1268]&m[1270]&m[1271]&m[1272]));
    m[1274] = (((m[638]&~m[1273]&~m[1275]&~m[1276]&~m[1277])|(~m[638]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(m[638]&m[1273]&~m[1275]&m[1276]&~m[1277])|(m[638]&~m[1273]&m[1275]&m[1276]&~m[1277])|(~m[638]&m[1273]&~m[1275]&~m[1276]&m[1277])|(~m[638]&~m[1273]&m[1275]&~m[1276]&m[1277])|(m[638]&m[1273]&m[1275]&~m[1276]&m[1277])|(~m[638]&m[1273]&m[1275]&m[1276]&m[1277]))&UnbiasedRNG[313])|((m[638]&~m[1273]&~m[1275]&m[1276]&~m[1277])|(~m[638]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[638]&~m[1273]&~m[1275]&~m[1276]&m[1277])|(m[638]&m[1273]&~m[1275]&~m[1276]&m[1277])|(m[638]&~m[1273]&m[1275]&~m[1276]&m[1277])|(~m[638]&~m[1273]&~m[1275]&m[1276]&m[1277])|(m[638]&~m[1273]&~m[1275]&m[1276]&m[1277])|(~m[638]&m[1273]&~m[1275]&m[1276]&m[1277])|(m[638]&m[1273]&~m[1275]&m[1276]&m[1277])|(~m[638]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[638]&~m[1273]&m[1275]&m[1276]&m[1277])|(m[638]&m[1273]&m[1275]&m[1276]&m[1277]));
    m[1279] = (((m[651]&~m[1278]&~m[1280]&~m[1281]&~m[1282])|(~m[651]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(m[651]&m[1278]&~m[1280]&m[1281]&~m[1282])|(m[651]&~m[1278]&m[1280]&m[1281]&~m[1282])|(~m[651]&m[1278]&~m[1280]&~m[1281]&m[1282])|(~m[651]&~m[1278]&m[1280]&~m[1281]&m[1282])|(m[651]&m[1278]&m[1280]&~m[1281]&m[1282])|(~m[651]&m[1278]&m[1280]&m[1281]&m[1282]))&UnbiasedRNG[314])|((m[651]&~m[1278]&~m[1280]&m[1281]&~m[1282])|(~m[651]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[651]&~m[1278]&~m[1280]&~m[1281]&m[1282])|(m[651]&m[1278]&~m[1280]&~m[1281]&m[1282])|(m[651]&~m[1278]&m[1280]&~m[1281]&m[1282])|(~m[651]&~m[1278]&~m[1280]&m[1281]&m[1282])|(m[651]&~m[1278]&~m[1280]&m[1281]&m[1282])|(~m[651]&m[1278]&~m[1280]&m[1281]&m[1282])|(m[651]&m[1278]&~m[1280]&m[1281]&m[1282])|(~m[651]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[651]&~m[1278]&m[1280]&m[1281]&m[1282])|(m[651]&m[1278]&m[1280]&m[1281]&m[1282]));
    m[1284] = (((m[664]&~m[1283]&~m[1285]&~m[1286]&~m[1287])|(~m[664]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(m[664]&m[1283]&~m[1285]&m[1286]&~m[1287])|(m[664]&~m[1283]&m[1285]&m[1286]&~m[1287])|(~m[664]&m[1283]&~m[1285]&~m[1286]&m[1287])|(~m[664]&~m[1283]&m[1285]&~m[1286]&m[1287])|(m[664]&m[1283]&m[1285]&~m[1286]&m[1287])|(~m[664]&m[1283]&m[1285]&m[1286]&m[1287]))&UnbiasedRNG[315])|((m[664]&~m[1283]&~m[1285]&m[1286]&~m[1287])|(~m[664]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[664]&~m[1283]&~m[1285]&~m[1286]&m[1287])|(m[664]&m[1283]&~m[1285]&~m[1286]&m[1287])|(m[664]&~m[1283]&m[1285]&~m[1286]&m[1287])|(~m[664]&~m[1283]&~m[1285]&m[1286]&m[1287])|(m[664]&~m[1283]&~m[1285]&m[1286]&m[1287])|(~m[664]&m[1283]&~m[1285]&m[1286]&m[1287])|(m[664]&m[1283]&~m[1285]&m[1286]&m[1287])|(~m[664]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[664]&~m[1283]&m[1285]&m[1286]&m[1287])|(m[664]&m[1283]&m[1285]&m[1286]&m[1287]));
    m[1289] = (((m[677]&~m[1288]&~m[1290]&~m[1291]&~m[1292])|(~m[677]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(m[677]&m[1288]&~m[1290]&m[1291]&~m[1292])|(m[677]&~m[1288]&m[1290]&m[1291]&~m[1292])|(~m[677]&m[1288]&~m[1290]&~m[1291]&m[1292])|(~m[677]&~m[1288]&m[1290]&~m[1291]&m[1292])|(m[677]&m[1288]&m[1290]&~m[1291]&m[1292])|(~m[677]&m[1288]&m[1290]&m[1291]&m[1292]))&UnbiasedRNG[316])|((m[677]&~m[1288]&~m[1290]&m[1291]&~m[1292])|(~m[677]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[677]&~m[1288]&~m[1290]&~m[1291]&m[1292])|(m[677]&m[1288]&~m[1290]&~m[1291]&m[1292])|(m[677]&~m[1288]&m[1290]&~m[1291]&m[1292])|(~m[677]&~m[1288]&~m[1290]&m[1291]&m[1292])|(m[677]&~m[1288]&~m[1290]&m[1291]&m[1292])|(~m[677]&m[1288]&~m[1290]&m[1291]&m[1292])|(m[677]&m[1288]&~m[1290]&m[1291]&m[1292])|(~m[677]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[677]&~m[1288]&m[1290]&m[1291]&m[1292])|(m[677]&m[1288]&m[1290]&m[1291]&m[1292]));
    m[1294] = (((m[690]&~m[1293]&~m[1295]&~m[1296]&~m[1297])|(~m[690]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(m[690]&m[1293]&~m[1295]&m[1296]&~m[1297])|(m[690]&~m[1293]&m[1295]&m[1296]&~m[1297])|(~m[690]&m[1293]&~m[1295]&~m[1296]&m[1297])|(~m[690]&~m[1293]&m[1295]&~m[1296]&m[1297])|(m[690]&m[1293]&m[1295]&~m[1296]&m[1297])|(~m[690]&m[1293]&m[1295]&m[1296]&m[1297]))&UnbiasedRNG[317])|((m[690]&~m[1293]&~m[1295]&m[1296]&~m[1297])|(~m[690]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[690]&~m[1293]&~m[1295]&~m[1296]&m[1297])|(m[690]&m[1293]&~m[1295]&~m[1296]&m[1297])|(m[690]&~m[1293]&m[1295]&~m[1296]&m[1297])|(~m[690]&~m[1293]&~m[1295]&m[1296]&m[1297])|(m[690]&~m[1293]&~m[1295]&m[1296]&m[1297])|(~m[690]&m[1293]&~m[1295]&m[1296]&m[1297])|(m[690]&m[1293]&~m[1295]&m[1296]&m[1297])|(~m[690]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[690]&~m[1293]&m[1295]&m[1296]&m[1297])|(m[690]&m[1293]&m[1295]&m[1296]&m[1297]));
    m[1299] = (((m[703]&~m[1298]&~m[1300]&~m[1301]&~m[1302])|(~m[703]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(m[703]&m[1298]&~m[1300]&m[1301]&~m[1302])|(m[703]&~m[1298]&m[1300]&m[1301]&~m[1302])|(~m[703]&m[1298]&~m[1300]&~m[1301]&m[1302])|(~m[703]&~m[1298]&m[1300]&~m[1301]&m[1302])|(m[703]&m[1298]&m[1300]&~m[1301]&m[1302])|(~m[703]&m[1298]&m[1300]&m[1301]&m[1302]))&UnbiasedRNG[318])|((m[703]&~m[1298]&~m[1300]&m[1301]&~m[1302])|(~m[703]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[703]&~m[1298]&~m[1300]&~m[1301]&m[1302])|(m[703]&m[1298]&~m[1300]&~m[1301]&m[1302])|(m[703]&~m[1298]&m[1300]&~m[1301]&m[1302])|(~m[703]&~m[1298]&~m[1300]&m[1301]&m[1302])|(m[703]&~m[1298]&~m[1300]&m[1301]&m[1302])|(~m[703]&m[1298]&~m[1300]&m[1301]&m[1302])|(m[703]&m[1298]&~m[1300]&m[1301]&m[1302])|(~m[703]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[703]&~m[1298]&m[1300]&m[1301]&m[1302])|(m[703]&m[1298]&m[1300]&m[1301]&m[1302]));
    m[1304] = (((m[716]&~m[1303]&~m[1305]&~m[1306]&~m[1307])|(~m[716]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(m[716]&m[1303]&~m[1305]&m[1306]&~m[1307])|(m[716]&~m[1303]&m[1305]&m[1306]&~m[1307])|(~m[716]&m[1303]&~m[1305]&~m[1306]&m[1307])|(~m[716]&~m[1303]&m[1305]&~m[1306]&m[1307])|(m[716]&m[1303]&m[1305]&~m[1306]&m[1307])|(~m[716]&m[1303]&m[1305]&m[1306]&m[1307]))&UnbiasedRNG[319])|((m[716]&~m[1303]&~m[1305]&m[1306]&~m[1307])|(~m[716]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[716]&~m[1303]&~m[1305]&~m[1306]&m[1307])|(m[716]&m[1303]&~m[1305]&~m[1306]&m[1307])|(m[716]&~m[1303]&m[1305]&~m[1306]&m[1307])|(~m[716]&~m[1303]&~m[1305]&m[1306]&m[1307])|(m[716]&~m[1303]&~m[1305]&m[1306]&m[1307])|(~m[716]&m[1303]&~m[1305]&m[1306]&m[1307])|(m[716]&m[1303]&~m[1305]&m[1306]&m[1307])|(~m[716]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[716]&~m[1303]&m[1305]&m[1306]&m[1307])|(m[716]&m[1303]&m[1305]&m[1306]&m[1307]));
    m[1309] = (((m[587]&~m[1308]&~m[1310]&~m[1311]&~m[1312])|(~m[587]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(m[587]&m[1308]&~m[1310]&m[1311]&~m[1312])|(m[587]&~m[1308]&m[1310]&m[1311]&~m[1312])|(~m[587]&m[1308]&~m[1310]&~m[1311]&m[1312])|(~m[587]&~m[1308]&m[1310]&~m[1311]&m[1312])|(m[587]&m[1308]&m[1310]&~m[1311]&m[1312])|(~m[587]&m[1308]&m[1310]&m[1311]&m[1312]))&UnbiasedRNG[320])|((m[587]&~m[1308]&~m[1310]&m[1311]&~m[1312])|(~m[587]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[587]&~m[1308]&~m[1310]&~m[1311]&m[1312])|(m[587]&m[1308]&~m[1310]&~m[1311]&m[1312])|(m[587]&~m[1308]&m[1310]&~m[1311]&m[1312])|(~m[587]&~m[1308]&~m[1310]&m[1311]&m[1312])|(m[587]&~m[1308]&~m[1310]&m[1311]&m[1312])|(~m[587]&m[1308]&~m[1310]&m[1311]&m[1312])|(m[587]&m[1308]&~m[1310]&m[1311]&m[1312])|(~m[587]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[587]&~m[1308]&m[1310]&m[1311]&m[1312])|(m[587]&m[1308]&m[1310]&m[1311]&m[1312]));
    m[1314] = (((m[600]&~m[1313]&~m[1315]&~m[1316]&~m[1317])|(~m[600]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(m[600]&m[1313]&~m[1315]&m[1316]&~m[1317])|(m[600]&~m[1313]&m[1315]&m[1316]&~m[1317])|(~m[600]&m[1313]&~m[1315]&~m[1316]&m[1317])|(~m[600]&~m[1313]&m[1315]&~m[1316]&m[1317])|(m[600]&m[1313]&m[1315]&~m[1316]&m[1317])|(~m[600]&m[1313]&m[1315]&m[1316]&m[1317]))&UnbiasedRNG[321])|((m[600]&~m[1313]&~m[1315]&m[1316]&~m[1317])|(~m[600]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[600]&~m[1313]&~m[1315]&~m[1316]&m[1317])|(m[600]&m[1313]&~m[1315]&~m[1316]&m[1317])|(m[600]&~m[1313]&m[1315]&~m[1316]&m[1317])|(~m[600]&~m[1313]&~m[1315]&m[1316]&m[1317])|(m[600]&~m[1313]&~m[1315]&m[1316]&m[1317])|(~m[600]&m[1313]&~m[1315]&m[1316]&m[1317])|(m[600]&m[1313]&~m[1315]&m[1316]&m[1317])|(~m[600]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[600]&~m[1313]&m[1315]&m[1316]&m[1317])|(m[600]&m[1313]&m[1315]&m[1316]&m[1317]));
    m[1319] = (((m[613]&~m[1318]&~m[1320]&~m[1321]&~m[1322])|(~m[613]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(m[613]&m[1318]&~m[1320]&m[1321]&~m[1322])|(m[613]&~m[1318]&m[1320]&m[1321]&~m[1322])|(~m[613]&m[1318]&~m[1320]&~m[1321]&m[1322])|(~m[613]&~m[1318]&m[1320]&~m[1321]&m[1322])|(m[613]&m[1318]&m[1320]&~m[1321]&m[1322])|(~m[613]&m[1318]&m[1320]&m[1321]&m[1322]))&UnbiasedRNG[322])|((m[613]&~m[1318]&~m[1320]&m[1321]&~m[1322])|(~m[613]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[613]&~m[1318]&~m[1320]&~m[1321]&m[1322])|(m[613]&m[1318]&~m[1320]&~m[1321]&m[1322])|(m[613]&~m[1318]&m[1320]&~m[1321]&m[1322])|(~m[613]&~m[1318]&~m[1320]&m[1321]&m[1322])|(m[613]&~m[1318]&~m[1320]&m[1321]&m[1322])|(~m[613]&m[1318]&~m[1320]&m[1321]&m[1322])|(m[613]&m[1318]&~m[1320]&m[1321]&m[1322])|(~m[613]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[613]&~m[1318]&m[1320]&m[1321]&m[1322])|(m[613]&m[1318]&m[1320]&m[1321]&m[1322]));
    m[1324] = (((m[626]&~m[1323]&~m[1325]&~m[1326]&~m[1327])|(~m[626]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(m[626]&m[1323]&~m[1325]&m[1326]&~m[1327])|(m[626]&~m[1323]&m[1325]&m[1326]&~m[1327])|(~m[626]&m[1323]&~m[1325]&~m[1326]&m[1327])|(~m[626]&~m[1323]&m[1325]&~m[1326]&m[1327])|(m[626]&m[1323]&m[1325]&~m[1326]&m[1327])|(~m[626]&m[1323]&m[1325]&m[1326]&m[1327]))&UnbiasedRNG[323])|((m[626]&~m[1323]&~m[1325]&m[1326]&~m[1327])|(~m[626]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[626]&~m[1323]&~m[1325]&~m[1326]&m[1327])|(m[626]&m[1323]&~m[1325]&~m[1326]&m[1327])|(m[626]&~m[1323]&m[1325]&~m[1326]&m[1327])|(~m[626]&~m[1323]&~m[1325]&m[1326]&m[1327])|(m[626]&~m[1323]&~m[1325]&m[1326]&m[1327])|(~m[626]&m[1323]&~m[1325]&m[1326]&m[1327])|(m[626]&m[1323]&~m[1325]&m[1326]&m[1327])|(~m[626]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[626]&~m[1323]&m[1325]&m[1326]&m[1327])|(m[626]&m[1323]&m[1325]&m[1326]&m[1327]));
    m[1329] = (((m[639]&~m[1328]&~m[1330]&~m[1331]&~m[1332])|(~m[639]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(m[639]&m[1328]&~m[1330]&m[1331]&~m[1332])|(m[639]&~m[1328]&m[1330]&m[1331]&~m[1332])|(~m[639]&m[1328]&~m[1330]&~m[1331]&m[1332])|(~m[639]&~m[1328]&m[1330]&~m[1331]&m[1332])|(m[639]&m[1328]&m[1330]&~m[1331]&m[1332])|(~m[639]&m[1328]&m[1330]&m[1331]&m[1332]))&UnbiasedRNG[324])|((m[639]&~m[1328]&~m[1330]&m[1331]&~m[1332])|(~m[639]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[639]&~m[1328]&~m[1330]&~m[1331]&m[1332])|(m[639]&m[1328]&~m[1330]&~m[1331]&m[1332])|(m[639]&~m[1328]&m[1330]&~m[1331]&m[1332])|(~m[639]&~m[1328]&~m[1330]&m[1331]&m[1332])|(m[639]&~m[1328]&~m[1330]&m[1331]&m[1332])|(~m[639]&m[1328]&~m[1330]&m[1331]&m[1332])|(m[639]&m[1328]&~m[1330]&m[1331]&m[1332])|(~m[639]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[639]&~m[1328]&m[1330]&m[1331]&m[1332])|(m[639]&m[1328]&m[1330]&m[1331]&m[1332]));
    m[1334] = (((m[652]&~m[1333]&~m[1335]&~m[1336]&~m[1337])|(~m[652]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(m[652]&m[1333]&~m[1335]&m[1336]&~m[1337])|(m[652]&~m[1333]&m[1335]&m[1336]&~m[1337])|(~m[652]&m[1333]&~m[1335]&~m[1336]&m[1337])|(~m[652]&~m[1333]&m[1335]&~m[1336]&m[1337])|(m[652]&m[1333]&m[1335]&~m[1336]&m[1337])|(~m[652]&m[1333]&m[1335]&m[1336]&m[1337]))&UnbiasedRNG[325])|((m[652]&~m[1333]&~m[1335]&m[1336]&~m[1337])|(~m[652]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[652]&~m[1333]&~m[1335]&~m[1336]&m[1337])|(m[652]&m[1333]&~m[1335]&~m[1336]&m[1337])|(m[652]&~m[1333]&m[1335]&~m[1336]&m[1337])|(~m[652]&~m[1333]&~m[1335]&m[1336]&m[1337])|(m[652]&~m[1333]&~m[1335]&m[1336]&m[1337])|(~m[652]&m[1333]&~m[1335]&m[1336]&m[1337])|(m[652]&m[1333]&~m[1335]&m[1336]&m[1337])|(~m[652]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[652]&~m[1333]&m[1335]&m[1336]&m[1337])|(m[652]&m[1333]&m[1335]&m[1336]&m[1337]));
    m[1339] = (((m[665]&~m[1338]&~m[1340]&~m[1341]&~m[1342])|(~m[665]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(m[665]&m[1338]&~m[1340]&m[1341]&~m[1342])|(m[665]&~m[1338]&m[1340]&m[1341]&~m[1342])|(~m[665]&m[1338]&~m[1340]&~m[1341]&m[1342])|(~m[665]&~m[1338]&m[1340]&~m[1341]&m[1342])|(m[665]&m[1338]&m[1340]&~m[1341]&m[1342])|(~m[665]&m[1338]&m[1340]&m[1341]&m[1342]))&UnbiasedRNG[326])|((m[665]&~m[1338]&~m[1340]&m[1341]&~m[1342])|(~m[665]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[665]&~m[1338]&~m[1340]&~m[1341]&m[1342])|(m[665]&m[1338]&~m[1340]&~m[1341]&m[1342])|(m[665]&~m[1338]&m[1340]&~m[1341]&m[1342])|(~m[665]&~m[1338]&~m[1340]&m[1341]&m[1342])|(m[665]&~m[1338]&~m[1340]&m[1341]&m[1342])|(~m[665]&m[1338]&~m[1340]&m[1341]&m[1342])|(m[665]&m[1338]&~m[1340]&m[1341]&m[1342])|(~m[665]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[665]&~m[1338]&m[1340]&m[1341]&m[1342])|(m[665]&m[1338]&m[1340]&m[1341]&m[1342]));
    m[1344] = (((m[678]&~m[1343]&~m[1345]&~m[1346]&~m[1347])|(~m[678]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(m[678]&m[1343]&~m[1345]&m[1346]&~m[1347])|(m[678]&~m[1343]&m[1345]&m[1346]&~m[1347])|(~m[678]&m[1343]&~m[1345]&~m[1346]&m[1347])|(~m[678]&~m[1343]&m[1345]&~m[1346]&m[1347])|(m[678]&m[1343]&m[1345]&~m[1346]&m[1347])|(~m[678]&m[1343]&m[1345]&m[1346]&m[1347]))&UnbiasedRNG[327])|((m[678]&~m[1343]&~m[1345]&m[1346]&~m[1347])|(~m[678]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[678]&~m[1343]&~m[1345]&~m[1346]&m[1347])|(m[678]&m[1343]&~m[1345]&~m[1346]&m[1347])|(m[678]&~m[1343]&m[1345]&~m[1346]&m[1347])|(~m[678]&~m[1343]&~m[1345]&m[1346]&m[1347])|(m[678]&~m[1343]&~m[1345]&m[1346]&m[1347])|(~m[678]&m[1343]&~m[1345]&m[1346]&m[1347])|(m[678]&m[1343]&~m[1345]&m[1346]&m[1347])|(~m[678]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[678]&~m[1343]&m[1345]&m[1346]&m[1347])|(m[678]&m[1343]&m[1345]&m[1346]&m[1347]));
    m[1349] = (((m[691]&~m[1348]&~m[1350]&~m[1351]&~m[1352])|(~m[691]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(m[691]&m[1348]&~m[1350]&m[1351]&~m[1352])|(m[691]&~m[1348]&m[1350]&m[1351]&~m[1352])|(~m[691]&m[1348]&~m[1350]&~m[1351]&m[1352])|(~m[691]&~m[1348]&m[1350]&~m[1351]&m[1352])|(m[691]&m[1348]&m[1350]&~m[1351]&m[1352])|(~m[691]&m[1348]&m[1350]&m[1351]&m[1352]))&UnbiasedRNG[328])|((m[691]&~m[1348]&~m[1350]&m[1351]&~m[1352])|(~m[691]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[691]&~m[1348]&~m[1350]&~m[1351]&m[1352])|(m[691]&m[1348]&~m[1350]&~m[1351]&m[1352])|(m[691]&~m[1348]&m[1350]&~m[1351]&m[1352])|(~m[691]&~m[1348]&~m[1350]&m[1351]&m[1352])|(m[691]&~m[1348]&~m[1350]&m[1351]&m[1352])|(~m[691]&m[1348]&~m[1350]&m[1351]&m[1352])|(m[691]&m[1348]&~m[1350]&m[1351]&m[1352])|(~m[691]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[691]&~m[1348]&m[1350]&m[1351]&m[1352])|(m[691]&m[1348]&m[1350]&m[1351]&m[1352]));
    m[1354] = (((m[704]&~m[1353]&~m[1355]&~m[1356]&~m[1357])|(~m[704]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(m[704]&m[1353]&~m[1355]&m[1356]&~m[1357])|(m[704]&~m[1353]&m[1355]&m[1356]&~m[1357])|(~m[704]&m[1353]&~m[1355]&~m[1356]&m[1357])|(~m[704]&~m[1353]&m[1355]&~m[1356]&m[1357])|(m[704]&m[1353]&m[1355]&~m[1356]&m[1357])|(~m[704]&m[1353]&m[1355]&m[1356]&m[1357]))&UnbiasedRNG[329])|((m[704]&~m[1353]&~m[1355]&m[1356]&~m[1357])|(~m[704]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[704]&~m[1353]&~m[1355]&~m[1356]&m[1357])|(m[704]&m[1353]&~m[1355]&~m[1356]&m[1357])|(m[704]&~m[1353]&m[1355]&~m[1356]&m[1357])|(~m[704]&~m[1353]&~m[1355]&m[1356]&m[1357])|(m[704]&~m[1353]&~m[1355]&m[1356]&m[1357])|(~m[704]&m[1353]&~m[1355]&m[1356]&m[1357])|(m[704]&m[1353]&~m[1355]&m[1356]&m[1357])|(~m[704]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[704]&~m[1353]&m[1355]&m[1356]&m[1357])|(m[704]&m[1353]&m[1355]&m[1356]&m[1357]));
    m[1359] = (((m[717]&~m[1358]&~m[1360]&~m[1361]&~m[1362])|(~m[717]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(m[717]&m[1358]&~m[1360]&m[1361]&~m[1362])|(m[717]&~m[1358]&m[1360]&m[1361]&~m[1362])|(~m[717]&m[1358]&~m[1360]&~m[1361]&m[1362])|(~m[717]&~m[1358]&m[1360]&~m[1361]&m[1362])|(m[717]&m[1358]&m[1360]&~m[1361]&m[1362])|(~m[717]&m[1358]&m[1360]&m[1361]&m[1362]))&UnbiasedRNG[330])|((m[717]&~m[1358]&~m[1360]&m[1361]&~m[1362])|(~m[717]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[717]&~m[1358]&~m[1360]&~m[1361]&m[1362])|(m[717]&m[1358]&~m[1360]&~m[1361]&m[1362])|(m[717]&~m[1358]&m[1360]&~m[1361]&m[1362])|(~m[717]&~m[1358]&~m[1360]&m[1361]&m[1362])|(m[717]&~m[1358]&~m[1360]&m[1361]&m[1362])|(~m[717]&m[1358]&~m[1360]&m[1361]&m[1362])|(m[717]&m[1358]&~m[1360]&m[1361]&m[1362])|(~m[717]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[717]&~m[1358]&m[1360]&m[1361]&m[1362])|(m[717]&m[1358]&m[1360]&m[1361]&m[1362]));
    m[1364] = (((m[601]&~m[1363]&~m[1365]&~m[1366]&~m[1367])|(~m[601]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(m[601]&m[1363]&~m[1365]&m[1366]&~m[1367])|(m[601]&~m[1363]&m[1365]&m[1366]&~m[1367])|(~m[601]&m[1363]&~m[1365]&~m[1366]&m[1367])|(~m[601]&~m[1363]&m[1365]&~m[1366]&m[1367])|(m[601]&m[1363]&m[1365]&~m[1366]&m[1367])|(~m[601]&m[1363]&m[1365]&m[1366]&m[1367]))&UnbiasedRNG[331])|((m[601]&~m[1363]&~m[1365]&m[1366]&~m[1367])|(~m[601]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[601]&~m[1363]&~m[1365]&~m[1366]&m[1367])|(m[601]&m[1363]&~m[1365]&~m[1366]&m[1367])|(m[601]&~m[1363]&m[1365]&~m[1366]&m[1367])|(~m[601]&~m[1363]&~m[1365]&m[1366]&m[1367])|(m[601]&~m[1363]&~m[1365]&m[1366]&m[1367])|(~m[601]&m[1363]&~m[1365]&m[1366]&m[1367])|(m[601]&m[1363]&~m[1365]&m[1366]&m[1367])|(~m[601]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[601]&~m[1363]&m[1365]&m[1366]&m[1367])|(m[601]&m[1363]&m[1365]&m[1366]&m[1367]));
    m[1369] = (((m[614]&~m[1368]&~m[1370]&~m[1371]&~m[1372])|(~m[614]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(m[614]&m[1368]&~m[1370]&m[1371]&~m[1372])|(m[614]&~m[1368]&m[1370]&m[1371]&~m[1372])|(~m[614]&m[1368]&~m[1370]&~m[1371]&m[1372])|(~m[614]&~m[1368]&m[1370]&~m[1371]&m[1372])|(m[614]&m[1368]&m[1370]&~m[1371]&m[1372])|(~m[614]&m[1368]&m[1370]&m[1371]&m[1372]))&UnbiasedRNG[332])|((m[614]&~m[1368]&~m[1370]&m[1371]&~m[1372])|(~m[614]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[614]&~m[1368]&~m[1370]&~m[1371]&m[1372])|(m[614]&m[1368]&~m[1370]&~m[1371]&m[1372])|(m[614]&~m[1368]&m[1370]&~m[1371]&m[1372])|(~m[614]&~m[1368]&~m[1370]&m[1371]&m[1372])|(m[614]&~m[1368]&~m[1370]&m[1371]&m[1372])|(~m[614]&m[1368]&~m[1370]&m[1371]&m[1372])|(m[614]&m[1368]&~m[1370]&m[1371]&m[1372])|(~m[614]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[614]&~m[1368]&m[1370]&m[1371]&m[1372])|(m[614]&m[1368]&m[1370]&m[1371]&m[1372]));
    m[1374] = (((m[627]&~m[1373]&~m[1375]&~m[1376]&~m[1377])|(~m[627]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(m[627]&m[1373]&~m[1375]&m[1376]&~m[1377])|(m[627]&~m[1373]&m[1375]&m[1376]&~m[1377])|(~m[627]&m[1373]&~m[1375]&~m[1376]&m[1377])|(~m[627]&~m[1373]&m[1375]&~m[1376]&m[1377])|(m[627]&m[1373]&m[1375]&~m[1376]&m[1377])|(~m[627]&m[1373]&m[1375]&m[1376]&m[1377]))&UnbiasedRNG[333])|((m[627]&~m[1373]&~m[1375]&m[1376]&~m[1377])|(~m[627]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[627]&~m[1373]&~m[1375]&~m[1376]&m[1377])|(m[627]&m[1373]&~m[1375]&~m[1376]&m[1377])|(m[627]&~m[1373]&m[1375]&~m[1376]&m[1377])|(~m[627]&~m[1373]&~m[1375]&m[1376]&m[1377])|(m[627]&~m[1373]&~m[1375]&m[1376]&m[1377])|(~m[627]&m[1373]&~m[1375]&m[1376]&m[1377])|(m[627]&m[1373]&~m[1375]&m[1376]&m[1377])|(~m[627]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[627]&~m[1373]&m[1375]&m[1376]&m[1377])|(m[627]&m[1373]&m[1375]&m[1376]&m[1377]));
    m[1379] = (((m[640]&~m[1378]&~m[1380]&~m[1381]&~m[1382])|(~m[640]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(m[640]&m[1378]&~m[1380]&m[1381]&~m[1382])|(m[640]&~m[1378]&m[1380]&m[1381]&~m[1382])|(~m[640]&m[1378]&~m[1380]&~m[1381]&m[1382])|(~m[640]&~m[1378]&m[1380]&~m[1381]&m[1382])|(m[640]&m[1378]&m[1380]&~m[1381]&m[1382])|(~m[640]&m[1378]&m[1380]&m[1381]&m[1382]))&UnbiasedRNG[334])|((m[640]&~m[1378]&~m[1380]&m[1381]&~m[1382])|(~m[640]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[640]&~m[1378]&~m[1380]&~m[1381]&m[1382])|(m[640]&m[1378]&~m[1380]&~m[1381]&m[1382])|(m[640]&~m[1378]&m[1380]&~m[1381]&m[1382])|(~m[640]&~m[1378]&~m[1380]&m[1381]&m[1382])|(m[640]&~m[1378]&~m[1380]&m[1381]&m[1382])|(~m[640]&m[1378]&~m[1380]&m[1381]&m[1382])|(m[640]&m[1378]&~m[1380]&m[1381]&m[1382])|(~m[640]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[640]&~m[1378]&m[1380]&m[1381]&m[1382])|(m[640]&m[1378]&m[1380]&m[1381]&m[1382]));
    m[1384] = (((m[653]&~m[1383]&~m[1385]&~m[1386]&~m[1387])|(~m[653]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(m[653]&m[1383]&~m[1385]&m[1386]&~m[1387])|(m[653]&~m[1383]&m[1385]&m[1386]&~m[1387])|(~m[653]&m[1383]&~m[1385]&~m[1386]&m[1387])|(~m[653]&~m[1383]&m[1385]&~m[1386]&m[1387])|(m[653]&m[1383]&m[1385]&~m[1386]&m[1387])|(~m[653]&m[1383]&m[1385]&m[1386]&m[1387]))&UnbiasedRNG[335])|((m[653]&~m[1383]&~m[1385]&m[1386]&~m[1387])|(~m[653]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[653]&~m[1383]&~m[1385]&~m[1386]&m[1387])|(m[653]&m[1383]&~m[1385]&~m[1386]&m[1387])|(m[653]&~m[1383]&m[1385]&~m[1386]&m[1387])|(~m[653]&~m[1383]&~m[1385]&m[1386]&m[1387])|(m[653]&~m[1383]&~m[1385]&m[1386]&m[1387])|(~m[653]&m[1383]&~m[1385]&m[1386]&m[1387])|(m[653]&m[1383]&~m[1385]&m[1386]&m[1387])|(~m[653]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[653]&~m[1383]&m[1385]&m[1386]&m[1387])|(m[653]&m[1383]&m[1385]&m[1386]&m[1387]));
    m[1389] = (((m[666]&~m[1388]&~m[1390]&~m[1391]&~m[1392])|(~m[666]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(m[666]&m[1388]&~m[1390]&m[1391]&~m[1392])|(m[666]&~m[1388]&m[1390]&m[1391]&~m[1392])|(~m[666]&m[1388]&~m[1390]&~m[1391]&m[1392])|(~m[666]&~m[1388]&m[1390]&~m[1391]&m[1392])|(m[666]&m[1388]&m[1390]&~m[1391]&m[1392])|(~m[666]&m[1388]&m[1390]&m[1391]&m[1392]))&UnbiasedRNG[336])|((m[666]&~m[1388]&~m[1390]&m[1391]&~m[1392])|(~m[666]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[666]&~m[1388]&~m[1390]&~m[1391]&m[1392])|(m[666]&m[1388]&~m[1390]&~m[1391]&m[1392])|(m[666]&~m[1388]&m[1390]&~m[1391]&m[1392])|(~m[666]&~m[1388]&~m[1390]&m[1391]&m[1392])|(m[666]&~m[1388]&~m[1390]&m[1391]&m[1392])|(~m[666]&m[1388]&~m[1390]&m[1391]&m[1392])|(m[666]&m[1388]&~m[1390]&m[1391]&m[1392])|(~m[666]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[666]&~m[1388]&m[1390]&m[1391]&m[1392])|(m[666]&m[1388]&m[1390]&m[1391]&m[1392]));
    m[1394] = (((m[679]&~m[1393]&~m[1395]&~m[1396]&~m[1397])|(~m[679]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(m[679]&m[1393]&~m[1395]&m[1396]&~m[1397])|(m[679]&~m[1393]&m[1395]&m[1396]&~m[1397])|(~m[679]&m[1393]&~m[1395]&~m[1396]&m[1397])|(~m[679]&~m[1393]&m[1395]&~m[1396]&m[1397])|(m[679]&m[1393]&m[1395]&~m[1396]&m[1397])|(~m[679]&m[1393]&m[1395]&m[1396]&m[1397]))&UnbiasedRNG[337])|((m[679]&~m[1393]&~m[1395]&m[1396]&~m[1397])|(~m[679]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[679]&~m[1393]&~m[1395]&~m[1396]&m[1397])|(m[679]&m[1393]&~m[1395]&~m[1396]&m[1397])|(m[679]&~m[1393]&m[1395]&~m[1396]&m[1397])|(~m[679]&~m[1393]&~m[1395]&m[1396]&m[1397])|(m[679]&~m[1393]&~m[1395]&m[1396]&m[1397])|(~m[679]&m[1393]&~m[1395]&m[1396]&m[1397])|(m[679]&m[1393]&~m[1395]&m[1396]&m[1397])|(~m[679]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[679]&~m[1393]&m[1395]&m[1396]&m[1397])|(m[679]&m[1393]&m[1395]&m[1396]&m[1397]));
    m[1399] = (((m[692]&~m[1398]&~m[1400]&~m[1401]&~m[1402])|(~m[692]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(m[692]&m[1398]&~m[1400]&m[1401]&~m[1402])|(m[692]&~m[1398]&m[1400]&m[1401]&~m[1402])|(~m[692]&m[1398]&~m[1400]&~m[1401]&m[1402])|(~m[692]&~m[1398]&m[1400]&~m[1401]&m[1402])|(m[692]&m[1398]&m[1400]&~m[1401]&m[1402])|(~m[692]&m[1398]&m[1400]&m[1401]&m[1402]))&UnbiasedRNG[338])|((m[692]&~m[1398]&~m[1400]&m[1401]&~m[1402])|(~m[692]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[692]&~m[1398]&~m[1400]&~m[1401]&m[1402])|(m[692]&m[1398]&~m[1400]&~m[1401]&m[1402])|(m[692]&~m[1398]&m[1400]&~m[1401]&m[1402])|(~m[692]&~m[1398]&~m[1400]&m[1401]&m[1402])|(m[692]&~m[1398]&~m[1400]&m[1401]&m[1402])|(~m[692]&m[1398]&~m[1400]&m[1401]&m[1402])|(m[692]&m[1398]&~m[1400]&m[1401]&m[1402])|(~m[692]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[692]&~m[1398]&m[1400]&m[1401]&m[1402])|(m[692]&m[1398]&m[1400]&m[1401]&m[1402]));
    m[1404] = (((m[705]&~m[1403]&~m[1405]&~m[1406]&~m[1407])|(~m[705]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(m[705]&m[1403]&~m[1405]&m[1406]&~m[1407])|(m[705]&~m[1403]&m[1405]&m[1406]&~m[1407])|(~m[705]&m[1403]&~m[1405]&~m[1406]&m[1407])|(~m[705]&~m[1403]&m[1405]&~m[1406]&m[1407])|(m[705]&m[1403]&m[1405]&~m[1406]&m[1407])|(~m[705]&m[1403]&m[1405]&m[1406]&m[1407]))&UnbiasedRNG[339])|((m[705]&~m[1403]&~m[1405]&m[1406]&~m[1407])|(~m[705]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[705]&~m[1403]&~m[1405]&~m[1406]&m[1407])|(m[705]&m[1403]&~m[1405]&~m[1406]&m[1407])|(m[705]&~m[1403]&m[1405]&~m[1406]&m[1407])|(~m[705]&~m[1403]&~m[1405]&m[1406]&m[1407])|(m[705]&~m[1403]&~m[1405]&m[1406]&m[1407])|(~m[705]&m[1403]&~m[1405]&m[1406]&m[1407])|(m[705]&m[1403]&~m[1405]&m[1406]&m[1407])|(~m[705]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[705]&~m[1403]&m[1405]&m[1406]&m[1407])|(m[705]&m[1403]&m[1405]&m[1406]&m[1407]));
    m[1409] = (((m[718]&~m[1408]&~m[1410]&~m[1411]&~m[1412])|(~m[718]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(m[718]&m[1408]&~m[1410]&m[1411]&~m[1412])|(m[718]&~m[1408]&m[1410]&m[1411]&~m[1412])|(~m[718]&m[1408]&~m[1410]&~m[1411]&m[1412])|(~m[718]&~m[1408]&m[1410]&~m[1411]&m[1412])|(m[718]&m[1408]&m[1410]&~m[1411]&m[1412])|(~m[718]&m[1408]&m[1410]&m[1411]&m[1412]))&UnbiasedRNG[340])|((m[718]&~m[1408]&~m[1410]&m[1411]&~m[1412])|(~m[718]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[718]&~m[1408]&~m[1410]&~m[1411]&m[1412])|(m[718]&m[1408]&~m[1410]&~m[1411]&m[1412])|(m[718]&~m[1408]&m[1410]&~m[1411]&m[1412])|(~m[718]&~m[1408]&~m[1410]&m[1411]&m[1412])|(m[718]&~m[1408]&~m[1410]&m[1411]&m[1412])|(~m[718]&m[1408]&~m[1410]&m[1411]&m[1412])|(m[718]&m[1408]&~m[1410]&m[1411]&m[1412])|(~m[718]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[718]&~m[1408]&m[1410]&m[1411]&m[1412])|(m[718]&m[1408]&m[1410]&m[1411]&m[1412]));
    m[1414] = (((m[615]&~m[1413]&~m[1415]&~m[1416]&~m[1417])|(~m[615]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(m[615]&m[1413]&~m[1415]&m[1416]&~m[1417])|(m[615]&~m[1413]&m[1415]&m[1416]&~m[1417])|(~m[615]&m[1413]&~m[1415]&~m[1416]&m[1417])|(~m[615]&~m[1413]&m[1415]&~m[1416]&m[1417])|(m[615]&m[1413]&m[1415]&~m[1416]&m[1417])|(~m[615]&m[1413]&m[1415]&m[1416]&m[1417]))&UnbiasedRNG[341])|((m[615]&~m[1413]&~m[1415]&m[1416]&~m[1417])|(~m[615]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[615]&~m[1413]&~m[1415]&~m[1416]&m[1417])|(m[615]&m[1413]&~m[1415]&~m[1416]&m[1417])|(m[615]&~m[1413]&m[1415]&~m[1416]&m[1417])|(~m[615]&~m[1413]&~m[1415]&m[1416]&m[1417])|(m[615]&~m[1413]&~m[1415]&m[1416]&m[1417])|(~m[615]&m[1413]&~m[1415]&m[1416]&m[1417])|(m[615]&m[1413]&~m[1415]&m[1416]&m[1417])|(~m[615]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[615]&~m[1413]&m[1415]&m[1416]&m[1417])|(m[615]&m[1413]&m[1415]&m[1416]&m[1417]));
    m[1419] = (((m[628]&~m[1418]&~m[1420]&~m[1421]&~m[1422])|(~m[628]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(m[628]&m[1418]&~m[1420]&m[1421]&~m[1422])|(m[628]&~m[1418]&m[1420]&m[1421]&~m[1422])|(~m[628]&m[1418]&~m[1420]&~m[1421]&m[1422])|(~m[628]&~m[1418]&m[1420]&~m[1421]&m[1422])|(m[628]&m[1418]&m[1420]&~m[1421]&m[1422])|(~m[628]&m[1418]&m[1420]&m[1421]&m[1422]))&UnbiasedRNG[342])|((m[628]&~m[1418]&~m[1420]&m[1421]&~m[1422])|(~m[628]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[628]&~m[1418]&~m[1420]&~m[1421]&m[1422])|(m[628]&m[1418]&~m[1420]&~m[1421]&m[1422])|(m[628]&~m[1418]&m[1420]&~m[1421]&m[1422])|(~m[628]&~m[1418]&~m[1420]&m[1421]&m[1422])|(m[628]&~m[1418]&~m[1420]&m[1421]&m[1422])|(~m[628]&m[1418]&~m[1420]&m[1421]&m[1422])|(m[628]&m[1418]&~m[1420]&m[1421]&m[1422])|(~m[628]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[628]&~m[1418]&m[1420]&m[1421]&m[1422])|(m[628]&m[1418]&m[1420]&m[1421]&m[1422]));
    m[1424] = (((m[641]&~m[1423]&~m[1425]&~m[1426]&~m[1427])|(~m[641]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(m[641]&m[1423]&~m[1425]&m[1426]&~m[1427])|(m[641]&~m[1423]&m[1425]&m[1426]&~m[1427])|(~m[641]&m[1423]&~m[1425]&~m[1426]&m[1427])|(~m[641]&~m[1423]&m[1425]&~m[1426]&m[1427])|(m[641]&m[1423]&m[1425]&~m[1426]&m[1427])|(~m[641]&m[1423]&m[1425]&m[1426]&m[1427]))&UnbiasedRNG[343])|((m[641]&~m[1423]&~m[1425]&m[1426]&~m[1427])|(~m[641]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[641]&~m[1423]&~m[1425]&~m[1426]&m[1427])|(m[641]&m[1423]&~m[1425]&~m[1426]&m[1427])|(m[641]&~m[1423]&m[1425]&~m[1426]&m[1427])|(~m[641]&~m[1423]&~m[1425]&m[1426]&m[1427])|(m[641]&~m[1423]&~m[1425]&m[1426]&m[1427])|(~m[641]&m[1423]&~m[1425]&m[1426]&m[1427])|(m[641]&m[1423]&~m[1425]&m[1426]&m[1427])|(~m[641]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[641]&~m[1423]&m[1425]&m[1426]&m[1427])|(m[641]&m[1423]&m[1425]&m[1426]&m[1427]));
    m[1429] = (((m[654]&~m[1428]&~m[1430]&~m[1431]&~m[1432])|(~m[654]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(m[654]&m[1428]&~m[1430]&m[1431]&~m[1432])|(m[654]&~m[1428]&m[1430]&m[1431]&~m[1432])|(~m[654]&m[1428]&~m[1430]&~m[1431]&m[1432])|(~m[654]&~m[1428]&m[1430]&~m[1431]&m[1432])|(m[654]&m[1428]&m[1430]&~m[1431]&m[1432])|(~m[654]&m[1428]&m[1430]&m[1431]&m[1432]))&UnbiasedRNG[344])|((m[654]&~m[1428]&~m[1430]&m[1431]&~m[1432])|(~m[654]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[654]&~m[1428]&~m[1430]&~m[1431]&m[1432])|(m[654]&m[1428]&~m[1430]&~m[1431]&m[1432])|(m[654]&~m[1428]&m[1430]&~m[1431]&m[1432])|(~m[654]&~m[1428]&~m[1430]&m[1431]&m[1432])|(m[654]&~m[1428]&~m[1430]&m[1431]&m[1432])|(~m[654]&m[1428]&~m[1430]&m[1431]&m[1432])|(m[654]&m[1428]&~m[1430]&m[1431]&m[1432])|(~m[654]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[654]&~m[1428]&m[1430]&m[1431]&m[1432])|(m[654]&m[1428]&m[1430]&m[1431]&m[1432]));
    m[1434] = (((m[667]&~m[1433]&~m[1435]&~m[1436]&~m[1437])|(~m[667]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(m[667]&m[1433]&~m[1435]&m[1436]&~m[1437])|(m[667]&~m[1433]&m[1435]&m[1436]&~m[1437])|(~m[667]&m[1433]&~m[1435]&~m[1436]&m[1437])|(~m[667]&~m[1433]&m[1435]&~m[1436]&m[1437])|(m[667]&m[1433]&m[1435]&~m[1436]&m[1437])|(~m[667]&m[1433]&m[1435]&m[1436]&m[1437]))&UnbiasedRNG[345])|((m[667]&~m[1433]&~m[1435]&m[1436]&~m[1437])|(~m[667]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[667]&~m[1433]&~m[1435]&~m[1436]&m[1437])|(m[667]&m[1433]&~m[1435]&~m[1436]&m[1437])|(m[667]&~m[1433]&m[1435]&~m[1436]&m[1437])|(~m[667]&~m[1433]&~m[1435]&m[1436]&m[1437])|(m[667]&~m[1433]&~m[1435]&m[1436]&m[1437])|(~m[667]&m[1433]&~m[1435]&m[1436]&m[1437])|(m[667]&m[1433]&~m[1435]&m[1436]&m[1437])|(~m[667]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[667]&~m[1433]&m[1435]&m[1436]&m[1437])|(m[667]&m[1433]&m[1435]&m[1436]&m[1437]));
    m[1439] = (((m[680]&~m[1438]&~m[1440]&~m[1441]&~m[1442])|(~m[680]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(m[680]&m[1438]&~m[1440]&m[1441]&~m[1442])|(m[680]&~m[1438]&m[1440]&m[1441]&~m[1442])|(~m[680]&m[1438]&~m[1440]&~m[1441]&m[1442])|(~m[680]&~m[1438]&m[1440]&~m[1441]&m[1442])|(m[680]&m[1438]&m[1440]&~m[1441]&m[1442])|(~m[680]&m[1438]&m[1440]&m[1441]&m[1442]))&UnbiasedRNG[346])|((m[680]&~m[1438]&~m[1440]&m[1441]&~m[1442])|(~m[680]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[680]&~m[1438]&~m[1440]&~m[1441]&m[1442])|(m[680]&m[1438]&~m[1440]&~m[1441]&m[1442])|(m[680]&~m[1438]&m[1440]&~m[1441]&m[1442])|(~m[680]&~m[1438]&~m[1440]&m[1441]&m[1442])|(m[680]&~m[1438]&~m[1440]&m[1441]&m[1442])|(~m[680]&m[1438]&~m[1440]&m[1441]&m[1442])|(m[680]&m[1438]&~m[1440]&m[1441]&m[1442])|(~m[680]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[680]&~m[1438]&m[1440]&m[1441]&m[1442])|(m[680]&m[1438]&m[1440]&m[1441]&m[1442]));
    m[1444] = (((m[693]&~m[1443]&~m[1445]&~m[1446]&~m[1447])|(~m[693]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(m[693]&m[1443]&~m[1445]&m[1446]&~m[1447])|(m[693]&~m[1443]&m[1445]&m[1446]&~m[1447])|(~m[693]&m[1443]&~m[1445]&~m[1446]&m[1447])|(~m[693]&~m[1443]&m[1445]&~m[1446]&m[1447])|(m[693]&m[1443]&m[1445]&~m[1446]&m[1447])|(~m[693]&m[1443]&m[1445]&m[1446]&m[1447]))&UnbiasedRNG[347])|((m[693]&~m[1443]&~m[1445]&m[1446]&~m[1447])|(~m[693]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[693]&~m[1443]&~m[1445]&~m[1446]&m[1447])|(m[693]&m[1443]&~m[1445]&~m[1446]&m[1447])|(m[693]&~m[1443]&m[1445]&~m[1446]&m[1447])|(~m[693]&~m[1443]&~m[1445]&m[1446]&m[1447])|(m[693]&~m[1443]&~m[1445]&m[1446]&m[1447])|(~m[693]&m[1443]&~m[1445]&m[1446]&m[1447])|(m[693]&m[1443]&~m[1445]&m[1446]&m[1447])|(~m[693]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[693]&~m[1443]&m[1445]&m[1446]&m[1447])|(m[693]&m[1443]&m[1445]&m[1446]&m[1447]));
    m[1449] = (((m[706]&~m[1448]&~m[1450]&~m[1451]&~m[1452])|(~m[706]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(m[706]&m[1448]&~m[1450]&m[1451]&~m[1452])|(m[706]&~m[1448]&m[1450]&m[1451]&~m[1452])|(~m[706]&m[1448]&~m[1450]&~m[1451]&m[1452])|(~m[706]&~m[1448]&m[1450]&~m[1451]&m[1452])|(m[706]&m[1448]&m[1450]&~m[1451]&m[1452])|(~m[706]&m[1448]&m[1450]&m[1451]&m[1452]))&UnbiasedRNG[348])|((m[706]&~m[1448]&~m[1450]&m[1451]&~m[1452])|(~m[706]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[706]&~m[1448]&~m[1450]&~m[1451]&m[1452])|(m[706]&m[1448]&~m[1450]&~m[1451]&m[1452])|(m[706]&~m[1448]&m[1450]&~m[1451]&m[1452])|(~m[706]&~m[1448]&~m[1450]&m[1451]&m[1452])|(m[706]&~m[1448]&~m[1450]&m[1451]&m[1452])|(~m[706]&m[1448]&~m[1450]&m[1451]&m[1452])|(m[706]&m[1448]&~m[1450]&m[1451]&m[1452])|(~m[706]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[706]&~m[1448]&m[1450]&m[1451]&m[1452])|(m[706]&m[1448]&m[1450]&m[1451]&m[1452]));
    m[1454] = (((m[719]&~m[1453]&~m[1455]&~m[1456]&~m[1457])|(~m[719]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(m[719]&m[1453]&~m[1455]&m[1456]&~m[1457])|(m[719]&~m[1453]&m[1455]&m[1456]&~m[1457])|(~m[719]&m[1453]&~m[1455]&~m[1456]&m[1457])|(~m[719]&~m[1453]&m[1455]&~m[1456]&m[1457])|(m[719]&m[1453]&m[1455]&~m[1456]&m[1457])|(~m[719]&m[1453]&m[1455]&m[1456]&m[1457]))&UnbiasedRNG[349])|((m[719]&~m[1453]&~m[1455]&m[1456]&~m[1457])|(~m[719]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[719]&~m[1453]&~m[1455]&~m[1456]&m[1457])|(m[719]&m[1453]&~m[1455]&~m[1456]&m[1457])|(m[719]&~m[1453]&m[1455]&~m[1456]&m[1457])|(~m[719]&~m[1453]&~m[1455]&m[1456]&m[1457])|(m[719]&~m[1453]&~m[1455]&m[1456]&m[1457])|(~m[719]&m[1453]&~m[1455]&m[1456]&m[1457])|(m[719]&m[1453]&~m[1455]&m[1456]&m[1457])|(~m[719]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[719]&~m[1453]&m[1455]&m[1456]&m[1457])|(m[719]&m[1453]&m[1455]&m[1456]&m[1457]));
    m[1459] = (((m[629]&~m[1458]&~m[1460]&~m[1461]&~m[1462])|(~m[629]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(m[629]&m[1458]&~m[1460]&m[1461]&~m[1462])|(m[629]&~m[1458]&m[1460]&m[1461]&~m[1462])|(~m[629]&m[1458]&~m[1460]&~m[1461]&m[1462])|(~m[629]&~m[1458]&m[1460]&~m[1461]&m[1462])|(m[629]&m[1458]&m[1460]&~m[1461]&m[1462])|(~m[629]&m[1458]&m[1460]&m[1461]&m[1462]))&UnbiasedRNG[350])|((m[629]&~m[1458]&~m[1460]&m[1461]&~m[1462])|(~m[629]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[629]&~m[1458]&~m[1460]&~m[1461]&m[1462])|(m[629]&m[1458]&~m[1460]&~m[1461]&m[1462])|(m[629]&~m[1458]&m[1460]&~m[1461]&m[1462])|(~m[629]&~m[1458]&~m[1460]&m[1461]&m[1462])|(m[629]&~m[1458]&~m[1460]&m[1461]&m[1462])|(~m[629]&m[1458]&~m[1460]&m[1461]&m[1462])|(m[629]&m[1458]&~m[1460]&m[1461]&m[1462])|(~m[629]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[629]&~m[1458]&m[1460]&m[1461]&m[1462])|(m[629]&m[1458]&m[1460]&m[1461]&m[1462]));
    m[1464] = (((m[642]&~m[1463]&~m[1465]&~m[1466]&~m[1467])|(~m[642]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(m[642]&m[1463]&~m[1465]&m[1466]&~m[1467])|(m[642]&~m[1463]&m[1465]&m[1466]&~m[1467])|(~m[642]&m[1463]&~m[1465]&~m[1466]&m[1467])|(~m[642]&~m[1463]&m[1465]&~m[1466]&m[1467])|(m[642]&m[1463]&m[1465]&~m[1466]&m[1467])|(~m[642]&m[1463]&m[1465]&m[1466]&m[1467]))&UnbiasedRNG[351])|((m[642]&~m[1463]&~m[1465]&m[1466]&~m[1467])|(~m[642]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[642]&~m[1463]&~m[1465]&~m[1466]&m[1467])|(m[642]&m[1463]&~m[1465]&~m[1466]&m[1467])|(m[642]&~m[1463]&m[1465]&~m[1466]&m[1467])|(~m[642]&~m[1463]&~m[1465]&m[1466]&m[1467])|(m[642]&~m[1463]&~m[1465]&m[1466]&m[1467])|(~m[642]&m[1463]&~m[1465]&m[1466]&m[1467])|(m[642]&m[1463]&~m[1465]&m[1466]&m[1467])|(~m[642]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[642]&~m[1463]&m[1465]&m[1466]&m[1467])|(m[642]&m[1463]&m[1465]&m[1466]&m[1467]));
    m[1469] = (((m[655]&~m[1468]&~m[1470]&~m[1471]&~m[1472])|(~m[655]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(m[655]&m[1468]&~m[1470]&m[1471]&~m[1472])|(m[655]&~m[1468]&m[1470]&m[1471]&~m[1472])|(~m[655]&m[1468]&~m[1470]&~m[1471]&m[1472])|(~m[655]&~m[1468]&m[1470]&~m[1471]&m[1472])|(m[655]&m[1468]&m[1470]&~m[1471]&m[1472])|(~m[655]&m[1468]&m[1470]&m[1471]&m[1472]))&UnbiasedRNG[352])|((m[655]&~m[1468]&~m[1470]&m[1471]&~m[1472])|(~m[655]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[655]&~m[1468]&~m[1470]&~m[1471]&m[1472])|(m[655]&m[1468]&~m[1470]&~m[1471]&m[1472])|(m[655]&~m[1468]&m[1470]&~m[1471]&m[1472])|(~m[655]&~m[1468]&~m[1470]&m[1471]&m[1472])|(m[655]&~m[1468]&~m[1470]&m[1471]&m[1472])|(~m[655]&m[1468]&~m[1470]&m[1471]&m[1472])|(m[655]&m[1468]&~m[1470]&m[1471]&m[1472])|(~m[655]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[655]&~m[1468]&m[1470]&m[1471]&m[1472])|(m[655]&m[1468]&m[1470]&m[1471]&m[1472]));
    m[1474] = (((m[668]&~m[1473]&~m[1475]&~m[1476]&~m[1477])|(~m[668]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(m[668]&m[1473]&~m[1475]&m[1476]&~m[1477])|(m[668]&~m[1473]&m[1475]&m[1476]&~m[1477])|(~m[668]&m[1473]&~m[1475]&~m[1476]&m[1477])|(~m[668]&~m[1473]&m[1475]&~m[1476]&m[1477])|(m[668]&m[1473]&m[1475]&~m[1476]&m[1477])|(~m[668]&m[1473]&m[1475]&m[1476]&m[1477]))&UnbiasedRNG[353])|((m[668]&~m[1473]&~m[1475]&m[1476]&~m[1477])|(~m[668]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[668]&~m[1473]&~m[1475]&~m[1476]&m[1477])|(m[668]&m[1473]&~m[1475]&~m[1476]&m[1477])|(m[668]&~m[1473]&m[1475]&~m[1476]&m[1477])|(~m[668]&~m[1473]&~m[1475]&m[1476]&m[1477])|(m[668]&~m[1473]&~m[1475]&m[1476]&m[1477])|(~m[668]&m[1473]&~m[1475]&m[1476]&m[1477])|(m[668]&m[1473]&~m[1475]&m[1476]&m[1477])|(~m[668]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[668]&~m[1473]&m[1475]&m[1476]&m[1477])|(m[668]&m[1473]&m[1475]&m[1476]&m[1477]));
    m[1479] = (((m[681]&~m[1478]&~m[1480]&~m[1481]&~m[1482])|(~m[681]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(m[681]&m[1478]&~m[1480]&m[1481]&~m[1482])|(m[681]&~m[1478]&m[1480]&m[1481]&~m[1482])|(~m[681]&m[1478]&~m[1480]&~m[1481]&m[1482])|(~m[681]&~m[1478]&m[1480]&~m[1481]&m[1482])|(m[681]&m[1478]&m[1480]&~m[1481]&m[1482])|(~m[681]&m[1478]&m[1480]&m[1481]&m[1482]))&UnbiasedRNG[354])|((m[681]&~m[1478]&~m[1480]&m[1481]&~m[1482])|(~m[681]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[681]&~m[1478]&~m[1480]&~m[1481]&m[1482])|(m[681]&m[1478]&~m[1480]&~m[1481]&m[1482])|(m[681]&~m[1478]&m[1480]&~m[1481]&m[1482])|(~m[681]&~m[1478]&~m[1480]&m[1481]&m[1482])|(m[681]&~m[1478]&~m[1480]&m[1481]&m[1482])|(~m[681]&m[1478]&~m[1480]&m[1481]&m[1482])|(m[681]&m[1478]&~m[1480]&m[1481]&m[1482])|(~m[681]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[681]&~m[1478]&m[1480]&m[1481]&m[1482])|(m[681]&m[1478]&m[1480]&m[1481]&m[1482]));
    m[1484] = (((m[694]&~m[1483]&~m[1485]&~m[1486]&~m[1487])|(~m[694]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(m[694]&m[1483]&~m[1485]&m[1486]&~m[1487])|(m[694]&~m[1483]&m[1485]&m[1486]&~m[1487])|(~m[694]&m[1483]&~m[1485]&~m[1486]&m[1487])|(~m[694]&~m[1483]&m[1485]&~m[1486]&m[1487])|(m[694]&m[1483]&m[1485]&~m[1486]&m[1487])|(~m[694]&m[1483]&m[1485]&m[1486]&m[1487]))&UnbiasedRNG[355])|((m[694]&~m[1483]&~m[1485]&m[1486]&~m[1487])|(~m[694]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[694]&~m[1483]&~m[1485]&~m[1486]&m[1487])|(m[694]&m[1483]&~m[1485]&~m[1486]&m[1487])|(m[694]&~m[1483]&m[1485]&~m[1486]&m[1487])|(~m[694]&~m[1483]&~m[1485]&m[1486]&m[1487])|(m[694]&~m[1483]&~m[1485]&m[1486]&m[1487])|(~m[694]&m[1483]&~m[1485]&m[1486]&m[1487])|(m[694]&m[1483]&~m[1485]&m[1486]&m[1487])|(~m[694]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[694]&~m[1483]&m[1485]&m[1486]&m[1487])|(m[694]&m[1483]&m[1485]&m[1486]&m[1487]));
    m[1489] = (((m[707]&~m[1488]&~m[1490]&~m[1491]&~m[1492])|(~m[707]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(m[707]&m[1488]&~m[1490]&m[1491]&~m[1492])|(m[707]&~m[1488]&m[1490]&m[1491]&~m[1492])|(~m[707]&m[1488]&~m[1490]&~m[1491]&m[1492])|(~m[707]&~m[1488]&m[1490]&~m[1491]&m[1492])|(m[707]&m[1488]&m[1490]&~m[1491]&m[1492])|(~m[707]&m[1488]&m[1490]&m[1491]&m[1492]))&UnbiasedRNG[356])|((m[707]&~m[1488]&~m[1490]&m[1491]&~m[1492])|(~m[707]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[707]&~m[1488]&~m[1490]&~m[1491]&m[1492])|(m[707]&m[1488]&~m[1490]&~m[1491]&m[1492])|(m[707]&~m[1488]&m[1490]&~m[1491]&m[1492])|(~m[707]&~m[1488]&~m[1490]&m[1491]&m[1492])|(m[707]&~m[1488]&~m[1490]&m[1491]&m[1492])|(~m[707]&m[1488]&~m[1490]&m[1491]&m[1492])|(m[707]&m[1488]&~m[1490]&m[1491]&m[1492])|(~m[707]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[707]&~m[1488]&m[1490]&m[1491]&m[1492])|(m[707]&m[1488]&m[1490]&m[1491]&m[1492]));
    m[1494] = (((m[720]&~m[1493]&~m[1495]&~m[1496]&~m[1497])|(~m[720]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(m[720]&m[1493]&~m[1495]&m[1496]&~m[1497])|(m[720]&~m[1493]&m[1495]&m[1496]&~m[1497])|(~m[720]&m[1493]&~m[1495]&~m[1496]&m[1497])|(~m[720]&~m[1493]&m[1495]&~m[1496]&m[1497])|(m[720]&m[1493]&m[1495]&~m[1496]&m[1497])|(~m[720]&m[1493]&m[1495]&m[1496]&m[1497]))&UnbiasedRNG[357])|((m[720]&~m[1493]&~m[1495]&m[1496]&~m[1497])|(~m[720]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[720]&~m[1493]&~m[1495]&~m[1496]&m[1497])|(m[720]&m[1493]&~m[1495]&~m[1496]&m[1497])|(m[720]&~m[1493]&m[1495]&~m[1496]&m[1497])|(~m[720]&~m[1493]&~m[1495]&m[1496]&m[1497])|(m[720]&~m[1493]&~m[1495]&m[1496]&m[1497])|(~m[720]&m[1493]&~m[1495]&m[1496]&m[1497])|(m[720]&m[1493]&~m[1495]&m[1496]&m[1497])|(~m[720]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[720]&~m[1493]&m[1495]&m[1496]&m[1497])|(m[720]&m[1493]&m[1495]&m[1496]&m[1497]));
    m[1499] = (((m[643]&~m[1498]&~m[1500]&~m[1501]&~m[1502])|(~m[643]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(m[643]&m[1498]&~m[1500]&m[1501]&~m[1502])|(m[643]&~m[1498]&m[1500]&m[1501]&~m[1502])|(~m[643]&m[1498]&~m[1500]&~m[1501]&m[1502])|(~m[643]&~m[1498]&m[1500]&~m[1501]&m[1502])|(m[643]&m[1498]&m[1500]&~m[1501]&m[1502])|(~m[643]&m[1498]&m[1500]&m[1501]&m[1502]))&UnbiasedRNG[358])|((m[643]&~m[1498]&~m[1500]&m[1501]&~m[1502])|(~m[643]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[643]&~m[1498]&~m[1500]&~m[1501]&m[1502])|(m[643]&m[1498]&~m[1500]&~m[1501]&m[1502])|(m[643]&~m[1498]&m[1500]&~m[1501]&m[1502])|(~m[643]&~m[1498]&~m[1500]&m[1501]&m[1502])|(m[643]&~m[1498]&~m[1500]&m[1501]&m[1502])|(~m[643]&m[1498]&~m[1500]&m[1501]&m[1502])|(m[643]&m[1498]&~m[1500]&m[1501]&m[1502])|(~m[643]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[643]&~m[1498]&m[1500]&m[1501]&m[1502])|(m[643]&m[1498]&m[1500]&m[1501]&m[1502]));
    m[1504] = (((m[656]&~m[1503]&~m[1505]&~m[1506]&~m[1507])|(~m[656]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(m[656]&m[1503]&~m[1505]&m[1506]&~m[1507])|(m[656]&~m[1503]&m[1505]&m[1506]&~m[1507])|(~m[656]&m[1503]&~m[1505]&~m[1506]&m[1507])|(~m[656]&~m[1503]&m[1505]&~m[1506]&m[1507])|(m[656]&m[1503]&m[1505]&~m[1506]&m[1507])|(~m[656]&m[1503]&m[1505]&m[1506]&m[1507]))&UnbiasedRNG[359])|((m[656]&~m[1503]&~m[1505]&m[1506]&~m[1507])|(~m[656]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[656]&~m[1503]&~m[1505]&~m[1506]&m[1507])|(m[656]&m[1503]&~m[1505]&~m[1506]&m[1507])|(m[656]&~m[1503]&m[1505]&~m[1506]&m[1507])|(~m[656]&~m[1503]&~m[1505]&m[1506]&m[1507])|(m[656]&~m[1503]&~m[1505]&m[1506]&m[1507])|(~m[656]&m[1503]&~m[1505]&m[1506]&m[1507])|(m[656]&m[1503]&~m[1505]&m[1506]&m[1507])|(~m[656]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[656]&~m[1503]&m[1505]&m[1506]&m[1507])|(m[656]&m[1503]&m[1505]&m[1506]&m[1507]));
    m[1509] = (((m[669]&~m[1508]&~m[1510]&~m[1511]&~m[1512])|(~m[669]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(m[669]&m[1508]&~m[1510]&m[1511]&~m[1512])|(m[669]&~m[1508]&m[1510]&m[1511]&~m[1512])|(~m[669]&m[1508]&~m[1510]&~m[1511]&m[1512])|(~m[669]&~m[1508]&m[1510]&~m[1511]&m[1512])|(m[669]&m[1508]&m[1510]&~m[1511]&m[1512])|(~m[669]&m[1508]&m[1510]&m[1511]&m[1512]))&UnbiasedRNG[360])|((m[669]&~m[1508]&~m[1510]&m[1511]&~m[1512])|(~m[669]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[669]&~m[1508]&~m[1510]&~m[1511]&m[1512])|(m[669]&m[1508]&~m[1510]&~m[1511]&m[1512])|(m[669]&~m[1508]&m[1510]&~m[1511]&m[1512])|(~m[669]&~m[1508]&~m[1510]&m[1511]&m[1512])|(m[669]&~m[1508]&~m[1510]&m[1511]&m[1512])|(~m[669]&m[1508]&~m[1510]&m[1511]&m[1512])|(m[669]&m[1508]&~m[1510]&m[1511]&m[1512])|(~m[669]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[669]&~m[1508]&m[1510]&m[1511]&m[1512])|(m[669]&m[1508]&m[1510]&m[1511]&m[1512]));
    m[1514] = (((m[682]&~m[1513]&~m[1515]&~m[1516]&~m[1517])|(~m[682]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(m[682]&m[1513]&~m[1515]&m[1516]&~m[1517])|(m[682]&~m[1513]&m[1515]&m[1516]&~m[1517])|(~m[682]&m[1513]&~m[1515]&~m[1516]&m[1517])|(~m[682]&~m[1513]&m[1515]&~m[1516]&m[1517])|(m[682]&m[1513]&m[1515]&~m[1516]&m[1517])|(~m[682]&m[1513]&m[1515]&m[1516]&m[1517]))&UnbiasedRNG[361])|((m[682]&~m[1513]&~m[1515]&m[1516]&~m[1517])|(~m[682]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[682]&~m[1513]&~m[1515]&~m[1516]&m[1517])|(m[682]&m[1513]&~m[1515]&~m[1516]&m[1517])|(m[682]&~m[1513]&m[1515]&~m[1516]&m[1517])|(~m[682]&~m[1513]&~m[1515]&m[1516]&m[1517])|(m[682]&~m[1513]&~m[1515]&m[1516]&m[1517])|(~m[682]&m[1513]&~m[1515]&m[1516]&m[1517])|(m[682]&m[1513]&~m[1515]&m[1516]&m[1517])|(~m[682]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[682]&~m[1513]&m[1515]&m[1516]&m[1517])|(m[682]&m[1513]&m[1515]&m[1516]&m[1517]));
    m[1519] = (((m[695]&~m[1518]&~m[1520]&~m[1521]&~m[1522])|(~m[695]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(m[695]&m[1518]&~m[1520]&m[1521]&~m[1522])|(m[695]&~m[1518]&m[1520]&m[1521]&~m[1522])|(~m[695]&m[1518]&~m[1520]&~m[1521]&m[1522])|(~m[695]&~m[1518]&m[1520]&~m[1521]&m[1522])|(m[695]&m[1518]&m[1520]&~m[1521]&m[1522])|(~m[695]&m[1518]&m[1520]&m[1521]&m[1522]))&UnbiasedRNG[362])|((m[695]&~m[1518]&~m[1520]&m[1521]&~m[1522])|(~m[695]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[695]&~m[1518]&~m[1520]&~m[1521]&m[1522])|(m[695]&m[1518]&~m[1520]&~m[1521]&m[1522])|(m[695]&~m[1518]&m[1520]&~m[1521]&m[1522])|(~m[695]&~m[1518]&~m[1520]&m[1521]&m[1522])|(m[695]&~m[1518]&~m[1520]&m[1521]&m[1522])|(~m[695]&m[1518]&~m[1520]&m[1521]&m[1522])|(m[695]&m[1518]&~m[1520]&m[1521]&m[1522])|(~m[695]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[695]&~m[1518]&m[1520]&m[1521]&m[1522])|(m[695]&m[1518]&m[1520]&m[1521]&m[1522]));
    m[1524] = (((m[708]&~m[1523]&~m[1525]&~m[1526]&~m[1527])|(~m[708]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(m[708]&m[1523]&~m[1525]&m[1526]&~m[1527])|(m[708]&~m[1523]&m[1525]&m[1526]&~m[1527])|(~m[708]&m[1523]&~m[1525]&~m[1526]&m[1527])|(~m[708]&~m[1523]&m[1525]&~m[1526]&m[1527])|(m[708]&m[1523]&m[1525]&~m[1526]&m[1527])|(~m[708]&m[1523]&m[1525]&m[1526]&m[1527]))&UnbiasedRNG[363])|((m[708]&~m[1523]&~m[1525]&m[1526]&~m[1527])|(~m[708]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[708]&~m[1523]&~m[1525]&~m[1526]&m[1527])|(m[708]&m[1523]&~m[1525]&~m[1526]&m[1527])|(m[708]&~m[1523]&m[1525]&~m[1526]&m[1527])|(~m[708]&~m[1523]&~m[1525]&m[1526]&m[1527])|(m[708]&~m[1523]&~m[1525]&m[1526]&m[1527])|(~m[708]&m[1523]&~m[1525]&m[1526]&m[1527])|(m[708]&m[1523]&~m[1525]&m[1526]&m[1527])|(~m[708]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[708]&~m[1523]&m[1525]&m[1526]&m[1527])|(m[708]&m[1523]&m[1525]&m[1526]&m[1527]));
    m[1529] = (((m[721]&~m[1528]&~m[1530]&~m[1531]&~m[1532])|(~m[721]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(m[721]&m[1528]&~m[1530]&m[1531]&~m[1532])|(m[721]&~m[1528]&m[1530]&m[1531]&~m[1532])|(~m[721]&m[1528]&~m[1530]&~m[1531]&m[1532])|(~m[721]&~m[1528]&m[1530]&~m[1531]&m[1532])|(m[721]&m[1528]&m[1530]&~m[1531]&m[1532])|(~m[721]&m[1528]&m[1530]&m[1531]&m[1532]))&UnbiasedRNG[364])|((m[721]&~m[1528]&~m[1530]&m[1531]&~m[1532])|(~m[721]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[721]&~m[1528]&~m[1530]&~m[1531]&m[1532])|(m[721]&m[1528]&~m[1530]&~m[1531]&m[1532])|(m[721]&~m[1528]&m[1530]&~m[1531]&m[1532])|(~m[721]&~m[1528]&~m[1530]&m[1531]&m[1532])|(m[721]&~m[1528]&~m[1530]&m[1531]&m[1532])|(~m[721]&m[1528]&~m[1530]&m[1531]&m[1532])|(m[721]&m[1528]&~m[1530]&m[1531]&m[1532])|(~m[721]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[721]&~m[1528]&m[1530]&m[1531]&m[1532])|(m[721]&m[1528]&m[1530]&m[1531]&m[1532]));
    m[1534] = (((m[657]&~m[1533]&~m[1535]&~m[1536]&~m[1537])|(~m[657]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(m[657]&m[1533]&~m[1535]&m[1536]&~m[1537])|(m[657]&~m[1533]&m[1535]&m[1536]&~m[1537])|(~m[657]&m[1533]&~m[1535]&~m[1536]&m[1537])|(~m[657]&~m[1533]&m[1535]&~m[1536]&m[1537])|(m[657]&m[1533]&m[1535]&~m[1536]&m[1537])|(~m[657]&m[1533]&m[1535]&m[1536]&m[1537]))&UnbiasedRNG[365])|((m[657]&~m[1533]&~m[1535]&m[1536]&~m[1537])|(~m[657]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[657]&~m[1533]&~m[1535]&~m[1536]&m[1537])|(m[657]&m[1533]&~m[1535]&~m[1536]&m[1537])|(m[657]&~m[1533]&m[1535]&~m[1536]&m[1537])|(~m[657]&~m[1533]&~m[1535]&m[1536]&m[1537])|(m[657]&~m[1533]&~m[1535]&m[1536]&m[1537])|(~m[657]&m[1533]&~m[1535]&m[1536]&m[1537])|(m[657]&m[1533]&~m[1535]&m[1536]&m[1537])|(~m[657]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[657]&~m[1533]&m[1535]&m[1536]&m[1537])|(m[657]&m[1533]&m[1535]&m[1536]&m[1537]));
    m[1539] = (((m[670]&~m[1538]&~m[1540]&~m[1541]&~m[1542])|(~m[670]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(m[670]&m[1538]&~m[1540]&m[1541]&~m[1542])|(m[670]&~m[1538]&m[1540]&m[1541]&~m[1542])|(~m[670]&m[1538]&~m[1540]&~m[1541]&m[1542])|(~m[670]&~m[1538]&m[1540]&~m[1541]&m[1542])|(m[670]&m[1538]&m[1540]&~m[1541]&m[1542])|(~m[670]&m[1538]&m[1540]&m[1541]&m[1542]))&UnbiasedRNG[366])|((m[670]&~m[1538]&~m[1540]&m[1541]&~m[1542])|(~m[670]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[670]&~m[1538]&~m[1540]&~m[1541]&m[1542])|(m[670]&m[1538]&~m[1540]&~m[1541]&m[1542])|(m[670]&~m[1538]&m[1540]&~m[1541]&m[1542])|(~m[670]&~m[1538]&~m[1540]&m[1541]&m[1542])|(m[670]&~m[1538]&~m[1540]&m[1541]&m[1542])|(~m[670]&m[1538]&~m[1540]&m[1541]&m[1542])|(m[670]&m[1538]&~m[1540]&m[1541]&m[1542])|(~m[670]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[670]&~m[1538]&m[1540]&m[1541]&m[1542])|(m[670]&m[1538]&m[1540]&m[1541]&m[1542]));
    m[1544] = (((m[683]&~m[1543]&~m[1545]&~m[1546]&~m[1547])|(~m[683]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(m[683]&m[1543]&~m[1545]&m[1546]&~m[1547])|(m[683]&~m[1543]&m[1545]&m[1546]&~m[1547])|(~m[683]&m[1543]&~m[1545]&~m[1546]&m[1547])|(~m[683]&~m[1543]&m[1545]&~m[1546]&m[1547])|(m[683]&m[1543]&m[1545]&~m[1546]&m[1547])|(~m[683]&m[1543]&m[1545]&m[1546]&m[1547]))&UnbiasedRNG[367])|((m[683]&~m[1543]&~m[1545]&m[1546]&~m[1547])|(~m[683]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[683]&~m[1543]&~m[1545]&~m[1546]&m[1547])|(m[683]&m[1543]&~m[1545]&~m[1546]&m[1547])|(m[683]&~m[1543]&m[1545]&~m[1546]&m[1547])|(~m[683]&~m[1543]&~m[1545]&m[1546]&m[1547])|(m[683]&~m[1543]&~m[1545]&m[1546]&m[1547])|(~m[683]&m[1543]&~m[1545]&m[1546]&m[1547])|(m[683]&m[1543]&~m[1545]&m[1546]&m[1547])|(~m[683]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[683]&~m[1543]&m[1545]&m[1546]&m[1547])|(m[683]&m[1543]&m[1545]&m[1546]&m[1547]));
    m[1549] = (((m[696]&~m[1548]&~m[1550]&~m[1551]&~m[1552])|(~m[696]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(m[696]&m[1548]&~m[1550]&m[1551]&~m[1552])|(m[696]&~m[1548]&m[1550]&m[1551]&~m[1552])|(~m[696]&m[1548]&~m[1550]&~m[1551]&m[1552])|(~m[696]&~m[1548]&m[1550]&~m[1551]&m[1552])|(m[696]&m[1548]&m[1550]&~m[1551]&m[1552])|(~m[696]&m[1548]&m[1550]&m[1551]&m[1552]))&UnbiasedRNG[368])|((m[696]&~m[1548]&~m[1550]&m[1551]&~m[1552])|(~m[696]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[696]&~m[1548]&~m[1550]&~m[1551]&m[1552])|(m[696]&m[1548]&~m[1550]&~m[1551]&m[1552])|(m[696]&~m[1548]&m[1550]&~m[1551]&m[1552])|(~m[696]&~m[1548]&~m[1550]&m[1551]&m[1552])|(m[696]&~m[1548]&~m[1550]&m[1551]&m[1552])|(~m[696]&m[1548]&~m[1550]&m[1551]&m[1552])|(m[696]&m[1548]&~m[1550]&m[1551]&m[1552])|(~m[696]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[696]&~m[1548]&m[1550]&m[1551]&m[1552])|(m[696]&m[1548]&m[1550]&m[1551]&m[1552]));
    m[1554] = (((m[709]&~m[1553]&~m[1555]&~m[1556]&~m[1557])|(~m[709]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(m[709]&m[1553]&~m[1555]&m[1556]&~m[1557])|(m[709]&~m[1553]&m[1555]&m[1556]&~m[1557])|(~m[709]&m[1553]&~m[1555]&~m[1556]&m[1557])|(~m[709]&~m[1553]&m[1555]&~m[1556]&m[1557])|(m[709]&m[1553]&m[1555]&~m[1556]&m[1557])|(~m[709]&m[1553]&m[1555]&m[1556]&m[1557]))&UnbiasedRNG[369])|((m[709]&~m[1553]&~m[1555]&m[1556]&~m[1557])|(~m[709]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[709]&~m[1553]&~m[1555]&~m[1556]&m[1557])|(m[709]&m[1553]&~m[1555]&~m[1556]&m[1557])|(m[709]&~m[1553]&m[1555]&~m[1556]&m[1557])|(~m[709]&~m[1553]&~m[1555]&m[1556]&m[1557])|(m[709]&~m[1553]&~m[1555]&m[1556]&m[1557])|(~m[709]&m[1553]&~m[1555]&m[1556]&m[1557])|(m[709]&m[1553]&~m[1555]&m[1556]&m[1557])|(~m[709]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[709]&~m[1553]&m[1555]&m[1556]&m[1557])|(m[709]&m[1553]&m[1555]&m[1556]&m[1557]));
    m[1559] = (((m[722]&~m[1558]&~m[1560]&~m[1561]&~m[1562])|(~m[722]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(m[722]&m[1558]&~m[1560]&m[1561]&~m[1562])|(m[722]&~m[1558]&m[1560]&m[1561]&~m[1562])|(~m[722]&m[1558]&~m[1560]&~m[1561]&m[1562])|(~m[722]&~m[1558]&m[1560]&~m[1561]&m[1562])|(m[722]&m[1558]&m[1560]&~m[1561]&m[1562])|(~m[722]&m[1558]&m[1560]&m[1561]&m[1562]))&UnbiasedRNG[370])|((m[722]&~m[1558]&~m[1560]&m[1561]&~m[1562])|(~m[722]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[722]&~m[1558]&~m[1560]&~m[1561]&m[1562])|(m[722]&m[1558]&~m[1560]&~m[1561]&m[1562])|(m[722]&~m[1558]&m[1560]&~m[1561]&m[1562])|(~m[722]&~m[1558]&~m[1560]&m[1561]&m[1562])|(m[722]&~m[1558]&~m[1560]&m[1561]&m[1562])|(~m[722]&m[1558]&~m[1560]&m[1561]&m[1562])|(m[722]&m[1558]&~m[1560]&m[1561]&m[1562])|(~m[722]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[722]&~m[1558]&m[1560]&m[1561]&m[1562])|(m[722]&m[1558]&m[1560]&m[1561]&m[1562]));
    m[1564] = (((m[671]&~m[1563]&~m[1565]&~m[1566]&~m[1567])|(~m[671]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(m[671]&m[1563]&~m[1565]&m[1566]&~m[1567])|(m[671]&~m[1563]&m[1565]&m[1566]&~m[1567])|(~m[671]&m[1563]&~m[1565]&~m[1566]&m[1567])|(~m[671]&~m[1563]&m[1565]&~m[1566]&m[1567])|(m[671]&m[1563]&m[1565]&~m[1566]&m[1567])|(~m[671]&m[1563]&m[1565]&m[1566]&m[1567]))&UnbiasedRNG[371])|((m[671]&~m[1563]&~m[1565]&m[1566]&~m[1567])|(~m[671]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[671]&~m[1563]&~m[1565]&~m[1566]&m[1567])|(m[671]&m[1563]&~m[1565]&~m[1566]&m[1567])|(m[671]&~m[1563]&m[1565]&~m[1566]&m[1567])|(~m[671]&~m[1563]&~m[1565]&m[1566]&m[1567])|(m[671]&~m[1563]&~m[1565]&m[1566]&m[1567])|(~m[671]&m[1563]&~m[1565]&m[1566]&m[1567])|(m[671]&m[1563]&~m[1565]&m[1566]&m[1567])|(~m[671]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[671]&~m[1563]&m[1565]&m[1566]&m[1567])|(m[671]&m[1563]&m[1565]&m[1566]&m[1567]));
    m[1569] = (((m[684]&~m[1568]&~m[1570]&~m[1571]&~m[1572])|(~m[684]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(m[684]&m[1568]&~m[1570]&m[1571]&~m[1572])|(m[684]&~m[1568]&m[1570]&m[1571]&~m[1572])|(~m[684]&m[1568]&~m[1570]&~m[1571]&m[1572])|(~m[684]&~m[1568]&m[1570]&~m[1571]&m[1572])|(m[684]&m[1568]&m[1570]&~m[1571]&m[1572])|(~m[684]&m[1568]&m[1570]&m[1571]&m[1572]))&UnbiasedRNG[372])|((m[684]&~m[1568]&~m[1570]&m[1571]&~m[1572])|(~m[684]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[684]&~m[1568]&~m[1570]&~m[1571]&m[1572])|(m[684]&m[1568]&~m[1570]&~m[1571]&m[1572])|(m[684]&~m[1568]&m[1570]&~m[1571]&m[1572])|(~m[684]&~m[1568]&~m[1570]&m[1571]&m[1572])|(m[684]&~m[1568]&~m[1570]&m[1571]&m[1572])|(~m[684]&m[1568]&~m[1570]&m[1571]&m[1572])|(m[684]&m[1568]&~m[1570]&m[1571]&m[1572])|(~m[684]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[684]&~m[1568]&m[1570]&m[1571]&m[1572])|(m[684]&m[1568]&m[1570]&m[1571]&m[1572]));
    m[1574] = (((m[697]&~m[1573]&~m[1575]&~m[1576]&~m[1577])|(~m[697]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(m[697]&m[1573]&~m[1575]&m[1576]&~m[1577])|(m[697]&~m[1573]&m[1575]&m[1576]&~m[1577])|(~m[697]&m[1573]&~m[1575]&~m[1576]&m[1577])|(~m[697]&~m[1573]&m[1575]&~m[1576]&m[1577])|(m[697]&m[1573]&m[1575]&~m[1576]&m[1577])|(~m[697]&m[1573]&m[1575]&m[1576]&m[1577]))&UnbiasedRNG[373])|((m[697]&~m[1573]&~m[1575]&m[1576]&~m[1577])|(~m[697]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[697]&~m[1573]&~m[1575]&~m[1576]&m[1577])|(m[697]&m[1573]&~m[1575]&~m[1576]&m[1577])|(m[697]&~m[1573]&m[1575]&~m[1576]&m[1577])|(~m[697]&~m[1573]&~m[1575]&m[1576]&m[1577])|(m[697]&~m[1573]&~m[1575]&m[1576]&m[1577])|(~m[697]&m[1573]&~m[1575]&m[1576]&m[1577])|(m[697]&m[1573]&~m[1575]&m[1576]&m[1577])|(~m[697]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[697]&~m[1573]&m[1575]&m[1576]&m[1577])|(m[697]&m[1573]&m[1575]&m[1576]&m[1577]));
    m[1579] = (((m[710]&~m[1578]&~m[1580]&~m[1581]&~m[1582])|(~m[710]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(m[710]&m[1578]&~m[1580]&m[1581]&~m[1582])|(m[710]&~m[1578]&m[1580]&m[1581]&~m[1582])|(~m[710]&m[1578]&~m[1580]&~m[1581]&m[1582])|(~m[710]&~m[1578]&m[1580]&~m[1581]&m[1582])|(m[710]&m[1578]&m[1580]&~m[1581]&m[1582])|(~m[710]&m[1578]&m[1580]&m[1581]&m[1582]))&UnbiasedRNG[374])|((m[710]&~m[1578]&~m[1580]&m[1581]&~m[1582])|(~m[710]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[710]&~m[1578]&~m[1580]&~m[1581]&m[1582])|(m[710]&m[1578]&~m[1580]&~m[1581]&m[1582])|(m[710]&~m[1578]&m[1580]&~m[1581]&m[1582])|(~m[710]&~m[1578]&~m[1580]&m[1581]&m[1582])|(m[710]&~m[1578]&~m[1580]&m[1581]&m[1582])|(~m[710]&m[1578]&~m[1580]&m[1581]&m[1582])|(m[710]&m[1578]&~m[1580]&m[1581]&m[1582])|(~m[710]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[710]&~m[1578]&m[1580]&m[1581]&m[1582])|(m[710]&m[1578]&m[1580]&m[1581]&m[1582]));
    m[1584] = (((m[723]&~m[1583]&~m[1585]&~m[1586]&~m[1587])|(~m[723]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(m[723]&m[1583]&~m[1585]&m[1586]&~m[1587])|(m[723]&~m[1583]&m[1585]&m[1586]&~m[1587])|(~m[723]&m[1583]&~m[1585]&~m[1586]&m[1587])|(~m[723]&~m[1583]&m[1585]&~m[1586]&m[1587])|(m[723]&m[1583]&m[1585]&~m[1586]&m[1587])|(~m[723]&m[1583]&m[1585]&m[1586]&m[1587]))&UnbiasedRNG[375])|((m[723]&~m[1583]&~m[1585]&m[1586]&~m[1587])|(~m[723]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[723]&~m[1583]&~m[1585]&~m[1586]&m[1587])|(m[723]&m[1583]&~m[1585]&~m[1586]&m[1587])|(m[723]&~m[1583]&m[1585]&~m[1586]&m[1587])|(~m[723]&~m[1583]&~m[1585]&m[1586]&m[1587])|(m[723]&~m[1583]&~m[1585]&m[1586]&m[1587])|(~m[723]&m[1583]&~m[1585]&m[1586]&m[1587])|(m[723]&m[1583]&~m[1585]&m[1586]&m[1587])|(~m[723]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[723]&~m[1583]&m[1585]&m[1586]&m[1587])|(m[723]&m[1583]&m[1585]&m[1586]&m[1587]));
    m[1589] = (((m[685]&~m[1588]&~m[1590]&~m[1591]&~m[1592])|(~m[685]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(m[685]&m[1588]&~m[1590]&m[1591]&~m[1592])|(m[685]&~m[1588]&m[1590]&m[1591]&~m[1592])|(~m[685]&m[1588]&~m[1590]&~m[1591]&m[1592])|(~m[685]&~m[1588]&m[1590]&~m[1591]&m[1592])|(m[685]&m[1588]&m[1590]&~m[1591]&m[1592])|(~m[685]&m[1588]&m[1590]&m[1591]&m[1592]))&UnbiasedRNG[376])|((m[685]&~m[1588]&~m[1590]&m[1591]&~m[1592])|(~m[685]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[685]&~m[1588]&~m[1590]&~m[1591]&m[1592])|(m[685]&m[1588]&~m[1590]&~m[1591]&m[1592])|(m[685]&~m[1588]&m[1590]&~m[1591]&m[1592])|(~m[685]&~m[1588]&~m[1590]&m[1591]&m[1592])|(m[685]&~m[1588]&~m[1590]&m[1591]&m[1592])|(~m[685]&m[1588]&~m[1590]&m[1591]&m[1592])|(m[685]&m[1588]&~m[1590]&m[1591]&m[1592])|(~m[685]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[685]&~m[1588]&m[1590]&m[1591]&m[1592])|(m[685]&m[1588]&m[1590]&m[1591]&m[1592]));
    m[1594] = (((m[698]&~m[1593]&~m[1595]&~m[1596]&~m[1597])|(~m[698]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(m[698]&m[1593]&~m[1595]&m[1596]&~m[1597])|(m[698]&~m[1593]&m[1595]&m[1596]&~m[1597])|(~m[698]&m[1593]&~m[1595]&~m[1596]&m[1597])|(~m[698]&~m[1593]&m[1595]&~m[1596]&m[1597])|(m[698]&m[1593]&m[1595]&~m[1596]&m[1597])|(~m[698]&m[1593]&m[1595]&m[1596]&m[1597]))&UnbiasedRNG[377])|((m[698]&~m[1593]&~m[1595]&m[1596]&~m[1597])|(~m[698]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[698]&~m[1593]&~m[1595]&~m[1596]&m[1597])|(m[698]&m[1593]&~m[1595]&~m[1596]&m[1597])|(m[698]&~m[1593]&m[1595]&~m[1596]&m[1597])|(~m[698]&~m[1593]&~m[1595]&m[1596]&m[1597])|(m[698]&~m[1593]&~m[1595]&m[1596]&m[1597])|(~m[698]&m[1593]&~m[1595]&m[1596]&m[1597])|(m[698]&m[1593]&~m[1595]&m[1596]&m[1597])|(~m[698]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[698]&~m[1593]&m[1595]&m[1596]&m[1597])|(m[698]&m[1593]&m[1595]&m[1596]&m[1597]));
    m[1599] = (((m[711]&~m[1598]&~m[1600]&~m[1601]&~m[1602])|(~m[711]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(m[711]&m[1598]&~m[1600]&m[1601]&~m[1602])|(m[711]&~m[1598]&m[1600]&m[1601]&~m[1602])|(~m[711]&m[1598]&~m[1600]&~m[1601]&m[1602])|(~m[711]&~m[1598]&m[1600]&~m[1601]&m[1602])|(m[711]&m[1598]&m[1600]&~m[1601]&m[1602])|(~m[711]&m[1598]&m[1600]&m[1601]&m[1602]))&UnbiasedRNG[378])|((m[711]&~m[1598]&~m[1600]&m[1601]&~m[1602])|(~m[711]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[711]&~m[1598]&~m[1600]&~m[1601]&m[1602])|(m[711]&m[1598]&~m[1600]&~m[1601]&m[1602])|(m[711]&~m[1598]&m[1600]&~m[1601]&m[1602])|(~m[711]&~m[1598]&~m[1600]&m[1601]&m[1602])|(m[711]&~m[1598]&~m[1600]&m[1601]&m[1602])|(~m[711]&m[1598]&~m[1600]&m[1601]&m[1602])|(m[711]&m[1598]&~m[1600]&m[1601]&m[1602])|(~m[711]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[711]&~m[1598]&m[1600]&m[1601]&m[1602])|(m[711]&m[1598]&m[1600]&m[1601]&m[1602]));
    m[1604] = (((m[724]&~m[1603]&~m[1605]&~m[1606]&~m[1607])|(~m[724]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(m[724]&m[1603]&~m[1605]&m[1606]&~m[1607])|(m[724]&~m[1603]&m[1605]&m[1606]&~m[1607])|(~m[724]&m[1603]&~m[1605]&~m[1606]&m[1607])|(~m[724]&~m[1603]&m[1605]&~m[1606]&m[1607])|(m[724]&m[1603]&m[1605]&~m[1606]&m[1607])|(~m[724]&m[1603]&m[1605]&m[1606]&m[1607]))&UnbiasedRNG[379])|((m[724]&~m[1603]&~m[1605]&m[1606]&~m[1607])|(~m[724]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[724]&~m[1603]&~m[1605]&~m[1606]&m[1607])|(m[724]&m[1603]&~m[1605]&~m[1606]&m[1607])|(m[724]&~m[1603]&m[1605]&~m[1606]&m[1607])|(~m[724]&~m[1603]&~m[1605]&m[1606]&m[1607])|(m[724]&~m[1603]&~m[1605]&m[1606]&m[1607])|(~m[724]&m[1603]&~m[1605]&m[1606]&m[1607])|(m[724]&m[1603]&~m[1605]&m[1606]&m[1607])|(~m[724]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[724]&~m[1603]&m[1605]&m[1606]&m[1607])|(m[724]&m[1603]&m[1605]&m[1606]&m[1607]));
    m[1609] = (((m[699]&~m[1608]&~m[1610]&~m[1611]&~m[1612])|(~m[699]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(m[699]&m[1608]&~m[1610]&m[1611]&~m[1612])|(m[699]&~m[1608]&m[1610]&m[1611]&~m[1612])|(~m[699]&m[1608]&~m[1610]&~m[1611]&m[1612])|(~m[699]&~m[1608]&m[1610]&~m[1611]&m[1612])|(m[699]&m[1608]&m[1610]&~m[1611]&m[1612])|(~m[699]&m[1608]&m[1610]&m[1611]&m[1612]))&UnbiasedRNG[380])|((m[699]&~m[1608]&~m[1610]&m[1611]&~m[1612])|(~m[699]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[699]&~m[1608]&~m[1610]&~m[1611]&m[1612])|(m[699]&m[1608]&~m[1610]&~m[1611]&m[1612])|(m[699]&~m[1608]&m[1610]&~m[1611]&m[1612])|(~m[699]&~m[1608]&~m[1610]&m[1611]&m[1612])|(m[699]&~m[1608]&~m[1610]&m[1611]&m[1612])|(~m[699]&m[1608]&~m[1610]&m[1611]&m[1612])|(m[699]&m[1608]&~m[1610]&m[1611]&m[1612])|(~m[699]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[699]&~m[1608]&m[1610]&m[1611]&m[1612])|(m[699]&m[1608]&m[1610]&m[1611]&m[1612]));
    m[1614] = (((m[712]&~m[1613]&~m[1615]&~m[1616]&~m[1617])|(~m[712]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(m[712]&m[1613]&~m[1615]&m[1616]&~m[1617])|(m[712]&~m[1613]&m[1615]&m[1616]&~m[1617])|(~m[712]&m[1613]&~m[1615]&~m[1616]&m[1617])|(~m[712]&~m[1613]&m[1615]&~m[1616]&m[1617])|(m[712]&m[1613]&m[1615]&~m[1616]&m[1617])|(~m[712]&m[1613]&m[1615]&m[1616]&m[1617]))&UnbiasedRNG[381])|((m[712]&~m[1613]&~m[1615]&m[1616]&~m[1617])|(~m[712]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[712]&~m[1613]&~m[1615]&~m[1616]&m[1617])|(m[712]&m[1613]&~m[1615]&~m[1616]&m[1617])|(m[712]&~m[1613]&m[1615]&~m[1616]&m[1617])|(~m[712]&~m[1613]&~m[1615]&m[1616]&m[1617])|(m[712]&~m[1613]&~m[1615]&m[1616]&m[1617])|(~m[712]&m[1613]&~m[1615]&m[1616]&m[1617])|(m[712]&m[1613]&~m[1615]&m[1616]&m[1617])|(~m[712]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[712]&~m[1613]&m[1615]&m[1616]&m[1617])|(m[712]&m[1613]&m[1615]&m[1616]&m[1617]));
    m[1619] = (((m[725]&~m[1618]&~m[1620]&~m[1621]&~m[1622])|(~m[725]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(m[725]&m[1618]&~m[1620]&m[1621]&~m[1622])|(m[725]&~m[1618]&m[1620]&m[1621]&~m[1622])|(~m[725]&m[1618]&~m[1620]&~m[1621]&m[1622])|(~m[725]&~m[1618]&m[1620]&~m[1621]&m[1622])|(m[725]&m[1618]&m[1620]&~m[1621]&m[1622])|(~m[725]&m[1618]&m[1620]&m[1621]&m[1622]))&UnbiasedRNG[382])|((m[725]&~m[1618]&~m[1620]&m[1621]&~m[1622])|(~m[725]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[725]&~m[1618]&~m[1620]&~m[1621]&m[1622])|(m[725]&m[1618]&~m[1620]&~m[1621]&m[1622])|(m[725]&~m[1618]&m[1620]&~m[1621]&m[1622])|(~m[725]&~m[1618]&~m[1620]&m[1621]&m[1622])|(m[725]&~m[1618]&~m[1620]&m[1621]&m[1622])|(~m[725]&m[1618]&~m[1620]&m[1621]&m[1622])|(m[725]&m[1618]&~m[1620]&m[1621]&m[1622])|(~m[725]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[725]&~m[1618]&m[1620]&m[1621]&m[1622])|(m[725]&m[1618]&m[1620]&m[1621]&m[1622]));
    m[1624] = (((m[713]&~m[1623]&~m[1625]&~m[1626]&~m[1627])|(~m[713]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(m[713]&m[1623]&~m[1625]&m[1626]&~m[1627])|(m[713]&~m[1623]&m[1625]&m[1626]&~m[1627])|(~m[713]&m[1623]&~m[1625]&~m[1626]&m[1627])|(~m[713]&~m[1623]&m[1625]&~m[1626]&m[1627])|(m[713]&m[1623]&m[1625]&~m[1626]&m[1627])|(~m[713]&m[1623]&m[1625]&m[1626]&m[1627]))&UnbiasedRNG[383])|((m[713]&~m[1623]&~m[1625]&m[1626]&~m[1627])|(~m[713]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[713]&~m[1623]&~m[1625]&~m[1626]&m[1627])|(m[713]&m[1623]&~m[1625]&~m[1626]&m[1627])|(m[713]&~m[1623]&m[1625]&~m[1626]&m[1627])|(~m[713]&~m[1623]&~m[1625]&m[1626]&m[1627])|(m[713]&~m[1623]&~m[1625]&m[1626]&m[1627])|(~m[713]&m[1623]&~m[1625]&m[1626]&m[1627])|(m[713]&m[1623]&~m[1625]&m[1626]&m[1627])|(~m[713]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[713]&~m[1623]&m[1625]&m[1626]&m[1627])|(m[713]&m[1623]&m[1625]&m[1626]&m[1627]));
    m[1629] = (((m[726]&~m[1628]&~m[1630]&~m[1631]&~m[1632])|(~m[726]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(m[726]&m[1628]&~m[1630]&m[1631]&~m[1632])|(m[726]&~m[1628]&m[1630]&m[1631]&~m[1632])|(~m[726]&m[1628]&~m[1630]&~m[1631]&m[1632])|(~m[726]&~m[1628]&m[1630]&~m[1631]&m[1632])|(m[726]&m[1628]&m[1630]&~m[1631]&m[1632])|(~m[726]&m[1628]&m[1630]&m[1631]&m[1632]))&UnbiasedRNG[384])|((m[726]&~m[1628]&~m[1630]&m[1631]&~m[1632])|(~m[726]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[726]&~m[1628]&~m[1630]&~m[1631]&m[1632])|(m[726]&m[1628]&~m[1630]&~m[1631]&m[1632])|(m[726]&~m[1628]&m[1630]&~m[1631]&m[1632])|(~m[726]&~m[1628]&~m[1630]&m[1631]&m[1632])|(m[726]&~m[1628]&~m[1630]&m[1631]&m[1632])|(~m[726]&m[1628]&~m[1630]&m[1631]&m[1632])|(m[726]&m[1628]&~m[1630]&m[1631]&m[1632])|(~m[726]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[726]&~m[1628]&m[1630]&m[1631]&m[1632])|(m[726]&m[1628]&m[1630]&m[1631]&m[1632]));
    m[1634] = (((m[727]&~m[1633]&~m[1635]&~m[1636]&~m[1637])|(~m[727]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(m[727]&m[1633]&~m[1635]&m[1636]&~m[1637])|(m[727]&~m[1633]&m[1635]&m[1636]&~m[1637])|(~m[727]&m[1633]&~m[1635]&~m[1636]&m[1637])|(~m[727]&~m[1633]&m[1635]&~m[1636]&m[1637])|(m[727]&m[1633]&m[1635]&~m[1636]&m[1637])|(~m[727]&m[1633]&m[1635]&m[1636]&m[1637]))&UnbiasedRNG[385])|((m[727]&~m[1633]&~m[1635]&m[1636]&~m[1637])|(~m[727]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[727]&~m[1633]&~m[1635]&~m[1636]&m[1637])|(m[727]&m[1633]&~m[1635]&~m[1636]&m[1637])|(m[727]&~m[1633]&m[1635]&~m[1636]&m[1637])|(~m[727]&~m[1633]&~m[1635]&m[1636]&m[1637])|(m[727]&~m[1633]&~m[1635]&m[1636]&m[1637])|(~m[727]&m[1633]&~m[1635]&m[1636]&m[1637])|(m[727]&m[1633]&~m[1635]&m[1636]&m[1637])|(~m[727]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[727]&~m[1633]&m[1635]&m[1636]&m[1637])|(m[727]&m[1633]&m[1635]&m[1636]&m[1637]));
end

always @(posedge color2_clk) begin
    m[336] = (((~m[42]&~m[140]&~m[532])|(m[42]&m[140]&~m[532]))&BiasedRNG[503])|(((m[42]&~m[140]&~m[532])|(~m[42]&m[140]&m[532]))&~BiasedRNG[503])|((~m[42]&~m[140]&m[532])|(m[42]&~m[140]&m[532])|(m[42]&m[140]&m[532]));
    m[337] = (((~m[42]&~m[154]&~m[533])|(m[42]&m[154]&~m[533]))&BiasedRNG[504])|(((m[42]&~m[154]&~m[533])|(~m[42]&m[154]&m[533]))&~BiasedRNG[504])|((~m[42]&~m[154]&m[533])|(m[42]&~m[154]&m[533])|(m[42]&m[154]&m[533]));
    m[338] = (((~m[98]&~m[168]&~m[534])|(m[98]&m[168]&~m[534]))&BiasedRNG[505])|(((m[98]&~m[168]&~m[534])|(~m[98]&m[168]&m[534]))&~BiasedRNG[505])|((~m[98]&~m[168]&m[534])|(m[98]&~m[168]&m[534])|(m[98]&m[168]&m[534]));
    m[339] = (((~m[98]&~m[182]&~m[535])|(m[98]&m[182]&~m[535]))&BiasedRNG[506])|(((m[98]&~m[182]&~m[535])|(~m[98]&m[182]&m[535]))&~BiasedRNG[506])|((~m[98]&~m[182]&m[535])|(m[98]&~m[182]&m[535])|(m[98]&m[182]&m[535]));
    m[340] = (((~m[98]&~m[196]&~m[536])|(m[98]&m[196]&~m[536]))&BiasedRNG[507])|(((m[98]&~m[196]&~m[536])|(~m[98]&m[196]&m[536]))&~BiasedRNG[507])|((~m[98]&~m[196]&m[536])|(m[98]&~m[196]&m[536])|(m[98]&m[196]&m[536]));
    m[341] = (((~m[98]&~m[210]&~m[537])|(m[98]&m[210]&~m[537]))&BiasedRNG[508])|(((m[98]&~m[210]&~m[537])|(~m[98]&m[210]&m[537]))&~BiasedRNG[508])|((~m[98]&~m[210]&m[537])|(m[98]&~m[210]&m[537])|(m[98]&m[210]&m[537]));
    m[350] = (((~m[43]&~m[141]&~m[546])|(m[43]&m[141]&~m[546]))&BiasedRNG[509])|(((m[43]&~m[141]&~m[546])|(~m[43]&m[141]&m[546]))&~BiasedRNG[509])|((~m[43]&~m[141]&m[546])|(m[43]&~m[141]&m[546])|(m[43]&m[141]&m[546]));
    m[351] = (((~m[43]&~m[155]&~m[547])|(m[43]&m[155]&~m[547]))&BiasedRNG[510])|(((m[43]&~m[155]&~m[547])|(~m[43]&m[155]&m[547]))&~BiasedRNG[510])|((~m[43]&~m[155]&m[547])|(m[43]&~m[155]&m[547])|(m[43]&m[155]&m[547]));
    m[352] = (((~m[101]&~m[169]&~m[548])|(m[101]&m[169]&~m[548]))&BiasedRNG[511])|(((m[101]&~m[169]&~m[548])|(~m[101]&m[169]&m[548]))&~BiasedRNG[511])|((~m[101]&~m[169]&m[548])|(m[101]&~m[169]&m[548])|(m[101]&m[169]&m[548]));
    m[353] = (((~m[101]&~m[183]&~m[549])|(m[101]&m[183]&~m[549]))&BiasedRNG[512])|(((m[101]&~m[183]&~m[549])|(~m[101]&m[183]&m[549]))&~BiasedRNG[512])|((~m[101]&~m[183]&m[549])|(m[101]&~m[183]&m[549])|(m[101]&m[183]&m[549]));
    m[354] = (((~m[101]&~m[197]&~m[550])|(m[101]&m[197]&~m[550]))&BiasedRNG[513])|(((m[101]&~m[197]&~m[550])|(~m[101]&m[197]&m[550]))&~BiasedRNG[513])|((~m[101]&~m[197]&m[550])|(m[101]&~m[197]&m[550])|(m[101]&m[197]&m[550]));
    m[355] = (((~m[101]&~m[211]&~m[551])|(m[101]&m[211]&~m[551]))&BiasedRNG[514])|(((m[101]&~m[211]&~m[551])|(~m[101]&m[211]&m[551]))&~BiasedRNG[514])|((~m[101]&~m[211]&m[551])|(m[101]&~m[211]&m[551])|(m[101]&m[211]&m[551]));
    m[364] = (((~m[44]&~m[142]&~m[560])|(m[44]&m[142]&~m[560]))&BiasedRNG[515])|(((m[44]&~m[142]&~m[560])|(~m[44]&m[142]&m[560]))&~BiasedRNG[515])|((~m[44]&~m[142]&m[560])|(m[44]&~m[142]&m[560])|(m[44]&m[142]&m[560]));
    m[365] = (((~m[44]&~m[156]&~m[561])|(m[44]&m[156]&~m[561]))&BiasedRNG[516])|(((m[44]&~m[156]&~m[561])|(~m[44]&m[156]&m[561]))&~BiasedRNG[516])|((~m[44]&~m[156]&m[561])|(m[44]&~m[156]&m[561])|(m[44]&m[156]&m[561]));
    m[366] = (((~m[104]&~m[170]&~m[562])|(m[104]&m[170]&~m[562]))&BiasedRNG[517])|(((m[104]&~m[170]&~m[562])|(~m[104]&m[170]&m[562]))&~BiasedRNG[517])|((~m[104]&~m[170]&m[562])|(m[104]&~m[170]&m[562])|(m[104]&m[170]&m[562]));
    m[367] = (((~m[104]&~m[184]&~m[563])|(m[104]&m[184]&~m[563]))&BiasedRNG[518])|(((m[104]&~m[184]&~m[563])|(~m[104]&m[184]&m[563]))&~BiasedRNG[518])|((~m[104]&~m[184]&m[563])|(m[104]&~m[184]&m[563])|(m[104]&m[184]&m[563]));
    m[368] = (((~m[104]&~m[198]&~m[564])|(m[104]&m[198]&~m[564]))&BiasedRNG[519])|(((m[104]&~m[198]&~m[564])|(~m[104]&m[198]&m[564]))&~BiasedRNG[519])|((~m[104]&~m[198]&m[564])|(m[104]&~m[198]&m[564])|(m[104]&m[198]&m[564]));
    m[369] = (((~m[104]&~m[212]&~m[565])|(m[104]&m[212]&~m[565]))&BiasedRNG[520])|(((m[104]&~m[212]&~m[565])|(~m[104]&m[212]&m[565]))&~BiasedRNG[520])|((~m[104]&~m[212]&m[565])|(m[104]&~m[212]&m[565])|(m[104]&m[212]&m[565]));
    m[378] = (((~m[45]&~m[143]&~m[574])|(m[45]&m[143]&~m[574]))&BiasedRNG[521])|(((m[45]&~m[143]&~m[574])|(~m[45]&m[143]&m[574]))&~BiasedRNG[521])|((~m[45]&~m[143]&m[574])|(m[45]&~m[143]&m[574])|(m[45]&m[143]&m[574]));
    m[379] = (((~m[45]&~m[157]&~m[575])|(m[45]&m[157]&~m[575]))&BiasedRNG[522])|(((m[45]&~m[157]&~m[575])|(~m[45]&m[157]&m[575]))&~BiasedRNG[522])|((~m[45]&~m[157]&m[575])|(m[45]&~m[157]&m[575])|(m[45]&m[157]&m[575]));
    m[380] = (((~m[107]&~m[171]&~m[576])|(m[107]&m[171]&~m[576]))&BiasedRNG[523])|(((m[107]&~m[171]&~m[576])|(~m[107]&m[171]&m[576]))&~BiasedRNG[523])|((~m[107]&~m[171]&m[576])|(m[107]&~m[171]&m[576])|(m[107]&m[171]&m[576]));
    m[381] = (((~m[107]&~m[185]&~m[577])|(m[107]&m[185]&~m[577]))&BiasedRNG[524])|(((m[107]&~m[185]&~m[577])|(~m[107]&m[185]&m[577]))&~BiasedRNG[524])|((~m[107]&~m[185]&m[577])|(m[107]&~m[185]&m[577])|(m[107]&m[185]&m[577]));
    m[382] = (((~m[107]&~m[199]&~m[578])|(m[107]&m[199]&~m[578]))&BiasedRNG[525])|(((m[107]&~m[199]&~m[578])|(~m[107]&m[199]&m[578]))&~BiasedRNG[525])|((~m[107]&~m[199]&m[578])|(m[107]&~m[199]&m[578])|(m[107]&m[199]&m[578]));
    m[383] = (((~m[107]&~m[213]&~m[579])|(m[107]&m[213]&~m[579]))&BiasedRNG[526])|(((m[107]&~m[213]&~m[579])|(~m[107]&m[213]&m[579]))&~BiasedRNG[526])|((~m[107]&~m[213]&m[579])|(m[107]&~m[213]&m[579])|(m[107]&m[213]&m[579]));
    m[392] = (((~m[46]&~m[144]&~m[588])|(m[46]&m[144]&~m[588]))&BiasedRNG[527])|(((m[46]&~m[144]&~m[588])|(~m[46]&m[144]&m[588]))&~BiasedRNG[527])|((~m[46]&~m[144]&m[588])|(m[46]&~m[144]&m[588])|(m[46]&m[144]&m[588]));
    m[393] = (((~m[46]&~m[158]&~m[589])|(m[46]&m[158]&~m[589]))&BiasedRNG[528])|(((m[46]&~m[158]&~m[589])|(~m[46]&m[158]&m[589]))&~BiasedRNG[528])|((~m[46]&~m[158]&m[589])|(m[46]&~m[158]&m[589])|(m[46]&m[158]&m[589]));
    m[394] = (((~m[110]&~m[172]&~m[590])|(m[110]&m[172]&~m[590]))&BiasedRNG[529])|(((m[110]&~m[172]&~m[590])|(~m[110]&m[172]&m[590]))&~BiasedRNG[529])|((~m[110]&~m[172]&m[590])|(m[110]&~m[172]&m[590])|(m[110]&m[172]&m[590]));
    m[395] = (((~m[110]&~m[186]&~m[591])|(m[110]&m[186]&~m[591]))&BiasedRNG[530])|(((m[110]&~m[186]&~m[591])|(~m[110]&m[186]&m[591]))&~BiasedRNG[530])|((~m[110]&~m[186]&m[591])|(m[110]&~m[186]&m[591])|(m[110]&m[186]&m[591]));
    m[396] = (((~m[110]&~m[200]&~m[592])|(m[110]&m[200]&~m[592]))&BiasedRNG[531])|(((m[110]&~m[200]&~m[592])|(~m[110]&m[200]&m[592]))&~BiasedRNG[531])|((~m[110]&~m[200]&m[592])|(m[110]&~m[200]&m[592])|(m[110]&m[200]&m[592]));
    m[397] = (((~m[110]&~m[214]&~m[593])|(m[110]&m[214]&~m[593]))&BiasedRNG[532])|(((m[110]&~m[214]&~m[593])|(~m[110]&m[214]&m[593]))&~BiasedRNG[532])|((~m[110]&~m[214]&m[593])|(m[110]&~m[214]&m[593])|(m[110]&m[214]&m[593]));
    m[406] = (((~m[47]&~m[145]&~m[602])|(m[47]&m[145]&~m[602]))&BiasedRNG[533])|(((m[47]&~m[145]&~m[602])|(~m[47]&m[145]&m[602]))&~BiasedRNG[533])|((~m[47]&~m[145]&m[602])|(m[47]&~m[145]&m[602])|(m[47]&m[145]&m[602]));
    m[407] = (((~m[47]&~m[159]&~m[603])|(m[47]&m[159]&~m[603]))&BiasedRNG[534])|(((m[47]&~m[159]&~m[603])|(~m[47]&m[159]&m[603]))&~BiasedRNG[534])|((~m[47]&~m[159]&m[603])|(m[47]&~m[159]&m[603])|(m[47]&m[159]&m[603]));
    m[408] = (((~m[113]&~m[173]&~m[604])|(m[113]&m[173]&~m[604]))&BiasedRNG[535])|(((m[113]&~m[173]&~m[604])|(~m[113]&m[173]&m[604]))&~BiasedRNG[535])|((~m[113]&~m[173]&m[604])|(m[113]&~m[173]&m[604])|(m[113]&m[173]&m[604]));
    m[409] = (((~m[113]&~m[187]&~m[605])|(m[113]&m[187]&~m[605]))&BiasedRNG[536])|(((m[113]&~m[187]&~m[605])|(~m[113]&m[187]&m[605]))&~BiasedRNG[536])|((~m[113]&~m[187]&m[605])|(m[113]&~m[187]&m[605])|(m[113]&m[187]&m[605]));
    m[410] = (((~m[113]&~m[201]&~m[606])|(m[113]&m[201]&~m[606]))&BiasedRNG[537])|(((m[113]&~m[201]&~m[606])|(~m[113]&m[201]&m[606]))&~BiasedRNG[537])|((~m[113]&~m[201]&m[606])|(m[113]&~m[201]&m[606])|(m[113]&m[201]&m[606]));
    m[411] = (((~m[113]&~m[215]&~m[607])|(m[113]&m[215]&~m[607]))&BiasedRNG[538])|(((m[113]&~m[215]&~m[607])|(~m[113]&m[215]&m[607]))&~BiasedRNG[538])|((~m[113]&~m[215]&m[607])|(m[113]&~m[215]&m[607])|(m[113]&m[215]&m[607]));
    m[426] = (((~m[117]&~m[230]&~m[622])|(m[117]&m[230]&~m[622]))&BiasedRNG[539])|(((m[117]&~m[230]&~m[622])|(~m[117]&m[230]&m[622]))&~BiasedRNG[539])|((~m[117]&~m[230]&m[622])|(m[117]&~m[230]&m[622])|(m[117]&m[230]&m[622]));
    m[427] = (((~m[117]&~m[244]&~m[623])|(m[117]&m[244]&~m[623]))&BiasedRNG[540])|(((m[117]&~m[244]&~m[623])|(~m[117]&m[244]&m[623]))&~BiasedRNG[540])|((~m[117]&~m[244]&m[623])|(m[117]&~m[244]&m[623])|(m[117]&m[244]&m[623]));
    m[428] = (((~m[117]&~m[258]&~m[624])|(m[117]&m[258]&~m[624]))&BiasedRNG[541])|(((m[117]&~m[258]&~m[624])|(~m[117]&m[258]&m[624]))&~BiasedRNG[541])|((~m[117]&~m[258]&m[624])|(m[117]&~m[258]&m[624])|(m[117]&m[258]&m[624]));
    m[429] = (((~m[117]&~m[272]&~m[625])|(m[117]&m[272]&~m[625]))&BiasedRNG[542])|(((m[117]&~m[272]&~m[625])|(~m[117]&m[272]&m[625]))&~BiasedRNG[542])|((~m[117]&~m[272]&m[625])|(m[117]&~m[272]&m[625])|(m[117]&m[272]&m[625]));
    m[430] = (((~m[118]&~m[286]&~m[626])|(m[118]&m[286]&~m[626]))&BiasedRNG[543])|(((m[118]&~m[286]&~m[626])|(~m[118]&m[286]&m[626]))&~BiasedRNG[543])|((~m[118]&~m[286]&m[626])|(m[118]&~m[286]&m[626])|(m[118]&m[286]&m[626]));
    m[431] = (((~m[118]&~m[300]&~m[627])|(m[118]&m[300]&~m[627]))&BiasedRNG[544])|(((m[118]&~m[300]&~m[627])|(~m[118]&m[300]&m[627]))&~BiasedRNG[544])|((~m[118]&~m[300]&m[627])|(m[118]&~m[300]&m[627])|(m[118]&m[300]&m[627]));
    m[432] = (((~m[118]&~m[314]&~m[628])|(m[118]&m[314]&~m[628]))&BiasedRNG[545])|(((m[118]&~m[314]&~m[628])|(~m[118]&m[314]&m[628]))&~BiasedRNG[545])|((~m[118]&~m[314]&m[628])|(m[118]&~m[314]&m[628])|(m[118]&m[314]&m[628]));
    m[433] = (((~m[118]&~m[328]&~m[629])|(m[118]&m[328]&~m[629]))&BiasedRNG[546])|(((m[118]&~m[328]&~m[629])|(~m[118]&m[328]&m[629]))&~BiasedRNG[546])|((~m[118]&~m[328]&m[629])|(m[118]&~m[328]&m[629])|(m[118]&m[328]&m[629]));
    m[440] = (((~m[120]&~m[231]&~m[636])|(m[120]&m[231]&~m[636]))&BiasedRNG[547])|(((m[120]&~m[231]&~m[636])|(~m[120]&m[231]&m[636]))&~BiasedRNG[547])|((~m[120]&~m[231]&m[636])|(m[120]&~m[231]&m[636])|(m[120]&m[231]&m[636]));
    m[441] = (((~m[120]&~m[245]&~m[637])|(m[120]&m[245]&~m[637]))&BiasedRNG[548])|(((m[120]&~m[245]&~m[637])|(~m[120]&m[245]&m[637]))&~BiasedRNG[548])|((~m[120]&~m[245]&m[637])|(m[120]&~m[245]&m[637])|(m[120]&m[245]&m[637]));
    m[442] = (((~m[120]&~m[259]&~m[638])|(m[120]&m[259]&~m[638]))&BiasedRNG[549])|(((m[120]&~m[259]&~m[638])|(~m[120]&m[259]&m[638]))&~BiasedRNG[549])|((~m[120]&~m[259]&m[638])|(m[120]&~m[259]&m[638])|(m[120]&m[259]&m[638]));
    m[443] = (((~m[120]&~m[273]&~m[639])|(m[120]&m[273]&~m[639]))&BiasedRNG[550])|(((m[120]&~m[273]&~m[639])|(~m[120]&m[273]&m[639]))&~BiasedRNG[550])|((~m[120]&~m[273]&m[639])|(m[120]&~m[273]&m[639])|(m[120]&m[273]&m[639]));
    m[444] = (((~m[121]&~m[287]&~m[640])|(m[121]&m[287]&~m[640]))&BiasedRNG[551])|(((m[121]&~m[287]&~m[640])|(~m[121]&m[287]&m[640]))&~BiasedRNG[551])|((~m[121]&~m[287]&m[640])|(m[121]&~m[287]&m[640])|(m[121]&m[287]&m[640]));
    m[445] = (((~m[121]&~m[301]&~m[641])|(m[121]&m[301]&~m[641]))&BiasedRNG[552])|(((m[121]&~m[301]&~m[641])|(~m[121]&m[301]&m[641]))&~BiasedRNG[552])|((~m[121]&~m[301]&m[641])|(m[121]&~m[301]&m[641])|(m[121]&m[301]&m[641]));
    m[446] = (((~m[121]&~m[315]&~m[642])|(m[121]&m[315]&~m[642]))&BiasedRNG[553])|(((m[121]&~m[315]&~m[642])|(~m[121]&m[315]&m[642]))&~BiasedRNG[553])|((~m[121]&~m[315]&m[642])|(m[121]&~m[315]&m[642])|(m[121]&m[315]&m[642]));
    m[447] = (((~m[121]&~m[329]&~m[643])|(m[121]&m[329]&~m[643]))&BiasedRNG[554])|(((m[121]&~m[329]&~m[643])|(~m[121]&m[329]&m[643]))&~BiasedRNG[554])|((~m[121]&~m[329]&m[643])|(m[121]&~m[329]&m[643])|(m[121]&m[329]&m[643]));
    m[454] = (((~m[123]&~m[232]&~m[650])|(m[123]&m[232]&~m[650]))&BiasedRNG[555])|(((m[123]&~m[232]&~m[650])|(~m[123]&m[232]&m[650]))&~BiasedRNG[555])|((~m[123]&~m[232]&m[650])|(m[123]&~m[232]&m[650])|(m[123]&m[232]&m[650]));
    m[455] = (((~m[123]&~m[246]&~m[651])|(m[123]&m[246]&~m[651]))&BiasedRNG[556])|(((m[123]&~m[246]&~m[651])|(~m[123]&m[246]&m[651]))&~BiasedRNG[556])|((~m[123]&~m[246]&m[651])|(m[123]&~m[246]&m[651])|(m[123]&m[246]&m[651]));
    m[456] = (((~m[123]&~m[260]&~m[652])|(m[123]&m[260]&~m[652]))&BiasedRNG[557])|(((m[123]&~m[260]&~m[652])|(~m[123]&m[260]&m[652]))&~BiasedRNG[557])|((~m[123]&~m[260]&m[652])|(m[123]&~m[260]&m[652])|(m[123]&m[260]&m[652]));
    m[457] = (((~m[123]&~m[274]&~m[653])|(m[123]&m[274]&~m[653]))&BiasedRNG[558])|(((m[123]&~m[274]&~m[653])|(~m[123]&m[274]&m[653]))&~BiasedRNG[558])|((~m[123]&~m[274]&m[653])|(m[123]&~m[274]&m[653])|(m[123]&m[274]&m[653]));
    m[458] = (((~m[124]&~m[288]&~m[654])|(m[124]&m[288]&~m[654]))&BiasedRNG[559])|(((m[124]&~m[288]&~m[654])|(~m[124]&m[288]&m[654]))&~BiasedRNG[559])|((~m[124]&~m[288]&m[654])|(m[124]&~m[288]&m[654])|(m[124]&m[288]&m[654]));
    m[459] = (((~m[124]&~m[302]&~m[655])|(m[124]&m[302]&~m[655]))&BiasedRNG[560])|(((m[124]&~m[302]&~m[655])|(~m[124]&m[302]&m[655]))&~BiasedRNG[560])|((~m[124]&~m[302]&m[655])|(m[124]&~m[302]&m[655])|(m[124]&m[302]&m[655]));
    m[460] = (((~m[124]&~m[316]&~m[656])|(m[124]&m[316]&~m[656]))&BiasedRNG[561])|(((m[124]&~m[316]&~m[656])|(~m[124]&m[316]&m[656]))&~BiasedRNG[561])|((~m[124]&~m[316]&m[656])|(m[124]&~m[316]&m[656])|(m[124]&m[316]&m[656]));
    m[461] = (((~m[124]&~m[330]&~m[657])|(m[124]&m[330]&~m[657]))&BiasedRNG[562])|(((m[124]&~m[330]&~m[657])|(~m[124]&m[330]&m[657]))&~BiasedRNG[562])|((~m[124]&~m[330]&m[657])|(m[124]&~m[330]&m[657])|(m[124]&m[330]&m[657]));
    m[468] = (((~m[126]&~m[233]&~m[664])|(m[126]&m[233]&~m[664]))&BiasedRNG[563])|(((m[126]&~m[233]&~m[664])|(~m[126]&m[233]&m[664]))&~BiasedRNG[563])|((~m[126]&~m[233]&m[664])|(m[126]&~m[233]&m[664])|(m[126]&m[233]&m[664]));
    m[469] = (((~m[126]&~m[247]&~m[665])|(m[126]&m[247]&~m[665]))&BiasedRNG[564])|(((m[126]&~m[247]&~m[665])|(~m[126]&m[247]&m[665]))&~BiasedRNG[564])|((~m[126]&~m[247]&m[665])|(m[126]&~m[247]&m[665])|(m[126]&m[247]&m[665]));
    m[470] = (((~m[126]&~m[261]&~m[666])|(m[126]&m[261]&~m[666]))&BiasedRNG[565])|(((m[126]&~m[261]&~m[666])|(~m[126]&m[261]&m[666]))&~BiasedRNG[565])|((~m[126]&~m[261]&m[666])|(m[126]&~m[261]&m[666])|(m[126]&m[261]&m[666]));
    m[471] = (((~m[126]&~m[275]&~m[667])|(m[126]&m[275]&~m[667]))&BiasedRNG[566])|(((m[126]&~m[275]&~m[667])|(~m[126]&m[275]&m[667]))&~BiasedRNG[566])|((~m[126]&~m[275]&m[667])|(m[126]&~m[275]&m[667])|(m[126]&m[275]&m[667]));
    m[472] = (((~m[127]&~m[289]&~m[668])|(m[127]&m[289]&~m[668]))&BiasedRNG[567])|(((m[127]&~m[289]&~m[668])|(~m[127]&m[289]&m[668]))&~BiasedRNG[567])|((~m[127]&~m[289]&m[668])|(m[127]&~m[289]&m[668])|(m[127]&m[289]&m[668]));
    m[473] = (((~m[127]&~m[303]&~m[669])|(m[127]&m[303]&~m[669]))&BiasedRNG[568])|(((m[127]&~m[303]&~m[669])|(~m[127]&m[303]&m[669]))&~BiasedRNG[568])|((~m[127]&~m[303]&m[669])|(m[127]&~m[303]&m[669])|(m[127]&m[303]&m[669]));
    m[474] = (((~m[127]&~m[317]&~m[670])|(m[127]&m[317]&~m[670]))&BiasedRNG[569])|(((m[127]&~m[317]&~m[670])|(~m[127]&m[317]&m[670]))&~BiasedRNG[569])|((~m[127]&~m[317]&m[670])|(m[127]&~m[317]&m[670])|(m[127]&m[317]&m[670]));
    m[475] = (((~m[127]&~m[331]&~m[671])|(m[127]&m[331]&~m[671]))&BiasedRNG[570])|(((m[127]&~m[331]&~m[671])|(~m[127]&m[331]&m[671]))&~BiasedRNG[570])|((~m[127]&~m[331]&m[671])|(m[127]&~m[331]&m[671])|(m[127]&m[331]&m[671]));
    m[482] = (((~m[129]&~m[234]&~m[678])|(m[129]&m[234]&~m[678]))&BiasedRNG[571])|(((m[129]&~m[234]&~m[678])|(~m[129]&m[234]&m[678]))&~BiasedRNG[571])|((~m[129]&~m[234]&m[678])|(m[129]&~m[234]&m[678])|(m[129]&m[234]&m[678]));
    m[483] = (((~m[129]&~m[248]&~m[679])|(m[129]&m[248]&~m[679]))&BiasedRNG[572])|(((m[129]&~m[248]&~m[679])|(~m[129]&m[248]&m[679]))&~BiasedRNG[572])|((~m[129]&~m[248]&m[679])|(m[129]&~m[248]&m[679])|(m[129]&m[248]&m[679]));
    m[484] = (((~m[129]&~m[262]&~m[680])|(m[129]&m[262]&~m[680]))&BiasedRNG[573])|(((m[129]&~m[262]&~m[680])|(~m[129]&m[262]&m[680]))&~BiasedRNG[573])|((~m[129]&~m[262]&m[680])|(m[129]&~m[262]&m[680])|(m[129]&m[262]&m[680]));
    m[485] = (((~m[129]&~m[276]&~m[681])|(m[129]&m[276]&~m[681]))&BiasedRNG[574])|(((m[129]&~m[276]&~m[681])|(~m[129]&m[276]&m[681]))&~BiasedRNG[574])|((~m[129]&~m[276]&m[681])|(m[129]&~m[276]&m[681])|(m[129]&m[276]&m[681]));
    m[486] = (((~m[130]&~m[290]&~m[682])|(m[130]&m[290]&~m[682]))&BiasedRNG[575])|(((m[130]&~m[290]&~m[682])|(~m[130]&m[290]&m[682]))&~BiasedRNG[575])|((~m[130]&~m[290]&m[682])|(m[130]&~m[290]&m[682])|(m[130]&m[290]&m[682]));
    m[487] = (((~m[130]&~m[304]&~m[683])|(m[130]&m[304]&~m[683]))&BiasedRNG[576])|(((m[130]&~m[304]&~m[683])|(~m[130]&m[304]&m[683]))&~BiasedRNG[576])|((~m[130]&~m[304]&m[683])|(m[130]&~m[304]&m[683])|(m[130]&m[304]&m[683]));
    m[488] = (((~m[130]&~m[318]&~m[684])|(m[130]&m[318]&~m[684]))&BiasedRNG[577])|(((m[130]&~m[318]&~m[684])|(~m[130]&m[318]&m[684]))&~BiasedRNG[577])|((~m[130]&~m[318]&m[684])|(m[130]&~m[318]&m[684])|(m[130]&m[318]&m[684]));
    m[489] = (((~m[130]&~m[332]&~m[685])|(m[130]&m[332]&~m[685]))&BiasedRNG[578])|(((m[130]&~m[332]&~m[685])|(~m[130]&m[332]&m[685]))&~BiasedRNG[578])|((~m[130]&~m[332]&m[685])|(m[130]&~m[332]&m[685])|(m[130]&m[332]&m[685]));
    m[496] = (((~m[132]&~m[235]&~m[692])|(m[132]&m[235]&~m[692]))&BiasedRNG[579])|(((m[132]&~m[235]&~m[692])|(~m[132]&m[235]&m[692]))&~BiasedRNG[579])|((~m[132]&~m[235]&m[692])|(m[132]&~m[235]&m[692])|(m[132]&m[235]&m[692]));
    m[497] = (((~m[132]&~m[249]&~m[693])|(m[132]&m[249]&~m[693]))&BiasedRNG[580])|(((m[132]&~m[249]&~m[693])|(~m[132]&m[249]&m[693]))&~BiasedRNG[580])|((~m[132]&~m[249]&m[693])|(m[132]&~m[249]&m[693])|(m[132]&m[249]&m[693]));
    m[498] = (((~m[132]&~m[263]&~m[694])|(m[132]&m[263]&~m[694]))&BiasedRNG[581])|(((m[132]&~m[263]&~m[694])|(~m[132]&m[263]&m[694]))&~BiasedRNG[581])|((~m[132]&~m[263]&m[694])|(m[132]&~m[263]&m[694])|(m[132]&m[263]&m[694]));
    m[499] = (((~m[132]&~m[277]&~m[695])|(m[132]&m[277]&~m[695]))&BiasedRNG[582])|(((m[132]&~m[277]&~m[695])|(~m[132]&m[277]&m[695]))&~BiasedRNG[582])|((~m[132]&~m[277]&m[695])|(m[132]&~m[277]&m[695])|(m[132]&m[277]&m[695]));
    m[500] = (((~m[133]&~m[291]&~m[696])|(m[133]&m[291]&~m[696]))&BiasedRNG[583])|(((m[133]&~m[291]&~m[696])|(~m[133]&m[291]&m[696]))&~BiasedRNG[583])|((~m[133]&~m[291]&m[696])|(m[133]&~m[291]&m[696])|(m[133]&m[291]&m[696]));
    m[501] = (((~m[133]&~m[305]&~m[697])|(m[133]&m[305]&~m[697]))&BiasedRNG[584])|(((m[133]&~m[305]&~m[697])|(~m[133]&m[305]&m[697]))&~BiasedRNG[584])|((~m[133]&~m[305]&m[697])|(m[133]&~m[305]&m[697])|(m[133]&m[305]&m[697]));
    m[502] = (((~m[133]&~m[319]&~m[698])|(m[133]&m[319]&~m[698]))&BiasedRNG[585])|(((m[133]&~m[319]&~m[698])|(~m[133]&m[319]&m[698]))&~BiasedRNG[585])|((~m[133]&~m[319]&m[698])|(m[133]&~m[319]&m[698])|(m[133]&m[319]&m[698]));
    m[503] = (((~m[133]&~m[333]&~m[699])|(m[133]&m[333]&~m[699]))&BiasedRNG[586])|(((m[133]&~m[333]&~m[699])|(~m[133]&m[333]&m[699]))&~BiasedRNG[586])|((~m[133]&~m[333]&m[699])|(m[133]&~m[333]&m[699])|(m[133]&m[333]&m[699]));
    m[510] = (((~m[135]&~m[236]&~m[706])|(m[135]&m[236]&~m[706]))&BiasedRNG[587])|(((m[135]&~m[236]&~m[706])|(~m[135]&m[236]&m[706]))&~BiasedRNG[587])|((~m[135]&~m[236]&m[706])|(m[135]&~m[236]&m[706])|(m[135]&m[236]&m[706]));
    m[511] = (((~m[135]&~m[250]&~m[707])|(m[135]&m[250]&~m[707]))&BiasedRNG[588])|(((m[135]&~m[250]&~m[707])|(~m[135]&m[250]&m[707]))&~BiasedRNG[588])|((~m[135]&~m[250]&m[707])|(m[135]&~m[250]&m[707])|(m[135]&m[250]&m[707]));
    m[512] = (((~m[135]&~m[264]&~m[708])|(m[135]&m[264]&~m[708]))&BiasedRNG[589])|(((m[135]&~m[264]&~m[708])|(~m[135]&m[264]&m[708]))&~BiasedRNG[589])|((~m[135]&~m[264]&m[708])|(m[135]&~m[264]&m[708])|(m[135]&m[264]&m[708]));
    m[513] = (((~m[135]&~m[278]&~m[709])|(m[135]&m[278]&~m[709]))&BiasedRNG[590])|(((m[135]&~m[278]&~m[709])|(~m[135]&m[278]&m[709]))&~BiasedRNG[590])|((~m[135]&~m[278]&m[709])|(m[135]&~m[278]&m[709])|(m[135]&m[278]&m[709]));
    m[514] = (((~m[136]&~m[292]&~m[710])|(m[136]&m[292]&~m[710]))&BiasedRNG[591])|(((m[136]&~m[292]&~m[710])|(~m[136]&m[292]&m[710]))&~BiasedRNG[591])|((~m[136]&~m[292]&m[710])|(m[136]&~m[292]&m[710])|(m[136]&m[292]&m[710]));
    m[515] = (((~m[136]&~m[306]&~m[711])|(m[136]&m[306]&~m[711]))&BiasedRNG[592])|(((m[136]&~m[306]&~m[711])|(~m[136]&m[306]&m[711]))&~BiasedRNG[592])|((~m[136]&~m[306]&m[711])|(m[136]&~m[306]&m[711])|(m[136]&m[306]&m[711]));
    m[516] = (((~m[136]&~m[320]&~m[712])|(m[136]&m[320]&~m[712]))&BiasedRNG[593])|(((m[136]&~m[320]&~m[712])|(~m[136]&m[320]&m[712]))&~BiasedRNG[593])|((~m[136]&~m[320]&m[712])|(m[136]&~m[320]&m[712])|(m[136]&m[320]&m[712]));
    m[517] = (((~m[136]&~m[334]&~m[713])|(m[136]&m[334]&~m[713]))&BiasedRNG[594])|(((m[136]&~m[334]&~m[713])|(~m[136]&m[334]&m[713]))&~BiasedRNG[594])|((~m[136]&~m[334]&m[713])|(m[136]&~m[334]&m[713])|(m[136]&m[334]&m[713]));
    m[524] = (((~m[138]&~m[237]&~m[720])|(m[138]&m[237]&~m[720]))&BiasedRNG[595])|(((m[138]&~m[237]&~m[720])|(~m[138]&m[237]&m[720]))&~BiasedRNG[595])|((~m[138]&~m[237]&m[720])|(m[138]&~m[237]&m[720])|(m[138]&m[237]&m[720]));
    m[525] = (((~m[138]&~m[251]&~m[721])|(m[138]&m[251]&~m[721]))&BiasedRNG[596])|(((m[138]&~m[251]&~m[721])|(~m[138]&m[251]&m[721]))&~BiasedRNG[596])|((~m[138]&~m[251]&m[721])|(m[138]&~m[251]&m[721])|(m[138]&m[251]&m[721]));
    m[526] = (((~m[138]&~m[265]&~m[722])|(m[138]&m[265]&~m[722]))&BiasedRNG[597])|(((m[138]&~m[265]&~m[722])|(~m[138]&m[265]&m[722]))&~BiasedRNG[597])|((~m[138]&~m[265]&m[722])|(m[138]&~m[265]&m[722])|(m[138]&m[265]&m[722]));
    m[527] = (((~m[138]&~m[279]&~m[723])|(m[138]&m[279]&~m[723]))&BiasedRNG[598])|(((m[138]&~m[279]&~m[723])|(~m[138]&m[279]&m[723]))&~BiasedRNG[598])|((~m[138]&~m[279]&m[723])|(m[138]&~m[279]&m[723])|(m[138]&m[279]&m[723]));
    m[528] = (((~m[139]&~m[293]&~m[724])|(m[139]&m[293]&~m[724]))&BiasedRNG[599])|(((m[139]&~m[293]&~m[724])|(~m[139]&m[293]&m[724]))&~BiasedRNG[599])|((~m[139]&~m[293]&m[724])|(m[139]&~m[293]&m[724])|(m[139]&m[293]&m[724]));
    m[529] = (((~m[139]&~m[307]&~m[725])|(m[139]&m[307]&~m[725]))&BiasedRNG[600])|(((m[139]&~m[307]&~m[725])|(~m[139]&m[307]&m[725]))&~BiasedRNG[600])|((~m[139]&~m[307]&m[725])|(m[139]&~m[307]&m[725])|(m[139]&m[307]&m[725]));
    m[530] = (((~m[139]&~m[321]&~m[726])|(m[139]&m[321]&~m[726]))&BiasedRNG[601])|(((m[139]&~m[321]&~m[726])|(~m[139]&m[321]&m[726]))&~BiasedRNG[601])|((~m[139]&~m[321]&m[726])|(m[139]&~m[321]&m[726])|(m[139]&m[321]&m[726]));
    m[531] = (((~m[139]&~m[335]&~m[727])|(m[139]&m[335]&~m[727]))&BiasedRNG[602])|(((m[139]&~m[335]&~m[727])|(~m[139]&m[335]&m[727]))&~BiasedRNG[602])|((~m[139]&~m[335]&m[727])|(m[139]&~m[335]&m[727])|(m[139]&m[335]&m[727]));
    m[538] = (((m[224]&~m[342]&m[803])|(~m[224]&m[342]&m[803]))&BiasedRNG[603])|(((m[224]&m[342]&~m[803]))&~BiasedRNG[603])|((m[224]&m[342]&m[803]));
    m[539] = (((m[238]&~m[343]&m[833])|(~m[238]&m[343]&m[833]))&BiasedRNG[604])|(((m[238]&m[343]&~m[833]))&~BiasedRNG[604])|((m[238]&m[343]&m[833]));
    m[540] = (((m[252]&~m[344]&m[868])|(~m[252]&m[344]&m[868]))&BiasedRNG[605])|(((m[252]&m[344]&~m[868]))&~BiasedRNG[605])|((m[252]&m[344]&m[868]));
    m[541] = (((m[266]&~m[345]&m[908])|(~m[266]&m[345]&m[908]))&BiasedRNG[606])|(((m[266]&m[345]&~m[908]))&~BiasedRNG[606])|((m[266]&m[345]&m[908]));
    m[542] = (((m[280]&~m[346]&m[953])|(~m[280]&m[346]&m[953]))&BiasedRNG[607])|(((m[280]&m[346]&~m[953]))&~BiasedRNG[607])|((m[280]&m[346]&m[953]));
    m[543] = (((m[294]&~m[347]&m[1003])|(~m[294]&m[347]&m[1003]))&BiasedRNG[608])|(((m[294]&m[347]&~m[1003]))&~BiasedRNG[608])|((m[294]&m[347]&m[1003]));
    m[544] = (((m[308]&~m[348]&m[1058])|(~m[308]&m[348]&m[1058]))&BiasedRNG[609])|(((m[308]&m[348]&~m[1058]))&~BiasedRNG[609])|((m[308]&m[348]&m[1058]));
    m[545] = (((m[322]&~m[349]&m[1118])|(~m[322]&m[349]&m[1118]))&BiasedRNG[610])|(((m[322]&m[349]&~m[1118]))&~BiasedRNG[610])|((m[322]&m[349]&m[1118]));
    m[552] = (((m[225]&~m[356]&m[834])|(~m[225]&m[356]&m[834]))&BiasedRNG[611])|(((m[225]&m[356]&~m[834]))&~BiasedRNG[611])|((m[225]&m[356]&m[834]));
    m[553] = (((m[239]&~m[357]&m[869])|(~m[239]&m[357]&m[869]))&BiasedRNG[612])|(((m[239]&m[357]&~m[869]))&~BiasedRNG[612])|((m[239]&m[357]&m[869]));
    m[554] = (((m[253]&~m[358]&m[909])|(~m[253]&m[358]&m[909]))&BiasedRNG[613])|(((m[253]&m[358]&~m[909]))&~BiasedRNG[613])|((m[253]&m[358]&m[909]));
    m[555] = (((m[267]&~m[359]&m[954])|(~m[267]&m[359]&m[954]))&BiasedRNG[614])|(((m[267]&m[359]&~m[954]))&~BiasedRNG[614])|((m[267]&m[359]&m[954]));
    m[556] = (((m[281]&~m[360]&m[1004])|(~m[281]&m[360]&m[1004]))&BiasedRNG[615])|(((m[281]&m[360]&~m[1004]))&~BiasedRNG[615])|((m[281]&m[360]&m[1004]));
    m[557] = (((m[295]&~m[361]&m[1059])|(~m[295]&m[361]&m[1059]))&BiasedRNG[616])|(((m[295]&m[361]&~m[1059]))&~BiasedRNG[616])|((m[295]&m[361]&m[1059]));
    m[558] = (((m[309]&~m[362]&m[1119])|(~m[309]&m[362]&m[1119]))&BiasedRNG[617])|(((m[309]&m[362]&~m[1119]))&~BiasedRNG[617])|((m[309]&m[362]&m[1119]));
    m[559] = (((m[323]&~m[363]&m[1184])|(~m[323]&m[363]&m[1184]))&BiasedRNG[618])|(((m[323]&m[363]&~m[1184]))&~BiasedRNG[618])|((m[323]&m[363]&m[1184]));
    m[566] = (((m[226]&~m[370]&m[874])|(~m[226]&m[370]&m[874]))&BiasedRNG[619])|(((m[226]&m[370]&~m[874]))&~BiasedRNG[619])|((m[226]&m[370]&m[874]));
    m[567] = (((m[240]&~m[371]&m[914])|(~m[240]&m[371]&m[914]))&BiasedRNG[620])|(((m[240]&m[371]&~m[914]))&~BiasedRNG[620])|((m[240]&m[371]&m[914]));
    m[568] = (((m[254]&~m[372]&m[959])|(~m[254]&m[372]&m[959]))&BiasedRNG[621])|(((m[254]&m[372]&~m[959]))&~BiasedRNG[621])|((m[254]&m[372]&m[959]));
    m[569] = (((m[268]&~m[373]&m[1009])|(~m[268]&m[373]&m[1009]))&BiasedRNG[622])|(((m[268]&m[373]&~m[1009]))&~BiasedRNG[622])|((m[268]&m[373]&m[1009]));
    m[570] = (((m[282]&~m[374]&m[1064])|(~m[282]&m[374]&m[1064]))&BiasedRNG[623])|(((m[282]&m[374]&~m[1064]))&~BiasedRNG[623])|((m[282]&m[374]&m[1064]));
    m[571] = (((m[296]&~m[375]&m[1124])|(~m[296]&m[375]&m[1124]))&BiasedRNG[624])|(((m[296]&m[375]&~m[1124]))&~BiasedRNG[624])|((m[296]&m[375]&m[1124]));
    m[572] = (((m[310]&~m[376]&m[1189])|(~m[310]&m[376]&m[1189]))&BiasedRNG[625])|(((m[310]&m[376]&~m[1189]))&~BiasedRNG[625])|((m[310]&m[376]&m[1189]));
    m[573] = (((m[324]&~m[377]&m[1249])|(~m[324]&m[377]&m[1249]))&BiasedRNG[626])|(((m[324]&m[377]&~m[1249]))&~BiasedRNG[626])|((m[324]&m[377]&m[1249]));
    m[580] = (((m[227]&~m[384]&m[919])|(~m[227]&m[384]&m[919]))&BiasedRNG[627])|(((m[227]&m[384]&~m[919]))&~BiasedRNG[627])|((m[227]&m[384]&m[919]));
    m[581] = (((m[241]&~m[385]&m[964])|(~m[241]&m[385]&m[964]))&BiasedRNG[628])|(((m[241]&m[385]&~m[964]))&~BiasedRNG[628])|((m[241]&m[385]&m[964]));
    m[582] = (((m[255]&~m[386]&m[1014])|(~m[255]&m[386]&m[1014]))&BiasedRNG[629])|(((m[255]&m[386]&~m[1014]))&~BiasedRNG[629])|((m[255]&m[386]&m[1014]));
    m[583] = (((m[269]&~m[387]&m[1069])|(~m[269]&m[387]&m[1069]))&BiasedRNG[630])|(((m[269]&m[387]&~m[1069]))&~BiasedRNG[630])|((m[269]&m[387]&m[1069]));
    m[584] = (((m[283]&~m[388]&m[1129])|(~m[283]&m[388]&m[1129]))&BiasedRNG[631])|(((m[283]&m[388]&~m[1129]))&~BiasedRNG[631])|((m[283]&m[388]&m[1129]));
    m[585] = (((m[297]&~m[389]&m[1194])|(~m[297]&m[389]&m[1194]))&BiasedRNG[632])|(((m[297]&m[389]&~m[1194]))&~BiasedRNG[632])|((m[297]&m[389]&m[1194]));
    m[586] = (((m[311]&~m[390]&m[1254])|(~m[311]&m[390]&m[1254]))&BiasedRNG[633])|(((m[311]&m[390]&~m[1254]))&~BiasedRNG[633])|((m[311]&m[390]&m[1254]));
    m[587] = (((m[325]&~m[391]&m[1309])|(~m[325]&m[391]&m[1309]))&BiasedRNG[634])|(((m[325]&m[391]&~m[1309]))&~BiasedRNG[634])|((m[325]&m[391]&m[1309]));
    m[594] = (((m[228]&~m[398]&m[969])|(~m[228]&m[398]&m[969]))&BiasedRNG[635])|(((m[228]&m[398]&~m[969]))&~BiasedRNG[635])|((m[228]&m[398]&m[969]));
    m[595] = (((m[242]&~m[399]&m[1019])|(~m[242]&m[399]&m[1019]))&BiasedRNG[636])|(((m[242]&m[399]&~m[1019]))&~BiasedRNG[636])|((m[242]&m[399]&m[1019]));
    m[596] = (((m[256]&~m[400]&m[1074])|(~m[256]&m[400]&m[1074]))&BiasedRNG[637])|(((m[256]&m[400]&~m[1074]))&~BiasedRNG[637])|((m[256]&m[400]&m[1074]));
    m[597] = (((m[270]&~m[401]&m[1134])|(~m[270]&m[401]&m[1134]))&BiasedRNG[638])|(((m[270]&m[401]&~m[1134]))&~BiasedRNG[638])|((m[270]&m[401]&m[1134]));
    m[598] = (((m[284]&~m[402]&m[1199])|(~m[284]&m[402]&m[1199]))&BiasedRNG[639])|(((m[284]&m[402]&~m[1199]))&~BiasedRNG[639])|((m[284]&m[402]&m[1199]));
    m[599] = (((m[298]&~m[403]&m[1259])|(~m[298]&m[403]&m[1259]))&BiasedRNG[640])|(((m[298]&m[403]&~m[1259]))&~BiasedRNG[640])|((m[298]&m[403]&m[1259]));
    m[600] = (((m[312]&~m[404]&m[1314])|(~m[312]&m[404]&m[1314]))&BiasedRNG[641])|(((m[312]&m[404]&~m[1314]))&~BiasedRNG[641])|((m[312]&m[404]&m[1314]));
    m[601] = (((m[326]&~m[405]&m[1364])|(~m[326]&m[405]&m[1364]))&BiasedRNG[642])|(((m[326]&m[405]&~m[1364]))&~BiasedRNG[642])|((m[326]&m[405]&m[1364]));
    m[608] = (((m[229]&~m[412]&m[1024])|(~m[229]&m[412]&m[1024]))&BiasedRNG[643])|(((m[229]&m[412]&~m[1024]))&~BiasedRNG[643])|((m[229]&m[412]&m[1024]));
    m[609] = (((m[243]&~m[413]&m[1079])|(~m[243]&m[413]&m[1079]))&BiasedRNG[644])|(((m[243]&m[413]&~m[1079]))&~BiasedRNG[644])|((m[243]&m[413]&m[1079]));
    m[610] = (((m[257]&~m[414]&m[1139])|(~m[257]&m[414]&m[1139]))&BiasedRNG[645])|(((m[257]&m[414]&~m[1139]))&~BiasedRNG[645])|((m[257]&m[414]&m[1139]));
    m[611] = (((m[271]&~m[415]&m[1204])|(~m[271]&m[415]&m[1204]))&BiasedRNG[646])|(((m[271]&m[415]&~m[1204]))&~BiasedRNG[646])|((m[271]&m[415]&m[1204]));
    m[612] = (((m[285]&~m[416]&m[1264])|(~m[285]&m[416]&m[1264]))&BiasedRNG[647])|(((m[285]&m[416]&~m[1264]))&~BiasedRNG[647])|((m[285]&m[416]&m[1264]));
    m[613] = (((m[299]&~m[417]&m[1319])|(~m[299]&m[417]&m[1319]))&BiasedRNG[648])|(((m[299]&m[417]&~m[1319]))&~BiasedRNG[648])|((m[299]&m[417]&m[1319]));
    m[614] = (((m[313]&~m[418]&m[1369])|(~m[313]&m[418]&m[1369]))&BiasedRNG[649])|(((m[313]&m[418]&~m[1369]))&~BiasedRNG[649])|((m[313]&m[418]&m[1369]));
    m[615] = (((m[327]&~m[419]&m[1414])|(~m[327]&m[419]&m[1414]))&BiasedRNG[650])|(((m[327]&m[419]&~m[1414]))&~BiasedRNG[650])|((m[327]&m[419]&m[1414]));
    m[616] = (((m[146]&~m[420]&m[829])|(~m[146]&m[420]&m[829]))&BiasedRNG[651])|(((m[146]&m[420]&~m[829]))&~BiasedRNG[651])|((m[146]&m[420]&m[829]));
    m[617] = (((m[160]&~m[421]&m[859])|(~m[160]&m[421]&m[859]))&BiasedRNG[652])|(((m[160]&m[421]&~m[859]))&~BiasedRNG[652])|((m[160]&m[421]&m[859]));
    m[618] = (((m[174]&~m[422]&m[894])|(~m[174]&m[422]&m[894]))&BiasedRNG[653])|(((m[174]&m[422]&~m[894]))&~BiasedRNG[653])|((m[174]&m[422]&m[894]));
    m[619] = (((m[188]&~m[423]&m[934])|(~m[188]&m[423]&m[934]))&BiasedRNG[654])|(((m[188]&m[423]&~m[934]))&~BiasedRNG[654])|((m[188]&m[423]&m[934]));
    m[620] = (((m[202]&~m[424]&m[979])|(~m[202]&m[424]&m[979]))&BiasedRNG[655])|(((m[202]&m[424]&~m[979]))&~BiasedRNG[655])|((m[202]&m[424]&m[979]));
    m[621] = (((m[216]&~m[425]&m[1029])|(~m[216]&m[425]&m[1029]))&BiasedRNG[656])|(((m[216]&m[425]&~m[1029]))&~BiasedRNG[656])|((m[216]&m[425]&m[1029]));
    m[630] = (((m[147]&~m[434]&m[864])|(~m[147]&m[434]&m[864]))&BiasedRNG[657])|(((m[147]&m[434]&~m[864]))&~BiasedRNG[657])|((m[147]&m[434]&m[864]));
    m[631] = (((m[161]&~m[435]&m[899])|(~m[161]&m[435]&m[899]))&BiasedRNG[658])|(((m[161]&m[435]&~m[899]))&~BiasedRNG[658])|((m[161]&m[435]&m[899]));
    m[632] = (((m[175]&~m[436]&m[939])|(~m[175]&m[436]&m[939]))&BiasedRNG[659])|(((m[175]&m[436]&~m[939]))&~BiasedRNG[659])|((m[175]&m[436]&m[939]));
    m[633] = (((m[189]&~m[437]&m[984])|(~m[189]&m[437]&m[984]))&BiasedRNG[660])|(((m[189]&m[437]&~m[984]))&~BiasedRNG[660])|((m[189]&m[437]&m[984]));
    m[634] = (((m[203]&~m[438]&m[1034])|(~m[203]&m[438]&m[1034]))&BiasedRNG[661])|(((m[203]&m[438]&~m[1034]))&~BiasedRNG[661])|((m[203]&m[438]&m[1034]));
    m[635] = (((m[217]&~m[439]&m[1089])|(~m[217]&m[439]&m[1089]))&BiasedRNG[662])|(((m[217]&m[439]&~m[1089]))&~BiasedRNG[662])|((m[217]&m[439]&m[1089]));
    m[644] = (((m[148]&~m[448]&m[904])|(~m[148]&m[448]&m[904]))&BiasedRNG[663])|(((m[148]&m[448]&~m[904]))&~BiasedRNG[663])|((m[148]&m[448]&m[904]));
    m[645] = (((m[162]&~m[449]&m[944])|(~m[162]&m[449]&m[944]))&BiasedRNG[664])|(((m[162]&m[449]&~m[944]))&~BiasedRNG[664])|((m[162]&m[449]&m[944]));
    m[646] = (((m[176]&~m[450]&m[989])|(~m[176]&m[450]&m[989]))&BiasedRNG[665])|(((m[176]&m[450]&~m[989]))&~BiasedRNG[665])|((m[176]&m[450]&m[989]));
    m[647] = (((m[190]&~m[451]&m[1039])|(~m[190]&m[451]&m[1039]))&BiasedRNG[666])|(((m[190]&m[451]&~m[1039]))&~BiasedRNG[666])|((m[190]&m[451]&m[1039]));
    m[648] = (((m[204]&~m[452]&m[1094])|(~m[204]&m[452]&m[1094]))&BiasedRNG[667])|(((m[204]&m[452]&~m[1094]))&~BiasedRNG[667])|((m[204]&m[452]&m[1094]));
    m[649] = (((m[218]&~m[453]&m[1154])|(~m[218]&m[453]&m[1154]))&BiasedRNG[668])|(((m[218]&m[453]&~m[1154]))&~BiasedRNG[668])|((m[218]&m[453]&m[1154]));
    m[658] = (((m[149]&~m[462]&m[949])|(~m[149]&m[462]&m[949]))&BiasedRNG[669])|(((m[149]&m[462]&~m[949]))&~BiasedRNG[669])|((m[149]&m[462]&m[949]));
    m[659] = (((m[163]&~m[463]&m[994])|(~m[163]&m[463]&m[994]))&BiasedRNG[670])|(((m[163]&m[463]&~m[994]))&~BiasedRNG[670])|((m[163]&m[463]&m[994]));
    m[660] = (((m[177]&~m[464]&m[1044])|(~m[177]&m[464]&m[1044]))&BiasedRNG[671])|(((m[177]&m[464]&~m[1044]))&~BiasedRNG[671])|((m[177]&m[464]&m[1044]));
    m[661] = (((m[191]&~m[465]&m[1099])|(~m[191]&m[465]&m[1099]))&BiasedRNG[672])|(((m[191]&m[465]&~m[1099]))&~BiasedRNG[672])|((m[191]&m[465]&m[1099]));
    m[662] = (((m[205]&~m[466]&m[1159])|(~m[205]&m[466]&m[1159]))&BiasedRNG[673])|(((m[205]&m[466]&~m[1159]))&~BiasedRNG[673])|((m[205]&m[466]&m[1159]));
    m[663] = (((m[219]&~m[467]&m[1224])|(~m[219]&m[467]&m[1224]))&BiasedRNG[674])|(((m[219]&m[467]&~m[1224]))&~BiasedRNG[674])|((m[219]&m[467]&m[1224]));
    m[672] = (((m[150]&~m[476]&m[999])|(~m[150]&m[476]&m[999]))&BiasedRNG[675])|(((m[150]&m[476]&~m[999]))&~BiasedRNG[675])|((m[150]&m[476]&m[999]));
    m[673] = (((m[164]&~m[477]&m[1049])|(~m[164]&m[477]&m[1049]))&BiasedRNG[676])|(((m[164]&m[477]&~m[1049]))&~BiasedRNG[676])|((m[164]&m[477]&m[1049]));
    m[674] = (((m[178]&~m[478]&m[1104])|(~m[178]&m[478]&m[1104]))&BiasedRNG[677])|(((m[178]&m[478]&~m[1104]))&~BiasedRNG[677])|((m[178]&m[478]&m[1104]));
    m[675] = (((m[192]&~m[479]&m[1164])|(~m[192]&m[479]&m[1164]))&BiasedRNG[678])|(((m[192]&m[479]&~m[1164]))&~BiasedRNG[678])|((m[192]&m[479]&m[1164]));
    m[676] = (((m[206]&~m[480]&m[1229])|(~m[206]&m[480]&m[1229]))&BiasedRNG[679])|(((m[206]&m[480]&~m[1229]))&~BiasedRNG[679])|((m[206]&m[480]&m[1229]));
    m[677] = (((m[220]&~m[481]&m[1289])|(~m[220]&m[481]&m[1289]))&BiasedRNG[680])|(((m[220]&m[481]&~m[1289]))&~BiasedRNG[680])|((m[220]&m[481]&m[1289]));
    m[686] = (((m[151]&~m[490]&m[1054])|(~m[151]&m[490]&m[1054]))&BiasedRNG[681])|(((m[151]&m[490]&~m[1054]))&~BiasedRNG[681])|((m[151]&m[490]&m[1054]));
    m[687] = (((m[165]&~m[491]&m[1109])|(~m[165]&m[491]&m[1109]))&BiasedRNG[682])|(((m[165]&m[491]&~m[1109]))&~BiasedRNG[682])|((m[165]&m[491]&m[1109]));
    m[688] = (((m[179]&~m[492]&m[1169])|(~m[179]&m[492]&m[1169]))&BiasedRNG[683])|(((m[179]&m[492]&~m[1169]))&~BiasedRNG[683])|((m[179]&m[492]&m[1169]));
    m[689] = (((m[193]&~m[493]&m[1234])|(~m[193]&m[493]&m[1234]))&BiasedRNG[684])|(((m[193]&m[493]&~m[1234]))&~BiasedRNG[684])|((m[193]&m[493]&m[1234]));
    m[690] = (((m[207]&~m[494]&m[1294])|(~m[207]&m[494]&m[1294]))&BiasedRNG[685])|(((m[207]&m[494]&~m[1294]))&~BiasedRNG[685])|((m[207]&m[494]&m[1294]));
    m[691] = (((m[221]&~m[495]&m[1349])|(~m[221]&m[495]&m[1349]))&BiasedRNG[686])|(((m[221]&m[495]&~m[1349]))&~BiasedRNG[686])|((m[221]&m[495]&m[1349]));
    m[700] = (((m[152]&~m[504]&m[1114])|(~m[152]&m[504]&m[1114]))&BiasedRNG[687])|(((m[152]&m[504]&~m[1114]))&~BiasedRNG[687])|((m[152]&m[504]&m[1114]));
    m[701] = (((m[166]&~m[505]&m[1174])|(~m[166]&m[505]&m[1174]))&BiasedRNG[688])|(((m[166]&m[505]&~m[1174]))&~BiasedRNG[688])|((m[166]&m[505]&m[1174]));
    m[702] = (((m[180]&~m[506]&m[1239])|(~m[180]&m[506]&m[1239]))&BiasedRNG[689])|(((m[180]&m[506]&~m[1239]))&~BiasedRNG[689])|((m[180]&m[506]&m[1239]));
    m[703] = (((m[194]&~m[507]&m[1299])|(~m[194]&m[507]&m[1299]))&BiasedRNG[690])|(((m[194]&m[507]&~m[1299]))&~BiasedRNG[690])|((m[194]&m[507]&m[1299]));
    m[704] = (((m[208]&~m[508]&m[1354])|(~m[208]&m[508]&m[1354]))&BiasedRNG[691])|(((m[208]&m[508]&~m[1354]))&~BiasedRNG[691])|((m[208]&m[508]&m[1354]));
    m[705] = (((m[222]&~m[509]&m[1404])|(~m[222]&m[509]&m[1404]))&BiasedRNG[692])|(((m[222]&m[509]&~m[1404]))&~BiasedRNG[692])|((m[222]&m[509]&m[1404]));
    m[714] = (((m[153]&~m[518]&m[1179])|(~m[153]&m[518]&m[1179]))&BiasedRNG[693])|(((m[153]&m[518]&~m[1179]))&~BiasedRNG[693])|((m[153]&m[518]&m[1179]));
    m[715] = (((m[167]&~m[519]&m[1244])|(~m[167]&m[519]&m[1244]))&BiasedRNG[694])|(((m[167]&m[519]&~m[1244]))&~BiasedRNG[694])|((m[167]&m[519]&m[1244]));
    m[716] = (((m[181]&~m[520]&m[1304])|(~m[181]&m[520]&m[1304]))&BiasedRNG[695])|(((m[181]&m[520]&~m[1304]))&~BiasedRNG[695])|((m[181]&m[520]&m[1304]));
    m[717] = (((m[195]&~m[521]&m[1359])|(~m[195]&m[521]&m[1359]))&BiasedRNG[696])|(((m[195]&m[521]&~m[1359]))&~BiasedRNG[696])|((m[195]&m[521]&m[1359]));
    m[718] = (((m[209]&~m[522]&m[1409])|(~m[209]&m[522]&m[1409]))&BiasedRNG[697])|(((m[209]&m[522]&~m[1409]))&~BiasedRNG[697])|((m[209]&m[522]&m[1409]));
    m[719] = (((m[223]&~m[523]&m[1454])|(~m[223]&m[523]&m[1454]))&BiasedRNG[698])|(((m[223]&m[523]&~m[1454]))&~BiasedRNG[698])|((m[223]&m[523]&m[1454]));
    m[729] = (((m[546]&~m[728]&~m[730]&~m[731]&~m[732])|(~m[546]&~m[728]&~m[730]&m[731]&~m[732])|(m[546]&m[728]&~m[730]&m[731]&~m[732])|(m[546]&~m[728]&m[730]&m[731]&~m[732])|(~m[546]&m[728]&~m[730]&~m[731]&m[732])|(~m[546]&~m[728]&m[730]&~m[731]&m[732])|(m[546]&m[728]&m[730]&~m[731]&m[732])|(~m[546]&m[728]&m[730]&m[731]&m[732]))&UnbiasedRNG[386])|((m[546]&~m[728]&~m[730]&m[731]&~m[732])|(~m[546]&~m[728]&~m[730]&~m[731]&m[732])|(m[546]&~m[728]&~m[730]&~m[731]&m[732])|(m[546]&m[728]&~m[730]&~m[731]&m[732])|(m[546]&~m[728]&m[730]&~m[731]&m[732])|(~m[546]&~m[728]&~m[730]&m[731]&m[732])|(m[546]&~m[728]&~m[730]&m[731]&m[732])|(~m[546]&m[728]&~m[730]&m[731]&m[732])|(m[546]&m[728]&~m[730]&m[731]&m[732])|(~m[546]&~m[728]&m[730]&m[731]&m[732])|(m[546]&~m[728]&m[730]&m[731]&m[732])|(m[546]&m[728]&m[730]&m[731]&m[732]));
    m[734] = (((m[547]&~m[733]&~m[735]&~m[736]&~m[737])|(~m[547]&~m[733]&~m[735]&m[736]&~m[737])|(m[547]&m[733]&~m[735]&m[736]&~m[737])|(m[547]&~m[733]&m[735]&m[736]&~m[737])|(~m[547]&m[733]&~m[735]&~m[736]&m[737])|(~m[547]&~m[733]&m[735]&~m[736]&m[737])|(m[547]&m[733]&m[735]&~m[736]&m[737])|(~m[547]&m[733]&m[735]&m[736]&m[737]))&UnbiasedRNG[387])|((m[547]&~m[733]&~m[735]&m[736]&~m[737])|(~m[547]&~m[733]&~m[735]&~m[736]&m[737])|(m[547]&~m[733]&~m[735]&~m[736]&m[737])|(m[547]&m[733]&~m[735]&~m[736]&m[737])|(m[547]&~m[733]&m[735]&~m[736]&m[737])|(~m[547]&~m[733]&~m[735]&m[736]&m[737])|(m[547]&~m[733]&~m[735]&m[736]&m[737])|(~m[547]&m[733]&~m[735]&m[736]&m[737])|(m[547]&m[733]&~m[735]&m[736]&m[737])|(~m[547]&~m[733]&m[735]&m[736]&m[737])|(m[547]&~m[733]&m[735]&m[736]&m[737])|(m[547]&m[733]&m[735]&m[736]&m[737]));
    m[739] = (((m[560]&~m[738]&~m[740]&~m[741]&~m[742])|(~m[560]&~m[738]&~m[740]&m[741]&~m[742])|(m[560]&m[738]&~m[740]&m[741]&~m[742])|(m[560]&~m[738]&m[740]&m[741]&~m[742])|(~m[560]&m[738]&~m[740]&~m[741]&m[742])|(~m[560]&~m[738]&m[740]&~m[741]&m[742])|(m[560]&m[738]&m[740]&~m[741]&m[742])|(~m[560]&m[738]&m[740]&m[741]&m[742]))&UnbiasedRNG[388])|((m[560]&~m[738]&~m[740]&m[741]&~m[742])|(~m[560]&~m[738]&~m[740]&~m[741]&m[742])|(m[560]&~m[738]&~m[740]&~m[741]&m[742])|(m[560]&m[738]&~m[740]&~m[741]&m[742])|(m[560]&~m[738]&m[740]&~m[741]&m[742])|(~m[560]&~m[738]&~m[740]&m[741]&m[742])|(m[560]&~m[738]&~m[740]&m[741]&m[742])|(~m[560]&m[738]&~m[740]&m[741]&m[742])|(m[560]&m[738]&~m[740]&m[741]&m[742])|(~m[560]&~m[738]&m[740]&m[741]&m[742])|(m[560]&~m[738]&m[740]&m[741]&m[742])|(m[560]&m[738]&m[740]&m[741]&m[742]));
    m[744] = (((m[548]&~m[743]&~m[745]&~m[746]&~m[747])|(~m[548]&~m[743]&~m[745]&m[746]&~m[747])|(m[548]&m[743]&~m[745]&m[746]&~m[747])|(m[548]&~m[743]&m[745]&m[746]&~m[747])|(~m[548]&m[743]&~m[745]&~m[746]&m[747])|(~m[548]&~m[743]&m[745]&~m[746]&m[747])|(m[548]&m[743]&m[745]&~m[746]&m[747])|(~m[548]&m[743]&m[745]&m[746]&m[747]))&UnbiasedRNG[389])|((m[548]&~m[743]&~m[745]&m[746]&~m[747])|(~m[548]&~m[743]&~m[745]&~m[746]&m[747])|(m[548]&~m[743]&~m[745]&~m[746]&m[747])|(m[548]&m[743]&~m[745]&~m[746]&m[747])|(m[548]&~m[743]&m[745]&~m[746]&m[747])|(~m[548]&~m[743]&~m[745]&m[746]&m[747])|(m[548]&~m[743]&~m[745]&m[746]&m[747])|(~m[548]&m[743]&~m[745]&m[746]&m[747])|(m[548]&m[743]&~m[745]&m[746]&m[747])|(~m[548]&~m[743]&m[745]&m[746]&m[747])|(m[548]&~m[743]&m[745]&m[746]&m[747])|(m[548]&m[743]&m[745]&m[746]&m[747]));
    m[749] = (((m[561]&~m[748]&~m[750]&~m[751]&~m[752])|(~m[561]&~m[748]&~m[750]&m[751]&~m[752])|(m[561]&m[748]&~m[750]&m[751]&~m[752])|(m[561]&~m[748]&m[750]&m[751]&~m[752])|(~m[561]&m[748]&~m[750]&~m[751]&m[752])|(~m[561]&~m[748]&m[750]&~m[751]&m[752])|(m[561]&m[748]&m[750]&~m[751]&m[752])|(~m[561]&m[748]&m[750]&m[751]&m[752]))&UnbiasedRNG[390])|((m[561]&~m[748]&~m[750]&m[751]&~m[752])|(~m[561]&~m[748]&~m[750]&~m[751]&m[752])|(m[561]&~m[748]&~m[750]&~m[751]&m[752])|(m[561]&m[748]&~m[750]&~m[751]&m[752])|(m[561]&~m[748]&m[750]&~m[751]&m[752])|(~m[561]&~m[748]&~m[750]&m[751]&m[752])|(m[561]&~m[748]&~m[750]&m[751]&m[752])|(~m[561]&m[748]&~m[750]&m[751]&m[752])|(m[561]&m[748]&~m[750]&m[751]&m[752])|(~m[561]&~m[748]&m[750]&m[751]&m[752])|(m[561]&~m[748]&m[750]&m[751]&m[752])|(m[561]&m[748]&m[750]&m[751]&m[752]));
    m[754] = (((m[574]&~m[753]&~m[755]&~m[756]&~m[757])|(~m[574]&~m[753]&~m[755]&m[756]&~m[757])|(m[574]&m[753]&~m[755]&m[756]&~m[757])|(m[574]&~m[753]&m[755]&m[756]&~m[757])|(~m[574]&m[753]&~m[755]&~m[756]&m[757])|(~m[574]&~m[753]&m[755]&~m[756]&m[757])|(m[574]&m[753]&m[755]&~m[756]&m[757])|(~m[574]&m[753]&m[755]&m[756]&m[757]))&UnbiasedRNG[391])|((m[574]&~m[753]&~m[755]&m[756]&~m[757])|(~m[574]&~m[753]&~m[755]&~m[756]&m[757])|(m[574]&~m[753]&~m[755]&~m[756]&m[757])|(m[574]&m[753]&~m[755]&~m[756]&m[757])|(m[574]&~m[753]&m[755]&~m[756]&m[757])|(~m[574]&~m[753]&~m[755]&m[756]&m[757])|(m[574]&~m[753]&~m[755]&m[756]&m[757])|(~m[574]&m[753]&~m[755]&m[756]&m[757])|(m[574]&m[753]&~m[755]&m[756]&m[757])|(~m[574]&~m[753]&m[755]&m[756]&m[757])|(m[574]&~m[753]&m[755]&m[756]&m[757])|(m[574]&m[753]&m[755]&m[756]&m[757]));
    m[759] = (((m[549]&~m[758]&~m[760]&~m[761]&~m[762])|(~m[549]&~m[758]&~m[760]&m[761]&~m[762])|(m[549]&m[758]&~m[760]&m[761]&~m[762])|(m[549]&~m[758]&m[760]&m[761]&~m[762])|(~m[549]&m[758]&~m[760]&~m[761]&m[762])|(~m[549]&~m[758]&m[760]&~m[761]&m[762])|(m[549]&m[758]&m[760]&~m[761]&m[762])|(~m[549]&m[758]&m[760]&m[761]&m[762]))&UnbiasedRNG[392])|((m[549]&~m[758]&~m[760]&m[761]&~m[762])|(~m[549]&~m[758]&~m[760]&~m[761]&m[762])|(m[549]&~m[758]&~m[760]&~m[761]&m[762])|(m[549]&m[758]&~m[760]&~m[761]&m[762])|(m[549]&~m[758]&m[760]&~m[761]&m[762])|(~m[549]&~m[758]&~m[760]&m[761]&m[762])|(m[549]&~m[758]&~m[760]&m[761]&m[762])|(~m[549]&m[758]&~m[760]&m[761]&m[762])|(m[549]&m[758]&~m[760]&m[761]&m[762])|(~m[549]&~m[758]&m[760]&m[761]&m[762])|(m[549]&~m[758]&m[760]&m[761]&m[762])|(m[549]&m[758]&m[760]&m[761]&m[762]));
    m[764] = (((m[562]&~m[763]&~m[765]&~m[766]&~m[767])|(~m[562]&~m[763]&~m[765]&m[766]&~m[767])|(m[562]&m[763]&~m[765]&m[766]&~m[767])|(m[562]&~m[763]&m[765]&m[766]&~m[767])|(~m[562]&m[763]&~m[765]&~m[766]&m[767])|(~m[562]&~m[763]&m[765]&~m[766]&m[767])|(m[562]&m[763]&m[765]&~m[766]&m[767])|(~m[562]&m[763]&m[765]&m[766]&m[767]))&UnbiasedRNG[393])|((m[562]&~m[763]&~m[765]&m[766]&~m[767])|(~m[562]&~m[763]&~m[765]&~m[766]&m[767])|(m[562]&~m[763]&~m[765]&~m[766]&m[767])|(m[562]&m[763]&~m[765]&~m[766]&m[767])|(m[562]&~m[763]&m[765]&~m[766]&m[767])|(~m[562]&~m[763]&~m[765]&m[766]&m[767])|(m[562]&~m[763]&~m[765]&m[766]&m[767])|(~m[562]&m[763]&~m[765]&m[766]&m[767])|(m[562]&m[763]&~m[765]&m[766]&m[767])|(~m[562]&~m[763]&m[765]&m[766]&m[767])|(m[562]&~m[763]&m[765]&m[766]&m[767])|(m[562]&m[763]&m[765]&m[766]&m[767]));
    m[769] = (((m[575]&~m[768]&~m[770]&~m[771]&~m[772])|(~m[575]&~m[768]&~m[770]&m[771]&~m[772])|(m[575]&m[768]&~m[770]&m[771]&~m[772])|(m[575]&~m[768]&m[770]&m[771]&~m[772])|(~m[575]&m[768]&~m[770]&~m[771]&m[772])|(~m[575]&~m[768]&m[770]&~m[771]&m[772])|(m[575]&m[768]&m[770]&~m[771]&m[772])|(~m[575]&m[768]&m[770]&m[771]&m[772]))&UnbiasedRNG[394])|((m[575]&~m[768]&~m[770]&m[771]&~m[772])|(~m[575]&~m[768]&~m[770]&~m[771]&m[772])|(m[575]&~m[768]&~m[770]&~m[771]&m[772])|(m[575]&m[768]&~m[770]&~m[771]&m[772])|(m[575]&~m[768]&m[770]&~m[771]&m[772])|(~m[575]&~m[768]&~m[770]&m[771]&m[772])|(m[575]&~m[768]&~m[770]&m[771]&m[772])|(~m[575]&m[768]&~m[770]&m[771]&m[772])|(m[575]&m[768]&~m[770]&m[771]&m[772])|(~m[575]&~m[768]&m[770]&m[771]&m[772])|(m[575]&~m[768]&m[770]&m[771]&m[772])|(m[575]&m[768]&m[770]&m[771]&m[772]));
    m[774] = (((m[588]&~m[773]&~m[775]&~m[776]&~m[777])|(~m[588]&~m[773]&~m[775]&m[776]&~m[777])|(m[588]&m[773]&~m[775]&m[776]&~m[777])|(m[588]&~m[773]&m[775]&m[776]&~m[777])|(~m[588]&m[773]&~m[775]&~m[776]&m[777])|(~m[588]&~m[773]&m[775]&~m[776]&m[777])|(m[588]&m[773]&m[775]&~m[776]&m[777])|(~m[588]&m[773]&m[775]&m[776]&m[777]))&UnbiasedRNG[395])|((m[588]&~m[773]&~m[775]&m[776]&~m[777])|(~m[588]&~m[773]&~m[775]&~m[776]&m[777])|(m[588]&~m[773]&~m[775]&~m[776]&m[777])|(m[588]&m[773]&~m[775]&~m[776]&m[777])|(m[588]&~m[773]&m[775]&~m[776]&m[777])|(~m[588]&~m[773]&~m[775]&m[776]&m[777])|(m[588]&~m[773]&~m[775]&m[776]&m[777])|(~m[588]&m[773]&~m[775]&m[776]&m[777])|(m[588]&m[773]&~m[775]&m[776]&m[777])|(~m[588]&~m[773]&m[775]&m[776]&m[777])|(m[588]&~m[773]&m[775]&m[776]&m[777])|(m[588]&m[773]&m[775]&m[776]&m[777]));
    m[779] = (((m[550]&~m[778]&~m[780]&~m[781]&~m[782])|(~m[550]&~m[778]&~m[780]&m[781]&~m[782])|(m[550]&m[778]&~m[780]&m[781]&~m[782])|(m[550]&~m[778]&m[780]&m[781]&~m[782])|(~m[550]&m[778]&~m[780]&~m[781]&m[782])|(~m[550]&~m[778]&m[780]&~m[781]&m[782])|(m[550]&m[778]&m[780]&~m[781]&m[782])|(~m[550]&m[778]&m[780]&m[781]&m[782]))&UnbiasedRNG[396])|((m[550]&~m[778]&~m[780]&m[781]&~m[782])|(~m[550]&~m[778]&~m[780]&~m[781]&m[782])|(m[550]&~m[778]&~m[780]&~m[781]&m[782])|(m[550]&m[778]&~m[780]&~m[781]&m[782])|(m[550]&~m[778]&m[780]&~m[781]&m[782])|(~m[550]&~m[778]&~m[780]&m[781]&m[782])|(m[550]&~m[778]&~m[780]&m[781]&m[782])|(~m[550]&m[778]&~m[780]&m[781]&m[782])|(m[550]&m[778]&~m[780]&m[781]&m[782])|(~m[550]&~m[778]&m[780]&m[781]&m[782])|(m[550]&~m[778]&m[780]&m[781]&m[782])|(m[550]&m[778]&m[780]&m[781]&m[782]));
    m[784] = (((m[563]&~m[783]&~m[785]&~m[786]&~m[787])|(~m[563]&~m[783]&~m[785]&m[786]&~m[787])|(m[563]&m[783]&~m[785]&m[786]&~m[787])|(m[563]&~m[783]&m[785]&m[786]&~m[787])|(~m[563]&m[783]&~m[785]&~m[786]&m[787])|(~m[563]&~m[783]&m[785]&~m[786]&m[787])|(m[563]&m[783]&m[785]&~m[786]&m[787])|(~m[563]&m[783]&m[785]&m[786]&m[787]))&UnbiasedRNG[397])|((m[563]&~m[783]&~m[785]&m[786]&~m[787])|(~m[563]&~m[783]&~m[785]&~m[786]&m[787])|(m[563]&~m[783]&~m[785]&~m[786]&m[787])|(m[563]&m[783]&~m[785]&~m[786]&m[787])|(m[563]&~m[783]&m[785]&~m[786]&m[787])|(~m[563]&~m[783]&~m[785]&m[786]&m[787])|(m[563]&~m[783]&~m[785]&m[786]&m[787])|(~m[563]&m[783]&~m[785]&m[786]&m[787])|(m[563]&m[783]&~m[785]&m[786]&m[787])|(~m[563]&~m[783]&m[785]&m[786]&m[787])|(m[563]&~m[783]&m[785]&m[786]&m[787])|(m[563]&m[783]&m[785]&m[786]&m[787]));
    m[789] = (((m[576]&~m[788]&~m[790]&~m[791]&~m[792])|(~m[576]&~m[788]&~m[790]&m[791]&~m[792])|(m[576]&m[788]&~m[790]&m[791]&~m[792])|(m[576]&~m[788]&m[790]&m[791]&~m[792])|(~m[576]&m[788]&~m[790]&~m[791]&m[792])|(~m[576]&~m[788]&m[790]&~m[791]&m[792])|(m[576]&m[788]&m[790]&~m[791]&m[792])|(~m[576]&m[788]&m[790]&m[791]&m[792]))&UnbiasedRNG[398])|((m[576]&~m[788]&~m[790]&m[791]&~m[792])|(~m[576]&~m[788]&~m[790]&~m[791]&m[792])|(m[576]&~m[788]&~m[790]&~m[791]&m[792])|(m[576]&m[788]&~m[790]&~m[791]&m[792])|(m[576]&~m[788]&m[790]&~m[791]&m[792])|(~m[576]&~m[788]&~m[790]&m[791]&m[792])|(m[576]&~m[788]&~m[790]&m[791]&m[792])|(~m[576]&m[788]&~m[790]&m[791]&m[792])|(m[576]&m[788]&~m[790]&m[791]&m[792])|(~m[576]&~m[788]&m[790]&m[791]&m[792])|(m[576]&~m[788]&m[790]&m[791]&m[792])|(m[576]&m[788]&m[790]&m[791]&m[792]));
    m[794] = (((m[589]&~m[793]&~m[795]&~m[796]&~m[797])|(~m[589]&~m[793]&~m[795]&m[796]&~m[797])|(m[589]&m[793]&~m[795]&m[796]&~m[797])|(m[589]&~m[793]&m[795]&m[796]&~m[797])|(~m[589]&m[793]&~m[795]&~m[796]&m[797])|(~m[589]&~m[793]&m[795]&~m[796]&m[797])|(m[589]&m[793]&m[795]&~m[796]&m[797])|(~m[589]&m[793]&m[795]&m[796]&m[797]))&UnbiasedRNG[399])|((m[589]&~m[793]&~m[795]&m[796]&~m[797])|(~m[589]&~m[793]&~m[795]&~m[796]&m[797])|(m[589]&~m[793]&~m[795]&~m[796]&m[797])|(m[589]&m[793]&~m[795]&~m[796]&m[797])|(m[589]&~m[793]&m[795]&~m[796]&m[797])|(~m[589]&~m[793]&~m[795]&m[796]&m[797])|(m[589]&~m[793]&~m[795]&m[796]&m[797])|(~m[589]&m[793]&~m[795]&m[796]&m[797])|(m[589]&m[793]&~m[795]&m[796]&m[797])|(~m[589]&~m[793]&m[795]&m[796]&m[797])|(m[589]&~m[793]&m[795]&m[796]&m[797])|(m[589]&m[793]&m[795]&m[796]&m[797]));
    m[799] = (((m[602]&~m[798]&~m[800]&~m[801]&~m[802])|(~m[602]&~m[798]&~m[800]&m[801]&~m[802])|(m[602]&m[798]&~m[800]&m[801]&~m[802])|(m[602]&~m[798]&m[800]&m[801]&~m[802])|(~m[602]&m[798]&~m[800]&~m[801]&m[802])|(~m[602]&~m[798]&m[800]&~m[801]&m[802])|(m[602]&m[798]&m[800]&~m[801]&m[802])|(~m[602]&m[798]&m[800]&m[801]&m[802]))&UnbiasedRNG[400])|((m[602]&~m[798]&~m[800]&m[801]&~m[802])|(~m[602]&~m[798]&~m[800]&~m[801]&m[802])|(m[602]&~m[798]&~m[800]&~m[801]&m[802])|(m[602]&m[798]&~m[800]&~m[801]&m[802])|(m[602]&~m[798]&m[800]&~m[801]&m[802])|(~m[602]&~m[798]&~m[800]&m[801]&m[802])|(m[602]&~m[798]&~m[800]&m[801]&m[802])|(~m[602]&m[798]&~m[800]&m[801]&m[802])|(m[602]&m[798]&~m[800]&m[801]&m[802])|(~m[602]&~m[798]&m[800]&m[801]&m[802])|(m[602]&~m[798]&m[800]&m[801]&m[802])|(m[602]&m[798]&m[800]&m[801]&m[802]));
    m[804] = (((m[551]&~m[803]&~m[805]&~m[806]&~m[807])|(~m[551]&~m[803]&~m[805]&m[806]&~m[807])|(m[551]&m[803]&~m[805]&m[806]&~m[807])|(m[551]&~m[803]&m[805]&m[806]&~m[807])|(~m[551]&m[803]&~m[805]&~m[806]&m[807])|(~m[551]&~m[803]&m[805]&~m[806]&m[807])|(m[551]&m[803]&m[805]&~m[806]&m[807])|(~m[551]&m[803]&m[805]&m[806]&m[807]))&UnbiasedRNG[401])|((m[551]&~m[803]&~m[805]&m[806]&~m[807])|(~m[551]&~m[803]&~m[805]&~m[806]&m[807])|(m[551]&~m[803]&~m[805]&~m[806]&m[807])|(m[551]&m[803]&~m[805]&~m[806]&m[807])|(m[551]&~m[803]&m[805]&~m[806]&m[807])|(~m[551]&~m[803]&~m[805]&m[806]&m[807])|(m[551]&~m[803]&~m[805]&m[806]&m[807])|(~m[551]&m[803]&~m[805]&m[806]&m[807])|(m[551]&m[803]&~m[805]&m[806]&m[807])|(~m[551]&~m[803]&m[805]&m[806]&m[807])|(m[551]&~m[803]&m[805]&m[806]&m[807])|(m[551]&m[803]&m[805]&m[806]&m[807]));
    m[809] = (((m[564]&~m[808]&~m[810]&~m[811]&~m[812])|(~m[564]&~m[808]&~m[810]&m[811]&~m[812])|(m[564]&m[808]&~m[810]&m[811]&~m[812])|(m[564]&~m[808]&m[810]&m[811]&~m[812])|(~m[564]&m[808]&~m[810]&~m[811]&m[812])|(~m[564]&~m[808]&m[810]&~m[811]&m[812])|(m[564]&m[808]&m[810]&~m[811]&m[812])|(~m[564]&m[808]&m[810]&m[811]&m[812]))&UnbiasedRNG[402])|((m[564]&~m[808]&~m[810]&m[811]&~m[812])|(~m[564]&~m[808]&~m[810]&~m[811]&m[812])|(m[564]&~m[808]&~m[810]&~m[811]&m[812])|(m[564]&m[808]&~m[810]&~m[811]&m[812])|(m[564]&~m[808]&m[810]&~m[811]&m[812])|(~m[564]&~m[808]&~m[810]&m[811]&m[812])|(m[564]&~m[808]&~m[810]&m[811]&m[812])|(~m[564]&m[808]&~m[810]&m[811]&m[812])|(m[564]&m[808]&~m[810]&m[811]&m[812])|(~m[564]&~m[808]&m[810]&m[811]&m[812])|(m[564]&~m[808]&m[810]&m[811]&m[812])|(m[564]&m[808]&m[810]&m[811]&m[812]));
    m[814] = (((m[577]&~m[813]&~m[815]&~m[816]&~m[817])|(~m[577]&~m[813]&~m[815]&m[816]&~m[817])|(m[577]&m[813]&~m[815]&m[816]&~m[817])|(m[577]&~m[813]&m[815]&m[816]&~m[817])|(~m[577]&m[813]&~m[815]&~m[816]&m[817])|(~m[577]&~m[813]&m[815]&~m[816]&m[817])|(m[577]&m[813]&m[815]&~m[816]&m[817])|(~m[577]&m[813]&m[815]&m[816]&m[817]))&UnbiasedRNG[403])|((m[577]&~m[813]&~m[815]&m[816]&~m[817])|(~m[577]&~m[813]&~m[815]&~m[816]&m[817])|(m[577]&~m[813]&~m[815]&~m[816]&m[817])|(m[577]&m[813]&~m[815]&~m[816]&m[817])|(m[577]&~m[813]&m[815]&~m[816]&m[817])|(~m[577]&~m[813]&~m[815]&m[816]&m[817])|(m[577]&~m[813]&~m[815]&m[816]&m[817])|(~m[577]&m[813]&~m[815]&m[816]&m[817])|(m[577]&m[813]&~m[815]&m[816]&m[817])|(~m[577]&~m[813]&m[815]&m[816]&m[817])|(m[577]&~m[813]&m[815]&m[816]&m[817])|(m[577]&m[813]&m[815]&m[816]&m[817]));
    m[819] = (((m[590]&~m[818]&~m[820]&~m[821]&~m[822])|(~m[590]&~m[818]&~m[820]&m[821]&~m[822])|(m[590]&m[818]&~m[820]&m[821]&~m[822])|(m[590]&~m[818]&m[820]&m[821]&~m[822])|(~m[590]&m[818]&~m[820]&~m[821]&m[822])|(~m[590]&~m[818]&m[820]&~m[821]&m[822])|(m[590]&m[818]&m[820]&~m[821]&m[822])|(~m[590]&m[818]&m[820]&m[821]&m[822]))&UnbiasedRNG[404])|((m[590]&~m[818]&~m[820]&m[821]&~m[822])|(~m[590]&~m[818]&~m[820]&~m[821]&m[822])|(m[590]&~m[818]&~m[820]&~m[821]&m[822])|(m[590]&m[818]&~m[820]&~m[821]&m[822])|(m[590]&~m[818]&m[820]&~m[821]&m[822])|(~m[590]&~m[818]&~m[820]&m[821]&m[822])|(m[590]&~m[818]&~m[820]&m[821]&m[822])|(~m[590]&m[818]&~m[820]&m[821]&m[822])|(m[590]&m[818]&~m[820]&m[821]&m[822])|(~m[590]&~m[818]&m[820]&m[821]&m[822])|(m[590]&~m[818]&m[820]&m[821]&m[822])|(m[590]&m[818]&m[820]&m[821]&m[822]));
    m[824] = (((m[603]&~m[823]&~m[825]&~m[826]&~m[827])|(~m[603]&~m[823]&~m[825]&m[826]&~m[827])|(m[603]&m[823]&~m[825]&m[826]&~m[827])|(m[603]&~m[823]&m[825]&m[826]&~m[827])|(~m[603]&m[823]&~m[825]&~m[826]&m[827])|(~m[603]&~m[823]&m[825]&~m[826]&m[827])|(m[603]&m[823]&m[825]&~m[826]&m[827])|(~m[603]&m[823]&m[825]&m[826]&m[827]))&UnbiasedRNG[405])|((m[603]&~m[823]&~m[825]&m[826]&~m[827])|(~m[603]&~m[823]&~m[825]&~m[826]&m[827])|(m[603]&~m[823]&~m[825]&~m[826]&m[827])|(m[603]&m[823]&~m[825]&~m[826]&m[827])|(m[603]&~m[823]&m[825]&~m[826]&m[827])|(~m[603]&~m[823]&~m[825]&m[826]&m[827])|(m[603]&~m[823]&~m[825]&m[826]&m[827])|(~m[603]&m[823]&~m[825]&m[826]&m[827])|(m[603]&m[823]&~m[825]&m[826]&m[827])|(~m[603]&~m[823]&m[825]&m[826]&m[827])|(m[603]&~m[823]&m[825]&m[826]&m[827])|(m[603]&m[823]&m[825]&m[826]&m[827]));
    m[835] = (((m[807]&~m[833]&~m[834]&~m[836]&~m[837])|(~m[807]&~m[833]&~m[834]&m[836]&~m[837])|(m[807]&m[833]&~m[834]&m[836]&~m[837])|(m[807]&~m[833]&m[834]&m[836]&~m[837])|(~m[807]&m[833]&~m[834]&~m[836]&m[837])|(~m[807]&~m[833]&m[834]&~m[836]&m[837])|(m[807]&m[833]&m[834]&~m[836]&m[837])|(~m[807]&m[833]&m[834]&m[836]&m[837]))&UnbiasedRNG[406])|((m[807]&~m[833]&~m[834]&m[836]&~m[837])|(~m[807]&~m[833]&~m[834]&~m[836]&m[837])|(m[807]&~m[833]&~m[834]&~m[836]&m[837])|(m[807]&m[833]&~m[834]&~m[836]&m[837])|(m[807]&~m[833]&m[834]&~m[836]&m[837])|(~m[807]&~m[833]&~m[834]&m[836]&m[837])|(m[807]&~m[833]&~m[834]&m[836]&m[837])|(~m[807]&m[833]&~m[834]&m[836]&m[837])|(m[807]&m[833]&~m[834]&m[836]&m[837])|(~m[807]&~m[833]&m[834]&m[836]&m[837])|(m[807]&~m[833]&m[834]&m[836]&m[837])|(m[807]&m[833]&m[834]&m[836]&m[837]));
    m[839] = (((m[565]&~m[838]&~m[840]&~m[841]&~m[842])|(~m[565]&~m[838]&~m[840]&m[841]&~m[842])|(m[565]&m[838]&~m[840]&m[841]&~m[842])|(m[565]&~m[838]&m[840]&m[841]&~m[842])|(~m[565]&m[838]&~m[840]&~m[841]&m[842])|(~m[565]&~m[838]&m[840]&~m[841]&m[842])|(m[565]&m[838]&m[840]&~m[841]&m[842])|(~m[565]&m[838]&m[840]&m[841]&m[842]))&UnbiasedRNG[407])|((m[565]&~m[838]&~m[840]&m[841]&~m[842])|(~m[565]&~m[838]&~m[840]&~m[841]&m[842])|(m[565]&~m[838]&~m[840]&~m[841]&m[842])|(m[565]&m[838]&~m[840]&~m[841]&m[842])|(m[565]&~m[838]&m[840]&~m[841]&m[842])|(~m[565]&~m[838]&~m[840]&m[841]&m[842])|(m[565]&~m[838]&~m[840]&m[841]&m[842])|(~m[565]&m[838]&~m[840]&m[841]&m[842])|(m[565]&m[838]&~m[840]&m[841]&m[842])|(~m[565]&~m[838]&m[840]&m[841]&m[842])|(m[565]&~m[838]&m[840]&m[841]&m[842])|(m[565]&m[838]&m[840]&m[841]&m[842]));
    m[844] = (((m[578]&~m[843]&~m[845]&~m[846]&~m[847])|(~m[578]&~m[843]&~m[845]&m[846]&~m[847])|(m[578]&m[843]&~m[845]&m[846]&~m[847])|(m[578]&~m[843]&m[845]&m[846]&~m[847])|(~m[578]&m[843]&~m[845]&~m[846]&m[847])|(~m[578]&~m[843]&m[845]&~m[846]&m[847])|(m[578]&m[843]&m[845]&~m[846]&m[847])|(~m[578]&m[843]&m[845]&m[846]&m[847]))&UnbiasedRNG[408])|((m[578]&~m[843]&~m[845]&m[846]&~m[847])|(~m[578]&~m[843]&~m[845]&~m[846]&m[847])|(m[578]&~m[843]&~m[845]&~m[846]&m[847])|(m[578]&m[843]&~m[845]&~m[846]&m[847])|(m[578]&~m[843]&m[845]&~m[846]&m[847])|(~m[578]&~m[843]&~m[845]&m[846]&m[847])|(m[578]&~m[843]&~m[845]&m[846]&m[847])|(~m[578]&m[843]&~m[845]&m[846]&m[847])|(m[578]&m[843]&~m[845]&m[846]&m[847])|(~m[578]&~m[843]&m[845]&m[846]&m[847])|(m[578]&~m[843]&m[845]&m[846]&m[847])|(m[578]&m[843]&m[845]&m[846]&m[847]));
    m[849] = (((m[591]&~m[848]&~m[850]&~m[851]&~m[852])|(~m[591]&~m[848]&~m[850]&m[851]&~m[852])|(m[591]&m[848]&~m[850]&m[851]&~m[852])|(m[591]&~m[848]&m[850]&m[851]&~m[852])|(~m[591]&m[848]&~m[850]&~m[851]&m[852])|(~m[591]&~m[848]&m[850]&~m[851]&m[852])|(m[591]&m[848]&m[850]&~m[851]&m[852])|(~m[591]&m[848]&m[850]&m[851]&m[852]))&UnbiasedRNG[409])|((m[591]&~m[848]&~m[850]&m[851]&~m[852])|(~m[591]&~m[848]&~m[850]&~m[851]&m[852])|(m[591]&~m[848]&~m[850]&~m[851]&m[852])|(m[591]&m[848]&~m[850]&~m[851]&m[852])|(m[591]&~m[848]&m[850]&~m[851]&m[852])|(~m[591]&~m[848]&~m[850]&m[851]&m[852])|(m[591]&~m[848]&~m[850]&m[851]&m[852])|(~m[591]&m[848]&~m[850]&m[851]&m[852])|(m[591]&m[848]&~m[850]&m[851]&m[852])|(~m[591]&~m[848]&m[850]&m[851]&m[852])|(m[591]&~m[848]&m[850]&m[851]&m[852])|(m[591]&m[848]&m[850]&m[851]&m[852]));
    m[854] = (((m[604]&~m[853]&~m[855]&~m[856]&~m[857])|(~m[604]&~m[853]&~m[855]&m[856]&~m[857])|(m[604]&m[853]&~m[855]&m[856]&~m[857])|(m[604]&~m[853]&m[855]&m[856]&~m[857])|(~m[604]&m[853]&~m[855]&~m[856]&m[857])|(~m[604]&~m[853]&m[855]&~m[856]&m[857])|(m[604]&m[853]&m[855]&~m[856]&m[857])|(~m[604]&m[853]&m[855]&m[856]&m[857]))&UnbiasedRNG[410])|((m[604]&~m[853]&~m[855]&m[856]&~m[857])|(~m[604]&~m[853]&~m[855]&~m[856]&m[857])|(m[604]&~m[853]&~m[855]&~m[856]&m[857])|(m[604]&m[853]&~m[855]&~m[856]&m[857])|(m[604]&~m[853]&m[855]&~m[856]&m[857])|(~m[604]&~m[853]&~m[855]&m[856]&m[857])|(m[604]&~m[853]&~m[855]&m[856]&m[857])|(~m[604]&m[853]&~m[855]&m[856]&m[857])|(m[604]&m[853]&~m[855]&m[856]&m[857])|(~m[604]&~m[853]&m[855]&m[856]&m[857])|(m[604]&~m[853]&m[855]&m[856]&m[857])|(m[604]&m[853]&m[855]&m[856]&m[857]));
    m[860] = (((m[832]&~m[858]&~m[859]&~m[861]&~m[862])|(~m[832]&~m[858]&~m[859]&m[861]&~m[862])|(m[832]&m[858]&~m[859]&m[861]&~m[862])|(m[832]&~m[858]&m[859]&m[861]&~m[862])|(~m[832]&m[858]&~m[859]&~m[861]&m[862])|(~m[832]&~m[858]&m[859]&~m[861]&m[862])|(m[832]&m[858]&m[859]&~m[861]&m[862])|(~m[832]&m[858]&m[859]&m[861]&m[862]))&UnbiasedRNG[411])|((m[832]&~m[858]&~m[859]&m[861]&~m[862])|(~m[832]&~m[858]&~m[859]&~m[861]&m[862])|(m[832]&~m[858]&~m[859]&~m[861]&m[862])|(m[832]&m[858]&~m[859]&~m[861]&m[862])|(m[832]&~m[858]&m[859]&~m[861]&m[862])|(~m[832]&~m[858]&~m[859]&m[861]&m[862])|(m[832]&~m[858]&~m[859]&m[861]&m[862])|(~m[832]&m[858]&~m[859]&m[861]&m[862])|(m[832]&m[858]&~m[859]&m[861]&m[862])|(~m[832]&~m[858]&m[859]&m[861]&m[862])|(m[832]&~m[858]&m[859]&m[861]&m[862])|(m[832]&m[858]&m[859]&m[861]&m[862]));
    m[870] = (((m[837]&~m[868]&~m[869]&~m[871]&~m[872])|(~m[837]&~m[868]&~m[869]&m[871]&~m[872])|(m[837]&m[868]&~m[869]&m[871]&~m[872])|(m[837]&~m[868]&m[869]&m[871]&~m[872])|(~m[837]&m[868]&~m[869]&~m[871]&m[872])|(~m[837]&~m[868]&m[869]&~m[871]&m[872])|(m[837]&m[868]&m[869]&~m[871]&m[872])|(~m[837]&m[868]&m[869]&m[871]&m[872]))&UnbiasedRNG[412])|((m[837]&~m[868]&~m[869]&m[871]&~m[872])|(~m[837]&~m[868]&~m[869]&~m[871]&m[872])|(m[837]&~m[868]&~m[869]&~m[871]&m[872])|(m[837]&m[868]&~m[869]&~m[871]&m[872])|(m[837]&~m[868]&m[869]&~m[871]&m[872])|(~m[837]&~m[868]&~m[869]&m[871]&m[872])|(m[837]&~m[868]&~m[869]&m[871]&m[872])|(~m[837]&m[868]&~m[869]&m[871]&m[872])|(m[837]&m[868]&~m[869]&m[871]&m[872])|(~m[837]&~m[868]&m[869]&m[871]&m[872])|(m[837]&~m[868]&m[869]&m[871]&m[872])|(m[837]&m[868]&m[869]&m[871]&m[872]));
    m[875] = (((m[842]&~m[873]&~m[874]&~m[876]&~m[877])|(~m[842]&~m[873]&~m[874]&m[876]&~m[877])|(m[842]&m[873]&~m[874]&m[876]&~m[877])|(m[842]&~m[873]&m[874]&m[876]&~m[877])|(~m[842]&m[873]&~m[874]&~m[876]&m[877])|(~m[842]&~m[873]&m[874]&~m[876]&m[877])|(m[842]&m[873]&m[874]&~m[876]&m[877])|(~m[842]&m[873]&m[874]&m[876]&m[877]))&UnbiasedRNG[413])|((m[842]&~m[873]&~m[874]&m[876]&~m[877])|(~m[842]&~m[873]&~m[874]&~m[876]&m[877])|(m[842]&~m[873]&~m[874]&~m[876]&m[877])|(m[842]&m[873]&~m[874]&~m[876]&m[877])|(m[842]&~m[873]&m[874]&~m[876]&m[877])|(~m[842]&~m[873]&~m[874]&m[876]&m[877])|(m[842]&~m[873]&~m[874]&m[876]&m[877])|(~m[842]&m[873]&~m[874]&m[876]&m[877])|(m[842]&m[873]&~m[874]&m[876]&m[877])|(~m[842]&~m[873]&m[874]&m[876]&m[877])|(m[842]&~m[873]&m[874]&m[876]&m[877])|(m[842]&m[873]&m[874]&m[876]&m[877]));
    m[879] = (((m[579]&~m[878]&~m[880]&~m[881]&~m[882])|(~m[579]&~m[878]&~m[880]&m[881]&~m[882])|(m[579]&m[878]&~m[880]&m[881]&~m[882])|(m[579]&~m[878]&m[880]&m[881]&~m[882])|(~m[579]&m[878]&~m[880]&~m[881]&m[882])|(~m[579]&~m[878]&m[880]&~m[881]&m[882])|(m[579]&m[878]&m[880]&~m[881]&m[882])|(~m[579]&m[878]&m[880]&m[881]&m[882]))&UnbiasedRNG[414])|((m[579]&~m[878]&~m[880]&m[881]&~m[882])|(~m[579]&~m[878]&~m[880]&~m[881]&m[882])|(m[579]&~m[878]&~m[880]&~m[881]&m[882])|(m[579]&m[878]&~m[880]&~m[881]&m[882])|(m[579]&~m[878]&m[880]&~m[881]&m[882])|(~m[579]&~m[878]&~m[880]&m[881]&m[882])|(m[579]&~m[878]&~m[880]&m[881]&m[882])|(~m[579]&m[878]&~m[880]&m[881]&m[882])|(m[579]&m[878]&~m[880]&m[881]&m[882])|(~m[579]&~m[878]&m[880]&m[881]&m[882])|(m[579]&~m[878]&m[880]&m[881]&m[882])|(m[579]&m[878]&m[880]&m[881]&m[882]));
    m[884] = (((m[592]&~m[883]&~m[885]&~m[886]&~m[887])|(~m[592]&~m[883]&~m[885]&m[886]&~m[887])|(m[592]&m[883]&~m[885]&m[886]&~m[887])|(m[592]&~m[883]&m[885]&m[886]&~m[887])|(~m[592]&m[883]&~m[885]&~m[886]&m[887])|(~m[592]&~m[883]&m[885]&~m[886]&m[887])|(m[592]&m[883]&m[885]&~m[886]&m[887])|(~m[592]&m[883]&m[885]&m[886]&m[887]))&UnbiasedRNG[415])|((m[592]&~m[883]&~m[885]&m[886]&~m[887])|(~m[592]&~m[883]&~m[885]&~m[886]&m[887])|(m[592]&~m[883]&~m[885]&~m[886]&m[887])|(m[592]&m[883]&~m[885]&~m[886]&m[887])|(m[592]&~m[883]&m[885]&~m[886]&m[887])|(~m[592]&~m[883]&~m[885]&m[886]&m[887])|(m[592]&~m[883]&~m[885]&m[886]&m[887])|(~m[592]&m[883]&~m[885]&m[886]&m[887])|(m[592]&m[883]&~m[885]&m[886]&m[887])|(~m[592]&~m[883]&m[885]&m[886]&m[887])|(m[592]&~m[883]&m[885]&m[886]&m[887])|(m[592]&m[883]&m[885]&m[886]&m[887]));
    m[889] = (((m[605]&~m[888]&~m[890]&~m[891]&~m[892])|(~m[605]&~m[888]&~m[890]&m[891]&~m[892])|(m[605]&m[888]&~m[890]&m[891]&~m[892])|(m[605]&~m[888]&m[890]&m[891]&~m[892])|(~m[605]&m[888]&~m[890]&~m[891]&m[892])|(~m[605]&~m[888]&m[890]&~m[891]&m[892])|(m[605]&m[888]&m[890]&~m[891]&m[892])|(~m[605]&m[888]&m[890]&m[891]&m[892]))&UnbiasedRNG[416])|((m[605]&~m[888]&~m[890]&m[891]&~m[892])|(~m[605]&~m[888]&~m[890]&~m[891]&m[892])|(m[605]&~m[888]&~m[890]&~m[891]&m[892])|(m[605]&m[888]&~m[890]&~m[891]&m[892])|(m[605]&~m[888]&m[890]&~m[891]&m[892])|(~m[605]&~m[888]&~m[890]&m[891]&m[892])|(m[605]&~m[888]&~m[890]&m[891]&m[892])|(~m[605]&m[888]&~m[890]&m[891]&m[892])|(m[605]&m[888]&~m[890]&m[891]&m[892])|(~m[605]&~m[888]&m[890]&m[891]&m[892])|(m[605]&~m[888]&m[890]&m[891]&m[892])|(m[605]&m[888]&m[890]&m[891]&m[892]));
    m[895] = (((m[862]&~m[893]&~m[894]&~m[896]&~m[897])|(~m[862]&~m[893]&~m[894]&m[896]&~m[897])|(m[862]&m[893]&~m[894]&m[896]&~m[897])|(m[862]&~m[893]&m[894]&m[896]&~m[897])|(~m[862]&m[893]&~m[894]&~m[896]&m[897])|(~m[862]&~m[893]&m[894]&~m[896]&m[897])|(m[862]&m[893]&m[894]&~m[896]&m[897])|(~m[862]&m[893]&m[894]&m[896]&m[897]))&UnbiasedRNG[417])|((m[862]&~m[893]&~m[894]&m[896]&~m[897])|(~m[862]&~m[893]&~m[894]&~m[896]&m[897])|(m[862]&~m[893]&~m[894]&~m[896]&m[897])|(m[862]&m[893]&~m[894]&~m[896]&m[897])|(m[862]&~m[893]&m[894]&~m[896]&m[897])|(~m[862]&~m[893]&~m[894]&m[896]&m[897])|(m[862]&~m[893]&~m[894]&m[896]&m[897])|(~m[862]&m[893]&~m[894]&m[896]&m[897])|(m[862]&m[893]&~m[894]&m[896]&m[897])|(~m[862]&~m[893]&m[894]&m[896]&m[897])|(m[862]&~m[893]&m[894]&m[896]&m[897])|(m[862]&m[893]&m[894]&m[896]&m[897]));
    m[900] = (((m[867]&~m[898]&~m[899]&~m[901]&~m[902])|(~m[867]&~m[898]&~m[899]&m[901]&~m[902])|(m[867]&m[898]&~m[899]&m[901]&~m[902])|(m[867]&~m[898]&m[899]&m[901]&~m[902])|(~m[867]&m[898]&~m[899]&~m[901]&m[902])|(~m[867]&~m[898]&m[899]&~m[901]&m[902])|(m[867]&m[898]&m[899]&~m[901]&m[902])|(~m[867]&m[898]&m[899]&m[901]&m[902]))&UnbiasedRNG[418])|((m[867]&~m[898]&~m[899]&m[901]&~m[902])|(~m[867]&~m[898]&~m[899]&~m[901]&m[902])|(m[867]&~m[898]&~m[899]&~m[901]&m[902])|(m[867]&m[898]&~m[899]&~m[901]&m[902])|(m[867]&~m[898]&m[899]&~m[901]&m[902])|(~m[867]&~m[898]&~m[899]&m[901]&m[902])|(m[867]&~m[898]&~m[899]&m[901]&m[902])|(~m[867]&m[898]&~m[899]&m[901]&m[902])|(m[867]&m[898]&~m[899]&m[901]&m[902])|(~m[867]&~m[898]&m[899]&m[901]&m[902])|(m[867]&~m[898]&m[899]&m[901]&m[902])|(m[867]&m[898]&m[899]&m[901]&m[902]));
    m[910] = (((m[872]&~m[908]&~m[909]&~m[911]&~m[912])|(~m[872]&~m[908]&~m[909]&m[911]&~m[912])|(m[872]&m[908]&~m[909]&m[911]&~m[912])|(m[872]&~m[908]&m[909]&m[911]&~m[912])|(~m[872]&m[908]&~m[909]&~m[911]&m[912])|(~m[872]&~m[908]&m[909]&~m[911]&m[912])|(m[872]&m[908]&m[909]&~m[911]&m[912])|(~m[872]&m[908]&m[909]&m[911]&m[912]))&UnbiasedRNG[419])|((m[872]&~m[908]&~m[909]&m[911]&~m[912])|(~m[872]&~m[908]&~m[909]&~m[911]&m[912])|(m[872]&~m[908]&~m[909]&~m[911]&m[912])|(m[872]&m[908]&~m[909]&~m[911]&m[912])|(m[872]&~m[908]&m[909]&~m[911]&m[912])|(~m[872]&~m[908]&~m[909]&m[911]&m[912])|(m[872]&~m[908]&~m[909]&m[911]&m[912])|(~m[872]&m[908]&~m[909]&m[911]&m[912])|(m[872]&m[908]&~m[909]&m[911]&m[912])|(~m[872]&~m[908]&m[909]&m[911]&m[912])|(m[872]&~m[908]&m[909]&m[911]&m[912])|(m[872]&m[908]&m[909]&m[911]&m[912]));
    m[915] = (((m[877]&~m[913]&~m[914]&~m[916]&~m[917])|(~m[877]&~m[913]&~m[914]&m[916]&~m[917])|(m[877]&m[913]&~m[914]&m[916]&~m[917])|(m[877]&~m[913]&m[914]&m[916]&~m[917])|(~m[877]&m[913]&~m[914]&~m[916]&m[917])|(~m[877]&~m[913]&m[914]&~m[916]&m[917])|(m[877]&m[913]&m[914]&~m[916]&m[917])|(~m[877]&m[913]&m[914]&m[916]&m[917]))&UnbiasedRNG[420])|((m[877]&~m[913]&~m[914]&m[916]&~m[917])|(~m[877]&~m[913]&~m[914]&~m[916]&m[917])|(m[877]&~m[913]&~m[914]&~m[916]&m[917])|(m[877]&m[913]&~m[914]&~m[916]&m[917])|(m[877]&~m[913]&m[914]&~m[916]&m[917])|(~m[877]&~m[913]&~m[914]&m[916]&m[917])|(m[877]&~m[913]&~m[914]&m[916]&m[917])|(~m[877]&m[913]&~m[914]&m[916]&m[917])|(m[877]&m[913]&~m[914]&m[916]&m[917])|(~m[877]&~m[913]&m[914]&m[916]&m[917])|(m[877]&~m[913]&m[914]&m[916]&m[917])|(m[877]&m[913]&m[914]&m[916]&m[917]));
    m[920] = (((m[882]&~m[918]&~m[919]&~m[921]&~m[922])|(~m[882]&~m[918]&~m[919]&m[921]&~m[922])|(m[882]&m[918]&~m[919]&m[921]&~m[922])|(m[882]&~m[918]&m[919]&m[921]&~m[922])|(~m[882]&m[918]&~m[919]&~m[921]&m[922])|(~m[882]&~m[918]&m[919]&~m[921]&m[922])|(m[882]&m[918]&m[919]&~m[921]&m[922])|(~m[882]&m[918]&m[919]&m[921]&m[922]))&UnbiasedRNG[421])|((m[882]&~m[918]&~m[919]&m[921]&~m[922])|(~m[882]&~m[918]&~m[919]&~m[921]&m[922])|(m[882]&~m[918]&~m[919]&~m[921]&m[922])|(m[882]&m[918]&~m[919]&~m[921]&m[922])|(m[882]&~m[918]&m[919]&~m[921]&m[922])|(~m[882]&~m[918]&~m[919]&m[921]&m[922])|(m[882]&~m[918]&~m[919]&m[921]&m[922])|(~m[882]&m[918]&~m[919]&m[921]&m[922])|(m[882]&m[918]&~m[919]&m[921]&m[922])|(~m[882]&~m[918]&m[919]&m[921]&m[922])|(m[882]&~m[918]&m[919]&m[921]&m[922])|(m[882]&m[918]&m[919]&m[921]&m[922]));
    m[924] = (((m[593]&~m[923]&~m[925]&~m[926]&~m[927])|(~m[593]&~m[923]&~m[925]&m[926]&~m[927])|(m[593]&m[923]&~m[925]&m[926]&~m[927])|(m[593]&~m[923]&m[925]&m[926]&~m[927])|(~m[593]&m[923]&~m[925]&~m[926]&m[927])|(~m[593]&~m[923]&m[925]&~m[926]&m[927])|(m[593]&m[923]&m[925]&~m[926]&m[927])|(~m[593]&m[923]&m[925]&m[926]&m[927]))&UnbiasedRNG[422])|((m[593]&~m[923]&~m[925]&m[926]&~m[927])|(~m[593]&~m[923]&~m[925]&~m[926]&m[927])|(m[593]&~m[923]&~m[925]&~m[926]&m[927])|(m[593]&m[923]&~m[925]&~m[926]&m[927])|(m[593]&~m[923]&m[925]&~m[926]&m[927])|(~m[593]&~m[923]&~m[925]&m[926]&m[927])|(m[593]&~m[923]&~m[925]&m[926]&m[927])|(~m[593]&m[923]&~m[925]&m[926]&m[927])|(m[593]&m[923]&~m[925]&m[926]&m[927])|(~m[593]&~m[923]&m[925]&m[926]&m[927])|(m[593]&~m[923]&m[925]&m[926]&m[927])|(m[593]&m[923]&m[925]&m[926]&m[927]));
    m[929] = (((m[606]&~m[928]&~m[930]&~m[931]&~m[932])|(~m[606]&~m[928]&~m[930]&m[931]&~m[932])|(m[606]&m[928]&~m[930]&m[931]&~m[932])|(m[606]&~m[928]&m[930]&m[931]&~m[932])|(~m[606]&m[928]&~m[930]&~m[931]&m[932])|(~m[606]&~m[928]&m[930]&~m[931]&m[932])|(m[606]&m[928]&m[930]&~m[931]&m[932])|(~m[606]&m[928]&m[930]&m[931]&m[932]))&UnbiasedRNG[423])|((m[606]&~m[928]&~m[930]&m[931]&~m[932])|(~m[606]&~m[928]&~m[930]&~m[931]&m[932])|(m[606]&~m[928]&~m[930]&~m[931]&m[932])|(m[606]&m[928]&~m[930]&~m[931]&m[932])|(m[606]&~m[928]&m[930]&~m[931]&m[932])|(~m[606]&~m[928]&~m[930]&m[931]&m[932])|(m[606]&~m[928]&~m[930]&m[931]&m[932])|(~m[606]&m[928]&~m[930]&m[931]&m[932])|(m[606]&m[928]&~m[930]&m[931]&m[932])|(~m[606]&~m[928]&m[930]&m[931]&m[932])|(m[606]&~m[928]&m[930]&m[931]&m[932])|(m[606]&m[928]&m[930]&m[931]&m[932]));
    m[935] = (((m[897]&~m[933]&~m[934]&~m[936]&~m[937])|(~m[897]&~m[933]&~m[934]&m[936]&~m[937])|(m[897]&m[933]&~m[934]&m[936]&~m[937])|(m[897]&~m[933]&m[934]&m[936]&~m[937])|(~m[897]&m[933]&~m[934]&~m[936]&m[937])|(~m[897]&~m[933]&m[934]&~m[936]&m[937])|(m[897]&m[933]&m[934]&~m[936]&m[937])|(~m[897]&m[933]&m[934]&m[936]&m[937]))&UnbiasedRNG[424])|((m[897]&~m[933]&~m[934]&m[936]&~m[937])|(~m[897]&~m[933]&~m[934]&~m[936]&m[937])|(m[897]&~m[933]&~m[934]&~m[936]&m[937])|(m[897]&m[933]&~m[934]&~m[936]&m[937])|(m[897]&~m[933]&m[934]&~m[936]&m[937])|(~m[897]&~m[933]&~m[934]&m[936]&m[937])|(m[897]&~m[933]&~m[934]&m[936]&m[937])|(~m[897]&m[933]&~m[934]&m[936]&m[937])|(m[897]&m[933]&~m[934]&m[936]&m[937])|(~m[897]&~m[933]&m[934]&m[936]&m[937])|(m[897]&~m[933]&m[934]&m[936]&m[937])|(m[897]&m[933]&m[934]&m[936]&m[937]));
    m[940] = (((m[902]&~m[938]&~m[939]&~m[941]&~m[942])|(~m[902]&~m[938]&~m[939]&m[941]&~m[942])|(m[902]&m[938]&~m[939]&m[941]&~m[942])|(m[902]&~m[938]&m[939]&m[941]&~m[942])|(~m[902]&m[938]&~m[939]&~m[941]&m[942])|(~m[902]&~m[938]&m[939]&~m[941]&m[942])|(m[902]&m[938]&m[939]&~m[941]&m[942])|(~m[902]&m[938]&m[939]&m[941]&m[942]))&UnbiasedRNG[425])|((m[902]&~m[938]&~m[939]&m[941]&~m[942])|(~m[902]&~m[938]&~m[939]&~m[941]&m[942])|(m[902]&~m[938]&~m[939]&~m[941]&m[942])|(m[902]&m[938]&~m[939]&~m[941]&m[942])|(m[902]&~m[938]&m[939]&~m[941]&m[942])|(~m[902]&~m[938]&~m[939]&m[941]&m[942])|(m[902]&~m[938]&~m[939]&m[941]&m[942])|(~m[902]&m[938]&~m[939]&m[941]&m[942])|(m[902]&m[938]&~m[939]&m[941]&m[942])|(~m[902]&~m[938]&m[939]&m[941]&m[942])|(m[902]&~m[938]&m[939]&m[941]&m[942])|(m[902]&m[938]&m[939]&m[941]&m[942]));
    m[945] = (((m[907]&~m[943]&~m[944]&~m[946]&~m[947])|(~m[907]&~m[943]&~m[944]&m[946]&~m[947])|(m[907]&m[943]&~m[944]&m[946]&~m[947])|(m[907]&~m[943]&m[944]&m[946]&~m[947])|(~m[907]&m[943]&~m[944]&~m[946]&m[947])|(~m[907]&~m[943]&m[944]&~m[946]&m[947])|(m[907]&m[943]&m[944]&~m[946]&m[947])|(~m[907]&m[943]&m[944]&m[946]&m[947]))&UnbiasedRNG[426])|((m[907]&~m[943]&~m[944]&m[946]&~m[947])|(~m[907]&~m[943]&~m[944]&~m[946]&m[947])|(m[907]&~m[943]&~m[944]&~m[946]&m[947])|(m[907]&m[943]&~m[944]&~m[946]&m[947])|(m[907]&~m[943]&m[944]&~m[946]&m[947])|(~m[907]&~m[943]&~m[944]&m[946]&m[947])|(m[907]&~m[943]&~m[944]&m[946]&m[947])|(~m[907]&m[943]&~m[944]&m[946]&m[947])|(m[907]&m[943]&~m[944]&m[946]&m[947])|(~m[907]&~m[943]&m[944]&m[946]&m[947])|(m[907]&~m[943]&m[944]&m[946]&m[947])|(m[907]&m[943]&m[944]&m[946]&m[947]));
    m[955] = (((m[912]&~m[953]&~m[954]&~m[956]&~m[957])|(~m[912]&~m[953]&~m[954]&m[956]&~m[957])|(m[912]&m[953]&~m[954]&m[956]&~m[957])|(m[912]&~m[953]&m[954]&m[956]&~m[957])|(~m[912]&m[953]&~m[954]&~m[956]&m[957])|(~m[912]&~m[953]&m[954]&~m[956]&m[957])|(m[912]&m[953]&m[954]&~m[956]&m[957])|(~m[912]&m[953]&m[954]&m[956]&m[957]))&UnbiasedRNG[427])|((m[912]&~m[953]&~m[954]&m[956]&~m[957])|(~m[912]&~m[953]&~m[954]&~m[956]&m[957])|(m[912]&~m[953]&~m[954]&~m[956]&m[957])|(m[912]&m[953]&~m[954]&~m[956]&m[957])|(m[912]&~m[953]&m[954]&~m[956]&m[957])|(~m[912]&~m[953]&~m[954]&m[956]&m[957])|(m[912]&~m[953]&~m[954]&m[956]&m[957])|(~m[912]&m[953]&~m[954]&m[956]&m[957])|(m[912]&m[953]&~m[954]&m[956]&m[957])|(~m[912]&~m[953]&m[954]&m[956]&m[957])|(m[912]&~m[953]&m[954]&m[956]&m[957])|(m[912]&m[953]&m[954]&m[956]&m[957]));
    m[960] = (((m[917]&~m[958]&~m[959]&~m[961]&~m[962])|(~m[917]&~m[958]&~m[959]&m[961]&~m[962])|(m[917]&m[958]&~m[959]&m[961]&~m[962])|(m[917]&~m[958]&m[959]&m[961]&~m[962])|(~m[917]&m[958]&~m[959]&~m[961]&m[962])|(~m[917]&~m[958]&m[959]&~m[961]&m[962])|(m[917]&m[958]&m[959]&~m[961]&m[962])|(~m[917]&m[958]&m[959]&m[961]&m[962]))&UnbiasedRNG[428])|((m[917]&~m[958]&~m[959]&m[961]&~m[962])|(~m[917]&~m[958]&~m[959]&~m[961]&m[962])|(m[917]&~m[958]&~m[959]&~m[961]&m[962])|(m[917]&m[958]&~m[959]&~m[961]&m[962])|(m[917]&~m[958]&m[959]&~m[961]&m[962])|(~m[917]&~m[958]&~m[959]&m[961]&m[962])|(m[917]&~m[958]&~m[959]&m[961]&m[962])|(~m[917]&m[958]&~m[959]&m[961]&m[962])|(m[917]&m[958]&~m[959]&m[961]&m[962])|(~m[917]&~m[958]&m[959]&m[961]&m[962])|(m[917]&~m[958]&m[959]&m[961]&m[962])|(m[917]&m[958]&m[959]&m[961]&m[962]));
    m[965] = (((m[922]&~m[963]&~m[964]&~m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&m[966]&~m[967])|(m[922]&m[963]&~m[964]&m[966]&~m[967])|(m[922]&~m[963]&m[964]&m[966]&~m[967])|(~m[922]&m[963]&~m[964]&~m[966]&m[967])|(~m[922]&~m[963]&m[964]&~m[966]&m[967])|(m[922]&m[963]&m[964]&~m[966]&m[967])|(~m[922]&m[963]&m[964]&m[966]&m[967]))&UnbiasedRNG[429])|((m[922]&~m[963]&~m[964]&m[966]&~m[967])|(~m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&~m[964]&~m[966]&m[967])|(m[922]&m[963]&~m[964]&~m[966]&m[967])|(m[922]&~m[963]&m[964]&~m[966]&m[967])|(~m[922]&~m[963]&~m[964]&m[966]&m[967])|(m[922]&~m[963]&~m[964]&m[966]&m[967])|(~m[922]&m[963]&~m[964]&m[966]&m[967])|(m[922]&m[963]&~m[964]&m[966]&m[967])|(~m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&~m[963]&m[964]&m[966]&m[967])|(m[922]&m[963]&m[964]&m[966]&m[967]));
    m[970] = (((m[927]&~m[968]&~m[969]&~m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&m[971]&~m[972])|(m[927]&m[968]&~m[969]&m[971]&~m[972])|(m[927]&~m[968]&m[969]&m[971]&~m[972])|(~m[927]&m[968]&~m[969]&~m[971]&m[972])|(~m[927]&~m[968]&m[969]&~m[971]&m[972])|(m[927]&m[968]&m[969]&~m[971]&m[972])|(~m[927]&m[968]&m[969]&m[971]&m[972]))&UnbiasedRNG[430])|((m[927]&~m[968]&~m[969]&m[971]&~m[972])|(~m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&~m[969]&~m[971]&m[972])|(m[927]&m[968]&~m[969]&~m[971]&m[972])|(m[927]&~m[968]&m[969]&~m[971]&m[972])|(~m[927]&~m[968]&~m[969]&m[971]&m[972])|(m[927]&~m[968]&~m[969]&m[971]&m[972])|(~m[927]&m[968]&~m[969]&m[971]&m[972])|(m[927]&m[968]&~m[969]&m[971]&m[972])|(~m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&~m[968]&m[969]&m[971]&m[972])|(m[927]&m[968]&m[969]&m[971]&m[972]));
    m[974] = (((m[607]&~m[973]&~m[975]&~m[976]&~m[977])|(~m[607]&~m[973]&~m[975]&m[976]&~m[977])|(m[607]&m[973]&~m[975]&m[976]&~m[977])|(m[607]&~m[973]&m[975]&m[976]&~m[977])|(~m[607]&m[973]&~m[975]&~m[976]&m[977])|(~m[607]&~m[973]&m[975]&~m[976]&m[977])|(m[607]&m[973]&m[975]&~m[976]&m[977])|(~m[607]&m[973]&m[975]&m[976]&m[977]))&UnbiasedRNG[431])|((m[607]&~m[973]&~m[975]&m[976]&~m[977])|(~m[607]&~m[973]&~m[975]&~m[976]&m[977])|(m[607]&~m[973]&~m[975]&~m[976]&m[977])|(m[607]&m[973]&~m[975]&~m[976]&m[977])|(m[607]&~m[973]&m[975]&~m[976]&m[977])|(~m[607]&~m[973]&~m[975]&m[976]&m[977])|(m[607]&~m[973]&~m[975]&m[976]&m[977])|(~m[607]&m[973]&~m[975]&m[976]&m[977])|(m[607]&m[973]&~m[975]&m[976]&m[977])|(~m[607]&~m[973]&m[975]&m[976]&m[977])|(m[607]&~m[973]&m[975]&m[976]&m[977])|(m[607]&m[973]&m[975]&m[976]&m[977]));
    m[980] = (((m[937]&~m[978]&~m[979]&~m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&m[981]&~m[982])|(m[937]&m[978]&~m[979]&m[981]&~m[982])|(m[937]&~m[978]&m[979]&m[981]&~m[982])|(~m[937]&m[978]&~m[979]&~m[981]&m[982])|(~m[937]&~m[978]&m[979]&~m[981]&m[982])|(m[937]&m[978]&m[979]&~m[981]&m[982])|(~m[937]&m[978]&m[979]&m[981]&m[982]))&UnbiasedRNG[432])|((m[937]&~m[978]&~m[979]&m[981]&~m[982])|(~m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&~m[979]&~m[981]&m[982])|(m[937]&m[978]&~m[979]&~m[981]&m[982])|(m[937]&~m[978]&m[979]&~m[981]&m[982])|(~m[937]&~m[978]&~m[979]&m[981]&m[982])|(m[937]&~m[978]&~m[979]&m[981]&m[982])|(~m[937]&m[978]&~m[979]&m[981]&m[982])|(m[937]&m[978]&~m[979]&m[981]&m[982])|(~m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&~m[978]&m[979]&m[981]&m[982])|(m[937]&m[978]&m[979]&m[981]&m[982]));
    m[985] = (((m[942]&~m[983]&~m[984]&~m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&m[986]&~m[987])|(m[942]&m[983]&~m[984]&m[986]&~m[987])|(m[942]&~m[983]&m[984]&m[986]&~m[987])|(~m[942]&m[983]&~m[984]&~m[986]&m[987])|(~m[942]&~m[983]&m[984]&~m[986]&m[987])|(m[942]&m[983]&m[984]&~m[986]&m[987])|(~m[942]&m[983]&m[984]&m[986]&m[987]))&UnbiasedRNG[433])|((m[942]&~m[983]&~m[984]&m[986]&~m[987])|(~m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&~m[984]&~m[986]&m[987])|(m[942]&m[983]&~m[984]&~m[986]&m[987])|(m[942]&~m[983]&m[984]&~m[986]&m[987])|(~m[942]&~m[983]&~m[984]&m[986]&m[987])|(m[942]&~m[983]&~m[984]&m[986]&m[987])|(~m[942]&m[983]&~m[984]&m[986]&m[987])|(m[942]&m[983]&~m[984]&m[986]&m[987])|(~m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&~m[983]&m[984]&m[986]&m[987])|(m[942]&m[983]&m[984]&m[986]&m[987]));
    m[990] = (((m[947]&~m[988]&~m[989]&~m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&m[991]&~m[992])|(m[947]&m[988]&~m[989]&m[991]&~m[992])|(m[947]&~m[988]&m[989]&m[991]&~m[992])|(~m[947]&m[988]&~m[989]&~m[991]&m[992])|(~m[947]&~m[988]&m[989]&~m[991]&m[992])|(m[947]&m[988]&m[989]&~m[991]&m[992])|(~m[947]&m[988]&m[989]&m[991]&m[992]))&UnbiasedRNG[434])|((m[947]&~m[988]&~m[989]&m[991]&~m[992])|(~m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&~m[989]&~m[991]&m[992])|(m[947]&m[988]&~m[989]&~m[991]&m[992])|(m[947]&~m[988]&m[989]&~m[991]&m[992])|(~m[947]&~m[988]&~m[989]&m[991]&m[992])|(m[947]&~m[988]&~m[989]&m[991]&m[992])|(~m[947]&m[988]&~m[989]&m[991]&m[992])|(m[947]&m[988]&~m[989]&m[991]&m[992])|(~m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&~m[988]&m[989]&m[991]&m[992])|(m[947]&m[988]&m[989]&m[991]&m[992]));
    m[995] = (((m[952]&~m[993]&~m[994]&~m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&m[996]&~m[997])|(m[952]&m[993]&~m[994]&m[996]&~m[997])|(m[952]&~m[993]&m[994]&m[996]&~m[997])|(~m[952]&m[993]&~m[994]&~m[996]&m[997])|(~m[952]&~m[993]&m[994]&~m[996]&m[997])|(m[952]&m[993]&m[994]&~m[996]&m[997])|(~m[952]&m[993]&m[994]&m[996]&m[997]))&UnbiasedRNG[435])|((m[952]&~m[993]&~m[994]&m[996]&~m[997])|(~m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&~m[994]&~m[996]&m[997])|(m[952]&m[993]&~m[994]&~m[996]&m[997])|(m[952]&~m[993]&m[994]&~m[996]&m[997])|(~m[952]&~m[993]&~m[994]&m[996]&m[997])|(m[952]&~m[993]&~m[994]&m[996]&m[997])|(~m[952]&m[993]&~m[994]&m[996]&m[997])|(m[952]&m[993]&~m[994]&m[996]&m[997])|(~m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&~m[993]&m[994]&m[996]&m[997])|(m[952]&m[993]&m[994]&m[996]&m[997]));
    m[1005] = (((m[957]&~m[1003]&~m[1004]&~m[1006]&~m[1007])|(~m[957]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(m[957]&m[1003]&~m[1004]&m[1006]&~m[1007])|(m[957]&~m[1003]&m[1004]&m[1006]&~m[1007])|(~m[957]&m[1003]&~m[1004]&~m[1006]&m[1007])|(~m[957]&~m[1003]&m[1004]&~m[1006]&m[1007])|(m[957]&m[1003]&m[1004]&~m[1006]&m[1007])|(~m[957]&m[1003]&m[1004]&m[1006]&m[1007]))&UnbiasedRNG[436])|((m[957]&~m[1003]&~m[1004]&m[1006]&~m[1007])|(~m[957]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[957]&~m[1003]&~m[1004]&~m[1006]&m[1007])|(m[957]&m[1003]&~m[1004]&~m[1006]&m[1007])|(m[957]&~m[1003]&m[1004]&~m[1006]&m[1007])|(~m[957]&~m[1003]&~m[1004]&m[1006]&m[1007])|(m[957]&~m[1003]&~m[1004]&m[1006]&m[1007])|(~m[957]&m[1003]&~m[1004]&m[1006]&m[1007])|(m[957]&m[1003]&~m[1004]&m[1006]&m[1007])|(~m[957]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[957]&~m[1003]&m[1004]&m[1006]&m[1007])|(m[957]&m[1003]&m[1004]&m[1006]&m[1007]));
    m[1010] = (((m[962]&~m[1008]&~m[1009]&~m[1011]&~m[1012])|(~m[962]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(m[962]&m[1008]&~m[1009]&m[1011]&~m[1012])|(m[962]&~m[1008]&m[1009]&m[1011]&~m[1012])|(~m[962]&m[1008]&~m[1009]&~m[1011]&m[1012])|(~m[962]&~m[1008]&m[1009]&~m[1011]&m[1012])|(m[962]&m[1008]&m[1009]&~m[1011]&m[1012])|(~m[962]&m[1008]&m[1009]&m[1011]&m[1012]))&UnbiasedRNG[437])|((m[962]&~m[1008]&~m[1009]&m[1011]&~m[1012])|(~m[962]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[962]&~m[1008]&~m[1009]&~m[1011]&m[1012])|(m[962]&m[1008]&~m[1009]&~m[1011]&m[1012])|(m[962]&~m[1008]&m[1009]&~m[1011]&m[1012])|(~m[962]&~m[1008]&~m[1009]&m[1011]&m[1012])|(m[962]&~m[1008]&~m[1009]&m[1011]&m[1012])|(~m[962]&m[1008]&~m[1009]&m[1011]&m[1012])|(m[962]&m[1008]&~m[1009]&m[1011]&m[1012])|(~m[962]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[962]&~m[1008]&m[1009]&m[1011]&m[1012])|(m[962]&m[1008]&m[1009]&m[1011]&m[1012]));
    m[1015] = (((m[967]&~m[1013]&~m[1014]&~m[1016]&~m[1017])|(~m[967]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(m[967]&m[1013]&~m[1014]&m[1016]&~m[1017])|(m[967]&~m[1013]&m[1014]&m[1016]&~m[1017])|(~m[967]&m[1013]&~m[1014]&~m[1016]&m[1017])|(~m[967]&~m[1013]&m[1014]&~m[1016]&m[1017])|(m[967]&m[1013]&m[1014]&~m[1016]&m[1017])|(~m[967]&m[1013]&m[1014]&m[1016]&m[1017]))&UnbiasedRNG[438])|((m[967]&~m[1013]&~m[1014]&m[1016]&~m[1017])|(~m[967]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[967]&~m[1013]&~m[1014]&~m[1016]&m[1017])|(m[967]&m[1013]&~m[1014]&~m[1016]&m[1017])|(m[967]&~m[1013]&m[1014]&~m[1016]&m[1017])|(~m[967]&~m[1013]&~m[1014]&m[1016]&m[1017])|(m[967]&~m[1013]&~m[1014]&m[1016]&m[1017])|(~m[967]&m[1013]&~m[1014]&m[1016]&m[1017])|(m[967]&m[1013]&~m[1014]&m[1016]&m[1017])|(~m[967]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[967]&~m[1013]&m[1014]&m[1016]&m[1017])|(m[967]&m[1013]&m[1014]&m[1016]&m[1017]));
    m[1020] = (((m[972]&~m[1018]&~m[1019]&~m[1021]&~m[1022])|(~m[972]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(m[972]&m[1018]&~m[1019]&m[1021]&~m[1022])|(m[972]&~m[1018]&m[1019]&m[1021]&~m[1022])|(~m[972]&m[1018]&~m[1019]&~m[1021]&m[1022])|(~m[972]&~m[1018]&m[1019]&~m[1021]&m[1022])|(m[972]&m[1018]&m[1019]&~m[1021]&m[1022])|(~m[972]&m[1018]&m[1019]&m[1021]&m[1022]))&UnbiasedRNG[439])|((m[972]&~m[1018]&~m[1019]&m[1021]&~m[1022])|(~m[972]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[972]&~m[1018]&~m[1019]&~m[1021]&m[1022])|(m[972]&m[1018]&~m[1019]&~m[1021]&m[1022])|(m[972]&~m[1018]&m[1019]&~m[1021]&m[1022])|(~m[972]&~m[1018]&~m[1019]&m[1021]&m[1022])|(m[972]&~m[1018]&~m[1019]&m[1021]&m[1022])|(~m[972]&m[1018]&~m[1019]&m[1021]&m[1022])|(m[972]&m[1018]&~m[1019]&m[1021]&m[1022])|(~m[972]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[972]&~m[1018]&m[1019]&m[1021]&m[1022])|(m[972]&m[1018]&m[1019]&m[1021]&m[1022]));
    m[1025] = (((m[977]&~m[1023]&~m[1024]&~m[1026]&~m[1027])|(~m[977]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(m[977]&m[1023]&~m[1024]&m[1026]&~m[1027])|(m[977]&~m[1023]&m[1024]&m[1026]&~m[1027])|(~m[977]&m[1023]&~m[1024]&~m[1026]&m[1027])|(~m[977]&~m[1023]&m[1024]&~m[1026]&m[1027])|(m[977]&m[1023]&m[1024]&~m[1026]&m[1027])|(~m[977]&m[1023]&m[1024]&m[1026]&m[1027]))&UnbiasedRNG[440])|((m[977]&~m[1023]&~m[1024]&m[1026]&~m[1027])|(~m[977]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[977]&~m[1023]&~m[1024]&~m[1026]&m[1027])|(m[977]&m[1023]&~m[1024]&~m[1026]&m[1027])|(m[977]&~m[1023]&m[1024]&~m[1026]&m[1027])|(~m[977]&~m[1023]&~m[1024]&m[1026]&m[1027])|(m[977]&~m[1023]&~m[1024]&m[1026]&m[1027])|(~m[977]&m[1023]&~m[1024]&m[1026]&m[1027])|(m[977]&m[1023]&~m[1024]&m[1026]&m[1027])|(~m[977]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[977]&~m[1023]&m[1024]&m[1026]&m[1027])|(m[977]&m[1023]&m[1024]&m[1026]&m[1027]));
    m[1030] = (((m[982]&~m[1028]&~m[1029]&~m[1031]&~m[1032])|(~m[982]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(m[982]&m[1028]&~m[1029]&m[1031]&~m[1032])|(m[982]&~m[1028]&m[1029]&m[1031]&~m[1032])|(~m[982]&m[1028]&~m[1029]&~m[1031]&m[1032])|(~m[982]&~m[1028]&m[1029]&~m[1031]&m[1032])|(m[982]&m[1028]&m[1029]&~m[1031]&m[1032])|(~m[982]&m[1028]&m[1029]&m[1031]&m[1032]))&UnbiasedRNG[441])|((m[982]&~m[1028]&~m[1029]&m[1031]&~m[1032])|(~m[982]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[982]&~m[1028]&~m[1029]&~m[1031]&m[1032])|(m[982]&m[1028]&~m[1029]&~m[1031]&m[1032])|(m[982]&~m[1028]&m[1029]&~m[1031]&m[1032])|(~m[982]&~m[1028]&~m[1029]&m[1031]&m[1032])|(m[982]&~m[1028]&~m[1029]&m[1031]&m[1032])|(~m[982]&m[1028]&~m[1029]&m[1031]&m[1032])|(m[982]&m[1028]&~m[1029]&m[1031]&m[1032])|(~m[982]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[982]&~m[1028]&m[1029]&m[1031]&m[1032])|(m[982]&m[1028]&m[1029]&m[1031]&m[1032]));
    m[1035] = (((m[987]&~m[1033]&~m[1034]&~m[1036]&~m[1037])|(~m[987]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(m[987]&m[1033]&~m[1034]&m[1036]&~m[1037])|(m[987]&~m[1033]&m[1034]&m[1036]&~m[1037])|(~m[987]&m[1033]&~m[1034]&~m[1036]&m[1037])|(~m[987]&~m[1033]&m[1034]&~m[1036]&m[1037])|(m[987]&m[1033]&m[1034]&~m[1036]&m[1037])|(~m[987]&m[1033]&m[1034]&m[1036]&m[1037]))&UnbiasedRNG[442])|((m[987]&~m[1033]&~m[1034]&m[1036]&~m[1037])|(~m[987]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[987]&~m[1033]&~m[1034]&~m[1036]&m[1037])|(m[987]&m[1033]&~m[1034]&~m[1036]&m[1037])|(m[987]&~m[1033]&m[1034]&~m[1036]&m[1037])|(~m[987]&~m[1033]&~m[1034]&m[1036]&m[1037])|(m[987]&~m[1033]&~m[1034]&m[1036]&m[1037])|(~m[987]&m[1033]&~m[1034]&m[1036]&m[1037])|(m[987]&m[1033]&~m[1034]&m[1036]&m[1037])|(~m[987]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[987]&~m[1033]&m[1034]&m[1036]&m[1037])|(m[987]&m[1033]&m[1034]&m[1036]&m[1037]));
    m[1040] = (((m[992]&~m[1038]&~m[1039]&~m[1041]&~m[1042])|(~m[992]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(m[992]&m[1038]&~m[1039]&m[1041]&~m[1042])|(m[992]&~m[1038]&m[1039]&m[1041]&~m[1042])|(~m[992]&m[1038]&~m[1039]&~m[1041]&m[1042])|(~m[992]&~m[1038]&m[1039]&~m[1041]&m[1042])|(m[992]&m[1038]&m[1039]&~m[1041]&m[1042])|(~m[992]&m[1038]&m[1039]&m[1041]&m[1042]))&UnbiasedRNG[443])|((m[992]&~m[1038]&~m[1039]&m[1041]&~m[1042])|(~m[992]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[992]&~m[1038]&~m[1039]&~m[1041]&m[1042])|(m[992]&m[1038]&~m[1039]&~m[1041]&m[1042])|(m[992]&~m[1038]&m[1039]&~m[1041]&m[1042])|(~m[992]&~m[1038]&~m[1039]&m[1041]&m[1042])|(m[992]&~m[1038]&~m[1039]&m[1041]&m[1042])|(~m[992]&m[1038]&~m[1039]&m[1041]&m[1042])|(m[992]&m[1038]&~m[1039]&m[1041]&m[1042])|(~m[992]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[992]&~m[1038]&m[1039]&m[1041]&m[1042])|(m[992]&m[1038]&m[1039]&m[1041]&m[1042]));
    m[1045] = (((m[997]&~m[1043]&~m[1044]&~m[1046]&~m[1047])|(~m[997]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(m[997]&m[1043]&~m[1044]&m[1046]&~m[1047])|(m[997]&~m[1043]&m[1044]&m[1046]&~m[1047])|(~m[997]&m[1043]&~m[1044]&~m[1046]&m[1047])|(~m[997]&~m[1043]&m[1044]&~m[1046]&m[1047])|(m[997]&m[1043]&m[1044]&~m[1046]&m[1047])|(~m[997]&m[1043]&m[1044]&m[1046]&m[1047]))&UnbiasedRNG[444])|((m[997]&~m[1043]&~m[1044]&m[1046]&~m[1047])|(~m[997]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[997]&~m[1043]&~m[1044]&~m[1046]&m[1047])|(m[997]&m[1043]&~m[1044]&~m[1046]&m[1047])|(m[997]&~m[1043]&m[1044]&~m[1046]&m[1047])|(~m[997]&~m[1043]&~m[1044]&m[1046]&m[1047])|(m[997]&~m[1043]&~m[1044]&m[1046]&m[1047])|(~m[997]&m[1043]&~m[1044]&m[1046]&m[1047])|(m[997]&m[1043]&~m[1044]&m[1046]&m[1047])|(~m[997]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[997]&~m[1043]&m[1044]&m[1046]&m[1047])|(m[997]&m[1043]&m[1044]&m[1046]&m[1047]));
    m[1050] = (((m[1002]&~m[1048]&~m[1049]&~m[1051]&~m[1052])|(~m[1002]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1002]&m[1048]&~m[1049]&m[1051]&~m[1052])|(m[1002]&~m[1048]&m[1049]&m[1051]&~m[1052])|(~m[1002]&m[1048]&~m[1049]&~m[1051]&m[1052])|(~m[1002]&~m[1048]&m[1049]&~m[1051]&m[1052])|(m[1002]&m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1002]&m[1048]&m[1049]&m[1051]&m[1052]))&UnbiasedRNG[445])|((m[1002]&~m[1048]&~m[1049]&m[1051]&~m[1052])|(~m[1002]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1002]&~m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1002]&m[1048]&~m[1049]&~m[1051]&m[1052])|(m[1002]&~m[1048]&m[1049]&~m[1051]&m[1052])|(~m[1002]&~m[1048]&~m[1049]&m[1051]&m[1052])|(m[1002]&~m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1002]&m[1048]&~m[1049]&m[1051]&m[1052])|(m[1002]&m[1048]&~m[1049]&m[1051]&m[1052])|(~m[1002]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1002]&~m[1048]&m[1049]&m[1051]&m[1052])|(m[1002]&m[1048]&m[1049]&m[1051]&m[1052]));
    m[1060] = (((m[1007]&~m[1058]&~m[1059]&~m[1061]&~m[1062])|(~m[1007]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1007]&m[1058]&~m[1059]&m[1061]&~m[1062])|(m[1007]&~m[1058]&m[1059]&m[1061]&~m[1062])|(~m[1007]&m[1058]&~m[1059]&~m[1061]&m[1062])|(~m[1007]&~m[1058]&m[1059]&~m[1061]&m[1062])|(m[1007]&m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1007]&m[1058]&m[1059]&m[1061]&m[1062]))&UnbiasedRNG[446])|((m[1007]&~m[1058]&~m[1059]&m[1061]&~m[1062])|(~m[1007]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1007]&~m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1007]&m[1058]&~m[1059]&~m[1061]&m[1062])|(m[1007]&~m[1058]&m[1059]&~m[1061]&m[1062])|(~m[1007]&~m[1058]&~m[1059]&m[1061]&m[1062])|(m[1007]&~m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1007]&m[1058]&~m[1059]&m[1061]&m[1062])|(m[1007]&m[1058]&~m[1059]&m[1061]&m[1062])|(~m[1007]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1007]&~m[1058]&m[1059]&m[1061]&m[1062])|(m[1007]&m[1058]&m[1059]&m[1061]&m[1062]));
    m[1065] = (((m[1012]&~m[1063]&~m[1064]&~m[1066]&~m[1067])|(~m[1012]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1012]&m[1063]&~m[1064]&m[1066]&~m[1067])|(m[1012]&~m[1063]&m[1064]&m[1066]&~m[1067])|(~m[1012]&m[1063]&~m[1064]&~m[1066]&m[1067])|(~m[1012]&~m[1063]&m[1064]&~m[1066]&m[1067])|(m[1012]&m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1012]&m[1063]&m[1064]&m[1066]&m[1067]))&UnbiasedRNG[447])|((m[1012]&~m[1063]&~m[1064]&m[1066]&~m[1067])|(~m[1012]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1012]&~m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1012]&m[1063]&~m[1064]&~m[1066]&m[1067])|(m[1012]&~m[1063]&m[1064]&~m[1066]&m[1067])|(~m[1012]&~m[1063]&~m[1064]&m[1066]&m[1067])|(m[1012]&~m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1012]&m[1063]&~m[1064]&m[1066]&m[1067])|(m[1012]&m[1063]&~m[1064]&m[1066]&m[1067])|(~m[1012]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1012]&~m[1063]&m[1064]&m[1066]&m[1067])|(m[1012]&m[1063]&m[1064]&m[1066]&m[1067]));
    m[1070] = (((m[1017]&~m[1068]&~m[1069]&~m[1071]&~m[1072])|(~m[1017]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1017]&m[1068]&~m[1069]&m[1071]&~m[1072])|(m[1017]&~m[1068]&m[1069]&m[1071]&~m[1072])|(~m[1017]&m[1068]&~m[1069]&~m[1071]&m[1072])|(~m[1017]&~m[1068]&m[1069]&~m[1071]&m[1072])|(m[1017]&m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1017]&m[1068]&m[1069]&m[1071]&m[1072]))&UnbiasedRNG[448])|((m[1017]&~m[1068]&~m[1069]&m[1071]&~m[1072])|(~m[1017]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1017]&~m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1017]&m[1068]&~m[1069]&~m[1071]&m[1072])|(m[1017]&~m[1068]&m[1069]&~m[1071]&m[1072])|(~m[1017]&~m[1068]&~m[1069]&m[1071]&m[1072])|(m[1017]&~m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1017]&m[1068]&~m[1069]&m[1071]&m[1072])|(m[1017]&m[1068]&~m[1069]&m[1071]&m[1072])|(~m[1017]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1017]&~m[1068]&m[1069]&m[1071]&m[1072])|(m[1017]&m[1068]&m[1069]&m[1071]&m[1072]));
    m[1075] = (((m[1022]&~m[1073]&~m[1074]&~m[1076]&~m[1077])|(~m[1022]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1022]&m[1073]&~m[1074]&m[1076]&~m[1077])|(m[1022]&~m[1073]&m[1074]&m[1076]&~m[1077])|(~m[1022]&m[1073]&~m[1074]&~m[1076]&m[1077])|(~m[1022]&~m[1073]&m[1074]&~m[1076]&m[1077])|(m[1022]&m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1022]&m[1073]&m[1074]&m[1076]&m[1077]))&UnbiasedRNG[449])|((m[1022]&~m[1073]&~m[1074]&m[1076]&~m[1077])|(~m[1022]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1022]&~m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1022]&m[1073]&~m[1074]&~m[1076]&m[1077])|(m[1022]&~m[1073]&m[1074]&~m[1076]&m[1077])|(~m[1022]&~m[1073]&~m[1074]&m[1076]&m[1077])|(m[1022]&~m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1022]&m[1073]&~m[1074]&m[1076]&m[1077])|(m[1022]&m[1073]&~m[1074]&m[1076]&m[1077])|(~m[1022]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1022]&~m[1073]&m[1074]&m[1076]&m[1077])|(m[1022]&m[1073]&m[1074]&m[1076]&m[1077]));
    m[1080] = (((m[1027]&~m[1078]&~m[1079]&~m[1081]&~m[1082])|(~m[1027]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1027]&m[1078]&~m[1079]&m[1081]&~m[1082])|(m[1027]&~m[1078]&m[1079]&m[1081]&~m[1082])|(~m[1027]&m[1078]&~m[1079]&~m[1081]&m[1082])|(~m[1027]&~m[1078]&m[1079]&~m[1081]&m[1082])|(m[1027]&m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1027]&m[1078]&m[1079]&m[1081]&m[1082]))&UnbiasedRNG[450])|((m[1027]&~m[1078]&~m[1079]&m[1081]&~m[1082])|(~m[1027]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1027]&~m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1027]&m[1078]&~m[1079]&~m[1081]&m[1082])|(m[1027]&~m[1078]&m[1079]&~m[1081]&m[1082])|(~m[1027]&~m[1078]&~m[1079]&m[1081]&m[1082])|(m[1027]&~m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1027]&m[1078]&~m[1079]&m[1081]&m[1082])|(m[1027]&m[1078]&~m[1079]&m[1081]&m[1082])|(~m[1027]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1027]&~m[1078]&m[1079]&m[1081]&m[1082])|(m[1027]&m[1078]&m[1079]&m[1081]&m[1082]));
    m[1085] = (((m[1032]&~m[1083]&~m[1084]&~m[1086]&~m[1087])|(~m[1032]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1032]&m[1083]&~m[1084]&m[1086]&~m[1087])|(m[1032]&~m[1083]&m[1084]&m[1086]&~m[1087])|(~m[1032]&m[1083]&~m[1084]&~m[1086]&m[1087])|(~m[1032]&~m[1083]&m[1084]&~m[1086]&m[1087])|(m[1032]&m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1032]&m[1083]&m[1084]&m[1086]&m[1087]))&UnbiasedRNG[451])|((m[1032]&~m[1083]&~m[1084]&m[1086]&~m[1087])|(~m[1032]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1032]&~m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1032]&m[1083]&~m[1084]&~m[1086]&m[1087])|(m[1032]&~m[1083]&m[1084]&~m[1086]&m[1087])|(~m[1032]&~m[1083]&~m[1084]&m[1086]&m[1087])|(m[1032]&~m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1032]&m[1083]&~m[1084]&m[1086]&m[1087])|(m[1032]&m[1083]&~m[1084]&m[1086]&m[1087])|(~m[1032]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1032]&~m[1083]&m[1084]&m[1086]&m[1087])|(m[1032]&m[1083]&m[1084]&m[1086]&m[1087]));
    m[1090] = (((m[1037]&~m[1088]&~m[1089]&~m[1091]&~m[1092])|(~m[1037]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1037]&m[1088]&~m[1089]&m[1091]&~m[1092])|(m[1037]&~m[1088]&m[1089]&m[1091]&~m[1092])|(~m[1037]&m[1088]&~m[1089]&~m[1091]&m[1092])|(~m[1037]&~m[1088]&m[1089]&~m[1091]&m[1092])|(m[1037]&m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1037]&m[1088]&m[1089]&m[1091]&m[1092]))&UnbiasedRNG[452])|((m[1037]&~m[1088]&~m[1089]&m[1091]&~m[1092])|(~m[1037]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1037]&~m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1037]&m[1088]&~m[1089]&~m[1091]&m[1092])|(m[1037]&~m[1088]&m[1089]&~m[1091]&m[1092])|(~m[1037]&~m[1088]&~m[1089]&m[1091]&m[1092])|(m[1037]&~m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1037]&m[1088]&~m[1089]&m[1091]&m[1092])|(m[1037]&m[1088]&~m[1089]&m[1091]&m[1092])|(~m[1037]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1037]&~m[1088]&m[1089]&m[1091]&m[1092])|(m[1037]&m[1088]&m[1089]&m[1091]&m[1092]));
    m[1095] = (((m[1042]&~m[1093]&~m[1094]&~m[1096]&~m[1097])|(~m[1042]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1042]&m[1093]&~m[1094]&m[1096]&~m[1097])|(m[1042]&~m[1093]&m[1094]&m[1096]&~m[1097])|(~m[1042]&m[1093]&~m[1094]&~m[1096]&m[1097])|(~m[1042]&~m[1093]&m[1094]&~m[1096]&m[1097])|(m[1042]&m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1042]&m[1093]&m[1094]&m[1096]&m[1097]))&UnbiasedRNG[453])|((m[1042]&~m[1093]&~m[1094]&m[1096]&~m[1097])|(~m[1042]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1042]&~m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1042]&m[1093]&~m[1094]&~m[1096]&m[1097])|(m[1042]&~m[1093]&m[1094]&~m[1096]&m[1097])|(~m[1042]&~m[1093]&~m[1094]&m[1096]&m[1097])|(m[1042]&~m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1042]&m[1093]&~m[1094]&m[1096]&m[1097])|(m[1042]&m[1093]&~m[1094]&m[1096]&m[1097])|(~m[1042]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1042]&~m[1093]&m[1094]&m[1096]&m[1097])|(m[1042]&m[1093]&m[1094]&m[1096]&m[1097]));
    m[1100] = (((m[1047]&~m[1098]&~m[1099]&~m[1101]&~m[1102])|(~m[1047]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1047]&m[1098]&~m[1099]&m[1101]&~m[1102])|(m[1047]&~m[1098]&m[1099]&m[1101]&~m[1102])|(~m[1047]&m[1098]&~m[1099]&~m[1101]&m[1102])|(~m[1047]&~m[1098]&m[1099]&~m[1101]&m[1102])|(m[1047]&m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1047]&m[1098]&m[1099]&m[1101]&m[1102]))&UnbiasedRNG[454])|((m[1047]&~m[1098]&~m[1099]&m[1101]&~m[1102])|(~m[1047]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1047]&~m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1047]&m[1098]&~m[1099]&~m[1101]&m[1102])|(m[1047]&~m[1098]&m[1099]&~m[1101]&m[1102])|(~m[1047]&~m[1098]&~m[1099]&m[1101]&m[1102])|(m[1047]&~m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1047]&m[1098]&~m[1099]&m[1101]&m[1102])|(m[1047]&m[1098]&~m[1099]&m[1101]&m[1102])|(~m[1047]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1047]&~m[1098]&m[1099]&m[1101]&m[1102])|(m[1047]&m[1098]&m[1099]&m[1101]&m[1102]));
    m[1105] = (((m[1052]&~m[1103]&~m[1104]&~m[1106]&~m[1107])|(~m[1052]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1052]&m[1103]&~m[1104]&m[1106]&~m[1107])|(m[1052]&~m[1103]&m[1104]&m[1106]&~m[1107])|(~m[1052]&m[1103]&~m[1104]&~m[1106]&m[1107])|(~m[1052]&~m[1103]&m[1104]&~m[1106]&m[1107])|(m[1052]&m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1052]&m[1103]&m[1104]&m[1106]&m[1107]))&UnbiasedRNG[455])|((m[1052]&~m[1103]&~m[1104]&m[1106]&~m[1107])|(~m[1052]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1052]&~m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1052]&m[1103]&~m[1104]&~m[1106]&m[1107])|(m[1052]&~m[1103]&m[1104]&~m[1106]&m[1107])|(~m[1052]&~m[1103]&~m[1104]&m[1106]&m[1107])|(m[1052]&~m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1052]&m[1103]&~m[1104]&m[1106]&m[1107])|(m[1052]&m[1103]&~m[1104]&m[1106]&m[1107])|(~m[1052]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1052]&~m[1103]&m[1104]&m[1106]&m[1107])|(m[1052]&m[1103]&m[1104]&m[1106]&m[1107]));
    m[1110] = (((m[1057]&~m[1108]&~m[1109]&~m[1111]&~m[1112])|(~m[1057]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1057]&m[1108]&~m[1109]&m[1111]&~m[1112])|(m[1057]&~m[1108]&m[1109]&m[1111]&~m[1112])|(~m[1057]&m[1108]&~m[1109]&~m[1111]&m[1112])|(~m[1057]&~m[1108]&m[1109]&~m[1111]&m[1112])|(m[1057]&m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1057]&m[1108]&m[1109]&m[1111]&m[1112]))&UnbiasedRNG[456])|((m[1057]&~m[1108]&~m[1109]&m[1111]&~m[1112])|(~m[1057]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1057]&~m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1057]&m[1108]&~m[1109]&~m[1111]&m[1112])|(m[1057]&~m[1108]&m[1109]&~m[1111]&m[1112])|(~m[1057]&~m[1108]&~m[1109]&m[1111]&m[1112])|(m[1057]&~m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1057]&m[1108]&~m[1109]&m[1111]&m[1112])|(m[1057]&m[1108]&~m[1109]&m[1111]&m[1112])|(~m[1057]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1057]&~m[1108]&m[1109]&m[1111]&m[1112])|(m[1057]&m[1108]&m[1109]&m[1111]&m[1112]));
    m[1120] = (((m[1062]&~m[1118]&~m[1119]&~m[1121]&~m[1122])|(~m[1062]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1062]&m[1118]&~m[1119]&m[1121]&~m[1122])|(m[1062]&~m[1118]&m[1119]&m[1121]&~m[1122])|(~m[1062]&m[1118]&~m[1119]&~m[1121]&m[1122])|(~m[1062]&~m[1118]&m[1119]&~m[1121]&m[1122])|(m[1062]&m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1062]&m[1118]&m[1119]&m[1121]&m[1122]))&UnbiasedRNG[457])|((m[1062]&~m[1118]&~m[1119]&m[1121]&~m[1122])|(~m[1062]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1062]&~m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1062]&m[1118]&~m[1119]&~m[1121]&m[1122])|(m[1062]&~m[1118]&m[1119]&~m[1121]&m[1122])|(~m[1062]&~m[1118]&~m[1119]&m[1121]&m[1122])|(m[1062]&~m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1062]&m[1118]&~m[1119]&m[1121]&m[1122])|(m[1062]&m[1118]&~m[1119]&m[1121]&m[1122])|(~m[1062]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1062]&~m[1118]&m[1119]&m[1121]&m[1122])|(m[1062]&m[1118]&m[1119]&m[1121]&m[1122]));
    m[1125] = (((m[1067]&~m[1123]&~m[1124]&~m[1126]&~m[1127])|(~m[1067]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1067]&m[1123]&~m[1124]&m[1126]&~m[1127])|(m[1067]&~m[1123]&m[1124]&m[1126]&~m[1127])|(~m[1067]&m[1123]&~m[1124]&~m[1126]&m[1127])|(~m[1067]&~m[1123]&m[1124]&~m[1126]&m[1127])|(m[1067]&m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1067]&m[1123]&m[1124]&m[1126]&m[1127]))&UnbiasedRNG[458])|((m[1067]&~m[1123]&~m[1124]&m[1126]&~m[1127])|(~m[1067]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1067]&~m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1067]&m[1123]&~m[1124]&~m[1126]&m[1127])|(m[1067]&~m[1123]&m[1124]&~m[1126]&m[1127])|(~m[1067]&~m[1123]&~m[1124]&m[1126]&m[1127])|(m[1067]&~m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1067]&m[1123]&~m[1124]&m[1126]&m[1127])|(m[1067]&m[1123]&~m[1124]&m[1126]&m[1127])|(~m[1067]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1067]&~m[1123]&m[1124]&m[1126]&m[1127])|(m[1067]&m[1123]&m[1124]&m[1126]&m[1127]));
    m[1130] = (((m[1072]&~m[1128]&~m[1129]&~m[1131]&~m[1132])|(~m[1072]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1072]&m[1128]&~m[1129]&m[1131]&~m[1132])|(m[1072]&~m[1128]&m[1129]&m[1131]&~m[1132])|(~m[1072]&m[1128]&~m[1129]&~m[1131]&m[1132])|(~m[1072]&~m[1128]&m[1129]&~m[1131]&m[1132])|(m[1072]&m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1072]&m[1128]&m[1129]&m[1131]&m[1132]))&UnbiasedRNG[459])|((m[1072]&~m[1128]&~m[1129]&m[1131]&~m[1132])|(~m[1072]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1072]&~m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1072]&m[1128]&~m[1129]&~m[1131]&m[1132])|(m[1072]&~m[1128]&m[1129]&~m[1131]&m[1132])|(~m[1072]&~m[1128]&~m[1129]&m[1131]&m[1132])|(m[1072]&~m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1072]&m[1128]&~m[1129]&m[1131]&m[1132])|(m[1072]&m[1128]&~m[1129]&m[1131]&m[1132])|(~m[1072]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1072]&~m[1128]&m[1129]&m[1131]&m[1132])|(m[1072]&m[1128]&m[1129]&m[1131]&m[1132]));
    m[1135] = (((m[1077]&~m[1133]&~m[1134]&~m[1136]&~m[1137])|(~m[1077]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1077]&m[1133]&~m[1134]&m[1136]&~m[1137])|(m[1077]&~m[1133]&m[1134]&m[1136]&~m[1137])|(~m[1077]&m[1133]&~m[1134]&~m[1136]&m[1137])|(~m[1077]&~m[1133]&m[1134]&~m[1136]&m[1137])|(m[1077]&m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1077]&m[1133]&m[1134]&m[1136]&m[1137]))&UnbiasedRNG[460])|((m[1077]&~m[1133]&~m[1134]&m[1136]&~m[1137])|(~m[1077]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1077]&~m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1077]&m[1133]&~m[1134]&~m[1136]&m[1137])|(m[1077]&~m[1133]&m[1134]&~m[1136]&m[1137])|(~m[1077]&~m[1133]&~m[1134]&m[1136]&m[1137])|(m[1077]&~m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1077]&m[1133]&~m[1134]&m[1136]&m[1137])|(m[1077]&m[1133]&~m[1134]&m[1136]&m[1137])|(~m[1077]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1077]&~m[1133]&m[1134]&m[1136]&m[1137])|(m[1077]&m[1133]&m[1134]&m[1136]&m[1137]));
    m[1140] = (((m[1082]&~m[1138]&~m[1139]&~m[1141]&~m[1142])|(~m[1082]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1082]&m[1138]&~m[1139]&m[1141]&~m[1142])|(m[1082]&~m[1138]&m[1139]&m[1141]&~m[1142])|(~m[1082]&m[1138]&~m[1139]&~m[1141]&m[1142])|(~m[1082]&~m[1138]&m[1139]&~m[1141]&m[1142])|(m[1082]&m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1082]&m[1138]&m[1139]&m[1141]&m[1142]))&UnbiasedRNG[461])|((m[1082]&~m[1138]&~m[1139]&m[1141]&~m[1142])|(~m[1082]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1082]&~m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1082]&m[1138]&~m[1139]&~m[1141]&m[1142])|(m[1082]&~m[1138]&m[1139]&~m[1141]&m[1142])|(~m[1082]&~m[1138]&~m[1139]&m[1141]&m[1142])|(m[1082]&~m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1082]&m[1138]&~m[1139]&m[1141]&m[1142])|(m[1082]&m[1138]&~m[1139]&m[1141]&m[1142])|(~m[1082]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1082]&~m[1138]&m[1139]&m[1141]&m[1142])|(m[1082]&m[1138]&m[1139]&m[1141]&m[1142]));
    m[1145] = (((m[1087]&~m[1143]&~m[1144]&~m[1146]&~m[1147])|(~m[1087]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1087]&m[1143]&~m[1144]&m[1146]&~m[1147])|(m[1087]&~m[1143]&m[1144]&m[1146]&~m[1147])|(~m[1087]&m[1143]&~m[1144]&~m[1146]&m[1147])|(~m[1087]&~m[1143]&m[1144]&~m[1146]&m[1147])|(m[1087]&m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1087]&m[1143]&m[1144]&m[1146]&m[1147]))&UnbiasedRNG[462])|((m[1087]&~m[1143]&~m[1144]&m[1146]&~m[1147])|(~m[1087]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1087]&~m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1087]&m[1143]&~m[1144]&~m[1146]&m[1147])|(m[1087]&~m[1143]&m[1144]&~m[1146]&m[1147])|(~m[1087]&~m[1143]&~m[1144]&m[1146]&m[1147])|(m[1087]&~m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1087]&m[1143]&~m[1144]&m[1146]&m[1147])|(m[1087]&m[1143]&~m[1144]&m[1146]&m[1147])|(~m[1087]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1087]&~m[1143]&m[1144]&m[1146]&m[1147])|(m[1087]&m[1143]&m[1144]&m[1146]&m[1147]));
    m[1150] = (((m[1092]&~m[1148]&~m[1149]&~m[1151]&~m[1152])|(~m[1092]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1092]&m[1148]&~m[1149]&m[1151]&~m[1152])|(m[1092]&~m[1148]&m[1149]&m[1151]&~m[1152])|(~m[1092]&m[1148]&~m[1149]&~m[1151]&m[1152])|(~m[1092]&~m[1148]&m[1149]&~m[1151]&m[1152])|(m[1092]&m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1092]&m[1148]&m[1149]&m[1151]&m[1152]))&UnbiasedRNG[463])|((m[1092]&~m[1148]&~m[1149]&m[1151]&~m[1152])|(~m[1092]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1092]&~m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1092]&m[1148]&~m[1149]&~m[1151]&m[1152])|(m[1092]&~m[1148]&m[1149]&~m[1151]&m[1152])|(~m[1092]&~m[1148]&~m[1149]&m[1151]&m[1152])|(m[1092]&~m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1092]&m[1148]&~m[1149]&m[1151]&m[1152])|(m[1092]&m[1148]&~m[1149]&m[1151]&m[1152])|(~m[1092]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1092]&~m[1148]&m[1149]&m[1151]&m[1152])|(m[1092]&m[1148]&m[1149]&m[1151]&m[1152]));
    m[1155] = (((m[1097]&~m[1153]&~m[1154]&~m[1156]&~m[1157])|(~m[1097]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1097]&m[1153]&~m[1154]&m[1156]&~m[1157])|(m[1097]&~m[1153]&m[1154]&m[1156]&~m[1157])|(~m[1097]&m[1153]&~m[1154]&~m[1156]&m[1157])|(~m[1097]&~m[1153]&m[1154]&~m[1156]&m[1157])|(m[1097]&m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1097]&m[1153]&m[1154]&m[1156]&m[1157]))&UnbiasedRNG[464])|((m[1097]&~m[1153]&~m[1154]&m[1156]&~m[1157])|(~m[1097]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1097]&~m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1097]&m[1153]&~m[1154]&~m[1156]&m[1157])|(m[1097]&~m[1153]&m[1154]&~m[1156]&m[1157])|(~m[1097]&~m[1153]&~m[1154]&m[1156]&m[1157])|(m[1097]&~m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1097]&m[1153]&~m[1154]&m[1156]&m[1157])|(m[1097]&m[1153]&~m[1154]&m[1156]&m[1157])|(~m[1097]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1097]&~m[1153]&m[1154]&m[1156]&m[1157])|(m[1097]&m[1153]&m[1154]&m[1156]&m[1157]));
    m[1160] = (((m[1102]&~m[1158]&~m[1159]&~m[1161]&~m[1162])|(~m[1102]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1102]&m[1158]&~m[1159]&m[1161]&~m[1162])|(m[1102]&~m[1158]&m[1159]&m[1161]&~m[1162])|(~m[1102]&m[1158]&~m[1159]&~m[1161]&m[1162])|(~m[1102]&~m[1158]&m[1159]&~m[1161]&m[1162])|(m[1102]&m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1102]&m[1158]&m[1159]&m[1161]&m[1162]))&UnbiasedRNG[465])|((m[1102]&~m[1158]&~m[1159]&m[1161]&~m[1162])|(~m[1102]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1102]&~m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1102]&m[1158]&~m[1159]&~m[1161]&m[1162])|(m[1102]&~m[1158]&m[1159]&~m[1161]&m[1162])|(~m[1102]&~m[1158]&~m[1159]&m[1161]&m[1162])|(m[1102]&~m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1102]&m[1158]&~m[1159]&m[1161]&m[1162])|(m[1102]&m[1158]&~m[1159]&m[1161]&m[1162])|(~m[1102]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1102]&~m[1158]&m[1159]&m[1161]&m[1162])|(m[1102]&m[1158]&m[1159]&m[1161]&m[1162]));
    m[1165] = (((m[1107]&~m[1163]&~m[1164]&~m[1166]&~m[1167])|(~m[1107]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1107]&m[1163]&~m[1164]&m[1166]&~m[1167])|(m[1107]&~m[1163]&m[1164]&m[1166]&~m[1167])|(~m[1107]&m[1163]&~m[1164]&~m[1166]&m[1167])|(~m[1107]&~m[1163]&m[1164]&~m[1166]&m[1167])|(m[1107]&m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1107]&m[1163]&m[1164]&m[1166]&m[1167]))&UnbiasedRNG[466])|((m[1107]&~m[1163]&~m[1164]&m[1166]&~m[1167])|(~m[1107]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1107]&~m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1107]&m[1163]&~m[1164]&~m[1166]&m[1167])|(m[1107]&~m[1163]&m[1164]&~m[1166]&m[1167])|(~m[1107]&~m[1163]&~m[1164]&m[1166]&m[1167])|(m[1107]&~m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1107]&m[1163]&~m[1164]&m[1166]&m[1167])|(m[1107]&m[1163]&~m[1164]&m[1166]&m[1167])|(~m[1107]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1107]&~m[1163]&m[1164]&m[1166]&m[1167])|(m[1107]&m[1163]&m[1164]&m[1166]&m[1167]));
    m[1170] = (((m[1112]&~m[1168]&~m[1169]&~m[1171]&~m[1172])|(~m[1112]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1112]&m[1168]&~m[1169]&m[1171]&~m[1172])|(m[1112]&~m[1168]&m[1169]&m[1171]&~m[1172])|(~m[1112]&m[1168]&~m[1169]&~m[1171]&m[1172])|(~m[1112]&~m[1168]&m[1169]&~m[1171]&m[1172])|(m[1112]&m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1112]&m[1168]&m[1169]&m[1171]&m[1172]))&UnbiasedRNG[467])|((m[1112]&~m[1168]&~m[1169]&m[1171]&~m[1172])|(~m[1112]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1112]&~m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1112]&m[1168]&~m[1169]&~m[1171]&m[1172])|(m[1112]&~m[1168]&m[1169]&~m[1171]&m[1172])|(~m[1112]&~m[1168]&~m[1169]&m[1171]&m[1172])|(m[1112]&~m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1112]&m[1168]&~m[1169]&m[1171]&m[1172])|(m[1112]&m[1168]&~m[1169]&m[1171]&m[1172])|(~m[1112]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1112]&~m[1168]&m[1169]&m[1171]&m[1172])|(m[1112]&m[1168]&m[1169]&m[1171]&m[1172]));
    m[1175] = (((m[1117]&~m[1173]&~m[1174]&~m[1176]&~m[1177])|(~m[1117]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1117]&m[1173]&~m[1174]&m[1176]&~m[1177])|(m[1117]&~m[1173]&m[1174]&m[1176]&~m[1177])|(~m[1117]&m[1173]&~m[1174]&~m[1176]&m[1177])|(~m[1117]&~m[1173]&m[1174]&~m[1176]&m[1177])|(m[1117]&m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1117]&m[1173]&m[1174]&m[1176]&m[1177]))&UnbiasedRNG[468])|((m[1117]&~m[1173]&~m[1174]&m[1176]&~m[1177])|(~m[1117]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1117]&~m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1117]&m[1173]&~m[1174]&~m[1176]&m[1177])|(m[1117]&~m[1173]&m[1174]&~m[1176]&m[1177])|(~m[1117]&~m[1173]&~m[1174]&m[1176]&m[1177])|(m[1117]&~m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1117]&m[1173]&~m[1174]&m[1176]&m[1177])|(m[1117]&m[1173]&~m[1174]&m[1176]&m[1177])|(~m[1117]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1117]&~m[1173]&m[1174]&m[1176]&m[1177])|(m[1117]&m[1173]&m[1174]&m[1176]&m[1177]));
    m[1185] = (((m[1122]&~m[1183]&~m[1184]&~m[1186]&~m[1187])|(~m[1122]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1122]&m[1183]&~m[1184]&m[1186]&~m[1187])|(m[1122]&~m[1183]&m[1184]&m[1186]&~m[1187])|(~m[1122]&m[1183]&~m[1184]&~m[1186]&m[1187])|(~m[1122]&~m[1183]&m[1184]&~m[1186]&m[1187])|(m[1122]&m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1122]&m[1183]&m[1184]&m[1186]&m[1187]))&UnbiasedRNG[469])|((m[1122]&~m[1183]&~m[1184]&m[1186]&~m[1187])|(~m[1122]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1122]&~m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1122]&m[1183]&~m[1184]&~m[1186]&m[1187])|(m[1122]&~m[1183]&m[1184]&~m[1186]&m[1187])|(~m[1122]&~m[1183]&~m[1184]&m[1186]&m[1187])|(m[1122]&~m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1122]&m[1183]&~m[1184]&m[1186]&m[1187])|(m[1122]&m[1183]&~m[1184]&m[1186]&m[1187])|(~m[1122]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1122]&~m[1183]&m[1184]&m[1186]&m[1187])|(m[1122]&m[1183]&m[1184]&m[1186]&m[1187]));
    m[1190] = (((m[1127]&~m[1188]&~m[1189]&~m[1191]&~m[1192])|(~m[1127]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1127]&m[1188]&~m[1189]&m[1191]&~m[1192])|(m[1127]&~m[1188]&m[1189]&m[1191]&~m[1192])|(~m[1127]&m[1188]&~m[1189]&~m[1191]&m[1192])|(~m[1127]&~m[1188]&m[1189]&~m[1191]&m[1192])|(m[1127]&m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1127]&m[1188]&m[1189]&m[1191]&m[1192]))&UnbiasedRNG[470])|((m[1127]&~m[1188]&~m[1189]&m[1191]&~m[1192])|(~m[1127]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1127]&~m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1127]&m[1188]&~m[1189]&~m[1191]&m[1192])|(m[1127]&~m[1188]&m[1189]&~m[1191]&m[1192])|(~m[1127]&~m[1188]&~m[1189]&m[1191]&m[1192])|(m[1127]&~m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1127]&m[1188]&~m[1189]&m[1191]&m[1192])|(m[1127]&m[1188]&~m[1189]&m[1191]&m[1192])|(~m[1127]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1127]&~m[1188]&m[1189]&m[1191]&m[1192])|(m[1127]&m[1188]&m[1189]&m[1191]&m[1192]));
    m[1195] = (((m[1132]&~m[1193]&~m[1194]&~m[1196]&~m[1197])|(~m[1132]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1132]&m[1193]&~m[1194]&m[1196]&~m[1197])|(m[1132]&~m[1193]&m[1194]&m[1196]&~m[1197])|(~m[1132]&m[1193]&~m[1194]&~m[1196]&m[1197])|(~m[1132]&~m[1193]&m[1194]&~m[1196]&m[1197])|(m[1132]&m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1132]&m[1193]&m[1194]&m[1196]&m[1197]))&UnbiasedRNG[471])|((m[1132]&~m[1193]&~m[1194]&m[1196]&~m[1197])|(~m[1132]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1132]&~m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1132]&m[1193]&~m[1194]&~m[1196]&m[1197])|(m[1132]&~m[1193]&m[1194]&~m[1196]&m[1197])|(~m[1132]&~m[1193]&~m[1194]&m[1196]&m[1197])|(m[1132]&~m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1132]&m[1193]&~m[1194]&m[1196]&m[1197])|(m[1132]&m[1193]&~m[1194]&m[1196]&m[1197])|(~m[1132]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1132]&~m[1193]&m[1194]&m[1196]&m[1197])|(m[1132]&m[1193]&m[1194]&m[1196]&m[1197]));
    m[1200] = (((m[1137]&~m[1198]&~m[1199]&~m[1201]&~m[1202])|(~m[1137]&~m[1198]&~m[1199]&m[1201]&~m[1202])|(m[1137]&m[1198]&~m[1199]&m[1201]&~m[1202])|(m[1137]&~m[1198]&m[1199]&m[1201]&~m[1202])|(~m[1137]&m[1198]&~m[1199]&~m[1201]&m[1202])|(~m[1137]&~m[1198]&m[1199]&~m[1201]&m[1202])|(m[1137]&m[1198]&m[1199]&~m[1201]&m[1202])|(~m[1137]&m[1198]&m[1199]&m[1201]&m[1202]))&UnbiasedRNG[472])|((m[1137]&~m[1198]&~m[1199]&m[1201]&~m[1202])|(~m[1137]&~m[1198]&~m[1199]&~m[1201]&m[1202])|(m[1137]&~m[1198]&~m[1199]&~m[1201]&m[1202])|(m[1137]&m[1198]&~m[1199]&~m[1201]&m[1202])|(m[1137]&~m[1198]&m[1199]&~m[1201]&m[1202])|(~m[1137]&~m[1198]&~m[1199]&m[1201]&m[1202])|(m[1137]&~m[1198]&~m[1199]&m[1201]&m[1202])|(~m[1137]&m[1198]&~m[1199]&m[1201]&m[1202])|(m[1137]&m[1198]&~m[1199]&m[1201]&m[1202])|(~m[1137]&~m[1198]&m[1199]&m[1201]&m[1202])|(m[1137]&~m[1198]&m[1199]&m[1201]&m[1202])|(m[1137]&m[1198]&m[1199]&m[1201]&m[1202]));
    m[1205] = (((m[1142]&~m[1203]&~m[1204]&~m[1206]&~m[1207])|(~m[1142]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1142]&m[1203]&~m[1204]&m[1206]&~m[1207])|(m[1142]&~m[1203]&m[1204]&m[1206]&~m[1207])|(~m[1142]&m[1203]&~m[1204]&~m[1206]&m[1207])|(~m[1142]&~m[1203]&m[1204]&~m[1206]&m[1207])|(m[1142]&m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1142]&m[1203]&m[1204]&m[1206]&m[1207]))&UnbiasedRNG[473])|((m[1142]&~m[1203]&~m[1204]&m[1206]&~m[1207])|(~m[1142]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1142]&~m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1142]&m[1203]&~m[1204]&~m[1206]&m[1207])|(m[1142]&~m[1203]&m[1204]&~m[1206]&m[1207])|(~m[1142]&~m[1203]&~m[1204]&m[1206]&m[1207])|(m[1142]&~m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1142]&m[1203]&~m[1204]&m[1206]&m[1207])|(m[1142]&m[1203]&~m[1204]&m[1206]&m[1207])|(~m[1142]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1142]&~m[1203]&m[1204]&m[1206]&m[1207])|(m[1142]&m[1203]&m[1204]&m[1206]&m[1207]));
    m[1210] = (((m[1147]&~m[1208]&~m[1209]&~m[1211]&~m[1212])|(~m[1147]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1147]&m[1208]&~m[1209]&m[1211]&~m[1212])|(m[1147]&~m[1208]&m[1209]&m[1211]&~m[1212])|(~m[1147]&m[1208]&~m[1209]&~m[1211]&m[1212])|(~m[1147]&~m[1208]&m[1209]&~m[1211]&m[1212])|(m[1147]&m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1147]&m[1208]&m[1209]&m[1211]&m[1212]))&UnbiasedRNG[474])|((m[1147]&~m[1208]&~m[1209]&m[1211]&~m[1212])|(~m[1147]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1147]&~m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1147]&m[1208]&~m[1209]&~m[1211]&m[1212])|(m[1147]&~m[1208]&m[1209]&~m[1211]&m[1212])|(~m[1147]&~m[1208]&~m[1209]&m[1211]&m[1212])|(m[1147]&~m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1147]&m[1208]&~m[1209]&m[1211]&m[1212])|(m[1147]&m[1208]&~m[1209]&m[1211]&m[1212])|(~m[1147]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1147]&~m[1208]&m[1209]&m[1211]&m[1212])|(m[1147]&m[1208]&m[1209]&m[1211]&m[1212]));
    m[1215] = (((m[1152]&~m[1213]&~m[1214]&~m[1216]&~m[1217])|(~m[1152]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1152]&m[1213]&~m[1214]&m[1216]&~m[1217])|(m[1152]&~m[1213]&m[1214]&m[1216]&~m[1217])|(~m[1152]&m[1213]&~m[1214]&~m[1216]&m[1217])|(~m[1152]&~m[1213]&m[1214]&~m[1216]&m[1217])|(m[1152]&m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1152]&m[1213]&m[1214]&m[1216]&m[1217]))&UnbiasedRNG[475])|((m[1152]&~m[1213]&~m[1214]&m[1216]&~m[1217])|(~m[1152]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1152]&~m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1152]&m[1213]&~m[1214]&~m[1216]&m[1217])|(m[1152]&~m[1213]&m[1214]&~m[1216]&m[1217])|(~m[1152]&~m[1213]&~m[1214]&m[1216]&m[1217])|(m[1152]&~m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1152]&m[1213]&~m[1214]&m[1216]&m[1217])|(m[1152]&m[1213]&~m[1214]&m[1216]&m[1217])|(~m[1152]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1152]&~m[1213]&m[1214]&m[1216]&m[1217])|(m[1152]&m[1213]&m[1214]&m[1216]&m[1217]));
    m[1220] = (((m[1157]&~m[1218]&~m[1219]&~m[1221]&~m[1222])|(~m[1157]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1157]&m[1218]&~m[1219]&m[1221]&~m[1222])|(m[1157]&~m[1218]&m[1219]&m[1221]&~m[1222])|(~m[1157]&m[1218]&~m[1219]&~m[1221]&m[1222])|(~m[1157]&~m[1218]&m[1219]&~m[1221]&m[1222])|(m[1157]&m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1157]&m[1218]&m[1219]&m[1221]&m[1222]))&UnbiasedRNG[476])|((m[1157]&~m[1218]&~m[1219]&m[1221]&~m[1222])|(~m[1157]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1157]&~m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1157]&m[1218]&~m[1219]&~m[1221]&m[1222])|(m[1157]&~m[1218]&m[1219]&~m[1221]&m[1222])|(~m[1157]&~m[1218]&~m[1219]&m[1221]&m[1222])|(m[1157]&~m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1157]&m[1218]&~m[1219]&m[1221]&m[1222])|(m[1157]&m[1218]&~m[1219]&m[1221]&m[1222])|(~m[1157]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1157]&~m[1218]&m[1219]&m[1221]&m[1222])|(m[1157]&m[1218]&m[1219]&m[1221]&m[1222]));
    m[1225] = (((m[1162]&~m[1223]&~m[1224]&~m[1226]&~m[1227])|(~m[1162]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1162]&m[1223]&~m[1224]&m[1226]&~m[1227])|(m[1162]&~m[1223]&m[1224]&m[1226]&~m[1227])|(~m[1162]&m[1223]&~m[1224]&~m[1226]&m[1227])|(~m[1162]&~m[1223]&m[1224]&~m[1226]&m[1227])|(m[1162]&m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1162]&m[1223]&m[1224]&m[1226]&m[1227]))&UnbiasedRNG[477])|((m[1162]&~m[1223]&~m[1224]&m[1226]&~m[1227])|(~m[1162]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1162]&~m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1162]&m[1223]&~m[1224]&~m[1226]&m[1227])|(m[1162]&~m[1223]&m[1224]&~m[1226]&m[1227])|(~m[1162]&~m[1223]&~m[1224]&m[1226]&m[1227])|(m[1162]&~m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1162]&m[1223]&~m[1224]&m[1226]&m[1227])|(m[1162]&m[1223]&~m[1224]&m[1226]&m[1227])|(~m[1162]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1162]&~m[1223]&m[1224]&m[1226]&m[1227])|(m[1162]&m[1223]&m[1224]&m[1226]&m[1227]));
    m[1230] = (((m[1167]&~m[1228]&~m[1229]&~m[1231]&~m[1232])|(~m[1167]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1167]&m[1228]&~m[1229]&m[1231]&~m[1232])|(m[1167]&~m[1228]&m[1229]&m[1231]&~m[1232])|(~m[1167]&m[1228]&~m[1229]&~m[1231]&m[1232])|(~m[1167]&~m[1228]&m[1229]&~m[1231]&m[1232])|(m[1167]&m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1167]&m[1228]&m[1229]&m[1231]&m[1232]))&UnbiasedRNG[478])|((m[1167]&~m[1228]&~m[1229]&m[1231]&~m[1232])|(~m[1167]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1167]&~m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1167]&m[1228]&~m[1229]&~m[1231]&m[1232])|(m[1167]&~m[1228]&m[1229]&~m[1231]&m[1232])|(~m[1167]&~m[1228]&~m[1229]&m[1231]&m[1232])|(m[1167]&~m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1167]&m[1228]&~m[1229]&m[1231]&m[1232])|(m[1167]&m[1228]&~m[1229]&m[1231]&m[1232])|(~m[1167]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1167]&~m[1228]&m[1229]&m[1231]&m[1232])|(m[1167]&m[1228]&m[1229]&m[1231]&m[1232]));
    m[1235] = (((m[1172]&~m[1233]&~m[1234]&~m[1236]&~m[1237])|(~m[1172]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1172]&m[1233]&~m[1234]&m[1236]&~m[1237])|(m[1172]&~m[1233]&m[1234]&m[1236]&~m[1237])|(~m[1172]&m[1233]&~m[1234]&~m[1236]&m[1237])|(~m[1172]&~m[1233]&m[1234]&~m[1236]&m[1237])|(m[1172]&m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1172]&m[1233]&m[1234]&m[1236]&m[1237]))&UnbiasedRNG[479])|((m[1172]&~m[1233]&~m[1234]&m[1236]&~m[1237])|(~m[1172]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1172]&~m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1172]&m[1233]&~m[1234]&~m[1236]&m[1237])|(m[1172]&~m[1233]&m[1234]&~m[1236]&m[1237])|(~m[1172]&~m[1233]&~m[1234]&m[1236]&m[1237])|(m[1172]&~m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1172]&m[1233]&~m[1234]&m[1236]&m[1237])|(m[1172]&m[1233]&~m[1234]&m[1236]&m[1237])|(~m[1172]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1172]&~m[1233]&m[1234]&m[1236]&m[1237])|(m[1172]&m[1233]&m[1234]&m[1236]&m[1237]));
    m[1240] = (((m[1177]&~m[1238]&~m[1239]&~m[1241]&~m[1242])|(~m[1177]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1177]&m[1238]&~m[1239]&m[1241]&~m[1242])|(m[1177]&~m[1238]&m[1239]&m[1241]&~m[1242])|(~m[1177]&m[1238]&~m[1239]&~m[1241]&m[1242])|(~m[1177]&~m[1238]&m[1239]&~m[1241]&m[1242])|(m[1177]&m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1177]&m[1238]&m[1239]&m[1241]&m[1242]))&UnbiasedRNG[480])|((m[1177]&~m[1238]&~m[1239]&m[1241]&~m[1242])|(~m[1177]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1177]&~m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1177]&m[1238]&~m[1239]&~m[1241]&m[1242])|(m[1177]&~m[1238]&m[1239]&~m[1241]&m[1242])|(~m[1177]&~m[1238]&~m[1239]&m[1241]&m[1242])|(m[1177]&~m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1177]&m[1238]&~m[1239]&m[1241]&m[1242])|(m[1177]&m[1238]&~m[1239]&m[1241]&m[1242])|(~m[1177]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1177]&~m[1238]&m[1239]&m[1241]&m[1242])|(m[1177]&m[1238]&m[1239]&m[1241]&m[1242]));
    m[1245] = (((m[1182]&~m[1243]&~m[1244]&~m[1246]&~m[1247])|(~m[1182]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1182]&m[1243]&~m[1244]&m[1246]&~m[1247])|(m[1182]&~m[1243]&m[1244]&m[1246]&~m[1247])|(~m[1182]&m[1243]&~m[1244]&~m[1246]&m[1247])|(~m[1182]&~m[1243]&m[1244]&~m[1246]&m[1247])|(m[1182]&m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1182]&m[1243]&m[1244]&m[1246]&m[1247]))&UnbiasedRNG[481])|((m[1182]&~m[1243]&~m[1244]&m[1246]&~m[1247])|(~m[1182]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1182]&~m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1182]&m[1243]&~m[1244]&~m[1246]&m[1247])|(m[1182]&~m[1243]&m[1244]&~m[1246]&m[1247])|(~m[1182]&~m[1243]&~m[1244]&m[1246]&m[1247])|(m[1182]&~m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1182]&m[1243]&~m[1244]&m[1246]&m[1247])|(m[1182]&m[1243]&~m[1244]&m[1246]&m[1247])|(~m[1182]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1182]&~m[1243]&m[1244]&m[1246]&m[1247])|(m[1182]&m[1243]&m[1244]&m[1246]&m[1247]));
    m[1250] = (((m[1192]&~m[1248]&~m[1249]&~m[1251]&~m[1252])|(~m[1192]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1192]&m[1248]&~m[1249]&m[1251]&~m[1252])|(m[1192]&~m[1248]&m[1249]&m[1251]&~m[1252])|(~m[1192]&m[1248]&~m[1249]&~m[1251]&m[1252])|(~m[1192]&~m[1248]&m[1249]&~m[1251]&m[1252])|(m[1192]&m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1192]&m[1248]&m[1249]&m[1251]&m[1252]))&UnbiasedRNG[482])|((m[1192]&~m[1248]&~m[1249]&m[1251]&~m[1252])|(~m[1192]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1192]&~m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1192]&m[1248]&~m[1249]&~m[1251]&m[1252])|(m[1192]&~m[1248]&m[1249]&~m[1251]&m[1252])|(~m[1192]&~m[1248]&~m[1249]&m[1251]&m[1252])|(m[1192]&~m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1192]&m[1248]&~m[1249]&m[1251]&m[1252])|(m[1192]&m[1248]&~m[1249]&m[1251]&m[1252])|(~m[1192]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1192]&~m[1248]&m[1249]&m[1251]&m[1252])|(m[1192]&m[1248]&m[1249]&m[1251]&m[1252]));
    m[1255] = (((m[1197]&~m[1253]&~m[1254]&~m[1256]&~m[1257])|(~m[1197]&~m[1253]&~m[1254]&m[1256]&~m[1257])|(m[1197]&m[1253]&~m[1254]&m[1256]&~m[1257])|(m[1197]&~m[1253]&m[1254]&m[1256]&~m[1257])|(~m[1197]&m[1253]&~m[1254]&~m[1256]&m[1257])|(~m[1197]&~m[1253]&m[1254]&~m[1256]&m[1257])|(m[1197]&m[1253]&m[1254]&~m[1256]&m[1257])|(~m[1197]&m[1253]&m[1254]&m[1256]&m[1257]))&UnbiasedRNG[483])|((m[1197]&~m[1253]&~m[1254]&m[1256]&~m[1257])|(~m[1197]&~m[1253]&~m[1254]&~m[1256]&m[1257])|(m[1197]&~m[1253]&~m[1254]&~m[1256]&m[1257])|(m[1197]&m[1253]&~m[1254]&~m[1256]&m[1257])|(m[1197]&~m[1253]&m[1254]&~m[1256]&m[1257])|(~m[1197]&~m[1253]&~m[1254]&m[1256]&m[1257])|(m[1197]&~m[1253]&~m[1254]&m[1256]&m[1257])|(~m[1197]&m[1253]&~m[1254]&m[1256]&m[1257])|(m[1197]&m[1253]&~m[1254]&m[1256]&m[1257])|(~m[1197]&~m[1253]&m[1254]&m[1256]&m[1257])|(m[1197]&~m[1253]&m[1254]&m[1256]&m[1257])|(m[1197]&m[1253]&m[1254]&m[1256]&m[1257]));
    m[1260] = (((m[1202]&~m[1258]&~m[1259]&~m[1261]&~m[1262])|(~m[1202]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1202]&m[1258]&~m[1259]&m[1261]&~m[1262])|(m[1202]&~m[1258]&m[1259]&m[1261]&~m[1262])|(~m[1202]&m[1258]&~m[1259]&~m[1261]&m[1262])|(~m[1202]&~m[1258]&m[1259]&~m[1261]&m[1262])|(m[1202]&m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1202]&m[1258]&m[1259]&m[1261]&m[1262]))&UnbiasedRNG[484])|((m[1202]&~m[1258]&~m[1259]&m[1261]&~m[1262])|(~m[1202]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1202]&~m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1202]&m[1258]&~m[1259]&~m[1261]&m[1262])|(m[1202]&~m[1258]&m[1259]&~m[1261]&m[1262])|(~m[1202]&~m[1258]&~m[1259]&m[1261]&m[1262])|(m[1202]&~m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1202]&m[1258]&~m[1259]&m[1261]&m[1262])|(m[1202]&m[1258]&~m[1259]&m[1261]&m[1262])|(~m[1202]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1202]&~m[1258]&m[1259]&m[1261]&m[1262])|(m[1202]&m[1258]&m[1259]&m[1261]&m[1262]));
    m[1265] = (((m[1207]&~m[1263]&~m[1264]&~m[1266]&~m[1267])|(~m[1207]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1207]&m[1263]&~m[1264]&m[1266]&~m[1267])|(m[1207]&~m[1263]&m[1264]&m[1266]&~m[1267])|(~m[1207]&m[1263]&~m[1264]&~m[1266]&m[1267])|(~m[1207]&~m[1263]&m[1264]&~m[1266]&m[1267])|(m[1207]&m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1207]&m[1263]&m[1264]&m[1266]&m[1267]))&UnbiasedRNG[485])|((m[1207]&~m[1263]&~m[1264]&m[1266]&~m[1267])|(~m[1207]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1207]&~m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1207]&m[1263]&~m[1264]&~m[1266]&m[1267])|(m[1207]&~m[1263]&m[1264]&~m[1266]&m[1267])|(~m[1207]&~m[1263]&~m[1264]&m[1266]&m[1267])|(m[1207]&~m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1207]&m[1263]&~m[1264]&m[1266]&m[1267])|(m[1207]&m[1263]&~m[1264]&m[1266]&m[1267])|(~m[1207]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1207]&~m[1263]&m[1264]&m[1266]&m[1267])|(m[1207]&m[1263]&m[1264]&m[1266]&m[1267]));
    m[1270] = (((m[1212]&~m[1268]&~m[1269]&~m[1271]&~m[1272])|(~m[1212]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1212]&m[1268]&~m[1269]&m[1271]&~m[1272])|(m[1212]&~m[1268]&m[1269]&m[1271]&~m[1272])|(~m[1212]&m[1268]&~m[1269]&~m[1271]&m[1272])|(~m[1212]&~m[1268]&m[1269]&~m[1271]&m[1272])|(m[1212]&m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1212]&m[1268]&m[1269]&m[1271]&m[1272]))&UnbiasedRNG[486])|((m[1212]&~m[1268]&~m[1269]&m[1271]&~m[1272])|(~m[1212]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1212]&~m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1212]&m[1268]&~m[1269]&~m[1271]&m[1272])|(m[1212]&~m[1268]&m[1269]&~m[1271]&m[1272])|(~m[1212]&~m[1268]&~m[1269]&m[1271]&m[1272])|(m[1212]&~m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1212]&m[1268]&~m[1269]&m[1271]&m[1272])|(m[1212]&m[1268]&~m[1269]&m[1271]&m[1272])|(~m[1212]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1212]&~m[1268]&m[1269]&m[1271]&m[1272])|(m[1212]&m[1268]&m[1269]&m[1271]&m[1272]));
    m[1275] = (((m[1217]&~m[1273]&~m[1274]&~m[1276]&~m[1277])|(~m[1217]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1217]&m[1273]&~m[1274]&m[1276]&~m[1277])|(m[1217]&~m[1273]&m[1274]&m[1276]&~m[1277])|(~m[1217]&m[1273]&~m[1274]&~m[1276]&m[1277])|(~m[1217]&~m[1273]&m[1274]&~m[1276]&m[1277])|(m[1217]&m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1217]&m[1273]&m[1274]&m[1276]&m[1277]))&UnbiasedRNG[487])|((m[1217]&~m[1273]&~m[1274]&m[1276]&~m[1277])|(~m[1217]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1217]&~m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1217]&m[1273]&~m[1274]&~m[1276]&m[1277])|(m[1217]&~m[1273]&m[1274]&~m[1276]&m[1277])|(~m[1217]&~m[1273]&~m[1274]&m[1276]&m[1277])|(m[1217]&~m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1217]&m[1273]&~m[1274]&m[1276]&m[1277])|(m[1217]&m[1273]&~m[1274]&m[1276]&m[1277])|(~m[1217]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1217]&~m[1273]&m[1274]&m[1276]&m[1277])|(m[1217]&m[1273]&m[1274]&m[1276]&m[1277]));
    m[1280] = (((m[1222]&~m[1278]&~m[1279]&~m[1281]&~m[1282])|(~m[1222]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1222]&m[1278]&~m[1279]&m[1281]&~m[1282])|(m[1222]&~m[1278]&m[1279]&m[1281]&~m[1282])|(~m[1222]&m[1278]&~m[1279]&~m[1281]&m[1282])|(~m[1222]&~m[1278]&m[1279]&~m[1281]&m[1282])|(m[1222]&m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1222]&m[1278]&m[1279]&m[1281]&m[1282]))&UnbiasedRNG[488])|((m[1222]&~m[1278]&~m[1279]&m[1281]&~m[1282])|(~m[1222]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1222]&~m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1222]&m[1278]&~m[1279]&~m[1281]&m[1282])|(m[1222]&~m[1278]&m[1279]&~m[1281]&m[1282])|(~m[1222]&~m[1278]&~m[1279]&m[1281]&m[1282])|(m[1222]&~m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1222]&m[1278]&~m[1279]&m[1281]&m[1282])|(m[1222]&m[1278]&~m[1279]&m[1281]&m[1282])|(~m[1222]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1222]&~m[1278]&m[1279]&m[1281]&m[1282])|(m[1222]&m[1278]&m[1279]&m[1281]&m[1282]));
    m[1285] = (((m[1227]&~m[1283]&~m[1284]&~m[1286]&~m[1287])|(~m[1227]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1227]&m[1283]&~m[1284]&m[1286]&~m[1287])|(m[1227]&~m[1283]&m[1284]&m[1286]&~m[1287])|(~m[1227]&m[1283]&~m[1284]&~m[1286]&m[1287])|(~m[1227]&~m[1283]&m[1284]&~m[1286]&m[1287])|(m[1227]&m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1227]&m[1283]&m[1284]&m[1286]&m[1287]))&UnbiasedRNG[489])|((m[1227]&~m[1283]&~m[1284]&m[1286]&~m[1287])|(~m[1227]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1227]&~m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1227]&m[1283]&~m[1284]&~m[1286]&m[1287])|(m[1227]&~m[1283]&m[1284]&~m[1286]&m[1287])|(~m[1227]&~m[1283]&~m[1284]&m[1286]&m[1287])|(m[1227]&~m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1227]&m[1283]&~m[1284]&m[1286]&m[1287])|(m[1227]&m[1283]&~m[1284]&m[1286]&m[1287])|(~m[1227]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1227]&~m[1283]&m[1284]&m[1286]&m[1287])|(m[1227]&m[1283]&m[1284]&m[1286]&m[1287]));
    m[1290] = (((m[1232]&~m[1288]&~m[1289]&~m[1291]&~m[1292])|(~m[1232]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1232]&m[1288]&~m[1289]&m[1291]&~m[1292])|(m[1232]&~m[1288]&m[1289]&m[1291]&~m[1292])|(~m[1232]&m[1288]&~m[1289]&~m[1291]&m[1292])|(~m[1232]&~m[1288]&m[1289]&~m[1291]&m[1292])|(m[1232]&m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1232]&m[1288]&m[1289]&m[1291]&m[1292]))&UnbiasedRNG[490])|((m[1232]&~m[1288]&~m[1289]&m[1291]&~m[1292])|(~m[1232]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1232]&~m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1232]&m[1288]&~m[1289]&~m[1291]&m[1292])|(m[1232]&~m[1288]&m[1289]&~m[1291]&m[1292])|(~m[1232]&~m[1288]&~m[1289]&m[1291]&m[1292])|(m[1232]&~m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1232]&m[1288]&~m[1289]&m[1291]&m[1292])|(m[1232]&m[1288]&~m[1289]&m[1291]&m[1292])|(~m[1232]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1232]&~m[1288]&m[1289]&m[1291]&m[1292])|(m[1232]&m[1288]&m[1289]&m[1291]&m[1292]));
    m[1295] = (((m[1237]&~m[1293]&~m[1294]&~m[1296]&~m[1297])|(~m[1237]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1237]&m[1293]&~m[1294]&m[1296]&~m[1297])|(m[1237]&~m[1293]&m[1294]&m[1296]&~m[1297])|(~m[1237]&m[1293]&~m[1294]&~m[1296]&m[1297])|(~m[1237]&~m[1293]&m[1294]&~m[1296]&m[1297])|(m[1237]&m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1237]&m[1293]&m[1294]&m[1296]&m[1297]))&UnbiasedRNG[491])|((m[1237]&~m[1293]&~m[1294]&m[1296]&~m[1297])|(~m[1237]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1237]&~m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1237]&m[1293]&~m[1294]&~m[1296]&m[1297])|(m[1237]&~m[1293]&m[1294]&~m[1296]&m[1297])|(~m[1237]&~m[1293]&~m[1294]&m[1296]&m[1297])|(m[1237]&~m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1237]&m[1293]&~m[1294]&m[1296]&m[1297])|(m[1237]&m[1293]&~m[1294]&m[1296]&m[1297])|(~m[1237]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1237]&~m[1293]&m[1294]&m[1296]&m[1297])|(m[1237]&m[1293]&m[1294]&m[1296]&m[1297]));
    m[1300] = (((m[1242]&~m[1298]&~m[1299]&~m[1301]&~m[1302])|(~m[1242]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1242]&m[1298]&~m[1299]&m[1301]&~m[1302])|(m[1242]&~m[1298]&m[1299]&m[1301]&~m[1302])|(~m[1242]&m[1298]&~m[1299]&~m[1301]&m[1302])|(~m[1242]&~m[1298]&m[1299]&~m[1301]&m[1302])|(m[1242]&m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1242]&m[1298]&m[1299]&m[1301]&m[1302]))&UnbiasedRNG[492])|((m[1242]&~m[1298]&~m[1299]&m[1301]&~m[1302])|(~m[1242]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1242]&~m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1242]&m[1298]&~m[1299]&~m[1301]&m[1302])|(m[1242]&~m[1298]&m[1299]&~m[1301]&m[1302])|(~m[1242]&~m[1298]&~m[1299]&m[1301]&m[1302])|(m[1242]&~m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1242]&m[1298]&~m[1299]&m[1301]&m[1302])|(m[1242]&m[1298]&~m[1299]&m[1301]&m[1302])|(~m[1242]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1242]&~m[1298]&m[1299]&m[1301]&m[1302])|(m[1242]&m[1298]&m[1299]&m[1301]&m[1302]));
    m[1305] = (((m[1247]&~m[1303]&~m[1304]&~m[1306]&~m[1307])|(~m[1247]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1247]&m[1303]&~m[1304]&m[1306]&~m[1307])|(m[1247]&~m[1303]&m[1304]&m[1306]&~m[1307])|(~m[1247]&m[1303]&~m[1304]&~m[1306]&m[1307])|(~m[1247]&~m[1303]&m[1304]&~m[1306]&m[1307])|(m[1247]&m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1247]&m[1303]&m[1304]&m[1306]&m[1307]))&UnbiasedRNG[493])|((m[1247]&~m[1303]&~m[1304]&m[1306]&~m[1307])|(~m[1247]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1247]&~m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1247]&m[1303]&~m[1304]&~m[1306]&m[1307])|(m[1247]&~m[1303]&m[1304]&~m[1306]&m[1307])|(~m[1247]&~m[1303]&~m[1304]&m[1306]&m[1307])|(m[1247]&~m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1247]&m[1303]&~m[1304]&m[1306]&m[1307])|(m[1247]&m[1303]&~m[1304]&m[1306]&m[1307])|(~m[1247]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1247]&~m[1303]&m[1304]&m[1306]&m[1307])|(m[1247]&m[1303]&m[1304]&m[1306]&m[1307]));
    m[1310] = (((m[1257]&~m[1308]&~m[1309]&~m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&~m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&~m[1312])|(~m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&m[1308]&m[1309]&m[1311]&m[1312]))&UnbiasedRNG[494])|((m[1257]&~m[1308]&~m[1309]&m[1311]&~m[1312])|(~m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&~m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&~m[1311]&m[1312])|(~m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&~m[1309]&m[1311]&m[1312])|(~m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&~m[1308]&m[1309]&m[1311]&m[1312])|(m[1257]&m[1308]&m[1309]&m[1311]&m[1312]));
    m[1315] = (((m[1262]&~m[1313]&~m[1314]&~m[1316]&~m[1317])|(~m[1262]&~m[1313]&~m[1314]&m[1316]&~m[1317])|(m[1262]&m[1313]&~m[1314]&m[1316]&~m[1317])|(m[1262]&~m[1313]&m[1314]&m[1316]&~m[1317])|(~m[1262]&m[1313]&~m[1314]&~m[1316]&m[1317])|(~m[1262]&~m[1313]&m[1314]&~m[1316]&m[1317])|(m[1262]&m[1313]&m[1314]&~m[1316]&m[1317])|(~m[1262]&m[1313]&m[1314]&m[1316]&m[1317]))&UnbiasedRNG[495])|((m[1262]&~m[1313]&~m[1314]&m[1316]&~m[1317])|(~m[1262]&~m[1313]&~m[1314]&~m[1316]&m[1317])|(m[1262]&~m[1313]&~m[1314]&~m[1316]&m[1317])|(m[1262]&m[1313]&~m[1314]&~m[1316]&m[1317])|(m[1262]&~m[1313]&m[1314]&~m[1316]&m[1317])|(~m[1262]&~m[1313]&~m[1314]&m[1316]&m[1317])|(m[1262]&~m[1313]&~m[1314]&m[1316]&m[1317])|(~m[1262]&m[1313]&~m[1314]&m[1316]&m[1317])|(m[1262]&m[1313]&~m[1314]&m[1316]&m[1317])|(~m[1262]&~m[1313]&m[1314]&m[1316]&m[1317])|(m[1262]&~m[1313]&m[1314]&m[1316]&m[1317])|(m[1262]&m[1313]&m[1314]&m[1316]&m[1317]));
    m[1320] = (((m[1267]&~m[1318]&~m[1319]&~m[1321]&~m[1322])|(~m[1267]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1267]&m[1318]&~m[1319]&m[1321]&~m[1322])|(m[1267]&~m[1318]&m[1319]&m[1321]&~m[1322])|(~m[1267]&m[1318]&~m[1319]&~m[1321]&m[1322])|(~m[1267]&~m[1318]&m[1319]&~m[1321]&m[1322])|(m[1267]&m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1267]&m[1318]&m[1319]&m[1321]&m[1322]))&UnbiasedRNG[496])|((m[1267]&~m[1318]&~m[1319]&m[1321]&~m[1322])|(~m[1267]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1267]&~m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1267]&m[1318]&~m[1319]&~m[1321]&m[1322])|(m[1267]&~m[1318]&m[1319]&~m[1321]&m[1322])|(~m[1267]&~m[1318]&~m[1319]&m[1321]&m[1322])|(m[1267]&~m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1267]&m[1318]&~m[1319]&m[1321]&m[1322])|(m[1267]&m[1318]&~m[1319]&m[1321]&m[1322])|(~m[1267]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1267]&~m[1318]&m[1319]&m[1321]&m[1322])|(m[1267]&m[1318]&m[1319]&m[1321]&m[1322]));
    m[1325] = (((m[1272]&~m[1323]&~m[1324]&~m[1326]&~m[1327])|(~m[1272]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1272]&m[1323]&~m[1324]&m[1326]&~m[1327])|(m[1272]&~m[1323]&m[1324]&m[1326]&~m[1327])|(~m[1272]&m[1323]&~m[1324]&~m[1326]&m[1327])|(~m[1272]&~m[1323]&m[1324]&~m[1326]&m[1327])|(m[1272]&m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1272]&m[1323]&m[1324]&m[1326]&m[1327]))&UnbiasedRNG[497])|((m[1272]&~m[1323]&~m[1324]&m[1326]&~m[1327])|(~m[1272]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1272]&~m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1272]&m[1323]&~m[1324]&~m[1326]&m[1327])|(m[1272]&~m[1323]&m[1324]&~m[1326]&m[1327])|(~m[1272]&~m[1323]&~m[1324]&m[1326]&m[1327])|(m[1272]&~m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1272]&m[1323]&~m[1324]&m[1326]&m[1327])|(m[1272]&m[1323]&~m[1324]&m[1326]&m[1327])|(~m[1272]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1272]&~m[1323]&m[1324]&m[1326]&m[1327])|(m[1272]&m[1323]&m[1324]&m[1326]&m[1327]));
    m[1330] = (((m[1277]&~m[1328]&~m[1329]&~m[1331]&~m[1332])|(~m[1277]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1277]&m[1328]&~m[1329]&m[1331]&~m[1332])|(m[1277]&~m[1328]&m[1329]&m[1331]&~m[1332])|(~m[1277]&m[1328]&~m[1329]&~m[1331]&m[1332])|(~m[1277]&~m[1328]&m[1329]&~m[1331]&m[1332])|(m[1277]&m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1277]&m[1328]&m[1329]&m[1331]&m[1332]))&UnbiasedRNG[498])|((m[1277]&~m[1328]&~m[1329]&m[1331]&~m[1332])|(~m[1277]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1277]&~m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1277]&m[1328]&~m[1329]&~m[1331]&m[1332])|(m[1277]&~m[1328]&m[1329]&~m[1331]&m[1332])|(~m[1277]&~m[1328]&~m[1329]&m[1331]&m[1332])|(m[1277]&~m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1277]&m[1328]&~m[1329]&m[1331]&m[1332])|(m[1277]&m[1328]&~m[1329]&m[1331]&m[1332])|(~m[1277]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1277]&~m[1328]&m[1329]&m[1331]&m[1332])|(m[1277]&m[1328]&m[1329]&m[1331]&m[1332]));
    m[1335] = (((m[1282]&~m[1333]&~m[1334]&~m[1336]&~m[1337])|(~m[1282]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1282]&m[1333]&~m[1334]&m[1336]&~m[1337])|(m[1282]&~m[1333]&m[1334]&m[1336]&~m[1337])|(~m[1282]&m[1333]&~m[1334]&~m[1336]&m[1337])|(~m[1282]&~m[1333]&m[1334]&~m[1336]&m[1337])|(m[1282]&m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1282]&m[1333]&m[1334]&m[1336]&m[1337]))&UnbiasedRNG[499])|((m[1282]&~m[1333]&~m[1334]&m[1336]&~m[1337])|(~m[1282]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1282]&~m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1282]&m[1333]&~m[1334]&~m[1336]&m[1337])|(m[1282]&~m[1333]&m[1334]&~m[1336]&m[1337])|(~m[1282]&~m[1333]&~m[1334]&m[1336]&m[1337])|(m[1282]&~m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1282]&m[1333]&~m[1334]&m[1336]&m[1337])|(m[1282]&m[1333]&~m[1334]&m[1336]&m[1337])|(~m[1282]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1282]&~m[1333]&m[1334]&m[1336]&m[1337])|(m[1282]&m[1333]&m[1334]&m[1336]&m[1337]));
    m[1340] = (((m[1287]&~m[1338]&~m[1339]&~m[1341]&~m[1342])|(~m[1287]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1287]&m[1338]&~m[1339]&m[1341]&~m[1342])|(m[1287]&~m[1338]&m[1339]&m[1341]&~m[1342])|(~m[1287]&m[1338]&~m[1339]&~m[1341]&m[1342])|(~m[1287]&~m[1338]&m[1339]&~m[1341]&m[1342])|(m[1287]&m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1287]&m[1338]&m[1339]&m[1341]&m[1342]))&UnbiasedRNG[500])|((m[1287]&~m[1338]&~m[1339]&m[1341]&~m[1342])|(~m[1287]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1287]&~m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1287]&m[1338]&~m[1339]&~m[1341]&m[1342])|(m[1287]&~m[1338]&m[1339]&~m[1341]&m[1342])|(~m[1287]&~m[1338]&~m[1339]&m[1341]&m[1342])|(m[1287]&~m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1287]&m[1338]&~m[1339]&m[1341]&m[1342])|(m[1287]&m[1338]&~m[1339]&m[1341]&m[1342])|(~m[1287]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1287]&~m[1338]&m[1339]&m[1341]&m[1342])|(m[1287]&m[1338]&m[1339]&m[1341]&m[1342]));
    m[1345] = (((m[1292]&~m[1343]&~m[1344]&~m[1346]&~m[1347])|(~m[1292]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1292]&m[1343]&~m[1344]&m[1346]&~m[1347])|(m[1292]&~m[1343]&m[1344]&m[1346]&~m[1347])|(~m[1292]&m[1343]&~m[1344]&~m[1346]&m[1347])|(~m[1292]&~m[1343]&m[1344]&~m[1346]&m[1347])|(m[1292]&m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1292]&m[1343]&m[1344]&m[1346]&m[1347]))&UnbiasedRNG[501])|((m[1292]&~m[1343]&~m[1344]&m[1346]&~m[1347])|(~m[1292]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1292]&~m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1292]&m[1343]&~m[1344]&~m[1346]&m[1347])|(m[1292]&~m[1343]&m[1344]&~m[1346]&m[1347])|(~m[1292]&~m[1343]&~m[1344]&m[1346]&m[1347])|(m[1292]&~m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1292]&m[1343]&~m[1344]&m[1346]&m[1347])|(m[1292]&m[1343]&~m[1344]&m[1346]&m[1347])|(~m[1292]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1292]&~m[1343]&m[1344]&m[1346]&m[1347])|(m[1292]&m[1343]&m[1344]&m[1346]&m[1347]));
    m[1350] = (((m[1297]&~m[1348]&~m[1349]&~m[1351]&~m[1352])|(~m[1297]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1297]&m[1348]&~m[1349]&m[1351]&~m[1352])|(m[1297]&~m[1348]&m[1349]&m[1351]&~m[1352])|(~m[1297]&m[1348]&~m[1349]&~m[1351]&m[1352])|(~m[1297]&~m[1348]&m[1349]&~m[1351]&m[1352])|(m[1297]&m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1297]&m[1348]&m[1349]&m[1351]&m[1352]))&UnbiasedRNG[502])|((m[1297]&~m[1348]&~m[1349]&m[1351]&~m[1352])|(~m[1297]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1297]&~m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1297]&m[1348]&~m[1349]&~m[1351]&m[1352])|(m[1297]&~m[1348]&m[1349]&~m[1351]&m[1352])|(~m[1297]&~m[1348]&~m[1349]&m[1351]&m[1352])|(m[1297]&~m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1297]&m[1348]&~m[1349]&m[1351]&m[1352])|(m[1297]&m[1348]&~m[1349]&m[1351]&m[1352])|(~m[1297]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1297]&~m[1348]&m[1349]&m[1351]&m[1352])|(m[1297]&m[1348]&m[1349]&m[1351]&m[1352]));
    m[1355] = (((m[1302]&~m[1353]&~m[1354]&~m[1356]&~m[1357])|(~m[1302]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1302]&m[1353]&~m[1354]&m[1356]&~m[1357])|(m[1302]&~m[1353]&m[1354]&m[1356]&~m[1357])|(~m[1302]&m[1353]&~m[1354]&~m[1356]&m[1357])|(~m[1302]&~m[1353]&m[1354]&~m[1356]&m[1357])|(m[1302]&m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1302]&m[1353]&m[1354]&m[1356]&m[1357]))&UnbiasedRNG[503])|((m[1302]&~m[1353]&~m[1354]&m[1356]&~m[1357])|(~m[1302]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1302]&~m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1302]&m[1353]&~m[1354]&~m[1356]&m[1357])|(m[1302]&~m[1353]&m[1354]&~m[1356]&m[1357])|(~m[1302]&~m[1353]&~m[1354]&m[1356]&m[1357])|(m[1302]&~m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1302]&m[1353]&~m[1354]&m[1356]&m[1357])|(m[1302]&m[1353]&~m[1354]&m[1356]&m[1357])|(~m[1302]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1302]&~m[1353]&m[1354]&m[1356]&m[1357])|(m[1302]&m[1353]&m[1354]&m[1356]&m[1357]));
    m[1360] = (((m[1307]&~m[1358]&~m[1359]&~m[1361]&~m[1362])|(~m[1307]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1307]&m[1358]&~m[1359]&m[1361]&~m[1362])|(m[1307]&~m[1358]&m[1359]&m[1361]&~m[1362])|(~m[1307]&m[1358]&~m[1359]&~m[1361]&m[1362])|(~m[1307]&~m[1358]&m[1359]&~m[1361]&m[1362])|(m[1307]&m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1307]&m[1358]&m[1359]&m[1361]&m[1362]))&UnbiasedRNG[504])|((m[1307]&~m[1358]&~m[1359]&m[1361]&~m[1362])|(~m[1307]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1307]&~m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1307]&m[1358]&~m[1359]&~m[1361]&m[1362])|(m[1307]&~m[1358]&m[1359]&~m[1361]&m[1362])|(~m[1307]&~m[1358]&~m[1359]&m[1361]&m[1362])|(m[1307]&~m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1307]&m[1358]&~m[1359]&m[1361]&m[1362])|(m[1307]&m[1358]&~m[1359]&m[1361]&m[1362])|(~m[1307]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1307]&~m[1358]&m[1359]&m[1361]&m[1362])|(m[1307]&m[1358]&m[1359]&m[1361]&m[1362]));
    m[1365] = (((m[1317]&~m[1363]&~m[1364]&~m[1366]&~m[1367])|(~m[1317]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1317]&m[1363]&~m[1364]&m[1366]&~m[1367])|(m[1317]&~m[1363]&m[1364]&m[1366]&~m[1367])|(~m[1317]&m[1363]&~m[1364]&~m[1366]&m[1367])|(~m[1317]&~m[1363]&m[1364]&~m[1366]&m[1367])|(m[1317]&m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1317]&m[1363]&m[1364]&m[1366]&m[1367]))&UnbiasedRNG[505])|((m[1317]&~m[1363]&~m[1364]&m[1366]&~m[1367])|(~m[1317]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1317]&~m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1317]&m[1363]&~m[1364]&~m[1366]&m[1367])|(m[1317]&~m[1363]&m[1364]&~m[1366]&m[1367])|(~m[1317]&~m[1363]&~m[1364]&m[1366]&m[1367])|(m[1317]&~m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1317]&m[1363]&~m[1364]&m[1366]&m[1367])|(m[1317]&m[1363]&~m[1364]&m[1366]&m[1367])|(~m[1317]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1317]&~m[1363]&m[1364]&m[1366]&m[1367])|(m[1317]&m[1363]&m[1364]&m[1366]&m[1367]));
    m[1370] = (((m[1322]&~m[1368]&~m[1369]&~m[1371]&~m[1372])|(~m[1322]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1322]&m[1368]&~m[1369]&m[1371]&~m[1372])|(m[1322]&~m[1368]&m[1369]&m[1371]&~m[1372])|(~m[1322]&m[1368]&~m[1369]&~m[1371]&m[1372])|(~m[1322]&~m[1368]&m[1369]&~m[1371]&m[1372])|(m[1322]&m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1322]&m[1368]&m[1369]&m[1371]&m[1372]))&UnbiasedRNG[506])|((m[1322]&~m[1368]&~m[1369]&m[1371]&~m[1372])|(~m[1322]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1322]&~m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1322]&m[1368]&~m[1369]&~m[1371]&m[1372])|(m[1322]&~m[1368]&m[1369]&~m[1371]&m[1372])|(~m[1322]&~m[1368]&~m[1369]&m[1371]&m[1372])|(m[1322]&~m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1322]&m[1368]&~m[1369]&m[1371]&m[1372])|(m[1322]&m[1368]&~m[1369]&m[1371]&m[1372])|(~m[1322]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1322]&~m[1368]&m[1369]&m[1371]&m[1372])|(m[1322]&m[1368]&m[1369]&m[1371]&m[1372]));
    m[1375] = (((m[1327]&~m[1373]&~m[1374]&~m[1376]&~m[1377])|(~m[1327]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1327]&m[1373]&~m[1374]&m[1376]&~m[1377])|(m[1327]&~m[1373]&m[1374]&m[1376]&~m[1377])|(~m[1327]&m[1373]&~m[1374]&~m[1376]&m[1377])|(~m[1327]&~m[1373]&m[1374]&~m[1376]&m[1377])|(m[1327]&m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1327]&m[1373]&m[1374]&m[1376]&m[1377]))&UnbiasedRNG[507])|((m[1327]&~m[1373]&~m[1374]&m[1376]&~m[1377])|(~m[1327]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1327]&~m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1327]&m[1373]&~m[1374]&~m[1376]&m[1377])|(m[1327]&~m[1373]&m[1374]&~m[1376]&m[1377])|(~m[1327]&~m[1373]&~m[1374]&m[1376]&m[1377])|(m[1327]&~m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1327]&m[1373]&~m[1374]&m[1376]&m[1377])|(m[1327]&m[1373]&~m[1374]&m[1376]&m[1377])|(~m[1327]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1327]&~m[1373]&m[1374]&m[1376]&m[1377])|(m[1327]&m[1373]&m[1374]&m[1376]&m[1377]));
    m[1380] = (((m[1332]&~m[1378]&~m[1379]&~m[1381]&~m[1382])|(~m[1332]&~m[1378]&~m[1379]&m[1381]&~m[1382])|(m[1332]&m[1378]&~m[1379]&m[1381]&~m[1382])|(m[1332]&~m[1378]&m[1379]&m[1381]&~m[1382])|(~m[1332]&m[1378]&~m[1379]&~m[1381]&m[1382])|(~m[1332]&~m[1378]&m[1379]&~m[1381]&m[1382])|(m[1332]&m[1378]&m[1379]&~m[1381]&m[1382])|(~m[1332]&m[1378]&m[1379]&m[1381]&m[1382]))&UnbiasedRNG[508])|((m[1332]&~m[1378]&~m[1379]&m[1381]&~m[1382])|(~m[1332]&~m[1378]&~m[1379]&~m[1381]&m[1382])|(m[1332]&~m[1378]&~m[1379]&~m[1381]&m[1382])|(m[1332]&m[1378]&~m[1379]&~m[1381]&m[1382])|(m[1332]&~m[1378]&m[1379]&~m[1381]&m[1382])|(~m[1332]&~m[1378]&~m[1379]&m[1381]&m[1382])|(m[1332]&~m[1378]&~m[1379]&m[1381]&m[1382])|(~m[1332]&m[1378]&~m[1379]&m[1381]&m[1382])|(m[1332]&m[1378]&~m[1379]&m[1381]&m[1382])|(~m[1332]&~m[1378]&m[1379]&m[1381]&m[1382])|(m[1332]&~m[1378]&m[1379]&m[1381]&m[1382])|(m[1332]&m[1378]&m[1379]&m[1381]&m[1382]));
    m[1385] = (((m[1337]&~m[1383]&~m[1384]&~m[1386]&~m[1387])|(~m[1337]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1337]&m[1383]&~m[1384]&m[1386]&~m[1387])|(m[1337]&~m[1383]&m[1384]&m[1386]&~m[1387])|(~m[1337]&m[1383]&~m[1384]&~m[1386]&m[1387])|(~m[1337]&~m[1383]&m[1384]&~m[1386]&m[1387])|(m[1337]&m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1337]&m[1383]&m[1384]&m[1386]&m[1387]))&UnbiasedRNG[509])|((m[1337]&~m[1383]&~m[1384]&m[1386]&~m[1387])|(~m[1337]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1337]&~m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1337]&m[1383]&~m[1384]&~m[1386]&m[1387])|(m[1337]&~m[1383]&m[1384]&~m[1386]&m[1387])|(~m[1337]&~m[1383]&~m[1384]&m[1386]&m[1387])|(m[1337]&~m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1337]&m[1383]&~m[1384]&m[1386]&m[1387])|(m[1337]&m[1383]&~m[1384]&m[1386]&m[1387])|(~m[1337]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1337]&~m[1383]&m[1384]&m[1386]&m[1387])|(m[1337]&m[1383]&m[1384]&m[1386]&m[1387]));
    m[1390] = (((m[1342]&~m[1388]&~m[1389]&~m[1391]&~m[1392])|(~m[1342]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1342]&m[1388]&~m[1389]&m[1391]&~m[1392])|(m[1342]&~m[1388]&m[1389]&m[1391]&~m[1392])|(~m[1342]&m[1388]&~m[1389]&~m[1391]&m[1392])|(~m[1342]&~m[1388]&m[1389]&~m[1391]&m[1392])|(m[1342]&m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1342]&m[1388]&m[1389]&m[1391]&m[1392]))&UnbiasedRNG[510])|((m[1342]&~m[1388]&~m[1389]&m[1391]&~m[1392])|(~m[1342]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1342]&~m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1342]&m[1388]&~m[1389]&~m[1391]&m[1392])|(m[1342]&~m[1388]&m[1389]&~m[1391]&m[1392])|(~m[1342]&~m[1388]&~m[1389]&m[1391]&m[1392])|(m[1342]&~m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1342]&m[1388]&~m[1389]&m[1391]&m[1392])|(m[1342]&m[1388]&~m[1389]&m[1391]&m[1392])|(~m[1342]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1342]&~m[1388]&m[1389]&m[1391]&m[1392])|(m[1342]&m[1388]&m[1389]&m[1391]&m[1392]));
    m[1395] = (((m[1347]&~m[1393]&~m[1394]&~m[1396]&~m[1397])|(~m[1347]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1347]&m[1393]&~m[1394]&m[1396]&~m[1397])|(m[1347]&~m[1393]&m[1394]&m[1396]&~m[1397])|(~m[1347]&m[1393]&~m[1394]&~m[1396]&m[1397])|(~m[1347]&~m[1393]&m[1394]&~m[1396]&m[1397])|(m[1347]&m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1347]&m[1393]&m[1394]&m[1396]&m[1397]))&UnbiasedRNG[511])|((m[1347]&~m[1393]&~m[1394]&m[1396]&~m[1397])|(~m[1347]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1347]&~m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1347]&m[1393]&~m[1394]&~m[1396]&m[1397])|(m[1347]&~m[1393]&m[1394]&~m[1396]&m[1397])|(~m[1347]&~m[1393]&~m[1394]&m[1396]&m[1397])|(m[1347]&~m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1347]&m[1393]&~m[1394]&m[1396]&m[1397])|(m[1347]&m[1393]&~m[1394]&m[1396]&m[1397])|(~m[1347]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1347]&~m[1393]&m[1394]&m[1396]&m[1397])|(m[1347]&m[1393]&m[1394]&m[1396]&m[1397]));
    m[1400] = (((m[1352]&~m[1398]&~m[1399]&~m[1401]&~m[1402])|(~m[1352]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1352]&m[1398]&~m[1399]&m[1401]&~m[1402])|(m[1352]&~m[1398]&m[1399]&m[1401]&~m[1402])|(~m[1352]&m[1398]&~m[1399]&~m[1401]&m[1402])|(~m[1352]&~m[1398]&m[1399]&~m[1401]&m[1402])|(m[1352]&m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1352]&m[1398]&m[1399]&m[1401]&m[1402]))&UnbiasedRNG[512])|((m[1352]&~m[1398]&~m[1399]&m[1401]&~m[1402])|(~m[1352]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1352]&~m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1352]&m[1398]&~m[1399]&~m[1401]&m[1402])|(m[1352]&~m[1398]&m[1399]&~m[1401]&m[1402])|(~m[1352]&~m[1398]&~m[1399]&m[1401]&m[1402])|(m[1352]&~m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1352]&m[1398]&~m[1399]&m[1401]&m[1402])|(m[1352]&m[1398]&~m[1399]&m[1401]&m[1402])|(~m[1352]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1352]&~m[1398]&m[1399]&m[1401]&m[1402])|(m[1352]&m[1398]&m[1399]&m[1401]&m[1402]));
    m[1405] = (((m[1357]&~m[1403]&~m[1404]&~m[1406]&~m[1407])|(~m[1357]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1357]&m[1403]&~m[1404]&m[1406]&~m[1407])|(m[1357]&~m[1403]&m[1404]&m[1406]&~m[1407])|(~m[1357]&m[1403]&~m[1404]&~m[1406]&m[1407])|(~m[1357]&~m[1403]&m[1404]&~m[1406]&m[1407])|(m[1357]&m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1357]&m[1403]&m[1404]&m[1406]&m[1407]))&UnbiasedRNG[513])|((m[1357]&~m[1403]&~m[1404]&m[1406]&~m[1407])|(~m[1357]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1357]&~m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1357]&m[1403]&~m[1404]&~m[1406]&m[1407])|(m[1357]&~m[1403]&m[1404]&~m[1406]&m[1407])|(~m[1357]&~m[1403]&~m[1404]&m[1406]&m[1407])|(m[1357]&~m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1357]&m[1403]&~m[1404]&m[1406]&m[1407])|(m[1357]&m[1403]&~m[1404]&m[1406]&m[1407])|(~m[1357]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1357]&~m[1403]&m[1404]&m[1406]&m[1407])|(m[1357]&m[1403]&m[1404]&m[1406]&m[1407]));
    m[1410] = (((m[1362]&~m[1408]&~m[1409]&~m[1411]&~m[1412])|(~m[1362]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1362]&m[1408]&~m[1409]&m[1411]&~m[1412])|(m[1362]&~m[1408]&m[1409]&m[1411]&~m[1412])|(~m[1362]&m[1408]&~m[1409]&~m[1411]&m[1412])|(~m[1362]&~m[1408]&m[1409]&~m[1411]&m[1412])|(m[1362]&m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1362]&m[1408]&m[1409]&m[1411]&m[1412]))&UnbiasedRNG[514])|((m[1362]&~m[1408]&~m[1409]&m[1411]&~m[1412])|(~m[1362]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1362]&~m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1362]&m[1408]&~m[1409]&~m[1411]&m[1412])|(m[1362]&~m[1408]&m[1409]&~m[1411]&m[1412])|(~m[1362]&~m[1408]&~m[1409]&m[1411]&m[1412])|(m[1362]&~m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1362]&m[1408]&~m[1409]&m[1411]&m[1412])|(m[1362]&m[1408]&~m[1409]&m[1411]&m[1412])|(~m[1362]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1362]&~m[1408]&m[1409]&m[1411]&m[1412])|(m[1362]&m[1408]&m[1409]&m[1411]&m[1412]));
    m[1415] = (((m[1372]&~m[1413]&~m[1414]&~m[1416]&~m[1417])|(~m[1372]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1372]&m[1413]&~m[1414]&m[1416]&~m[1417])|(m[1372]&~m[1413]&m[1414]&m[1416]&~m[1417])|(~m[1372]&m[1413]&~m[1414]&~m[1416]&m[1417])|(~m[1372]&~m[1413]&m[1414]&~m[1416]&m[1417])|(m[1372]&m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1372]&m[1413]&m[1414]&m[1416]&m[1417]))&UnbiasedRNG[515])|((m[1372]&~m[1413]&~m[1414]&m[1416]&~m[1417])|(~m[1372]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1372]&~m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1372]&m[1413]&~m[1414]&~m[1416]&m[1417])|(m[1372]&~m[1413]&m[1414]&~m[1416]&m[1417])|(~m[1372]&~m[1413]&~m[1414]&m[1416]&m[1417])|(m[1372]&~m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1372]&m[1413]&~m[1414]&m[1416]&m[1417])|(m[1372]&m[1413]&~m[1414]&m[1416]&m[1417])|(~m[1372]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1372]&~m[1413]&m[1414]&m[1416]&m[1417])|(m[1372]&m[1413]&m[1414]&m[1416]&m[1417]));
    m[1420] = (((m[1377]&~m[1418]&~m[1419]&~m[1421]&~m[1422])|(~m[1377]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1377]&m[1418]&~m[1419]&m[1421]&~m[1422])|(m[1377]&~m[1418]&m[1419]&m[1421]&~m[1422])|(~m[1377]&m[1418]&~m[1419]&~m[1421]&m[1422])|(~m[1377]&~m[1418]&m[1419]&~m[1421]&m[1422])|(m[1377]&m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1377]&m[1418]&m[1419]&m[1421]&m[1422]))&UnbiasedRNG[516])|((m[1377]&~m[1418]&~m[1419]&m[1421]&~m[1422])|(~m[1377]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1377]&~m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1377]&m[1418]&~m[1419]&~m[1421]&m[1422])|(m[1377]&~m[1418]&m[1419]&~m[1421]&m[1422])|(~m[1377]&~m[1418]&~m[1419]&m[1421]&m[1422])|(m[1377]&~m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1377]&m[1418]&~m[1419]&m[1421]&m[1422])|(m[1377]&m[1418]&~m[1419]&m[1421]&m[1422])|(~m[1377]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1377]&~m[1418]&m[1419]&m[1421]&m[1422])|(m[1377]&m[1418]&m[1419]&m[1421]&m[1422]));
    m[1425] = (((m[1382]&~m[1423]&~m[1424]&~m[1426]&~m[1427])|(~m[1382]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1382]&m[1423]&~m[1424]&m[1426]&~m[1427])|(m[1382]&~m[1423]&m[1424]&m[1426]&~m[1427])|(~m[1382]&m[1423]&~m[1424]&~m[1426]&m[1427])|(~m[1382]&~m[1423]&m[1424]&~m[1426]&m[1427])|(m[1382]&m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1382]&m[1423]&m[1424]&m[1426]&m[1427]))&UnbiasedRNG[517])|((m[1382]&~m[1423]&~m[1424]&m[1426]&~m[1427])|(~m[1382]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1382]&~m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1382]&m[1423]&~m[1424]&~m[1426]&m[1427])|(m[1382]&~m[1423]&m[1424]&~m[1426]&m[1427])|(~m[1382]&~m[1423]&~m[1424]&m[1426]&m[1427])|(m[1382]&~m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1382]&m[1423]&~m[1424]&m[1426]&m[1427])|(m[1382]&m[1423]&~m[1424]&m[1426]&m[1427])|(~m[1382]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1382]&~m[1423]&m[1424]&m[1426]&m[1427])|(m[1382]&m[1423]&m[1424]&m[1426]&m[1427]));
    m[1430] = (((m[1387]&~m[1428]&~m[1429]&~m[1431]&~m[1432])|(~m[1387]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1387]&m[1428]&~m[1429]&m[1431]&~m[1432])|(m[1387]&~m[1428]&m[1429]&m[1431]&~m[1432])|(~m[1387]&m[1428]&~m[1429]&~m[1431]&m[1432])|(~m[1387]&~m[1428]&m[1429]&~m[1431]&m[1432])|(m[1387]&m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1387]&m[1428]&m[1429]&m[1431]&m[1432]))&UnbiasedRNG[518])|((m[1387]&~m[1428]&~m[1429]&m[1431]&~m[1432])|(~m[1387]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1387]&~m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1387]&m[1428]&~m[1429]&~m[1431]&m[1432])|(m[1387]&~m[1428]&m[1429]&~m[1431]&m[1432])|(~m[1387]&~m[1428]&~m[1429]&m[1431]&m[1432])|(m[1387]&~m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1387]&m[1428]&~m[1429]&m[1431]&m[1432])|(m[1387]&m[1428]&~m[1429]&m[1431]&m[1432])|(~m[1387]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1387]&~m[1428]&m[1429]&m[1431]&m[1432])|(m[1387]&m[1428]&m[1429]&m[1431]&m[1432]));
    m[1435] = (((m[1392]&~m[1433]&~m[1434]&~m[1436]&~m[1437])|(~m[1392]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1392]&m[1433]&~m[1434]&m[1436]&~m[1437])|(m[1392]&~m[1433]&m[1434]&m[1436]&~m[1437])|(~m[1392]&m[1433]&~m[1434]&~m[1436]&m[1437])|(~m[1392]&~m[1433]&m[1434]&~m[1436]&m[1437])|(m[1392]&m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1392]&m[1433]&m[1434]&m[1436]&m[1437]))&UnbiasedRNG[519])|((m[1392]&~m[1433]&~m[1434]&m[1436]&~m[1437])|(~m[1392]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1392]&~m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1392]&m[1433]&~m[1434]&~m[1436]&m[1437])|(m[1392]&~m[1433]&m[1434]&~m[1436]&m[1437])|(~m[1392]&~m[1433]&~m[1434]&m[1436]&m[1437])|(m[1392]&~m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1392]&m[1433]&~m[1434]&m[1436]&m[1437])|(m[1392]&m[1433]&~m[1434]&m[1436]&m[1437])|(~m[1392]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1392]&~m[1433]&m[1434]&m[1436]&m[1437])|(m[1392]&m[1433]&m[1434]&m[1436]&m[1437]));
    m[1440] = (((m[1397]&~m[1438]&~m[1439]&~m[1441]&~m[1442])|(~m[1397]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1397]&m[1438]&~m[1439]&m[1441]&~m[1442])|(m[1397]&~m[1438]&m[1439]&m[1441]&~m[1442])|(~m[1397]&m[1438]&~m[1439]&~m[1441]&m[1442])|(~m[1397]&~m[1438]&m[1439]&~m[1441]&m[1442])|(m[1397]&m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1397]&m[1438]&m[1439]&m[1441]&m[1442]))&UnbiasedRNG[520])|((m[1397]&~m[1438]&~m[1439]&m[1441]&~m[1442])|(~m[1397]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1397]&~m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1397]&m[1438]&~m[1439]&~m[1441]&m[1442])|(m[1397]&~m[1438]&m[1439]&~m[1441]&m[1442])|(~m[1397]&~m[1438]&~m[1439]&m[1441]&m[1442])|(m[1397]&~m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1397]&m[1438]&~m[1439]&m[1441]&m[1442])|(m[1397]&m[1438]&~m[1439]&m[1441]&m[1442])|(~m[1397]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1397]&~m[1438]&m[1439]&m[1441]&m[1442])|(m[1397]&m[1438]&m[1439]&m[1441]&m[1442]));
    m[1445] = (((m[1402]&~m[1443]&~m[1444]&~m[1446]&~m[1447])|(~m[1402]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1402]&m[1443]&~m[1444]&m[1446]&~m[1447])|(m[1402]&~m[1443]&m[1444]&m[1446]&~m[1447])|(~m[1402]&m[1443]&~m[1444]&~m[1446]&m[1447])|(~m[1402]&~m[1443]&m[1444]&~m[1446]&m[1447])|(m[1402]&m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1402]&m[1443]&m[1444]&m[1446]&m[1447]))&UnbiasedRNG[521])|((m[1402]&~m[1443]&~m[1444]&m[1446]&~m[1447])|(~m[1402]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1402]&~m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1402]&m[1443]&~m[1444]&~m[1446]&m[1447])|(m[1402]&~m[1443]&m[1444]&~m[1446]&m[1447])|(~m[1402]&~m[1443]&~m[1444]&m[1446]&m[1447])|(m[1402]&~m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1402]&m[1443]&~m[1444]&m[1446]&m[1447])|(m[1402]&m[1443]&~m[1444]&m[1446]&m[1447])|(~m[1402]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1402]&~m[1443]&m[1444]&m[1446]&m[1447])|(m[1402]&m[1443]&m[1444]&m[1446]&m[1447]));
    m[1450] = (((m[1407]&~m[1448]&~m[1449]&~m[1451]&~m[1452])|(~m[1407]&~m[1448]&~m[1449]&m[1451]&~m[1452])|(m[1407]&m[1448]&~m[1449]&m[1451]&~m[1452])|(m[1407]&~m[1448]&m[1449]&m[1451]&~m[1452])|(~m[1407]&m[1448]&~m[1449]&~m[1451]&m[1452])|(~m[1407]&~m[1448]&m[1449]&~m[1451]&m[1452])|(m[1407]&m[1448]&m[1449]&~m[1451]&m[1452])|(~m[1407]&m[1448]&m[1449]&m[1451]&m[1452]))&UnbiasedRNG[522])|((m[1407]&~m[1448]&~m[1449]&m[1451]&~m[1452])|(~m[1407]&~m[1448]&~m[1449]&~m[1451]&m[1452])|(m[1407]&~m[1448]&~m[1449]&~m[1451]&m[1452])|(m[1407]&m[1448]&~m[1449]&~m[1451]&m[1452])|(m[1407]&~m[1448]&m[1449]&~m[1451]&m[1452])|(~m[1407]&~m[1448]&~m[1449]&m[1451]&m[1452])|(m[1407]&~m[1448]&~m[1449]&m[1451]&m[1452])|(~m[1407]&m[1448]&~m[1449]&m[1451]&m[1452])|(m[1407]&m[1448]&~m[1449]&m[1451]&m[1452])|(~m[1407]&~m[1448]&m[1449]&m[1451]&m[1452])|(m[1407]&~m[1448]&m[1449]&m[1451]&m[1452])|(m[1407]&m[1448]&m[1449]&m[1451]&m[1452]));
    m[1455] = (((m[1412]&~m[1453]&~m[1454]&~m[1456]&~m[1457])|(~m[1412]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1412]&m[1453]&~m[1454]&m[1456]&~m[1457])|(m[1412]&~m[1453]&m[1454]&m[1456]&~m[1457])|(~m[1412]&m[1453]&~m[1454]&~m[1456]&m[1457])|(~m[1412]&~m[1453]&m[1454]&~m[1456]&m[1457])|(m[1412]&m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1412]&m[1453]&m[1454]&m[1456]&m[1457]))&UnbiasedRNG[523])|((m[1412]&~m[1453]&~m[1454]&m[1456]&~m[1457])|(~m[1412]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1412]&~m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1412]&m[1453]&~m[1454]&~m[1456]&m[1457])|(m[1412]&~m[1453]&m[1454]&~m[1456]&m[1457])|(~m[1412]&~m[1453]&~m[1454]&m[1456]&m[1457])|(m[1412]&~m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1412]&m[1453]&~m[1454]&m[1456]&m[1457])|(m[1412]&m[1453]&~m[1454]&m[1456]&m[1457])|(~m[1412]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1412]&~m[1453]&m[1454]&m[1456]&m[1457])|(m[1412]&m[1453]&m[1454]&m[1456]&m[1457]));
    m[1460] = (((m[1422]&~m[1458]&~m[1459]&~m[1461]&~m[1462])|(~m[1422]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1422]&m[1458]&~m[1459]&m[1461]&~m[1462])|(m[1422]&~m[1458]&m[1459]&m[1461]&~m[1462])|(~m[1422]&m[1458]&~m[1459]&~m[1461]&m[1462])|(~m[1422]&~m[1458]&m[1459]&~m[1461]&m[1462])|(m[1422]&m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1422]&m[1458]&m[1459]&m[1461]&m[1462]))&UnbiasedRNG[524])|((m[1422]&~m[1458]&~m[1459]&m[1461]&~m[1462])|(~m[1422]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1422]&~m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1422]&m[1458]&~m[1459]&~m[1461]&m[1462])|(m[1422]&~m[1458]&m[1459]&~m[1461]&m[1462])|(~m[1422]&~m[1458]&~m[1459]&m[1461]&m[1462])|(m[1422]&~m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1422]&m[1458]&~m[1459]&m[1461]&m[1462])|(m[1422]&m[1458]&~m[1459]&m[1461]&m[1462])|(~m[1422]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1422]&~m[1458]&m[1459]&m[1461]&m[1462])|(m[1422]&m[1458]&m[1459]&m[1461]&m[1462]));
    m[1465] = (((m[1427]&~m[1463]&~m[1464]&~m[1466]&~m[1467])|(~m[1427]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1427]&m[1463]&~m[1464]&m[1466]&~m[1467])|(m[1427]&~m[1463]&m[1464]&m[1466]&~m[1467])|(~m[1427]&m[1463]&~m[1464]&~m[1466]&m[1467])|(~m[1427]&~m[1463]&m[1464]&~m[1466]&m[1467])|(m[1427]&m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1427]&m[1463]&m[1464]&m[1466]&m[1467]))&UnbiasedRNG[525])|((m[1427]&~m[1463]&~m[1464]&m[1466]&~m[1467])|(~m[1427]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1427]&~m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1427]&m[1463]&~m[1464]&~m[1466]&m[1467])|(m[1427]&~m[1463]&m[1464]&~m[1466]&m[1467])|(~m[1427]&~m[1463]&~m[1464]&m[1466]&m[1467])|(m[1427]&~m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1427]&m[1463]&~m[1464]&m[1466]&m[1467])|(m[1427]&m[1463]&~m[1464]&m[1466]&m[1467])|(~m[1427]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1427]&~m[1463]&m[1464]&m[1466]&m[1467])|(m[1427]&m[1463]&m[1464]&m[1466]&m[1467]));
    m[1470] = (((m[1432]&~m[1468]&~m[1469]&~m[1471]&~m[1472])|(~m[1432]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1432]&m[1468]&~m[1469]&m[1471]&~m[1472])|(m[1432]&~m[1468]&m[1469]&m[1471]&~m[1472])|(~m[1432]&m[1468]&~m[1469]&~m[1471]&m[1472])|(~m[1432]&~m[1468]&m[1469]&~m[1471]&m[1472])|(m[1432]&m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1432]&m[1468]&m[1469]&m[1471]&m[1472]))&UnbiasedRNG[526])|((m[1432]&~m[1468]&~m[1469]&m[1471]&~m[1472])|(~m[1432]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1432]&~m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1432]&m[1468]&~m[1469]&~m[1471]&m[1472])|(m[1432]&~m[1468]&m[1469]&~m[1471]&m[1472])|(~m[1432]&~m[1468]&~m[1469]&m[1471]&m[1472])|(m[1432]&~m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1432]&m[1468]&~m[1469]&m[1471]&m[1472])|(m[1432]&m[1468]&~m[1469]&m[1471]&m[1472])|(~m[1432]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1432]&~m[1468]&m[1469]&m[1471]&m[1472])|(m[1432]&m[1468]&m[1469]&m[1471]&m[1472]));
    m[1475] = (((m[1437]&~m[1473]&~m[1474]&~m[1476]&~m[1477])|(~m[1437]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1437]&m[1473]&~m[1474]&m[1476]&~m[1477])|(m[1437]&~m[1473]&m[1474]&m[1476]&~m[1477])|(~m[1437]&m[1473]&~m[1474]&~m[1476]&m[1477])|(~m[1437]&~m[1473]&m[1474]&~m[1476]&m[1477])|(m[1437]&m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1437]&m[1473]&m[1474]&m[1476]&m[1477]))&UnbiasedRNG[527])|((m[1437]&~m[1473]&~m[1474]&m[1476]&~m[1477])|(~m[1437]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1437]&~m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1437]&m[1473]&~m[1474]&~m[1476]&m[1477])|(m[1437]&~m[1473]&m[1474]&~m[1476]&m[1477])|(~m[1437]&~m[1473]&~m[1474]&m[1476]&m[1477])|(m[1437]&~m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1437]&m[1473]&~m[1474]&m[1476]&m[1477])|(m[1437]&m[1473]&~m[1474]&m[1476]&m[1477])|(~m[1437]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1437]&~m[1473]&m[1474]&m[1476]&m[1477])|(m[1437]&m[1473]&m[1474]&m[1476]&m[1477]));
    m[1480] = (((m[1442]&~m[1478]&~m[1479]&~m[1481]&~m[1482])|(~m[1442]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1442]&m[1478]&~m[1479]&m[1481]&~m[1482])|(m[1442]&~m[1478]&m[1479]&m[1481]&~m[1482])|(~m[1442]&m[1478]&~m[1479]&~m[1481]&m[1482])|(~m[1442]&~m[1478]&m[1479]&~m[1481]&m[1482])|(m[1442]&m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1442]&m[1478]&m[1479]&m[1481]&m[1482]))&UnbiasedRNG[528])|((m[1442]&~m[1478]&~m[1479]&m[1481]&~m[1482])|(~m[1442]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1442]&~m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1442]&m[1478]&~m[1479]&~m[1481]&m[1482])|(m[1442]&~m[1478]&m[1479]&~m[1481]&m[1482])|(~m[1442]&~m[1478]&~m[1479]&m[1481]&m[1482])|(m[1442]&~m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1442]&m[1478]&~m[1479]&m[1481]&m[1482])|(m[1442]&m[1478]&~m[1479]&m[1481]&m[1482])|(~m[1442]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1442]&~m[1478]&m[1479]&m[1481]&m[1482])|(m[1442]&m[1478]&m[1479]&m[1481]&m[1482]));
    m[1485] = (((m[1447]&~m[1483]&~m[1484]&~m[1486]&~m[1487])|(~m[1447]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1447]&m[1483]&~m[1484]&m[1486]&~m[1487])|(m[1447]&~m[1483]&m[1484]&m[1486]&~m[1487])|(~m[1447]&m[1483]&~m[1484]&~m[1486]&m[1487])|(~m[1447]&~m[1483]&m[1484]&~m[1486]&m[1487])|(m[1447]&m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1447]&m[1483]&m[1484]&m[1486]&m[1487]))&UnbiasedRNG[529])|((m[1447]&~m[1483]&~m[1484]&m[1486]&~m[1487])|(~m[1447]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1447]&~m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1447]&m[1483]&~m[1484]&~m[1486]&m[1487])|(m[1447]&~m[1483]&m[1484]&~m[1486]&m[1487])|(~m[1447]&~m[1483]&~m[1484]&m[1486]&m[1487])|(m[1447]&~m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1447]&m[1483]&~m[1484]&m[1486]&m[1487])|(m[1447]&m[1483]&~m[1484]&m[1486]&m[1487])|(~m[1447]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1447]&~m[1483]&m[1484]&m[1486]&m[1487])|(m[1447]&m[1483]&m[1484]&m[1486]&m[1487]));
    m[1490] = (((m[1452]&~m[1488]&~m[1489]&~m[1491]&~m[1492])|(~m[1452]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1452]&m[1488]&~m[1489]&m[1491]&~m[1492])|(m[1452]&~m[1488]&m[1489]&m[1491]&~m[1492])|(~m[1452]&m[1488]&~m[1489]&~m[1491]&m[1492])|(~m[1452]&~m[1488]&m[1489]&~m[1491]&m[1492])|(m[1452]&m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1452]&m[1488]&m[1489]&m[1491]&m[1492]))&UnbiasedRNG[530])|((m[1452]&~m[1488]&~m[1489]&m[1491]&~m[1492])|(~m[1452]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1452]&~m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1452]&m[1488]&~m[1489]&~m[1491]&m[1492])|(m[1452]&~m[1488]&m[1489]&~m[1491]&m[1492])|(~m[1452]&~m[1488]&~m[1489]&m[1491]&m[1492])|(m[1452]&~m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1452]&m[1488]&~m[1489]&m[1491]&m[1492])|(m[1452]&m[1488]&~m[1489]&m[1491]&m[1492])|(~m[1452]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1452]&~m[1488]&m[1489]&m[1491]&m[1492])|(m[1452]&m[1488]&m[1489]&m[1491]&m[1492]));
    m[1495] = (((m[1457]&~m[1493]&~m[1494]&~m[1496]&~m[1497])|(~m[1457]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1457]&m[1493]&~m[1494]&m[1496]&~m[1497])|(m[1457]&~m[1493]&m[1494]&m[1496]&~m[1497])|(~m[1457]&m[1493]&~m[1494]&~m[1496]&m[1497])|(~m[1457]&~m[1493]&m[1494]&~m[1496]&m[1497])|(m[1457]&m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1457]&m[1493]&m[1494]&m[1496]&m[1497]))&UnbiasedRNG[531])|((m[1457]&~m[1493]&~m[1494]&m[1496]&~m[1497])|(~m[1457]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1457]&~m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1457]&m[1493]&~m[1494]&~m[1496]&m[1497])|(m[1457]&~m[1493]&m[1494]&~m[1496]&m[1497])|(~m[1457]&~m[1493]&~m[1494]&m[1496]&m[1497])|(m[1457]&~m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1457]&m[1493]&~m[1494]&m[1496]&m[1497])|(m[1457]&m[1493]&~m[1494]&m[1496]&m[1497])|(~m[1457]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1457]&~m[1493]&m[1494]&m[1496]&m[1497])|(m[1457]&m[1493]&m[1494]&m[1496]&m[1497]));
    m[1500] = (((m[1467]&~m[1498]&~m[1499]&~m[1501]&~m[1502])|(~m[1467]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1467]&m[1498]&~m[1499]&m[1501]&~m[1502])|(m[1467]&~m[1498]&m[1499]&m[1501]&~m[1502])|(~m[1467]&m[1498]&~m[1499]&~m[1501]&m[1502])|(~m[1467]&~m[1498]&m[1499]&~m[1501]&m[1502])|(m[1467]&m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1467]&m[1498]&m[1499]&m[1501]&m[1502]))&UnbiasedRNG[532])|((m[1467]&~m[1498]&~m[1499]&m[1501]&~m[1502])|(~m[1467]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1467]&~m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1467]&m[1498]&~m[1499]&~m[1501]&m[1502])|(m[1467]&~m[1498]&m[1499]&~m[1501]&m[1502])|(~m[1467]&~m[1498]&~m[1499]&m[1501]&m[1502])|(m[1467]&~m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1467]&m[1498]&~m[1499]&m[1501]&m[1502])|(m[1467]&m[1498]&~m[1499]&m[1501]&m[1502])|(~m[1467]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1467]&~m[1498]&m[1499]&m[1501]&m[1502])|(m[1467]&m[1498]&m[1499]&m[1501]&m[1502]));
    m[1505] = (((m[1472]&~m[1503]&~m[1504]&~m[1506]&~m[1507])|(~m[1472]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1472]&m[1503]&~m[1504]&m[1506]&~m[1507])|(m[1472]&~m[1503]&m[1504]&m[1506]&~m[1507])|(~m[1472]&m[1503]&~m[1504]&~m[1506]&m[1507])|(~m[1472]&~m[1503]&m[1504]&~m[1506]&m[1507])|(m[1472]&m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1472]&m[1503]&m[1504]&m[1506]&m[1507]))&UnbiasedRNG[533])|((m[1472]&~m[1503]&~m[1504]&m[1506]&~m[1507])|(~m[1472]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1472]&~m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1472]&m[1503]&~m[1504]&~m[1506]&m[1507])|(m[1472]&~m[1503]&m[1504]&~m[1506]&m[1507])|(~m[1472]&~m[1503]&~m[1504]&m[1506]&m[1507])|(m[1472]&~m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1472]&m[1503]&~m[1504]&m[1506]&m[1507])|(m[1472]&m[1503]&~m[1504]&m[1506]&m[1507])|(~m[1472]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1472]&~m[1503]&m[1504]&m[1506]&m[1507])|(m[1472]&m[1503]&m[1504]&m[1506]&m[1507]));
    m[1510] = (((m[1477]&~m[1508]&~m[1509]&~m[1511]&~m[1512])|(~m[1477]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1477]&m[1508]&~m[1509]&m[1511]&~m[1512])|(m[1477]&~m[1508]&m[1509]&m[1511]&~m[1512])|(~m[1477]&m[1508]&~m[1509]&~m[1511]&m[1512])|(~m[1477]&~m[1508]&m[1509]&~m[1511]&m[1512])|(m[1477]&m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1477]&m[1508]&m[1509]&m[1511]&m[1512]))&UnbiasedRNG[534])|((m[1477]&~m[1508]&~m[1509]&m[1511]&~m[1512])|(~m[1477]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1477]&~m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1477]&m[1508]&~m[1509]&~m[1511]&m[1512])|(m[1477]&~m[1508]&m[1509]&~m[1511]&m[1512])|(~m[1477]&~m[1508]&~m[1509]&m[1511]&m[1512])|(m[1477]&~m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1477]&m[1508]&~m[1509]&m[1511]&m[1512])|(m[1477]&m[1508]&~m[1509]&m[1511]&m[1512])|(~m[1477]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1477]&~m[1508]&m[1509]&m[1511]&m[1512])|(m[1477]&m[1508]&m[1509]&m[1511]&m[1512]));
    m[1515] = (((m[1482]&~m[1513]&~m[1514]&~m[1516]&~m[1517])|(~m[1482]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1482]&m[1513]&~m[1514]&m[1516]&~m[1517])|(m[1482]&~m[1513]&m[1514]&m[1516]&~m[1517])|(~m[1482]&m[1513]&~m[1514]&~m[1516]&m[1517])|(~m[1482]&~m[1513]&m[1514]&~m[1516]&m[1517])|(m[1482]&m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1482]&m[1513]&m[1514]&m[1516]&m[1517]))&UnbiasedRNG[535])|((m[1482]&~m[1513]&~m[1514]&m[1516]&~m[1517])|(~m[1482]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1482]&~m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1482]&m[1513]&~m[1514]&~m[1516]&m[1517])|(m[1482]&~m[1513]&m[1514]&~m[1516]&m[1517])|(~m[1482]&~m[1513]&~m[1514]&m[1516]&m[1517])|(m[1482]&~m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1482]&m[1513]&~m[1514]&m[1516]&m[1517])|(m[1482]&m[1513]&~m[1514]&m[1516]&m[1517])|(~m[1482]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1482]&~m[1513]&m[1514]&m[1516]&m[1517])|(m[1482]&m[1513]&m[1514]&m[1516]&m[1517]));
    m[1520] = (((m[1487]&~m[1518]&~m[1519]&~m[1521]&~m[1522])|(~m[1487]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1487]&m[1518]&~m[1519]&m[1521]&~m[1522])|(m[1487]&~m[1518]&m[1519]&m[1521]&~m[1522])|(~m[1487]&m[1518]&~m[1519]&~m[1521]&m[1522])|(~m[1487]&~m[1518]&m[1519]&~m[1521]&m[1522])|(m[1487]&m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1487]&m[1518]&m[1519]&m[1521]&m[1522]))&UnbiasedRNG[536])|((m[1487]&~m[1518]&~m[1519]&m[1521]&~m[1522])|(~m[1487]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1487]&~m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1487]&m[1518]&~m[1519]&~m[1521]&m[1522])|(m[1487]&~m[1518]&m[1519]&~m[1521]&m[1522])|(~m[1487]&~m[1518]&~m[1519]&m[1521]&m[1522])|(m[1487]&~m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1487]&m[1518]&~m[1519]&m[1521]&m[1522])|(m[1487]&m[1518]&~m[1519]&m[1521]&m[1522])|(~m[1487]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1487]&~m[1518]&m[1519]&m[1521]&m[1522])|(m[1487]&m[1518]&m[1519]&m[1521]&m[1522]));
    m[1525] = (((m[1492]&~m[1523]&~m[1524]&~m[1526]&~m[1527])|(~m[1492]&~m[1523]&~m[1524]&m[1526]&~m[1527])|(m[1492]&m[1523]&~m[1524]&m[1526]&~m[1527])|(m[1492]&~m[1523]&m[1524]&m[1526]&~m[1527])|(~m[1492]&m[1523]&~m[1524]&~m[1526]&m[1527])|(~m[1492]&~m[1523]&m[1524]&~m[1526]&m[1527])|(m[1492]&m[1523]&m[1524]&~m[1526]&m[1527])|(~m[1492]&m[1523]&m[1524]&m[1526]&m[1527]))&UnbiasedRNG[537])|((m[1492]&~m[1523]&~m[1524]&m[1526]&~m[1527])|(~m[1492]&~m[1523]&~m[1524]&~m[1526]&m[1527])|(m[1492]&~m[1523]&~m[1524]&~m[1526]&m[1527])|(m[1492]&m[1523]&~m[1524]&~m[1526]&m[1527])|(m[1492]&~m[1523]&m[1524]&~m[1526]&m[1527])|(~m[1492]&~m[1523]&~m[1524]&m[1526]&m[1527])|(m[1492]&~m[1523]&~m[1524]&m[1526]&m[1527])|(~m[1492]&m[1523]&~m[1524]&m[1526]&m[1527])|(m[1492]&m[1523]&~m[1524]&m[1526]&m[1527])|(~m[1492]&~m[1523]&m[1524]&m[1526]&m[1527])|(m[1492]&~m[1523]&m[1524]&m[1526]&m[1527])|(m[1492]&m[1523]&m[1524]&m[1526]&m[1527]));
    m[1530] = (((m[1497]&~m[1528]&~m[1529]&~m[1531]&~m[1532])|(~m[1497]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1497]&m[1528]&~m[1529]&m[1531]&~m[1532])|(m[1497]&~m[1528]&m[1529]&m[1531]&~m[1532])|(~m[1497]&m[1528]&~m[1529]&~m[1531]&m[1532])|(~m[1497]&~m[1528]&m[1529]&~m[1531]&m[1532])|(m[1497]&m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1497]&m[1528]&m[1529]&m[1531]&m[1532]))&UnbiasedRNG[538])|((m[1497]&~m[1528]&~m[1529]&m[1531]&~m[1532])|(~m[1497]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1497]&~m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1497]&m[1528]&~m[1529]&~m[1531]&m[1532])|(m[1497]&~m[1528]&m[1529]&~m[1531]&m[1532])|(~m[1497]&~m[1528]&~m[1529]&m[1531]&m[1532])|(m[1497]&~m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1497]&m[1528]&~m[1529]&m[1531]&m[1532])|(m[1497]&m[1528]&~m[1529]&m[1531]&m[1532])|(~m[1497]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1497]&~m[1528]&m[1529]&m[1531]&m[1532])|(m[1497]&m[1528]&m[1529]&m[1531]&m[1532]));
    m[1535] = (((m[1507]&~m[1533]&~m[1534]&~m[1536]&~m[1537])|(~m[1507]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1507]&m[1533]&~m[1534]&m[1536]&~m[1537])|(m[1507]&~m[1533]&m[1534]&m[1536]&~m[1537])|(~m[1507]&m[1533]&~m[1534]&~m[1536]&m[1537])|(~m[1507]&~m[1533]&m[1534]&~m[1536]&m[1537])|(m[1507]&m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1507]&m[1533]&m[1534]&m[1536]&m[1537]))&UnbiasedRNG[539])|((m[1507]&~m[1533]&~m[1534]&m[1536]&~m[1537])|(~m[1507]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1507]&~m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1507]&m[1533]&~m[1534]&~m[1536]&m[1537])|(m[1507]&~m[1533]&m[1534]&~m[1536]&m[1537])|(~m[1507]&~m[1533]&~m[1534]&m[1536]&m[1537])|(m[1507]&~m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1507]&m[1533]&~m[1534]&m[1536]&m[1537])|(m[1507]&m[1533]&~m[1534]&m[1536]&m[1537])|(~m[1507]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1507]&~m[1533]&m[1534]&m[1536]&m[1537])|(m[1507]&m[1533]&m[1534]&m[1536]&m[1537]));
    m[1540] = (((m[1512]&~m[1538]&~m[1539]&~m[1541]&~m[1542])|(~m[1512]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1512]&m[1538]&~m[1539]&m[1541]&~m[1542])|(m[1512]&~m[1538]&m[1539]&m[1541]&~m[1542])|(~m[1512]&m[1538]&~m[1539]&~m[1541]&m[1542])|(~m[1512]&~m[1538]&m[1539]&~m[1541]&m[1542])|(m[1512]&m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1512]&m[1538]&m[1539]&m[1541]&m[1542]))&UnbiasedRNG[540])|((m[1512]&~m[1538]&~m[1539]&m[1541]&~m[1542])|(~m[1512]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1512]&~m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1512]&m[1538]&~m[1539]&~m[1541]&m[1542])|(m[1512]&~m[1538]&m[1539]&~m[1541]&m[1542])|(~m[1512]&~m[1538]&~m[1539]&m[1541]&m[1542])|(m[1512]&~m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1512]&m[1538]&~m[1539]&m[1541]&m[1542])|(m[1512]&m[1538]&~m[1539]&m[1541]&m[1542])|(~m[1512]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1512]&~m[1538]&m[1539]&m[1541]&m[1542])|(m[1512]&m[1538]&m[1539]&m[1541]&m[1542]));
    m[1545] = (((m[1517]&~m[1543]&~m[1544]&~m[1546]&~m[1547])|(~m[1517]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1517]&m[1543]&~m[1544]&m[1546]&~m[1547])|(m[1517]&~m[1543]&m[1544]&m[1546]&~m[1547])|(~m[1517]&m[1543]&~m[1544]&~m[1546]&m[1547])|(~m[1517]&~m[1543]&m[1544]&~m[1546]&m[1547])|(m[1517]&m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1517]&m[1543]&m[1544]&m[1546]&m[1547]))&UnbiasedRNG[541])|((m[1517]&~m[1543]&~m[1544]&m[1546]&~m[1547])|(~m[1517]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1517]&~m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1517]&m[1543]&~m[1544]&~m[1546]&m[1547])|(m[1517]&~m[1543]&m[1544]&~m[1546]&m[1547])|(~m[1517]&~m[1543]&~m[1544]&m[1546]&m[1547])|(m[1517]&~m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1517]&m[1543]&~m[1544]&m[1546]&m[1547])|(m[1517]&m[1543]&~m[1544]&m[1546]&m[1547])|(~m[1517]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1517]&~m[1543]&m[1544]&m[1546]&m[1547])|(m[1517]&m[1543]&m[1544]&m[1546]&m[1547]));
    m[1550] = (((m[1522]&~m[1548]&~m[1549]&~m[1551]&~m[1552])|(~m[1522]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1522]&m[1548]&~m[1549]&m[1551]&~m[1552])|(m[1522]&~m[1548]&m[1549]&m[1551]&~m[1552])|(~m[1522]&m[1548]&~m[1549]&~m[1551]&m[1552])|(~m[1522]&~m[1548]&m[1549]&~m[1551]&m[1552])|(m[1522]&m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1522]&m[1548]&m[1549]&m[1551]&m[1552]))&UnbiasedRNG[542])|((m[1522]&~m[1548]&~m[1549]&m[1551]&~m[1552])|(~m[1522]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1522]&~m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1522]&m[1548]&~m[1549]&~m[1551]&m[1552])|(m[1522]&~m[1548]&m[1549]&~m[1551]&m[1552])|(~m[1522]&~m[1548]&~m[1549]&m[1551]&m[1552])|(m[1522]&~m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1522]&m[1548]&~m[1549]&m[1551]&m[1552])|(m[1522]&m[1548]&~m[1549]&m[1551]&m[1552])|(~m[1522]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1522]&~m[1548]&m[1549]&m[1551]&m[1552])|(m[1522]&m[1548]&m[1549]&m[1551]&m[1552]));
    m[1555] = (((m[1527]&~m[1553]&~m[1554]&~m[1556]&~m[1557])|(~m[1527]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1527]&m[1553]&~m[1554]&m[1556]&~m[1557])|(m[1527]&~m[1553]&m[1554]&m[1556]&~m[1557])|(~m[1527]&m[1553]&~m[1554]&~m[1556]&m[1557])|(~m[1527]&~m[1553]&m[1554]&~m[1556]&m[1557])|(m[1527]&m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1527]&m[1553]&m[1554]&m[1556]&m[1557]))&UnbiasedRNG[543])|((m[1527]&~m[1553]&~m[1554]&m[1556]&~m[1557])|(~m[1527]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1527]&~m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1527]&m[1553]&~m[1554]&~m[1556]&m[1557])|(m[1527]&~m[1553]&m[1554]&~m[1556]&m[1557])|(~m[1527]&~m[1553]&~m[1554]&m[1556]&m[1557])|(m[1527]&~m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1527]&m[1553]&~m[1554]&m[1556]&m[1557])|(m[1527]&m[1553]&~m[1554]&m[1556]&m[1557])|(~m[1527]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1527]&~m[1553]&m[1554]&m[1556]&m[1557])|(m[1527]&m[1553]&m[1554]&m[1556]&m[1557]));
    m[1560] = (((m[1532]&~m[1558]&~m[1559]&~m[1561]&~m[1562])|(~m[1532]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1532]&m[1558]&~m[1559]&m[1561]&~m[1562])|(m[1532]&~m[1558]&m[1559]&m[1561]&~m[1562])|(~m[1532]&m[1558]&~m[1559]&~m[1561]&m[1562])|(~m[1532]&~m[1558]&m[1559]&~m[1561]&m[1562])|(m[1532]&m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1532]&m[1558]&m[1559]&m[1561]&m[1562]))&UnbiasedRNG[544])|((m[1532]&~m[1558]&~m[1559]&m[1561]&~m[1562])|(~m[1532]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1532]&~m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1532]&m[1558]&~m[1559]&~m[1561]&m[1562])|(m[1532]&~m[1558]&m[1559]&~m[1561]&m[1562])|(~m[1532]&~m[1558]&~m[1559]&m[1561]&m[1562])|(m[1532]&~m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1532]&m[1558]&~m[1559]&m[1561]&m[1562])|(m[1532]&m[1558]&~m[1559]&m[1561]&m[1562])|(~m[1532]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1532]&~m[1558]&m[1559]&m[1561]&m[1562])|(m[1532]&m[1558]&m[1559]&m[1561]&m[1562]));
    m[1565] = (((m[1542]&~m[1563]&~m[1564]&~m[1566]&~m[1567])|(~m[1542]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1542]&m[1563]&~m[1564]&m[1566]&~m[1567])|(m[1542]&~m[1563]&m[1564]&m[1566]&~m[1567])|(~m[1542]&m[1563]&~m[1564]&~m[1566]&m[1567])|(~m[1542]&~m[1563]&m[1564]&~m[1566]&m[1567])|(m[1542]&m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1542]&m[1563]&m[1564]&m[1566]&m[1567]))&UnbiasedRNG[545])|((m[1542]&~m[1563]&~m[1564]&m[1566]&~m[1567])|(~m[1542]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1542]&~m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1542]&m[1563]&~m[1564]&~m[1566]&m[1567])|(m[1542]&~m[1563]&m[1564]&~m[1566]&m[1567])|(~m[1542]&~m[1563]&~m[1564]&m[1566]&m[1567])|(m[1542]&~m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1542]&m[1563]&~m[1564]&m[1566]&m[1567])|(m[1542]&m[1563]&~m[1564]&m[1566]&m[1567])|(~m[1542]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1542]&~m[1563]&m[1564]&m[1566]&m[1567])|(m[1542]&m[1563]&m[1564]&m[1566]&m[1567]));
    m[1570] = (((m[1547]&~m[1568]&~m[1569]&~m[1571]&~m[1572])|(~m[1547]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1547]&m[1568]&~m[1569]&m[1571]&~m[1572])|(m[1547]&~m[1568]&m[1569]&m[1571]&~m[1572])|(~m[1547]&m[1568]&~m[1569]&~m[1571]&m[1572])|(~m[1547]&~m[1568]&m[1569]&~m[1571]&m[1572])|(m[1547]&m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1547]&m[1568]&m[1569]&m[1571]&m[1572]))&UnbiasedRNG[546])|((m[1547]&~m[1568]&~m[1569]&m[1571]&~m[1572])|(~m[1547]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1547]&~m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1547]&m[1568]&~m[1569]&~m[1571]&m[1572])|(m[1547]&~m[1568]&m[1569]&~m[1571]&m[1572])|(~m[1547]&~m[1568]&~m[1569]&m[1571]&m[1572])|(m[1547]&~m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1547]&m[1568]&~m[1569]&m[1571]&m[1572])|(m[1547]&m[1568]&~m[1569]&m[1571]&m[1572])|(~m[1547]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1547]&~m[1568]&m[1569]&m[1571]&m[1572])|(m[1547]&m[1568]&m[1569]&m[1571]&m[1572]));
    m[1575] = (((m[1552]&~m[1573]&~m[1574]&~m[1576]&~m[1577])|(~m[1552]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1552]&m[1573]&~m[1574]&m[1576]&~m[1577])|(m[1552]&~m[1573]&m[1574]&m[1576]&~m[1577])|(~m[1552]&m[1573]&~m[1574]&~m[1576]&m[1577])|(~m[1552]&~m[1573]&m[1574]&~m[1576]&m[1577])|(m[1552]&m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1552]&m[1573]&m[1574]&m[1576]&m[1577]))&UnbiasedRNG[547])|((m[1552]&~m[1573]&~m[1574]&m[1576]&~m[1577])|(~m[1552]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1552]&~m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1552]&m[1573]&~m[1574]&~m[1576]&m[1577])|(m[1552]&~m[1573]&m[1574]&~m[1576]&m[1577])|(~m[1552]&~m[1573]&~m[1574]&m[1576]&m[1577])|(m[1552]&~m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1552]&m[1573]&~m[1574]&m[1576]&m[1577])|(m[1552]&m[1573]&~m[1574]&m[1576]&m[1577])|(~m[1552]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1552]&~m[1573]&m[1574]&m[1576]&m[1577])|(m[1552]&m[1573]&m[1574]&m[1576]&m[1577]));
    m[1580] = (((m[1557]&~m[1578]&~m[1579]&~m[1581]&~m[1582])|(~m[1557]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1557]&m[1578]&~m[1579]&m[1581]&~m[1582])|(m[1557]&~m[1578]&m[1579]&m[1581]&~m[1582])|(~m[1557]&m[1578]&~m[1579]&~m[1581]&m[1582])|(~m[1557]&~m[1578]&m[1579]&~m[1581]&m[1582])|(m[1557]&m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1557]&m[1578]&m[1579]&m[1581]&m[1582]))&UnbiasedRNG[548])|((m[1557]&~m[1578]&~m[1579]&m[1581]&~m[1582])|(~m[1557]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1557]&~m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1557]&m[1578]&~m[1579]&~m[1581]&m[1582])|(m[1557]&~m[1578]&m[1579]&~m[1581]&m[1582])|(~m[1557]&~m[1578]&~m[1579]&m[1581]&m[1582])|(m[1557]&~m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1557]&m[1578]&~m[1579]&m[1581]&m[1582])|(m[1557]&m[1578]&~m[1579]&m[1581]&m[1582])|(~m[1557]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1557]&~m[1578]&m[1579]&m[1581]&m[1582])|(m[1557]&m[1578]&m[1579]&m[1581]&m[1582]));
    m[1585] = (((m[1562]&~m[1583]&~m[1584]&~m[1586]&~m[1587])|(~m[1562]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1562]&m[1583]&~m[1584]&m[1586]&~m[1587])|(m[1562]&~m[1583]&m[1584]&m[1586]&~m[1587])|(~m[1562]&m[1583]&~m[1584]&~m[1586]&m[1587])|(~m[1562]&~m[1583]&m[1584]&~m[1586]&m[1587])|(m[1562]&m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1562]&m[1583]&m[1584]&m[1586]&m[1587]))&UnbiasedRNG[549])|((m[1562]&~m[1583]&~m[1584]&m[1586]&~m[1587])|(~m[1562]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1562]&~m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1562]&m[1583]&~m[1584]&~m[1586]&m[1587])|(m[1562]&~m[1583]&m[1584]&~m[1586]&m[1587])|(~m[1562]&~m[1583]&~m[1584]&m[1586]&m[1587])|(m[1562]&~m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1562]&m[1583]&~m[1584]&m[1586]&m[1587])|(m[1562]&m[1583]&~m[1584]&m[1586]&m[1587])|(~m[1562]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1562]&~m[1583]&m[1584]&m[1586]&m[1587])|(m[1562]&m[1583]&m[1584]&m[1586]&m[1587]));
    m[1590] = (((m[1572]&~m[1588]&~m[1589]&~m[1591]&~m[1592])|(~m[1572]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1572]&m[1588]&~m[1589]&m[1591]&~m[1592])|(m[1572]&~m[1588]&m[1589]&m[1591]&~m[1592])|(~m[1572]&m[1588]&~m[1589]&~m[1591]&m[1592])|(~m[1572]&~m[1588]&m[1589]&~m[1591]&m[1592])|(m[1572]&m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1572]&m[1588]&m[1589]&m[1591]&m[1592]))&UnbiasedRNG[550])|((m[1572]&~m[1588]&~m[1589]&m[1591]&~m[1592])|(~m[1572]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1572]&~m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1572]&m[1588]&~m[1589]&~m[1591]&m[1592])|(m[1572]&~m[1588]&m[1589]&~m[1591]&m[1592])|(~m[1572]&~m[1588]&~m[1589]&m[1591]&m[1592])|(m[1572]&~m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1572]&m[1588]&~m[1589]&m[1591]&m[1592])|(m[1572]&m[1588]&~m[1589]&m[1591]&m[1592])|(~m[1572]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1572]&~m[1588]&m[1589]&m[1591]&m[1592])|(m[1572]&m[1588]&m[1589]&m[1591]&m[1592]));
    m[1595] = (((m[1577]&~m[1593]&~m[1594]&~m[1596]&~m[1597])|(~m[1577]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1577]&m[1593]&~m[1594]&m[1596]&~m[1597])|(m[1577]&~m[1593]&m[1594]&m[1596]&~m[1597])|(~m[1577]&m[1593]&~m[1594]&~m[1596]&m[1597])|(~m[1577]&~m[1593]&m[1594]&~m[1596]&m[1597])|(m[1577]&m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1577]&m[1593]&m[1594]&m[1596]&m[1597]))&UnbiasedRNG[551])|((m[1577]&~m[1593]&~m[1594]&m[1596]&~m[1597])|(~m[1577]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1577]&~m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1577]&m[1593]&~m[1594]&~m[1596]&m[1597])|(m[1577]&~m[1593]&m[1594]&~m[1596]&m[1597])|(~m[1577]&~m[1593]&~m[1594]&m[1596]&m[1597])|(m[1577]&~m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1577]&m[1593]&~m[1594]&m[1596]&m[1597])|(m[1577]&m[1593]&~m[1594]&m[1596]&m[1597])|(~m[1577]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1577]&~m[1593]&m[1594]&m[1596]&m[1597])|(m[1577]&m[1593]&m[1594]&m[1596]&m[1597]));
    m[1600] = (((m[1582]&~m[1598]&~m[1599]&~m[1601]&~m[1602])|(~m[1582]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1582]&m[1598]&~m[1599]&m[1601]&~m[1602])|(m[1582]&~m[1598]&m[1599]&m[1601]&~m[1602])|(~m[1582]&m[1598]&~m[1599]&~m[1601]&m[1602])|(~m[1582]&~m[1598]&m[1599]&~m[1601]&m[1602])|(m[1582]&m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1582]&m[1598]&m[1599]&m[1601]&m[1602]))&UnbiasedRNG[552])|((m[1582]&~m[1598]&~m[1599]&m[1601]&~m[1602])|(~m[1582]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1582]&~m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1582]&m[1598]&~m[1599]&~m[1601]&m[1602])|(m[1582]&~m[1598]&m[1599]&~m[1601]&m[1602])|(~m[1582]&~m[1598]&~m[1599]&m[1601]&m[1602])|(m[1582]&~m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1582]&m[1598]&~m[1599]&m[1601]&m[1602])|(m[1582]&m[1598]&~m[1599]&m[1601]&m[1602])|(~m[1582]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1582]&~m[1598]&m[1599]&m[1601]&m[1602])|(m[1582]&m[1598]&m[1599]&m[1601]&m[1602]));
    m[1605] = (((m[1587]&~m[1603]&~m[1604]&~m[1606]&~m[1607])|(~m[1587]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1587]&m[1603]&~m[1604]&m[1606]&~m[1607])|(m[1587]&~m[1603]&m[1604]&m[1606]&~m[1607])|(~m[1587]&m[1603]&~m[1604]&~m[1606]&m[1607])|(~m[1587]&~m[1603]&m[1604]&~m[1606]&m[1607])|(m[1587]&m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1587]&m[1603]&m[1604]&m[1606]&m[1607]))&UnbiasedRNG[553])|((m[1587]&~m[1603]&~m[1604]&m[1606]&~m[1607])|(~m[1587]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1587]&~m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1587]&m[1603]&~m[1604]&~m[1606]&m[1607])|(m[1587]&~m[1603]&m[1604]&~m[1606]&m[1607])|(~m[1587]&~m[1603]&~m[1604]&m[1606]&m[1607])|(m[1587]&~m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1587]&m[1603]&~m[1604]&m[1606]&m[1607])|(m[1587]&m[1603]&~m[1604]&m[1606]&m[1607])|(~m[1587]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1587]&~m[1603]&m[1604]&m[1606]&m[1607])|(m[1587]&m[1603]&m[1604]&m[1606]&m[1607]));
    m[1610] = (((m[1597]&~m[1608]&~m[1609]&~m[1611]&~m[1612])|(~m[1597]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1597]&m[1608]&~m[1609]&m[1611]&~m[1612])|(m[1597]&~m[1608]&m[1609]&m[1611]&~m[1612])|(~m[1597]&m[1608]&~m[1609]&~m[1611]&m[1612])|(~m[1597]&~m[1608]&m[1609]&~m[1611]&m[1612])|(m[1597]&m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1597]&m[1608]&m[1609]&m[1611]&m[1612]))&UnbiasedRNG[554])|((m[1597]&~m[1608]&~m[1609]&m[1611]&~m[1612])|(~m[1597]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1597]&~m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1597]&m[1608]&~m[1609]&~m[1611]&m[1612])|(m[1597]&~m[1608]&m[1609]&~m[1611]&m[1612])|(~m[1597]&~m[1608]&~m[1609]&m[1611]&m[1612])|(m[1597]&~m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1597]&m[1608]&~m[1609]&m[1611]&m[1612])|(m[1597]&m[1608]&~m[1609]&m[1611]&m[1612])|(~m[1597]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1597]&~m[1608]&m[1609]&m[1611]&m[1612])|(m[1597]&m[1608]&m[1609]&m[1611]&m[1612]));
    m[1615] = (((m[1602]&~m[1613]&~m[1614]&~m[1616]&~m[1617])|(~m[1602]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1602]&m[1613]&~m[1614]&m[1616]&~m[1617])|(m[1602]&~m[1613]&m[1614]&m[1616]&~m[1617])|(~m[1602]&m[1613]&~m[1614]&~m[1616]&m[1617])|(~m[1602]&~m[1613]&m[1614]&~m[1616]&m[1617])|(m[1602]&m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1602]&m[1613]&m[1614]&m[1616]&m[1617]))&UnbiasedRNG[555])|((m[1602]&~m[1613]&~m[1614]&m[1616]&~m[1617])|(~m[1602]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1602]&~m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1602]&m[1613]&~m[1614]&~m[1616]&m[1617])|(m[1602]&~m[1613]&m[1614]&~m[1616]&m[1617])|(~m[1602]&~m[1613]&~m[1614]&m[1616]&m[1617])|(m[1602]&~m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1602]&m[1613]&~m[1614]&m[1616]&m[1617])|(m[1602]&m[1613]&~m[1614]&m[1616]&m[1617])|(~m[1602]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1602]&~m[1613]&m[1614]&m[1616]&m[1617])|(m[1602]&m[1613]&m[1614]&m[1616]&m[1617]));
    m[1620] = (((m[1607]&~m[1618]&~m[1619]&~m[1621]&~m[1622])|(~m[1607]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1607]&m[1618]&~m[1619]&m[1621]&~m[1622])|(m[1607]&~m[1618]&m[1619]&m[1621]&~m[1622])|(~m[1607]&m[1618]&~m[1619]&~m[1621]&m[1622])|(~m[1607]&~m[1618]&m[1619]&~m[1621]&m[1622])|(m[1607]&m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1607]&m[1618]&m[1619]&m[1621]&m[1622]))&UnbiasedRNG[556])|((m[1607]&~m[1618]&~m[1619]&m[1621]&~m[1622])|(~m[1607]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1607]&~m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1607]&m[1618]&~m[1619]&~m[1621]&m[1622])|(m[1607]&~m[1618]&m[1619]&~m[1621]&m[1622])|(~m[1607]&~m[1618]&~m[1619]&m[1621]&m[1622])|(m[1607]&~m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1607]&m[1618]&~m[1619]&m[1621]&m[1622])|(m[1607]&m[1618]&~m[1619]&m[1621]&m[1622])|(~m[1607]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1607]&~m[1618]&m[1619]&m[1621]&m[1622])|(m[1607]&m[1618]&m[1619]&m[1621]&m[1622]));
    m[1625] = (((m[1617]&~m[1623]&~m[1624]&~m[1626]&~m[1627])|(~m[1617]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1617]&m[1623]&~m[1624]&m[1626]&~m[1627])|(m[1617]&~m[1623]&m[1624]&m[1626]&~m[1627])|(~m[1617]&m[1623]&~m[1624]&~m[1626]&m[1627])|(~m[1617]&~m[1623]&m[1624]&~m[1626]&m[1627])|(m[1617]&m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1617]&m[1623]&m[1624]&m[1626]&m[1627]))&UnbiasedRNG[557])|((m[1617]&~m[1623]&~m[1624]&m[1626]&~m[1627])|(~m[1617]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1617]&~m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1617]&m[1623]&~m[1624]&~m[1626]&m[1627])|(m[1617]&~m[1623]&m[1624]&~m[1626]&m[1627])|(~m[1617]&~m[1623]&~m[1624]&m[1626]&m[1627])|(m[1617]&~m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1617]&m[1623]&~m[1624]&m[1626]&m[1627])|(m[1617]&m[1623]&~m[1624]&m[1626]&m[1627])|(~m[1617]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1617]&~m[1623]&m[1624]&m[1626]&m[1627])|(m[1617]&m[1623]&m[1624]&m[1626]&m[1627]));
    m[1630] = (((m[1622]&~m[1628]&~m[1629]&~m[1631]&~m[1632])|(~m[1622]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1622]&m[1628]&~m[1629]&m[1631]&~m[1632])|(m[1622]&~m[1628]&m[1629]&m[1631]&~m[1632])|(~m[1622]&m[1628]&~m[1629]&~m[1631]&m[1632])|(~m[1622]&~m[1628]&m[1629]&~m[1631]&m[1632])|(m[1622]&m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1622]&m[1628]&m[1629]&m[1631]&m[1632]))&UnbiasedRNG[558])|((m[1622]&~m[1628]&~m[1629]&m[1631]&~m[1632])|(~m[1622]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1622]&~m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1622]&m[1628]&~m[1629]&~m[1631]&m[1632])|(m[1622]&~m[1628]&m[1629]&~m[1631]&m[1632])|(~m[1622]&~m[1628]&~m[1629]&m[1631]&m[1632])|(m[1622]&~m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1622]&m[1628]&~m[1629]&m[1631]&m[1632])|(m[1622]&m[1628]&~m[1629]&m[1631]&m[1632])|(~m[1622]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1622]&~m[1628]&m[1629]&m[1631]&m[1632])|(m[1622]&m[1628]&m[1629]&m[1631]&m[1632]));
    m[1635] = (((m[1632]&~m[1633]&~m[1634]&~m[1636]&~m[1637])|(~m[1632]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1632]&m[1633]&~m[1634]&m[1636]&~m[1637])|(m[1632]&~m[1633]&m[1634]&m[1636]&~m[1637])|(~m[1632]&m[1633]&~m[1634]&~m[1636]&m[1637])|(~m[1632]&~m[1633]&m[1634]&~m[1636]&m[1637])|(m[1632]&m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1632]&m[1633]&m[1634]&m[1636]&m[1637]))&UnbiasedRNG[559])|((m[1632]&~m[1633]&~m[1634]&m[1636]&~m[1637])|(~m[1632]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1632]&~m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1632]&m[1633]&~m[1634]&~m[1636]&m[1637])|(m[1632]&~m[1633]&m[1634]&~m[1636]&m[1637])|(~m[1632]&~m[1633]&~m[1634]&m[1636]&m[1637])|(m[1632]&~m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1632]&m[1633]&~m[1634]&m[1636]&m[1637])|(m[1632]&m[1633]&~m[1634]&m[1636]&m[1637])|(~m[1632]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1632]&~m[1633]&m[1634]&m[1636]&m[1637])|(m[1632]&m[1633]&m[1634]&m[1636]&m[1637]));
end

always @(posedge color3_clk) begin
    m[736] = (((m[733]&~m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&m[734]&~m[735]&~m[737]&~m[738])|(~m[733]&~m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&m[737]&~m[738])|(~m[733]&~m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&m[737]&m[738])|(m[733]&~m[734]&m[735]&m[737]&m[738])|(~m[733]&m[734]&m[735]&m[737]&m[738]))&UnbiasedRNG[560])|((m[733]&m[734]&~m[735]&~m[737]&~m[738])|(m[733]&~m[734]&m[735]&~m[737]&~m[738])|(~m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&m[734]&m[735]&~m[737]&~m[738])|(m[733]&~m[734]&~m[735]&~m[737]&m[738])|(~m[733]&m[734]&~m[735]&~m[737]&m[738])|(m[733]&m[734]&~m[735]&~m[737]&m[738])|(~m[733]&~m[734]&m[735]&~m[737]&m[738])|(m[733]&~m[734]&m[735]&~m[737]&m[738])|(~m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&~m[737]&m[738])|(m[733]&m[734]&m[735]&m[737]&m[738]));
    m[746] = (((m[743]&~m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&m[744]&~m[745]&~m[747]&~m[748])|(~m[743]&~m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&m[747]&~m[748])|(~m[743]&~m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&m[747]&m[748])|(m[743]&~m[744]&m[745]&m[747]&m[748])|(~m[743]&m[744]&m[745]&m[747]&m[748]))&UnbiasedRNG[561])|((m[743]&m[744]&~m[745]&~m[747]&~m[748])|(m[743]&~m[744]&m[745]&~m[747]&~m[748])|(~m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&m[744]&m[745]&~m[747]&~m[748])|(m[743]&~m[744]&~m[745]&~m[747]&m[748])|(~m[743]&m[744]&~m[745]&~m[747]&m[748])|(m[743]&m[744]&~m[745]&~m[747]&m[748])|(~m[743]&~m[744]&m[745]&~m[747]&m[748])|(m[743]&~m[744]&m[745]&~m[747]&m[748])|(~m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&~m[747]&m[748])|(m[743]&m[744]&m[745]&m[747]&m[748]));
    m[751] = (((m[748]&~m[749]&~m[750]&~m[752]&~m[753])|(~m[748]&m[749]&~m[750]&~m[752]&~m[753])|(~m[748]&~m[749]&m[750]&~m[752]&~m[753])|(m[748]&m[749]&m[750]&m[752]&~m[753])|(~m[748]&~m[749]&~m[750]&~m[752]&m[753])|(m[748]&m[749]&~m[750]&m[752]&m[753])|(m[748]&~m[749]&m[750]&m[752]&m[753])|(~m[748]&m[749]&m[750]&m[752]&m[753]))&UnbiasedRNG[562])|((m[748]&m[749]&~m[750]&~m[752]&~m[753])|(m[748]&~m[749]&m[750]&~m[752]&~m[753])|(~m[748]&m[749]&m[750]&~m[752]&~m[753])|(m[748]&m[749]&m[750]&~m[752]&~m[753])|(m[748]&~m[749]&~m[750]&~m[752]&m[753])|(~m[748]&m[749]&~m[750]&~m[752]&m[753])|(m[748]&m[749]&~m[750]&~m[752]&m[753])|(~m[748]&~m[749]&m[750]&~m[752]&m[753])|(m[748]&~m[749]&m[750]&~m[752]&m[753])|(~m[748]&m[749]&m[750]&~m[752]&m[753])|(m[748]&m[749]&m[750]&~m[752]&m[753])|(m[748]&m[749]&m[750]&m[752]&m[753]));
    m[761] = (((m[758]&~m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&m[759]&~m[760]&~m[762]&~m[763])|(~m[758]&~m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&m[762]&~m[763])|(~m[758]&~m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&m[762]&m[763])|(m[758]&~m[759]&m[760]&m[762]&m[763])|(~m[758]&m[759]&m[760]&m[762]&m[763]))&UnbiasedRNG[563])|((m[758]&m[759]&~m[760]&~m[762]&~m[763])|(m[758]&~m[759]&m[760]&~m[762]&~m[763])|(~m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&m[759]&m[760]&~m[762]&~m[763])|(m[758]&~m[759]&~m[760]&~m[762]&m[763])|(~m[758]&m[759]&~m[760]&~m[762]&m[763])|(m[758]&m[759]&~m[760]&~m[762]&m[763])|(~m[758]&~m[759]&m[760]&~m[762]&m[763])|(m[758]&~m[759]&m[760]&~m[762]&m[763])|(~m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&~m[762]&m[763])|(m[758]&m[759]&m[760]&m[762]&m[763]));
    m[766] = (((m[763]&~m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&m[764]&~m[765]&~m[767]&~m[768])|(~m[763]&~m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&m[767]&~m[768])|(~m[763]&~m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&m[767]&m[768])|(m[763]&~m[764]&m[765]&m[767]&m[768])|(~m[763]&m[764]&m[765]&m[767]&m[768]))&UnbiasedRNG[564])|((m[763]&m[764]&~m[765]&~m[767]&~m[768])|(m[763]&~m[764]&m[765]&~m[767]&~m[768])|(~m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&m[764]&m[765]&~m[767]&~m[768])|(m[763]&~m[764]&~m[765]&~m[767]&m[768])|(~m[763]&m[764]&~m[765]&~m[767]&m[768])|(m[763]&m[764]&~m[765]&~m[767]&m[768])|(~m[763]&~m[764]&m[765]&~m[767]&m[768])|(m[763]&~m[764]&m[765]&~m[767]&m[768])|(~m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&~m[767]&m[768])|(m[763]&m[764]&m[765]&m[767]&m[768]));
    m[771] = (((m[768]&~m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&m[769]&~m[770]&~m[772]&~m[773])|(~m[768]&~m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&m[772]&~m[773])|(~m[768]&~m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&m[772]&m[773])|(m[768]&~m[769]&m[770]&m[772]&m[773])|(~m[768]&m[769]&m[770]&m[772]&m[773]))&UnbiasedRNG[565])|((m[768]&m[769]&~m[770]&~m[772]&~m[773])|(m[768]&~m[769]&m[770]&~m[772]&~m[773])|(~m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&m[769]&m[770]&~m[772]&~m[773])|(m[768]&~m[769]&~m[770]&~m[772]&m[773])|(~m[768]&m[769]&~m[770]&~m[772]&m[773])|(m[768]&m[769]&~m[770]&~m[772]&m[773])|(~m[768]&~m[769]&m[770]&~m[772]&m[773])|(m[768]&~m[769]&m[770]&~m[772]&m[773])|(~m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&~m[772]&m[773])|(m[768]&m[769]&m[770]&m[772]&m[773]));
    m[781] = (((m[778]&~m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&m[779]&~m[780]&~m[782]&~m[783])|(~m[778]&~m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&m[782]&~m[783])|(~m[778]&~m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&m[782]&m[783])|(m[778]&~m[779]&m[780]&m[782]&m[783])|(~m[778]&m[779]&m[780]&m[782]&m[783]))&UnbiasedRNG[566])|((m[778]&m[779]&~m[780]&~m[782]&~m[783])|(m[778]&~m[779]&m[780]&~m[782]&~m[783])|(~m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&m[779]&m[780]&~m[782]&~m[783])|(m[778]&~m[779]&~m[780]&~m[782]&m[783])|(~m[778]&m[779]&~m[780]&~m[782]&m[783])|(m[778]&m[779]&~m[780]&~m[782]&m[783])|(~m[778]&~m[779]&m[780]&~m[782]&m[783])|(m[778]&~m[779]&m[780]&~m[782]&m[783])|(~m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&~m[782]&m[783])|(m[778]&m[779]&m[780]&m[782]&m[783]));
    m[786] = (((m[783]&~m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&m[784]&~m[785]&~m[787]&~m[788])|(~m[783]&~m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&m[787]&~m[788])|(~m[783]&~m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&m[787]&m[788])|(m[783]&~m[784]&m[785]&m[787]&m[788])|(~m[783]&m[784]&m[785]&m[787]&m[788]))&UnbiasedRNG[567])|((m[783]&m[784]&~m[785]&~m[787]&~m[788])|(m[783]&~m[784]&m[785]&~m[787]&~m[788])|(~m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&m[784]&m[785]&~m[787]&~m[788])|(m[783]&~m[784]&~m[785]&~m[787]&m[788])|(~m[783]&m[784]&~m[785]&~m[787]&m[788])|(m[783]&m[784]&~m[785]&~m[787]&m[788])|(~m[783]&~m[784]&m[785]&~m[787]&m[788])|(m[783]&~m[784]&m[785]&~m[787]&m[788])|(~m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&~m[787]&m[788])|(m[783]&m[784]&m[785]&m[787]&m[788]));
    m[791] = (((m[788]&~m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&m[789]&~m[790]&~m[792]&~m[793])|(~m[788]&~m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&m[792]&~m[793])|(~m[788]&~m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&m[792]&m[793])|(m[788]&~m[789]&m[790]&m[792]&m[793])|(~m[788]&m[789]&m[790]&m[792]&m[793]))&UnbiasedRNG[568])|((m[788]&m[789]&~m[790]&~m[792]&~m[793])|(m[788]&~m[789]&m[790]&~m[792]&~m[793])|(~m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&m[789]&m[790]&~m[792]&~m[793])|(m[788]&~m[789]&~m[790]&~m[792]&m[793])|(~m[788]&m[789]&~m[790]&~m[792]&m[793])|(m[788]&m[789]&~m[790]&~m[792]&m[793])|(~m[788]&~m[789]&m[790]&~m[792]&m[793])|(m[788]&~m[789]&m[790]&~m[792]&m[793])|(~m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&~m[792]&m[793])|(m[788]&m[789]&m[790]&m[792]&m[793]));
    m[796] = (((m[793]&~m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&m[794]&~m[795]&~m[797]&~m[798])|(~m[793]&~m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&m[797]&~m[798])|(~m[793]&~m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&m[797]&m[798])|(m[793]&~m[794]&m[795]&m[797]&m[798])|(~m[793]&m[794]&m[795]&m[797]&m[798]))&UnbiasedRNG[569])|((m[793]&m[794]&~m[795]&~m[797]&~m[798])|(m[793]&~m[794]&m[795]&~m[797]&~m[798])|(~m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&m[794]&m[795]&~m[797]&~m[798])|(m[793]&~m[794]&~m[795]&~m[797]&m[798])|(~m[793]&m[794]&~m[795]&~m[797]&m[798])|(m[793]&m[794]&~m[795]&~m[797]&m[798])|(~m[793]&~m[794]&m[795]&~m[797]&m[798])|(m[793]&~m[794]&m[795]&~m[797]&m[798])|(~m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&~m[797]&m[798])|(m[793]&m[794]&m[795]&m[797]&m[798]));
    m[806] = (((m[803]&~m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&m[804]&~m[805]&~m[807]&~m[808])|(~m[803]&~m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&m[807]&~m[808])|(~m[803]&~m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&m[807]&m[808])|(m[803]&~m[804]&m[805]&m[807]&m[808])|(~m[803]&m[804]&m[805]&m[807]&m[808]))&UnbiasedRNG[570])|((m[803]&m[804]&~m[805]&~m[807]&~m[808])|(m[803]&~m[804]&m[805]&~m[807]&~m[808])|(~m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&m[804]&m[805]&~m[807]&~m[808])|(m[803]&~m[804]&~m[805]&~m[807]&m[808])|(~m[803]&m[804]&~m[805]&~m[807]&m[808])|(m[803]&m[804]&~m[805]&~m[807]&m[808])|(~m[803]&~m[804]&m[805]&~m[807]&m[808])|(m[803]&~m[804]&m[805]&~m[807]&m[808])|(~m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&~m[807]&m[808])|(m[803]&m[804]&m[805]&m[807]&m[808]));
    m[811] = (((m[808]&~m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&m[809]&~m[810]&~m[812]&~m[813])|(~m[808]&~m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&m[812]&~m[813])|(~m[808]&~m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&m[812]&m[813])|(m[808]&~m[809]&m[810]&m[812]&m[813])|(~m[808]&m[809]&m[810]&m[812]&m[813]))&UnbiasedRNG[571])|((m[808]&m[809]&~m[810]&~m[812]&~m[813])|(m[808]&~m[809]&m[810]&~m[812]&~m[813])|(~m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&m[809]&m[810]&~m[812]&~m[813])|(m[808]&~m[809]&~m[810]&~m[812]&m[813])|(~m[808]&m[809]&~m[810]&~m[812]&m[813])|(m[808]&m[809]&~m[810]&~m[812]&m[813])|(~m[808]&~m[809]&m[810]&~m[812]&m[813])|(m[808]&~m[809]&m[810]&~m[812]&m[813])|(~m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&~m[812]&m[813])|(m[808]&m[809]&m[810]&m[812]&m[813]));
    m[816] = (((m[813]&~m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&m[814]&~m[815]&~m[817]&~m[818])|(~m[813]&~m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&m[817]&~m[818])|(~m[813]&~m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&m[817]&m[818])|(m[813]&~m[814]&m[815]&m[817]&m[818])|(~m[813]&m[814]&m[815]&m[817]&m[818]))&UnbiasedRNG[572])|((m[813]&m[814]&~m[815]&~m[817]&~m[818])|(m[813]&~m[814]&m[815]&~m[817]&~m[818])|(~m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&m[814]&m[815]&~m[817]&~m[818])|(m[813]&~m[814]&~m[815]&~m[817]&m[818])|(~m[813]&m[814]&~m[815]&~m[817]&m[818])|(m[813]&m[814]&~m[815]&~m[817]&m[818])|(~m[813]&~m[814]&m[815]&~m[817]&m[818])|(m[813]&~m[814]&m[815]&~m[817]&m[818])|(~m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&~m[817]&m[818])|(m[813]&m[814]&m[815]&m[817]&m[818]));
    m[821] = (((m[818]&~m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&m[819]&~m[820]&~m[822]&~m[823])|(~m[818]&~m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&m[822]&~m[823])|(~m[818]&~m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&m[822]&m[823])|(m[818]&~m[819]&m[820]&m[822]&m[823])|(~m[818]&m[819]&m[820]&m[822]&m[823]))&UnbiasedRNG[573])|((m[818]&m[819]&~m[820]&~m[822]&~m[823])|(m[818]&~m[819]&m[820]&~m[822]&~m[823])|(~m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&m[819]&m[820]&~m[822]&~m[823])|(m[818]&~m[819]&~m[820]&~m[822]&m[823])|(~m[818]&m[819]&~m[820]&~m[822]&m[823])|(m[818]&m[819]&~m[820]&~m[822]&m[823])|(~m[818]&~m[819]&m[820]&~m[822]&m[823])|(m[818]&~m[819]&m[820]&~m[822]&m[823])|(~m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&~m[822]&m[823])|(m[818]&m[819]&m[820]&m[822]&m[823]));
    m[826] = (((m[823]&~m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&m[824]&~m[825]&~m[827]&~m[828])|(~m[823]&~m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&m[827]&~m[828])|(~m[823]&~m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&m[827]&m[828])|(m[823]&~m[824]&m[825]&m[827]&m[828])|(~m[823]&m[824]&m[825]&m[827]&m[828]))&UnbiasedRNG[574])|((m[823]&m[824]&~m[825]&~m[827]&~m[828])|(m[823]&~m[824]&m[825]&~m[827]&~m[828])|(~m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&m[824]&m[825]&~m[827]&~m[828])|(m[823]&~m[824]&~m[825]&~m[827]&m[828])|(~m[823]&m[824]&~m[825]&~m[827]&m[828])|(m[823]&m[824]&~m[825]&~m[827]&m[828])|(~m[823]&~m[824]&m[825]&~m[827]&m[828])|(m[823]&~m[824]&m[825]&~m[827]&m[828])|(~m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&~m[827]&m[828])|(m[823]&m[824]&m[825]&m[827]&m[828]));
    m[836] = (((m[833]&~m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&m[834]&~m[835]&~m[837]&~m[838])|(~m[833]&~m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&m[837]&~m[838])|(~m[833]&~m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&m[837]&m[838])|(m[833]&~m[834]&m[835]&m[837]&m[838])|(~m[833]&m[834]&m[835]&m[837]&m[838]))&UnbiasedRNG[575])|((m[833]&m[834]&~m[835]&~m[837]&~m[838])|(m[833]&~m[834]&m[835]&~m[837]&~m[838])|(~m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&m[834]&m[835]&~m[837]&~m[838])|(m[833]&~m[834]&~m[835]&~m[837]&m[838])|(~m[833]&m[834]&~m[835]&~m[837]&m[838])|(m[833]&m[834]&~m[835]&~m[837]&m[838])|(~m[833]&~m[834]&m[835]&~m[837]&m[838])|(m[833]&~m[834]&m[835]&~m[837]&m[838])|(~m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&~m[837]&m[838])|(m[833]&m[834]&m[835]&m[837]&m[838]));
    m[841] = (((m[838]&~m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&m[839]&~m[840]&~m[842]&~m[843])|(~m[838]&~m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&m[842]&~m[843])|(~m[838]&~m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&m[842]&m[843])|(m[838]&~m[839]&m[840]&m[842]&m[843])|(~m[838]&m[839]&m[840]&m[842]&m[843]))&UnbiasedRNG[576])|((m[838]&m[839]&~m[840]&~m[842]&~m[843])|(m[838]&~m[839]&m[840]&~m[842]&~m[843])|(~m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&m[839]&m[840]&~m[842]&~m[843])|(m[838]&~m[839]&~m[840]&~m[842]&m[843])|(~m[838]&m[839]&~m[840]&~m[842]&m[843])|(m[838]&m[839]&~m[840]&~m[842]&m[843])|(~m[838]&~m[839]&m[840]&~m[842]&m[843])|(m[838]&~m[839]&m[840]&~m[842]&m[843])|(~m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&~m[842]&m[843])|(m[838]&m[839]&m[840]&m[842]&m[843]));
    m[846] = (((m[843]&~m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&m[844]&~m[845]&~m[847]&~m[848])|(~m[843]&~m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&m[847]&~m[848])|(~m[843]&~m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&m[847]&m[848])|(m[843]&~m[844]&m[845]&m[847]&m[848])|(~m[843]&m[844]&m[845]&m[847]&m[848]))&UnbiasedRNG[577])|((m[843]&m[844]&~m[845]&~m[847]&~m[848])|(m[843]&~m[844]&m[845]&~m[847]&~m[848])|(~m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&m[844]&m[845]&~m[847]&~m[848])|(m[843]&~m[844]&~m[845]&~m[847]&m[848])|(~m[843]&m[844]&~m[845]&~m[847]&m[848])|(m[843]&m[844]&~m[845]&~m[847]&m[848])|(~m[843]&~m[844]&m[845]&~m[847]&m[848])|(m[843]&~m[844]&m[845]&~m[847]&m[848])|(~m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&~m[847]&m[848])|(m[843]&m[844]&m[845]&m[847]&m[848]));
    m[851] = (((m[848]&~m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&m[849]&~m[850]&~m[852]&~m[853])|(~m[848]&~m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&m[852]&~m[853])|(~m[848]&~m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&m[852]&m[853])|(m[848]&~m[849]&m[850]&m[852]&m[853])|(~m[848]&m[849]&m[850]&m[852]&m[853]))&UnbiasedRNG[578])|((m[848]&m[849]&~m[850]&~m[852]&~m[853])|(m[848]&~m[849]&m[850]&~m[852]&~m[853])|(~m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&m[849]&m[850]&~m[852]&~m[853])|(m[848]&~m[849]&~m[850]&~m[852]&m[853])|(~m[848]&m[849]&~m[850]&~m[852]&m[853])|(m[848]&m[849]&~m[850]&~m[852]&m[853])|(~m[848]&~m[849]&m[850]&~m[852]&m[853])|(m[848]&~m[849]&m[850]&~m[852]&m[853])|(~m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&~m[852]&m[853])|(m[848]&m[849]&m[850]&m[852]&m[853]));
    m[856] = (((m[853]&~m[854]&~m[855]&~m[857]&~m[858])|(~m[853]&m[854]&~m[855]&~m[857]&~m[858])|(~m[853]&~m[854]&m[855]&~m[857]&~m[858])|(m[853]&m[854]&m[855]&m[857]&~m[858])|(~m[853]&~m[854]&~m[855]&~m[857]&m[858])|(m[853]&m[854]&~m[855]&m[857]&m[858])|(m[853]&~m[854]&m[855]&m[857]&m[858])|(~m[853]&m[854]&m[855]&m[857]&m[858]))&UnbiasedRNG[579])|((m[853]&m[854]&~m[855]&~m[857]&~m[858])|(m[853]&~m[854]&m[855]&~m[857]&~m[858])|(~m[853]&m[854]&m[855]&~m[857]&~m[858])|(m[853]&m[854]&m[855]&~m[857]&~m[858])|(m[853]&~m[854]&~m[855]&~m[857]&m[858])|(~m[853]&m[854]&~m[855]&~m[857]&m[858])|(m[853]&m[854]&~m[855]&~m[857]&m[858])|(~m[853]&~m[854]&m[855]&~m[857]&m[858])|(m[853]&~m[854]&m[855]&~m[857]&m[858])|(~m[853]&m[854]&m[855]&~m[857]&m[858])|(m[853]&m[854]&m[855]&~m[857]&m[858])|(m[853]&m[854]&m[855]&m[857]&m[858]));
    m[861] = (((m[858]&~m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&m[859]&~m[860]&~m[862]&~m[863])|(~m[858]&~m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&m[862]&~m[863])|(~m[858]&~m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&m[862]&m[863])|(m[858]&~m[859]&m[860]&m[862]&m[863])|(~m[858]&m[859]&m[860]&m[862]&m[863]))&UnbiasedRNG[580])|((m[858]&m[859]&~m[860]&~m[862]&~m[863])|(m[858]&~m[859]&m[860]&~m[862]&~m[863])|(~m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&m[859]&m[860]&~m[862]&~m[863])|(m[858]&~m[859]&~m[860]&~m[862]&m[863])|(~m[858]&m[859]&~m[860]&~m[862]&m[863])|(m[858]&m[859]&~m[860]&~m[862]&m[863])|(~m[858]&~m[859]&m[860]&~m[862]&m[863])|(m[858]&~m[859]&m[860]&~m[862]&m[863])|(~m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&~m[862]&m[863])|(m[858]&m[859]&m[860]&m[862]&m[863]));
    m[871] = (((m[868]&~m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&m[869]&~m[870]&~m[872]&~m[873])|(~m[868]&~m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&m[872]&~m[873])|(~m[868]&~m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&m[872]&m[873])|(m[868]&~m[869]&m[870]&m[872]&m[873])|(~m[868]&m[869]&m[870]&m[872]&m[873]))&UnbiasedRNG[581])|((m[868]&m[869]&~m[870]&~m[872]&~m[873])|(m[868]&~m[869]&m[870]&~m[872]&~m[873])|(~m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&m[869]&m[870]&~m[872]&~m[873])|(m[868]&~m[869]&~m[870]&~m[872]&m[873])|(~m[868]&m[869]&~m[870]&~m[872]&m[873])|(m[868]&m[869]&~m[870]&~m[872]&m[873])|(~m[868]&~m[869]&m[870]&~m[872]&m[873])|(m[868]&~m[869]&m[870]&~m[872]&m[873])|(~m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&~m[872]&m[873])|(m[868]&m[869]&m[870]&m[872]&m[873]));
    m[876] = (((m[873]&~m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&m[874]&~m[875]&~m[877]&~m[878])|(~m[873]&~m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&m[877]&~m[878])|(~m[873]&~m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&m[877]&m[878])|(m[873]&~m[874]&m[875]&m[877]&m[878])|(~m[873]&m[874]&m[875]&m[877]&m[878]))&UnbiasedRNG[582])|((m[873]&m[874]&~m[875]&~m[877]&~m[878])|(m[873]&~m[874]&m[875]&~m[877]&~m[878])|(~m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&m[874]&m[875]&~m[877]&~m[878])|(m[873]&~m[874]&~m[875]&~m[877]&m[878])|(~m[873]&m[874]&~m[875]&~m[877]&m[878])|(m[873]&m[874]&~m[875]&~m[877]&m[878])|(~m[873]&~m[874]&m[875]&~m[877]&m[878])|(m[873]&~m[874]&m[875]&~m[877]&m[878])|(~m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&~m[877]&m[878])|(m[873]&m[874]&m[875]&m[877]&m[878]));
    m[881] = (((m[878]&~m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&m[879]&~m[880]&~m[882]&~m[883])|(~m[878]&~m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&m[882]&~m[883])|(~m[878]&~m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&m[882]&m[883])|(m[878]&~m[879]&m[880]&m[882]&m[883])|(~m[878]&m[879]&m[880]&m[882]&m[883]))&UnbiasedRNG[583])|((m[878]&m[879]&~m[880]&~m[882]&~m[883])|(m[878]&~m[879]&m[880]&~m[882]&~m[883])|(~m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&m[879]&m[880]&~m[882]&~m[883])|(m[878]&~m[879]&~m[880]&~m[882]&m[883])|(~m[878]&m[879]&~m[880]&~m[882]&m[883])|(m[878]&m[879]&~m[880]&~m[882]&m[883])|(~m[878]&~m[879]&m[880]&~m[882]&m[883])|(m[878]&~m[879]&m[880]&~m[882]&m[883])|(~m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&~m[882]&m[883])|(m[878]&m[879]&m[880]&m[882]&m[883]));
    m[886] = (((m[883]&~m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&m[884]&~m[885]&~m[887]&~m[888])|(~m[883]&~m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&m[887]&~m[888])|(~m[883]&~m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&m[887]&m[888])|(m[883]&~m[884]&m[885]&m[887]&m[888])|(~m[883]&m[884]&m[885]&m[887]&m[888]))&UnbiasedRNG[584])|((m[883]&m[884]&~m[885]&~m[887]&~m[888])|(m[883]&~m[884]&m[885]&~m[887]&~m[888])|(~m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&m[884]&m[885]&~m[887]&~m[888])|(m[883]&~m[884]&~m[885]&~m[887]&m[888])|(~m[883]&m[884]&~m[885]&~m[887]&m[888])|(m[883]&m[884]&~m[885]&~m[887]&m[888])|(~m[883]&~m[884]&m[885]&~m[887]&m[888])|(m[883]&~m[884]&m[885]&~m[887]&m[888])|(~m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&~m[887]&m[888])|(m[883]&m[884]&m[885]&m[887]&m[888]));
    m[891] = (((m[888]&~m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&m[889]&~m[890]&~m[892]&~m[893])|(~m[888]&~m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&m[892]&~m[893])|(~m[888]&~m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&m[892]&m[893])|(m[888]&~m[889]&m[890]&m[892]&m[893])|(~m[888]&m[889]&m[890]&m[892]&m[893]))&UnbiasedRNG[585])|((m[888]&m[889]&~m[890]&~m[892]&~m[893])|(m[888]&~m[889]&m[890]&~m[892]&~m[893])|(~m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&m[889]&m[890]&~m[892]&~m[893])|(m[888]&~m[889]&~m[890]&~m[892]&m[893])|(~m[888]&m[889]&~m[890]&~m[892]&m[893])|(m[888]&m[889]&~m[890]&~m[892]&m[893])|(~m[888]&~m[889]&m[890]&~m[892]&m[893])|(m[888]&~m[889]&m[890]&~m[892]&m[893])|(~m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&~m[892]&m[893])|(m[888]&m[889]&m[890]&m[892]&m[893]));
    m[896] = (((m[893]&~m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&m[894]&~m[895]&~m[897]&~m[898])|(~m[893]&~m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&m[897]&~m[898])|(~m[893]&~m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&m[897]&m[898])|(m[893]&~m[894]&m[895]&m[897]&m[898])|(~m[893]&m[894]&m[895]&m[897]&m[898]))&UnbiasedRNG[586])|((m[893]&m[894]&~m[895]&~m[897]&~m[898])|(m[893]&~m[894]&m[895]&~m[897]&~m[898])|(~m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&m[894]&m[895]&~m[897]&~m[898])|(m[893]&~m[894]&~m[895]&~m[897]&m[898])|(~m[893]&m[894]&~m[895]&~m[897]&m[898])|(m[893]&m[894]&~m[895]&~m[897]&m[898])|(~m[893]&~m[894]&m[895]&~m[897]&m[898])|(m[893]&~m[894]&m[895]&~m[897]&m[898])|(~m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&~m[897]&m[898])|(m[893]&m[894]&m[895]&m[897]&m[898]));
    m[901] = (((m[898]&~m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&m[899]&~m[900]&~m[902]&~m[903])|(~m[898]&~m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&m[902]&~m[903])|(~m[898]&~m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&m[902]&m[903])|(m[898]&~m[899]&m[900]&m[902]&m[903])|(~m[898]&m[899]&m[900]&m[902]&m[903]))&UnbiasedRNG[587])|((m[898]&m[899]&~m[900]&~m[902]&~m[903])|(m[898]&~m[899]&m[900]&~m[902]&~m[903])|(~m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&m[899]&m[900]&~m[902]&~m[903])|(m[898]&~m[899]&~m[900]&~m[902]&m[903])|(~m[898]&m[899]&~m[900]&~m[902]&m[903])|(m[898]&m[899]&~m[900]&~m[902]&m[903])|(~m[898]&~m[899]&m[900]&~m[902]&m[903])|(m[898]&~m[899]&m[900]&~m[902]&m[903])|(~m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&~m[902]&m[903])|(m[898]&m[899]&m[900]&m[902]&m[903]));
    m[911] = (((m[908]&~m[909]&~m[910]&~m[912]&~m[913])|(~m[908]&m[909]&~m[910]&~m[912]&~m[913])|(~m[908]&~m[909]&m[910]&~m[912]&~m[913])|(m[908]&m[909]&m[910]&m[912]&~m[913])|(~m[908]&~m[909]&~m[910]&~m[912]&m[913])|(m[908]&m[909]&~m[910]&m[912]&m[913])|(m[908]&~m[909]&m[910]&m[912]&m[913])|(~m[908]&m[909]&m[910]&m[912]&m[913]))&UnbiasedRNG[588])|((m[908]&m[909]&~m[910]&~m[912]&~m[913])|(m[908]&~m[909]&m[910]&~m[912]&~m[913])|(~m[908]&m[909]&m[910]&~m[912]&~m[913])|(m[908]&m[909]&m[910]&~m[912]&~m[913])|(m[908]&~m[909]&~m[910]&~m[912]&m[913])|(~m[908]&m[909]&~m[910]&~m[912]&m[913])|(m[908]&m[909]&~m[910]&~m[912]&m[913])|(~m[908]&~m[909]&m[910]&~m[912]&m[913])|(m[908]&~m[909]&m[910]&~m[912]&m[913])|(~m[908]&m[909]&m[910]&~m[912]&m[913])|(m[908]&m[909]&m[910]&~m[912]&m[913])|(m[908]&m[909]&m[910]&m[912]&m[913]));
    m[916] = (((m[913]&~m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&m[914]&~m[915]&~m[917]&~m[918])|(~m[913]&~m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&m[917]&~m[918])|(~m[913]&~m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&m[917]&m[918])|(m[913]&~m[914]&m[915]&m[917]&m[918])|(~m[913]&m[914]&m[915]&m[917]&m[918]))&UnbiasedRNG[589])|((m[913]&m[914]&~m[915]&~m[917]&~m[918])|(m[913]&~m[914]&m[915]&~m[917]&~m[918])|(~m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&m[914]&m[915]&~m[917]&~m[918])|(m[913]&~m[914]&~m[915]&~m[917]&m[918])|(~m[913]&m[914]&~m[915]&~m[917]&m[918])|(m[913]&m[914]&~m[915]&~m[917]&m[918])|(~m[913]&~m[914]&m[915]&~m[917]&m[918])|(m[913]&~m[914]&m[915]&~m[917]&m[918])|(~m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&~m[917]&m[918])|(m[913]&m[914]&m[915]&m[917]&m[918]));
    m[921] = (((m[918]&~m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&m[919]&~m[920]&~m[922]&~m[923])|(~m[918]&~m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&m[922]&~m[923])|(~m[918]&~m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&m[922]&m[923])|(m[918]&~m[919]&m[920]&m[922]&m[923])|(~m[918]&m[919]&m[920]&m[922]&m[923]))&UnbiasedRNG[590])|((m[918]&m[919]&~m[920]&~m[922]&~m[923])|(m[918]&~m[919]&m[920]&~m[922]&~m[923])|(~m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&m[919]&m[920]&~m[922]&~m[923])|(m[918]&~m[919]&~m[920]&~m[922]&m[923])|(~m[918]&m[919]&~m[920]&~m[922]&m[923])|(m[918]&m[919]&~m[920]&~m[922]&m[923])|(~m[918]&~m[919]&m[920]&~m[922]&m[923])|(m[918]&~m[919]&m[920]&~m[922]&m[923])|(~m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&~m[922]&m[923])|(m[918]&m[919]&m[920]&m[922]&m[923]));
    m[926] = (((m[923]&~m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&m[924]&~m[925]&~m[927]&~m[928])|(~m[923]&~m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&m[927]&~m[928])|(~m[923]&~m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&m[927]&m[928])|(m[923]&~m[924]&m[925]&m[927]&m[928])|(~m[923]&m[924]&m[925]&m[927]&m[928]))&UnbiasedRNG[591])|((m[923]&m[924]&~m[925]&~m[927]&~m[928])|(m[923]&~m[924]&m[925]&~m[927]&~m[928])|(~m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&m[924]&m[925]&~m[927]&~m[928])|(m[923]&~m[924]&~m[925]&~m[927]&m[928])|(~m[923]&m[924]&~m[925]&~m[927]&m[928])|(m[923]&m[924]&~m[925]&~m[927]&m[928])|(~m[923]&~m[924]&m[925]&~m[927]&m[928])|(m[923]&~m[924]&m[925]&~m[927]&m[928])|(~m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&~m[927]&m[928])|(m[923]&m[924]&m[925]&m[927]&m[928]));
    m[931] = (((m[928]&~m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&m[929]&~m[930]&~m[932]&~m[933])|(~m[928]&~m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&m[932]&~m[933])|(~m[928]&~m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&m[932]&m[933])|(m[928]&~m[929]&m[930]&m[932]&m[933])|(~m[928]&m[929]&m[930]&m[932]&m[933]))&UnbiasedRNG[592])|((m[928]&m[929]&~m[930]&~m[932]&~m[933])|(m[928]&~m[929]&m[930]&~m[932]&~m[933])|(~m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&m[929]&m[930]&~m[932]&~m[933])|(m[928]&~m[929]&~m[930]&~m[932]&m[933])|(~m[928]&m[929]&~m[930]&~m[932]&m[933])|(m[928]&m[929]&~m[930]&~m[932]&m[933])|(~m[928]&~m[929]&m[930]&~m[932]&m[933])|(m[928]&~m[929]&m[930]&~m[932]&m[933])|(~m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&~m[932]&m[933])|(m[928]&m[929]&m[930]&m[932]&m[933]));
    m[936] = (((m[933]&~m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&m[934]&~m[935]&~m[937]&~m[938])|(~m[933]&~m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&m[937]&~m[938])|(~m[933]&~m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&m[937]&m[938])|(m[933]&~m[934]&m[935]&m[937]&m[938])|(~m[933]&m[934]&m[935]&m[937]&m[938]))&UnbiasedRNG[593])|((m[933]&m[934]&~m[935]&~m[937]&~m[938])|(m[933]&~m[934]&m[935]&~m[937]&~m[938])|(~m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&m[934]&m[935]&~m[937]&~m[938])|(m[933]&~m[934]&~m[935]&~m[937]&m[938])|(~m[933]&m[934]&~m[935]&~m[937]&m[938])|(m[933]&m[934]&~m[935]&~m[937]&m[938])|(~m[933]&~m[934]&m[935]&~m[937]&m[938])|(m[933]&~m[934]&m[935]&~m[937]&m[938])|(~m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&~m[937]&m[938])|(m[933]&m[934]&m[935]&m[937]&m[938]));
    m[941] = (((m[938]&~m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&m[939]&~m[940]&~m[942]&~m[943])|(~m[938]&~m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&m[942]&~m[943])|(~m[938]&~m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&m[942]&m[943])|(m[938]&~m[939]&m[940]&m[942]&m[943])|(~m[938]&m[939]&m[940]&m[942]&m[943]))&UnbiasedRNG[594])|((m[938]&m[939]&~m[940]&~m[942]&~m[943])|(m[938]&~m[939]&m[940]&~m[942]&~m[943])|(~m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&m[939]&m[940]&~m[942]&~m[943])|(m[938]&~m[939]&~m[940]&~m[942]&m[943])|(~m[938]&m[939]&~m[940]&~m[942]&m[943])|(m[938]&m[939]&~m[940]&~m[942]&m[943])|(~m[938]&~m[939]&m[940]&~m[942]&m[943])|(m[938]&~m[939]&m[940]&~m[942]&m[943])|(~m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&~m[942]&m[943])|(m[938]&m[939]&m[940]&m[942]&m[943]));
    m[946] = (((m[943]&~m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&m[944]&~m[945]&~m[947]&~m[948])|(~m[943]&~m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&m[947]&~m[948])|(~m[943]&~m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&m[947]&m[948])|(m[943]&~m[944]&m[945]&m[947]&m[948])|(~m[943]&m[944]&m[945]&m[947]&m[948]))&UnbiasedRNG[595])|((m[943]&m[944]&~m[945]&~m[947]&~m[948])|(m[943]&~m[944]&m[945]&~m[947]&~m[948])|(~m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&m[944]&m[945]&~m[947]&~m[948])|(m[943]&~m[944]&~m[945]&~m[947]&m[948])|(~m[943]&m[944]&~m[945]&~m[947]&m[948])|(m[943]&m[944]&~m[945]&~m[947]&m[948])|(~m[943]&~m[944]&m[945]&~m[947]&m[948])|(m[943]&~m[944]&m[945]&~m[947]&m[948])|(~m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&~m[947]&m[948])|(m[943]&m[944]&m[945]&m[947]&m[948]));
    m[956] = (((m[953]&~m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&m[954]&~m[955]&~m[957]&~m[958])|(~m[953]&~m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&m[957]&~m[958])|(~m[953]&~m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&m[957]&m[958])|(m[953]&~m[954]&m[955]&m[957]&m[958])|(~m[953]&m[954]&m[955]&m[957]&m[958]))&UnbiasedRNG[596])|((m[953]&m[954]&~m[955]&~m[957]&~m[958])|(m[953]&~m[954]&m[955]&~m[957]&~m[958])|(~m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&m[954]&m[955]&~m[957]&~m[958])|(m[953]&~m[954]&~m[955]&~m[957]&m[958])|(~m[953]&m[954]&~m[955]&~m[957]&m[958])|(m[953]&m[954]&~m[955]&~m[957]&m[958])|(~m[953]&~m[954]&m[955]&~m[957]&m[958])|(m[953]&~m[954]&m[955]&~m[957]&m[958])|(~m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&~m[957]&m[958])|(m[953]&m[954]&m[955]&m[957]&m[958]));
    m[961] = (((m[958]&~m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&m[959]&~m[960]&~m[962]&~m[963])|(~m[958]&~m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&m[962]&~m[963])|(~m[958]&~m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&m[962]&m[963])|(m[958]&~m[959]&m[960]&m[962]&m[963])|(~m[958]&m[959]&m[960]&m[962]&m[963]))&UnbiasedRNG[597])|((m[958]&m[959]&~m[960]&~m[962]&~m[963])|(m[958]&~m[959]&m[960]&~m[962]&~m[963])|(~m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&m[959]&m[960]&~m[962]&~m[963])|(m[958]&~m[959]&~m[960]&~m[962]&m[963])|(~m[958]&m[959]&~m[960]&~m[962]&m[963])|(m[958]&m[959]&~m[960]&~m[962]&m[963])|(~m[958]&~m[959]&m[960]&~m[962]&m[963])|(m[958]&~m[959]&m[960]&~m[962]&m[963])|(~m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&~m[962]&m[963])|(m[958]&m[959]&m[960]&m[962]&m[963]));
    m[966] = (((m[963]&~m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&m[964]&~m[965]&~m[967]&~m[968])|(~m[963]&~m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&m[967]&~m[968])|(~m[963]&~m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&m[967]&m[968])|(m[963]&~m[964]&m[965]&m[967]&m[968])|(~m[963]&m[964]&m[965]&m[967]&m[968]))&UnbiasedRNG[598])|((m[963]&m[964]&~m[965]&~m[967]&~m[968])|(m[963]&~m[964]&m[965]&~m[967]&~m[968])|(~m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&m[964]&m[965]&~m[967]&~m[968])|(m[963]&~m[964]&~m[965]&~m[967]&m[968])|(~m[963]&m[964]&~m[965]&~m[967]&m[968])|(m[963]&m[964]&~m[965]&~m[967]&m[968])|(~m[963]&~m[964]&m[965]&~m[967]&m[968])|(m[963]&~m[964]&m[965]&~m[967]&m[968])|(~m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&~m[967]&m[968])|(m[963]&m[964]&m[965]&m[967]&m[968]));
    m[971] = (((m[968]&~m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&m[969]&~m[970]&~m[972]&~m[973])|(~m[968]&~m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&m[972]&~m[973])|(~m[968]&~m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&m[972]&m[973])|(m[968]&~m[969]&m[970]&m[972]&m[973])|(~m[968]&m[969]&m[970]&m[972]&m[973]))&UnbiasedRNG[599])|((m[968]&m[969]&~m[970]&~m[972]&~m[973])|(m[968]&~m[969]&m[970]&~m[972]&~m[973])|(~m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&m[969]&m[970]&~m[972]&~m[973])|(m[968]&~m[969]&~m[970]&~m[972]&m[973])|(~m[968]&m[969]&~m[970]&~m[972]&m[973])|(m[968]&m[969]&~m[970]&~m[972]&m[973])|(~m[968]&~m[969]&m[970]&~m[972]&m[973])|(m[968]&~m[969]&m[970]&~m[972]&m[973])|(~m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&~m[972]&m[973])|(m[968]&m[969]&m[970]&m[972]&m[973]));
    m[976] = (((m[973]&~m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&m[974]&~m[975]&~m[977]&~m[978])|(~m[973]&~m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&m[977]&~m[978])|(~m[973]&~m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&m[977]&m[978])|(m[973]&~m[974]&m[975]&m[977]&m[978])|(~m[973]&m[974]&m[975]&m[977]&m[978]))&UnbiasedRNG[600])|((m[973]&m[974]&~m[975]&~m[977]&~m[978])|(m[973]&~m[974]&m[975]&~m[977]&~m[978])|(~m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&m[974]&m[975]&~m[977]&~m[978])|(m[973]&~m[974]&~m[975]&~m[977]&m[978])|(~m[973]&m[974]&~m[975]&~m[977]&m[978])|(m[973]&m[974]&~m[975]&~m[977]&m[978])|(~m[973]&~m[974]&m[975]&~m[977]&m[978])|(m[973]&~m[974]&m[975]&~m[977]&m[978])|(~m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&~m[977]&m[978])|(m[973]&m[974]&m[975]&m[977]&m[978]));
    m[981] = (((m[978]&~m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&m[979]&~m[980]&~m[982]&~m[983])|(~m[978]&~m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&m[982]&~m[983])|(~m[978]&~m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&m[982]&m[983])|(m[978]&~m[979]&m[980]&m[982]&m[983])|(~m[978]&m[979]&m[980]&m[982]&m[983]))&UnbiasedRNG[601])|((m[978]&m[979]&~m[980]&~m[982]&~m[983])|(m[978]&~m[979]&m[980]&~m[982]&~m[983])|(~m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&m[979]&m[980]&~m[982]&~m[983])|(m[978]&~m[979]&~m[980]&~m[982]&m[983])|(~m[978]&m[979]&~m[980]&~m[982]&m[983])|(m[978]&m[979]&~m[980]&~m[982]&m[983])|(~m[978]&~m[979]&m[980]&~m[982]&m[983])|(m[978]&~m[979]&m[980]&~m[982]&m[983])|(~m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&~m[982]&m[983])|(m[978]&m[979]&m[980]&m[982]&m[983]));
    m[986] = (((m[983]&~m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&m[984]&~m[985]&~m[987]&~m[988])|(~m[983]&~m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&m[987]&~m[988])|(~m[983]&~m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&m[987]&m[988])|(m[983]&~m[984]&m[985]&m[987]&m[988])|(~m[983]&m[984]&m[985]&m[987]&m[988]))&UnbiasedRNG[602])|((m[983]&m[984]&~m[985]&~m[987]&~m[988])|(m[983]&~m[984]&m[985]&~m[987]&~m[988])|(~m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&m[984]&m[985]&~m[987]&~m[988])|(m[983]&~m[984]&~m[985]&~m[987]&m[988])|(~m[983]&m[984]&~m[985]&~m[987]&m[988])|(m[983]&m[984]&~m[985]&~m[987]&m[988])|(~m[983]&~m[984]&m[985]&~m[987]&m[988])|(m[983]&~m[984]&m[985]&~m[987]&m[988])|(~m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&~m[987]&m[988])|(m[983]&m[984]&m[985]&m[987]&m[988]));
    m[991] = (((m[988]&~m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&m[989]&~m[990]&~m[992]&~m[993])|(~m[988]&~m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&m[992]&~m[993])|(~m[988]&~m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&m[992]&m[993])|(m[988]&~m[989]&m[990]&m[992]&m[993])|(~m[988]&m[989]&m[990]&m[992]&m[993]))&UnbiasedRNG[603])|((m[988]&m[989]&~m[990]&~m[992]&~m[993])|(m[988]&~m[989]&m[990]&~m[992]&~m[993])|(~m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&m[989]&m[990]&~m[992]&~m[993])|(m[988]&~m[989]&~m[990]&~m[992]&m[993])|(~m[988]&m[989]&~m[990]&~m[992]&m[993])|(m[988]&m[989]&~m[990]&~m[992]&m[993])|(~m[988]&~m[989]&m[990]&~m[992]&m[993])|(m[988]&~m[989]&m[990]&~m[992]&m[993])|(~m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&~m[992]&m[993])|(m[988]&m[989]&m[990]&m[992]&m[993]));
    m[996] = (((m[993]&~m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&m[994]&~m[995]&~m[997]&~m[998])|(~m[993]&~m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&m[997]&~m[998])|(~m[993]&~m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&m[997]&m[998])|(m[993]&~m[994]&m[995]&m[997]&m[998])|(~m[993]&m[994]&m[995]&m[997]&m[998]))&UnbiasedRNG[604])|((m[993]&m[994]&~m[995]&~m[997]&~m[998])|(m[993]&~m[994]&m[995]&~m[997]&~m[998])|(~m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&m[994]&m[995]&~m[997]&~m[998])|(m[993]&~m[994]&~m[995]&~m[997]&m[998])|(~m[993]&m[994]&~m[995]&~m[997]&m[998])|(m[993]&m[994]&~m[995]&~m[997]&m[998])|(~m[993]&~m[994]&m[995]&~m[997]&m[998])|(m[993]&~m[994]&m[995]&~m[997]&m[998])|(~m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&~m[997]&m[998])|(m[993]&m[994]&m[995]&m[997]&m[998]));
    m[1006] = (((m[1003]&~m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&~m[1008])|(~m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&m[1007]&m[1008]))&UnbiasedRNG[605])|((m[1003]&m[1004]&~m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&~m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&~m[1008])|(m[1003]&~m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&~m[1005]&~m[1007]&m[1008])|(~m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&~m[1004]&m[1005]&~m[1007]&m[1008])|(~m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&~m[1007]&m[1008])|(m[1003]&m[1004]&m[1005]&m[1007]&m[1008]));
    m[1011] = (((m[1008]&~m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&~m[1013])|(~m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&m[1012]&m[1013]))&UnbiasedRNG[606])|((m[1008]&m[1009]&~m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&~m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&~m[1013])|(m[1008]&~m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&~m[1010]&~m[1012]&m[1013])|(~m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&~m[1009]&m[1010]&~m[1012]&m[1013])|(~m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&~m[1012]&m[1013])|(m[1008]&m[1009]&m[1010]&m[1012]&m[1013]));
    m[1016] = (((m[1013]&~m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&~m[1018])|(~m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&m[1017]&m[1018]))&UnbiasedRNG[607])|((m[1013]&m[1014]&~m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&~m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&~m[1018])|(m[1013]&~m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&~m[1015]&~m[1017]&m[1018])|(~m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&~m[1014]&m[1015]&~m[1017]&m[1018])|(~m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&~m[1017]&m[1018])|(m[1013]&m[1014]&m[1015]&m[1017]&m[1018]));
    m[1021] = (((m[1018]&~m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&~m[1023])|(~m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&m[1022]&m[1023]))&UnbiasedRNG[608])|((m[1018]&m[1019]&~m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&~m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&~m[1023])|(m[1018]&~m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&~m[1020]&~m[1022]&m[1023])|(~m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&~m[1019]&m[1020]&~m[1022]&m[1023])|(~m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&~m[1022]&m[1023])|(m[1018]&m[1019]&m[1020]&m[1022]&m[1023]));
    m[1026] = (((m[1023]&~m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&~m[1028])|(~m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&m[1027]&m[1028]))&UnbiasedRNG[609])|((m[1023]&m[1024]&~m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&~m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&~m[1028])|(m[1023]&~m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&~m[1025]&~m[1027]&m[1028])|(~m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&~m[1024]&m[1025]&~m[1027]&m[1028])|(~m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&~m[1027]&m[1028])|(m[1023]&m[1024]&m[1025]&m[1027]&m[1028]));
    m[1031] = (((m[1028]&~m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&~m[1033])|(~m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&m[1032]&m[1033]))&UnbiasedRNG[610])|((m[1028]&m[1029]&~m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&~m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&~m[1033])|(m[1028]&~m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&~m[1030]&~m[1032]&m[1033])|(~m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&~m[1029]&m[1030]&~m[1032]&m[1033])|(~m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&~m[1032]&m[1033])|(m[1028]&m[1029]&m[1030]&m[1032]&m[1033]));
    m[1036] = (((m[1033]&~m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&~m[1038])|(~m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&m[1037]&m[1038]))&UnbiasedRNG[611])|((m[1033]&m[1034]&~m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&~m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&~m[1038])|(m[1033]&~m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&~m[1035]&~m[1037]&m[1038])|(~m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&~m[1034]&m[1035]&~m[1037]&m[1038])|(~m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&~m[1037]&m[1038])|(m[1033]&m[1034]&m[1035]&m[1037]&m[1038]));
    m[1041] = (((m[1038]&~m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&~m[1043])|(~m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&m[1042]&m[1043]))&UnbiasedRNG[612])|((m[1038]&m[1039]&~m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&~m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&~m[1043])|(m[1038]&~m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&~m[1040]&~m[1042]&m[1043])|(~m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&~m[1039]&m[1040]&~m[1042]&m[1043])|(~m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&~m[1042]&m[1043])|(m[1038]&m[1039]&m[1040]&m[1042]&m[1043]));
    m[1046] = (((m[1043]&~m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&~m[1048])|(~m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&m[1047]&m[1048]))&UnbiasedRNG[613])|((m[1043]&m[1044]&~m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&~m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&~m[1048])|(m[1043]&~m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&~m[1045]&~m[1047]&m[1048])|(~m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&~m[1044]&m[1045]&~m[1047]&m[1048])|(~m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&~m[1047]&m[1048])|(m[1043]&m[1044]&m[1045]&m[1047]&m[1048]));
    m[1051] = (((m[1048]&~m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&~m[1053])|(~m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&m[1052]&m[1053]))&UnbiasedRNG[614])|((m[1048]&m[1049]&~m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&~m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&~m[1053])|(m[1048]&~m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&~m[1050]&~m[1052]&m[1053])|(~m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&~m[1049]&m[1050]&~m[1052]&m[1053])|(~m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&~m[1052]&m[1053])|(m[1048]&m[1049]&m[1050]&m[1052]&m[1053]));
    m[1061] = (((m[1058]&~m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&~m[1063])|(~m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&m[1062]&m[1063]))&UnbiasedRNG[615])|((m[1058]&m[1059]&~m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&~m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&~m[1063])|(m[1058]&~m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&~m[1060]&~m[1062]&m[1063])|(~m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&~m[1059]&m[1060]&~m[1062]&m[1063])|(~m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&~m[1062]&m[1063])|(m[1058]&m[1059]&m[1060]&m[1062]&m[1063]));
    m[1066] = (((m[1063]&~m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&~m[1068])|(~m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&m[1067]&m[1068]))&UnbiasedRNG[616])|((m[1063]&m[1064]&~m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&~m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&~m[1068])|(m[1063]&~m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&~m[1065]&~m[1067]&m[1068])|(~m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&~m[1064]&m[1065]&~m[1067]&m[1068])|(~m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&~m[1067]&m[1068])|(m[1063]&m[1064]&m[1065]&m[1067]&m[1068]));
    m[1071] = (((m[1068]&~m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&~m[1073])|(~m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&m[1072]&m[1073]))&UnbiasedRNG[617])|((m[1068]&m[1069]&~m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&~m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&~m[1073])|(m[1068]&~m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&~m[1070]&~m[1072]&m[1073])|(~m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&~m[1069]&m[1070]&~m[1072]&m[1073])|(~m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&~m[1072]&m[1073])|(m[1068]&m[1069]&m[1070]&m[1072]&m[1073]));
    m[1076] = (((m[1073]&~m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&~m[1078])|(~m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&m[1077]&m[1078]))&UnbiasedRNG[618])|((m[1073]&m[1074]&~m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&~m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&~m[1078])|(m[1073]&~m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&~m[1075]&~m[1077]&m[1078])|(~m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&~m[1074]&m[1075]&~m[1077]&m[1078])|(~m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&~m[1077]&m[1078])|(m[1073]&m[1074]&m[1075]&m[1077]&m[1078]));
    m[1081] = (((m[1078]&~m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&~m[1083])|(~m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&m[1082]&m[1083]))&UnbiasedRNG[619])|((m[1078]&m[1079]&~m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&~m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&~m[1083])|(m[1078]&~m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&~m[1080]&~m[1082]&m[1083])|(~m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&~m[1079]&m[1080]&~m[1082]&m[1083])|(~m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&~m[1082]&m[1083])|(m[1078]&m[1079]&m[1080]&m[1082]&m[1083]));
    m[1086] = (((m[1083]&~m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&~m[1088])|(~m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&m[1087]&m[1088]))&UnbiasedRNG[620])|((m[1083]&m[1084]&~m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&~m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&~m[1088])|(m[1083]&~m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&~m[1085]&~m[1087]&m[1088])|(~m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&~m[1084]&m[1085]&~m[1087]&m[1088])|(~m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&~m[1087]&m[1088])|(m[1083]&m[1084]&m[1085]&m[1087]&m[1088]));
    m[1091] = (((m[1088]&~m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&~m[1093])|(~m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&m[1092]&m[1093]))&UnbiasedRNG[621])|((m[1088]&m[1089]&~m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&~m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&~m[1093])|(m[1088]&~m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&~m[1090]&~m[1092]&m[1093])|(~m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&~m[1089]&m[1090]&~m[1092]&m[1093])|(~m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&~m[1092]&m[1093])|(m[1088]&m[1089]&m[1090]&m[1092]&m[1093]));
    m[1096] = (((m[1093]&~m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&~m[1098])|(~m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&m[1097]&m[1098]))&UnbiasedRNG[622])|((m[1093]&m[1094]&~m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&~m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&~m[1098])|(m[1093]&~m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&~m[1095]&~m[1097]&m[1098])|(~m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&~m[1094]&m[1095]&~m[1097]&m[1098])|(~m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&~m[1097]&m[1098])|(m[1093]&m[1094]&m[1095]&m[1097]&m[1098]));
    m[1101] = (((m[1098]&~m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&~m[1103])|(~m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&m[1102]&m[1103]))&UnbiasedRNG[623])|((m[1098]&m[1099]&~m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&~m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&~m[1103])|(m[1098]&~m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&~m[1100]&~m[1102]&m[1103])|(~m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&~m[1099]&m[1100]&~m[1102]&m[1103])|(~m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&~m[1102]&m[1103])|(m[1098]&m[1099]&m[1100]&m[1102]&m[1103]));
    m[1106] = (((m[1103]&~m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&~m[1108])|(~m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&m[1107]&m[1108]))&UnbiasedRNG[624])|((m[1103]&m[1104]&~m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&~m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&~m[1108])|(m[1103]&~m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&~m[1105]&~m[1107]&m[1108])|(~m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&~m[1104]&m[1105]&~m[1107]&m[1108])|(~m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&~m[1107]&m[1108])|(m[1103]&m[1104]&m[1105]&m[1107]&m[1108]));
    m[1111] = (((m[1108]&~m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&~m[1113])|(~m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&m[1112]&m[1113]))&UnbiasedRNG[625])|((m[1108]&m[1109]&~m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&~m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&~m[1113])|(m[1108]&~m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&~m[1110]&~m[1112]&m[1113])|(~m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&~m[1109]&m[1110]&~m[1112]&m[1113])|(~m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&~m[1112]&m[1113])|(m[1108]&m[1109]&m[1110]&m[1112]&m[1113]));
    m[1121] = (((m[1118]&~m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&~m[1123])|(~m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&m[1122]&m[1123]))&UnbiasedRNG[626])|((m[1118]&m[1119]&~m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&~m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&~m[1123])|(m[1118]&~m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&~m[1120]&~m[1122]&m[1123])|(~m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&~m[1119]&m[1120]&~m[1122]&m[1123])|(~m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&~m[1122]&m[1123])|(m[1118]&m[1119]&m[1120]&m[1122]&m[1123]));
    m[1126] = (((m[1123]&~m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&~m[1128])|(~m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&m[1127]&m[1128]))&UnbiasedRNG[627])|((m[1123]&m[1124]&~m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&~m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&~m[1128])|(m[1123]&~m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&~m[1125]&~m[1127]&m[1128])|(~m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&~m[1124]&m[1125]&~m[1127]&m[1128])|(~m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&~m[1127]&m[1128])|(m[1123]&m[1124]&m[1125]&m[1127]&m[1128]));
    m[1131] = (((m[1128]&~m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&~m[1133])|(~m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&m[1132]&m[1133]))&UnbiasedRNG[628])|((m[1128]&m[1129]&~m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&~m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&~m[1133])|(m[1128]&~m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&~m[1130]&~m[1132]&m[1133])|(~m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&~m[1129]&m[1130]&~m[1132]&m[1133])|(~m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&~m[1132]&m[1133])|(m[1128]&m[1129]&m[1130]&m[1132]&m[1133]));
    m[1136] = (((m[1133]&~m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&~m[1138])|(~m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&m[1137]&m[1138]))&UnbiasedRNG[629])|((m[1133]&m[1134]&~m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&~m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&~m[1138])|(m[1133]&~m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&~m[1135]&~m[1137]&m[1138])|(~m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&~m[1134]&m[1135]&~m[1137]&m[1138])|(~m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&~m[1137]&m[1138])|(m[1133]&m[1134]&m[1135]&m[1137]&m[1138]));
    m[1141] = (((m[1138]&~m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&~m[1143])|(~m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&m[1142]&m[1143]))&UnbiasedRNG[630])|((m[1138]&m[1139]&~m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&~m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&~m[1143])|(m[1138]&~m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&~m[1140]&~m[1142]&m[1143])|(~m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&~m[1139]&m[1140]&~m[1142]&m[1143])|(~m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&~m[1142]&m[1143])|(m[1138]&m[1139]&m[1140]&m[1142]&m[1143]));
    m[1146] = (((m[1143]&~m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&~m[1148])|(~m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&m[1147]&m[1148]))&UnbiasedRNG[631])|((m[1143]&m[1144]&~m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&~m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&~m[1148])|(m[1143]&~m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&~m[1145]&~m[1147]&m[1148])|(~m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&~m[1144]&m[1145]&~m[1147]&m[1148])|(~m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&~m[1147]&m[1148])|(m[1143]&m[1144]&m[1145]&m[1147]&m[1148]));
    m[1151] = (((m[1148]&~m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&~m[1153])|(~m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&m[1152]&m[1153]))&UnbiasedRNG[632])|((m[1148]&m[1149]&~m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&~m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&~m[1153])|(m[1148]&~m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&~m[1150]&~m[1152]&m[1153])|(~m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&~m[1149]&m[1150]&~m[1152]&m[1153])|(~m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&~m[1152]&m[1153])|(m[1148]&m[1149]&m[1150]&m[1152]&m[1153]));
    m[1156] = (((m[1153]&~m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&~m[1158])|(~m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&m[1157]&m[1158]))&UnbiasedRNG[633])|((m[1153]&m[1154]&~m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&~m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&~m[1158])|(m[1153]&~m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&~m[1155]&~m[1157]&m[1158])|(~m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&~m[1154]&m[1155]&~m[1157]&m[1158])|(~m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&~m[1157]&m[1158])|(m[1153]&m[1154]&m[1155]&m[1157]&m[1158]));
    m[1161] = (((m[1158]&~m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&~m[1163])|(~m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&m[1162]&m[1163]))&UnbiasedRNG[634])|((m[1158]&m[1159]&~m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&~m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&~m[1163])|(m[1158]&~m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&~m[1160]&~m[1162]&m[1163])|(~m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&~m[1159]&m[1160]&~m[1162]&m[1163])|(~m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&~m[1162]&m[1163])|(m[1158]&m[1159]&m[1160]&m[1162]&m[1163]));
    m[1166] = (((m[1163]&~m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&~m[1168])|(~m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&m[1167]&m[1168]))&UnbiasedRNG[635])|((m[1163]&m[1164]&~m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&~m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&~m[1168])|(m[1163]&~m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&~m[1165]&~m[1167]&m[1168])|(~m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&~m[1164]&m[1165]&~m[1167]&m[1168])|(~m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&~m[1167]&m[1168])|(m[1163]&m[1164]&m[1165]&m[1167]&m[1168]));
    m[1171] = (((m[1168]&~m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&~m[1173])|(~m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&m[1172]&m[1173]))&UnbiasedRNG[636])|((m[1168]&m[1169]&~m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&~m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&~m[1173])|(m[1168]&~m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&~m[1170]&~m[1172]&m[1173])|(~m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&~m[1169]&m[1170]&~m[1172]&m[1173])|(~m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&~m[1172]&m[1173])|(m[1168]&m[1169]&m[1170]&m[1172]&m[1173]));
    m[1176] = (((m[1173]&~m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&~m[1178])|(~m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&m[1177]&m[1178]))&UnbiasedRNG[637])|((m[1173]&m[1174]&~m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&~m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&~m[1178])|(m[1173]&~m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&~m[1175]&~m[1177]&m[1178])|(~m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&~m[1174]&m[1175]&~m[1177]&m[1178])|(~m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&~m[1177]&m[1178])|(m[1173]&m[1174]&m[1175]&m[1177]&m[1178]));
    m[1186] = (((m[1183]&~m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&~m[1188])|(~m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&m[1187]&m[1188]))&UnbiasedRNG[638])|((m[1183]&m[1184]&~m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&~m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&~m[1188])|(m[1183]&~m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&~m[1185]&~m[1187]&m[1188])|(~m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&~m[1184]&m[1185]&~m[1187]&m[1188])|(~m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&~m[1187]&m[1188])|(m[1183]&m[1184]&m[1185]&m[1187]&m[1188]));
    m[1191] = (((m[1188]&~m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&~m[1193])|(~m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&m[1192]&m[1193]))&UnbiasedRNG[639])|((m[1188]&m[1189]&~m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&~m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&~m[1193])|(m[1188]&~m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&~m[1190]&~m[1192]&m[1193])|(~m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&~m[1189]&m[1190]&~m[1192]&m[1193])|(~m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&~m[1192]&m[1193])|(m[1188]&m[1189]&m[1190]&m[1192]&m[1193]));
    m[1196] = (((m[1193]&~m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&~m[1198])|(~m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&m[1197]&m[1198]))&UnbiasedRNG[640])|((m[1193]&m[1194]&~m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&~m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&~m[1198])|(m[1193]&~m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&~m[1195]&~m[1197]&m[1198])|(~m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&~m[1194]&m[1195]&~m[1197]&m[1198])|(~m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&~m[1197]&m[1198])|(m[1193]&m[1194]&m[1195]&m[1197]&m[1198]));
    m[1201] = (((m[1198]&~m[1199]&~m[1200]&~m[1202]&~m[1203])|(~m[1198]&m[1199]&~m[1200]&~m[1202]&~m[1203])|(~m[1198]&~m[1199]&m[1200]&~m[1202]&~m[1203])|(m[1198]&m[1199]&m[1200]&m[1202]&~m[1203])|(~m[1198]&~m[1199]&~m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&~m[1200]&m[1202]&m[1203])|(m[1198]&~m[1199]&m[1200]&m[1202]&m[1203])|(~m[1198]&m[1199]&m[1200]&m[1202]&m[1203]))&UnbiasedRNG[641])|((m[1198]&m[1199]&~m[1200]&~m[1202]&~m[1203])|(m[1198]&~m[1199]&m[1200]&~m[1202]&~m[1203])|(~m[1198]&m[1199]&m[1200]&~m[1202]&~m[1203])|(m[1198]&m[1199]&m[1200]&~m[1202]&~m[1203])|(m[1198]&~m[1199]&~m[1200]&~m[1202]&m[1203])|(~m[1198]&m[1199]&~m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&~m[1200]&~m[1202]&m[1203])|(~m[1198]&~m[1199]&m[1200]&~m[1202]&m[1203])|(m[1198]&~m[1199]&m[1200]&~m[1202]&m[1203])|(~m[1198]&m[1199]&m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&m[1200]&~m[1202]&m[1203])|(m[1198]&m[1199]&m[1200]&m[1202]&m[1203]));
    m[1206] = (((m[1203]&~m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&~m[1208])|(~m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&m[1207]&m[1208]))&UnbiasedRNG[642])|((m[1203]&m[1204]&~m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&~m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&~m[1208])|(m[1203]&~m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&~m[1205]&~m[1207]&m[1208])|(~m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&~m[1204]&m[1205]&~m[1207]&m[1208])|(~m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&~m[1207]&m[1208])|(m[1203]&m[1204]&m[1205]&m[1207]&m[1208]));
    m[1211] = (((m[1208]&~m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&~m[1213])|(~m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&m[1212]&m[1213]))&UnbiasedRNG[643])|((m[1208]&m[1209]&~m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&~m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&~m[1213])|(m[1208]&~m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&~m[1210]&~m[1212]&m[1213])|(~m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&~m[1209]&m[1210]&~m[1212]&m[1213])|(~m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&~m[1212]&m[1213])|(m[1208]&m[1209]&m[1210]&m[1212]&m[1213]));
    m[1216] = (((m[1213]&~m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&~m[1218])|(~m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&m[1217]&m[1218]))&UnbiasedRNG[644])|((m[1213]&m[1214]&~m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&~m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&~m[1218])|(m[1213]&~m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&~m[1215]&~m[1217]&m[1218])|(~m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&~m[1214]&m[1215]&~m[1217]&m[1218])|(~m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&~m[1217]&m[1218])|(m[1213]&m[1214]&m[1215]&m[1217]&m[1218]));
    m[1221] = (((m[1218]&~m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&~m[1223])|(~m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&m[1222]&m[1223]))&UnbiasedRNG[645])|((m[1218]&m[1219]&~m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&~m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&~m[1223])|(m[1218]&~m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&~m[1220]&~m[1222]&m[1223])|(~m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&~m[1219]&m[1220]&~m[1222]&m[1223])|(~m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&~m[1222]&m[1223])|(m[1218]&m[1219]&m[1220]&m[1222]&m[1223]));
    m[1226] = (((m[1223]&~m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&~m[1228])|(~m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&m[1227]&m[1228]))&UnbiasedRNG[646])|((m[1223]&m[1224]&~m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&~m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&~m[1228])|(m[1223]&~m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&~m[1225]&~m[1227]&m[1228])|(~m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&~m[1224]&m[1225]&~m[1227]&m[1228])|(~m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&~m[1227]&m[1228])|(m[1223]&m[1224]&m[1225]&m[1227]&m[1228]));
    m[1231] = (((m[1228]&~m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&~m[1233])|(~m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&m[1232]&m[1233]))&UnbiasedRNG[647])|((m[1228]&m[1229]&~m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&~m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&~m[1233])|(m[1228]&~m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&~m[1230]&~m[1232]&m[1233])|(~m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&~m[1229]&m[1230]&~m[1232]&m[1233])|(~m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&~m[1232]&m[1233])|(m[1228]&m[1229]&m[1230]&m[1232]&m[1233]));
    m[1236] = (((m[1233]&~m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&~m[1238])|(~m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&m[1237]&m[1238]))&UnbiasedRNG[648])|((m[1233]&m[1234]&~m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&~m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&~m[1238])|(m[1233]&~m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&~m[1235]&~m[1237]&m[1238])|(~m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&~m[1234]&m[1235]&~m[1237]&m[1238])|(~m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&~m[1237]&m[1238])|(m[1233]&m[1234]&m[1235]&m[1237]&m[1238]));
    m[1241] = (((m[1238]&~m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&~m[1243])|(~m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&m[1242]&m[1243]))&UnbiasedRNG[649])|((m[1238]&m[1239]&~m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&~m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&~m[1243])|(m[1238]&~m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&~m[1240]&~m[1242]&m[1243])|(~m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&~m[1239]&m[1240]&~m[1242]&m[1243])|(~m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&~m[1242]&m[1243])|(m[1238]&m[1239]&m[1240]&m[1242]&m[1243]));
    m[1251] = (((m[1248]&~m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&~m[1253])|(~m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&m[1252]&m[1253]))&UnbiasedRNG[650])|((m[1248]&m[1249]&~m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&~m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&~m[1253])|(m[1248]&~m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&~m[1250]&~m[1252]&m[1253])|(~m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&~m[1249]&m[1250]&~m[1252]&m[1253])|(~m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&~m[1252]&m[1253])|(m[1248]&m[1249]&m[1250]&m[1252]&m[1253]));
    m[1256] = (((m[1253]&~m[1254]&~m[1255]&~m[1257]&~m[1258])|(~m[1253]&m[1254]&~m[1255]&~m[1257]&~m[1258])|(~m[1253]&~m[1254]&m[1255]&~m[1257]&~m[1258])|(m[1253]&m[1254]&m[1255]&m[1257]&~m[1258])|(~m[1253]&~m[1254]&~m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&~m[1255]&m[1257]&m[1258])|(m[1253]&~m[1254]&m[1255]&m[1257]&m[1258])|(~m[1253]&m[1254]&m[1255]&m[1257]&m[1258]))&UnbiasedRNG[651])|((m[1253]&m[1254]&~m[1255]&~m[1257]&~m[1258])|(m[1253]&~m[1254]&m[1255]&~m[1257]&~m[1258])|(~m[1253]&m[1254]&m[1255]&~m[1257]&~m[1258])|(m[1253]&m[1254]&m[1255]&~m[1257]&~m[1258])|(m[1253]&~m[1254]&~m[1255]&~m[1257]&m[1258])|(~m[1253]&m[1254]&~m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&~m[1255]&~m[1257]&m[1258])|(~m[1253]&~m[1254]&m[1255]&~m[1257]&m[1258])|(m[1253]&~m[1254]&m[1255]&~m[1257]&m[1258])|(~m[1253]&m[1254]&m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&m[1255]&~m[1257]&m[1258])|(m[1253]&m[1254]&m[1255]&m[1257]&m[1258]));
    m[1261] = (((m[1258]&~m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&~m[1263])|(~m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&m[1262]&m[1263]))&UnbiasedRNG[652])|((m[1258]&m[1259]&~m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&~m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&~m[1263])|(m[1258]&~m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&~m[1260]&~m[1262]&m[1263])|(~m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&~m[1259]&m[1260]&~m[1262]&m[1263])|(~m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&~m[1262]&m[1263])|(m[1258]&m[1259]&m[1260]&m[1262]&m[1263]));
    m[1266] = (((m[1263]&~m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&~m[1268])|(~m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&m[1267]&m[1268]))&UnbiasedRNG[653])|((m[1263]&m[1264]&~m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&~m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&~m[1268])|(m[1263]&~m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&~m[1265]&~m[1267]&m[1268])|(~m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&~m[1264]&m[1265]&~m[1267]&m[1268])|(~m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&~m[1267]&m[1268])|(m[1263]&m[1264]&m[1265]&m[1267]&m[1268]));
    m[1271] = (((m[1268]&~m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&~m[1273])|(~m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&m[1272]&m[1273]))&UnbiasedRNG[654])|((m[1268]&m[1269]&~m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&~m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&~m[1273])|(m[1268]&~m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&~m[1270]&~m[1272]&m[1273])|(~m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&~m[1269]&m[1270]&~m[1272]&m[1273])|(~m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&~m[1272]&m[1273])|(m[1268]&m[1269]&m[1270]&m[1272]&m[1273]));
    m[1276] = (((m[1273]&~m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&~m[1278])|(~m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&m[1277]&m[1278]))&UnbiasedRNG[655])|((m[1273]&m[1274]&~m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&~m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&~m[1278])|(m[1273]&~m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&~m[1275]&~m[1277]&m[1278])|(~m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&~m[1274]&m[1275]&~m[1277]&m[1278])|(~m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&~m[1277]&m[1278])|(m[1273]&m[1274]&m[1275]&m[1277]&m[1278]));
    m[1281] = (((m[1278]&~m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&~m[1283])|(~m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&m[1282]&m[1283]))&UnbiasedRNG[656])|((m[1278]&m[1279]&~m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&~m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&~m[1283])|(m[1278]&~m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&~m[1280]&~m[1282]&m[1283])|(~m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&~m[1279]&m[1280]&~m[1282]&m[1283])|(~m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&~m[1282]&m[1283])|(m[1278]&m[1279]&m[1280]&m[1282]&m[1283]));
    m[1286] = (((m[1283]&~m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&~m[1288])|(~m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&m[1287]&m[1288]))&UnbiasedRNG[657])|((m[1283]&m[1284]&~m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&~m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&~m[1288])|(m[1283]&~m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&~m[1285]&~m[1287]&m[1288])|(~m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&~m[1284]&m[1285]&~m[1287]&m[1288])|(~m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&~m[1287]&m[1288])|(m[1283]&m[1284]&m[1285]&m[1287]&m[1288]));
    m[1291] = (((m[1288]&~m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&~m[1293])|(~m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&m[1292]&m[1293]))&UnbiasedRNG[658])|((m[1288]&m[1289]&~m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&~m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&~m[1293])|(m[1288]&~m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&~m[1290]&~m[1292]&m[1293])|(~m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&~m[1289]&m[1290]&~m[1292]&m[1293])|(~m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&~m[1292]&m[1293])|(m[1288]&m[1289]&m[1290]&m[1292]&m[1293]));
    m[1296] = (((m[1293]&~m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&~m[1298])|(~m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&m[1297]&m[1298]))&UnbiasedRNG[659])|((m[1293]&m[1294]&~m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&~m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&~m[1298])|(m[1293]&~m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&~m[1295]&~m[1297]&m[1298])|(~m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&~m[1294]&m[1295]&~m[1297]&m[1298])|(~m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&~m[1297]&m[1298])|(m[1293]&m[1294]&m[1295]&m[1297]&m[1298]));
    m[1301] = (((m[1298]&~m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&~m[1303])|(~m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&m[1302]&m[1303]))&UnbiasedRNG[660])|((m[1298]&m[1299]&~m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&~m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&~m[1303])|(m[1298]&~m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&~m[1300]&~m[1302]&m[1303])|(~m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&~m[1299]&m[1300]&~m[1302]&m[1303])|(~m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&~m[1302]&m[1303])|(m[1298]&m[1299]&m[1300]&m[1302]&m[1303]));
    m[1311] = (((m[1308]&~m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&~m[1313])|(~m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&m[1312]&m[1313]))&UnbiasedRNG[661])|((m[1308]&m[1309]&~m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&~m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&~m[1313])|(m[1308]&~m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&~m[1310]&~m[1312]&m[1313])|(~m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&~m[1309]&m[1310]&~m[1312]&m[1313])|(~m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&~m[1312]&m[1313])|(m[1308]&m[1309]&m[1310]&m[1312]&m[1313]));
    m[1316] = (((m[1313]&~m[1314]&~m[1315]&~m[1317]&~m[1318])|(~m[1313]&m[1314]&~m[1315]&~m[1317]&~m[1318])|(~m[1313]&~m[1314]&m[1315]&~m[1317]&~m[1318])|(m[1313]&m[1314]&m[1315]&m[1317]&~m[1318])|(~m[1313]&~m[1314]&~m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&~m[1315]&m[1317]&m[1318])|(m[1313]&~m[1314]&m[1315]&m[1317]&m[1318])|(~m[1313]&m[1314]&m[1315]&m[1317]&m[1318]))&UnbiasedRNG[662])|((m[1313]&m[1314]&~m[1315]&~m[1317]&~m[1318])|(m[1313]&~m[1314]&m[1315]&~m[1317]&~m[1318])|(~m[1313]&m[1314]&m[1315]&~m[1317]&~m[1318])|(m[1313]&m[1314]&m[1315]&~m[1317]&~m[1318])|(m[1313]&~m[1314]&~m[1315]&~m[1317]&m[1318])|(~m[1313]&m[1314]&~m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&~m[1315]&~m[1317]&m[1318])|(~m[1313]&~m[1314]&m[1315]&~m[1317]&m[1318])|(m[1313]&~m[1314]&m[1315]&~m[1317]&m[1318])|(~m[1313]&m[1314]&m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&m[1315]&~m[1317]&m[1318])|(m[1313]&m[1314]&m[1315]&m[1317]&m[1318]));
    m[1321] = (((m[1318]&~m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&~m[1323])|(~m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&m[1322]&m[1323]))&UnbiasedRNG[663])|((m[1318]&m[1319]&~m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&~m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&~m[1323])|(m[1318]&~m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&~m[1320]&~m[1322]&m[1323])|(~m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&~m[1319]&m[1320]&~m[1322]&m[1323])|(~m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&~m[1322]&m[1323])|(m[1318]&m[1319]&m[1320]&m[1322]&m[1323]));
    m[1326] = (((m[1323]&~m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&~m[1328])|(~m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&m[1327]&m[1328]))&UnbiasedRNG[664])|((m[1323]&m[1324]&~m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&~m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&~m[1328])|(m[1323]&~m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&~m[1325]&~m[1327]&m[1328])|(~m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&~m[1324]&m[1325]&~m[1327]&m[1328])|(~m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&~m[1327]&m[1328])|(m[1323]&m[1324]&m[1325]&m[1327]&m[1328]));
    m[1331] = (((m[1328]&~m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&~m[1333])|(~m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&m[1332]&m[1333]))&UnbiasedRNG[665])|((m[1328]&m[1329]&~m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&~m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&~m[1333])|(m[1328]&~m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&~m[1330]&~m[1332]&m[1333])|(~m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&~m[1329]&m[1330]&~m[1332]&m[1333])|(~m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&~m[1332]&m[1333])|(m[1328]&m[1329]&m[1330]&m[1332]&m[1333]));
    m[1336] = (((m[1333]&~m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&~m[1338])|(~m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&m[1337]&m[1338]))&UnbiasedRNG[666])|((m[1333]&m[1334]&~m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&~m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&~m[1338])|(m[1333]&~m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&~m[1335]&~m[1337]&m[1338])|(~m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&~m[1334]&m[1335]&~m[1337]&m[1338])|(~m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&~m[1337]&m[1338])|(m[1333]&m[1334]&m[1335]&m[1337]&m[1338]));
    m[1341] = (((m[1338]&~m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&~m[1343])|(~m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&m[1342]&m[1343]))&UnbiasedRNG[667])|((m[1338]&m[1339]&~m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&~m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&~m[1343])|(m[1338]&~m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&~m[1340]&~m[1342]&m[1343])|(~m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&~m[1339]&m[1340]&~m[1342]&m[1343])|(~m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&~m[1342]&m[1343])|(m[1338]&m[1339]&m[1340]&m[1342]&m[1343]));
    m[1346] = (((m[1343]&~m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&~m[1348])|(~m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&m[1347]&m[1348]))&UnbiasedRNG[668])|((m[1343]&m[1344]&~m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&~m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&~m[1348])|(m[1343]&~m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&~m[1345]&~m[1347]&m[1348])|(~m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&~m[1344]&m[1345]&~m[1347]&m[1348])|(~m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&~m[1347]&m[1348])|(m[1343]&m[1344]&m[1345]&m[1347]&m[1348]));
    m[1351] = (((m[1348]&~m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&~m[1353])|(~m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&m[1352]&m[1353]))&UnbiasedRNG[669])|((m[1348]&m[1349]&~m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&~m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&~m[1353])|(m[1348]&~m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&~m[1350]&~m[1352]&m[1353])|(~m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&~m[1349]&m[1350]&~m[1352]&m[1353])|(~m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&~m[1352]&m[1353])|(m[1348]&m[1349]&m[1350]&m[1352]&m[1353]));
    m[1356] = (((m[1353]&~m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&~m[1358])|(~m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&m[1357]&m[1358]))&UnbiasedRNG[670])|((m[1353]&m[1354]&~m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&~m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&~m[1358])|(m[1353]&~m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&~m[1355]&~m[1357]&m[1358])|(~m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&~m[1354]&m[1355]&~m[1357]&m[1358])|(~m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&~m[1357]&m[1358])|(m[1353]&m[1354]&m[1355]&m[1357]&m[1358]));
    m[1366] = (((m[1363]&~m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&~m[1368])|(~m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&m[1367]&m[1368]))&UnbiasedRNG[671])|((m[1363]&m[1364]&~m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&~m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&~m[1368])|(m[1363]&~m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&~m[1365]&~m[1367]&m[1368])|(~m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&~m[1364]&m[1365]&~m[1367]&m[1368])|(~m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&~m[1367]&m[1368])|(m[1363]&m[1364]&m[1365]&m[1367]&m[1368]));
    m[1371] = (((m[1368]&~m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&~m[1373])|(~m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&m[1372]&m[1373]))&UnbiasedRNG[672])|((m[1368]&m[1369]&~m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&~m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&~m[1373])|(m[1368]&~m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&~m[1370]&~m[1372]&m[1373])|(~m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&~m[1369]&m[1370]&~m[1372]&m[1373])|(~m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&~m[1372]&m[1373])|(m[1368]&m[1369]&m[1370]&m[1372]&m[1373]));
    m[1376] = (((m[1373]&~m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&~m[1378])|(~m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&m[1377]&m[1378]))&UnbiasedRNG[673])|((m[1373]&m[1374]&~m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&~m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&~m[1378])|(m[1373]&~m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&~m[1375]&~m[1377]&m[1378])|(~m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&~m[1374]&m[1375]&~m[1377]&m[1378])|(~m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&~m[1377]&m[1378])|(m[1373]&m[1374]&m[1375]&m[1377]&m[1378]));
    m[1381] = (((m[1378]&~m[1379]&~m[1380]&~m[1382]&~m[1383])|(~m[1378]&m[1379]&~m[1380]&~m[1382]&~m[1383])|(~m[1378]&~m[1379]&m[1380]&~m[1382]&~m[1383])|(m[1378]&m[1379]&m[1380]&m[1382]&~m[1383])|(~m[1378]&~m[1379]&~m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&~m[1380]&m[1382]&m[1383])|(m[1378]&~m[1379]&m[1380]&m[1382]&m[1383])|(~m[1378]&m[1379]&m[1380]&m[1382]&m[1383]))&UnbiasedRNG[674])|((m[1378]&m[1379]&~m[1380]&~m[1382]&~m[1383])|(m[1378]&~m[1379]&m[1380]&~m[1382]&~m[1383])|(~m[1378]&m[1379]&m[1380]&~m[1382]&~m[1383])|(m[1378]&m[1379]&m[1380]&~m[1382]&~m[1383])|(m[1378]&~m[1379]&~m[1380]&~m[1382]&m[1383])|(~m[1378]&m[1379]&~m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&~m[1380]&~m[1382]&m[1383])|(~m[1378]&~m[1379]&m[1380]&~m[1382]&m[1383])|(m[1378]&~m[1379]&m[1380]&~m[1382]&m[1383])|(~m[1378]&m[1379]&m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&m[1380]&~m[1382]&m[1383])|(m[1378]&m[1379]&m[1380]&m[1382]&m[1383]));
    m[1386] = (((m[1383]&~m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&~m[1388])|(~m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&m[1387]&m[1388]))&UnbiasedRNG[675])|((m[1383]&m[1384]&~m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&~m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&~m[1388])|(m[1383]&~m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&~m[1385]&~m[1387]&m[1388])|(~m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&~m[1384]&m[1385]&~m[1387]&m[1388])|(~m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&~m[1387]&m[1388])|(m[1383]&m[1384]&m[1385]&m[1387]&m[1388]));
    m[1391] = (((m[1388]&~m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&~m[1393])|(~m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&m[1392]&m[1393]))&UnbiasedRNG[676])|((m[1388]&m[1389]&~m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&~m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&~m[1393])|(m[1388]&~m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&~m[1390]&~m[1392]&m[1393])|(~m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&~m[1389]&m[1390]&~m[1392]&m[1393])|(~m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&~m[1392]&m[1393])|(m[1388]&m[1389]&m[1390]&m[1392]&m[1393]));
    m[1396] = (((m[1393]&~m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&~m[1398])|(~m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&m[1397]&m[1398]))&UnbiasedRNG[677])|((m[1393]&m[1394]&~m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&~m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&~m[1398])|(m[1393]&~m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&~m[1395]&~m[1397]&m[1398])|(~m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&~m[1394]&m[1395]&~m[1397]&m[1398])|(~m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&~m[1397]&m[1398])|(m[1393]&m[1394]&m[1395]&m[1397]&m[1398]));
    m[1401] = (((m[1398]&~m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&~m[1403])|(~m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&m[1402]&m[1403]))&UnbiasedRNG[678])|((m[1398]&m[1399]&~m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&~m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&~m[1403])|(m[1398]&~m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&~m[1400]&~m[1402]&m[1403])|(~m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&~m[1399]&m[1400]&~m[1402]&m[1403])|(~m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&~m[1402]&m[1403])|(m[1398]&m[1399]&m[1400]&m[1402]&m[1403]));
    m[1406] = (((m[1403]&~m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&~m[1408])|(~m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&m[1407]&m[1408]))&UnbiasedRNG[679])|((m[1403]&m[1404]&~m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&~m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&~m[1408])|(m[1403]&~m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&~m[1405]&~m[1407]&m[1408])|(~m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&~m[1404]&m[1405]&~m[1407]&m[1408])|(~m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&~m[1407]&m[1408])|(m[1403]&m[1404]&m[1405]&m[1407]&m[1408]));
    m[1416] = (((m[1413]&~m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&~m[1418])|(~m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&m[1417]&m[1418]))&UnbiasedRNG[680])|((m[1413]&m[1414]&~m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&~m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&~m[1418])|(m[1413]&~m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&~m[1415]&~m[1417]&m[1418])|(~m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&~m[1414]&m[1415]&~m[1417]&m[1418])|(~m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&~m[1417]&m[1418])|(m[1413]&m[1414]&m[1415]&m[1417]&m[1418]));
    m[1421] = (((m[1418]&~m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&~m[1423])|(~m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&m[1422]&m[1423]))&UnbiasedRNG[681])|((m[1418]&m[1419]&~m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&~m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&~m[1423])|(m[1418]&~m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&~m[1420]&~m[1422]&m[1423])|(~m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&~m[1419]&m[1420]&~m[1422]&m[1423])|(~m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&~m[1422]&m[1423])|(m[1418]&m[1419]&m[1420]&m[1422]&m[1423]));
    m[1426] = (((m[1423]&~m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&~m[1428])|(~m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&m[1427]&m[1428]))&UnbiasedRNG[682])|((m[1423]&m[1424]&~m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&~m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&~m[1428])|(m[1423]&~m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&~m[1425]&~m[1427]&m[1428])|(~m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&~m[1424]&m[1425]&~m[1427]&m[1428])|(~m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&~m[1427]&m[1428])|(m[1423]&m[1424]&m[1425]&m[1427]&m[1428]));
    m[1431] = (((m[1428]&~m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&~m[1433])|(~m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&m[1432]&m[1433]))&UnbiasedRNG[683])|((m[1428]&m[1429]&~m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&~m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&~m[1433])|(m[1428]&~m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&~m[1430]&~m[1432]&m[1433])|(~m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&~m[1429]&m[1430]&~m[1432]&m[1433])|(~m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&~m[1432]&m[1433])|(m[1428]&m[1429]&m[1430]&m[1432]&m[1433]));
    m[1436] = (((m[1433]&~m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&~m[1438])|(~m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&m[1437]&m[1438]))&UnbiasedRNG[684])|((m[1433]&m[1434]&~m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&~m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&~m[1438])|(m[1433]&~m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&~m[1435]&~m[1437]&m[1438])|(~m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&~m[1434]&m[1435]&~m[1437]&m[1438])|(~m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&~m[1437]&m[1438])|(m[1433]&m[1434]&m[1435]&m[1437]&m[1438]));
    m[1441] = (((m[1438]&~m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&~m[1443])|(~m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&m[1442]&m[1443]))&UnbiasedRNG[685])|((m[1438]&m[1439]&~m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&~m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&~m[1443])|(m[1438]&~m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&~m[1440]&~m[1442]&m[1443])|(~m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&~m[1439]&m[1440]&~m[1442]&m[1443])|(~m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&~m[1442]&m[1443])|(m[1438]&m[1439]&m[1440]&m[1442]&m[1443]));
    m[1446] = (((m[1443]&~m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&~m[1448])|(~m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&m[1447]&m[1448]))&UnbiasedRNG[686])|((m[1443]&m[1444]&~m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&~m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&~m[1448])|(m[1443]&~m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&~m[1445]&~m[1447]&m[1448])|(~m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&~m[1444]&m[1445]&~m[1447]&m[1448])|(~m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&~m[1447]&m[1448])|(m[1443]&m[1444]&m[1445]&m[1447]&m[1448]));
    m[1451] = (((m[1448]&~m[1449]&~m[1450]&~m[1452]&~m[1453])|(~m[1448]&m[1449]&~m[1450]&~m[1452]&~m[1453])|(~m[1448]&~m[1449]&m[1450]&~m[1452]&~m[1453])|(m[1448]&m[1449]&m[1450]&m[1452]&~m[1453])|(~m[1448]&~m[1449]&~m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&~m[1450]&m[1452]&m[1453])|(m[1448]&~m[1449]&m[1450]&m[1452]&m[1453])|(~m[1448]&m[1449]&m[1450]&m[1452]&m[1453]))&UnbiasedRNG[687])|((m[1448]&m[1449]&~m[1450]&~m[1452]&~m[1453])|(m[1448]&~m[1449]&m[1450]&~m[1452]&~m[1453])|(~m[1448]&m[1449]&m[1450]&~m[1452]&~m[1453])|(m[1448]&m[1449]&m[1450]&~m[1452]&~m[1453])|(m[1448]&~m[1449]&~m[1450]&~m[1452]&m[1453])|(~m[1448]&m[1449]&~m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&~m[1450]&~m[1452]&m[1453])|(~m[1448]&~m[1449]&m[1450]&~m[1452]&m[1453])|(m[1448]&~m[1449]&m[1450]&~m[1452]&m[1453])|(~m[1448]&m[1449]&m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&m[1450]&~m[1452]&m[1453])|(m[1448]&m[1449]&m[1450]&m[1452]&m[1453]));
    m[1461] = (((m[1458]&~m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&~m[1463])|(~m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&m[1462]&m[1463]))&UnbiasedRNG[688])|((m[1458]&m[1459]&~m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&~m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&~m[1463])|(m[1458]&~m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&~m[1460]&~m[1462]&m[1463])|(~m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&~m[1459]&m[1460]&~m[1462]&m[1463])|(~m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&~m[1462]&m[1463])|(m[1458]&m[1459]&m[1460]&m[1462]&m[1463]));
    m[1466] = (((m[1463]&~m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&~m[1468])|(~m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&m[1467]&m[1468]))&UnbiasedRNG[689])|((m[1463]&m[1464]&~m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&~m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&~m[1468])|(m[1463]&~m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&~m[1465]&~m[1467]&m[1468])|(~m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&~m[1464]&m[1465]&~m[1467]&m[1468])|(~m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&~m[1467]&m[1468])|(m[1463]&m[1464]&m[1465]&m[1467]&m[1468]));
    m[1471] = (((m[1468]&~m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&~m[1473])|(~m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&m[1472]&m[1473]))&UnbiasedRNG[690])|((m[1468]&m[1469]&~m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&~m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&~m[1473])|(m[1468]&~m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&~m[1470]&~m[1472]&m[1473])|(~m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&~m[1469]&m[1470]&~m[1472]&m[1473])|(~m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&~m[1472]&m[1473])|(m[1468]&m[1469]&m[1470]&m[1472]&m[1473]));
    m[1476] = (((m[1473]&~m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&~m[1478])|(~m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&m[1477]&m[1478]))&UnbiasedRNG[691])|((m[1473]&m[1474]&~m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&~m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&~m[1478])|(m[1473]&~m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&~m[1475]&~m[1477]&m[1478])|(~m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&~m[1474]&m[1475]&~m[1477]&m[1478])|(~m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&~m[1477]&m[1478])|(m[1473]&m[1474]&m[1475]&m[1477]&m[1478]));
    m[1481] = (((m[1478]&~m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&~m[1483])|(~m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&m[1482]&m[1483]))&UnbiasedRNG[692])|((m[1478]&m[1479]&~m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&~m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&~m[1483])|(m[1478]&~m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&~m[1480]&~m[1482]&m[1483])|(~m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&~m[1479]&m[1480]&~m[1482]&m[1483])|(~m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&~m[1482]&m[1483])|(m[1478]&m[1479]&m[1480]&m[1482]&m[1483]));
    m[1486] = (((m[1483]&~m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&~m[1488])|(~m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&m[1487]&m[1488]))&UnbiasedRNG[693])|((m[1483]&m[1484]&~m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&~m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&~m[1488])|(m[1483]&~m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&~m[1485]&~m[1487]&m[1488])|(~m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&~m[1484]&m[1485]&~m[1487]&m[1488])|(~m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&~m[1487]&m[1488])|(m[1483]&m[1484]&m[1485]&m[1487]&m[1488]));
    m[1491] = (((m[1488]&~m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&~m[1493])|(~m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&m[1492]&m[1493]))&UnbiasedRNG[694])|((m[1488]&m[1489]&~m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&~m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&~m[1493])|(m[1488]&~m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&~m[1490]&~m[1492]&m[1493])|(~m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&~m[1489]&m[1490]&~m[1492]&m[1493])|(~m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&~m[1492]&m[1493])|(m[1488]&m[1489]&m[1490]&m[1492]&m[1493]));
    m[1501] = (((m[1498]&~m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&~m[1503])|(~m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&m[1502]&m[1503]))&UnbiasedRNG[695])|((m[1498]&m[1499]&~m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&~m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&~m[1503])|(m[1498]&~m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&~m[1500]&~m[1502]&m[1503])|(~m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&~m[1499]&m[1500]&~m[1502]&m[1503])|(~m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&~m[1502]&m[1503])|(m[1498]&m[1499]&m[1500]&m[1502]&m[1503]));
    m[1506] = (((m[1503]&~m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&~m[1508])|(~m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&m[1507]&m[1508]))&UnbiasedRNG[696])|((m[1503]&m[1504]&~m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&~m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&~m[1508])|(m[1503]&~m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&~m[1505]&~m[1507]&m[1508])|(~m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&~m[1504]&m[1505]&~m[1507]&m[1508])|(~m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&~m[1507]&m[1508])|(m[1503]&m[1504]&m[1505]&m[1507]&m[1508]));
    m[1511] = (((m[1508]&~m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&~m[1513])|(~m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&m[1512]&m[1513]))&UnbiasedRNG[697])|((m[1508]&m[1509]&~m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&~m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&~m[1513])|(m[1508]&~m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&~m[1510]&~m[1512]&m[1513])|(~m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&~m[1509]&m[1510]&~m[1512]&m[1513])|(~m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&~m[1512]&m[1513])|(m[1508]&m[1509]&m[1510]&m[1512]&m[1513]));
    m[1516] = (((m[1513]&~m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&~m[1518])|(~m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&m[1517]&m[1518]))&UnbiasedRNG[698])|((m[1513]&m[1514]&~m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&~m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&~m[1518])|(m[1513]&~m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&~m[1515]&~m[1517]&m[1518])|(~m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&~m[1514]&m[1515]&~m[1517]&m[1518])|(~m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&~m[1517]&m[1518])|(m[1513]&m[1514]&m[1515]&m[1517]&m[1518]));
    m[1521] = (((m[1518]&~m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&~m[1523])|(~m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&m[1522]&m[1523]))&UnbiasedRNG[699])|((m[1518]&m[1519]&~m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&~m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&~m[1523])|(m[1518]&~m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&~m[1520]&~m[1522]&m[1523])|(~m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&~m[1519]&m[1520]&~m[1522]&m[1523])|(~m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&~m[1522]&m[1523])|(m[1518]&m[1519]&m[1520]&m[1522]&m[1523]));
    m[1526] = (((m[1523]&~m[1524]&~m[1525]&~m[1527]&~m[1528])|(~m[1523]&m[1524]&~m[1525]&~m[1527]&~m[1528])|(~m[1523]&~m[1524]&m[1525]&~m[1527]&~m[1528])|(m[1523]&m[1524]&m[1525]&m[1527]&~m[1528])|(~m[1523]&~m[1524]&~m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&~m[1525]&m[1527]&m[1528])|(m[1523]&~m[1524]&m[1525]&m[1527]&m[1528])|(~m[1523]&m[1524]&m[1525]&m[1527]&m[1528]))&UnbiasedRNG[700])|((m[1523]&m[1524]&~m[1525]&~m[1527]&~m[1528])|(m[1523]&~m[1524]&m[1525]&~m[1527]&~m[1528])|(~m[1523]&m[1524]&m[1525]&~m[1527]&~m[1528])|(m[1523]&m[1524]&m[1525]&~m[1527]&~m[1528])|(m[1523]&~m[1524]&~m[1525]&~m[1527]&m[1528])|(~m[1523]&m[1524]&~m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&~m[1525]&~m[1527]&m[1528])|(~m[1523]&~m[1524]&m[1525]&~m[1527]&m[1528])|(m[1523]&~m[1524]&m[1525]&~m[1527]&m[1528])|(~m[1523]&m[1524]&m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&m[1525]&~m[1527]&m[1528])|(m[1523]&m[1524]&m[1525]&m[1527]&m[1528]));
    m[1536] = (((m[1533]&~m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&~m[1538])|(~m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&m[1537]&m[1538]))&UnbiasedRNG[701])|((m[1533]&m[1534]&~m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&~m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&~m[1538])|(m[1533]&~m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&~m[1535]&~m[1537]&m[1538])|(~m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&~m[1534]&m[1535]&~m[1537]&m[1538])|(~m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&~m[1537]&m[1538])|(m[1533]&m[1534]&m[1535]&m[1537]&m[1538]));
    m[1541] = (((m[1538]&~m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&~m[1543])|(~m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&m[1542]&m[1543]))&UnbiasedRNG[702])|((m[1538]&m[1539]&~m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&~m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&~m[1543])|(m[1538]&~m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&~m[1540]&~m[1542]&m[1543])|(~m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&~m[1539]&m[1540]&~m[1542]&m[1543])|(~m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&~m[1542]&m[1543])|(m[1538]&m[1539]&m[1540]&m[1542]&m[1543]));
    m[1546] = (((m[1543]&~m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&~m[1548])|(~m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&m[1547]&m[1548]))&UnbiasedRNG[703])|((m[1543]&m[1544]&~m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&~m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&~m[1548])|(m[1543]&~m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&~m[1545]&~m[1547]&m[1548])|(~m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&~m[1544]&m[1545]&~m[1547]&m[1548])|(~m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&~m[1547]&m[1548])|(m[1543]&m[1544]&m[1545]&m[1547]&m[1548]));
    m[1551] = (((m[1548]&~m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&~m[1553])|(~m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&m[1552]&m[1553]))&UnbiasedRNG[704])|((m[1548]&m[1549]&~m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&~m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&~m[1553])|(m[1548]&~m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&~m[1550]&~m[1552]&m[1553])|(~m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&~m[1549]&m[1550]&~m[1552]&m[1553])|(~m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&~m[1552]&m[1553])|(m[1548]&m[1549]&m[1550]&m[1552]&m[1553]));
    m[1556] = (((m[1553]&~m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&~m[1558])|(~m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&m[1557]&m[1558]))&UnbiasedRNG[705])|((m[1553]&m[1554]&~m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&~m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&~m[1558])|(m[1553]&~m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&~m[1555]&~m[1557]&m[1558])|(~m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&~m[1554]&m[1555]&~m[1557]&m[1558])|(~m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&~m[1557]&m[1558])|(m[1553]&m[1554]&m[1555]&m[1557]&m[1558]));
    m[1566] = (((m[1563]&~m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&~m[1568])|(~m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&m[1567]&m[1568]))&UnbiasedRNG[706])|((m[1563]&m[1564]&~m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&~m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&~m[1568])|(m[1563]&~m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&~m[1565]&~m[1567]&m[1568])|(~m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&~m[1564]&m[1565]&~m[1567]&m[1568])|(~m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&~m[1567]&m[1568])|(m[1563]&m[1564]&m[1565]&m[1567]&m[1568]));
    m[1571] = (((m[1568]&~m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&~m[1573])|(~m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&m[1572]&m[1573]))&UnbiasedRNG[707])|((m[1568]&m[1569]&~m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&~m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&~m[1573])|(m[1568]&~m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&~m[1570]&~m[1572]&m[1573])|(~m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&~m[1569]&m[1570]&~m[1572]&m[1573])|(~m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&~m[1572]&m[1573])|(m[1568]&m[1569]&m[1570]&m[1572]&m[1573]));
    m[1576] = (((m[1573]&~m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&~m[1578])|(~m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&m[1577]&m[1578]))&UnbiasedRNG[708])|((m[1573]&m[1574]&~m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&~m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&~m[1578])|(m[1573]&~m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&~m[1575]&~m[1577]&m[1578])|(~m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&~m[1574]&m[1575]&~m[1577]&m[1578])|(~m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&~m[1577]&m[1578])|(m[1573]&m[1574]&m[1575]&m[1577]&m[1578]));
    m[1581] = (((m[1578]&~m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&~m[1583])|(~m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&m[1582]&m[1583]))&UnbiasedRNG[709])|((m[1578]&m[1579]&~m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&~m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&~m[1583])|(m[1578]&~m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&~m[1580]&~m[1582]&m[1583])|(~m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&~m[1579]&m[1580]&~m[1582]&m[1583])|(~m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&~m[1582]&m[1583])|(m[1578]&m[1579]&m[1580]&m[1582]&m[1583]));
    m[1591] = (((m[1588]&~m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&~m[1593])|(~m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&m[1592]&m[1593]))&UnbiasedRNG[710])|((m[1588]&m[1589]&~m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&~m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&~m[1593])|(m[1588]&~m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&~m[1590]&~m[1592]&m[1593])|(~m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&~m[1589]&m[1590]&~m[1592]&m[1593])|(~m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&~m[1592]&m[1593])|(m[1588]&m[1589]&m[1590]&m[1592]&m[1593]));
    m[1596] = (((m[1593]&~m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&~m[1598])|(~m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&m[1597]&m[1598]))&UnbiasedRNG[711])|((m[1593]&m[1594]&~m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&~m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&~m[1598])|(m[1593]&~m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&~m[1595]&~m[1597]&m[1598])|(~m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&~m[1594]&m[1595]&~m[1597]&m[1598])|(~m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&~m[1597]&m[1598])|(m[1593]&m[1594]&m[1595]&m[1597]&m[1598]));
    m[1601] = (((m[1598]&~m[1599]&~m[1600]&~m[1602]&~m[1603])|(~m[1598]&m[1599]&~m[1600]&~m[1602]&~m[1603])|(~m[1598]&~m[1599]&m[1600]&~m[1602]&~m[1603])|(m[1598]&m[1599]&m[1600]&m[1602]&~m[1603])|(~m[1598]&~m[1599]&~m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&~m[1600]&m[1602]&m[1603])|(m[1598]&~m[1599]&m[1600]&m[1602]&m[1603])|(~m[1598]&m[1599]&m[1600]&m[1602]&m[1603]))&UnbiasedRNG[712])|((m[1598]&m[1599]&~m[1600]&~m[1602]&~m[1603])|(m[1598]&~m[1599]&m[1600]&~m[1602]&~m[1603])|(~m[1598]&m[1599]&m[1600]&~m[1602]&~m[1603])|(m[1598]&m[1599]&m[1600]&~m[1602]&~m[1603])|(m[1598]&~m[1599]&~m[1600]&~m[1602]&m[1603])|(~m[1598]&m[1599]&~m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&~m[1600]&~m[1602]&m[1603])|(~m[1598]&~m[1599]&m[1600]&~m[1602]&m[1603])|(m[1598]&~m[1599]&m[1600]&~m[1602]&m[1603])|(~m[1598]&m[1599]&m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&m[1600]&~m[1602]&m[1603])|(m[1598]&m[1599]&m[1600]&m[1602]&m[1603]));
    m[1611] = (((m[1608]&~m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&~m[1613])|(~m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&m[1612]&m[1613]))&UnbiasedRNG[713])|((m[1608]&m[1609]&~m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&~m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&~m[1613])|(m[1608]&~m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&~m[1610]&~m[1612]&m[1613])|(~m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&~m[1609]&m[1610]&~m[1612]&m[1613])|(~m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&~m[1612]&m[1613])|(m[1608]&m[1609]&m[1610]&m[1612]&m[1613]));
    m[1616] = (((m[1613]&~m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&~m[1618])|(~m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&m[1617]&m[1618]))&UnbiasedRNG[714])|((m[1613]&m[1614]&~m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&~m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&~m[1618])|(m[1613]&~m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&~m[1615]&~m[1617]&m[1618])|(~m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&~m[1614]&m[1615]&~m[1617]&m[1618])|(~m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&~m[1617]&m[1618])|(m[1613]&m[1614]&m[1615]&m[1617]&m[1618]));
    m[1626] = (((m[1623]&~m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&~m[1628])|(~m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&m[1627]&m[1628]))&UnbiasedRNG[715])|((m[1623]&m[1624]&~m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&~m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&~m[1628])|(m[1623]&~m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&~m[1625]&~m[1627]&m[1628])|(~m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&~m[1624]&m[1625]&~m[1627]&m[1628])|(~m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&~m[1627]&m[1628])|(m[1623]&m[1624]&m[1625]&m[1627]&m[1628]));
end

always @(posedge color4_clk) begin
    m[732] = (((m[728]&~m[729]&~m[730]&~m[731]&~m[735])|(~m[728]&m[729]&~m[730]&~m[731]&~m[735])|(~m[728]&~m[729]&m[730]&~m[731]&~m[735])|(m[728]&m[729]&~m[730]&m[731]&~m[735])|(m[728]&~m[729]&m[730]&m[731]&~m[735])|(~m[728]&m[729]&m[730]&m[731]&~m[735]))&BiasedRNG[699])|(((m[728]&~m[729]&~m[730]&~m[731]&m[735])|(~m[728]&m[729]&~m[730]&~m[731]&m[735])|(~m[728]&~m[729]&m[730]&~m[731]&m[735])|(m[728]&m[729]&~m[730]&m[731]&m[735])|(m[728]&~m[729]&m[730]&m[731]&m[735])|(~m[728]&m[729]&m[730]&m[731]&m[735]))&~BiasedRNG[699])|((m[728]&m[729]&~m[730]&~m[731]&~m[735])|(m[728]&~m[729]&m[730]&~m[731]&~m[735])|(~m[728]&m[729]&m[730]&~m[731]&~m[735])|(m[728]&m[729]&m[730]&~m[731]&~m[735])|(m[728]&m[729]&m[730]&m[731]&~m[735])|(m[728]&m[729]&~m[730]&~m[731]&m[735])|(m[728]&~m[729]&m[730]&~m[731]&m[735])|(~m[728]&m[729]&m[730]&~m[731]&m[735])|(m[728]&m[729]&m[730]&~m[731]&m[735])|(m[728]&m[729]&m[730]&m[731]&m[735]));
    m[737] = (((m[733]&~m[734]&~m[735]&~m[736]&~m[745])|(~m[733]&m[734]&~m[735]&~m[736]&~m[745])|(~m[733]&~m[734]&m[735]&~m[736]&~m[745])|(m[733]&m[734]&~m[735]&m[736]&~m[745])|(m[733]&~m[734]&m[735]&m[736]&~m[745])|(~m[733]&m[734]&m[735]&m[736]&~m[745]))&BiasedRNG[700])|(((m[733]&~m[734]&~m[735]&~m[736]&m[745])|(~m[733]&m[734]&~m[735]&~m[736]&m[745])|(~m[733]&~m[734]&m[735]&~m[736]&m[745])|(m[733]&m[734]&~m[735]&m[736]&m[745])|(m[733]&~m[734]&m[735]&m[736]&m[745])|(~m[733]&m[734]&m[735]&m[736]&m[745]))&~BiasedRNG[700])|((m[733]&m[734]&~m[735]&~m[736]&~m[745])|(m[733]&~m[734]&m[735]&~m[736]&~m[745])|(~m[733]&m[734]&m[735]&~m[736]&~m[745])|(m[733]&m[734]&m[735]&~m[736]&~m[745])|(m[733]&m[734]&m[735]&m[736]&~m[745])|(m[733]&m[734]&~m[735]&~m[736]&m[745])|(m[733]&~m[734]&m[735]&~m[736]&m[745])|(~m[733]&m[734]&m[735]&~m[736]&m[745])|(m[733]&m[734]&m[735]&~m[736]&m[745])|(m[733]&m[734]&m[735]&m[736]&m[745]));
    m[742] = (((m[738]&~m[739]&~m[740]&~m[741]&~m[750])|(~m[738]&m[739]&~m[740]&~m[741]&~m[750])|(~m[738]&~m[739]&m[740]&~m[741]&~m[750])|(m[738]&m[739]&~m[740]&m[741]&~m[750])|(m[738]&~m[739]&m[740]&m[741]&~m[750])|(~m[738]&m[739]&m[740]&m[741]&~m[750]))&BiasedRNG[701])|(((m[738]&~m[739]&~m[740]&~m[741]&m[750])|(~m[738]&m[739]&~m[740]&~m[741]&m[750])|(~m[738]&~m[739]&m[740]&~m[741]&m[750])|(m[738]&m[739]&~m[740]&m[741]&m[750])|(m[738]&~m[739]&m[740]&m[741]&m[750])|(~m[738]&m[739]&m[740]&m[741]&m[750]))&~BiasedRNG[701])|((m[738]&m[739]&~m[740]&~m[741]&~m[750])|(m[738]&~m[739]&m[740]&~m[741]&~m[750])|(~m[738]&m[739]&m[740]&~m[741]&~m[750])|(m[738]&m[739]&m[740]&~m[741]&~m[750])|(m[738]&m[739]&m[740]&m[741]&~m[750])|(m[738]&m[739]&~m[740]&~m[741]&m[750])|(m[738]&~m[739]&m[740]&~m[741]&m[750])|(~m[738]&m[739]&m[740]&~m[741]&m[750])|(m[738]&m[739]&m[740]&~m[741]&m[750])|(m[738]&m[739]&m[740]&m[741]&m[750]));
    m[747] = (((m[743]&~m[744]&~m[745]&~m[746]&~m[760])|(~m[743]&m[744]&~m[745]&~m[746]&~m[760])|(~m[743]&~m[744]&m[745]&~m[746]&~m[760])|(m[743]&m[744]&~m[745]&m[746]&~m[760])|(m[743]&~m[744]&m[745]&m[746]&~m[760])|(~m[743]&m[744]&m[745]&m[746]&~m[760]))&BiasedRNG[702])|(((m[743]&~m[744]&~m[745]&~m[746]&m[760])|(~m[743]&m[744]&~m[745]&~m[746]&m[760])|(~m[743]&~m[744]&m[745]&~m[746]&m[760])|(m[743]&m[744]&~m[745]&m[746]&m[760])|(m[743]&~m[744]&m[745]&m[746]&m[760])|(~m[743]&m[744]&m[745]&m[746]&m[760]))&~BiasedRNG[702])|((m[743]&m[744]&~m[745]&~m[746]&~m[760])|(m[743]&~m[744]&m[745]&~m[746]&~m[760])|(~m[743]&m[744]&m[745]&~m[746]&~m[760])|(m[743]&m[744]&m[745]&~m[746]&~m[760])|(m[743]&m[744]&m[745]&m[746]&~m[760])|(m[743]&m[744]&~m[745]&~m[746]&m[760])|(m[743]&~m[744]&m[745]&~m[746]&m[760])|(~m[743]&m[744]&m[745]&~m[746]&m[760])|(m[743]&m[744]&m[745]&~m[746]&m[760])|(m[743]&m[744]&m[745]&m[746]&m[760]));
    m[752] = (((m[748]&~m[749]&~m[750]&~m[751]&~m[765])|(~m[748]&m[749]&~m[750]&~m[751]&~m[765])|(~m[748]&~m[749]&m[750]&~m[751]&~m[765])|(m[748]&m[749]&~m[750]&m[751]&~m[765])|(m[748]&~m[749]&m[750]&m[751]&~m[765])|(~m[748]&m[749]&m[750]&m[751]&~m[765]))&BiasedRNG[703])|(((m[748]&~m[749]&~m[750]&~m[751]&m[765])|(~m[748]&m[749]&~m[750]&~m[751]&m[765])|(~m[748]&~m[749]&m[750]&~m[751]&m[765])|(m[748]&m[749]&~m[750]&m[751]&m[765])|(m[748]&~m[749]&m[750]&m[751]&m[765])|(~m[748]&m[749]&m[750]&m[751]&m[765]))&~BiasedRNG[703])|((m[748]&m[749]&~m[750]&~m[751]&~m[765])|(m[748]&~m[749]&m[750]&~m[751]&~m[765])|(~m[748]&m[749]&m[750]&~m[751]&~m[765])|(m[748]&m[749]&m[750]&~m[751]&~m[765])|(m[748]&m[749]&m[750]&m[751]&~m[765])|(m[748]&m[749]&~m[750]&~m[751]&m[765])|(m[748]&~m[749]&m[750]&~m[751]&m[765])|(~m[748]&m[749]&m[750]&~m[751]&m[765])|(m[748]&m[749]&m[750]&~m[751]&m[765])|(m[748]&m[749]&m[750]&m[751]&m[765]));
    m[757] = (((m[753]&~m[754]&~m[755]&~m[756]&~m[770])|(~m[753]&m[754]&~m[755]&~m[756]&~m[770])|(~m[753]&~m[754]&m[755]&~m[756]&~m[770])|(m[753]&m[754]&~m[755]&m[756]&~m[770])|(m[753]&~m[754]&m[755]&m[756]&~m[770])|(~m[753]&m[754]&m[755]&m[756]&~m[770]))&BiasedRNG[704])|(((m[753]&~m[754]&~m[755]&~m[756]&m[770])|(~m[753]&m[754]&~m[755]&~m[756]&m[770])|(~m[753]&~m[754]&m[755]&~m[756]&m[770])|(m[753]&m[754]&~m[755]&m[756]&m[770])|(m[753]&~m[754]&m[755]&m[756]&m[770])|(~m[753]&m[754]&m[755]&m[756]&m[770]))&~BiasedRNG[704])|((m[753]&m[754]&~m[755]&~m[756]&~m[770])|(m[753]&~m[754]&m[755]&~m[756]&~m[770])|(~m[753]&m[754]&m[755]&~m[756]&~m[770])|(m[753]&m[754]&m[755]&~m[756]&~m[770])|(m[753]&m[754]&m[755]&m[756]&~m[770])|(m[753]&m[754]&~m[755]&~m[756]&m[770])|(m[753]&~m[754]&m[755]&~m[756]&m[770])|(~m[753]&m[754]&m[755]&~m[756]&m[770])|(m[753]&m[754]&m[755]&~m[756]&m[770])|(m[753]&m[754]&m[755]&m[756]&m[770]));
    m[762] = (((m[758]&~m[759]&~m[760]&~m[761]&~m[780])|(~m[758]&m[759]&~m[760]&~m[761]&~m[780])|(~m[758]&~m[759]&m[760]&~m[761]&~m[780])|(m[758]&m[759]&~m[760]&m[761]&~m[780])|(m[758]&~m[759]&m[760]&m[761]&~m[780])|(~m[758]&m[759]&m[760]&m[761]&~m[780]))&BiasedRNG[705])|(((m[758]&~m[759]&~m[760]&~m[761]&m[780])|(~m[758]&m[759]&~m[760]&~m[761]&m[780])|(~m[758]&~m[759]&m[760]&~m[761]&m[780])|(m[758]&m[759]&~m[760]&m[761]&m[780])|(m[758]&~m[759]&m[760]&m[761]&m[780])|(~m[758]&m[759]&m[760]&m[761]&m[780]))&~BiasedRNG[705])|((m[758]&m[759]&~m[760]&~m[761]&~m[780])|(m[758]&~m[759]&m[760]&~m[761]&~m[780])|(~m[758]&m[759]&m[760]&~m[761]&~m[780])|(m[758]&m[759]&m[760]&~m[761]&~m[780])|(m[758]&m[759]&m[760]&m[761]&~m[780])|(m[758]&m[759]&~m[760]&~m[761]&m[780])|(m[758]&~m[759]&m[760]&~m[761]&m[780])|(~m[758]&m[759]&m[760]&~m[761]&m[780])|(m[758]&m[759]&m[760]&~m[761]&m[780])|(m[758]&m[759]&m[760]&m[761]&m[780]));
    m[767] = (((m[763]&~m[764]&~m[765]&~m[766]&~m[785])|(~m[763]&m[764]&~m[765]&~m[766]&~m[785])|(~m[763]&~m[764]&m[765]&~m[766]&~m[785])|(m[763]&m[764]&~m[765]&m[766]&~m[785])|(m[763]&~m[764]&m[765]&m[766]&~m[785])|(~m[763]&m[764]&m[765]&m[766]&~m[785]))&BiasedRNG[706])|(((m[763]&~m[764]&~m[765]&~m[766]&m[785])|(~m[763]&m[764]&~m[765]&~m[766]&m[785])|(~m[763]&~m[764]&m[765]&~m[766]&m[785])|(m[763]&m[764]&~m[765]&m[766]&m[785])|(m[763]&~m[764]&m[765]&m[766]&m[785])|(~m[763]&m[764]&m[765]&m[766]&m[785]))&~BiasedRNG[706])|((m[763]&m[764]&~m[765]&~m[766]&~m[785])|(m[763]&~m[764]&m[765]&~m[766]&~m[785])|(~m[763]&m[764]&m[765]&~m[766]&~m[785])|(m[763]&m[764]&m[765]&~m[766]&~m[785])|(m[763]&m[764]&m[765]&m[766]&~m[785])|(m[763]&m[764]&~m[765]&~m[766]&m[785])|(m[763]&~m[764]&m[765]&~m[766]&m[785])|(~m[763]&m[764]&m[765]&~m[766]&m[785])|(m[763]&m[764]&m[765]&~m[766]&m[785])|(m[763]&m[764]&m[765]&m[766]&m[785]));
    m[772] = (((m[768]&~m[769]&~m[770]&~m[771]&~m[790])|(~m[768]&m[769]&~m[770]&~m[771]&~m[790])|(~m[768]&~m[769]&m[770]&~m[771]&~m[790])|(m[768]&m[769]&~m[770]&m[771]&~m[790])|(m[768]&~m[769]&m[770]&m[771]&~m[790])|(~m[768]&m[769]&m[770]&m[771]&~m[790]))&BiasedRNG[707])|(((m[768]&~m[769]&~m[770]&~m[771]&m[790])|(~m[768]&m[769]&~m[770]&~m[771]&m[790])|(~m[768]&~m[769]&m[770]&~m[771]&m[790])|(m[768]&m[769]&~m[770]&m[771]&m[790])|(m[768]&~m[769]&m[770]&m[771]&m[790])|(~m[768]&m[769]&m[770]&m[771]&m[790]))&~BiasedRNG[707])|((m[768]&m[769]&~m[770]&~m[771]&~m[790])|(m[768]&~m[769]&m[770]&~m[771]&~m[790])|(~m[768]&m[769]&m[770]&~m[771]&~m[790])|(m[768]&m[769]&m[770]&~m[771]&~m[790])|(m[768]&m[769]&m[770]&m[771]&~m[790])|(m[768]&m[769]&~m[770]&~m[771]&m[790])|(m[768]&~m[769]&m[770]&~m[771]&m[790])|(~m[768]&m[769]&m[770]&~m[771]&m[790])|(m[768]&m[769]&m[770]&~m[771]&m[790])|(m[768]&m[769]&m[770]&m[771]&m[790]));
    m[777] = (((m[773]&~m[774]&~m[775]&~m[776]&~m[795])|(~m[773]&m[774]&~m[775]&~m[776]&~m[795])|(~m[773]&~m[774]&m[775]&~m[776]&~m[795])|(m[773]&m[774]&~m[775]&m[776]&~m[795])|(m[773]&~m[774]&m[775]&m[776]&~m[795])|(~m[773]&m[774]&m[775]&m[776]&~m[795]))&BiasedRNG[708])|(((m[773]&~m[774]&~m[775]&~m[776]&m[795])|(~m[773]&m[774]&~m[775]&~m[776]&m[795])|(~m[773]&~m[774]&m[775]&~m[776]&m[795])|(m[773]&m[774]&~m[775]&m[776]&m[795])|(m[773]&~m[774]&m[775]&m[776]&m[795])|(~m[773]&m[774]&m[775]&m[776]&m[795]))&~BiasedRNG[708])|((m[773]&m[774]&~m[775]&~m[776]&~m[795])|(m[773]&~m[774]&m[775]&~m[776]&~m[795])|(~m[773]&m[774]&m[775]&~m[776]&~m[795])|(m[773]&m[774]&m[775]&~m[776]&~m[795])|(m[773]&m[774]&m[775]&m[776]&~m[795])|(m[773]&m[774]&~m[775]&~m[776]&m[795])|(m[773]&~m[774]&m[775]&~m[776]&m[795])|(~m[773]&m[774]&m[775]&~m[776]&m[795])|(m[773]&m[774]&m[775]&~m[776]&m[795])|(m[773]&m[774]&m[775]&m[776]&m[795]));
    m[782] = (((m[778]&~m[779]&~m[780]&~m[781]&~m[805])|(~m[778]&m[779]&~m[780]&~m[781]&~m[805])|(~m[778]&~m[779]&m[780]&~m[781]&~m[805])|(m[778]&m[779]&~m[780]&m[781]&~m[805])|(m[778]&~m[779]&m[780]&m[781]&~m[805])|(~m[778]&m[779]&m[780]&m[781]&~m[805]))&BiasedRNG[709])|(((m[778]&~m[779]&~m[780]&~m[781]&m[805])|(~m[778]&m[779]&~m[780]&~m[781]&m[805])|(~m[778]&~m[779]&m[780]&~m[781]&m[805])|(m[778]&m[779]&~m[780]&m[781]&m[805])|(m[778]&~m[779]&m[780]&m[781]&m[805])|(~m[778]&m[779]&m[780]&m[781]&m[805]))&~BiasedRNG[709])|((m[778]&m[779]&~m[780]&~m[781]&~m[805])|(m[778]&~m[779]&m[780]&~m[781]&~m[805])|(~m[778]&m[779]&m[780]&~m[781]&~m[805])|(m[778]&m[779]&m[780]&~m[781]&~m[805])|(m[778]&m[779]&m[780]&m[781]&~m[805])|(m[778]&m[779]&~m[780]&~m[781]&m[805])|(m[778]&~m[779]&m[780]&~m[781]&m[805])|(~m[778]&m[779]&m[780]&~m[781]&m[805])|(m[778]&m[779]&m[780]&~m[781]&m[805])|(m[778]&m[779]&m[780]&m[781]&m[805]));
    m[787] = (((m[783]&~m[784]&~m[785]&~m[786]&~m[810])|(~m[783]&m[784]&~m[785]&~m[786]&~m[810])|(~m[783]&~m[784]&m[785]&~m[786]&~m[810])|(m[783]&m[784]&~m[785]&m[786]&~m[810])|(m[783]&~m[784]&m[785]&m[786]&~m[810])|(~m[783]&m[784]&m[785]&m[786]&~m[810]))&BiasedRNG[710])|(((m[783]&~m[784]&~m[785]&~m[786]&m[810])|(~m[783]&m[784]&~m[785]&~m[786]&m[810])|(~m[783]&~m[784]&m[785]&~m[786]&m[810])|(m[783]&m[784]&~m[785]&m[786]&m[810])|(m[783]&~m[784]&m[785]&m[786]&m[810])|(~m[783]&m[784]&m[785]&m[786]&m[810]))&~BiasedRNG[710])|((m[783]&m[784]&~m[785]&~m[786]&~m[810])|(m[783]&~m[784]&m[785]&~m[786]&~m[810])|(~m[783]&m[784]&m[785]&~m[786]&~m[810])|(m[783]&m[784]&m[785]&~m[786]&~m[810])|(m[783]&m[784]&m[785]&m[786]&~m[810])|(m[783]&m[784]&~m[785]&~m[786]&m[810])|(m[783]&~m[784]&m[785]&~m[786]&m[810])|(~m[783]&m[784]&m[785]&~m[786]&m[810])|(m[783]&m[784]&m[785]&~m[786]&m[810])|(m[783]&m[784]&m[785]&m[786]&m[810]));
    m[792] = (((m[788]&~m[789]&~m[790]&~m[791]&~m[815])|(~m[788]&m[789]&~m[790]&~m[791]&~m[815])|(~m[788]&~m[789]&m[790]&~m[791]&~m[815])|(m[788]&m[789]&~m[790]&m[791]&~m[815])|(m[788]&~m[789]&m[790]&m[791]&~m[815])|(~m[788]&m[789]&m[790]&m[791]&~m[815]))&BiasedRNG[711])|(((m[788]&~m[789]&~m[790]&~m[791]&m[815])|(~m[788]&m[789]&~m[790]&~m[791]&m[815])|(~m[788]&~m[789]&m[790]&~m[791]&m[815])|(m[788]&m[789]&~m[790]&m[791]&m[815])|(m[788]&~m[789]&m[790]&m[791]&m[815])|(~m[788]&m[789]&m[790]&m[791]&m[815]))&~BiasedRNG[711])|((m[788]&m[789]&~m[790]&~m[791]&~m[815])|(m[788]&~m[789]&m[790]&~m[791]&~m[815])|(~m[788]&m[789]&m[790]&~m[791]&~m[815])|(m[788]&m[789]&m[790]&~m[791]&~m[815])|(m[788]&m[789]&m[790]&m[791]&~m[815])|(m[788]&m[789]&~m[790]&~m[791]&m[815])|(m[788]&~m[789]&m[790]&~m[791]&m[815])|(~m[788]&m[789]&m[790]&~m[791]&m[815])|(m[788]&m[789]&m[790]&~m[791]&m[815])|(m[788]&m[789]&m[790]&m[791]&m[815]));
    m[797] = (((m[793]&~m[794]&~m[795]&~m[796]&~m[820])|(~m[793]&m[794]&~m[795]&~m[796]&~m[820])|(~m[793]&~m[794]&m[795]&~m[796]&~m[820])|(m[793]&m[794]&~m[795]&m[796]&~m[820])|(m[793]&~m[794]&m[795]&m[796]&~m[820])|(~m[793]&m[794]&m[795]&m[796]&~m[820]))&BiasedRNG[712])|(((m[793]&~m[794]&~m[795]&~m[796]&m[820])|(~m[793]&m[794]&~m[795]&~m[796]&m[820])|(~m[793]&~m[794]&m[795]&~m[796]&m[820])|(m[793]&m[794]&~m[795]&m[796]&m[820])|(m[793]&~m[794]&m[795]&m[796]&m[820])|(~m[793]&m[794]&m[795]&m[796]&m[820]))&~BiasedRNG[712])|((m[793]&m[794]&~m[795]&~m[796]&~m[820])|(m[793]&~m[794]&m[795]&~m[796]&~m[820])|(~m[793]&m[794]&m[795]&~m[796]&~m[820])|(m[793]&m[794]&m[795]&~m[796]&~m[820])|(m[793]&m[794]&m[795]&m[796]&~m[820])|(m[793]&m[794]&~m[795]&~m[796]&m[820])|(m[793]&~m[794]&m[795]&~m[796]&m[820])|(~m[793]&m[794]&m[795]&~m[796]&m[820])|(m[793]&m[794]&m[795]&~m[796]&m[820])|(m[793]&m[794]&m[795]&m[796]&m[820]));
    m[802] = (((m[798]&~m[799]&~m[800]&~m[801]&~m[825])|(~m[798]&m[799]&~m[800]&~m[801]&~m[825])|(~m[798]&~m[799]&m[800]&~m[801]&~m[825])|(m[798]&m[799]&~m[800]&m[801]&~m[825])|(m[798]&~m[799]&m[800]&m[801]&~m[825])|(~m[798]&m[799]&m[800]&m[801]&~m[825]))&BiasedRNG[713])|(((m[798]&~m[799]&~m[800]&~m[801]&m[825])|(~m[798]&m[799]&~m[800]&~m[801]&m[825])|(~m[798]&~m[799]&m[800]&~m[801]&m[825])|(m[798]&m[799]&~m[800]&m[801]&m[825])|(m[798]&~m[799]&m[800]&m[801]&m[825])|(~m[798]&m[799]&m[800]&m[801]&m[825]))&~BiasedRNG[713])|((m[798]&m[799]&~m[800]&~m[801]&~m[825])|(m[798]&~m[799]&m[800]&~m[801]&~m[825])|(~m[798]&m[799]&m[800]&~m[801]&~m[825])|(m[798]&m[799]&m[800]&~m[801]&~m[825])|(m[798]&m[799]&m[800]&m[801]&~m[825])|(m[798]&m[799]&~m[800]&~m[801]&m[825])|(m[798]&~m[799]&m[800]&~m[801]&m[825])|(~m[798]&m[799]&m[800]&~m[801]&m[825])|(m[798]&m[799]&m[800]&~m[801]&m[825])|(m[798]&m[799]&m[800]&m[801]&m[825]));
    m[807] = (((m[803]&~m[804]&~m[805]&~m[806]&~m[835])|(~m[803]&m[804]&~m[805]&~m[806]&~m[835])|(~m[803]&~m[804]&m[805]&~m[806]&~m[835])|(m[803]&m[804]&~m[805]&m[806]&~m[835])|(m[803]&~m[804]&m[805]&m[806]&~m[835])|(~m[803]&m[804]&m[805]&m[806]&~m[835]))&BiasedRNG[714])|(((m[803]&~m[804]&~m[805]&~m[806]&m[835])|(~m[803]&m[804]&~m[805]&~m[806]&m[835])|(~m[803]&~m[804]&m[805]&~m[806]&m[835])|(m[803]&m[804]&~m[805]&m[806]&m[835])|(m[803]&~m[804]&m[805]&m[806]&m[835])|(~m[803]&m[804]&m[805]&m[806]&m[835]))&~BiasedRNG[714])|((m[803]&m[804]&~m[805]&~m[806]&~m[835])|(m[803]&~m[804]&m[805]&~m[806]&~m[835])|(~m[803]&m[804]&m[805]&~m[806]&~m[835])|(m[803]&m[804]&m[805]&~m[806]&~m[835])|(m[803]&m[804]&m[805]&m[806]&~m[835])|(m[803]&m[804]&~m[805]&~m[806]&m[835])|(m[803]&~m[804]&m[805]&~m[806]&m[835])|(~m[803]&m[804]&m[805]&~m[806]&m[835])|(m[803]&m[804]&m[805]&~m[806]&m[835])|(m[803]&m[804]&m[805]&m[806]&m[835]));
    m[812] = (((m[808]&~m[809]&~m[810]&~m[811]&~m[840])|(~m[808]&m[809]&~m[810]&~m[811]&~m[840])|(~m[808]&~m[809]&m[810]&~m[811]&~m[840])|(m[808]&m[809]&~m[810]&m[811]&~m[840])|(m[808]&~m[809]&m[810]&m[811]&~m[840])|(~m[808]&m[809]&m[810]&m[811]&~m[840]))&BiasedRNG[715])|(((m[808]&~m[809]&~m[810]&~m[811]&m[840])|(~m[808]&m[809]&~m[810]&~m[811]&m[840])|(~m[808]&~m[809]&m[810]&~m[811]&m[840])|(m[808]&m[809]&~m[810]&m[811]&m[840])|(m[808]&~m[809]&m[810]&m[811]&m[840])|(~m[808]&m[809]&m[810]&m[811]&m[840]))&~BiasedRNG[715])|((m[808]&m[809]&~m[810]&~m[811]&~m[840])|(m[808]&~m[809]&m[810]&~m[811]&~m[840])|(~m[808]&m[809]&m[810]&~m[811]&~m[840])|(m[808]&m[809]&m[810]&~m[811]&~m[840])|(m[808]&m[809]&m[810]&m[811]&~m[840])|(m[808]&m[809]&~m[810]&~m[811]&m[840])|(m[808]&~m[809]&m[810]&~m[811]&m[840])|(~m[808]&m[809]&m[810]&~m[811]&m[840])|(m[808]&m[809]&m[810]&~m[811]&m[840])|(m[808]&m[809]&m[810]&m[811]&m[840]));
    m[817] = (((m[813]&~m[814]&~m[815]&~m[816]&~m[845])|(~m[813]&m[814]&~m[815]&~m[816]&~m[845])|(~m[813]&~m[814]&m[815]&~m[816]&~m[845])|(m[813]&m[814]&~m[815]&m[816]&~m[845])|(m[813]&~m[814]&m[815]&m[816]&~m[845])|(~m[813]&m[814]&m[815]&m[816]&~m[845]))&BiasedRNG[716])|(((m[813]&~m[814]&~m[815]&~m[816]&m[845])|(~m[813]&m[814]&~m[815]&~m[816]&m[845])|(~m[813]&~m[814]&m[815]&~m[816]&m[845])|(m[813]&m[814]&~m[815]&m[816]&m[845])|(m[813]&~m[814]&m[815]&m[816]&m[845])|(~m[813]&m[814]&m[815]&m[816]&m[845]))&~BiasedRNG[716])|((m[813]&m[814]&~m[815]&~m[816]&~m[845])|(m[813]&~m[814]&m[815]&~m[816]&~m[845])|(~m[813]&m[814]&m[815]&~m[816]&~m[845])|(m[813]&m[814]&m[815]&~m[816]&~m[845])|(m[813]&m[814]&m[815]&m[816]&~m[845])|(m[813]&m[814]&~m[815]&~m[816]&m[845])|(m[813]&~m[814]&m[815]&~m[816]&m[845])|(~m[813]&m[814]&m[815]&~m[816]&m[845])|(m[813]&m[814]&m[815]&~m[816]&m[845])|(m[813]&m[814]&m[815]&m[816]&m[845]));
    m[822] = (((m[818]&~m[819]&~m[820]&~m[821]&~m[850])|(~m[818]&m[819]&~m[820]&~m[821]&~m[850])|(~m[818]&~m[819]&m[820]&~m[821]&~m[850])|(m[818]&m[819]&~m[820]&m[821]&~m[850])|(m[818]&~m[819]&m[820]&m[821]&~m[850])|(~m[818]&m[819]&m[820]&m[821]&~m[850]))&BiasedRNG[717])|(((m[818]&~m[819]&~m[820]&~m[821]&m[850])|(~m[818]&m[819]&~m[820]&~m[821]&m[850])|(~m[818]&~m[819]&m[820]&~m[821]&m[850])|(m[818]&m[819]&~m[820]&m[821]&m[850])|(m[818]&~m[819]&m[820]&m[821]&m[850])|(~m[818]&m[819]&m[820]&m[821]&m[850]))&~BiasedRNG[717])|((m[818]&m[819]&~m[820]&~m[821]&~m[850])|(m[818]&~m[819]&m[820]&~m[821]&~m[850])|(~m[818]&m[819]&m[820]&~m[821]&~m[850])|(m[818]&m[819]&m[820]&~m[821]&~m[850])|(m[818]&m[819]&m[820]&m[821]&~m[850])|(m[818]&m[819]&~m[820]&~m[821]&m[850])|(m[818]&~m[819]&m[820]&~m[821]&m[850])|(~m[818]&m[819]&m[820]&~m[821]&m[850])|(m[818]&m[819]&m[820]&~m[821]&m[850])|(m[818]&m[819]&m[820]&m[821]&m[850]));
    m[827] = (((m[823]&~m[824]&~m[825]&~m[826]&~m[855])|(~m[823]&m[824]&~m[825]&~m[826]&~m[855])|(~m[823]&~m[824]&m[825]&~m[826]&~m[855])|(m[823]&m[824]&~m[825]&m[826]&~m[855])|(m[823]&~m[824]&m[825]&m[826]&~m[855])|(~m[823]&m[824]&m[825]&m[826]&~m[855]))&BiasedRNG[718])|(((m[823]&~m[824]&~m[825]&~m[826]&m[855])|(~m[823]&m[824]&~m[825]&~m[826]&m[855])|(~m[823]&~m[824]&m[825]&~m[826]&m[855])|(m[823]&m[824]&~m[825]&m[826]&m[855])|(m[823]&~m[824]&m[825]&m[826]&m[855])|(~m[823]&m[824]&m[825]&m[826]&m[855]))&~BiasedRNG[718])|((m[823]&m[824]&~m[825]&~m[826]&~m[855])|(m[823]&~m[824]&m[825]&~m[826]&~m[855])|(~m[823]&m[824]&m[825]&~m[826]&~m[855])|(m[823]&m[824]&m[825]&~m[826]&~m[855])|(m[823]&m[824]&m[825]&m[826]&~m[855])|(m[823]&m[824]&~m[825]&~m[826]&m[855])|(m[823]&~m[824]&m[825]&~m[826]&m[855])|(~m[823]&m[824]&m[825]&~m[826]&m[855])|(m[823]&m[824]&m[825]&~m[826]&m[855])|(m[823]&m[824]&m[825]&m[826]&m[855]));
    m[832] = (((m[828]&~m[829]&~m[830]&~m[831]&~m[860])|(~m[828]&m[829]&~m[830]&~m[831]&~m[860])|(~m[828]&~m[829]&m[830]&~m[831]&~m[860])|(m[828]&m[829]&~m[830]&m[831]&~m[860])|(m[828]&~m[829]&m[830]&m[831]&~m[860])|(~m[828]&m[829]&m[830]&m[831]&~m[860]))&BiasedRNG[719])|(((m[828]&~m[829]&~m[830]&~m[831]&m[860])|(~m[828]&m[829]&~m[830]&~m[831]&m[860])|(~m[828]&~m[829]&m[830]&~m[831]&m[860])|(m[828]&m[829]&~m[830]&m[831]&m[860])|(m[828]&~m[829]&m[830]&m[831]&m[860])|(~m[828]&m[829]&m[830]&m[831]&m[860]))&~BiasedRNG[719])|((m[828]&m[829]&~m[830]&~m[831]&~m[860])|(m[828]&~m[829]&m[830]&~m[831]&~m[860])|(~m[828]&m[829]&m[830]&~m[831]&~m[860])|(m[828]&m[829]&m[830]&~m[831]&~m[860])|(m[828]&m[829]&m[830]&m[831]&~m[860])|(m[828]&m[829]&~m[830]&~m[831]&m[860])|(m[828]&~m[829]&m[830]&~m[831]&m[860])|(~m[828]&m[829]&m[830]&~m[831]&m[860])|(m[828]&m[829]&m[830]&~m[831]&m[860])|(m[828]&m[829]&m[830]&m[831]&m[860]));
    m[837] = (((m[833]&~m[834]&~m[835]&~m[836]&~m[870])|(~m[833]&m[834]&~m[835]&~m[836]&~m[870])|(~m[833]&~m[834]&m[835]&~m[836]&~m[870])|(m[833]&m[834]&~m[835]&m[836]&~m[870])|(m[833]&~m[834]&m[835]&m[836]&~m[870])|(~m[833]&m[834]&m[835]&m[836]&~m[870]))&BiasedRNG[720])|(((m[833]&~m[834]&~m[835]&~m[836]&m[870])|(~m[833]&m[834]&~m[835]&~m[836]&m[870])|(~m[833]&~m[834]&m[835]&~m[836]&m[870])|(m[833]&m[834]&~m[835]&m[836]&m[870])|(m[833]&~m[834]&m[835]&m[836]&m[870])|(~m[833]&m[834]&m[835]&m[836]&m[870]))&~BiasedRNG[720])|((m[833]&m[834]&~m[835]&~m[836]&~m[870])|(m[833]&~m[834]&m[835]&~m[836]&~m[870])|(~m[833]&m[834]&m[835]&~m[836]&~m[870])|(m[833]&m[834]&m[835]&~m[836]&~m[870])|(m[833]&m[834]&m[835]&m[836]&~m[870])|(m[833]&m[834]&~m[835]&~m[836]&m[870])|(m[833]&~m[834]&m[835]&~m[836]&m[870])|(~m[833]&m[834]&m[835]&~m[836]&m[870])|(m[833]&m[834]&m[835]&~m[836]&m[870])|(m[833]&m[834]&m[835]&m[836]&m[870]));
    m[842] = (((m[838]&~m[839]&~m[840]&~m[841]&~m[875])|(~m[838]&m[839]&~m[840]&~m[841]&~m[875])|(~m[838]&~m[839]&m[840]&~m[841]&~m[875])|(m[838]&m[839]&~m[840]&m[841]&~m[875])|(m[838]&~m[839]&m[840]&m[841]&~m[875])|(~m[838]&m[839]&m[840]&m[841]&~m[875]))&BiasedRNG[721])|(((m[838]&~m[839]&~m[840]&~m[841]&m[875])|(~m[838]&m[839]&~m[840]&~m[841]&m[875])|(~m[838]&~m[839]&m[840]&~m[841]&m[875])|(m[838]&m[839]&~m[840]&m[841]&m[875])|(m[838]&~m[839]&m[840]&m[841]&m[875])|(~m[838]&m[839]&m[840]&m[841]&m[875]))&~BiasedRNG[721])|((m[838]&m[839]&~m[840]&~m[841]&~m[875])|(m[838]&~m[839]&m[840]&~m[841]&~m[875])|(~m[838]&m[839]&m[840]&~m[841]&~m[875])|(m[838]&m[839]&m[840]&~m[841]&~m[875])|(m[838]&m[839]&m[840]&m[841]&~m[875])|(m[838]&m[839]&~m[840]&~m[841]&m[875])|(m[838]&~m[839]&m[840]&~m[841]&m[875])|(~m[838]&m[839]&m[840]&~m[841]&m[875])|(m[838]&m[839]&m[840]&~m[841]&m[875])|(m[838]&m[839]&m[840]&m[841]&m[875]));
    m[847] = (((m[843]&~m[844]&~m[845]&~m[846]&~m[880])|(~m[843]&m[844]&~m[845]&~m[846]&~m[880])|(~m[843]&~m[844]&m[845]&~m[846]&~m[880])|(m[843]&m[844]&~m[845]&m[846]&~m[880])|(m[843]&~m[844]&m[845]&m[846]&~m[880])|(~m[843]&m[844]&m[845]&m[846]&~m[880]))&BiasedRNG[722])|(((m[843]&~m[844]&~m[845]&~m[846]&m[880])|(~m[843]&m[844]&~m[845]&~m[846]&m[880])|(~m[843]&~m[844]&m[845]&~m[846]&m[880])|(m[843]&m[844]&~m[845]&m[846]&m[880])|(m[843]&~m[844]&m[845]&m[846]&m[880])|(~m[843]&m[844]&m[845]&m[846]&m[880]))&~BiasedRNG[722])|((m[843]&m[844]&~m[845]&~m[846]&~m[880])|(m[843]&~m[844]&m[845]&~m[846]&~m[880])|(~m[843]&m[844]&m[845]&~m[846]&~m[880])|(m[843]&m[844]&m[845]&~m[846]&~m[880])|(m[843]&m[844]&m[845]&m[846]&~m[880])|(m[843]&m[844]&~m[845]&~m[846]&m[880])|(m[843]&~m[844]&m[845]&~m[846]&m[880])|(~m[843]&m[844]&m[845]&~m[846]&m[880])|(m[843]&m[844]&m[845]&~m[846]&m[880])|(m[843]&m[844]&m[845]&m[846]&m[880]));
    m[852] = (((m[848]&~m[849]&~m[850]&~m[851]&~m[885])|(~m[848]&m[849]&~m[850]&~m[851]&~m[885])|(~m[848]&~m[849]&m[850]&~m[851]&~m[885])|(m[848]&m[849]&~m[850]&m[851]&~m[885])|(m[848]&~m[849]&m[850]&m[851]&~m[885])|(~m[848]&m[849]&m[850]&m[851]&~m[885]))&BiasedRNG[723])|(((m[848]&~m[849]&~m[850]&~m[851]&m[885])|(~m[848]&m[849]&~m[850]&~m[851]&m[885])|(~m[848]&~m[849]&m[850]&~m[851]&m[885])|(m[848]&m[849]&~m[850]&m[851]&m[885])|(m[848]&~m[849]&m[850]&m[851]&m[885])|(~m[848]&m[849]&m[850]&m[851]&m[885]))&~BiasedRNG[723])|((m[848]&m[849]&~m[850]&~m[851]&~m[885])|(m[848]&~m[849]&m[850]&~m[851]&~m[885])|(~m[848]&m[849]&m[850]&~m[851]&~m[885])|(m[848]&m[849]&m[850]&~m[851]&~m[885])|(m[848]&m[849]&m[850]&m[851]&~m[885])|(m[848]&m[849]&~m[850]&~m[851]&m[885])|(m[848]&~m[849]&m[850]&~m[851]&m[885])|(~m[848]&m[849]&m[850]&~m[851]&m[885])|(m[848]&m[849]&m[850]&~m[851]&m[885])|(m[848]&m[849]&m[850]&m[851]&m[885]));
    m[857] = (((m[853]&~m[854]&~m[855]&~m[856]&~m[890])|(~m[853]&m[854]&~m[855]&~m[856]&~m[890])|(~m[853]&~m[854]&m[855]&~m[856]&~m[890])|(m[853]&m[854]&~m[855]&m[856]&~m[890])|(m[853]&~m[854]&m[855]&m[856]&~m[890])|(~m[853]&m[854]&m[855]&m[856]&~m[890]))&BiasedRNG[724])|(((m[853]&~m[854]&~m[855]&~m[856]&m[890])|(~m[853]&m[854]&~m[855]&~m[856]&m[890])|(~m[853]&~m[854]&m[855]&~m[856]&m[890])|(m[853]&m[854]&~m[855]&m[856]&m[890])|(m[853]&~m[854]&m[855]&m[856]&m[890])|(~m[853]&m[854]&m[855]&m[856]&m[890]))&~BiasedRNG[724])|((m[853]&m[854]&~m[855]&~m[856]&~m[890])|(m[853]&~m[854]&m[855]&~m[856]&~m[890])|(~m[853]&m[854]&m[855]&~m[856]&~m[890])|(m[853]&m[854]&m[855]&~m[856]&~m[890])|(m[853]&m[854]&m[855]&m[856]&~m[890])|(m[853]&m[854]&~m[855]&~m[856]&m[890])|(m[853]&~m[854]&m[855]&~m[856]&m[890])|(~m[853]&m[854]&m[855]&~m[856]&m[890])|(m[853]&m[854]&m[855]&~m[856]&m[890])|(m[853]&m[854]&m[855]&m[856]&m[890]));
    m[862] = (((m[858]&~m[859]&~m[860]&~m[861]&~m[895])|(~m[858]&m[859]&~m[860]&~m[861]&~m[895])|(~m[858]&~m[859]&m[860]&~m[861]&~m[895])|(m[858]&m[859]&~m[860]&m[861]&~m[895])|(m[858]&~m[859]&m[860]&m[861]&~m[895])|(~m[858]&m[859]&m[860]&m[861]&~m[895]))&BiasedRNG[725])|(((m[858]&~m[859]&~m[860]&~m[861]&m[895])|(~m[858]&m[859]&~m[860]&~m[861]&m[895])|(~m[858]&~m[859]&m[860]&~m[861]&m[895])|(m[858]&m[859]&~m[860]&m[861]&m[895])|(m[858]&~m[859]&m[860]&m[861]&m[895])|(~m[858]&m[859]&m[860]&m[861]&m[895]))&~BiasedRNG[725])|((m[858]&m[859]&~m[860]&~m[861]&~m[895])|(m[858]&~m[859]&m[860]&~m[861]&~m[895])|(~m[858]&m[859]&m[860]&~m[861]&~m[895])|(m[858]&m[859]&m[860]&~m[861]&~m[895])|(m[858]&m[859]&m[860]&m[861]&~m[895])|(m[858]&m[859]&~m[860]&~m[861]&m[895])|(m[858]&~m[859]&m[860]&~m[861]&m[895])|(~m[858]&m[859]&m[860]&~m[861]&m[895])|(m[858]&m[859]&m[860]&~m[861]&m[895])|(m[858]&m[859]&m[860]&m[861]&m[895]));
    m[867] = (((m[863]&~m[864]&~m[865]&~m[866]&~m[900])|(~m[863]&m[864]&~m[865]&~m[866]&~m[900])|(~m[863]&~m[864]&m[865]&~m[866]&~m[900])|(m[863]&m[864]&~m[865]&m[866]&~m[900])|(m[863]&~m[864]&m[865]&m[866]&~m[900])|(~m[863]&m[864]&m[865]&m[866]&~m[900]))&BiasedRNG[726])|(((m[863]&~m[864]&~m[865]&~m[866]&m[900])|(~m[863]&m[864]&~m[865]&~m[866]&m[900])|(~m[863]&~m[864]&m[865]&~m[866]&m[900])|(m[863]&m[864]&~m[865]&m[866]&m[900])|(m[863]&~m[864]&m[865]&m[866]&m[900])|(~m[863]&m[864]&m[865]&m[866]&m[900]))&~BiasedRNG[726])|((m[863]&m[864]&~m[865]&~m[866]&~m[900])|(m[863]&~m[864]&m[865]&~m[866]&~m[900])|(~m[863]&m[864]&m[865]&~m[866]&~m[900])|(m[863]&m[864]&m[865]&~m[866]&~m[900])|(m[863]&m[864]&m[865]&m[866]&~m[900])|(m[863]&m[864]&~m[865]&~m[866]&m[900])|(m[863]&~m[864]&m[865]&~m[866]&m[900])|(~m[863]&m[864]&m[865]&~m[866]&m[900])|(m[863]&m[864]&m[865]&~m[866]&m[900])|(m[863]&m[864]&m[865]&m[866]&m[900]));
    m[872] = (((m[868]&~m[869]&~m[870]&~m[871]&~m[910])|(~m[868]&m[869]&~m[870]&~m[871]&~m[910])|(~m[868]&~m[869]&m[870]&~m[871]&~m[910])|(m[868]&m[869]&~m[870]&m[871]&~m[910])|(m[868]&~m[869]&m[870]&m[871]&~m[910])|(~m[868]&m[869]&m[870]&m[871]&~m[910]))&BiasedRNG[727])|(((m[868]&~m[869]&~m[870]&~m[871]&m[910])|(~m[868]&m[869]&~m[870]&~m[871]&m[910])|(~m[868]&~m[869]&m[870]&~m[871]&m[910])|(m[868]&m[869]&~m[870]&m[871]&m[910])|(m[868]&~m[869]&m[870]&m[871]&m[910])|(~m[868]&m[869]&m[870]&m[871]&m[910]))&~BiasedRNG[727])|((m[868]&m[869]&~m[870]&~m[871]&~m[910])|(m[868]&~m[869]&m[870]&~m[871]&~m[910])|(~m[868]&m[869]&m[870]&~m[871]&~m[910])|(m[868]&m[869]&m[870]&~m[871]&~m[910])|(m[868]&m[869]&m[870]&m[871]&~m[910])|(m[868]&m[869]&~m[870]&~m[871]&m[910])|(m[868]&~m[869]&m[870]&~m[871]&m[910])|(~m[868]&m[869]&m[870]&~m[871]&m[910])|(m[868]&m[869]&m[870]&~m[871]&m[910])|(m[868]&m[869]&m[870]&m[871]&m[910]));
    m[877] = (((m[873]&~m[874]&~m[875]&~m[876]&~m[915])|(~m[873]&m[874]&~m[875]&~m[876]&~m[915])|(~m[873]&~m[874]&m[875]&~m[876]&~m[915])|(m[873]&m[874]&~m[875]&m[876]&~m[915])|(m[873]&~m[874]&m[875]&m[876]&~m[915])|(~m[873]&m[874]&m[875]&m[876]&~m[915]))&BiasedRNG[728])|(((m[873]&~m[874]&~m[875]&~m[876]&m[915])|(~m[873]&m[874]&~m[875]&~m[876]&m[915])|(~m[873]&~m[874]&m[875]&~m[876]&m[915])|(m[873]&m[874]&~m[875]&m[876]&m[915])|(m[873]&~m[874]&m[875]&m[876]&m[915])|(~m[873]&m[874]&m[875]&m[876]&m[915]))&~BiasedRNG[728])|((m[873]&m[874]&~m[875]&~m[876]&~m[915])|(m[873]&~m[874]&m[875]&~m[876]&~m[915])|(~m[873]&m[874]&m[875]&~m[876]&~m[915])|(m[873]&m[874]&m[875]&~m[876]&~m[915])|(m[873]&m[874]&m[875]&m[876]&~m[915])|(m[873]&m[874]&~m[875]&~m[876]&m[915])|(m[873]&~m[874]&m[875]&~m[876]&m[915])|(~m[873]&m[874]&m[875]&~m[876]&m[915])|(m[873]&m[874]&m[875]&~m[876]&m[915])|(m[873]&m[874]&m[875]&m[876]&m[915]));
    m[882] = (((m[878]&~m[879]&~m[880]&~m[881]&~m[920])|(~m[878]&m[879]&~m[880]&~m[881]&~m[920])|(~m[878]&~m[879]&m[880]&~m[881]&~m[920])|(m[878]&m[879]&~m[880]&m[881]&~m[920])|(m[878]&~m[879]&m[880]&m[881]&~m[920])|(~m[878]&m[879]&m[880]&m[881]&~m[920]))&BiasedRNG[729])|(((m[878]&~m[879]&~m[880]&~m[881]&m[920])|(~m[878]&m[879]&~m[880]&~m[881]&m[920])|(~m[878]&~m[879]&m[880]&~m[881]&m[920])|(m[878]&m[879]&~m[880]&m[881]&m[920])|(m[878]&~m[879]&m[880]&m[881]&m[920])|(~m[878]&m[879]&m[880]&m[881]&m[920]))&~BiasedRNG[729])|((m[878]&m[879]&~m[880]&~m[881]&~m[920])|(m[878]&~m[879]&m[880]&~m[881]&~m[920])|(~m[878]&m[879]&m[880]&~m[881]&~m[920])|(m[878]&m[879]&m[880]&~m[881]&~m[920])|(m[878]&m[879]&m[880]&m[881]&~m[920])|(m[878]&m[879]&~m[880]&~m[881]&m[920])|(m[878]&~m[879]&m[880]&~m[881]&m[920])|(~m[878]&m[879]&m[880]&~m[881]&m[920])|(m[878]&m[879]&m[880]&~m[881]&m[920])|(m[878]&m[879]&m[880]&m[881]&m[920]));
    m[887] = (((m[883]&~m[884]&~m[885]&~m[886]&~m[925])|(~m[883]&m[884]&~m[885]&~m[886]&~m[925])|(~m[883]&~m[884]&m[885]&~m[886]&~m[925])|(m[883]&m[884]&~m[885]&m[886]&~m[925])|(m[883]&~m[884]&m[885]&m[886]&~m[925])|(~m[883]&m[884]&m[885]&m[886]&~m[925]))&BiasedRNG[730])|(((m[883]&~m[884]&~m[885]&~m[886]&m[925])|(~m[883]&m[884]&~m[885]&~m[886]&m[925])|(~m[883]&~m[884]&m[885]&~m[886]&m[925])|(m[883]&m[884]&~m[885]&m[886]&m[925])|(m[883]&~m[884]&m[885]&m[886]&m[925])|(~m[883]&m[884]&m[885]&m[886]&m[925]))&~BiasedRNG[730])|((m[883]&m[884]&~m[885]&~m[886]&~m[925])|(m[883]&~m[884]&m[885]&~m[886]&~m[925])|(~m[883]&m[884]&m[885]&~m[886]&~m[925])|(m[883]&m[884]&m[885]&~m[886]&~m[925])|(m[883]&m[884]&m[885]&m[886]&~m[925])|(m[883]&m[884]&~m[885]&~m[886]&m[925])|(m[883]&~m[884]&m[885]&~m[886]&m[925])|(~m[883]&m[884]&m[885]&~m[886]&m[925])|(m[883]&m[884]&m[885]&~m[886]&m[925])|(m[883]&m[884]&m[885]&m[886]&m[925]));
    m[892] = (((m[888]&~m[889]&~m[890]&~m[891]&~m[930])|(~m[888]&m[889]&~m[890]&~m[891]&~m[930])|(~m[888]&~m[889]&m[890]&~m[891]&~m[930])|(m[888]&m[889]&~m[890]&m[891]&~m[930])|(m[888]&~m[889]&m[890]&m[891]&~m[930])|(~m[888]&m[889]&m[890]&m[891]&~m[930]))&BiasedRNG[731])|(((m[888]&~m[889]&~m[890]&~m[891]&m[930])|(~m[888]&m[889]&~m[890]&~m[891]&m[930])|(~m[888]&~m[889]&m[890]&~m[891]&m[930])|(m[888]&m[889]&~m[890]&m[891]&m[930])|(m[888]&~m[889]&m[890]&m[891]&m[930])|(~m[888]&m[889]&m[890]&m[891]&m[930]))&~BiasedRNG[731])|((m[888]&m[889]&~m[890]&~m[891]&~m[930])|(m[888]&~m[889]&m[890]&~m[891]&~m[930])|(~m[888]&m[889]&m[890]&~m[891]&~m[930])|(m[888]&m[889]&m[890]&~m[891]&~m[930])|(m[888]&m[889]&m[890]&m[891]&~m[930])|(m[888]&m[889]&~m[890]&~m[891]&m[930])|(m[888]&~m[889]&m[890]&~m[891]&m[930])|(~m[888]&m[889]&m[890]&~m[891]&m[930])|(m[888]&m[889]&m[890]&~m[891]&m[930])|(m[888]&m[889]&m[890]&m[891]&m[930]));
    m[897] = (((m[893]&~m[894]&~m[895]&~m[896]&~m[935])|(~m[893]&m[894]&~m[895]&~m[896]&~m[935])|(~m[893]&~m[894]&m[895]&~m[896]&~m[935])|(m[893]&m[894]&~m[895]&m[896]&~m[935])|(m[893]&~m[894]&m[895]&m[896]&~m[935])|(~m[893]&m[894]&m[895]&m[896]&~m[935]))&BiasedRNG[732])|(((m[893]&~m[894]&~m[895]&~m[896]&m[935])|(~m[893]&m[894]&~m[895]&~m[896]&m[935])|(~m[893]&~m[894]&m[895]&~m[896]&m[935])|(m[893]&m[894]&~m[895]&m[896]&m[935])|(m[893]&~m[894]&m[895]&m[896]&m[935])|(~m[893]&m[894]&m[895]&m[896]&m[935]))&~BiasedRNG[732])|((m[893]&m[894]&~m[895]&~m[896]&~m[935])|(m[893]&~m[894]&m[895]&~m[896]&~m[935])|(~m[893]&m[894]&m[895]&~m[896]&~m[935])|(m[893]&m[894]&m[895]&~m[896]&~m[935])|(m[893]&m[894]&m[895]&m[896]&~m[935])|(m[893]&m[894]&~m[895]&~m[896]&m[935])|(m[893]&~m[894]&m[895]&~m[896]&m[935])|(~m[893]&m[894]&m[895]&~m[896]&m[935])|(m[893]&m[894]&m[895]&~m[896]&m[935])|(m[893]&m[894]&m[895]&m[896]&m[935]));
    m[902] = (((m[898]&~m[899]&~m[900]&~m[901]&~m[940])|(~m[898]&m[899]&~m[900]&~m[901]&~m[940])|(~m[898]&~m[899]&m[900]&~m[901]&~m[940])|(m[898]&m[899]&~m[900]&m[901]&~m[940])|(m[898]&~m[899]&m[900]&m[901]&~m[940])|(~m[898]&m[899]&m[900]&m[901]&~m[940]))&BiasedRNG[733])|(((m[898]&~m[899]&~m[900]&~m[901]&m[940])|(~m[898]&m[899]&~m[900]&~m[901]&m[940])|(~m[898]&~m[899]&m[900]&~m[901]&m[940])|(m[898]&m[899]&~m[900]&m[901]&m[940])|(m[898]&~m[899]&m[900]&m[901]&m[940])|(~m[898]&m[899]&m[900]&m[901]&m[940]))&~BiasedRNG[733])|((m[898]&m[899]&~m[900]&~m[901]&~m[940])|(m[898]&~m[899]&m[900]&~m[901]&~m[940])|(~m[898]&m[899]&m[900]&~m[901]&~m[940])|(m[898]&m[899]&m[900]&~m[901]&~m[940])|(m[898]&m[899]&m[900]&m[901]&~m[940])|(m[898]&m[899]&~m[900]&~m[901]&m[940])|(m[898]&~m[899]&m[900]&~m[901]&m[940])|(~m[898]&m[899]&m[900]&~m[901]&m[940])|(m[898]&m[899]&m[900]&~m[901]&m[940])|(m[898]&m[899]&m[900]&m[901]&m[940]));
    m[907] = (((m[903]&~m[904]&~m[905]&~m[906]&~m[945])|(~m[903]&m[904]&~m[905]&~m[906]&~m[945])|(~m[903]&~m[904]&m[905]&~m[906]&~m[945])|(m[903]&m[904]&~m[905]&m[906]&~m[945])|(m[903]&~m[904]&m[905]&m[906]&~m[945])|(~m[903]&m[904]&m[905]&m[906]&~m[945]))&BiasedRNG[734])|(((m[903]&~m[904]&~m[905]&~m[906]&m[945])|(~m[903]&m[904]&~m[905]&~m[906]&m[945])|(~m[903]&~m[904]&m[905]&~m[906]&m[945])|(m[903]&m[904]&~m[905]&m[906]&m[945])|(m[903]&~m[904]&m[905]&m[906]&m[945])|(~m[903]&m[904]&m[905]&m[906]&m[945]))&~BiasedRNG[734])|((m[903]&m[904]&~m[905]&~m[906]&~m[945])|(m[903]&~m[904]&m[905]&~m[906]&~m[945])|(~m[903]&m[904]&m[905]&~m[906]&~m[945])|(m[903]&m[904]&m[905]&~m[906]&~m[945])|(m[903]&m[904]&m[905]&m[906]&~m[945])|(m[903]&m[904]&~m[905]&~m[906]&m[945])|(m[903]&~m[904]&m[905]&~m[906]&m[945])|(~m[903]&m[904]&m[905]&~m[906]&m[945])|(m[903]&m[904]&m[905]&~m[906]&m[945])|(m[903]&m[904]&m[905]&m[906]&m[945]));
    m[912] = (((m[908]&~m[909]&~m[910]&~m[911]&~m[955])|(~m[908]&m[909]&~m[910]&~m[911]&~m[955])|(~m[908]&~m[909]&m[910]&~m[911]&~m[955])|(m[908]&m[909]&~m[910]&m[911]&~m[955])|(m[908]&~m[909]&m[910]&m[911]&~m[955])|(~m[908]&m[909]&m[910]&m[911]&~m[955]))&BiasedRNG[735])|(((m[908]&~m[909]&~m[910]&~m[911]&m[955])|(~m[908]&m[909]&~m[910]&~m[911]&m[955])|(~m[908]&~m[909]&m[910]&~m[911]&m[955])|(m[908]&m[909]&~m[910]&m[911]&m[955])|(m[908]&~m[909]&m[910]&m[911]&m[955])|(~m[908]&m[909]&m[910]&m[911]&m[955]))&~BiasedRNG[735])|((m[908]&m[909]&~m[910]&~m[911]&~m[955])|(m[908]&~m[909]&m[910]&~m[911]&~m[955])|(~m[908]&m[909]&m[910]&~m[911]&~m[955])|(m[908]&m[909]&m[910]&~m[911]&~m[955])|(m[908]&m[909]&m[910]&m[911]&~m[955])|(m[908]&m[909]&~m[910]&~m[911]&m[955])|(m[908]&~m[909]&m[910]&~m[911]&m[955])|(~m[908]&m[909]&m[910]&~m[911]&m[955])|(m[908]&m[909]&m[910]&~m[911]&m[955])|(m[908]&m[909]&m[910]&m[911]&m[955]));
    m[917] = (((m[913]&~m[914]&~m[915]&~m[916]&~m[960])|(~m[913]&m[914]&~m[915]&~m[916]&~m[960])|(~m[913]&~m[914]&m[915]&~m[916]&~m[960])|(m[913]&m[914]&~m[915]&m[916]&~m[960])|(m[913]&~m[914]&m[915]&m[916]&~m[960])|(~m[913]&m[914]&m[915]&m[916]&~m[960]))&BiasedRNG[736])|(((m[913]&~m[914]&~m[915]&~m[916]&m[960])|(~m[913]&m[914]&~m[915]&~m[916]&m[960])|(~m[913]&~m[914]&m[915]&~m[916]&m[960])|(m[913]&m[914]&~m[915]&m[916]&m[960])|(m[913]&~m[914]&m[915]&m[916]&m[960])|(~m[913]&m[914]&m[915]&m[916]&m[960]))&~BiasedRNG[736])|((m[913]&m[914]&~m[915]&~m[916]&~m[960])|(m[913]&~m[914]&m[915]&~m[916]&~m[960])|(~m[913]&m[914]&m[915]&~m[916]&~m[960])|(m[913]&m[914]&m[915]&~m[916]&~m[960])|(m[913]&m[914]&m[915]&m[916]&~m[960])|(m[913]&m[914]&~m[915]&~m[916]&m[960])|(m[913]&~m[914]&m[915]&~m[916]&m[960])|(~m[913]&m[914]&m[915]&~m[916]&m[960])|(m[913]&m[914]&m[915]&~m[916]&m[960])|(m[913]&m[914]&m[915]&m[916]&m[960]));
    m[922] = (((m[918]&~m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&m[919]&~m[920]&~m[921]&~m[965])|(~m[918]&~m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&~m[920]&m[921]&~m[965])|(m[918]&~m[919]&m[920]&m[921]&~m[965])|(~m[918]&m[919]&m[920]&m[921]&~m[965]))&BiasedRNG[737])|(((m[918]&~m[919]&~m[920]&~m[921]&m[965])|(~m[918]&m[919]&~m[920]&~m[921]&m[965])|(~m[918]&~m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&~m[920]&m[921]&m[965])|(m[918]&~m[919]&m[920]&m[921]&m[965])|(~m[918]&m[919]&m[920]&m[921]&m[965]))&~BiasedRNG[737])|((m[918]&m[919]&~m[920]&~m[921]&~m[965])|(m[918]&~m[919]&m[920]&~m[921]&~m[965])|(~m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&~m[921]&~m[965])|(m[918]&m[919]&m[920]&m[921]&~m[965])|(m[918]&m[919]&~m[920]&~m[921]&m[965])|(m[918]&~m[919]&m[920]&~m[921]&m[965])|(~m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&~m[921]&m[965])|(m[918]&m[919]&m[920]&m[921]&m[965]));
    m[927] = (((m[923]&~m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&m[924]&~m[925]&~m[926]&~m[970])|(~m[923]&~m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&~m[925]&m[926]&~m[970])|(m[923]&~m[924]&m[925]&m[926]&~m[970])|(~m[923]&m[924]&m[925]&m[926]&~m[970]))&BiasedRNG[738])|(((m[923]&~m[924]&~m[925]&~m[926]&m[970])|(~m[923]&m[924]&~m[925]&~m[926]&m[970])|(~m[923]&~m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&~m[925]&m[926]&m[970])|(m[923]&~m[924]&m[925]&m[926]&m[970])|(~m[923]&m[924]&m[925]&m[926]&m[970]))&~BiasedRNG[738])|((m[923]&m[924]&~m[925]&~m[926]&~m[970])|(m[923]&~m[924]&m[925]&~m[926]&~m[970])|(~m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&~m[926]&~m[970])|(m[923]&m[924]&m[925]&m[926]&~m[970])|(m[923]&m[924]&~m[925]&~m[926]&m[970])|(m[923]&~m[924]&m[925]&~m[926]&m[970])|(~m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&~m[926]&m[970])|(m[923]&m[924]&m[925]&m[926]&m[970]));
    m[932] = (((m[928]&~m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&m[929]&~m[930]&~m[931]&~m[975])|(~m[928]&~m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&~m[930]&m[931]&~m[975])|(m[928]&~m[929]&m[930]&m[931]&~m[975])|(~m[928]&m[929]&m[930]&m[931]&~m[975]))&BiasedRNG[739])|(((m[928]&~m[929]&~m[930]&~m[931]&m[975])|(~m[928]&m[929]&~m[930]&~m[931]&m[975])|(~m[928]&~m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&~m[930]&m[931]&m[975])|(m[928]&~m[929]&m[930]&m[931]&m[975])|(~m[928]&m[929]&m[930]&m[931]&m[975]))&~BiasedRNG[739])|((m[928]&m[929]&~m[930]&~m[931]&~m[975])|(m[928]&~m[929]&m[930]&~m[931]&~m[975])|(~m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&~m[931]&~m[975])|(m[928]&m[929]&m[930]&m[931]&~m[975])|(m[928]&m[929]&~m[930]&~m[931]&m[975])|(m[928]&~m[929]&m[930]&~m[931]&m[975])|(~m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&~m[931]&m[975])|(m[928]&m[929]&m[930]&m[931]&m[975]));
    m[937] = (((m[933]&~m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&m[934]&~m[935]&~m[936]&~m[980])|(~m[933]&~m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&~m[935]&m[936]&~m[980])|(m[933]&~m[934]&m[935]&m[936]&~m[980])|(~m[933]&m[934]&m[935]&m[936]&~m[980]))&BiasedRNG[740])|(((m[933]&~m[934]&~m[935]&~m[936]&m[980])|(~m[933]&m[934]&~m[935]&~m[936]&m[980])|(~m[933]&~m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&~m[935]&m[936]&m[980])|(m[933]&~m[934]&m[935]&m[936]&m[980])|(~m[933]&m[934]&m[935]&m[936]&m[980]))&~BiasedRNG[740])|((m[933]&m[934]&~m[935]&~m[936]&~m[980])|(m[933]&~m[934]&m[935]&~m[936]&~m[980])|(~m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&~m[936]&~m[980])|(m[933]&m[934]&m[935]&m[936]&~m[980])|(m[933]&m[934]&~m[935]&~m[936]&m[980])|(m[933]&~m[934]&m[935]&~m[936]&m[980])|(~m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&~m[936]&m[980])|(m[933]&m[934]&m[935]&m[936]&m[980]));
    m[942] = (((m[938]&~m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&m[939]&~m[940]&~m[941]&~m[985])|(~m[938]&~m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&~m[940]&m[941]&~m[985])|(m[938]&~m[939]&m[940]&m[941]&~m[985])|(~m[938]&m[939]&m[940]&m[941]&~m[985]))&BiasedRNG[741])|(((m[938]&~m[939]&~m[940]&~m[941]&m[985])|(~m[938]&m[939]&~m[940]&~m[941]&m[985])|(~m[938]&~m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&~m[940]&m[941]&m[985])|(m[938]&~m[939]&m[940]&m[941]&m[985])|(~m[938]&m[939]&m[940]&m[941]&m[985]))&~BiasedRNG[741])|((m[938]&m[939]&~m[940]&~m[941]&~m[985])|(m[938]&~m[939]&m[940]&~m[941]&~m[985])|(~m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&~m[941]&~m[985])|(m[938]&m[939]&m[940]&m[941]&~m[985])|(m[938]&m[939]&~m[940]&~m[941]&m[985])|(m[938]&~m[939]&m[940]&~m[941]&m[985])|(~m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&~m[941]&m[985])|(m[938]&m[939]&m[940]&m[941]&m[985]));
    m[947] = (((m[943]&~m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&m[944]&~m[945]&~m[946]&~m[990])|(~m[943]&~m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&~m[945]&m[946]&~m[990])|(m[943]&~m[944]&m[945]&m[946]&~m[990])|(~m[943]&m[944]&m[945]&m[946]&~m[990]))&BiasedRNG[742])|(((m[943]&~m[944]&~m[945]&~m[946]&m[990])|(~m[943]&m[944]&~m[945]&~m[946]&m[990])|(~m[943]&~m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&~m[945]&m[946]&m[990])|(m[943]&~m[944]&m[945]&m[946]&m[990])|(~m[943]&m[944]&m[945]&m[946]&m[990]))&~BiasedRNG[742])|((m[943]&m[944]&~m[945]&~m[946]&~m[990])|(m[943]&~m[944]&m[945]&~m[946]&~m[990])|(~m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&~m[946]&~m[990])|(m[943]&m[944]&m[945]&m[946]&~m[990])|(m[943]&m[944]&~m[945]&~m[946]&m[990])|(m[943]&~m[944]&m[945]&~m[946]&m[990])|(~m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&~m[946]&m[990])|(m[943]&m[944]&m[945]&m[946]&m[990]));
    m[952] = (((m[948]&~m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&m[949]&~m[950]&~m[951]&~m[995])|(~m[948]&~m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&~m[950]&m[951]&~m[995])|(m[948]&~m[949]&m[950]&m[951]&~m[995])|(~m[948]&m[949]&m[950]&m[951]&~m[995]))&BiasedRNG[743])|(((m[948]&~m[949]&~m[950]&~m[951]&m[995])|(~m[948]&m[949]&~m[950]&~m[951]&m[995])|(~m[948]&~m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&~m[950]&m[951]&m[995])|(m[948]&~m[949]&m[950]&m[951]&m[995])|(~m[948]&m[949]&m[950]&m[951]&m[995]))&~BiasedRNG[743])|((m[948]&m[949]&~m[950]&~m[951]&~m[995])|(m[948]&~m[949]&m[950]&~m[951]&~m[995])|(~m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&~m[951]&~m[995])|(m[948]&m[949]&m[950]&m[951]&~m[995])|(m[948]&m[949]&~m[950]&~m[951]&m[995])|(m[948]&~m[949]&m[950]&~m[951]&m[995])|(~m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&~m[951]&m[995])|(m[948]&m[949]&m[950]&m[951]&m[995]));
    m[957] = (((m[953]&~m[954]&~m[955]&~m[956]&~m[1005])|(~m[953]&m[954]&~m[955]&~m[956]&~m[1005])|(~m[953]&~m[954]&m[955]&~m[956]&~m[1005])|(m[953]&m[954]&~m[955]&m[956]&~m[1005])|(m[953]&~m[954]&m[955]&m[956]&~m[1005])|(~m[953]&m[954]&m[955]&m[956]&~m[1005]))&BiasedRNG[744])|(((m[953]&~m[954]&~m[955]&~m[956]&m[1005])|(~m[953]&m[954]&~m[955]&~m[956]&m[1005])|(~m[953]&~m[954]&m[955]&~m[956]&m[1005])|(m[953]&m[954]&~m[955]&m[956]&m[1005])|(m[953]&~m[954]&m[955]&m[956]&m[1005])|(~m[953]&m[954]&m[955]&m[956]&m[1005]))&~BiasedRNG[744])|((m[953]&m[954]&~m[955]&~m[956]&~m[1005])|(m[953]&~m[954]&m[955]&~m[956]&~m[1005])|(~m[953]&m[954]&m[955]&~m[956]&~m[1005])|(m[953]&m[954]&m[955]&~m[956]&~m[1005])|(m[953]&m[954]&m[955]&m[956]&~m[1005])|(m[953]&m[954]&~m[955]&~m[956]&m[1005])|(m[953]&~m[954]&m[955]&~m[956]&m[1005])|(~m[953]&m[954]&m[955]&~m[956]&m[1005])|(m[953]&m[954]&m[955]&~m[956]&m[1005])|(m[953]&m[954]&m[955]&m[956]&m[1005]));
    m[962] = (((m[958]&~m[959]&~m[960]&~m[961]&~m[1010])|(~m[958]&m[959]&~m[960]&~m[961]&~m[1010])|(~m[958]&~m[959]&m[960]&~m[961]&~m[1010])|(m[958]&m[959]&~m[960]&m[961]&~m[1010])|(m[958]&~m[959]&m[960]&m[961]&~m[1010])|(~m[958]&m[959]&m[960]&m[961]&~m[1010]))&BiasedRNG[745])|(((m[958]&~m[959]&~m[960]&~m[961]&m[1010])|(~m[958]&m[959]&~m[960]&~m[961]&m[1010])|(~m[958]&~m[959]&m[960]&~m[961]&m[1010])|(m[958]&m[959]&~m[960]&m[961]&m[1010])|(m[958]&~m[959]&m[960]&m[961]&m[1010])|(~m[958]&m[959]&m[960]&m[961]&m[1010]))&~BiasedRNG[745])|((m[958]&m[959]&~m[960]&~m[961]&~m[1010])|(m[958]&~m[959]&m[960]&~m[961]&~m[1010])|(~m[958]&m[959]&m[960]&~m[961]&~m[1010])|(m[958]&m[959]&m[960]&~m[961]&~m[1010])|(m[958]&m[959]&m[960]&m[961]&~m[1010])|(m[958]&m[959]&~m[960]&~m[961]&m[1010])|(m[958]&~m[959]&m[960]&~m[961]&m[1010])|(~m[958]&m[959]&m[960]&~m[961]&m[1010])|(m[958]&m[959]&m[960]&~m[961]&m[1010])|(m[958]&m[959]&m[960]&m[961]&m[1010]));
    m[967] = (((m[963]&~m[964]&~m[965]&~m[966]&~m[1015])|(~m[963]&m[964]&~m[965]&~m[966]&~m[1015])|(~m[963]&~m[964]&m[965]&~m[966]&~m[1015])|(m[963]&m[964]&~m[965]&m[966]&~m[1015])|(m[963]&~m[964]&m[965]&m[966]&~m[1015])|(~m[963]&m[964]&m[965]&m[966]&~m[1015]))&BiasedRNG[746])|(((m[963]&~m[964]&~m[965]&~m[966]&m[1015])|(~m[963]&m[964]&~m[965]&~m[966]&m[1015])|(~m[963]&~m[964]&m[965]&~m[966]&m[1015])|(m[963]&m[964]&~m[965]&m[966]&m[1015])|(m[963]&~m[964]&m[965]&m[966]&m[1015])|(~m[963]&m[964]&m[965]&m[966]&m[1015]))&~BiasedRNG[746])|((m[963]&m[964]&~m[965]&~m[966]&~m[1015])|(m[963]&~m[964]&m[965]&~m[966]&~m[1015])|(~m[963]&m[964]&m[965]&~m[966]&~m[1015])|(m[963]&m[964]&m[965]&~m[966]&~m[1015])|(m[963]&m[964]&m[965]&m[966]&~m[1015])|(m[963]&m[964]&~m[965]&~m[966]&m[1015])|(m[963]&~m[964]&m[965]&~m[966]&m[1015])|(~m[963]&m[964]&m[965]&~m[966]&m[1015])|(m[963]&m[964]&m[965]&~m[966]&m[1015])|(m[963]&m[964]&m[965]&m[966]&m[1015]));
    m[972] = (((m[968]&~m[969]&~m[970]&~m[971]&~m[1020])|(~m[968]&m[969]&~m[970]&~m[971]&~m[1020])|(~m[968]&~m[969]&m[970]&~m[971]&~m[1020])|(m[968]&m[969]&~m[970]&m[971]&~m[1020])|(m[968]&~m[969]&m[970]&m[971]&~m[1020])|(~m[968]&m[969]&m[970]&m[971]&~m[1020]))&BiasedRNG[747])|(((m[968]&~m[969]&~m[970]&~m[971]&m[1020])|(~m[968]&m[969]&~m[970]&~m[971]&m[1020])|(~m[968]&~m[969]&m[970]&~m[971]&m[1020])|(m[968]&m[969]&~m[970]&m[971]&m[1020])|(m[968]&~m[969]&m[970]&m[971]&m[1020])|(~m[968]&m[969]&m[970]&m[971]&m[1020]))&~BiasedRNG[747])|((m[968]&m[969]&~m[970]&~m[971]&~m[1020])|(m[968]&~m[969]&m[970]&~m[971]&~m[1020])|(~m[968]&m[969]&m[970]&~m[971]&~m[1020])|(m[968]&m[969]&m[970]&~m[971]&~m[1020])|(m[968]&m[969]&m[970]&m[971]&~m[1020])|(m[968]&m[969]&~m[970]&~m[971]&m[1020])|(m[968]&~m[969]&m[970]&~m[971]&m[1020])|(~m[968]&m[969]&m[970]&~m[971]&m[1020])|(m[968]&m[969]&m[970]&~m[971]&m[1020])|(m[968]&m[969]&m[970]&m[971]&m[1020]));
    m[977] = (((m[973]&~m[974]&~m[975]&~m[976]&~m[1025])|(~m[973]&m[974]&~m[975]&~m[976]&~m[1025])|(~m[973]&~m[974]&m[975]&~m[976]&~m[1025])|(m[973]&m[974]&~m[975]&m[976]&~m[1025])|(m[973]&~m[974]&m[975]&m[976]&~m[1025])|(~m[973]&m[974]&m[975]&m[976]&~m[1025]))&BiasedRNG[748])|(((m[973]&~m[974]&~m[975]&~m[976]&m[1025])|(~m[973]&m[974]&~m[975]&~m[976]&m[1025])|(~m[973]&~m[974]&m[975]&~m[976]&m[1025])|(m[973]&m[974]&~m[975]&m[976]&m[1025])|(m[973]&~m[974]&m[975]&m[976]&m[1025])|(~m[973]&m[974]&m[975]&m[976]&m[1025]))&~BiasedRNG[748])|((m[973]&m[974]&~m[975]&~m[976]&~m[1025])|(m[973]&~m[974]&m[975]&~m[976]&~m[1025])|(~m[973]&m[974]&m[975]&~m[976]&~m[1025])|(m[973]&m[974]&m[975]&~m[976]&~m[1025])|(m[973]&m[974]&m[975]&m[976]&~m[1025])|(m[973]&m[974]&~m[975]&~m[976]&m[1025])|(m[973]&~m[974]&m[975]&~m[976]&m[1025])|(~m[973]&m[974]&m[975]&~m[976]&m[1025])|(m[973]&m[974]&m[975]&~m[976]&m[1025])|(m[973]&m[974]&m[975]&m[976]&m[1025]));
    m[982] = (((m[978]&~m[979]&~m[980]&~m[981]&~m[1030])|(~m[978]&m[979]&~m[980]&~m[981]&~m[1030])|(~m[978]&~m[979]&m[980]&~m[981]&~m[1030])|(m[978]&m[979]&~m[980]&m[981]&~m[1030])|(m[978]&~m[979]&m[980]&m[981]&~m[1030])|(~m[978]&m[979]&m[980]&m[981]&~m[1030]))&BiasedRNG[749])|(((m[978]&~m[979]&~m[980]&~m[981]&m[1030])|(~m[978]&m[979]&~m[980]&~m[981]&m[1030])|(~m[978]&~m[979]&m[980]&~m[981]&m[1030])|(m[978]&m[979]&~m[980]&m[981]&m[1030])|(m[978]&~m[979]&m[980]&m[981]&m[1030])|(~m[978]&m[979]&m[980]&m[981]&m[1030]))&~BiasedRNG[749])|((m[978]&m[979]&~m[980]&~m[981]&~m[1030])|(m[978]&~m[979]&m[980]&~m[981]&~m[1030])|(~m[978]&m[979]&m[980]&~m[981]&~m[1030])|(m[978]&m[979]&m[980]&~m[981]&~m[1030])|(m[978]&m[979]&m[980]&m[981]&~m[1030])|(m[978]&m[979]&~m[980]&~m[981]&m[1030])|(m[978]&~m[979]&m[980]&~m[981]&m[1030])|(~m[978]&m[979]&m[980]&~m[981]&m[1030])|(m[978]&m[979]&m[980]&~m[981]&m[1030])|(m[978]&m[979]&m[980]&m[981]&m[1030]));
    m[987] = (((m[983]&~m[984]&~m[985]&~m[986]&~m[1035])|(~m[983]&m[984]&~m[985]&~m[986]&~m[1035])|(~m[983]&~m[984]&m[985]&~m[986]&~m[1035])|(m[983]&m[984]&~m[985]&m[986]&~m[1035])|(m[983]&~m[984]&m[985]&m[986]&~m[1035])|(~m[983]&m[984]&m[985]&m[986]&~m[1035]))&BiasedRNG[750])|(((m[983]&~m[984]&~m[985]&~m[986]&m[1035])|(~m[983]&m[984]&~m[985]&~m[986]&m[1035])|(~m[983]&~m[984]&m[985]&~m[986]&m[1035])|(m[983]&m[984]&~m[985]&m[986]&m[1035])|(m[983]&~m[984]&m[985]&m[986]&m[1035])|(~m[983]&m[984]&m[985]&m[986]&m[1035]))&~BiasedRNG[750])|((m[983]&m[984]&~m[985]&~m[986]&~m[1035])|(m[983]&~m[984]&m[985]&~m[986]&~m[1035])|(~m[983]&m[984]&m[985]&~m[986]&~m[1035])|(m[983]&m[984]&m[985]&~m[986]&~m[1035])|(m[983]&m[984]&m[985]&m[986]&~m[1035])|(m[983]&m[984]&~m[985]&~m[986]&m[1035])|(m[983]&~m[984]&m[985]&~m[986]&m[1035])|(~m[983]&m[984]&m[985]&~m[986]&m[1035])|(m[983]&m[984]&m[985]&~m[986]&m[1035])|(m[983]&m[984]&m[985]&m[986]&m[1035]));
    m[992] = (((m[988]&~m[989]&~m[990]&~m[991]&~m[1040])|(~m[988]&m[989]&~m[990]&~m[991]&~m[1040])|(~m[988]&~m[989]&m[990]&~m[991]&~m[1040])|(m[988]&m[989]&~m[990]&m[991]&~m[1040])|(m[988]&~m[989]&m[990]&m[991]&~m[1040])|(~m[988]&m[989]&m[990]&m[991]&~m[1040]))&BiasedRNG[751])|(((m[988]&~m[989]&~m[990]&~m[991]&m[1040])|(~m[988]&m[989]&~m[990]&~m[991]&m[1040])|(~m[988]&~m[989]&m[990]&~m[991]&m[1040])|(m[988]&m[989]&~m[990]&m[991]&m[1040])|(m[988]&~m[989]&m[990]&m[991]&m[1040])|(~m[988]&m[989]&m[990]&m[991]&m[1040]))&~BiasedRNG[751])|((m[988]&m[989]&~m[990]&~m[991]&~m[1040])|(m[988]&~m[989]&m[990]&~m[991]&~m[1040])|(~m[988]&m[989]&m[990]&~m[991]&~m[1040])|(m[988]&m[989]&m[990]&~m[991]&~m[1040])|(m[988]&m[989]&m[990]&m[991]&~m[1040])|(m[988]&m[989]&~m[990]&~m[991]&m[1040])|(m[988]&~m[989]&m[990]&~m[991]&m[1040])|(~m[988]&m[989]&m[990]&~m[991]&m[1040])|(m[988]&m[989]&m[990]&~m[991]&m[1040])|(m[988]&m[989]&m[990]&m[991]&m[1040]));
    m[997] = (((m[993]&~m[994]&~m[995]&~m[996]&~m[1045])|(~m[993]&m[994]&~m[995]&~m[996]&~m[1045])|(~m[993]&~m[994]&m[995]&~m[996]&~m[1045])|(m[993]&m[994]&~m[995]&m[996]&~m[1045])|(m[993]&~m[994]&m[995]&m[996]&~m[1045])|(~m[993]&m[994]&m[995]&m[996]&~m[1045]))&BiasedRNG[752])|(((m[993]&~m[994]&~m[995]&~m[996]&m[1045])|(~m[993]&m[994]&~m[995]&~m[996]&m[1045])|(~m[993]&~m[994]&m[995]&~m[996]&m[1045])|(m[993]&m[994]&~m[995]&m[996]&m[1045])|(m[993]&~m[994]&m[995]&m[996]&m[1045])|(~m[993]&m[994]&m[995]&m[996]&m[1045]))&~BiasedRNG[752])|((m[993]&m[994]&~m[995]&~m[996]&~m[1045])|(m[993]&~m[994]&m[995]&~m[996]&~m[1045])|(~m[993]&m[994]&m[995]&~m[996]&~m[1045])|(m[993]&m[994]&m[995]&~m[996]&~m[1045])|(m[993]&m[994]&m[995]&m[996]&~m[1045])|(m[993]&m[994]&~m[995]&~m[996]&m[1045])|(m[993]&~m[994]&m[995]&~m[996]&m[1045])|(~m[993]&m[994]&m[995]&~m[996]&m[1045])|(m[993]&m[994]&m[995]&~m[996]&m[1045])|(m[993]&m[994]&m[995]&m[996]&m[1045]));
    m[1002] = (((m[998]&~m[999]&~m[1000]&~m[1001]&~m[1050])|(~m[998]&m[999]&~m[1000]&~m[1001]&~m[1050])|(~m[998]&~m[999]&m[1000]&~m[1001]&~m[1050])|(m[998]&m[999]&~m[1000]&m[1001]&~m[1050])|(m[998]&~m[999]&m[1000]&m[1001]&~m[1050])|(~m[998]&m[999]&m[1000]&m[1001]&~m[1050]))&BiasedRNG[753])|(((m[998]&~m[999]&~m[1000]&~m[1001]&m[1050])|(~m[998]&m[999]&~m[1000]&~m[1001]&m[1050])|(~m[998]&~m[999]&m[1000]&~m[1001]&m[1050])|(m[998]&m[999]&~m[1000]&m[1001]&m[1050])|(m[998]&~m[999]&m[1000]&m[1001]&m[1050])|(~m[998]&m[999]&m[1000]&m[1001]&m[1050]))&~BiasedRNG[753])|((m[998]&m[999]&~m[1000]&~m[1001]&~m[1050])|(m[998]&~m[999]&m[1000]&~m[1001]&~m[1050])|(~m[998]&m[999]&m[1000]&~m[1001]&~m[1050])|(m[998]&m[999]&m[1000]&~m[1001]&~m[1050])|(m[998]&m[999]&m[1000]&m[1001]&~m[1050])|(m[998]&m[999]&~m[1000]&~m[1001]&m[1050])|(m[998]&~m[999]&m[1000]&~m[1001]&m[1050])|(~m[998]&m[999]&m[1000]&~m[1001]&m[1050])|(m[998]&m[999]&m[1000]&~m[1001]&m[1050])|(m[998]&m[999]&m[1000]&m[1001]&m[1050]));
    m[1007] = (((m[1003]&~m[1004]&~m[1005]&~m[1006]&~m[1060])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1060])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1060])|(m[1003]&m[1004]&~m[1005]&m[1006]&~m[1060])|(m[1003]&~m[1004]&m[1005]&m[1006]&~m[1060])|(~m[1003]&m[1004]&m[1005]&m[1006]&~m[1060]))&BiasedRNG[754])|(((m[1003]&~m[1004]&~m[1005]&~m[1006]&m[1060])|(~m[1003]&m[1004]&~m[1005]&~m[1006]&m[1060])|(~m[1003]&~m[1004]&m[1005]&~m[1006]&m[1060])|(m[1003]&m[1004]&~m[1005]&m[1006]&m[1060])|(m[1003]&~m[1004]&m[1005]&m[1006]&m[1060])|(~m[1003]&m[1004]&m[1005]&m[1006]&m[1060]))&~BiasedRNG[754])|((m[1003]&m[1004]&~m[1005]&~m[1006]&~m[1060])|(m[1003]&~m[1004]&m[1005]&~m[1006]&~m[1060])|(~m[1003]&m[1004]&m[1005]&~m[1006]&~m[1060])|(m[1003]&m[1004]&m[1005]&~m[1006]&~m[1060])|(m[1003]&m[1004]&m[1005]&m[1006]&~m[1060])|(m[1003]&m[1004]&~m[1005]&~m[1006]&m[1060])|(m[1003]&~m[1004]&m[1005]&~m[1006]&m[1060])|(~m[1003]&m[1004]&m[1005]&~m[1006]&m[1060])|(m[1003]&m[1004]&m[1005]&~m[1006]&m[1060])|(m[1003]&m[1004]&m[1005]&m[1006]&m[1060]));
    m[1012] = (((m[1008]&~m[1009]&~m[1010]&~m[1011]&~m[1065])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1065])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1065])|(m[1008]&m[1009]&~m[1010]&m[1011]&~m[1065])|(m[1008]&~m[1009]&m[1010]&m[1011]&~m[1065])|(~m[1008]&m[1009]&m[1010]&m[1011]&~m[1065]))&BiasedRNG[755])|(((m[1008]&~m[1009]&~m[1010]&~m[1011]&m[1065])|(~m[1008]&m[1009]&~m[1010]&~m[1011]&m[1065])|(~m[1008]&~m[1009]&m[1010]&~m[1011]&m[1065])|(m[1008]&m[1009]&~m[1010]&m[1011]&m[1065])|(m[1008]&~m[1009]&m[1010]&m[1011]&m[1065])|(~m[1008]&m[1009]&m[1010]&m[1011]&m[1065]))&~BiasedRNG[755])|((m[1008]&m[1009]&~m[1010]&~m[1011]&~m[1065])|(m[1008]&~m[1009]&m[1010]&~m[1011]&~m[1065])|(~m[1008]&m[1009]&m[1010]&~m[1011]&~m[1065])|(m[1008]&m[1009]&m[1010]&~m[1011]&~m[1065])|(m[1008]&m[1009]&m[1010]&m[1011]&~m[1065])|(m[1008]&m[1009]&~m[1010]&~m[1011]&m[1065])|(m[1008]&~m[1009]&m[1010]&~m[1011]&m[1065])|(~m[1008]&m[1009]&m[1010]&~m[1011]&m[1065])|(m[1008]&m[1009]&m[1010]&~m[1011]&m[1065])|(m[1008]&m[1009]&m[1010]&m[1011]&m[1065]));
    m[1017] = (((m[1013]&~m[1014]&~m[1015]&~m[1016]&~m[1070])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1070])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1070])|(m[1013]&m[1014]&~m[1015]&m[1016]&~m[1070])|(m[1013]&~m[1014]&m[1015]&m[1016]&~m[1070])|(~m[1013]&m[1014]&m[1015]&m[1016]&~m[1070]))&BiasedRNG[756])|(((m[1013]&~m[1014]&~m[1015]&~m[1016]&m[1070])|(~m[1013]&m[1014]&~m[1015]&~m[1016]&m[1070])|(~m[1013]&~m[1014]&m[1015]&~m[1016]&m[1070])|(m[1013]&m[1014]&~m[1015]&m[1016]&m[1070])|(m[1013]&~m[1014]&m[1015]&m[1016]&m[1070])|(~m[1013]&m[1014]&m[1015]&m[1016]&m[1070]))&~BiasedRNG[756])|((m[1013]&m[1014]&~m[1015]&~m[1016]&~m[1070])|(m[1013]&~m[1014]&m[1015]&~m[1016]&~m[1070])|(~m[1013]&m[1014]&m[1015]&~m[1016]&~m[1070])|(m[1013]&m[1014]&m[1015]&~m[1016]&~m[1070])|(m[1013]&m[1014]&m[1015]&m[1016]&~m[1070])|(m[1013]&m[1014]&~m[1015]&~m[1016]&m[1070])|(m[1013]&~m[1014]&m[1015]&~m[1016]&m[1070])|(~m[1013]&m[1014]&m[1015]&~m[1016]&m[1070])|(m[1013]&m[1014]&m[1015]&~m[1016]&m[1070])|(m[1013]&m[1014]&m[1015]&m[1016]&m[1070]));
    m[1022] = (((m[1018]&~m[1019]&~m[1020]&~m[1021]&~m[1075])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1075])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1075])|(m[1018]&m[1019]&~m[1020]&m[1021]&~m[1075])|(m[1018]&~m[1019]&m[1020]&m[1021]&~m[1075])|(~m[1018]&m[1019]&m[1020]&m[1021]&~m[1075]))&BiasedRNG[757])|(((m[1018]&~m[1019]&~m[1020]&~m[1021]&m[1075])|(~m[1018]&m[1019]&~m[1020]&~m[1021]&m[1075])|(~m[1018]&~m[1019]&m[1020]&~m[1021]&m[1075])|(m[1018]&m[1019]&~m[1020]&m[1021]&m[1075])|(m[1018]&~m[1019]&m[1020]&m[1021]&m[1075])|(~m[1018]&m[1019]&m[1020]&m[1021]&m[1075]))&~BiasedRNG[757])|((m[1018]&m[1019]&~m[1020]&~m[1021]&~m[1075])|(m[1018]&~m[1019]&m[1020]&~m[1021]&~m[1075])|(~m[1018]&m[1019]&m[1020]&~m[1021]&~m[1075])|(m[1018]&m[1019]&m[1020]&~m[1021]&~m[1075])|(m[1018]&m[1019]&m[1020]&m[1021]&~m[1075])|(m[1018]&m[1019]&~m[1020]&~m[1021]&m[1075])|(m[1018]&~m[1019]&m[1020]&~m[1021]&m[1075])|(~m[1018]&m[1019]&m[1020]&~m[1021]&m[1075])|(m[1018]&m[1019]&m[1020]&~m[1021]&m[1075])|(m[1018]&m[1019]&m[1020]&m[1021]&m[1075]));
    m[1027] = (((m[1023]&~m[1024]&~m[1025]&~m[1026]&~m[1080])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1080])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1080])|(m[1023]&m[1024]&~m[1025]&m[1026]&~m[1080])|(m[1023]&~m[1024]&m[1025]&m[1026]&~m[1080])|(~m[1023]&m[1024]&m[1025]&m[1026]&~m[1080]))&BiasedRNG[758])|(((m[1023]&~m[1024]&~m[1025]&~m[1026]&m[1080])|(~m[1023]&m[1024]&~m[1025]&~m[1026]&m[1080])|(~m[1023]&~m[1024]&m[1025]&~m[1026]&m[1080])|(m[1023]&m[1024]&~m[1025]&m[1026]&m[1080])|(m[1023]&~m[1024]&m[1025]&m[1026]&m[1080])|(~m[1023]&m[1024]&m[1025]&m[1026]&m[1080]))&~BiasedRNG[758])|((m[1023]&m[1024]&~m[1025]&~m[1026]&~m[1080])|(m[1023]&~m[1024]&m[1025]&~m[1026]&~m[1080])|(~m[1023]&m[1024]&m[1025]&~m[1026]&~m[1080])|(m[1023]&m[1024]&m[1025]&~m[1026]&~m[1080])|(m[1023]&m[1024]&m[1025]&m[1026]&~m[1080])|(m[1023]&m[1024]&~m[1025]&~m[1026]&m[1080])|(m[1023]&~m[1024]&m[1025]&~m[1026]&m[1080])|(~m[1023]&m[1024]&m[1025]&~m[1026]&m[1080])|(m[1023]&m[1024]&m[1025]&~m[1026]&m[1080])|(m[1023]&m[1024]&m[1025]&m[1026]&m[1080]));
    m[1032] = (((m[1028]&~m[1029]&~m[1030]&~m[1031]&~m[1085])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1085])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1085])|(m[1028]&m[1029]&~m[1030]&m[1031]&~m[1085])|(m[1028]&~m[1029]&m[1030]&m[1031]&~m[1085])|(~m[1028]&m[1029]&m[1030]&m[1031]&~m[1085]))&BiasedRNG[759])|(((m[1028]&~m[1029]&~m[1030]&~m[1031]&m[1085])|(~m[1028]&m[1029]&~m[1030]&~m[1031]&m[1085])|(~m[1028]&~m[1029]&m[1030]&~m[1031]&m[1085])|(m[1028]&m[1029]&~m[1030]&m[1031]&m[1085])|(m[1028]&~m[1029]&m[1030]&m[1031]&m[1085])|(~m[1028]&m[1029]&m[1030]&m[1031]&m[1085]))&~BiasedRNG[759])|((m[1028]&m[1029]&~m[1030]&~m[1031]&~m[1085])|(m[1028]&~m[1029]&m[1030]&~m[1031]&~m[1085])|(~m[1028]&m[1029]&m[1030]&~m[1031]&~m[1085])|(m[1028]&m[1029]&m[1030]&~m[1031]&~m[1085])|(m[1028]&m[1029]&m[1030]&m[1031]&~m[1085])|(m[1028]&m[1029]&~m[1030]&~m[1031]&m[1085])|(m[1028]&~m[1029]&m[1030]&~m[1031]&m[1085])|(~m[1028]&m[1029]&m[1030]&~m[1031]&m[1085])|(m[1028]&m[1029]&m[1030]&~m[1031]&m[1085])|(m[1028]&m[1029]&m[1030]&m[1031]&m[1085]));
    m[1037] = (((m[1033]&~m[1034]&~m[1035]&~m[1036]&~m[1090])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1090])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1090])|(m[1033]&m[1034]&~m[1035]&m[1036]&~m[1090])|(m[1033]&~m[1034]&m[1035]&m[1036]&~m[1090])|(~m[1033]&m[1034]&m[1035]&m[1036]&~m[1090]))&BiasedRNG[760])|(((m[1033]&~m[1034]&~m[1035]&~m[1036]&m[1090])|(~m[1033]&m[1034]&~m[1035]&~m[1036]&m[1090])|(~m[1033]&~m[1034]&m[1035]&~m[1036]&m[1090])|(m[1033]&m[1034]&~m[1035]&m[1036]&m[1090])|(m[1033]&~m[1034]&m[1035]&m[1036]&m[1090])|(~m[1033]&m[1034]&m[1035]&m[1036]&m[1090]))&~BiasedRNG[760])|((m[1033]&m[1034]&~m[1035]&~m[1036]&~m[1090])|(m[1033]&~m[1034]&m[1035]&~m[1036]&~m[1090])|(~m[1033]&m[1034]&m[1035]&~m[1036]&~m[1090])|(m[1033]&m[1034]&m[1035]&~m[1036]&~m[1090])|(m[1033]&m[1034]&m[1035]&m[1036]&~m[1090])|(m[1033]&m[1034]&~m[1035]&~m[1036]&m[1090])|(m[1033]&~m[1034]&m[1035]&~m[1036]&m[1090])|(~m[1033]&m[1034]&m[1035]&~m[1036]&m[1090])|(m[1033]&m[1034]&m[1035]&~m[1036]&m[1090])|(m[1033]&m[1034]&m[1035]&m[1036]&m[1090]));
    m[1042] = (((m[1038]&~m[1039]&~m[1040]&~m[1041]&~m[1095])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1095])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1095])|(m[1038]&m[1039]&~m[1040]&m[1041]&~m[1095])|(m[1038]&~m[1039]&m[1040]&m[1041]&~m[1095])|(~m[1038]&m[1039]&m[1040]&m[1041]&~m[1095]))&BiasedRNG[761])|(((m[1038]&~m[1039]&~m[1040]&~m[1041]&m[1095])|(~m[1038]&m[1039]&~m[1040]&~m[1041]&m[1095])|(~m[1038]&~m[1039]&m[1040]&~m[1041]&m[1095])|(m[1038]&m[1039]&~m[1040]&m[1041]&m[1095])|(m[1038]&~m[1039]&m[1040]&m[1041]&m[1095])|(~m[1038]&m[1039]&m[1040]&m[1041]&m[1095]))&~BiasedRNG[761])|((m[1038]&m[1039]&~m[1040]&~m[1041]&~m[1095])|(m[1038]&~m[1039]&m[1040]&~m[1041]&~m[1095])|(~m[1038]&m[1039]&m[1040]&~m[1041]&~m[1095])|(m[1038]&m[1039]&m[1040]&~m[1041]&~m[1095])|(m[1038]&m[1039]&m[1040]&m[1041]&~m[1095])|(m[1038]&m[1039]&~m[1040]&~m[1041]&m[1095])|(m[1038]&~m[1039]&m[1040]&~m[1041]&m[1095])|(~m[1038]&m[1039]&m[1040]&~m[1041]&m[1095])|(m[1038]&m[1039]&m[1040]&~m[1041]&m[1095])|(m[1038]&m[1039]&m[1040]&m[1041]&m[1095]));
    m[1047] = (((m[1043]&~m[1044]&~m[1045]&~m[1046]&~m[1100])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1100])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1100])|(m[1043]&m[1044]&~m[1045]&m[1046]&~m[1100])|(m[1043]&~m[1044]&m[1045]&m[1046]&~m[1100])|(~m[1043]&m[1044]&m[1045]&m[1046]&~m[1100]))&BiasedRNG[762])|(((m[1043]&~m[1044]&~m[1045]&~m[1046]&m[1100])|(~m[1043]&m[1044]&~m[1045]&~m[1046]&m[1100])|(~m[1043]&~m[1044]&m[1045]&~m[1046]&m[1100])|(m[1043]&m[1044]&~m[1045]&m[1046]&m[1100])|(m[1043]&~m[1044]&m[1045]&m[1046]&m[1100])|(~m[1043]&m[1044]&m[1045]&m[1046]&m[1100]))&~BiasedRNG[762])|((m[1043]&m[1044]&~m[1045]&~m[1046]&~m[1100])|(m[1043]&~m[1044]&m[1045]&~m[1046]&~m[1100])|(~m[1043]&m[1044]&m[1045]&~m[1046]&~m[1100])|(m[1043]&m[1044]&m[1045]&~m[1046]&~m[1100])|(m[1043]&m[1044]&m[1045]&m[1046]&~m[1100])|(m[1043]&m[1044]&~m[1045]&~m[1046]&m[1100])|(m[1043]&~m[1044]&m[1045]&~m[1046]&m[1100])|(~m[1043]&m[1044]&m[1045]&~m[1046]&m[1100])|(m[1043]&m[1044]&m[1045]&~m[1046]&m[1100])|(m[1043]&m[1044]&m[1045]&m[1046]&m[1100]));
    m[1052] = (((m[1048]&~m[1049]&~m[1050]&~m[1051]&~m[1105])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1105])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1105])|(m[1048]&m[1049]&~m[1050]&m[1051]&~m[1105])|(m[1048]&~m[1049]&m[1050]&m[1051]&~m[1105])|(~m[1048]&m[1049]&m[1050]&m[1051]&~m[1105]))&BiasedRNG[763])|(((m[1048]&~m[1049]&~m[1050]&~m[1051]&m[1105])|(~m[1048]&m[1049]&~m[1050]&~m[1051]&m[1105])|(~m[1048]&~m[1049]&m[1050]&~m[1051]&m[1105])|(m[1048]&m[1049]&~m[1050]&m[1051]&m[1105])|(m[1048]&~m[1049]&m[1050]&m[1051]&m[1105])|(~m[1048]&m[1049]&m[1050]&m[1051]&m[1105]))&~BiasedRNG[763])|((m[1048]&m[1049]&~m[1050]&~m[1051]&~m[1105])|(m[1048]&~m[1049]&m[1050]&~m[1051]&~m[1105])|(~m[1048]&m[1049]&m[1050]&~m[1051]&~m[1105])|(m[1048]&m[1049]&m[1050]&~m[1051]&~m[1105])|(m[1048]&m[1049]&m[1050]&m[1051]&~m[1105])|(m[1048]&m[1049]&~m[1050]&~m[1051]&m[1105])|(m[1048]&~m[1049]&m[1050]&~m[1051]&m[1105])|(~m[1048]&m[1049]&m[1050]&~m[1051]&m[1105])|(m[1048]&m[1049]&m[1050]&~m[1051]&m[1105])|(m[1048]&m[1049]&m[1050]&m[1051]&m[1105]));
    m[1057] = (((m[1053]&~m[1054]&~m[1055]&~m[1056]&~m[1110])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1110])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1110])|(m[1053]&m[1054]&~m[1055]&m[1056]&~m[1110])|(m[1053]&~m[1054]&m[1055]&m[1056]&~m[1110])|(~m[1053]&m[1054]&m[1055]&m[1056]&~m[1110]))&BiasedRNG[764])|(((m[1053]&~m[1054]&~m[1055]&~m[1056]&m[1110])|(~m[1053]&m[1054]&~m[1055]&~m[1056]&m[1110])|(~m[1053]&~m[1054]&m[1055]&~m[1056]&m[1110])|(m[1053]&m[1054]&~m[1055]&m[1056]&m[1110])|(m[1053]&~m[1054]&m[1055]&m[1056]&m[1110])|(~m[1053]&m[1054]&m[1055]&m[1056]&m[1110]))&~BiasedRNG[764])|((m[1053]&m[1054]&~m[1055]&~m[1056]&~m[1110])|(m[1053]&~m[1054]&m[1055]&~m[1056]&~m[1110])|(~m[1053]&m[1054]&m[1055]&~m[1056]&~m[1110])|(m[1053]&m[1054]&m[1055]&~m[1056]&~m[1110])|(m[1053]&m[1054]&m[1055]&m[1056]&~m[1110])|(m[1053]&m[1054]&~m[1055]&~m[1056]&m[1110])|(m[1053]&~m[1054]&m[1055]&~m[1056]&m[1110])|(~m[1053]&m[1054]&m[1055]&~m[1056]&m[1110])|(m[1053]&m[1054]&m[1055]&~m[1056]&m[1110])|(m[1053]&m[1054]&m[1055]&m[1056]&m[1110]));
    m[1062] = (((m[1058]&~m[1059]&~m[1060]&~m[1061]&~m[1120])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1120])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1120])|(m[1058]&m[1059]&~m[1060]&m[1061]&~m[1120])|(m[1058]&~m[1059]&m[1060]&m[1061]&~m[1120])|(~m[1058]&m[1059]&m[1060]&m[1061]&~m[1120]))&BiasedRNG[765])|(((m[1058]&~m[1059]&~m[1060]&~m[1061]&m[1120])|(~m[1058]&m[1059]&~m[1060]&~m[1061]&m[1120])|(~m[1058]&~m[1059]&m[1060]&~m[1061]&m[1120])|(m[1058]&m[1059]&~m[1060]&m[1061]&m[1120])|(m[1058]&~m[1059]&m[1060]&m[1061]&m[1120])|(~m[1058]&m[1059]&m[1060]&m[1061]&m[1120]))&~BiasedRNG[765])|((m[1058]&m[1059]&~m[1060]&~m[1061]&~m[1120])|(m[1058]&~m[1059]&m[1060]&~m[1061]&~m[1120])|(~m[1058]&m[1059]&m[1060]&~m[1061]&~m[1120])|(m[1058]&m[1059]&m[1060]&~m[1061]&~m[1120])|(m[1058]&m[1059]&m[1060]&m[1061]&~m[1120])|(m[1058]&m[1059]&~m[1060]&~m[1061]&m[1120])|(m[1058]&~m[1059]&m[1060]&~m[1061]&m[1120])|(~m[1058]&m[1059]&m[1060]&~m[1061]&m[1120])|(m[1058]&m[1059]&m[1060]&~m[1061]&m[1120])|(m[1058]&m[1059]&m[1060]&m[1061]&m[1120]));
    m[1067] = (((m[1063]&~m[1064]&~m[1065]&~m[1066]&~m[1125])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1125])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1125])|(m[1063]&m[1064]&~m[1065]&m[1066]&~m[1125])|(m[1063]&~m[1064]&m[1065]&m[1066]&~m[1125])|(~m[1063]&m[1064]&m[1065]&m[1066]&~m[1125]))&BiasedRNG[766])|(((m[1063]&~m[1064]&~m[1065]&~m[1066]&m[1125])|(~m[1063]&m[1064]&~m[1065]&~m[1066]&m[1125])|(~m[1063]&~m[1064]&m[1065]&~m[1066]&m[1125])|(m[1063]&m[1064]&~m[1065]&m[1066]&m[1125])|(m[1063]&~m[1064]&m[1065]&m[1066]&m[1125])|(~m[1063]&m[1064]&m[1065]&m[1066]&m[1125]))&~BiasedRNG[766])|((m[1063]&m[1064]&~m[1065]&~m[1066]&~m[1125])|(m[1063]&~m[1064]&m[1065]&~m[1066]&~m[1125])|(~m[1063]&m[1064]&m[1065]&~m[1066]&~m[1125])|(m[1063]&m[1064]&m[1065]&~m[1066]&~m[1125])|(m[1063]&m[1064]&m[1065]&m[1066]&~m[1125])|(m[1063]&m[1064]&~m[1065]&~m[1066]&m[1125])|(m[1063]&~m[1064]&m[1065]&~m[1066]&m[1125])|(~m[1063]&m[1064]&m[1065]&~m[1066]&m[1125])|(m[1063]&m[1064]&m[1065]&~m[1066]&m[1125])|(m[1063]&m[1064]&m[1065]&m[1066]&m[1125]));
    m[1072] = (((m[1068]&~m[1069]&~m[1070]&~m[1071]&~m[1130])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1130])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1130])|(m[1068]&m[1069]&~m[1070]&m[1071]&~m[1130])|(m[1068]&~m[1069]&m[1070]&m[1071]&~m[1130])|(~m[1068]&m[1069]&m[1070]&m[1071]&~m[1130]))&BiasedRNG[767])|(((m[1068]&~m[1069]&~m[1070]&~m[1071]&m[1130])|(~m[1068]&m[1069]&~m[1070]&~m[1071]&m[1130])|(~m[1068]&~m[1069]&m[1070]&~m[1071]&m[1130])|(m[1068]&m[1069]&~m[1070]&m[1071]&m[1130])|(m[1068]&~m[1069]&m[1070]&m[1071]&m[1130])|(~m[1068]&m[1069]&m[1070]&m[1071]&m[1130]))&~BiasedRNG[767])|((m[1068]&m[1069]&~m[1070]&~m[1071]&~m[1130])|(m[1068]&~m[1069]&m[1070]&~m[1071]&~m[1130])|(~m[1068]&m[1069]&m[1070]&~m[1071]&~m[1130])|(m[1068]&m[1069]&m[1070]&~m[1071]&~m[1130])|(m[1068]&m[1069]&m[1070]&m[1071]&~m[1130])|(m[1068]&m[1069]&~m[1070]&~m[1071]&m[1130])|(m[1068]&~m[1069]&m[1070]&~m[1071]&m[1130])|(~m[1068]&m[1069]&m[1070]&~m[1071]&m[1130])|(m[1068]&m[1069]&m[1070]&~m[1071]&m[1130])|(m[1068]&m[1069]&m[1070]&m[1071]&m[1130]));
    m[1077] = (((m[1073]&~m[1074]&~m[1075]&~m[1076]&~m[1135])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1135])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1135])|(m[1073]&m[1074]&~m[1075]&m[1076]&~m[1135])|(m[1073]&~m[1074]&m[1075]&m[1076]&~m[1135])|(~m[1073]&m[1074]&m[1075]&m[1076]&~m[1135]))&BiasedRNG[768])|(((m[1073]&~m[1074]&~m[1075]&~m[1076]&m[1135])|(~m[1073]&m[1074]&~m[1075]&~m[1076]&m[1135])|(~m[1073]&~m[1074]&m[1075]&~m[1076]&m[1135])|(m[1073]&m[1074]&~m[1075]&m[1076]&m[1135])|(m[1073]&~m[1074]&m[1075]&m[1076]&m[1135])|(~m[1073]&m[1074]&m[1075]&m[1076]&m[1135]))&~BiasedRNG[768])|((m[1073]&m[1074]&~m[1075]&~m[1076]&~m[1135])|(m[1073]&~m[1074]&m[1075]&~m[1076]&~m[1135])|(~m[1073]&m[1074]&m[1075]&~m[1076]&~m[1135])|(m[1073]&m[1074]&m[1075]&~m[1076]&~m[1135])|(m[1073]&m[1074]&m[1075]&m[1076]&~m[1135])|(m[1073]&m[1074]&~m[1075]&~m[1076]&m[1135])|(m[1073]&~m[1074]&m[1075]&~m[1076]&m[1135])|(~m[1073]&m[1074]&m[1075]&~m[1076]&m[1135])|(m[1073]&m[1074]&m[1075]&~m[1076]&m[1135])|(m[1073]&m[1074]&m[1075]&m[1076]&m[1135]));
    m[1082] = (((m[1078]&~m[1079]&~m[1080]&~m[1081]&~m[1140])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1140])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1140])|(m[1078]&m[1079]&~m[1080]&m[1081]&~m[1140])|(m[1078]&~m[1079]&m[1080]&m[1081]&~m[1140])|(~m[1078]&m[1079]&m[1080]&m[1081]&~m[1140]))&BiasedRNG[769])|(((m[1078]&~m[1079]&~m[1080]&~m[1081]&m[1140])|(~m[1078]&m[1079]&~m[1080]&~m[1081]&m[1140])|(~m[1078]&~m[1079]&m[1080]&~m[1081]&m[1140])|(m[1078]&m[1079]&~m[1080]&m[1081]&m[1140])|(m[1078]&~m[1079]&m[1080]&m[1081]&m[1140])|(~m[1078]&m[1079]&m[1080]&m[1081]&m[1140]))&~BiasedRNG[769])|((m[1078]&m[1079]&~m[1080]&~m[1081]&~m[1140])|(m[1078]&~m[1079]&m[1080]&~m[1081]&~m[1140])|(~m[1078]&m[1079]&m[1080]&~m[1081]&~m[1140])|(m[1078]&m[1079]&m[1080]&~m[1081]&~m[1140])|(m[1078]&m[1079]&m[1080]&m[1081]&~m[1140])|(m[1078]&m[1079]&~m[1080]&~m[1081]&m[1140])|(m[1078]&~m[1079]&m[1080]&~m[1081]&m[1140])|(~m[1078]&m[1079]&m[1080]&~m[1081]&m[1140])|(m[1078]&m[1079]&m[1080]&~m[1081]&m[1140])|(m[1078]&m[1079]&m[1080]&m[1081]&m[1140]));
    m[1087] = (((m[1083]&~m[1084]&~m[1085]&~m[1086]&~m[1145])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1145])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1145])|(m[1083]&m[1084]&~m[1085]&m[1086]&~m[1145])|(m[1083]&~m[1084]&m[1085]&m[1086]&~m[1145])|(~m[1083]&m[1084]&m[1085]&m[1086]&~m[1145]))&BiasedRNG[770])|(((m[1083]&~m[1084]&~m[1085]&~m[1086]&m[1145])|(~m[1083]&m[1084]&~m[1085]&~m[1086]&m[1145])|(~m[1083]&~m[1084]&m[1085]&~m[1086]&m[1145])|(m[1083]&m[1084]&~m[1085]&m[1086]&m[1145])|(m[1083]&~m[1084]&m[1085]&m[1086]&m[1145])|(~m[1083]&m[1084]&m[1085]&m[1086]&m[1145]))&~BiasedRNG[770])|((m[1083]&m[1084]&~m[1085]&~m[1086]&~m[1145])|(m[1083]&~m[1084]&m[1085]&~m[1086]&~m[1145])|(~m[1083]&m[1084]&m[1085]&~m[1086]&~m[1145])|(m[1083]&m[1084]&m[1085]&~m[1086]&~m[1145])|(m[1083]&m[1084]&m[1085]&m[1086]&~m[1145])|(m[1083]&m[1084]&~m[1085]&~m[1086]&m[1145])|(m[1083]&~m[1084]&m[1085]&~m[1086]&m[1145])|(~m[1083]&m[1084]&m[1085]&~m[1086]&m[1145])|(m[1083]&m[1084]&m[1085]&~m[1086]&m[1145])|(m[1083]&m[1084]&m[1085]&m[1086]&m[1145]));
    m[1092] = (((m[1088]&~m[1089]&~m[1090]&~m[1091]&~m[1150])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1150])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1150])|(m[1088]&m[1089]&~m[1090]&m[1091]&~m[1150])|(m[1088]&~m[1089]&m[1090]&m[1091]&~m[1150])|(~m[1088]&m[1089]&m[1090]&m[1091]&~m[1150]))&BiasedRNG[771])|(((m[1088]&~m[1089]&~m[1090]&~m[1091]&m[1150])|(~m[1088]&m[1089]&~m[1090]&~m[1091]&m[1150])|(~m[1088]&~m[1089]&m[1090]&~m[1091]&m[1150])|(m[1088]&m[1089]&~m[1090]&m[1091]&m[1150])|(m[1088]&~m[1089]&m[1090]&m[1091]&m[1150])|(~m[1088]&m[1089]&m[1090]&m[1091]&m[1150]))&~BiasedRNG[771])|((m[1088]&m[1089]&~m[1090]&~m[1091]&~m[1150])|(m[1088]&~m[1089]&m[1090]&~m[1091]&~m[1150])|(~m[1088]&m[1089]&m[1090]&~m[1091]&~m[1150])|(m[1088]&m[1089]&m[1090]&~m[1091]&~m[1150])|(m[1088]&m[1089]&m[1090]&m[1091]&~m[1150])|(m[1088]&m[1089]&~m[1090]&~m[1091]&m[1150])|(m[1088]&~m[1089]&m[1090]&~m[1091]&m[1150])|(~m[1088]&m[1089]&m[1090]&~m[1091]&m[1150])|(m[1088]&m[1089]&m[1090]&~m[1091]&m[1150])|(m[1088]&m[1089]&m[1090]&m[1091]&m[1150]));
    m[1097] = (((m[1093]&~m[1094]&~m[1095]&~m[1096]&~m[1155])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1155])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1155])|(m[1093]&m[1094]&~m[1095]&m[1096]&~m[1155])|(m[1093]&~m[1094]&m[1095]&m[1096]&~m[1155])|(~m[1093]&m[1094]&m[1095]&m[1096]&~m[1155]))&BiasedRNG[772])|(((m[1093]&~m[1094]&~m[1095]&~m[1096]&m[1155])|(~m[1093]&m[1094]&~m[1095]&~m[1096]&m[1155])|(~m[1093]&~m[1094]&m[1095]&~m[1096]&m[1155])|(m[1093]&m[1094]&~m[1095]&m[1096]&m[1155])|(m[1093]&~m[1094]&m[1095]&m[1096]&m[1155])|(~m[1093]&m[1094]&m[1095]&m[1096]&m[1155]))&~BiasedRNG[772])|((m[1093]&m[1094]&~m[1095]&~m[1096]&~m[1155])|(m[1093]&~m[1094]&m[1095]&~m[1096]&~m[1155])|(~m[1093]&m[1094]&m[1095]&~m[1096]&~m[1155])|(m[1093]&m[1094]&m[1095]&~m[1096]&~m[1155])|(m[1093]&m[1094]&m[1095]&m[1096]&~m[1155])|(m[1093]&m[1094]&~m[1095]&~m[1096]&m[1155])|(m[1093]&~m[1094]&m[1095]&~m[1096]&m[1155])|(~m[1093]&m[1094]&m[1095]&~m[1096]&m[1155])|(m[1093]&m[1094]&m[1095]&~m[1096]&m[1155])|(m[1093]&m[1094]&m[1095]&m[1096]&m[1155]));
    m[1102] = (((m[1098]&~m[1099]&~m[1100]&~m[1101]&~m[1160])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1160])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1160])|(m[1098]&m[1099]&~m[1100]&m[1101]&~m[1160])|(m[1098]&~m[1099]&m[1100]&m[1101]&~m[1160])|(~m[1098]&m[1099]&m[1100]&m[1101]&~m[1160]))&BiasedRNG[773])|(((m[1098]&~m[1099]&~m[1100]&~m[1101]&m[1160])|(~m[1098]&m[1099]&~m[1100]&~m[1101]&m[1160])|(~m[1098]&~m[1099]&m[1100]&~m[1101]&m[1160])|(m[1098]&m[1099]&~m[1100]&m[1101]&m[1160])|(m[1098]&~m[1099]&m[1100]&m[1101]&m[1160])|(~m[1098]&m[1099]&m[1100]&m[1101]&m[1160]))&~BiasedRNG[773])|((m[1098]&m[1099]&~m[1100]&~m[1101]&~m[1160])|(m[1098]&~m[1099]&m[1100]&~m[1101]&~m[1160])|(~m[1098]&m[1099]&m[1100]&~m[1101]&~m[1160])|(m[1098]&m[1099]&m[1100]&~m[1101]&~m[1160])|(m[1098]&m[1099]&m[1100]&m[1101]&~m[1160])|(m[1098]&m[1099]&~m[1100]&~m[1101]&m[1160])|(m[1098]&~m[1099]&m[1100]&~m[1101]&m[1160])|(~m[1098]&m[1099]&m[1100]&~m[1101]&m[1160])|(m[1098]&m[1099]&m[1100]&~m[1101]&m[1160])|(m[1098]&m[1099]&m[1100]&m[1101]&m[1160]));
    m[1107] = (((m[1103]&~m[1104]&~m[1105]&~m[1106]&~m[1165])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1165])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1165])|(m[1103]&m[1104]&~m[1105]&m[1106]&~m[1165])|(m[1103]&~m[1104]&m[1105]&m[1106]&~m[1165])|(~m[1103]&m[1104]&m[1105]&m[1106]&~m[1165]))&BiasedRNG[774])|(((m[1103]&~m[1104]&~m[1105]&~m[1106]&m[1165])|(~m[1103]&m[1104]&~m[1105]&~m[1106]&m[1165])|(~m[1103]&~m[1104]&m[1105]&~m[1106]&m[1165])|(m[1103]&m[1104]&~m[1105]&m[1106]&m[1165])|(m[1103]&~m[1104]&m[1105]&m[1106]&m[1165])|(~m[1103]&m[1104]&m[1105]&m[1106]&m[1165]))&~BiasedRNG[774])|((m[1103]&m[1104]&~m[1105]&~m[1106]&~m[1165])|(m[1103]&~m[1104]&m[1105]&~m[1106]&~m[1165])|(~m[1103]&m[1104]&m[1105]&~m[1106]&~m[1165])|(m[1103]&m[1104]&m[1105]&~m[1106]&~m[1165])|(m[1103]&m[1104]&m[1105]&m[1106]&~m[1165])|(m[1103]&m[1104]&~m[1105]&~m[1106]&m[1165])|(m[1103]&~m[1104]&m[1105]&~m[1106]&m[1165])|(~m[1103]&m[1104]&m[1105]&~m[1106]&m[1165])|(m[1103]&m[1104]&m[1105]&~m[1106]&m[1165])|(m[1103]&m[1104]&m[1105]&m[1106]&m[1165]));
    m[1112] = (((m[1108]&~m[1109]&~m[1110]&~m[1111]&~m[1170])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1170])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1170])|(m[1108]&m[1109]&~m[1110]&m[1111]&~m[1170])|(m[1108]&~m[1109]&m[1110]&m[1111]&~m[1170])|(~m[1108]&m[1109]&m[1110]&m[1111]&~m[1170]))&BiasedRNG[775])|(((m[1108]&~m[1109]&~m[1110]&~m[1111]&m[1170])|(~m[1108]&m[1109]&~m[1110]&~m[1111]&m[1170])|(~m[1108]&~m[1109]&m[1110]&~m[1111]&m[1170])|(m[1108]&m[1109]&~m[1110]&m[1111]&m[1170])|(m[1108]&~m[1109]&m[1110]&m[1111]&m[1170])|(~m[1108]&m[1109]&m[1110]&m[1111]&m[1170]))&~BiasedRNG[775])|((m[1108]&m[1109]&~m[1110]&~m[1111]&~m[1170])|(m[1108]&~m[1109]&m[1110]&~m[1111]&~m[1170])|(~m[1108]&m[1109]&m[1110]&~m[1111]&~m[1170])|(m[1108]&m[1109]&m[1110]&~m[1111]&~m[1170])|(m[1108]&m[1109]&m[1110]&m[1111]&~m[1170])|(m[1108]&m[1109]&~m[1110]&~m[1111]&m[1170])|(m[1108]&~m[1109]&m[1110]&~m[1111]&m[1170])|(~m[1108]&m[1109]&m[1110]&~m[1111]&m[1170])|(m[1108]&m[1109]&m[1110]&~m[1111]&m[1170])|(m[1108]&m[1109]&m[1110]&m[1111]&m[1170]));
    m[1117] = (((m[1113]&~m[1114]&~m[1115]&~m[1116]&~m[1175])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1175])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1175])|(m[1113]&m[1114]&~m[1115]&m[1116]&~m[1175])|(m[1113]&~m[1114]&m[1115]&m[1116]&~m[1175])|(~m[1113]&m[1114]&m[1115]&m[1116]&~m[1175]))&BiasedRNG[776])|(((m[1113]&~m[1114]&~m[1115]&~m[1116]&m[1175])|(~m[1113]&m[1114]&~m[1115]&~m[1116]&m[1175])|(~m[1113]&~m[1114]&m[1115]&~m[1116]&m[1175])|(m[1113]&m[1114]&~m[1115]&m[1116]&m[1175])|(m[1113]&~m[1114]&m[1115]&m[1116]&m[1175])|(~m[1113]&m[1114]&m[1115]&m[1116]&m[1175]))&~BiasedRNG[776])|((m[1113]&m[1114]&~m[1115]&~m[1116]&~m[1175])|(m[1113]&~m[1114]&m[1115]&~m[1116]&~m[1175])|(~m[1113]&m[1114]&m[1115]&~m[1116]&~m[1175])|(m[1113]&m[1114]&m[1115]&~m[1116]&~m[1175])|(m[1113]&m[1114]&m[1115]&m[1116]&~m[1175])|(m[1113]&m[1114]&~m[1115]&~m[1116]&m[1175])|(m[1113]&~m[1114]&m[1115]&~m[1116]&m[1175])|(~m[1113]&m[1114]&m[1115]&~m[1116]&m[1175])|(m[1113]&m[1114]&m[1115]&~m[1116]&m[1175])|(m[1113]&m[1114]&m[1115]&m[1116]&m[1175]));
    m[1122] = (((m[1118]&~m[1119]&~m[1120]&~m[1121]&~m[1185])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1185])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1185])|(m[1118]&m[1119]&~m[1120]&m[1121]&~m[1185])|(m[1118]&~m[1119]&m[1120]&m[1121]&~m[1185])|(~m[1118]&m[1119]&m[1120]&m[1121]&~m[1185]))&BiasedRNG[777])|(((m[1118]&~m[1119]&~m[1120]&~m[1121]&m[1185])|(~m[1118]&m[1119]&~m[1120]&~m[1121]&m[1185])|(~m[1118]&~m[1119]&m[1120]&~m[1121]&m[1185])|(m[1118]&m[1119]&~m[1120]&m[1121]&m[1185])|(m[1118]&~m[1119]&m[1120]&m[1121]&m[1185])|(~m[1118]&m[1119]&m[1120]&m[1121]&m[1185]))&~BiasedRNG[777])|((m[1118]&m[1119]&~m[1120]&~m[1121]&~m[1185])|(m[1118]&~m[1119]&m[1120]&~m[1121]&~m[1185])|(~m[1118]&m[1119]&m[1120]&~m[1121]&~m[1185])|(m[1118]&m[1119]&m[1120]&~m[1121]&~m[1185])|(m[1118]&m[1119]&m[1120]&m[1121]&~m[1185])|(m[1118]&m[1119]&~m[1120]&~m[1121]&m[1185])|(m[1118]&~m[1119]&m[1120]&~m[1121]&m[1185])|(~m[1118]&m[1119]&m[1120]&~m[1121]&m[1185])|(m[1118]&m[1119]&m[1120]&~m[1121]&m[1185])|(m[1118]&m[1119]&m[1120]&m[1121]&m[1185]));
    m[1127] = (((m[1123]&~m[1124]&~m[1125]&~m[1126]&~m[1190])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1190])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1190])|(m[1123]&m[1124]&~m[1125]&m[1126]&~m[1190])|(m[1123]&~m[1124]&m[1125]&m[1126]&~m[1190])|(~m[1123]&m[1124]&m[1125]&m[1126]&~m[1190]))&BiasedRNG[778])|(((m[1123]&~m[1124]&~m[1125]&~m[1126]&m[1190])|(~m[1123]&m[1124]&~m[1125]&~m[1126]&m[1190])|(~m[1123]&~m[1124]&m[1125]&~m[1126]&m[1190])|(m[1123]&m[1124]&~m[1125]&m[1126]&m[1190])|(m[1123]&~m[1124]&m[1125]&m[1126]&m[1190])|(~m[1123]&m[1124]&m[1125]&m[1126]&m[1190]))&~BiasedRNG[778])|((m[1123]&m[1124]&~m[1125]&~m[1126]&~m[1190])|(m[1123]&~m[1124]&m[1125]&~m[1126]&~m[1190])|(~m[1123]&m[1124]&m[1125]&~m[1126]&~m[1190])|(m[1123]&m[1124]&m[1125]&~m[1126]&~m[1190])|(m[1123]&m[1124]&m[1125]&m[1126]&~m[1190])|(m[1123]&m[1124]&~m[1125]&~m[1126]&m[1190])|(m[1123]&~m[1124]&m[1125]&~m[1126]&m[1190])|(~m[1123]&m[1124]&m[1125]&~m[1126]&m[1190])|(m[1123]&m[1124]&m[1125]&~m[1126]&m[1190])|(m[1123]&m[1124]&m[1125]&m[1126]&m[1190]));
    m[1132] = (((m[1128]&~m[1129]&~m[1130]&~m[1131]&~m[1195])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1195])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1195])|(m[1128]&m[1129]&~m[1130]&m[1131]&~m[1195])|(m[1128]&~m[1129]&m[1130]&m[1131]&~m[1195])|(~m[1128]&m[1129]&m[1130]&m[1131]&~m[1195]))&BiasedRNG[779])|(((m[1128]&~m[1129]&~m[1130]&~m[1131]&m[1195])|(~m[1128]&m[1129]&~m[1130]&~m[1131]&m[1195])|(~m[1128]&~m[1129]&m[1130]&~m[1131]&m[1195])|(m[1128]&m[1129]&~m[1130]&m[1131]&m[1195])|(m[1128]&~m[1129]&m[1130]&m[1131]&m[1195])|(~m[1128]&m[1129]&m[1130]&m[1131]&m[1195]))&~BiasedRNG[779])|((m[1128]&m[1129]&~m[1130]&~m[1131]&~m[1195])|(m[1128]&~m[1129]&m[1130]&~m[1131]&~m[1195])|(~m[1128]&m[1129]&m[1130]&~m[1131]&~m[1195])|(m[1128]&m[1129]&m[1130]&~m[1131]&~m[1195])|(m[1128]&m[1129]&m[1130]&m[1131]&~m[1195])|(m[1128]&m[1129]&~m[1130]&~m[1131]&m[1195])|(m[1128]&~m[1129]&m[1130]&~m[1131]&m[1195])|(~m[1128]&m[1129]&m[1130]&~m[1131]&m[1195])|(m[1128]&m[1129]&m[1130]&~m[1131]&m[1195])|(m[1128]&m[1129]&m[1130]&m[1131]&m[1195]));
    m[1137] = (((m[1133]&~m[1134]&~m[1135]&~m[1136]&~m[1200])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1200])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1200])|(m[1133]&m[1134]&~m[1135]&m[1136]&~m[1200])|(m[1133]&~m[1134]&m[1135]&m[1136]&~m[1200])|(~m[1133]&m[1134]&m[1135]&m[1136]&~m[1200]))&BiasedRNG[780])|(((m[1133]&~m[1134]&~m[1135]&~m[1136]&m[1200])|(~m[1133]&m[1134]&~m[1135]&~m[1136]&m[1200])|(~m[1133]&~m[1134]&m[1135]&~m[1136]&m[1200])|(m[1133]&m[1134]&~m[1135]&m[1136]&m[1200])|(m[1133]&~m[1134]&m[1135]&m[1136]&m[1200])|(~m[1133]&m[1134]&m[1135]&m[1136]&m[1200]))&~BiasedRNG[780])|((m[1133]&m[1134]&~m[1135]&~m[1136]&~m[1200])|(m[1133]&~m[1134]&m[1135]&~m[1136]&~m[1200])|(~m[1133]&m[1134]&m[1135]&~m[1136]&~m[1200])|(m[1133]&m[1134]&m[1135]&~m[1136]&~m[1200])|(m[1133]&m[1134]&m[1135]&m[1136]&~m[1200])|(m[1133]&m[1134]&~m[1135]&~m[1136]&m[1200])|(m[1133]&~m[1134]&m[1135]&~m[1136]&m[1200])|(~m[1133]&m[1134]&m[1135]&~m[1136]&m[1200])|(m[1133]&m[1134]&m[1135]&~m[1136]&m[1200])|(m[1133]&m[1134]&m[1135]&m[1136]&m[1200]));
    m[1142] = (((m[1138]&~m[1139]&~m[1140]&~m[1141]&~m[1205])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1205])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1205])|(m[1138]&m[1139]&~m[1140]&m[1141]&~m[1205])|(m[1138]&~m[1139]&m[1140]&m[1141]&~m[1205])|(~m[1138]&m[1139]&m[1140]&m[1141]&~m[1205]))&BiasedRNG[781])|(((m[1138]&~m[1139]&~m[1140]&~m[1141]&m[1205])|(~m[1138]&m[1139]&~m[1140]&~m[1141]&m[1205])|(~m[1138]&~m[1139]&m[1140]&~m[1141]&m[1205])|(m[1138]&m[1139]&~m[1140]&m[1141]&m[1205])|(m[1138]&~m[1139]&m[1140]&m[1141]&m[1205])|(~m[1138]&m[1139]&m[1140]&m[1141]&m[1205]))&~BiasedRNG[781])|((m[1138]&m[1139]&~m[1140]&~m[1141]&~m[1205])|(m[1138]&~m[1139]&m[1140]&~m[1141]&~m[1205])|(~m[1138]&m[1139]&m[1140]&~m[1141]&~m[1205])|(m[1138]&m[1139]&m[1140]&~m[1141]&~m[1205])|(m[1138]&m[1139]&m[1140]&m[1141]&~m[1205])|(m[1138]&m[1139]&~m[1140]&~m[1141]&m[1205])|(m[1138]&~m[1139]&m[1140]&~m[1141]&m[1205])|(~m[1138]&m[1139]&m[1140]&~m[1141]&m[1205])|(m[1138]&m[1139]&m[1140]&~m[1141]&m[1205])|(m[1138]&m[1139]&m[1140]&m[1141]&m[1205]));
    m[1147] = (((m[1143]&~m[1144]&~m[1145]&~m[1146]&~m[1210])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1210])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1210])|(m[1143]&m[1144]&~m[1145]&m[1146]&~m[1210])|(m[1143]&~m[1144]&m[1145]&m[1146]&~m[1210])|(~m[1143]&m[1144]&m[1145]&m[1146]&~m[1210]))&BiasedRNG[782])|(((m[1143]&~m[1144]&~m[1145]&~m[1146]&m[1210])|(~m[1143]&m[1144]&~m[1145]&~m[1146]&m[1210])|(~m[1143]&~m[1144]&m[1145]&~m[1146]&m[1210])|(m[1143]&m[1144]&~m[1145]&m[1146]&m[1210])|(m[1143]&~m[1144]&m[1145]&m[1146]&m[1210])|(~m[1143]&m[1144]&m[1145]&m[1146]&m[1210]))&~BiasedRNG[782])|((m[1143]&m[1144]&~m[1145]&~m[1146]&~m[1210])|(m[1143]&~m[1144]&m[1145]&~m[1146]&~m[1210])|(~m[1143]&m[1144]&m[1145]&~m[1146]&~m[1210])|(m[1143]&m[1144]&m[1145]&~m[1146]&~m[1210])|(m[1143]&m[1144]&m[1145]&m[1146]&~m[1210])|(m[1143]&m[1144]&~m[1145]&~m[1146]&m[1210])|(m[1143]&~m[1144]&m[1145]&~m[1146]&m[1210])|(~m[1143]&m[1144]&m[1145]&~m[1146]&m[1210])|(m[1143]&m[1144]&m[1145]&~m[1146]&m[1210])|(m[1143]&m[1144]&m[1145]&m[1146]&m[1210]));
    m[1152] = (((m[1148]&~m[1149]&~m[1150]&~m[1151]&~m[1215])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1215])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1215])|(m[1148]&m[1149]&~m[1150]&m[1151]&~m[1215])|(m[1148]&~m[1149]&m[1150]&m[1151]&~m[1215])|(~m[1148]&m[1149]&m[1150]&m[1151]&~m[1215]))&BiasedRNG[783])|(((m[1148]&~m[1149]&~m[1150]&~m[1151]&m[1215])|(~m[1148]&m[1149]&~m[1150]&~m[1151]&m[1215])|(~m[1148]&~m[1149]&m[1150]&~m[1151]&m[1215])|(m[1148]&m[1149]&~m[1150]&m[1151]&m[1215])|(m[1148]&~m[1149]&m[1150]&m[1151]&m[1215])|(~m[1148]&m[1149]&m[1150]&m[1151]&m[1215]))&~BiasedRNG[783])|((m[1148]&m[1149]&~m[1150]&~m[1151]&~m[1215])|(m[1148]&~m[1149]&m[1150]&~m[1151]&~m[1215])|(~m[1148]&m[1149]&m[1150]&~m[1151]&~m[1215])|(m[1148]&m[1149]&m[1150]&~m[1151]&~m[1215])|(m[1148]&m[1149]&m[1150]&m[1151]&~m[1215])|(m[1148]&m[1149]&~m[1150]&~m[1151]&m[1215])|(m[1148]&~m[1149]&m[1150]&~m[1151]&m[1215])|(~m[1148]&m[1149]&m[1150]&~m[1151]&m[1215])|(m[1148]&m[1149]&m[1150]&~m[1151]&m[1215])|(m[1148]&m[1149]&m[1150]&m[1151]&m[1215]));
    m[1157] = (((m[1153]&~m[1154]&~m[1155]&~m[1156]&~m[1220])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1220])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1220])|(m[1153]&m[1154]&~m[1155]&m[1156]&~m[1220])|(m[1153]&~m[1154]&m[1155]&m[1156]&~m[1220])|(~m[1153]&m[1154]&m[1155]&m[1156]&~m[1220]))&BiasedRNG[784])|(((m[1153]&~m[1154]&~m[1155]&~m[1156]&m[1220])|(~m[1153]&m[1154]&~m[1155]&~m[1156]&m[1220])|(~m[1153]&~m[1154]&m[1155]&~m[1156]&m[1220])|(m[1153]&m[1154]&~m[1155]&m[1156]&m[1220])|(m[1153]&~m[1154]&m[1155]&m[1156]&m[1220])|(~m[1153]&m[1154]&m[1155]&m[1156]&m[1220]))&~BiasedRNG[784])|((m[1153]&m[1154]&~m[1155]&~m[1156]&~m[1220])|(m[1153]&~m[1154]&m[1155]&~m[1156]&~m[1220])|(~m[1153]&m[1154]&m[1155]&~m[1156]&~m[1220])|(m[1153]&m[1154]&m[1155]&~m[1156]&~m[1220])|(m[1153]&m[1154]&m[1155]&m[1156]&~m[1220])|(m[1153]&m[1154]&~m[1155]&~m[1156]&m[1220])|(m[1153]&~m[1154]&m[1155]&~m[1156]&m[1220])|(~m[1153]&m[1154]&m[1155]&~m[1156]&m[1220])|(m[1153]&m[1154]&m[1155]&~m[1156]&m[1220])|(m[1153]&m[1154]&m[1155]&m[1156]&m[1220]));
    m[1162] = (((m[1158]&~m[1159]&~m[1160]&~m[1161]&~m[1225])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1225])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1225])|(m[1158]&m[1159]&~m[1160]&m[1161]&~m[1225])|(m[1158]&~m[1159]&m[1160]&m[1161]&~m[1225])|(~m[1158]&m[1159]&m[1160]&m[1161]&~m[1225]))&BiasedRNG[785])|(((m[1158]&~m[1159]&~m[1160]&~m[1161]&m[1225])|(~m[1158]&m[1159]&~m[1160]&~m[1161]&m[1225])|(~m[1158]&~m[1159]&m[1160]&~m[1161]&m[1225])|(m[1158]&m[1159]&~m[1160]&m[1161]&m[1225])|(m[1158]&~m[1159]&m[1160]&m[1161]&m[1225])|(~m[1158]&m[1159]&m[1160]&m[1161]&m[1225]))&~BiasedRNG[785])|((m[1158]&m[1159]&~m[1160]&~m[1161]&~m[1225])|(m[1158]&~m[1159]&m[1160]&~m[1161]&~m[1225])|(~m[1158]&m[1159]&m[1160]&~m[1161]&~m[1225])|(m[1158]&m[1159]&m[1160]&~m[1161]&~m[1225])|(m[1158]&m[1159]&m[1160]&m[1161]&~m[1225])|(m[1158]&m[1159]&~m[1160]&~m[1161]&m[1225])|(m[1158]&~m[1159]&m[1160]&~m[1161]&m[1225])|(~m[1158]&m[1159]&m[1160]&~m[1161]&m[1225])|(m[1158]&m[1159]&m[1160]&~m[1161]&m[1225])|(m[1158]&m[1159]&m[1160]&m[1161]&m[1225]));
    m[1167] = (((m[1163]&~m[1164]&~m[1165]&~m[1166]&~m[1230])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1230])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1230])|(m[1163]&m[1164]&~m[1165]&m[1166]&~m[1230])|(m[1163]&~m[1164]&m[1165]&m[1166]&~m[1230])|(~m[1163]&m[1164]&m[1165]&m[1166]&~m[1230]))&BiasedRNG[786])|(((m[1163]&~m[1164]&~m[1165]&~m[1166]&m[1230])|(~m[1163]&m[1164]&~m[1165]&~m[1166]&m[1230])|(~m[1163]&~m[1164]&m[1165]&~m[1166]&m[1230])|(m[1163]&m[1164]&~m[1165]&m[1166]&m[1230])|(m[1163]&~m[1164]&m[1165]&m[1166]&m[1230])|(~m[1163]&m[1164]&m[1165]&m[1166]&m[1230]))&~BiasedRNG[786])|((m[1163]&m[1164]&~m[1165]&~m[1166]&~m[1230])|(m[1163]&~m[1164]&m[1165]&~m[1166]&~m[1230])|(~m[1163]&m[1164]&m[1165]&~m[1166]&~m[1230])|(m[1163]&m[1164]&m[1165]&~m[1166]&~m[1230])|(m[1163]&m[1164]&m[1165]&m[1166]&~m[1230])|(m[1163]&m[1164]&~m[1165]&~m[1166]&m[1230])|(m[1163]&~m[1164]&m[1165]&~m[1166]&m[1230])|(~m[1163]&m[1164]&m[1165]&~m[1166]&m[1230])|(m[1163]&m[1164]&m[1165]&~m[1166]&m[1230])|(m[1163]&m[1164]&m[1165]&m[1166]&m[1230]));
    m[1172] = (((m[1168]&~m[1169]&~m[1170]&~m[1171]&~m[1235])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1235])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1235])|(m[1168]&m[1169]&~m[1170]&m[1171]&~m[1235])|(m[1168]&~m[1169]&m[1170]&m[1171]&~m[1235])|(~m[1168]&m[1169]&m[1170]&m[1171]&~m[1235]))&BiasedRNG[787])|(((m[1168]&~m[1169]&~m[1170]&~m[1171]&m[1235])|(~m[1168]&m[1169]&~m[1170]&~m[1171]&m[1235])|(~m[1168]&~m[1169]&m[1170]&~m[1171]&m[1235])|(m[1168]&m[1169]&~m[1170]&m[1171]&m[1235])|(m[1168]&~m[1169]&m[1170]&m[1171]&m[1235])|(~m[1168]&m[1169]&m[1170]&m[1171]&m[1235]))&~BiasedRNG[787])|((m[1168]&m[1169]&~m[1170]&~m[1171]&~m[1235])|(m[1168]&~m[1169]&m[1170]&~m[1171]&~m[1235])|(~m[1168]&m[1169]&m[1170]&~m[1171]&~m[1235])|(m[1168]&m[1169]&m[1170]&~m[1171]&~m[1235])|(m[1168]&m[1169]&m[1170]&m[1171]&~m[1235])|(m[1168]&m[1169]&~m[1170]&~m[1171]&m[1235])|(m[1168]&~m[1169]&m[1170]&~m[1171]&m[1235])|(~m[1168]&m[1169]&m[1170]&~m[1171]&m[1235])|(m[1168]&m[1169]&m[1170]&~m[1171]&m[1235])|(m[1168]&m[1169]&m[1170]&m[1171]&m[1235]));
    m[1177] = (((m[1173]&~m[1174]&~m[1175]&~m[1176]&~m[1240])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1240])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1240])|(m[1173]&m[1174]&~m[1175]&m[1176]&~m[1240])|(m[1173]&~m[1174]&m[1175]&m[1176]&~m[1240])|(~m[1173]&m[1174]&m[1175]&m[1176]&~m[1240]))&BiasedRNG[788])|(((m[1173]&~m[1174]&~m[1175]&~m[1176]&m[1240])|(~m[1173]&m[1174]&~m[1175]&~m[1176]&m[1240])|(~m[1173]&~m[1174]&m[1175]&~m[1176]&m[1240])|(m[1173]&m[1174]&~m[1175]&m[1176]&m[1240])|(m[1173]&~m[1174]&m[1175]&m[1176]&m[1240])|(~m[1173]&m[1174]&m[1175]&m[1176]&m[1240]))&~BiasedRNG[788])|((m[1173]&m[1174]&~m[1175]&~m[1176]&~m[1240])|(m[1173]&~m[1174]&m[1175]&~m[1176]&~m[1240])|(~m[1173]&m[1174]&m[1175]&~m[1176]&~m[1240])|(m[1173]&m[1174]&m[1175]&~m[1176]&~m[1240])|(m[1173]&m[1174]&m[1175]&m[1176]&~m[1240])|(m[1173]&m[1174]&~m[1175]&~m[1176]&m[1240])|(m[1173]&~m[1174]&m[1175]&~m[1176]&m[1240])|(~m[1173]&m[1174]&m[1175]&~m[1176]&m[1240])|(m[1173]&m[1174]&m[1175]&~m[1176]&m[1240])|(m[1173]&m[1174]&m[1175]&m[1176]&m[1240]));
    m[1182] = (((m[1178]&~m[1179]&~m[1180]&~m[1181]&~m[1245])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1245])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1245])|(m[1178]&m[1179]&~m[1180]&m[1181]&~m[1245])|(m[1178]&~m[1179]&m[1180]&m[1181]&~m[1245])|(~m[1178]&m[1179]&m[1180]&m[1181]&~m[1245]))&BiasedRNG[789])|(((m[1178]&~m[1179]&~m[1180]&~m[1181]&m[1245])|(~m[1178]&m[1179]&~m[1180]&~m[1181]&m[1245])|(~m[1178]&~m[1179]&m[1180]&~m[1181]&m[1245])|(m[1178]&m[1179]&~m[1180]&m[1181]&m[1245])|(m[1178]&~m[1179]&m[1180]&m[1181]&m[1245])|(~m[1178]&m[1179]&m[1180]&m[1181]&m[1245]))&~BiasedRNG[789])|((m[1178]&m[1179]&~m[1180]&~m[1181]&~m[1245])|(m[1178]&~m[1179]&m[1180]&~m[1181]&~m[1245])|(~m[1178]&m[1179]&m[1180]&~m[1181]&~m[1245])|(m[1178]&m[1179]&m[1180]&~m[1181]&~m[1245])|(m[1178]&m[1179]&m[1180]&m[1181]&~m[1245])|(m[1178]&m[1179]&~m[1180]&~m[1181]&m[1245])|(m[1178]&~m[1179]&m[1180]&~m[1181]&m[1245])|(~m[1178]&m[1179]&m[1180]&~m[1181]&m[1245])|(m[1178]&m[1179]&m[1180]&~m[1181]&m[1245])|(m[1178]&m[1179]&m[1180]&m[1181]&m[1245]));
    m[1187] = (((m[1183]&~m[1184]&~m[1185]&~m[1186]&~m[1248])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1248])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1248])|(m[1183]&m[1184]&~m[1185]&m[1186]&~m[1248])|(m[1183]&~m[1184]&m[1185]&m[1186]&~m[1248])|(~m[1183]&m[1184]&m[1185]&m[1186]&~m[1248]))&BiasedRNG[790])|(((m[1183]&~m[1184]&~m[1185]&~m[1186]&m[1248])|(~m[1183]&m[1184]&~m[1185]&~m[1186]&m[1248])|(~m[1183]&~m[1184]&m[1185]&~m[1186]&m[1248])|(m[1183]&m[1184]&~m[1185]&m[1186]&m[1248])|(m[1183]&~m[1184]&m[1185]&m[1186]&m[1248])|(~m[1183]&m[1184]&m[1185]&m[1186]&m[1248]))&~BiasedRNG[790])|((m[1183]&m[1184]&~m[1185]&~m[1186]&~m[1248])|(m[1183]&~m[1184]&m[1185]&~m[1186]&~m[1248])|(~m[1183]&m[1184]&m[1185]&~m[1186]&~m[1248])|(m[1183]&m[1184]&m[1185]&~m[1186]&~m[1248])|(m[1183]&m[1184]&m[1185]&m[1186]&~m[1248])|(m[1183]&m[1184]&~m[1185]&~m[1186]&m[1248])|(m[1183]&~m[1184]&m[1185]&~m[1186]&m[1248])|(~m[1183]&m[1184]&m[1185]&~m[1186]&m[1248])|(m[1183]&m[1184]&m[1185]&~m[1186]&m[1248])|(m[1183]&m[1184]&m[1185]&m[1186]&m[1248]));
    m[1192] = (((m[1188]&~m[1189]&~m[1190]&~m[1191]&~m[1250])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1250])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1250])|(m[1188]&m[1189]&~m[1190]&m[1191]&~m[1250])|(m[1188]&~m[1189]&m[1190]&m[1191]&~m[1250])|(~m[1188]&m[1189]&m[1190]&m[1191]&~m[1250]))&BiasedRNG[791])|(((m[1188]&~m[1189]&~m[1190]&~m[1191]&m[1250])|(~m[1188]&m[1189]&~m[1190]&~m[1191]&m[1250])|(~m[1188]&~m[1189]&m[1190]&~m[1191]&m[1250])|(m[1188]&m[1189]&~m[1190]&m[1191]&m[1250])|(m[1188]&~m[1189]&m[1190]&m[1191]&m[1250])|(~m[1188]&m[1189]&m[1190]&m[1191]&m[1250]))&~BiasedRNG[791])|((m[1188]&m[1189]&~m[1190]&~m[1191]&~m[1250])|(m[1188]&~m[1189]&m[1190]&~m[1191]&~m[1250])|(~m[1188]&m[1189]&m[1190]&~m[1191]&~m[1250])|(m[1188]&m[1189]&m[1190]&~m[1191]&~m[1250])|(m[1188]&m[1189]&m[1190]&m[1191]&~m[1250])|(m[1188]&m[1189]&~m[1190]&~m[1191]&m[1250])|(m[1188]&~m[1189]&m[1190]&~m[1191]&m[1250])|(~m[1188]&m[1189]&m[1190]&~m[1191]&m[1250])|(m[1188]&m[1189]&m[1190]&~m[1191]&m[1250])|(m[1188]&m[1189]&m[1190]&m[1191]&m[1250]));
    m[1197] = (((m[1193]&~m[1194]&~m[1195]&~m[1196]&~m[1255])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1255])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1255])|(m[1193]&m[1194]&~m[1195]&m[1196]&~m[1255])|(m[1193]&~m[1194]&m[1195]&m[1196]&~m[1255])|(~m[1193]&m[1194]&m[1195]&m[1196]&~m[1255]))&BiasedRNG[792])|(((m[1193]&~m[1194]&~m[1195]&~m[1196]&m[1255])|(~m[1193]&m[1194]&~m[1195]&~m[1196]&m[1255])|(~m[1193]&~m[1194]&m[1195]&~m[1196]&m[1255])|(m[1193]&m[1194]&~m[1195]&m[1196]&m[1255])|(m[1193]&~m[1194]&m[1195]&m[1196]&m[1255])|(~m[1193]&m[1194]&m[1195]&m[1196]&m[1255]))&~BiasedRNG[792])|((m[1193]&m[1194]&~m[1195]&~m[1196]&~m[1255])|(m[1193]&~m[1194]&m[1195]&~m[1196]&~m[1255])|(~m[1193]&m[1194]&m[1195]&~m[1196]&~m[1255])|(m[1193]&m[1194]&m[1195]&~m[1196]&~m[1255])|(m[1193]&m[1194]&m[1195]&m[1196]&~m[1255])|(m[1193]&m[1194]&~m[1195]&~m[1196]&m[1255])|(m[1193]&~m[1194]&m[1195]&~m[1196]&m[1255])|(~m[1193]&m[1194]&m[1195]&~m[1196]&m[1255])|(m[1193]&m[1194]&m[1195]&~m[1196]&m[1255])|(m[1193]&m[1194]&m[1195]&m[1196]&m[1255]));
    m[1202] = (((m[1198]&~m[1199]&~m[1200]&~m[1201]&~m[1260])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1260])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1260])|(m[1198]&m[1199]&~m[1200]&m[1201]&~m[1260])|(m[1198]&~m[1199]&m[1200]&m[1201]&~m[1260])|(~m[1198]&m[1199]&m[1200]&m[1201]&~m[1260]))&BiasedRNG[793])|(((m[1198]&~m[1199]&~m[1200]&~m[1201]&m[1260])|(~m[1198]&m[1199]&~m[1200]&~m[1201]&m[1260])|(~m[1198]&~m[1199]&m[1200]&~m[1201]&m[1260])|(m[1198]&m[1199]&~m[1200]&m[1201]&m[1260])|(m[1198]&~m[1199]&m[1200]&m[1201]&m[1260])|(~m[1198]&m[1199]&m[1200]&m[1201]&m[1260]))&~BiasedRNG[793])|((m[1198]&m[1199]&~m[1200]&~m[1201]&~m[1260])|(m[1198]&~m[1199]&m[1200]&~m[1201]&~m[1260])|(~m[1198]&m[1199]&m[1200]&~m[1201]&~m[1260])|(m[1198]&m[1199]&m[1200]&~m[1201]&~m[1260])|(m[1198]&m[1199]&m[1200]&m[1201]&~m[1260])|(m[1198]&m[1199]&~m[1200]&~m[1201]&m[1260])|(m[1198]&~m[1199]&m[1200]&~m[1201]&m[1260])|(~m[1198]&m[1199]&m[1200]&~m[1201]&m[1260])|(m[1198]&m[1199]&m[1200]&~m[1201]&m[1260])|(m[1198]&m[1199]&m[1200]&m[1201]&m[1260]));
    m[1207] = (((m[1203]&~m[1204]&~m[1205]&~m[1206]&~m[1265])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1265])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1265])|(m[1203]&m[1204]&~m[1205]&m[1206]&~m[1265])|(m[1203]&~m[1204]&m[1205]&m[1206]&~m[1265])|(~m[1203]&m[1204]&m[1205]&m[1206]&~m[1265]))&BiasedRNG[794])|(((m[1203]&~m[1204]&~m[1205]&~m[1206]&m[1265])|(~m[1203]&m[1204]&~m[1205]&~m[1206]&m[1265])|(~m[1203]&~m[1204]&m[1205]&~m[1206]&m[1265])|(m[1203]&m[1204]&~m[1205]&m[1206]&m[1265])|(m[1203]&~m[1204]&m[1205]&m[1206]&m[1265])|(~m[1203]&m[1204]&m[1205]&m[1206]&m[1265]))&~BiasedRNG[794])|((m[1203]&m[1204]&~m[1205]&~m[1206]&~m[1265])|(m[1203]&~m[1204]&m[1205]&~m[1206]&~m[1265])|(~m[1203]&m[1204]&m[1205]&~m[1206]&~m[1265])|(m[1203]&m[1204]&m[1205]&~m[1206]&~m[1265])|(m[1203]&m[1204]&m[1205]&m[1206]&~m[1265])|(m[1203]&m[1204]&~m[1205]&~m[1206]&m[1265])|(m[1203]&~m[1204]&m[1205]&~m[1206]&m[1265])|(~m[1203]&m[1204]&m[1205]&~m[1206]&m[1265])|(m[1203]&m[1204]&m[1205]&~m[1206]&m[1265])|(m[1203]&m[1204]&m[1205]&m[1206]&m[1265]));
    m[1212] = (((m[1208]&~m[1209]&~m[1210]&~m[1211]&~m[1270])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1270])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1270])|(m[1208]&m[1209]&~m[1210]&m[1211]&~m[1270])|(m[1208]&~m[1209]&m[1210]&m[1211]&~m[1270])|(~m[1208]&m[1209]&m[1210]&m[1211]&~m[1270]))&BiasedRNG[795])|(((m[1208]&~m[1209]&~m[1210]&~m[1211]&m[1270])|(~m[1208]&m[1209]&~m[1210]&~m[1211]&m[1270])|(~m[1208]&~m[1209]&m[1210]&~m[1211]&m[1270])|(m[1208]&m[1209]&~m[1210]&m[1211]&m[1270])|(m[1208]&~m[1209]&m[1210]&m[1211]&m[1270])|(~m[1208]&m[1209]&m[1210]&m[1211]&m[1270]))&~BiasedRNG[795])|((m[1208]&m[1209]&~m[1210]&~m[1211]&~m[1270])|(m[1208]&~m[1209]&m[1210]&~m[1211]&~m[1270])|(~m[1208]&m[1209]&m[1210]&~m[1211]&~m[1270])|(m[1208]&m[1209]&m[1210]&~m[1211]&~m[1270])|(m[1208]&m[1209]&m[1210]&m[1211]&~m[1270])|(m[1208]&m[1209]&~m[1210]&~m[1211]&m[1270])|(m[1208]&~m[1209]&m[1210]&~m[1211]&m[1270])|(~m[1208]&m[1209]&m[1210]&~m[1211]&m[1270])|(m[1208]&m[1209]&m[1210]&~m[1211]&m[1270])|(m[1208]&m[1209]&m[1210]&m[1211]&m[1270]));
    m[1217] = (((m[1213]&~m[1214]&~m[1215]&~m[1216]&~m[1275])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1275])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1275])|(m[1213]&m[1214]&~m[1215]&m[1216]&~m[1275])|(m[1213]&~m[1214]&m[1215]&m[1216]&~m[1275])|(~m[1213]&m[1214]&m[1215]&m[1216]&~m[1275]))&BiasedRNG[796])|(((m[1213]&~m[1214]&~m[1215]&~m[1216]&m[1275])|(~m[1213]&m[1214]&~m[1215]&~m[1216]&m[1275])|(~m[1213]&~m[1214]&m[1215]&~m[1216]&m[1275])|(m[1213]&m[1214]&~m[1215]&m[1216]&m[1275])|(m[1213]&~m[1214]&m[1215]&m[1216]&m[1275])|(~m[1213]&m[1214]&m[1215]&m[1216]&m[1275]))&~BiasedRNG[796])|((m[1213]&m[1214]&~m[1215]&~m[1216]&~m[1275])|(m[1213]&~m[1214]&m[1215]&~m[1216]&~m[1275])|(~m[1213]&m[1214]&m[1215]&~m[1216]&~m[1275])|(m[1213]&m[1214]&m[1215]&~m[1216]&~m[1275])|(m[1213]&m[1214]&m[1215]&m[1216]&~m[1275])|(m[1213]&m[1214]&~m[1215]&~m[1216]&m[1275])|(m[1213]&~m[1214]&m[1215]&~m[1216]&m[1275])|(~m[1213]&m[1214]&m[1215]&~m[1216]&m[1275])|(m[1213]&m[1214]&m[1215]&~m[1216]&m[1275])|(m[1213]&m[1214]&m[1215]&m[1216]&m[1275]));
    m[1222] = (((m[1218]&~m[1219]&~m[1220]&~m[1221]&~m[1280])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1280])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1280])|(m[1218]&m[1219]&~m[1220]&m[1221]&~m[1280])|(m[1218]&~m[1219]&m[1220]&m[1221]&~m[1280])|(~m[1218]&m[1219]&m[1220]&m[1221]&~m[1280]))&BiasedRNG[797])|(((m[1218]&~m[1219]&~m[1220]&~m[1221]&m[1280])|(~m[1218]&m[1219]&~m[1220]&~m[1221]&m[1280])|(~m[1218]&~m[1219]&m[1220]&~m[1221]&m[1280])|(m[1218]&m[1219]&~m[1220]&m[1221]&m[1280])|(m[1218]&~m[1219]&m[1220]&m[1221]&m[1280])|(~m[1218]&m[1219]&m[1220]&m[1221]&m[1280]))&~BiasedRNG[797])|((m[1218]&m[1219]&~m[1220]&~m[1221]&~m[1280])|(m[1218]&~m[1219]&m[1220]&~m[1221]&~m[1280])|(~m[1218]&m[1219]&m[1220]&~m[1221]&~m[1280])|(m[1218]&m[1219]&m[1220]&~m[1221]&~m[1280])|(m[1218]&m[1219]&m[1220]&m[1221]&~m[1280])|(m[1218]&m[1219]&~m[1220]&~m[1221]&m[1280])|(m[1218]&~m[1219]&m[1220]&~m[1221]&m[1280])|(~m[1218]&m[1219]&m[1220]&~m[1221]&m[1280])|(m[1218]&m[1219]&m[1220]&~m[1221]&m[1280])|(m[1218]&m[1219]&m[1220]&m[1221]&m[1280]));
    m[1227] = (((m[1223]&~m[1224]&~m[1225]&~m[1226]&~m[1285])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1285])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1285])|(m[1223]&m[1224]&~m[1225]&m[1226]&~m[1285])|(m[1223]&~m[1224]&m[1225]&m[1226]&~m[1285])|(~m[1223]&m[1224]&m[1225]&m[1226]&~m[1285]))&BiasedRNG[798])|(((m[1223]&~m[1224]&~m[1225]&~m[1226]&m[1285])|(~m[1223]&m[1224]&~m[1225]&~m[1226]&m[1285])|(~m[1223]&~m[1224]&m[1225]&~m[1226]&m[1285])|(m[1223]&m[1224]&~m[1225]&m[1226]&m[1285])|(m[1223]&~m[1224]&m[1225]&m[1226]&m[1285])|(~m[1223]&m[1224]&m[1225]&m[1226]&m[1285]))&~BiasedRNG[798])|((m[1223]&m[1224]&~m[1225]&~m[1226]&~m[1285])|(m[1223]&~m[1224]&m[1225]&~m[1226]&~m[1285])|(~m[1223]&m[1224]&m[1225]&~m[1226]&~m[1285])|(m[1223]&m[1224]&m[1225]&~m[1226]&~m[1285])|(m[1223]&m[1224]&m[1225]&m[1226]&~m[1285])|(m[1223]&m[1224]&~m[1225]&~m[1226]&m[1285])|(m[1223]&~m[1224]&m[1225]&~m[1226]&m[1285])|(~m[1223]&m[1224]&m[1225]&~m[1226]&m[1285])|(m[1223]&m[1224]&m[1225]&~m[1226]&m[1285])|(m[1223]&m[1224]&m[1225]&m[1226]&m[1285]));
    m[1232] = (((m[1228]&~m[1229]&~m[1230]&~m[1231]&~m[1290])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1290])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1290])|(m[1228]&m[1229]&~m[1230]&m[1231]&~m[1290])|(m[1228]&~m[1229]&m[1230]&m[1231]&~m[1290])|(~m[1228]&m[1229]&m[1230]&m[1231]&~m[1290]))&BiasedRNG[799])|(((m[1228]&~m[1229]&~m[1230]&~m[1231]&m[1290])|(~m[1228]&m[1229]&~m[1230]&~m[1231]&m[1290])|(~m[1228]&~m[1229]&m[1230]&~m[1231]&m[1290])|(m[1228]&m[1229]&~m[1230]&m[1231]&m[1290])|(m[1228]&~m[1229]&m[1230]&m[1231]&m[1290])|(~m[1228]&m[1229]&m[1230]&m[1231]&m[1290]))&~BiasedRNG[799])|((m[1228]&m[1229]&~m[1230]&~m[1231]&~m[1290])|(m[1228]&~m[1229]&m[1230]&~m[1231]&~m[1290])|(~m[1228]&m[1229]&m[1230]&~m[1231]&~m[1290])|(m[1228]&m[1229]&m[1230]&~m[1231]&~m[1290])|(m[1228]&m[1229]&m[1230]&m[1231]&~m[1290])|(m[1228]&m[1229]&~m[1230]&~m[1231]&m[1290])|(m[1228]&~m[1229]&m[1230]&~m[1231]&m[1290])|(~m[1228]&m[1229]&m[1230]&~m[1231]&m[1290])|(m[1228]&m[1229]&m[1230]&~m[1231]&m[1290])|(m[1228]&m[1229]&m[1230]&m[1231]&m[1290]));
    m[1237] = (((m[1233]&~m[1234]&~m[1235]&~m[1236]&~m[1295])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1295])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1295])|(m[1233]&m[1234]&~m[1235]&m[1236]&~m[1295])|(m[1233]&~m[1234]&m[1235]&m[1236]&~m[1295])|(~m[1233]&m[1234]&m[1235]&m[1236]&~m[1295]))&BiasedRNG[800])|(((m[1233]&~m[1234]&~m[1235]&~m[1236]&m[1295])|(~m[1233]&m[1234]&~m[1235]&~m[1236]&m[1295])|(~m[1233]&~m[1234]&m[1235]&~m[1236]&m[1295])|(m[1233]&m[1234]&~m[1235]&m[1236]&m[1295])|(m[1233]&~m[1234]&m[1235]&m[1236]&m[1295])|(~m[1233]&m[1234]&m[1235]&m[1236]&m[1295]))&~BiasedRNG[800])|((m[1233]&m[1234]&~m[1235]&~m[1236]&~m[1295])|(m[1233]&~m[1234]&m[1235]&~m[1236]&~m[1295])|(~m[1233]&m[1234]&m[1235]&~m[1236]&~m[1295])|(m[1233]&m[1234]&m[1235]&~m[1236]&~m[1295])|(m[1233]&m[1234]&m[1235]&m[1236]&~m[1295])|(m[1233]&m[1234]&~m[1235]&~m[1236]&m[1295])|(m[1233]&~m[1234]&m[1235]&~m[1236]&m[1295])|(~m[1233]&m[1234]&m[1235]&~m[1236]&m[1295])|(m[1233]&m[1234]&m[1235]&~m[1236]&m[1295])|(m[1233]&m[1234]&m[1235]&m[1236]&m[1295]));
    m[1242] = (((m[1238]&~m[1239]&~m[1240]&~m[1241]&~m[1300])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1300])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1300])|(m[1238]&m[1239]&~m[1240]&m[1241]&~m[1300])|(m[1238]&~m[1239]&m[1240]&m[1241]&~m[1300])|(~m[1238]&m[1239]&m[1240]&m[1241]&~m[1300]))&BiasedRNG[801])|(((m[1238]&~m[1239]&~m[1240]&~m[1241]&m[1300])|(~m[1238]&m[1239]&~m[1240]&~m[1241]&m[1300])|(~m[1238]&~m[1239]&m[1240]&~m[1241]&m[1300])|(m[1238]&m[1239]&~m[1240]&m[1241]&m[1300])|(m[1238]&~m[1239]&m[1240]&m[1241]&m[1300])|(~m[1238]&m[1239]&m[1240]&m[1241]&m[1300]))&~BiasedRNG[801])|((m[1238]&m[1239]&~m[1240]&~m[1241]&~m[1300])|(m[1238]&~m[1239]&m[1240]&~m[1241]&~m[1300])|(~m[1238]&m[1239]&m[1240]&~m[1241]&~m[1300])|(m[1238]&m[1239]&m[1240]&~m[1241]&~m[1300])|(m[1238]&m[1239]&m[1240]&m[1241]&~m[1300])|(m[1238]&m[1239]&~m[1240]&~m[1241]&m[1300])|(m[1238]&~m[1239]&m[1240]&~m[1241]&m[1300])|(~m[1238]&m[1239]&m[1240]&~m[1241]&m[1300])|(m[1238]&m[1239]&m[1240]&~m[1241]&m[1300])|(m[1238]&m[1239]&m[1240]&m[1241]&m[1300]));
    m[1247] = (((m[1243]&~m[1244]&~m[1245]&~m[1246]&~m[1305])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1305])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1305])|(m[1243]&m[1244]&~m[1245]&m[1246]&~m[1305])|(m[1243]&~m[1244]&m[1245]&m[1246]&~m[1305])|(~m[1243]&m[1244]&m[1245]&m[1246]&~m[1305]))&BiasedRNG[802])|(((m[1243]&~m[1244]&~m[1245]&~m[1246]&m[1305])|(~m[1243]&m[1244]&~m[1245]&~m[1246]&m[1305])|(~m[1243]&~m[1244]&m[1245]&~m[1246]&m[1305])|(m[1243]&m[1244]&~m[1245]&m[1246]&m[1305])|(m[1243]&~m[1244]&m[1245]&m[1246]&m[1305])|(~m[1243]&m[1244]&m[1245]&m[1246]&m[1305]))&~BiasedRNG[802])|((m[1243]&m[1244]&~m[1245]&~m[1246]&~m[1305])|(m[1243]&~m[1244]&m[1245]&~m[1246]&~m[1305])|(~m[1243]&m[1244]&m[1245]&~m[1246]&~m[1305])|(m[1243]&m[1244]&m[1245]&~m[1246]&~m[1305])|(m[1243]&m[1244]&m[1245]&m[1246]&~m[1305])|(m[1243]&m[1244]&~m[1245]&~m[1246]&m[1305])|(m[1243]&~m[1244]&m[1245]&~m[1246]&m[1305])|(~m[1243]&m[1244]&m[1245]&~m[1246]&m[1305])|(m[1243]&m[1244]&m[1245]&~m[1246]&m[1305])|(m[1243]&m[1244]&m[1245]&m[1246]&m[1305]));
    m[1252] = (((m[1248]&~m[1249]&~m[1250]&~m[1251]&~m[1308])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1308])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1308])|(m[1248]&m[1249]&~m[1250]&m[1251]&~m[1308])|(m[1248]&~m[1249]&m[1250]&m[1251]&~m[1308])|(~m[1248]&m[1249]&m[1250]&m[1251]&~m[1308]))&BiasedRNG[803])|(((m[1248]&~m[1249]&~m[1250]&~m[1251]&m[1308])|(~m[1248]&m[1249]&~m[1250]&~m[1251]&m[1308])|(~m[1248]&~m[1249]&m[1250]&~m[1251]&m[1308])|(m[1248]&m[1249]&~m[1250]&m[1251]&m[1308])|(m[1248]&~m[1249]&m[1250]&m[1251]&m[1308])|(~m[1248]&m[1249]&m[1250]&m[1251]&m[1308]))&~BiasedRNG[803])|((m[1248]&m[1249]&~m[1250]&~m[1251]&~m[1308])|(m[1248]&~m[1249]&m[1250]&~m[1251]&~m[1308])|(~m[1248]&m[1249]&m[1250]&~m[1251]&~m[1308])|(m[1248]&m[1249]&m[1250]&~m[1251]&~m[1308])|(m[1248]&m[1249]&m[1250]&m[1251]&~m[1308])|(m[1248]&m[1249]&~m[1250]&~m[1251]&m[1308])|(m[1248]&~m[1249]&m[1250]&~m[1251]&m[1308])|(~m[1248]&m[1249]&m[1250]&~m[1251]&m[1308])|(m[1248]&m[1249]&m[1250]&~m[1251]&m[1308])|(m[1248]&m[1249]&m[1250]&m[1251]&m[1308]));
    m[1257] = (((m[1253]&~m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&~m[1310]))&BiasedRNG[804])|(((m[1253]&~m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(~m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&~m[1255]&m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&m[1256]&m[1310]))&~BiasedRNG[804])|((m[1253]&m[1254]&~m[1255]&~m[1256]&~m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&~m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&~m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&~m[1310])|(m[1253]&m[1254]&~m[1255]&~m[1256]&m[1310])|(m[1253]&~m[1254]&m[1255]&~m[1256]&m[1310])|(~m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&~m[1256]&m[1310])|(m[1253]&m[1254]&m[1255]&m[1256]&m[1310]));
    m[1262] = (((m[1258]&~m[1259]&~m[1260]&~m[1261]&~m[1315])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1315])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1315])|(m[1258]&m[1259]&~m[1260]&m[1261]&~m[1315])|(m[1258]&~m[1259]&m[1260]&m[1261]&~m[1315])|(~m[1258]&m[1259]&m[1260]&m[1261]&~m[1315]))&BiasedRNG[805])|(((m[1258]&~m[1259]&~m[1260]&~m[1261]&m[1315])|(~m[1258]&m[1259]&~m[1260]&~m[1261]&m[1315])|(~m[1258]&~m[1259]&m[1260]&~m[1261]&m[1315])|(m[1258]&m[1259]&~m[1260]&m[1261]&m[1315])|(m[1258]&~m[1259]&m[1260]&m[1261]&m[1315])|(~m[1258]&m[1259]&m[1260]&m[1261]&m[1315]))&~BiasedRNG[805])|((m[1258]&m[1259]&~m[1260]&~m[1261]&~m[1315])|(m[1258]&~m[1259]&m[1260]&~m[1261]&~m[1315])|(~m[1258]&m[1259]&m[1260]&~m[1261]&~m[1315])|(m[1258]&m[1259]&m[1260]&~m[1261]&~m[1315])|(m[1258]&m[1259]&m[1260]&m[1261]&~m[1315])|(m[1258]&m[1259]&~m[1260]&~m[1261]&m[1315])|(m[1258]&~m[1259]&m[1260]&~m[1261]&m[1315])|(~m[1258]&m[1259]&m[1260]&~m[1261]&m[1315])|(m[1258]&m[1259]&m[1260]&~m[1261]&m[1315])|(m[1258]&m[1259]&m[1260]&m[1261]&m[1315]));
    m[1267] = (((m[1263]&~m[1264]&~m[1265]&~m[1266]&~m[1320])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1320])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1320])|(m[1263]&m[1264]&~m[1265]&m[1266]&~m[1320])|(m[1263]&~m[1264]&m[1265]&m[1266]&~m[1320])|(~m[1263]&m[1264]&m[1265]&m[1266]&~m[1320]))&BiasedRNG[806])|(((m[1263]&~m[1264]&~m[1265]&~m[1266]&m[1320])|(~m[1263]&m[1264]&~m[1265]&~m[1266]&m[1320])|(~m[1263]&~m[1264]&m[1265]&~m[1266]&m[1320])|(m[1263]&m[1264]&~m[1265]&m[1266]&m[1320])|(m[1263]&~m[1264]&m[1265]&m[1266]&m[1320])|(~m[1263]&m[1264]&m[1265]&m[1266]&m[1320]))&~BiasedRNG[806])|((m[1263]&m[1264]&~m[1265]&~m[1266]&~m[1320])|(m[1263]&~m[1264]&m[1265]&~m[1266]&~m[1320])|(~m[1263]&m[1264]&m[1265]&~m[1266]&~m[1320])|(m[1263]&m[1264]&m[1265]&~m[1266]&~m[1320])|(m[1263]&m[1264]&m[1265]&m[1266]&~m[1320])|(m[1263]&m[1264]&~m[1265]&~m[1266]&m[1320])|(m[1263]&~m[1264]&m[1265]&~m[1266]&m[1320])|(~m[1263]&m[1264]&m[1265]&~m[1266]&m[1320])|(m[1263]&m[1264]&m[1265]&~m[1266]&m[1320])|(m[1263]&m[1264]&m[1265]&m[1266]&m[1320]));
    m[1272] = (((m[1268]&~m[1269]&~m[1270]&~m[1271]&~m[1325])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1325])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1325])|(m[1268]&m[1269]&~m[1270]&m[1271]&~m[1325])|(m[1268]&~m[1269]&m[1270]&m[1271]&~m[1325])|(~m[1268]&m[1269]&m[1270]&m[1271]&~m[1325]))&BiasedRNG[807])|(((m[1268]&~m[1269]&~m[1270]&~m[1271]&m[1325])|(~m[1268]&m[1269]&~m[1270]&~m[1271]&m[1325])|(~m[1268]&~m[1269]&m[1270]&~m[1271]&m[1325])|(m[1268]&m[1269]&~m[1270]&m[1271]&m[1325])|(m[1268]&~m[1269]&m[1270]&m[1271]&m[1325])|(~m[1268]&m[1269]&m[1270]&m[1271]&m[1325]))&~BiasedRNG[807])|((m[1268]&m[1269]&~m[1270]&~m[1271]&~m[1325])|(m[1268]&~m[1269]&m[1270]&~m[1271]&~m[1325])|(~m[1268]&m[1269]&m[1270]&~m[1271]&~m[1325])|(m[1268]&m[1269]&m[1270]&~m[1271]&~m[1325])|(m[1268]&m[1269]&m[1270]&m[1271]&~m[1325])|(m[1268]&m[1269]&~m[1270]&~m[1271]&m[1325])|(m[1268]&~m[1269]&m[1270]&~m[1271]&m[1325])|(~m[1268]&m[1269]&m[1270]&~m[1271]&m[1325])|(m[1268]&m[1269]&m[1270]&~m[1271]&m[1325])|(m[1268]&m[1269]&m[1270]&m[1271]&m[1325]));
    m[1277] = (((m[1273]&~m[1274]&~m[1275]&~m[1276]&~m[1330])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1330])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1330])|(m[1273]&m[1274]&~m[1275]&m[1276]&~m[1330])|(m[1273]&~m[1274]&m[1275]&m[1276]&~m[1330])|(~m[1273]&m[1274]&m[1275]&m[1276]&~m[1330]))&BiasedRNG[808])|(((m[1273]&~m[1274]&~m[1275]&~m[1276]&m[1330])|(~m[1273]&m[1274]&~m[1275]&~m[1276]&m[1330])|(~m[1273]&~m[1274]&m[1275]&~m[1276]&m[1330])|(m[1273]&m[1274]&~m[1275]&m[1276]&m[1330])|(m[1273]&~m[1274]&m[1275]&m[1276]&m[1330])|(~m[1273]&m[1274]&m[1275]&m[1276]&m[1330]))&~BiasedRNG[808])|((m[1273]&m[1274]&~m[1275]&~m[1276]&~m[1330])|(m[1273]&~m[1274]&m[1275]&~m[1276]&~m[1330])|(~m[1273]&m[1274]&m[1275]&~m[1276]&~m[1330])|(m[1273]&m[1274]&m[1275]&~m[1276]&~m[1330])|(m[1273]&m[1274]&m[1275]&m[1276]&~m[1330])|(m[1273]&m[1274]&~m[1275]&~m[1276]&m[1330])|(m[1273]&~m[1274]&m[1275]&~m[1276]&m[1330])|(~m[1273]&m[1274]&m[1275]&~m[1276]&m[1330])|(m[1273]&m[1274]&m[1275]&~m[1276]&m[1330])|(m[1273]&m[1274]&m[1275]&m[1276]&m[1330]));
    m[1282] = (((m[1278]&~m[1279]&~m[1280]&~m[1281]&~m[1335])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1335])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1335])|(m[1278]&m[1279]&~m[1280]&m[1281]&~m[1335])|(m[1278]&~m[1279]&m[1280]&m[1281]&~m[1335])|(~m[1278]&m[1279]&m[1280]&m[1281]&~m[1335]))&BiasedRNG[809])|(((m[1278]&~m[1279]&~m[1280]&~m[1281]&m[1335])|(~m[1278]&m[1279]&~m[1280]&~m[1281]&m[1335])|(~m[1278]&~m[1279]&m[1280]&~m[1281]&m[1335])|(m[1278]&m[1279]&~m[1280]&m[1281]&m[1335])|(m[1278]&~m[1279]&m[1280]&m[1281]&m[1335])|(~m[1278]&m[1279]&m[1280]&m[1281]&m[1335]))&~BiasedRNG[809])|((m[1278]&m[1279]&~m[1280]&~m[1281]&~m[1335])|(m[1278]&~m[1279]&m[1280]&~m[1281]&~m[1335])|(~m[1278]&m[1279]&m[1280]&~m[1281]&~m[1335])|(m[1278]&m[1279]&m[1280]&~m[1281]&~m[1335])|(m[1278]&m[1279]&m[1280]&m[1281]&~m[1335])|(m[1278]&m[1279]&~m[1280]&~m[1281]&m[1335])|(m[1278]&~m[1279]&m[1280]&~m[1281]&m[1335])|(~m[1278]&m[1279]&m[1280]&~m[1281]&m[1335])|(m[1278]&m[1279]&m[1280]&~m[1281]&m[1335])|(m[1278]&m[1279]&m[1280]&m[1281]&m[1335]));
    m[1287] = (((m[1283]&~m[1284]&~m[1285]&~m[1286]&~m[1340])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1340])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1340])|(m[1283]&m[1284]&~m[1285]&m[1286]&~m[1340])|(m[1283]&~m[1284]&m[1285]&m[1286]&~m[1340])|(~m[1283]&m[1284]&m[1285]&m[1286]&~m[1340]))&BiasedRNG[810])|(((m[1283]&~m[1284]&~m[1285]&~m[1286]&m[1340])|(~m[1283]&m[1284]&~m[1285]&~m[1286]&m[1340])|(~m[1283]&~m[1284]&m[1285]&~m[1286]&m[1340])|(m[1283]&m[1284]&~m[1285]&m[1286]&m[1340])|(m[1283]&~m[1284]&m[1285]&m[1286]&m[1340])|(~m[1283]&m[1284]&m[1285]&m[1286]&m[1340]))&~BiasedRNG[810])|((m[1283]&m[1284]&~m[1285]&~m[1286]&~m[1340])|(m[1283]&~m[1284]&m[1285]&~m[1286]&~m[1340])|(~m[1283]&m[1284]&m[1285]&~m[1286]&~m[1340])|(m[1283]&m[1284]&m[1285]&~m[1286]&~m[1340])|(m[1283]&m[1284]&m[1285]&m[1286]&~m[1340])|(m[1283]&m[1284]&~m[1285]&~m[1286]&m[1340])|(m[1283]&~m[1284]&m[1285]&~m[1286]&m[1340])|(~m[1283]&m[1284]&m[1285]&~m[1286]&m[1340])|(m[1283]&m[1284]&m[1285]&~m[1286]&m[1340])|(m[1283]&m[1284]&m[1285]&m[1286]&m[1340]));
    m[1292] = (((m[1288]&~m[1289]&~m[1290]&~m[1291]&~m[1345])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1345])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1345])|(m[1288]&m[1289]&~m[1290]&m[1291]&~m[1345])|(m[1288]&~m[1289]&m[1290]&m[1291]&~m[1345])|(~m[1288]&m[1289]&m[1290]&m[1291]&~m[1345]))&BiasedRNG[811])|(((m[1288]&~m[1289]&~m[1290]&~m[1291]&m[1345])|(~m[1288]&m[1289]&~m[1290]&~m[1291]&m[1345])|(~m[1288]&~m[1289]&m[1290]&~m[1291]&m[1345])|(m[1288]&m[1289]&~m[1290]&m[1291]&m[1345])|(m[1288]&~m[1289]&m[1290]&m[1291]&m[1345])|(~m[1288]&m[1289]&m[1290]&m[1291]&m[1345]))&~BiasedRNG[811])|((m[1288]&m[1289]&~m[1290]&~m[1291]&~m[1345])|(m[1288]&~m[1289]&m[1290]&~m[1291]&~m[1345])|(~m[1288]&m[1289]&m[1290]&~m[1291]&~m[1345])|(m[1288]&m[1289]&m[1290]&~m[1291]&~m[1345])|(m[1288]&m[1289]&m[1290]&m[1291]&~m[1345])|(m[1288]&m[1289]&~m[1290]&~m[1291]&m[1345])|(m[1288]&~m[1289]&m[1290]&~m[1291]&m[1345])|(~m[1288]&m[1289]&m[1290]&~m[1291]&m[1345])|(m[1288]&m[1289]&m[1290]&~m[1291]&m[1345])|(m[1288]&m[1289]&m[1290]&m[1291]&m[1345]));
    m[1297] = (((m[1293]&~m[1294]&~m[1295]&~m[1296]&~m[1350])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1350])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1350])|(m[1293]&m[1294]&~m[1295]&m[1296]&~m[1350])|(m[1293]&~m[1294]&m[1295]&m[1296]&~m[1350])|(~m[1293]&m[1294]&m[1295]&m[1296]&~m[1350]))&BiasedRNG[812])|(((m[1293]&~m[1294]&~m[1295]&~m[1296]&m[1350])|(~m[1293]&m[1294]&~m[1295]&~m[1296]&m[1350])|(~m[1293]&~m[1294]&m[1295]&~m[1296]&m[1350])|(m[1293]&m[1294]&~m[1295]&m[1296]&m[1350])|(m[1293]&~m[1294]&m[1295]&m[1296]&m[1350])|(~m[1293]&m[1294]&m[1295]&m[1296]&m[1350]))&~BiasedRNG[812])|((m[1293]&m[1294]&~m[1295]&~m[1296]&~m[1350])|(m[1293]&~m[1294]&m[1295]&~m[1296]&~m[1350])|(~m[1293]&m[1294]&m[1295]&~m[1296]&~m[1350])|(m[1293]&m[1294]&m[1295]&~m[1296]&~m[1350])|(m[1293]&m[1294]&m[1295]&m[1296]&~m[1350])|(m[1293]&m[1294]&~m[1295]&~m[1296]&m[1350])|(m[1293]&~m[1294]&m[1295]&~m[1296]&m[1350])|(~m[1293]&m[1294]&m[1295]&~m[1296]&m[1350])|(m[1293]&m[1294]&m[1295]&~m[1296]&m[1350])|(m[1293]&m[1294]&m[1295]&m[1296]&m[1350]));
    m[1302] = (((m[1298]&~m[1299]&~m[1300]&~m[1301]&~m[1355])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1355])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1355])|(m[1298]&m[1299]&~m[1300]&m[1301]&~m[1355])|(m[1298]&~m[1299]&m[1300]&m[1301]&~m[1355])|(~m[1298]&m[1299]&m[1300]&m[1301]&~m[1355]))&BiasedRNG[813])|(((m[1298]&~m[1299]&~m[1300]&~m[1301]&m[1355])|(~m[1298]&m[1299]&~m[1300]&~m[1301]&m[1355])|(~m[1298]&~m[1299]&m[1300]&~m[1301]&m[1355])|(m[1298]&m[1299]&~m[1300]&m[1301]&m[1355])|(m[1298]&~m[1299]&m[1300]&m[1301]&m[1355])|(~m[1298]&m[1299]&m[1300]&m[1301]&m[1355]))&~BiasedRNG[813])|((m[1298]&m[1299]&~m[1300]&~m[1301]&~m[1355])|(m[1298]&~m[1299]&m[1300]&~m[1301]&~m[1355])|(~m[1298]&m[1299]&m[1300]&~m[1301]&~m[1355])|(m[1298]&m[1299]&m[1300]&~m[1301]&~m[1355])|(m[1298]&m[1299]&m[1300]&m[1301]&~m[1355])|(m[1298]&m[1299]&~m[1300]&~m[1301]&m[1355])|(m[1298]&~m[1299]&m[1300]&~m[1301]&m[1355])|(~m[1298]&m[1299]&m[1300]&~m[1301]&m[1355])|(m[1298]&m[1299]&m[1300]&~m[1301]&m[1355])|(m[1298]&m[1299]&m[1300]&m[1301]&m[1355]));
    m[1307] = (((m[1303]&~m[1304]&~m[1305]&~m[1306]&~m[1360])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1360])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1360])|(m[1303]&m[1304]&~m[1305]&m[1306]&~m[1360])|(m[1303]&~m[1304]&m[1305]&m[1306]&~m[1360])|(~m[1303]&m[1304]&m[1305]&m[1306]&~m[1360]))&BiasedRNG[814])|(((m[1303]&~m[1304]&~m[1305]&~m[1306]&m[1360])|(~m[1303]&m[1304]&~m[1305]&~m[1306]&m[1360])|(~m[1303]&~m[1304]&m[1305]&~m[1306]&m[1360])|(m[1303]&m[1304]&~m[1305]&m[1306]&m[1360])|(m[1303]&~m[1304]&m[1305]&m[1306]&m[1360])|(~m[1303]&m[1304]&m[1305]&m[1306]&m[1360]))&~BiasedRNG[814])|((m[1303]&m[1304]&~m[1305]&~m[1306]&~m[1360])|(m[1303]&~m[1304]&m[1305]&~m[1306]&~m[1360])|(~m[1303]&m[1304]&m[1305]&~m[1306]&~m[1360])|(m[1303]&m[1304]&m[1305]&~m[1306]&~m[1360])|(m[1303]&m[1304]&m[1305]&m[1306]&~m[1360])|(m[1303]&m[1304]&~m[1305]&~m[1306]&m[1360])|(m[1303]&~m[1304]&m[1305]&~m[1306]&m[1360])|(~m[1303]&m[1304]&m[1305]&~m[1306]&m[1360])|(m[1303]&m[1304]&m[1305]&~m[1306]&m[1360])|(m[1303]&m[1304]&m[1305]&m[1306]&m[1360]));
    m[1312] = (((m[1308]&~m[1309]&~m[1310]&~m[1311]&~m[1363])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1363])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1363])|(m[1308]&m[1309]&~m[1310]&m[1311]&~m[1363])|(m[1308]&~m[1309]&m[1310]&m[1311]&~m[1363])|(~m[1308]&m[1309]&m[1310]&m[1311]&~m[1363]))&BiasedRNG[815])|(((m[1308]&~m[1309]&~m[1310]&~m[1311]&m[1363])|(~m[1308]&m[1309]&~m[1310]&~m[1311]&m[1363])|(~m[1308]&~m[1309]&m[1310]&~m[1311]&m[1363])|(m[1308]&m[1309]&~m[1310]&m[1311]&m[1363])|(m[1308]&~m[1309]&m[1310]&m[1311]&m[1363])|(~m[1308]&m[1309]&m[1310]&m[1311]&m[1363]))&~BiasedRNG[815])|((m[1308]&m[1309]&~m[1310]&~m[1311]&~m[1363])|(m[1308]&~m[1309]&m[1310]&~m[1311]&~m[1363])|(~m[1308]&m[1309]&m[1310]&~m[1311]&~m[1363])|(m[1308]&m[1309]&m[1310]&~m[1311]&~m[1363])|(m[1308]&m[1309]&m[1310]&m[1311]&~m[1363])|(m[1308]&m[1309]&~m[1310]&~m[1311]&m[1363])|(m[1308]&~m[1309]&m[1310]&~m[1311]&m[1363])|(~m[1308]&m[1309]&m[1310]&~m[1311]&m[1363])|(m[1308]&m[1309]&m[1310]&~m[1311]&m[1363])|(m[1308]&m[1309]&m[1310]&m[1311]&m[1363]));
    m[1317] = (((m[1313]&~m[1314]&~m[1315]&~m[1316]&~m[1365])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1365])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1365])|(m[1313]&m[1314]&~m[1315]&m[1316]&~m[1365])|(m[1313]&~m[1314]&m[1315]&m[1316]&~m[1365])|(~m[1313]&m[1314]&m[1315]&m[1316]&~m[1365]))&BiasedRNG[816])|(((m[1313]&~m[1314]&~m[1315]&~m[1316]&m[1365])|(~m[1313]&m[1314]&~m[1315]&~m[1316]&m[1365])|(~m[1313]&~m[1314]&m[1315]&~m[1316]&m[1365])|(m[1313]&m[1314]&~m[1315]&m[1316]&m[1365])|(m[1313]&~m[1314]&m[1315]&m[1316]&m[1365])|(~m[1313]&m[1314]&m[1315]&m[1316]&m[1365]))&~BiasedRNG[816])|((m[1313]&m[1314]&~m[1315]&~m[1316]&~m[1365])|(m[1313]&~m[1314]&m[1315]&~m[1316]&~m[1365])|(~m[1313]&m[1314]&m[1315]&~m[1316]&~m[1365])|(m[1313]&m[1314]&m[1315]&~m[1316]&~m[1365])|(m[1313]&m[1314]&m[1315]&m[1316]&~m[1365])|(m[1313]&m[1314]&~m[1315]&~m[1316]&m[1365])|(m[1313]&~m[1314]&m[1315]&~m[1316]&m[1365])|(~m[1313]&m[1314]&m[1315]&~m[1316]&m[1365])|(m[1313]&m[1314]&m[1315]&~m[1316]&m[1365])|(m[1313]&m[1314]&m[1315]&m[1316]&m[1365]));
    m[1322] = (((m[1318]&~m[1319]&~m[1320]&~m[1321]&~m[1370])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1370])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1370])|(m[1318]&m[1319]&~m[1320]&m[1321]&~m[1370])|(m[1318]&~m[1319]&m[1320]&m[1321]&~m[1370])|(~m[1318]&m[1319]&m[1320]&m[1321]&~m[1370]))&BiasedRNG[817])|(((m[1318]&~m[1319]&~m[1320]&~m[1321]&m[1370])|(~m[1318]&m[1319]&~m[1320]&~m[1321]&m[1370])|(~m[1318]&~m[1319]&m[1320]&~m[1321]&m[1370])|(m[1318]&m[1319]&~m[1320]&m[1321]&m[1370])|(m[1318]&~m[1319]&m[1320]&m[1321]&m[1370])|(~m[1318]&m[1319]&m[1320]&m[1321]&m[1370]))&~BiasedRNG[817])|((m[1318]&m[1319]&~m[1320]&~m[1321]&~m[1370])|(m[1318]&~m[1319]&m[1320]&~m[1321]&~m[1370])|(~m[1318]&m[1319]&m[1320]&~m[1321]&~m[1370])|(m[1318]&m[1319]&m[1320]&~m[1321]&~m[1370])|(m[1318]&m[1319]&m[1320]&m[1321]&~m[1370])|(m[1318]&m[1319]&~m[1320]&~m[1321]&m[1370])|(m[1318]&~m[1319]&m[1320]&~m[1321]&m[1370])|(~m[1318]&m[1319]&m[1320]&~m[1321]&m[1370])|(m[1318]&m[1319]&m[1320]&~m[1321]&m[1370])|(m[1318]&m[1319]&m[1320]&m[1321]&m[1370]));
    m[1327] = (((m[1323]&~m[1324]&~m[1325]&~m[1326]&~m[1375])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1375])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1375])|(m[1323]&m[1324]&~m[1325]&m[1326]&~m[1375])|(m[1323]&~m[1324]&m[1325]&m[1326]&~m[1375])|(~m[1323]&m[1324]&m[1325]&m[1326]&~m[1375]))&BiasedRNG[818])|(((m[1323]&~m[1324]&~m[1325]&~m[1326]&m[1375])|(~m[1323]&m[1324]&~m[1325]&~m[1326]&m[1375])|(~m[1323]&~m[1324]&m[1325]&~m[1326]&m[1375])|(m[1323]&m[1324]&~m[1325]&m[1326]&m[1375])|(m[1323]&~m[1324]&m[1325]&m[1326]&m[1375])|(~m[1323]&m[1324]&m[1325]&m[1326]&m[1375]))&~BiasedRNG[818])|((m[1323]&m[1324]&~m[1325]&~m[1326]&~m[1375])|(m[1323]&~m[1324]&m[1325]&~m[1326]&~m[1375])|(~m[1323]&m[1324]&m[1325]&~m[1326]&~m[1375])|(m[1323]&m[1324]&m[1325]&~m[1326]&~m[1375])|(m[1323]&m[1324]&m[1325]&m[1326]&~m[1375])|(m[1323]&m[1324]&~m[1325]&~m[1326]&m[1375])|(m[1323]&~m[1324]&m[1325]&~m[1326]&m[1375])|(~m[1323]&m[1324]&m[1325]&~m[1326]&m[1375])|(m[1323]&m[1324]&m[1325]&~m[1326]&m[1375])|(m[1323]&m[1324]&m[1325]&m[1326]&m[1375]));
    m[1332] = (((m[1328]&~m[1329]&~m[1330]&~m[1331]&~m[1380])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1380])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1380])|(m[1328]&m[1329]&~m[1330]&m[1331]&~m[1380])|(m[1328]&~m[1329]&m[1330]&m[1331]&~m[1380])|(~m[1328]&m[1329]&m[1330]&m[1331]&~m[1380]))&BiasedRNG[819])|(((m[1328]&~m[1329]&~m[1330]&~m[1331]&m[1380])|(~m[1328]&m[1329]&~m[1330]&~m[1331]&m[1380])|(~m[1328]&~m[1329]&m[1330]&~m[1331]&m[1380])|(m[1328]&m[1329]&~m[1330]&m[1331]&m[1380])|(m[1328]&~m[1329]&m[1330]&m[1331]&m[1380])|(~m[1328]&m[1329]&m[1330]&m[1331]&m[1380]))&~BiasedRNG[819])|((m[1328]&m[1329]&~m[1330]&~m[1331]&~m[1380])|(m[1328]&~m[1329]&m[1330]&~m[1331]&~m[1380])|(~m[1328]&m[1329]&m[1330]&~m[1331]&~m[1380])|(m[1328]&m[1329]&m[1330]&~m[1331]&~m[1380])|(m[1328]&m[1329]&m[1330]&m[1331]&~m[1380])|(m[1328]&m[1329]&~m[1330]&~m[1331]&m[1380])|(m[1328]&~m[1329]&m[1330]&~m[1331]&m[1380])|(~m[1328]&m[1329]&m[1330]&~m[1331]&m[1380])|(m[1328]&m[1329]&m[1330]&~m[1331]&m[1380])|(m[1328]&m[1329]&m[1330]&m[1331]&m[1380]));
    m[1337] = (((m[1333]&~m[1334]&~m[1335]&~m[1336]&~m[1385])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1385])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1385])|(m[1333]&m[1334]&~m[1335]&m[1336]&~m[1385])|(m[1333]&~m[1334]&m[1335]&m[1336]&~m[1385])|(~m[1333]&m[1334]&m[1335]&m[1336]&~m[1385]))&BiasedRNG[820])|(((m[1333]&~m[1334]&~m[1335]&~m[1336]&m[1385])|(~m[1333]&m[1334]&~m[1335]&~m[1336]&m[1385])|(~m[1333]&~m[1334]&m[1335]&~m[1336]&m[1385])|(m[1333]&m[1334]&~m[1335]&m[1336]&m[1385])|(m[1333]&~m[1334]&m[1335]&m[1336]&m[1385])|(~m[1333]&m[1334]&m[1335]&m[1336]&m[1385]))&~BiasedRNG[820])|((m[1333]&m[1334]&~m[1335]&~m[1336]&~m[1385])|(m[1333]&~m[1334]&m[1335]&~m[1336]&~m[1385])|(~m[1333]&m[1334]&m[1335]&~m[1336]&~m[1385])|(m[1333]&m[1334]&m[1335]&~m[1336]&~m[1385])|(m[1333]&m[1334]&m[1335]&m[1336]&~m[1385])|(m[1333]&m[1334]&~m[1335]&~m[1336]&m[1385])|(m[1333]&~m[1334]&m[1335]&~m[1336]&m[1385])|(~m[1333]&m[1334]&m[1335]&~m[1336]&m[1385])|(m[1333]&m[1334]&m[1335]&~m[1336]&m[1385])|(m[1333]&m[1334]&m[1335]&m[1336]&m[1385]));
    m[1342] = (((m[1338]&~m[1339]&~m[1340]&~m[1341]&~m[1390])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1390])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1390])|(m[1338]&m[1339]&~m[1340]&m[1341]&~m[1390])|(m[1338]&~m[1339]&m[1340]&m[1341]&~m[1390])|(~m[1338]&m[1339]&m[1340]&m[1341]&~m[1390]))&BiasedRNG[821])|(((m[1338]&~m[1339]&~m[1340]&~m[1341]&m[1390])|(~m[1338]&m[1339]&~m[1340]&~m[1341]&m[1390])|(~m[1338]&~m[1339]&m[1340]&~m[1341]&m[1390])|(m[1338]&m[1339]&~m[1340]&m[1341]&m[1390])|(m[1338]&~m[1339]&m[1340]&m[1341]&m[1390])|(~m[1338]&m[1339]&m[1340]&m[1341]&m[1390]))&~BiasedRNG[821])|((m[1338]&m[1339]&~m[1340]&~m[1341]&~m[1390])|(m[1338]&~m[1339]&m[1340]&~m[1341]&~m[1390])|(~m[1338]&m[1339]&m[1340]&~m[1341]&~m[1390])|(m[1338]&m[1339]&m[1340]&~m[1341]&~m[1390])|(m[1338]&m[1339]&m[1340]&m[1341]&~m[1390])|(m[1338]&m[1339]&~m[1340]&~m[1341]&m[1390])|(m[1338]&~m[1339]&m[1340]&~m[1341]&m[1390])|(~m[1338]&m[1339]&m[1340]&~m[1341]&m[1390])|(m[1338]&m[1339]&m[1340]&~m[1341]&m[1390])|(m[1338]&m[1339]&m[1340]&m[1341]&m[1390]));
    m[1347] = (((m[1343]&~m[1344]&~m[1345]&~m[1346]&~m[1395])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1395])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1395])|(m[1343]&m[1344]&~m[1345]&m[1346]&~m[1395])|(m[1343]&~m[1344]&m[1345]&m[1346]&~m[1395])|(~m[1343]&m[1344]&m[1345]&m[1346]&~m[1395]))&BiasedRNG[822])|(((m[1343]&~m[1344]&~m[1345]&~m[1346]&m[1395])|(~m[1343]&m[1344]&~m[1345]&~m[1346]&m[1395])|(~m[1343]&~m[1344]&m[1345]&~m[1346]&m[1395])|(m[1343]&m[1344]&~m[1345]&m[1346]&m[1395])|(m[1343]&~m[1344]&m[1345]&m[1346]&m[1395])|(~m[1343]&m[1344]&m[1345]&m[1346]&m[1395]))&~BiasedRNG[822])|((m[1343]&m[1344]&~m[1345]&~m[1346]&~m[1395])|(m[1343]&~m[1344]&m[1345]&~m[1346]&~m[1395])|(~m[1343]&m[1344]&m[1345]&~m[1346]&~m[1395])|(m[1343]&m[1344]&m[1345]&~m[1346]&~m[1395])|(m[1343]&m[1344]&m[1345]&m[1346]&~m[1395])|(m[1343]&m[1344]&~m[1345]&~m[1346]&m[1395])|(m[1343]&~m[1344]&m[1345]&~m[1346]&m[1395])|(~m[1343]&m[1344]&m[1345]&~m[1346]&m[1395])|(m[1343]&m[1344]&m[1345]&~m[1346]&m[1395])|(m[1343]&m[1344]&m[1345]&m[1346]&m[1395]));
    m[1352] = (((m[1348]&~m[1349]&~m[1350]&~m[1351]&~m[1400])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1400])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1400])|(m[1348]&m[1349]&~m[1350]&m[1351]&~m[1400])|(m[1348]&~m[1349]&m[1350]&m[1351]&~m[1400])|(~m[1348]&m[1349]&m[1350]&m[1351]&~m[1400]))&BiasedRNG[823])|(((m[1348]&~m[1349]&~m[1350]&~m[1351]&m[1400])|(~m[1348]&m[1349]&~m[1350]&~m[1351]&m[1400])|(~m[1348]&~m[1349]&m[1350]&~m[1351]&m[1400])|(m[1348]&m[1349]&~m[1350]&m[1351]&m[1400])|(m[1348]&~m[1349]&m[1350]&m[1351]&m[1400])|(~m[1348]&m[1349]&m[1350]&m[1351]&m[1400]))&~BiasedRNG[823])|((m[1348]&m[1349]&~m[1350]&~m[1351]&~m[1400])|(m[1348]&~m[1349]&m[1350]&~m[1351]&~m[1400])|(~m[1348]&m[1349]&m[1350]&~m[1351]&~m[1400])|(m[1348]&m[1349]&m[1350]&~m[1351]&~m[1400])|(m[1348]&m[1349]&m[1350]&m[1351]&~m[1400])|(m[1348]&m[1349]&~m[1350]&~m[1351]&m[1400])|(m[1348]&~m[1349]&m[1350]&~m[1351]&m[1400])|(~m[1348]&m[1349]&m[1350]&~m[1351]&m[1400])|(m[1348]&m[1349]&m[1350]&~m[1351]&m[1400])|(m[1348]&m[1349]&m[1350]&m[1351]&m[1400]));
    m[1357] = (((m[1353]&~m[1354]&~m[1355]&~m[1356]&~m[1405])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1405])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1405])|(m[1353]&m[1354]&~m[1355]&m[1356]&~m[1405])|(m[1353]&~m[1354]&m[1355]&m[1356]&~m[1405])|(~m[1353]&m[1354]&m[1355]&m[1356]&~m[1405]))&BiasedRNG[824])|(((m[1353]&~m[1354]&~m[1355]&~m[1356]&m[1405])|(~m[1353]&m[1354]&~m[1355]&~m[1356]&m[1405])|(~m[1353]&~m[1354]&m[1355]&~m[1356]&m[1405])|(m[1353]&m[1354]&~m[1355]&m[1356]&m[1405])|(m[1353]&~m[1354]&m[1355]&m[1356]&m[1405])|(~m[1353]&m[1354]&m[1355]&m[1356]&m[1405]))&~BiasedRNG[824])|((m[1353]&m[1354]&~m[1355]&~m[1356]&~m[1405])|(m[1353]&~m[1354]&m[1355]&~m[1356]&~m[1405])|(~m[1353]&m[1354]&m[1355]&~m[1356]&~m[1405])|(m[1353]&m[1354]&m[1355]&~m[1356]&~m[1405])|(m[1353]&m[1354]&m[1355]&m[1356]&~m[1405])|(m[1353]&m[1354]&~m[1355]&~m[1356]&m[1405])|(m[1353]&~m[1354]&m[1355]&~m[1356]&m[1405])|(~m[1353]&m[1354]&m[1355]&~m[1356]&m[1405])|(m[1353]&m[1354]&m[1355]&~m[1356]&m[1405])|(m[1353]&m[1354]&m[1355]&m[1356]&m[1405]));
    m[1362] = (((m[1358]&~m[1359]&~m[1360]&~m[1361]&~m[1410])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1410])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1410])|(m[1358]&m[1359]&~m[1360]&m[1361]&~m[1410])|(m[1358]&~m[1359]&m[1360]&m[1361]&~m[1410])|(~m[1358]&m[1359]&m[1360]&m[1361]&~m[1410]))&BiasedRNG[825])|(((m[1358]&~m[1359]&~m[1360]&~m[1361]&m[1410])|(~m[1358]&m[1359]&~m[1360]&~m[1361]&m[1410])|(~m[1358]&~m[1359]&m[1360]&~m[1361]&m[1410])|(m[1358]&m[1359]&~m[1360]&m[1361]&m[1410])|(m[1358]&~m[1359]&m[1360]&m[1361]&m[1410])|(~m[1358]&m[1359]&m[1360]&m[1361]&m[1410]))&~BiasedRNG[825])|((m[1358]&m[1359]&~m[1360]&~m[1361]&~m[1410])|(m[1358]&~m[1359]&m[1360]&~m[1361]&~m[1410])|(~m[1358]&m[1359]&m[1360]&~m[1361]&~m[1410])|(m[1358]&m[1359]&m[1360]&~m[1361]&~m[1410])|(m[1358]&m[1359]&m[1360]&m[1361]&~m[1410])|(m[1358]&m[1359]&~m[1360]&~m[1361]&m[1410])|(m[1358]&~m[1359]&m[1360]&~m[1361]&m[1410])|(~m[1358]&m[1359]&m[1360]&~m[1361]&m[1410])|(m[1358]&m[1359]&m[1360]&~m[1361]&m[1410])|(m[1358]&m[1359]&m[1360]&m[1361]&m[1410]));
    m[1367] = (((m[1363]&~m[1364]&~m[1365]&~m[1366]&~m[1413])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1413])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1413])|(m[1363]&m[1364]&~m[1365]&m[1366]&~m[1413])|(m[1363]&~m[1364]&m[1365]&m[1366]&~m[1413])|(~m[1363]&m[1364]&m[1365]&m[1366]&~m[1413]))&BiasedRNG[826])|(((m[1363]&~m[1364]&~m[1365]&~m[1366]&m[1413])|(~m[1363]&m[1364]&~m[1365]&~m[1366]&m[1413])|(~m[1363]&~m[1364]&m[1365]&~m[1366]&m[1413])|(m[1363]&m[1364]&~m[1365]&m[1366]&m[1413])|(m[1363]&~m[1364]&m[1365]&m[1366]&m[1413])|(~m[1363]&m[1364]&m[1365]&m[1366]&m[1413]))&~BiasedRNG[826])|((m[1363]&m[1364]&~m[1365]&~m[1366]&~m[1413])|(m[1363]&~m[1364]&m[1365]&~m[1366]&~m[1413])|(~m[1363]&m[1364]&m[1365]&~m[1366]&~m[1413])|(m[1363]&m[1364]&m[1365]&~m[1366]&~m[1413])|(m[1363]&m[1364]&m[1365]&m[1366]&~m[1413])|(m[1363]&m[1364]&~m[1365]&~m[1366]&m[1413])|(m[1363]&~m[1364]&m[1365]&~m[1366]&m[1413])|(~m[1363]&m[1364]&m[1365]&~m[1366]&m[1413])|(m[1363]&m[1364]&m[1365]&~m[1366]&m[1413])|(m[1363]&m[1364]&m[1365]&m[1366]&m[1413]));
    m[1372] = (((m[1368]&~m[1369]&~m[1370]&~m[1371]&~m[1415])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1415])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1415])|(m[1368]&m[1369]&~m[1370]&m[1371]&~m[1415])|(m[1368]&~m[1369]&m[1370]&m[1371]&~m[1415])|(~m[1368]&m[1369]&m[1370]&m[1371]&~m[1415]))&BiasedRNG[827])|(((m[1368]&~m[1369]&~m[1370]&~m[1371]&m[1415])|(~m[1368]&m[1369]&~m[1370]&~m[1371]&m[1415])|(~m[1368]&~m[1369]&m[1370]&~m[1371]&m[1415])|(m[1368]&m[1369]&~m[1370]&m[1371]&m[1415])|(m[1368]&~m[1369]&m[1370]&m[1371]&m[1415])|(~m[1368]&m[1369]&m[1370]&m[1371]&m[1415]))&~BiasedRNG[827])|((m[1368]&m[1369]&~m[1370]&~m[1371]&~m[1415])|(m[1368]&~m[1369]&m[1370]&~m[1371]&~m[1415])|(~m[1368]&m[1369]&m[1370]&~m[1371]&~m[1415])|(m[1368]&m[1369]&m[1370]&~m[1371]&~m[1415])|(m[1368]&m[1369]&m[1370]&m[1371]&~m[1415])|(m[1368]&m[1369]&~m[1370]&~m[1371]&m[1415])|(m[1368]&~m[1369]&m[1370]&~m[1371]&m[1415])|(~m[1368]&m[1369]&m[1370]&~m[1371]&m[1415])|(m[1368]&m[1369]&m[1370]&~m[1371]&m[1415])|(m[1368]&m[1369]&m[1370]&m[1371]&m[1415]));
    m[1377] = (((m[1373]&~m[1374]&~m[1375]&~m[1376]&~m[1420])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1420])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1420])|(m[1373]&m[1374]&~m[1375]&m[1376]&~m[1420])|(m[1373]&~m[1374]&m[1375]&m[1376]&~m[1420])|(~m[1373]&m[1374]&m[1375]&m[1376]&~m[1420]))&BiasedRNG[828])|(((m[1373]&~m[1374]&~m[1375]&~m[1376]&m[1420])|(~m[1373]&m[1374]&~m[1375]&~m[1376]&m[1420])|(~m[1373]&~m[1374]&m[1375]&~m[1376]&m[1420])|(m[1373]&m[1374]&~m[1375]&m[1376]&m[1420])|(m[1373]&~m[1374]&m[1375]&m[1376]&m[1420])|(~m[1373]&m[1374]&m[1375]&m[1376]&m[1420]))&~BiasedRNG[828])|((m[1373]&m[1374]&~m[1375]&~m[1376]&~m[1420])|(m[1373]&~m[1374]&m[1375]&~m[1376]&~m[1420])|(~m[1373]&m[1374]&m[1375]&~m[1376]&~m[1420])|(m[1373]&m[1374]&m[1375]&~m[1376]&~m[1420])|(m[1373]&m[1374]&m[1375]&m[1376]&~m[1420])|(m[1373]&m[1374]&~m[1375]&~m[1376]&m[1420])|(m[1373]&~m[1374]&m[1375]&~m[1376]&m[1420])|(~m[1373]&m[1374]&m[1375]&~m[1376]&m[1420])|(m[1373]&m[1374]&m[1375]&~m[1376]&m[1420])|(m[1373]&m[1374]&m[1375]&m[1376]&m[1420]));
    m[1382] = (((m[1378]&~m[1379]&~m[1380]&~m[1381]&~m[1425])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1425])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1425])|(m[1378]&m[1379]&~m[1380]&m[1381]&~m[1425])|(m[1378]&~m[1379]&m[1380]&m[1381]&~m[1425])|(~m[1378]&m[1379]&m[1380]&m[1381]&~m[1425]))&BiasedRNG[829])|(((m[1378]&~m[1379]&~m[1380]&~m[1381]&m[1425])|(~m[1378]&m[1379]&~m[1380]&~m[1381]&m[1425])|(~m[1378]&~m[1379]&m[1380]&~m[1381]&m[1425])|(m[1378]&m[1379]&~m[1380]&m[1381]&m[1425])|(m[1378]&~m[1379]&m[1380]&m[1381]&m[1425])|(~m[1378]&m[1379]&m[1380]&m[1381]&m[1425]))&~BiasedRNG[829])|((m[1378]&m[1379]&~m[1380]&~m[1381]&~m[1425])|(m[1378]&~m[1379]&m[1380]&~m[1381]&~m[1425])|(~m[1378]&m[1379]&m[1380]&~m[1381]&~m[1425])|(m[1378]&m[1379]&m[1380]&~m[1381]&~m[1425])|(m[1378]&m[1379]&m[1380]&m[1381]&~m[1425])|(m[1378]&m[1379]&~m[1380]&~m[1381]&m[1425])|(m[1378]&~m[1379]&m[1380]&~m[1381]&m[1425])|(~m[1378]&m[1379]&m[1380]&~m[1381]&m[1425])|(m[1378]&m[1379]&m[1380]&~m[1381]&m[1425])|(m[1378]&m[1379]&m[1380]&m[1381]&m[1425]));
    m[1387] = (((m[1383]&~m[1384]&~m[1385]&~m[1386]&~m[1430])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1430])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1430])|(m[1383]&m[1384]&~m[1385]&m[1386]&~m[1430])|(m[1383]&~m[1384]&m[1385]&m[1386]&~m[1430])|(~m[1383]&m[1384]&m[1385]&m[1386]&~m[1430]))&BiasedRNG[830])|(((m[1383]&~m[1384]&~m[1385]&~m[1386]&m[1430])|(~m[1383]&m[1384]&~m[1385]&~m[1386]&m[1430])|(~m[1383]&~m[1384]&m[1385]&~m[1386]&m[1430])|(m[1383]&m[1384]&~m[1385]&m[1386]&m[1430])|(m[1383]&~m[1384]&m[1385]&m[1386]&m[1430])|(~m[1383]&m[1384]&m[1385]&m[1386]&m[1430]))&~BiasedRNG[830])|((m[1383]&m[1384]&~m[1385]&~m[1386]&~m[1430])|(m[1383]&~m[1384]&m[1385]&~m[1386]&~m[1430])|(~m[1383]&m[1384]&m[1385]&~m[1386]&~m[1430])|(m[1383]&m[1384]&m[1385]&~m[1386]&~m[1430])|(m[1383]&m[1384]&m[1385]&m[1386]&~m[1430])|(m[1383]&m[1384]&~m[1385]&~m[1386]&m[1430])|(m[1383]&~m[1384]&m[1385]&~m[1386]&m[1430])|(~m[1383]&m[1384]&m[1385]&~m[1386]&m[1430])|(m[1383]&m[1384]&m[1385]&~m[1386]&m[1430])|(m[1383]&m[1384]&m[1385]&m[1386]&m[1430]));
    m[1392] = (((m[1388]&~m[1389]&~m[1390]&~m[1391]&~m[1435])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1435])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1435])|(m[1388]&m[1389]&~m[1390]&m[1391]&~m[1435])|(m[1388]&~m[1389]&m[1390]&m[1391]&~m[1435])|(~m[1388]&m[1389]&m[1390]&m[1391]&~m[1435]))&BiasedRNG[831])|(((m[1388]&~m[1389]&~m[1390]&~m[1391]&m[1435])|(~m[1388]&m[1389]&~m[1390]&~m[1391]&m[1435])|(~m[1388]&~m[1389]&m[1390]&~m[1391]&m[1435])|(m[1388]&m[1389]&~m[1390]&m[1391]&m[1435])|(m[1388]&~m[1389]&m[1390]&m[1391]&m[1435])|(~m[1388]&m[1389]&m[1390]&m[1391]&m[1435]))&~BiasedRNG[831])|((m[1388]&m[1389]&~m[1390]&~m[1391]&~m[1435])|(m[1388]&~m[1389]&m[1390]&~m[1391]&~m[1435])|(~m[1388]&m[1389]&m[1390]&~m[1391]&~m[1435])|(m[1388]&m[1389]&m[1390]&~m[1391]&~m[1435])|(m[1388]&m[1389]&m[1390]&m[1391]&~m[1435])|(m[1388]&m[1389]&~m[1390]&~m[1391]&m[1435])|(m[1388]&~m[1389]&m[1390]&~m[1391]&m[1435])|(~m[1388]&m[1389]&m[1390]&~m[1391]&m[1435])|(m[1388]&m[1389]&m[1390]&~m[1391]&m[1435])|(m[1388]&m[1389]&m[1390]&m[1391]&m[1435]));
    m[1397] = (((m[1393]&~m[1394]&~m[1395]&~m[1396]&~m[1440])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1440])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1440])|(m[1393]&m[1394]&~m[1395]&m[1396]&~m[1440])|(m[1393]&~m[1394]&m[1395]&m[1396]&~m[1440])|(~m[1393]&m[1394]&m[1395]&m[1396]&~m[1440]))&BiasedRNG[832])|(((m[1393]&~m[1394]&~m[1395]&~m[1396]&m[1440])|(~m[1393]&m[1394]&~m[1395]&~m[1396]&m[1440])|(~m[1393]&~m[1394]&m[1395]&~m[1396]&m[1440])|(m[1393]&m[1394]&~m[1395]&m[1396]&m[1440])|(m[1393]&~m[1394]&m[1395]&m[1396]&m[1440])|(~m[1393]&m[1394]&m[1395]&m[1396]&m[1440]))&~BiasedRNG[832])|((m[1393]&m[1394]&~m[1395]&~m[1396]&~m[1440])|(m[1393]&~m[1394]&m[1395]&~m[1396]&~m[1440])|(~m[1393]&m[1394]&m[1395]&~m[1396]&~m[1440])|(m[1393]&m[1394]&m[1395]&~m[1396]&~m[1440])|(m[1393]&m[1394]&m[1395]&m[1396]&~m[1440])|(m[1393]&m[1394]&~m[1395]&~m[1396]&m[1440])|(m[1393]&~m[1394]&m[1395]&~m[1396]&m[1440])|(~m[1393]&m[1394]&m[1395]&~m[1396]&m[1440])|(m[1393]&m[1394]&m[1395]&~m[1396]&m[1440])|(m[1393]&m[1394]&m[1395]&m[1396]&m[1440]));
    m[1402] = (((m[1398]&~m[1399]&~m[1400]&~m[1401]&~m[1445])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1445])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1445])|(m[1398]&m[1399]&~m[1400]&m[1401]&~m[1445])|(m[1398]&~m[1399]&m[1400]&m[1401]&~m[1445])|(~m[1398]&m[1399]&m[1400]&m[1401]&~m[1445]))&BiasedRNG[833])|(((m[1398]&~m[1399]&~m[1400]&~m[1401]&m[1445])|(~m[1398]&m[1399]&~m[1400]&~m[1401]&m[1445])|(~m[1398]&~m[1399]&m[1400]&~m[1401]&m[1445])|(m[1398]&m[1399]&~m[1400]&m[1401]&m[1445])|(m[1398]&~m[1399]&m[1400]&m[1401]&m[1445])|(~m[1398]&m[1399]&m[1400]&m[1401]&m[1445]))&~BiasedRNG[833])|((m[1398]&m[1399]&~m[1400]&~m[1401]&~m[1445])|(m[1398]&~m[1399]&m[1400]&~m[1401]&~m[1445])|(~m[1398]&m[1399]&m[1400]&~m[1401]&~m[1445])|(m[1398]&m[1399]&m[1400]&~m[1401]&~m[1445])|(m[1398]&m[1399]&m[1400]&m[1401]&~m[1445])|(m[1398]&m[1399]&~m[1400]&~m[1401]&m[1445])|(m[1398]&~m[1399]&m[1400]&~m[1401]&m[1445])|(~m[1398]&m[1399]&m[1400]&~m[1401]&m[1445])|(m[1398]&m[1399]&m[1400]&~m[1401]&m[1445])|(m[1398]&m[1399]&m[1400]&m[1401]&m[1445]));
    m[1407] = (((m[1403]&~m[1404]&~m[1405]&~m[1406]&~m[1450])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1450])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1450])|(m[1403]&m[1404]&~m[1405]&m[1406]&~m[1450])|(m[1403]&~m[1404]&m[1405]&m[1406]&~m[1450])|(~m[1403]&m[1404]&m[1405]&m[1406]&~m[1450]))&BiasedRNG[834])|(((m[1403]&~m[1404]&~m[1405]&~m[1406]&m[1450])|(~m[1403]&m[1404]&~m[1405]&~m[1406]&m[1450])|(~m[1403]&~m[1404]&m[1405]&~m[1406]&m[1450])|(m[1403]&m[1404]&~m[1405]&m[1406]&m[1450])|(m[1403]&~m[1404]&m[1405]&m[1406]&m[1450])|(~m[1403]&m[1404]&m[1405]&m[1406]&m[1450]))&~BiasedRNG[834])|((m[1403]&m[1404]&~m[1405]&~m[1406]&~m[1450])|(m[1403]&~m[1404]&m[1405]&~m[1406]&~m[1450])|(~m[1403]&m[1404]&m[1405]&~m[1406]&~m[1450])|(m[1403]&m[1404]&m[1405]&~m[1406]&~m[1450])|(m[1403]&m[1404]&m[1405]&m[1406]&~m[1450])|(m[1403]&m[1404]&~m[1405]&~m[1406]&m[1450])|(m[1403]&~m[1404]&m[1405]&~m[1406]&m[1450])|(~m[1403]&m[1404]&m[1405]&~m[1406]&m[1450])|(m[1403]&m[1404]&m[1405]&~m[1406]&m[1450])|(m[1403]&m[1404]&m[1405]&m[1406]&m[1450]));
    m[1412] = (((m[1408]&~m[1409]&~m[1410]&~m[1411]&~m[1455])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1455])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1455])|(m[1408]&m[1409]&~m[1410]&m[1411]&~m[1455])|(m[1408]&~m[1409]&m[1410]&m[1411]&~m[1455])|(~m[1408]&m[1409]&m[1410]&m[1411]&~m[1455]))&BiasedRNG[835])|(((m[1408]&~m[1409]&~m[1410]&~m[1411]&m[1455])|(~m[1408]&m[1409]&~m[1410]&~m[1411]&m[1455])|(~m[1408]&~m[1409]&m[1410]&~m[1411]&m[1455])|(m[1408]&m[1409]&~m[1410]&m[1411]&m[1455])|(m[1408]&~m[1409]&m[1410]&m[1411]&m[1455])|(~m[1408]&m[1409]&m[1410]&m[1411]&m[1455]))&~BiasedRNG[835])|((m[1408]&m[1409]&~m[1410]&~m[1411]&~m[1455])|(m[1408]&~m[1409]&m[1410]&~m[1411]&~m[1455])|(~m[1408]&m[1409]&m[1410]&~m[1411]&~m[1455])|(m[1408]&m[1409]&m[1410]&~m[1411]&~m[1455])|(m[1408]&m[1409]&m[1410]&m[1411]&~m[1455])|(m[1408]&m[1409]&~m[1410]&~m[1411]&m[1455])|(m[1408]&~m[1409]&m[1410]&~m[1411]&m[1455])|(~m[1408]&m[1409]&m[1410]&~m[1411]&m[1455])|(m[1408]&m[1409]&m[1410]&~m[1411]&m[1455])|(m[1408]&m[1409]&m[1410]&m[1411]&m[1455]));
    m[1417] = (((m[1413]&~m[1414]&~m[1415]&~m[1416]&~m[1458])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1458])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1458])|(m[1413]&m[1414]&~m[1415]&m[1416]&~m[1458])|(m[1413]&~m[1414]&m[1415]&m[1416]&~m[1458])|(~m[1413]&m[1414]&m[1415]&m[1416]&~m[1458]))&BiasedRNG[836])|(((m[1413]&~m[1414]&~m[1415]&~m[1416]&m[1458])|(~m[1413]&m[1414]&~m[1415]&~m[1416]&m[1458])|(~m[1413]&~m[1414]&m[1415]&~m[1416]&m[1458])|(m[1413]&m[1414]&~m[1415]&m[1416]&m[1458])|(m[1413]&~m[1414]&m[1415]&m[1416]&m[1458])|(~m[1413]&m[1414]&m[1415]&m[1416]&m[1458]))&~BiasedRNG[836])|((m[1413]&m[1414]&~m[1415]&~m[1416]&~m[1458])|(m[1413]&~m[1414]&m[1415]&~m[1416]&~m[1458])|(~m[1413]&m[1414]&m[1415]&~m[1416]&~m[1458])|(m[1413]&m[1414]&m[1415]&~m[1416]&~m[1458])|(m[1413]&m[1414]&m[1415]&m[1416]&~m[1458])|(m[1413]&m[1414]&~m[1415]&~m[1416]&m[1458])|(m[1413]&~m[1414]&m[1415]&~m[1416]&m[1458])|(~m[1413]&m[1414]&m[1415]&~m[1416]&m[1458])|(m[1413]&m[1414]&m[1415]&~m[1416]&m[1458])|(m[1413]&m[1414]&m[1415]&m[1416]&m[1458]));
    m[1422] = (((m[1418]&~m[1419]&~m[1420]&~m[1421]&~m[1460])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1460])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1460])|(m[1418]&m[1419]&~m[1420]&m[1421]&~m[1460])|(m[1418]&~m[1419]&m[1420]&m[1421]&~m[1460])|(~m[1418]&m[1419]&m[1420]&m[1421]&~m[1460]))&BiasedRNG[837])|(((m[1418]&~m[1419]&~m[1420]&~m[1421]&m[1460])|(~m[1418]&m[1419]&~m[1420]&~m[1421]&m[1460])|(~m[1418]&~m[1419]&m[1420]&~m[1421]&m[1460])|(m[1418]&m[1419]&~m[1420]&m[1421]&m[1460])|(m[1418]&~m[1419]&m[1420]&m[1421]&m[1460])|(~m[1418]&m[1419]&m[1420]&m[1421]&m[1460]))&~BiasedRNG[837])|((m[1418]&m[1419]&~m[1420]&~m[1421]&~m[1460])|(m[1418]&~m[1419]&m[1420]&~m[1421]&~m[1460])|(~m[1418]&m[1419]&m[1420]&~m[1421]&~m[1460])|(m[1418]&m[1419]&m[1420]&~m[1421]&~m[1460])|(m[1418]&m[1419]&m[1420]&m[1421]&~m[1460])|(m[1418]&m[1419]&~m[1420]&~m[1421]&m[1460])|(m[1418]&~m[1419]&m[1420]&~m[1421]&m[1460])|(~m[1418]&m[1419]&m[1420]&~m[1421]&m[1460])|(m[1418]&m[1419]&m[1420]&~m[1421]&m[1460])|(m[1418]&m[1419]&m[1420]&m[1421]&m[1460]));
    m[1427] = (((m[1423]&~m[1424]&~m[1425]&~m[1426]&~m[1465])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1465])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1465])|(m[1423]&m[1424]&~m[1425]&m[1426]&~m[1465])|(m[1423]&~m[1424]&m[1425]&m[1426]&~m[1465])|(~m[1423]&m[1424]&m[1425]&m[1426]&~m[1465]))&BiasedRNG[838])|(((m[1423]&~m[1424]&~m[1425]&~m[1426]&m[1465])|(~m[1423]&m[1424]&~m[1425]&~m[1426]&m[1465])|(~m[1423]&~m[1424]&m[1425]&~m[1426]&m[1465])|(m[1423]&m[1424]&~m[1425]&m[1426]&m[1465])|(m[1423]&~m[1424]&m[1425]&m[1426]&m[1465])|(~m[1423]&m[1424]&m[1425]&m[1426]&m[1465]))&~BiasedRNG[838])|((m[1423]&m[1424]&~m[1425]&~m[1426]&~m[1465])|(m[1423]&~m[1424]&m[1425]&~m[1426]&~m[1465])|(~m[1423]&m[1424]&m[1425]&~m[1426]&~m[1465])|(m[1423]&m[1424]&m[1425]&~m[1426]&~m[1465])|(m[1423]&m[1424]&m[1425]&m[1426]&~m[1465])|(m[1423]&m[1424]&~m[1425]&~m[1426]&m[1465])|(m[1423]&~m[1424]&m[1425]&~m[1426]&m[1465])|(~m[1423]&m[1424]&m[1425]&~m[1426]&m[1465])|(m[1423]&m[1424]&m[1425]&~m[1426]&m[1465])|(m[1423]&m[1424]&m[1425]&m[1426]&m[1465]));
    m[1432] = (((m[1428]&~m[1429]&~m[1430]&~m[1431]&~m[1470])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1470])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1470])|(m[1428]&m[1429]&~m[1430]&m[1431]&~m[1470])|(m[1428]&~m[1429]&m[1430]&m[1431]&~m[1470])|(~m[1428]&m[1429]&m[1430]&m[1431]&~m[1470]))&BiasedRNG[839])|(((m[1428]&~m[1429]&~m[1430]&~m[1431]&m[1470])|(~m[1428]&m[1429]&~m[1430]&~m[1431]&m[1470])|(~m[1428]&~m[1429]&m[1430]&~m[1431]&m[1470])|(m[1428]&m[1429]&~m[1430]&m[1431]&m[1470])|(m[1428]&~m[1429]&m[1430]&m[1431]&m[1470])|(~m[1428]&m[1429]&m[1430]&m[1431]&m[1470]))&~BiasedRNG[839])|((m[1428]&m[1429]&~m[1430]&~m[1431]&~m[1470])|(m[1428]&~m[1429]&m[1430]&~m[1431]&~m[1470])|(~m[1428]&m[1429]&m[1430]&~m[1431]&~m[1470])|(m[1428]&m[1429]&m[1430]&~m[1431]&~m[1470])|(m[1428]&m[1429]&m[1430]&m[1431]&~m[1470])|(m[1428]&m[1429]&~m[1430]&~m[1431]&m[1470])|(m[1428]&~m[1429]&m[1430]&~m[1431]&m[1470])|(~m[1428]&m[1429]&m[1430]&~m[1431]&m[1470])|(m[1428]&m[1429]&m[1430]&~m[1431]&m[1470])|(m[1428]&m[1429]&m[1430]&m[1431]&m[1470]));
    m[1437] = (((m[1433]&~m[1434]&~m[1435]&~m[1436]&~m[1475])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1475])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1475])|(m[1433]&m[1434]&~m[1435]&m[1436]&~m[1475])|(m[1433]&~m[1434]&m[1435]&m[1436]&~m[1475])|(~m[1433]&m[1434]&m[1435]&m[1436]&~m[1475]))&BiasedRNG[840])|(((m[1433]&~m[1434]&~m[1435]&~m[1436]&m[1475])|(~m[1433]&m[1434]&~m[1435]&~m[1436]&m[1475])|(~m[1433]&~m[1434]&m[1435]&~m[1436]&m[1475])|(m[1433]&m[1434]&~m[1435]&m[1436]&m[1475])|(m[1433]&~m[1434]&m[1435]&m[1436]&m[1475])|(~m[1433]&m[1434]&m[1435]&m[1436]&m[1475]))&~BiasedRNG[840])|((m[1433]&m[1434]&~m[1435]&~m[1436]&~m[1475])|(m[1433]&~m[1434]&m[1435]&~m[1436]&~m[1475])|(~m[1433]&m[1434]&m[1435]&~m[1436]&~m[1475])|(m[1433]&m[1434]&m[1435]&~m[1436]&~m[1475])|(m[1433]&m[1434]&m[1435]&m[1436]&~m[1475])|(m[1433]&m[1434]&~m[1435]&~m[1436]&m[1475])|(m[1433]&~m[1434]&m[1435]&~m[1436]&m[1475])|(~m[1433]&m[1434]&m[1435]&~m[1436]&m[1475])|(m[1433]&m[1434]&m[1435]&~m[1436]&m[1475])|(m[1433]&m[1434]&m[1435]&m[1436]&m[1475]));
    m[1442] = (((m[1438]&~m[1439]&~m[1440]&~m[1441]&~m[1480])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1480])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1480])|(m[1438]&m[1439]&~m[1440]&m[1441]&~m[1480])|(m[1438]&~m[1439]&m[1440]&m[1441]&~m[1480])|(~m[1438]&m[1439]&m[1440]&m[1441]&~m[1480]))&BiasedRNG[841])|(((m[1438]&~m[1439]&~m[1440]&~m[1441]&m[1480])|(~m[1438]&m[1439]&~m[1440]&~m[1441]&m[1480])|(~m[1438]&~m[1439]&m[1440]&~m[1441]&m[1480])|(m[1438]&m[1439]&~m[1440]&m[1441]&m[1480])|(m[1438]&~m[1439]&m[1440]&m[1441]&m[1480])|(~m[1438]&m[1439]&m[1440]&m[1441]&m[1480]))&~BiasedRNG[841])|((m[1438]&m[1439]&~m[1440]&~m[1441]&~m[1480])|(m[1438]&~m[1439]&m[1440]&~m[1441]&~m[1480])|(~m[1438]&m[1439]&m[1440]&~m[1441]&~m[1480])|(m[1438]&m[1439]&m[1440]&~m[1441]&~m[1480])|(m[1438]&m[1439]&m[1440]&m[1441]&~m[1480])|(m[1438]&m[1439]&~m[1440]&~m[1441]&m[1480])|(m[1438]&~m[1439]&m[1440]&~m[1441]&m[1480])|(~m[1438]&m[1439]&m[1440]&~m[1441]&m[1480])|(m[1438]&m[1439]&m[1440]&~m[1441]&m[1480])|(m[1438]&m[1439]&m[1440]&m[1441]&m[1480]));
    m[1447] = (((m[1443]&~m[1444]&~m[1445]&~m[1446]&~m[1485])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1485])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1485])|(m[1443]&m[1444]&~m[1445]&m[1446]&~m[1485])|(m[1443]&~m[1444]&m[1445]&m[1446]&~m[1485])|(~m[1443]&m[1444]&m[1445]&m[1446]&~m[1485]))&BiasedRNG[842])|(((m[1443]&~m[1444]&~m[1445]&~m[1446]&m[1485])|(~m[1443]&m[1444]&~m[1445]&~m[1446]&m[1485])|(~m[1443]&~m[1444]&m[1445]&~m[1446]&m[1485])|(m[1443]&m[1444]&~m[1445]&m[1446]&m[1485])|(m[1443]&~m[1444]&m[1445]&m[1446]&m[1485])|(~m[1443]&m[1444]&m[1445]&m[1446]&m[1485]))&~BiasedRNG[842])|((m[1443]&m[1444]&~m[1445]&~m[1446]&~m[1485])|(m[1443]&~m[1444]&m[1445]&~m[1446]&~m[1485])|(~m[1443]&m[1444]&m[1445]&~m[1446]&~m[1485])|(m[1443]&m[1444]&m[1445]&~m[1446]&~m[1485])|(m[1443]&m[1444]&m[1445]&m[1446]&~m[1485])|(m[1443]&m[1444]&~m[1445]&~m[1446]&m[1485])|(m[1443]&~m[1444]&m[1445]&~m[1446]&m[1485])|(~m[1443]&m[1444]&m[1445]&~m[1446]&m[1485])|(m[1443]&m[1444]&m[1445]&~m[1446]&m[1485])|(m[1443]&m[1444]&m[1445]&m[1446]&m[1485]));
    m[1452] = (((m[1448]&~m[1449]&~m[1450]&~m[1451]&~m[1490])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1490])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1490])|(m[1448]&m[1449]&~m[1450]&m[1451]&~m[1490])|(m[1448]&~m[1449]&m[1450]&m[1451]&~m[1490])|(~m[1448]&m[1449]&m[1450]&m[1451]&~m[1490]))&BiasedRNG[843])|(((m[1448]&~m[1449]&~m[1450]&~m[1451]&m[1490])|(~m[1448]&m[1449]&~m[1450]&~m[1451]&m[1490])|(~m[1448]&~m[1449]&m[1450]&~m[1451]&m[1490])|(m[1448]&m[1449]&~m[1450]&m[1451]&m[1490])|(m[1448]&~m[1449]&m[1450]&m[1451]&m[1490])|(~m[1448]&m[1449]&m[1450]&m[1451]&m[1490]))&~BiasedRNG[843])|((m[1448]&m[1449]&~m[1450]&~m[1451]&~m[1490])|(m[1448]&~m[1449]&m[1450]&~m[1451]&~m[1490])|(~m[1448]&m[1449]&m[1450]&~m[1451]&~m[1490])|(m[1448]&m[1449]&m[1450]&~m[1451]&~m[1490])|(m[1448]&m[1449]&m[1450]&m[1451]&~m[1490])|(m[1448]&m[1449]&~m[1450]&~m[1451]&m[1490])|(m[1448]&~m[1449]&m[1450]&~m[1451]&m[1490])|(~m[1448]&m[1449]&m[1450]&~m[1451]&m[1490])|(m[1448]&m[1449]&m[1450]&~m[1451]&m[1490])|(m[1448]&m[1449]&m[1450]&m[1451]&m[1490]));
    m[1457] = (((m[1453]&~m[1454]&~m[1455]&~m[1456]&~m[1495])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1495])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1495])|(m[1453]&m[1454]&~m[1455]&m[1456]&~m[1495])|(m[1453]&~m[1454]&m[1455]&m[1456]&~m[1495])|(~m[1453]&m[1454]&m[1455]&m[1456]&~m[1495]))&BiasedRNG[844])|(((m[1453]&~m[1454]&~m[1455]&~m[1456]&m[1495])|(~m[1453]&m[1454]&~m[1455]&~m[1456]&m[1495])|(~m[1453]&~m[1454]&m[1455]&~m[1456]&m[1495])|(m[1453]&m[1454]&~m[1455]&m[1456]&m[1495])|(m[1453]&~m[1454]&m[1455]&m[1456]&m[1495])|(~m[1453]&m[1454]&m[1455]&m[1456]&m[1495]))&~BiasedRNG[844])|((m[1453]&m[1454]&~m[1455]&~m[1456]&~m[1495])|(m[1453]&~m[1454]&m[1455]&~m[1456]&~m[1495])|(~m[1453]&m[1454]&m[1455]&~m[1456]&~m[1495])|(m[1453]&m[1454]&m[1455]&~m[1456]&~m[1495])|(m[1453]&m[1454]&m[1455]&m[1456]&~m[1495])|(m[1453]&m[1454]&~m[1455]&~m[1456]&m[1495])|(m[1453]&~m[1454]&m[1455]&~m[1456]&m[1495])|(~m[1453]&m[1454]&m[1455]&~m[1456]&m[1495])|(m[1453]&m[1454]&m[1455]&~m[1456]&m[1495])|(m[1453]&m[1454]&m[1455]&m[1456]&m[1495]));
    m[1462] = (((m[1458]&~m[1459]&~m[1460]&~m[1461]&~m[1498])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1498])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1498])|(m[1458]&m[1459]&~m[1460]&m[1461]&~m[1498])|(m[1458]&~m[1459]&m[1460]&m[1461]&~m[1498])|(~m[1458]&m[1459]&m[1460]&m[1461]&~m[1498]))&BiasedRNG[845])|(((m[1458]&~m[1459]&~m[1460]&~m[1461]&m[1498])|(~m[1458]&m[1459]&~m[1460]&~m[1461]&m[1498])|(~m[1458]&~m[1459]&m[1460]&~m[1461]&m[1498])|(m[1458]&m[1459]&~m[1460]&m[1461]&m[1498])|(m[1458]&~m[1459]&m[1460]&m[1461]&m[1498])|(~m[1458]&m[1459]&m[1460]&m[1461]&m[1498]))&~BiasedRNG[845])|((m[1458]&m[1459]&~m[1460]&~m[1461]&~m[1498])|(m[1458]&~m[1459]&m[1460]&~m[1461]&~m[1498])|(~m[1458]&m[1459]&m[1460]&~m[1461]&~m[1498])|(m[1458]&m[1459]&m[1460]&~m[1461]&~m[1498])|(m[1458]&m[1459]&m[1460]&m[1461]&~m[1498])|(m[1458]&m[1459]&~m[1460]&~m[1461]&m[1498])|(m[1458]&~m[1459]&m[1460]&~m[1461]&m[1498])|(~m[1458]&m[1459]&m[1460]&~m[1461]&m[1498])|(m[1458]&m[1459]&m[1460]&~m[1461]&m[1498])|(m[1458]&m[1459]&m[1460]&m[1461]&m[1498]));
    m[1467] = (((m[1463]&~m[1464]&~m[1465]&~m[1466]&~m[1500])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1500])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1500])|(m[1463]&m[1464]&~m[1465]&m[1466]&~m[1500])|(m[1463]&~m[1464]&m[1465]&m[1466]&~m[1500])|(~m[1463]&m[1464]&m[1465]&m[1466]&~m[1500]))&BiasedRNG[846])|(((m[1463]&~m[1464]&~m[1465]&~m[1466]&m[1500])|(~m[1463]&m[1464]&~m[1465]&~m[1466]&m[1500])|(~m[1463]&~m[1464]&m[1465]&~m[1466]&m[1500])|(m[1463]&m[1464]&~m[1465]&m[1466]&m[1500])|(m[1463]&~m[1464]&m[1465]&m[1466]&m[1500])|(~m[1463]&m[1464]&m[1465]&m[1466]&m[1500]))&~BiasedRNG[846])|((m[1463]&m[1464]&~m[1465]&~m[1466]&~m[1500])|(m[1463]&~m[1464]&m[1465]&~m[1466]&~m[1500])|(~m[1463]&m[1464]&m[1465]&~m[1466]&~m[1500])|(m[1463]&m[1464]&m[1465]&~m[1466]&~m[1500])|(m[1463]&m[1464]&m[1465]&m[1466]&~m[1500])|(m[1463]&m[1464]&~m[1465]&~m[1466]&m[1500])|(m[1463]&~m[1464]&m[1465]&~m[1466]&m[1500])|(~m[1463]&m[1464]&m[1465]&~m[1466]&m[1500])|(m[1463]&m[1464]&m[1465]&~m[1466]&m[1500])|(m[1463]&m[1464]&m[1465]&m[1466]&m[1500]));
    m[1472] = (((m[1468]&~m[1469]&~m[1470]&~m[1471]&~m[1505])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1505])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1505])|(m[1468]&m[1469]&~m[1470]&m[1471]&~m[1505])|(m[1468]&~m[1469]&m[1470]&m[1471]&~m[1505])|(~m[1468]&m[1469]&m[1470]&m[1471]&~m[1505]))&BiasedRNG[847])|(((m[1468]&~m[1469]&~m[1470]&~m[1471]&m[1505])|(~m[1468]&m[1469]&~m[1470]&~m[1471]&m[1505])|(~m[1468]&~m[1469]&m[1470]&~m[1471]&m[1505])|(m[1468]&m[1469]&~m[1470]&m[1471]&m[1505])|(m[1468]&~m[1469]&m[1470]&m[1471]&m[1505])|(~m[1468]&m[1469]&m[1470]&m[1471]&m[1505]))&~BiasedRNG[847])|((m[1468]&m[1469]&~m[1470]&~m[1471]&~m[1505])|(m[1468]&~m[1469]&m[1470]&~m[1471]&~m[1505])|(~m[1468]&m[1469]&m[1470]&~m[1471]&~m[1505])|(m[1468]&m[1469]&m[1470]&~m[1471]&~m[1505])|(m[1468]&m[1469]&m[1470]&m[1471]&~m[1505])|(m[1468]&m[1469]&~m[1470]&~m[1471]&m[1505])|(m[1468]&~m[1469]&m[1470]&~m[1471]&m[1505])|(~m[1468]&m[1469]&m[1470]&~m[1471]&m[1505])|(m[1468]&m[1469]&m[1470]&~m[1471]&m[1505])|(m[1468]&m[1469]&m[1470]&m[1471]&m[1505]));
    m[1477] = (((m[1473]&~m[1474]&~m[1475]&~m[1476]&~m[1510])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1510])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1510])|(m[1473]&m[1474]&~m[1475]&m[1476]&~m[1510])|(m[1473]&~m[1474]&m[1475]&m[1476]&~m[1510])|(~m[1473]&m[1474]&m[1475]&m[1476]&~m[1510]))&BiasedRNG[848])|(((m[1473]&~m[1474]&~m[1475]&~m[1476]&m[1510])|(~m[1473]&m[1474]&~m[1475]&~m[1476]&m[1510])|(~m[1473]&~m[1474]&m[1475]&~m[1476]&m[1510])|(m[1473]&m[1474]&~m[1475]&m[1476]&m[1510])|(m[1473]&~m[1474]&m[1475]&m[1476]&m[1510])|(~m[1473]&m[1474]&m[1475]&m[1476]&m[1510]))&~BiasedRNG[848])|((m[1473]&m[1474]&~m[1475]&~m[1476]&~m[1510])|(m[1473]&~m[1474]&m[1475]&~m[1476]&~m[1510])|(~m[1473]&m[1474]&m[1475]&~m[1476]&~m[1510])|(m[1473]&m[1474]&m[1475]&~m[1476]&~m[1510])|(m[1473]&m[1474]&m[1475]&m[1476]&~m[1510])|(m[1473]&m[1474]&~m[1475]&~m[1476]&m[1510])|(m[1473]&~m[1474]&m[1475]&~m[1476]&m[1510])|(~m[1473]&m[1474]&m[1475]&~m[1476]&m[1510])|(m[1473]&m[1474]&m[1475]&~m[1476]&m[1510])|(m[1473]&m[1474]&m[1475]&m[1476]&m[1510]));
    m[1482] = (((m[1478]&~m[1479]&~m[1480]&~m[1481]&~m[1515])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1515])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1515])|(m[1478]&m[1479]&~m[1480]&m[1481]&~m[1515])|(m[1478]&~m[1479]&m[1480]&m[1481]&~m[1515])|(~m[1478]&m[1479]&m[1480]&m[1481]&~m[1515]))&BiasedRNG[849])|(((m[1478]&~m[1479]&~m[1480]&~m[1481]&m[1515])|(~m[1478]&m[1479]&~m[1480]&~m[1481]&m[1515])|(~m[1478]&~m[1479]&m[1480]&~m[1481]&m[1515])|(m[1478]&m[1479]&~m[1480]&m[1481]&m[1515])|(m[1478]&~m[1479]&m[1480]&m[1481]&m[1515])|(~m[1478]&m[1479]&m[1480]&m[1481]&m[1515]))&~BiasedRNG[849])|((m[1478]&m[1479]&~m[1480]&~m[1481]&~m[1515])|(m[1478]&~m[1479]&m[1480]&~m[1481]&~m[1515])|(~m[1478]&m[1479]&m[1480]&~m[1481]&~m[1515])|(m[1478]&m[1479]&m[1480]&~m[1481]&~m[1515])|(m[1478]&m[1479]&m[1480]&m[1481]&~m[1515])|(m[1478]&m[1479]&~m[1480]&~m[1481]&m[1515])|(m[1478]&~m[1479]&m[1480]&~m[1481]&m[1515])|(~m[1478]&m[1479]&m[1480]&~m[1481]&m[1515])|(m[1478]&m[1479]&m[1480]&~m[1481]&m[1515])|(m[1478]&m[1479]&m[1480]&m[1481]&m[1515]));
    m[1487] = (((m[1483]&~m[1484]&~m[1485]&~m[1486]&~m[1520])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1520])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1520])|(m[1483]&m[1484]&~m[1485]&m[1486]&~m[1520])|(m[1483]&~m[1484]&m[1485]&m[1486]&~m[1520])|(~m[1483]&m[1484]&m[1485]&m[1486]&~m[1520]))&BiasedRNG[850])|(((m[1483]&~m[1484]&~m[1485]&~m[1486]&m[1520])|(~m[1483]&m[1484]&~m[1485]&~m[1486]&m[1520])|(~m[1483]&~m[1484]&m[1485]&~m[1486]&m[1520])|(m[1483]&m[1484]&~m[1485]&m[1486]&m[1520])|(m[1483]&~m[1484]&m[1485]&m[1486]&m[1520])|(~m[1483]&m[1484]&m[1485]&m[1486]&m[1520]))&~BiasedRNG[850])|((m[1483]&m[1484]&~m[1485]&~m[1486]&~m[1520])|(m[1483]&~m[1484]&m[1485]&~m[1486]&~m[1520])|(~m[1483]&m[1484]&m[1485]&~m[1486]&~m[1520])|(m[1483]&m[1484]&m[1485]&~m[1486]&~m[1520])|(m[1483]&m[1484]&m[1485]&m[1486]&~m[1520])|(m[1483]&m[1484]&~m[1485]&~m[1486]&m[1520])|(m[1483]&~m[1484]&m[1485]&~m[1486]&m[1520])|(~m[1483]&m[1484]&m[1485]&~m[1486]&m[1520])|(m[1483]&m[1484]&m[1485]&~m[1486]&m[1520])|(m[1483]&m[1484]&m[1485]&m[1486]&m[1520]));
    m[1492] = (((m[1488]&~m[1489]&~m[1490]&~m[1491]&~m[1525])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1525])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1525])|(m[1488]&m[1489]&~m[1490]&m[1491]&~m[1525])|(m[1488]&~m[1489]&m[1490]&m[1491]&~m[1525])|(~m[1488]&m[1489]&m[1490]&m[1491]&~m[1525]))&BiasedRNG[851])|(((m[1488]&~m[1489]&~m[1490]&~m[1491]&m[1525])|(~m[1488]&m[1489]&~m[1490]&~m[1491]&m[1525])|(~m[1488]&~m[1489]&m[1490]&~m[1491]&m[1525])|(m[1488]&m[1489]&~m[1490]&m[1491]&m[1525])|(m[1488]&~m[1489]&m[1490]&m[1491]&m[1525])|(~m[1488]&m[1489]&m[1490]&m[1491]&m[1525]))&~BiasedRNG[851])|((m[1488]&m[1489]&~m[1490]&~m[1491]&~m[1525])|(m[1488]&~m[1489]&m[1490]&~m[1491]&~m[1525])|(~m[1488]&m[1489]&m[1490]&~m[1491]&~m[1525])|(m[1488]&m[1489]&m[1490]&~m[1491]&~m[1525])|(m[1488]&m[1489]&m[1490]&m[1491]&~m[1525])|(m[1488]&m[1489]&~m[1490]&~m[1491]&m[1525])|(m[1488]&~m[1489]&m[1490]&~m[1491]&m[1525])|(~m[1488]&m[1489]&m[1490]&~m[1491]&m[1525])|(m[1488]&m[1489]&m[1490]&~m[1491]&m[1525])|(m[1488]&m[1489]&m[1490]&m[1491]&m[1525]));
    m[1497] = (((m[1493]&~m[1494]&~m[1495]&~m[1496]&~m[1530])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1530])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1530])|(m[1493]&m[1494]&~m[1495]&m[1496]&~m[1530])|(m[1493]&~m[1494]&m[1495]&m[1496]&~m[1530])|(~m[1493]&m[1494]&m[1495]&m[1496]&~m[1530]))&BiasedRNG[852])|(((m[1493]&~m[1494]&~m[1495]&~m[1496]&m[1530])|(~m[1493]&m[1494]&~m[1495]&~m[1496]&m[1530])|(~m[1493]&~m[1494]&m[1495]&~m[1496]&m[1530])|(m[1493]&m[1494]&~m[1495]&m[1496]&m[1530])|(m[1493]&~m[1494]&m[1495]&m[1496]&m[1530])|(~m[1493]&m[1494]&m[1495]&m[1496]&m[1530]))&~BiasedRNG[852])|((m[1493]&m[1494]&~m[1495]&~m[1496]&~m[1530])|(m[1493]&~m[1494]&m[1495]&~m[1496]&~m[1530])|(~m[1493]&m[1494]&m[1495]&~m[1496]&~m[1530])|(m[1493]&m[1494]&m[1495]&~m[1496]&~m[1530])|(m[1493]&m[1494]&m[1495]&m[1496]&~m[1530])|(m[1493]&m[1494]&~m[1495]&~m[1496]&m[1530])|(m[1493]&~m[1494]&m[1495]&~m[1496]&m[1530])|(~m[1493]&m[1494]&m[1495]&~m[1496]&m[1530])|(m[1493]&m[1494]&m[1495]&~m[1496]&m[1530])|(m[1493]&m[1494]&m[1495]&m[1496]&m[1530]));
    m[1502] = (((m[1498]&~m[1499]&~m[1500]&~m[1501]&~m[1533])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1533])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1533])|(m[1498]&m[1499]&~m[1500]&m[1501]&~m[1533])|(m[1498]&~m[1499]&m[1500]&m[1501]&~m[1533])|(~m[1498]&m[1499]&m[1500]&m[1501]&~m[1533]))&BiasedRNG[853])|(((m[1498]&~m[1499]&~m[1500]&~m[1501]&m[1533])|(~m[1498]&m[1499]&~m[1500]&~m[1501]&m[1533])|(~m[1498]&~m[1499]&m[1500]&~m[1501]&m[1533])|(m[1498]&m[1499]&~m[1500]&m[1501]&m[1533])|(m[1498]&~m[1499]&m[1500]&m[1501]&m[1533])|(~m[1498]&m[1499]&m[1500]&m[1501]&m[1533]))&~BiasedRNG[853])|((m[1498]&m[1499]&~m[1500]&~m[1501]&~m[1533])|(m[1498]&~m[1499]&m[1500]&~m[1501]&~m[1533])|(~m[1498]&m[1499]&m[1500]&~m[1501]&~m[1533])|(m[1498]&m[1499]&m[1500]&~m[1501]&~m[1533])|(m[1498]&m[1499]&m[1500]&m[1501]&~m[1533])|(m[1498]&m[1499]&~m[1500]&~m[1501]&m[1533])|(m[1498]&~m[1499]&m[1500]&~m[1501]&m[1533])|(~m[1498]&m[1499]&m[1500]&~m[1501]&m[1533])|(m[1498]&m[1499]&m[1500]&~m[1501]&m[1533])|(m[1498]&m[1499]&m[1500]&m[1501]&m[1533]));
    m[1507] = (((m[1503]&~m[1504]&~m[1505]&~m[1506]&~m[1535])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1535])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1535])|(m[1503]&m[1504]&~m[1505]&m[1506]&~m[1535])|(m[1503]&~m[1504]&m[1505]&m[1506]&~m[1535])|(~m[1503]&m[1504]&m[1505]&m[1506]&~m[1535]))&BiasedRNG[854])|(((m[1503]&~m[1504]&~m[1505]&~m[1506]&m[1535])|(~m[1503]&m[1504]&~m[1505]&~m[1506]&m[1535])|(~m[1503]&~m[1504]&m[1505]&~m[1506]&m[1535])|(m[1503]&m[1504]&~m[1505]&m[1506]&m[1535])|(m[1503]&~m[1504]&m[1505]&m[1506]&m[1535])|(~m[1503]&m[1504]&m[1505]&m[1506]&m[1535]))&~BiasedRNG[854])|((m[1503]&m[1504]&~m[1505]&~m[1506]&~m[1535])|(m[1503]&~m[1504]&m[1505]&~m[1506]&~m[1535])|(~m[1503]&m[1504]&m[1505]&~m[1506]&~m[1535])|(m[1503]&m[1504]&m[1505]&~m[1506]&~m[1535])|(m[1503]&m[1504]&m[1505]&m[1506]&~m[1535])|(m[1503]&m[1504]&~m[1505]&~m[1506]&m[1535])|(m[1503]&~m[1504]&m[1505]&~m[1506]&m[1535])|(~m[1503]&m[1504]&m[1505]&~m[1506]&m[1535])|(m[1503]&m[1504]&m[1505]&~m[1506]&m[1535])|(m[1503]&m[1504]&m[1505]&m[1506]&m[1535]));
    m[1512] = (((m[1508]&~m[1509]&~m[1510]&~m[1511]&~m[1540])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1540])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1540])|(m[1508]&m[1509]&~m[1510]&m[1511]&~m[1540])|(m[1508]&~m[1509]&m[1510]&m[1511]&~m[1540])|(~m[1508]&m[1509]&m[1510]&m[1511]&~m[1540]))&BiasedRNG[855])|(((m[1508]&~m[1509]&~m[1510]&~m[1511]&m[1540])|(~m[1508]&m[1509]&~m[1510]&~m[1511]&m[1540])|(~m[1508]&~m[1509]&m[1510]&~m[1511]&m[1540])|(m[1508]&m[1509]&~m[1510]&m[1511]&m[1540])|(m[1508]&~m[1509]&m[1510]&m[1511]&m[1540])|(~m[1508]&m[1509]&m[1510]&m[1511]&m[1540]))&~BiasedRNG[855])|((m[1508]&m[1509]&~m[1510]&~m[1511]&~m[1540])|(m[1508]&~m[1509]&m[1510]&~m[1511]&~m[1540])|(~m[1508]&m[1509]&m[1510]&~m[1511]&~m[1540])|(m[1508]&m[1509]&m[1510]&~m[1511]&~m[1540])|(m[1508]&m[1509]&m[1510]&m[1511]&~m[1540])|(m[1508]&m[1509]&~m[1510]&~m[1511]&m[1540])|(m[1508]&~m[1509]&m[1510]&~m[1511]&m[1540])|(~m[1508]&m[1509]&m[1510]&~m[1511]&m[1540])|(m[1508]&m[1509]&m[1510]&~m[1511]&m[1540])|(m[1508]&m[1509]&m[1510]&m[1511]&m[1540]));
    m[1517] = (((m[1513]&~m[1514]&~m[1515]&~m[1516]&~m[1545])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1545])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1545])|(m[1513]&m[1514]&~m[1515]&m[1516]&~m[1545])|(m[1513]&~m[1514]&m[1515]&m[1516]&~m[1545])|(~m[1513]&m[1514]&m[1515]&m[1516]&~m[1545]))&BiasedRNG[856])|(((m[1513]&~m[1514]&~m[1515]&~m[1516]&m[1545])|(~m[1513]&m[1514]&~m[1515]&~m[1516]&m[1545])|(~m[1513]&~m[1514]&m[1515]&~m[1516]&m[1545])|(m[1513]&m[1514]&~m[1515]&m[1516]&m[1545])|(m[1513]&~m[1514]&m[1515]&m[1516]&m[1545])|(~m[1513]&m[1514]&m[1515]&m[1516]&m[1545]))&~BiasedRNG[856])|((m[1513]&m[1514]&~m[1515]&~m[1516]&~m[1545])|(m[1513]&~m[1514]&m[1515]&~m[1516]&~m[1545])|(~m[1513]&m[1514]&m[1515]&~m[1516]&~m[1545])|(m[1513]&m[1514]&m[1515]&~m[1516]&~m[1545])|(m[1513]&m[1514]&m[1515]&m[1516]&~m[1545])|(m[1513]&m[1514]&~m[1515]&~m[1516]&m[1545])|(m[1513]&~m[1514]&m[1515]&~m[1516]&m[1545])|(~m[1513]&m[1514]&m[1515]&~m[1516]&m[1545])|(m[1513]&m[1514]&m[1515]&~m[1516]&m[1545])|(m[1513]&m[1514]&m[1515]&m[1516]&m[1545]));
    m[1522] = (((m[1518]&~m[1519]&~m[1520]&~m[1521]&~m[1550])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1550])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1550])|(m[1518]&m[1519]&~m[1520]&m[1521]&~m[1550])|(m[1518]&~m[1519]&m[1520]&m[1521]&~m[1550])|(~m[1518]&m[1519]&m[1520]&m[1521]&~m[1550]))&BiasedRNG[857])|(((m[1518]&~m[1519]&~m[1520]&~m[1521]&m[1550])|(~m[1518]&m[1519]&~m[1520]&~m[1521]&m[1550])|(~m[1518]&~m[1519]&m[1520]&~m[1521]&m[1550])|(m[1518]&m[1519]&~m[1520]&m[1521]&m[1550])|(m[1518]&~m[1519]&m[1520]&m[1521]&m[1550])|(~m[1518]&m[1519]&m[1520]&m[1521]&m[1550]))&~BiasedRNG[857])|((m[1518]&m[1519]&~m[1520]&~m[1521]&~m[1550])|(m[1518]&~m[1519]&m[1520]&~m[1521]&~m[1550])|(~m[1518]&m[1519]&m[1520]&~m[1521]&~m[1550])|(m[1518]&m[1519]&m[1520]&~m[1521]&~m[1550])|(m[1518]&m[1519]&m[1520]&m[1521]&~m[1550])|(m[1518]&m[1519]&~m[1520]&~m[1521]&m[1550])|(m[1518]&~m[1519]&m[1520]&~m[1521]&m[1550])|(~m[1518]&m[1519]&m[1520]&~m[1521]&m[1550])|(m[1518]&m[1519]&m[1520]&~m[1521]&m[1550])|(m[1518]&m[1519]&m[1520]&m[1521]&m[1550]));
    m[1527] = (((m[1523]&~m[1524]&~m[1525]&~m[1526]&~m[1555])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1555])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1555])|(m[1523]&m[1524]&~m[1525]&m[1526]&~m[1555])|(m[1523]&~m[1524]&m[1525]&m[1526]&~m[1555])|(~m[1523]&m[1524]&m[1525]&m[1526]&~m[1555]))&BiasedRNG[858])|(((m[1523]&~m[1524]&~m[1525]&~m[1526]&m[1555])|(~m[1523]&m[1524]&~m[1525]&~m[1526]&m[1555])|(~m[1523]&~m[1524]&m[1525]&~m[1526]&m[1555])|(m[1523]&m[1524]&~m[1525]&m[1526]&m[1555])|(m[1523]&~m[1524]&m[1525]&m[1526]&m[1555])|(~m[1523]&m[1524]&m[1525]&m[1526]&m[1555]))&~BiasedRNG[858])|((m[1523]&m[1524]&~m[1525]&~m[1526]&~m[1555])|(m[1523]&~m[1524]&m[1525]&~m[1526]&~m[1555])|(~m[1523]&m[1524]&m[1525]&~m[1526]&~m[1555])|(m[1523]&m[1524]&m[1525]&~m[1526]&~m[1555])|(m[1523]&m[1524]&m[1525]&m[1526]&~m[1555])|(m[1523]&m[1524]&~m[1525]&~m[1526]&m[1555])|(m[1523]&~m[1524]&m[1525]&~m[1526]&m[1555])|(~m[1523]&m[1524]&m[1525]&~m[1526]&m[1555])|(m[1523]&m[1524]&m[1525]&~m[1526]&m[1555])|(m[1523]&m[1524]&m[1525]&m[1526]&m[1555]));
    m[1532] = (((m[1528]&~m[1529]&~m[1530]&~m[1531]&~m[1560])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1560])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1560])|(m[1528]&m[1529]&~m[1530]&m[1531]&~m[1560])|(m[1528]&~m[1529]&m[1530]&m[1531]&~m[1560])|(~m[1528]&m[1529]&m[1530]&m[1531]&~m[1560]))&BiasedRNG[859])|(((m[1528]&~m[1529]&~m[1530]&~m[1531]&m[1560])|(~m[1528]&m[1529]&~m[1530]&~m[1531]&m[1560])|(~m[1528]&~m[1529]&m[1530]&~m[1531]&m[1560])|(m[1528]&m[1529]&~m[1530]&m[1531]&m[1560])|(m[1528]&~m[1529]&m[1530]&m[1531]&m[1560])|(~m[1528]&m[1529]&m[1530]&m[1531]&m[1560]))&~BiasedRNG[859])|((m[1528]&m[1529]&~m[1530]&~m[1531]&~m[1560])|(m[1528]&~m[1529]&m[1530]&~m[1531]&~m[1560])|(~m[1528]&m[1529]&m[1530]&~m[1531]&~m[1560])|(m[1528]&m[1529]&m[1530]&~m[1531]&~m[1560])|(m[1528]&m[1529]&m[1530]&m[1531]&~m[1560])|(m[1528]&m[1529]&~m[1530]&~m[1531]&m[1560])|(m[1528]&~m[1529]&m[1530]&~m[1531]&m[1560])|(~m[1528]&m[1529]&m[1530]&~m[1531]&m[1560])|(m[1528]&m[1529]&m[1530]&~m[1531]&m[1560])|(m[1528]&m[1529]&m[1530]&m[1531]&m[1560]));
    m[1537] = (((m[1533]&~m[1534]&~m[1535]&~m[1536]&~m[1563])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1563])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1563])|(m[1533]&m[1534]&~m[1535]&m[1536]&~m[1563])|(m[1533]&~m[1534]&m[1535]&m[1536]&~m[1563])|(~m[1533]&m[1534]&m[1535]&m[1536]&~m[1563]))&BiasedRNG[860])|(((m[1533]&~m[1534]&~m[1535]&~m[1536]&m[1563])|(~m[1533]&m[1534]&~m[1535]&~m[1536]&m[1563])|(~m[1533]&~m[1534]&m[1535]&~m[1536]&m[1563])|(m[1533]&m[1534]&~m[1535]&m[1536]&m[1563])|(m[1533]&~m[1534]&m[1535]&m[1536]&m[1563])|(~m[1533]&m[1534]&m[1535]&m[1536]&m[1563]))&~BiasedRNG[860])|((m[1533]&m[1534]&~m[1535]&~m[1536]&~m[1563])|(m[1533]&~m[1534]&m[1535]&~m[1536]&~m[1563])|(~m[1533]&m[1534]&m[1535]&~m[1536]&~m[1563])|(m[1533]&m[1534]&m[1535]&~m[1536]&~m[1563])|(m[1533]&m[1534]&m[1535]&m[1536]&~m[1563])|(m[1533]&m[1534]&~m[1535]&~m[1536]&m[1563])|(m[1533]&~m[1534]&m[1535]&~m[1536]&m[1563])|(~m[1533]&m[1534]&m[1535]&~m[1536]&m[1563])|(m[1533]&m[1534]&m[1535]&~m[1536]&m[1563])|(m[1533]&m[1534]&m[1535]&m[1536]&m[1563]));
    m[1542] = (((m[1538]&~m[1539]&~m[1540]&~m[1541]&~m[1565])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1565])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1565])|(m[1538]&m[1539]&~m[1540]&m[1541]&~m[1565])|(m[1538]&~m[1539]&m[1540]&m[1541]&~m[1565])|(~m[1538]&m[1539]&m[1540]&m[1541]&~m[1565]))&BiasedRNG[861])|(((m[1538]&~m[1539]&~m[1540]&~m[1541]&m[1565])|(~m[1538]&m[1539]&~m[1540]&~m[1541]&m[1565])|(~m[1538]&~m[1539]&m[1540]&~m[1541]&m[1565])|(m[1538]&m[1539]&~m[1540]&m[1541]&m[1565])|(m[1538]&~m[1539]&m[1540]&m[1541]&m[1565])|(~m[1538]&m[1539]&m[1540]&m[1541]&m[1565]))&~BiasedRNG[861])|((m[1538]&m[1539]&~m[1540]&~m[1541]&~m[1565])|(m[1538]&~m[1539]&m[1540]&~m[1541]&~m[1565])|(~m[1538]&m[1539]&m[1540]&~m[1541]&~m[1565])|(m[1538]&m[1539]&m[1540]&~m[1541]&~m[1565])|(m[1538]&m[1539]&m[1540]&m[1541]&~m[1565])|(m[1538]&m[1539]&~m[1540]&~m[1541]&m[1565])|(m[1538]&~m[1539]&m[1540]&~m[1541]&m[1565])|(~m[1538]&m[1539]&m[1540]&~m[1541]&m[1565])|(m[1538]&m[1539]&m[1540]&~m[1541]&m[1565])|(m[1538]&m[1539]&m[1540]&m[1541]&m[1565]));
    m[1547] = (((m[1543]&~m[1544]&~m[1545]&~m[1546]&~m[1570])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1570])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1570])|(m[1543]&m[1544]&~m[1545]&m[1546]&~m[1570])|(m[1543]&~m[1544]&m[1545]&m[1546]&~m[1570])|(~m[1543]&m[1544]&m[1545]&m[1546]&~m[1570]))&BiasedRNG[862])|(((m[1543]&~m[1544]&~m[1545]&~m[1546]&m[1570])|(~m[1543]&m[1544]&~m[1545]&~m[1546]&m[1570])|(~m[1543]&~m[1544]&m[1545]&~m[1546]&m[1570])|(m[1543]&m[1544]&~m[1545]&m[1546]&m[1570])|(m[1543]&~m[1544]&m[1545]&m[1546]&m[1570])|(~m[1543]&m[1544]&m[1545]&m[1546]&m[1570]))&~BiasedRNG[862])|((m[1543]&m[1544]&~m[1545]&~m[1546]&~m[1570])|(m[1543]&~m[1544]&m[1545]&~m[1546]&~m[1570])|(~m[1543]&m[1544]&m[1545]&~m[1546]&~m[1570])|(m[1543]&m[1544]&m[1545]&~m[1546]&~m[1570])|(m[1543]&m[1544]&m[1545]&m[1546]&~m[1570])|(m[1543]&m[1544]&~m[1545]&~m[1546]&m[1570])|(m[1543]&~m[1544]&m[1545]&~m[1546]&m[1570])|(~m[1543]&m[1544]&m[1545]&~m[1546]&m[1570])|(m[1543]&m[1544]&m[1545]&~m[1546]&m[1570])|(m[1543]&m[1544]&m[1545]&m[1546]&m[1570]));
    m[1552] = (((m[1548]&~m[1549]&~m[1550]&~m[1551]&~m[1575])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1575])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1575])|(m[1548]&m[1549]&~m[1550]&m[1551]&~m[1575])|(m[1548]&~m[1549]&m[1550]&m[1551]&~m[1575])|(~m[1548]&m[1549]&m[1550]&m[1551]&~m[1575]))&BiasedRNG[863])|(((m[1548]&~m[1549]&~m[1550]&~m[1551]&m[1575])|(~m[1548]&m[1549]&~m[1550]&~m[1551]&m[1575])|(~m[1548]&~m[1549]&m[1550]&~m[1551]&m[1575])|(m[1548]&m[1549]&~m[1550]&m[1551]&m[1575])|(m[1548]&~m[1549]&m[1550]&m[1551]&m[1575])|(~m[1548]&m[1549]&m[1550]&m[1551]&m[1575]))&~BiasedRNG[863])|((m[1548]&m[1549]&~m[1550]&~m[1551]&~m[1575])|(m[1548]&~m[1549]&m[1550]&~m[1551]&~m[1575])|(~m[1548]&m[1549]&m[1550]&~m[1551]&~m[1575])|(m[1548]&m[1549]&m[1550]&~m[1551]&~m[1575])|(m[1548]&m[1549]&m[1550]&m[1551]&~m[1575])|(m[1548]&m[1549]&~m[1550]&~m[1551]&m[1575])|(m[1548]&~m[1549]&m[1550]&~m[1551]&m[1575])|(~m[1548]&m[1549]&m[1550]&~m[1551]&m[1575])|(m[1548]&m[1549]&m[1550]&~m[1551]&m[1575])|(m[1548]&m[1549]&m[1550]&m[1551]&m[1575]));
    m[1557] = (((m[1553]&~m[1554]&~m[1555]&~m[1556]&~m[1580])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1580])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1580])|(m[1553]&m[1554]&~m[1555]&m[1556]&~m[1580])|(m[1553]&~m[1554]&m[1555]&m[1556]&~m[1580])|(~m[1553]&m[1554]&m[1555]&m[1556]&~m[1580]))&BiasedRNG[864])|(((m[1553]&~m[1554]&~m[1555]&~m[1556]&m[1580])|(~m[1553]&m[1554]&~m[1555]&~m[1556]&m[1580])|(~m[1553]&~m[1554]&m[1555]&~m[1556]&m[1580])|(m[1553]&m[1554]&~m[1555]&m[1556]&m[1580])|(m[1553]&~m[1554]&m[1555]&m[1556]&m[1580])|(~m[1553]&m[1554]&m[1555]&m[1556]&m[1580]))&~BiasedRNG[864])|((m[1553]&m[1554]&~m[1555]&~m[1556]&~m[1580])|(m[1553]&~m[1554]&m[1555]&~m[1556]&~m[1580])|(~m[1553]&m[1554]&m[1555]&~m[1556]&~m[1580])|(m[1553]&m[1554]&m[1555]&~m[1556]&~m[1580])|(m[1553]&m[1554]&m[1555]&m[1556]&~m[1580])|(m[1553]&m[1554]&~m[1555]&~m[1556]&m[1580])|(m[1553]&~m[1554]&m[1555]&~m[1556]&m[1580])|(~m[1553]&m[1554]&m[1555]&~m[1556]&m[1580])|(m[1553]&m[1554]&m[1555]&~m[1556]&m[1580])|(m[1553]&m[1554]&m[1555]&m[1556]&m[1580]));
    m[1562] = (((m[1558]&~m[1559]&~m[1560]&~m[1561]&~m[1585])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1585])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1585])|(m[1558]&m[1559]&~m[1560]&m[1561]&~m[1585])|(m[1558]&~m[1559]&m[1560]&m[1561]&~m[1585])|(~m[1558]&m[1559]&m[1560]&m[1561]&~m[1585]))&BiasedRNG[865])|(((m[1558]&~m[1559]&~m[1560]&~m[1561]&m[1585])|(~m[1558]&m[1559]&~m[1560]&~m[1561]&m[1585])|(~m[1558]&~m[1559]&m[1560]&~m[1561]&m[1585])|(m[1558]&m[1559]&~m[1560]&m[1561]&m[1585])|(m[1558]&~m[1559]&m[1560]&m[1561]&m[1585])|(~m[1558]&m[1559]&m[1560]&m[1561]&m[1585]))&~BiasedRNG[865])|((m[1558]&m[1559]&~m[1560]&~m[1561]&~m[1585])|(m[1558]&~m[1559]&m[1560]&~m[1561]&~m[1585])|(~m[1558]&m[1559]&m[1560]&~m[1561]&~m[1585])|(m[1558]&m[1559]&m[1560]&~m[1561]&~m[1585])|(m[1558]&m[1559]&m[1560]&m[1561]&~m[1585])|(m[1558]&m[1559]&~m[1560]&~m[1561]&m[1585])|(m[1558]&~m[1559]&m[1560]&~m[1561]&m[1585])|(~m[1558]&m[1559]&m[1560]&~m[1561]&m[1585])|(m[1558]&m[1559]&m[1560]&~m[1561]&m[1585])|(m[1558]&m[1559]&m[1560]&m[1561]&m[1585]));
    m[1567] = (((m[1563]&~m[1564]&~m[1565]&~m[1566]&~m[1588])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1588])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1588])|(m[1563]&m[1564]&~m[1565]&m[1566]&~m[1588])|(m[1563]&~m[1564]&m[1565]&m[1566]&~m[1588])|(~m[1563]&m[1564]&m[1565]&m[1566]&~m[1588]))&BiasedRNG[866])|(((m[1563]&~m[1564]&~m[1565]&~m[1566]&m[1588])|(~m[1563]&m[1564]&~m[1565]&~m[1566]&m[1588])|(~m[1563]&~m[1564]&m[1565]&~m[1566]&m[1588])|(m[1563]&m[1564]&~m[1565]&m[1566]&m[1588])|(m[1563]&~m[1564]&m[1565]&m[1566]&m[1588])|(~m[1563]&m[1564]&m[1565]&m[1566]&m[1588]))&~BiasedRNG[866])|((m[1563]&m[1564]&~m[1565]&~m[1566]&~m[1588])|(m[1563]&~m[1564]&m[1565]&~m[1566]&~m[1588])|(~m[1563]&m[1564]&m[1565]&~m[1566]&~m[1588])|(m[1563]&m[1564]&m[1565]&~m[1566]&~m[1588])|(m[1563]&m[1564]&m[1565]&m[1566]&~m[1588])|(m[1563]&m[1564]&~m[1565]&~m[1566]&m[1588])|(m[1563]&~m[1564]&m[1565]&~m[1566]&m[1588])|(~m[1563]&m[1564]&m[1565]&~m[1566]&m[1588])|(m[1563]&m[1564]&m[1565]&~m[1566]&m[1588])|(m[1563]&m[1564]&m[1565]&m[1566]&m[1588]));
    m[1572] = (((m[1568]&~m[1569]&~m[1570]&~m[1571]&~m[1590])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1590])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1590])|(m[1568]&m[1569]&~m[1570]&m[1571]&~m[1590])|(m[1568]&~m[1569]&m[1570]&m[1571]&~m[1590])|(~m[1568]&m[1569]&m[1570]&m[1571]&~m[1590]))&BiasedRNG[867])|(((m[1568]&~m[1569]&~m[1570]&~m[1571]&m[1590])|(~m[1568]&m[1569]&~m[1570]&~m[1571]&m[1590])|(~m[1568]&~m[1569]&m[1570]&~m[1571]&m[1590])|(m[1568]&m[1569]&~m[1570]&m[1571]&m[1590])|(m[1568]&~m[1569]&m[1570]&m[1571]&m[1590])|(~m[1568]&m[1569]&m[1570]&m[1571]&m[1590]))&~BiasedRNG[867])|((m[1568]&m[1569]&~m[1570]&~m[1571]&~m[1590])|(m[1568]&~m[1569]&m[1570]&~m[1571]&~m[1590])|(~m[1568]&m[1569]&m[1570]&~m[1571]&~m[1590])|(m[1568]&m[1569]&m[1570]&~m[1571]&~m[1590])|(m[1568]&m[1569]&m[1570]&m[1571]&~m[1590])|(m[1568]&m[1569]&~m[1570]&~m[1571]&m[1590])|(m[1568]&~m[1569]&m[1570]&~m[1571]&m[1590])|(~m[1568]&m[1569]&m[1570]&~m[1571]&m[1590])|(m[1568]&m[1569]&m[1570]&~m[1571]&m[1590])|(m[1568]&m[1569]&m[1570]&m[1571]&m[1590]));
    m[1577] = (((m[1573]&~m[1574]&~m[1575]&~m[1576]&~m[1595])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1595])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1595])|(m[1573]&m[1574]&~m[1575]&m[1576]&~m[1595])|(m[1573]&~m[1574]&m[1575]&m[1576]&~m[1595])|(~m[1573]&m[1574]&m[1575]&m[1576]&~m[1595]))&BiasedRNG[868])|(((m[1573]&~m[1574]&~m[1575]&~m[1576]&m[1595])|(~m[1573]&m[1574]&~m[1575]&~m[1576]&m[1595])|(~m[1573]&~m[1574]&m[1575]&~m[1576]&m[1595])|(m[1573]&m[1574]&~m[1575]&m[1576]&m[1595])|(m[1573]&~m[1574]&m[1575]&m[1576]&m[1595])|(~m[1573]&m[1574]&m[1575]&m[1576]&m[1595]))&~BiasedRNG[868])|((m[1573]&m[1574]&~m[1575]&~m[1576]&~m[1595])|(m[1573]&~m[1574]&m[1575]&~m[1576]&~m[1595])|(~m[1573]&m[1574]&m[1575]&~m[1576]&~m[1595])|(m[1573]&m[1574]&m[1575]&~m[1576]&~m[1595])|(m[1573]&m[1574]&m[1575]&m[1576]&~m[1595])|(m[1573]&m[1574]&~m[1575]&~m[1576]&m[1595])|(m[1573]&~m[1574]&m[1575]&~m[1576]&m[1595])|(~m[1573]&m[1574]&m[1575]&~m[1576]&m[1595])|(m[1573]&m[1574]&m[1575]&~m[1576]&m[1595])|(m[1573]&m[1574]&m[1575]&m[1576]&m[1595]));
    m[1582] = (((m[1578]&~m[1579]&~m[1580]&~m[1581]&~m[1600])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1600])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1600])|(m[1578]&m[1579]&~m[1580]&m[1581]&~m[1600])|(m[1578]&~m[1579]&m[1580]&m[1581]&~m[1600])|(~m[1578]&m[1579]&m[1580]&m[1581]&~m[1600]))&BiasedRNG[869])|(((m[1578]&~m[1579]&~m[1580]&~m[1581]&m[1600])|(~m[1578]&m[1579]&~m[1580]&~m[1581]&m[1600])|(~m[1578]&~m[1579]&m[1580]&~m[1581]&m[1600])|(m[1578]&m[1579]&~m[1580]&m[1581]&m[1600])|(m[1578]&~m[1579]&m[1580]&m[1581]&m[1600])|(~m[1578]&m[1579]&m[1580]&m[1581]&m[1600]))&~BiasedRNG[869])|((m[1578]&m[1579]&~m[1580]&~m[1581]&~m[1600])|(m[1578]&~m[1579]&m[1580]&~m[1581]&~m[1600])|(~m[1578]&m[1579]&m[1580]&~m[1581]&~m[1600])|(m[1578]&m[1579]&m[1580]&~m[1581]&~m[1600])|(m[1578]&m[1579]&m[1580]&m[1581]&~m[1600])|(m[1578]&m[1579]&~m[1580]&~m[1581]&m[1600])|(m[1578]&~m[1579]&m[1580]&~m[1581]&m[1600])|(~m[1578]&m[1579]&m[1580]&~m[1581]&m[1600])|(m[1578]&m[1579]&m[1580]&~m[1581]&m[1600])|(m[1578]&m[1579]&m[1580]&m[1581]&m[1600]));
    m[1587] = (((m[1583]&~m[1584]&~m[1585]&~m[1586]&~m[1605])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1605])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1605])|(m[1583]&m[1584]&~m[1585]&m[1586]&~m[1605])|(m[1583]&~m[1584]&m[1585]&m[1586]&~m[1605])|(~m[1583]&m[1584]&m[1585]&m[1586]&~m[1605]))&BiasedRNG[870])|(((m[1583]&~m[1584]&~m[1585]&~m[1586]&m[1605])|(~m[1583]&m[1584]&~m[1585]&~m[1586]&m[1605])|(~m[1583]&~m[1584]&m[1585]&~m[1586]&m[1605])|(m[1583]&m[1584]&~m[1585]&m[1586]&m[1605])|(m[1583]&~m[1584]&m[1585]&m[1586]&m[1605])|(~m[1583]&m[1584]&m[1585]&m[1586]&m[1605]))&~BiasedRNG[870])|((m[1583]&m[1584]&~m[1585]&~m[1586]&~m[1605])|(m[1583]&~m[1584]&m[1585]&~m[1586]&~m[1605])|(~m[1583]&m[1584]&m[1585]&~m[1586]&~m[1605])|(m[1583]&m[1584]&m[1585]&~m[1586]&~m[1605])|(m[1583]&m[1584]&m[1585]&m[1586]&~m[1605])|(m[1583]&m[1584]&~m[1585]&~m[1586]&m[1605])|(m[1583]&~m[1584]&m[1585]&~m[1586]&m[1605])|(~m[1583]&m[1584]&m[1585]&~m[1586]&m[1605])|(m[1583]&m[1584]&m[1585]&~m[1586]&m[1605])|(m[1583]&m[1584]&m[1585]&m[1586]&m[1605]));
    m[1592] = (((m[1588]&~m[1589]&~m[1590]&~m[1591]&~m[1608])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1608])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1608])|(m[1588]&m[1589]&~m[1590]&m[1591]&~m[1608])|(m[1588]&~m[1589]&m[1590]&m[1591]&~m[1608])|(~m[1588]&m[1589]&m[1590]&m[1591]&~m[1608]))&BiasedRNG[871])|(((m[1588]&~m[1589]&~m[1590]&~m[1591]&m[1608])|(~m[1588]&m[1589]&~m[1590]&~m[1591]&m[1608])|(~m[1588]&~m[1589]&m[1590]&~m[1591]&m[1608])|(m[1588]&m[1589]&~m[1590]&m[1591]&m[1608])|(m[1588]&~m[1589]&m[1590]&m[1591]&m[1608])|(~m[1588]&m[1589]&m[1590]&m[1591]&m[1608]))&~BiasedRNG[871])|((m[1588]&m[1589]&~m[1590]&~m[1591]&~m[1608])|(m[1588]&~m[1589]&m[1590]&~m[1591]&~m[1608])|(~m[1588]&m[1589]&m[1590]&~m[1591]&~m[1608])|(m[1588]&m[1589]&m[1590]&~m[1591]&~m[1608])|(m[1588]&m[1589]&m[1590]&m[1591]&~m[1608])|(m[1588]&m[1589]&~m[1590]&~m[1591]&m[1608])|(m[1588]&~m[1589]&m[1590]&~m[1591]&m[1608])|(~m[1588]&m[1589]&m[1590]&~m[1591]&m[1608])|(m[1588]&m[1589]&m[1590]&~m[1591]&m[1608])|(m[1588]&m[1589]&m[1590]&m[1591]&m[1608]));
    m[1597] = (((m[1593]&~m[1594]&~m[1595]&~m[1596]&~m[1610])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1610])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1610])|(m[1593]&m[1594]&~m[1595]&m[1596]&~m[1610])|(m[1593]&~m[1594]&m[1595]&m[1596]&~m[1610])|(~m[1593]&m[1594]&m[1595]&m[1596]&~m[1610]))&BiasedRNG[872])|(((m[1593]&~m[1594]&~m[1595]&~m[1596]&m[1610])|(~m[1593]&m[1594]&~m[1595]&~m[1596]&m[1610])|(~m[1593]&~m[1594]&m[1595]&~m[1596]&m[1610])|(m[1593]&m[1594]&~m[1595]&m[1596]&m[1610])|(m[1593]&~m[1594]&m[1595]&m[1596]&m[1610])|(~m[1593]&m[1594]&m[1595]&m[1596]&m[1610]))&~BiasedRNG[872])|((m[1593]&m[1594]&~m[1595]&~m[1596]&~m[1610])|(m[1593]&~m[1594]&m[1595]&~m[1596]&~m[1610])|(~m[1593]&m[1594]&m[1595]&~m[1596]&~m[1610])|(m[1593]&m[1594]&m[1595]&~m[1596]&~m[1610])|(m[1593]&m[1594]&m[1595]&m[1596]&~m[1610])|(m[1593]&m[1594]&~m[1595]&~m[1596]&m[1610])|(m[1593]&~m[1594]&m[1595]&~m[1596]&m[1610])|(~m[1593]&m[1594]&m[1595]&~m[1596]&m[1610])|(m[1593]&m[1594]&m[1595]&~m[1596]&m[1610])|(m[1593]&m[1594]&m[1595]&m[1596]&m[1610]));
    m[1602] = (((m[1598]&~m[1599]&~m[1600]&~m[1601]&~m[1615])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1615])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1615])|(m[1598]&m[1599]&~m[1600]&m[1601]&~m[1615])|(m[1598]&~m[1599]&m[1600]&m[1601]&~m[1615])|(~m[1598]&m[1599]&m[1600]&m[1601]&~m[1615]))&BiasedRNG[873])|(((m[1598]&~m[1599]&~m[1600]&~m[1601]&m[1615])|(~m[1598]&m[1599]&~m[1600]&~m[1601]&m[1615])|(~m[1598]&~m[1599]&m[1600]&~m[1601]&m[1615])|(m[1598]&m[1599]&~m[1600]&m[1601]&m[1615])|(m[1598]&~m[1599]&m[1600]&m[1601]&m[1615])|(~m[1598]&m[1599]&m[1600]&m[1601]&m[1615]))&~BiasedRNG[873])|((m[1598]&m[1599]&~m[1600]&~m[1601]&~m[1615])|(m[1598]&~m[1599]&m[1600]&~m[1601]&~m[1615])|(~m[1598]&m[1599]&m[1600]&~m[1601]&~m[1615])|(m[1598]&m[1599]&m[1600]&~m[1601]&~m[1615])|(m[1598]&m[1599]&m[1600]&m[1601]&~m[1615])|(m[1598]&m[1599]&~m[1600]&~m[1601]&m[1615])|(m[1598]&~m[1599]&m[1600]&~m[1601]&m[1615])|(~m[1598]&m[1599]&m[1600]&~m[1601]&m[1615])|(m[1598]&m[1599]&m[1600]&~m[1601]&m[1615])|(m[1598]&m[1599]&m[1600]&m[1601]&m[1615]));
    m[1607] = (((m[1603]&~m[1604]&~m[1605]&~m[1606]&~m[1620])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1620])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1620])|(m[1603]&m[1604]&~m[1605]&m[1606]&~m[1620])|(m[1603]&~m[1604]&m[1605]&m[1606]&~m[1620])|(~m[1603]&m[1604]&m[1605]&m[1606]&~m[1620]))&BiasedRNG[874])|(((m[1603]&~m[1604]&~m[1605]&~m[1606]&m[1620])|(~m[1603]&m[1604]&~m[1605]&~m[1606]&m[1620])|(~m[1603]&~m[1604]&m[1605]&~m[1606]&m[1620])|(m[1603]&m[1604]&~m[1605]&m[1606]&m[1620])|(m[1603]&~m[1604]&m[1605]&m[1606]&m[1620])|(~m[1603]&m[1604]&m[1605]&m[1606]&m[1620]))&~BiasedRNG[874])|((m[1603]&m[1604]&~m[1605]&~m[1606]&~m[1620])|(m[1603]&~m[1604]&m[1605]&~m[1606]&~m[1620])|(~m[1603]&m[1604]&m[1605]&~m[1606]&~m[1620])|(m[1603]&m[1604]&m[1605]&~m[1606]&~m[1620])|(m[1603]&m[1604]&m[1605]&m[1606]&~m[1620])|(m[1603]&m[1604]&~m[1605]&~m[1606]&m[1620])|(m[1603]&~m[1604]&m[1605]&~m[1606]&m[1620])|(~m[1603]&m[1604]&m[1605]&~m[1606]&m[1620])|(m[1603]&m[1604]&m[1605]&~m[1606]&m[1620])|(m[1603]&m[1604]&m[1605]&m[1606]&m[1620]));
    m[1612] = (((m[1608]&~m[1609]&~m[1610]&~m[1611]&~m[1623])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1623])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1623])|(m[1608]&m[1609]&~m[1610]&m[1611]&~m[1623])|(m[1608]&~m[1609]&m[1610]&m[1611]&~m[1623])|(~m[1608]&m[1609]&m[1610]&m[1611]&~m[1623]))&BiasedRNG[875])|(((m[1608]&~m[1609]&~m[1610]&~m[1611]&m[1623])|(~m[1608]&m[1609]&~m[1610]&~m[1611]&m[1623])|(~m[1608]&~m[1609]&m[1610]&~m[1611]&m[1623])|(m[1608]&m[1609]&~m[1610]&m[1611]&m[1623])|(m[1608]&~m[1609]&m[1610]&m[1611]&m[1623])|(~m[1608]&m[1609]&m[1610]&m[1611]&m[1623]))&~BiasedRNG[875])|((m[1608]&m[1609]&~m[1610]&~m[1611]&~m[1623])|(m[1608]&~m[1609]&m[1610]&~m[1611]&~m[1623])|(~m[1608]&m[1609]&m[1610]&~m[1611]&~m[1623])|(m[1608]&m[1609]&m[1610]&~m[1611]&~m[1623])|(m[1608]&m[1609]&m[1610]&m[1611]&~m[1623])|(m[1608]&m[1609]&~m[1610]&~m[1611]&m[1623])|(m[1608]&~m[1609]&m[1610]&~m[1611]&m[1623])|(~m[1608]&m[1609]&m[1610]&~m[1611]&m[1623])|(m[1608]&m[1609]&m[1610]&~m[1611]&m[1623])|(m[1608]&m[1609]&m[1610]&m[1611]&m[1623]));
    m[1617] = (((m[1613]&~m[1614]&~m[1615]&~m[1616]&~m[1625])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1625])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1625])|(m[1613]&m[1614]&~m[1615]&m[1616]&~m[1625])|(m[1613]&~m[1614]&m[1615]&m[1616]&~m[1625])|(~m[1613]&m[1614]&m[1615]&m[1616]&~m[1625]))&BiasedRNG[876])|(((m[1613]&~m[1614]&~m[1615]&~m[1616]&m[1625])|(~m[1613]&m[1614]&~m[1615]&~m[1616]&m[1625])|(~m[1613]&~m[1614]&m[1615]&~m[1616]&m[1625])|(m[1613]&m[1614]&~m[1615]&m[1616]&m[1625])|(m[1613]&~m[1614]&m[1615]&m[1616]&m[1625])|(~m[1613]&m[1614]&m[1615]&m[1616]&m[1625]))&~BiasedRNG[876])|((m[1613]&m[1614]&~m[1615]&~m[1616]&~m[1625])|(m[1613]&~m[1614]&m[1615]&~m[1616]&~m[1625])|(~m[1613]&m[1614]&m[1615]&~m[1616]&~m[1625])|(m[1613]&m[1614]&m[1615]&~m[1616]&~m[1625])|(m[1613]&m[1614]&m[1615]&m[1616]&~m[1625])|(m[1613]&m[1614]&~m[1615]&~m[1616]&m[1625])|(m[1613]&~m[1614]&m[1615]&~m[1616]&m[1625])|(~m[1613]&m[1614]&m[1615]&~m[1616]&m[1625])|(m[1613]&m[1614]&m[1615]&~m[1616]&m[1625])|(m[1613]&m[1614]&m[1615]&m[1616]&m[1625]));
    m[1622] = (((m[1618]&~m[1619]&~m[1620]&~m[1621]&~m[1630])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1630])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1630])|(m[1618]&m[1619]&~m[1620]&m[1621]&~m[1630])|(m[1618]&~m[1619]&m[1620]&m[1621]&~m[1630])|(~m[1618]&m[1619]&m[1620]&m[1621]&~m[1630]))&BiasedRNG[877])|(((m[1618]&~m[1619]&~m[1620]&~m[1621]&m[1630])|(~m[1618]&m[1619]&~m[1620]&~m[1621]&m[1630])|(~m[1618]&~m[1619]&m[1620]&~m[1621]&m[1630])|(m[1618]&m[1619]&~m[1620]&m[1621]&m[1630])|(m[1618]&~m[1619]&m[1620]&m[1621]&m[1630])|(~m[1618]&m[1619]&m[1620]&m[1621]&m[1630]))&~BiasedRNG[877])|((m[1618]&m[1619]&~m[1620]&~m[1621]&~m[1630])|(m[1618]&~m[1619]&m[1620]&~m[1621]&~m[1630])|(~m[1618]&m[1619]&m[1620]&~m[1621]&~m[1630])|(m[1618]&m[1619]&m[1620]&~m[1621]&~m[1630])|(m[1618]&m[1619]&m[1620]&m[1621]&~m[1630])|(m[1618]&m[1619]&~m[1620]&~m[1621]&m[1630])|(m[1618]&~m[1619]&m[1620]&~m[1621]&m[1630])|(~m[1618]&m[1619]&m[1620]&~m[1621]&m[1630])|(m[1618]&m[1619]&m[1620]&~m[1621]&m[1630])|(m[1618]&m[1619]&m[1620]&m[1621]&m[1630]));
    m[1627] = (((m[1623]&~m[1624]&~m[1625]&~m[1626]&~m[1633])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1633])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1633])|(m[1623]&m[1624]&~m[1625]&m[1626]&~m[1633])|(m[1623]&~m[1624]&m[1625]&m[1626]&~m[1633])|(~m[1623]&m[1624]&m[1625]&m[1626]&~m[1633]))&BiasedRNG[878])|(((m[1623]&~m[1624]&~m[1625]&~m[1626]&m[1633])|(~m[1623]&m[1624]&~m[1625]&~m[1626]&m[1633])|(~m[1623]&~m[1624]&m[1625]&~m[1626]&m[1633])|(m[1623]&m[1624]&~m[1625]&m[1626]&m[1633])|(m[1623]&~m[1624]&m[1625]&m[1626]&m[1633])|(~m[1623]&m[1624]&m[1625]&m[1626]&m[1633]))&~BiasedRNG[878])|((m[1623]&m[1624]&~m[1625]&~m[1626]&~m[1633])|(m[1623]&~m[1624]&m[1625]&~m[1626]&~m[1633])|(~m[1623]&m[1624]&m[1625]&~m[1626]&~m[1633])|(m[1623]&m[1624]&m[1625]&~m[1626]&~m[1633])|(m[1623]&m[1624]&m[1625]&m[1626]&~m[1633])|(m[1623]&m[1624]&~m[1625]&~m[1626]&m[1633])|(m[1623]&~m[1624]&m[1625]&~m[1626]&m[1633])|(~m[1623]&m[1624]&m[1625]&~m[1626]&m[1633])|(m[1623]&m[1624]&m[1625]&~m[1626]&m[1633])|(m[1623]&m[1624]&m[1625]&m[1626]&m[1633]));
    m[1632] = (((m[1628]&~m[1629]&~m[1630]&~m[1631]&~m[1635])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1635])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1635])|(m[1628]&m[1629]&~m[1630]&m[1631]&~m[1635])|(m[1628]&~m[1629]&m[1630]&m[1631]&~m[1635])|(~m[1628]&m[1629]&m[1630]&m[1631]&~m[1635]))&BiasedRNG[879])|(((m[1628]&~m[1629]&~m[1630]&~m[1631]&m[1635])|(~m[1628]&m[1629]&~m[1630]&~m[1631]&m[1635])|(~m[1628]&~m[1629]&m[1630]&~m[1631]&m[1635])|(m[1628]&m[1629]&~m[1630]&m[1631]&m[1635])|(m[1628]&~m[1629]&m[1630]&m[1631]&m[1635])|(~m[1628]&m[1629]&m[1630]&m[1631]&m[1635]))&~BiasedRNG[879])|((m[1628]&m[1629]&~m[1630]&~m[1631]&~m[1635])|(m[1628]&~m[1629]&m[1630]&~m[1631]&~m[1635])|(~m[1628]&m[1629]&m[1630]&~m[1631]&~m[1635])|(m[1628]&m[1629]&m[1630]&~m[1631]&~m[1635])|(m[1628]&m[1629]&m[1630]&m[1631]&~m[1635])|(m[1628]&m[1629]&~m[1630]&~m[1631]&m[1635])|(m[1628]&~m[1629]&m[1630]&~m[1631]&m[1635])|(~m[1628]&m[1629]&m[1630]&~m[1631]&m[1635])|(m[1628]&m[1629]&m[1630]&~m[1631]&m[1635])|(m[1628]&m[1629]&m[1630]&m[1631]&m[1635]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[363]&LFSRcolor0[298]&LFSRcolor0[936]&LFSRcolor0[658]);
    BiasedRNG[1] = (LFSRcolor0[1093]&LFSRcolor0[88]&LFSRcolor0[356]&LFSRcolor0[1238]);
    BiasedRNG[2] = (LFSRcolor0[1148]&LFSRcolor0[1181]&LFSRcolor0[1124]&LFSRcolor0[779]);
    BiasedRNG[3] = (LFSRcolor0[250]&LFSRcolor0[671]&LFSRcolor0[1186]&LFSRcolor0[1138]);
    BiasedRNG[4] = (LFSRcolor0[786]&LFSRcolor0[952]&LFSRcolor0[36]&LFSRcolor0[1139]);
    BiasedRNG[5] = (LFSRcolor0[1231]&LFSRcolor0[752]&LFSRcolor0[252]&LFSRcolor0[1241]);
    BiasedRNG[6] = (LFSRcolor0[555]&LFSRcolor0[83]&LFSRcolor0[736]&LFSRcolor0[552]);
    BiasedRNG[7] = (LFSRcolor0[239]&LFSRcolor0[1218]&LFSRcolor0[243]&LFSRcolor0[1092]);
    BiasedRNG[8] = (LFSRcolor0[1179]&LFSRcolor0[311]&LFSRcolor0[1078]&LFSRcolor0[314]);
    BiasedRNG[9] = (LFSRcolor0[1017]&LFSRcolor0[430]&LFSRcolor0[509]&LFSRcolor0[2]);
    BiasedRNG[10] = (LFSRcolor0[582]&LFSRcolor0[516]&LFSRcolor0[1228]&LFSRcolor0[1065]);
    BiasedRNG[11] = (LFSRcolor0[1192]&LFSRcolor0[107]&LFSRcolor0[875]&LFSRcolor0[829]);
    BiasedRNG[12] = (LFSRcolor0[256]&LFSRcolor0[847]&LFSRcolor0[484]&LFSRcolor0[1006]);
    BiasedRNG[13] = (LFSRcolor0[319]&LFSRcolor0[905]&LFSRcolor0[370]&LFSRcolor0[260]);
    BiasedRNG[14] = (LFSRcolor0[290]&LFSRcolor0[755]&LFSRcolor0[104]&LFSRcolor0[638]);
    BiasedRNG[15] = (LFSRcolor0[605]&LFSRcolor0[1167]&LFSRcolor0[1100]&LFSRcolor0[1025]);
    BiasedRNG[16] = (LFSRcolor0[659]&LFSRcolor0[1088]&LFSRcolor0[482]&LFSRcolor0[58]);
    BiasedRNG[17] = (LFSRcolor0[954]&LFSRcolor0[322]&LFSRcolor0[425]&LFSRcolor0[420]);
    BiasedRNG[18] = (LFSRcolor0[1170]&LFSRcolor0[1068]&LFSRcolor0[1205]&LFSRcolor0[297]);
    BiasedRNG[19] = (LFSRcolor0[728]&LFSRcolor0[277]&LFSRcolor0[825]&LFSRcolor0[1197]);
    BiasedRNG[20] = (LFSRcolor0[567]&LFSRcolor0[75]&LFSRcolor0[139]&LFSRcolor0[496]);
    BiasedRNG[21] = (LFSRcolor0[108]&LFSRcolor0[1109]&LFSRcolor0[553]&LFSRcolor0[1115]);
    BiasedRNG[22] = (LFSRcolor0[70]&LFSRcolor0[933]&LFSRcolor0[398]&LFSRcolor0[307]);
    BiasedRNG[23] = (LFSRcolor0[473]&LFSRcolor0[368]&LFSRcolor0[569]&LFSRcolor0[554]);
    BiasedRNG[24] = (LFSRcolor0[153]&LFSRcolor0[741]&LFSRcolor0[455]&LFSRcolor0[523]);
    BiasedRNG[25] = (LFSRcolor0[561]&LFSRcolor0[1145]&LFSRcolor0[393]&LFSRcolor0[427]);
    BiasedRNG[26] = (LFSRcolor0[633]&LFSRcolor0[456]&LFSRcolor0[1097]&LFSRcolor0[38]);
    BiasedRNG[27] = (LFSRcolor0[1158]&LFSRcolor0[1057]&LFSRcolor0[498]&LFSRcolor0[780]);
    BiasedRNG[28] = (LFSRcolor0[914]&LFSRcolor0[709]&LFSRcolor0[890]&LFSRcolor0[406]);
    BiasedRNG[29] = (LFSRcolor0[62]&LFSRcolor0[255]&LFSRcolor0[1028]&LFSRcolor0[804]);
    BiasedRNG[30] = (LFSRcolor0[179]&LFSRcolor0[1004]&LFSRcolor0[388]&LFSRcolor0[852]);
    BiasedRNG[31] = (LFSRcolor0[1162]&LFSRcolor0[968]&LFSRcolor0[1011]&LFSRcolor0[1103]);
    BiasedRNG[32] = (LFSRcolor0[771]&LFSRcolor0[846]&LFSRcolor0[807]&LFSRcolor0[904]);
    BiasedRNG[33] = (LFSRcolor0[941]&LFSRcolor0[327]&LFSRcolor0[114]&LFSRcolor0[886]);
    BiasedRNG[34] = (LFSRcolor0[992]&LFSRcolor0[703]&LFSRcolor0[5]&LFSRcolor0[787]);
    BiasedRNG[35] = (LFSRcolor0[160]&LFSRcolor0[1082]&LFSRcolor0[810]&LFSRcolor0[879]);
    BiasedRNG[36] = (LFSRcolor0[1049]&LFSRcolor0[9]&LFSRcolor0[1074]&LFSRcolor0[365]);
    BiasedRNG[37] = (LFSRcolor0[1116]&LFSRcolor0[740]&LFSRcolor0[585]&LFSRcolor0[720]);
    BiasedRNG[38] = (LFSRcolor0[1120]&LFSRcolor0[73]&LFSRcolor0[537]&LFSRcolor0[293]);
    BiasedRNG[39] = (LFSRcolor0[340]&LFSRcolor0[919]&LFSRcolor0[188]&LFSRcolor0[839]);
    BiasedRNG[40] = (LFSRcolor0[1154]&LFSRcolor0[405]&LFSRcolor0[991]&LFSRcolor0[283]);
    BiasedRNG[41] = (LFSRcolor0[102]&LFSRcolor0[799]&LFSRcolor0[421]&LFSRcolor0[538]);
    BiasedRNG[42] = (LFSRcolor0[1083]&LFSRcolor0[1053]&LFSRcolor0[15]&LFSRcolor0[274]);
    BiasedRNG[43] = (LFSRcolor0[940]&LFSRcolor0[1194]&LFSRcolor0[996]&LFSRcolor0[956]);
    BiasedRNG[44] = (LFSRcolor0[19]&LFSRcolor0[560]&LFSRcolor0[828]&LFSRcolor0[920]);
    BiasedRNG[45] = (LFSRcolor0[611]&LFSRcolor0[749]&LFSRcolor0[1079]&LFSRcolor0[201]);
    BiasedRNG[46] = (LFSRcolor0[445]&LFSRcolor0[573]&LFSRcolor0[602]&LFSRcolor0[359]);
    BiasedRNG[47] = (LFSRcolor0[483]&LFSRcolor0[721]&LFSRcolor0[1224]&LFSRcolor0[614]);
    BiasedRNG[48] = (LFSRcolor0[105]&LFSRcolor0[299]&LFSRcolor0[598]&LFSRcolor0[254]);
    BiasedRNG[49] = (LFSRcolor0[40]&LFSRcolor0[262]&LFSRcolor0[1214]&LFSRcolor0[637]);
    BiasedRNG[50] = (LFSRcolor0[630]&LFSRcolor0[942]&LFSRcolor0[883]&LFSRcolor0[873]);
    BiasedRNG[51] = (LFSRcolor0[120]&LFSRcolor0[690]&LFSRcolor0[216]&LFSRcolor0[46]);
    BiasedRNG[52] = (LFSRcolor0[1202]&LFSRcolor0[699]&LFSRcolor0[305]&LFSRcolor0[1012]);
    BiasedRNG[53] = (LFSRcolor0[915]&LFSRcolor0[203]&LFSRcolor0[337]&LFSRcolor0[115]);
    BiasedRNG[54] = (LFSRcolor0[384]&LFSRcolor0[676]&LFSRcolor0[619]&LFSRcolor0[589]);
    BiasedRNG[55] = (LFSRcolor0[148]&LFSRcolor0[1211]&LFSRcolor0[494]&LFSRcolor0[970]);
    BiasedRNG[56] = (LFSRcolor0[836]&LFSRcolor0[449]&LFSRcolor0[411]&LFSRcolor0[190]);
    BiasedRNG[57] = (LFSRcolor0[651]&LFSRcolor0[231]&LFSRcolor0[833]&LFSRcolor0[387]);
    BiasedRNG[58] = (LFSRcolor0[784]&LFSRcolor0[600]&LFSRcolor0[60]&LFSRcolor0[127]);
    BiasedRNG[59] = (LFSRcolor0[535]&LFSRcolor0[1042]&LFSRcolor0[581]&LFSRcolor0[524]);
    BiasedRNG[60] = (LFSRcolor0[1]&LFSRcolor0[907]&LFSRcolor0[1140]&LFSRcolor0[1182]);
    BiasedRNG[61] = (LFSRcolor0[512]&LFSRcolor0[962]&LFSRcolor0[367]&LFSRcolor0[1062]);
    BiasedRNG[62] = (LFSRcolor0[301]&LFSRcolor0[6]&LFSRcolor0[325]&LFSRcolor0[1066]);
    BiasedRNG[63] = (LFSRcolor0[410]&LFSRcolor0[574]&LFSRcolor0[69]&LFSRcolor0[528]);
    BiasedRNG[64] = (LFSRcolor0[1052]&LFSRcolor0[1204]&LFSRcolor0[1054]&LFSRcolor0[385]);
    BiasedRNG[65] = (LFSRcolor0[767]&LFSRcolor0[680]&LFSRcolor0[916]&LFSRcolor0[931]);
    BiasedRNG[66] = (LFSRcolor0[897]&LFSRcolor0[296]&LFSRcolor0[966]&LFSRcolor0[1173]);
    BiasedRNG[67] = (LFSRcolor0[362]&LFSRcolor0[544]&LFSRcolor0[475]&LFSRcolor0[1047]);
    BiasedRNG[68] = (LFSRcolor0[1221]&LFSRcolor0[171]&LFSRcolor0[90]&LFSRcolor0[241]);
    BiasedRNG[69] = (LFSRcolor0[55]&LFSRcolor0[577]&LFSRcolor0[742]&LFSRcolor0[267]);
    BiasedRNG[70] = (LFSRcolor0[714]&LFSRcolor0[71]&LFSRcolor0[1075]&LFSRcolor0[811]);
    BiasedRNG[71] = (LFSRcolor0[1022]&LFSRcolor0[1178]&LFSRcolor0[1149]&LFSRcolor0[923]);
    BiasedRNG[72] = (LFSRcolor0[51]&LFSRcolor0[717]&LFSRcolor0[335]&LFSRcolor0[200]);
    BiasedRNG[73] = (LFSRcolor0[838]&LFSRcolor0[565]&LFSRcolor0[608]&LFSRcolor0[1152]);
    BiasedRNG[74] = (LFSRcolor0[280]&LFSRcolor0[677]&LFSRcolor0[353]&LFSRcolor0[437]);
    BiasedRNG[75] = (LFSRcolor0[782]&LFSRcolor0[949]&LFSRcolor0[1073]&LFSRcolor0[30]);
    BiasedRNG[76] = (LFSRcolor0[612]&LFSRcolor0[622]&LFSRcolor0[237]&LFSRcolor0[818]);
    BiasedRNG[77] = (LFSRcolor0[716]&LFSRcolor0[497]&LFSRcolor0[236]&LFSRcolor0[912]);
    BiasedRNG[78] = (LFSRcolor0[711]&LFSRcolor0[350]&LFSRcolor0[1037]&LFSRcolor0[1039]);
    BiasedRNG[79] = (LFSRcolor0[447]&LFSRcolor0[14]&LFSRcolor0[673]&LFSRcolor0[1201]);
    BiasedRNG[80] = (LFSRcolor0[1196]&LFSRcolor0[621]&LFSRcolor0[1085]&LFSRcolor0[814]);
    BiasedRNG[81] = (LFSRcolor0[24]&LFSRcolor0[464]&LFSRcolor0[840]&LFSRcolor0[226]);
    BiasedRNG[82] = (LFSRcolor0[750]&LFSRcolor0[681]&LFSRcolor0[294]&LFSRcolor0[450]);
    BiasedRNG[83] = (LFSRcolor0[719]&LFSRcolor0[881]&LFSRcolor0[1005]&LFSRcolor0[998]);
    BiasedRNG[84] = (LFSRcolor0[76]&LFSRcolor0[1029]&LFSRcolor0[366]&LFSRcolor0[877]);
    BiasedRNG[85] = (LFSRcolor0[1081]&LFSRcolor0[1018]&LFSRcolor0[901]&LFSRcolor0[331]);
    BiasedRNG[86] = (LFSRcolor0[479]&LFSRcolor0[287]&LFSRcolor0[234]&LFSRcolor0[391]);
    BiasedRNG[87] = (LFSRcolor0[110]&LFSRcolor0[380]&LFSRcolor0[689]&LFSRcolor0[888]);
    BiasedRNG[88] = (LFSRcolor0[371]&LFSRcolor0[729]&LFSRcolor0[109]&LFSRcolor0[31]);
    BiasedRNG[89] = (LFSRcolor0[540]&LFSRcolor0[369]&LFSRcolor0[209]&LFSRcolor0[1234]);
    BiasedRNG[90] = (LFSRcolor0[1077]&LFSRcolor0[909]&LFSRcolor0[1142]&LFSRcolor0[1106]);
    BiasedRNG[91] = (LFSRcolor0[522]&LFSRcolor0[328]&LFSRcolor0[557]&LFSRcolor0[98]);
    BiasedRNG[92] = (LFSRcolor0[609]&LFSRcolor0[126]&LFSRcolor0[155]&LFSRcolor0[64]);
    BiasedRNG[93] = (LFSRcolor0[1209]&LFSRcolor0[871]&LFSRcolor0[636]&LFSRcolor0[656]);
    BiasedRNG[94] = (LFSRcolor0[32]&LFSRcolor0[352]&LFSRcolor0[49]&LFSRcolor0[422]);
    BiasedRNG[95] = (LFSRcolor0[419]&LFSRcolor0[520]&LFSRcolor0[1183]&LFSRcolor0[18]);
    BiasedRNG[96] = (LFSRcolor0[310]&LFSRcolor0[63]&LFSRcolor0[649]&LFSRcolor0[1208]);
    BiasedRNG[97] = (LFSRcolor0[228]&LFSRcolor0[543]&LFSRcolor0[896]&LFSRcolor0[809]);
    BiasedRNG[98] = (LFSRcolor0[669]&LFSRcolor0[590]&LFSRcolor0[986]&LFSRcolor0[1177]);
    BiasedRNG[99] = (LFSRcolor0[383]&LFSRcolor0[858]&LFSRcolor0[791]&LFSRcolor0[308]);
    BiasedRNG[100] = (LFSRcolor0[639]&LFSRcolor0[329]&LFSRcolor0[181]&LFSRcolor0[400]);
    BiasedRNG[101] = (LFSRcolor0[263]&LFSRcolor0[128]&LFSRcolor0[972]&LFSRcolor0[929]);
    BiasedRNG[102] = (LFSRcolor0[1021]&LFSRcolor0[1061]&LFSRcolor0[951]&LFSRcolor0[541]);
    BiasedRNG[103] = (LFSRcolor0[477]&LFSRcolor0[1090]&LFSRcolor0[627]&LFSRcolor0[358]);
    BiasedRNG[104] = (LFSRcolor0[817]&LFSRcolor0[648]&LFSRcolor0[618]&LFSRcolor0[513]);
    BiasedRNG[105] = (LFSRcolor0[733]&LFSRcolor0[978]&LFSRcolor0[660]&LFSRcolor0[924]);
    BiasedRNG[106] = (LFSRcolor0[158]&LFSRcolor0[195]&LFSRcolor0[253]&LFSRcolor0[932]);
    BiasedRNG[107] = (LFSRcolor0[969]&LFSRcolor0[654]&LFSRcolor0[603]&LFSRcolor0[424]);
    BiasedRNG[108] = (LFSRcolor0[382]&LFSRcolor0[1095]&LFSRcolor0[693]&LFSRcolor0[684]);
    BiasedRNG[109] = (LFSRcolor0[1003]&LFSRcolor0[150]&LFSRcolor0[152]&LFSRcolor0[610]);
    BiasedRNG[110] = (LFSRcolor0[270]&LFSRcolor0[316]&LFSRcolor0[822]&LFSRcolor0[312]);
    BiasedRNG[111] = (LFSRcolor0[59]&LFSRcolor0[562]&LFSRcolor0[657]&LFSRcolor0[413]);
    BiasedRNG[112] = (LFSRcolor0[26]&LFSRcolor0[103]&LFSRcolor0[180]&LFSRcolor0[173]);
    BiasedRNG[113] = (LFSRcolor0[94]&LFSRcolor0[855]&LFSRcolor0[223]&LFSRcolor0[1096]);
    BiasedRNG[114] = (LFSRcolor0[506]&LFSRcolor0[922]&LFSRcolor0[157]&LFSRcolor0[136]);
    BiasedRNG[115] = (LFSRcolor0[416]&LFSRcolor0[798]&LFSRcolor0[42]&LFSRcolor0[860]);
    BiasedRNG[116] = (LFSRcolor0[159]&LFSRcolor0[392]&LFSRcolor0[950]&LFSRcolor0[1195]);
    BiasedRNG[117] = (LFSRcolor0[439]&LFSRcolor0[662]&LFSRcolor0[485]&LFSRcolor0[230]);
    BiasedRNG[118] = (LFSRcolor0[1185]&LFSRcolor0[959]&LFSRcolor0[975]&LFSRcolor0[377]);
    BiasedRNG[119] = (LFSRcolor0[1180]&LFSRcolor0[961]&LFSRcolor0[233]&LFSRcolor0[1153]);
    BiasedRNG[120] = (LFSRcolor0[1189]&LFSRcolor0[1001]&LFSRcolor0[318]&LFSRcolor0[935]);
    BiasedRNG[121] = (LFSRcolor0[1110]&LFSRcolor0[644]&LFSRcolor0[759]&LFSRcolor0[534]);
    BiasedRNG[122] = (LFSRcolor0[1024]&LFSRcolor0[227]&LFSRcolor0[1122]&LFSRcolor0[596]);
    BiasedRNG[123] = (LFSRcolor0[606]&LFSRcolor0[185]&LFSRcolor0[501]&LFSRcolor0[696]);
    BiasedRNG[124] = (LFSRcolor0[960]&LFSRcolor0[550]&LFSRcolor0[511]&LFSRcolor0[221]);
    BiasedRNG[125] = (LFSRcolor0[588]&LFSRcolor0[232]&LFSRcolor0[313]&LFSRcolor0[191]);
    BiasedRNG[126] = (LFSRcolor0[859]&LFSRcolor0[792]&LFSRcolor0[121]&LFSRcolor0[462]);
    BiasedRNG[127] = (LFSRcolor0[1020]&LFSRcolor0[624]&LFSRcolor0[379]&LFSRcolor0[184]);
    BiasedRNG[128] = (LFSRcolor0[1107]&LFSRcolor0[1150]&LFSRcolor0[438]&LFSRcolor0[112]);
    BiasedRNG[129] = (LFSRcolor0[142]&LFSRcolor0[404]&LFSRcolor0[172]&LFSRcolor0[35]);
    BiasedRNG[130] = (LFSRcolor0[551]&LFSRcolor0[1098]&LFSRcolor0[1227]&LFSRcolor0[176]);
    BiasedRNG[131] = (LFSRcolor0[646]&LFSRcolor0[687]&LFSRcolor0[701]&LFSRcolor0[495]);
    BiasedRNG[132] = (LFSRcolor0[134]&LFSRcolor0[911]&LFSRcolor0[758]&LFSRcolor0[1127]);
    BiasedRNG[133] = (LFSRcolor0[343]&LFSRcolor0[917]&LFSRcolor0[1069]&LFSRcolor0[169]);
    BiasedRNG[134] = (LFSRcolor0[682]&LFSRcolor0[1118]&LFSRcolor0[212]&LFSRcolor0[830]);
    BiasedRNG[135] = (LFSRcolor0[880]&LFSRcolor0[481]&LFSRcolor0[154]&LFSRcolor0[202]);
    BiasedRNG[136] = (LFSRcolor0[955]&LFSRcolor0[1147]&LFSRcolor0[113]&LFSRcolor0[685]);
    BiasedRNG[137] = (LFSRcolor0[198]&LFSRcolor0[514]&LFSRcolor0[468]&LFSRcolor0[900]);
    BiasedRNG[138] = (LFSRcolor0[238]&LFSRcolor0[478]&LFSRcolor0[751]&LFSRcolor0[499]);
    BiasedRNG[139] = (LFSRcolor0[1113]&LFSRcolor0[1191]&LFSRcolor0[351]&LFSRcolor0[339]);
    BiasedRNG[140] = (LFSRcolor0[793]&LFSRcolor0[1156]&LFSRcolor0[774]&LFSRcolor0[765]);
    BiasedRNG[141] = (LFSRcolor0[217]&LFSRcolor0[208]&LFSRcolor0[640]&LFSRcolor0[597]);
    BiasedRNG[142] = (LFSRcolor0[225]&LFSRcolor0[579]&LFSRcolor0[632]&LFSRcolor0[889]);
    BiasedRNG[143] = (LFSRcolor0[937]&LFSRcolor0[620]&LFSRcolor0[219]&LFSRcolor0[373]);
    BiasedRNG[144] = (LFSRcolor0[162]&LFSRcolor0[66]&LFSRcolor0[835]&LFSRcolor0[1215]);
    BiasedRNG[145] = (LFSRcolor0[725]&LFSRcolor0[876]&LFSRcolor0[1161]&LFSRcolor0[207]);
    BiasedRNG[146] = (LFSRcolor0[634]&LFSRcolor0[1217]&LFSRcolor0[796]&LFSRcolor0[823]);
    BiasedRNG[147] = (LFSRcolor0[347]&LFSRcolor0[264]&LFSRcolor0[434]&LFSRcolor0[1033]);
    BiasedRNG[148] = (LFSRcolor0[278]&LFSRcolor0[276]&LFSRcolor0[702]&LFSRcolor0[458]);
    BiasedRNG[149] = (LFSRcolor0[1203]&LFSRcolor0[125]&LFSRcolor0[317]&LFSRcolor0[451]);
    BiasedRNG[150] = (LFSRcolor0[586]&LFSRcolor0[525]&LFSRcolor0[1131]&LFSRcolor0[500]);
    BiasedRNG[151] = (LFSRcolor0[472]&LFSRcolor0[240]&LFSRcolor0[164]&LFSRcolor0[707]);
    BiasedRNG[152] = (LFSRcolor0[53]&LFSRcolor0[133]&LFSRcolor0[23]&LFSRcolor0[1134]);
    BiasedRNG[153] = (LFSRcolor0[993]&LFSRcolor0[1094]&LFSRcolor0[724]&LFSRcolor0[539]);
    BiasedRNG[154] = (LFSRcolor0[1126]&LFSRcolor0[258]&LFSRcolor0[1200]&LFSRcolor0[1121]);
    BiasedRNG[155] = (LFSRcolor0[86]&LFSRcolor0[893]&LFSRcolor0[376]&LFSRcolor0[739]);
    BiasedRNG[156] = (LFSRcolor0[747]&LFSRcolor0[1143]&LFSRcolor0[426]&LFSRcolor0[613]);
    BiasedRNG[157] = (LFSRcolor0[926]&LFSRcolor0[938]&LFSRcolor0[891]&LFSRcolor0[519]);
    BiasedRNG[158] = (LFSRcolor0[849]&LFSRcolor0[504]&LFSRcolor0[894]&LFSRcolor0[570]);
    BiasedRNG[159] = (LFSRcolor0[781]&LFSRcolor0[229]&LFSRcolor0[939]&LFSRcolor0[402]);
    BiasedRNG[160] = (LFSRcolor0[546]&LFSRcolor0[291]&LFSRcolor0[403]&LFSRcolor0[138]);
    BiasedRNG[161] = (LFSRcolor0[1163]&LFSRcolor0[1036]&LFSRcolor0[443]&LFSRcolor0[448]);
    BiasedRNG[162] = (LFSRcolor0[27]&LFSRcolor0[333]&LFSRcolor0[33]&LFSRcolor0[1104]);
    BiasedRNG[163] = (LFSRcolor0[770]&LFSRcolor0[418]&LFSRcolor0[41]&LFSRcolor0[442]);
    BiasedRNG[164] = (LFSRcolor0[145]&LFSRcolor0[204]&LFSRcolor0[1045]&LFSRcolor0[688]);
    BiasedRNG[165] = (LFSRcolor0[166]&LFSRcolor0[50]&LFSRcolor0[865]&LFSRcolor0[987]);
    BiasedRNG[166] = (LFSRcolor0[979]&LFSRcolor0[783]&LFSRcolor0[321]&LFSRcolor0[132]);
    BiasedRNG[167] = (LFSRcolor0[446]&LFSRcolor0[211]&LFSRcolor0[22]&LFSRcolor0[872]);
    BiasedRNG[168] = (LFSRcolor0[776]&LFSRcolor0[1240]&LFSRcolor0[206]&LFSRcolor0[271]);
    BiasedRNG[169] = (LFSRcolor0[1133]&LFSRcolor0[1184]&LFSRcolor0[1051]&LFSRcolor0[1019]);
    BiasedRNG[170] = (LFSRcolor0[819]&LFSRcolor0[921]&LFSRcolor0[576]&LFSRcolor0[1026]);
    BiasedRNG[171] = (LFSRcolor0[186]&LFSRcolor0[99]&LFSRcolor0[934]&LFSRcolor0[338]);
    BiasedRNG[172] = (LFSRcolor0[1239]&LFSRcolor0[1060]&LFSRcolor0[74]&LFSRcolor0[163]);
    BiasedRNG[173] = (LFSRcolor0[1114]&LFSRcolor0[718]&LFSRcolor0[801]&LFSRcolor0[397]);
    BiasedRNG[174] = (LFSRcolor0[726]&LFSRcolor0[559]&LFSRcolor0[899]&LFSRcolor0[183]);
    BiasedRNG[175] = (LFSRcolor0[655]&LFSRcolor0[853]&LFSRcolor0[1174]&LFSRcolor0[16]);
    BiasedRNG[176] = (LFSRcolor0[678]&LFSRcolor0[295]&LFSRcolor0[547]&LFSRcolor0[1015]);
    BiasedRNG[177] = (LFSRcolor0[344]&LFSRcolor0[389]&LFSRcolor0[268]&LFSRcolor0[1207]);
    BiasedRNG[178] = (LFSRcolor0[25]&LFSRcolor0[686]&LFSRcolor0[1035]&LFSRcolor0[587]);
    BiasedRNG[179] = (LFSRcolor0[526]&LFSRcolor0[1137]&LFSRcolor0[831]&LFSRcolor0[762]);
    BiasedRNG[180] = (LFSRcolor0[1089]&LFSRcolor0[769]&LFSRcolor0[408]&LFSRcolor0[43]);
    BiasedRNG[181] = (LFSRcolor0[775]&LFSRcolor0[471]&LFSRcolor0[1151]&LFSRcolor0[244]);
    BiasedRNG[182] = (LFSRcolor0[77]&LFSRcolor0[1190]&LFSRcolor0[592]&LFSRcolor0[628]);
    BiasedRNG[183] = (LFSRcolor0[815]&LFSRcolor0[575]&LFSRcolor0[1187]&LFSRcolor0[275]);
    BiasedRNG[184] = (LFSRcolor0[44]&LFSRcolor0[1169]&LFSRcolor0[187]&LFSRcolor0[753]);
    BiasedRNG[185] = (LFSRcolor0[510]&LFSRcolor0[558]&LFSRcolor0[863]&LFSRcolor0[963]);
    BiasedRNG[186] = (LFSRcolor0[861]&LFSRcolor0[257]&LFSRcolor0[245]&LFSRcolor0[583]);
    BiasedRNG[187] = (LFSRcolor0[1076]&LFSRcolor0[1188]&LFSRcolor0[816]&LFSRcolor0[1159]);
    BiasedRNG[188] = (LFSRcolor0[466]&LFSRcolor0[884]&LFSRcolor0[144]&LFSRcolor0[39]);
    BiasedRNG[189] = (LFSRcolor0[668]&LFSRcolor0[214]&LFSRcolor0[415]&LFSRcolor0[556]);
    BiasedRNG[190] = (LFSRcolor0[625]&LFSRcolor0[1119]&LFSRcolor0[93]&LFSRcolor0[3]);
    BiasedRNG[191] = (LFSRcolor0[867]&LFSRcolor0[84]&LFSRcolor0[10]&LFSRcolor0[265]);
    BiasedRNG[192] = (LFSRcolor0[976]&LFSRcolor0[820]&LFSRcolor0[731]&LFSRcolor0[870]);
    BiasedRNG[193] = (LFSRcolor0[119]&LFSRcolor0[13]&LFSRcolor0[1056]&LFSRcolor0[210]);
    BiasedRNG[194] = (LFSRcolor0[763]&LFSRcolor0[354]&LFSRcolor0[545]&LFSRcolor0[251]);
    BiasedRNG[195] = (LFSRcolor0[386]&LFSRcolor0[222]&LFSRcolor0[248]&LFSRcolor0[571]);
    BiasedRNG[196] = (LFSRcolor0[1144]&LFSRcolor0[1070]&LFSRcolor0[985]&LFSRcolor0[533]);
    BiasedRNG[197] = (LFSRcolor0[679]&LFSRcolor0[947]&LFSRcolor0[432]&LFSRcolor0[381]);
    BiasedRNG[198] = (LFSRcolor0[281]&LFSRcolor0[697]&LFSRcolor0[177]&LFSRcolor0[396]);
    BiasedRNG[199] = (LFSRcolor0[97]&LFSRcolor0[977]&LFSRcolor0[61]&LFSRcolor0[452]);
    BiasedRNG[200] = (LFSRcolor0[518]&LFSRcolor0[665]&LFSRcolor0[360]&LFSRcolor0[111]);
    BiasedRNG[201] = (LFSRcolor0[663]&LFSRcolor0[11]&LFSRcolor0[37]&LFSRcolor0[832]);
    BiasedRNG[202] = (LFSRcolor0[436]&LFSRcolor0[1027]&LFSRcolor0[96]&LFSRcolor0[1123]);
    BiasedRNG[203] = (LFSRcolor0[56]&LFSRcolor0[745]&LFSRcolor0[507]&LFSRcolor0[395]);
    BiasedRNG[204] = (LFSRcolor0[953]&LFSRcolor0[635]&LFSRcolor0[995]&LFSRcolor0[994]);
    BiasedRNG[205] = (LFSRcolor0[910]&LFSRcolor0[666]&LFSRcolor0[1091]&LFSRcolor0[300]);
    BiasedRNG[206] = (LFSRcolor0[643]&LFSRcolor0[944]&LFSRcolor0[957]&LFSRcolor0[790]);
    BiasedRNG[207] = (LFSRcolor0[515]&LFSRcolor0[945]&LFSRcolor0[282]&LFSRcolor0[151]);
    BiasedRNG[208] = (LFSRcolor0[641]&LFSRcolor0[694]&LFSRcolor0[118]&LFSRcolor0[269]);
    BiasedRNG[209] = (LFSRcolor0[593]&LFSRcolor0[542]&LFSRcolor0[675]&LFSRcolor0[1125]);
    BiasedRNG[210] = (LFSRcolor0[892]&LFSRcolor0[981]&LFSRcolor0[664]&LFSRcolor0[626]);
    BiasedRNG[211] = (LFSRcolor0[869]&LFSRcolor0[326]&LFSRcolor0[286]&LFSRcolor0[259]);
    BiasedRNG[212] = (LFSRcolor0[469]&LFSRcolor0[652]&LFSRcolor0[984]&LFSRcolor0[47]);
    BiasedRNG[213] = (LFSRcolor0[761]&LFSRcolor0[722]&LFSRcolor0[401]&LFSRcolor0[617]);
    BiasedRNG[214] = (LFSRcolor0[723]&LFSRcolor0[1160]&LFSRcolor0[399]&LFSRcolor0[12]);
    BiasedRNG[215] = (LFSRcolor0[1084]&LFSRcolor0[895]&LFSRcolor0[1031]&LFSRcolor0[1132]);
    BiasedRNG[216] = (LFSRcolor0[1155]&LFSRcolor0[1130]&LFSRcolor0[82]&LFSRcolor0[444]);
    BiasedRNG[217] = (LFSRcolor0[304]&LFSRcolor0[130]&LFSRcolor0[140]&LFSRcolor0[744]);
    BiasedRNG[218] = (LFSRcolor0[599]&LFSRcolor0[460]&LFSRcolor0[357]&LFSRcolor0[149]);
    BiasedRNG[219] = (LFSRcolor0[997]&LFSRcolor0[490]&LFSRcolor0[943]&LFSRcolor0[530]);
    BiasedRNG[220] = (LFSRcolor0[194]&LFSRcolor0[8]&LFSRcolor0[868]&LFSRcolor0[302]);
    BiasedRNG[221] = (LFSRcolor0[616]&LFSRcolor0[330]&LFSRcolor0[715]&LFSRcolor0[824]);
    BiasedRNG[222] = (LFSRcolor0[488]&LFSRcolor0[1199]&LFSRcolor0[568]&LFSRcolor0[1059]);
    BiasedRNG[223] = (LFSRcolor0[1168]&LFSRcolor0[7]&LFSRcolor0[748]&LFSRcolor0[925]);
    BiasedRNG[224] = (LFSRcolor0[727]&LFSRcolor0[197]&LFSRcolor0[52]&LFSRcolor0[135]);
    BiasedRNG[225] = (LFSRcolor0[843]&LFSRcolor0[795]&LFSRcolor0[372]&LFSRcolor0[361]);
    BiasedRNG[226] = (LFSRcolor0[1229]&LFSRcolor0[320]&LFSRcolor0[242]&LFSRcolor0[1112]);
    BiasedRNG[227] = (LFSRcolor0[266]&LFSRcolor0[493]&LFSRcolor0[487]&LFSRcolor0[887]);
    BiasedRNG[228] = (LFSRcolor0[117]&LFSRcolor0[80]&LFSRcolor0[1016]&LFSRcolor0[465]);
    BiasedRNG[229] = (LFSRcolor0[1030]&LFSRcolor0[958]&LFSRcolor0[1172]&LFSRcolor0[182]);
    BiasedRNG[230] = (LFSRcolor0[1193]&LFSRcolor0[178]&LFSRcolor0[980]&LFSRcolor0[454]);
    BiasedRNG[231] = (LFSRcolor0[989]&LFSRcolor0[218]&LFSRcolor0[670]&LFSRcolor0[854]);
    BiasedRNG[232] = (LFSRcolor0[348]&LFSRcolor0[1040]&LFSRcolor0[1063]&LFSRcolor0[650]);
    BiasedRNG[233] = (LFSRcolor0[1222]&LFSRcolor0[168]&LFSRcolor0[549]&LFSRcolor0[193]);
    BiasedRNG[234] = (LFSRcolor0[414]&LFSRcolor0[973]&LFSRcolor0[374]&LFSRcolor0[913]);
    BiasedRNG[235] = (LFSRcolor0[1038]&LFSRcolor0[355]&LFSRcolor0[131]&LFSRcolor0[834]);
    BiasedRNG[236] = (LFSRcolor0[967]&LFSRcolor0[502]&LFSRcolor0[143]&LFSRcolor0[808]);
    BiasedRNG[237] = (LFSRcolor0[1223]&LFSRcolor0[441]&LFSRcolor0[428]&LFSRcolor0[595]);
    BiasedRNG[238] = (LFSRcolor0[491]&LFSRcolor0[521]&LFSRcolor0[453]&LFSRcolor0[1050]);
    BiasedRNG[239] = (LFSRcolor0[1232]&LFSRcolor0[457]&LFSRcolor0[766]&LFSRcolor0[850]);
    BiasedRNG[240] = (LFSRcolor0[578]&LFSRcolor0[346]&LFSRcolor0[72]&LFSRcolor0[1233]);
    BiasedRNG[241] = (LFSRcolor0[764]&LFSRcolor0[584]&LFSRcolor0[1226]&LFSRcolor0[756]);
    BiasedRNG[242] = (LFSRcolor0[273]&LFSRcolor0[803]&LFSRcolor0[288]&LFSRcolor0[235]);
    BiasedRNG[243] = (LFSRcolor0[1225]&LFSRcolor0[4]&LFSRcolor0[101]&LFSRcolor0[440]);
    BiasedRNG[244] = (LFSRcolor0[738]&LFSRcolor0[812]&LFSRcolor0[862]&LFSRcolor0[563]);
    BiasedRNG[245] = (LFSRcolor0[390]&LFSRcolor0[754]&LFSRcolor0[45]&LFSRcolor0[1080]);
    BiasedRNG[246] = (LFSRcolor0[566]&LFSRcolor0[137]&LFSRcolor0[1010]&LFSRcolor0[805]);
    BiasedRNG[247] = (LFSRcolor0[1171]&LFSRcolor0[517]&LFSRcolor0[730]&LFSRcolor0[303]);
    BiasedRNG[248] = (LFSRcolor0[292]&LFSRcolor0[1013]&LFSRcolor0[735]&LFSRcolor0[48]);
    BiasedRNG[249] = (LFSRcolor0[167]&LFSRcolor0[844]&LFSRcolor0[1212]&LFSRcolor0[189]);
    BiasedRNG[250] = (LFSRcolor0[990]&LFSRcolor0[480]&LFSRcolor0[1014]&LFSRcolor0[34]);
    BiasedRNG[251] = (LFSRcolor0[334]&LFSRcolor0[285]&LFSRcolor0[661]&LFSRcolor0[192]);
    UnbiasedRNG[0] = LFSRcolor0[423];
    UnbiasedRNG[1] = LFSRcolor0[20];
    UnbiasedRNG[2] = LFSRcolor0[246];
    UnbiasedRNG[3] = LFSRcolor0[746];
    UnbiasedRNG[4] = LFSRcolor0[505];
    UnbiasedRNG[5] = LFSRcolor0[706];
    UnbiasedRNG[6] = LFSRcolor0[813];
    UnbiasedRNG[7] = LFSRcolor0[1041];
    UnbiasedRNG[8] = LFSRcolor0[122];
    UnbiasedRNG[9] = LFSRcolor0[906];
    UnbiasedRNG[10] = LFSRcolor0[531];
    UnbiasedRNG[11] = LFSRcolor0[508];
    UnbiasedRNG[12] = LFSRcolor0[737];
    UnbiasedRNG[13] = LFSRcolor0[467];
    UnbiasedRNG[14] = LFSRcolor0[349];
    UnbiasedRNG[15] = LFSRcolor0[1064];
    UnbiasedRNG[16] = LFSRcolor0[324];
    UnbiasedRNG[17] = LFSRcolor0[856];
    UnbiasedRNG[18] = LFSRcolor0[647];
    UnbiasedRNG[19] = LFSRcolor0[1000];
    UnbiasedRNG[20] = LFSRcolor0[417];
    UnbiasedRNG[21] = LFSRcolor0[772];
    UnbiasedRNG[22] = LFSRcolor0[548];
    UnbiasedRNG[23] = LFSRcolor0[1164];
    UnbiasedRNG[24] = LFSRcolor0[708];
    UnbiasedRNG[25] = LFSRcolor0[89];
    UnbiasedRNG[26] = LFSRcolor0[802];
    UnbiasedRNG[27] = LFSRcolor0[1099];
    UnbiasedRNG[28] = LFSRcolor0[691];
    UnbiasedRNG[29] = LFSRcolor0[864];
    UnbiasedRNG[30] = LFSRcolor0[170];
    UnbiasedRNG[31] = LFSRcolor0[874];
    UnbiasedRNG[32] = LFSRcolor0[215];
    UnbiasedRNG[33] = LFSRcolor0[1111];
    UnbiasedRNG[34] = LFSRcolor0[213];
    UnbiasedRNG[35] = LFSRcolor0[653];
    UnbiasedRNG[36] = LFSRcolor0[851];
    UnbiasedRNG[37] = LFSRcolor0[1128];
    UnbiasedRNG[38] = LFSRcolor0[734];
    UnbiasedRNG[39] = LFSRcolor0[988];
    UnbiasedRNG[40] = LFSRcolor0[1237];
    UnbiasedRNG[41] = LFSRcolor0[79];
    UnbiasedRNG[42] = LFSRcolor0[760];
    UnbiasedRNG[43] = LFSRcolor0[1117];
    UnbiasedRNG[44] = LFSRcolor0[1136];
    UnbiasedRNG[45] = LFSRcolor0[928];
    UnbiasedRNG[46] = LFSRcolor0[247];
    UnbiasedRNG[47] = LFSRcolor0[489];
    UnbiasedRNG[48] = LFSRcolor0[332];
    UnbiasedRNG[49] = LFSRcolor0[964];
    UnbiasedRNG[50] = LFSRcolor0[1044];
    UnbiasedRNG[51] = LFSRcolor0[1046];
    UnbiasedRNG[52] = LFSRcolor0[394];
    UnbiasedRNG[53] = LFSRcolor0[1230];
    UnbiasedRNG[54] = LFSRcolor0[1206];
    UnbiasedRNG[55] = LFSRcolor0[1176];
    UnbiasedRNG[56] = LFSRcolor0[17];
    UnbiasedRNG[57] = LFSRcolor0[174];
    UnbiasedRNG[58] = LFSRcolor0[785];
    UnbiasedRNG[59] = LFSRcolor0[794];
    UnbiasedRNG[60] = LFSRcolor0[279];
    UnbiasedRNG[61] = LFSRcolor0[407];
    UnbiasedRNG[62] = LFSRcolor0[1032];
    UnbiasedRNG[63] = LFSRcolor0[965];
    UnbiasedRNG[64] = LFSRcolor0[409];
    UnbiasedRNG[65] = LFSRcolor0[196];
    UnbiasedRNG[66] = LFSRcolor0[129];
    UnbiasedRNG[67] = LFSRcolor0[800];
    UnbiasedRNG[68] = LFSRcolor0[623];
    UnbiasedRNG[69] = LFSRcolor0[92];
    UnbiasedRNG[70] = LFSRcolor0[604];
    UnbiasedRNG[71] = LFSRcolor0[672];
    UnbiasedRNG[72] = LFSRcolor0[826];
    UnbiasedRNG[73] = LFSRcolor0[156];
    UnbiasedRNG[74] = LFSRcolor0[1086];
    UnbiasedRNG[75] = LFSRcolor0[364];
    UnbiasedRNG[76] = LFSRcolor0[848];
    UnbiasedRNG[77] = LFSRcolor0[866];
    UnbiasedRNG[78] = LFSRcolor0[463];
    UnbiasedRNG[79] = LFSRcolor0[141];
    UnbiasedRNG[80] = LFSRcolor0[433];
    UnbiasedRNG[81] = LFSRcolor0[1165];
    UnbiasedRNG[82] = LFSRcolor0[580];
    UnbiasedRNG[83] = LFSRcolor0[683];
    UnbiasedRNG[84] = LFSRcolor0[165];
    UnbiasedRNG[85] = LFSRcolor0[1048];
    UnbiasedRNG[86] = LFSRcolor0[983];
    UnbiasedRNG[87] = LFSRcolor0[342];
    UnbiasedRNG[88] = LFSRcolor0[806];
    UnbiasedRNG[89] = LFSRcolor0[81];
    UnbiasedRNG[90] = LFSRcolor0[470];
    UnbiasedRNG[91] = LFSRcolor0[645];
    UnbiasedRNG[92] = LFSRcolor0[199];
    UnbiasedRNG[93] = LFSRcolor0[797];
    UnbiasedRNG[94] = LFSRcolor0[971];
    UnbiasedRNG[95] = LFSRcolor0[21];
    UnbiasedRNG[96] = LFSRcolor0[712];
    UnbiasedRNG[97] = LFSRcolor0[878];
    UnbiasedRNG[98] = LFSRcolor0[674];
    UnbiasedRNG[99] = LFSRcolor0[67];
    UnbiasedRNG[100] = LFSRcolor0[284];
    UnbiasedRNG[101] = LFSRcolor0[1210];
    UnbiasedRNG[102] = LFSRcolor0[885];
    UnbiasedRNG[103] = LFSRcolor0[1002];
    UnbiasedRNG[104] = LFSRcolor0[903];
    UnbiasedRNG[105] = LFSRcolor0[1071];
    UnbiasedRNG[106] = LFSRcolor0[1157];
    UnbiasedRNG[107] = LFSRcolor0[474];
    UnbiasedRNG[108] = LFSRcolor0[572];
    UnbiasedRNG[109] = LFSRcolor0[1105];
    UnbiasedRNG[110] = LFSRcolor0[123];
    UnbiasedRNG[111] = LFSRcolor0[1034];
    UnbiasedRNG[112] = LFSRcolor0[930];
    UnbiasedRNG[113] = LFSRcolor0[345];
    UnbiasedRNG[114] = LFSRcolor0[768];
    UnbiasedRNG[115] = LFSRcolor0[459];
    UnbiasedRNG[116] = LFSRcolor0[1166];
    UnbiasedRNG[117] = LFSRcolor0[841];
    UnbiasedRNG[118] = LFSRcolor0[821];
    UnbiasedRNG[119] = LFSRcolor0[57];
    UnbiasedRNG[120] = LFSRcolor0[908];
    UnbiasedRNG[121] = LFSRcolor0[837];
    UnbiasedRNG[122] = LFSRcolor0[777];
    UnbiasedRNG[123] = LFSRcolor0[289];
    UnbiasedRNG[124] = LFSRcolor0[116];
    UnbiasedRNG[125] = LFSRcolor0[667];
    UnbiasedRNG[126] = LFSRcolor0[336];
    UnbiasedRNG[127] = LFSRcolor0[982];
    UnbiasedRNG[128] = LFSRcolor0[527];
    UnbiasedRNG[129] = LFSRcolor0[205];
    UnbiasedRNG[130] = LFSRcolor0[1141];
    UnbiasedRNG[131] = LFSRcolor0[842];
    UnbiasedRNG[132] = LFSRcolor0[378];
    UnbiasedRNG[133] = LFSRcolor0[124];
    UnbiasedRNG[134] = LFSRcolor0[68];
    UnbiasedRNG[135] = LFSRcolor0[315];
    UnbiasedRNG[136] = LFSRcolor0[220];
    UnbiasedRNG[137] = LFSRcolor0[857];
    UnbiasedRNG[138] = LFSRcolor0[1067];
    UnbiasedRNG[139] = LFSRcolor0[743];
    UnbiasedRNG[140] = LFSRcolor0[529];
    UnbiasedRNG[141] = LFSRcolor0[827];
    UnbiasedRNG[142] = LFSRcolor0[788];
    UnbiasedRNG[143] = LFSRcolor0[91];
    UnbiasedRNG[144] = LFSRcolor0[106];
    UnbiasedRNG[145] = LFSRcolor0[341];
    UnbiasedRNG[146] = LFSRcolor0[146];
    UnbiasedRNG[147] = LFSRcolor0[732];
    UnbiasedRNG[148] = LFSRcolor0[591];
    UnbiasedRNG[149] = LFSRcolor0[1236];
    UnbiasedRNG[150] = LFSRcolor0[1235];
    UnbiasedRNG[151] = LFSRcolor0[323];
    UnbiasedRNG[152] = LFSRcolor0[700];
    UnbiasedRNG[153] = LFSRcolor0[773];
    UnbiasedRNG[154] = LFSRcolor0[882];
    UnbiasedRNG[155] = LFSRcolor0[147];
    UnbiasedRNG[156] = LFSRcolor0[1135];
    UnbiasedRNG[157] = LFSRcolor0[692];
    UnbiasedRNG[158] = LFSRcolor0[1009];
    UnbiasedRNG[159] = LFSRcolor0[431];
    UnbiasedRNG[160] = LFSRcolor0[1129];
    UnbiasedRNG[161] = LFSRcolor0[486];
    UnbiasedRNG[162] = LFSRcolor0[78];
    UnbiasedRNG[163] = LFSRcolor0[175];
    UnbiasedRNG[164] = LFSRcolor0[375];
    UnbiasedRNG[165] = LFSRcolor0[698];
    UnbiasedRNG[166] = LFSRcolor0[435];
    UnbiasedRNG[167] = LFSRcolor0[607];
    UnbiasedRNG[168] = LFSRcolor0[1102];
    UnbiasedRNG[169] = LFSRcolor0[898];
    UnbiasedRNG[170] = LFSRcolor0[476];
    UnbiasedRNG[171] = LFSRcolor0[87];
    UnbiasedRNG[172] = LFSRcolor0[503];
    UnbiasedRNG[173] = LFSRcolor0[1058];
    UnbiasedRNG[174] = LFSRcolor0[918];
    UnbiasedRNG[175] = LFSRcolor0[629];
    UnbiasedRNG[176] = LFSRcolor0[1101];
    UnbiasedRNG[177] = LFSRcolor0[642];
    UnbiasedRNG[178] = LFSRcolor0[100];
    UnbiasedRNG[179] = LFSRcolor0[946];
    UnbiasedRNG[180] = LFSRcolor0[54];
    UnbiasedRNG[181] = LFSRcolor0[1213];
    UnbiasedRNG[182] = LFSRcolor0[1146];
    UnbiasedRNG[183] = LFSRcolor0[710];
    UnbiasedRNG[184] = LFSRcolor0[1043];
    UnbiasedRNG[185] = LFSRcolor0[1055];
    UnbiasedRNG[186] = LFSRcolor0[1108];
    UnbiasedRNG[187] = LFSRcolor0[1008];
    UnbiasedRNG[188] = LFSRcolor0[564];
    UnbiasedRNG[189] = LFSRcolor0[224];
    UnbiasedRNG[190] = LFSRcolor0[789];
    UnbiasedRNG[191] = LFSRcolor0[65];
    UnbiasedRNG[192] = LFSRcolor0[1220];
    UnbiasedRNG[193] = LFSRcolor0[309];
    UnbiasedRNG[194] = LFSRcolor0[532];
    UnbiasedRNG[195] = LFSRcolor0[1175];
    UnbiasedRNG[196] = LFSRcolor0[999];
    UnbiasedRNG[197] = LFSRcolor0[429];
    UnbiasedRNG[198] = LFSRcolor0[412];
    UnbiasedRNG[199] = LFSRcolor0[272];
    UnbiasedRNG[200] = LFSRcolor0[902];
    UnbiasedRNG[201] = LFSRcolor0[1216];
    UnbiasedRNG[202] = LFSRcolor0[0];
    UnbiasedRNG[203] = LFSRcolor0[461];
    UnbiasedRNG[204] = LFSRcolor0[601];
    UnbiasedRNG[205] = LFSRcolor0[705];
    UnbiasedRNG[206] = LFSRcolor0[704];
    UnbiasedRNG[207] = LFSRcolor0[1219];
    UnbiasedRNG[208] = LFSRcolor0[1198];
end

always @(posedge color0_clk) begin
    BiasedRNG[252] = (LFSRcolor1[304]&LFSRcolor1[360]&LFSRcolor1[1106]&LFSRcolor1[513]);
    BiasedRNG[253] = (LFSRcolor1[263]&LFSRcolor1[268]&LFSRcolor1[557]&LFSRcolor1[761]);
    BiasedRNG[254] = (LFSRcolor1[717]&LFSRcolor1[517]&LFSRcolor1[456]&LFSRcolor1[973]);
    BiasedRNG[255] = (LFSRcolor1[965]&LFSRcolor1[375]&LFSRcolor1[695]&LFSRcolor1[587]);
    BiasedRNG[256] = (LFSRcolor1[994]&LFSRcolor1[368]&LFSRcolor1[1049]&LFSRcolor1[802]);
    BiasedRNG[257] = (LFSRcolor1[525]&LFSRcolor1[831]&LFSRcolor1[852]&LFSRcolor1[112]);
    BiasedRNG[258] = (LFSRcolor1[668]&LFSRcolor1[483]&LFSRcolor1[716]&LFSRcolor1[433]);
    BiasedRNG[259] = (LFSRcolor1[825]&LFSRcolor1[756]&LFSRcolor1[816]&LFSRcolor1[390]);
    BiasedRNG[260] = (LFSRcolor1[77]&LFSRcolor1[1180]&LFSRcolor1[1104]&LFSRcolor1[738]);
    BiasedRNG[261] = (LFSRcolor1[70]&LFSRcolor1[235]&LFSRcolor1[697]&LFSRcolor1[206]);
    BiasedRNG[262] = (LFSRcolor1[219]&LFSRcolor1[934]&LFSRcolor1[552]&LFSRcolor1[735]);
    BiasedRNG[263] = (LFSRcolor1[150]&LFSRcolor1[277]&LFSRcolor1[956]&LFSRcolor1[937]);
    BiasedRNG[264] = (LFSRcolor1[622]&LFSRcolor1[1146]&LFSRcolor1[699]&LFSRcolor1[575]);
    BiasedRNG[265] = (LFSRcolor1[174]&LFSRcolor1[907]&LFSRcolor1[187]&LFSRcolor1[1073]);
    BiasedRNG[266] = (LFSRcolor1[527]&LFSRcolor1[156]&LFSRcolor1[630]&LFSRcolor1[922]);
    BiasedRNG[267] = (LFSRcolor1[20]&LFSRcolor1[100]&LFSRcolor1[157]&LFSRcolor1[447]);
    BiasedRNG[268] = (LFSRcolor1[32]&LFSRcolor1[1051]&LFSRcolor1[1076]&LFSRcolor1[336]);
    BiasedRNG[269] = (LFSRcolor1[801]&LFSRcolor1[679]&LFSRcolor1[786]&LFSRcolor1[496]);
    BiasedRNG[270] = (LFSRcolor1[538]&LFSRcolor1[615]&LFSRcolor1[777]&LFSRcolor1[216]);
    BiasedRNG[271] = (LFSRcolor1[993]&LFSRcolor1[896]&LFSRcolor1[388]&LFSRcolor1[69]);
    BiasedRNG[272] = (LFSRcolor1[95]&LFSRcolor1[602]&LFSRcolor1[395]&LFSRcolor1[689]);
    BiasedRNG[273] = (LFSRcolor1[1096]&LFSRcolor1[1166]&LFSRcolor1[259]&LFSRcolor1[1005]);
    BiasedRNG[274] = (LFSRcolor1[901]&LFSRcolor1[265]&LFSRcolor1[1010]&LFSRcolor1[1002]);
    BiasedRNG[275] = (LFSRcolor1[539]&LFSRcolor1[505]&LFSRcolor1[252]&LFSRcolor1[325]);
    BiasedRNG[276] = (LFSRcolor1[1009]&LFSRcolor1[814]&LFSRcolor1[136]&LFSRcolor1[149]);
    BiasedRNG[277] = (LFSRcolor1[534]&LFSRcolor1[1056]&LFSRcolor1[789]&LFSRcolor1[308]);
    BiasedRNG[278] = (LFSRcolor1[611]&LFSRcolor1[427]&LFSRcolor1[613]&LFSRcolor1[260]);
    BiasedRNG[279] = (LFSRcolor1[46]&LFSRcolor1[908]&LFSRcolor1[970]&LFSRcolor1[102]);
    BiasedRNG[280] = (LFSRcolor1[1047]&LFSRcolor1[1178]&LFSRcolor1[628]&LFSRcolor1[551]);
    BiasedRNG[281] = (LFSRcolor1[72]&LFSRcolor1[1082]&LFSRcolor1[410]&LFSRcolor1[126]);
    BiasedRNG[282] = (LFSRcolor1[929]&LFSRcolor1[196]&LFSRcolor1[846]&LFSRcolor1[197]);
    BiasedRNG[283] = (LFSRcolor1[221]&LFSRcolor1[439]&LFSRcolor1[14]&LFSRcolor1[512]);
    BiasedRNG[284] = (LFSRcolor1[921]&LFSRcolor1[598]&LFSRcolor1[807]&LFSRcolor1[25]);
    BiasedRNG[285] = (LFSRcolor1[230]&LFSRcolor1[1]&LFSRcolor1[838]&LFSRcolor1[317]);
    BiasedRNG[286] = (LFSRcolor1[741]&LFSRcolor1[1130]&LFSRcolor1[680]&LFSRcolor1[114]);
    BiasedRNG[287] = (LFSRcolor1[573]&LFSRcolor1[1000]&LFSRcolor1[339]&LFSRcolor1[683]);
    BiasedRNG[288] = (LFSRcolor1[272]&LFSRcolor1[324]&LFSRcolor1[38]&LFSRcolor1[725]);
    BiasedRNG[289] = (LFSRcolor1[763]&LFSRcolor1[548]&LFSRcolor1[736]&LFSRcolor1[782]);
    BiasedRNG[290] = (LFSRcolor1[26]&LFSRcolor1[231]&LFSRcolor1[918]&LFSRcolor1[1025]);
    BiasedRNG[291] = (LFSRcolor1[347]&LFSRcolor1[982]&LFSRcolor1[58]&LFSRcolor1[132]);
    BiasedRNG[292] = (LFSRcolor1[1156]&LFSRcolor1[652]&LFSRcolor1[1041]&LFSRcolor1[1108]);
    BiasedRNG[293] = (LFSRcolor1[490]&LFSRcolor1[341]&LFSRcolor1[869]&LFSRcolor1[969]);
    BiasedRNG[294] = (LFSRcolor1[391]&LFSRcolor1[240]&LFSRcolor1[1048]&LFSRcolor1[64]);
    BiasedRNG[295] = (LFSRcolor1[37]&LFSRcolor1[808]&LFSRcolor1[979]&LFSRcolor1[1147]);
    BiasedRNG[296] = (LFSRcolor1[262]&LFSRcolor1[627]&LFSRcolor1[599]&LFSRcolor1[634]);
    BiasedRNG[297] = (LFSRcolor1[608]&LFSRcolor1[733]&LFSRcolor1[1081]&LFSRcolor1[530]);
    BiasedRNG[298] = (LFSRcolor1[919]&LFSRcolor1[83]&LFSRcolor1[104]&LFSRcolor1[729]);
    BiasedRNG[299] = (LFSRcolor1[1125]&LFSRcolor1[238]&LFSRcolor1[387]&LFSRcolor1[579]);
    BiasedRNG[300] = (LFSRcolor1[89]&LFSRcolor1[1139]&LFSRcolor1[1113]&LFSRcolor1[6]);
    BiasedRNG[301] = (LFSRcolor1[87]&LFSRcolor1[361]&LFSRcolor1[1007]&LFSRcolor1[809]);
    BiasedRNG[302] = (LFSRcolor1[312]&LFSRcolor1[392]&LFSRcolor1[402]&LFSRcolor1[228]);
    BiasedRNG[303] = (LFSRcolor1[559]&LFSRcolor1[314]&LFSRcolor1[643]&LFSRcolor1[642]);
    BiasedRNG[304] = (LFSRcolor1[435]&LFSRcolor1[254]&LFSRcolor1[181]&LFSRcolor1[549]);
    BiasedRNG[305] = (LFSRcolor1[631]&LFSRcolor1[463]&LFSRcolor1[894]&LFSRcolor1[567]);
    BiasedRNG[306] = (LFSRcolor1[843]&LFSRcolor1[337]&LFSRcolor1[620]&LFSRcolor1[185]);
    BiasedRNG[307] = (LFSRcolor1[526]&LFSRcolor1[172]&LFSRcolor1[1022]&LFSRcolor1[590]);
    BiasedRNG[308] = (LFSRcolor1[797]&LFSRcolor1[676]&LFSRcolor1[464]&LFSRcolor1[203]);
    BiasedRNG[309] = (LFSRcolor1[974]&LFSRcolor1[1114]&LFSRcolor1[52]&LFSRcolor1[438]);
    BiasedRNG[310] = (LFSRcolor1[1061]&LFSRcolor1[398]&LFSRcolor1[775]&LFSRcolor1[233]);
    BiasedRNG[311] = (LFSRcolor1[1018]&LFSRcolor1[218]&LFSRcolor1[237]&LFSRcolor1[887]);
    BiasedRNG[312] = (LFSRcolor1[718]&LFSRcolor1[61]&LFSRcolor1[1074]&LFSRcolor1[207]);
    BiasedRNG[313] = (LFSRcolor1[1179]&LFSRcolor1[633]&LFSRcolor1[712]&LFSRcolor1[619]);
    BiasedRNG[314] = (LFSRcolor1[857]&LFSRcolor1[847]&LFSRcolor1[616]&LFSRcolor1[201]);
    BiasedRNG[315] = (LFSRcolor1[374]&LFSRcolor1[1110]&LFSRcolor1[980]&LFSRcolor1[1191]);
    BiasedRNG[316] = (LFSRcolor1[140]&LFSRcolor1[721]&LFSRcolor1[499]&LFSRcolor1[1088]);
    BiasedRNG[317] = (LFSRcolor1[798]&LFSRcolor1[1059]&LFSRcolor1[1085]&LFSRcolor1[1115]);
    BiasedRNG[318] = (LFSRcolor1[576]&LFSRcolor1[161]&LFSRcolor1[988]&LFSRcolor1[376]);
    BiasedRNG[319] = (LFSRcolor1[222]&LFSRcolor1[188]&LFSRcolor1[179]&LFSRcolor1[1079]);
    BiasedRNG[320] = (LFSRcolor1[572]&LFSRcolor1[90]&LFSRcolor1[758]&LFSRcolor1[355]);
    BiasedRNG[321] = (LFSRcolor1[830]&LFSRcolor1[691]&LFSRcolor1[365]&LFSRcolor1[139]);
    BiasedRNG[322] = (LFSRcolor1[1121]&LFSRcolor1[470]&LFSRcolor1[243]&LFSRcolor1[940]);
    BiasedRNG[323] = (LFSRcolor1[476]&LFSRcolor1[737]&LFSRcolor1[609]&LFSRcolor1[1087]);
    BiasedRNG[324] = (LFSRcolor1[205]&LFSRcolor1[770]&LFSRcolor1[446]&LFSRcolor1[767]);
    BiasedRNG[325] = (LFSRcolor1[369]&LFSRcolor1[1168]&LFSRcolor1[183]&LFSRcolor1[635]);
    BiasedRNG[326] = (LFSRcolor1[1013]&LFSRcolor1[791]&LFSRcolor1[1117]&LFSRcolor1[867]);
    BiasedRNG[327] = (LFSRcolor1[593]&LFSRcolor1[531]&LFSRcolor1[1095]&LFSRcolor1[556]);
    BiasedRNG[328] = (LFSRcolor1[851]&LFSRcolor1[332]&LFSRcolor1[455]&LFSRcolor1[794]);
    BiasedRNG[329] = (LFSRcolor1[436]&LFSRcolor1[878]&LFSRcolor1[954]&LFSRcolor1[759]);
    BiasedRNG[330] = (LFSRcolor1[1099]&LFSRcolor1[560]&LFSRcolor1[708]&LFSRcolor1[316]);
    BiasedRNG[331] = (LFSRcolor1[674]&LFSRcolor1[1071]&LFSRcolor1[309]&LFSRcolor1[21]);
    BiasedRNG[332] = (LFSRcolor1[1158]&LFSRcolor1[773]&LFSRcolor1[577]&LFSRcolor1[251]);
    BiasedRNG[333] = (LFSRcolor1[292]&LFSRcolor1[601]&LFSRcolor1[923]&LFSRcolor1[764]);
    BiasedRNG[334] = (LFSRcolor1[440]&LFSRcolor1[768]&LFSRcolor1[184]&LFSRcolor1[778]);
    BiasedRNG[335] = (LFSRcolor1[389]&LFSRcolor1[202]&LFSRcolor1[650]&LFSRcolor1[790]);
    BiasedRNG[336] = (LFSRcolor1[494]&LFSRcolor1[968]&LFSRcolor1[424]&LFSRcolor1[1003]);
    BiasedRNG[337] = (LFSRcolor1[34]&LFSRcolor1[193]&LFSRcolor1[298]&LFSRcolor1[171]);
    BiasedRNG[338] = (LFSRcolor1[78]&LFSRcolor1[130]&LFSRcolor1[595]&LFSRcolor1[753]);
    BiasedRNG[339] = (LFSRcolor1[192]&LFSRcolor1[748]&LFSRcolor1[367]&LFSRcolor1[282]);
    BiasedRNG[340] = (LFSRcolor1[714]&LFSRcolor1[62]&LFSRcolor1[561]&LFSRcolor1[176]);
    BiasedRNG[341] = (LFSRcolor1[1089]&LFSRcolor1[82]&LFSRcolor1[844]&LFSRcolor1[227]);
    BiasedRNG[342] = (LFSRcolor1[429]&LFSRcolor1[811]&LFSRcolor1[854]&LFSRcolor1[465]);
    BiasedRNG[343] = (LFSRcolor1[3]&LFSRcolor1[845]&LFSRcolor1[574]&LFSRcolor1[881]);
    BiasedRNG[344] = (LFSRcolor1[1145]&LFSRcolor1[755]&LFSRcolor1[480]&LFSRcolor1[366]);
    BiasedRNG[345] = (LFSRcolor1[1140]&LFSRcolor1[752]&LFSRcolor1[264]&LFSRcolor1[295]);
    BiasedRNG[346] = (LFSRcolor1[999]&LFSRcolor1[134]&LFSRcolor1[978]&LFSRcolor1[484]);
    BiasedRNG[347] = (LFSRcolor1[884]&LFSRcolor1[315]&LFSRcolor1[564]&LFSRcolor1[431]);
    BiasedRNG[348] = (LFSRcolor1[1066]&LFSRcolor1[865]&LFSRcolor1[888]&LFSRcolor1[938]);
    BiasedRNG[349] = (LFSRcolor1[545]&LFSRcolor1[459]&LFSRcolor1[747]&LFSRcolor1[1046]);
    BiasedRNG[350] = (LFSRcolor1[396]&LFSRcolor1[849]&LFSRcolor1[1029]&LFSRcolor1[507]);
    BiasedRNG[351] = (LFSRcolor1[866]&LFSRcolor1[473]&LFSRcolor1[124]&LFSRcolor1[48]);
    BiasedRNG[352] = (LFSRcolor1[895]&LFSRcolor1[144]&LFSRcolor1[677]&LFSRcolor1[899]);
    BiasedRNG[353] = (LFSRcolor1[10]&LFSRcolor1[143]&LFSRcolor1[111]&LFSRcolor1[175]);
    BiasedRNG[354] = (LFSRcolor1[460]&LFSRcolor1[353]&LFSRcolor1[301]&LFSRcolor1[302]);
    BiasedRNG[355] = (LFSRcolor1[1163]&LFSRcolor1[1173]&LFSRcolor1[1050]&LFSRcolor1[930]);
    BiasedRNG[356] = (LFSRcolor1[698]&LFSRcolor1[1015]&LFSRcolor1[1080]&LFSRcolor1[358]);
    BiasedRNG[357] = (LFSRcolor1[1053]&LFSRcolor1[663]&LFSRcolor1[727]&LFSRcolor1[364]);
    BiasedRNG[358] = (LFSRcolor1[1111]&LFSRcolor1[1052]&LFSRcolor1[253]&LFSRcolor1[510]);
    BiasedRNG[359] = (LFSRcolor1[774]&LFSRcolor1[269]&LFSRcolor1[542]&LFSRcolor1[106]);
    BiasedRNG[360] = (LFSRcolor1[720]&LFSRcolor1[730]&LFSRcolor1[1045]&LFSRcolor1[672]);
    BiasedRNG[361] = (LFSRcolor1[329]&LFSRcolor1[297]&LFSRcolor1[582]&LFSRcolor1[750]);
    BiasedRNG[362] = (LFSRcolor1[874]&LFSRcolor1[322]&LFSRcolor1[294]&LFSRcolor1[1075]);
    BiasedRNG[363] = (LFSRcolor1[226]&LFSRcolor1[278]&LFSRcolor1[863]&LFSRcolor1[989]);
    BiasedRNG[364] = (LFSRcolor1[664]&LFSRcolor1[220]&LFSRcolor1[142]&LFSRcolor1[1164]);
    BiasedRNG[365] = (LFSRcolor1[653]&LFSRcolor1[271]&LFSRcolor1[624]&LFSRcolor1[853]);
    BiasedRNG[366] = (LFSRcolor1[79]&LFSRcolor1[502]&LFSRcolor1[732]&LFSRcolor1[67]);
    BiasedRNG[367] = (LFSRcolor1[17]&LFSRcolor1[122]&LFSRcolor1[955]&LFSRcolor1[370]);
    BiasedRNG[368] = (LFSRcolor1[701]&LFSRcolor1[1165]&LFSRcolor1[519]&LFSRcolor1[73]);
    BiasedRNG[369] = (LFSRcolor1[117]&LFSRcolor1[1062]&LFSRcolor1[804]&LFSRcolor1[518]);
    BiasedRNG[370] = (LFSRcolor1[267]&LFSRcolor1[600]&LFSRcolor1[909]&LFSRcolor1[357]);
    BiasedRNG[371] = (LFSRcolor1[877]&LFSRcolor1[275]&LFSRcolor1[1141]&LFSRcolor1[327]);
    BiasedRNG[372] = (LFSRcolor1[581]&LFSRcolor1[1167]&LFSRcolor1[76]&LFSRcolor1[246]);
    BiasedRNG[373] = (LFSRcolor1[163]&LFSRcolor1[409]&LFSRcolor1[133]&LFSRcolor1[98]);
    BiasedRNG[374] = (LFSRcolor1[647]&LFSRcolor1[585]&LFSRcolor1[660]&LFSRcolor1[638]);
    BiasedRNG[375] = (LFSRcolor1[318]&LFSRcolor1[461]&LFSRcolor1[898]&LFSRcolor1[1069]);
    BiasedRNG[376] = (LFSRcolor1[1177]&LFSRcolor1[1054]&LFSRcolor1[42]&LFSRcolor1[783]);
    BiasedRNG[377] = (LFSRcolor1[710]&LFSRcolor1[964]&LFSRcolor1[148]&LFSRcolor1[565]);
    BiasedRNG[378] = (LFSRcolor1[356]&LFSRcolor1[925]&LFSRcolor1[1036]&LFSRcolor1[850]);
    BiasedRNG[379] = (LFSRcolor1[408]&LFSRcolor1[1183]&LFSRcolor1[864]&LFSRcolor1[1078]);
    BiasedRNG[380] = (LFSRcolor1[607]&LFSRcolor1[11]&LFSRcolor1[51]&LFSRcolor1[23]);
    BiasedRNG[381] = (LFSRcolor1[30]&LFSRcolor1[855]&LFSRcolor1[771]&LFSRcolor1[234]);
    BiasedRNG[382] = (LFSRcolor1[1148]&LFSRcolor1[953]&LFSRcolor1[757]&LFSRcolor1[746]);
    BiasedRNG[383] = (LFSRcolor1[669]&LFSRcolor1[784]&LFSRcolor1[500]&LFSRcolor1[165]);
    BiasedRNG[384] = (LFSRcolor1[40]&LFSRcolor1[281]&LFSRcolor1[84]&LFSRcolor1[787]);
    BiasedRNG[385] = (LFSRcolor1[917]&LFSRcolor1[214]&LFSRcolor1[836]&LFSRcolor1[803]);
    BiasedRNG[386] = (LFSRcolor1[180]&LFSRcolor1[286]&LFSRcolor1[769]&LFSRcolor1[612]);
    BiasedRNG[387] = (LFSRcolor1[949]&LFSRcolor1[1154]&LFSRcolor1[1094]&LFSRcolor1[256]);
    BiasedRNG[388] = (LFSRcolor1[451]&LFSRcolor1[509]&LFSRcolor1[1188]&LFSRcolor1[1157]);
    BiasedRNG[389] = (LFSRcolor1[153]&LFSRcolor1[529]&LFSRcolor1[1030]&LFSRcolor1[967]);
    BiasedRNG[390] = (LFSRcolor1[1037]&LFSRcolor1[481]&LFSRcolor1[306]&LFSRcolor1[333]);
    BiasedRNG[391] = (LFSRcolor1[859]&LFSRcolor1[1162]&LFSRcolor1[478]&LFSRcolor1[430]);
    BiasedRNG[392] = (LFSRcolor1[562]&LFSRcolor1[96]&LFSRcolor1[837]&LFSRcolor1[501]);
    BiasedRNG[393] = (LFSRcolor1[709]&LFSRcolor1[121]&LFSRcolor1[65]&LFSRcolor1[734]);
    BiasedRNG[394] = (LFSRcolor1[707]&LFSRcolor1[544]&LFSRcolor1[467]&LFSRcolor1[702]);
    BiasedRNG[395] = (LFSRcolor1[1017]&LFSRcolor1[245]&LFSRcolor1[145]&LFSRcolor1[570]);
    BiasedRNG[396] = (LFSRcolor1[870]&LFSRcolor1[550]&LFSRcolor1[359]&LFSRcolor1[486]);
    BiasedRNG[397] = (LFSRcolor1[406]&LFSRcolor1[536]&LFSRcolor1[723]&LFSRcolor1[1070]);
    BiasedRNG[398] = (LFSRcolor1[662]&LFSRcolor1[810]&LFSRcolor1[806]&LFSRcolor1[532]);
    BiasedRNG[399] = (LFSRcolor1[19]&LFSRcolor1[403]&LFSRcolor1[313]&LFSRcolor1[841]);
    BiasedRNG[400] = (LFSRcolor1[694]&LFSRcolor1[1011]&LFSRcolor1[833]&LFSRcolor1[445]);
    BiasedRNG[401] = (LFSRcolor1[35]&LFSRcolor1[167]&LFSRcolor1[421]&LFSRcolor1[1169]);
    BiasedRNG[402] = (LFSRcolor1[742]&LFSRcolor1[832]&LFSRcolor1[1027]&LFSRcolor1[670]);
    BiasedRNG[403] = (LFSRcolor1[1176]&LFSRcolor1[86]&LFSRcolor1[1186]&LFSRcolor1[495]);
    BiasedRNG[404] = (LFSRcolor1[434]&LFSRcolor1[745]&LFSRcolor1[80]&LFSRcolor1[303]);
    BiasedRNG[405] = (LFSRcolor1[382]&LFSRcolor1[43]&LFSRcolor1[1135]&LFSRcolor1[726]);
    BiasedRNG[406] = (LFSRcolor1[1063]&LFSRcolor1[199]&LFSRcolor1[453]&LFSRcolor1[16]);
    BiasedRNG[407] = (LFSRcolor1[553]&LFSRcolor1[59]&LFSRcolor1[941]&LFSRcolor1[681]);
    BiasedRNG[408] = (LFSRcolor1[232]&LFSRcolor1[125]&LFSRcolor1[897]&LFSRcolor1[442]);
    BiasedRNG[409] = (LFSRcolor1[997]&LFSRcolor1[673]&LFSRcolor1[31]&LFSRcolor1[944]);
    BiasedRNG[410] = (LFSRcolor1[152]&LFSRcolor1[1004]&LFSRcolor1[0]&LFSRcolor1[649]);
    BiasedRNG[411] = (LFSRcolor1[1109]&LFSRcolor1[1097]&LFSRcolor1[210]&LFSRcolor1[284]);
    BiasedRNG[412] = (LFSRcolor1[984]&LFSRcolor1[131]&LFSRcolor1[972]&LFSRcolor1[18]);
    BiasedRNG[413] = (LFSRcolor1[818]&LFSRcolor1[189]&LFSRcolor1[300]&LFSRcolor1[340]);
    BiasedRNG[414] = (LFSRcolor1[1044]&LFSRcolor1[173]&LFSRcolor1[443]&LFSRcolor1[886]);
    BiasedRNG[415] = (LFSRcolor1[1038]&LFSRcolor1[154]&LFSRcolor1[648]&LFSRcolor1[349]);
    BiasedRNG[416] = (LFSRcolor1[475]&LFSRcolor1[249]&LFSRcolor1[346]&LFSRcolor1[822]);
    BiasedRNG[417] = (LFSRcolor1[289]&LFSRcolor1[554]&LFSRcolor1[876]&LFSRcolor1[916]);
    BiasedRNG[418] = (LFSRcolor1[1077]&LFSRcolor1[428]&LFSRcolor1[60]&LFSRcolor1[1153]);
    BiasedRNG[419] = (LFSRcolor1[110]&LFSRcolor1[120]&LFSRcolor1[950]&LFSRcolor1[880]);
    BiasedRNG[420] = (LFSRcolor1[799]&LFSRcolor1[785]&LFSRcolor1[779]&LFSRcolor1[75]);
    BiasedRNG[421] = (LFSRcolor1[488]&LFSRcolor1[939]&LFSRcolor1[812]&LFSRcolor1[1040]);
    BiasedRNG[422] = (LFSRcolor1[158]&LFSRcolor1[657]&LFSRcolor1[1142]&LFSRcolor1[618]);
    BiasedRNG[423] = (LFSRcolor1[1102]&LFSRcolor1[93]&LFSRcolor1[705]&LFSRcolor1[1187]);
    BiasedRNG[424] = (LFSRcolor1[273]&LFSRcolor1[1086]&LFSRcolor1[305]&LFSRcolor1[454]);
    BiasedRNG[425] = (LFSRcolor1[200]&LFSRcolor1[378]&LFSRcolor1[521]&LFSRcolor1[471]);
    BiasedRNG[426] = (LFSRcolor1[910]&LFSRcolor1[36]&LFSRcolor1[1001]&LFSRcolor1[856]);
    BiasedRNG[427] = (LFSRcolor1[22]&LFSRcolor1[414]&LFSRcolor1[780]&LFSRcolor1[9]);
    BiasedRNG[428] = (LFSRcolor1[450]&LFSRcolor1[393]&LFSRcolor1[212]&LFSRcolor1[686]);
    BiasedRNG[429] = (LFSRcolor1[94]&LFSRcolor1[693]&LFSRcolor1[963]&LFSRcolor1[946]);
    BiasedRNG[430] = (LFSRcolor1[474]&LFSRcolor1[28]&LFSRcolor1[377]&LFSRcolor1[477]);
    BiasedRNG[431] = (LFSRcolor1[528]&LFSRcolor1[626]&LFSRcolor1[99]&LFSRcolor1[1084]);
    BiasedRNG[432] = (LFSRcolor1[497]&LFSRcolor1[1112]&LFSRcolor1[108]&LFSRcolor1[45]);
    BiasedRNG[433] = (LFSRcolor1[250]&LFSRcolor1[147]&LFSRcolor1[604]&LFSRcolor1[920]);
    BiasedRNG[434] = (LFSRcolor1[1119]&LFSRcolor1[728]&LFSRcolor1[1192]&LFSRcolor1[688]);
    BiasedRNG[435] = (LFSRcolor1[990]&LFSRcolor1[912]&LFSRcolor1[614]&LFSRcolor1[546]);
    BiasedRNG[436] = (LFSRcolor1[580]&LFSRcolor1[330]&LFSRcolor1[690]&LFSRcolor1[606]);
    BiasedRNG[437] = (LFSRcolor1[1120]&LFSRcolor1[326]&LFSRcolor1[904]&LFSRcolor1[224]);
    BiasedRNG[438] = (LFSRcolor1[871]&LFSRcolor1[715]&LFSRcolor1[826]&LFSRcolor1[151]);
    BiasedRNG[439] = (LFSRcolor1[1136]&LFSRcolor1[283]&LFSRcolor1[821]&LFSRcolor1[135]);
    BiasedRNG[440] = (LFSRcolor1[828]&LFSRcolor1[762]&LFSRcolor1[1189]&LFSRcolor1[655]);
    BiasedRNG[441] = (LFSRcolor1[522]&LFSRcolor1[889]&LFSRcolor1[489]&LFSRcolor1[101]);
    BiasedRNG[442] = (LFSRcolor1[1060]&LFSRcolor1[636]&LFSRcolor1[319]&LFSRcolor1[744]);
    BiasedRNG[443] = (LFSRcolor1[675]&LFSRcolor1[432]&LFSRcolor1[1185]&LFSRcolor1[417]);
    BiasedRNG[444] = (LFSRcolor1[842]&LFSRcolor1[827]&LFSRcolor1[33]&LFSRcolor1[74]);
    BiasedRNG[445] = (LFSRcolor1[860]&LFSRcolor1[623]&LFSRcolor1[49]&LFSRcolor1[1144]);
    BiasedRNG[446] = (LFSRcolor1[665]&LFSRcolor1[53]&LFSRcolor1[1127]&LFSRcolor1[986]);
    BiasedRNG[447] = (LFSRcolor1[363]&LFSRcolor1[146]&LFSRcolor1[1016]&LFSRcolor1[1131]);
    BiasedRNG[448] = (LFSRcolor1[1181]&LFSRcolor1[947]&LFSRcolor1[731]&LFSRcolor1[7]);
    BiasedRNG[449] = (LFSRcolor1[217]&LFSRcolor1[523]&LFSRcolor1[129]&LFSRcolor1[41]);
    BiasedRNG[450] = (LFSRcolor1[795]&LFSRcolor1[1123]&LFSRcolor1[823]&LFSRcolor1[584]);
    BiasedRNG[451] = (LFSRcolor1[765]&LFSRcolor1[1161]&LFSRcolor1[1026]&LFSRcolor1[503]);
    BiasedRNG[452] = (LFSRcolor1[160]&LFSRcolor1[914]&LFSRcolor1[380]&LFSRcolor1[137]);
    BiasedRNG[453] = (LFSRcolor1[1031]&LFSRcolor1[211]&LFSRcolor1[942]&LFSRcolor1[639]);
    BiasedRNG[454] = (LFSRcolor1[1184]&LFSRcolor1[426]&LFSRcolor1[405]&LFSRcolor1[362]);
    BiasedRNG[455] = (LFSRcolor1[103]&LFSRcolor1[419]&LFSRcolor1[713]&LFSRcolor1[63]);
    BiasedRNG[456] = (LFSRcolor1[208]&LFSRcolor1[170]&LFSRcolor1[397]&LFSRcolor1[1012]);
    BiasedRNG[457] = (LFSRcolor1[81]&LFSRcolor1[383]&LFSRcolor1[1032]&LFSRcolor1[819]);
    BiasedRNG[458] = (LFSRcolor1[274]&LFSRcolor1[569]&LFSRcolor1[998]&LFSRcolor1[583]);
    BiasedRNG[459] = (LFSRcolor1[645]&LFSRcolor1[992]&LFSRcolor1[338]&LFSRcolor1[1190]);
    BiasedRNG[460] = (LFSRcolor1[879]&LFSRcolor1[1152]&LFSRcolor1[159]&LFSRcolor1[113]);
    BiasedRNG[461] = (LFSRcolor1[498]&LFSRcolor1[893]&LFSRcolor1[1129]&LFSRcolor1[905]);
    BiasedRNG[462] = (LFSRcolor1[1100]&LFSRcolor1[441]&LFSRcolor1[971]&LFSRcolor1[961]);
    BiasedRNG[463] = (LFSRcolor1[566]&LFSRcolor1[423]&LFSRcolor1[592]&LFSRcolor1[469]);
    BiasedRNG[464] = (LFSRcolor1[666]&LFSRcolor1[724]&LFSRcolor1[394]&LFSRcolor1[781]);
    BiasedRNG[465] = (LFSRcolor1[1021]&LFSRcolor1[164]&LFSRcolor1[520]&LFSRcolor1[661]);
    BiasedRNG[466] = (LFSRcolor1[1107]&LFSRcolor1[640]&LFSRcolor1[511]&LFSRcolor1[482]);
    BiasedRNG[467] = (LFSRcolor1[411]&LFSRcolor1[632]&LFSRcolor1[400]&LFSRcolor1[1065]);
    BiasedRNG[468] = (LFSRcolor1[817]&LFSRcolor1[625]&LFSRcolor1[1093]&LFSRcolor1[911]);
    BiasedRNG[469] = (LFSRcolor1[996]&LFSRcolor1[1103]&LFSRcolor1[987]&LFSRcolor1[524]);
    BiasedRNG[470] = (LFSRcolor1[547]&LFSRcolor1[47]&LFSRcolor1[535]&LFSRcolor1[873]);
    BiasedRNG[471] = (LFSRcolor1[1134]&LFSRcolor1[288]&LFSRcolor1[91]&LFSRcolor1[223]);
    BiasedRNG[472] = (LFSRcolor1[504]&LFSRcolor1[351]&LFSRcolor1[379]&LFSRcolor1[1151]);
    BiasedRNG[473] = (LFSRcolor1[533]&LFSRcolor1[682]&LFSRcolor1[687]&LFSRcolor1[617]);
    BiasedRNG[474] = (LFSRcolor1[485]&LFSRcolor1[307]&LFSRcolor1[343]&LFSRcolor1[586]);
    BiasedRNG[475] = (LFSRcolor1[412]&LFSRcolor1[105]&LFSRcolor1[335]&LFSRcolor1[119]);
    BiasedRNG[476] = (LFSRcolor1[15]&LFSRcolor1[1195]&LFSRcolor1[568]&LFSRcolor1[966]);
    BiasedRNG[477] = (LFSRcolor1[516]&LFSRcolor1[678]&LFSRcolor1[890]&LFSRcolor1[711]);
    BiasedRNG[478] = (LFSRcolor1[399]&LFSRcolor1[558]&LFSRcolor1[492]&LFSRcolor1[248]);
    BiasedRNG[479] = (LFSRcolor1[279]&LFSRcolor1[514]&LFSRcolor1[241]&LFSRcolor1[71]);
    BiasedRNG[480] = (LFSRcolor1[168]&LFSRcolor1[141]&LFSRcolor1[646]&LFSRcolor1[299]);
    BiasedRNG[481] = (LFSRcolor1[792]&LFSRcolor1[5]&LFSRcolor1[515]&LFSRcolor1[350]);
    BiasedRNG[482] = (LFSRcolor1[169]&LFSRcolor1[1068]&LFSRcolor1[1132]&LFSRcolor1[981]);
    BiasedRNG[483] = (LFSRcolor1[861]&LFSRcolor1[457]&LFSRcolor1[594]&LFSRcolor1[1138]);
    BiasedRNG[484] = (LFSRcolor1[413]&LFSRcolor1[1137]&LFSRcolor1[591]&LFSRcolor1[692]);
    BiasedRNG[485] = (LFSRcolor1[1023]&LFSRcolor1[882]&LFSRcolor1[578]&LFSRcolor1[213]);
    BiasedRNG[486] = (LFSRcolor1[541]&LFSRcolor1[700]&LFSRcolor1[386]&LFSRcolor1[719]);
    BiasedRNG[487] = (LFSRcolor1[1024]&LFSRcolor1[766]&LFSRcolor1[915]&LFSRcolor1[1055]);
    BiasedRNG[488] = (LFSRcolor1[1020]&LFSRcolor1[229]&LFSRcolor1[109]&LFSRcolor1[491]);
    BiasedRNG[489] = (LFSRcolor1[537]&LFSRcolor1[24]&LFSRcolor1[1034]&LFSRcolor1[1019]);
    BiasedRNG[490] = (LFSRcolor1[820]&LFSRcolor1[416]&LFSRcolor1[788]&LFSRcolor1[739]);
    BiasedRNG[491] = (LFSRcolor1[128]&LFSRcolor1[373]&LFSRcolor1[805]&LFSRcolor1[466]);
    BiasedRNG[492] = (LFSRcolor1[667]&LFSRcolor1[66]&LFSRcolor1[116]&LFSRcolor1[858]);
    BiasedRNG[493] = (LFSRcolor1[829]&LFSRcolor1[751]&LFSRcolor1[437]&LFSRcolor1[493]);
    BiasedRNG[494] = (LFSRcolor1[596]&LFSRcolor1[945]&LFSRcolor1[107]&LFSRcolor1[462]);
    BiasedRNG[495] = (LFSRcolor1[321]&LFSRcolor1[815]&LFSRcolor1[958]&LFSRcolor1[540]);
    BiasedRNG[496] = (LFSRcolor1[848]&LFSRcolor1[50]&LFSRcolor1[1035]&LFSRcolor1[995]);
    BiasedRNG[497] = (LFSRcolor1[1006]&LFSRcolor1[872]&LFSRcolor1[749]&LFSRcolor1[885]);
    BiasedRNG[498] = (LFSRcolor1[928]&LFSRcolor1[588]&LFSRcolor1[891]&LFSRcolor1[276]);
    BiasedRNG[499] = (LFSRcolor1[824]&LFSRcolor1[354]&LFSRcolor1[204]&LFSRcolor1[166]);
    BiasedRNG[500] = (LFSRcolor1[178]&LFSRcolor1[97]&LFSRcolor1[685]&LFSRcolor1[936]);
    BiasedRNG[501] = (LFSRcolor1[44]&LFSRcolor1[458]&LFSRcolor1[868]&LFSRcolor1[266]);
    BiasedRNG[502] = (LFSRcolor1[415]&LFSRcolor1[385]&LFSRcolor1[311]&LFSRcolor1[1172]);
    UnbiasedRNG[209] = LFSRcolor1[310];
    UnbiasedRNG[210] = LFSRcolor1[244];
    UnbiasedRNG[211] = LFSRcolor1[1171];
    UnbiasedRNG[212] = LFSRcolor1[258];
    UnbiasedRNG[213] = LFSRcolor1[1159];
    UnbiasedRNG[214] = LFSRcolor1[754];
    UnbiasedRNG[215] = LFSRcolor1[1170];
    UnbiasedRNG[216] = LFSRcolor1[597];
    UnbiasedRNG[217] = LFSRcolor1[1033];
    UnbiasedRNG[218] = LFSRcolor1[621];
    UnbiasedRNG[219] = LFSRcolor1[407];
    UnbiasedRNG[220] = LFSRcolor1[903];
    UnbiasedRNG[221] = LFSRcolor1[1008];
    UnbiasedRNG[222] = LFSRcolor1[931];
    UnbiasedRNG[223] = LFSRcolor1[659];
    UnbiasedRNG[224] = LFSRcolor1[706];
    UnbiasedRNG[225] = LFSRcolor1[285];
    UnbiasedRNG[226] = LFSRcolor1[975];
    UnbiasedRNG[227] = LFSRcolor1[209];
    UnbiasedRNG[228] = LFSRcolor1[1193];
    UnbiasedRNG[229] = LFSRcolor1[123];
    UnbiasedRNG[230] = LFSRcolor1[983];
    UnbiasedRNG[231] = LFSRcolor1[1101];
    UnbiasedRNG[232] = LFSRcolor1[177];
    UnbiasedRNG[233] = LFSRcolor1[472];
    UnbiasedRNG[234] = LFSRcolor1[1155];
    UnbiasedRNG[235] = LFSRcolor1[948];
    UnbiasedRNG[236] = LFSRcolor1[344];
    UnbiasedRNG[237] = LFSRcolor1[444];
    UnbiasedRNG[238] = LFSRcolor1[242];
    UnbiasedRNG[239] = LFSRcolor1[1043];
    UnbiasedRNG[240] = LFSRcolor1[1042];
    UnbiasedRNG[241] = LFSRcolor1[293];
    UnbiasedRNG[242] = LFSRcolor1[722];
    UnbiasedRNG[243] = LFSRcolor1[704];
    UnbiasedRNG[244] = LFSRcolor1[875];
    UnbiasedRNG[245] = LFSRcolor1[420];
    UnbiasedRNG[246] = LFSRcolor1[138];
    UnbiasedRNG[247] = LFSRcolor1[605];
    UnbiasedRNG[248] = LFSRcolor1[1116];
    UnbiasedRNG[249] = LFSRcolor1[236];
    UnbiasedRNG[250] = LFSRcolor1[55];
    UnbiasedRNG[251] = LFSRcolor1[1105];
    UnbiasedRNG[252] = LFSRcolor1[449];
    UnbiasedRNG[253] = LFSRcolor1[239];
    UnbiasedRNG[254] = LFSRcolor1[331];
    UnbiasedRNG[255] = LFSRcolor1[1064];
    UnbiasedRNG[256] = LFSRcolor1[215];
    UnbiasedRNG[257] = LFSRcolor1[12];
    UnbiasedRNG[258] = LFSRcolor1[985];
    UnbiasedRNG[259] = LFSRcolor1[883];
    UnbiasedRNG[260] = LFSRcolor1[793];
    UnbiasedRNG[261] = LFSRcolor1[913];
    UnbiasedRNG[262] = LFSRcolor1[182];
    UnbiasedRNG[263] = LFSRcolor1[261];
    UnbiasedRNG[264] = LFSRcolor1[1083];
    UnbiasedRNG[265] = LFSRcolor1[603];
    UnbiasedRNG[266] = LFSRcolor1[834];
    UnbiasedRNG[267] = LFSRcolor1[1091];
    UnbiasedRNG[268] = LFSRcolor1[800];
    UnbiasedRNG[269] = LFSRcolor1[696];
    UnbiasedRNG[270] = LFSRcolor1[54];
    UnbiasedRNG[271] = LFSRcolor1[906];
    UnbiasedRNG[272] = LFSRcolor1[418];
    UnbiasedRNG[273] = LFSRcolor1[296];
    UnbiasedRNG[274] = LFSRcolor1[951];
    UnbiasedRNG[275] = LFSRcolor1[772];
    UnbiasedRNG[276] = LFSRcolor1[1028];
    UnbiasedRNG[277] = LFSRcolor1[1039];
    UnbiasedRNG[278] = LFSRcolor1[637];
    UnbiasedRNG[279] = LFSRcolor1[563];
    UnbiasedRNG[280] = LFSRcolor1[1126];
    UnbiasedRNG[281] = LFSRcolor1[977];
    UnbiasedRNG[282] = LFSRcolor1[1149];
    UnbiasedRNG[283] = LFSRcolor1[656];
    UnbiasedRNG[284] = LFSRcolor1[345];
    UnbiasedRNG[285] = LFSRcolor1[932];
    UnbiasedRNG[286] = LFSRcolor1[813];
    UnbiasedRNG[287] = LFSRcolor1[372];
    UnbiasedRNG[288] = LFSRcolor1[1067];
    UnbiasedRNG[289] = LFSRcolor1[760];
    UnbiasedRNG[290] = LFSRcolor1[658];
    UnbiasedRNG[291] = LFSRcolor1[127];
    UnbiasedRNG[292] = LFSRcolor1[629];
    UnbiasedRNG[293] = LFSRcolor1[644];
    UnbiasedRNG[294] = LFSRcolor1[555];
    UnbiasedRNG[295] = LFSRcolor1[291];
    UnbiasedRNG[296] = LFSRcolor1[840];
    UnbiasedRNG[297] = LFSRcolor1[641];
    UnbiasedRNG[298] = LFSRcolor1[684];
    UnbiasedRNG[299] = LFSRcolor1[1092];
    UnbiasedRNG[300] = LFSRcolor1[651];
    UnbiasedRNG[301] = LFSRcolor1[926];
    UnbiasedRNG[302] = LFSRcolor1[703];
    UnbiasedRNG[303] = LFSRcolor1[8];
    UnbiasedRNG[304] = LFSRcolor1[371];
    UnbiasedRNG[305] = LFSRcolor1[933];
    UnbiasedRNG[306] = LFSRcolor1[13];
    UnbiasedRNG[307] = LFSRcolor1[654];
    UnbiasedRNG[308] = LFSRcolor1[194];
    UnbiasedRNG[309] = LFSRcolor1[1128];
    UnbiasedRNG[310] = LFSRcolor1[1118];
    UnbiasedRNG[311] = LFSRcolor1[960];
    UnbiasedRNG[312] = LFSRcolor1[927];
    UnbiasedRNG[313] = LFSRcolor1[487];
    UnbiasedRNG[314] = LFSRcolor1[957];
    UnbiasedRNG[315] = LFSRcolor1[1124];
    UnbiasedRNG[316] = LFSRcolor1[862];
    UnbiasedRNG[317] = LFSRcolor1[1058];
    UnbiasedRNG[318] = LFSRcolor1[835];
    UnbiasedRNG[319] = LFSRcolor1[186];
    UnbiasedRNG[320] = LFSRcolor1[198];
    UnbiasedRNG[321] = LFSRcolor1[68];
    UnbiasedRNG[322] = LFSRcolor1[900];
    UnbiasedRNG[323] = LFSRcolor1[328];
    UnbiasedRNG[324] = LFSRcolor1[270];
    UnbiasedRNG[325] = LFSRcolor1[571];
    UnbiasedRNG[326] = LFSRcolor1[404];
    UnbiasedRNG[327] = LFSRcolor1[796];
    UnbiasedRNG[328] = LFSRcolor1[839];
    UnbiasedRNG[329] = LFSRcolor1[115];
    UnbiasedRNG[330] = LFSRcolor1[935];
    UnbiasedRNG[331] = LFSRcolor1[401];
    UnbiasedRNG[332] = LFSRcolor1[290];
    UnbiasedRNG[333] = LFSRcolor1[323];
    UnbiasedRNG[334] = LFSRcolor1[776];
    UnbiasedRNG[335] = LFSRcolor1[943];
    UnbiasedRNG[336] = LFSRcolor1[1133];
    UnbiasedRNG[337] = LFSRcolor1[902];
    UnbiasedRNG[338] = LFSRcolor1[952];
    UnbiasedRNG[339] = LFSRcolor1[976];
    UnbiasedRNG[340] = LFSRcolor1[92];
    UnbiasedRNG[341] = LFSRcolor1[508];
    UnbiasedRNG[342] = LFSRcolor1[452];
    UnbiasedRNG[343] = LFSRcolor1[1150];
    UnbiasedRNG[344] = LFSRcolor1[1194];
    UnbiasedRNG[345] = LFSRcolor1[255];
    UnbiasedRNG[346] = LFSRcolor1[671];
    UnbiasedRNG[347] = LFSRcolor1[85];
    UnbiasedRNG[348] = LFSRcolor1[287];
    UnbiasedRNG[349] = LFSRcolor1[381];
    UnbiasedRNG[350] = LFSRcolor1[342];
    UnbiasedRNG[351] = LFSRcolor1[1098];
    UnbiasedRNG[352] = LFSRcolor1[589];
    UnbiasedRNG[353] = LFSRcolor1[88];
    UnbiasedRNG[354] = LFSRcolor1[962];
    UnbiasedRNG[355] = LFSRcolor1[155];
    UnbiasedRNG[356] = LFSRcolor1[334];
    UnbiasedRNG[357] = LFSRcolor1[743];
    UnbiasedRNG[358] = LFSRcolor1[190];
    UnbiasedRNG[359] = LFSRcolor1[39];
    UnbiasedRNG[360] = LFSRcolor1[1174];
    UnbiasedRNG[361] = LFSRcolor1[1057];
    UnbiasedRNG[362] = LFSRcolor1[348];
    UnbiasedRNG[363] = LFSRcolor1[991];
    UnbiasedRNG[364] = LFSRcolor1[506];
    UnbiasedRNG[365] = LFSRcolor1[448];
    UnbiasedRNG[366] = LFSRcolor1[191];
    UnbiasedRNG[367] = LFSRcolor1[162];
    UnbiasedRNG[368] = LFSRcolor1[195];
    UnbiasedRNG[369] = LFSRcolor1[740];
    UnbiasedRNG[370] = LFSRcolor1[1090];
    UnbiasedRNG[371] = LFSRcolor1[543];
    UnbiasedRNG[372] = LFSRcolor1[2];
    UnbiasedRNG[373] = LFSRcolor1[257];
    UnbiasedRNG[374] = LFSRcolor1[56];
    UnbiasedRNG[375] = LFSRcolor1[118];
    UnbiasedRNG[376] = LFSRcolor1[29];
    UnbiasedRNG[377] = LFSRcolor1[4];
    UnbiasedRNG[378] = LFSRcolor1[479];
    UnbiasedRNG[379] = LFSRcolor1[1160];
    UnbiasedRNG[380] = LFSRcolor1[280];
    UnbiasedRNG[381] = LFSRcolor1[384];
    UnbiasedRNG[382] = LFSRcolor1[352];
    UnbiasedRNG[383] = LFSRcolor1[247];
    UnbiasedRNG[384] = LFSRcolor1[892];
    UnbiasedRNG[385] = LFSRcolor1[422];
end

always @(posedge color1_clk) begin
    BiasedRNG[503] = (LFSRcolor2[706]&LFSRcolor2[932]&LFSRcolor2[658]&LFSRcolor2[117]);
    BiasedRNG[504] = (LFSRcolor2[812]&LFSRcolor2[729]&LFSRcolor2[251]&LFSRcolor2[310]);
    BiasedRNG[505] = (LFSRcolor2[496]&LFSRcolor2[542]&LFSRcolor2[488]&LFSRcolor2[578]);
    BiasedRNG[506] = (LFSRcolor2[635]&LFSRcolor2[197]&LFSRcolor2[500]&LFSRcolor2[770]);
    BiasedRNG[507] = (LFSRcolor2[851]&LFSRcolor2[568]&LFSRcolor2[59]&LFSRcolor2[247]);
    BiasedRNG[508] = (LFSRcolor2[92]&LFSRcolor2[725]&LFSRcolor2[81]&LFSRcolor2[847]);
    BiasedRNG[509] = (LFSRcolor2[203]&LFSRcolor2[96]&LFSRcolor2[576]&LFSRcolor2[107]);
    BiasedRNG[510] = (LFSRcolor2[227]&LFSRcolor2[631]&LFSRcolor2[917]&LFSRcolor2[487]);
    BiasedRNG[511] = (LFSRcolor2[905]&LFSRcolor2[718]&LFSRcolor2[611]&LFSRcolor2[938]);
    BiasedRNG[512] = (LFSRcolor2[7]&LFSRcolor2[595]&LFSRcolor2[46]&LFSRcolor2[777]);
    BiasedRNG[513] = (LFSRcolor2[243]&LFSRcolor2[530]&LFSRcolor2[538]&LFSRcolor2[510]);
    BiasedRNG[514] = (LFSRcolor2[387]&LFSRcolor2[583]&LFSRcolor2[385]&LFSRcolor2[226]);
    BiasedRNG[515] = (LFSRcolor2[79]&LFSRcolor2[775]&LFSRcolor2[460]&LFSRcolor2[318]);
    BiasedRNG[516] = (LFSRcolor2[41]&LFSRcolor2[25]&LFSRcolor2[432]&LFSRcolor2[813]);
    BiasedRNG[517] = (LFSRcolor2[624]&LFSRcolor2[957]&LFSRcolor2[669]&LFSRcolor2[850]);
    BiasedRNG[518] = (LFSRcolor2[228]&LFSRcolor2[914]&LFSRcolor2[731]&LFSRcolor2[116]);
    BiasedRNG[519] = (LFSRcolor2[605]&LFSRcolor2[807]&LFSRcolor2[489]&LFSRcolor2[527]);
    BiasedRNG[520] = (LFSRcolor2[463]&LFSRcolor2[443]&LFSRcolor2[627]&LFSRcolor2[152]);
    BiasedRNG[521] = (LFSRcolor2[505]&LFSRcolor2[588]&LFSRcolor2[214]&LFSRcolor2[467]);
    BiasedRNG[522] = (LFSRcolor2[415]&LFSRcolor2[963]&LFSRcolor2[19]&LFSRcolor2[926]);
    BiasedRNG[523] = (LFSRcolor2[283]&LFSRcolor2[535]&LFSRcolor2[295]&LFSRcolor2[659]);
    BiasedRNG[524] = (LFSRcolor2[862]&LFSRcolor2[778]&LFSRcolor2[419]&LFSRcolor2[185]);
    BiasedRNG[525] = (LFSRcolor2[177]&LFSRcolor2[787]&LFSRcolor2[786]&LFSRcolor2[934]);
    BiasedRNG[526] = (LFSRcolor2[908]&LFSRcolor2[918]&LFSRcolor2[162]&LFSRcolor2[38]);
    BiasedRNG[527] = (LFSRcolor2[698]&LFSRcolor2[766]&LFSRcolor2[114]&LFSRcolor2[49]);
    BiasedRNG[528] = (LFSRcolor2[546]&LFSRcolor2[520]&LFSRcolor2[100]&LFSRcolor2[35]);
    BiasedRNG[529] = (LFSRcolor2[883]&LFSRcolor2[414]&LFSRcolor2[94]&LFSRcolor2[187]);
    BiasedRNG[530] = (LFSRcolor2[321]&LFSRcolor2[964]&LFSRcolor2[276]&LFSRcolor2[916]);
    BiasedRNG[531] = (LFSRcolor2[449]&LFSRcolor2[286]&LFSRcolor2[367]&LFSRcolor2[944]);
    BiasedRNG[532] = (LFSRcolor2[896]&LFSRcolor2[167]&LFSRcolor2[597]&LFSRcolor2[62]);
    BiasedRNG[533] = (LFSRcolor2[362]&LFSRcolor2[893]&LFSRcolor2[333]&LFSRcolor2[477]);
    BiasedRNG[534] = (LFSRcolor2[231]&LFSRcolor2[131]&LFSRcolor2[40]&LFSRcolor2[223]);
    BiasedRNG[535] = (LFSRcolor2[547]&LFSRcolor2[532]&LFSRcolor2[80]&LFSRcolor2[651]);
    BiasedRNG[536] = (LFSRcolor2[765]&LFSRcolor2[182]&LFSRcolor2[349]&LFSRcolor2[345]);
    BiasedRNG[537] = (LFSRcolor2[585]&LFSRcolor2[895]&LFSRcolor2[269]&LFSRcolor2[143]);
    BiasedRNG[538] = (LFSRcolor2[374]&LFSRcolor2[159]&LFSRcolor2[347]&LFSRcolor2[313]);
    BiasedRNG[539] = (LFSRcolor2[302]&LFSRcolor2[685]&LFSRcolor2[907]&LFSRcolor2[561]);
    BiasedRNG[540] = (LFSRcolor2[697]&LFSRcolor2[453]&LFSRcolor2[93]&LFSRcolor2[327]);
    BiasedRNG[541] = (LFSRcolor2[260]&LFSRcolor2[202]&LFSRcolor2[300]&LFSRcolor2[853]);
    BiasedRNG[542] = (LFSRcolor2[480]&LFSRcolor2[626]&LFSRcolor2[475]&LFSRcolor2[4]);
    BiasedRNG[543] = (LFSRcolor2[816]&LFSRcolor2[402]&LFSRcolor2[495]&LFSRcolor2[240]);
    BiasedRNG[544] = (LFSRcolor2[579]&LFSRcolor2[346]&LFSRcolor2[910]&LFSRcolor2[137]);
    BiasedRNG[545] = (LFSRcolor2[222]&LFSRcolor2[656]&LFSRcolor2[359]&LFSRcolor2[852]);
    BiasedRNG[546] = (LFSRcolor2[254]&LFSRcolor2[391]&LFSRcolor2[193]&LFSRcolor2[9]);
    BiasedRNG[547] = (LFSRcolor2[21]&LFSRcolor2[919]&LFSRcolor2[365]&LFSRcolor2[95]);
    BiasedRNG[548] = (LFSRcolor2[408]&LFSRcolor2[44]&LFSRcolor2[1]&LFSRcolor2[544]);
    BiasedRNG[549] = (LFSRcolor2[838]&LFSRcolor2[573]&LFSRcolor2[471]&LFSRcolor2[672]);
    BiasedRNG[550] = (LFSRcolor2[78]&LFSRcolor2[22]&LFSRcolor2[702]&LFSRcolor2[762]);
    BiasedRNG[551] = (LFSRcolor2[829]&LFSRcolor2[550]&LFSRcolor2[737]&LFSRcolor2[634]);
    BiasedRNG[552] = (LFSRcolor2[504]&LFSRcolor2[363]&LFSRcolor2[750]&LFSRcolor2[229]);
    BiasedRNG[553] = (LFSRcolor2[653]&LFSRcolor2[430]&LFSRcolor2[366]&LFSRcolor2[519]);
    BiasedRNG[554] = (LFSRcolor2[413]&LFSRcolor2[219]&LFSRcolor2[435]&LFSRcolor2[929]);
    BiasedRNG[555] = (LFSRcolor2[275]&LFSRcolor2[873]&LFSRcolor2[484]&LFSRcolor2[288]);
    BiasedRNG[556] = (LFSRcolor2[90]&LFSRcolor2[861]&LFSRcolor2[736]&LFSRcolor2[600]);
    BiasedRNG[557] = (LFSRcolor2[841]&LFSRcolor2[171]&LFSRcolor2[705]&LFSRcolor2[297]);
    BiasedRNG[558] = (LFSRcolor2[562]&LFSRcolor2[213]&LFSRcolor2[921]&LFSRcolor2[678]);
    BiasedRNG[559] = (LFSRcolor2[65]&LFSRcolor2[749]&LFSRcolor2[590]&LFSRcolor2[582]);
    BiasedRNG[560] = (LFSRcolor2[632]&LFSRcolor2[709]&LFSRcolor2[48]&LFSRcolor2[72]);
    BiasedRNG[561] = (LFSRcolor2[294]&LFSRcolor2[422]&LFSRcolor2[784]&LFSRcolor2[328]);
    BiasedRNG[562] = (LFSRcolor2[405]&LFSRcolor2[891]&LFSRcolor2[8]&LFSRcolor2[936]);
    BiasedRNG[563] = (LFSRcolor2[221]&LFSRcolor2[132]&LFSRcolor2[450]&LFSRcolor2[139]);
    BiasedRNG[564] = (LFSRcolor2[403]&LFSRcolor2[781]&LFSRcolor2[864]&LFSRcolor2[45]);
    BiasedRNG[565] = (LFSRcolor2[623]&LFSRcolor2[503]&LFSRcolor2[559]&LFSRcolor2[198]);
    BiasedRNG[566] = (LFSRcolor2[311]&LFSRcolor2[596]&LFSRcolor2[879]&LFSRcolor2[343]);
    BiasedRNG[567] = (LFSRcolor2[526]&LFSRcolor2[20]&LFSRcolor2[869]&LFSRcolor2[512]);
    BiasedRNG[568] = (LFSRcolor2[289]&LFSRcolor2[312]&LFSRcolor2[67]&LFSRcolor2[820]);
    BiasedRNG[569] = (LFSRcolor2[109]&LFSRcolor2[60]&LFSRcolor2[639]&LFSRcolor2[833]);
    BiasedRNG[570] = (LFSRcolor2[75]&LFSRcolor2[522]&LFSRcolor2[170]&LFSRcolor2[560]);
    BiasedRNG[571] = (LFSRcolor2[12]&LFSRcolor2[800]&LFSRcolor2[695]&LFSRcolor2[335]);
    BiasedRNG[572] = (LFSRcolor2[734]&LFSRcolor2[947]&LFSRcolor2[620]&LFSRcolor2[429]);
    BiasedRNG[573] = (LFSRcolor2[101]&LFSRcolor2[466]&LFSRcolor2[662]&LFSRcolor2[148]);
    BiasedRNG[574] = (LFSRcolor2[353]&LFSRcolor2[395]&LFSRcolor2[806]&LFSRcolor2[446]);
    BiasedRNG[575] = (LFSRcolor2[790]&LFSRcolor2[299]&LFSRcolor2[404]&LFSRcolor2[281]);
    BiasedRNG[576] = (LFSRcolor2[665]&LFSRcolor2[523]&LFSRcolor2[375]&LFSRcolor2[715]);
    BiasedRNG[577] = (LFSRcolor2[144]&LFSRcolor2[180]&LFSRcolor2[188]&LFSRcolor2[215]);
    BiasedRNG[578] = (LFSRcolor2[931]&LFSRcolor2[845]&LFSRcolor2[558]&LFSRcolor2[748]);
    BiasedRNG[579] = (LFSRcolor2[710]&LFSRcolor2[580]&LFSRcolor2[370]&LFSRcolor2[315]);
    BiasedRNG[580] = (LFSRcolor2[106]&LFSRcolor2[324]&LFSRcolor2[298]&LFSRcolor2[53]);
    BiasedRNG[581] = (LFSRcolor2[880]&LFSRcolor2[716]&LFSRcolor2[468]&LFSRcolor2[531]);
    BiasedRNG[582] = (LFSRcolor2[804]&LFSRcolor2[97]&LFSRcolor2[423]&LFSRcolor2[86]);
    BiasedRNG[583] = (LFSRcolor2[184]&LFSRcolor2[273]&LFSRcolor2[733]&LFSRcolor2[890]);
    BiasedRNG[584] = (LFSRcolor2[619]&LFSRcolor2[872]&LFSRcolor2[911]&LFSRcolor2[553]);
    BiasedRNG[585] = (LFSRcolor2[145]&LFSRcolor2[201]&LFSRcolor2[108]&LFSRcolor2[577]);
    BiasedRNG[586] = (LFSRcolor2[473]&LFSRcolor2[629]&LFSRcolor2[501]&LFSRcolor2[661]);
    BiasedRNG[587] = (LFSRcolor2[2]&LFSRcolor2[211]&LFSRcolor2[431]&LFSRcolor2[909]);
    BiasedRNG[588] = (LFSRcolor2[616]&LFSRcolor2[352]&LFSRcolor2[54]&LFSRcolor2[416]);
    BiasedRNG[589] = (LFSRcolor2[452]&LFSRcolor2[875]&LFSRcolor2[615]&LFSRcolor2[955]);
    BiasedRNG[590] = (LFSRcolor2[566]&LFSRcolor2[440]&LFSRcolor2[842]&LFSRcolor2[952]);
    BiasedRNG[591] = (LFSRcolor2[448]&LFSRcolor2[802]&LFSRcolor2[621]&LFSRcolor2[115]);
    BiasedRNG[592] = (LFSRcolor2[768]&LFSRcolor2[205]&LFSRcolor2[545]&LFSRcolor2[863]);
    BiasedRNG[593] = (LFSRcolor2[220]&LFSRcolor2[757]&LFSRcolor2[871]&LFSRcolor2[158]);
    BiasedRNG[594] = (LFSRcolor2[758]&LFSRcolor2[55]&LFSRcolor2[613]&LFSRcolor2[401]);
    BiasedRNG[595] = (LFSRcolor2[950]&LFSRcolor2[348]&LFSRcolor2[478]&LFSRcolor2[498]);
    BiasedRNG[596] = (LFSRcolor2[688]&LFSRcolor2[386]&LFSRcolor2[309]&LFSRcolor2[506]);
    BiasedRNG[597] = (LFSRcolor2[56]&LFSRcolor2[14]&LFSRcolor2[64]&LFSRcolor2[303]);
    BiasedRNG[598] = (LFSRcolor2[361]&LFSRcolor2[52]&LFSRcolor2[47]&LFSRcolor2[27]);
    BiasedRNG[599] = (LFSRcolor2[848]&LFSRcolor2[540]&LFSRcolor2[743]&LFSRcolor2[956]);
    BiasedRNG[600] = (LFSRcolor2[599]&LFSRcolor2[33]&LFSRcolor2[785]&LFSRcolor2[617]);
    BiasedRNG[601] = (LFSRcolor2[886]&LFSRcolor2[824]&LFSRcolor2[937]&LFSRcolor2[690]);
    BiasedRNG[602] = (LFSRcolor2[885]&LFSRcolor2[655]&LFSRcolor2[279]&LFSRcolor2[83]);
    BiasedRNG[603] = (LFSRcolor2[713]&LFSRcolor2[252]&LFSRcolor2[154]&LFSRcolor2[141]);
    BiasedRNG[604] = (LFSRcolor2[774]&LFSRcolor2[741]&LFSRcolor2[293]&LFSRcolor2[337]);
    BiasedRNG[605] = (LFSRcolor2[814]&LFSRcolor2[456]&LFSRcolor2[657]&LFSRcolor2[663]);
    BiasedRNG[606] = (LFSRcolor2[803]&LFSRcolor2[514]&LFSRcolor2[822]&LFSRcolor2[884]);
    BiasedRNG[607] = (LFSRcolor2[320]&LFSRcolor2[818]&LFSRcolor2[857]&LFSRcolor2[767]);
    BiasedRNG[608] = (LFSRcolor2[157]&LFSRcolor2[483]&LFSRcolor2[434]&LFSRcolor2[207]);
    BiasedRNG[609] = (LFSRcolor2[127]&LFSRcolor2[461]&LFSRcolor2[296]&LFSRcolor2[459]);
    BiasedRNG[610] = (LFSRcolor2[282]&LFSRcolor2[537]&LFSRcolor2[277]&LFSRcolor2[485]);
    BiasedRNG[611] = (LFSRcolor2[727]&LFSRcolor2[682]&LFSRcolor2[248]&LFSRcolor2[751]);
    BiasedRNG[612] = (LFSRcolor2[301]&LFSRcolor2[134]&LFSRcolor2[250]&LFSRcolor2[556]);
    BiasedRNG[613] = (LFSRcolor2[445]&LFSRcolor2[607]&LFSRcolor2[959]&LFSRcolor2[826]);
    BiasedRNG[614] = (LFSRcolor2[858]&LFSRcolor2[225]&LFSRcolor2[149]&LFSRcolor2[670]);
    BiasedRNG[615] = (LFSRcolor2[719]&LFSRcolor2[51]&LFSRcolor2[614]&LFSRcolor2[645]);
    BiasedRNG[616] = (LFSRcolor2[381]&LFSRcolor2[633]&LFSRcolor2[140]&LFSRcolor2[465]);
    BiasedRNG[617] = (LFSRcolor2[364]&LFSRcolor2[592]&LFSRcolor2[161]&LFSRcolor2[754]);
    BiasedRNG[618] = (LFSRcolor2[923]&LFSRcolor2[482]&LFSRcolor2[458]&LFSRcolor2[671]);
    BiasedRNG[619] = (LFSRcolor2[711]&LFSRcolor2[948]&LFSRcolor2[797]&LFSRcolor2[439]);
    BiasedRNG[620] = (LFSRcolor2[726]&LFSRcolor2[0]&LFSRcolor2[855]&LFSRcolor2[266]);
    BiasedRNG[621] = (LFSRcolor2[712]&LFSRcolor2[509]&LFSRcolor2[261]&LFSRcolor2[334]);
    BiasedRNG[622] = (LFSRcolor2[245]&LFSRcolor2[369]&LFSRcolor2[70]&LFSRcolor2[832]);
    BiasedRNG[623] = (LFSRcolor2[942]&LFSRcolor2[121]&LFSRcolor2[591]&LFSRcolor2[341]);
    BiasedRNG[624] = (LFSRcolor2[330]&LFSRcolor2[181]&LFSRcolor2[776]&LFSRcolor2[105]);
    BiasedRNG[625] = (LFSRcolor2[941]&LFSRcolor2[771]&LFSRcolor2[168]&LFSRcolor2[87]);
    BiasedRNG[626] = (LFSRcolor2[37]&LFSRcolor2[878]&LFSRcolor2[606]&LFSRcolor2[76]);
    BiasedRNG[627] = (LFSRcolor2[191]&LFSRcolor2[263]&LFSRcolor2[628]&LFSRcolor2[319]);
    BiasedRNG[628] = (LFSRcolor2[256]&LFSRcolor2[508]&LFSRcolor2[692]&LFSRcolor2[102]);
    BiasedRNG[629] = (LFSRcolor2[732]&LFSRcolor2[253]&LFSRcolor2[696]&LFSRcolor2[856]);
    BiasedRNG[630] = (LFSRcolor2[773]&LFSRcolor2[454]&LFSRcolor2[217]&LFSRcolor2[764]);
    BiasedRNG[631] = (LFSRcolor2[499]&LFSRcolor2[808]&LFSRcolor2[830]&LFSRcolor2[939]);
    BiasedRNG[632] = (LFSRcolor2[15]&LFSRcolor2[133]&LFSRcolor2[208]&LFSRcolor2[630]);
    BiasedRNG[633] = (LFSRcolor2[233]&LFSRcolor2[280]&LFSRcolor2[828]&LFSRcolor2[641]);
    BiasedRNG[634] = (LFSRcolor2[742]&LFSRcolor2[23]&LFSRcolor2[780]&LFSRcolor2[237]);
    BiasedRNG[635] = (LFSRcolor2[481]&LFSRcolor2[746]&LFSRcolor2[867]&LFSRcolor2[194]);
    BiasedRNG[636] = (LFSRcolor2[528]&LFSRcolor2[612]&LFSRcolor2[469]&LFSRcolor2[572]);
    BiasedRNG[637] = (LFSRcolor2[472]&LFSRcolor2[444]&LFSRcolor2[410]&LFSRcolor2[239]);
    BiasedRNG[638] = (LFSRcolor2[694]&LFSRcolor2[940]&LFSRcolor2[292]&LFSRcolor2[342]);
    BiasedRNG[639] = (LFSRcolor2[759]&LFSRcolor2[383]&LFSRcolor2[664]&LFSRcolor2[428]);
    BiasedRNG[640] = (LFSRcolor2[112]&LFSRcolor2[209]&LFSRcolor2[753]&LFSRcolor2[949]);
    BiasedRNG[641] = (LFSRcolor2[146]&LFSRcolor2[809]&LFSRcolor2[418]&LFSRcolor2[11]);
    BiasedRNG[642] = (LFSRcolor2[426]&LFSRcolor2[329]&LFSRcolor2[644]&LFSRcolor2[464]);
    BiasedRNG[643] = (LFSRcolor2[189]&LFSRcolor2[350]&LFSRcolor2[61]&LFSRcolor2[474]);
    BiasedRNG[644] = (LFSRcolor2[160]&LFSRcolor2[604]&LFSRcolor2[147]&LFSRcolor2[16]);
    BiasedRNG[645] = (LFSRcolor2[516]&LFSRcolor2[174]&LFSRcolor2[760]&LFSRcolor2[336]);
    BiasedRNG[646] = (LFSRcolor2[278]&LFSRcolor2[224]&LFSRcolor2[881]&LFSRcolor2[799]);
    BiasedRNG[647] = (LFSRcolor2[823]&LFSRcolor2[642]&LFSRcolor2[411]&LFSRcolor2[843]);
    BiasedRNG[648] = (LFSRcolor2[723]&LFSRcolor2[539]&LFSRcolor2[259]&LFSRcolor2[340]);
    BiasedRNG[649] = (LFSRcolor2[10]&LFSRcolor2[906]&LFSRcolor2[849]&LFSRcolor2[548]);
    BiasedRNG[650] = (LFSRcolor2[920]&LFSRcolor2[314]&LFSRcolor2[894]&LFSRcolor2[587]);
    BiasedRNG[651] = (LFSRcolor2[491]&LFSRcolor2[390]&LFSRcolor2[637]&LFSRcolor2[887]);
    BiasedRNG[652] = (LFSRcolor2[877]&LFSRcolor2[68]&LFSRcolor2[668]&LFSRcolor2[305]);
    BiasedRNG[653] = (LFSRcolor2[840]&LFSRcolor2[190]&LFSRcolor2[186]&LFSRcolor2[424]);
    BiasedRNG[654] = (LFSRcolor2[339]&LFSRcolor2[494]&LFSRcolor2[772]&LFSRcolor2[821]);
    BiasedRNG[655] = (LFSRcolor2[667]&LFSRcolor2[122]&LFSRcolor2[647]&LFSRcolor2[264]);
    BiasedRNG[656] = (LFSRcolor2[782]&LFSRcolor2[589]&LFSRcolor2[486]&LFSRcolor2[246]);
    BiasedRNG[657] = (LFSRcolor2[608]&LFSRcolor2[274]&LFSRcolor2[151]&LFSRcolor2[192]);
    BiasedRNG[658] = (LFSRcolor2[675]&LFSRcolor2[925]&LFSRcolor2[172]&LFSRcolor2[551]);
    BiasedRNG[659] = (LFSRcolor2[763]&LFSRcolor2[129]&LFSRcolor2[793]&LFSRcolor2[831]);
    BiasedRNG[660] = (LFSRcolor2[156]&LFSRcolor2[372]&LFSRcolor2[32]&LFSRcolor2[846]);
    BiasedRNG[661] = (LFSRcolor2[502]&LFSRcolor2[358]&LFSRcolor2[317]&LFSRcolor2[603]);
    BiasedRNG[662] = (LFSRcolor2[447]&LFSRcolor2[91]&LFSRcolor2[962]&LFSRcolor2[427]);
    BiasedRNG[663] = (LFSRcolor2[643]&LFSRcolor2[399]&LFSRcolor2[110]&LFSRcolor2[801]);
    BiasedRNG[664] = (LFSRcolor2[638]&LFSRcolor2[543]&LFSRcolor2[679]&LFSRcolor2[730]);
    BiasedRNG[665] = (LFSRcolor2[451]&LFSRcolor2[837]&LFSRcolor2[701]&LFSRcolor2[844]);
    BiasedRNG[666] = (LFSRcolor2[834]&LFSRcolor2[351]&LFSRcolor2[874]&LFSRcolor2[882]);
    BiasedRNG[667] = (LFSRcolor2[338]&LFSRcolor2[610]&LFSRcolor2[625]&LFSRcolor2[457]);
    BiasedRNG[668] = (LFSRcolor2[735]&LFSRcolor2[142]&LFSRcolor2[493]&LFSRcolor2[534]);
    BiasedRNG[669] = (LFSRcolor2[574]&LFSRcolor2[900]&LFSRcolor2[307]&LFSRcolor2[722]);
    BiasedRNG[670] = (LFSRcolor2[699]&LFSRcolor2[707]&LFSRcolor2[123]&LFSRcolor2[721]);
    BiasedRNG[671] = (LFSRcolor2[511]&LFSRcolor2[552]&LFSRcolor2[680]&LFSRcolor2[128]);
    BiasedRNG[672] = (LFSRcolor2[622]&LFSRcolor2[779]&LFSRcolor2[316]&LFSRcolor2[961]);
    BiasedRNG[673] = (LFSRcolor2[870]&LFSRcolor2[104]&LFSRcolor2[331]&LFSRcolor2[63]);
    BiasedRNG[674] = (LFSRcolor2[943]&LFSRcolor2[77]&LFSRcolor2[71]&LFSRcolor2[584]);
    BiasedRNG[675] = (LFSRcolor2[249]&LFSRcolor2[517]&LFSRcolor2[238]&LFSRcolor2[555]);
    BiasedRNG[676] = (LFSRcolor2[953]&LFSRcolor2[88]&LFSRcolor2[618]&LFSRcolor2[571]);
    BiasedRNG[677] = (LFSRcolor2[396]&LFSRcolor2[904]&LFSRcolor2[636]&LFSRcolor2[355]);
    BiasedRNG[678] = (LFSRcolor2[113]&LFSRcolor2[379]&LFSRcolor2[125]&LFSRcolor2[389]);
    BiasedRNG[679] = (LFSRcolor2[406]&LFSRcolor2[744]&LFSRcolor2[34]&LFSRcolor2[507]);
    BiasedRNG[680] = (LFSRcolor2[598]&LFSRcolor2[586]&LFSRcolor2[135]&LFSRcolor2[946]);
    BiasedRNG[681] = (LFSRcolor2[176]&LFSRcolor2[179]&LFSRcolor2[57]&LFSRcolor2[103]);
    BiasedRNG[682] = (LFSRcolor2[924]&LFSRcolor2[234]&LFSRcolor2[541]&LFSRcolor2[792]);
    BiasedRNG[683] = (LFSRcolor2[788]&LFSRcolor2[684]&LFSRcolor2[794]&LFSRcolor2[601]);
    BiasedRNG[684] = (LFSRcolor2[136]&LFSRcolor2[344]&LFSRcolor2[533]&LFSRcolor2[204]);
    BiasedRNG[685] = (LFSRcolor2[490]&LFSRcolor2[839]&LFSRcolor2[236]&LFSRcolor2[438]);
    BiasedRNG[686] = (LFSRcolor2[6]&LFSRcolor2[235]&LFSRcolor2[752]&LFSRcolor2[82]);
    BiasedRNG[687] = (LFSRcolor2[756]&LFSRcolor2[479]&LFSRcolor2[332]&LFSRcolor2[210]);
    BiasedRNG[688] = (LFSRcolor2[433]&LFSRcolor2[594]&LFSRcolor2[724]&LFSRcolor2[284]);
    BiasedRNG[689] = (LFSRcolor2[84]&LFSRcolor2[796]&LFSRcolor2[196]&LFSRcolor2[257]);
    BiasedRNG[690] = (LFSRcolor2[686]&LFSRcolor2[287]&LFSRcolor2[912]&LFSRcolor2[195]);
    BiasedRNG[691] = (LFSRcolor2[388]&LFSRcolor2[549]&LFSRcolor2[441]&LFSRcolor2[897]);
    BiasedRNG[692] = (LFSRcolor2[704]&LFSRcolor2[31]&LFSRcolor2[462]&LFSRcolor2[5]);
    BiasedRNG[693] = (LFSRcolor2[119]&LFSRcolor2[425]&LFSRcolor2[360]&LFSRcolor2[581]);
    BiasedRNG[694] = (LFSRcolor2[681]&LFSRcolor2[126]&LFSRcolor2[903]&LFSRcolor2[717]);
    BiasedRNG[695] = (LFSRcolor2[960]&LFSRcolor2[898]&LFSRcolor2[384]&LFSRcolor2[28]);
    BiasedRNG[696] = (LFSRcolor2[36]&LFSRcolor2[755]&LFSRcolor2[421]&LFSRcolor2[199]);
    BiasedRNG[697] = (LFSRcolor2[178]&LFSRcolor2[738]&LFSRcolor2[165]&LFSRcolor2[529]);
    BiasedRNG[698] = (LFSRcolor2[728]&LFSRcolor2[308]&LFSRcolor2[536]&LFSRcolor2[761]);
    UnbiasedRNG[386] = LFSRcolor2[640];
    UnbiasedRNG[387] = LFSRcolor2[646];
    UnbiasedRNG[388] = LFSRcolor2[954];
    UnbiasedRNG[389] = LFSRcolor2[860];
    UnbiasedRNG[390] = LFSRcolor2[50];
    UnbiasedRNG[391] = LFSRcolor2[745];
    UnbiasedRNG[392] = LFSRcolor2[889];
    UnbiasedRNG[393] = LFSRcolor2[255];
    UnbiasedRNG[394] = LFSRcolor2[3];
    UnbiasedRNG[395] = LFSRcolor2[827];
    UnbiasedRNG[396] = LFSRcolor2[322];
    UnbiasedRNG[397] = LFSRcolor2[267];
    UnbiasedRNG[398] = LFSRcolor2[442];
    UnbiasedRNG[399] = LFSRcolor2[865];
    UnbiasedRNG[400] = LFSRcolor2[118];
    UnbiasedRNG[401] = LFSRcolor2[377];
    UnbiasedRNG[402] = LFSRcolor2[654];
    UnbiasedRNG[403] = LFSRcolor2[652];
    UnbiasedRNG[404] = LFSRcolor2[935];
    UnbiasedRNG[405] = LFSRcolor2[693];
    UnbiasedRNG[406] = LFSRcolor2[687];
    UnbiasedRNG[407] = LFSRcolor2[789];
    UnbiasedRNG[408] = LFSRcolor2[524];
    UnbiasedRNG[409] = LFSRcolor2[703];
    UnbiasedRNG[410] = LFSRcolor2[554];
    UnbiasedRNG[411] = LFSRcolor2[164];
    UnbiasedRNG[412] = LFSRcolor2[564];
    UnbiasedRNG[413] = LFSRcolor2[700];
    UnbiasedRNG[414] = LFSRcolor2[945];
    UnbiasedRNG[415] = LFSRcolor2[29];
    UnbiasedRNG[416] = LFSRcolor2[138];
    UnbiasedRNG[417] = LFSRcolor2[492];
    UnbiasedRNG[418] = LFSRcolor2[373];
    UnbiasedRNG[419] = LFSRcolor2[356];
    UnbiasedRNG[420] = LFSRcolor2[437];
    UnbiasedRNG[421] = LFSRcolor2[674];
    UnbiasedRNG[422] = LFSRcolor2[739];
    UnbiasedRNG[423] = LFSRcolor2[376];
    UnbiasedRNG[424] = LFSRcolor2[89];
    UnbiasedRNG[425] = LFSRcolor2[304];
    UnbiasedRNG[426] = LFSRcolor2[163];
    UnbiasedRNG[427] = LFSRcolor2[169];
    UnbiasedRNG[428] = LFSRcolor2[928];
    UnbiasedRNG[429] = LFSRcolor2[380];
    UnbiasedRNG[430] = LFSRcolor2[150];
    UnbiasedRNG[431] = LFSRcolor2[73];
    UnbiasedRNG[432] = LFSRcolor2[265];
    UnbiasedRNG[433] = LFSRcolor2[677];
    UnbiasedRNG[434] = LFSRcolor2[888];
    UnbiasedRNG[435] = LFSRcolor2[378];
    UnbiasedRNG[436] = LFSRcolor2[98];
    UnbiasedRNG[437] = LFSRcolor2[183];
    UnbiasedRNG[438] = LFSRcolor2[155];
    UnbiasedRNG[439] = LFSRcolor2[306];
    UnbiasedRNG[440] = LFSRcolor2[525];
    UnbiasedRNG[441] = LFSRcolor2[902];
    UnbiasedRNG[442] = LFSRcolor2[951];
    UnbiasedRNG[443] = LFSRcolor2[99];
    UnbiasedRNG[444] = LFSRcolor2[609];
    UnbiasedRNG[445] = LFSRcolor2[913];
    UnbiasedRNG[446] = LFSRcolor2[39];
    UnbiasedRNG[447] = LFSRcolor2[436];
    UnbiasedRNG[448] = LFSRcolor2[930];
    UnbiasedRNG[449] = LFSRcolor2[206];
    UnbiasedRNG[450] = LFSRcolor2[567];
    UnbiasedRNG[451] = LFSRcolor2[409];
    UnbiasedRNG[452] = LFSRcolor2[676];
    UnbiasedRNG[453] = LFSRcolor2[400];
    UnbiasedRNG[454] = LFSRcolor2[368];
    UnbiasedRNG[455] = LFSRcolor2[382];
    UnbiasedRNG[456] = LFSRcolor2[291];
    UnbiasedRNG[457] = LFSRcolor2[258];
    UnbiasedRNG[458] = LFSRcolor2[18];
    UnbiasedRNG[459] = LFSRcolor2[470];
    UnbiasedRNG[460] = LFSRcolor2[24];
    UnbiasedRNG[461] = LFSRcolor2[120];
    UnbiasedRNG[462] = LFSRcolor2[859];
    UnbiasedRNG[463] = LFSRcolor2[868];
    UnbiasedRNG[464] = LFSRcolor2[836];
    UnbiasedRNG[465] = LFSRcolor2[854];
    UnbiasedRNG[466] = LFSRcolor2[866];
    UnbiasedRNG[467] = LFSRcolor2[232];
    UnbiasedRNG[468] = LFSRcolor2[769];
    UnbiasedRNG[469] = LFSRcolor2[69];
    UnbiasedRNG[470] = LFSRcolor2[43];
    UnbiasedRNG[471] = LFSRcolor2[805];
    UnbiasedRNG[472] = LFSRcolor2[593];
    UnbiasedRNG[473] = LFSRcolor2[602];
    UnbiasedRNG[474] = LFSRcolor2[212];
    UnbiasedRNG[475] = LFSRcolor2[270];
    UnbiasedRNG[476] = LFSRcolor2[819];
    UnbiasedRNG[477] = LFSRcolor2[268];
    UnbiasedRNG[478] = LFSRcolor2[26];
    UnbiasedRNG[479] = LFSRcolor2[398];
    UnbiasedRNG[480] = LFSRcolor2[166];
    UnbiasedRNG[481] = LFSRcolor2[455];
    UnbiasedRNG[482] = LFSRcolor2[476];
    UnbiasedRNG[483] = LFSRcolor2[892];
    UnbiasedRNG[484] = LFSRcolor2[783];
    UnbiasedRNG[485] = LFSRcolor2[153];
    UnbiasedRNG[486] = LFSRcolor2[272];
    UnbiasedRNG[487] = LFSRcolor2[513];
    UnbiasedRNG[488] = LFSRcolor2[124];
    UnbiasedRNG[489] = LFSRcolor2[575];
    UnbiasedRNG[490] = LFSRcolor2[392];
    UnbiasedRNG[491] = LFSRcolor2[111];
    UnbiasedRNG[492] = LFSRcolor2[835];
    UnbiasedRNG[493] = LFSRcolor2[130];
    UnbiasedRNG[494] = LFSRcolor2[42];
    UnbiasedRNG[495] = LFSRcolor2[747];
    UnbiasedRNG[496] = LFSRcolor2[230];
    UnbiasedRNG[497] = LFSRcolor2[394];
    UnbiasedRNG[498] = LFSRcolor2[740];
    UnbiasedRNG[499] = LFSRcolor2[412];
    UnbiasedRNG[500] = LFSRcolor2[708];
    UnbiasedRNG[501] = LFSRcolor2[262];
    UnbiasedRNG[502] = LFSRcolor2[173];
    UnbiasedRNG[503] = LFSRcolor2[915];
    UnbiasedRNG[504] = LFSRcolor2[689];
    UnbiasedRNG[505] = LFSRcolor2[557];
    UnbiasedRNG[506] = LFSRcolor2[660];
    UnbiasedRNG[507] = LFSRcolor2[200];
    UnbiasedRNG[508] = LFSRcolor2[810];
    UnbiasedRNG[509] = LFSRcolor2[795];
    UnbiasedRNG[510] = LFSRcolor2[17];
    UnbiasedRNG[511] = LFSRcolor2[901];
    UnbiasedRNG[512] = LFSRcolor2[326];
    UnbiasedRNG[513] = LFSRcolor2[285];
    UnbiasedRNG[514] = LFSRcolor2[241];
    UnbiasedRNG[515] = LFSRcolor2[927];
    UnbiasedRNG[516] = LFSRcolor2[933];
    UnbiasedRNG[517] = LFSRcolor2[791];
    UnbiasedRNG[518] = LFSRcolor2[354];
    UnbiasedRNG[519] = LFSRcolor2[648];
    UnbiasedRNG[520] = LFSRcolor2[271];
    UnbiasedRNG[521] = LFSRcolor2[30];
    UnbiasedRNG[522] = LFSRcolor2[563];
    UnbiasedRNG[523] = LFSRcolor2[798];
    UnbiasedRNG[524] = LFSRcolor2[817];
    UnbiasedRNG[525] = LFSRcolor2[570];
    UnbiasedRNG[526] = LFSRcolor2[325];
    UnbiasedRNG[527] = LFSRcolor2[649];
    UnbiasedRNG[528] = LFSRcolor2[825];
    UnbiasedRNG[529] = LFSRcolor2[85];
    UnbiasedRNG[530] = LFSRcolor2[666];
    UnbiasedRNG[531] = LFSRcolor2[515];
    UnbiasedRNG[532] = LFSRcolor2[13];
    UnbiasedRNG[533] = LFSRcolor2[74];
    UnbiasedRNG[534] = LFSRcolor2[569];
    UnbiasedRNG[535] = LFSRcolor2[175];
    UnbiasedRNG[536] = LFSRcolor2[420];
    UnbiasedRNG[537] = LFSRcolor2[417];
    UnbiasedRNG[538] = LFSRcolor2[407];
    UnbiasedRNG[539] = LFSRcolor2[714];
    UnbiasedRNG[540] = LFSRcolor2[811];
    UnbiasedRNG[541] = LFSRcolor2[876];
    UnbiasedRNG[542] = LFSRcolor2[965];
    UnbiasedRNG[543] = LFSRcolor2[565];
    UnbiasedRNG[544] = LFSRcolor2[521];
    UnbiasedRNG[545] = LFSRcolor2[899];
    UnbiasedRNG[546] = LFSRcolor2[371];
    UnbiasedRNG[547] = LFSRcolor2[815];
    UnbiasedRNG[548] = LFSRcolor2[290];
    UnbiasedRNG[549] = LFSRcolor2[397];
    UnbiasedRNG[550] = LFSRcolor2[518];
    UnbiasedRNG[551] = LFSRcolor2[958];
    UnbiasedRNG[552] = LFSRcolor2[58];
    UnbiasedRNG[553] = LFSRcolor2[673];
    UnbiasedRNG[554] = LFSRcolor2[218];
    UnbiasedRNG[555] = LFSRcolor2[922];
    UnbiasedRNG[556] = LFSRcolor2[357];
    UnbiasedRNG[557] = LFSRcolor2[683];
    UnbiasedRNG[558] = LFSRcolor2[393];
    UnbiasedRNG[559] = LFSRcolor2[691];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[560] = LFSRcolor3[181];
    UnbiasedRNG[561] = LFSRcolor3[52];
    UnbiasedRNG[562] = LFSRcolor3[72];
    UnbiasedRNG[563] = LFSRcolor3[179];
    UnbiasedRNG[564] = LFSRcolor3[67];
    UnbiasedRNG[565] = LFSRcolor3[73];
    UnbiasedRNG[566] = LFSRcolor3[119];
    UnbiasedRNG[567] = LFSRcolor3[160];
    UnbiasedRNG[568] = LFSRcolor3[112];
    UnbiasedRNG[569] = LFSRcolor3[8];
    UnbiasedRNG[570] = LFSRcolor3[25];
    UnbiasedRNG[571] = LFSRcolor3[77];
    UnbiasedRNG[572] = LFSRcolor3[138];
    UnbiasedRNG[573] = LFSRcolor3[50];
    UnbiasedRNG[574] = LFSRcolor3[123];
    UnbiasedRNG[575] = LFSRcolor3[90];
    UnbiasedRNG[576] = LFSRcolor3[163];
    UnbiasedRNG[577] = LFSRcolor3[58];
    UnbiasedRNG[578] = LFSRcolor3[86];
    UnbiasedRNG[579] = LFSRcolor3[13];
    UnbiasedRNG[580] = LFSRcolor3[131];
    UnbiasedRNG[581] = LFSRcolor3[99];
    UnbiasedRNG[582] = LFSRcolor3[155];
    UnbiasedRNG[583] = LFSRcolor3[41];
    UnbiasedRNG[584] = LFSRcolor3[165];
    UnbiasedRNG[585] = LFSRcolor3[92];
    UnbiasedRNG[586] = LFSRcolor3[122];
    UnbiasedRNG[587] = LFSRcolor3[48];
    UnbiasedRNG[588] = LFSRcolor3[148];
    UnbiasedRNG[589] = LFSRcolor3[100];
    UnbiasedRNG[590] = LFSRcolor3[101];
    UnbiasedRNG[591] = LFSRcolor3[115];
    UnbiasedRNG[592] = LFSRcolor3[87];
    UnbiasedRNG[593] = LFSRcolor3[95];
    UnbiasedRNG[594] = LFSRcolor3[59];
    UnbiasedRNG[595] = LFSRcolor3[121];
    UnbiasedRNG[596] = LFSRcolor3[140];
    UnbiasedRNG[597] = LFSRcolor3[117];
    UnbiasedRNG[598] = LFSRcolor3[16];
    UnbiasedRNG[599] = LFSRcolor3[142];
    UnbiasedRNG[600] = LFSRcolor3[169];
    UnbiasedRNG[601] = LFSRcolor3[27];
    UnbiasedRNG[602] = LFSRcolor3[45];
    UnbiasedRNG[603] = LFSRcolor3[109];
    UnbiasedRNG[604] = LFSRcolor3[137];
    UnbiasedRNG[605] = LFSRcolor3[103];
    UnbiasedRNG[606] = LFSRcolor3[128];
    UnbiasedRNG[607] = LFSRcolor3[180];
    UnbiasedRNG[608] = LFSRcolor3[150];
    UnbiasedRNG[609] = LFSRcolor3[66];
    UnbiasedRNG[610] = LFSRcolor3[154];
    UnbiasedRNG[611] = LFSRcolor3[91];
    UnbiasedRNG[612] = LFSRcolor3[113];
    UnbiasedRNG[613] = LFSRcolor3[170];
    UnbiasedRNG[614] = LFSRcolor3[108];
    UnbiasedRNG[615] = LFSRcolor3[102];
    UnbiasedRNG[616] = LFSRcolor3[30];
    UnbiasedRNG[617] = LFSRcolor3[85];
    UnbiasedRNG[618] = LFSRcolor3[146];
    UnbiasedRNG[619] = LFSRcolor3[141];
    UnbiasedRNG[620] = LFSRcolor3[98];
    UnbiasedRNG[621] = LFSRcolor3[152];
    UnbiasedRNG[622] = LFSRcolor3[54];
    UnbiasedRNG[623] = LFSRcolor3[20];
    UnbiasedRNG[624] = LFSRcolor3[133];
    UnbiasedRNG[625] = LFSRcolor3[147];
    UnbiasedRNG[626] = LFSRcolor3[105];
    UnbiasedRNG[627] = LFSRcolor3[183];
    UnbiasedRNG[628] = LFSRcolor3[166];
    UnbiasedRNG[629] = LFSRcolor3[29];
    UnbiasedRNG[630] = LFSRcolor3[82];
    UnbiasedRNG[631] = LFSRcolor3[47];
    UnbiasedRNG[632] = LFSRcolor3[173];
    UnbiasedRNG[633] = LFSRcolor3[158];
    UnbiasedRNG[634] = LFSRcolor3[56];
    UnbiasedRNG[635] = LFSRcolor3[74];
    UnbiasedRNG[636] = LFSRcolor3[11];
    UnbiasedRNG[637] = LFSRcolor3[65];
    UnbiasedRNG[638] = LFSRcolor3[84];
    UnbiasedRNG[639] = LFSRcolor3[18];
    UnbiasedRNG[640] = LFSRcolor3[26];
    UnbiasedRNG[641] = LFSRcolor3[42];
    UnbiasedRNG[642] = LFSRcolor3[40];
    UnbiasedRNG[643] = LFSRcolor3[110];
    UnbiasedRNG[644] = LFSRcolor3[93];
    UnbiasedRNG[645] = LFSRcolor3[167];
    UnbiasedRNG[646] = LFSRcolor3[36];
    UnbiasedRNG[647] = LFSRcolor3[28];
    UnbiasedRNG[648] = LFSRcolor3[7];
    UnbiasedRNG[649] = LFSRcolor3[53];
    UnbiasedRNG[650] = LFSRcolor3[156];
    UnbiasedRNG[651] = LFSRcolor3[168];
    UnbiasedRNG[652] = LFSRcolor3[38];
    UnbiasedRNG[653] = LFSRcolor3[9];
    UnbiasedRNG[654] = LFSRcolor3[125];
    UnbiasedRNG[655] = LFSRcolor3[69];
    UnbiasedRNG[656] = LFSRcolor3[136];
    UnbiasedRNG[657] = LFSRcolor3[1];
    UnbiasedRNG[658] = LFSRcolor3[23];
    UnbiasedRNG[659] = LFSRcolor3[132];
    UnbiasedRNG[660] = LFSRcolor3[171];
    UnbiasedRNG[661] = LFSRcolor3[143];
    UnbiasedRNG[662] = LFSRcolor3[62];
    UnbiasedRNG[663] = LFSRcolor3[4];
    UnbiasedRNG[664] = LFSRcolor3[97];
    UnbiasedRNG[665] = LFSRcolor3[114];
    UnbiasedRNG[666] = LFSRcolor3[106];
    UnbiasedRNG[667] = LFSRcolor3[22];
    UnbiasedRNG[668] = LFSRcolor3[172];
    UnbiasedRNG[669] = LFSRcolor3[89];
    UnbiasedRNG[670] = LFSRcolor3[17];
    UnbiasedRNG[671] = LFSRcolor3[116];
    UnbiasedRNG[672] = LFSRcolor3[57];
    UnbiasedRNG[673] = LFSRcolor3[5];
    UnbiasedRNG[674] = LFSRcolor3[60];
    UnbiasedRNG[675] = LFSRcolor3[157];
    UnbiasedRNG[676] = LFSRcolor3[81];
    UnbiasedRNG[677] = LFSRcolor3[126];
    UnbiasedRNG[678] = LFSRcolor3[177];
    UnbiasedRNG[679] = LFSRcolor3[43];
    UnbiasedRNG[680] = LFSRcolor3[0];
    UnbiasedRNG[681] = LFSRcolor3[46];
    UnbiasedRNG[682] = LFSRcolor3[32];
    UnbiasedRNG[683] = LFSRcolor3[178];
    UnbiasedRNG[684] = LFSRcolor3[124];
    UnbiasedRNG[685] = LFSRcolor3[49];
    UnbiasedRNG[686] = LFSRcolor3[75];
    UnbiasedRNG[687] = LFSRcolor3[78];
    UnbiasedRNG[688] = LFSRcolor3[12];
    UnbiasedRNG[689] = LFSRcolor3[144];
    UnbiasedRNG[690] = LFSRcolor3[83];
    UnbiasedRNG[691] = LFSRcolor3[159];
    UnbiasedRNG[692] = LFSRcolor3[139];
    UnbiasedRNG[693] = LFSRcolor3[21];
    UnbiasedRNG[694] = LFSRcolor3[39];
    UnbiasedRNG[695] = LFSRcolor3[182];
    UnbiasedRNG[696] = LFSRcolor3[175];
    UnbiasedRNG[697] = LFSRcolor3[33];
    UnbiasedRNG[698] = LFSRcolor3[149];
    UnbiasedRNG[699] = LFSRcolor3[107];
    UnbiasedRNG[700] = LFSRcolor3[88];
    UnbiasedRNG[701] = LFSRcolor3[120];
    UnbiasedRNG[702] = LFSRcolor3[64];
    UnbiasedRNG[703] = LFSRcolor3[104];
    UnbiasedRNG[704] = LFSRcolor3[134];
    UnbiasedRNG[705] = LFSRcolor3[68];
    UnbiasedRNG[706] = LFSRcolor3[6];
    UnbiasedRNG[707] = LFSRcolor3[24];
    UnbiasedRNG[708] = LFSRcolor3[135];
    UnbiasedRNG[709] = LFSRcolor3[55];
    UnbiasedRNG[710] = LFSRcolor3[51];
    UnbiasedRNG[711] = LFSRcolor3[44];
    UnbiasedRNG[712] = LFSRcolor3[130];
    UnbiasedRNG[713] = LFSRcolor3[111];
    UnbiasedRNG[714] = LFSRcolor3[80];
    UnbiasedRNG[715] = LFSRcolor3[129];
end

always @(posedge color3_clk) begin
    BiasedRNG[699] = (LFSRcolor4[565]&LFSRcolor4[355]&LFSRcolor4[552]&LFSRcolor4[143]);
    BiasedRNG[700] = (LFSRcolor4[379]&LFSRcolor4[696]&LFSRcolor4[673]&LFSRcolor4[286]);
    BiasedRNG[701] = (LFSRcolor4[373]&LFSRcolor4[566]&LFSRcolor4[251]&LFSRcolor4[233]);
    BiasedRNG[702] = (LFSRcolor4[638]&LFSRcolor4[325]&LFSRcolor4[370]&LFSRcolor4[322]);
    BiasedRNG[703] = (LFSRcolor4[343]&LFSRcolor4[64]&LFSRcolor4[18]&LFSRcolor4[328]);
    BiasedRNG[704] = (LFSRcolor4[78]&LFSRcolor4[114]&LFSRcolor4[241]&LFSRcolor4[734]);
    BiasedRNG[705] = (LFSRcolor4[530]&LFSRcolor4[96]&LFSRcolor4[634]&LFSRcolor4[48]);
    BiasedRNG[706] = (LFSRcolor4[319]&LFSRcolor4[177]&LFSRcolor4[641]&LFSRcolor4[37]);
    BiasedRNG[707] = (LFSRcolor4[452]&LFSRcolor4[60]&LFSRcolor4[400]&LFSRcolor4[548]);
    BiasedRNG[708] = (LFSRcolor4[213]&LFSRcolor4[396]&LFSRcolor4[75]&LFSRcolor4[682]);
    BiasedRNG[709] = (LFSRcolor4[165]&LFSRcolor4[722]&LFSRcolor4[480]&LFSRcolor4[395]);
    BiasedRNG[710] = (LFSRcolor4[365]&LFSRcolor4[523]&LFSRcolor4[637]&LFSRcolor4[372]);
    BiasedRNG[711] = (LFSRcolor4[600]&LFSRcolor4[147]&LFSRcolor4[31]&LFSRcolor4[290]);
    BiasedRNG[712] = (LFSRcolor4[567]&LFSRcolor4[270]&LFSRcolor4[598]&LFSRcolor4[304]);
    BiasedRNG[713] = (LFSRcolor4[464]&LFSRcolor4[446]&LFSRcolor4[525]&LFSRcolor4[9]);
    BiasedRNG[714] = (LFSRcolor4[606]&LFSRcolor4[594]&LFSRcolor4[675]&LFSRcolor4[592]);
    BiasedRNG[715] = (LFSRcolor4[735]&LFSRcolor4[698]&LFSRcolor4[426]&LFSRcolor4[133]);
    BiasedRNG[716] = (LFSRcolor4[482]&LFSRcolor4[429]&LFSRcolor4[701]&LFSRcolor4[403]);
    BiasedRNG[717] = (LFSRcolor4[170]&LFSRcolor4[351]&LFSRcolor4[148]&LFSRcolor4[691]);
    BiasedRNG[718] = (LFSRcolor4[616]&LFSRcolor4[444]&LFSRcolor4[115]&LFSRcolor4[484]);
    BiasedRNG[719] = (LFSRcolor4[625]&LFSRcolor4[498]&LFSRcolor4[221]&LFSRcolor4[236]);
    BiasedRNG[720] = (LFSRcolor4[128]&LFSRcolor4[601]&LFSRcolor4[469]&LFSRcolor4[225]);
    BiasedRNG[721] = (LFSRcolor4[680]&LFSRcolor4[724]&LFSRcolor4[88]&LFSRcolor4[551]);
    BiasedRNG[722] = (LFSRcolor4[65]&LFSRcolor4[36]&LFSRcolor4[714]&LFSRcolor4[561]);
    BiasedRNG[723] = (LFSRcolor4[649]&LFSRcolor4[553]&LFSRcolor4[399]&LFSRcolor4[67]);
    BiasedRNG[724] = (LFSRcolor4[635]&LFSRcolor4[222]&LFSRcolor4[347]&LFSRcolor4[175]);
    BiasedRNG[725] = (LFSRcolor4[99]&LFSRcolor4[292]&LFSRcolor4[66]&LFSRcolor4[423]);
    BiasedRNG[726] = (LFSRcolor4[49]&LFSRcolor4[22]&LFSRcolor4[459]&LFSRcolor4[575]);
    BiasedRNG[727] = (LFSRcolor4[214]&LFSRcolor4[334]&LFSRcolor4[652]&LFSRcolor4[136]);
    BiasedRNG[728] = (LFSRcolor4[310]&LFSRcolor4[371]&LFSRcolor4[55]&LFSRcolor4[492]);
    BiasedRNG[729] = (LFSRcolor4[367]&LFSRcolor4[458]&LFSRcolor4[103]&LFSRcolor4[534]);
    BiasedRNG[730] = (LFSRcolor4[257]&LFSRcolor4[242]&LFSRcolor4[437]&LFSRcolor4[585]);
    BiasedRNG[731] = (LFSRcolor4[248]&LFSRcolor4[249]&LFSRcolor4[234]&LFSRcolor4[260]);
    BiasedRNG[732] = (LFSRcolor4[188]&LFSRcolor4[359]&LFSRcolor4[411]&LFSRcolor4[685]);
    BiasedRNG[733] = (LFSRcolor4[59]&LFSRcolor4[700]&LFSRcolor4[382]&LFSRcolor4[481]);
    BiasedRNG[734] = (LFSRcolor4[718]&LFSRcolor4[172]&LFSRcolor4[406]&LFSRcolor4[483]);
    BiasedRNG[735] = (LFSRcolor4[211]&LFSRcolor4[666]&LFSRcolor4[667]&LFSRcolor4[267]);
    BiasedRNG[736] = (LFSRcolor4[279]&LFSRcolor4[421]&LFSRcolor4[563]&LFSRcolor4[58]);
    BiasedRNG[737] = (LFSRcolor4[644]&LFSRcolor4[79]&LFSRcolor4[564]&LFSRcolor4[72]);
    BiasedRNG[738] = (LFSRcolor4[107]&LFSRcolor4[204]&LFSRcolor4[179]&LFSRcolor4[116]);
    BiasedRNG[739] = (LFSRcolor4[721]&LFSRcolor4[576]&LFSRcolor4[521]&LFSRcolor4[187]);
    BiasedRNG[740] = (LFSRcolor4[2]&LFSRcolor4[124]&LFSRcolor4[300]&LFSRcolor4[81]);
    BiasedRNG[741] = (LFSRcolor4[475]&LFSRcolor4[610]&LFSRcolor4[160]&LFSRcolor4[53]);
    BiasedRNG[742] = (LFSRcolor4[393]&LFSRcolor4[456]&LFSRcolor4[380]&LFSRcolor4[486]);
    BiasedRNG[743] = (LFSRcolor4[268]&LFSRcolor4[418]&LFSRcolor4[320]&LFSRcolor4[584]);
    BiasedRNG[744] = (LFSRcolor4[419]&LFSRcolor4[569]&LFSRcolor4[608]&LFSRcolor4[568]);
    BiasedRNG[745] = (LFSRcolor4[369]&LFSRcolor4[683]&LFSRcolor4[298]&LFSRcolor4[368]);
    BiasedRNG[746] = (LFSRcolor4[195]&LFSRcolor4[583]&LFSRcolor4[476]&LFSRcolor4[23]);
    BiasedRNG[747] = (LFSRcolor4[25]&LFSRcolor4[388]&LFSRcolor4[16]&LFSRcolor4[163]);
    BiasedRNG[748] = (LFSRcolor4[274]&LFSRcolor4[436]&LFSRcolor4[89]&LFSRcolor4[4]);
    BiasedRNG[749] = (LFSRcolor4[636]&LFSRcolor4[604]&LFSRcolor4[424]&LFSRcolor4[428]);
    BiasedRNG[750] = (LFSRcolor4[439]&LFSRcolor4[11]&LFSRcolor4[206]&LFSRcolor4[408]);
    BiasedRNG[751] = (LFSRcolor4[40]&LFSRcolor4[330]&LFSRcolor4[176]&LFSRcolor4[264]);
    BiasedRNG[752] = (LFSRcolor4[282]&LFSRcolor4[231]&LFSRcolor4[285]&LFSRcolor4[515]);
    BiasedRNG[753] = (LFSRcolor4[398]&LFSRcolor4[599]&LFSRcolor4[445]&LFSRcolor4[173]);
    BiasedRNG[754] = (LFSRcolor4[291]&LFSRcolor4[385]&LFSRcolor4[357]&LFSRcolor4[517]);
    BiasedRNG[755] = (LFSRcolor4[500]&LFSRcolor4[478]&LFSRcolor4[202]&LFSRcolor4[725]);
    BiasedRNG[756] = (LFSRcolor4[412]&LFSRcolor4[117]&LFSRcolor4[348]&LFSRcolor4[485]);
    BiasedRNG[757] = (LFSRcolor4[581]&LFSRcolor4[27]&LFSRcolor4[3]&LFSRcolor4[197]);
    BiasedRNG[758] = (LFSRcolor4[146]&LFSRcolor4[528]&LFSRcolor4[615]&LFSRcolor4[390]);
    BiasedRNG[759] = (LFSRcolor4[12]&LFSRcolor4[127]&LFSRcolor4[702]&LFSRcolor4[0]);
    BiasedRNG[760] = (LFSRcolor4[326]&LFSRcolor4[559]&LFSRcolor4[296]&LFSRcolor4[681]);
    BiasedRNG[761] = (LFSRcolor4[230]&LFSRcolor4[461]&LFSRcolor4[654]&LFSRcolor4[121]);
    BiasedRNG[762] = (LFSRcolor4[438]&LFSRcolor4[74]&LFSRcolor4[502]&LFSRcolor4[684]);
    BiasedRNG[763] = (LFSRcolor4[134]&LFSRcolor4[589]&LFSRcolor4[465]&LFSRcolor4[180]);
    BiasedRNG[764] = (LFSRcolor4[674]&LFSRcolor4[162]&LFSRcolor4[582]&LFSRcolor4[76]);
    BiasedRNG[765] = (LFSRcolor4[468]&LFSRcolor4[317]&LFSRcolor4[715]&LFSRcolor4[470]);
    BiasedRNG[766] = (LFSRcolor4[658]&LFSRcolor4[207]&LFSRcolor4[572]&LFSRcolor4[405]);
    BiasedRNG[767] = (LFSRcolor4[97]&LFSRcolor4[100]&LFSRcolor4[556]&LFSRcolor4[98]);
    BiasedRNG[768] = (LFSRcolor4[453]&LFSRcolor4[87]&LFSRcolor4[588]&LFSRcolor4[297]);
    BiasedRNG[769] = (LFSRcolor4[352]&LFSRcolor4[535]&LFSRcolor4[137]&LFSRcolor4[30]);
    BiasedRNG[770] = (LFSRcolor4[686]&LFSRcolor4[276]&LFSRcolor4[497]&LFSRcolor4[20]);
    BiasedRNG[771] = (LFSRcolor4[295]&LFSRcolor4[256]&LFSRcolor4[273]&LFSRcolor4[110]);
    BiasedRNG[772] = (LFSRcolor4[460]&LFSRcolor4[194]&LFSRcolor4[672]&LFSRcolor4[178]);
    BiasedRNG[773] = (LFSRcolor4[32]&LFSRcolor4[693]&LFSRcolor4[104]&LFSRcolor4[159]);
    BiasedRNG[774] = (LFSRcolor4[191]&LFSRcolor4[259]&LFSRcolor4[245]&LFSRcolor4[156]);
    BiasedRNG[775] = (LFSRcolor4[655]&LFSRcolor4[663]&LFSRcolor4[474]&LFSRcolor4[183]);
    BiasedRNG[776] = (LFSRcolor4[41]&LFSRcolor4[47]&LFSRcolor4[547]&LFSRcolor4[210]);
    BiasedRNG[777] = (LFSRcolor4[171]&LFSRcolor4[669]&LFSRcolor4[494]&LFSRcolor4[537]);
    BiasedRNG[778] = (LFSRcolor4[85]&LFSRcolor4[612]&LFSRcolor4[263]&LFSRcolor4[730]);
    BiasedRNG[779] = (LFSRcolor4[21]&LFSRcolor4[512]&LFSRcolor4[374]&LFSRcolor4[450]);
    BiasedRNG[780] = (LFSRcolor4[192]&LFSRcolor4[624]&LFSRcolor4[154]&LFSRcolor4[299]);
    BiasedRNG[781] = (LFSRcolor4[209]&LFSRcolor4[294]&LFSRcolor4[653]&LFSRcolor4[414]);
    BiasedRNG[782] = (LFSRcolor4[253]&LFSRcolor4[284]&LFSRcolor4[350]&LFSRcolor4[316]);
    BiasedRNG[783] = (LFSRcolor4[410]&LFSRcolor4[224]&LFSRcolor4[45]&LFSRcolor4[473]);
    BiasedRNG[784] = (LFSRcolor4[323]&LFSRcolor4[327]&LFSRcolor4[135]&LFSRcolor4[643]);
    BiasedRNG[785] = (LFSRcolor4[269]&LFSRcolor4[455]&LFSRcolor4[590]&LFSRcolor4[511]);
    BiasedRNG[786] = (LFSRcolor4[471]&LFSRcolor4[454]&LFSRcolor4[70]&LFSRcolor4[558]);
    BiasedRNG[787] = (LFSRcolor4[315]&LFSRcolor4[540]&LFSRcolor4[8]&LFSRcolor4[544]);
    BiasedRNG[788] = (LFSRcolor4[630]&LFSRcolor4[657]&LFSRcolor4[93]&LFSRcolor4[626]);
    BiasedRNG[789] = (LFSRcolor4[167]&LFSRcolor4[198]&LFSRcolor4[308]&LFSRcolor4[490]);
    BiasedRNG[790] = (LFSRcolor4[605]&LFSRcolor4[441]&LFSRcolor4[442]&LFSRcolor4[587]);
    BiasedRNG[791] = (LFSRcolor4[13]&LFSRcolor4[506]&LFSRcolor4[420]&LFSRcolor4[168]);
    BiasedRNG[792] = (LFSRcolor4[609]&LFSRcolor4[536]&LFSRcolor4[150]&LFSRcolor4[151]);
    BiasedRNG[793] = (LFSRcolor4[695]&LFSRcolor4[218]&LFSRcolor4[337]&LFSRcolor4[189]);
    BiasedRNG[794] = (LFSRcolor4[522]&LFSRcolor4[705]&LFSRcolor4[247]&LFSRcolor4[280]);
    BiasedRNG[795] = (LFSRcolor4[220]&LFSRcolor4[434]&LFSRcolor4[240]&LFSRcolor4[223]);
    BiasedRNG[796] = (LFSRcolor4[340]&LFSRcolor4[613]&LFSRcolor4[34]&LFSRcolor4[694]);
    BiasedRNG[797] = (LFSRcolor4[24]&LFSRcolor4[622]&LFSRcolor4[250]&LFSRcolor4[278]);
    BiasedRNG[798] = (LFSRcolor4[467]&LFSRcolor4[707]&LFSRcolor4[621]&LFSRcolor4[560]);
    BiasedRNG[799] = (LFSRcolor4[35]&LFSRcolor4[313]&LFSRcolor4[662]&LFSRcolor4[112]);
    BiasedRNG[800] = (LFSRcolor4[541]&LFSRcolor4[728]&LFSRcolor4[462]&LFSRcolor4[447]);
    BiasedRNG[801] = (LFSRcolor4[90]&LFSRcolor4[538]&LFSRcolor4[432]&LFSRcolor4[733]);
    BiasedRNG[802] = (LFSRcolor4[309]&LFSRcolor4[157]&LFSRcolor4[384]&LFSRcolor4[692]);
    BiasedRNG[803] = (LFSRcolor4[266]&LFSRcolor4[697]&LFSRcolor4[356]&LFSRcolor4[201]);
    BiasedRNG[804] = (LFSRcolor4[43]&LFSRcolor4[125]&LFSRcolor4[443]&LFSRcolor4[519]);
    BiasedRNG[805] = (LFSRcolor4[332]&LFSRcolor4[129]&LFSRcolor4[10]&LFSRcolor4[226]);
    BiasedRNG[806] = (LFSRcolor4[578]&LFSRcolor4[91]&LFSRcolor4[346]&LFSRcolor4[311]);
    BiasedRNG[807] = (LFSRcolor4[574]&LFSRcolor4[533]&LFSRcolor4[407]&LFSRcolor4[149]);
    BiasedRNG[808] = (LFSRcolor4[174]&LFSRcolor4[417]&LFSRcolor4[61]&LFSRcolor4[628]);
    BiasedRNG[809] = (LFSRcolor4[50]&LFSRcolor4[394]&LFSRcolor4[26]&LFSRcolor4[83]);
    BiasedRNG[810] = (LFSRcolor4[56]&LFSRcolor4[397]&LFSRcolor4[329]&LFSRcolor4[381]);
    BiasedRNG[811] = (LFSRcolor4[562]&LFSRcolor4[678]&LFSRcolor4[262]&LFSRcolor4[573]);
    BiasedRNG[812] = (LFSRcolor4[451]&LFSRcolor4[113]&LFSRcolor4[401]&LFSRcolor4[472]);
    BiasedRNG[813] = (LFSRcolor4[647]&LFSRcolor4[496]&LFSRcolor4[277]&LFSRcolor4[688]);
    BiasedRNG[814] = (LFSRcolor4[489]&LFSRcolor4[513]&LFSRcolor4[161]&LFSRcolor4[595]);
    BiasedRNG[815] = (LFSRcolor4[306]&LFSRcolor4[668]&LFSRcolor4[677]&LFSRcolor4[440]);
    BiasedRNG[816] = (LFSRcolor4[169]&LFSRcolor4[690]&LFSRcolor4[314]&LFSRcolor4[554]);
    BiasedRNG[817] = (LFSRcolor4[729]&LFSRcolor4[664]&LFSRcolor4[131]&LFSRcolor4[363]);
    BiasedRNG[818] = (LFSRcolor4[670]&LFSRcolor4[618]&LFSRcolor4[46]&LFSRcolor4[122]);
    BiasedRNG[819] = (LFSRcolor4[504]&LFSRcolor4[166]&LFSRcolor4[660]&LFSRcolor4[5]);
    BiasedRNG[820] = (LFSRcolor4[518]&LFSRcolor4[620]&LFSRcolor4[69]&LFSRcolor4[181]);
    BiasedRNG[821] = (LFSRcolor4[52]&LFSRcolor4[193]&LFSRcolor4[708]&LFSRcolor4[203]);
    BiasedRNG[822] = (LFSRcolor4[435]&LFSRcolor4[501]&LFSRcolor4[243]&LFSRcolor4[237]);
    BiasedRNG[823] = (LFSRcolor4[336]&LFSRcolor4[699]&LFSRcolor4[244]&LFSRcolor4[510]);
    BiasedRNG[824] = (LFSRcolor4[550]&LFSRcolor4[466]&LFSRcolor4[524]&LFSRcolor4[366]);
    BiasedRNG[825] = (LFSRcolor4[255]&LFSRcolor4[331]&LFSRcolor4[338]&LFSRcolor4[703]);
    BiasedRNG[826] = (LFSRcolor4[717]&LFSRcolor4[709]&LFSRcolor4[57]&LFSRcolor4[318]);
    BiasedRNG[827] = (LFSRcolor4[409]&LFSRcolor4[415]&LFSRcolor4[15]&LFSRcolor4[487]);
    BiasedRNG[828] = (LFSRcolor4[145]&LFSRcolor4[427]&LFSRcolor4[305]&LFSRcolor4[182]);
    BiasedRNG[829] = (LFSRcolor4[84]&LFSRcolor4[503]&LFSRcolor4[42]&LFSRcolor4[650]);
    BiasedRNG[830] = (LFSRcolor4[593]&LFSRcolor4[579]&LFSRcolor4[391]&LFSRcolor4[158]);
    BiasedRNG[831] = (LFSRcolor4[520]&LFSRcolor4[542]&LFSRcolor4[596]&LFSRcolor4[252]);
    BiasedRNG[832] = (LFSRcolor4[586]&LFSRcolor4[1]&LFSRcolor4[102]&LFSRcolor4[153]);
    BiasedRNG[833] = (LFSRcolor4[293]&LFSRcolor4[505]&LFSRcolor4[499]&LFSRcolor4[479]);
    BiasedRNG[834] = (LFSRcolor4[283]&LFSRcolor4[378]&LFSRcolor4[186]&LFSRcolor4[543]);
    BiasedRNG[835] = (LFSRcolor4[108]&LFSRcolor4[632]&LFSRcolor4[358]&LFSRcolor4[62]);
    BiasedRNG[836] = (LFSRcolor4[642]&LFSRcolor4[353]&LFSRcolor4[545]&LFSRcolor4[17]);
    BiasedRNG[837] = (LFSRcolor4[577]&LFSRcolor4[416]&LFSRcolor4[246]&LFSRcolor4[342]);
    BiasedRNG[838] = (LFSRcolor4[404]&LFSRcolor4[28]&LFSRcolor4[271]&LFSRcolor4[387]);
    BiasedRNG[839] = (LFSRcolor4[611]&LFSRcolor4[265]&LFSRcolor4[208]&LFSRcolor4[646]);
    BiasedRNG[840] = (LFSRcolor4[33]&LFSRcolor4[341]&LFSRcolor4[711]&LFSRcolor4[671]);
    BiasedRNG[841] = (LFSRcolor4[488]&LFSRcolor4[14]&LFSRcolor4[539]&LFSRcolor4[94]);
    BiasedRNG[842] = (LFSRcolor4[706]&LFSRcolor4[190]&LFSRcolor4[603]&LFSRcolor4[200]);
    BiasedRNG[843] = (LFSRcolor4[448]&LFSRcolor4[591]&LFSRcolor4[716]&LFSRcolor4[376]);
    BiasedRNG[844] = (LFSRcolor4[235]&LFSRcolor4[324]&LFSRcolor4[73]&LFSRcolor4[123]);
    BiasedRNG[845] = (LFSRcolor4[77]&LFSRcolor4[212]&LFSRcolor4[44]&LFSRcolor4[288]);
    BiasedRNG[846] = (LFSRcolor4[732]&LFSRcolor4[720]&LFSRcolor4[155]&LFSRcolor4[345]);
    BiasedRNG[847] = (LFSRcolor4[354]&LFSRcolor4[509]&LFSRcolor4[723]&LFSRcolor4[639]);
    BiasedRNG[848] = (LFSRcolor4[109]&LFSRcolor4[51]&LFSRcolor4[333]&LFSRcolor4[7]);
    BiasedRNG[849] = (LFSRcolor4[713]&LFSRcolor4[130]&LFSRcolor4[659]&LFSRcolor4[144]);
    BiasedRNG[850] = (LFSRcolor4[312]&LFSRcolor4[719]&LFSRcolor4[120]&LFSRcolor4[287]);
    BiasedRNG[851] = (LFSRcolor4[138]&LFSRcolor4[629]&LFSRcolor4[710]&LFSRcolor4[199]);
    BiasedRNG[852] = (LFSRcolor4[95]&LFSRcolor4[661]&LFSRcolor4[164]&LFSRcolor4[19]);
    BiasedRNG[853] = (LFSRcolor4[80]&LFSRcolor4[516]&LFSRcolor4[238]&LFSRcolor4[139]);
    BiasedRNG[854] = (LFSRcolor4[665]&LFSRcolor4[726]&LFSRcolor4[71]&LFSRcolor4[526]);
    BiasedRNG[855] = (LFSRcolor4[361]&LFSRcolor4[571]&LFSRcolor4[531]&LFSRcolor4[228]);
    BiasedRNG[856] = (LFSRcolor4[570]&LFSRcolor4[689]&LFSRcolor4[216]&LFSRcolor4[232]);
    BiasedRNG[857] = (LFSRcolor4[457]&LFSRcolor4[514]&LFSRcolor4[532]&LFSRcolor4[555]);
    BiasedRNG[858] = (LFSRcolor4[431]&LFSRcolor4[335]&LFSRcolor4[731]&LFSRcolor4[607]);
    BiasedRNG[859] = (LFSRcolor4[425]&LFSRcolor4[491]&LFSRcolor4[54]&LFSRcolor4[184]);
    BiasedRNG[860] = (LFSRcolor4[205]&LFSRcolor4[449]&LFSRcolor4[339]&LFSRcolor4[648]);
    BiasedRNG[861] = (LFSRcolor4[619]&LFSRcolor4[152]&LFSRcolor4[254]&LFSRcolor4[349]);
    BiasedRNG[862] = (LFSRcolor4[413]&LFSRcolor4[344]&LFSRcolor4[727]&LFSRcolor4[141]);
    BiasedRNG[863] = (LFSRcolor4[640]&LFSRcolor4[106]&LFSRcolor4[383]&LFSRcolor4[433]);
    BiasedRNG[864] = (LFSRcolor4[215]&LFSRcolor4[557]&LFSRcolor4[651]&LFSRcolor4[614]);
    BiasedRNG[865] = (LFSRcolor4[196]&LFSRcolor4[392]&LFSRcolor4[422]&LFSRcolor4[623]);
    BiasedRNG[866] = (LFSRcolor4[377]&LFSRcolor4[111]&LFSRcolor4[493]&LFSRcolor4[360]);
    BiasedRNG[867] = (LFSRcolor4[627]&LFSRcolor4[289]&LFSRcolor4[507]&LFSRcolor4[6]);
    BiasedRNG[868] = (LFSRcolor4[39]&LFSRcolor4[389]&LFSRcolor4[386]&LFSRcolor4[86]);
    BiasedRNG[869] = (LFSRcolor4[119]&LFSRcolor4[92]&LFSRcolor4[258]&LFSRcolor4[321]);
    BiasedRNG[870] = (LFSRcolor4[430]&LFSRcolor4[82]&LFSRcolor4[239]&LFSRcolor4[307]);
    BiasedRNG[871] = (LFSRcolor4[140]&LFSRcolor4[219]&LFSRcolor4[633]&LFSRcolor4[301]);
    BiasedRNG[872] = (LFSRcolor4[272]&LFSRcolor4[229]&LFSRcolor4[118]&LFSRcolor4[546]);
    BiasedRNG[873] = (LFSRcolor4[549]&LFSRcolor4[402]&LFSRcolor4[508]&LFSRcolor4[676]);
    BiasedRNG[874] = (LFSRcolor4[68]&LFSRcolor4[217]&LFSRcolor4[185]&LFSRcolor4[645]);
    BiasedRNG[875] = (LFSRcolor4[477]&LFSRcolor4[105]&LFSRcolor4[227]&LFSRcolor4[712]);
    BiasedRNG[876] = (LFSRcolor4[29]&LFSRcolor4[302]&LFSRcolor4[364]&LFSRcolor4[529]);
    BiasedRNG[877] = (LFSRcolor4[63]&LFSRcolor4[463]&LFSRcolor4[362]&LFSRcolor4[38]);
    BiasedRNG[878] = (LFSRcolor4[602]&LFSRcolor4[303]&LFSRcolor4[527]&LFSRcolor4[679]);
    BiasedRNG[879] = (LFSRcolor4[495]&LFSRcolor4[687]&LFSRcolor4[261]&LFSRcolor4[617]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule