//Generated automatically via 'Gen_VerilogRunTilDone_LFSR_3-25.ipynb python code'

`timescale 1ns / 1ps

module main(
    input SYS_CLK_100M_P,
    input SYS_CLK_100M_N,
    output W_LED_0,
    output W_LED_1,
    output W_LED_2,
    output W_LED_3
    );

wire sample_clk;
wire color0_clk;
wire color1_clk;
wire color2_clk;
wire color3_clk;
wire color4_clk;
reg [31:0] counter;
initial counter = 32'b0;
reg [15:0] solution;
reg solution_flag;
initial solution_flag = 1'b0;
reg failure;
initial failure = 1'b0;
wire [367:0] LFSRcolor0;
wire [459:0] LFSRcolor1;
wire [321:0] LFSRcolor2;
wire [45:0] LFSRcolor3;
wire [229:0] LFSRcolor4;
reg [277:0] BiasedRNG;       //For I=+/-1 cases
reg [217:0] UnbiasedRNG;   //For I=0 cases
reg [0:519] m;
//To keep from synthesizing away:
assign W_LED_0=m[0];
assign W_LED_1=m[1];
assign W_LED_2=failure;
assign W_LED_3=solution_flag;

//Initialize the system for Reverse operation:
initial m[176] = 1'b1;
initial m[243] = 1'b0;
initial m[253] = 1'b0;
initial m[268] = 1'b1;
initial m[288] = 1'b1;
initial m[313] = 1'b0;
initial m[343] = 1'b1;
initial m[378] = 1'b0;
initial m[413] = 1'b1;
initial m[443] = 1'b1;
initial m[468] = 1'b0;
initial m[488] = 1'b1;
initial m[503] = 1'b1;
initial m[513] = 1'b0;
initial m[518] = 1'b1;
initial m[519] = 1'b1;

//Initialize the PBits clamped to zero:
initial m[242] = 1'b0;
initial m[252] = 1'b0;
initial m[267] = 1'b0;
initial m[287] = 1'b0;
initial m[312] = 1'b0;
initial m[342] = 1'b0;
initial m[377] = 1'b0;
initial m[380] = 1'b0;

//Generate the pseudo-entropy source:
lfsr #(.seed(46'b0010110111100101000000011010101100110100010101)) LFSR0_0(.LFSRregister(LFSRcolor0[45:0]),.clk(sample_clk));
lfsr #(.seed(46'b0011110000101011000110100000101011100100010011)) LFSR0_1(.LFSRregister(LFSRcolor0[91:46]),.clk(sample_clk));
lfsr #(.seed(46'b1100001101001100000011110100110010101011010011)) LFSR0_2(.LFSRregister(LFSRcolor0[137:92]),.clk(sample_clk));
lfsr #(.seed(46'b0100111000010101111101001000000000111010100010)) LFSR0_3(.LFSRregister(LFSRcolor0[183:138]),.clk(sample_clk));
lfsr #(.seed(46'b1000101000100100110001110001110111001101010101)) LFSR0_4(.LFSRregister(LFSRcolor0[229:184]),.clk(sample_clk));
lfsr #(.seed(46'b1101010011111111100111000000011001000110100101)) LFSR0_5(.LFSRregister(LFSRcolor0[275:230]),.clk(sample_clk));
lfsr #(.seed(46'b0100000110011000011001111000110101001100111110)) LFSR0_6(.LFSRregister(LFSRcolor0[321:276]),.clk(sample_clk));
lfsr #(.seed(46'b1111110011011001001000001010101010001001110011)) LFSR0_7(.LFSRregister(LFSRcolor0[367:322]),.clk(sample_clk));
lfsr #(.seed(46'b1100100010000000011010100011010010111100011101)) LFSR1_0(.LFSRregister(LFSRcolor1[45:0]),.clk(color0_clk));
lfsr #(.seed(46'b0001011001010101100110011010101101101101011011)) LFSR1_1(.LFSRregister(LFSRcolor1[91:46]),.clk(color0_clk));
lfsr #(.seed(46'b0101111110001010010110110011111101010000110010)) LFSR1_2(.LFSRregister(LFSRcolor1[137:92]),.clk(color0_clk));
lfsr #(.seed(46'b0100111010001000011000110111111101111011010010)) LFSR1_3(.LFSRregister(LFSRcolor1[183:138]),.clk(color0_clk));
lfsr #(.seed(46'b1100011111110010011110010010001110100000101100)) LFSR1_4(.LFSRregister(LFSRcolor1[229:184]),.clk(color0_clk));
lfsr #(.seed(46'b1110110000100001111100001101000111011001110101)) LFSR1_5(.LFSRregister(LFSRcolor1[275:230]),.clk(color0_clk));
lfsr #(.seed(46'b0001100011010010001010011100010011101101100000)) LFSR1_6(.LFSRregister(LFSRcolor1[321:276]),.clk(color0_clk));
lfsr #(.seed(46'b0011111110000000111000111101000000010100101010)) LFSR1_7(.LFSRregister(LFSRcolor1[367:322]),.clk(color0_clk));
lfsr #(.seed(46'b0000011000011111110001001001110110001010101101)) LFSR1_8(.LFSRregister(LFSRcolor1[413:368]),.clk(color0_clk));
lfsr #(.seed(46'b0010001010011010010011001010001010001110001001)) LFSR1_9(.LFSRregister(LFSRcolor1[459:414]),.clk(color0_clk));
lfsr #(.seed(46'b1010100010010011101010110110001100000101100101)) LFSR2_0(.LFSRregister(LFSRcolor2[45:0]),.clk(color1_clk));
lfsr #(.seed(46'b0001000011101001111111000001001010010000000010)) LFSR2_1(.LFSRregister(LFSRcolor2[91:46]),.clk(color1_clk));
lfsr #(.seed(46'b1011001001111000101101111101100011110111111011)) LFSR2_2(.LFSRregister(LFSRcolor2[137:92]),.clk(color1_clk));
lfsr #(.seed(46'b1010100101010101001100110101001110000101100000)) LFSR2_3(.LFSRregister(LFSRcolor2[183:138]),.clk(color1_clk));
lfsr #(.seed(46'b0010000011111010001011001010110010010000110101)) LFSR2_4(.LFSRregister(LFSRcolor2[229:184]),.clk(color1_clk));
lfsr #(.seed(46'b0101011001111101100101110111011001011101100110)) LFSR2_5(.LFSRregister(LFSRcolor2[275:230]),.clk(color1_clk));
lfsr #(.seed(46'b0111010000000110010111000001001000011010110100)) LFSR2_6(.LFSRregister(LFSRcolor2[321:276]),.clk(color1_clk));
lfsr #(.seed(46'b1000101111101011011101101111011010001101010010)) LFSR3_0(.LFSRregister(LFSRcolor3[45:0]),.clk(color2_clk));
lfsr #(.seed(46'b0110001010001001001100010011111110110010011001)) LFSR4_0(.LFSRregister(LFSRcolor4[45:0]),.clk(color3_clk));
lfsr #(.seed(46'b1100111101110100111101110110001111011100110001)) LFSR4_1(.LFSRregister(LFSRcolor4[91:46]),.clk(color3_clk));
lfsr #(.seed(46'b1100101000011101011010110010001000010110101110)) LFSR4_2(.LFSRregister(LFSRcolor4[137:92]),.clk(color3_clk));
lfsr #(.seed(46'b0100111011100100011111000101011100101010101010)) LFSR4_3(.LFSRregister(LFSRcolor4[183:138]),.clk(color3_clk));
lfsr #(.seed(46'b1010110100100011110000000101010101100001100001)) LFSR4_4(.LFSRregister(LFSRcolor4[229:184]),.clk(color3_clk));

//Set the initial state of unclamped m to random bits:
initial m[0] = 0;
initial m[1] = 1;
initial m[2] = 0;
initial m[3] = 0;
initial m[4] = 0;
initial m[5] = 1;
initial m[6] = 1;
initial m[7] = 1;
initial m[8] = 0;
initial m[9] = 0;
initial m[10] = 0;
initial m[11] = 1;
initial m[12] = 0;
initial m[13] = 0;
initial m[14] = 0;
initial m[15] = 0;
initial m[16] = 0;
initial m[17] = 1;
initial m[18] = 0;
initial m[19] = 1;
initial m[20] = 0;
initial m[21] = 1;
initial m[22] = 0;
initial m[23] = 1;
initial m[24] = 1;
initial m[25] = 0;
initial m[26] = 0;
initial m[27] = 1;
initial m[28] = 0;
initial m[29] = 1;
initial m[30] = 0;
initial m[31] = 0;
initial m[32] = 0;
initial m[33] = 1;
initial m[34] = 1;
initial m[35] = 1;
initial m[36] = 1;
initial m[37] = 1;
initial m[38] = 0;
initial m[39] = 1;
initial m[40] = 0;
initial m[41] = 0;
initial m[42] = 0;
initial m[43] = 0;
initial m[44] = 0;
initial m[45] = 0;
initial m[46] = 1;
initial m[47] = 0;
initial m[48] = 0;
initial m[49] = 0;
initial m[50] = 1;
initial m[51] = 0;
initial m[52] = 1;
initial m[53] = 1;
initial m[54] = 1;
initial m[55] = 0;
initial m[56] = 0;
initial m[57] = 0;
initial m[58] = 0;
initial m[59] = 1;
initial m[60] = 0;
initial m[61] = 0;
initial m[62] = 0;
initial m[63] = 1;
initial m[64] = 0;
initial m[65] = 1;
initial m[66] = 0;
initial m[67] = 1;
initial m[68] = 0;
initial m[69] = 1;
initial m[70] = 0;
initial m[71] = 1;
initial m[72] = 1;
initial m[73] = 1;
initial m[74] = 0;
initial m[75] = 0;
initial m[76] = 1;
initial m[77] = 1;
initial m[78] = 1;
initial m[79] = 1;
initial m[80] = 1;
initial m[81] = 0;
initial m[82] = 1;
initial m[83] = 1;
initial m[84] = 0;
initial m[85] = 1;
initial m[86] = 0;
initial m[87] = 0;
initial m[88] = 1;
initial m[89] = 0;
initial m[90] = 0;
initial m[91] = 1;
initial m[92] = 1;
initial m[93] = 1;
initial m[94] = 0;
initial m[95] = 0;
initial m[96] = 1;
initial m[97] = 0;
initial m[98] = 0;
initial m[99] = 1;
initial m[100] = 0;
initial m[101] = 1;
initial m[102] = 0;
initial m[103] = 1;
initial m[104] = 0;
initial m[105] = 0;
initial m[106] = 1;
initial m[107] = 1;
initial m[108] = 1;
initial m[109] = 0;
initial m[110] = 1;
initial m[111] = 0;
initial m[112] = 0;
initial m[113] = 1;
initial m[114] = 0;
initial m[115] = 0;
initial m[116] = 0;
initial m[117] = 0;
initial m[118] = 1;
initial m[119] = 1;
initial m[120] = 1;
initial m[121] = 0;
initial m[122] = 0;
initial m[123] = 1;
initial m[124] = 1;
initial m[125] = 1;
initial m[126] = 0;
initial m[127] = 0;
initial m[128] = 0;
initial m[129] = 0;
initial m[130] = 0;
initial m[131] = 0;
initial m[132] = 1;
initial m[133] = 0;
initial m[134] = 1;
initial m[135] = 0;
initial m[136] = 1;
initial m[137] = 1;
initial m[138] = 1;
initial m[139] = 0;
initial m[140] = 1;
initial m[141] = 0;
initial m[142] = 1;
initial m[143] = 0;
initial m[144] = 1;
initial m[145] = 0;
initial m[146] = 1;
initial m[147] = 1;
initial m[148] = 0;
initial m[149] = 1;
initial m[150] = 0;
initial m[151] = 0;
initial m[152] = 1;
initial m[153] = 1;
initial m[154] = 1;
initial m[155] = 0;
initial m[156] = 0;
initial m[157] = 0;
initial m[158] = 0;
initial m[159] = 1;
initial m[160] = 0;
initial m[161] = 0;
initial m[162] = 1;
initial m[163] = 1;
initial m[164] = 0;
initial m[165] = 1;
initial m[166] = 1;
initial m[167] = 0;
initial m[168] = 1;
initial m[169] = 1;
initial m[170] = 0;
initial m[171] = 0;
initial m[172] = 1;
initial m[173] = 1;
initial m[174] = 0;
initial m[175] = 0;
initial m[177] = 1;
initial m[178] = 1;
initial m[179] = 1;
initial m[180] = 1;
initial m[181] = 0;
initial m[182] = 0;
initial m[183] = 1;
initial m[184] = 1;
initial m[185] = 0;
initial m[186] = 1;
initial m[187] = 1;
initial m[188] = 0;
initial m[189] = 1;
initial m[190] = 1;
initial m[191] = 1;
initial m[192] = 0;
initial m[193] = 0;
initial m[194] = 1;
initial m[195] = 0;
initial m[196] = 0;
initial m[197] = 1;
initial m[198] = 0;
initial m[199] = 0;
initial m[200] = 1;
initial m[201] = 1;
initial m[202] = 0;
initial m[203] = 0;
initial m[204] = 1;
initial m[205] = 1;
initial m[206] = 1;
initial m[207] = 0;
initial m[208] = 1;
initial m[209] = 1;
initial m[210] = 0;
initial m[211] = 1;
initial m[212] = 1;
initial m[213] = 0;
initial m[214] = 1;
initial m[215] = 1;
initial m[216] = 1;
initial m[217] = 0;
initial m[218] = 1;
initial m[219] = 1;
initial m[220] = 0;
initial m[221] = 1;
initial m[222] = 1;
initial m[223] = 0;
initial m[224] = 0;
initial m[225] = 0;
initial m[226] = 0;
initial m[227] = 1;
initial m[228] = 1;
initial m[229] = 0;
initial m[230] = 1;
initial m[231] = 0;
initial m[232] = 1;
initial m[233] = 1;
initial m[234] = 1;
initial m[235] = 0;
initial m[236] = 1;
initial m[237] = 0;
initial m[238] = 1;
initial m[239] = 0;
initial m[240] = 0;
initial m[241] = 0;
initial m[244] = 0;
initial m[245] = 0;
initial m[246] = 1;
initial m[247] = 0;
initial m[248] = 0;
initial m[249] = 1;
initial m[250] = 0;
initial m[251] = 1;
initial m[254] = 1;
initial m[255] = 1;
initial m[256] = 1;
initial m[257] = 1;
initial m[258] = 0;
initial m[259] = 1;
initial m[260] = 1;
initial m[261] = 1;
initial m[262] = 1;
initial m[263] = 0;
initial m[264] = 0;
initial m[265] = 1;
initial m[266] = 0;
initial m[269] = 1;
initial m[270] = 0;
initial m[271] = 1;
initial m[272] = 0;
initial m[273] = 0;
initial m[274] = 0;
initial m[275] = 1;
initial m[276] = 1;
initial m[277] = 1;
initial m[278] = 1;
initial m[279] = 0;
initial m[280] = 1;
initial m[281] = 1;
initial m[282] = 1;
initial m[283] = 1;
initial m[284] = 0;
initial m[285] = 1;
initial m[286] = 0;
initial m[289] = 1;
initial m[290] = 1;
initial m[291] = 1;
initial m[292] = 0;
initial m[293] = 0;
initial m[294] = 0;
initial m[295] = 0;
initial m[296] = 1;
initial m[297] = 1;
initial m[298] = 1;
initial m[299] = 1;
initial m[300] = 1;
initial m[301] = 0;
initial m[302] = 0;
initial m[303] = 0;
initial m[304] = 0;
initial m[305] = 1;
initial m[306] = 0;
initial m[307] = 1;
initial m[308] = 0;
initial m[309] = 0;
initial m[310] = 1;
initial m[311] = 1;
initial m[314] = 0;
initial m[315] = 0;
initial m[316] = 0;
initial m[317] = 1;
initial m[318] = 0;
initial m[319] = 1;
initial m[320] = 1;
initial m[321] = 1;
initial m[322] = 0;
initial m[323] = 1;
initial m[324] = 0;
initial m[325] = 1;
initial m[326] = 0;
initial m[327] = 1;
initial m[328] = 1;
initial m[329] = 1;
initial m[330] = 1;
initial m[331] = 1;
initial m[332] = 0;
initial m[333] = 0;
initial m[334] = 1;
initial m[335] = 1;
initial m[336] = 1;
initial m[337] = 0;
initial m[338] = 0;
initial m[339] = 1;
initial m[340] = 1;
initial m[341] = 1;
initial m[344] = 1;
initial m[345] = 1;
initial m[346] = 0;
initial m[347] = 1;
initial m[348] = 0;
initial m[349] = 0;
initial m[350] = 1;
initial m[351] = 1;
initial m[352] = 1;
initial m[353] = 0;
initial m[354] = 0;
initial m[355] = 0;
initial m[356] = 0;
initial m[357] = 0;
initial m[358] = 1;
initial m[359] = 1;
initial m[360] = 0;
initial m[361] = 1;
initial m[362] = 0;
initial m[363] = 0;
initial m[364] = 0;
initial m[365] = 1;
initial m[366] = 1;
initial m[367] = 0;
initial m[368] = 1;
initial m[369] = 0;
initial m[370] = 1;
initial m[371] = 1;
initial m[372] = 0;
initial m[373] = 1;
initial m[374] = 1;
initial m[375] = 1;
initial m[376] = 0;
initial m[379] = 1;
initial m[381] = 1;
initial m[382] = 1;
initial m[383] = 1;
initial m[384] = 1;
initial m[385] = 0;
initial m[386] = 0;
initial m[387] = 1;
initial m[388] = 0;
initial m[389] = 0;
initial m[390] = 1;
initial m[391] = 1;
initial m[392] = 1;
initial m[393] = 1;
initial m[394] = 1;
initial m[395] = 0;
initial m[396] = 1;
initial m[397] = 1;
initial m[398] = 0;
initial m[399] = 0;
initial m[400] = 1;
initial m[401] = 0;
initial m[402] = 1;
initial m[403] = 1;
initial m[404] = 0;
initial m[405] = 0;
initial m[406] = 1;
initial m[407] = 0;
initial m[408] = 0;
initial m[409] = 0;
initial m[410] = 0;
initial m[411] = 0;
initial m[412] = 1;
initial m[414] = 0;
initial m[415] = 1;
initial m[416] = 1;
initial m[417] = 0;
initial m[418] = 0;
initial m[419] = 1;
initial m[420] = 1;
initial m[421] = 1;
initial m[422] = 1;
initial m[423] = 1;
initial m[424] = 0;
initial m[425] = 0;
initial m[426] = 1;
initial m[427] = 1;
initial m[428] = 0;
initial m[429] = 1;
initial m[430] = 0;
initial m[431] = 1;
initial m[432] = 0;
initial m[433] = 0;
initial m[434] = 1;
initial m[435] = 1;
initial m[436] = 1;
initial m[437] = 1;
initial m[438] = 1;
initial m[439] = 1;
initial m[440] = 1;
initial m[441] = 1;
initial m[442] = 0;
initial m[444] = 0;
initial m[445] = 0;
initial m[446] = 1;
initial m[447] = 1;
initial m[448] = 1;
initial m[449] = 0;
initial m[450] = 0;
initial m[451] = 0;
initial m[452] = 0;
initial m[453] = 0;
initial m[454] = 0;
initial m[455] = 1;
initial m[456] = 0;
initial m[457] = 1;
initial m[458] = 1;
initial m[459] = 1;
initial m[460] = 1;
initial m[461] = 1;
initial m[462] = 1;
initial m[463] = 1;
initial m[464] = 0;
initial m[465] = 1;
initial m[466] = 1;
initial m[467] = 1;
initial m[469] = 0;
initial m[470] = 0;
initial m[471] = 1;
initial m[472] = 0;
initial m[473] = 0;
initial m[474] = 1;
initial m[475] = 1;
initial m[476] = 1;
initial m[477] = 1;
initial m[478] = 0;
initial m[479] = 0;
initial m[480] = 0;
initial m[481] = 0;
initial m[482] = 0;
initial m[483] = 0;
initial m[484] = 0;
initial m[485] = 0;
initial m[486] = 1;
initial m[487] = 1;
initial m[489] = 1;
initial m[490] = 0;
initial m[491] = 1;
initial m[492] = 1;
initial m[493] = 0;
initial m[494] = 0;
initial m[495] = 1;
initial m[496] = 1;
initial m[497] = 1;
initial m[498] = 1;
initial m[499] = 1;
initial m[500] = 1;
initial m[501] = 1;
initial m[502] = 0;
initial m[504] = 0;
initial m[505] = 0;
initial m[506] = 1;
initial m[507] = 1;
initial m[508] = 1;
initial m[509] = 1;
initial m[510] = 1;
initial m[511] = 0;
initial m[512] = 1;
initial m[514] = 0;
initial m[515] = 0;
initial m[516] = 1;
initial m[517] = 1;

//Check if the factor state matches the product state:
always @(posedge sample_clk) begin
    solution = {m[7],m[6],m[5],m[4],m[3],m[2],m[1],m[0]}*{m[15],m[14],m[13],m[12],m[11],m[10],m[9],m[8]};
end

always @(negedge sample_clk) begin
    if (solution == 16'b1101101101011001)
        solution_flag = 1'b1;
    else begin
        if (counter==32'b11111111111111111111111111111111) begin
            failure = 1'b1;
        end else
            counter = counter + 32'b1;
    end
end

//Update the outputs by color:
always @(posedge color0_clk) begin
    m[0] = (((m[16]&~m[17])|(~m[16]&m[17]))&UnbiasedRNG[0])|((m[16]&m[17]));
    m[1] = (((m[18]&~m[19])|(~m[18]&m[19]))&UnbiasedRNG[1])|((m[18]&m[19]));
    m[2] = (((m[20]&~m[21])|(~m[20]&m[21]))&UnbiasedRNG[2])|((m[20]&m[21]));
    m[3] = (((m[22]&~m[23])|(~m[22]&m[23]))&UnbiasedRNG[3])|((m[22]&m[23]));
    m[4] = (((m[24]&~m[25])|(~m[24]&m[25]))&UnbiasedRNG[4])|((m[24]&m[25]));
    m[5] = (((m[26]&~m[27])|(~m[26]&m[27]))&UnbiasedRNG[5])|((m[26]&m[27]));
    m[6] = (((m[28]&~m[29])|(~m[28]&m[29]))&UnbiasedRNG[6])|((m[28]&m[29]));
    m[7] = (((m[30]&~m[31])|(~m[30]&m[31]))&UnbiasedRNG[7])|((m[30]&m[31]));
    m[8] = (((m[32]&~m[33])|(~m[32]&m[33]))&UnbiasedRNG[8])|((m[32]&m[33]));
    m[9] = (((m[34]&~m[35])|(~m[34]&m[35]))&UnbiasedRNG[9])|((m[34]&m[35]));
    m[10] = (((m[36]&~m[37])|(~m[36]&m[37]))&UnbiasedRNG[10])|((m[36]&m[37]));
    m[11] = (((m[38]&~m[39])|(~m[38]&m[39]))&UnbiasedRNG[11])|((m[38]&m[39]));
    m[12] = (((m[40]&~m[41])|(~m[40]&m[41]))&UnbiasedRNG[12])|((m[40]&m[41]));
    m[13] = (((m[42]&~m[43])|(~m[42]&m[43]))&UnbiasedRNG[13])|((m[42]&m[43]));
    m[14] = (((m[44]&~m[45])|(~m[44]&m[45]))&UnbiasedRNG[14])|((m[44]&m[45]));
    m[15] = (((m[46]&~m[47])|(~m[46]&m[47]))&UnbiasedRNG[15])|((m[46]&m[47]));
    m[48] = (((~m[16]&~m[112]&~m[176])|(m[16]&m[112]&~m[176]))&BiasedRNG[0])|(((m[16]&~m[112]&~m[176])|(~m[16]&m[112]&m[176]))&~BiasedRNG[0])|((~m[16]&~m[112]&m[176])|(m[16]&~m[112]&m[176])|(m[16]&m[112]&m[176]));
    m[49] = (((~m[16]&~m[120]&~m[184])|(m[16]&m[120]&~m[184]))&BiasedRNG[1])|(((m[16]&~m[120]&~m[184])|(~m[16]&m[120]&m[184]))&~BiasedRNG[1])|((~m[16]&~m[120]&m[184])|(m[16]&~m[120]&m[184])|(m[16]&m[120]&m[184]));
    m[50] = (((~m[16]&~m[128]&~m[192])|(m[16]&m[128]&~m[192]))&BiasedRNG[2])|(((m[16]&~m[128]&~m[192])|(~m[16]&m[128]&m[192]))&~BiasedRNG[2])|((~m[16]&~m[128]&m[192])|(m[16]&~m[128]&m[192])|(m[16]&m[128]&m[192]));
    m[51] = (((~m[16]&~m[136]&~m[200])|(m[16]&m[136]&~m[200]))&BiasedRNG[3])|(((m[16]&~m[136]&~m[200])|(~m[16]&m[136]&m[200]))&~BiasedRNG[3])|((~m[16]&~m[136]&m[200])|(m[16]&~m[136]&m[200])|(m[16]&m[136]&m[200]));
    m[52] = (((~m[17]&~m[144]&~m[208])|(m[17]&m[144]&~m[208]))&BiasedRNG[4])|(((m[17]&~m[144]&~m[208])|(~m[17]&m[144]&m[208]))&~BiasedRNG[4])|((~m[17]&~m[144]&m[208])|(m[17]&~m[144]&m[208])|(m[17]&m[144]&m[208]));
    m[53] = (((~m[17]&~m[152]&~m[216])|(m[17]&m[152]&~m[216]))&BiasedRNG[5])|(((m[17]&~m[152]&~m[216])|(~m[17]&m[152]&m[216]))&~BiasedRNG[5])|((~m[17]&~m[152]&m[216])|(m[17]&~m[152]&m[216])|(m[17]&m[152]&m[216]));
    m[54] = (((~m[17]&~m[160]&~m[224])|(m[17]&m[160]&~m[224]))&BiasedRNG[6])|(((m[17]&~m[160]&~m[224])|(~m[17]&m[160]&m[224]))&~BiasedRNG[6])|((~m[17]&~m[160]&m[224])|(m[17]&~m[160]&m[224])|(m[17]&m[160]&m[224]));
    m[55] = (((~m[17]&~m[168]&~m[232])|(m[17]&m[168]&~m[232]))&BiasedRNG[7])|(((m[17]&~m[168]&~m[232])|(~m[17]&m[168]&m[232]))&~BiasedRNG[7])|((~m[17]&~m[168]&m[232])|(m[17]&~m[168]&m[232])|(m[17]&m[168]&m[232]));
    m[56] = (((~m[18]&~m[113]&~m[177])|(m[18]&m[113]&~m[177]))&BiasedRNG[8])|(((m[18]&~m[113]&~m[177])|(~m[18]&m[113]&m[177]))&~BiasedRNG[8])|((~m[18]&~m[113]&m[177])|(m[18]&~m[113]&m[177])|(m[18]&m[113]&m[177]));
    m[57] = (((~m[18]&~m[121]&~m[185])|(m[18]&m[121]&~m[185]))&BiasedRNG[9])|(((m[18]&~m[121]&~m[185])|(~m[18]&m[121]&m[185]))&~BiasedRNG[9])|((~m[18]&~m[121]&m[185])|(m[18]&~m[121]&m[185])|(m[18]&m[121]&m[185]));
    m[58] = (((~m[18]&~m[129]&~m[193])|(m[18]&m[129]&~m[193]))&BiasedRNG[10])|(((m[18]&~m[129]&~m[193])|(~m[18]&m[129]&m[193]))&~BiasedRNG[10])|((~m[18]&~m[129]&m[193])|(m[18]&~m[129]&m[193])|(m[18]&m[129]&m[193]));
    m[59] = (((~m[18]&~m[137]&~m[201])|(m[18]&m[137]&~m[201]))&BiasedRNG[11])|(((m[18]&~m[137]&~m[201])|(~m[18]&m[137]&m[201]))&~BiasedRNG[11])|((~m[18]&~m[137]&m[201])|(m[18]&~m[137]&m[201])|(m[18]&m[137]&m[201]));
    m[60] = (((~m[19]&~m[145]&~m[209])|(m[19]&m[145]&~m[209]))&BiasedRNG[12])|(((m[19]&~m[145]&~m[209])|(~m[19]&m[145]&m[209]))&~BiasedRNG[12])|((~m[19]&~m[145]&m[209])|(m[19]&~m[145]&m[209])|(m[19]&m[145]&m[209]));
    m[61] = (((~m[19]&~m[153]&~m[217])|(m[19]&m[153]&~m[217]))&BiasedRNG[13])|(((m[19]&~m[153]&~m[217])|(~m[19]&m[153]&m[217]))&~BiasedRNG[13])|((~m[19]&~m[153]&m[217])|(m[19]&~m[153]&m[217])|(m[19]&m[153]&m[217]));
    m[62] = (((~m[19]&~m[161]&~m[225])|(m[19]&m[161]&~m[225]))&BiasedRNG[14])|(((m[19]&~m[161]&~m[225])|(~m[19]&m[161]&m[225]))&~BiasedRNG[14])|((~m[19]&~m[161]&m[225])|(m[19]&~m[161]&m[225])|(m[19]&m[161]&m[225]));
    m[63] = (((~m[19]&~m[169]&~m[233])|(m[19]&m[169]&~m[233]))&BiasedRNG[15])|(((m[19]&~m[169]&~m[233])|(~m[19]&m[169]&m[233]))&~BiasedRNG[15])|((~m[19]&~m[169]&m[233])|(m[19]&~m[169]&m[233])|(m[19]&m[169]&m[233]));
    m[64] = (((~m[20]&~m[114]&~m[178])|(m[20]&m[114]&~m[178]))&BiasedRNG[16])|(((m[20]&~m[114]&~m[178])|(~m[20]&m[114]&m[178]))&~BiasedRNG[16])|((~m[20]&~m[114]&m[178])|(m[20]&~m[114]&m[178])|(m[20]&m[114]&m[178]));
    m[65] = (((~m[20]&~m[122]&~m[186])|(m[20]&m[122]&~m[186]))&BiasedRNG[17])|(((m[20]&~m[122]&~m[186])|(~m[20]&m[122]&m[186]))&~BiasedRNG[17])|((~m[20]&~m[122]&m[186])|(m[20]&~m[122]&m[186])|(m[20]&m[122]&m[186]));
    m[66] = (((~m[20]&~m[130]&~m[194])|(m[20]&m[130]&~m[194]))&BiasedRNG[18])|(((m[20]&~m[130]&~m[194])|(~m[20]&m[130]&m[194]))&~BiasedRNG[18])|((~m[20]&~m[130]&m[194])|(m[20]&~m[130]&m[194])|(m[20]&m[130]&m[194]));
    m[67] = (((~m[20]&~m[138]&~m[202])|(m[20]&m[138]&~m[202]))&BiasedRNG[19])|(((m[20]&~m[138]&~m[202])|(~m[20]&m[138]&m[202]))&~BiasedRNG[19])|((~m[20]&~m[138]&m[202])|(m[20]&~m[138]&m[202])|(m[20]&m[138]&m[202]));
    m[68] = (((~m[21]&~m[146]&~m[210])|(m[21]&m[146]&~m[210]))&BiasedRNG[20])|(((m[21]&~m[146]&~m[210])|(~m[21]&m[146]&m[210]))&~BiasedRNG[20])|((~m[21]&~m[146]&m[210])|(m[21]&~m[146]&m[210])|(m[21]&m[146]&m[210]));
    m[69] = (((~m[21]&~m[154]&~m[218])|(m[21]&m[154]&~m[218]))&BiasedRNG[21])|(((m[21]&~m[154]&~m[218])|(~m[21]&m[154]&m[218]))&~BiasedRNG[21])|((~m[21]&~m[154]&m[218])|(m[21]&~m[154]&m[218])|(m[21]&m[154]&m[218]));
    m[70] = (((~m[21]&~m[162]&~m[226])|(m[21]&m[162]&~m[226]))&BiasedRNG[22])|(((m[21]&~m[162]&~m[226])|(~m[21]&m[162]&m[226]))&~BiasedRNG[22])|((~m[21]&~m[162]&m[226])|(m[21]&~m[162]&m[226])|(m[21]&m[162]&m[226]));
    m[71] = (((~m[21]&~m[170]&~m[234])|(m[21]&m[170]&~m[234]))&BiasedRNG[23])|(((m[21]&~m[170]&~m[234])|(~m[21]&m[170]&m[234]))&~BiasedRNG[23])|((~m[21]&~m[170]&m[234])|(m[21]&~m[170]&m[234])|(m[21]&m[170]&m[234]));
    m[72] = (((~m[22]&~m[115]&~m[179])|(m[22]&m[115]&~m[179]))&BiasedRNG[24])|(((m[22]&~m[115]&~m[179])|(~m[22]&m[115]&m[179]))&~BiasedRNG[24])|((~m[22]&~m[115]&m[179])|(m[22]&~m[115]&m[179])|(m[22]&m[115]&m[179]));
    m[73] = (((~m[22]&~m[123]&~m[187])|(m[22]&m[123]&~m[187]))&BiasedRNG[25])|(((m[22]&~m[123]&~m[187])|(~m[22]&m[123]&m[187]))&~BiasedRNG[25])|((~m[22]&~m[123]&m[187])|(m[22]&~m[123]&m[187])|(m[22]&m[123]&m[187]));
    m[74] = (((~m[22]&~m[131]&~m[195])|(m[22]&m[131]&~m[195]))&BiasedRNG[26])|(((m[22]&~m[131]&~m[195])|(~m[22]&m[131]&m[195]))&~BiasedRNG[26])|((~m[22]&~m[131]&m[195])|(m[22]&~m[131]&m[195])|(m[22]&m[131]&m[195]));
    m[75] = (((~m[22]&~m[139]&~m[203])|(m[22]&m[139]&~m[203]))&BiasedRNG[27])|(((m[22]&~m[139]&~m[203])|(~m[22]&m[139]&m[203]))&~BiasedRNG[27])|((~m[22]&~m[139]&m[203])|(m[22]&~m[139]&m[203])|(m[22]&m[139]&m[203]));
    m[76] = (((~m[23]&~m[147]&~m[211])|(m[23]&m[147]&~m[211]))&BiasedRNG[28])|(((m[23]&~m[147]&~m[211])|(~m[23]&m[147]&m[211]))&~BiasedRNG[28])|((~m[23]&~m[147]&m[211])|(m[23]&~m[147]&m[211])|(m[23]&m[147]&m[211]));
    m[77] = (((~m[23]&~m[155]&~m[219])|(m[23]&m[155]&~m[219]))&BiasedRNG[29])|(((m[23]&~m[155]&~m[219])|(~m[23]&m[155]&m[219]))&~BiasedRNG[29])|((~m[23]&~m[155]&m[219])|(m[23]&~m[155]&m[219])|(m[23]&m[155]&m[219]));
    m[78] = (((~m[23]&~m[163]&~m[227])|(m[23]&m[163]&~m[227]))&BiasedRNG[30])|(((m[23]&~m[163]&~m[227])|(~m[23]&m[163]&m[227]))&~BiasedRNG[30])|((~m[23]&~m[163]&m[227])|(m[23]&~m[163]&m[227])|(m[23]&m[163]&m[227]));
    m[79] = (((~m[23]&~m[171]&~m[235])|(m[23]&m[171]&~m[235]))&BiasedRNG[31])|(((m[23]&~m[171]&~m[235])|(~m[23]&m[171]&m[235]))&~BiasedRNG[31])|((~m[23]&~m[171]&m[235])|(m[23]&~m[171]&m[235])|(m[23]&m[171]&m[235]));
    m[80] = (((~m[24]&~m[116]&~m[180])|(m[24]&m[116]&~m[180]))&BiasedRNG[32])|(((m[24]&~m[116]&~m[180])|(~m[24]&m[116]&m[180]))&~BiasedRNG[32])|((~m[24]&~m[116]&m[180])|(m[24]&~m[116]&m[180])|(m[24]&m[116]&m[180]));
    m[81] = (((~m[24]&~m[124]&~m[188])|(m[24]&m[124]&~m[188]))&BiasedRNG[33])|(((m[24]&~m[124]&~m[188])|(~m[24]&m[124]&m[188]))&~BiasedRNG[33])|((~m[24]&~m[124]&m[188])|(m[24]&~m[124]&m[188])|(m[24]&m[124]&m[188]));
    m[82] = (((~m[24]&~m[132]&~m[196])|(m[24]&m[132]&~m[196]))&BiasedRNG[34])|(((m[24]&~m[132]&~m[196])|(~m[24]&m[132]&m[196]))&~BiasedRNG[34])|((~m[24]&~m[132]&m[196])|(m[24]&~m[132]&m[196])|(m[24]&m[132]&m[196]));
    m[83] = (((~m[24]&~m[140]&~m[204])|(m[24]&m[140]&~m[204]))&BiasedRNG[35])|(((m[24]&~m[140]&~m[204])|(~m[24]&m[140]&m[204]))&~BiasedRNG[35])|((~m[24]&~m[140]&m[204])|(m[24]&~m[140]&m[204])|(m[24]&m[140]&m[204]));
    m[84] = (((~m[25]&~m[148]&~m[212])|(m[25]&m[148]&~m[212]))&BiasedRNG[36])|(((m[25]&~m[148]&~m[212])|(~m[25]&m[148]&m[212]))&~BiasedRNG[36])|((~m[25]&~m[148]&m[212])|(m[25]&~m[148]&m[212])|(m[25]&m[148]&m[212]));
    m[85] = (((~m[25]&~m[156]&~m[220])|(m[25]&m[156]&~m[220]))&BiasedRNG[37])|(((m[25]&~m[156]&~m[220])|(~m[25]&m[156]&m[220]))&~BiasedRNG[37])|((~m[25]&~m[156]&m[220])|(m[25]&~m[156]&m[220])|(m[25]&m[156]&m[220]));
    m[86] = (((~m[25]&~m[164]&~m[228])|(m[25]&m[164]&~m[228]))&BiasedRNG[38])|(((m[25]&~m[164]&~m[228])|(~m[25]&m[164]&m[228]))&~BiasedRNG[38])|((~m[25]&~m[164]&m[228])|(m[25]&~m[164]&m[228])|(m[25]&m[164]&m[228]));
    m[87] = (((~m[25]&~m[172]&~m[236])|(m[25]&m[172]&~m[236]))&BiasedRNG[39])|(((m[25]&~m[172]&~m[236])|(~m[25]&m[172]&m[236]))&~BiasedRNG[39])|((~m[25]&~m[172]&m[236])|(m[25]&~m[172]&m[236])|(m[25]&m[172]&m[236]));
    m[88] = (((~m[26]&~m[117]&~m[181])|(m[26]&m[117]&~m[181]))&BiasedRNG[40])|(((m[26]&~m[117]&~m[181])|(~m[26]&m[117]&m[181]))&~BiasedRNG[40])|((~m[26]&~m[117]&m[181])|(m[26]&~m[117]&m[181])|(m[26]&m[117]&m[181]));
    m[89] = (((~m[26]&~m[125]&~m[189])|(m[26]&m[125]&~m[189]))&BiasedRNG[41])|(((m[26]&~m[125]&~m[189])|(~m[26]&m[125]&m[189]))&~BiasedRNG[41])|((~m[26]&~m[125]&m[189])|(m[26]&~m[125]&m[189])|(m[26]&m[125]&m[189]));
    m[90] = (((~m[26]&~m[133]&~m[197])|(m[26]&m[133]&~m[197]))&BiasedRNG[42])|(((m[26]&~m[133]&~m[197])|(~m[26]&m[133]&m[197]))&~BiasedRNG[42])|((~m[26]&~m[133]&m[197])|(m[26]&~m[133]&m[197])|(m[26]&m[133]&m[197]));
    m[91] = (((~m[26]&~m[141]&~m[205])|(m[26]&m[141]&~m[205]))&BiasedRNG[43])|(((m[26]&~m[141]&~m[205])|(~m[26]&m[141]&m[205]))&~BiasedRNG[43])|((~m[26]&~m[141]&m[205])|(m[26]&~m[141]&m[205])|(m[26]&m[141]&m[205]));
    m[92] = (((~m[27]&~m[149]&~m[213])|(m[27]&m[149]&~m[213]))&BiasedRNG[44])|(((m[27]&~m[149]&~m[213])|(~m[27]&m[149]&m[213]))&~BiasedRNG[44])|((~m[27]&~m[149]&m[213])|(m[27]&~m[149]&m[213])|(m[27]&m[149]&m[213]));
    m[93] = (((~m[27]&~m[157]&~m[221])|(m[27]&m[157]&~m[221]))&BiasedRNG[45])|(((m[27]&~m[157]&~m[221])|(~m[27]&m[157]&m[221]))&~BiasedRNG[45])|((~m[27]&~m[157]&m[221])|(m[27]&~m[157]&m[221])|(m[27]&m[157]&m[221]));
    m[94] = (((~m[27]&~m[165]&~m[229])|(m[27]&m[165]&~m[229]))&BiasedRNG[46])|(((m[27]&~m[165]&~m[229])|(~m[27]&m[165]&m[229]))&~BiasedRNG[46])|((~m[27]&~m[165]&m[229])|(m[27]&~m[165]&m[229])|(m[27]&m[165]&m[229]));
    m[95] = (((~m[27]&~m[173]&~m[237])|(m[27]&m[173]&~m[237]))&BiasedRNG[47])|(((m[27]&~m[173]&~m[237])|(~m[27]&m[173]&m[237]))&~BiasedRNG[47])|((~m[27]&~m[173]&m[237])|(m[27]&~m[173]&m[237])|(m[27]&m[173]&m[237]));
    m[96] = (((~m[28]&~m[118]&~m[182])|(m[28]&m[118]&~m[182]))&BiasedRNG[48])|(((m[28]&~m[118]&~m[182])|(~m[28]&m[118]&m[182]))&~BiasedRNG[48])|((~m[28]&~m[118]&m[182])|(m[28]&~m[118]&m[182])|(m[28]&m[118]&m[182]));
    m[97] = (((~m[28]&~m[126]&~m[190])|(m[28]&m[126]&~m[190]))&BiasedRNG[49])|(((m[28]&~m[126]&~m[190])|(~m[28]&m[126]&m[190]))&~BiasedRNG[49])|((~m[28]&~m[126]&m[190])|(m[28]&~m[126]&m[190])|(m[28]&m[126]&m[190]));
    m[98] = (((~m[28]&~m[134]&~m[198])|(m[28]&m[134]&~m[198]))&BiasedRNG[50])|(((m[28]&~m[134]&~m[198])|(~m[28]&m[134]&m[198]))&~BiasedRNG[50])|((~m[28]&~m[134]&m[198])|(m[28]&~m[134]&m[198])|(m[28]&m[134]&m[198]));
    m[99] = (((~m[28]&~m[142]&~m[206])|(m[28]&m[142]&~m[206]))&BiasedRNG[51])|(((m[28]&~m[142]&~m[206])|(~m[28]&m[142]&m[206]))&~BiasedRNG[51])|((~m[28]&~m[142]&m[206])|(m[28]&~m[142]&m[206])|(m[28]&m[142]&m[206]));
    m[100] = (((~m[29]&~m[150]&~m[214])|(m[29]&m[150]&~m[214]))&BiasedRNG[52])|(((m[29]&~m[150]&~m[214])|(~m[29]&m[150]&m[214]))&~BiasedRNG[52])|((~m[29]&~m[150]&m[214])|(m[29]&~m[150]&m[214])|(m[29]&m[150]&m[214]));
    m[101] = (((~m[29]&~m[158]&~m[222])|(m[29]&m[158]&~m[222]))&BiasedRNG[53])|(((m[29]&~m[158]&~m[222])|(~m[29]&m[158]&m[222]))&~BiasedRNG[53])|((~m[29]&~m[158]&m[222])|(m[29]&~m[158]&m[222])|(m[29]&m[158]&m[222]));
    m[102] = (((~m[29]&~m[166]&~m[230])|(m[29]&m[166]&~m[230]))&BiasedRNG[54])|(((m[29]&~m[166]&~m[230])|(~m[29]&m[166]&m[230]))&~BiasedRNG[54])|((~m[29]&~m[166]&m[230])|(m[29]&~m[166]&m[230])|(m[29]&m[166]&m[230]));
    m[103] = (((~m[29]&~m[174]&~m[238])|(m[29]&m[174]&~m[238]))&BiasedRNG[55])|(((m[29]&~m[174]&~m[238])|(~m[29]&m[174]&m[238]))&~BiasedRNG[55])|((~m[29]&~m[174]&m[238])|(m[29]&~m[174]&m[238])|(m[29]&m[174]&m[238]));
    m[104] = (((~m[30]&~m[119]&~m[183])|(m[30]&m[119]&~m[183]))&BiasedRNG[56])|(((m[30]&~m[119]&~m[183])|(~m[30]&m[119]&m[183]))&~BiasedRNG[56])|((~m[30]&~m[119]&m[183])|(m[30]&~m[119]&m[183])|(m[30]&m[119]&m[183]));
    m[105] = (((~m[30]&~m[127]&~m[191])|(m[30]&m[127]&~m[191]))&BiasedRNG[57])|(((m[30]&~m[127]&~m[191])|(~m[30]&m[127]&m[191]))&~BiasedRNG[57])|((~m[30]&~m[127]&m[191])|(m[30]&~m[127]&m[191])|(m[30]&m[127]&m[191]));
    m[106] = (((~m[30]&~m[135]&~m[199])|(m[30]&m[135]&~m[199]))&BiasedRNG[58])|(((m[30]&~m[135]&~m[199])|(~m[30]&m[135]&m[199]))&~BiasedRNG[58])|((~m[30]&~m[135]&m[199])|(m[30]&~m[135]&m[199])|(m[30]&m[135]&m[199]));
    m[107] = (((~m[30]&~m[143]&~m[207])|(m[30]&m[143]&~m[207]))&BiasedRNG[59])|(((m[30]&~m[143]&~m[207])|(~m[30]&m[143]&m[207]))&~BiasedRNG[59])|((~m[30]&~m[143]&m[207])|(m[30]&~m[143]&m[207])|(m[30]&m[143]&m[207]));
    m[108] = (((~m[31]&~m[151]&~m[215])|(m[31]&m[151]&~m[215]))&BiasedRNG[60])|(((m[31]&~m[151]&~m[215])|(~m[31]&m[151]&m[215]))&~BiasedRNG[60])|((~m[31]&~m[151]&m[215])|(m[31]&~m[151]&m[215])|(m[31]&m[151]&m[215]));
    m[109] = (((~m[31]&~m[159]&~m[223])|(m[31]&m[159]&~m[223]))&BiasedRNG[61])|(((m[31]&~m[159]&~m[223])|(~m[31]&m[159]&m[223]))&~BiasedRNG[61])|((~m[31]&~m[159]&m[223])|(m[31]&~m[159]&m[223])|(m[31]&m[159]&m[223]));
    m[110] = (((~m[31]&~m[167]&~m[231])|(m[31]&m[167]&~m[231]))&BiasedRNG[62])|(((m[31]&~m[167]&~m[231])|(~m[31]&m[167]&m[231]))&~BiasedRNG[62])|((~m[31]&~m[167]&m[231])|(m[31]&~m[167]&m[231])|(m[31]&m[167]&m[231]));
    m[111] = (((~m[31]&~m[175]&~m[239])|(m[31]&m[175]&~m[239]))&BiasedRNG[63])|(((m[31]&~m[175]&~m[239])|(~m[31]&m[175]&m[239]))&~BiasedRNG[63])|((~m[31]&~m[175]&m[239])|(m[31]&~m[175]&m[239])|(m[31]&m[175]&m[239]));
    m[240] = (((m[177]&~m[241]&~m[242]&~m[243]&~m[244])|(~m[177]&~m[241]&~m[242]&m[243]&~m[244])|(m[177]&m[241]&~m[242]&m[243]&~m[244])|(m[177]&~m[241]&m[242]&m[243]&~m[244])|(~m[177]&m[241]&~m[242]&~m[243]&m[244])|(~m[177]&~m[241]&m[242]&~m[243]&m[244])|(m[177]&m[241]&m[242]&~m[243]&m[244])|(~m[177]&m[241]&m[242]&m[243]&m[244]))&UnbiasedRNG[16])|((m[177]&~m[241]&~m[242]&m[243]&~m[244])|(~m[177]&~m[241]&~m[242]&~m[243]&m[244])|(m[177]&~m[241]&~m[242]&~m[243]&m[244])|(m[177]&m[241]&~m[242]&~m[243]&m[244])|(m[177]&~m[241]&m[242]&~m[243]&m[244])|(~m[177]&~m[241]&~m[242]&m[243]&m[244])|(m[177]&~m[241]&~m[242]&m[243]&m[244])|(~m[177]&m[241]&~m[242]&m[243]&m[244])|(m[177]&m[241]&~m[242]&m[243]&m[244])|(~m[177]&~m[241]&m[242]&m[243]&m[244])|(m[177]&~m[241]&m[242]&m[243]&m[244])|(m[177]&m[241]&m[242]&m[243]&m[244]));
    m[245] = (((m[178]&~m[246]&~m[247]&~m[248]&~m[249])|(~m[178]&~m[246]&~m[247]&m[248]&~m[249])|(m[178]&m[246]&~m[247]&m[248]&~m[249])|(m[178]&~m[246]&m[247]&m[248]&~m[249])|(~m[178]&m[246]&~m[247]&~m[248]&m[249])|(~m[178]&~m[246]&m[247]&~m[248]&m[249])|(m[178]&m[246]&m[247]&~m[248]&m[249])|(~m[178]&m[246]&m[247]&m[248]&m[249]))&UnbiasedRNG[17])|((m[178]&~m[246]&~m[247]&m[248]&~m[249])|(~m[178]&~m[246]&~m[247]&~m[248]&m[249])|(m[178]&~m[246]&~m[247]&~m[248]&m[249])|(m[178]&m[246]&~m[247]&~m[248]&m[249])|(m[178]&~m[246]&m[247]&~m[248]&m[249])|(~m[178]&~m[246]&~m[247]&m[248]&m[249])|(m[178]&~m[246]&~m[247]&m[248]&m[249])|(~m[178]&m[246]&~m[247]&m[248]&m[249])|(m[178]&m[246]&~m[247]&m[248]&m[249])|(~m[178]&~m[246]&m[247]&m[248]&m[249])|(m[178]&~m[246]&m[247]&m[248]&m[249])|(m[178]&m[246]&m[247]&m[248]&m[249]));
    m[250] = (((m[248]&~m[251]&~m[252]&~m[253]&~m[254])|(~m[248]&~m[251]&~m[252]&m[253]&~m[254])|(m[248]&m[251]&~m[252]&m[253]&~m[254])|(m[248]&~m[251]&m[252]&m[253]&~m[254])|(~m[248]&m[251]&~m[252]&~m[253]&m[254])|(~m[248]&~m[251]&m[252]&~m[253]&m[254])|(m[248]&m[251]&m[252]&~m[253]&m[254])|(~m[248]&m[251]&m[252]&m[253]&m[254]))&UnbiasedRNG[18])|((m[248]&~m[251]&~m[252]&m[253]&~m[254])|(~m[248]&~m[251]&~m[252]&~m[253]&m[254])|(m[248]&~m[251]&~m[252]&~m[253]&m[254])|(m[248]&m[251]&~m[252]&~m[253]&m[254])|(m[248]&~m[251]&m[252]&~m[253]&m[254])|(~m[248]&~m[251]&~m[252]&m[253]&m[254])|(m[248]&~m[251]&~m[252]&m[253]&m[254])|(~m[248]&m[251]&~m[252]&m[253]&m[254])|(m[248]&m[251]&~m[252]&m[253]&m[254])|(~m[248]&~m[251]&m[252]&m[253]&m[254])|(m[248]&~m[251]&m[252]&m[253]&m[254])|(m[248]&m[251]&m[252]&m[253]&m[254]));
    m[255] = (((m[179]&~m[256]&~m[257]&~m[258]&~m[259])|(~m[179]&~m[256]&~m[257]&m[258]&~m[259])|(m[179]&m[256]&~m[257]&m[258]&~m[259])|(m[179]&~m[256]&m[257]&m[258]&~m[259])|(~m[179]&m[256]&~m[257]&~m[258]&m[259])|(~m[179]&~m[256]&m[257]&~m[258]&m[259])|(m[179]&m[256]&m[257]&~m[258]&m[259])|(~m[179]&m[256]&m[257]&m[258]&m[259]))&UnbiasedRNG[19])|((m[179]&~m[256]&~m[257]&m[258]&~m[259])|(~m[179]&~m[256]&~m[257]&~m[258]&m[259])|(m[179]&~m[256]&~m[257]&~m[258]&m[259])|(m[179]&m[256]&~m[257]&~m[258]&m[259])|(m[179]&~m[256]&m[257]&~m[258]&m[259])|(~m[179]&~m[256]&~m[257]&m[258]&m[259])|(m[179]&~m[256]&~m[257]&m[258]&m[259])|(~m[179]&m[256]&~m[257]&m[258]&m[259])|(m[179]&m[256]&~m[257]&m[258]&m[259])|(~m[179]&~m[256]&m[257]&m[258]&m[259])|(m[179]&~m[256]&m[257]&m[258]&m[259])|(m[179]&m[256]&m[257]&m[258]&m[259]));
    m[260] = (((m[258]&~m[261]&~m[262]&~m[263]&~m[264])|(~m[258]&~m[261]&~m[262]&m[263]&~m[264])|(m[258]&m[261]&~m[262]&m[263]&~m[264])|(m[258]&~m[261]&m[262]&m[263]&~m[264])|(~m[258]&m[261]&~m[262]&~m[263]&m[264])|(~m[258]&~m[261]&m[262]&~m[263]&m[264])|(m[258]&m[261]&m[262]&~m[263]&m[264])|(~m[258]&m[261]&m[262]&m[263]&m[264]))&UnbiasedRNG[20])|((m[258]&~m[261]&~m[262]&m[263]&~m[264])|(~m[258]&~m[261]&~m[262]&~m[263]&m[264])|(m[258]&~m[261]&~m[262]&~m[263]&m[264])|(m[258]&m[261]&~m[262]&~m[263]&m[264])|(m[258]&~m[261]&m[262]&~m[263]&m[264])|(~m[258]&~m[261]&~m[262]&m[263]&m[264])|(m[258]&~m[261]&~m[262]&m[263]&m[264])|(~m[258]&m[261]&~m[262]&m[263]&m[264])|(m[258]&m[261]&~m[262]&m[263]&m[264])|(~m[258]&~m[261]&m[262]&m[263]&m[264])|(m[258]&~m[261]&m[262]&m[263]&m[264])|(m[258]&m[261]&m[262]&m[263]&m[264]));
    m[265] = (((m[263]&~m[266]&~m[267]&~m[268]&~m[269])|(~m[263]&~m[266]&~m[267]&m[268]&~m[269])|(m[263]&m[266]&~m[267]&m[268]&~m[269])|(m[263]&~m[266]&m[267]&m[268]&~m[269])|(~m[263]&m[266]&~m[267]&~m[268]&m[269])|(~m[263]&~m[266]&m[267]&~m[268]&m[269])|(m[263]&m[266]&m[267]&~m[268]&m[269])|(~m[263]&m[266]&m[267]&m[268]&m[269]))&UnbiasedRNG[21])|((m[263]&~m[266]&~m[267]&m[268]&~m[269])|(~m[263]&~m[266]&~m[267]&~m[268]&m[269])|(m[263]&~m[266]&~m[267]&~m[268]&m[269])|(m[263]&m[266]&~m[267]&~m[268]&m[269])|(m[263]&~m[266]&m[267]&~m[268]&m[269])|(~m[263]&~m[266]&~m[267]&m[268]&m[269])|(m[263]&~m[266]&~m[267]&m[268]&m[269])|(~m[263]&m[266]&~m[267]&m[268]&m[269])|(m[263]&m[266]&~m[267]&m[268]&m[269])|(~m[263]&~m[266]&m[267]&m[268]&m[269])|(m[263]&~m[266]&m[267]&m[268]&m[269])|(m[263]&m[266]&m[267]&m[268]&m[269]));
    m[270] = (((m[180]&~m[271]&~m[272]&~m[273]&~m[274])|(~m[180]&~m[271]&~m[272]&m[273]&~m[274])|(m[180]&m[271]&~m[272]&m[273]&~m[274])|(m[180]&~m[271]&m[272]&m[273]&~m[274])|(~m[180]&m[271]&~m[272]&~m[273]&m[274])|(~m[180]&~m[271]&m[272]&~m[273]&m[274])|(m[180]&m[271]&m[272]&~m[273]&m[274])|(~m[180]&m[271]&m[272]&m[273]&m[274]))&UnbiasedRNG[22])|((m[180]&~m[271]&~m[272]&m[273]&~m[274])|(~m[180]&~m[271]&~m[272]&~m[273]&m[274])|(m[180]&~m[271]&~m[272]&~m[273]&m[274])|(m[180]&m[271]&~m[272]&~m[273]&m[274])|(m[180]&~m[271]&m[272]&~m[273]&m[274])|(~m[180]&~m[271]&~m[272]&m[273]&m[274])|(m[180]&~m[271]&~m[272]&m[273]&m[274])|(~m[180]&m[271]&~m[272]&m[273]&m[274])|(m[180]&m[271]&~m[272]&m[273]&m[274])|(~m[180]&~m[271]&m[272]&m[273]&m[274])|(m[180]&~m[271]&m[272]&m[273]&m[274])|(m[180]&m[271]&m[272]&m[273]&m[274]));
    m[275] = (((m[273]&~m[276]&~m[277]&~m[278]&~m[279])|(~m[273]&~m[276]&~m[277]&m[278]&~m[279])|(m[273]&m[276]&~m[277]&m[278]&~m[279])|(m[273]&~m[276]&m[277]&m[278]&~m[279])|(~m[273]&m[276]&~m[277]&~m[278]&m[279])|(~m[273]&~m[276]&m[277]&~m[278]&m[279])|(m[273]&m[276]&m[277]&~m[278]&m[279])|(~m[273]&m[276]&m[277]&m[278]&m[279]))&UnbiasedRNG[23])|((m[273]&~m[276]&~m[277]&m[278]&~m[279])|(~m[273]&~m[276]&~m[277]&~m[278]&m[279])|(m[273]&~m[276]&~m[277]&~m[278]&m[279])|(m[273]&m[276]&~m[277]&~m[278]&m[279])|(m[273]&~m[276]&m[277]&~m[278]&m[279])|(~m[273]&~m[276]&~m[277]&m[278]&m[279])|(m[273]&~m[276]&~m[277]&m[278]&m[279])|(~m[273]&m[276]&~m[277]&m[278]&m[279])|(m[273]&m[276]&~m[277]&m[278]&m[279])|(~m[273]&~m[276]&m[277]&m[278]&m[279])|(m[273]&~m[276]&m[277]&m[278]&m[279])|(m[273]&m[276]&m[277]&m[278]&m[279]));
    m[280] = (((m[278]&~m[281]&~m[282]&~m[283]&~m[284])|(~m[278]&~m[281]&~m[282]&m[283]&~m[284])|(m[278]&m[281]&~m[282]&m[283]&~m[284])|(m[278]&~m[281]&m[282]&m[283]&~m[284])|(~m[278]&m[281]&~m[282]&~m[283]&m[284])|(~m[278]&~m[281]&m[282]&~m[283]&m[284])|(m[278]&m[281]&m[282]&~m[283]&m[284])|(~m[278]&m[281]&m[282]&m[283]&m[284]))&UnbiasedRNG[24])|((m[278]&~m[281]&~m[282]&m[283]&~m[284])|(~m[278]&~m[281]&~m[282]&~m[283]&m[284])|(m[278]&~m[281]&~m[282]&~m[283]&m[284])|(m[278]&m[281]&~m[282]&~m[283]&m[284])|(m[278]&~m[281]&m[282]&~m[283]&m[284])|(~m[278]&~m[281]&~m[282]&m[283]&m[284])|(m[278]&~m[281]&~m[282]&m[283]&m[284])|(~m[278]&m[281]&~m[282]&m[283]&m[284])|(m[278]&m[281]&~m[282]&m[283]&m[284])|(~m[278]&~m[281]&m[282]&m[283]&m[284])|(m[278]&~m[281]&m[282]&m[283]&m[284])|(m[278]&m[281]&m[282]&m[283]&m[284]));
    m[285] = (((m[283]&~m[286]&~m[287]&~m[288]&~m[289])|(~m[283]&~m[286]&~m[287]&m[288]&~m[289])|(m[283]&m[286]&~m[287]&m[288]&~m[289])|(m[283]&~m[286]&m[287]&m[288]&~m[289])|(~m[283]&m[286]&~m[287]&~m[288]&m[289])|(~m[283]&~m[286]&m[287]&~m[288]&m[289])|(m[283]&m[286]&m[287]&~m[288]&m[289])|(~m[283]&m[286]&m[287]&m[288]&m[289]))&UnbiasedRNG[25])|((m[283]&~m[286]&~m[287]&m[288]&~m[289])|(~m[283]&~m[286]&~m[287]&~m[288]&m[289])|(m[283]&~m[286]&~m[287]&~m[288]&m[289])|(m[283]&m[286]&~m[287]&~m[288]&m[289])|(m[283]&~m[286]&m[287]&~m[288]&m[289])|(~m[283]&~m[286]&~m[287]&m[288]&m[289])|(m[283]&~m[286]&~m[287]&m[288]&m[289])|(~m[283]&m[286]&~m[287]&m[288]&m[289])|(m[283]&m[286]&~m[287]&m[288]&m[289])|(~m[283]&~m[286]&m[287]&m[288]&m[289])|(m[283]&~m[286]&m[287]&m[288]&m[289])|(m[283]&m[286]&m[287]&m[288]&m[289]));
    m[290] = (((m[181]&~m[291]&~m[292]&~m[293]&~m[294])|(~m[181]&~m[291]&~m[292]&m[293]&~m[294])|(m[181]&m[291]&~m[292]&m[293]&~m[294])|(m[181]&~m[291]&m[292]&m[293]&~m[294])|(~m[181]&m[291]&~m[292]&~m[293]&m[294])|(~m[181]&~m[291]&m[292]&~m[293]&m[294])|(m[181]&m[291]&m[292]&~m[293]&m[294])|(~m[181]&m[291]&m[292]&m[293]&m[294]))&UnbiasedRNG[26])|((m[181]&~m[291]&~m[292]&m[293]&~m[294])|(~m[181]&~m[291]&~m[292]&~m[293]&m[294])|(m[181]&~m[291]&~m[292]&~m[293]&m[294])|(m[181]&m[291]&~m[292]&~m[293]&m[294])|(m[181]&~m[291]&m[292]&~m[293]&m[294])|(~m[181]&~m[291]&~m[292]&m[293]&m[294])|(m[181]&~m[291]&~m[292]&m[293]&m[294])|(~m[181]&m[291]&~m[292]&m[293]&m[294])|(m[181]&m[291]&~m[292]&m[293]&m[294])|(~m[181]&~m[291]&m[292]&m[293]&m[294])|(m[181]&~m[291]&m[292]&m[293]&m[294])|(m[181]&m[291]&m[292]&m[293]&m[294]));
    m[295] = (((m[293]&~m[296]&~m[297]&~m[298]&~m[299])|(~m[293]&~m[296]&~m[297]&m[298]&~m[299])|(m[293]&m[296]&~m[297]&m[298]&~m[299])|(m[293]&~m[296]&m[297]&m[298]&~m[299])|(~m[293]&m[296]&~m[297]&~m[298]&m[299])|(~m[293]&~m[296]&m[297]&~m[298]&m[299])|(m[293]&m[296]&m[297]&~m[298]&m[299])|(~m[293]&m[296]&m[297]&m[298]&m[299]))&UnbiasedRNG[27])|((m[293]&~m[296]&~m[297]&m[298]&~m[299])|(~m[293]&~m[296]&~m[297]&~m[298]&m[299])|(m[293]&~m[296]&~m[297]&~m[298]&m[299])|(m[293]&m[296]&~m[297]&~m[298]&m[299])|(m[293]&~m[296]&m[297]&~m[298]&m[299])|(~m[293]&~m[296]&~m[297]&m[298]&m[299])|(m[293]&~m[296]&~m[297]&m[298]&m[299])|(~m[293]&m[296]&~m[297]&m[298]&m[299])|(m[293]&m[296]&~m[297]&m[298]&m[299])|(~m[293]&~m[296]&m[297]&m[298]&m[299])|(m[293]&~m[296]&m[297]&m[298]&m[299])|(m[293]&m[296]&m[297]&m[298]&m[299]));
    m[300] = (((m[298]&~m[301]&~m[302]&~m[303]&~m[304])|(~m[298]&~m[301]&~m[302]&m[303]&~m[304])|(m[298]&m[301]&~m[302]&m[303]&~m[304])|(m[298]&~m[301]&m[302]&m[303]&~m[304])|(~m[298]&m[301]&~m[302]&~m[303]&m[304])|(~m[298]&~m[301]&m[302]&~m[303]&m[304])|(m[298]&m[301]&m[302]&~m[303]&m[304])|(~m[298]&m[301]&m[302]&m[303]&m[304]))&UnbiasedRNG[28])|((m[298]&~m[301]&~m[302]&m[303]&~m[304])|(~m[298]&~m[301]&~m[302]&~m[303]&m[304])|(m[298]&~m[301]&~m[302]&~m[303]&m[304])|(m[298]&m[301]&~m[302]&~m[303]&m[304])|(m[298]&~m[301]&m[302]&~m[303]&m[304])|(~m[298]&~m[301]&~m[302]&m[303]&m[304])|(m[298]&~m[301]&~m[302]&m[303]&m[304])|(~m[298]&m[301]&~m[302]&m[303]&m[304])|(m[298]&m[301]&~m[302]&m[303]&m[304])|(~m[298]&~m[301]&m[302]&m[303]&m[304])|(m[298]&~m[301]&m[302]&m[303]&m[304])|(m[298]&m[301]&m[302]&m[303]&m[304]));
    m[305] = (((m[303]&~m[306]&~m[307]&~m[308]&~m[309])|(~m[303]&~m[306]&~m[307]&m[308]&~m[309])|(m[303]&m[306]&~m[307]&m[308]&~m[309])|(m[303]&~m[306]&m[307]&m[308]&~m[309])|(~m[303]&m[306]&~m[307]&~m[308]&m[309])|(~m[303]&~m[306]&m[307]&~m[308]&m[309])|(m[303]&m[306]&m[307]&~m[308]&m[309])|(~m[303]&m[306]&m[307]&m[308]&m[309]))&UnbiasedRNG[29])|((m[303]&~m[306]&~m[307]&m[308]&~m[309])|(~m[303]&~m[306]&~m[307]&~m[308]&m[309])|(m[303]&~m[306]&~m[307]&~m[308]&m[309])|(m[303]&m[306]&~m[307]&~m[308]&m[309])|(m[303]&~m[306]&m[307]&~m[308]&m[309])|(~m[303]&~m[306]&~m[307]&m[308]&m[309])|(m[303]&~m[306]&~m[307]&m[308]&m[309])|(~m[303]&m[306]&~m[307]&m[308]&m[309])|(m[303]&m[306]&~m[307]&m[308]&m[309])|(~m[303]&~m[306]&m[307]&m[308]&m[309])|(m[303]&~m[306]&m[307]&m[308]&m[309])|(m[303]&m[306]&m[307]&m[308]&m[309]));
    m[310] = (((m[308]&~m[311]&~m[312]&~m[313]&~m[314])|(~m[308]&~m[311]&~m[312]&m[313]&~m[314])|(m[308]&m[311]&~m[312]&m[313]&~m[314])|(m[308]&~m[311]&m[312]&m[313]&~m[314])|(~m[308]&m[311]&~m[312]&~m[313]&m[314])|(~m[308]&~m[311]&m[312]&~m[313]&m[314])|(m[308]&m[311]&m[312]&~m[313]&m[314])|(~m[308]&m[311]&m[312]&m[313]&m[314]))&UnbiasedRNG[30])|((m[308]&~m[311]&~m[312]&m[313]&~m[314])|(~m[308]&~m[311]&~m[312]&~m[313]&m[314])|(m[308]&~m[311]&~m[312]&~m[313]&m[314])|(m[308]&m[311]&~m[312]&~m[313]&m[314])|(m[308]&~m[311]&m[312]&~m[313]&m[314])|(~m[308]&~m[311]&~m[312]&m[313]&m[314])|(m[308]&~m[311]&~m[312]&m[313]&m[314])|(~m[308]&m[311]&~m[312]&m[313]&m[314])|(m[308]&m[311]&~m[312]&m[313]&m[314])|(~m[308]&~m[311]&m[312]&m[313]&m[314])|(m[308]&~m[311]&m[312]&m[313]&m[314])|(m[308]&m[311]&m[312]&m[313]&m[314]));
    m[315] = (((m[182]&~m[316]&~m[317]&~m[318]&~m[319])|(~m[182]&~m[316]&~m[317]&m[318]&~m[319])|(m[182]&m[316]&~m[317]&m[318]&~m[319])|(m[182]&~m[316]&m[317]&m[318]&~m[319])|(~m[182]&m[316]&~m[317]&~m[318]&m[319])|(~m[182]&~m[316]&m[317]&~m[318]&m[319])|(m[182]&m[316]&m[317]&~m[318]&m[319])|(~m[182]&m[316]&m[317]&m[318]&m[319]))&UnbiasedRNG[31])|((m[182]&~m[316]&~m[317]&m[318]&~m[319])|(~m[182]&~m[316]&~m[317]&~m[318]&m[319])|(m[182]&~m[316]&~m[317]&~m[318]&m[319])|(m[182]&m[316]&~m[317]&~m[318]&m[319])|(m[182]&~m[316]&m[317]&~m[318]&m[319])|(~m[182]&~m[316]&~m[317]&m[318]&m[319])|(m[182]&~m[316]&~m[317]&m[318]&m[319])|(~m[182]&m[316]&~m[317]&m[318]&m[319])|(m[182]&m[316]&~m[317]&m[318]&m[319])|(~m[182]&~m[316]&m[317]&m[318]&m[319])|(m[182]&~m[316]&m[317]&m[318]&m[319])|(m[182]&m[316]&m[317]&m[318]&m[319]));
    m[320] = (((m[318]&~m[321]&~m[322]&~m[323]&~m[324])|(~m[318]&~m[321]&~m[322]&m[323]&~m[324])|(m[318]&m[321]&~m[322]&m[323]&~m[324])|(m[318]&~m[321]&m[322]&m[323]&~m[324])|(~m[318]&m[321]&~m[322]&~m[323]&m[324])|(~m[318]&~m[321]&m[322]&~m[323]&m[324])|(m[318]&m[321]&m[322]&~m[323]&m[324])|(~m[318]&m[321]&m[322]&m[323]&m[324]))&UnbiasedRNG[32])|((m[318]&~m[321]&~m[322]&m[323]&~m[324])|(~m[318]&~m[321]&~m[322]&~m[323]&m[324])|(m[318]&~m[321]&~m[322]&~m[323]&m[324])|(m[318]&m[321]&~m[322]&~m[323]&m[324])|(m[318]&~m[321]&m[322]&~m[323]&m[324])|(~m[318]&~m[321]&~m[322]&m[323]&m[324])|(m[318]&~m[321]&~m[322]&m[323]&m[324])|(~m[318]&m[321]&~m[322]&m[323]&m[324])|(m[318]&m[321]&~m[322]&m[323]&m[324])|(~m[318]&~m[321]&m[322]&m[323]&m[324])|(m[318]&~m[321]&m[322]&m[323]&m[324])|(m[318]&m[321]&m[322]&m[323]&m[324]));
    m[325] = (((m[323]&~m[326]&~m[327]&~m[328]&~m[329])|(~m[323]&~m[326]&~m[327]&m[328]&~m[329])|(m[323]&m[326]&~m[327]&m[328]&~m[329])|(m[323]&~m[326]&m[327]&m[328]&~m[329])|(~m[323]&m[326]&~m[327]&~m[328]&m[329])|(~m[323]&~m[326]&m[327]&~m[328]&m[329])|(m[323]&m[326]&m[327]&~m[328]&m[329])|(~m[323]&m[326]&m[327]&m[328]&m[329]))&UnbiasedRNG[33])|((m[323]&~m[326]&~m[327]&m[328]&~m[329])|(~m[323]&~m[326]&~m[327]&~m[328]&m[329])|(m[323]&~m[326]&~m[327]&~m[328]&m[329])|(m[323]&m[326]&~m[327]&~m[328]&m[329])|(m[323]&~m[326]&m[327]&~m[328]&m[329])|(~m[323]&~m[326]&~m[327]&m[328]&m[329])|(m[323]&~m[326]&~m[327]&m[328]&m[329])|(~m[323]&m[326]&~m[327]&m[328]&m[329])|(m[323]&m[326]&~m[327]&m[328]&m[329])|(~m[323]&~m[326]&m[327]&m[328]&m[329])|(m[323]&~m[326]&m[327]&m[328]&m[329])|(m[323]&m[326]&m[327]&m[328]&m[329]));
    m[330] = (((m[328]&~m[331]&~m[332]&~m[333]&~m[334])|(~m[328]&~m[331]&~m[332]&m[333]&~m[334])|(m[328]&m[331]&~m[332]&m[333]&~m[334])|(m[328]&~m[331]&m[332]&m[333]&~m[334])|(~m[328]&m[331]&~m[332]&~m[333]&m[334])|(~m[328]&~m[331]&m[332]&~m[333]&m[334])|(m[328]&m[331]&m[332]&~m[333]&m[334])|(~m[328]&m[331]&m[332]&m[333]&m[334]))&UnbiasedRNG[34])|((m[328]&~m[331]&~m[332]&m[333]&~m[334])|(~m[328]&~m[331]&~m[332]&~m[333]&m[334])|(m[328]&~m[331]&~m[332]&~m[333]&m[334])|(m[328]&m[331]&~m[332]&~m[333]&m[334])|(m[328]&~m[331]&m[332]&~m[333]&m[334])|(~m[328]&~m[331]&~m[332]&m[333]&m[334])|(m[328]&~m[331]&~m[332]&m[333]&m[334])|(~m[328]&m[331]&~m[332]&m[333]&m[334])|(m[328]&m[331]&~m[332]&m[333]&m[334])|(~m[328]&~m[331]&m[332]&m[333]&m[334])|(m[328]&~m[331]&m[332]&m[333]&m[334])|(m[328]&m[331]&m[332]&m[333]&m[334]));
    m[335] = (((m[333]&~m[336]&~m[337]&~m[338]&~m[339])|(~m[333]&~m[336]&~m[337]&m[338]&~m[339])|(m[333]&m[336]&~m[337]&m[338]&~m[339])|(m[333]&~m[336]&m[337]&m[338]&~m[339])|(~m[333]&m[336]&~m[337]&~m[338]&m[339])|(~m[333]&~m[336]&m[337]&~m[338]&m[339])|(m[333]&m[336]&m[337]&~m[338]&m[339])|(~m[333]&m[336]&m[337]&m[338]&m[339]))&UnbiasedRNG[35])|((m[333]&~m[336]&~m[337]&m[338]&~m[339])|(~m[333]&~m[336]&~m[337]&~m[338]&m[339])|(m[333]&~m[336]&~m[337]&~m[338]&m[339])|(m[333]&m[336]&~m[337]&~m[338]&m[339])|(m[333]&~m[336]&m[337]&~m[338]&m[339])|(~m[333]&~m[336]&~m[337]&m[338]&m[339])|(m[333]&~m[336]&~m[337]&m[338]&m[339])|(~m[333]&m[336]&~m[337]&m[338]&m[339])|(m[333]&m[336]&~m[337]&m[338]&m[339])|(~m[333]&~m[336]&m[337]&m[338]&m[339])|(m[333]&~m[336]&m[337]&m[338]&m[339])|(m[333]&m[336]&m[337]&m[338]&m[339]));
    m[340] = (((m[338]&~m[341]&~m[342]&~m[343]&~m[344])|(~m[338]&~m[341]&~m[342]&m[343]&~m[344])|(m[338]&m[341]&~m[342]&m[343]&~m[344])|(m[338]&~m[341]&m[342]&m[343]&~m[344])|(~m[338]&m[341]&~m[342]&~m[343]&m[344])|(~m[338]&~m[341]&m[342]&~m[343]&m[344])|(m[338]&m[341]&m[342]&~m[343]&m[344])|(~m[338]&m[341]&m[342]&m[343]&m[344]))&UnbiasedRNG[36])|((m[338]&~m[341]&~m[342]&m[343]&~m[344])|(~m[338]&~m[341]&~m[342]&~m[343]&m[344])|(m[338]&~m[341]&~m[342]&~m[343]&m[344])|(m[338]&m[341]&~m[342]&~m[343]&m[344])|(m[338]&~m[341]&m[342]&~m[343]&m[344])|(~m[338]&~m[341]&~m[342]&m[343]&m[344])|(m[338]&~m[341]&~m[342]&m[343]&m[344])|(~m[338]&m[341]&~m[342]&m[343]&m[344])|(m[338]&m[341]&~m[342]&m[343]&m[344])|(~m[338]&~m[341]&m[342]&m[343]&m[344])|(m[338]&~m[341]&m[342]&m[343]&m[344])|(m[338]&m[341]&m[342]&m[343]&m[344]));
    m[345] = (((m[183]&~m[346]&~m[347]&~m[348]&~m[349])|(~m[183]&~m[346]&~m[347]&m[348]&~m[349])|(m[183]&m[346]&~m[347]&m[348]&~m[349])|(m[183]&~m[346]&m[347]&m[348]&~m[349])|(~m[183]&m[346]&~m[347]&~m[348]&m[349])|(~m[183]&~m[346]&m[347]&~m[348]&m[349])|(m[183]&m[346]&m[347]&~m[348]&m[349])|(~m[183]&m[346]&m[347]&m[348]&m[349]))&UnbiasedRNG[37])|((m[183]&~m[346]&~m[347]&m[348]&~m[349])|(~m[183]&~m[346]&~m[347]&~m[348]&m[349])|(m[183]&~m[346]&~m[347]&~m[348]&m[349])|(m[183]&m[346]&~m[347]&~m[348]&m[349])|(m[183]&~m[346]&m[347]&~m[348]&m[349])|(~m[183]&~m[346]&~m[347]&m[348]&m[349])|(m[183]&~m[346]&~m[347]&m[348]&m[349])|(~m[183]&m[346]&~m[347]&m[348]&m[349])|(m[183]&m[346]&~m[347]&m[348]&m[349])|(~m[183]&~m[346]&m[347]&m[348]&m[349])|(m[183]&~m[346]&m[347]&m[348]&m[349])|(m[183]&m[346]&m[347]&m[348]&m[349]));
    m[350] = (((m[348]&~m[351]&~m[352]&~m[353]&~m[354])|(~m[348]&~m[351]&~m[352]&m[353]&~m[354])|(m[348]&m[351]&~m[352]&m[353]&~m[354])|(m[348]&~m[351]&m[352]&m[353]&~m[354])|(~m[348]&m[351]&~m[352]&~m[353]&m[354])|(~m[348]&~m[351]&m[352]&~m[353]&m[354])|(m[348]&m[351]&m[352]&~m[353]&m[354])|(~m[348]&m[351]&m[352]&m[353]&m[354]))&UnbiasedRNG[38])|((m[348]&~m[351]&~m[352]&m[353]&~m[354])|(~m[348]&~m[351]&~m[352]&~m[353]&m[354])|(m[348]&~m[351]&~m[352]&~m[353]&m[354])|(m[348]&m[351]&~m[352]&~m[353]&m[354])|(m[348]&~m[351]&m[352]&~m[353]&m[354])|(~m[348]&~m[351]&~m[352]&m[353]&m[354])|(m[348]&~m[351]&~m[352]&m[353]&m[354])|(~m[348]&m[351]&~m[352]&m[353]&m[354])|(m[348]&m[351]&~m[352]&m[353]&m[354])|(~m[348]&~m[351]&m[352]&m[353]&m[354])|(m[348]&~m[351]&m[352]&m[353]&m[354])|(m[348]&m[351]&m[352]&m[353]&m[354]));
    m[355] = (((m[353]&~m[356]&~m[357]&~m[358]&~m[359])|(~m[353]&~m[356]&~m[357]&m[358]&~m[359])|(m[353]&m[356]&~m[357]&m[358]&~m[359])|(m[353]&~m[356]&m[357]&m[358]&~m[359])|(~m[353]&m[356]&~m[357]&~m[358]&m[359])|(~m[353]&~m[356]&m[357]&~m[358]&m[359])|(m[353]&m[356]&m[357]&~m[358]&m[359])|(~m[353]&m[356]&m[357]&m[358]&m[359]))&UnbiasedRNG[39])|((m[353]&~m[356]&~m[357]&m[358]&~m[359])|(~m[353]&~m[356]&~m[357]&~m[358]&m[359])|(m[353]&~m[356]&~m[357]&~m[358]&m[359])|(m[353]&m[356]&~m[357]&~m[358]&m[359])|(m[353]&~m[356]&m[357]&~m[358]&m[359])|(~m[353]&~m[356]&~m[357]&m[358]&m[359])|(m[353]&~m[356]&~m[357]&m[358]&m[359])|(~m[353]&m[356]&~m[357]&m[358]&m[359])|(m[353]&m[356]&~m[357]&m[358]&m[359])|(~m[353]&~m[356]&m[357]&m[358]&m[359])|(m[353]&~m[356]&m[357]&m[358]&m[359])|(m[353]&m[356]&m[357]&m[358]&m[359]));
    m[360] = (((m[358]&~m[361]&~m[362]&~m[363]&~m[364])|(~m[358]&~m[361]&~m[362]&m[363]&~m[364])|(m[358]&m[361]&~m[362]&m[363]&~m[364])|(m[358]&~m[361]&m[362]&m[363]&~m[364])|(~m[358]&m[361]&~m[362]&~m[363]&m[364])|(~m[358]&~m[361]&m[362]&~m[363]&m[364])|(m[358]&m[361]&m[362]&~m[363]&m[364])|(~m[358]&m[361]&m[362]&m[363]&m[364]))&UnbiasedRNG[40])|((m[358]&~m[361]&~m[362]&m[363]&~m[364])|(~m[358]&~m[361]&~m[362]&~m[363]&m[364])|(m[358]&~m[361]&~m[362]&~m[363]&m[364])|(m[358]&m[361]&~m[362]&~m[363]&m[364])|(m[358]&~m[361]&m[362]&~m[363]&m[364])|(~m[358]&~m[361]&~m[362]&m[363]&m[364])|(m[358]&~m[361]&~m[362]&m[363]&m[364])|(~m[358]&m[361]&~m[362]&m[363]&m[364])|(m[358]&m[361]&~m[362]&m[363]&m[364])|(~m[358]&~m[361]&m[362]&m[363]&m[364])|(m[358]&~m[361]&m[362]&m[363]&m[364])|(m[358]&m[361]&m[362]&m[363]&m[364]));
    m[365] = (((m[363]&~m[366]&~m[367]&~m[368]&~m[369])|(~m[363]&~m[366]&~m[367]&m[368]&~m[369])|(m[363]&m[366]&~m[367]&m[368]&~m[369])|(m[363]&~m[366]&m[367]&m[368]&~m[369])|(~m[363]&m[366]&~m[367]&~m[368]&m[369])|(~m[363]&~m[366]&m[367]&~m[368]&m[369])|(m[363]&m[366]&m[367]&~m[368]&m[369])|(~m[363]&m[366]&m[367]&m[368]&m[369]))&UnbiasedRNG[41])|((m[363]&~m[366]&~m[367]&m[368]&~m[369])|(~m[363]&~m[366]&~m[367]&~m[368]&m[369])|(m[363]&~m[366]&~m[367]&~m[368]&m[369])|(m[363]&m[366]&~m[367]&~m[368]&m[369])|(m[363]&~m[366]&m[367]&~m[368]&m[369])|(~m[363]&~m[366]&~m[367]&m[368]&m[369])|(m[363]&~m[366]&~m[367]&m[368]&m[369])|(~m[363]&m[366]&~m[367]&m[368]&m[369])|(m[363]&m[366]&~m[367]&m[368]&m[369])|(~m[363]&~m[366]&m[367]&m[368]&m[369])|(m[363]&~m[366]&m[367]&m[368]&m[369])|(m[363]&m[366]&m[367]&m[368]&m[369]));
    m[370] = (((m[368]&~m[371]&~m[372]&~m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&m[373]&~m[374])|(m[368]&m[371]&~m[372]&m[373]&~m[374])|(m[368]&~m[371]&m[372]&m[373]&~m[374])|(~m[368]&m[371]&~m[372]&~m[373]&m[374])|(~m[368]&~m[371]&m[372]&~m[373]&m[374])|(m[368]&m[371]&m[372]&~m[373]&m[374])|(~m[368]&m[371]&m[372]&m[373]&m[374]))&UnbiasedRNG[42])|((m[368]&~m[371]&~m[372]&m[373]&~m[374])|(~m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&~m[372]&~m[373]&m[374])|(m[368]&m[371]&~m[372]&~m[373]&m[374])|(m[368]&~m[371]&m[372]&~m[373]&m[374])|(~m[368]&~m[371]&~m[372]&m[373]&m[374])|(m[368]&~m[371]&~m[372]&m[373]&m[374])|(~m[368]&m[371]&~m[372]&m[373]&m[374])|(m[368]&m[371]&~m[372]&m[373]&m[374])|(~m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&~m[371]&m[372]&m[373]&m[374])|(m[368]&m[371]&m[372]&m[373]&m[374]));
    m[375] = (((m[373]&~m[376]&~m[377]&~m[378]&~m[379])|(~m[373]&~m[376]&~m[377]&m[378]&~m[379])|(m[373]&m[376]&~m[377]&m[378]&~m[379])|(m[373]&~m[376]&m[377]&m[378]&~m[379])|(~m[373]&m[376]&~m[377]&~m[378]&m[379])|(~m[373]&~m[376]&m[377]&~m[378]&m[379])|(m[373]&m[376]&m[377]&~m[378]&m[379])|(~m[373]&m[376]&m[377]&m[378]&m[379]))&UnbiasedRNG[43])|((m[373]&~m[376]&~m[377]&m[378]&~m[379])|(~m[373]&~m[376]&~m[377]&~m[378]&m[379])|(m[373]&~m[376]&~m[377]&~m[378]&m[379])|(m[373]&m[376]&~m[377]&~m[378]&m[379])|(m[373]&~m[376]&m[377]&~m[378]&m[379])|(~m[373]&~m[376]&~m[377]&m[378]&m[379])|(m[373]&~m[376]&~m[377]&m[378]&m[379])|(~m[373]&m[376]&~m[377]&m[378]&m[379])|(m[373]&m[376]&~m[377]&m[378]&m[379])|(~m[373]&~m[376]&m[377]&m[378]&m[379])|(m[373]&~m[376]&m[377]&m[378]&m[379])|(m[373]&m[376]&m[377]&m[378]&m[379]));
    m[385] = (((m[383]&~m[386]&~m[387]&~m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&m[388]&~m[389])|(m[383]&m[386]&~m[387]&m[388]&~m[389])|(m[383]&~m[386]&m[387]&m[388]&~m[389])|(~m[383]&m[386]&~m[387]&~m[388]&m[389])|(~m[383]&~m[386]&m[387]&~m[388]&m[389])|(m[383]&m[386]&m[387]&~m[388]&m[389])|(~m[383]&m[386]&m[387]&m[388]&m[389]))&UnbiasedRNG[44])|((m[383]&~m[386]&~m[387]&m[388]&~m[389])|(~m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&~m[387]&~m[388]&m[389])|(m[383]&m[386]&~m[387]&~m[388]&m[389])|(m[383]&~m[386]&m[387]&~m[388]&m[389])|(~m[383]&~m[386]&~m[387]&m[388]&m[389])|(m[383]&~m[386]&~m[387]&m[388]&m[389])|(~m[383]&m[386]&~m[387]&m[388]&m[389])|(m[383]&m[386]&~m[387]&m[388]&m[389])|(~m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&~m[386]&m[387]&m[388]&m[389])|(m[383]&m[386]&m[387]&m[388]&m[389]));
    m[390] = (((m[388]&~m[391]&~m[392]&~m[393]&~m[394])|(~m[388]&~m[391]&~m[392]&m[393]&~m[394])|(m[388]&m[391]&~m[392]&m[393]&~m[394])|(m[388]&~m[391]&m[392]&m[393]&~m[394])|(~m[388]&m[391]&~m[392]&~m[393]&m[394])|(~m[388]&~m[391]&m[392]&~m[393]&m[394])|(m[388]&m[391]&m[392]&~m[393]&m[394])|(~m[388]&m[391]&m[392]&m[393]&m[394]))&UnbiasedRNG[45])|((m[388]&~m[391]&~m[392]&m[393]&~m[394])|(~m[388]&~m[391]&~m[392]&~m[393]&m[394])|(m[388]&~m[391]&~m[392]&~m[393]&m[394])|(m[388]&m[391]&~m[392]&~m[393]&m[394])|(m[388]&~m[391]&m[392]&~m[393]&m[394])|(~m[388]&~m[391]&~m[392]&m[393]&m[394])|(m[388]&~m[391]&~m[392]&m[393]&m[394])|(~m[388]&m[391]&~m[392]&m[393]&m[394])|(m[388]&m[391]&~m[392]&m[393]&m[394])|(~m[388]&~m[391]&m[392]&m[393]&m[394])|(m[388]&~m[391]&m[392]&m[393]&m[394])|(m[388]&m[391]&m[392]&m[393]&m[394]));
    m[395] = (((m[393]&~m[396]&~m[397]&~m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&m[398]&~m[399])|(m[393]&m[396]&~m[397]&m[398]&~m[399])|(m[393]&~m[396]&m[397]&m[398]&~m[399])|(~m[393]&m[396]&~m[397]&~m[398]&m[399])|(~m[393]&~m[396]&m[397]&~m[398]&m[399])|(m[393]&m[396]&m[397]&~m[398]&m[399])|(~m[393]&m[396]&m[397]&m[398]&m[399]))&UnbiasedRNG[46])|((m[393]&~m[396]&~m[397]&m[398]&~m[399])|(~m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&~m[397]&~m[398]&m[399])|(m[393]&m[396]&~m[397]&~m[398]&m[399])|(m[393]&~m[396]&m[397]&~m[398]&m[399])|(~m[393]&~m[396]&~m[397]&m[398]&m[399])|(m[393]&~m[396]&~m[397]&m[398]&m[399])|(~m[393]&m[396]&~m[397]&m[398]&m[399])|(m[393]&m[396]&~m[397]&m[398]&m[399])|(~m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&~m[396]&m[397]&m[398]&m[399])|(m[393]&m[396]&m[397]&m[398]&m[399]));
    m[400] = (((m[398]&~m[401]&~m[402]&~m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&m[403]&~m[404])|(m[398]&m[401]&~m[402]&m[403]&~m[404])|(m[398]&~m[401]&m[402]&m[403]&~m[404])|(~m[398]&m[401]&~m[402]&~m[403]&m[404])|(~m[398]&~m[401]&m[402]&~m[403]&m[404])|(m[398]&m[401]&m[402]&~m[403]&m[404])|(~m[398]&m[401]&m[402]&m[403]&m[404]))&UnbiasedRNG[47])|((m[398]&~m[401]&~m[402]&m[403]&~m[404])|(~m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&~m[402]&~m[403]&m[404])|(m[398]&m[401]&~m[402]&~m[403]&m[404])|(m[398]&~m[401]&m[402]&~m[403]&m[404])|(~m[398]&~m[401]&~m[402]&m[403]&m[404])|(m[398]&~m[401]&~m[402]&m[403]&m[404])|(~m[398]&m[401]&~m[402]&m[403]&m[404])|(m[398]&m[401]&~m[402]&m[403]&m[404])|(~m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&~m[401]&m[402]&m[403]&m[404])|(m[398]&m[401]&m[402]&m[403]&m[404]));
    m[405] = (((m[403]&~m[406]&~m[407]&~m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&m[408]&~m[409])|(m[403]&m[406]&~m[407]&m[408]&~m[409])|(m[403]&~m[406]&m[407]&m[408]&~m[409])|(~m[403]&m[406]&~m[407]&~m[408]&m[409])|(~m[403]&~m[406]&m[407]&~m[408]&m[409])|(m[403]&m[406]&m[407]&~m[408]&m[409])|(~m[403]&m[406]&m[407]&m[408]&m[409]))&UnbiasedRNG[48])|((m[403]&~m[406]&~m[407]&m[408]&~m[409])|(~m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&~m[407]&~m[408]&m[409])|(m[403]&m[406]&~m[407]&~m[408]&m[409])|(m[403]&~m[406]&m[407]&~m[408]&m[409])|(~m[403]&~m[406]&~m[407]&m[408]&m[409])|(m[403]&~m[406]&~m[407]&m[408]&m[409])|(~m[403]&m[406]&~m[407]&m[408]&m[409])|(m[403]&m[406]&~m[407]&m[408]&m[409])|(~m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&~m[406]&m[407]&m[408]&m[409])|(m[403]&m[406]&m[407]&m[408]&m[409]));
    m[410] = (((m[408]&~m[411]&~m[412]&~m[413]&~m[414])|(~m[408]&~m[411]&~m[412]&m[413]&~m[414])|(m[408]&m[411]&~m[412]&m[413]&~m[414])|(m[408]&~m[411]&m[412]&m[413]&~m[414])|(~m[408]&m[411]&~m[412]&~m[413]&m[414])|(~m[408]&~m[411]&m[412]&~m[413]&m[414])|(m[408]&m[411]&m[412]&~m[413]&m[414])|(~m[408]&m[411]&m[412]&m[413]&m[414]))&UnbiasedRNG[49])|((m[408]&~m[411]&~m[412]&m[413]&~m[414])|(~m[408]&~m[411]&~m[412]&~m[413]&m[414])|(m[408]&~m[411]&~m[412]&~m[413]&m[414])|(m[408]&m[411]&~m[412]&~m[413]&m[414])|(m[408]&~m[411]&m[412]&~m[413]&m[414])|(~m[408]&~m[411]&~m[412]&m[413]&m[414])|(m[408]&~m[411]&~m[412]&m[413]&m[414])|(~m[408]&m[411]&~m[412]&m[413]&m[414])|(m[408]&m[411]&~m[412]&m[413]&m[414])|(~m[408]&~m[411]&m[412]&m[413]&m[414])|(m[408]&~m[411]&m[412]&m[413]&m[414])|(m[408]&m[411]&m[412]&m[413]&m[414]));
    m[415] = (((m[384]&~m[416]&~m[417]&~m[418]&~m[419])|(~m[384]&~m[416]&~m[417]&m[418]&~m[419])|(m[384]&m[416]&~m[417]&m[418]&~m[419])|(m[384]&~m[416]&m[417]&m[418]&~m[419])|(~m[384]&m[416]&~m[417]&~m[418]&m[419])|(~m[384]&~m[416]&m[417]&~m[418]&m[419])|(m[384]&m[416]&m[417]&~m[418]&m[419])|(~m[384]&m[416]&m[417]&m[418]&m[419]))&UnbiasedRNG[50])|((m[384]&~m[416]&~m[417]&m[418]&~m[419])|(~m[384]&~m[416]&~m[417]&~m[418]&m[419])|(m[384]&~m[416]&~m[417]&~m[418]&m[419])|(m[384]&m[416]&~m[417]&~m[418]&m[419])|(m[384]&~m[416]&m[417]&~m[418]&m[419])|(~m[384]&~m[416]&~m[417]&m[418]&m[419])|(m[384]&~m[416]&~m[417]&m[418]&m[419])|(~m[384]&m[416]&~m[417]&m[418]&m[419])|(m[384]&m[416]&~m[417]&m[418]&m[419])|(~m[384]&~m[416]&m[417]&m[418]&m[419])|(m[384]&~m[416]&m[417]&m[418]&m[419])|(m[384]&m[416]&m[417]&m[418]&m[419]));
    m[420] = (((m[418]&~m[421]&~m[422]&~m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&m[423]&~m[424])|(m[418]&m[421]&~m[422]&m[423]&~m[424])|(m[418]&~m[421]&m[422]&m[423]&~m[424])|(~m[418]&m[421]&~m[422]&~m[423]&m[424])|(~m[418]&~m[421]&m[422]&~m[423]&m[424])|(m[418]&m[421]&m[422]&~m[423]&m[424])|(~m[418]&m[421]&m[422]&m[423]&m[424]))&UnbiasedRNG[51])|((m[418]&~m[421]&~m[422]&m[423]&~m[424])|(~m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&~m[422]&~m[423]&m[424])|(m[418]&m[421]&~m[422]&~m[423]&m[424])|(m[418]&~m[421]&m[422]&~m[423]&m[424])|(~m[418]&~m[421]&~m[422]&m[423]&m[424])|(m[418]&~m[421]&~m[422]&m[423]&m[424])|(~m[418]&m[421]&~m[422]&m[423]&m[424])|(m[418]&m[421]&~m[422]&m[423]&m[424])|(~m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&~m[421]&m[422]&m[423]&m[424])|(m[418]&m[421]&m[422]&m[423]&m[424]));
    m[425] = (((m[423]&~m[426]&~m[427]&~m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&m[428]&~m[429])|(m[423]&m[426]&~m[427]&m[428]&~m[429])|(m[423]&~m[426]&m[427]&m[428]&~m[429])|(~m[423]&m[426]&~m[427]&~m[428]&m[429])|(~m[423]&~m[426]&m[427]&~m[428]&m[429])|(m[423]&m[426]&m[427]&~m[428]&m[429])|(~m[423]&m[426]&m[427]&m[428]&m[429]))&UnbiasedRNG[52])|((m[423]&~m[426]&~m[427]&m[428]&~m[429])|(~m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&~m[427]&~m[428]&m[429])|(m[423]&m[426]&~m[427]&~m[428]&m[429])|(m[423]&~m[426]&m[427]&~m[428]&m[429])|(~m[423]&~m[426]&~m[427]&m[428]&m[429])|(m[423]&~m[426]&~m[427]&m[428]&m[429])|(~m[423]&m[426]&~m[427]&m[428]&m[429])|(m[423]&m[426]&~m[427]&m[428]&m[429])|(~m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&~m[426]&m[427]&m[428]&m[429])|(m[423]&m[426]&m[427]&m[428]&m[429]));
    m[430] = (((m[428]&~m[431]&~m[432]&~m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&m[433]&~m[434])|(m[428]&m[431]&~m[432]&m[433]&~m[434])|(m[428]&~m[431]&m[432]&m[433]&~m[434])|(~m[428]&m[431]&~m[432]&~m[433]&m[434])|(~m[428]&~m[431]&m[432]&~m[433]&m[434])|(m[428]&m[431]&m[432]&~m[433]&m[434])|(~m[428]&m[431]&m[432]&m[433]&m[434]))&UnbiasedRNG[53])|((m[428]&~m[431]&~m[432]&m[433]&~m[434])|(~m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&~m[432]&~m[433]&m[434])|(m[428]&m[431]&~m[432]&~m[433]&m[434])|(m[428]&~m[431]&m[432]&~m[433]&m[434])|(~m[428]&~m[431]&~m[432]&m[433]&m[434])|(m[428]&~m[431]&~m[432]&m[433]&m[434])|(~m[428]&m[431]&~m[432]&m[433]&m[434])|(m[428]&m[431]&~m[432]&m[433]&m[434])|(~m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&~m[431]&m[432]&m[433]&m[434])|(m[428]&m[431]&m[432]&m[433]&m[434]));
    m[435] = (((m[433]&~m[436]&~m[437]&~m[438]&~m[439])|(~m[433]&~m[436]&~m[437]&m[438]&~m[439])|(m[433]&m[436]&~m[437]&m[438]&~m[439])|(m[433]&~m[436]&m[437]&m[438]&~m[439])|(~m[433]&m[436]&~m[437]&~m[438]&m[439])|(~m[433]&~m[436]&m[437]&~m[438]&m[439])|(m[433]&m[436]&m[437]&~m[438]&m[439])|(~m[433]&m[436]&m[437]&m[438]&m[439]))&UnbiasedRNG[54])|((m[433]&~m[436]&~m[437]&m[438]&~m[439])|(~m[433]&~m[436]&~m[437]&~m[438]&m[439])|(m[433]&~m[436]&~m[437]&~m[438]&m[439])|(m[433]&m[436]&~m[437]&~m[438]&m[439])|(m[433]&~m[436]&m[437]&~m[438]&m[439])|(~m[433]&~m[436]&~m[437]&m[438]&m[439])|(m[433]&~m[436]&~m[437]&m[438]&m[439])|(~m[433]&m[436]&~m[437]&m[438]&m[439])|(m[433]&m[436]&~m[437]&m[438]&m[439])|(~m[433]&~m[436]&m[437]&m[438]&m[439])|(m[433]&~m[436]&m[437]&m[438]&m[439])|(m[433]&m[436]&m[437]&m[438]&m[439]));
    m[440] = (((m[438]&~m[441]&~m[442]&~m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&m[443]&~m[444])|(m[438]&m[441]&~m[442]&m[443]&~m[444])|(m[438]&~m[441]&m[442]&m[443]&~m[444])|(~m[438]&m[441]&~m[442]&~m[443]&m[444])|(~m[438]&~m[441]&m[442]&~m[443]&m[444])|(m[438]&m[441]&m[442]&~m[443]&m[444])|(~m[438]&m[441]&m[442]&m[443]&m[444]))&UnbiasedRNG[55])|((m[438]&~m[441]&~m[442]&m[443]&~m[444])|(~m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&~m[442]&~m[443]&m[444])|(m[438]&m[441]&~m[442]&~m[443]&m[444])|(m[438]&~m[441]&m[442]&~m[443]&m[444])|(~m[438]&~m[441]&~m[442]&m[443]&m[444])|(m[438]&~m[441]&~m[442]&m[443]&m[444])|(~m[438]&m[441]&~m[442]&m[443]&m[444])|(m[438]&m[441]&~m[442]&m[443]&m[444])|(~m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&~m[441]&m[442]&m[443]&m[444])|(m[438]&m[441]&m[442]&m[443]&m[444]));
    m[445] = (((m[419]&~m[446]&~m[447]&~m[448]&~m[449])|(~m[419]&~m[446]&~m[447]&m[448]&~m[449])|(m[419]&m[446]&~m[447]&m[448]&~m[449])|(m[419]&~m[446]&m[447]&m[448]&~m[449])|(~m[419]&m[446]&~m[447]&~m[448]&m[449])|(~m[419]&~m[446]&m[447]&~m[448]&m[449])|(m[419]&m[446]&m[447]&~m[448]&m[449])|(~m[419]&m[446]&m[447]&m[448]&m[449]))&UnbiasedRNG[56])|((m[419]&~m[446]&~m[447]&m[448]&~m[449])|(~m[419]&~m[446]&~m[447]&~m[448]&m[449])|(m[419]&~m[446]&~m[447]&~m[448]&m[449])|(m[419]&m[446]&~m[447]&~m[448]&m[449])|(m[419]&~m[446]&m[447]&~m[448]&m[449])|(~m[419]&~m[446]&~m[447]&m[448]&m[449])|(m[419]&~m[446]&~m[447]&m[448]&m[449])|(~m[419]&m[446]&~m[447]&m[448]&m[449])|(m[419]&m[446]&~m[447]&m[448]&m[449])|(~m[419]&~m[446]&m[447]&m[448]&m[449])|(m[419]&~m[446]&m[447]&m[448]&m[449])|(m[419]&m[446]&m[447]&m[448]&m[449]));
    m[450] = (((m[448]&~m[451]&~m[452]&~m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&m[453]&~m[454])|(m[448]&m[451]&~m[452]&m[453]&~m[454])|(m[448]&~m[451]&m[452]&m[453]&~m[454])|(~m[448]&m[451]&~m[452]&~m[453]&m[454])|(~m[448]&~m[451]&m[452]&~m[453]&m[454])|(m[448]&m[451]&m[452]&~m[453]&m[454])|(~m[448]&m[451]&m[452]&m[453]&m[454]))&UnbiasedRNG[57])|((m[448]&~m[451]&~m[452]&m[453]&~m[454])|(~m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&~m[452]&~m[453]&m[454])|(m[448]&m[451]&~m[452]&~m[453]&m[454])|(m[448]&~m[451]&m[452]&~m[453]&m[454])|(~m[448]&~m[451]&~m[452]&m[453]&m[454])|(m[448]&~m[451]&~m[452]&m[453]&m[454])|(~m[448]&m[451]&~m[452]&m[453]&m[454])|(m[448]&m[451]&~m[452]&m[453]&m[454])|(~m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&~m[451]&m[452]&m[453]&m[454])|(m[448]&m[451]&m[452]&m[453]&m[454]));
    m[455] = (((m[453]&~m[456]&~m[457]&~m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&m[458]&~m[459])|(m[453]&m[456]&~m[457]&m[458]&~m[459])|(m[453]&~m[456]&m[457]&m[458]&~m[459])|(~m[453]&m[456]&~m[457]&~m[458]&m[459])|(~m[453]&~m[456]&m[457]&~m[458]&m[459])|(m[453]&m[456]&m[457]&~m[458]&m[459])|(~m[453]&m[456]&m[457]&m[458]&m[459]))&UnbiasedRNG[58])|((m[453]&~m[456]&~m[457]&m[458]&~m[459])|(~m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&~m[457]&~m[458]&m[459])|(m[453]&m[456]&~m[457]&~m[458]&m[459])|(m[453]&~m[456]&m[457]&~m[458]&m[459])|(~m[453]&~m[456]&~m[457]&m[458]&m[459])|(m[453]&~m[456]&~m[457]&m[458]&m[459])|(~m[453]&m[456]&~m[457]&m[458]&m[459])|(m[453]&m[456]&~m[457]&m[458]&m[459])|(~m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&~m[456]&m[457]&m[458]&m[459])|(m[453]&m[456]&m[457]&m[458]&m[459]));
    m[460] = (((m[458]&~m[461]&~m[462]&~m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&m[463]&~m[464])|(m[458]&m[461]&~m[462]&m[463]&~m[464])|(m[458]&~m[461]&m[462]&m[463]&~m[464])|(~m[458]&m[461]&~m[462]&~m[463]&m[464])|(~m[458]&~m[461]&m[462]&~m[463]&m[464])|(m[458]&m[461]&m[462]&~m[463]&m[464])|(~m[458]&m[461]&m[462]&m[463]&m[464]))&UnbiasedRNG[59])|((m[458]&~m[461]&~m[462]&m[463]&~m[464])|(~m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&~m[462]&~m[463]&m[464])|(m[458]&m[461]&~m[462]&~m[463]&m[464])|(m[458]&~m[461]&m[462]&~m[463]&m[464])|(~m[458]&~m[461]&~m[462]&m[463]&m[464])|(m[458]&~m[461]&~m[462]&m[463]&m[464])|(~m[458]&m[461]&~m[462]&m[463]&m[464])|(m[458]&m[461]&~m[462]&m[463]&m[464])|(~m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&~m[461]&m[462]&m[463]&m[464])|(m[458]&m[461]&m[462]&m[463]&m[464]));
    m[465] = (((m[463]&~m[466]&~m[467]&~m[468]&~m[469])|(~m[463]&~m[466]&~m[467]&m[468]&~m[469])|(m[463]&m[466]&~m[467]&m[468]&~m[469])|(m[463]&~m[466]&m[467]&m[468]&~m[469])|(~m[463]&m[466]&~m[467]&~m[468]&m[469])|(~m[463]&~m[466]&m[467]&~m[468]&m[469])|(m[463]&m[466]&m[467]&~m[468]&m[469])|(~m[463]&m[466]&m[467]&m[468]&m[469]))&UnbiasedRNG[60])|((m[463]&~m[466]&~m[467]&m[468]&~m[469])|(~m[463]&~m[466]&~m[467]&~m[468]&m[469])|(m[463]&~m[466]&~m[467]&~m[468]&m[469])|(m[463]&m[466]&~m[467]&~m[468]&m[469])|(m[463]&~m[466]&m[467]&~m[468]&m[469])|(~m[463]&~m[466]&~m[467]&m[468]&m[469])|(m[463]&~m[466]&~m[467]&m[468]&m[469])|(~m[463]&m[466]&~m[467]&m[468]&m[469])|(m[463]&m[466]&~m[467]&m[468]&m[469])|(~m[463]&~m[466]&m[467]&m[468]&m[469])|(m[463]&~m[466]&m[467]&m[468]&m[469])|(m[463]&m[466]&m[467]&m[468]&m[469]));
    m[470] = (((m[449]&~m[471]&~m[472]&~m[473]&~m[474])|(~m[449]&~m[471]&~m[472]&m[473]&~m[474])|(m[449]&m[471]&~m[472]&m[473]&~m[474])|(m[449]&~m[471]&m[472]&m[473]&~m[474])|(~m[449]&m[471]&~m[472]&~m[473]&m[474])|(~m[449]&~m[471]&m[472]&~m[473]&m[474])|(m[449]&m[471]&m[472]&~m[473]&m[474])|(~m[449]&m[471]&m[472]&m[473]&m[474]))&UnbiasedRNG[61])|((m[449]&~m[471]&~m[472]&m[473]&~m[474])|(~m[449]&~m[471]&~m[472]&~m[473]&m[474])|(m[449]&~m[471]&~m[472]&~m[473]&m[474])|(m[449]&m[471]&~m[472]&~m[473]&m[474])|(m[449]&~m[471]&m[472]&~m[473]&m[474])|(~m[449]&~m[471]&~m[472]&m[473]&m[474])|(m[449]&~m[471]&~m[472]&m[473]&m[474])|(~m[449]&m[471]&~m[472]&m[473]&m[474])|(m[449]&m[471]&~m[472]&m[473]&m[474])|(~m[449]&~m[471]&m[472]&m[473]&m[474])|(m[449]&~m[471]&m[472]&m[473]&m[474])|(m[449]&m[471]&m[472]&m[473]&m[474]));
    m[475] = (((m[473]&~m[476]&~m[477]&~m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&m[478]&~m[479])|(m[473]&m[476]&~m[477]&m[478]&~m[479])|(m[473]&~m[476]&m[477]&m[478]&~m[479])|(~m[473]&m[476]&~m[477]&~m[478]&m[479])|(~m[473]&~m[476]&m[477]&~m[478]&m[479])|(m[473]&m[476]&m[477]&~m[478]&m[479])|(~m[473]&m[476]&m[477]&m[478]&m[479]))&UnbiasedRNG[62])|((m[473]&~m[476]&~m[477]&m[478]&~m[479])|(~m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&~m[477]&~m[478]&m[479])|(m[473]&m[476]&~m[477]&~m[478]&m[479])|(m[473]&~m[476]&m[477]&~m[478]&m[479])|(~m[473]&~m[476]&~m[477]&m[478]&m[479])|(m[473]&~m[476]&~m[477]&m[478]&m[479])|(~m[473]&m[476]&~m[477]&m[478]&m[479])|(m[473]&m[476]&~m[477]&m[478]&m[479])|(~m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&~m[476]&m[477]&m[478]&m[479])|(m[473]&m[476]&m[477]&m[478]&m[479]));
    m[480] = (((m[478]&~m[481]&~m[482]&~m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&m[483]&~m[484])|(m[478]&m[481]&~m[482]&m[483]&~m[484])|(m[478]&~m[481]&m[482]&m[483]&~m[484])|(~m[478]&m[481]&~m[482]&~m[483]&m[484])|(~m[478]&~m[481]&m[482]&~m[483]&m[484])|(m[478]&m[481]&m[482]&~m[483]&m[484])|(~m[478]&m[481]&m[482]&m[483]&m[484]))&UnbiasedRNG[63])|((m[478]&~m[481]&~m[482]&m[483]&~m[484])|(~m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&~m[482]&~m[483]&m[484])|(m[478]&m[481]&~m[482]&~m[483]&m[484])|(m[478]&~m[481]&m[482]&~m[483]&m[484])|(~m[478]&~m[481]&~m[482]&m[483]&m[484])|(m[478]&~m[481]&~m[482]&m[483]&m[484])|(~m[478]&m[481]&~m[482]&m[483]&m[484])|(m[478]&m[481]&~m[482]&m[483]&m[484])|(~m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&~m[481]&m[482]&m[483]&m[484])|(m[478]&m[481]&m[482]&m[483]&m[484]));
    m[485] = (((m[483]&~m[486]&~m[487]&~m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&m[488]&~m[489])|(m[483]&m[486]&~m[487]&m[488]&~m[489])|(m[483]&~m[486]&m[487]&m[488]&~m[489])|(~m[483]&m[486]&~m[487]&~m[488]&m[489])|(~m[483]&~m[486]&m[487]&~m[488]&m[489])|(m[483]&m[486]&m[487]&~m[488]&m[489])|(~m[483]&m[486]&m[487]&m[488]&m[489]))&UnbiasedRNG[64])|((m[483]&~m[486]&~m[487]&m[488]&~m[489])|(~m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&~m[487]&~m[488]&m[489])|(m[483]&m[486]&~m[487]&~m[488]&m[489])|(m[483]&~m[486]&m[487]&~m[488]&m[489])|(~m[483]&~m[486]&~m[487]&m[488]&m[489])|(m[483]&~m[486]&~m[487]&m[488]&m[489])|(~m[483]&m[486]&~m[487]&m[488]&m[489])|(m[483]&m[486]&~m[487]&m[488]&m[489])|(~m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&~m[486]&m[487]&m[488]&m[489])|(m[483]&m[486]&m[487]&m[488]&m[489]));
    m[490] = (((m[474]&~m[491]&~m[492]&~m[493]&~m[494])|(~m[474]&~m[491]&~m[492]&m[493]&~m[494])|(m[474]&m[491]&~m[492]&m[493]&~m[494])|(m[474]&~m[491]&m[492]&m[493]&~m[494])|(~m[474]&m[491]&~m[492]&~m[493]&m[494])|(~m[474]&~m[491]&m[492]&~m[493]&m[494])|(m[474]&m[491]&m[492]&~m[493]&m[494])|(~m[474]&m[491]&m[492]&m[493]&m[494]))&UnbiasedRNG[65])|((m[474]&~m[491]&~m[492]&m[493]&~m[494])|(~m[474]&~m[491]&~m[492]&~m[493]&m[494])|(m[474]&~m[491]&~m[492]&~m[493]&m[494])|(m[474]&m[491]&~m[492]&~m[493]&m[494])|(m[474]&~m[491]&m[492]&~m[493]&m[494])|(~m[474]&~m[491]&~m[492]&m[493]&m[494])|(m[474]&~m[491]&~m[492]&m[493]&m[494])|(~m[474]&m[491]&~m[492]&m[493]&m[494])|(m[474]&m[491]&~m[492]&m[493]&m[494])|(~m[474]&~m[491]&m[492]&m[493]&m[494])|(m[474]&~m[491]&m[492]&m[493]&m[494])|(m[474]&m[491]&m[492]&m[493]&m[494]));
    m[495] = (((m[493]&~m[496]&~m[497]&~m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&m[498]&~m[499])|(m[493]&m[496]&~m[497]&m[498]&~m[499])|(m[493]&~m[496]&m[497]&m[498]&~m[499])|(~m[493]&m[496]&~m[497]&~m[498]&m[499])|(~m[493]&~m[496]&m[497]&~m[498]&m[499])|(m[493]&m[496]&m[497]&~m[498]&m[499])|(~m[493]&m[496]&m[497]&m[498]&m[499]))&UnbiasedRNG[66])|((m[493]&~m[496]&~m[497]&m[498]&~m[499])|(~m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&~m[497]&~m[498]&m[499])|(m[493]&m[496]&~m[497]&~m[498]&m[499])|(m[493]&~m[496]&m[497]&~m[498]&m[499])|(~m[493]&~m[496]&~m[497]&m[498]&m[499])|(m[493]&~m[496]&~m[497]&m[498]&m[499])|(~m[493]&m[496]&~m[497]&m[498]&m[499])|(m[493]&m[496]&~m[497]&m[498]&m[499])|(~m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&~m[496]&m[497]&m[498]&m[499])|(m[493]&m[496]&m[497]&m[498]&m[499]));
    m[500] = (((m[498]&~m[501]&~m[502]&~m[503]&~m[504])|(~m[498]&~m[501]&~m[502]&m[503]&~m[504])|(m[498]&m[501]&~m[502]&m[503]&~m[504])|(m[498]&~m[501]&m[502]&m[503]&~m[504])|(~m[498]&m[501]&~m[502]&~m[503]&m[504])|(~m[498]&~m[501]&m[502]&~m[503]&m[504])|(m[498]&m[501]&m[502]&~m[503]&m[504])|(~m[498]&m[501]&m[502]&m[503]&m[504]))&UnbiasedRNG[67])|((m[498]&~m[501]&~m[502]&m[503]&~m[504])|(~m[498]&~m[501]&~m[502]&~m[503]&m[504])|(m[498]&~m[501]&~m[502]&~m[503]&m[504])|(m[498]&m[501]&~m[502]&~m[503]&m[504])|(m[498]&~m[501]&m[502]&~m[503]&m[504])|(~m[498]&~m[501]&~m[502]&m[503]&m[504])|(m[498]&~m[501]&~m[502]&m[503]&m[504])|(~m[498]&m[501]&~m[502]&m[503]&m[504])|(m[498]&m[501]&~m[502]&m[503]&m[504])|(~m[498]&~m[501]&m[502]&m[503]&m[504])|(m[498]&~m[501]&m[502]&m[503]&m[504])|(m[498]&m[501]&m[502]&m[503]&m[504]));
    m[505] = (((m[494]&~m[506]&~m[507]&~m[508]&~m[509])|(~m[494]&~m[506]&~m[507]&m[508]&~m[509])|(m[494]&m[506]&~m[507]&m[508]&~m[509])|(m[494]&~m[506]&m[507]&m[508]&~m[509])|(~m[494]&m[506]&~m[507]&~m[508]&m[509])|(~m[494]&~m[506]&m[507]&~m[508]&m[509])|(m[494]&m[506]&m[507]&~m[508]&m[509])|(~m[494]&m[506]&m[507]&m[508]&m[509]))&UnbiasedRNG[68])|((m[494]&~m[506]&~m[507]&m[508]&~m[509])|(~m[494]&~m[506]&~m[507]&~m[508]&m[509])|(m[494]&~m[506]&~m[507]&~m[508]&m[509])|(m[494]&m[506]&~m[507]&~m[508]&m[509])|(m[494]&~m[506]&m[507]&~m[508]&m[509])|(~m[494]&~m[506]&~m[507]&m[508]&m[509])|(m[494]&~m[506]&~m[507]&m[508]&m[509])|(~m[494]&m[506]&~m[507]&m[508]&m[509])|(m[494]&m[506]&~m[507]&m[508]&m[509])|(~m[494]&~m[506]&m[507]&m[508]&m[509])|(m[494]&~m[506]&m[507]&m[508]&m[509])|(m[494]&m[506]&m[507]&m[508]&m[509]));
    m[510] = (((m[508]&~m[511]&~m[512]&~m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&m[513]&~m[514])|(m[508]&m[511]&~m[512]&m[513]&~m[514])|(m[508]&~m[511]&m[512]&m[513]&~m[514])|(~m[508]&m[511]&~m[512]&~m[513]&m[514])|(~m[508]&~m[511]&m[512]&~m[513]&m[514])|(m[508]&m[511]&m[512]&~m[513]&m[514])|(~m[508]&m[511]&m[512]&m[513]&m[514]))&UnbiasedRNG[69])|((m[508]&~m[511]&~m[512]&m[513]&~m[514])|(~m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&~m[512]&~m[513]&m[514])|(m[508]&m[511]&~m[512]&~m[513]&m[514])|(m[508]&~m[511]&m[512]&~m[513]&m[514])|(~m[508]&~m[511]&~m[512]&m[513]&m[514])|(m[508]&~m[511]&~m[512]&m[513]&m[514])|(~m[508]&m[511]&~m[512]&m[513]&m[514])|(m[508]&m[511]&~m[512]&m[513]&m[514])|(~m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&~m[511]&m[512]&m[513]&m[514])|(m[508]&m[511]&m[512]&m[513]&m[514]));
    m[515] = (((m[509]&~m[516]&~m[517]&~m[518]&~m[519])|(~m[509]&~m[516]&~m[517]&m[518]&~m[519])|(m[509]&m[516]&~m[517]&m[518]&~m[519])|(m[509]&~m[516]&m[517]&m[518]&~m[519])|(~m[509]&m[516]&~m[517]&~m[518]&m[519])|(~m[509]&~m[516]&m[517]&~m[518]&m[519])|(m[509]&m[516]&m[517]&~m[518]&m[519])|(~m[509]&m[516]&m[517]&m[518]&m[519]))&UnbiasedRNG[70])|((m[509]&~m[516]&~m[517]&m[518]&~m[519])|(~m[509]&~m[516]&~m[517]&~m[518]&m[519])|(m[509]&~m[516]&~m[517]&~m[518]&m[519])|(m[509]&m[516]&~m[517]&~m[518]&m[519])|(m[509]&~m[516]&m[517]&~m[518]&m[519])|(~m[509]&~m[516]&~m[517]&m[518]&m[519])|(m[509]&~m[516]&~m[517]&m[518]&m[519])|(~m[509]&m[516]&~m[517]&m[518]&m[519])|(m[509]&m[516]&~m[517]&m[518]&m[519])|(~m[509]&~m[516]&m[517]&m[518]&m[519])|(m[509]&~m[516]&m[517]&m[518]&m[519])|(m[509]&m[516]&m[517]&m[518]&m[519]));
end

always @(posedge color1_clk) begin
    m[16] = (((m[0]&m[48]&~m[49]&~m[50]&~m[51])|(m[0]&~m[48]&m[49]&~m[50]&~m[51])|(~m[0]&m[48]&m[49]&~m[50]&~m[51])|(m[0]&~m[48]&~m[49]&m[50]&~m[51])|(~m[0]&m[48]&~m[49]&m[50]&~m[51])|(~m[0]&~m[48]&m[49]&m[50]&~m[51])|(m[0]&~m[48]&~m[49]&~m[50]&m[51])|(~m[0]&m[48]&~m[49]&~m[50]&m[51])|(~m[0]&~m[48]&m[49]&~m[50]&m[51])|(~m[0]&~m[48]&~m[49]&m[50]&m[51]))&BiasedRNG[64])|(((m[0]&m[48]&m[49]&~m[50]&~m[51])|(m[0]&m[48]&~m[49]&m[50]&~m[51])|(m[0]&~m[48]&m[49]&m[50]&~m[51])|(~m[0]&m[48]&m[49]&m[50]&~m[51])|(m[0]&m[48]&~m[49]&~m[50]&m[51])|(m[0]&~m[48]&m[49]&~m[50]&m[51])|(~m[0]&m[48]&m[49]&~m[50]&m[51])|(m[0]&~m[48]&~m[49]&m[50]&m[51])|(~m[0]&m[48]&~m[49]&m[50]&m[51])|(~m[0]&~m[48]&m[49]&m[50]&m[51]))&~BiasedRNG[64])|((m[0]&m[48]&m[49]&m[50]&~m[51])|(m[0]&m[48]&m[49]&~m[50]&m[51])|(m[0]&m[48]&~m[49]&m[50]&m[51])|(m[0]&~m[48]&m[49]&m[50]&m[51])|(~m[0]&m[48]&m[49]&m[50]&m[51])|(m[0]&m[48]&m[49]&m[50]&m[51]));
    m[17] = (((m[0]&m[52]&~m[53]&~m[54]&~m[55])|(m[0]&~m[52]&m[53]&~m[54]&~m[55])|(~m[0]&m[52]&m[53]&~m[54]&~m[55])|(m[0]&~m[52]&~m[53]&m[54]&~m[55])|(~m[0]&m[52]&~m[53]&m[54]&~m[55])|(~m[0]&~m[52]&m[53]&m[54]&~m[55])|(m[0]&~m[52]&~m[53]&~m[54]&m[55])|(~m[0]&m[52]&~m[53]&~m[54]&m[55])|(~m[0]&~m[52]&m[53]&~m[54]&m[55])|(~m[0]&~m[52]&~m[53]&m[54]&m[55]))&BiasedRNG[65])|(((m[0]&m[52]&m[53]&~m[54]&~m[55])|(m[0]&m[52]&~m[53]&m[54]&~m[55])|(m[0]&~m[52]&m[53]&m[54]&~m[55])|(~m[0]&m[52]&m[53]&m[54]&~m[55])|(m[0]&m[52]&~m[53]&~m[54]&m[55])|(m[0]&~m[52]&m[53]&~m[54]&m[55])|(~m[0]&m[52]&m[53]&~m[54]&m[55])|(m[0]&~m[52]&~m[53]&m[54]&m[55])|(~m[0]&m[52]&~m[53]&m[54]&m[55])|(~m[0]&~m[52]&m[53]&m[54]&m[55]))&~BiasedRNG[65])|((m[0]&m[52]&m[53]&m[54]&~m[55])|(m[0]&m[52]&m[53]&~m[54]&m[55])|(m[0]&m[52]&~m[53]&m[54]&m[55])|(m[0]&~m[52]&m[53]&m[54]&m[55])|(~m[0]&m[52]&m[53]&m[54]&m[55])|(m[0]&m[52]&m[53]&m[54]&m[55]));
    m[18] = (((m[1]&m[56]&~m[57]&~m[58]&~m[59])|(m[1]&~m[56]&m[57]&~m[58]&~m[59])|(~m[1]&m[56]&m[57]&~m[58]&~m[59])|(m[1]&~m[56]&~m[57]&m[58]&~m[59])|(~m[1]&m[56]&~m[57]&m[58]&~m[59])|(~m[1]&~m[56]&m[57]&m[58]&~m[59])|(m[1]&~m[56]&~m[57]&~m[58]&m[59])|(~m[1]&m[56]&~m[57]&~m[58]&m[59])|(~m[1]&~m[56]&m[57]&~m[58]&m[59])|(~m[1]&~m[56]&~m[57]&m[58]&m[59]))&BiasedRNG[66])|(((m[1]&m[56]&m[57]&~m[58]&~m[59])|(m[1]&m[56]&~m[57]&m[58]&~m[59])|(m[1]&~m[56]&m[57]&m[58]&~m[59])|(~m[1]&m[56]&m[57]&m[58]&~m[59])|(m[1]&m[56]&~m[57]&~m[58]&m[59])|(m[1]&~m[56]&m[57]&~m[58]&m[59])|(~m[1]&m[56]&m[57]&~m[58]&m[59])|(m[1]&~m[56]&~m[57]&m[58]&m[59])|(~m[1]&m[56]&~m[57]&m[58]&m[59])|(~m[1]&~m[56]&m[57]&m[58]&m[59]))&~BiasedRNG[66])|((m[1]&m[56]&m[57]&m[58]&~m[59])|(m[1]&m[56]&m[57]&~m[58]&m[59])|(m[1]&m[56]&~m[57]&m[58]&m[59])|(m[1]&~m[56]&m[57]&m[58]&m[59])|(~m[1]&m[56]&m[57]&m[58]&m[59])|(m[1]&m[56]&m[57]&m[58]&m[59]));
    m[19] = (((m[1]&m[60]&~m[61]&~m[62]&~m[63])|(m[1]&~m[60]&m[61]&~m[62]&~m[63])|(~m[1]&m[60]&m[61]&~m[62]&~m[63])|(m[1]&~m[60]&~m[61]&m[62]&~m[63])|(~m[1]&m[60]&~m[61]&m[62]&~m[63])|(~m[1]&~m[60]&m[61]&m[62]&~m[63])|(m[1]&~m[60]&~m[61]&~m[62]&m[63])|(~m[1]&m[60]&~m[61]&~m[62]&m[63])|(~m[1]&~m[60]&m[61]&~m[62]&m[63])|(~m[1]&~m[60]&~m[61]&m[62]&m[63]))&BiasedRNG[67])|(((m[1]&m[60]&m[61]&~m[62]&~m[63])|(m[1]&m[60]&~m[61]&m[62]&~m[63])|(m[1]&~m[60]&m[61]&m[62]&~m[63])|(~m[1]&m[60]&m[61]&m[62]&~m[63])|(m[1]&m[60]&~m[61]&~m[62]&m[63])|(m[1]&~m[60]&m[61]&~m[62]&m[63])|(~m[1]&m[60]&m[61]&~m[62]&m[63])|(m[1]&~m[60]&~m[61]&m[62]&m[63])|(~m[1]&m[60]&~m[61]&m[62]&m[63])|(~m[1]&~m[60]&m[61]&m[62]&m[63]))&~BiasedRNG[67])|((m[1]&m[60]&m[61]&m[62]&~m[63])|(m[1]&m[60]&m[61]&~m[62]&m[63])|(m[1]&m[60]&~m[61]&m[62]&m[63])|(m[1]&~m[60]&m[61]&m[62]&m[63])|(~m[1]&m[60]&m[61]&m[62]&m[63])|(m[1]&m[60]&m[61]&m[62]&m[63]));
    m[20] = (((m[2]&m[64]&~m[65]&~m[66]&~m[67])|(m[2]&~m[64]&m[65]&~m[66]&~m[67])|(~m[2]&m[64]&m[65]&~m[66]&~m[67])|(m[2]&~m[64]&~m[65]&m[66]&~m[67])|(~m[2]&m[64]&~m[65]&m[66]&~m[67])|(~m[2]&~m[64]&m[65]&m[66]&~m[67])|(m[2]&~m[64]&~m[65]&~m[66]&m[67])|(~m[2]&m[64]&~m[65]&~m[66]&m[67])|(~m[2]&~m[64]&m[65]&~m[66]&m[67])|(~m[2]&~m[64]&~m[65]&m[66]&m[67]))&BiasedRNG[68])|(((m[2]&m[64]&m[65]&~m[66]&~m[67])|(m[2]&m[64]&~m[65]&m[66]&~m[67])|(m[2]&~m[64]&m[65]&m[66]&~m[67])|(~m[2]&m[64]&m[65]&m[66]&~m[67])|(m[2]&m[64]&~m[65]&~m[66]&m[67])|(m[2]&~m[64]&m[65]&~m[66]&m[67])|(~m[2]&m[64]&m[65]&~m[66]&m[67])|(m[2]&~m[64]&~m[65]&m[66]&m[67])|(~m[2]&m[64]&~m[65]&m[66]&m[67])|(~m[2]&~m[64]&m[65]&m[66]&m[67]))&~BiasedRNG[68])|((m[2]&m[64]&m[65]&m[66]&~m[67])|(m[2]&m[64]&m[65]&~m[66]&m[67])|(m[2]&m[64]&~m[65]&m[66]&m[67])|(m[2]&~m[64]&m[65]&m[66]&m[67])|(~m[2]&m[64]&m[65]&m[66]&m[67])|(m[2]&m[64]&m[65]&m[66]&m[67]));
    m[21] = (((m[2]&m[68]&~m[69]&~m[70]&~m[71])|(m[2]&~m[68]&m[69]&~m[70]&~m[71])|(~m[2]&m[68]&m[69]&~m[70]&~m[71])|(m[2]&~m[68]&~m[69]&m[70]&~m[71])|(~m[2]&m[68]&~m[69]&m[70]&~m[71])|(~m[2]&~m[68]&m[69]&m[70]&~m[71])|(m[2]&~m[68]&~m[69]&~m[70]&m[71])|(~m[2]&m[68]&~m[69]&~m[70]&m[71])|(~m[2]&~m[68]&m[69]&~m[70]&m[71])|(~m[2]&~m[68]&~m[69]&m[70]&m[71]))&BiasedRNG[69])|(((m[2]&m[68]&m[69]&~m[70]&~m[71])|(m[2]&m[68]&~m[69]&m[70]&~m[71])|(m[2]&~m[68]&m[69]&m[70]&~m[71])|(~m[2]&m[68]&m[69]&m[70]&~m[71])|(m[2]&m[68]&~m[69]&~m[70]&m[71])|(m[2]&~m[68]&m[69]&~m[70]&m[71])|(~m[2]&m[68]&m[69]&~m[70]&m[71])|(m[2]&~m[68]&~m[69]&m[70]&m[71])|(~m[2]&m[68]&~m[69]&m[70]&m[71])|(~m[2]&~m[68]&m[69]&m[70]&m[71]))&~BiasedRNG[69])|((m[2]&m[68]&m[69]&m[70]&~m[71])|(m[2]&m[68]&m[69]&~m[70]&m[71])|(m[2]&m[68]&~m[69]&m[70]&m[71])|(m[2]&~m[68]&m[69]&m[70]&m[71])|(~m[2]&m[68]&m[69]&m[70]&m[71])|(m[2]&m[68]&m[69]&m[70]&m[71]));
    m[22] = (((m[3]&m[72]&~m[73]&~m[74]&~m[75])|(m[3]&~m[72]&m[73]&~m[74]&~m[75])|(~m[3]&m[72]&m[73]&~m[74]&~m[75])|(m[3]&~m[72]&~m[73]&m[74]&~m[75])|(~m[3]&m[72]&~m[73]&m[74]&~m[75])|(~m[3]&~m[72]&m[73]&m[74]&~m[75])|(m[3]&~m[72]&~m[73]&~m[74]&m[75])|(~m[3]&m[72]&~m[73]&~m[74]&m[75])|(~m[3]&~m[72]&m[73]&~m[74]&m[75])|(~m[3]&~m[72]&~m[73]&m[74]&m[75]))&BiasedRNG[70])|(((m[3]&m[72]&m[73]&~m[74]&~m[75])|(m[3]&m[72]&~m[73]&m[74]&~m[75])|(m[3]&~m[72]&m[73]&m[74]&~m[75])|(~m[3]&m[72]&m[73]&m[74]&~m[75])|(m[3]&m[72]&~m[73]&~m[74]&m[75])|(m[3]&~m[72]&m[73]&~m[74]&m[75])|(~m[3]&m[72]&m[73]&~m[74]&m[75])|(m[3]&~m[72]&~m[73]&m[74]&m[75])|(~m[3]&m[72]&~m[73]&m[74]&m[75])|(~m[3]&~m[72]&m[73]&m[74]&m[75]))&~BiasedRNG[70])|((m[3]&m[72]&m[73]&m[74]&~m[75])|(m[3]&m[72]&m[73]&~m[74]&m[75])|(m[3]&m[72]&~m[73]&m[74]&m[75])|(m[3]&~m[72]&m[73]&m[74]&m[75])|(~m[3]&m[72]&m[73]&m[74]&m[75])|(m[3]&m[72]&m[73]&m[74]&m[75]));
    m[23] = (((m[3]&m[76]&~m[77]&~m[78]&~m[79])|(m[3]&~m[76]&m[77]&~m[78]&~m[79])|(~m[3]&m[76]&m[77]&~m[78]&~m[79])|(m[3]&~m[76]&~m[77]&m[78]&~m[79])|(~m[3]&m[76]&~m[77]&m[78]&~m[79])|(~m[3]&~m[76]&m[77]&m[78]&~m[79])|(m[3]&~m[76]&~m[77]&~m[78]&m[79])|(~m[3]&m[76]&~m[77]&~m[78]&m[79])|(~m[3]&~m[76]&m[77]&~m[78]&m[79])|(~m[3]&~m[76]&~m[77]&m[78]&m[79]))&BiasedRNG[71])|(((m[3]&m[76]&m[77]&~m[78]&~m[79])|(m[3]&m[76]&~m[77]&m[78]&~m[79])|(m[3]&~m[76]&m[77]&m[78]&~m[79])|(~m[3]&m[76]&m[77]&m[78]&~m[79])|(m[3]&m[76]&~m[77]&~m[78]&m[79])|(m[3]&~m[76]&m[77]&~m[78]&m[79])|(~m[3]&m[76]&m[77]&~m[78]&m[79])|(m[3]&~m[76]&~m[77]&m[78]&m[79])|(~m[3]&m[76]&~m[77]&m[78]&m[79])|(~m[3]&~m[76]&m[77]&m[78]&m[79]))&~BiasedRNG[71])|((m[3]&m[76]&m[77]&m[78]&~m[79])|(m[3]&m[76]&m[77]&~m[78]&m[79])|(m[3]&m[76]&~m[77]&m[78]&m[79])|(m[3]&~m[76]&m[77]&m[78]&m[79])|(~m[3]&m[76]&m[77]&m[78]&m[79])|(m[3]&m[76]&m[77]&m[78]&m[79]));
    m[24] = (((m[4]&m[80]&~m[81]&~m[82]&~m[83])|(m[4]&~m[80]&m[81]&~m[82]&~m[83])|(~m[4]&m[80]&m[81]&~m[82]&~m[83])|(m[4]&~m[80]&~m[81]&m[82]&~m[83])|(~m[4]&m[80]&~m[81]&m[82]&~m[83])|(~m[4]&~m[80]&m[81]&m[82]&~m[83])|(m[4]&~m[80]&~m[81]&~m[82]&m[83])|(~m[4]&m[80]&~m[81]&~m[82]&m[83])|(~m[4]&~m[80]&m[81]&~m[82]&m[83])|(~m[4]&~m[80]&~m[81]&m[82]&m[83]))&BiasedRNG[72])|(((m[4]&m[80]&m[81]&~m[82]&~m[83])|(m[4]&m[80]&~m[81]&m[82]&~m[83])|(m[4]&~m[80]&m[81]&m[82]&~m[83])|(~m[4]&m[80]&m[81]&m[82]&~m[83])|(m[4]&m[80]&~m[81]&~m[82]&m[83])|(m[4]&~m[80]&m[81]&~m[82]&m[83])|(~m[4]&m[80]&m[81]&~m[82]&m[83])|(m[4]&~m[80]&~m[81]&m[82]&m[83])|(~m[4]&m[80]&~m[81]&m[82]&m[83])|(~m[4]&~m[80]&m[81]&m[82]&m[83]))&~BiasedRNG[72])|((m[4]&m[80]&m[81]&m[82]&~m[83])|(m[4]&m[80]&m[81]&~m[82]&m[83])|(m[4]&m[80]&~m[81]&m[82]&m[83])|(m[4]&~m[80]&m[81]&m[82]&m[83])|(~m[4]&m[80]&m[81]&m[82]&m[83])|(m[4]&m[80]&m[81]&m[82]&m[83]));
    m[25] = (((m[4]&m[84]&~m[85]&~m[86]&~m[87])|(m[4]&~m[84]&m[85]&~m[86]&~m[87])|(~m[4]&m[84]&m[85]&~m[86]&~m[87])|(m[4]&~m[84]&~m[85]&m[86]&~m[87])|(~m[4]&m[84]&~m[85]&m[86]&~m[87])|(~m[4]&~m[84]&m[85]&m[86]&~m[87])|(m[4]&~m[84]&~m[85]&~m[86]&m[87])|(~m[4]&m[84]&~m[85]&~m[86]&m[87])|(~m[4]&~m[84]&m[85]&~m[86]&m[87])|(~m[4]&~m[84]&~m[85]&m[86]&m[87]))&BiasedRNG[73])|(((m[4]&m[84]&m[85]&~m[86]&~m[87])|(m[4]&m[84]&~m[85]&m[86]&~m[87])|(m[4]&~m[84]&m[85]&m[86]&~m[87])|(~m[4]&m[84]&m[85]&m[86]&~m[87])|(m[4]&m[84]&~m[85]&~m[86]&m[87])|(m[4]&~m[84]&m[85]&~m[86]&m[87])|(~m[4]&m[84]&m[85]&~m[86]&m[87])|(m[4]&~m[84]&~m[85]&m[86]&m[87])|(~m[4]&m[84]&~m[85]&m[86]&m[87])|(~m[4]&~m[84]&m[85]&m[86]&m[87]))&~BiasedRNG[73])|((m[4]&m[84]&m[85]&m[86]&~m[87])|(m[4]&m[84]&m[85]&~m[86]&m[87])|(m[4]&m[84]&~m[85]&m[86]&m[87])|(m[4]&~m[84]&m[85]&m[86]&m[87])|(~m[4]&m[84]&m[85]&m[86]&m[87])|(m[4]&m[84]&m[85]&m[86]&m[87]));
    m[26] = (((m[5]&m[88]&~m[89]&~m[90]&~m[91])|(m[5]&~m[88]&m[89]&~m[90]&~m[91])|(~m[5]&m[88]&m[89]&~m[90]&~m[91])|(m[5]&~m[88]&~m[89]&m[90]&~m[91])|(~m[5]&m[88]&~m[89]&m[90]&~m[91])|(~m[5]&~m[88]&m[89]&m[90]&~m[91])|(m[5]&~m[88]&~m[89]&~m[90]&m[91])|(~m[5]&m[88]&~m[89]&~m[90]&m[91])|(~m[5]&~m[88]&m[89]&~m[90]&m[91])|(~m[5]&~m[88]&~m[89]&m[90]&m[91]))&BiasedRNG[74])|(((m[5]&m[88]&m[89]&~m[90]&~m[91])|(m[5]&m[88]&~m[89]&m[90]&~m[91])|(m[5]&~m[88]&m[89]&m[90]&~m[91])|(~m[5]&m[88]&m[89]&m[90]&~m[91])|(m[5]&m[88]&~m[89]&~m[90]&m[91])|(m[5]&~m[88]&m[89]&~m[90]&m[91])|(~m[5]&m[88]&m[89]&~m[90]&m[91])|(m[5]&~m[88]&~m[89]&m[90]&m[91])|(~m[5]&m[88]&~m[89]&m[90]&m[91])|(~m[5]&~m[88]&m[89]&m[90]&m[91]))&~BiasedRNG[74])|((m[5]&m[88]&m[89]&m[90]&~m[91])|(m[5]&m[88]&m[89]&~m[90]&m[91])|(m[5]&m[88]&~m[89]&m[90]&m[91])|(m[5]&~m[88]&m[89]&m[90]&m[91])|(~m[5]&m[88]&m[89]&m[90]&m[91])|(m[5]&m[88]&m[89]&m[90]&m[91]));
    m[27] = (((m[5]&m[92]&~m[93]&~m[94]&~m[95])|(m[5]&~m[92]&m[93]&~m[94]&~m[95])|(~m[5]&m[92]&m[93]&~m[94]&~m[95])|(m[5]&~m[92]&~m[93]&m[94]&~m[95])|(~m[5]&m[92]&~m[93]&m[94]&~m[95])|(~m[5]&~m[92]&m[93]&m[94]&~m[95])|(m[5]&~m[92]&~m[93]&~m[94]&m[95])|(~m[5]&m[92]&~m[93]&~m[94]&m[95])|(~m[5]&~m[92]&m[93]&~m[94]&m[95])|(~m[5]&~m[92]&~m[93]&m[94]&m[95]))&BiasedRNG[75])|(((m[5]&m[92]&m[93]&~m[94]&~m[95])|(m[5]&m[92]&~m[93]&m[94]&~m[95])|(m[5]&~m[92]&m[93]&m[94]&~m[95])|(~m[5]&m[92]&m[93]&m[94]&~m[95])|(m[5]&m[92]&~m[93]&~m[94]&m[95])|(m[5]&~m[92]&m[93]&~m[94]&m[95])|(~m[5]&m[92]&m[93]&~m[94]&m[95])|(m[5]&~m[92]&~m[93]&m[94]&m[95])|(~m[5]&m[92]&~m[93]&m[94]&m[95])|(~m[5]&~m[92]&m[93]&m[94]&m[95]))&~BiasedRNG[75])|((m[5]&m[92]&m[93]&m[94]&~m[95])|(m[5]&m[92]&m[93]&~m[94]&m[95])|(m[5]&m[92]&~m[93]&m[94]&m[95])|(m[5]&~m[92]&m[93]&m[94]&m[95])|(~m[5]&m[92]&m[93]&m[94]&m[95])|(m[5]&m[92]&m[93]&m[94]&m[95]));
    m[28] = (((m[6]&m[96]&~m[97]&~m[98]&~m[99])|(m[6]&~m[96]&m[97]&~m[98]&~m[99])|(~m[6]&m[96]&m[97]&~m[98]&~m[99])|(m[6]&~m[96]&~m[97]&m[98]&~m[99])|(~m[6]&m[96]&~m[97]&m[98]&~m[99])|(~m[6]&~m[96]&m[97]&m[98]&~m[99])|(m[6]&~m[96]&~m[97]&~m[98]&m[99])|(~m[6]&m[96]&~m[97]&~m[98]&m[99])|(~m[6]&~m[96]&m[97]&~m[98]&m[99])|(~m[6]&~m[96]&~m[97]&m[98]&m[99]))&BiasedRNG[76])|(((m[6]&m[96]&m[97]&~m[98]&~m[99])|(m[6]&m[96]&~m[97]&m[98]&~m[99])|(m[6]&~m[96]&m[97]&m[98]&~m[99])|(~m[6]&m[96]&m[97]&m[98]&~m[99])|(m[6]&m[96]&~m[97]&~m[98]&m[99])|(m[6]&~m[96]&m[97]&~m[98]&m[99])|(~m[6]&m[96]&m[97]&~m[98]&m[99])|(m[6]&~m[96]&~m[97]&m[98]&m[99])|(~m[6]&m[96]&~m[97]&m[98]&m[99])|(~m[6]&~m[96]&m[97]&m[98]&m[99]))&~BiasedRNG[76])|((m[6]&m[96]&m[97]&m[98]&~m[99])|(m[6]&m[96]&m[97]&~m[98]&m[99])|(m[6]&m[96]&~m[97]&m[98]&m[99])|(m[6]&~m[96]&m[97]&m[98]&m[99])|(~m[6]&m[96]&m[97]&m[98]&m[99])|(m[6]&m[96]&m[97]&m[98]&m[99]));
    m[29] = (((m[6]&m[100]&~m[101]&~m[102]&~m[103])|(m[6]&~m[100]&m[101]&~m[102]&~m[103])|(~m[6]&m[100]&m[101]&~m[102]&~m[103])|(m[6]&~m[100]&~m[101]&m[102]&~m[103])|(~m[6]&m[100]&~m[101]&m[102]&~m[103])|(~m[6]&~m[100]&m[101]&m[102]&~m[103])|(m[6]&~m[100]&~m[101]&~m[102]&m[103])|(~m[6]&m[100]&~m[101]&~m[102]&m[103])|(~m[6]&~m[100]&m[101]&~m[102]&m[103])|(~m[6]&~m[100]&~m[101]&m[102]&m[103]))&BiasedRNG[77])|(((m[6]&m[100]&m[101]&~m[102]&~m[103])|(m[6]&m[100]&~m[101]&m[102]&~m[103])|(m[6]&~m[100]&m[101]&m[102]&~m[103])|(~m[6]&m[100]&m[101]&m[102]&~m[103])|(m[6]&m[100]&~m[101]&~m[102]&m[103])|(m[6]&~m[100]&m[101]&~m[102]&m[103])|(~m[6]&m[100]&m[101]&~m[102]&m[103])|(m[6]&~m[100]&~m[101]&m[102]&m[103])|(~m[6]&m[100]&~m[101]&m[102]&m[103])|(~m[6]&~m[100]&m[101]&m[102]&m[103]))&~BiasedRNG[77])|((m[6]&m[100]&m[101]&m[102]&~m[103])|(m[6]&m[100]&m[101]&~m[102]&m[103])|(m[6]&m[100]&~m[101]&m[102]&m[103])|(m[6]&~m[100]&m[101]&m[102]&m[103])|(~m[6]&m[100]&m[101]&m[102]&m[103])|(m[6]&m[100]&m[101]&m[102]&m[103]));
    m[30] = (((m[7]&m[104]&~m[105]&~m[106]&~m[107])|(m[7]&~m[104]&m[105]&~m[106]&~m[107])|(~m[7]&m[104]&m[105]&~m[106]&~m[107])|(m[7]&~m[104]&~m[105]&m[106]&~m[107])|(~m[7]&m[104]&~m[105]&m[106]&~m[107])|(~m[7]&~m[104]&m[105]&m[106]&~m[107])|(m[7]&~m[104]&~m[105]&~m[106]&m[107])|(~m[7]&m[104]&~m[105]&~m[106]&m[107])|(~m[7]&~m[104]&m[105]&~m[106]&m[107])|(~m[7]&~m[104]&~m[105]&m[106]&m[107]))&BiasedRNG[78])|(((m[7]&m[104]&m[105]&~m[106]&~m[107])|(m[7]&m[104]&~m[105]&m[106]&~m[107])|(m[7]&~m[104]&m[105]&m[106]&~m[107])|(~m[7]&m[104]&m[105]&m[106]&~m[107])|(m[7]&m[104]&~m[105]&~m[106]&m[107])|(m[7]&~m[104]&m[105]&~m[106]&m[107])|(~m[7]&m[104]&m[105]&~m[106]&m[107])|(m[7]&~m[104]&~m[105]&m[106]&m[107])|(~m[7]&m[104]&~m[105]&m[106]&m[107])|(~m[7]&~m[104]&m[105]&m[106]&m[107]))&~BiasedRNG[78])|((m[7]&m[104]&m[105]&m[106]&~m[107])|(m[7]&m[104]&m[105]&~m[106]&m[107])|(m[7]&m[104]&~m[105]&m[106]&m[107])|(m[7]&~m[104]&m[105]&m[106]&m[107])|(~m[7]&m[104]&m[105]&m[106]&m[107])|(m[7]&m[104]&m[105]&m[106]&m[107]));
    m[31] = (((m[7]&m[108]&~m[109]&~m[110]&~m[111])|(m[7]&~m[108]&m[109]&~m[110]&~m[111])|(~m[7]&m[108]&m[109]&~m[110]&~m[111])|(m[7]&~m[108]&~m[109]&m[110]&~m[111])|(~m[7]&m[108]&~m[109]&m[110]&~m[111])|(~m[7]&~m[108]&m[109]&m[110]&~m[111])|(m[7]&~m[108]&~m[109]&~m[110]&m[111])|(~m[7]&m[108]&~m[109]&~m[110]&m[111])|(~m[7]&~m[108]&m[109]&~m[110]&m[111])|(~m[7]&~m[108]&~m[109]&m[110]&m[111]))&BiasedRNG[79])|(((m[7]&m[108]&m[109]&~m[110]&~m[111])|(m[7]&m[108]&~m[109]&m[110]&~m[111])|(m[7]&~m[108]&m[109]&m[110]&~m[111])|(~m[7]&m[108]&m[109]&m[110]&~m[111])|(m[7]&m[108]&~m[109]&~m[110]&m[111])|(m[7]&~m[108]&m[109]&~m[110]&m[111])|(~m[7]&m[108]&m[109]&~m[110]&m[111])|(m[7]&~m[108]&~m[109]&m[110]&m[111])|(~m[7]&m[108]&~m[109]&m[110]&m[111])|(~m[7]&~m[108]&m[109]&m[110]&m[111]))&~BiasedRNG[79])|((m[7]&m[108]&m[109]&m[110]&~m[111])|(m[7]&m[108]&m[109]&~m[110]&m[111])|(m[7]&m[108]&~m[109]&m[110]&m[111])|(m[7]&~m[108]&m[109]&m[110]&m[111])|(~m[7]&m[108]&m[109]&m[110]&m[111])|(m[7]&m[108]&m[109]&m[110]&m[111]));
    m[32] = (((m[8]&m[112]&~m[113]&~m[114]&~m[115])|(m[8]&~m[112]&m[113]&~m[114]&~m[115])|(~m[8]&m[112]&m[113]&~m[114]&~m[115])|(m[8]&~m[112]&~m[113]&m[114]&~m[115])|(~m[8]&m[112]&~m[113]&m[114]&~m[115])|(~m[8]&~m[112]&m[113]&m[114]&~m[115])|(m[8]&~m[112]&~m[113]&~m[114]&m[115])|(~m[8]&m[112]&~m[113]&~m[114]&m[115])|(~m[8]&~m[112]&m[113]&~m[114]&m[115])|(~m[8]&~m[112]&~m[113]&m[114]&m[115]))&BiasedRNG[80])|(((m[8]&m[112]&m[113]&~m[114]&~m[115])|(m[8]&m[112]&~m[113]&m[114]&~m[115])|(m[8]&~m[112]&m[113]&m[114]&~m[115])|(~m[8]&m[112]&m[113]&m[114]&~m[115])|(m[8]&m[112]&~m[113]&~m[114]&m[115])|(m[8]&~m[112]&m[113]&~m[114]&m[115])|(~m[8]&m[112]&m[113]&~m[114]&m[115])|(m[8]&~m[112]&~m[113]&m[114]&m[115])|(~m[8]&m[112]&~m[113]&m[114]&m[115])|(~m[8]&~m[112]&m[113]&m[114]&m[115]))&~BiasedRNG[80])|((m[8]&m[112]&m[113]&m[114]&~m[115])|(m[8]&m[112]&m[113]&~m[114]&m[115])|(m[8]&m[112]&~m[113]&m[114]&m[115])|(m[8]&~m[112]&m[113]&m[114]&m[115])|(~m[8]&m[112]&m[113]&m[114]&m[115])|(m[8]&m[112]&m[113]&m[114]&m[115]));
    m[33] = (((m[8]&m[116]&~m[117]&~m[118]&~m[119])|(m[8]&~m[116]&m[117]&~m[118]&~m[119])|(~m[8]&m[116]&m[117]&~m[118]&~m[119])|(m[8]&~m[116]&~m[117]&m[118]&~m[119])|(~m[8]&m[116]&~m[117]&m[118]&~m[119])|(~m[8]&~m[116]&m[117]&m[118]&~m[119])|(m[8]&~m[116]&~m[117]&~m[118]&m[119])|(~m[8]&m[116]&~m[117]&~m[118]&m[119])|(~m[8]&~m[116]&m[117]&~m[118]&m[119])|(~m[8]&~m[116]&~m[117]&m[118]&m[119]))&BiasedRNG[81])|(((m[8]&m[116]&m[117]&~m[118]&~m[119])|(m[8]&m[116]&~m[117]&m[118]&~m[119])|(m[8]&~m[116]&m[117]&m[118]&~m[119])|(~m[8]&m[116]&m[117]&m[118]&~m[119])|(m[8]&m[116]&~m[117]&~m[118]&m[119])|(m[8]&~m[116]&m[117]&~m[118]&m[119])|(~m[8]&m[116]&m[117]&~m[118]&m[119])|(m[8]&~m[116]&~m[117]&m[118]&m[119])|(~m[8]&m[116]&~m[117]&m[118]&m[119])|(~m[8]&~m[116]&m[117]&m[118]&m[119]))&~BiasedRNG[81])|((m[8]&m[116]&m[117]&m[118]&~m[119])|(m[8]&m[116]&m[117]&~m[118]&m[119])|(m[8]&m[116]&~m[117]&m[118]&m[119])|(m[8]&~m[116]&m[117]&m[118]&m[119])|(~m[8]&m[116]&m[117]&m[118]&m[119])|(m[8]&m[116]&m[117]&m[118]&m[119]));
    m[34] = (((m[9]&m[120]&~m[121]&~m[122]&~m[123])|(m[9]&~m[120]&m[121]&~m[122]&~m[123])|(~m[9]&m[120]&m[121]&~m[122]&~m[123])|(m[9]&~m[120]&~m[121]&m[122]&~m[123])|(~m[9]&m[120]&~m[121]&m[122]&~m[123])|(~m[9]&~m[120]&m[121]&m[122]&~m[123])|(m[9]&~m[120]&~m[121]&~m[122]&m[123])|(~m[9]&m[120]&~m[121]&~m[122]&m[123])|(~m[9]&~m[120]&m[121]&~m[122]&m[123])|(~m[9]&~m[120]&~m[121]&m[122]&m[123]))&BiasedRNG[82])|(((m[9]&m[120]&m[121]&~m[122]&~m[123])|(m[9]&m[120]&~m[121]&m[122]&~m[123])|(m[9]&~m[120]&m[121]&m[122]&~m[123])|(~m[9]&m[120]&m[121]&m[122]&~m[123])|(m[9]&m[120]&~m[121]&~m[122]&m[123])|(m[9]&~m[120]&m[121]&~m[122]&m[123])|(~m[9]&m[120]&m[121]&~m[122]&m[123])|(m[9]&~m[120]&~m[121]&m[122]&m[123])|(~m[9]&m[120]&~m[121]&m[122]&m[123])|(~m[9]&~m[120]&m[121]&m[122]&m[123]))&~BiasedRNG[82])|((m[9]&m[120]&m[121]&m[122]&~m[123])|(m[9]&m[120]&m[121]&~m[122]&m[123])|(m[9]&m[120]&~m[121]&m[122]&m[123])|(m[9]&~m[120]&m[121]&m[122]&m[123])|(~m[9]&m[120]&m[121]&m[122]&m[123])|(m[9]&m[120]&m[121]&m[122]&m[123]));
    m[35] = (((m[9]&m[124]&~m[125]&~m[126]&~m[127])|(m[9]&~m[124]&m[125]&~m[126]&~m[127])|(~m[9]&m[124]&m[125]&~m[126]&~m[127])|(m[9]&~m[124]&~m[125]&m[126]&~m[127])|(~m[9]&m[124]&~m[125]&m[126]&~m[127])|(~m[9]&~m[124]&m[125]&m[126]&~m[127])|(m[9]&~m[124]&~m[125]&~m[126]&m[127])|(~m[9]&m[124]&~m[125]&~m[126]&m[127])|(~m[9]&~m[124]&m[125]&~m[126]&m[127])|(~m[9]&~m[124]&~m[125]&m[126]&m[127]))&BiasedRNG[83])|(((m[9]&m[124]&m[125]&~m[126]&~m[127])|(m[9]&m[124]&~m[125]&m[126]&~m[127])|(m[9]&~m[124]&m[125]&m[126]&~m[127])|(~m[9]&m[124]&m[125]&m[126]&~m[127])|(m[9]&m[124]&~m[125]&~m[126]&m[127])|(m[9]&~m[124]&m[125]&~m[126]&m[127])|(~m[9]&m[124]&m[125]&~m[126]&m[127])|(m[9]&~m[124]&~m[125]&m[126]&m[127])|(~m[9]&m[124]&~m[125]&m[126]&m[127])|(~m[9]&~m[124]&m[125]&m[126]&m[127]))&~BiasedRNG[83])|((m[9]&m[124]&m[125]&m[126]&~m[127])|(m[9]&m[124]&m[125]&~m[126]&m[127])|(m[9]&m[124]&~m[125]&m[126]&m[127])|(m[9]&~m[124]&m[125]&m[126]&m[127])|(~m[9]&m[124]&m[125]&m[126]&m[127])|(m[9]&m[124]&m[125]&m[126]&m[127]));
    m[36] = (((m[10]&m[128]&~m[129]&~m[130]&~m[131])|(m[10]&~m[128]&m[129]&~m[130]&~m[131])|(~m[10]&m[128]&m[129]&~m[130]&~m[131])|(m[10]&~m[128]&~m[129]&m[130]&~m[131])|(~m[10]&m[128]&~m[129]&m[130]&~m[131])|(~m[10]&~m[128]&m[129]&m[130]&~m[131])|(m[10]&~m[128]&~m[129]&~m[130]&m[131])|(~m[10]&m[128]&~m[129]&~m[130]&m[131])|(~m[10]&~m[128]&m[129]&~m[130]&m[131])|(~m[10]&~m[128]&~m[129]&m[130]&m[131]))&BiasedRNG[84])|(((m[10]&m[128]&m[129]&~m[130]&~m[131])|(m[10]&m[128]&~m[129]&m[130]&~m[131])|(m[10]&~m[128]&m[129]&m[130]&~m[131])|(~m[10]&m[128]&m[129]&m[130]&~m[131])|(m[10]&m[128]&~m[129]&~m[130]&m[131])|(m[10]&~m[128]&m[129]&~m[130]&m[131])|(~m[10]&m[128]&m[129]&~m[130]&m[131])|(m[10]&~m[128]&~m[129]&m[130]&m[131])|(~m[10]&m[128]&~m[129]&m[130]&m[131])|(~m[10]&~m[128]&m[129]&m[130]&m[131]))&~BiasedRNG[84])|((m[10]&m[128]&m[129]&m[130]&~m[131])|(m[10]&m[128]&m[129]&~m[130]&m[131])|(m[10]&m[128]&~m[129]&m[130]&m[131])|(m[10]&~m[128]&m[129]&m[130]&m[131])|(~m[10]&m[128]&m[129]&m[130]&m[131])|(m[10]&m[128]&m[129]&m[130]&m[131]));
    m[37] = (((m[10]&m[132]&~m[133]&~m[134]&~m[135])|(m[10]&~m[132]&m[133]&~m[134]&~m[135])|(~m[10]&m[132]&m[133]&~m[134]&~m[135])|(m[10]&~m[132]&~m[133]&m[134]&~m[135])|(~m[10]&m[132]&~m[133]&m[134]&~m[135])|(~m[10]&~m[132]&m[133]&m[134]&~m[135])|(m[10]&~m[132]&~m[133]&~m[134]&m[135])|(~m[10]&m[132]&~m[133]&~m[134]&m[135])|(~m[10]&~m[132]&m[133]&~m[134]&m[135])|(~m[10]&~m[132]&~m[133]&m[134]&m[135]))&BiasedRNG[85])|(((m[10]&m[132]&m[133]&~m[134]&~m[135])|(m[10]&m[132]&~m[133]&m[134]&~m[135])|(m[10]&~m[132]&m[133]&m[134]&~m[135])|(~m[10]&m[132]&m[133]&m[134]&~m[135])|(m[10]&m[132]&~m[133]&~m[134]&m[135])|(m[10]&~m[132]&m[133]&~m[134]&m[135])|(~m[10]&m[132]&m[133]&~m[134]&m[135])|(m[10]&~m[132]&~m[133]&m[134]&m[135])|(~m[10]&m[132]&~m[133]&m[134]&m[135])|(~m[10]&~m[132]&m[133]&m[134]&m[135]))&~BiasedRNG[85])|((m[10]&m[132]&m[133]&m[134]&~m[135])|(m[10]&m[132]&m[133]&~m[134]&m[135])|(m[10]&m[132]&~m[133]&m[134]&m[135])|(m[10]&~m[132]&m[133]&m[134]&m[135])|(~m[10]&m[132]&m[133]&m[134]&m[135])|(m[10]&m[132]&m[133]&m[134]&m[135]));
    m[38] = (((m[11]&m[136]&~m[137]&~m[138]&~m[139])|(m[11]&~m[136]&m[137]&~m[138]&~m[139])|(~m[11]&m[136]&m[137]&~m[138]&~m[139])|(m[11]&~m[136]&~m[137]&m[138]&~m[139])|(~m[11]&m[136]&~m[137]&m[138]&~m[139])|(~m[11]&~m[136]&m[137]&m[138]&~m[139])|(m[11]&~m[136]&~m[137]&~m[138]&m[139])|(~m[11]&m[136]&~m[137]&~m[138]&m[139])|(~m[11]&~m[136]&m[137]&~m[138]&m[139])|(~m[11]&~m[136]&~m[137]&m[138]&m[139]))&BiasedRNG[86])|(((m[11]&m[136]&m[137]&~m[138]&~m[139])|(m[11]&m[136]&~m[137]&m[138]&~m[139])|(m[11]&~m[136]&m[137]&m[138]&~m[139])|(~m[11]&m[136]&m[137]&m[138]&~m[139])|(m[11]&m[136]&~m[137]&~m[138]&m[139])|(m[11]&~m[136]&m[137]&~m[138]&m[139])|(~m[11]&m[136]&m[137]&~m[138]&m[139])|(m[11]&~m[136]&~m[137]&m[138]&m[139])|(~m[11]&m[136]&~m[137]&m[138]&m[139])|(~m[11]&~m[136]&m[137]&m[138]&m[139]))&~BiasedRNG[86])|((m[11]&m[136]&m[137]&m[138]&~m[139])|(m[11]&m[136]&m[137]&~m[138]&m[139])|(m[11]&m[136]&~m[137]&m[138]&m[139])|(m[11]&~m[136]&m[137]&m[138]&m[139])|(~m[11]&m[136]&m[137]&m[138]&m[139])|(m[11]&m[136]&m[137]&m[138]&m[139]));
    m[39] = (((m[11]&m[140]&~m[141]&~m[142]&~m[143])|(m[11]&~m[140]&m[141]&~m[142]&~m[143])|(~m[11]&m[140]&m[141]&~m[142]&~m[143])|(m[11]&~m[140]&~m[141]&m[142]&~m[143])|(~m[11]&m[140]&~m[141]&m[142]&~m[143])|(~m[11]&~m[140]&m[141]&m[142]&~m[143])|(m[11]&~m[140]&~m[141]&~m[142]&m[143])|(~m[11]&m[140]&~m[141]&~m[142]&m[143])|(~m[11]&~m[140]&m[141]&~m[142]&m[143])|(~m[11]&~m[140]&~m[141]&m[142]&m[143]))&BiasedRNG[87])|(((m[11]&m[140]&m[141]&~m[142]&~m[143])|(m[11]&m[140]&~m[141]&m[142]&~m[143])|(m[11]&~m[140]&m[141]&m[142]&~m[143])|(~m[11]&m[140]&m[141]&m[142]&~m[143])|(m[11]&m[140]&~m[141]&~m[142]&m[143])|(m[11]&~m[140]&m[141]&~m[142]&m[143])|(~m[11]&m[140]&m[141]&~m[142]&m[143])|(m[11]&~m[140]&~m[141]&m[142]&m[143])|(~m[11]&m[140]&~m[141]&m[142]&m[143])|(~m[11]&~m[140]&m[141]&m[142]&m[143]))&~BiasedRNG[87])|((m[11]&m[140]&m[141]&m[142]&~m[143])|(m[11]&m[140]&m[141]&~m[142]&m[143])|(m[11]&m[140]&~m[141]&m[142]&m[143])|(m[11]&~m[140]&m[141]&m[142]&m[143])|(~m[11]&m[140]&m[141]&m[142]&m[143])|(m[11]&m[140]&m[141]&m[142]&m[143]));
    m[40] = (((m[12]&m[144]&~m[145]&~m[146]&~m[147])|(m[12]&~m[144]&m[145]&~m[146]&~m[147])|(~m[12]&m[144]&m[145]&~m[146]&~m[147])|(m[12]&~m[144]&~m[145]&m[146]&~m[147])|(~m[12]&m[144]&~m[145]&m[146]&~m[147])|(~m[12]&~m[144]&m[145]&m[146]&~m[147])|(m[12]&~m[144]&~m[145]&~m[146]&m[147])|(~m[12]&m[144]&~m[145]&~m[146]&m[147])|(~m[12]&~m[144]&m[145]&~m[146]&m[147])|(~m[12]&~m[144]&~m[145]&m[146]&m[147]))&BiasedRNG[88])|(((m[12]&m[144]&m[145]&~m[146]&~m[147])|(m[12]&m[144]&~m[145]&m[146]&~m[147])|(m[12]&~m[144]&m[145]&m[146]&~m[147])|(~m[12]&m[144]&m[145]&m[146]&~m[147])|(m[12]&m[144]&~m[145]&~m[146]&m[147])|(m[12]&~m[144]&m[145]&~m[146]&m[147])|(~m[12]&m[144]&m[145]&~m[146]&m[147])|(m[12]&~m[144]&~m[145]&m[146]&m[147])|(~m[12]&m[144]&~m[145]&m[146]&m[147])|(~m[12]&~m[144]&m[145]&m[146]&m[147]))&~BiasedRNG[88])|((m[12]&m[144]&m[145]&m[146]&~m[147])|(m[12]&m[144]&m[145]&~m[146]&m[147])|(m[12]&m[144]&~m[145]&m[146]&m[147])|(m[12]&~m[144]&m[145]&m[146]&m[147])|(~m[12]&m[144]&m[145]&m[146]&m[147])|(m[12]&m[144]&m[145]&m[146]&m[147]));
    m[41] = (((m[12]&m[148]&~m[149]&~m[150]&~m[151])|(m[12]&~m[148]&m[149]&~m[150]&~m[151])|(~m[12]&m[148]&m[149]&~m[150]&~m[151])|(m[12]&~m[148]&~m[149]&m[150]&~m[151])|(~m[12]&m[148]&~m[149]&m[150]&~m[151])|(~m[12]&~m[148]&m[149]&m[150]&~m[151])|(m[12]&~m[148]&~m[149]&~m[150]&m[151])|(~m[12]&m[148]&~m[149]&~m[150]&m[151])|(~m[12]&~m[148]&m[149]&~m[150]&m[151])|(~m[12]&~m[148]&~m[149]&m[150]&m[151]))&BiasedRNG[89])|(((m[12]&m[148]&m[149]&~m[150]&~m[151])|(m[12]&m[148]&~m[149]&m[150]&~m[151])|(m[12]&~m[148]&m[149]&m[150]&~m[151])|(~m[12]&m[148]&m[149]&m[150]&~m[151])|(m[12]&m[148]&~m[149]&~m[150]&m[151])|(m[12]&~m[148]&m[149]&~m[150]&m[151])|(~m[12]&m[148]&m[149]&~m[150]&m[151])|(m[12]&~m[148]&~m[149]&m[150]&m[151])|(~m[12]&m[148]&~m[149]&m[150]&m[151])|(~m[12]&~m[148]&m[149]&m[150]&m[151]))&~BiasedRNG[89])|((m[12]&m[148]&m[149]&m[150]&~m[151])|(m[12]&m[148]&m[149]&~m[150]&m[151])|(m[12]&m[148]&~m[149]&m[150]&m[151])|(m[12]&~m[148]&m[149]&m[150]&m[151])|(~m[12]&m[148]&m[149]&m[150]&m[151])|(m[12]&m[148]&m[149]&m[150]&m[151]));
    m[42] = (((m[13]&m[152]&~m[153]&~m[154]&~m[155])|(m[13]&~m[152]&m[153]&~m[154]&~m[155])|(~m[13]&m[152]&m[153]&~m[154]&~m[155])|(m[13]&~m[152]&~m[153]&m[154]&~m[155])|(~m[13]&m[152]&~m[153]&m[154]&~m[155])|(~m[13]&~m[152]&m[153]&m[154]&~m[155])|(m[13]&~m[152]&~m[153]&~m[154]&m[155])|(~m[13]&m[152]&~m[153]&~m[154]&m[155])|(~m[13]&~m[152]&m[153]&~m[154]&m[155])|(~m[13]&~m[152]&~m[153]&m[154]&m[155]))&BiasedRNG[90])|(((m[13]&m[152]&m[153]&~m[154]&~m[155])|(m[13]&m[152]&~m[153]&m[154]&~m[155])|(m[13]&~m[152]&m[153]&m[154]&~m[155])|(~m[13]&m[152]&m[153]&m[154]&~m[155])|(m[13]&m[152]&~m[153]&~m[154]&m[155])|(m[13]&~m[152]&m[153]&~m[154]&m[155])|(~m[13]&m[152]&m[153]&~m[154]&m[155])|(m[13]&~m[152]&~m[153]&m[154]&m[155])|(~m[13]&m[152]&~m[153]&m[154]&m[155])|(~m[13]&~m[152]&m[153]&m[154]&m[155]))&~BiasedRNG[90])|((m[13]&m[152]&m[153]&m[154]&~m[155])|(m[13]&m[152]&m[153]&~m[154]&m[155])|(m[13]&m[152]&~m[153]&m[154]&m[155])|(m[13]&~m[152]&m[153]&m[154]&m[155])|(~m[13]&m[152]&m[153]&m[154]&m[155])|(m[13]&m[152]&m[153]&m[154]&m[155]));
    m[43] = (((m[13]&m[156]&~m[157]&~m[158]&~m[159])|(m[13]&~m[156]&m[157]&~m[158]&~m[159])|(~m[13]&m[156]&m[157]&~m[158]&~m[159])|(m[13]&~m[156]&~m[157]&m[158]&~m[159])|(~m[13]&m[156]&~m[157]&m[158]&~m[159])|(~m[13]&~m[156]&m[157]&m[158]&~m[159])|(m[13]&~m[156]&~m[157]&~m[158]&m[159])|(~m[13]&m[156]&~m[157]&~m[158]&m[159])|(~m[13]&~m[156]&m[157]&~m[158]&m[159])|(~m[13]&~m[156]&~m[157]&m[158]&m[159]))&BiasedRNG[91])|(((m[13]&m[156]&m[157]&~m[158]&~m[159])|(m[13]&m[156]&~m[157]&m[158]&~m[159])|(m[13]&~m[156]&m[157]&m[158]&~m[159])|(~m[13]&m[156]&m[157]&m[158]&~m[159])|(m[13]&m[156]&~m[157]&~m[158]&m[159])|(m[13]&~m[156]&m[157]&~m[158]&m[159])|(~m[13]&m[156]&m[157]&~m[158]&m[159])|(m[13]&~m[156]&~m[157]&m[158]&m[159])|(~m[13]&m[156]&~m[157]&m[158]&m[159])|(~m[13]&~m[156]&m[157]&m[158]&m[159]))&~BiasedRNG[91])|((m[13]&m[156]&m[157]&m[158]&~m[159])|(m[13]&m[156]&m[157]&~m[158]&m[159])|(m[13]&m[156]&~m[157]&m[158]&m[159])|(m[13]&~m[156]&m[157]&m[158]&m[159])|(~m[13]&m[156]&m[157]&m[158]&m[159])|(m[13]&m[156]&m[157]&m[158]&m[159]));
    m[44] = (((m[14]&m[160]&~m[161]&~m[162]&~m[163])|(m[14]&~m[160]&m[161]&~m[162]&~m[163])|(~m[14]&m[160]&m[161]&~m[162]&~m[163])|(m[14]&~m[160]&~m[161]&m[162]&~m[163])|(~m[14]&m[160]&~m[161]&m[162]&~m[163])|(~m[14]&~m[160]&m[161]&m[162]&~m[163])|(m[14]&~m[160]&~m[161]&~m[162]&m[163])|(~m[14]&m[160]&~m[161]&~m[162]&m[163])|(~m[14]&~m[160]&m[161]&~m[162]&m[163])|(~m[14]&~m[160]&~m[161]&m[162]&m[163]))&BiasedRNG[92])|(((m[14]&m[160]&m[161]&~m[162]&~m[163])|(m[14]&m[160]&~m[161]&m[162]&~m[163])|(m[14]&~m[160]&m[161]&m[162]&~m[163])|(~m[14]&m[160]&m[161]&m[162]&~m[163])|(m[14]&m[160]&~m[161]&~m[162]&m[163])|(m[14]&~m[160]&m[161]&~m[162]&m[163])|(~m[14]&m[160]&m[161]&~m[162]&m[163])|(m[14]&~m[160]&~m[161]&m[162]&m[163])|(~m[14]&m[160]&~m[161]&m[162]&m[163])|(~m[14]&~m[160]&m[161]&m[162]&m[163]))&~BiasedRNG[92])|((m[14]&m[160]&m[161]&m[162]&~m[163])|(m[14]&m[160]&m[161]&~m[162]&m[163])|(m[14]&m[160]&~m[161]&m[162]&m[163])|(m[14]&~m[160]&m[161]&m[162]&m[163])|(~m[14]&m[160]&m[161]&m[162]&m[163])|(m[14]&m[160]&m[161]&m[162]&m[163]));
    m[45] = (((m[14]&m[164]&~m[165]&~m[166]&~m[167])|(m[14]&~m[164]&m[165]&~m[166]&~m[167])|(~m[14]&m[164]&m[165]&~m[166]&~m[167])|(m[14]&~m[164]&~m[165]&m[166]&~m[167])|(~m[14]&m[164]&~m[165]&m[166]&~m[167])|(~m[14]&~m[164]&m[165]&m[166]&~m[167])|(m[14]&~m[164]&~m[165]&~m[166]&m[167])|(~m[14]&m[164]&~m[165]&~m[166]&m[167])|(~m[14]&~m[164]&m[165]&~m[166]&m[167])|(~m[14]&~m[164]&~m[165]&m[166]&m[167]))&BiasedRNG[93])|(((m[14]&m[164]&m[165]&~m[166]&~m[167])|(m[14]&m[164]&~m[165]&m[166]&~m[167])|(m[14]&~m[164]&m[165]&m[166]&~m[167])|(~m[14]&m[164]&m[165]&m[166]&~m[167])|(m[14]&m[164]&~m[165]&~m[166]&m[167])|(m[14]&~m[164]&m[165]&~m[166]&m[167])|(~m[14]&m[164]&m[165]&~m[166]&m[167])|(m[14]&~m[164]&~m[165]&m[166]&m[167])|(~m[14]&m[164]&~m[165]&m[166]&m[167])|(~m[14]&~m[164]&m[165]&m[166]&m[167]))&~BiasedRNG[93])|((m[14]&m[164]&m[165]&m[166]&~m[167])|(m[14]&m[164]&m[165]&~m[166]&m[167])|(m[14]&m[164]&~m[165]&m[166]&m[167])|(m[14]&~m[164]&m[165]&m[166]&m[167])|(~m[14]&m[164]&m[165]&m[166]&m[167])|(m[14]&m[164]&m[165]&m[166]&m[167]));
    m[46] = (((m[15]&m[168]&~m[169]&~m[170]&~m[171])|(m[15]&~m[168]&m[169]&~m[170]&~m[171])|(~m[15]&m[168]&m[169]&~m[170]&~m[171])|(m[15]&~m[168]&~m[169]&m[170]&~m[171])|(~m[15]&m[168]&~m[169]&m[170]&~m[171])|(~m[15]&~m[168]&m[169]&m[170]&~m[171])|(m[15]&~m[168]&~m[169]&~m[170]&m[171])|(~m[15]&m[168]&~m[169]&~m[170]&m[171])|(~m[15]&~m[168]&m[169]&~m[170]&m[171])|(~m[15]&~m[168]&~m[169]&m[170]&m[171]))&BiasedRNG[94])|(((m[15]&m[168]&m[169]&~m[170]&~m[171])|(m[15]&m[168]&~m[169]&m[170]&~m[171])|(m[15]&~m[168]&m[169]&m[170]&~m[171])|(~m[15]&m[168]&m[169]&m[170]&~m[171])|(m[15]&m[168]&~m[169]&~m[170]&m[171])|(m[15]&~m[168]&m[169]&~m[170]&m[171])|(~m[15]&m[168]&m[169]&~m[170]&m[171])|(m[15]&~m[168]&~m[169]&m[170]&m[171])|(~m[15]&m[168]&~m[169]&m[170]&m[171])|(~m[15]&~m[168]&m[169]&m[170]&m[171]))&~BiasedRNG[94])|((m[15]&m[168]&m[169]&m[170]&~m[171])|(m[15]&m[168]&m[169]&~m[170]&m[171])|(m[15]&m[168]&~m[169]&m[170]&m[171])|(m[15]&~m[168]&m[169]&m[170]&m[171])|(~m[15]&m[168]&m[169]&m[170]&m[171])|(m[15]&m[168]&m[169]&m[170]&m[171]));
    m[47] = (((m[15]&m[172]&~m[173]&~m[174]&~m[175])|(m[15]&~m[172]&m[173]&~m[174]&~m[175])|(~m[15]&m[172]&m[173]&~m[174]&~m[175])|(m[15]&~m[172]&~m[173]&m[174]&~m[175])|(~m[15]&m[172]&~m[173]&m[174]&~m[175])|(~m[15]&~m[172]&m[173]&m[174]&~m[175])|(m[15]&~m[172]&~m[173]&~m[174]&m[175])|(~m[15]&m[172]&~m[173]&~m[174]&m[175])|(~m[15]&~m[172]&m[173]&~m[174]&m[175])|(~m[15]&~m[172]&~m[173]&m[174]&m[175]))&BiasedRNG[95])|(((m[15]&m[172]&m[173]&~m[174]&~m[175])|(m[15]&m[172]&~m[173]&m[174]&~m[175])|(m[15]&~m[172]&m[173]&m[174]&~m[175])|(~m[15]&m[172]&m[173]&m[174]&~m[175])|(m[15]&m[172]&~m[173]&~m[174]&m[175])|(m[15]&~m[172]&m[173]&~m[174]&m[175])|(~m[15]&m[172]&m[173]&~m[174]&m[175])|(m[15]&~m[172]&~m[173]&m[174]&m[175])|(~m[15]&m[172]&~m[173]&m[174]&m[175])|(~m[15]&~m[172]&m[173]&m[174]&m[175]))&~BiasedRNG[95])|((m[15]&m[172]&m[173]&m[174]&~m[175])|(m[15]&m[172]&m[173]&~m[174]&m[175])|(m[15]&m[172]&~m[173]&m[174]&m[175])|(m[15]&~m[172]&m[173]&m[174]&m[175])|(~m[15]&m[172]&m[173]&m[174]&m[175])|(m[15]&m[172]&m[173]&m[174]&m[175]));
    m[177] = (((m[56]&~m[113]&m[240])|(~m[56]&m[113]&m[240]))&BiasedRNG[96])|(((m[56]&m[113]&~m[240]))&~BiasedRNG[96])|((m[56]&m[113]&m[240]));
    m[178] = (((m[64]&~m[114]&m[245])|(~m[64]&m[114]&m[245]))&BiasedRNG[97])|(((m[64]&m[114]&~m[245]))&~BiasedRNG[97])|((m[64]&m[114]&m[245]));
    m[179] = (((m[72]&~m[115]&m[255])|(~m[72]&m[115]&m[255]))&BiasedRNG[98])|(((m[72]&m[115]&~m[255]))&~BiasedRNG[98])|((m[72]&m[115]&m[255]));
    m[180] = (((m[80]&~m[116]&m[270])|(~m[80]&m[116]&m[270]))&BiasedRNG[99])|(((m[80]&m[116]&~m[270]))&~BiasedRNG[99])|((m[80]&m[116]&m[270]));
    m[181] = (((m[88]&~m[117]&m[290])|(~m[88]&m[117]&m[290]))&BiasedRNG[100])|(((m[88]&m[117]&~m[290]))&~BiasedRNG[100])|((m[88]&m[117]&m[290]));
    m[182] = (((m[96]&~m[118]&m[315])|(~m[96]&m[118]&m[315]))&BiasedRNG[101])|(((m[96]&m[118]&~m[315]))&~BiasedRNG[101])|((m[96]&m[118]&m[315]));
    m[183] = (((m[104]&~m[119]&m[345])|(~m[104]&m[119]&m[345]))&BiasedRNG[102])|(((m[104]&m[119]&~m[345]))&~BiasedRNG[102])|((m[104]&m[119]&m[345]));
    m[184] = (((m[49]&~m[120]&m[241])|(~m[49]&m[120]&m[241]))&BiasedRNG[103])|(((m[49]&m[120]&~m[241]))&~BiasedRNG[103])|((m[49]&m[120]&m[241]));
    m[185] = (((m[57]&~m[121]&m[246])|(~m[57]&m[121]&m[246]))&BiasedRNG[104])|(((m[57]&m[121]&~m[246]))&~BiasedRNG[104])|((m[57]&m[121]&m[246]));
    m[186] = (((m[65]&~m[122]&m[256])|(~m[65]&m[122]&m[256]))&BiasedRNG[105])|(((m[65]&m[122]&~m[256]))&~BiasedRNG[105])|((m[65]&m[122]&m[256]));
    m[187] = (((m[73]&~m[123]&m[271])|(~m[73]&m[123]&m[271]))&BiasedRNG[106])|(((m[73]&m[123]&~m[271]))&~BiasedRNG[106])|((m[73]&m[123]&m[271]));
    m[188] = (((m[81]&~m[124]&m[291])|(~m[81]&m[124]&m[291]))&BiasedRNG[107])|(((m[81]&m[124]&~m[291]))&~BiasedRNG[107])|((m[81]&m[124]&m[291]));
    m[189] = (((m[89]&~m[125]&m[316])|(~m[89]&m[125]&m[316]))&BiasedRNG[108])|(((m[89]&m[125]&~m[316]))&~BiasedRNG[108])|((m[89]&m[125]&m[316]));
    m[190] = (((m[97]&~m[126]&m[346])|(~m[97]&m[126]&m[346]))&BiasedRNG[109])|(((m[97]&m[126]&~m[346]))&~BiasedRNG[109])|((m[97]&m[126]&m[346]));
    m[191] = (((m[105]&~m[127]&m[381])|(~m[105]&m[127]&m[381]))&BiasedRNG[110])|(((m[105]&m[127]&~m[381]))&~BiasedRNG[110])|((m[105]&m[127]&m[381]));
    m[192] = (((m[50]&~m[128]&m[251])|(~m[50]&m[128]&m[251]))&BiasedRNG[111])|(((m[50]&m[128]&~m[251]))&~BiasedRNG[111])|((m[50]&m[128]&m[251]));
    m[193] = (((m[58]&~m[129]&m[261])|(~m[58]&m[129]&m[261]))&BiasedRNG[112])|(((m[58]&m[129]&~m[261]))&~BiasedRNG[112])|((m[58]&m[129]&m[261]));
    m[194] = (((m[66]&~m[130]&m[276])|(~m[66]&m[130]&m[276]))&BiasedRNG[113])|(((m[66]&m[130]&~m[276]))&~BiasedRNG[113])|((m[66]&m[130]&m[276]));
    m[195] = (((m[74]&~m[131]&m[296])|(~m[74]&m[131]&m[296]))&BiasedRNG[114])|(((m[74]&m[131]&~m[296]))&~BiasedRNG[114])|((m[74]&m[131]&m[296]));
    m[196] = (((m[82]&~m[132]&m[321])|(~m[82]&m[132]&m[321]))&BiasedRNG[115])|(((m[82]&m[132]&~m[321]))&~BiasedRNG[115])|((m[82]&m[132]&m[321]));
    m[197] = (((m[90]&~m[133]&m[351])|(~m[90]&m[133]&m[351]))&BiasedRNG[116])|(((m[90]&m[133]&~m[351]))&~BiasedRNG[116])|((m[90]&m[133]&m[351]));
    m[198] = (((m[98]&~m[134]&m[386])|(~m[98]&m[134]&m[386]))&BiasedRNG[117])|(((m[98]&m[134]&~m[386]))&~BiasedRNG[117])|((m[98]&m[134]&m[386]));
    m[199] = (((m[106]&~m[135]&m[416])|(~m[106]&m[135]&m[416]))&BiasedRNG[118])|(((m[106]&m[135]&~m[416]))&~BiasedRNG[118])|((m[106]&m[135]&m[416]));
    m[200] = (((m[51]&~m[136]&m[266])|(~m[51]&m[136]&m[266]))&BiasedRNG[119])|(((m[51]&m[136]&~m[266]))&~BiasedRNG[119])|((m[51]&m[136]&m[266]));
    m[201] = (((m[59]&~m[137]&m[281])|(~m[59]&m[137]&m[281]))&BiasedRNG[120])|(((m[59]&m[137]&~m[281]))&~BiasedRNG[120])|((m[59]&m[137]&m[281]));
    m[202] = (((m[67]&~m[138]&m[301])|(~m[67]&m[138]&m[301]))&BiasedRNG[121])|(((m[67]&m[138]&~m[301]))&~BiasedRNG[121])|((m[67]&m[138]&m[301]));
    m[203] = (((m[75]&~m[139]&m[326])|(~m[75]&m[139]&m[326]))&BiasedRNG[122])|(((m[75]&m[139]&~m[326]))&~BiasedRNG[122])|((m[75]&m[139]&m[326]));
    m[204] = (((m[83]&~m[140]&m[356])|(~m[83]&m[140]&m[356]))&BiasedRNG[123])|(((m[83]&m[140]&~m[356]))&~BiasedRNG[123])|((m[83]&m[140]&m[356]));
    m[205] = (((m[91]&~m[141]&m[391])|(~m[91]&m[141]&m[391]))&BiasedRNG[124])|(((m[91]&m[141]&~m[391]))&~BiasedRNG[124])|((m[91]&m[141]&m[391]));
    m[206] = (((m[99]&~m[142]&m[421])|(~m[99]&m[142]&m[421]))&BiasedRNG[125])|(((m[99]&m[142]&~m[421]))&~BiasedRNG[125])|((m[99]&m[142]&m[421]));
    m[207] = (((m[107]&~m[143]&m[446])|(~m[107]&m[143]&m[446]))&BiasedRNG[126])|(((m[107]&m[143]&~m[446]))&~BiasedRNG[126])|((m[107]&m[143]&m[446]));
    m[208] = (((m[52]&~m[144]&m[286])|(~m[52]&m[144]&m[286]))&BiasedRNG[127])|(((m[52]&m[144]&~m[286]))&~BiasedRNG[127])|((m[52]&m[144]&m[286]));
    m[209] = (((m[60]&~m[145]&m[306])|(~m[60]&m[145]&m[306]))&BiasedRNG[128])|(((m[60]&m[145]&~m[306]))&~BiasedRNG[128])|((m[60]&m[145]&m[306]));
    m[210] = (((m[68]&~m[146]&m[331])|(~m[68]&m[146]&m[331]))&BiasedRNG[129])|(((m[68]&m[146]&~m[331]))&~BiasedRNG[129])|((m[68]&m[146]&m[331]));
    m[211] = (((m[76]&~m[147]&m[361])|(~m[76]&m[147]&m[361]))&BiasedRNG[130])|(((m[76]&m[147]&~m[361]))&~BiasedRNG[130])|((m[76]&m[147]&m[361]));
    m[212] = (((m[84]&~m[148]&m[396])|(~m[84]&m[148]&m[396]))&BiasedRNG[131])|(((m[84]&m[148]&~m[396]))&~BiasedRNG[131])|((m[84]&m[148]&m[396]));
    m[213] = (((m[92]&~m[149]&m[426])|(~m[92]&m[149]&m[426]))&BiasedRNG[132])|(((m[92]&m[149]&~m[426]))&~BiasedRNG[132])|((m[92]&m[149]&m[426]));
    m[214] = (((m[100]&~m[150]&m[451])|(~m[100]&m[150]&m[451]))&BiasedRNG[133])|(((m[100]&m[150]&~m[451]))&~BiasedRNG[133])|((m[100]&m[150]&m[451]));
    m[215] = (((m[108]&~m[151]&m[471])|(~m[108]&m[151]&m[471]))&BiasedRNG[134])|(((m[108]&m[151]&~m[471]))&~BiasedRNG[134])|((m[108]&m[151]&m[471]));
    m[216] = (((m[53]&~m[152]&m[311])|(~m[53]&m[152]&m[311]))&BiasedRNG[135])|(((m[53]&m[152]&~m[311]))&~BiasedRNG[135])|((m[53]&m[152]&m[311]));
    m[217] = (((m[61]&~m[153]&m[336])|(~m[61]&m[153]&m[336]))&BiasedRNG[136])|(((m[61]&m[153]&~m[336]))&~BiasedRNG[136])|((m[61]&m[153]&m[336]));
    m[218] = (((m[69]&~m[154]&m[366])|(~m[69]&m[154]&m[366]))&BiasedRNG[137])|(((m[69]&m[154]&~m[366]))&~BiasedRNG[137])|((m[69]&m[154]&m[366]));
    m[219] = (((m[77]&~m[155]&m[401])|(~m[77]&m[155]&m[401]))&BiasedRNG[138])|(((m[77]&m[155]&~m[401]))&~BiasedRNG[138])|((m[77]&m[155]&m[401]));
    m[220] = (((m[85]&~m[156]&m[431])|(~m[85]&m[156]&m[431]))&BiasedRNG[139])|(((m[85]&m[156]&~m[431]))&~BiasedRNG[139])|((m[85]&m[156]&m[431]));
    m[221] = (((m[93]&~m[157]&m[456])|(~m[93]&m[157]&m[456]))&BiasedRNG[140])|(((m[93]&m[157]&~m[456]))&~BiasedRNG[140])|((m[93]&m[157]&m[456]));
    m[222] = (((m[101]&~m[158]&m[476])|(~m[101]&m[158]&m[476]))&BiasedRNG[141])|(((m[101]&m[158]&~m[476]))&~BiasedRNG[141])|((m[101]&m[158]&m[476]));
    m[223] = (((m[109]&~m[159]&m[491])|(~m[109]&m[159]&m[491]))&BiasedRNG[142])|(((m[109]&m[159]&~m[491]))&~BiasedRNG[142])|((m[109]&m[159]&m[491]));
    m[224] = (((m[54]&~m[160]&m[341])|(~m[54]&m[160]&m[341]))&BiasedRNG[143])|(((m[54]&m[160]&~m[341]))&~BiasedRNG[143])|((m[54]&m[160]&m[341]));
    m[225] = (((m[62]&~m[161]&m[371])|(~m[62]&m[161]&m[371]))&BiasedRNG[144])|(((m[62]&m[161]&~m[371]))&~BiasedRNG[144])|((m[62]&m[161]&m[371]));
    m[226] = (((m[70]&~m[162]&m[406])|(~m[70]&m[162]&m[406]))&BiasedRNG[145])|(((m[70]&m[162]&~m[406]))&~BiasedRNG[145])|((m[70]&m[162]&m[406]));
    m[227] = (((m[78]&~m[163]&m[436])|(~m[78]&m[163]&m[436]))&BiasedRNG[146])|(((m[78]&m[163]&~m[436]))&~BiasedRNG[146])|((m[78]&m[163]&m[436]));
    m[228] = (((m[86]&~m[164]&m[461])|(~m[86]&m[164]&m[461]))&BiasedRNG[147])|(((m[86]&m[164]&~m[461]))&~BiasedRNG[147])|((m[86]&m[164]&m[461]));
    m[229] = (((m[94]&~m[165]&m[481])|(~m[94]&m[165]&m[481]))&BiasedRNG[148])|(((m[94]&m[165]&~m[481]))&~BiasedRNG[148])|((m[94]&m[165]&m[481]));
    m[230] = (((m[102]&~m[166]&m[496])|(~m[102]&m[166]&m[496]))&BiasedRNG[149])|(((m[102]&m[166]&~m[496]))&~BiasedRNG[149])|((m[102]&m[166]&m[496]));
    m[231] = (((m[110]&~m[167]&m[506])|(~m[110]&m[167]&m[506]))&BiasedRNG[150])|(((m[110]&m[167]&~m[506]))&~BiasedRNG[150])|((m[110]&m[167]&m[506]));
    m[232] = (((m[55]&~m[168]&m[376])|(~m[55]&m[168]&m[376]))&BiasedRNG[151])|(((m[55]&m[168]&~m[376]))&~BiasedRNG[151])|((m[55]&m[168]&m[376]));
    m[233] = (((m[63]&~m[169]&m[411])|(~m[63]&m[169]&m[411]))&BiasedRNG[152])|(((m[63]&m[169]&~m[411]))&~BiasedRNG[152])|((m[63]&m[169]&m[411]));
    m[234] = (((m[71]&~m[170]&m[441])|(~m[71]&m[170]&m[441]))&BiasedRNG[153])|(((m[71]&m[170]&~m[441]))&~BiasedRNG[153])|((m[71]&m[170]&m[441]));
    m[235] = (((m[79]&~m[171]&m[466])|(~m[79]&m[171]&m[466]))&BiasedRNG[154])|(((m[79]&m[171]&~m[466]))&~BiasedRNG[154])|((m[79]&m[171]&m[466]));
    m[236] = (((m[87]&~m[172]&m[486])|(~m[87]&m[172]&m[486]))&BiasedRNG[155])|(((m[87]&m[172]&~m[486]))&~BiasedRNG[155])|((m[87]&m[172]&m[486]));
    m[237] = (((m[95]&~m[173]&m[501])|(~m[95]&m[173]&m[501]))&BiasedRNG[156])|(((m[95]&m[173]&~m[501]))&~BiasedRNG[156])|((m[95]&m[173]&m[501]));
    m[238] = (((m[103]&~m[174]&m[511])|(~m[103]&m[174]&m[511]))&BiasedRNG[157])|(((m[103]&m[174]&~m[511]))&~BiasedRNG[157])|((m[103]&m[174]&m[511]));
    m[239] = (((m[111]&~m[175]&m[516])|(~m[111]&m[175]&m[516]))&BiasedRNG[158])|(((m[111]&m[175]&~m[516]))&~BiasedRNG[158])|((m[111]&m[175]&m[516]));
    m[247] = (((m[244]&~m[245]&~m[246]&~m[248]&~m[249])|(~m[244]&~m[245]&~m[246]&m[248]&~m[249])|(m[244]&m[245]&~m[246]&m[248]&~m[249])|(m[244]&~m[245]&m[246]&m[248]&~m[249])|(~m[244]&m[245]&~m[246]&~m[248]&m[249])|(~m[244]&~m[245]&m[246]&~m[248]&m[249])|(m[244]&m[245]&m[246]&~m[248]&m[249])|(~m[244]&m[245]&m[246]&m[248]&m[249]))&UnbiasedRNG[71])|((m[244]&~m[245]&~m[246]&m[248]&~m[249])|(~m[244]&~m[245]&~m[246]&~m[248]&m[249])|(m[244]&~m[245]&~m[246]&~m[248]&m[249])|(m[244]&m[245]&~m[246]&~m[248]&m[249])|(m[244]&~m[245]&m[246]&~m[248]&m[249])|(~m[244]&~m[245]&~m[246]&m[248]&m[249])|(m[244]&~m[245]&~m[246]&m[248]&m[249])|(~m[244]&m[245]&~m[246]&m[248]&m[249])|(m[244]&m[245]&~m[246]&m[248]&m[249])|(~m[244]&~m[245]&m[246]&m[248]&m[249])|(m[244]&~m[245]&m[246]&m[248]&m[249])|(m[244]&m[245]&m[246]&m[248]&m[249]));
    m[257] = (((m[249]&~m[255]&~m[256]&~m[258]&~m[259])|(~m[249]&~m[255]&~m[256]&m[258]&~m[259])|(m[249]&m[255]&~m[256]&m[258]&~m[259])|(m[249]&~m[255]&m[256]&m[258]&~m[259])|(~m[249]&m[255]&~m[256]&~m[258]&m[259])|(~m[249]&~m[255]&m[256]&~m[258]&m[259])|(m[249]&m[255]&m[256]&~m[258]&m[259])|(~m[249]&m[255]&m[256]&m[258]&m[259]))&UnbiasedRNG[72])|((m[249]&~m[255]&~m[256]&m[258]&~m[259])|(~m[249]&~m[255]&~m[256]&~m[258]&m[259])|(m[249]&~m[255]&~m[256]&~m[258]&m[259])|(m[249]&m[255]&~m[256]&~m[258]&m[259])|(m[249]&~m[255]&m[256]&~m[258]&m[259])|(~m[249]&~m[255]&~m[256]&m[258]&m[259])|(m[249]&~m[255]&~m[256]&m[258]&m[259])|(~m[249]&m[255]&~m[256]&m[258]&m[259])|(m[249]&m[255]&~m[256]&m[258]&m[259])|(~m[249]&~m[255]&m[256]&m[258]&m[259])|(m[249]&~m[255]&m[256]&m[258]&m[259])|(m[249]&m[255]&m[256]&m[258]&m[259]));
    m[262] = (((m[254]&~m[260]&~m[261]&~m[263]&~m[264])|(~m[254]&~m[260]&~m[261]&m[263]&~m[264])|(m[254]&m[260]&~m[261]&m[263]&~m[264])|(m[254]&~m[260]&m[261]&m[263]&~m[264])|(~m[254]&m[260]&~m[261]&~m[263]&m[264])|(~m[254]&~m[260]&m[261]&~m[263]&m[264])|(m[254]&m[260]&m[261]&~m[263]&m[264])|(~m[254]&m[260]&m[261]&m[263]&m[264]))&UnbiasedRNG[73])|((m[254]&~m[260]&~m[261]&m[263]&~m[264])|(~m[254]&~m[260]&~m[261]&~m[263]&m[264])|(m[254]&~m[260]&~m[261]&~m[263]&m[264])|(m[254]&m[260]&~m[261]&~m[263]&m[264])|(m[254]&~m[260]&m[261]&~m[263]&m[264])|(~m[254]&~m[260]&~m[261]&m[263]&m[264])|(m[254]&~m[260]&~m[261]&m[263]&m[264])|(~m[254]&m[260]&~m[261]&m[263]&m[264])|(m[254]&m[260]&~m[261]&m[263]&m[264])|(~m[254]&~m[260]&m[261]&m[263]&m[264])|(m[254]&~m[260]&m[261]&m[263]&m[264])|(m[254]&m[260]&m[261]&m[263]&m[264]));
    m[272] = (((m[259]&~m[270]&~m[271]&~m[273]&~m[274])|(~m[259]&~m[270]&~m[271]&m[273]&~m[274])|(m[259]&m[270]&~m[271]&m[273]&~m[274])|(m[259]&~m[270]&m[271]&m[273]&~m[274])|(~m[259]&m[270]&~m[271]&~m[273]&m[274])|(~m[259]&~m[270]&m[271]&~m[273]&m[274])|(m[259]&m[270]&m[271]&~m[273]&m[274])|(~m[259]&m[270]&m[271]&m[273]&m[274]))&UnbiasedRNG[74])|((m[259]&~m[270]&~m[271]&m[273]&~m[274])|(~m[259]&~m[270]&~m[271]&~m[273]&m[274])|(m[259]&~m[270]&~m[271]&~m[273]&m[274])|(m[259]&m[270]&~m[271]&~m[273]&m[274])|(m[259]&~m[270]&m[271]&~m[273]&m[274])|(~m[259]&~m[270]&~m[271]&m[273]&m[274])|(m[259]&~m[270]&~m[271]&m[273]&m[274])|(~m[259]&m[270]&~m[271]&m[273]&m[274])|(m[259]&m[270]&~m[271]&m[273]&m[274])|(~m[259]&~m[270]&m[271]&m[273]&m[274])|(m[259]&~m[270]&m[271]&m[273]&m[274])|(m[259]&m[270]&m[271]&m[273]&m[274]));
    m[277] = (((m[264]&~m[275]&~m[276]&~m[278]&~m[279])|(~m[264]&~m[275]&~m[276]&m[278]&~m[279])|(m[264]&m[275]&~m[276]&m[278]&~m[279])|(m[264]&~m[275]&m[276]&m[278]&~m[279])|(~m[264]&m[275]&~m[276]&~m[278]&m[279])|(~m[264]&~m[275]&m[276]&~m[278]&m[279])|(m[264]&m[275]&m[276]&~m[278]&m[279])|(~m[264]&m[275]&m[276]&m[278]&m[279]))&UnbiasedRNG[75])|((m[264]&~m[275]&~m[276]&m[278]&~m[279])|(~m[264]&~m[275]&~m[276]&~m[278]&m[279])|(m[264]&~m[275]&~m[276]&~m[278]&m[279])|(m[264]&m[275]&~m[276]&~m[278]&m[279])|(m[264]&~m[275]&m[276]&~m[278]&m[279])|(~m[264]&~m[275]&~m[276]&m[278]&m[279])|(m[264]&~m[275]&~m[276]&m[278]&m[279])|(~m[264]&m[275]&~m[276]&m[278]&m[279])|(m[264]&m[275]&~m[276]&m[278]&m[279])|(~m[264]&~m[275]&m[276]&m[278]&m[279])|(m[264]&~m[275]&m[276]&m[278]&m[279])|(m[264]&m[275]&m[276]&m[278]&m[279]));
    m[282] = (((m[269]&~m[280]&~m[281]&~m[283]&~m[284])|(~m[269]&~m[280]&~m[281]&m[283]&~m[284])|(m[269]&m[280]&~m[281]&m[283]&~m[284])|(m[269]&~m[280]&m[281]&m[283]&~m[284])|(~m[269]&m[280]&~m[281]&~m[283]&m[284])|(~m[269]&~m[280]&m[281]&~m[283]&m[284])|(m[269]&m[280]&m[281]&~m[283]&m[284])|(~m[269]&m[280]&m[281]&m[283]&m[284]))&UnbiasedRNG[76])|((m[269]&~m[280]&~m[281]&m[283]&~m[284])|(~m[269]&~m[280]&~m[281]&~m[283]&m[284])|(m[269]&~m[280]&~m[281]&~m[283]&m[284])|(m[269]&m[280]&~m[281]&~m[283]&m[284])|(m[269]&~m[280]&m[281]&~m[283]&m[284])|(~m[269]&~m[280]&~m[281]&m[283]&m[284])|(m[269]&~m[280]&~m[281]&m[283]&m[284])|(~m[269]&m[280]&~m[281]&m[283]&m[284])|(m[269]&m[280]&~m[281]&m[283]&m[284])|(~m[269]&~m[280]&m[281]&m[283]&m[284])|(m[269]&~m[280]&m[281]&m[283]&m[284])|(m[269]&m[280]&m[281]&m[283]&m[284]));
    m[292] = (((m[274]&~m[290]&~m[291]&~m[293]&~m[294])|(~m[274]&~m[290]&~m[291]&m[293]&~m[294])|(m[274]&m[290]&~m[291]&m[293]&~m[294])|(m[274]&~m[290]&m[291]&m[293]&~m[294])|(~m[274]&m[290]&~m[291]&~m[293]&m[294])|(~m[274]&~m[290]&m[291]&~m[293]&m[294])|(m[274]&m[290]&m[291]&~m[293]&m[294])|(~m[274]&m[290]&m[291]&m[293]&m[294]))&UnbiasedRNG[77])|((m[274]&~m[290]&~m[291]&m[293]&~m[294])|(~m[274]&~m[290]&~m[291]&~m[293]&m[294])|(m[274]&~m[290]&~m[291]&~m[293]&m[294])|(m[274]&m[290]&~m[291]&~m[293]&m[294])|(m[274]&~m[290]&m[291]&~m[293]&m[294])|(~m[274]&~m[290]&~m[291]&m[293]&m[294])|(m[274]&~m[290]&~m[291]&m[293]&m[294])|(~m[274]&m[290]&~m[291]&m[293]&m[294])|(m[274]&m[290]&~m[291]&m[293]&m[294])|(~m[274]&~m[290]&m[291]&m[293]&m[294])|(m[274]&~m[290]&m[291]&m[293]&m[294])|(m[274]&m[290]&m[291]&m[293]&m[294]));
    m[297] = (((m[279]&~m[295]&~m[296]&~m[298]&~m[299])|(~m[279]&~m[295]&~m[296]&m[298]&~m[299])|(m[279]&m[295]&~m[296]&m[298]&~m[299])|(m[279]&~m[295]&m[296]&m[298]&~m[299])|(~m[279]&m[295]&~m[296]&~m[298]&m[299])|(~m[279]&~m[295]&m[296]&~m[298]&m[299])|(m[279]&m[295]&m[296]&~m[298]&m[299])|(~m[279]&m[295]&m[296]&m[298]&m[299]))&UnbiasedRNG[78])|((m[279]&~m[295]&~m[296]&m[298]&~m[299])|(~m[279]&~m[295]&~m[296]&~m[298]&m[299])|(m[279]&~m[295]&~m[296]&~m[298]&m[299])|(m[279]&m[295]&~m[296]&~m[298]&m[299])|(m[279]&~m[295]&m[296]&~m[298]&m[299])|(~m[279]&~m[295]&~m[296]&m[298]&m[299])|(m[279]&~m[295]&~m[296]&m[298]&m[299])|(~m[279]&m[295]&~m[296]&m[298]&m[299])|(m[279]&m[295]&~m[296]&m[298]&m[299])|(~m[279]&~m[295]&m[296]&m[298]&m[299])|(m[279]&~m[295]&m[296]&m[298]&m[299])|(m[279]&m[295]&m[296]&m[298]&m[299]));
    m[302] = (((m[284]&~m[300]&~m[301]&~m[303]&~m[304])|(~m[284]&~m[300]&~m[301]&m[303]&~m[304])|(m[284]&m[300]&~m[301]&m[303]&~m[304])|(m[284]&~m[300]&m[301]&m[303]&~m[304])|(~m[284]&m[300]&~m[301]&~m[303]&m[304])|(~m[284]&~m[300]&m[301]&~m[303]&m[304])|(m[284]&m[300]&m[301]&~m[303]&m[304])|(~m[284]&m[300]&m[301]&m[303]&m[304]))&UnbiasedRNG[79])|((m[284]&~m[300]&~m[301]&m[303]&~m[304])|(~m[284]&~m[300]&~m[301]&~m[303]&m[304])|(m[284]&~m[300]&~m[301]&~m[303]&m[304])|(m[284]&m[300]&~m[301]&~m[303]&m[304])|(m[284]&~m[300]&m[301]&~m[303]&m[304])|(~m[284]&~m[300]&~m[301]&m[303]&m[304])|(m[284]&~m[300]&~m[301]&m[303]&m[304])|(~m[284]&m[300]&~m[301]&m[303]&m[304])|(m[284]&m[300]&~m[301]&m[303]&m[304])|(~m[284]&~m[300]&m[301]&m[303]&m[304])|(m[284]&~m[300]&m[301]&m[303]&m[304])|(m[284]&m[300]&m[301]&m[303]&m[304]));
    m[307] = (((m[289]&~m[305]&~m[306]&~m[308]&~m[309])|(~m[289]&~m[305]&~m[306]&m[308]&~m[309])|(m[289]&m[305]&~m[306]&m[308]&~m[309])|(m[289]&~m[305]&m[306]&m[308]&~m[309])|(~m[289]&m[305]&~m[306]&~m[308]&m[309])|(~m[289]&~m[305]&m[306]&~m[308]&m[309])|(m[289]&m[305]&m[306]&~m[308]&m[309])|(~m[289]&m[305]&m[306]&m[308]&m[309]))&UnbiasedRNG[80])|((m[289]&~m[305]&~m[306]&m[308]&~m[309])|(~m[289]&~m[305]&~m[306]&~m[308]&m[309])|(m[289]&~m[305]&~m[306]&~m[308]&m[309])|(m[289]&m[305]&~m[306]&~m[308]&m[309])|(m[289]&~m[305]&m[306]&~m[308]&m[309])|(~m[289]&~m[305]&~m[306]&m[308]&m[309])|(m[289]&~m[305]&~m[306]&m[308]&m[309])|(~m[289]&m[305]&~m[306]&m[308]&m[309])|(m[289]&m[305]&~m[306]&m[308]&m[309])|(~m[289]&~m[305]&m[306]&m[308]&m[309])|(m[289]&~m[305]&m[306]&m[308]&m[309])|(m[289]&m[305]&m[306]&m[308]&m[309]));
    m[317] = (((m[294]&~m[315]&~m[316]&~m[318]&~m[319])|(~m[294]&~m[315]&~m[316]&m[318]&~m[319])|(m[294]&m[315]&~m[316]&m[318]&~m[319])|(m[294]&~m[315]&m[316]&m[318]&~m[319])|(~m[294]&m[315]&~m[316]&~m[318]&m[319])|(~m[294]&~m[315]&m[316]&~m[318]&m[319])|(m[294]&m[315]&m[316]&~m[318]&m[319])|(~m[294]&m[315]&m[316]&m[318]&m[319]))&UnbiasedRNG[81])|((m[294]&~m[315]&~m[316]&m[318]&~m[319])|(~m[294]&~m[315]&~m[316]&~m[318]&m[319])|(m[294]&~m[315]&~m[316]&~m[318]&m[319])|(m[294]&m[315]&~m[316]&~m[318]&m[319])|(m[294]&~m[315]&m[316]&~m[318]&m[319])|(~m[294]&~m[315]&~m[316]&m[318]&m[319])|(m[294]&~m[315]&~m[316]&m[318]&m[319])|(~m[294]&m[315]&~m[316]&m[318]&m[319])|(m[294]&m[315]&~m[316]&m[318]&m[319])|(~m[294]&~m[315]&m[316]&m[318]&m[319])|(m[294]&~m[315]&m[316]&m[318]&m[319])|(m[294]&m[315]&m[316]&m[318]&m[319]));
    m[322] = (((m[299]&~m[320]&~m[321]&~m[323]&~m[324])|(~m[299]&~m[320]&~m[321]&m[323]&~m[324])|(m[299]&m[320]&~m[321]&m[323]&~m[324])|(m[299]&~m[320]&m[321]&m[323]&~m[324])|(~m[299]&m[320]&~m[321]&~m[323]&m[324])|(~m[299]&~m[320]&m[321]&~m[323]&m[324])|(m[299]&m[320]&m[321]&~m[323]&m[324])|(~m[299]&m[320]&m[321]&m[323]&m[324]))&UnbiasedRNG[82])|((m[299]&~m[320]&~m[321]&m[323]&~m[324])|(~m[299]&~m[320]&~m[321]&~m[323]&m[324])|(m[299]&~m[320]&~m[321]&~m[323]&m[324])|(m[299]&m[320]&~m[321]&~m[323]&m[324])|(m[299]&~m[320]&m[321]&~m[323]&m[324])|(~m[299]&~m[320]&~m[321]&m[323]&m[324])|(m[299]&~m[320]&~m[321]&m[323]&m[324])|(~m[299]&m[320]&~m[321]&m[323]&m[324])|(m[299]&m[320]&~m[321]&m[323]&m[324])|(~m[299]&~m[320]&m[321]&m[323]&m[324])|(m[299]&~m[320]&m[321]&m[323]&m[324])|(m[299]&m[320]&m[321]&m[323]&m[324]));
    m[327] = (((m[304]&~m[325]&~m[326]&~m[328]&~m[329])|(~m[304]&~m[325]&~m[326]&m[328]&~m[329])|(m[304]&m[325]&~m[326]&m[328]&~m[329])|(m[304]&~m[325]&m[326]&m[328]&~m[329])|(~m[304]&m[325]&~m[326]&~m[328]&m[329])|(~m[304]&~m[325]&m[326]&~m[328]&m[329])|(m[304]&m[325]&m[326]&~m[328]&m[329])|(~m[304]&m[325]&m[326]&m[328]&m[329]))&UnbiasedRNG[83])|((m[304]&~m[325]&~m[326]&m[328]&~m[329])|(~m[304]&~m[325]&~m[326]&~m[328]&m[329])|(m[304]&~m[325]&~m[326]&~m[328]&m[329])|(m[304]&m[325]&~m[326]&~m[328]&m[329])|(m[304]&~m[325]&m[326]&~m[328]&m[329])|(~m[304]&~m[325]&~m[326]&m[328]&m[329])|(m[304]&~m[325]&~m[326]&m[328]&m[329])|(~m[304]&m[325]&~m[326]&m[328]&m[329])|(m[304]&m[325]&~m[326]&m[328]&m[329])|(~m[304]&~m[325]&m[326]&m[328]&m[329])|(m[304]&~m[325]&m[326]&m[328]&m[329])|(m[304]&m[325]&m[326]&m[328]&m[329]));
    m[332] = (((m[309]&~m[330]&~m[331]&~m[333]&~m[334])|(~m[309]&~m[330]&~m[331]&m[333]&~m[334])|(m[309]&m[330]&~m[331]&m[333]&~m[334])|(m[309]&~m[330]&m[331]&m[333]&~m[334])|(~m[309]&m[330]&~m[331]&~m[333]&m[334])|(~m[309]&~m[330]&m[331]&~m[333]&m[334])|(m[309]&m[330]&m[331]&~m[333]&m[334])|(~m[309]&m[330]&m[331]&m[333]&m[334]))&UnbiasedRNG[84])|((m[309]&~m[330]&~m[331]&m[333]&~m[334])|(~m[309]&~m[330]&~m[331]&~m[333]&m[334])|(m[309]&~m[330]&~m[331]&~m[333]&m[334])|(m[309]&m[330]&~m[331]&~m[333]&m[334])|(m[309]&~m[330]&m[331]&~m[333]&m[334])|(~m[309]&~m[330]&~m[331]&m[333]&m[334])|(m[309]&~m[330]&~m[331]&m[333]&m[334])|(~m[309]&m[330]&~m[331]&m[333]&m[334])|(m[309]&m[330]&~m[331]&m[333]&m[334])|(~m[309]&~m[330]&m[331]&m[333]&m[334])|(m[309]&~m[330]&m[331]&m[333]&m[334])|(m[309]&m[330]&m[331]&m[333]&m[334]));
    m[337] = (((m[314]&~m[335]&~m[336]&~m[338]&~m[339])|(~m[314]&~m[335]&~m[336]&m[338]&~m[339])|(m[314]&m[335]&~m[336]&m[338]&~m[339])|(m[314]&~m[335]&m[336]&m[338]&~m[339])|(~m[314]&m[335]&~m[336]&~m[338]&m[339])|(~m[314]&~m[335]&m[336]&~m[338]&m[339])|(m[314]&m[335]&m[336]&~m[338]&m[339])|(~m[314]&m[335]&m[336]&m[338]&m[339]))&UnbiasedRNG[85])|((m[314]&~m[335]&~m[336]&m[338]&~m[339])|(~m[314]&~m[335]&~m[336]&~m[338]&m[339])|(m[314]&~m[335]&~m[336]&~m[338]&m[339])|(m[314]&m[335]&~m[336]&~m[338]&m[339])|(m[314]&~m[335]&m[336]&~m[338]&m[339])|(~m[314]&~m[335]&~m[336]&m[338]&m[339])|(m[314]&~m[335]&~m[336]&m[338]&m[339])|(~m[314]&m[335]&~m[336]&m[338]&m[339])|(m[314]&m[335]&~m[336]&m[338]&m[339])|(~m[314]&~m[335]&m[336]&m[338]&m[339])|(m[314]&~m[335]&m[336]&m[338]&m[339])|(m[314]&m[335]&m[336]&m[338]&m[339]));
    m[347] = (((m[319]&~m[345]&~m[346]&~m[348]&~m[349])|(~m[319]&~m[345]&~m[346]&m[348]&~m[349])|(m[319]&m[345]&~m[346]&m[348]&~m[349])|(m[319]&~m[345]&m[346]&m[348]&~m[349])|(~m[319]&m[345]&~m[346]&~m[348]&m[349])|(~m[319]&~m[345]&m[346]&~m[348]&m[349])|(m[319]&m[345]&m[346]&~m[348]&m[349])|(~m[319]&m[345]&m[346]&m[348]&m[349]))&UnbiasedRNG[86])|((m[319]&~m[345]&~m[346]&m[348]&~m[349])|(~m[319]&~m[345]&~m[346]&~m[348]&m[349])|(m[319]&~m[345]&~m[346]&~m[348]&m[349])|(m[319]&m[345]&~m[346]&~m[348]&m[349])|(m[319]&~m[345]&m[346]&~m[348]&m[349])|(~m[319]&~m[345]&~m[346]&m[348]&m[349])|(m[319]&~m[345]&~m[346]&m[348]&m[349])|(~m[319]&m[345]&~m[346]&m[348]&m[349])|(m[319]&m[345]&~m[346]&m[348]&m[349])|(~m[319]&~m[345]&m[346]&m[348]&m[349])|(m[319]&~m[345]&m[346]&m[348]&m[349])|(m[319]&m[345]&m[346]&m[348]&m[349]));
    m[352] = (((m[324]&~m[350]&~m[351]&~m[353]&~m[354])|(~m[324]&~m[350]&~m[351]&m[353]&~m[354])|(m[324]&m[350]&~m[351]&m[353]&~m[354])|(m[324]&~m[350]&m[351]&m[353]&~m[354])|(~m[324]&m[350]&~m[351]&~m[353]&m[354])|(~m[324]&~m[350]&m[351]&~m[353]&m[354])|(m[324]&m[350]&m[351]&~m[353]&m[354])|(~m[324]&m[350]&m[351]&m[353]&m[354]))&UnbiasedRNG[87])|((m[324]&~m[350]&~m[351]&m[353]&~m[354])|(~m[324]&~m[350]&~m[351]&~m[353]&m[354])|(m[324]&~m[350]&~m[351]&~m[353]&m[354])|(m[324]&m[350]&~m[351]&~m[353]&m[354])|(m[324]&~m[350]&m[351]&~m[353]&m[354])|(~m[324]&~m[350]&~m[351]&m[353]&m[354])|(m[324]&~m[350]&~m[351]&m[353]&m[354])|(~m[324]&m[350]&~m[351]&m[353]&m[354])|(m[324]&m[350]&~m[351]&m[353]&m[354])|(~m[324]&~m[350]&m[351]&m[353]&m[354])|(m[324]&~m[350]&m[351]&m[353]&m[354])|(m[324]&m[350]&m[351]&m[353]&m[354]));
    m[357] = (((m[329]&~m[355]&~m[356]&~m[358]&~m[359])|(~m[329]&~m[355]&~m[356]&m[358]&~m[359])|(m[329]&m[355]&~m[356]&m[358]&~m[359])|(m[329]&~m[355]&m[356]&m[358]&~m[359])|(~m[329]&m[355]&~m[356]&~m[358]&m[359])|(~m[329]&~m[355]&m[356]&~m[358]&m[359])|(m[329]&m[355]&m[356]&~m[358]&m[359])|(~m[329]&m[355]&m[356]&m[358]&m[359]))&UnbiasedRNG[88])|((m[329]&~m[355]&~m[356]&m[358]&~m[359])|(~m[329]&~m[355]&~m[356]&~m[358]&m[359])|(m[329]&~m[355]&~m[356]&~m[358]&m[359])|(m[329]&m[355]&~m[356]&~m[358]&m[359])|(m[329]&~m[355]&m[356]&~m[358]&m[359])|(~m[329]&~m[355]&~m[356]&m[358]&m[359])|(m[329]&~m[355]&~m[356]&m[358]&m[359])|(~m[329]&m[355]&~m[356]&m[358]&m[359])|(m[329]&m[355]&~m[356]&m[358]&m[359])|(~m[329]&~m[355]&m[356]&m[358]&m[359])|(m[329]&~m[355]&m[356]&m[358]&m[359])|(m[329]&m[355]&m[356]&m[358]&m[359]));
    m[362] = (((m[334]&~m[360]&~m[361]&~m[363]&~m[364])|(~m[334]&~m[360]&~m[361]&m[363]&~m[364])|(m[334]&m[360]&~m[361]&m[363]&~m[364])|(m[334]&~m[360]&m[361]&m[363]&~m[364])|(~m[334]&m[360]&~m[361]&~m[363]&m[364])|(~m[334]&~m[360]&m[361]&~m[363]&m[364])|(m[334]&m[360]&m[361]&~m[363]&m[364])|(~m[334]&m[360]&m[361]&m[363]&m[364]))&UnbiasedRNG[89])|((m[334]&~m[360]&~m[361]&m[363]&~m[364])|(~m[334]&~m[360]&~m[361]&~m[363]&m[364])|(m[334]&~m[360]&~m[361]&~m[363]&m[364])|(m[334]&m[360]&~m[361]&~m[363]&m[364])|(m[334]&~m[360]&m[361]&~m[363]&m[364])|(~m[334]&~m[360]&~m[361]&m[363]&m[364])|(m[334]&~m[360]&~m[361]&m[363]&m[364])|(~m[334]&m[360]&~m[361]&m[363]&m[364])|(m[334]&m[360]&~m[361]&m[363]&m[364])|(~m[334]&~m[360]&m[361]&m[363]&m[364])|(m[334]&~m[360]&m[361]&m[363]&m[364])|(m[334]&m[360]&m[361]&m[363]&m[364]));
    m[367] = (((m[339]&~m[365]&~m[366]&~m[368]&~m[369])|(~m[339]&~m[365]&~m[366]&m[368]&~m[369])|(m[339]&m[365]&~m[366]&m[368]&~m[369])|(m[339]&~m[365]&m[366]&m[368]&~m[369])|(~m[339]&m[365]&~m[366]&~m[368]&m[369])|(~m[339]&~m[365]&m[366]&~m[368]&m[369])|(m[339]&m[365]&m[366]&~m[368]&m[369])|(~m[339]&m[365]&m[366]&m[368]&m[369]))&UnbiasedRNG[90])|((m[339]&~m[365]&~m[366]&m[368]&~m[369])|(~m[339]&~m[365]&~m[366]&~m[368]&m[369])|(m[339]&~m[365]&~m[366]&~m[368]&m[369])|(m[339]&m[365]&~m[366]&~m[368]&m[369])|(m[339]&~m[365]&m[366]&~m[368]&m[369])|(~m[339]&~m[365]&~m[366]&m[368]&m[369])|(m[339]&~m[365]&~m[366]&m[368]&m[369])|(~m[339]&m[365]&~m[366]&m[368]&m[369])|(m[339]&m[365]&~m[366]&m[368]&m[369])|(~m[339]&~m[365]&m[366]&m[368]&m[369])|(m[339]&~m[365]&m[366]&m[368]&m[369])|(m[339]&m[365]&m[366]&m[368]&m[369]));
    m[372] = (((m[344]&~m[370]&~m[371]&~m[373]&~m[374])|(~m[344]&~m[370]&~m[371]&m[373]&~m[374])|(m[344]&m[370]&~m[371]&m[373]&~m[374])|(m[344]&~m[370]&m[371]&m[373]&~m[374])|(~m[344]&m[370]&~m[371]&~m[373]&m[374])|(~m[344]&~m[370]&m[371]&~m[373]&m[374])|(m[344]&m[370]&m[371]&~m[373]&m[374])|(~m[344]&m[370]&m[371]&m[373]&m[374]))&UnbiasedRNG[91])|((m[344]&~m[370]&~m[371]&m[373]&~m[374])|(~m[344]&~m[370]&~m[371]&~m[373]&m[374])|(m[344]&~m[370]&~m[371]&~m[373]&m[374])|(m[344]&m[370]&~m[371]&~m[373]&m[374])|(m[344]&~m[370]&m[371]&~m[373]&m[374])|(~m[344]&~m[370]&~m[371]&m[373]&m[374])|(m[344]&~m[370]&~m[371]&m[373]&m[374])|(~m[344]&m[370]&~m[371]&m[373]&m[374])|(m[344]&m[370]&~m[371]&m[373]&m[374])|(~m[344]&~m[370]&m[371]&m[373]&m[374])|(m[344]&~m[370]&m[371]&m[373]&m[374])|(m[344]&m[370]&m[371]&m[373]&m[374]));
    m[382] = (((m[349]&~m[380]&~m[381]&~m[383]&~m[384])|(~m[349]&~m[380]&~m[381]&m[383]&~m[384])|(m[349]&m[380]&~m[381]&m[383]&~m[384])|(m[349]&~m[380]&m[381]&m[383]&~m[384])|(~m[349]&m[380]&~m[381]&~m[383]&m[384])|(~m[349]&~m[380]&m[381]&~m[383]&m[384])|(m[349]&m[380]&m[381]&~m[383]&m[384])|(~m[349]&m[380]&m[381]&m[383]&m[384]))&UnbiasedRNG[92])|((m[349]&~m[380]&~m[381]&m[383]&~m[384])|(~m[349]&~m[380]&~m[381]&~m[383]&m[384])|(m[349]&~m[380]&~m[381]&~m[383]&m[384])|(m[349]&m[380]&~m[381]&~m[383]&m[384])|(m[349]&~m[380]&m[381]&~m[383]&m[384])|(~m[349]&~m[380]&~m[381]&m[383]&m[384])|(m[349]&~m[380]&~m[381]&m[383]&m[384])|(~m[349]&m[380]&~m[381]&m[383]&m[384])|(m[349]&m[380]&~m[381]&m[383]&m[384])|(~m[349]&~m[380]&m[381]&m[383]&m[384])|(m[349]&~m[380]&m[381]&m[383]&m[384])|(m[349]&m[380]&m[381]&m[383]&m[384]));
    m[387] = (((m[354]&~m[385]&~m[386]&~m[388]&~m[389])|(~m[354]&~m[385]&~m[386]&m[388]&~m[389])|(m[354]&m[385]&~m[386]&m[388]&~m[389])|(m[354]&~m[385]&m[386]&m[388]&~m[389])|(~m[354]&m[385]&~m[386]&~m[388]&m[389])|(~m[354]&~m[385]&m[386]&~m[388]&m[389])|(m[354]&m[385]&m[386]&~m[388]&m[389])|(~m[354]&m[385]&m[386]&m[388]&m[389]))&UnbiasedRNG[93])|((m[354]&~m[385]&~m[386]&m[388]&~m[389])|(~m[354]&~m[385]&~m[386]&~m[388]&m[389])|(m[354]&~m[385]&~m[386]&~m[388]&m[389])|(m[354]&m[385]&~m[386]&~m[388]&m[389])|(m[354]&~m[385]&m[386]&~m[388]&m[389])|(~m[354]&~m[385]&~m[386]&m[388]&m[389])|(m[354]&~m[385]&~m[386]&m[388]&m[389])|(~m[354]&m[385]&~m[386]&m[388]&m[389])|(m[354]&m[385]&~m[386]&m[388]&m[389])|(~m[354]&~m[385]&m[386]&m[388]&m[389])|(m[354]&~m[385]&m[386]&m[388]&m[389])|(m[354]&m[385]&m[386]&m[388]&m[389]));
    m[392] = (((m[359]&~m[390]&~m[391]&~m[393]&~m[394])|(~m[359]&~m[390]&~m[391]&m[393]&~m[394])|(m[359]&m[390]&~m[391]&m[393]&~m[394])|(m[359]&~m[390]&m[391]&m[393]&~m[394])|(~m[359]&m[390]&~m[391]&~m[393]&m[394])|(~m[359]&~m[390]&m[391]&~m[393]&m[394])|(m[359]&m[390]&m[391]&~m[393]&m[394])|(~m[359]&m[390]&m[391]&m[393]&m[394]))&UnbiasedRNG[94])|((m[359]&~m[390]&~m[391]&m[393]&~m[394])|(~m[359]&~m[390]&~m[391]&~m[393]&m[394])|(m[359]&~m[390]&~m[391]&~m[393]&m[394])|(m[359]&m[390]&~m[391]&~m[393]&m[394])|(m[359]&~m[390]&m[391]&~m[393]&m[394])|(~m[359]&~m[390]&~m[391]&m[393]&m[394])|(m[359]&~m[390]&~m[391]&m[393]&m[394])|(~m[359]&m[390]&~m[391]&m[393]&m[394])|(m[359]&m[390]&~m[391]&m[393]&m[394])|(~m[359]&~m[390]&m[391]&m[393]&m[394])|(m[359]&~m[390]&m[391]&m[393]&m[394])|(m[359]&m[390]&m[391]&m[393]&m[394]));
    m[397] = (((m[364]&~m[395]&~m[396]&~m[398]&~m[399])|(~m[364]&~m[395]&~m[396]&m[398]&~m[399])|(m[364]&m[395]&~m[396]&m[398]&~m[399])|(m[364]&~m[395]&m[396]&m[398]&~m[399])|(~m[364]&m[395]&~m[396]&~m[398]&m[399])|(~m[364]&~m[395]&m[396]&~m[398]&m[399])|(m[364]&m[395]&m[396]&~m[398]&m[399])|(~m[364]&m[395]&m[396]&m[398]&m[399]))&UnbiasedRNG[95])|((m[364]&~m[395]&~m[396]&m[398]&~m[399])|(~m[364]&~m[395]&~m[396]&~m[398]&m[399])|(m[364]&~m[395]&~m[396]&~m[398]&m[399])|(m[364]&m[395]&~m[396]&~m[398]&m[399])|(m[364]&~m[395]&m[396]&~m[398]&m[399])|(~m[364]&~m[395]&~m[396]&m[398]&m[399])|(m[364]&~m[395]&~m[396]&m[398]&m[399])|(~m[364]&m[395]&~m[396]&m[398]&m[399])|(m[364]&m[395]&~m[396]&m[398]&m[399])|(~m[364]&~m[395]&m[396]&m[398]&m[399])|(m[364]&~m[395]&m[396]&m[398]&m[399])|(m[364]&m[395]&m[396]&m[398]&m[399]));
    m[402] = (((m[369]&~m[400]&~m[401]&~m[403]&~m[404])|(~m[369]&~m[400]&~m[401]&m[403]&~m[404])|(m[369]&m[400]&~m[401]&m[403]&~m[404])|(m[369]&~m[400]&m[401]&m[403]&~m[404])|(~m[369]&m[400]&~m[401]&~m[403]&m[404])|(~m[369]&~m[400]&m[401]&~m[403]&m[404])|(m[369]&m[400]&m[401]&~m[403]&m[404])|(~m[369]&m[400]&m[401]&m[403]&m[404]))&UnbiasedRNG[96])|((m[369]&~m[400]&~m[401]&m[403]&~m[404])|(~m[369]&~m[400]&~m[401]&~m[403]&m[404])|(m[369]&~m[400]&~m[401]&~m[403]&m[404])|(m[369]&m[400]&~m[401]&~m[403]&m[404])|(m[369]&~m[400]&m[401]&~m[403]&m[404])|(~m[369]&~m[400]&~m[401]&m[403]&m[404])|(m[369]&~m[400]&~m[401]&m[403]&m[404])|(~m[369]&m[400]&~m[401]&m[403]&m[404])|(m[369]&m[400]&~m[401]&m[403]&m[404])|(~m[369]&~m[400]&m[401]&m[403]&m[404])|(m[369]&~m[400]&m[401]&m[403]&m[404])|(m[369]&m[400]&m[401]&m[403]&m[404]));
    m[407] = (((m[374]&~m[405]&~m[406]&~m[408]&~m[409])|(~m[374]&~m[405]&~m[406]&m[408]&~m[409])|(m[374]&m[405]&~m[406]&m[408]&~m[409])|(m[374]&~m[405]&m[406]&m[408]&~m[409])|(~m[374]&m[405]&~m[406]&~m[408]&m[409])|(~m[374]&~m[405]&m[406]&~m[408]&m[409])|(m[374]&m[405]&m[406]&~m[408]&m[409])|(~m[374]&m[405]&m[406]&m[408]&m[409]))&UnbiasedRNG[97])|((m[374]&~m[405]&~m[406]&m[408]&~m[409])|(~m[374]&~m[405]&~m[406]&~m[408]&m[409])|(m[374]&~m[405]&~m[406]&~m[408]&m[409])|(m[374]&m[405]&~m[406]&~m[408]&m[409])|(m[374]&~m[405]&m[406]&~m[408]&m[409])|(~m[374]&~m[405]&~m[406]&m[408]&m[409])|(m[374]&~m[405]&~m[406]&m[408]&m[409])|(~m[374]&m[405]&~m[406]&m[408]&m[409])|(m[374]&m[405]&~m[406]&m[408]&m[409])|(~m[374]&~m[405]&m[406]&m[408]&m[409])|(m[374]&~m[405]&m[406]&m[408]&m[409])|(m[374]&m[405]&m[406]&m[408]&m[409]));
    m[412] = (((m[379]&~m[410]&~m[411]&~m[413]&~m[414])|(~m[379]&~m[410]&~m[411]&m[413]&~m[414])|(m[379]&m[410]&~m[411]&m[413]&~m[414])|(m[379]&~m[410]&m[411]&m[413]&~m[414])|(~m[379]&m[410]&~m[411]&~m[413]&m[414])|(~m[379]&~m[410]&m[411]&~m[413]&m[414])|(m[379]&m[410]&m[411]&~m[413]&m[414])|(~m[379]&m[410]&m[411]&m[413]&m[414]))&UnbiasedRNG[98])|((m[379]&~m[410]&~m[411]&m[413]&~m[414])|(~m[379]&~m[410]&~m[411]&~m[413]&m[414])|(m[379]&~m[410]&~m[411]&~m[413]&m[414])|(m[379]&m[410]&~m[411]&~m[413]&m[414])|(m[379]&~m[410]&m[411]&~m[413]&m[414])|(~m[379]&~m[410]&~m[411]&m[413]&m[414])|(m[379]&~m[410]&~m[411]&m[413]&m[414])|(~m[379]&m[410]&~m[411]&m[413]&m[414])|(m[379]&m[410]&~m[411]&m[413]&m[414])|(~m[379]&~m[410]&m[411]&m[413]&m[414])|(m[379]&~m[410]&m[411]&m[413]&m[414])|(m[379]&m[410]&m[411]&m[413]&m[414]));
    m[417] = (((m[389]&~m[415]&~m[416]&~m[418]&~m[419])|(~m[389]&~m[415]&~m[416]&m[418]&~m[419])|(m[389]&m[415]&~m[416]&m[418]&~m[419])|(m[389]&~m[415]&m[416]&m[418]&~m[419])|(~m[389]&m[415]&~m[416]&~m[418]&m[419])|(~m[389]&~m[415]&m[416]&~m[418]&m[419])|(m[389]&m[415]&m[416]&~m[418]&m[419])|(~m[389]&m[415]&m[416]&m[418]&m[419]))&UnbiasedRNG[99])|((m[389]&~m[415]&~m[416]&m[418]&~m[419])|(~m[389]&~m[415]&~m[416]&~m[418]&m[419])|(m[389]&~m[415]&~m[416]&~m[418]&m[419])|(m[389]&m[415]&~m[416]&~m[418]&m[419])|(m[389]&~m[415]&m[416]&~m[418]&m[419])|(~m[389]&~m[415]&~m[416]&m[418]&m[419])|(m[389]&~m[415]&~m[416]&m[418]&m[419])|(~m[389]&m[415]&~m[416]&m[418]&m[419])|(m[389]&m[415]&~m[416]&m[418]&m[419])|(~m[389]&~m[415]&m[416]&m[418]&m[419])|(m[389]&~m[415]&m[416]&m[418]&m[419])|(m[389]&m[415]&m[416]&m[418]&m[419]));
    m[422] = (((m[394]&~m[420]&~m[421]&~m[423]&~m[424])|(~m[394]&~m[420]&~m[421]&m[423]&~m[424])|(m[394]&m[420]&~m[421]&m[423]&~m[424])|(m[394]&~m[420]&m[421]&m[423]&~m[424])|(~m[394]&m[420]&~m[421]&~m[423]&m[424])|(~m[394]&~m[420]&m[421]&~m[423]&m[424])|(m[394]&m[420]&m[421]&~m[423]&m[424])|(~m[394]&m[420]&m[421]&m[423]&m[424]))&UnbiasedRNG[100])|((m[394]&~m[420]&~m[421]&m[423]&~m[424])|(~m[394]&~m[420]&~m[421]&~m[423]&m[424])|(m[394]&~m[420]&~m[421]&~m[423]&m[424])|(m[394]&m[420]&~m[421]&~m[423]&m[424])|(m[394]&~m[420]&m[421]&~m[423]&m[424])|(~m[394]&~m[420]&~m[421]&m[423]&m[424])|(m[394]&~m[420]&~m[421]&m[423]&m[424])|(~m[394]&m[420]&~m[421]&m[423]&m[424])|(m[394]&m[420]&~m[421]&m[423]&m[424])|(~m[394]&~m[420]&m[421]&m[423]&m[424])|(m[394]&~m[420]&m[421]&m[423]&m[424])|(m[394]&m[420]&m[421]&m[423]&m[424]));
    m[427] = (((m[399]&~m[425]&~m[426]&~m[428]&~m[429])|(~m[399]&~m[425]&~m[426]&m[428]&~m[429])|(m[399]&m[425]&~m[426]&m[428]&~m[429])|(m[399]&~m[425]&m[426]&m[428]&~m[429])|(~m[399]&m[425]&~m[426]&~m[428]&m[429])|(~m[399]&~m[425]&m[426]&~m[428]&m[429])|(m[399]&m[425]&m[426]&~m[428]&m[429])|(~m[399]&m[425]&m[426]&m[428]&m[429]))&UnbiasedRNG[101])|((m[399]&~m[425]&~m[426]&m[428]&~m[429])|(~m[399]&~m[425]&~m[426]&~m[428]&m[429])|(m[399]&~m[425]&~m[426]&~m[428]&m[429])|(m[399]&m[425]&~m[426]&~m[428]&m[429])|(m[399]&~m[425]&m[426]&~m[428]&m[429])|(~m[399]&~m[425]&~m[426]&m[428]&m[429])|(m[399]&~m[425]&~m[426]&m[428]&m[429])|(~m[399]&m[425]&~m[426]&m[428]&m[429])|(m[399]&m[425]&~m[426]&m[428]&m[429])|(~m[399]&~m[425]&m[426]&m[428]&m[429])|(m[399]&~m[425]&m[426]&m[428]&m[429])|(m[399]&m[425]&m[426]&m[428]&m[429]));
    m[432] = (((m[404]&~m[430]&~m[431]&~m[433]&~m[434])|(~m[404]&~m[430]&~m[431]&m[433]&~m[434])|(m[404]&m[430]&~m[431]&m[433]&~m[434])|(m[404]&~m[430]&m[431]&m[433]&~m[434])|(~m[404]&m[430]&~m[431]&~m[433]&m[434])|(~m[404]&~m[430]&m[431]&~m[433]&m[434])|(m[404]&m[430]&m[431]&~m[433]&m[434])|(~m[404]&m[430]&m[431]&m[433]&m[434]))&UnbiasedRNG[102])|((m[404]&~m[430]&~m[431]&m[433]&~m[434])|(~m[404]&~m[430]&~m[431]&~m[433]&m[434])|(m[404]&~m[430]&~m[431]&~m[433]&m[434])|(m[404]&m[430]&~m[431]&~m[433]&m[434])|(m[404]&~m[430]&m[431]&~m[433]&m[434])|(~m[404]&~m[430]&~m[431]&m[433]&m[434])|(m[404]&~m[430]&~m[431]&m[433]&m[434])|(~m[404]&m[430]&~m[431]&m[433]&m[434])|(m[404]&m[430]&~m[431]&m[433]&m[434])|(~m[404]&~m[430]&m[431]&m[433]&m[434])|(m[404]&~m[430]&m[431]&m[433]&m[434])|(m[404]&m[430]&m[431]&m[433]&m[434]));
    m[437] = (((m[409]&~m[435]&~m[436]&~m[438]&~m[439])|(~m[409]&~m[435]&~m[436]&m[438]&~m[439])|(m[409]&m[435]&~m[436]&m[438]&~m[439])|(m[409]&~m[435]&m[436]&m[438]&~m[439])|(~m[409]&m[435]&~m[436]&~m[438]&m[439])|(~m[409]&~m[435]&m[436]&~m[438]&m[439])|(m[409]&m[435]&m[436]&~m[438]&m[439])|(~m[409]&m[435]&m[436]&m[438]&m[439]))&UnbiasedRNG[103])|((m[409]&~m[435]&~m[436]&m[438]&~m[439])|(~m[409]&~m[435]&~m[436]&~m[438]&m[439])|(m[409]&~m[435]&~m[436]&~m[438]&m[439])|(m[409]&m[435]&~m[436]&~m[438]&m[439])|(m[409]&~m[435]&m[436]&~m[438]&m[439])|(~m[409]&~m[435]&~m[436]&m[438]&m[439])|(m[409]&~m[435]&~m[436]&m[438]&m[439])|(~m[409]&m[435]&~m[436]&m[438]&m[439])|(m[409]&m[435]&~m[436]&m[438]&m[439])|(~m[409]&~m[435]&m[436]&m[438]&m[439])|(m[409]&~m[435]&m[436]&m[438]&m[439])|(m[409]&m[435]&m[436]&m[438]&m[439]));
    m[442] = (((m[414]&~m[440]&~m[441]&~m[443]&~m[444])|(~m[414]&~m[440]&~m[441]&m[443]&~m[444])|(m[414]&m[440]&~m[441]&m[443]&~m[444])|(m[414]&~m[440]&m[441]&m[443]&~m[444])|(~m[414]&m[440]&~m[441]&~m[443]&m[444])|(~m[414]&~m[440]&m[441]&~m[443]&m[444])|(m[414]&m[440]&m[441]&~m[443]&m[444])|(~m[414]&m[440]&m[441]&m[443]&m[444]))&UnbiasedRNG[104])|((m[414]&~m[440]&~m[441]&m[443]&~m[444])|(~m[414]&~m[440]&~m[441]&~m[443]&m[444])|(m[414]&~m[440]&~m[441]&~m[443]&m[444])|(m[414]&m[440]&~m[441]&~m[443]&m[444])|(m[414]&~m[440]&m[441]&~m[443]&m[444])|(~m[414]&~m[440]&~m[441]&m[443]&m[444])|(m[414]&~m[440]&~m[441]&m[443]&m[444])|(~m[414]&m[440]&~m[441]&m[443]&m[444])|(m[414]&m[440]&~m[441]&m[443]&m[444])|(~m[414]&~m[440]&m[441]&m[443]&m[444])|(m[414]&~m[440]&m[441]&m[443]&m[444])|(m[414]&m[440]&m[441]&m[443]&m[444]));
    m[447] = (((m[424]&~m[445]&~m[446]&~m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&m[448]&~m[449])|(m[424]&m[445]&~m[446]&m[448]&~m[449])|(m[424]&~m[445]&m[446]&m[448]&~m[449])|(~m[424]&m[445]&~m[446]&~m[448]&m[449])|(~m[424]&~m[445]&m[446]&~m[448]&m[449])|(m[424]&m[445]&m[446]&~m[448]&m[449])|(~m[424]&m[445]&m[446]&m[448]&m[449]))&UnbiasedRNG[105])|((m[424]&~m[445]&~m[446]&m[448]&~m[449])|(~m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&~m[446]&~m[448]&m[449])|(m[424]&m[445]&~m[446]&~m[448]&m[449])|(m[424]&~m[445]&m[446]&~m[448]&m[449])|(~m[424]&~m[445]&~m[446]&m[448]&m[449])|(m[424]&~m[445]&~m[446]&m[448]&m[449])|(~m[424]&m[445]&~m[446]&m[448]&m[449])|(m[424]&m[445]&~m[446]&m[448]&m[449])|(~m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&~m[445]&m[446]&m[448]&m[449])|(m[424]&m[445]&m[446]&m[448]&m[449]));
    m[452] = (((m[429]&~m[450]&~m[451]&~m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&m[453]&~m[454])|(m[429]&m[450]&~m[451]&m[453]&~m[454])|(m[429]&~m[450]&m[451]&m[453]&~m[454])|(~m[429]&m[450]&~m[451]&~m[453]&m[454])|(~m[429]&~m[450]&m[451]&~m[453]&m[454])|(m[429]&m[450]&m[451]&~m[453]&m[454])|(~m[429]&m[450]&m[451]&m[453]&m[454]))&UnbiasedRNG[106])|((m[429]&~m[450]&~m[451]&m[453]&~m[454])|(~m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&~m[451]&~m[453]&m[454])|(m[429]&m[450]&~m[451]&~m[453]&m[454])|(m[429]&~m[450]&m[451]&~m[453]&m[454])|(~m[429]&~m[450]&~m[451]&m[453]&m[454])|(m[429]&~m[450]&~m[451]&m[453]&m[454])|(~m[429]&m[450]&~m[451]&m[453]&m[454])|(m[429]&m[450]&~m[451]&m[453]&m[454])|(~m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&~m[450]&m[451]&m[453]&m[454])|(m[429]&m[450]&m[451]&m[453]&m[454]));
    m[457] = (((m[434]&~m[455]&~m[456]&~m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&m[458]&~m[459])|(m[434]&m[455]&~m[456]&m[458]&~m[459])|(m[434]&~m[455]&m[456]&m[458]&~m[459])|(~m[434]&m[455]&~m[456]&~m[458]&m[459])|(~m[434]&~m[455]&m[456]&~m[458]&m[459])|(m[434]&m[455]&m[456]&~m[458]&m[459])|(~m[434]&m[455]&m[456]&m[458]&m[459]))&UnbiasedRNG[107])|((m[434]&~m[455]&~m[456]&m[458]&~m[459])|(~m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&~m[456]&~m[458]&m[459])|(m[434]&m[455]&~m[456]&~m[458]&m[459])|(m[434]&~m[455]&m[456]&~m[458]&m[459])|(~m[434]&~m[455]&~m[456]&m[458]&m[459])|(m[434]&~m[455]&~m[456]&m[458]&m[459])|(~m[434]&m[455]&~m[456]&m[458]&m[459])|(m[434]&m[455]&~m[456]&m[458]&m[459])|(~m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&~m[455]&m[456]&m[458]&m[459])|(m[434]&m[455]&m[456]&m[458]&m[459]));
    m[462] = (((m[439]&~m[460]&~m[461]&~m[463]&~m[464])|(~m[439]&~m[460]&~m[461]&m[463]&~m[464])|(m[439]&m[460]&~m[461]&m[463]&~m[464])|(m[439]&~m[460]&m[461]&m[463]&~m[464])|(~m[439]&m[460]&~m[461]&~m[463]&m[464])|(~m[439]&~m[460]&m[461]&~m[463]&m[464])|(m[439]&m[460]&m[461]&~m[463]&m[464])|(~m[439]&m[460]&m[461]&m[463]&m[464]))&UnbiasedRNG[108])|((m[439]&~m[460]&~m[461]&m[463]&~m[464])|(~m[439]&~m[460]&~m[461]&~m[463]&m[464])|(m[439]&~m[460]&~m[461]&~m[463]&m[464])|(m[439]&m[460]&~m[461]&~m[463]&m[464])|(m[439]&~m[460]&m[461]&~m[463]&m[464])|(~m[439]&~m[460]&~m[461]&m[463]&m[464])|(m[439]&~m[460]&~m[461]&m[463]&m[464])|(~m[439]&m[460]&~m[461]&m[463]&m[464])|(m[439]&m[460]&~m[461]&m[463]&m[464])|(~m[439]&~m[460]&m[461]&m[463]&m[464])|(m[439]&~m[460]&m[461]&m[463]&m[464])|(m[439]&m[460]&m[461]&m[463]&m[464]));
    m[467] = (((m[444]&~m[465]&~m[466]&~m[468]&~m[469])|(~m[444]&~m[465]&~m[466]&m[468]&~m[469])|(m[444]&m[465]&~m[466]&m[468]&~m[469])|(m[444]&~m[465]&m[466]&m[468]&~m[469])|(~m[444]&m[465]&~m[466]&~m[468]&m[469])|(~m[444]&~m[465]&m[466]&~m[468]&m[469])|(m[444]&m[465]&m[466]&~m[468]&m[469])|(~m[444]&m[465]&m[466]&m[468]&m[469]))&UnbiasedRNG[109])|((m[444]&~m[465]&~m[466]&m[468]&~m[469])|(~m[444]&~m[465]&~m[466]&~m[468]&m[469])|(m[444]&~m[465]&~m[466]&~m[468]&m[469])|(m[444]&m[465]&~m[466]&~m[468]&m[469])|(m[444]&~m[465]&m[466]&~m[468]&m[469])|(~m[444]&~m[465]&~m[466]&m[468]&m[469])|(m[444]&~m[465]&~m[466]&m[468]&m[469])|(~m[444]&m[465]&~m[466]&m[468]&m[469])|(m[444]&m[465]&~m[466]&m[468]&m[469])|(~m[444]&~m[465]&m[466]&m[468]&m[469])|(m[444]&~m[465]&m[466]&m[468]&m[469])|(m[444]&m[465]&m[466]&m[468]&m[469]));
    m[472] = (((m[454]&~m[470]&~m[471]&~m[473]&~m[474])|(~m[454]&~m[470]&~m[471]&m[473]&~m[474])|(m[454]&m[470]&~m[471]&m[473]&~m[474])|(m[454]&~m[470]&m[471]&m[473]&~m[474])|(~m[454]&m[470]&~m[471]&~m[473]&m[474])|(~m[454]&~m[470]&m[471]&~m[473]&m[474])|(m[454]&m[470]&m[471]&~m[473]&m[474])|(~m[454]&m[470]&m[471]&m[473]&m[474]))&UnbiasedRNG[110])|((m[454]&~m[470]&~m[471]&m[473]&~m[474])|(~m[454]&~m[470]&~m[471]&~m[473]&m[474])|(m[454]&~m[470]&~m[471]&~m[473]&m[474])|(m[454]&m[470]&~m[471]&~m[473]&m[474])|(m[454]&~m[470]&m[471]&~m[473]&m[474])|(~m[454]&~m[470]&~m[471]&m[473]&m[474])|(m[454]&~m[470]&~m[471]&m[473]&m[474])|(~m[454]&m[470]&~m[471]&m[473]&m[474])|(m[454]&m[470]&~m[471]&m[473]&m[474])|(~m[454]&~m[470]&m[471]&m[473]&m[474])|(m[454]&~m[470]&m[471]&m[473]&m[474])|(m[454]&m[470]&m[471]&m[473]&m[474]));
    m[477] = (((m[459]&~m[475]&~m[476]&~m[478]&~m[479])|(~m[459]&~m[475]&~m[476]&m[478]&~m[479])|(m[459]&m[475]&~m[476]&m[478]&~m[479])|(m[459]&~m[475]&m[476]&m[478]&~m[479])|(~m[459]&m[475]&~m[476]&~m[478]&m[479])|(~m[459]&~m[475]&m[476]&~m[478]&m[479])|(m[459]&m[475]&m[476]&~m[478]&m[479])|(~m[459]&m[475]&m[476]&m[478]&m[479]))&UnbiasedRNG[111])|((m[459]&~m[475]&~m[476]&m[478]&~m[479])|(~m[459]&~m[475]&~m[476]&~m[478]&m[479])|(m[459]&~m[475]&~m[476]&~m[478]&m[479])|(m[459]&m[475]&~m[476]&~m[478]&m[479])|(m[459]&~m[475]&m[476]&~m[478]&m[479])|(~m[459]&~m[475]&~m[476]&m[478]&m[479])|(m[459]&~m[475]&~m[476]&m[478]&m[479])|(~m[459]&m[475]&~m[476]&m[478]&m[479])|(m[459]&m[475]&~m[476]&m[478]&m[479])|(~m[459]&~m[475]&m[476]&m[478]&m[479])|(m[459]&~m[475]&m[476]&m[478]&m[479])|(m[459]&m[475]&m[476]&m[478]&m[479]));
    m[482] = (((m[464]&~m[480]&~m[481]&~m[483]&~m[484])|(~m[464]&~m[480]&~m[481]&m[483]&~m[484])|(m[464]&m[480]&~m[481]&m[483]&~m[484])|(m[464]&~m[480]&m[481]&m[483]&~m[484])|(~m[464]&m[480]&~m[481]&~m[483]&m[484])|(~m[464]&~m[480]&m[481]&~m[483]&m[484])|(m[464]&m[480]&m[481]&~m[483]&m[484])|(~m[464]&m[480]&m[481]&m[483]&m[484]))&UnbiasedRNG[112])|((m[464]&~m[480]&~m[481]&m[483]&~m[484])|(~m[464]&~m[480]&~m[481]&~m[483]&m[484])|(m[464]&~m[480]&~m[481]&~m[483]&m[484])|(m[464]&m[480]&~m[481]&~m[483]&m[484])|(m[464]&~m[480]&m[481]&~m[483]&m[484])|(~m[464]&~m[480]&~m[481]&m[483]&m[484])|(m[464]&~m[480]&~m[481]&m[483]&m[484])|(~m[464]&m[480]&~m[481]&m[483]&m[484])|(m[464]&m[480]&~m[481]&m[483]&m[484])|(~m[464]&~m[480]&m[481]&m[483]&m[484])|(m[464]&~m[480]&m[481]&m[483]&m[484])|(m[464]&m[480]&m[481]&m[483]&m[484]));
    m[487] = (((m[469]&~m[485]&~m[486]&~m[488]&~m[489])|(~m[469]&~m[485]&~m[486]&m[488]&~m[489])|(m[469]&m[485]&~m[486]&m[488]&~m[489])|(m[469]&~m[485]&m[486]&m[488]&~m[489])|(~m[469]&m[485]&~m[486]&~m[488]&m[489])|(~m[469]&~m[485]&m[486]&~m[488]&m[489])|(m[469]&m[485]&m[486]&~m[488]&m[489])|(~m[469]&m[485]&m[486]&m[488]&m[489]))&UnbiasedRNG[113])|((m[469]&~m[485]&~m[486]&m[488]&~m[489])|(~m[469]&~m[485]&~m[486]&~m[488]&m[489])|(m[469]&~m[485]&~m[486]&~m[488]&m[489])|(m[469]&m[485]&~m[486]&~m[488]&m[489])|(m[469]&~m[485]&m[486]&~m[488]&m[489])|(~m[469]&~m[485]&~m[486]&m[488]&m[489])|(m[469]&~m[485]&~m[486]&m[488]&m[489])|(~m[469]&m[485]&~m[486]&m[488]&m[489])|(m[469]&m[485]&~m[486]&m[488]&m[489])|(~m[469]&~m[485]&m[486]&m[488]&m[489])|(m[469]&~m[485]&m[486]&m[488]&m[489])|(m[469]&m[485]&m[486]&m[488]&m[489]));
    m[492] = (((m[479]&~m[490]&~m[491]&~m[493]&~m[494])|(~m[479]&~m[490]&~m[491]&m[493]&~m[494])|(m[479]&m[490]&~m[491]&m[493]&~m[494])|(m[479]&~m[490]&m[491]&m[493]&~m[494])|(~m[479]&m[490]&~m[491]&~m[493]&m[494])|(~m[479]&~m[490]&m[491]&~m[493]&m[494])|(m[479]&m[490]&m[491]&~m[493]&m[494])|(~m[479]&m[490]&m[491]&m[493]&m[494]))&UnbiasedRNG[114])|((m[479]&~m[490]&~m[491]&m[493]&~m[494])|(~m[479]&~m[490]&~m[491]&~m[493]&m[494])|(m[479]&~m[490]&~m[491]&~m[493]&m[494])|(m[479]&m[490]&~m[491]&~m[493]&m[494])|(m[479]&~m[490]&m[491]&~m[493]&m[494])|(~m[479]&~m[490]&~m[491]&m[493]&m[494])|(m[479]&~m[490]&~m[491]&m[493]&m[494])|(~m[479]&m[490]&~m[491]&m[493]&m[494])|(m[479]&m[490]&~m[491]&m[493]&m[494])|(~m[479]&~m[490]&m[491]&m[493]&m[494])|(m[479]&~m[490]&m[491]&m[493]&m[494])|(m[479]&m[490]&m[491]&m[493]&m[494]));
    m[497] = (((m[484]&~m[495]&~m[496]&~m[498]&~m[499])|(~m[484]&~m[495]&~m[496]&m[498]&~m[499])|(m[484]&m[495]&~m[496]&m[498]&~m[499])|(m[484]&~m[495]&m[496]&m[498]&~m[499])|(~m[484]&m[495]&~m[496]&~m[498]&m[499])|(~m[484]&~m[495]&m[496]&~m[498]&m[499])|(m[484]&m[495]&m[496]&~m[498]&m[499])|(~m[484]&m[495]&m[496]&m[498]&m[499]))&UnbiasedRNG[115])|((m[484]&~m[495]&~m[496]&m[498]&~m[499])|(~m[484]&~m[495]&~m[496]&~m[498]&m[499])|(m[484]&~m[495]&~m[496]&~m[498]&m[499])|(m[484]&m[495]&~m[496]&~m[498]&m[499])|(m[484]&~m[495]&m[496]&~m[498]&m[499])|(~m[484]&~m[495]&~m[496]&m[498]&m[499])|(m[484]&~m[495]&~m[496]&m[498]&m[499])|(~m[484]&m[495]&~m[496]&m[498]&m[499])|(m[484]&m[495]&~m[496]&m[498]&m[499])|(~m[484]&~m[495]&m[496]&m[498]&m[499])|(m[484]&~m[495]&m[496]&m[498]&m[499])|(m[484]&m[495]&m[496]&m[498]&m[499]));
    m[502] = (((m[489]&~m[500]&~m[501]&~m[503]&~m[504])|(~m[489]&~m[500]&~m[501]&m[503]&~m[504])|(m[489]&m[500]&~m[501]&m[503]&~m[504])|(m[489]&~m[500]&m[501]&m[503]&~m[504])|(~m[489]&m[500]&~m[501]&~m[503]&m[504])|(~m[489]&~m[500]&m[501]&~m[503]&m[504])|(m[489]&m[500]&m[501]&~m[503]&m[504])|(~m[489]&m[500]&m[501]&m[503]&m[504]))&UnbiasedRNG[116])|((m[489]&~m[500]&~m[501]&m[503]&~m[504])|(~m[489]&~m[500]&~m[501]&~m[503]&m[504])|(m[489]&~m[500]&~m[501]&~m[503]&m[504])|(m[489]&m[500]&~m[501]&~m[503]&m[504])|(m[489]&~m[500]&m[501]&~m[503]&m[504])|(~m[489]&~m[500]&~m[501]&m[503]&m[504])|(m[489]&~m[500]&~m[501]&m[503]&m[504])|(~m[489]&m[500]&~m[501]&m[503]&m[504])|(m[489]&m[500]&~m[501]&m[503]&m[504])|(~m[489]&~m[500]&m[501]&m[503]&m[504])|(m[489]&~m[500]&m[501]&m[503]&m[504])|(m[489]&m[500]&m[501]&m[503]&m[504]));
    m[507] = (((m[499]&~m[505]&~m[506]&~m[508]&~m[509])|(~m[499]&~m[505]&~m[506]&m[508]&~m[509])|(m[499]&m[505]&~m[506]&m[508]&~m[509])|(m[499]&~m[505]&m[506]&m[508]&~m[509])|(~m[499]&m[505]&~m[506]&~m[508]&m[509])|(~m[499]&~m[505]&m[506]&~m[508]&m[509])|(m[499]&m[505]&m[506]&~m[508]&m[509])|(~m[499]&m[505]&m[506]&m[508]&m[509]))&UnbiasedRNG[117])|((m[499]&~m[505]&~m[506]&m[508]&~m[509])|(~m[499]&~m[505]&~m[506]&~m[508]&m[509])|(m[499]&~m[505]&~m[506]&~m[508]&m[509])|(m[499]&m[505]&~m[506]&~m[508]&m[509])|(m[499]&~m[505]&m[506]&~m[508]&m[509])|(~m[499]&~m[505]&~m[506]&m[508]&m[509])|(m[499]&~m[505]&~m[506]&m[508]&m[509])|(~m[499]&m[505]&~m[506]&m[508]&m[509])|(m[499]&m[505]&~m[506]&m[508]&m[509])|(~m[499]&~m[505]&m[506]&m[508]&m[509])|(m[499]&~m[505]&m[506]&m[508]&m[509])|(m[499]&m[505]&m[506]&m[508]&m[509]));
    m[512] = (((m[504]&~m[510]&~m[511]&~m[513]&~m[514])|(~m[504]&~m[510]&~m[511]&m[513]&~m[514])|(m[504]&m[510]&~m[511]&m[513]&~m[514])|(m[504]&~m[510]&m[511]&m[513]&~m[514])|(~m[504]&m[510]&~m[511]&~m[513]&m[514])|(~m[504]&~m[510]&m[511]&~m[513]&m[514])|(m[504]&m[510]&m[511]&~m[513]&m[514])|(~m[504]&m[510]&m[511]&m[513]&m[514]))&UnbiasedRNG[118])|((m[504]&~m[510]&~m[511]&m[513]&~m[514])|(~m[504]&~m[510]&~m[511]&~m[513]&m[514])|(m[504]&~m[510]&~m[511]&~m[513]&m[514])|(m[504]&m[510]&~m[511]&~m[513]&m[514])|(m[504]&~m[510]&m[511]&~m[513]&m[514])|(~m[504]&~m[510]&~m[511]&m[513]&m[514])|(m[504]&~m[510]&~m[511]&m[513]&m[514])|(~m[504]&m[510]&~m[511]&m[513]&m[514])|(m[504]&m[510]&~m[511]&m[513]&m[514])|(~m[504]&~m[510]&m[511]&m[513]&m[514])|(m[504]&~m[510]&m[511]&m[513]&m[514])|(m[504]&m[510]&m[511]&m[513]&m[514]));
    m[517] = (((m[514]&~m[515]&~m[516]&~m[518]&~m[519])|(~m[514]&~m[515]&~m[516]&m[518]&~m[519])|(m[514]&m[515]&~m[516]&m[518]&~m[519])|(m[514]&~m[515]&m[516]&m[518]&~m[519])|(~m[514]&m[515]&~m[516]&~m[518]&m[519])|(~m[514]&~m[515]&m[516]&~m[518]&m[519])|(m[514]&m[515]&m[516]&~m[518]&m[519])|(~m[514]&m[515]&m[516]&m[518]&m[519]))&UnbiasedRNG[119])|((m[514]&~m[515]&~m[516]&m[518]&~m[519])|(~m[514]&~m[515]&~m[516]&~m[518]&m[519])|(m[514]&~m[515]&~m[516]&~m[518]&m[519])|(m[514]&m[515]&~m[516]&~m[518]&m[519])|(m[514]&~m[515]&m[516]&~m[518]&m[519])|(~m[514]&~m[515]&~m[516]&m[518]&m[519])|(m[514]&~m[515]&~m[516]&m[518]&m[519])|(~m[514]&m[515]&~m[516]&m[518]&m[519])|(m[514]&m[515]&~m[516]&m[518]&m[519])|(~m[514]&~m[515]&m[516]&m[518]&m[519])|(m[514]&~m[515]&m[516]&m[518]&m[519])|(m[514]&m[515]&m[516]&m[518]&m[519]));
end

always @(posedge color2_clk) begin
    m[112] = (((~m[32]&~m[48]&~m[176])|(m[32]&m[48]&~m[176]))&BiasedRNG[159])|(((m[32]&~m[48]&~m[176])|(~m[32]&m[48]&m[176]))&~BiasedRNG[159])|((~m[32]&~m[48]&m[176])|(m[32]&~m[48]&m[176])|(m[32]&m[48]&m[176]));
    m[113] = (((~m[32]&~m[56]&~m[177])|(m[32]&m[56]&~m[177]))&BiasedRNG[160])|(((m[32]&~m[56]&~m[177])|(~m[32]&m[56]&m[177]))&~BiasedRNG[160])|((~m[32]&~m[56]&m[177])|(m[32]&~m[56]&m[177])|(m[32]&m[56]&m[177]));
    m[114] = (((~m[32]&~m[64]&~m[178])|(m[32]&m[64]&~m[178]))&BiasedRNG[161])|(((m[32]&~m[64]&~m[178])|(~m[32]&m[64]&m[178]))&~BiasedRNG[161])|((~m[32]&~m[64]&m[178])|(m[32]&~m[64]&m[178])|(m[32]&m[64]&m[178]));
    m[115] = (((~m[32]&~m[72]&~m[179])|(m[32]&m[72]&~m[179]))&BiasedRNG[162])|(((m[32]&~m[72]&~m[179])|(~m[32]&m[72]&m[179]))&~BiasedRNG[162])|((~m[32]&~m[72]&m[179])|(m[32]&~m[72]&m[179])|(m[32]&m[72]&m[179]));
    m[116] = (((~m[33]&~m[80]&~m[180])|(m[33]&m[80]&~m[180]))&BiasedRNG[163])|(((m[33]&~m[80]&~m[180])|(~m[33]&m[80]&m[180]))&~BiasedRNG[163])|((~m[33]&~m[80]&m[180])|(m[33]&~m[80]&m[180])|(m[33]&m[80]&m[180]));
    m[117] = (((~m[33]&~m[88]&~m[181])|(m[33]&m[88]&~m[181]))&BiasedRNG[164])|(((m[33]&~m[88]&~m[181])|(~m[33]&m[88]&m[181]))&~BiasedRNG[164])|((~m[33]&~m[88]&m[181])|(m[33]&~m[88]&m[181])|(m[33]&m[88]&m[181]));
    m[118] = (((~m[33]&~m[96]&~m[182])|(m[33]&m[96]&~m[182]))&BiasedRNG[165])|(((m[33]&~m[96]&~m[182])|(~m[33]&m[96]&m[182]))&~BiasedRNG[165])|((~m[33]&~m[96]&m[182])|(m[33]&~m[96]&m[182])|(m[33]&m[96]&m[182]));
    m[119] = (((~m[33]&~m[104]&~m[183])|(m[33]&m[104]&~m[183]))&BiasedRNG[166])|(((m[33]&~m[104]&~m[183])|(~m[33]&m[104]&m[183]))&~BiasedRNG[166])|((~m[33]&~m[104]&m[183])|(m[33]&~m[104]&m[183])|(m[33]&m[104]&m[183]));
    m[120] = (((~m[34]&~m[49]&~m[184])|(m[34]&m[49]&~m[184]))&BiasedRNG[167])|(((m[34]&~m[49]&~m[184])|(~m[34]&m[49]&m[184]))&~BiasedRNG[167])|((~m[34]&~m[49]&m[184])|(m[34]&~m[49]&m[184])|(m[34]&m[49]&m[184]));
    m[121] = (((~m[34]&~m[57]&~m[185])|(m[34]&m[57]&~m[185]))&BiasedRNG[168])|(((m[34]&~m[57]&~m[185])|(~m[34]&m[57]&m[185]))&~BiasedRNG[168])|((~m[34]&~m[57]&m[185])|(m[34]&~m[57]&m[185])|(m[34]&m[57]&m[185]));
    m[122] = (((~m[34]&~m[65]&~m[186])|(m[34]&m[65]&~m[186]))&BiasedRNG[169])|(((m[34]&~m[65]&~m[186])|(~m[34]&m[65]&m[186]))&~BiasedRNG[169])|((~m[34]&~m[65]&m[186])|(m[34]&~m[65]&m[186])|(m[34]&m[65]&m[186]));
    m[123] = (((~m[34]&~m[73]&~m[187])|(m[34]&m[73]&~m[187]))&BiasedRNG[170])|(((m[34]&~m[73]&~m[187])|(~m[34]&m[73]&m[187]))&~BiasedRNG[170])|((~m[34]&~m[73]&m[187])|(m[34]&~m[73]&m[187])|(m[34]&m[73]&m[187]));
    m[124] = (((~m[35]&~m[81]&~m[188])|(m[35]&m[81]&~m[188]))&BiasedRNG[171])|(((m[35]&~m[81]&~m[188])|(~m[35]&m[81]&m[188]))&~BiasedRNG[171])|((~m[35]&~m[81]&m[188])|(m[35]&~m[81]&m[188])|(m[35]&m[81]&m[188]));
    m[125] = (((~m[35]&~m[89]&~m[189])|(m[35]&m[89]&~m[189]))&BiasedRNG[172])|(((m[35]&~m[89]&~m[189])|(~m[35]&m[89]&m[189]))&~BiasedRNG[172])|((~m[35]&~m[89]&m[189])|(m[35]&~m[89]&m[189])|(m[35]&m[89]&m[189]));
    m[126] = (((~m[35]&~m[97]&~m[190])|(m[35]&m[97]&~m[190]))&BiasedRNG[173])|(((m[35]&~m[97]&~m[190])|(~m[35]&m[97]&m[190]))&~BiasedRNG[173])|((~m[35]&~m[97]&m[190])|(m[35]&~m[97]&m[190])|(m[35]&m[97]&m[190]));
    m[127] = (((~m[35]&~m[105]&~m[191])|(m[35]&m[105]&~m[191]))&BiasedRNG[174])|(((m[35]&~m[105]&~m[191])|(~m[35]&m[105]&m[191]))&~BiasedRNG[174])|((~m[35]&~m[105]&m[191])|(m[35]&~m[105]&m[191])|(m[35]&m[105]&m[191]));
    m[128] = (((~m[36]&~m[50]&~m[192])|(m[36]&m[50]&~m[192]))&BiasedRNG[175])|(((m[36]&~m[50]&~m[192])|(~m[36]&m[50]&m[192]))&~BiasedRNG[175])|((~m[36]&~m[50]&m[192])|(m[36]&~m[50]&m[192])|(m[36]&m[50]&m[192]));
    m[129] = (((~m[36]&~m[58]&~m[193])|(m[36]&m[58]&~m[193]))&BiasedRNG[176])|(((m[36]&~m[58]&~m[193])|(~m[36]&m[58]&m[193]))&~BiasedRNG[176])|((~m[36]&~m[58]&m[193])|(m[36]&~m[58]&m[193])|(m[36]&m[58]&m[193]));
    m[130] = (((~m[36]&~m[66]&~m[194])|(m[36]&m[66]&~m[194]))&BiasedRNG[177])|(((m[36]&~m[66]&~m[194])|(~m[36]&m[66]&m[194]))&~BiasedRNG[177])|((~m[36]&~m[66]&m[194])|(m[36]&~m[66]&m[194])|(m[36]&m[66]&m[194]));
    m[131] = (((~m[36]&~m[74]&~m[195])|(m[36]&m[74]&~m[195]))&BiasedRNG[178])|(((m[36]&~m[74]&~m[195])|(~m[36]&m[74]&m[195]))&~BiasedRNG[178])|((~m[36]&~m[74]&m[195])|(m[36]&~m[74]&m[195])|(m[36]&m[74]&m[195]));
    m[132] = (((~m[37]&~m[82]&~m[196])|(m[37]&m[82]&~m[196]))&BiasedRNG[179])|(((m[37]&~m[82]&~m[196])|(~m[37]&m[82]&m[196]))&~BiasedRNG[179])|((~m[37]&~m[82]&m[196])|(m[37]&~m[82]&m[196])|(m[37]&m[82]&m[196]));
    m[133] = (((~m[37]&~m[90]&~m[197])|(m[37]&m[90]&~m[197]))&BiasedRNG[180])|(((m[37]&~m[90]&~m[197])|(~m[37]&m[90]&m[197]))&~BiasedRNG[180])|((~m[37]&~m[90]&m[197])|(m[37]&~m[90]&m[197])|(m[37]&m[90]&m[197]));
    m[134] = (((~m[37]&~m[98]&~m[198])|(m[37]&m[98]&~m[198]))&BiasedRNG[181])|(((m[37]&~m[98]&~m[198])|(~m[37]&m[98]&m[198]))&~BiasedRNG[181])|((~m[37]&~m[98]&m[198])|(m[37]&~m[98]&m[198])|(m[37]&m[98]&m[198]));
    m[135] = (((~m[37]&~m[106]&~m[199])|(m[37]&m[106]&~m[199]))&BiasedRNG[182])|(((m[37]&~m[106]&~m[199])|(~m[37]&m[106]&m[199]))&~BiasedRNG[182])|((~m[37]&~m[106]&m[199])|(m[37]&~m[106]&m[199])|(m[37]&m[106]&m[199]));
    m[136] = (((~m[38]&~m[51]&~m[200])|(m[38]&m[51]&~m[200]))&BiasedRNG[183])|(((m[38]&~m[51]&~m[200])|(~m[38]&m[51]&m[200]))&~BiasedRNG[183])|((~m[38]&~m[51]&m[200])|(m[38]&~m[51]&m[200])|(m[38]&m[51]&m[200]));
    m[137] = (((~m[38]&~m[59]&~m[201])|(m[38]&m[59]&~m[201]))&BiasedRNG[184])|(((m[38]&~m[59]&~m[201])|(~m[38]&m[59]&m[201]))&~BiasedRNG[184])|((~m[38]&~m[59]&m[201])|(m[38]&~m[59]&m[201])|(m[38]&m[59]&m[201]));
    m[138] = (((~m[38]&~m[67]&~m[202])|(m[38]&m[67]&~m[202]))&BiasedRNG[185])|(((m[38]&~m[67]&~m[202])|(~m[38]&m[67]&m[202]))&~BiasedRNG[185])|((~m[38]&~m[67]&m[202])|(m[38]&~m[67]&m[202])|(m[38]&m[67]&m[202]));
    m[139] = (((~m[38]&~m[75]&~m[203])|(m[38]&m[75]&~m[203]))&BiasedRNG[186])|(((m[38]&~m[75]&~m[203])|(~m[38]&m[75]&m[203]))&~BiasedRNG[186])|((~m[38]&~m[75]&m[203])|(m[38]&~m[75]&m[203])|(m[38]&m[75]&m[203]));
    m[140] = (((~m[39]&~m[83]&~m[204])|(m[39]&m[83]&~m[204]))&BiasedRNG[187])|(((m[39]&~m[83]&~m[204])|(~m[39]&m[83]&m[204]))&~BiasedRNG[187])|((~m[39]&~m[83]&m[204])|(m[39]&~m[83]&m[204])|(m[39]&m[83]&m[204]));
    m[141] = (((~m[39]&~m[91]&~m[205])|(m[39]&m[91]&~m[205]))&BiasedRNG[188])|(((m[39]&~m[91]&~m[205])|(~m[39]&m[91]&m[205]))&~BiasedRNG[188])|((~m[39]&~m[91]&m[205])|(m[39]&~m[91]&m[205])|(m[39]&m[91]&m[205]));
    m[142] = (((~m[39]&~m[99]&~m[206])|(m[39]&m[99]&~m[206]))&BiasedRNG[189])|(((m[39]&~m[99]&~m[206])|(~m[39]&m[99]&m[206]))&~BiasedRNG[189])|((~m[39]&~m[99]&m[206])|(m[39]&~m[99]&m[206])|(m[39]&m[99]&m[206]));
    m[143] = (((~m[39]&~m[107]&~m[207])|(m[39]&m[107]&~m[207]))&BiasedRNG[190])|(((m[39]&~m[107]&~m[207])|(~m[39]&m[107]&m[207]))&~BiasedRNG[190])|((~m[39]&~m[107]&m[207])|(m[39]&~m[107]&m[207])|(m[39]&m[107]&m[207]));
    m[144] = (((~m[40]&~m[52]&~m[208])|(m[40]&m[52]&~m[208]))&BiasedRNG[191])|(((m[40]&~m[52]&~m[208])|(~m[40]&m[52]&m[208]))&~BiasedRNG[191])|((~m[40]&~m[52]&m[208])|(m[40]&~m[52]&m[208])|(m[40]&m[52]&m[208]));
    m[145] = (((~m[40]&~m[60]&~m[209])|(m[40]&m[60]&~m[209]))&BiasedRNG[192])|(((m[40]&~m[60]&~m[209])|(~m[40]&m[60]&m[209]))&~BiasedRNG[192])|((~m[40]&~m[60]&m[209])|(m[40]&~m[60]&m[209])|(m[40]&m[60]&m[209]));
    m[146] = (((~m[40]&~m[68]&~m[210])|(m[40]&m[68]&~m[210]))&BiasedRNG[193])|(((m[40]&~m[68]&~m[210])|(~m[40]&m[68]&m[210]))&~BiasedRNG[193])|((~m[40]&~m[68]&m[210])|(m[40]&~m[68]&m[210])|(m[40]&m[68]&m[210]));
    m[147] = (((~m[40]&~m[76]&~m[211])|(m[40]&m[76]&~m[211]))&BiasedRNG[194])|(((m[40]&~m[76]&~m[211])|(~m[40]&m[76]&m[211]))&~BiasedRNG[194])|((~m[40]&~m[76]&m[211])|(m[40]&~m[76]&m[211])|(m[40]&m[76]&m[211]));
    m[148] = (((~m[41]&~m[84]&~m[212])|(m[41]&m[84]&~m[212]))&BiasedRNG[195])|(((m[41]&~m[84]&~m[212])|(~m[41]&m[84]&m[212]))&~BiasedRNG[195])|((~m[41]&~m[84]&m[212])|(m[41]&~m[84]&m[212])|(m[41]&m[84]&m[212]));
    m[149] = (((~m[41]&~m[92]&~m[213])|(m[41]&m[92]&~m[213]))&BiasedRNG[196])|(((m[41]&~m[92]&~m[213])|(~m[41]&m[92]&m[213]))&~BiasedRNG[196])|((~m[41]&~m[92]&m[213])|(m[41]&~m[92]&m[213])|(m[41]&m[92]&m[213]));
    m[150] = (((~m[41]&~m[100]&~m[214])|(m[41]&m[100]&~m[214]))&BiasedRNG[197])|(((m[41]&~m[100]&~m[214])|(~m[41]&m[100]&m[214]))&~BiasedRNG[197])|((~m[41]&~m[100]&m[214])|(m[41]&~m[100]&m[214])|(m[41]&m[100]&m[214]));
    m[151] = (((~m[41]&~m[108]&~m[215])|(m[41]&m[108]&~m[215]))&BiasedRNG[198])|(((m[41]&~m[108]&~m[215])|(~m[41]&m[108]&m[215]))&~BiasedRNG[198])|((~m[41]&~m[108]&m[215])|(m[41]&~m[108]&m[215])|(m[41]&m[108]&m[215]));
    m[152] = (((~m[42]&~m[53]&~m[216])|(m[42]&m[53]&~m[216]))&BiasedRNG[199])|(((m[42]&~m[53]&~m[216])|(~m[42]&m[53]&m[216]))&~BiasedRNG[199])|((~m[42]&~m[53]&m[216])|(m[42]&~m[53]&m[216])|(m[42]&m[53]&m[216]));
    m[153] = (((~m[42]&~m[61]&~m[217])|(m[42]&m[61]&~m[217]))&BiasedRNG[200])|(((m[42]&~m[61]&~m[217])|(~m[42]&m[61]&m[217]))&~BiasedRNG[200])|((~m[42]&~m[61]&m[217])|(m[42]&~m[61]&m[217])|(m[42]&m[61]&m[217]));
    m[154] = (((~m[42]&~m[69]&~m[218])|(m[42]&m[69]&~m[218]))&BiasedRNG[201])|(((m[42]&~m[69]&~m[218])|(~m[42]&m[69]&m[218]))&~BiasedRNG[201])|((~m[42]&~m[69]&m[218])|(m[42]&~m[69]&m[218])|(m[42]&m[69]&m[218]));
    m[155] = (((~m[42]&~m[77]&~m[219])|(m[42]&m[77]&~m[219]))&BiasedRNG[202])|(((m[42]&~m[77]&~m[219])|(~m[42]&m[77]&m[219]))&~BiasedRNG[202])|((~m[42]&~m[77]&m[219])|(m[42]&~m[77]&m[219])|(m[42]&m[77]&m[219]));
    m[156] = (((~m[43]&~m[85]&~m[220])|(m[43]&m[85]&~m[220]))&BiasedRNG[203])|(((m[43]&~m[85]&~m[220])|(~m[43]&m[85]&m[220]))&~BiasedRNG[203])|((~m[43]&~m[85]&m[220])|(m[43]&~m[85]&m[220])|(m[43]&m[85]&m[220]));
    m[157] = (((~m[43]&~m[93]&~m[221])|(m[43]&m[93]&~m[221]))&BiasedRNG[204])|(((m[43]&~m[93]&~m[221])|(~m[43]&m[93]&m[221]))&~BiasedRNG[204])|((~m[43]&~m[93]&m[221])|(m[43]&~m[93]&m[221])|(m[43]&m[93]&m[221]));
    m[158] = (((~m[43]&~m[101]&~m[222])|(m[43]&m[101]&~m[222]))&BiasedRNG[205])|(((m[43]&~m[101]&~m[222])|(~m[43]&m[101]&m[222]))&~BiasedRNG[205])|((~m[43]&~m[101]&m[222])|(m[43]&~m[101]&m[222])|(m[43]&m[101]&m[222]));
    m[159] = (((~m[43]&~m[109]&~m[223])|(m[43]&m[109]&~m[223]))&BiasedRNG[206])|(((m[43]&~m[109]&~m[223])|(~m[43]&m[109]&m[223]))&~BiasedRNG[206])|((~m[43]&~m[109]&m[223])|(m[43]&~m[109]&m[223])|(m[43]&m[109]&m[223]));
    m[160] = (((~m[44]&~m[54]&~m[224])|(m[44]&m[54]&~m[224]))&BiasedRNG[207])|(((m[44]&~m[54]&~m[224])|(~m[44]&m[54]&m[224]))&~BiasedRNG[207])|((~m[44]&~m[54]&m[224])|(m[44]&~m[54]&m[224])|(m[44]&m[54]&m[224]));
    m[161] = (((~m[44]&~m[62]&~m[225])|(m[44]&m[62]&~m[225]))&BiasedRNG[208])|(((m[44]&~m[62]&~m[225])|(~m[44]&m[62]&m[225]))&~BiasedRNG[208])|((~m[44]&~m[62]&m[225])|(m[44]&~m[62]&m[225])|(m[44]&m[62]&m[225]));
    m[162] = (((~m[44]&~m[70]&~m[226])|(m[44]&m[70]&~m[226]))&BiasedRNG[209])|(((m[44]&~m[70]&~m[226])|(~m[44]&m[70]&m[226]))&~BiasedRNG[209])|((~m[44]&~m[70]&m[226])|(m[44]&~m[70]&m[226])|(m[44]&m[70]&m[226]));
    m[163] = (((~m[44]&~m[78]&~m[227])|(m[44]&m[78]&~m[227]))&BiasedRNG[210])|(((m[44]&~m[78]&~m[227])|(~m[44]&m[78]&m[227]))&~BiasedRNG[210])|((~m[44]&~m[78]&m[227])|(m[44]&~m[78]&m[227])|(m[44]&m[78]&m[227]));
    m[164] = (((~m[45]&~m[86]&~m[228])|(m[45]&m[86]&~m[228]))&BiasedRNG[211])|(((m[45]&~m[86]&~m[228])|(~m[45]&m[86]&m[228]))&~BiasedRNG[211])|((~m[45]&~m[86]&m[228])|(m[45]&~m[86]&m[228])|(m[45]&m[86]&m[228]));
    m[165] = (((~m[45]&~m[94]&~m[229])|(m[45]&m[94]&~m[229]))&BiasedRNG[212])|(((m[45]&~m[94]&~m[229])|(~m[45]&m[94]&m[229]))&~BiasedRNG[212])|((~m[45]&~m[94]&m[229])|(m[45]&~m[94]&m[229])|(m[45]&m[94]&m[229]));
    m[166] = (((~m[45]&~m[102]&~m[230])|(m[45]&m[102]&~m[230]))&BiasedRNG[213])|(((m[45]&~m[102]&~m[230])|(~m[45]&m[102]&m[230]))&~BiasedRNG[213])|((~m[45]&~m[102]&m[230])|(m[45]&~m[102]&m[230])|(m[45]&m[102]&m[230]));
    m[167] = (((~m[45]&~m[110]&~m[231])|(m[45]&m[110]&~m[231]))&BiasedRNG[214])|(((m[45]&~m[110]&~m[231])|(~m[45]&m[110]&m[231]))&~BiasedRNG[214])|((~m[45]&~m[110]&m[231])|(m[45]&~m[110]&m[231])|(m[45]&m[110]&m[231]));
    m[168] = (((~m[46]&~m[55]&~m[232])|(m[46]&m[55]&~m[232]))&BiasedRNG[215])|(((m[46]&~m[55]&~m[232])|(~m[46]&m[55]&m[232]))&~BiasedRNG[215])|((~m[46]&~m[55]&m[232])|(m[46]&~m[55]&m[232])|(m[46]&m[55]&m[232]));
    m[169] = (((~m[46]&~m[63]&~m[233])|(m[46]&m[63]&~m[233]))&BiasedRNG[216])|(((m[46]&~m[63]&~m[233])|(~m[46]&m[63]&m[233]))&~BiasedRNG[216])|((~m[46]&~m[63]&m[233])|(m[46]&~m[63]&m[233])|(m[46]&m[63]&m[233]));
    m[170] = (((~m[46]&~m[71]&~m[234])|(m[46]&m[71]&~m[234]))&BiasedRNG[217])|(((m[46]&~m[71]&~m[234])|(~m[46]&m[71]&m[234]))&~BiasedRNG[217])|((~m[46]&~m[71]&m[234])|(m[46]&~m[71]&m[234])|(m[46]&m[71]&m[234]));
    m[171] = (((~m[46]&~m[79]&~m[235])|(m[46]&m[79]&~m[235]))&BiasedRNG[218])|(((m[46]&~m[79]&~m[235])|(~m[46]&m[79]&m[235]))&~BiasedRNG[218])|((~m[46]&~m[79]&m[235])|(m[46]&~m[79]&m[235])|(m[46]&m[79]&m[235]));
    m[172] = (((~m[47]&~m[87]&~m[236])|(m[47]&m[87]&~m[236]))&BiasedRNG[219])|(((m[47]&~m[87]&~m[236])|(~m[47]&m[87]&m[236]))&~BiasedRNG[219])|((~m[47]&~m[87]&m[236])|(m[47]&~m[87]&m[236])|(m[47]&m[87]&m[236]));
    m[173] = (((~m[47]&~m[95]&~m[237])|(m[47]&m[95]&~m[237]))&BiasedRNG[220])|(((m[47]&~m[95]&~m[237])|(~m[47]&m[95]&m[237]))&~BiasedRNG[220])|((~m[47]&~m[95]&m[237])|(m[47]&~m[95]&m[237])|(m[47]&m[95]&m[237]));
    m[174] = (((~m[47]&~m[103]&~m[238])|(m[47]&m[103]&~m[238]))&BiasedRNG[221])|(((m[47]&~m[103]&~m[238])|(~m[47]&m[103]&m[238]))&~BiasedRNG[221])|((~m[47]&~m[103]&m[238])|(m[47]&~m[103]&m[238])|(m[47]&m[103]&m[238]));
    m[175] = (((~m[47]&~m[111]&~m[239])|(m[47]&m[111]&~m[239]))&BiasedRNG[222])|(((m[47]&~m[111]&~m[239])|(~m[47]&m[111]&m[239]))&~BiasedRNG[222])|((~m[47]&~m[111]&m[239])|(m[47]&~m[111]&m[239])|(m[47]&m[111]&m[239]));
    m[241] = (((m[184]&~m[240]&~m[242]&~m[243]&~m[244])|(~m[184]&~m[240]&~m[242]&m[243]&~m[244])|(m[184]&m[240]&~m[242]&m[243]&~m[244])|(m[184]&~m[240]&m[242]&m[243]&~m[244])|(~m[184]&m[240]&~m[242]&~m[243]&m[244])|(~m[184]&~m[240]&m[242]&~m[243]&m[244])|(m[184]&m[240]&m[242]&~m[243]&m[244])|(~m[184]&m[240]&m[242]&m[243]&m[244]))&UnbiasedRNG[120])|((m[184]&~m[240]&~m[242]&m[243]&~m[244])|(~m[184]&~m[240]&~m[242]&~m[243]&m[244])|(m[184]&~m[240]&~m[242]&~m[243]&m[244])|(m[184]&m[240]&~m[242]&~m[243]&m[244])|(m[184]&~m[240]&m[242]&~m[243]&m[244])|(~m[184]&~m[240]&~m[242]&m[243]&m[244])|(m[184]&~m[240]&~m[242]&m[243]&m[244])|(~m[184]&m[240]&~m[242]&m[243]&m[244])|(m[184]&m[240]&~m[242]&m[243]&m[244])|(~m[184]&~m[240]&m[242]&m[243]&m[244])|(m[184]&~m[240]&m[242]&m[243]&m[244])|(m[184]&m[240]&m[242]&m[243]&m[244]));
    m[246] = (((m[185]&~m[245]&~m[247]&~m[248]&~m[249])|(~m[185]&~m[245]&~m[247]&m[248]&~m[249])|(m[185]&m[245]&~m[247]&m[248]&~m[249])|(m[185]&~m[245]&m[247]&m[248]&~m[249])|(~m[185]&m[245]&~m[247]&~m[248]&m[249])|(~m[185]&~m[245]&m[247]&~m[248]&m[249])|(m[185]&m[245]&m[247]&~m[248]&m[249])|(~m[185]&m[245]&m[247]&m[248]&m[249]))&UnbiasedRNG[121])|((m[185]&~m[245]&~m[247]&m[248]&~m[249])|(~m[185]&~m[245]&~m[247]&~m[248]&m[249])|(m[185]&~m[245]&~m[247]&~m[248]&m[249])|(m[185]&m[245]&~m[247]&~m[248]&m[249])|(m[185]&~m[245]&m[247]&~m[248]&m[249])|(~m[185]&~m[245]&~m[247]&m[248]&m[249])|(m[185]&~m[245]&~m[247]&m[248]&m[249])|(~m[185]&m[245]&~m[247]&m[248]&m[249])|(m[185]&m[245]&~m[247]&m[248]&m[249])|(~m[185]&~m[245]&m[247]&m[248]&m[249])|(m[185]&~m[245]&m[247]&m[248]&m[249])|(m[185]&m[245]&m[247]&m[248]&m[249]));
    m[251] = (((m[192]&~m[250]&~m[252]&~m[253]&~m[254])|(~m[192]&~m[250]&~m[252]&m[253]&~m[254])|(m[192]&m[250]&~m[252]&m[253]&~m[254])|(m[192]&~m[250]&m[252]&m[253]&~m[254])|(~m[192]&m[250]&~m[252]&~m[253]&m[254])|(~m[192]&~m[250]&m[252]&~m[253]&m[254])|(m[192]&m[250]&m[252]&~m[253]&m[254])|(~m[192]&m[250]&m[252]&m[253]&m[254]))&UnbiasedRNG[122])|((m[192]&~m[250]&~m[252]&m[253]&~m[254])|(~m[192]&~m[250]&~m[252]&~m[253]&m[254])|(m[192]&~m[250]&~m[252]&~m[253]&m[254])|(m[192]&m[250]&~m[252]&~m[253]&m[254])|(m[192]&~m[250]&m[252]&~m[253]&m[254])|(~m[192]&~m[250]&~m[252]&m[253]&m[254])|(m[192]&~m[250]&~m[252]&m[253]&m[254])|(~m[192]&m[250]&~m[252]&m[253]&m[254])|(m[192]&m[250]&~m[252]&m[253]&m[254])|(~m[192]&~m[250]&m[252]&m[253]&m[254])|(m[192]&~m[250]&m[252]&m[253]&m[254])|(m[192]&m[250]&m[252]&m[253]&m[254]));
    m[256] = (((m[186]&~m[255]&~m[257]&~m[258]&~m[259])|(~m[186]&~m[255]&~m[257]&m[258]&~m[259])|(m[186]&m[255]&~m[257]&m[258]&~m[259])|(m[186]&~m[255]&m[257]&m[258]&~m[259])|(~m[186]&m[255]&~m[257]&~m[258]&m[259])|(~m[186]&~m[255]&m[257]&~m[258]&m[259])|(m[186]&m[255]&m[257]&~m[258]&m[259])|(~m[186]&m[255]&m[257]&m[258]&m[259]))&UnbiasedRNG[123])|((m[186]&~m[255]&~m[257]&m[258]&~m[259])|(~m[186]&~m[255]&~m[257]&~m[258]&m[259])|(m[186]&~m[255]&~m[257]&~m[258]&m[259])|(m[186]&m[255]&~m[257]&~m[258]&m[259])|(m[186]&~m[255]&m[257]&~m[258]&m[259])|(~m[186]&~m[255]&~m[257]&m[258]&m[259])|(m[186]&~m[255]&~m[257]&m[258]&m[259])|(~m[186]&m[255]&~m[257]&m[258]&m[259])|(m[186]&m[255]&~m[257]&m[258]&m[259])|(~m[186]&~m[255]&m[257]&m[258]&m[259])|(m[186]&~m[255]&m[257]&m[258]&m[259])|(m[186]&m[255]&m[257]&m[258]&m[259]));
    m[261] = (((m[193]&~m[260]&~m[262]&~m[263]&~m[264])|(~m[193]&~m[260]&~m[262]&m[263]&~m[264])|(m[193]&m[260]&~m[262]&m[263]&~m[264])|(m[193]&~m[260]&m[262]&m[263]&~m[264])|(~m[193]&m[260]&~m[262]&~m[263]&m[264])|(~m[193]&~m[260]&m[262]&~m[263]&m[264])|(m[193]&m[260]&m[262]&~m[263]&m[264])|(~m[193]&m[260]&m[262]&m[263]&m[264]))&UnbiasedRNG[124])|((m[193]&~m[260]&~m[262]&m[263]&~m[264])|(~m[193]&~m[260]&~m[262]&~m[263]&m[264])|(m[193]&~m[260]&~m[262]&~m[263]&m[264])|(m[193]&m[260]&~m[262]&~m[263]&m[264])|(m[193]&~m[260]&m[262]&~m[263]&m[264])|(~m[193]&~m[260]&~m[262]&m[263]&m[264])|(m[193]&~m[260]&~m[262]&m[263]&m[264])|(~m[193]&m[260]&~m[262]&m[263]&m[264])|(m[193]&m[260]&~m[262]&m[263]&m[264])|(~m[193]&~m[260]&m[262]&m[263]&m[264])|(m[193]&~m[260]&m[262]&m[263]&m[264])|(m[193]&m[260]&m[262]&m[263]&m[264]));
    m[266] = (((m[200]&~m[265]&~m[267]&~m[268]&~m[269])|(~m[200]&~m[265]&~m[267]&m[268]&~m[269])|(m[200]&m[265]&~m[267]&m[268]&~m[269])|(m[200]&~m[265]&m[267]&m[268]&~m[269])|(~m[200]&m[265]&~m[267]&~m[268]&m[269])|(~m[200]&~m[265]&m[267]&~m[268]&m[269])|(m[200]&m[265]&m[267]&~m[268]&m[269])|(~m[200]&m[265]&m[267]&m[268]&m[269]))&UnbiasedRNG[125])|((m[200]&~m[265]&~m[267]&m[268]&~m[269])|(~m[200]&~m[265]&~m[267]&~m[268]&m[269])|(m[200]&~m[265]&~m[267]&~m[268]&m[269])|(m[200]&m[265]&~m[267]&~m[268]&m[269])|(m[200]&~m[265]&m[267]&~m[268]&m[269])|(~m[200]&~m[265]&~m[267]&m[268]&m[269])|(m[200]&~m[265]&~m[267]&m[268]&m[269])|(~m[200]&m[265]&~m[267]&m[268]&m[269])|(m[200]&m[265]&~m[267]&m[268]&m[269])|(~m[200]&~m[265]&m[267]&m[268]&m[269])|(m[200]&~m[265]&m[267]&m[268]&m[269])|(m[200]&m[265]&m[267]&m[268]&m[269]));
    m[271] = (((m[187]&~m[270]&~m[272]&~m[273]&~m[274])|(~m[187]&~m[270]&~m[272]&m[273]&~m[274])|(m[187]&m[270]&~m[272]&m[273]&~m[274])|(m[187]&~m[270]&m[272]&m[273]&~m[274])|(~m[187]&m[270]&~m[272]&~m[273]&m[274])|(~m[187]&~m[270]&m[272]&~m[273]&m[274])|(m[187]&m[270]&m[272]&~m[273]&m[274])|(~m[187]&m[270]&m[272]&m[273]&m[274]))&UnbiasedRNG[126])|((m[187]&~m[270]&~m[272]&m[273]&~m[274])|(~m[187]&~m[270]&~m[272]&~m[273]&m[274])|(m[187]&~m[270]&~m[272]&~m[273]&m[274])|(m[187]&m[270]&~m[272]&~m[273]&m[274])|(m[187]&~m[270]&m[272]&~m[273]&m[274])|(~m[187]&~m[270]&~m[272]&m[273]&m[274])|(m[187]&~m[270]&~m[272]&m[273]&m[274])|(~m[187]&m[270]&~m[272]&m[273]&m[274])|(m[187]&m[270]&~m[272]&m[273]&m[274])|(~m[187]&~m[270]&m[272]&m[273]&m[274])|(m[187]&~m[270]&m[272]&m[273]&m[274])|(m[187]&m[270]&m[272]&m[273]&m[274]));
    m[276] = (((m[194]&~m[275]&~m[277]&~m[278]&~m[279])|(~m[194]&~m[275]&~m[277]&m[278]&~m[279])|(m[194]&m[275]&~m[277]&m[278]&~m[279])|(m[194]&~m[275]&m[277]&m[278]&~m[279])|(~m[194]&m[275]&~m[277]&~m[278]&m[279])|(~m[194]&~m[275]&m[277]&~m[278]&m[279])|(m[194]&m[275]&m[277]&~m[278]&m[279])|(~m[194]&m[275]&m[277]&m[278]&m[279]))&UnbiasedRNG[127])|((m[194]&~m[275]&~m[277]&m[278]&~m[279])|(~m[194]&~m[275]&~m[277]&~m[278]&m[279])|(m[194]&~m[275]&~m[277]&~m[278]&m[279])|(m[194]&m[275]&~m[277]&~m[278]&m[279])|(m[194]&~m[275]&m[277]&~m[278]&m[279])|(~m[194]&~m[275]&~m[277]&m[278]&m[279])|(m[194]&~m[275]&~m[277]&m[278]&m[279])|(~m[194]&m[275]&~m[277]&m[278]&m[279])|(m[194]&m[275]&~m[277]&m[278]&m[279])|(~m[194]&~m[275]&m[277]&m[278]&m[279])|(m[194]&~m[275]&m[277]&m[278]&m[279])|(m[194]&m[275]&m[277]&m[278]&m[279]));
    m[281] = (((m[201]&~m[280]&~m[282]&~m[283]&~m[284])|(~m[201]&~m[280]&~m[282]&m[283]&~m[284])|(m[201]&m[280]&~m[282]&m[283]&~m[284])|(m[201]&~m[280]&m[282]&m[283]&~m[284])|(~m[201]&m[280]&~m[282]&~m[283]&m[284])|(~m[201]&~m[280]&m[282]&~m[283]&m[284])|(m[201]&m[280]&m[282]&~m[283]&m[284])|(~m[201]&m[280]&m[282]&m[283]&m[284]))&UnbiasedRNG[128])|((m[201]&~m[280]&~m[282]&m[283]&~m[284])|(~m[201]&~m[280]&~m[282]&~m[283]&m[284])|(m[201]&~m[280]&~m[282]&~m[283]&m[284])|(m[201]&m[280]&~m[282]&~m[283]&m[284])|(m[201]&~m[280]&m[282]&~m[283]&m[284])|(~m[201]&~m[280]&~m[282]&m[283]&m[284])|(m[201]&~m[280]&~m[282]&m[283]&m[284])|(~m[201]&m[280]&~m[282]&m[283]&m[284])|(m[201]&m[280]&~m[282]&m[283]&m[284])|(~m[201]&~m[280]&m[282]&m[283]&m[284])|(m[201]&~m[280]&m[282]&m[283]&m[284])|(m[201]&m[280]&m[282]&m[283]&m[284]));
    m[286] = (((m[208]&~m[285]&~m[287]&~m[288]&~m[289])|(~m[208]&~m[285]&~m[287]&m[288]&~m[289])|(m[208]&m[285]&~m[287]&m[288]&~m[289])|(m[208]&~m[285]&m[287]&m[288]&~m[289])|(~m[208]&m[285]&~m[287]&~m[288]&m[289])|(~m[208]&~m[285]&m[287]&~m[288]&m[289])|(m[208]&m[285]&m[287]&~m[288]&m[289])|(~m[208]&m[285]&m[287]&m[288]&m[289]))&UnbiasedRNG[129])|((m[208]&~m[285]&~m[287]&m[288]&~m[289])|(~m[208]&~m[285]&~m[287]&~m[288]&m[289])|(m[208]&~m[285]&~m[287]&~m[288]&m[289])|(m[208]&m[285]&~m[287]&~m[288]&m[289])|(m[208]&~m[285]&m[287]&~m[288]&m[289])|(~m[208]&~m[285]&~m[287]&m[288]&m[289])|(m[208]&~m[285]&~m[287]&m[288]&m[289])|(~m[208]&m[285]&~m[287]&m[288]&m[289])|(m[208]&m[285]&~m[287]&m[288]&m[289])|(~m[208]&~m[285]&m[287]&m[288]&m[289])|(m[208]&~m[285]&m[287]&m[288]&m[289])|(m[208]&m[285]&m[287]&m[288]&m[289]));
    m[291] = (((m[188]&~m[290]&~m[292]&~m[293]&~m[294])|(~m[188]&~m[290]&~m[292]&m[293]&~m[294])|(m[188]&m[290]&~m[292]&m[293]&~m[294])|(m[188]&~m[290]&m[292]&m[293]&~m[294])|(~m[188]&m[290]&~m[292]&~m[293]&m[294])|(~m[188]&~m[290]&m[292]&~m[293]&m[294])|(m[188]&m[290]&m[292]&~m[293]&m[294])|(~m[188]&m[290]&m[292]&m[293]&m[294]))&UnbiasedRNG[130])|((m[188]&~m[290]&~m[292]&m[293]&~m[294])|(~m[188]&~m[290]&~m[292]&~m[293]&m[294])|(m[188]&~m[290]&~m[292]&~m[293]&m[294])|(m[188]&m[290]&~m[292]&~m[293]&m[294])|(m[188]&~m[290]&m[292]&~m[293]&m[294])|(~m[188]&~m[290]&~m[292]&m[293]&m[294])|(m[188]&~m[290]&~m[292]&m[293]&m[294])|(~m[188]&m[290]&~m[292]&m[293]&m[294])|(m[188]&m[290]&~m[292]&m[293]&m[294])|(~m[188]&~m[290]&m[292]&m[293]&m[294])|(m[188]&~m[290]&m[292]&m[293]&m[294])|(m[188]&m[290]&m[292]&m[293]&m[294]));
    m[296] = (((m[195]&~m[295]&~m[297]&~m[298]&~m[299])|(~m[195]&~m[295]&~m[297]&m[298]&~m[299])|(m[195]&m[295]&~m[297]&m[298]&~m[299])|(m[195]&~m[295]&m[297]&m[298]&~m[299])|(~m[195]&m[295]&~m[297]&~m[298]&m[299])|(~m[195]&~m[295]&m[297]&~m[298]&m[299])|(m[195]&m[295]&m[297]&~m[298]&m[299])|(~m[195]&m[295]&m[297]&m[298]&m[299]))&UnbiasedRNG[131])|((m[195]&~m[295]&~m[297]&m[298]&~m[299])|(~m[195]&~m[295]&~m[297]&~m[298]&m[299])|(m[195]&~m[295]&~m[297]&~m[298]&m[299])|(m[195]&m[295]&~m[297]&~m[298]&m[299])|(m[195]&~m[295]&m[297]&~m[298]&m[299])|(~m[195]&~m[295]&~m[297]&m[298]&m[299])|(m[195]&~m[295]&~m[297]&m[298]&m[299])|(~m[195]&m[295]&~m[297]&m[298]&m[299])|(m[195]&m[295]&~m[297]&m[298]&m[299])|(~m[195]&~m[295]&m[297]&m[298]&m[299])|(m[195]&~m[295]&m[297]&m[298]&m[299])|(m[195]&m[295]&m[297]&m[298]&m[299]));
    m[301] = (((m[202]&~m[300]&~m[302]&~m[303]&~m[304])|(~m[202]&~m[300]&~m[302]&m[303]&~m[304])|(m[202]&m[300]&~m[302]&m[303]&~m[304])|(m[202]&~m[300]&m[302]&m[303]&~m[304])|(~m[202]&m[300]&~m[302]&~m[303]&m[304])|(~m[202]&~m[300]&m[302]&~m[303]&m[304])|(m[202]&m[300]&m[302]&~m[303]&m[304])|(~m[202]&m[300]&m[302]&m[303]&m[304]))&UnbiasedRNG[132])|((m[202]&~m[300]&~m[302]&m[303]&~m[304])|(~m[202]&~m[300]&~m[302]&~m[303]&m[304])|(m[202]&~m[300]&~m[302]&~m[303]&m[304])|(m[202]&m[300]&~m[302]&~m[303]&m[304])|(m[202]&~m[300]&m[302]&~m[303]&m[304])|(~m[202]&~m[300]&~m[302]&m[303]&m[304])|(m[202]&~m[300]&~m[302]&m[303]&m[304])|(~m[202]&m[300]&~m[302]&m[303]&m[304])|(m[202]&m[300]&~m[302]&m[303]&m[304])|(~m[202]&~m[300]&m[302]&m[303]&m[304])|(m[202]&~m[300]&m[302]&m[303]&m[304])|(m[202]&m[300]&m[302]&m[303]&m[304]));
    m[306] = (((m[209]&~m[305]&~m[307]&~m[308]&~m[309])|(~m[209]&~m[305]&~m[307]&m[308]&~m[309])|(m[209]&m[305]&~m[307]&m[308]&~m[309])|(m[209]&~m[305]&m[307]&m[308]&~m[309])|(~m[209]&m[305]&~m[307]&~m[308]&m[309])|(~m[209]&~m[305]&m[307]&~m[308]&m[309])|(m[209]&m[305]&m[307]&~m[308]&m[309])|(~m[209]&m[305]&m[307]&m[308]&m[309]))&UnbiasedRNG[133])|((m[209]&~m[305]&~m[307]&m[308]&~m[309])|(~m[209]&~m[305]&~m[307]&~m[308]&m[309])|(m[209]&~m[305]&~m[307]&~m[308]&m[309])|(m[209]&m[305]&~m[307]&~m[308]&m[309])|(m[209]&~m[305]&m[307]&~m[308]&m[309])|(~m[209]&~m[305]&~m[307]&m[308]&m[309])|(m[209]&~m[305]&~m[307]&m[308]&m[309])|(~m[209]&m[305]&~m[307]&m[308]&m[309])|(m[209]&m[305]&~m[307]&m[308]&m[309])|(~m[209]&~m[305]&m[307]&m[308]&m[309])|(m[209]&~m[305]&m[307]&m[308]&m[309])|(m[209]&m[305]&m[307]&m[308]&m[309]));
    m[311] = (((m[216]&~m[310]&~m[312]&~m[313]&~m[314])|(~m[216]&~m[310]&~m[312]&m[313]&~m[314])|(m[216]&m[310]&~m[312]&m[313]&~m[314])|(m[216]&~m[310]&m[312]&m[313]&~m[314])|(~m[216]&m[310]&~m[312]&~m[313]&m[314])|(~m[216]&~m[310]&m[312]&~m[313]&m[314])|(m[216]&m[310]&m[312]&~m[313]&m[314])|(~m[216]&m[310]&m[312]&m[313]&m[314]))&UnbiasedRNG[134])|((m[216]&~m[310]&~m[312]&m[313]&~m[314])|(~m[216]&~m[310]&~m[312]&~m[313]&m[314])|(m[216]&~m[310]&~m[312]&~m[313]&m[314])|(m[216]&m[310]&~m[312]&~m[313]&m[314])|(m[216]&~m[310]&m[312]&~m[313]&m[314])|(~m[216]&~m[310]&~m[312]&m[313]&m[314])|(m[216]&~m[310]&~m[312]&m[313]&m[314])|(~m[216]&m[310]&~m[312]&m[313]&m[314])|(m[216]&m[310]&~m[312]&m[313]&m[314])|(~m[216]&~m[310]&m[312]&m[313]&m[314])|(m[216]&~m[310]&m[312]&m[313]&m[314])|(m[216]&m[310]&m[312]&m[313]&m[314]));
    m[316] = (((m[189]&~m[315]&~m[317]&~m[318]&~m[319])|(~m[189]&~m[315]&~m[317]&m[318]&~m[319])|(m[189]&m[315]&~m[317]&m[318]&~m[319])|(m[189]&~m[315]&m[317]&m[318]&~m[319])|(~m[189]&m[315]&~m[317]&~m[318]&m[319])|(~m[189]&~m[315]&m[317]&~m[318]&m[319])|(m[189]&m[315]&m[317]&~m[318]&m[319])|(~m[189]&m[315]&m[317]&m[318]&m[319]))&UnbiasedRNG[135])|((m[189]&~m[315]&~m[317]&m[318]&~m[319])|(~m[189]&~m[315]&~m[317]&~m[318]&m[319])|(m[189]&~m[315]&~m[317]&~m[318]&m[319])|(m[189]&m[315]&~m[317]&~m[318]&m[319])|(m[189]&~m[315]&m[317]&~m[318]&m[319])|(~m[189]&~m[315]&~m[317]&m[318]&m[319])|(m[189]&~m[315]&~m[317]&m[318]&m[319])|(~m[189]&m[315]&~m[317]&m[318]&m[319])|(m[189]&m[315]&~m[317]&m[318]&m[319])|(~m[189]&~m[315]&m[317]&m[318]&m[319])|(m[189]&~m[315]&m[317]&m[318]&m[319])|(m[189]&m[315]&m[317]&m[318]&m[319]));
    m[321] = (((m[196]&~m[320]&~m[322]&~m[323]&~m[324])|(~m[196]&~m[320]&~m[322]&m[323]&~m[324])|(m[196]&m[320]&~m[322]&m[323]&~m[324])|(m[196]&~m[320]&m[322]&m[323]&~m[324])|(~m[196]&m[320]&~m[322]&~m[323]&m[324])|(~m[196]&~m[320]&m[322]&~m[323]&m[324])|(m[196]&m[320]&m[322]&~m[323]&m[324])|(~m[196]&m[320]&m[322]&m[323]&m[324]))&UnbiasedRNG[136])|((m[196]&~m[320]&~m[322]&m[323]&~m[324])|(~m[196]&~m[320]&~m[322]&~m[323]&m[324])|(m[196]&~m[320]&~m[322]&~m[323]&m[324])|(m[196]&m[320]&~m[322]&~m[323]&m[324])|(m[196]&~m[320]&m[322]&~m[323]&m[324])|(~m[196]&~m[320]&~m[322]&m[323]&m[324])|(m[196]&~m[320]&~m[322]&m[323]&m[324])|(~m[196]&m[320]&~m[322]&m[323]&m[324])|(m[196]&m[320]&~m[322]&m[323]&m[324])|(~m[196]&~m[320]&m[322]&m[323]&m[324])|(m[196]&~m[320]&m[322]&m[323]&m[324])|(m[196]&m[320]&m[322]&m[323]&m[324]));
    m[326] = (((m[203]&~m[325]&~m[327]&~m[328]&~m[329])|(~m[203]&~m[325]&~m[327]&m[328]&~m[329])|(m[203]&m[325]&~m[327]&m[328]&~m[329])|(m[203]&~m[325]&m[327]&m[328]&~m[329])|(~m[203]&m[325]&~m[327]&~m[328]&m[329])|(~m[203]&~m[325]&m[327]&~m[328]&m[329])|(m[203]&m[325]&m[327]&~m[328]&m[329])|(~m[203]&m[325]&m[327]&m[328]&m[329]))&UnbiasedRNG[137])|((m[203]&~m[325]&~m[327]&m[328]&~m[329])|(~m[203]&~m[325]&~m[327]&~m[328]&m[329])|(m[203]&~m[325]&~m[327]&~m[328]&m[329])|(m[203]&m[325]&~m[327]&~m[328]&m[329])|(m[203]&~m[325]&m[327]&~m[328]&m[329])|(~m[203]&~m[325]&~m[327]&m[328]&m[329])|(m[203]&~m[325]&~m[327]&m[328]&m[329])|(~m[203]&m[325]&~m[327]&m[328]&m[329])|(m[203]&m[325]&~m[327]&m[328]&m[329])|(~m[203]&~m[325]&m[327]&m[328]&m[329])|(m[203]&~m[325]&m[327]&m[328]&m[329])|(m[203]&m[325]&m[327]&m[328]&m[329]));
    m[331] = (((m[210]&~m[330]&~m[332]&~m[333]&~m[334])|(~m[210]&~m[330]&~m[332]&m[333]&~m[334])|(m[210]&m[330]&~m[332]&m[333]&~m[334])|(m[210]&~m[330]&m[332]&m[333]&~m[334])|(~m[210]&m[330]&~m[332]&~m[333]&m[334])|(~m[210]&~m[330]&m[332]&~m[333]&m[334])|(m[210]&m[330]&m[332]&~m[333]&m[334])|(~m[210]&m[330]&m[332]&m[333]&m[334]))&UnbiasedRNG[138])|((m[210]&~m[330]&~m[332]&m[333]&~m[334])|(~m[210]&~m[330]&~m[332]&~m[333]&m[334])|(m[210]&~m[330]&~m[332]&~m[333]&m[334])|(m[210]&m[330]&~m[332]&~m[333]&m[334])|(m[210]&~m[330]&m[332]&~m[333]&m[334])|(~m[210]&~m[330]&~m[332]&m[333]&m[334])|(m[210]&~m[330]&~m[332]&m[333]&m[334])|(~m[210]&m[330]&~m[332]&m[333]&m[334])|(m[210]&m[330]&~m[332]&m[333]&m[334])|(~m[210]&~m[330]&m[332]&m[333]&m[334])|(m[210]&~m[330]&m[332]&m[333]&m[334])|(m[210]&m[330]&m[332]&m[333]&m[334]));
    m[336] = (((m[217]&~m[335]&~m[337]&~m[338]&~m[339])|(~m[217]&~m[335]&~m[337]&m[338]&~m[339])|(m[217]&m[335]&~m[337]&m[338]&~m[339])|(m[217]&~m[335]&m[337]&m[338]&~m[339])|(~m[217]&m[335]&~m[337]&~m[338]&m[339])|(~m[217]&~m[335]&m[337]&~m[338]&m[339])|(m[217]&m[335]&m[337]&~m[338]&m[339])|(~m[217]&m[335]&m[337]&m[338]&m[339]))&UnbiasedRNG[139])|((m[217]&~m[335]&~m[337]&m[338]&~m[339])|(~m[217]&~m[335]&~m[337]&~m[338]&m[339])|(m[217]&~m[335]&~m[337]&~m[338]&m[339])|(m[217]&m[335]&~m[337]&~m[338]&m[339])|(m[217]&~m[335]&m[337]&~m[338]&m[339])|(~m[217]&~m[335]&~m[337]&m[338]&m[339])|(m[217]&~m[335]&~m[337]&m[338]&m[339])|(~m[217]&m[335]&~m[337]&m[338]&m[339])|(m[217]&m[335]&~m[337]&m[338]&m[339])|(~m[217]&~m[335]&m[337]&m[338]&m[339])|(m[217]&~m[335]&m[337]&m[338]&m[339])|(m[217]&m[335]&m[337]&m[338]&m[339]));
    m[341] = (((m[224]&~m[340]&~m[342]&~m[343]&~m[344])|(~m[224]&~m[340]&~m[342]&m[343]&~m[344])|(m[224]&m[340]&~m[342]&m[343]&~m[344])|(m[224]&~m[340]&m[342]&m[343]&~m[344])|(~m[224]&m[340]&~m[342]&~m[343]&m[344])|(~m[224]&~m[340]&m[342]&~m[343]&m[344])|(m[224]&m[340]&m[342]&~m[343]&m[344])|(~m[224]&m[340]&m[342]&m[343]&m[344]))&UnbiasedRNG[140])|((m[224]&~m[340]&~m[342]&m[343]&~m[344])|(~m[224]&~m[340]&~m[342]&~m[343]&m[344])|(m[224]&~m[340]&~m[342]&~m[343]&m[344])|(m[224]&m[340]&~m[342]&~m[343]&m[344])|(m[224]&~m[340]&m[342]&~m[343]&m[344])|(~m[224]&~m[340]&~m[342]&m[343]&m[344])|(m[224]&~m[340]&~m[342]&m[343]&m[344])|(~m[224]&m[340]&~m[342]&m[343]&m[344])|(m[224]&m[340]&~m[342]&m[343]&m[344])|(~m[224]&~m[340]&m[342]&m[343]&m[344])|(m[224]&~m[340]&m[342]&m[343]&m[344])|(m[224]&m[340]&m[342]&m[343]&m[344]));
    m[346] = (((m[190]&~m[345]&~m[347]&~m[348]&~m[349])|(~m[190]&~m[345]&~m[347]&m[348]&~m[349])|(m[190]&m[345]&~m[347]&m[348]&~m[349])|(m[190]&~m[345]&m[347]&m[348]&~m[349])|(~m[190]&m[345]&~m[347]&~m[348]&m[349])|(~m[190]&~m[345]&m[347]&~m[348]&m[349])|(m[190]&m[345]&m[347]&~m[348]&m[349])|(~m[190]&m[345]&m[347]&m[348]&m[349]))&UnbiasedRNG[141])|((m[190]&~m[345]&~m[347]&m[348]&~m[349])|(~m[190]&~m[345]&~m[347]&~m[348]&m[349])|(m[190]&~m[345]&~m[347]&~m[348]&m[349])|(m[190]&m[345]&~m[347]&~m[348]&m[349])|(m[190]&~m[345]&m[347]&~m[348]&m[349])|(~m[190]&~m[345]&~m[347]&m[348]&m[349])|(m[190]&~m[345]&~m[347]&m[348]&m[349])|(~m[190]&m[345]&~m[347]&m[348]&m[349])|(m[190]&m[345]&~m[347]&m[348]&m[349])|(~m[190]&~m[345]&m[347]&m[348]&m[349])|(m[190]&~m[345]&m[347]&m[348]&m[349])|(m[190]&m[345]&m[347]&m[348]&m[349]));
    m[351] = (((m[197]&~m[350]&~m[352]&~m[353]&~m[354])|(~m[197]&~m[350]&~m[352]&m[353]&~m[354])|(m[197]&m[350]&~m[352]&m[353]&~m[354])|(m[197]&~m[350]&m[352]&m[353]&~m[354])|(~m[197]&m[350]&~m[352]&~m[353]&m[354])|(~m[197]&~m[350]&m[352]&~m[353]&m[354])|(m[197]&m[350]&m[352]&~m[353]&m[354])|(~m[197]&m[350]&m[352]&m[353]&m[354]))&UnbiasedRNG[142])|((m[197]&~m[350]&~m[352]&m[353]&~m[354])|(~m[197]&~m[350]&~m[352]&~m[353]&m[354])|(m[197]&~m[350]&~m[352]&~m[353]&m[354])|(m[197]&m[350]&~m[352]&~m[353]&m[354])|(m[197]&~m[350]&m[352]&~m[353]&m[354])|(~m[197]&~m[350]&~m[352]&m[353]&m[354])|(m[197]&~m[350]&~m[352]&m[353]&m[354])|(~m[197]&m[350]&~m[352]&m[353]&m[354])|(m[197]&m[350]&~m[352]&m[353]&m[354])|(~m[197]&~m[350]&m[352]&m[353]&m[354])|(m[197]&~m[350]&m[352]&m[353]&m[354])|(m[197]&m[350]&m[352]&m[353]&m[354]));
    m[356] = (((m[204]&~m[355]&~m[357]&~m[358]&~m[359])|(~m[204]&~m[355]&~m[357]&m[358]&~m[359])|(m[204]&m[355]&~m[357]&m[358]&~m[359])|(m[204]&~m[355]&m[357]&m[358]&~m[359])|(~m[204]&m[355]&~m[357]&~m[358]&m[359])|(~m[204]&~m[355]&m[357]&~m[358]&m[359])|(m[204]&m[355]&m[357]&~m[358]&m[359])|(~m[204]&m[355]&m[357]&m[358]&m[359]))&UnbiasedRNG[143])|((m[204]&~m[355]&~m[357]&m[358]&~m[359])|(~m[204]&~m[355]&~m[357]&~m[358]&m[359])|(m[204]&~m[355]&~m[357]&~m[358]&m[359])|(m[204]&m[355]&~m[357]&~m[358]&m[359])|(m[204]&~m[355]&m[357]&~m[358]&m[359])|(~m[204]&~m[355]&~m[357]&m[358]&m[359])|(m[204]&~m[355]&~m[357]&m[358]&m[359])|(~m[204]&m[355]&~m[357]&m[358]&m[359])|(m[204]&m[355]&~m[357]&m[358]&m[359])|(~m[204]&~m[355]&m[357]&m[358]&m[359])|(m[204]&~m[355]&m[357]&m[358]&m[359])|(m[204]&m[355]&m[357]&m[358]&m[359]));
    m[361] = (((m[211]&~m[360]&~m[362]&~m[363]&~m[364])|(~m[211]&~m[360]&~m[362]&m[363]&~m[364])|(m[211]&m[360]&~m[362]&m[363]&~m[364])|(m[211]&~m[360]&m[362]&m[363]&~m[364])|(~m[211]&m[360]&~m[362]&~m[363]&m[364])|(~m[211]&~m[360]&m[362]&~m[363]&m[364])|(m[211]&m[360]&m[362]&~m[363]&m[364])|(~m[211]&m[360]&m[362]&m[363]&m[364]))&UnbiasedRNG[144])|((m[211]&~m[360]&~m[362]&m[363]&~m[364])|(~m[211]&~m[360]&~m[362]&~m[363]&m[364])|(m[211]&~m[360]&~m[362]&~m[363]&m[364])|(m[211]&m[360]&~m[362]&~m[363]&m[364])|(m[211]&~m[360]&m[362]&~m[363]&m[364])|(~m[211]&~m[360]&~m[362]&m[363]&m[364])|(m[211]&~m[360]&~m[362]&m[363]&m[364])|(~m[211]&m[360]&~m[362]&m[363]&m[364])|(m[211]&m[360]&~m[362]&m[363]&m[364])|(~m[211]&~m[360]&m[362]&m[363]&m[364])|(m[211]&~m[360]&m[362]&m[363]&m[364])|(m[211]&m[360]&m[362]&m[363]&m[364]));
    m[366] = (((m[218]&~m[365]&~m[367]&~m[368]&~m[369])|(~m[218]&~m[365]&~m[367]&m[368]&~m[369])|(m[218]&m[365]&~m[367]&m[368]&~m[369])|(m[218]&~m[365]&m[367]&m[368]&~m[369])|(~m[218]&m[365]&~m[367]&~m[368]&m[369])|(~m[218]&~m[365]&m[367]&~m[368]&m[369])|(m[218]&m[365]&m[367]&~m[368]&m[369])|(~m[218]&m[365]&m[367]&m[368]&m[369]))&UnbiasedRNG[145])|((m[218]&~m[365]&~m[367]&m[368]&~m[369])|(~m[218]&~m[365]&~m[367]&~m[368]&m[369])|(m[218]&~m[365]&~m[367]&~m[368]&m[369])|(m[218]&m[365]&~m[367]&~m[368]&m[369])|(m[218]&~m[365]&m[367]&~m[368]&m[369])|(~m[218]&~m[365]&~m[367]&m[368]&m[369])|(m[218]&~m[365]&~m[367]&m[368]&m[369])|(~m[218]&m[365]&~m[367]&m[368]&m[369])|(m[218]&m[365]&~m[367]&m[368]&m[369])|(~m[218]&~m[365]&m[367]&m[368]&m[369])|(m[218]&~m[365]&m[367]&m[368]&m[369])|(m[218]&m[365]&m[367]&m[368]&m[369]));
    m[371] = (((m[225]&~m[370]&~m[372]&~m[373]&~m[374])|(~m[225]&~m[370]&~m[372]&m[373]&~m[374])|(m[225]&m[370]&~m[372]&m[373]&~m[374])|(m[225]&~m[370]&m[372]&m[373]&~m[374])|(~m[225]&m[370]&~m[372]&~m[373]&m[374])|(~m[225]&~m[370]&m[372]&~m[373]&m[374])|(m[225]&m[370]&m[372]&~m[373]&m[374])|(~m[225]&m[370]&m[372]&m[373]&m[374]))&UnbiasedRNG[146])|((m[225]&~m[370]&~m[372]&m[373]&~m[374])|(~m[225]&~m[370]&~m[372]&~m[373]&m[374])|(m[225]&~m[370]&~m[372]&~m[373]&m[374])|(m[225]&m[370]&~m[372]&~m[373]&m[374])|(m[225]&~m[370]&m[372]&~m[373]&m[374])|(~m[225]&~m[370]&~m[372]&m[373]&m[374])|(m[225]&~m[370]&~m[372]&m[373]&m[374])|(~m[225]&m[370]&~m[372]&m[373]&m[374])|(m[225]&m[370]&~m[372]&m[373]&m[374])|(~m[225]&~m[370]&m[372]&m[373]&m[374])|(m[225]&~m[370]&m[372]&m[373]&m[374])|(m[225]&m[370]&m[372]&m[373]&m[374]));
    m[376] = (((m[232]&~m[375]&~m[377]&~m[378]&~m[379])|(~m[232]&~m[375]&~m[377]&m[378]&~m[379])|(m[232]&m[375]&~m[377]&m[378]&~m[379])|(m[232]&~m[375]&m[377]&m[378]&~m[379])|(~m[232]&m[375]&~m[377]&~m[378]&m[379])|(~m[232]&~m[375]&m[377]&~m[378]&m[379])|(m[232]&m[375]&m[377]&~m[378]&m[379])|(~m[232]&m[375]&m[377]&m[378]&m[379]))&UnbiasedRNG[147])|((m[232]&~m[375]&~m[377]&m[378]&~m[379])|(~m[232]&~m[375]&~m[377]&~m[378]&m[379])|(m[232]&~m[375]&~m[377]&~m[378]&m[379])|(m[232]&m[375]&~m[377]&~m[378]&m[379])|(m[232]&~m[375]&m[377]&~m[378]&m[379])|(~m[232]&~m[375]&~m[377]&m[378]&m[379])|(m[232]&~m[375]&~m[377]&m[378]&m[379])|(~m[232]&m[375]&~m[377]&m[378]&m[379])|(m[232]&m[375]&~m[377]&m[378]&m[379])|(~m[232]&~m[375]&m[377]&m[378]&m[379])|(m[232]&~m[375]&m[377]&m[378]&m[379])|(m[232]&m[375]&m[377]&m[378]&m[379]));
    m[381] = (((m[191]&~m[380]&~m[382]&~m[383]&~m[384])|(~m[191]&~m[380]&~m[382]&m[383]&~m[384])|(m[191]&m[380]&~m[382]&m[383]&~m[384])|(m[191]&~m[380]&m[382]&m[383]&~m[384])|(~m[191]&m[380]&~m[382]&~m[383]&m[384])|(~m[191]&~m[380]&m[382]&~m[383]&m[384])|(m[191]&m[380]&m[382]&~m[383]&m[384])|(~m[191]&m[380]&m[382]&m[383]&m[384]))&UnbiasedRNG[148])|((m[191]&~m[380]&~m[382]&m[383]&~m[384])|(~m[191]&~m[380]&~m[382]&~m[383]&m[384])|(m[191]&~m[380]&~m[382]&~m[383]&m[384])|(m[191]&m[380]&~m[382]&~m[383]&m[384])|(m[191]&~m[380]&m[382]&~m[383]&m[384])|(~m[191]&~m[380]&~m[382]&m[383]&m[384])|(m[191]&~m[380]&~m[382]&m[383]&m[384])|(~m[191]&m[380]&~m[382]&m[383]&m[384])|(m[191]&m[380]&~m[382]&m[383]&m[384])|(~m[191]&~m[380]&m[382]&m[383]&m[384])|(m[191]&~m[380]&m[382]&m[383]&m[384])|(m[191]&m[380]&m[382]&m[383]&m[384]));
    m[386] = (((m[198]&~m[385]&~m[387]&~m[388]&~m[389])|(~m[198]&~m[385]&~m[387]&m[388]&~m[389])|(m[198]&m[385]&~m[387]&m[388]&~m[389])|(m[198]&~m[385]&m[387]&m[388]&~m[389])|(~m[198]&m[385]&~m[387]&~m[388]&m[389])|(~m[198]&~m[385]&m[387]&~m[388]&m[389])|(m[198]&m[385]&m[387]&~m[388]&m[389])|(~m[198]&m[385]&m[387]&m[388]&m[389]))&UnbiasedRNG[149])|((m[198]&~m[385]&~m[387]&m[388]&~m[389])|(~m[198]&~m[385]&~m[387]&~m[388]&m[389])|(m[198]&~m[385]&~m[387]&~m[388]&m[389])|(m[198]&m[385]&~m[387]&~m[388]&m[389])|(m[198]&~m[385]&m[387]&~m[388]&m[389])|(~m[198]&~m[385]&~m[387]&m[388]&m[389])|(m[198]&~m[385]&~m[387]&m[388]&m[389])|(~m[198]&m[385]&~m[387]&m[388]&m[389])|(m[198]&m[385]&~m[387]&m[388]&m[389])|(~m[198]&~m[385]&m[387]&m[388]&m[389])|(m[198]&~m[385]&m[387]&m[388]&m[389])|(m[198]&m[385]&m[387]&m[388]&m[389]));
    m[391] = (((m[205]&~m[390]&~m[392]&~m[393]&~m[394])|(~m[205]&~m[390]&~m[392]&m[393]&~m[394])|(m[205]&m[390]&~m[392]&m[393]&~m[394])|(m[205]&~m[390]&m[392]&m[393]&~m[394])|(~m[205]&m[390]&~m[392]&~m[393]&m[394])|(~m[205]&~m[390]&m[392]&~m[393]&m[394])|(m[205]&m[390]&m[392]&~m[393]&m[394])|(~m[205]&m[390]&m[392]&m[393]&m[394]))&UnbiasedRNG[150])|((m[205]&~m[390]&~m[392]&m[393]&~m[394])|(~m[205]&~m[390]&~m[392]&~m[393]&m[394])|(m[205]&~m[390]&~m[392]&~m[393]&m[394])|(m[205]&m[390]&~m[392]&~m[393]&m[394])|(m[205]&~m[390]&m[392]&~m[393]&m[394])|(~m[205]&~m[390]&~m[392]&m[393]&m[394])|(m[205]&~m[390]&~m[392]&m[393]&m[394])|(~m[205]&m[390]&~m[392]&m[393]&m[394])|(m[205]&m[390]&~m[392]&m[393]&m[394])|(~m[205]&~m[390]&m[392]&m[393]&m[394])|(m[205]&~m[390]&m[392]&m[393]&m[394])|(m[205]&m[390]&m[392]&m[393]&m[394]));
    m[396] = (((m[212]&~m[395]&~m[397]&~m[398]&~m[399])|(~m[212]&~m[395]&~m[397]&m[398]&~m[399])|(m[212]&m[395]&~m[397]&m[398]&~m[399])|(m[212]&~m[395]&m[397]&m[398]&~m[399])|(~m[212]&m[395]&~m[397]&~m[398]&m[399])|(~m[212]&~m[395]&m[397]&~m[398]&m[399])|(m[212]&m[395]&m[397]&~m[398]&m[399])|(~m[212]&m[395]&m[397]&m[398]&m[399]))&UnbiasedRNG[151])|((m[212]&~m[395]&~m[397]&m[398]&~m[399])|(~m[212]&~m[395]&~m[397]&~m[398]&m[399])|(m[212]&~m[395]&~m[397]&~m[398]&m[399])|(m[212]&m[395]&~m[397]&~m[398]&m[399])|(m[212]&~m[395]&m[397]&~m[398]&m[399])|(~m[212]&~m[395]&~m[397]&m[398]&m[399])|(m[212]&~m[395]&~m[397]&m[398]&m[399])|(~m[212]&m[395]&~m[397]&m[398]&m[399])|(m[212]&m[395]&~m[397]&m[398]&m[399])|(~m[212]&~m[395]&m[397]&m[398]&m[399])|(m[212]&~m[395]&m[397]&m[398]&m[399])|(m[212]&m[395]&m[397]&m[398]&m[399]));
    m[401] = (((m[219]&~m[400]&~m[402]&~m[403]&~m[404])|(~m[219]&~m[400]&~m[402]&m[403]&~m[404])|(m[219]&m[400]&~m[402]&m[403]&~m[404])|(m[219]&~m[400]&m[402]&m[403]&~m[404])|(~m[219]&m[400]&~m[402]&~m[403]&m[404])|(~m[219]&~m[400]&m[402]&~m[403]&m[404])|(m[219]&m[400]&m[402]&~m[403]&m[404])|(~m[219]&m[400]&m[402]&m[403]&m[404]))&UnbiasedRNG[152])|((m[219]&~m[400]&~m[402]&m[403]&~m[404])|(~m[219]&~m[400]&~m[402]&~m[403]&m[404])|(m[219]&~m[400]&~m[402]&~m[403]&m[404])|(m[219]&m[400]&~m[402]&~m[403]&m[404])|(m[219]&~m[400]&m[402]&~m[403]&m[404])|(~m[219]&~m[400]&~m[402]&m[403]&m[404])|(m[219]&~m[400]&~m[402]&m[403]&m[404])|(~m[219]&m[400]&~m[402]&m[403]&m[404])|(m[219]&m[400]&~m[402]&m[403]&m[404])|(~m[219]&~m[400]&m[402]&m[403]&m[404])|(m[219]&~m[400]&m[402]&m[403]&m[404])|(m[219]&m[400]&m[402]&m[403]&m[404]));
    m[406] = (((m[226]&~m[405]&~m[407]&~m[408]&~m[409])|(~m[226]&~m[405]&~m[407]&m[408]&~m[409])|(m[226]&m[405]&~m[407]&m[408]&~m[409])|(m[226]&~m[405]&m[407]&m[408]&~m[409])|(~m[226]&m[405]&~m[407]&~m[408]&m[409])|(~m[226]&~m[405]&m[407]&~m[408]&m[409])|(m[226]&m[405]&m[407]&~m[408]&m[409])|(~m[226]&m[405]&m[407]&m[408]&m[409]))&UnbiasedRNG[153])|((m[226]&~m[405]&~m[407]&m[408]&~m[409])|(~m[226]&~m[405]&~m[407]&~m[408]&m[409])|(m[226]&~m[405]&~m[407]&~m[408]&m[409])|(m[226]&m[405]&~m[407]&~m[408]&m[409])|(m[226]&~m[405]&m[407]&~m[408]&m[409])|(~m[226]&~m[405]&~m[407]&m[408]&m[409])|(m[226]&~m[405]&~m[407]&m[408]&m[409])|(~m[226]&m[405]&~m[407]&m[408]&m[409])|(m[226]&m[405]&~m[407]&m[408]&m[409])|(~m[226]&~m[405]&m[407]&m[408]&m[409])|(m[226]&~m[405]&m[407]&m[408]&m[409])|(m[226]&m[405]&m[407]&m[408]&m[409]));
    m[411] = (((m[233]&~m[410]&~m[412]&~m[413]&~m[414])|(~m[233]&~m[410]&~m[412]&m[413]&~m[414])|(m[233]&m[410]&~m[412]&m[413]&~m[414])|(m[233]&~m[410]&m[412]&m[413]&~m[414])|(~m[233]&m[410]&~m[412]&~m[413]&m[414])|(~m[233]&~m[410]&m[412]&~m[413]&m[414])|(m[233]&m[410]&m[412]&~m[413]&m[414])|(~m[233]&m[410]&m[412]&m[413]&m[414]))&UnbiasedRNG[154])|((m[233]&~m[410]&~m[412]&m[413]&~m[414])|(~m[233]&~m[410]&~m[412]&~m[413]&m[414])|(m[233]&~m[410]&~m[412]&~m[413]&m[414])|(m[233]&m[410]&~m[412]&~m[413]&m[414])|(m[233]&~m[410]&m[412]&~m[413]&m[414])|(~m[233]&~m[410]&~m[412]&m[413]&m[414])|(m[233]&~m[410]&~m[412]&m[413]&m[414])|(~m[233]&m[410]&~m[412]&m[413]&m[414])|(m[233]&m[410]&~m[412]&m[413]&m[414])|(~m[233]&~m[410]&m[412]&m[413]&m[414])|(m[233]&~m[410]&m[412]&m[413]&m[414])|(m[233]&m[410]&m[412]&m[413]&m[414]));
    m[416] = (((m[199]&~m[415]&~m[417]&~m[418]&~m[419])|(~m[199]&~m[415]&~m[417]&m[418]&~m[419])|(m[199]&m[415]&~m[417]&m[418]&~m[419])|(m[199]&~m[415]&m[417]&m[418]&~m[419])|(~m[199]&m[415]&~m[417]&~m[418]&m[419])|(~m[199]&~m[415]&m[417]&~m[418]&m[419])|(m[199]&m[415]&m[417]&~m[418]&m[419])|(~m[199]&m[415]&m[417]&m[418]&m[419]))&UnbiasedRNG[155])|((m[199]&~m[415]&~m[417]&m[418]&~m[419])|(~m[199]&~m[415]&~m[417]&~m[418]&m[419])|(m[199]&~m[415]&~m[417]&~m[418]&m[419])|(m[199]&m[415]&~m[417]&~m[418]&m[419])|(m[199]&~m[415]&m[417]&~m[418]&m[419])|(~m[199]&~m[415]&~m[417]&m[418]&m[419])|(m[199]&~m[415]&~m[417]&m[418]&m[419])|(~m[199]&m[415]&~m[417]&m[418]&m[419])|(m[199]&m[415]&~m[417]&m[418]&m[419])|(~m[199]&~m[415]&m[417]&m[418]&m[419])|(m[199]&~m[415]&m[417]&m[418]&m[419])|(m[199]&m[415]&m[417]&m[418]&m[419]));
    m[421] = (((m[206]&~m[420]&~m[422]&~m[423]&~m[424])|(~m[206]&~m[420]&~m[422]&m[423]&~m[424])|(m[206]&m[420]&~m[422]&m[423]&~m[424])|(m[206]&~m[420]&m[422]&m[423]&~m[424])|(~m[206]&m[420]&~m[422]&~m[423]&m[424])|(~m[206]&~m[420]&m[422]&~m[423]&m[424])|(m[206]&m[420]&m[422]&~m[423]&m[424])|(~m[206]&m[420]&m[422]&m[423]&m[424]))&UnbiasedRNG[156])|((m[206]&~m[420]&~m[422]&m[423]&~m[424])|(~m[206]&~m[420]&~m[422]&~m[423]&m[424])|(m[206]&~m[420]&~m[422]&~m[423]&m[424])|(m[206]&m[420]&~m[422]&~m[423]&m[424])|(m[206]&~m[420]&m[422]&~m[423]&m[424])|(~m[206]&~m[420]&~m[422]&m[423]&m[424])|(m[206]&~m[420]&~m[422]&m[423]&m[424])|(~m[206]&m[420]&~m[422]&m[423]&m[424])|(m[206]&m[420]&~m[422]&m[423]&m[424])|(~m[206]&~m[420]&m[422]&m[423]&m[424])|(m[206]&~m[420]&m[422]&m[423]&m[424])|(m[206]&m[420]&m[422]&m[423]&m[424]));
    m[426] = (((m[213]&~m[425]&~m[427]&~m[428]&~m[429])|(~m[213]&~m[425]&~m[427]&m[428]&~m[429])|(m[213]&m[425]&~m[427]&m[428]&~m[429])|(m[213]&~m[425]&m[427]&m[428]&~m[429])|(~m[213]&m[425]&~m[427]&~m[428]&m[429])|(~m[213]&~m[425]&m[427]&~m[428]&m[429])|(m[213]&m[425]&m[427]&~m[428]&m[429])|(~m[213]&m[425]&m[427]&m[428]&m[429]))&UnbiasedRNG[157])|((m[213]&~m[425]&~m[427]&m[428]&~m[429])|(~m[213]&~m[425]&~m[427]&~m[428]&m[429])|(m[213]&~m[425]&~m[427]&~m[428]&m[429])|(m[213]&m[425]&~m[427]&~m[428]&m[429])|(m[213]&~m[425]&m[427]&~m[428]&m[429])|(~m[213]&~m[425]&~m[427]&m[428]&m[429])|(m[213]&~m[425]&~m[427]&m[428]&m[429])|(~m[213]&m[425]&~m[427]&m[428]&m[429])|(m[213]&m[425]&~m[427]&m[428]&m[429])|(~m[213]&~m[425]&m[427]&m[428]&m[429])|(m[213]&~m[425]&m[427]&m[428]&m[429])|(m[213]&m[425]&m[427]&m[428]&m[429]));
    m[431] = (((m[220]&~m[430]&~m[432]&~m[433]&~m[434])|(~m[220]&~m[430]&~m[432]&m[433]&~m[434])|(m[220]&m[430]&~m[432]&m[433]&~m[434])|(m[220]&~m[430]&m[432]&m[433]&~m[434])|(~m[220]&m[430]&~m[432]&~m[433]&m[434])|(~m[220]&~m[430]&m[432]&~m[433]&m[434])|(m[220]&m[430]&m[432]&~m[433]&m[434])|(~m[220]&m[430]&m[432]&m[433]&m[434]))&UnbiasedRNG[158])|((m[220]&~m[430]&~m[432]&m[433]&~m[434])|(~m[220]&~m[430]&~m[432]&~m[433]&m[434])|(m[220]&~m[430]&~m[432]&~m[433]&m[434])|(m[220]&m[430]&~m[432]&~m[433]&m[434])|(m[220]&~m[430]&m[432]&~m[433]&m[434])|(~m[220]&~m[430]&~m[432]&m[433]&m[434])|(m[220]&~m[430]&~m[432]&m[433]&m[434])|(~m[220]&m[430]&~m[432]&m[433]&m[434])|(m[220]&m[430]&~m[432]&m[433]&m[434])|(~m[220]&~m[430]&m[432]&m[433]&m[434])|(m[220]&~m[430]&m[432]&m[433]&m[434])|(m[220]&m[430]&m[432]&m[433]&m[434]));
    m[436] = (((m[227]&~m[435]&~m[437]&~m[438]&~m[439])|(~m[227]&~m[435]&~m[437]&m[438]&~m[439])|(m[227]&m[435]&~m[437]&m[438]&~m[439])|(m[227]&~m[435]&m[437]&m[438]&~m[439])|(~m[227]&m[435]&~m[437]&~m[438]&m[439])|(~m[227]&~m[435]&m[437]&~m[438]&m[439])|(m[227]&m[435]&m[437]&~m[438]&m[439])|(~m[227]&m[435]&m[437]&m[438]&m[439]))&UnbiasedRNG[159])|((m[227]&~m[435]&~m[437]&m[438]&~m[439])|(~m[227]&~m[435]&~m[437]&~m[438]&m[439])|(m[227]&~m[435]&~m[437]&~m[438]&m[439])|(m[227]&m[435]&~m[437]&~m[438]&m[439])|(m[227]&~m[435]&m[437]&~m[438]&m[439])|(~m[227]&~m[435]&~m[437]&m[438]&m[439])|(m[227]&~m[435]&~m[437]&m[438]&m[439])|(~m[227]&m[435]&~m[437]&m[438]&m[439])|(m[227]&m[435]&~m[437]&m[438]&m[439])|(~m[227]&~m[435]&m[437]&m[438]&m[439])|(m[227]&~m[435]&m[437]&m[438]&m[439])|(m[227]&m[435]&m[437]&m[438]&m[439]));
    m[441] = (((m[234]&~m[440]&~m[442]&~m[443]&~m[444])|(~m[234]&~m[440]&~m[442]&m[443]&~m[444])|(m[234]&m[440]&~m[442]&m[443]&~m[444])|(m[234]&~m[440]&m[442]&m[443]&~m[444])|(~m[234]&m[440]&~m[442]&~m[443]&m[444])|(~m[234]&~m[440]&m[442]&~m[443]&m[444])|(m[234]&m[440]&m[442]&~m[443]&m[444])|(~m[234]&m[440]&m[442]&m[443]&m[444]))&UnbiasedRNG[160])|((m[234]&~m[440]&~m[442]&m[443]&~m[444])|(~m[234]&~m[440]&~m[442]&~m[443]&m[444])|(m[234]&~m[440]&~m[442]&~m[443]&m[444])|(m[234]&m[440]&~m[442]&~m[443]&m[444])|(m[234]&~m[440]&m[442]&~m[443]&m[444])|(~m[234]&~m[440]&~m[442]&m[443]&m[444])|(m[234]&~m[440]&~m[442]&m[443]&m[444])|(~m[234]&m[440]&~m[442]&m[443]&m[444])|(m[234]&m[440]&~m[442]&m[443]&m[444])|(~m[234]&~m[440]&m[442]&m[443]&m[444])|(m[234]&~m[440]&m[442]&m[443]&m[444])|(m[234]&m[440]&m[442]&m[443]&m[444]));
    m[446] = (((m[207]&~m[445]&~m[447]&~m[448]&~m[449])|(~m[207]&~m[445]&~m[447]&m[448]&~m[449])|(m[207]&m[445]&~m[447]&m[448]&~m[449])|(m[207]&~m[445]&m[447]&m[448]&~m[449])|(~m[207]&m[445]&~m[447]&~m[448]&m[449])|(~m[207]&~m[445]&m[447]&~m[448]&m[449])|(m[207]&m[445]&m[447]&~m[448]&m[449])|(~m[207]&m[445]&m[447]&m[448]&m[449]))&UnbiasedRNG[161])|((m[207]&~m[445]&~m[447]&m[448]&~m[449])|(~m[207]&~m[445]&~m[447]&~m[448]&m[449])|(m[207]&~m[445]&~m[447]&~m[448]&m[449])|(m[207]&m[445]&~m[447]&~m[448]&m[449])|(m[207]&~m[445]&m[447]&~m[448]&m[449])|(~m[207]&~m[445]&~m[447]&m[448]&m[449])|(m[207]&~m[445]&~m[447]&m[448]&m[449])|(~m[207]&m[445]&~m[447]&m[448]&m[449])|(m[207]&m[445]&~m[447]&m[448]&m[449])|(~m[207]&~m[445]&m[447]&m[448]&m[449])|(m[207]&~m[445]&m[447]&m[448]&m[449])|(m[207]&m[445]&m[447]&m[448]&m[449]));
    m[451] = (((m[214]&~m[450]&~m[452]&~m[453]&~m[454])|(~m[214]&~m[450]&~m[452]&m[453]&~m[454])|(m[214]&m[450]&~m[452]&m[453]&~m[454])|(m[214]&~m[450]&m[452]&m[453]&~m[454])|(~m[214]&m[450]&~m[452]&~m[453]&m[454])|(~m[214]&~m[450]&m[452]&~m[453]&m[454])|(m[214]&m[450]&m[452]&~m[453]&m[454])|(~m[214]&m[450]&m[452]&m[453]&m[454]))&UnbiasedRNG[162])|((m[214]&~m[450]&~m[452]&m[453]&~m[454])|(~m[214]&~m[450]&~m[452]&~m[453]&m[454])|(m[214]&~m[450]&~m[452]&~m[453]&m[454])|(m[214]&m[450]&~m[452]&~m[453]&m[454])|(m[214]&~m[450]&m[452]&~m[453]&m[454])|(~m[214]&~m[450]&~m[452]&m[453]&m[454])|(m[214]&~m[450]&~m[452]&m[453]&m[454])|(~m[214]&m[450]&~m[452]&m[453]&m[454])|(m[214]&m[450]&~m[452]&m[453]&m[454])|(~m[214]&~m[450]&m[452]&m[453]&m[454])|(m[214]&~m[450]&m[452]&m[453]&m[454])|(m[214]&m[450]&m[452]&m[453]&m[454]));
    m[456] = (((m[221]&~m[455]&~m[457]&~m[458]&~m[459])|(~m[221]&~m[455]&~m[457]&m[458]&~m[459])|(m[221]&m[455]&~m[457]&m[458]&~m[459])|(m[221]&~m[455]&m[457]&m[458]&~m[459])|(~m[221]&m[455]&~m[457]&~m[458]&m[459])|(~m[221]&~m[455]&m[457]&~m[458]&m[459])|(m[221]&m[455]&m[457]&~m[458]&m[459])|(~m[221]&m[455]&m[457]&m[458]&m[459]))&UnbiasedRNG[163])|((m[221]&~m[455]&~m[457]&m[458]&~m[459])|(~m[221]&~m[455]&~m[457]&~m[458]&m[459])|(m[221]&~m[455]&~m[457]&~m[458]&m[459])|(m[221]&m[455]&~m[457]&~m[458]&m[459])|(m[221]&~m[455]&m[457]&~m[458]&m[459])|(~m[221]&~m[455]&~m[457]&m[458]&m[459])|(m[221]&~m[455]&~m[457]&m[458]&m[459])|(~m[221]&m[455]&~m[457]&m[458]&m[459])|(m[221]&m[455]&~m[457]&m[458]&m[459])|(~m[221]&~m[455]&m[457]&m[458]&m[459])|(m[221]&~m[455]&m[457]&m[458]&m[459])|(m[221]&m[455]&m[457]&m[458]&m[459]));
    m[461] = (((m[228]&~m[460]&~m[462]&~m[463]&~m[464])|(~m[228]&~m[460]&~m[462]&m[463]&~m[464])|(m[228]&m[460]&~m[462]&m[463]&~m[464])|(m[228]&~m[460]&m[462]&m[463]&~m[464])|(~m[228]&m[460]&~m[462]&~m[463]&m[464])|(~m[228]&~m[460]&m[462]&~m[463]&m[464])|(m[228]&m[460]&m[462]&~m[463]&m[464])|(~m[228]&m[460]&m[462]&m[463]&m[464]))&UnbiasedRNG[164])|((m[228]&~m[460]&~m[462]&m[463]&~m[464])|(~m[228]&~m[460]&~m[462]&~m[463]&m[464])|(m[228]&~m[460]&~m[462]&~m[463]&m[464])|(m[228]&m[460]&~m[462]&~m[463]&m[464])|(m[228]&~m[460]&m[462]&~m[463]&m[464])|(~m[228]&~m[460]&~m[462]&m[463]&m[464])|(m[228]&~m[460]&~m[462]&m[463]&m[464])|(~m[228]&m[460]&~m[462]&m[463]&m[464])|(m[228]&m[460]&~m[462]&m[463]&m[464])|(~m[228]&~m[460]&m[462]&m[463]&m[464])|(m[228]&~m[460]&m[462]&m[463]&m[464])|(m[228]&m[460]&m[462]&m[463]&m[464]));
    m[466] = (((m[235]&~m[465]&~m[467]&~m[468]&~m[469])|(~m[235]&~m[465]&~m[467]&m[468]&~m[469])|(m[235]&m[465]&~m[467]&m[468]&~m[469])|(m[235]&~m[465]&m[467]&m[468]&~m[469])|(~m[235]&m[465]&~m[467]&~m[468]&m[469])|(~m[235]&~m[465]&m[467]&~m[468]&m[469])|(m[235]&m[465]&m[467]&~m[468]&m[469])|(~m[235]&m[465]&m[467]&m[468]&m[469]))&UnbiasedRNG[165])|((m[235]&~m[465]&~m[467]&m[468]&~m[469])|(~m[235]&~m[465]&~m[467]&~m[468]&m[469])|(m[235]&~m[465]&~m[467]&~m[468]&m[469])|(m[235]&m[465]&~m[467]&~m[468]&m[469])|(m[235]&~m[465]&m[467]&~m[468]&m[469])|(~m[235]&~m[465]&~m[467]&m[468]&m[469])|(m[235]&~m[465]&~m[467]&m[468]&m[469])|(~m[235]&m[465]&~m[467]&m[468]&m[469])|(m[235]&m[465]&~m[467]&m[468]&m[469])|(~m[235]&~m[465]&m[467]&m[468]&m[469])|(m[235]&~m[465]&m[467]&m[468]&m[469])|(m[235]&m[465]&m[467]&m[468]&m[469]));
    m[471] = (((m[215]&~m[470]&~m[472]&~m[473]&~m[474])|(~m[215]&~m[470]&~m[472]&m[473]&~m[474])|(m[215]&m[470]&~m[472]&m[473]&~m[474])|(m[215]&~m[470]&m[472]&m[473]&~m[474])|(~m[215]&m[470]&~m[472]&~m[473]&m[474])|(~m[215]&~m[470]&m[472]&~m[473]&m[474])|(m[215]&m[470]&m[472]&~m[473]&m[474])|(~m[215]&m[470]&m[472]&m[473]&m[474]))&UnbiasedRNG[166])|((m[215]&~m[470]&~m[472]&m[473]&~m[474])|(~m[215]&~m[470]&~m[472]&~m[473]&m[474])|(m[215]&~m[470]&~m[472]&~m[473]&m[474])|(m[215]&m[470]&~m[472]&~m[473]&m[474])|(m[215]&~m[470]&m[472]&~m[473]&m[474])|(~m[215]&~m[470]&~m[472]&m[473]&m[474])|(m[215]&~m[470]&~m[472]&m[473]&m[474])|(~m[215]&m[470]&~m[472]&m[473]&m[474])|(m[215]&m[470]&~m[472]&m[473]&m[474])|(~m[215]&~m[470]&m[472]&m[473]&m[474])|(m[215]&~m[470]&m[472]&m[473]&m[474])|(m[215]&m[470]&m[472]&m[473]&m[474]));
    m[476] = (((m[222]&~m[475]&~m[477]&~m[478]&~m[479])|(~m[222]&~m[475]&~m[477]&m[478]&~m[479])|(m[222]&m[475]&~m[477]&m[478]&~m[479])|(m[222]&~m[475]&m[477]&m[478]&~m[479])|(~m[222]&m[475]&~m[477]&~m[478]&m[479])|(~m[222]&~m[475]&m[477]&~m[478]&m[479])|(m[222]&m[475]&m[477]&~m[478]&m[479])|(~m[222]&m[475]&m[477]&m[478]&m[479]))&UnbiasedRNG[167])|((m[222]&~m[475]&~m[477]&m[478]&~m[479])|(~m[222]&~m[475]&~m[477]&~m[478]&m[479])|(m[222]&~m[475]&~m[477]&~m[478]&m[479])|(m[222]&m[475]&~m[477]&~m[478]&m[479])|(m[222]&~m[475]&m[477]&~m[478]&m[479])|(~m[222]&~m[475]&~m[477]&m[478]&m[479])|(m[222]&~m[475]&~m[477]&m[478]&m[479])|(~m[222]&m[475]&~m[477]&m[478]&m[479])|(m[222]&m[475]&~m[477]&m[478]&m[479])|(~m[222]&~m[475]&m[477]&m[478]&m[479])|(m[222]&~m[475]&m[477]&m[478]&m[479])|(m[222]&m[475]&m[477]&m[478]&m[479]));
    m[481] = (((m[229]&~m[480]&~m[482]&~m[483]&~m[484])|(~m[229]&~m[480]&~m[482]&m[483]&~m[484])|(m[229]&m[480]&~m[482]&m[483]&~m[484])|(m[229]&~m[480]&m[482]&m[483]&~m[484])|(~m[229]&m[480]&~m[482]&~m[483]&m[484])|(~m[229]&~m[480]&m[482]&~m[483]&m[484])|(m[229]&m[480]&m[482]&~m[483]&m[484])|(~m[229]&m[480]&m[482]&m[483]&m[484]))&UnbiasedRNG[168])|((m[229]&~m[480]&~m[482]&m[483]&~m[484])|(~m[229]&~m[480]&~m[482]&~m[483]&m[484])|(m[229]&~m[480]&~m[482]&~m[483]&m[484])|(m[229]&m[480]&~m[482]&~m[483]&m[484])|(m[229]&~m[480]&m[482]&~m[483]&m[484])|(~m[229]&~m[480]&~m[482]&m[483]&m[484])|(m[229]&~m[480]&~m[482]&m[483]&m[484])|(~m[229]&m[480]&~m[482]&m[483]&m[484])|(m[229]&m[480]&~m[482]&m[483]&m[484])|(~m[229]&~m[480]&m[482]&m[483]&m[484])|(m[229]&~m[480]&m[482]&m[483]&m[484])|(m[229]&m[480]&m[482]&m[483]&m[484]));
    m[486] = (((m[236]&~m[485]&~m[487]&~m[488]&~m[489])|(~m[236]&~m[485]&~m[487]&m[488]&~m[489])|(m[236]&m[485]&~m[487]&m[488]&~m[489])|(m[236]&~m[485]&m[487]&m[488]&~m[489])|(~m[236]&m[485]&~m[487]&~m[488]&m[489])|(~m[236]&~m[485]&m[487]&~m[488]&m[489])|(m[236]&m[485]&m[487]&~m[488]&m[489])|(~m[236]&m[485]&m[487]&m[488]&m[489]))&UnbiasedRNG[169])|((m[236]&~m[485]&~m[487]&m[488]&~m[489])|(~m[236]&~m[485]&~m[487]&~m[488]&m[489])|(m[236]&~m[485]&~m[487]&~m[488]&m[489])|(m[236]&m[485]&~m[487]&~m[488]&m[489])|(m[236]&~m[485]&m[487]&~m[488]&m[489])|(~m[236]&~m[485]&~m[487]&m[488]&m[489])|(m[236]&~m[485]&~m[487]&m[488]&m[489])|(~m[236]&m[485]&~m[487]&m[488]&m[489])|(m[236]&m[485]&~m[487]&m[488]&m[489])|(~m[236]&~m[485]&m[487]&m[488]&m[489])|(m[236]&~m[485]&m[487]&m[488]&m[489])|(m[236]&m[485]&m[487]&m[488]&m[489]));
    m[491] = (((m[223]&~m[490]&~m[492]&~m[493]&~m[494])|(~m[223]&~m[490]&~m[492]&m[493]&~m[494])|(m[223]&m[490]&~m[492]&m[493]&~m[494])|(m[223]&~m[490]&m[492]&m[493]&~m[494])|(~m[223]&m[490]&~m[492]&~m[493]&m[494])|(~m[223]&~m[490]&m[492]&~m[493]&m[494])|(m[223]&m[490]&m[492]&~m[493]&m[494])|(~m[223]&m[490]&m[492]&m[493]&m[494]))&UnbiasedRNG[170])|((m[223]&~m[490]&~m[492]&m[493]&~m[494])|(~m[223]&~m[490]&~m[492]&~m[493]&m[494])|(m[223]&~m[490]&~m[492]&~m[493]&m[494])|(m[223]&m[490]&~m[492]&~m[493]&m[494])|(m[223]&~m[490]&m[492]&~m[493]&m[494])|(~m[223]&~m[490]&~m[492]&m[493]&m[494])|(m[223]&~m[490]&~m[492]&m[493]&m[494])|(~m[223]&m[490]&~m[492]&m[493]&m[494])|(m[223]&m[490]&~m[492]&m[493]&m[494])|(~m[223]&~m[490]&m[492]&m[493]&m[494])|(m[223]&~m[490]&m[492]&m[493]&m[494])|(m[223]&m[490]&m[492]&m[493]&m[494]));
    m[496] = (((m[230]&~m[495]&~m[497]&~m[498]&~m[499])|(~m[230]&~m[495]&~m[497]&m[498]&~m[499])|(m[230]&m[495]&~m[497]&m[498]&~m[499])|(m[230]&~m[495]&m[497]&m[498]&~m[499])|(~m[230]&m[495]&~m[497]&~m[498]&m[499])|(~m[230]&~m[495]&m[497]&~m[498]&m[499])|(m[230]&m[495]&m[497]&~m[498]&m[499])|(~m[230]&m[495]&m[497]&m[498]&m[499]))&UnbiasedRNG[171])|((m[230]&~m[495]&~m[497]&m[498]&~m[499])|(~m[230]&~m[495]&~m[497]&~m[498]&m[499])|(m[230]&~m[495]&~m[497]&~m[498]&m[499])|(m[230]&m[495]&~m[497]&~m[498]&m[499])|(m[230]&~m[495]&m[497]&~m[498]&m[499])|(~m[230]&~m[495]&~m[497]&m[498]&m[499])|(m[230]&~m[495]&~m[497]&m[498]&m[499])|(~m[230]&m[495]&~m[497]&m[498]&m[499])|(m[230]&m[495]&~m[497]&m[498]&m[499])|(~m[230]&~m[495]&m[497]&m[498]&m[499])|(m[230]&~m[495]&m[497]&m[498]&m[499])|(m[230]&m[495]&m[497]&m[498]&m[499]));
    m[501] = (((m[237]&~m[500]&~m[502]&~m[503]&~m[504])|(~m[237]&~m[500]&~m[502]&m[503]&~m[504])|(m[237]&m[500]&~m[502]&m[503]&~m[504])|(m[237]&~m[500]&m[502]&m[503]&~m[504])|(~m[237]&m[500]&~m[502]&~m[503]&m[504])|(~m[237]&~m[500]&m[502]&~m[503]&m[504])|(m[237]&m[500]&m[502]&~m[503]&m[504])|(~m[237]&m[500]&m[502]&m[503]&m[504]))&UnbiasedRNG[172])|((m[237]&~m[500]&~m[502]&m[503]&~m[504])|(~m[237]&~m[500]&~m[502]&~m[503]&m[504])|(m[237]&~m[500]&~m[502]&~m[503]&m[504])|(m[237]&m[500]&~m[502]&~m[503]&m[504])|(m[237]&~m[500]&m[502]&~m[503]&m[504])|(~m[237]&~m[500]&~m[502]&m[503]&m[504])|(m[237]&~m[500]&~m[502]&m[503]&m[504])|(~m[237]&m[500]&~m[502]&m[503]&m[504])|(m[237]&m[500]&~m[502]&m[503]&m[504])|(~m[237]&~m[500]&m[502]&m[503]&m[504])|(m[237]&~m[500]&m[502]&m[503]&m[504])|(m[237]&m[500]&m[502]&m[503]&m[504]));
    m[506] = (((m[231]&~m[505]&~m[507]&~m[508]&~m[509])|(~m[231]&~m[505]&~m[507]&m[508]&~m[509])|(m[231]&m[505]&~m[507]&m[508]&~m[509])|(m[231]&~m[505]&m[507]&m[508]&~m[509])|(~m[231]&m[505]&~m[507]&~m[508]&m[509])|(~m[231]&~m[505]&m[507]&~m[508]&m[509])|(m[231]&m[505]&m[507]&~m[508]&m[509])|(~m[231]&m[505]&m[507]&m[508]&m[509]))&UnbiasedRNG[173])|((m[231]&~m[505]&~m[507]&m[508]&~m[509])|(~m[231]&~m[505]&~m[507]&~m[508]&m[509])|(m[231]&~m[505]&~m[507]&~m[508]&m[509])|(m[231]&m[505]&~m[507]&~m[508]&m[509])|(m[231]&~m[505]&m[507]&~m[508]&m[509])|(~m[231]&~m[505]&~m[507]&m[508]&m[509])|(m[231]&~m[505]&~m[507]&m[508]&m[509])|(~m[231]&m[505]&~m[507]&m[508]&m[509])|(m[231]&m[505]&~m[507]&m[508]&m[509])|(~m[231]&~m[505]&m[507]&m[508]&m[509])|(m[231]&~m[505]&m[507]&m[508]&m[509])|(m[231]&m[505]&m[507]&m[508]&m[509]));
    m[511] = (((m[238]&~m[510]&~m[512]&~m[513]&~m[514])|(~m[238]&~m[510]&~m[512]&m[513]&~m[514])|(m[238]&m[510]&~m[512]&m[513]&~m[514])|(m[238]&~m[510]&m[512]&m[513]&~m[514])|(~m[238]&m[510]&~m[512]&~m[513]&m[514])|(~m[238]&~m[510]&m[512]&~m[513]&m[514])|(m[238]&m[510]&m[512]&~m[513]&m[514])|(~m[238]&m[510]&m[512]&m[513]&m[514]))&UnbiasedRNG[174])|((m[238]&~m[510]&~m[512]&m[513]&~m[514])|(~m[238]&~m[510]&~m[512]&~m[513]&m[514])|(m[238]&~m[510]&~m[512]&~m[513]&m[514])|(m[238]&m[510]&~m[512]&~m[513]&m[514])|(m[238]&~m[510]&m[512]&~m[513]&m[514])|(~m[238]&~m[510]&~m[512]&m[513]&m[514])|(m[238]&~m[510]&~m[512]&m[513]&m[514])|(~m[238]&m[510]&~m[512]&m[513]&m[514])|(m[238]&m[510]&~m[512]&m[513]&m[514])|(~m[238]&~m[510]&m[512]&m[513]&m[514])|(m[238]&~m[510]&m[512]&m[513]&m[514])|(m[238]&m[510]&m[512]&m[513]&m[514]));
    m[516] = (((m[239]&~m[515]&~m[517]&~m[518]&~m[519])|(~m[239]&~m[515]&~m[517]&m[518]&~m[519])|(m[239]&m[515]&~m[517]&m[518]&~m[519])|(m[239]&~m[515]&m[517]&m[518]&~m[519])|(~m[239]&m[515]&~m[517]&~m[518]&m[519])|(~m[239]&~m[515]&m[517]&~m[518]&m[519])|(m[239]&m[515]&m[517]&~m[518]&m[519])|(~m[239]&m[515]&m[517]&m[518]&m[519]))&UnbiasedRNG[175])|((m[239]&~m[515]&~m[517]&m[518]&~m[519])|(~m[239]&~m[515]&~m[517]&~m[518]&m[519])|(m[239]&~m[515]&~m[517]&~m[518]&m[519])|(m[239]&m[515]&~m[517]&~m[518]&m[519])|(m[239]&~m[515]&m[517]&~m[518]&m[519])|(~m[239]&~m[515]&~m[517]&m[518]&m[519])|(m[239]&~m[515]&~m[517]&m[518]&m[519])|(~m[239]&m[515]&~m[517]&m[518]&m[519])|(m[239]&m[515]&~m[517]&m[518]&m[519])|(~m[239]&~m[515]&m[517]&m[518]&m[519])|(m[239]&~m[515]&m[517]&m[518]&m[519])|(m[239]&m[515]&m[517]&m[518]&m[519]));
end

always @(posedge color3_clk) begin
    m[248] = (((m[245]&~m[246]&~m[247]&~m[249]&~m[250])|(~m[245]&m[246]&~m[247]&~m[249]&~m[250])|(~m[245]&~m[246]&m[247]&~m[249]&~m[250])|(m[245]&m[246]&m[247]&m[249]&~m[250])|(~m[245]&~m[246]&~m[247]&~m[249]&m[250])|(m[245]&m[246]&~m[247]&m[249]&m[250])|(m[245]&~m[246]&m[247]&m[249]&m[250])|(~m[245]&m[246]&m[247]&m[249]&m[250]))&UnbiasedRNG[176])|((m[245]&m[246]&~m[247]&~m[249]&~m[250])|(m[245]&~m[246]&m[247]&~m[249]&~m[250])|(~m[245]&m[246]&m[247]&~m[249]&~m[250])|(m[245]&m[246]&m[247]&~m[249]&~m[250])|(m[245]&~m[246]&~m[247]&~m[249]&m[250])|(~m[245]&m[246]&~m[247]&~m[249]&m[250])|(m[245]&m[246]&~m[247]&~m[249]&m[250])|(~m[245]&~m[246]&m[247]&~m[249]&m[250])|(m[245]&~m[246]&m[247]&~m[249]&m[250])|(~m[245]&m[246]&m[247]&~m[249]&m[250])|(m[245]&m[246]&m[247]&~m[249]&m[250])|(m[245]&m[246]&m[247]&m[249]&m[250]));
    m[258] = (((m[255]&~m[256]&~m[257]&~m[259]&~m[260])|(~m[255]&m[256]&~m[257]&~m[259]&~m[260])|(~m[255]&~m[256]&m[257]&~m[259]&~m[260])|(m[255]&m[256]&m[257]&m[259]&~m[260])|(~m[255]&~m[256]&~m[257]&~m[259]&m[260])|(m[255]&m[256]&~m[257]&m[259]&m[260])|(m[255]&~m[256]&m[257]&m[259]&m[260])|(~m[255]&m[256]&m[257]&m[259]&m[260]))&UnbiasedRNG[177])|((m[255]&m[256]&~m[257]&~m[259]&~m[260])|(m[255]&~m[256]&m[257]&~m[259]&~m[260])|(~m[255]&m[256]&m[257]&~m[259]&~m[260])|(m[255]&m[256]&m[257]&~m[259]&~m[260])|(m[255]&~m[256]&~m[257]&~m[259]&m[260])|(~m[255]&m[256]&~m[257]&~m[259]&m[260])|(m[255]&m[256]&~m[257]&~m[259]&m[260])|(~m[255]&~m[256]&m[257]&~m[259]&m[260])|(m[255]&~m[256]&m[257]&~m[259]&m[260])|(~m[255]&m[256]&m[257]&~m[259]&m[260])|(m[255]&m[256]&m[257]&~m[259]&m[260])|(m[255]&m[256]&m[257]&m[259]&m[260]));
    m[263] = (((m[260]&~m[261]&~m[262]&~m[264]&~m[265])|(~m[260]&m[261]&~m[262]&~m[264]&~m[265])|(~m[260]&~m[261]&m[262]&~m[264]&~m[265])|(m[260]&m[261]&m[262]&m[264]&~m[265])|(~m[260]&~m[261]&~m[262]&~m[264]&m[265])|(m[260]&m[261]&~m[262]&m[264]&m[265])|(m[260]&~m[261]&m[262]&m[264]&m[265])|(~m[260]&m[261]&m[262]&m[264]&m[265]))&UnbiasedRNG[178])|((m[260]&m[261]&~m[262]&~m[264]&~m[265])|(m[260]&~m[261]&m[262]&~m[264]&~m[265])|(~m[260]&m[261]&m[262]&~m[264]&~m[265])|(m[260]&m[261]&m[262]&~m[264]&~m[265])|(m[260]&~m[261]&~m[262]&~m[264]&m[265])|(~m[260]&m[261]&~m[262]&~m[264]&m[265])|(m[260]&m[261]&~m[262]&~m[264]&m[265])|(~m[260]&~m[261]&m[262]&~m[264]&m[265])|(m[260]&~m[261]&m[262]&~m[264]&m[265])|(~m[260]&m[261]&m[262]&~m[264]&m[265])|(m[260]&m[261]&m[262]&~m[264]&m[265])|(m[260]&m[261]&m[262]&m[264]&m[265]));
    m[273] = (((m[270]&~m[271]&~m[272]&~m[274]&~m[275])|(~m[270]&m[271]&~m[272]&~m[274]&~m[275])|(~m[270]&~m[271]&m[272]&~m[274]&~m[275])|(m[270]&m[271]&m[272]&m[274]&~m[275])|(~m[270]&~m[271]&~m[272]&~m[274]&m[275])|(m[270]&m[271]&~m[272]&m[274]&m[275])|(m[270]&~m[271]&m[272]&m[274]&m[275])|(~m[270]&m[271]&m[272]&m[274]&m[275]))&UnbiasedRNG[179])|((m[270]&m[271]&~m[272]&~m[274]&~m[275])|(m[270]&~m[271]&m[272]&~m[274]&~m[275])|(~m[270]&m[271]&m[272]&~m[274]&~m[275])|(m[270]&m[271]&m[272]&~m[274]&~m[275])|(m[270]&~m[271]&~m[272]&~m[274]&m[275])|(~m[270]&m[271]&~m[272]&~m[274]&m[275])|(m[270]&m[271]&~m[272]&~m[274]&m[275])|(~m[270]&~m[271]&m[272]&~m[274]&m[275])|(m[270]&~m[271]&m[272]&~m[274]&m[275])|(~m[270]&m[271]&m[272]&~m[274]&m[275])|(m[270]&m[271]&m[272]&~m[274]&m[275])|(m[270]&m[271]&m[272]&m[274]&m[275]));
    m[278] = (((m[275]&~m[276]&~m[277]&~m[279]&~m[280])|(~m[275]&m[276]&~m[277]&~m[279]&~m[280])|(~m[275]&~m[276]&m[277]&~m[279]&~m[280])|(m[275]&m[276]&m[277]&m[279]&~m[280])|(~m[275]&~m[276]&~m[277]&~m[279]&m[280])|(m[275]&m[276]&~m[277]&m[279]&m[280])|(m[275]&~m[276]&m[277]&m[279]&m[280])|(~m[275]&m[276]&m[277]&m[279]&m[280]))&UnbiasedRNG[180])|((m[275]&m[276]&~m[277]&~m[279]&~m[280])|(m[275]&~m[276]&m[277]&~m[279]&~m[280])|(~m[275]&m[276]&m[277]&~m[279]&~m[280])|(m[275]&m[276]&m[277]&~m[279]&~m[280])|(m[275]&~m[276]&~m[277]&~m[279]&m[280])|(~m[275]&m[276]&~m[277]&~m[279]&m[280])|(m[275]&m[276]&~m[277]&~m[279]&m[280])|(~m[275]&~m[276]&m[277]&~m[279]&m[280])|(m[275]&~m[276]&m[277]&~m[279]&m[280])|(~m[275]&m[276]&m[277]&~m[279]&m[280])|(m[275]&m[276]&m[277]&~m[279]&m[280])|(m[275]&m[276]&m[277]&m[279]&m[280]));
    m[283] = (((m[280]&~m[281]&~m[282]&~m[284]&~m[285])|(~m[280]&m[281]&~m[282]&~m[284]&~m[285])|(~m[280]&~m[281]&m[282]&~m[284]&~m[285])|(m[280]&m[281]&m[282]&m[284]&~m[285])|(~m[280]&~m[281]&~m[282]&~m[284]&m[285])|(m[280]&m[281]&~m[282]&m[284]&m[285])|(m[280]&~m[281]&m[282]&m[284]&m[285])|(~m[280]&m[281]&m[282]&m[284]&m[285]))&UnbiasedRNG[181])|((m[280]&m[281]&~m[282]&~m[284]&~m[285])|(m[280]&~m[281]&m[282]&~m[284]&~m[285])|(~m[280]&m[281]&m[282]&~m[284]&~m[285])|(m[280]&m[281]&m[282]&~m[284]&~m[285])|(m[280]&~m[281]&~m[282]&~m[284]&m[285])|(~m[280]&m[281]&~m[282]&~m[284]&m[285])|(m[280]&m[281]&~m[282]&~m[284]&m[285])|(~m[280]&~m[281]&m[282]&~m[284]&m[285])|(m[280]&~m[281]&m[282]&~m[284]&m[285])|(~m[280]&m[281]&m[282]&~m[284]&m[285])|(m[280]&m[281]&m[282]&~m[284]&m[285])|(m[280]&m[281]&m[282]&m[284]&m[285]));
    m[293] = (((m[290]&~m[291]&~m[292]&~m[294]&~m[295])|(~m[290]&m[291]&~m[292]&~m[294]&~m[295])|(~m[290]&~m[291]&m[292]&~m[294]&~m[295])|(m[290]&m[291]&m[292]&m[294]&~m[295])|(~m[290]&~m[291]&~m[292]&~m[294]&m[295])|(m[290]&m[291]&~m[292]&m[294]&m[295])|(m[290]&~m[291]&m[292]&m[294]&m[295])|(~m[290]&m[291]&m[292]&m[294]&m[295]))&UnbiasedRNG[182])|((m[290]&m[291]&~m[292]&~m[294]&~m[295])|(m[290]&~m[291]&m[292]&~m[294]&~m[295])|(~m[290]&m[291]&m[292]&~m[294]&~m[295])|(m[290]&m[291]&m[292]&~m[294]&~m[295])|(m[290]&~m[291]&~m[292]&~m[294]&m[295])|(~m[290]&m[291]&~m[292]&~m[294]&m[295])|(m[290]&m[291]&~m[292]&~m[294]&m[295])|(~m[290]&~m[291]&m[292]&~m[294]&m[295])|(m[290]&~m[291]&m[292]&~m[294]&m[295])|(~m[290]&m[291]&m[292]&~m[294]&m[295])|(m[290]&m[291]&m[292]&~m[294]&m[295])|(m[290]&m[291]&m[292]&m[294]&m[295]));
    m[298] = (((m[295]&~m[296]&~m[297]&~m[299]&~m[300])|(~m[295]&m[296]&~m[297]&~m[299]&~m[300])|(~m[295]&~m[296]&m[297]&~m[299]&~m[300])|(m[295]&m[296]&m[297]&m[299]&~m[300])|(~m[295]&~m[296]&~m[297]&~m[299]&m[300])|(m[295]&m[296]&~m[297]&m[299]&m[300])|(m[295]&~m[296]&m[297]&m[299]&m[300])|(~m[295]&m[296]&m[297]&m[299]&m[300]))&UnbiasedRNG[183])|((m[295]&m[296]&~m[297]&~m[299]&~m[300])|(m[295]&~m[296]&m[297]&~m[299]&~m[300])|(~m[295]&m[296]&m[297]&~m[299]&~m[300])|(m[295]&m[296]&m[297]&~m[299]&~m[300])|(m[295]&~m[296]&~m[297]&~m[299]&m[300])|(~m[295]&m[296]&~m[297]&~m[299]&m[300])|(m[295]&m[296]&~m[297]&~m[299]&m[300])|(~m[295]&~m[296]&m[297]&~m[299]&m[300])|(m[295]&~m[296]&m[297]&~m[299]&m[300])|(~m[295]&m[296]&m[297]&~m[299]&m[300])|(m[295]&m[296]&m[297]&~m[299]&m[300])|(m[295]&m[296]&m[297]&m[299]&m[300]));
    m[303] = (((m[300]&~m[301]&~m[302]&~m[304]&~m[305])|(~m[300]&m[301]&~m[302]&~m[304]&~m[305])|(~m[300]&~m[301]&m[302]&~m[304]&~m[305])|(m[300]&m[301]&m[302]&m[304]&~m[305])|(~m[300]&~m[301]&~m[302]&~m[304]&m[305])|(m[300]&m[301]&~m[302]&m[304]&m[305])|(m[300]&~m[301]&m[302]&m[304]&m[305])|(~m[300]&m[301]&m[302]&m[304]&m[305]))&UnbiasedRNG[184])|((m[300]&m[301]&~m[302]&~m[304]&~m[305])|(m[300]&~m[301]&m[302]&~m[304]&~m[305])|(~m[300]&m[301]&m[302]&~m[304]&~m[305])|(m[300]&m[301]&m[302]&~m[304]&~m[305])|(m[300]&~m[301]&~m[302]&~m[304]&m[305])|(~m[300]&m[301]&~m[302]&~m[304]&m[305])|(m[300]&m[301]&~m[302]&~m[304]&m[305])|(~m[300]&~m[301]&m[302]&~m[304]&m[305])|(m[300]&~m[301]&m[302]&~m[304]&m[305])|(~m[300]&m[301]&m[302]&~m[304]&m[305])|(m[300]&m[301]&m[302]&~m[304]&m[305])|(m[300]&m[301]&m[302]&m[304]&m[305]));
    m[308] = (((m[305]&~m[306]&~m[307]&~m[309]&~m[310])|(~m[305]&m[306]&~m[307]&~m[309]&~m[310])|(~m[305]&~m[306]&m[307]&~m[309]&~m[310])|(m[305]&m[306]&m[307]&m[309]&~m[310])|(~m[305]&~m[306]&~m[307]&~m[309]&m[310])|(m[305]&m[306]&~m[307]&m[309]&m[310])|(m[305]&~m[306]&m[307]&m[309]&m[310])|(~m[305]&m[306]&m[307]&m[309]&m[310]))&UnbiasedRNG[185])|((m[305]&m[306]&~m[307]&~m[309]&~m[310])|(m[305]&~m[306]&m[307]&~m[309]&~m[310])|(~m[305]&m[306]&m[307]&~m[309]&~m[310])|(m[305]&m[306]&m[307]&~m[309]&~m[310])|(m[305]&~m[306]&~m[307]&~m[309]&m[310])|(~m[305]&m[306]&~m[307]&~m[309]&m[310])|(m[305]&m[306]&~m[307]&~m[309]&m[310])|(~m[305]&~m[306]&m[307]&~m[309]&m[310])|(m[305]&~m[306]&m[307]&~m[309]&m[310])|(~m[305]&m[306]&m[307]&~m[309]&m[310])|(m[305]&m[306]&m[307]&~m[309]&m[310])|(m[305]&m[306]&m[307]&m[309]&m[310]));
    m[318] = (((m[315]&~m[316]&~m[317]&~m[319]&~m[320])|(~m[315]&m[316]&~m[317]&~m[319]&~m[320])|(~m[315]&~m[316]&m[317]&~m[319]&~m[320])|(m[315]&m[316]&m[317]&m[319]&~m[320])|(~m[315]&~m[316]&~m[317]&~m[319]&m[320])|(m[315]&m[316]&~m[317]&m[319]&m[320])|(m[315]&~m[316]&m[317]&m[319]&m[320])|(~m[315]&m[316]&m[317]&m[319]&m[320]))&UnbiasedRNG[186])|((m[315]&m[316]&~m[317]&~m[319]&~m[320])|(m[315]&~m[316]&m[317]&~m[319]&~m[320])|(~m[315]&m[316]&m[317]&~m[319]&~m[320])|(m[315]&m[316]&m[317]&~m[319]&~m[320])|(m[315]&~m[316]&~m[317]&~m[319]&m[320])|(~m[315]&m[316]&~m[317]&~m[319]&m[320])|(m[315]&m[316]&~m[317]&~m[319]&m[320])|(~m[315]&~m[316]&m[317]&~m[319]&m[320])|(m[315]&~m[316]&m[317]&~m[319]&m[320])|(~m[315]&m[316]&m[317]&~m[319]&m[320])|(m[315]&m[316]&m[317]&~m[319]&m[320])|(m[315]&m[316]&m[317]&m[319]&m[320]));
    m[323] = (((m[320]&~m[321]&~m[322]&~m[324]&~m[325])|(~m[320]&m[321]&~m[322]&~m[324]&~m[325])|(~m[320]&~m[321]&m[322]&~m[324]&~m[325])|(m[320]&m[321]&m[322]&m[324]&~m[325])|(~m[320]&~m[321]&~m[322]&~m[324]&m[325])|(m[320]&m[321]&~m[322]&m[324]&m[325])|(m[320]&~m[321]&m[322]&m[324]&m[325])|(~m[320]&m[321]&m[322]&m[324]&m[325]))&UnbiasedRNG[187])|((m[320]&m[321]&~m[322]&~m[324]&~m[325])|(m[320]&~m[321]&m[322]&~m[324]&~m[325])|(~m[320]&m[321]&m[322]&~m[324]&~m[325])|(m[320]&m[321]&m[322]&~m[324]&~m[325])|(m[320]&~m[321]&~m[322]&~m[324]&m[325])|(~m[320]&m[321]&~m[322]&~m[324]&m[325])|(m[320]&m[321]&~m[322]&~m[324]&m[325])|(~m[320]&~m[321]&m[322]&~m[324]&m[325])|(m[320]&~m[321]&m[322]&~m[324]&m[325])|(~m[320]&m[321]&m[322]&~m[324]&m[325])|(m[320]&m[321]&m[322]&~m[324]&m[325])|(m[320]&m[321]&m[322]&m[324]&m[325]));
    m[328] = (((m[325]&~m[326]&~m[327]&~m[329]&~m[330])|(~m[325]&m[326]&~m[327]&~m[329]&~m[330])|(~m[325]&~m[326]&m[327]&~m[329]&~m[330])|(m[325]&m[326]&m[327]&m[329]&~m[330])|(~m[325]&~m[326]&~m[327]&~m[329]&m[330])|(m[325]&m[326]&~m[327]&m[329]&m[330])|(m[325]&~m[326]&m[327]&m[329]&m[330])|(~m[325]&m[326]&m[327]&m[329]&m[330]))&UnbiasedRNG[188])|((m[325]&m[326]&~m[327]&~m[329]&~m[330])|(m[325]&~m[326]&m[327]&~m[329]&~m[330])|(~m[325]&m[326]&m[327]&~m[329]&~m[330])|(m[325]&m[326]&m[327]&~m[329]&~m[330])|(m[325]&~m[326]&~m[327]&~m[329]&m[330])|(~m[325]&m[326]&~m[327]&~m[329]&m[330])|(m[325]&m[326]&~m[327]&~m[329]&m[330])|(~m[325]&~m[326]&m[327]&~m[329]&m[330])|(m[325]&~m[326]&m[327]&~m[329]&m[330])|(~m[325]&m[326]&m[327]&~m[329]&m[330])|(m[325]&m[326]&m[327]&~m[329]&m[330])|(m[325]&m[326]&m[327]&m[329]&m[330]));
    m[333] = (((m[330]&~m[331]&~m[332]&~m[334]&~m[335])|(~m[330]&m[331]&~m[332]&~m[334]&~m[335])|(~m[330]&~m[331]&m[332]&~m[334]&~m[335])|(m[330]&m[331]&m[332]&m[334]&~m[335])|(~m[330]&~m[331]&~m[332]&~m[334]&m[335])|(m[330]&m[331]&~m[332]&m[334]&m[335])|(m[330]&~m[331]&m[332]&m[334]&m[335])|(~m[330]&m[331]&m[332]&m[334]&m[335]))&UnbiasedRNG[189])|((m[330]&m[331]&~m[332]&~m[334]&~m[335])|(m[330]&~m[331]&m[332]&~m[334]&~m[335])|(~m[330]&m[331]&m[332]&~m[334]&~m[335])|(m[330]&m[331]&m[332]&~m[334]&~m[335])|(m[330]&~m[331]&~m[332]&~m[334]&m[335])|(~m[330]&m[331]&~m[332]&~m[334]&m[335])|(m[330]&m[331]&~m[332]&~m[334]&m[335])|(~m[330]&~m[331]&m[332]&~m[334]&m[335])|(m[330]&~m[331]&m[332]&~m[334]&m[335])|(~m[330]&m[331]&m[332]&~m[334]&m[335])|(m[330]&m[331]&m[332]&~m[334]&m[335])|(m[330]&m[331]&m[332]&m[334]&m[335]));
    m[338] = (((m[335]&~m[336]&~m[337]&~m[339]&~m[340])|(~m[335]&m[336]&~m[337]&~m[339]&~m[340])|(~m[335]&~m[336]&m[337]&~m[339]&~m[340])|(m[335]&m[336]&m[337]&m[339]&~m[340])|(~m[335]&~m[336]&~m[337]&~m[339]&m[340])|(m[335]&m[336]&~m[337]&m[339]&m[340])|(m[335]&~m[336]&m[337]&m[339]&m[340])|(~m[335]&m[336]&m[337]&m[339]&m[340]))&UnbiasedRNG[190])|((m[335]&m[336]&~m[337]&~m[339]&~m[340])|(m[335]&~m[336]&m[337]&~m[339]&~m[340])|(~m[335]&m[336]&m[337]&~m[339]&~m[340])|(m[335]&m[336]&m[337]&~m[339]&~m[340])|(m[335]&~m[336]&~m[337]&~m[339]&m[340])|(~m[335]&m[336]&~m[337]&~m[339]&m[340])|(m[335]&m[336]&~m[337]&~m[339]&m[340])|(~m[335]&~m[336]&m[337]&~m[339]&m[340])|(m[335]&~m[336]&m[337]&~m[339]&m[340])|(~m[335]&m[336]&m[337]&~m[339]&m[340])|(m[335]&m[336]&m[337]&~m[339]&m[340])|(m[335]&m[336]&m[337]&m[339]&m[340]));
    m[348] = (((m[345]&~m[346]&~m[347]&~m[349]&~m[350])|(~m[345]&m[346]&~m[347]&~m[349]&~m[350])|(~m[345]&~m[346]&m[347]&~m[349]&~m[350])|(m[345]&m[346]&m[347]&m[349]&~m[350])|(~m[345]&~m[346]&~m[347]&~m[349]&m[350])|(m[345]&m[346]&~m[347]&m[349]&m[350])|(m[345]&~m[346]&m[347]&m[349]&m[350])|(~m[345]&m[346]&m[347]&m[349]&m[350]))&UnbiasedRNG[191])|((m[345]&m[346]&~m[347]&~m[349]&~m[350])|(m[345]&~m[346]&m[347]&~m[349]&~m[350])|(~m[345]&m[346]&m[347]&~m[349]&~m[350])|(m[345]&m[346]&m[347]&~m[349]&~m[350])|(m[345]&~m[346]&~m[347]&~m[349]&m[350])|(~m[345]&m[346]&~m[347]&~m[349]&m[350])|(m[345]&m[346]&~m[347]&~m[349]&m[350])|(~m[345]&~m[346]&m[347]&~m[349]&m[350])|(m[345]&~m[346]&m[347]&~m[349]&m[350])|(~m[345]&m[346]&m[347]&~m[349]&m[350])|(m[345]&m[346]&m[347]&~m[349]&m[350])|(m[345]&m[346]&m[347]&m[349]&m[350]));
    m[353] = (((m[350]&~m[351]&~m[352]&~m[354]&~m[355])|(~m[350]&m[351]&~m[352]&~m[354]&~m[355])|(~m[350]&~m[351]&m[352]&~m[354]&~m[355])|(m[350]&m[351]&m[352]&m[354]&~m[355])|(~m[350]&~m[351]&~m[352]&~m[354]&m[355])|(m[350]&m[351]&~m[352]&m[354]&m[355])|(m[350]&~m[351]&m[352]&m[354]&m[355])|(~m[350]&m[351]&m[352]&m[354]&m[355]))&UnbiasedRNG[192])|((m[350]&m[351]&~m[352]&~m[354]&~m[355])|(m[350]&~m[351]&m[352]&~m[354]&~m[355])|(~m[350]&m[351]&m[352]&~m[354]&~m[355])|(m[350]&m[351]&m[352]&~m[354]&~m[355])|(m[350]&~m[351]&~m[352]&~m[354]&m[355])|(~m[350]&m[351]&~m[352]&~m[354]&m[355])|(m[350]&m[351]&~m[352]&~m[354]&m[355])|(~m[350]&~m[351]&m[352]&~m[354]&m[355])|(m[350]&~m[351]&m[352]&~m[354]&m[355])|(~m[350]&m[351]&m[352]&~m[354]&m[355])|(m[350]&m[351]&m[352]&~m[354]&m[355])|(m[350]&m[351]&m[352]&m[354]&m[355]));
    m[358] = (((m[355]&~m[356]&~m[357]&~m[359]&~m[360])|(~m[355]&m[356]&~m[357]&~m[359]&~m[360])|(~m[355]&~m[356]&m[357]&~m[359]&~m[360])|(m[355]&m[356]&m[357]&m[359]&~m[360])|(~m[355]&~m[356]&~m[357]&~m[359]&m[360])|(m[355]&m[356]&~m[357]&m[359]&m[360])|(m[355]&~m[356]&m[357]&m[359]&m[360])|(~m[355]&m[356]&m[357]&m[359]&m[360]))&UnbiasedRNG[193])|((m[355]&m[356]&~m[357]&~m[359]&~m[360])|(m[355]&~m[356]&m[357]&~m[359]&~m[360])|(~m[355]&m[356]&m[357]&~m[359]&~m[360])|(m[355]&m[356]&m[357]&~m[359]&~m[360])|(m[355]&~m[356]&~m[357]&~m[359]&m[360])|(~m[355]&m[356]&~m[357]&~m[359]&m[360])|(m[355]&m[356]&~m[357]&~m[359]&m[360])|(~m[355]&~m[356]&m[357]&~m[359]&m[360])|(m[355]&~m[356]&m[357]&~m[359]&m[360])|(~m[355]&m[356]&m[357]&~m[359]&m[360])|(m[355]&m[356]&m[357]&~m[359]&m[360])|(m[355]&m[356]&m[357]&m[359]&m[360]));
    m[363] = (((m[360]&~m[361]&~m[362]&~m[364]&~m[365])|(~m[360]&m[361]&~m[362]&~m[364]&~m[365])|(~m[360]&~m[361]&m[362]&~m[364]&~m[365])|(m[360]&m[361]&m[362]&m[364]&~m[365])|(~m[360]&~m[361]&~m[362]&~m[364]&m[365])|(m[360]&m[361]&~m[362]&m[364]&m[365])|(m[360]&~m[361]&m[362]&m[364]&m[365])|(~m[360]&m[361]&m[362]&m[364]&m[365]))&UnbiasedRNG[194])|((m[360]&m[361]&~m[362]&~m[364]&~m[365])|(m[360]&~m[361]&m[362]&~m[364]&~m[365])|(~m[360]&m[361]&m[362]&~m[364]&~m[365])|(m[360]&m[361]&m[362]&~m[364]&~m[365])|(m[360]&~m[361]&~m[362]&~m[364]&m[365])|(~m[360]&m[361]&~m[362]&~m[364]&m[365])|(m[360]&m[361]&~m[362]&~m[364]&m[365])|(~m[360]&~m[361]&m[362]&~m[364]&m[365])|(m[360]&~m[361]&m[362]&~m[364]&m[365])|(~m[360]&m[361]&m[362]&~m[364]&m[365])|(m[360]&m[361]&m[362]&~m[364]&m[365])|(m[360]&m[361]&m[362]&m[364]&m[365]));
    m[368] = (((m[365]&~m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&m[366]&~m[367]&~m[369]&~m[370])|(~m[365]&~m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&m[369]&~m[370])|(~m[365]&~m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&m[369]&m[370])|(m[365]&~m[366]&m[367]&m[369]&m[370])|(~m[365]&m[366]&m[367]&m[369]&m[370]))&UnbiasedRNG[195])|((m[365]&m[366]&~m[367]&~m[369]&~m[370])|(m[365]&~m[366]&m[367]&~m[369]&~m[370])|(~m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&m[366]&m[367]&~m[369]&~m[370])|(m[365]&~m[366]&~m[367]&~m[369]&m[370])|(~m[365]&m[366]&~m[367]&~m[369]&m[370])|(m[365]&m[366]&~m[367]&~m[369]&m[370])|(~m[365]&~m[366]&m[367]&~m[369]&m[370])|(m[365]&~m[366]&m[367]&~m[369]&m[370])|(~m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&~m[369]&m[370])|(m[365]&m[366]&m[367]&m[369]&m[370]));
    m[373] = (((m[370]&~m[371]&~m[372]&~m[374]&~m[375])|(~m[370]&m[371]&~m[372]&~m[374]&~m[375])|(~m[370]&~m[371]&m[372]&~m[374]&~m[375])|(m[370]&m[371]&m[372]&m[374]&~m[375])|(~m[370]&~m[371]&~m[372]&~m[374]&m[375])|(m[370]&m[371]&~m[372]&m[374]&m[375])|(m[370]&~m[371]&m[372]&m[374]&m[375])|(~m[370]&m[371]&m[372]&m[374]&m[375]))&UnbiasedRNG[196])|((m[370]&m[371]&~m[372]&~m[374]&~m[375])|(m[370]&~m[371]&m[372]&~m[374]&~m[375])|(~m[370]&m[371]&m[372]&~m[374]&~m[375])|(m[370]&m[371]&m[372]&~m[374]&~m[375])|(m[370]&~m[371]&~m[372]&~m[374]&m[375])|(~m[370]&m[371]&~m[372]&~m[374]&m[375])|(m[370]&m[371]&~m[372]&~m[374]&m[375])|(~m[370]&~m[371]&m[372]&~m[374]&m[375])|(m[370]&~m[371]&m[372]&~m[374]&m[375])|(~m[370]&m[371]&m[372]&~m[374]&m[375])|(m[370]&m[371]&m[372]&~m[374]&m[375])|(m[370]&m[371]&m[372]&m[374]&m[375]));
    m[383] = (((m[380]&~m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&m[381]&~m[382]&~m[384]&~m[385])|(~m[380]&~m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&m[384]&~m[385])|(~m[380]&~m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&m[384]&m[385])|(m[380]&~m[381]&m[382]&m[384]&m[385])|(~m[380]&m[381]&m[382]&m[384]&m[385]))&UnbiasedRNG[197])|((m[380]&m[381]&~m[382]&~m[384]&~m[385])|(m[380]&~m[381]&m[382]&~m[384]&~m[385])|(~m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&m[381]&m[382]&~m[384]&~m[385])|(m[380]&~m[381]&~m[382]&~m[384]&m[385])|(~m[380]&m[381]&~m[382]&~m[384]&m[385])|(m[380]&m[381]&~m[382]&~m[384]&m[385])|(~m[380]&~m[381]&m[382]&~m[384]&m[385])|(m[380]&~m[381]&m[382]&~m[384]&m[385])|(~m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&~m[384]&m[385])|(m[380]&m[381]&m[382]&m[384]&m[385]));
    m[388] = (((m[385]&~m[386]&~m[387]&~m[389]&~m[390])|(~m[385]&m[386]&~m[387]&~m[389]&~m[390])|(~m[385]&~m[386]&m[387]&~m[389]&~m[390])|(m[385]&m[386]&m[387]&m[389]&~m[390])|(~m[385]&~m[386]&~m[387]&~m[389]&m[390])|(m[385]&m[386]&~m[387]&m[389]&m[390])|(m[385]&~m[386]&m[387]&m[389]&m[390])|(~m[385]&m[386]&m[387]&m[389]&m[390]))&UnbiasedRNG[198])|((m[385]&m[386]&~m[387]&~m[389]&~m[390])|(m[385]&~m[386]&m[387]&~m[389]&~m[390])|(~m[385]&m[386]&m[387]&~m[389]&~m[390])|(m[385]&m[386]&m[387]&~m[389]&~m[390])|(m[385]&~m[386]&~m[387]&~m[389]&m[390])|(~m[385]&m[386]&~m[387]&~m[389]&m[390])|(m[385]&m[386]&~m[387]&~m[389]&m[390])|(~m[385]&~m[386]&m[387]&~m[389]&m[390])|(m[385]&~m[386]&m[387]&~m[389]&m[390])|(~m[385]&m[386]&m[387]&~m[389]&m[390])|(m[385]&m[386]&m[387]&~m[389]&m[390])|(m[385]&m[386]&m[387]&m[389]&m[390]));
    m[393] = (((m[390]&~m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&m[391]&~m[392]&~m[394]&~m[395])|(~m[390]&~m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&m[394]&~m[395])|(~m[390]&~m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&m[394]&m[395])|(m[390]&~m[391]&m[392]&m[394]&m[395])|(~m[390]&m[391]&m[392]&m[394]&m[395]))&UnbiasedRNG[199])|((m[390]&m[391]&~m[392]&~m[394]&~m[395])|(m[390]&~m[391]&m[392]&~m[394]&~m[395])|(~m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&m[391]&m[392]&~m[394]&~m[395])|(m[390]&~m[391]&~m[392]&~m[394]&m[395])|(~m[390]&m[391]&~m[392]&~m[394]&m[395])|(m[390]&m[391]&~m[392]&~m[394]&m[395])|(~m[390]&~m[391]&m[392]&~m[394]&m[395])|(m[390]&~m[391]&m[392]&~m[394]&m[395])|(~m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&~m[394]&m[395])|(m[390]&m[391]&m[392]&m[394]&m[395]));
    m[398] = (((m[395]&~m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&m[396]&~m[397]&~m[399]&~m[400])|(~m[395]&~m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&m[399]&~m[400])|(~m[395]&~m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&m[399]&m[400])|(m[395]&~m[396]&m[397]&m[399]&m[400])|(~m[395]&m[396]&m[397]&m[399]&m[400]))&UnbiasedRNG[200])|((m[395]&m[396]&~m[397]&~m[399]&~m[400])|(m[395]&~m[396]&m[397]&~m[399]&~m[400])|(~m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&m[396]&m[397]&~m[399]&~m[400])|(m[395]&~m[396]&~m[397]&~m[399]&m[400])|(~m[395]&m[396]&~m[397]&~m[399]&m[400])|(m[395]&m[396]&~m[397]&~m[399]&m[400])|(~m[395]&~m[396]&m[397]&~m[399]&m[400])|(m[395]&~m[396]&m[397]&~m[399]&m[400])|(~m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&~m[399]&m[400])|(m[395]&m[396]&m[397]&m[399]&m[400]));
    m[403] = (((m[400]&~m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&m[401]&~m[402]&~m[404]&~m[405])|(~m[400]&~m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&m[404]&~m[405])|(~m[400]&~m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&m[404]&m[405])|(m[400]&~m[401]&m[402]&m[404]&m[405])|(~m[400]&m[401]&m[402]&m[404]&m[405]))&UnbiasedRNG[201])|((m[400]&m[401]&~m[402]&~m[404]&~m[405])|(m[400]&~m[401]&m[402]&~m[404]&~m[405])|(~m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&m[401]&m[402]&~m[404]&~m[405])|(m[400]&~m[401]&~m[402]&~m[404]&m[405])|(~m[400]&m[401]&~m[402]&~m[404]&m[405])|(m[400]&m[401]&~m[402]&~m[404]&m[405])|(~m[400]&~m[401]&m[402]&~m[404]&m[405])|(m[400]&~m[401]&m[402]&~m[404]&m[405])|(~m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&~m[404]&m[405])|(m[400]&m[401]&m[402]&m[404]&m[405]));
    m[408] = (((m[405]&~m[406]&~m[407]&~m[409]&~m[410])|(~m[405]&m[406]&~m[407]&~m[409]&~m[410])|(~m[405]&~m[406]&m[407]&~m[409]&~m[410])|(m[405]&m[406]&m[407]&m[409]&~m[410])|(~m[405]&~m[406]&~m[407]&~m[409]&m[410])|(m[405]&m[406]&~m[407]&m[409]&m[410])|(m[405]&~m[406]&m[407]&m[409]&m[410])|(~m[405]&m[406]&m[407]&m[409]&m[410]))&UnbiasedRNG[202])|((m[405]&m[406]&~m[407]&~m[409]&~m[410])|(m[405]&~m[406]&m[407]&~m[409]&~m[410])|(~m[405]&m[406]&m[407]&~m[409]&~m[410])|(m[405]&m[406]&m[407]&~m[409]&~m[410])|(m[405]&~m[406]&~m[407]&~m[409]&m[410])|(~m[405]&m[406]&~m[407]&~m[409]&m[410])|(m[405]&m[406]&~m[407]&~m[409]&m[410])|(~m[405]&~m[406]&m[407]&~m[409]&m[410])|(m[405]&~m[406]&m[407]&~m[409]&m[410])|(~m[405]&m[406]&m[407]&~m[409]&m[410])|(m[405]&m[406]&m[407]&~m[409]&m[410])|(m[405]&m[406]&m[407]&m[409]&m[410]));
    m[418] = (((m[415]&~m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&m[416]&~m[417]&~m[419]&~m[420])|(~m[415]&~m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&m[419]&~m[420])|(~m[415]&~m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&m[419]&m[420])|(m[415]&~m[416]&m[417]&m[419]&m[420])|(~m[415]&m[416]&m[417]&m[419]&m[420]))&UnbiasedRNG[203])|((m[415]&m[416]&~m[417]&~m[419]&~m[420])|(m[415]&~m[416]&m[417]&~m[419]&~m[420])|(~m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&m[416]&m[417]&~m[419]&~m[420])|(m[415]&~m[416]&~m[417]&~m[419]&m[420])|(~m[415]&m[416]&~m[417]&~m[419]&m[420])|(m[415]&m[416]&~m[417]&~m[419]&m[420])|(~m[415]&~m[416]&m[417]&~m[419]&m[420])|(m[415]&~m[416]&m[417]&~m[419]&m[420])|(~m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&~m[419]&m[420])|(m[415]&m[416]&m[417]&m[419]&m[420]));
    m[423] = (((m[420]&~m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&m[421]&~m[422]&~m[424]&~m[425])|(~m[420]&~m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&m[424]&~m[425])|(~m[420]&~m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&m[424]&m[425])|(m[420]&~m[421]&m[422]&m[424]&m[425])|(~m[420]&m[421]&m[422]&m[424]&m[425]))&UnbiasedRNG[204])|((m[420]&m[421]&~m[422]&~m[424]&~m[425])|(m[420]&~m[421]&m[422]&~m[424]&~m[425])|(~m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&m[421]&m[422]&~m[424]&~m[425])|(m[420]&~m[421]&~m[422]&~m[424]&m[425])|(~m[420]&m[421]&~m[422]&~m[424]&m[425])|(m[420]&m[421]&~m[422]&~m[424]&m[425])|(~m[420]&~m[421]&m[422]&~m[424]&m[425])|(m[420]&~m[421]&m[422]&~m[424]&m[425])|(~m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&~m[424]&m[425])|(m[420]&m[421]&m[422]&m[424]&m[425]));
    m[428] = (((m[425]&~m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&m[426]&~m[427]&~m[429]&~m[430])|(~m[425]&~m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&m[429]&~m[430])|(~m[425]&~m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&m[429]&m[430])|(m[425]&~m[426]&m[427]&m[429]&m[430])|(~m[425]&m[426]&m[427]&m[429]&m[430]))&UnbiasedRNG[205])|((m[425]&m[426]&~m[427]&~m[429]&~m[430])|(m[425]&~m[426]&m[427]&~m[429]&~m[430])|(~m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&m[426]&m[427]&~m[429]&~m[430])|(m[425]&~m[426]&~m[427]&~m[429]&m[430])|(~m[425]&m[426]&~m[427]&~m[429]&m[430])|(m[425]&m[426]&~m[427]&~m[429]&m[430])|(~m[425]&~m[426]&m[427]&~m[429]&m[430])|(m[425]&~m[426]&m[427]&~m[429]&m[430])|(~m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&~m[429]&m[430])|(m[425]&m[426]&m[427]&m[429]&m[430]));
    m[433] = (((m[430]&~m[431]&~m[432]&~m[434]&~m[435])|(~m[430]&m[431]&~m[432]&~m[434]&~m[435])|(~m[430]&~m[431]&m[432]&~m[434]&~m[435])|(m[430]&m[431]&m[432]&m[434]&~m[435])|(~m[430]&~m[431]&~m[432]&~m[434]&m[435])|(m[430]&m[431]&~m[432]&m[434]&m[435])|(m[430]&~m[431]&m[432]&m[434]&m[435])|(~m[430]&m[431]&m[432]&m[434]&m[435]))&UnbiasedRNG[206])|((m[430]&m[431]&~m[432]&~m[434]&~m[435])|(m[430]&~m[431]&m[432]&~m[434]&~m[435])|(~m[430]&m[431]&m[432]&~m[434]&~m[435])|(m[430]&m[431]&m[432]&~m[434]&~m[435])|(m[430]&~m[431]&~m[432]&~m[434]&m[435])|(~m[430]&m[431]&~m[432]&~m[434]&m[435])|(m[430]&m[431]&~m[432]&~m[434]&m[435])|(~m[430]&~m[431]&m[432]&~m[434]&m[435])|(m[430]&~m[431]&m[432]&~m[434]&m[435])|(~m[430]&m[431]&m[432]&~m[434]&m[435])|(m[430]&m[431]&m[432]&~m[434]&m[435])|(m[430]&m[431]&m[432]&m[434]&m[435]));
    m[438] = (((m[435]&~m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&m[436]&~m[437]&~m[439]&~m[440])|(~m[435]&~m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&m[439]&~m[440])|(~m[435]&~m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&m[439]&m[440])|(m[435]&~m[436]&m[437]&m[439]&m[440])|(~m[435]&m[436]&m[437]&m[439]&m[440]))&UnbiasedRNG[207])|((m[435]&m[436]&~m[437]&~m[439]&~m[440])|(m[435]&~m[436]&m[437]&~m[439]&~m[440])|(~m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&m[436]&m[437]&~m[439]&~m[440])|(m[435]&~m[436]&~m[437]&~m[439]&m[440])|(~m[435]&m[436]&~m[437]&~m[439]&m[440])|(m[435]&m[436]&~m[437]&~m[439]&m[440])|(~m[435]&~m[436]&m[437]&~m[439]&m[440])|(m[435]&~m[436]&m[437]&~m[439]&m[440])|(~m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&~m[439]&m[440])|(m[435]&m[436]&m[437]&m[439]&m[440]));
    m[448] = (((m[445]&~m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&m[446]&~m[447]&~m[449]&~m[450])|(~m[445]&~m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&m[449]&~m[450])|(~m[445]&~m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&m[449]&m[450])|(m[445]&~m[446]&m[447]&m[449]&m[450])|(~m[445]&m[446]&m[447]&m[449]&m[450]))&UnbiasedRNG[208])|((m[445]&m[446]&~m[447]&~m[449]&~m[450])|(m[445]&~m[446]&m[447]&~m[449]&~m[450])|(~m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&m[446]&m[447]&~m[449]&~m[450])|(m[445]&~m[446]&~m[447]&~m[449]&m[450])|(~m[445]&m[446]&~m[447]&~m[449]&m[450])|(m[445]&m[446]&~m[447]&~m[449]&m[450])|(~m[445]&~m[446]&m[447]&~m[449]&m[450])|(m[445]&~m[446]&m[447]&~m[449]&m[450])|(~m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&~m[449]&m[450])|(m[445]&m[446]&m[447]&m[449]&m[450]));
    m[453] = (((m[450]&~m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&m[451]&~m[452]&~m[454]&~m[455])|(~m[450]&~m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&m[454]&~m[455])|(~m[450]&~m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&m[454]&m[455])|(m[450]&~m[451]&m[452]&m[454]&m[455])|(~m[450]&m[451]&m[452]&m[454]&m[455]))&UnbiasedRNG[209])|((m[450]&m[451]&~m[452]&~m[454]&~m[455])|(m[450]&~m[451]&m[452]&~m[454]&~m[455])|(~m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&m[451]&m[452]&~m[454]&~m[455])|(m[450]&~m[451]&~m[452]&~m[454]&m[455])|(~m[450]&m[451]&~m[452]&~m[454]&m[455])|(m[450]&m[451]&~m[452]&~m[454]&m[455])|(~m[450]&~m[451]&m[452]&~m[454]&m[455])|(m[450]&~m[451]&m[452]&~m[454]&m[455])|(~m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&~m[454]&m[455])|(m[450]&m[451]&m[452]&m[454]&m[455]));
    m[458] = (((m[455]&~m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&m[456]&~m[457]&~m[459]&~m[460])|(~m[455]&~m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&m[459]&~m[460])|(~m[455]&~m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&m[459]&m[460])|(m[455]&~m[456]&m[457]&m[459]&m[460])|(~m[455]&m[456]&m[457]&m[459]&m[460]))&UnbiasedRNG[210])|((m[455]&m[456]&~m[457]&~m[459]&~m[460])|(m[455]&~m[456]&m[457]&~m[459]&~m[460])|(~m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&m[456]&m[457]&~m[459]&~m[460])|(m[455]&~m[456]&~m[457]&~m[459]&m[460])|(~m[455]&m[456]&~m[457]&~m[459]&m[460])|(m[455]&m[456]&~m[457]&~m[459]&m[460])|(~m[455]&~m[456]&m[457]&~m[459]&m[460])|(m[455]&~m[456]&m[457]&~m[459]&m[460])|(~m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&~m[459]&m[460])|(m[455]&m[456]&m[457]&m[459]&m[460]));
    m[463] = (((m[460]&~m[461]&~m[462]&~m[464]&~m[465])|(~m[460]&m[461]&~m[462]&~m[464]&~m[465])|(~m[460]&~m[461]&m[462]&~m[464]&~m[465])|(m[460]&m[461]&m[462]&m[464]&~m[465])|(~m[460]&~m[461]&~m[462]&~m[464]&m[465])|(m[460]&m[461]&~m[462]&m[464]&m[465])|(m[460]&~m[461]&m[462]&m[464]&m[465])|(~m[460]&m[461]&m[462]&m[464]&m[465]))&UnbiasedRNG[211])|((m[460]&m[461]&~m[462]&~m[464]&~m[465])|(m[460]&~m[461]&m[462]&~m[464]&~m[465])|(~m[460]&m[461]&m[462]&~m[464]&~m[465])|(m[460]&m[461]&m[462]&~m[464]&~m[465])|(m[460]&~m[461]&~m[462]&~m[464]&m[465])|(~m[460]&m[461]&~m[462]&~m[464]&m[465])|(m[460]&m[461]&~m[462]&~m[464]&m[465])|(~m[460]&~m[461]&m[462]&~m[464]&m[465])|(m[460]&~m[461]&m[462]&~m[464]&m[465])|(~m[460]&m[461]&m[462]&~m[464]&m[465])|(m[460]&m[461]&m[462]&~m[464]&m[465])|(m[460]&m[461]&m[462]&m[464]&m[465]));
    m[473] = (((m[470]&~m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&m[471]&~m[472]&~m[474]&~m[475])|(~m[470]&~m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&m[474]&~m[475])|(~m[470]&~m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&m[474]&m[475])|(m[470]&~m[471]&m[472]&m[474]&m[475])|(~m[470]&m[471]&m[472]&m[474]&m[475]))&UnbiasedRNG[212])|((m[470]&m[471]&~m[472]&~m[474]&~m[475])|(m[470]&~m[471]&m[472]&~m[474]&~m[475])|(~m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&m[471]&m[472]&~m[474]&~m[475])|(m[470]&~m[471]&~m[472]&~m[474]&m[475])|(~m[470]&m[471]&~m[472]&~m[474]&m[475])|(m[470]&m[471]&~m[472]&~m[474]&m[475])|(~m[470]&~m[471]&m[472]&~m[474]&m[475])|(m[470]&~m[471]&m[472]&~m[474]&m[475])|(~m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&~m[474]&m[475])|(m[470]&m[471]&m[472]&m[474]&m[475]));
    m[478] = (((m[475]&~m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&m[476]&~m[477]&~m[479]&~m[480])|(~m[475]&~m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&m[479]&~m[480])|(~m[475]&~m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&m[479]&m[480])|(m[475]&~m[476]&m[477]&m[479]&m[480])|(~m[475]&m[476]&m[477]&m[479]&m[480]))&UnbiasedRNG[213])|((m[475]&m[476]&~m[477]&~m[479]&~m[480])|(m[475]&~m[476]&m[477]&~m[479]&~m[480])|(~m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&m[476]&m[477]&~m[479]&~m[480])|(m[475]&~m[476]&~m[477]&~m[479]&m[480])|(~m[475]&m[476]&~m[477]&~m[479]&m[480])|(m[475]&m[476]&~m[477]&~m[479]&m[480])|(~m[475]&~m[476]&m[477]&~m[479]&m[480])|(m[475]&~m[476]&m[477]&~m[479]&m[480])|(~m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&~m[479]&m[480])|(m[475]&m[476]&m[477]&m[479]&m[480]));
    m[483] = (((m[480]&~m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&m[481]&~m[482]&~m[484]&~m[485])|(~m[480]&~m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&m[484]&~m[485])|(~m[480]&~m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&m[484]&m[485])|(m[480]&~m[481]&m[482]&m[484]&m[485])|(~m[480]&m[481]&m[482]&m[484]&m[485]))&UnbiasedRNG[214])|((m[480]&m[481]&~m[482]&~m[484]&~m[485])|(m[480]&~m[481]&m[482]&~m[484]&~m[485])|(~m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&m[481]&m[482]&~m[484]&~m[485])|(m[480]&~m[481]&~m[482]&~m[484]&m[485])|(~m[480]&m[481]&~m[482]&~m[484]&m[485])|(m[480]&m[481]&~m[482]&~m[484]&m[485])|(~m[480]&~m[481]&m[482]&~m[484]&m[485])|(m[480]&~m[481]&m[482]&~m[484]&m[485])|(~m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&~m[484]&m[485])|(m[480]&m[481]&m[482]&m[484]&m[485]));
    m[493] = (((m[490]&~m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&m[491]&~m[492]&~m[494]&~m[495])|(~m[490]&~m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&m[494]&~m[495])|(~m[490]&~m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&m[494]&m[495])|(m[490]&~m[491]&m[492]&m[494]&m[495])|(~m[490]&m[491]&m[492]&m[494]&m[495]))&UnbiasedRNG[215])|((m[490]&m[491]&~m[492]&~m[494]&~m[495])|(m[490]&~m[491]&m[492]&~m[494]&~m[495])|(~m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&m[491]&m[492]&~m[494]&~m[495])|(m[490]&~m[491]&~m[492]&~m[494]&m[495])|(~m[490]&m[491]&~m[492]&~m[494]&m[495])|(m[490]&m[491]&~m[492]&~m[494]&m[495])|(~m[490]&~m[491]&m[492]&~m[494]&m[495])|(m[490]&~m[491]&m[492]&~m[494]&m[495])|(~m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&~m[494]&m[495])|(m[490]&m[491]&m[492]&m[494]&m[495]));
    m[498] = (((m[495]&~m[496]&~m[497]&~m[499]&~m[500])|(~m[495]&m[496]&~m[497]&~m[499]&~m[500])|(~m[495]&~m[496]&m[497]&~m[499]&~m[500])|(m[495]&m[496]&m[497]&m[499]&~m[500])|(~m[495]&~m[496]&~m[497]&~m[499]&m[500])|(m[495]&m[496]&~m[497]&m[499]&m[500])|(m[495]&~m[496]&m[497]&m[499]&m[500])|(~m[495]&m[496]&m[497]&m[499]&m[500]))&UnbiasedRNG[216])|((m[495]&m[496]&~m[497]&~m[499]&~m[500])|(m[495]&~m[496]&m[497]&~m[499]&~m[500])|(~m[495]&m[496]&m[497]&~m[499]&~m[500])|(m[495]&m[496]&m[497]&~m[499]&~m[500])|(m[495]&~m[496]&~m[497]&~m[499]&m[500])|(~m[495]&m[496]&~m[497]&~m[499]&m[500])|(m[495]&m[496]&~m[497]&~m[499]&m[500])|(~m[495]&~m[496]&m[497]&~m[499]&m[500])|(m[495]&~m[496]&m[497]&~m[499]&m[500])|(~m[495]&m[496]&m[497]&~m[499]&m[500])|(m[495]&m[496]&m[497]&~m[499]&m[500])|(m[495]&m[496]&m[497]&m[499]&m[500]));
    m[508] = (((m[505]&~m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&m[506]&~m[507]&~m[509]&~m[510])|(~m[505]&~m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&m[509]&~m[510])|(~m[505]&~m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&m[509]&m[510])|(m[505]&~m[506]&m[507]&m[509]&m[510])|(~m[505]&m[506]&m[507]&m[509]&m[510]))&UnbiasedRNG[217])|((m[505]&m[506]&~m[507]&~m[509]&~m[510])|(m[505]&~m[506]&m[507]&~m[509]&~m[510])|(~m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&m[506]&m[507]&~m[509]&~m[510])|(m[505]&~m[506]&~m[507]&~m[509]&m[510])|(~m[505]&m[506]&~m[507]&~m[509]&m[510])|(m[505]&m[506]&~m[507]&~m[509]&m[510])|(~m[505]&~m[506]&m[507]&~m[509]&m[510])|(m[505]&~m[506]&m[507]&~m[509]&m[510])|(~m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&~m[509]&m[510])|(m[505]&m[506]&m[507]&m[509]&m[510]));
end

always @(posedge color4_clk) begin
    m[244] = (((m[240]&~m[241]&~m[242]&~m[243]&~m[247])|(~m[240]&m[241]&~m[242]&~m[243]&~m[247])|(~m[240]&~m[241]&m[242]&~m[243]&~m[247])|(m[240]&m[241]&~m[242]&m[243]&~m[247])|(m[240]&~m[241]&m[242]&m[243]&~m[247])|(~m[240]&m[241]&m[242]&m[243]&~m[247]))&BiasedRNG[223])|(((m[240]&~m[241]&~m[242]&~m[243]&m[247])|(~m[240]&m[241]&~m[242]&~m[243]&m[247])|(~m[240]&~m[241]&m[242]&~m[243]&m[247])|(m[240]&m[241]&~m[242]&m[243]&m[247])|(m[240]&~m[241]&m[242]&m[243]&m[247])|(~m[240]&m[241]&m[242]&m[243]&m[247]))&~BiasedRNG[223])|((m[240]&m[241]&~m[242]&~m[243]&~m[247])|(m[240]&~m[241]&m[242]&~m[243]&~m[247])|(~m[240]&m[241]&m[242]&~m[243]&~m[247])|(m[240]&m[241]&m[242]&~m[243]&~m[247])|(m[240]&m[241]&m[242]&m[243]&~m[247])|(m[240]&m[241]&~m[242]&~m[243]&m[247])|(m[240]&~m[241]&m[242]&~m[243]&m[247])|(~m[240]&m[241]&m[242]&~m[243]&m[247])|(m[240]&m[241]&m[242]&~m[243]&m[247])|(m[240]&m[241]&m[242]&m[243]&m[247]));
    m[249] = (((m[245]&~m[246]&~m[247]&~m[248]&~m[257])|(~m[245]&m[246]&~m[247]&~m[248]&~m[257])|(~m[245]&~m[246]&m[247]&~m[248]&~m[257])|(m[245]&m[246]&~m[247]&m[248]&~m[257])|(m[245]&~m[246]&m[247]&m[248]&~m[257])|(~m[245]&m[246]&m[247]&m[248]&~m[257]))&BiasedRNG[224])|(((m[245]&~m[246]&~m[247]&~m[248]&m[257])|(~m[245]&m[246]&~m[247]&~m[248]&m[257])|(~m[245]&~m[246]&m[247]&~m[248]&m[257])|(m[245]&m[246]&~m[247]&m[248]&m[257])|(m[245]&~m[246]&m[247]&m[248]&m[257])|(~m[245]&m[246]&m[247]&m[248]&m[257]))&~BiasedRNG[224])|((m[245]&m[246]&~m[247]&~m[248]&~m[257])|(m[245]&~m[246]&m[247]&~m[248]&~m[257])|(~m[245]&m[246]&m[247]&~m[248]&~m[257])|(m[245]&m[246]&m[247]&~m[248]&~m[257])|(m[245]&m[246]&m[247]&m[248]&~m[257])|(m[245]&m[246]&~m[247]&~m[248]&m[257])|(m[245]&~m[246]&m[247]&~m[248]&m[257])|(~m[245]&m[246]&m[247]&~m[248]&m[257])|(m[245]&m[246]&m[247]&~m[248]&m[257])|(m[245]&m[246]&m[247]&m[248]&m[257]));
    m[254] = (((m[250]&~m[251]&~m[252]&~m[253]&~m[262])|(~m[250]&m[251]&~m[252]&~m[253]&~m[262])|(~m[250]&~m[251]&m[252]&~m[253]&~m[262])|(m[250]&m[251]&~m[252]&m[253]&~m[262])|(m[250]&~m[251]&m[252]&m[253]&~m[262])|(~m[250]&m[251]&m[252]&m[253]&~m[262]))&BiasedRNG[225])|(((m[250]&~m[251]&~m[252]&~m[253]&m[262])|(~m[250]&m[251]&~m[252]&~m[253]&m[262])|(~m[250]&~m[251]&m[252]&~m[253]&m[262])|(m[250]&m[251]&~m[252]&m[253]&m[262])|(m[250]&~m[251]&m[252]&m[253]&m[262])|(~m[250]&m[251]&m[252]&m[253]&m[262]))&~BiasedRNG[225])|((m[250]&m[251]&~m[252]&~m[253]&~m[262])|(m[250]&~m[251]&m[252]&~m[253]&~m[262])|(~m[250]&m[251]&m[252]&~m[253]&~m[262])|(m[250]&m[251]&m[252]&~m[253]&~m[262])|(m[250]&m[251]&m[252]&m[253]&~m[262])|(m[250]&m[251]&~m[252]&~m[253]&m[262])|(m[250]&~m[251]&m[252]&~m[253]&m[262])|(~m[250]&m[251]&m[252]&~m[253]&m[262])|(m[250]&m[251]&m[252]&~m[253]&m[262])|(m[250]&m[251]&m[252]&m[253]&m[262]));
    m[259] = (((m[255]&~m[256]&~m[257]&~m[258]&~m[272])|(~m[255]&m[256]&~m[257]&~m[258]&~m[272])|(~m[255]&~m[256]&m[257]&~m[258]&~m[272])|(m[255]&m[256]&~m[257]&m[258]&~m[272])|(m[255]&~m[256]&m[257]&m[258]&~m[272])|(~m[255]&m[256]&m[257]&m[258]&~m[272]))&BiasedRNG[226])|(((m[255]&~m[256]&~m[257]&~m[258]&m[272])|(~m[255]&m[256]&~m[257]&~m[258]&m[272])|(~m[255]&~m[256]&m[257]&~m[258]&m[272])|(m[255]&m[256]&~m[257]&m[258]&m[272])|(m[255]&~m[256]&m[257]&m[258]&m[272])|(~m[255]&m[256]&m[257]&m[258]&m[272]))&~BiasedRNG[226])|((m[255]&m[256]&~m[257]&~m[258]&~m[272])|(m[255]&~m[256]&m[257]&~m[258]&~m[272])|(~m[255]&m[256]&m[257]&~m[258]&~m[272])|(m[255]&m[256]&m[257]&~m[258]&~m[272])|(m[255]&m[256]&m[257]&m[258]&~m[272])|(m[255]&m[256]&~m[257]&~m[258]&m[272])|(m[255]&~m[256]&m[257]&~m[258]&m[272])|(~m[255]&m[256]&m[257]&~m[258]&m[272])|(m[255]&m[256]&m[257]&~m[258]&m[272])|(m[255]&m[256]&m[257]&m[258]&m[272]));
    m[264] = (((m[260]&~m[261]&~m[262]&~m[263]&~m[277])|(~m[260]&m[261]&~m[262]&~m[263]&~m[277])|(~m[260]&~m[261]&m[262]&~m[263]&~m[277])|(m[260]&m[261]&~m[262]&m[263]&~m[277])|(m[260]&~m[261]&m[262]&m[263]&~m[277])|(~m[260]&m[261]&m[262]&m[263]&~m[277]))&BiasedRNG[227])|(((m[260]&~m[261]&~m[262]&~m[263]&m[277])|(~m[260]&m[261]&~m[262]&~m[263]&m[277])|(~m[260]&~m[261]&m[262]&~m[263]&m[277])|(m[260]&m[261]&~m[262]&m[263]&m[277])|(m[260]&~m[261]&m[262]&m[263]&m[277])|(~m[260]&m[261]&m[262]&m[263]&m[277]))&~BiasedRNG[227])|((m[260]&m[261]&~m[262]&~m[263]&~m[277])|(m[260]&~m[261]&m[262]&~m[263]&~m[277])|(~m[260]&m[261]&m[262]&~m[263]&~m[277])|(m[260]&m[261]&m[262]&~m[263]&~m[277])|(m[260]&m[261]&m[262]&m[263]&~m[277])|(m[260]&m[261]&~m[262]&~m[263]&m[277])|(m[260]&~m[261]&m[262]&~m[263]&m[277])|(~m[260]&m[261]&m[262]&~m[263]&m[277])|(m[260]&m[261]&m[262]&~m[263]&m[277])|(m[260]&m[261]&m[262]&m[263]&m[277]));
    m[269] = (((m[265]&~m[266]&~m[267]&~m[268]&~m[282])|(~m[265]&m[266]&~m[267]&~m[268]&~m[282])|(~m[265]&~m[266]&m[267]&~m[268]&~m[282])|(m[265]&m[266]&~m[267]&m[268]&~m[282])|(m[265]&~m[266]&m[267]&m[268]&~m[282])|(~m[265]&m[266]&m[267]&m[268]&~m[282]))&BiasedRNG[228])|(((m[265]&~m[266]&~m[267]&~m[268]&m[282])|(~m[265]&m[266]&~m[267]&~m[268]&m[282])|(~m[265]&~m[266]&m[267]&~m[268]&m[282])|(m[265]&m[266]&~m[267]&m[268]&m[282])|(m[265]&~m[266]&m[267]&m[268]&m[282])|(~m[265]&m[266]&m[267]&m[268]&m[282]))&~BiasedRNG[228])|((m[265]&m[266]&~m[267]&~m[268]&~m[282])|(m[265]&~m[266]&m[267]&~m[268]&~m[282])|(~m[265]&m[266]&m[267]&~m[268]&~m[282])|(m[265]&m[266]&m[267]&~m[268]&~m[282])|(m[265]&m[266]&m[267]&m[268]&~m[282])|(m[265]&m[266]&~m[267]&~m[268]&m[282])|(m[265]&~m[266]&m[267]&~m[268]&m[282])|(~m[265]&m[266]&m[267]&~m[268]&m[282])|(m[265]&m[266]&m[267]&~m[268]&m[282])|(m[265]&m[266]&m[267]&m[268]&m[282]));
    m[274] = (((m[270]&~m[271]&~m[272]&~m[273]&~m[292])|(~m[270]&m[271]&~m[272]&~m[273]&~m[292])|(~m[270]&~m[271]&m[272]&~m[273]&~m[292])|(m[270]&m[271]&~m[272]&m[273]&~m[292])|(m[270]&~m[271]&m[272]&m[273]&~m[292])|(~m[270]&m[271]&m[272]&m[273]&~m[292]))&BiasedRNG[229])|(((m[270]&~m[271]&~m[272]&~m[273]&m[292])|(~m[270]&m[271]&~m[272]&~m[273]&m[292])|(~m[270]&~m[271]&m[272]&~m[273]&m[292])|(m[270]&m[271]&~m[272]&m[273]&m[292])|(m[270]&~m[271]&m[272]&m[273]&m[292])|(~m[270]&m[271]&m[272]&m[273]&m[292]))&~BiasedRNG[229])|((m[270]&m[271]&~m[272]&~m[273]&~m[292])|(m[270]&~m[271]&m[272]&~m[273]&~m[292])|(~m[270]&m[271]&m[272]&~m[273]&~m[292])|(m[270]&m[271]&m[272]&~m[273]&~m[292])|(m[270]&m[271]&m[272]&m[273]&~m[292])|(m[270]&m[271]&~m[272]&~m[273]&m[292])|(m[270]&~m[271]&m[272]&~m[273]&m[292])|(~m[270]&m[271]&m[272]&~m[273]&m[292])|(m[270]&m[271]&m[272]&~m[273]&m[292])|(m[270]&m[271]&m[272]&m[273]&m[292]));
    m[279] = (((m[275]&~m[276]&~m[277]&~m[278]&~m[297])|(~m[275]&m[276]&~m[277]&~m[278]&~m[297])|(~m[275]&~m[276]&m[277]&~m[278]&~m[297])|(m[275]&m[276]&~m[277]&m[278]&~m[297])|(m[275]&~m[276]&m[277]&m[278]&~m[297])|(~m[275]&m[276]&m[277]&m[278]&~m[297]))&BiasedRNG[230])|(((m[275]&~m[276]&~m[277]&~m[278]&m[297])|(~m[275]&m[276]&~m[277]&~m[278]&m[297])|(~m[275]&~m[276]&m[277]&~m[278]&m[297])|(m[275]&m[276]&~m[277]&m[278]&m[297])|(m[275]&~m[276]&m[277]&m[278]&m[297])|(~m[275]&m[276]&m[277]&m[278]&m[297]))&~BiasedRNG[230])|((m[275]&m[276]&~m[277]&~m[278]&~m[297])|(m[275]&~m[276]&m[277]&~m[278]&~m[297])|(~m[275]&m[276]&m[277]&~m[278]&~m[297])|(m[275]&m[276]&m[277]&~m[278]&~m[297])|(m[275]&m[276]&m[277]&m[278]&~m[297])|(m[275]&m[276]&~m[277]&~m[278]&m[297])|(m[275]&~m[276]&m[277]&~m[278]&m[297])|(~m[275]&m[276]&m[277]&~m[278]&m[297])|(m[275]&m[276]&m[277]&~m[278]&m[297])|(m[275]&m[276]&m[277]&m[278]&m[297]));
    m[284] = (((m[280]&~m[281]&~m[282]&~m[283]&~m[302])|(~m[280]&m[281]&~m[282]&~m[283]&~m[302])|(~m[280]&~m[281]&m[282]&~m[283]&~m[302])|(m[280]&m[281]&~m[282]&m[283]&~m[302])|(m[280]&~m[281]&m[282]&m[283]&~m[302])|(~m[280]&m[281]&m[282]&m[283]&~m[302]))&BiasedRNG[231])|(((m[280]&~m[281]&~m[282]&~m[283]&m[302])|(~m[280]&m[281]&~m[282]&~m[283]&m[302])|(~m[280]&~m[281]&m[282]&~m[283]&m[302])|(m[280]&m[281]&~m[282]&m[283]&m[302])|(m[280]&~m[281]&m[282]&m[283]&m[302])|(~m[280]&m[281]&m[282]&m[283]&m[302]))&~BiasedRNG[231])|((m[280]&m[281]&~m[282]&~m[283]&~m[302])|(m[280]&~m[281]&m[282]&~m[283]&~m[302])|(~m[280]&m[281]&m[282]&~m[283]&~m[302])|(m[280]&m[281]&m[282]&~m[283]&~m[302])|(m[280]&m[281]&m[282]&m[283]&~m[302])|(m[280]&m[281]&~m[282]&~m[283]&m[302])|(m[280]&~m[281]&m[282]&~m[283]&m[302])|(~m[280]&m[281]&m[282]&~m[283]&m[302])|(m[280]&m[281]&m[282]&~m[283]&m[302])|(m[280]&m[281]&m[282]&m[283]&m[302]));
    m[289] = (((m[285]&~m[286]&~m[287]&~m[288]&~m[307])|(~m[285]&m[286]&~m[287]&~m[288]&~m[307])|(~m[285]&~m[286]&m[287]&~m[288]&~m[307])|(m[285]&m[286]&~m[287]&m[288]&~m[307])|(m[285]&~m[286]&m[287]&m[288]&~m[307])|(~m[285]&m[286]&m[287]&m[288]&~m[307]))&BiasedRNG[232])|(((m[285]&~m[286]&~m[287]&~m[288]&m[307])|(~m[285]&m[286]&~m[287]&~m[288]&m[307])|(~m[285]&~m[286]&m[287]&~m[288]&m[307])|(m[285]&m[286]&~m[287]&m[288]&m[307])|(m[285]&~m[286]&m[287]&m[288]&m[307])|(~m[285]&m[286]&m[287]&m[288]&m[307]))&~BiasedRNG[232])|((m[285]&m[286]&~m[287]&~m[288]&~m[307])|(m[285]&~m[286]&m[287]&~m[288]&~m[307])|(~m[285]&m[286]&m[287]&~m[288]&~m[307])|(m[285]&m[286]&m[287]&~m[288]&~m[307])|(m[285]&m[286]&m[287]&m[288]&~m[307])|(m[285]&m[286]&~m[287]&~m[288]&m[307])|(m[285]&~m[286]&m[287]&~m[288]&m[307])|(~m[285]&m[286]&m[287]&~m[288]&m[307])|(m[285]&m[286]&m[287]&~m[288]&m[307])|(m[285]&m[286]&m[287]&m[288]&m[307]));
    m[294] = (((m[290]&~m[291]&~m[292]&~m[293]&~m[317])|(~m[290]&m[291]&~m[292]&~m[293]&~m[317])|(~m[290]&~m[291]&m[292]&~m[293]&~m[317])|(m[290]&m[291]&~m[292]&m[293]&~m[317])|(m[290]&~m[291]&m[292]&m[293]&~m[317])|(~m[290]&m[291]&m[292]&m[293]&~m[317]))&BiasedRNG[233])|(((m[290]&~m[291]&~m[292]&~m[293]&m[317])|(~m[290]&m[291]&~m[292]&~m[293]&m[317])|(~m[290]&~m[291]&m[292]&~m[293]&m[317])|(m[290]&m[291]&~m[292]&m[293]&m[317])|(m[290]&~m[291]&m[292]&m[293]&m[317])|(~m[290]&m[291]&m[292]&m[293]&m[317]))&~BiasedRNG[233])|((m[290]&m[291]&~m[292]&~m[293]&~m[317])|(m[290]&~m[291]&m[292]&~m[293]&~m[317])|(~m[290]&m[291]&m[292]&~m[293]&~m[317])|(m[290]&m[291]&m[292]&~m[293]&~m[317])|(m[290]&m[291]&m[292]&m[293]&~m[317])|(m[290]&m[291]&~m[292]&~m[293]&m[317])|(m[290]&~m[291]&m[292]&~m[293]&m[317])|(~m[290]&m[291]&m[292]&~m[293]&m[317])|(m[290]&m[291]&m[292]&~m[293]&m[317])|(m[290]&m[291]&m[292]&m[293]&m[317]));
    m[299] = (((m[295]&~m[296]&~m[297]&~m[298]&~m[322])|(~m[295]&m[296]&~m[297]&~m[298]&~m[322])|(~m[295]&~m[296]&m[297]&~m[298]&~m[322])|(m[295]&m[296]&~m[297]&m[298]&~m[322])|(m[295]&~m[296]&m[297]&m[298]&~m[322])|(~m[295]&m[296]&m[297]&m[298]&~m[322]))&BiasedRNG[234])|(((m[295]&~m[296]&~m[297]&~m[298]&m[322])|(~m[295]&m[296]&~m[297]&~m[298]&m[322])|(~m[295]&~m[296]&m[297]&~m[298]&m[322])|(m[295]&m[296]&~m[297]&m[298]&m[322])|(m[295]&~m[296]&m[297]&m[298]&m[322])|(~m[295]&m[296]&m[297]&m[298]&m[322]))&~BiasedRNG[234])|((m[295]&m[296]&~m[297]&~m[298]&~m[322])|(m[295]&~m[296]&m[297]&~m[298]&~m[322])|(~m[295]&m[296]&m[297]&~m[298]&~m[322])|(m[295]&m[296]&m[297]&~m[298]&~m[322])|(m[295]&m[296]&m[297]&m[298]&~m[322])|(m[295]&m[296]&~m[297]&~m[298]&m[322])|(m[295]&~m[296]&m[297]&~m[298]&m[322])|(~m[295]&m[296]&m[297]&~m[298]&m[322])|(m[295]&m[296]&m[297]&~m[298]&m[322])|(m[295]&m[296]&m[297]&m[298]&m[322]));
    m[304] = (((m[300]&~m[301]&~m[302]&~m[303]&~m[327])|(~m[300]&m[301]&~m[302]&~m[303]&~m[327])|(~m[300]&~m[301]&m[302]&~m[303]&~m[327])|(m[300]&m[301]&~m[302]&m[303]&~m[327])|(m[300]&~m[301]&m[302]&m[303]&~m[327])|(~m[300]&m[301]&m[302]&m[303]&~m[327]))&BiasedRNG[235])|(((m[300]&~m[301]&~m[302]&~m[303]&m[327])|(~m[300]&m[301]&~m[302]&~m[303]&m[327])|(~m[300]&~m[301]&m[302]&~m[303]&m[327])|(m[300]&m[301]&~m[302]&m[303]&m[327])|(m[300]&~m[301]&m[302]&m[303]&m[327])|(~m[300]&m[301]&m[302]&m[303]&m[327]))&~BiasedRNG[235])|((m[300]&m[301]&~m[302]&~m[303]&~m[327])|(m[300]&~m[301]&m[302]&~m[303]&~m[327])|(~m[300]&m[301]&m[302]&~m[303]&~m[327])|(m[300]&m[301]&m[302]&~m[303]&~m[327])|(m[300]&m[301]&m[302]&m[303]&~m[327])|(m[300]&m[301]&~m[302]&~m[303]&m[327])|(m[300]&~m[301]&m[302]&~m[303]&m[327])|(~m[300]&m[301]&m[302]&~m[303]&m[327])|(m[300]&m[301]&m[302]&~m[303]&m[327])|(m[300]&m[301]&m[302]&m[303]&m[327]));
    m[309] = (((m[305]&~m[306]&~m[307]&~m[308]&~m[332])|(~m[305]&m[306]&~m[307]&~m[308]&~m[332])|(~m[305]&~m[306]&m[307]&~m[308]&~m[332])|(m[305]&m[306]&~m[307]&m[308]&~m[332])|(m[305]&~m[306]&m[307]&m[308]&~m[332])|(~m[305]&m[306]&m[307]&m[308]&~m[332]))&BiasedRNG[236])|(((m[305]&~m[306]&~m[307]&~m[308]&m[332])|(~m[305]&m[306]&~m[307]&~m[308]&m[332])|(~m[305]&~m[306]&m[307]&~m[308]&m[332])|(m[305]&m[306]&~m[307]&m[308]&m[332])|(m[305]&~m[306]&m[307]&m[308]&m[332])|(~m[305]&m[306]&m[307]&m[308]&m[332]))&~BiasedRNG[236])|((m[305]&m[306]&~m[307]&~m[308]&~m[332])|(m[305]&~m[306]&m[307]&~m[308]&~m[332])|(~m[305]&m[306]&m[307]&~m[308]&~m[332])|(m[305]&m[306]&m[307]&~m[308]&~m[332])|(m[305]&m[306]&m[307]&m[308]&~m[332])|(m[305]&m[306]&~m[307]&~m[308]&m[332])|(m[305]&~m[306]&m[307]&~m[308]&m[332])|(~m[305]&m[306]&m[307]&~m[308]&m[332])|(m[305]&m[306]&m[307]&~m[308]&m[332])|(m[305]&m[306]&m[307]&m[308]&m[332]));
    m[314] = (((m[310]&~m[311]&~m[312]&~m[313]&~m[337])|(~m[310]&m[311]&~m[312]&~m[313]&~m[337])|(~m[310]&~m[311]&m[312]&~m[313]&~m[337])|(m[310]&m[311]&~m[312]&m[313]&~m[337])|(m[310]&~m[311]&m[312]&m[313]&~m[337])|(~m[310]&m[311]&m[312]&m[313]&~m[337]))&BiasedRNG[237])|(((m[310]&~m[311]&~m[312]&~m[313]&m[337])|(~m[310]&m[311]&~m[312]&~m[313]&m[337])|(~m[310]&~m[311]&m[312]&~m[313]&m[337])|(m[310]&m[311]&~m[312]&m[313]&m[337])|(m[310]&~m[311]&m[312]&m[313]&m[337])|(~m[310]&m[311]&m[312]&m[313]&m[337]))&~BiasedRNG[237])|((m[310]&m[311]&~m[312]&~m[313]&~m[337])|(m[310]&~m[311]&m[312]&~m[313]&~m[337])|(~m[310]&m[311]&m[312]&~m[313]&~m[337])|(m[310]&m[311]&m[312]&~m[313]&~m[337])|(m[310]&m[311]&m[312]&m[313]&~m[337])|(m[310]&m[311]&~m[312]&~m[313]&m[337])|(m[310]&~m[311]&m[312]&~m[313]&m[337])|(~m[310]&m[311]&m[312]&~m[313]&m[337])|(m[310]&m[311]&m[312]&~m[313]&m[337])|(m[310]&m[311]&m[312]&m[313]&m[337]));
    m[319] = (((m[315]&~m[316]&~m[317]&~m[318]&~m[347])|(~m[315]&m[316]&~m[317]&~m[318]&~m[347])|(~m[315]&~m[316]&m[317]&~m[318]&~m[347])|(m[315]&m[316]&~m[317]&m[318]&~m[347])|(m[315]&~m[316]&m[317]&m[318]&~m[347])|(~m[315]&m[316]&m[317]&m[318]&~m[347]))&BiasedRNG[238])|(((m[315]&~m[316]&~m[317]&~m[318]&m[347])|(~m[315]&m[316]&~m[317]&~m[318]&m[347])|(~m[315]&~m[316]&m[317]&~m[318]&m[347])|(m[315]&m[316]&~m[317]&m[318]&m[347])|(m[315]&~m[316]&m[317]&m[318]&m[347])|(~m[315]&m[316]&m[317]&m[318]&m[347]))&~BiasedRNG[238])|((m[315]&m[316]&~m[317]&~m[318]&~m[347])|(m[315]&~m[316]&m[317]&~m[318]&~m[347])|(~m[315]&m[316]&m[317]&~m[318]&~m[347])|(m[315]&m[316]&m[317]&~m[318]&~m[347])|(m[315]&m[316]&m[317]&m[318]&~m[347])|(m[315]&m[316]&~m[317]&~m[318]&m[347])|(m[315]&~m[316]&m[317]&~m[318]&m[347])|(~m[315]&m[316]&m[317]&~m[318]&m[347])|(m[315]&m[316]&m[317]&~m[318]&m[347])|(m[315]&m[316]&m[317]&m[318]&m[347]));
    m[324] = (((m[320]&~m[321]&~m[322]&~m[323]&~m[352])|(~m[320]&m[321]&~m[322]&~m[323]&~m[352])|(~m[320]&~m[321]&m[322]&~m[323]&~m[352])|(m[320]&m[321]&~m[322]&m[323]&~m[352])|(m[320]&~m[321]&m[322]&m[323]&~m[352])|(~m[320]&m[321]&m[322]&m[323]&~m[352]))&BiasedRNG[239])|(((m[320]&~m[321]&~m[322]&~m[323]&m[352])|(~m[320]&m[321]&~m[322]&~m[323]&m[352])|(~m[320]&~m[321]&m[322]&~m[323]&m[352])|(m[320]&m[321]&~m[322]&m[323]&m[352])|(m[320]&~m[321]&m[322]&m[323]&m[352])|(~m[320]&m[321]&m[322]&m[323]&m[352]))&~BiasedRNG[239])|((m[320]&m[321]&~m[322]&~m[323]&~m[352])|(m[320]&~m[321]&m[322]&~m[323]&~m[352])|(~m[320]&m[321]&m[322]&~m[323]&~m[352])|(m[320]&m[321]&m[322]&~m[323]&~m[352])|(m[320]&m[321]&m[322]&m[323]&~m[352])|(m[320]&m[321]&~m[322]&~m[323]&m[352])|(m[320]&~m[321]&m[322]&~m[323]&m[352])|(~m[320]&m[321]&m[322]&~m[323]&m[352])|(m[320]&m[321]&m[322]&~m[323]&m[352])|(m[320]&m[321]&m[322]&m[323]&m[352]));
    m[329] = (((m[325]&~m[326]&~m[327]&~m[328]&~m[357])|(~m[325]&m[326]&~m[327]&~m[328]&~m[357])|(~m[325]&~m[326]&m[327]&~m[328]&~m[357])|(m[325]&m[326]&~m[327]&m[328]&~m[357])|(m[325]&~m[326]&m[327]&m[328]&~m[357])|(~m[325]&m[326]&m[327]&m[328]&~m[357]))&BiasedRNG[240])|(((m[325]&~m[326]&~m[327]&~m[328]&m[357])|(~m[325]&m[326]&~m[327]&~m[328]&m[357])|(~m[325]&~m[326]&m[327]&~m[328]&m[357])|(m[325]&m[326]&~m[327]&m[328]&m[357])|(m[325]&~m[326]&m[327]&m[328]&m[357])|(~m[325]&m[326]&m[327]&m[328]&m[357]))&~BiasedRNG[240])|((m[325]&m[326]&~m[327]&~m[328]&~m[357])|(m[325]&~m[326]&m[327]&~m[328]&~m[357])|(~m[325]&m[326]&m[327]&~m[328]&~m[357])|(m[325]&m[326]&m[327]&~m[328]&~m[357])|(m[325]&m[326]&m[327]&m[328]&~m[357])|(m[325]&m[326]&~m[327]&~m[328]&m[357])|(m[325]&~m[326]&m[327]&~m[328]&m[357])|(~m[325]&m[326]&m[327]&~m[328]&m[357])|(m[325]&m[326]&m[327]&~m[328]&m[357])|(m[325]&m[326]&m[327]&m[328]&m[357]));
    m[334] = (((m[330]&~m[331]&~m[332]&~m[333]&~m[362])|(~m[330]&m[331]&~m[332]&~m[333]&~m[362])|(~m[330]&~m[331]&m[332]&~m[333]&~m[362])|(m[330]&m[331]&~m[332]&m[333]&~m[362])|(m[330]&~m[331]&m[332]&m[333]&~m[362])|(~m[330]&m[331]&m[332]&m[333]&~m[362]))&BiasedRNG[241])|(((m[330]&~m[331]&~m[332]&~m[333]&m[362])|(~m[330]&m[331]&~m[332]&~m[333]&m[362])|(~m[330]&~m[331]&m[332]&~m[333]&m[362])|(m[330]&m[331]&~m[332]&m[333]&m[362])|(m[330]&~m[331]&m[332]&m[333]&m[362])|(~m[330]&m[331]&m[332]&m[333]&m[362]))&~BiasedRNG[241])|((m[330]&m[331]&~m[332]&~m[333]&~m[362])|(m[330]&~m[331]&m[332]&~m[333]&~m[362])|(~m[330]&m[331]&m[332]&~m[333]&~m[362])|(m[330]&m[331]&m[332]&~m[333]&~m[362])|(m[330]&m[331]&m[332]&m[333]&~m[362])|(m[330]&m[331]&~m[332]&~m[333]&m[362])|(m[330]&~m[331]&m[332]&~m[333]&m[362])|(~m[330]&m[331]&m[332]&~m[333]&m[362])|(m[330]&m[331]&m[332]&~m[333]&m[362])|(m[330]&m[331]&m[332]&m[333]&m[362]));
    m[339] = (((m[335]&~m[336]&~m[337]&~m[338]&~m[367])|(~m[335]&m[336]&~m[337]&~m[338]&~m[367])|(~m[335]&~m[336]&m[337]&~m[338]&~m[367])|(m[335]&m[336]&~m[337]&m[338]&~m[367])|(m[335]&~m[336]&m[337]&m[338]&~m[367])|(~m[335]&m[336]&m[337]&m[338]&~m[367]))&BiasedRNG[242])|(((m[335]&~m[336]&~m[337]&~m[338]&m[367])|(~m[335]&m[336]&~m[337]&~m[338]&m[367])|(~m[335]&~m[336]&m[337]&~m[338]&m[367])|(m[335]&m[336]&~m[337]&m[338]&m[367])|(m[335]&~m[336]&m[337]&m[338]&m[367])|(~m[335]&m[336]&m[337]&m[338]&m[367]))&~BiasedRNG[242])|((m[335]&m[336]&~m[337]&~m[338]&~m[367])|(m[335]&~m[336]&m[337]&~m[338]&~m[367])|(~m[335]&m[336]&m[337]&~m[338]&~m[367])|(m[335]&m[336]&m[337]&~m[338]&~m[367])|(m[335]&m[336]&m[337]&m[338]&~m[367])|(m[335]&m[336]&~m[337]&~m[338]&m[367])|(m[335]&~m[336]&m[337]&~m[338]&m[367])|(~m[335]&m[336]&m[337]&~m[338]&m[367])|(m[335]&m[336]&m[337]&~m[338]&m[367])|(m[335]&m[336]&m[337]&m[338]&m[367]));
    m[344] = (((m[340]&~m[341]&~m[342]&~m[343]&~m[372])|(~m[340]&m[341]&~m[342]&~m[343]&~m[372])|(~m[340]&~m[341]&m[342]&~m[343]&~m[372])|(m[340]&m[341]&~m[342]&m[343]&~m[372])|(m[340]&~m[341]&m[342]&m[343]&~m[372])|(~m[340]&m[341]&m[342]&m[343]&~m[372]))&BiasedRNG[243])|(((m[340]&~m[341]&~m[342]&~m[343]&m[372])|(~m[340]&m[341]&~m[342]&~m[343]&m[372])|(~m[340]&~m[341]&m[342]&~m[343]&m[372])|(m[340]&m[341]&~m[342]&m[343]&m[372])|(m[340]&~m[341]&m[342]&m[343]&m[372])|(~m[340]&m[341]&m[342]&m[343]&m[372]))&~BiasedRNG[243])|((m[340]&m[341]&~m[342]&~m[343]&~m[372])|(m[340]&~m[341]&m[342]&~m[343]&~m[372])|(~m[340]&m[341]&m[342]&~m[343]&~m[372])|(m[340]&m[341]&m[342]&~m[343]&~m[372])|(m[340]&m[341]&m[342]&m[343]&~m[372])|(m[340]&m[341]&~m[342]&~m[343]&m[372])|(m[340]&~m[341]&m[342]&~m[343]&m[372])|(~m[340]&m[341]&m[342]&~m[343]&m[372])|(m[340]&m[341]&m[342]&~m[343]&m[372])|(m[340]&m[341]&m[342]&m[343]&m[372]));
    m[349] = (((m[345]&~m[346]&~m[347]&~m[348]&~m[382])|(~m[345]&m[346]&~m[347]&~m[348]&~m[382])|(~m[345]&~m[346]&m[347]&~m[348]&~m[382])|(m[345]&m[346]&~m[347]&m[348]&~m[382])|(m[345]&~m[346]&m[347]&m[348]&~m[382])|(~m[345]&m[346]&m[347]&m[348]&~m[382]))&BiasedRNG[244])|(((m[345]&~m[346]&~m[347]&~m[348]&m[382])|(~m[345]&m[346]&~m[347]&~m[348]&m[382])|(~m[345]&~m[346]&m[347]&~m[348]&m[382])|(m[345]&m[346]&~m[347]&m[348]&m[382])|(m[345]&~m[346]&m[347]&m[348]&m[382])|(~m[345]&m[346]&m[347]&m[348]&m[382]))&~BiasedRNG[244])|((m[345]&m[346]&~m[347]&~m[348]&~m[382])|(m[345]&~m[346]&m[347]&~m[348]&~m[382])|(~m[345]&m[346]&m[347]&~m[348]&~m[382])|(m[345]&m[346]&m[347]&~m[348]&~m[382])|(m[345]&m[346]&m[347]&m[348]&~m[382])|(m[345]&m[346]&~m[347]&~m[348]&m[382])|(m[345]&~m[346]&m[347]&~m[348]&m[382])|(~m[345]&m[346]&m[347]&~m[348]&m[382])|(m[345]&m[346]&m[347]&~m[348]&m[382])|(m[345]&m[346]&m[347]&m[348]&m[382]));
    m[354] = (((m[350]&~m[351]&~m[352]&~m[353]&~m[387])|(~m[350]&m[351]&~m[352]&~m[353]&~m[387])|(~m[350]&~m[351]&m[352]&~m[353]&~m[387])|(m[350]&m[351]&~m[352]&m[353]&~m[387])|(m[350]&~m[351]&m[352]&m[353]&~m[387])|(~m[350]&m[351]&m[352]&m[353]&~m[387]))&BiasedRNG[245])|(((m[350]&~m[351]&~m[352]&~m[353]&m[387])|(~m[350]&m[351]&~m[352]&~m[353]&m[387])|(~m[350]&~m[351]&m[352]&~m[353]&m[387])|(m[350]&m[351]&~m[352]&m[353]&m[387])|(m[350]&~m[351]&m[352]&m[353]&m[387])|(~m[350]&m[351]&m[352]&m[353]&m[387]))&~BiasedRNG[245])|((m[350]&m[351]&~m[352]&~m[353]&~m[387])|(m[350]&~m[351]&m[352]&~m[353]&~m[387])|(~m[350]&m[351]&m[352]&~m[353]&~m[387])|(m[350]&m[351]&m[352]&~m[353]&~m[387])|(m[350]&m[351]&m[352]&m[353]&~m[387])|(m[350]&m[351]&~m[352]&~m[353]&m[387])|(m[350]&~m[351]&m[352]&~m[353]&m[387])|(~m[350]&m[351]&m[352]&~m[353]&m[387])|(m[350]&m[351]&m[352]&~m[353]&m[387])|(m[350]&m[351]&m[352]&m[353]&m[387]));
    m[359] = (((m[355]&~m[356]&~m[357]&~m[358]&~m[392])|(~m[355]&m[356]&~m[357]&~m[358]&~m[392])|(~m[355]&~m[356]&m[357]&~m[358]&~m[392])|(m[355]&m[356]&~m[357]&m[358]&~m[392])|(m[355]&~m[356]&m[357]&m[358]&~m[392])|(~m[355]&m[356]&m[357]&m[358]&~m[392]))&BiasedRNG[246])|(((m[355]&~m[356]&~m[357]&~m[358]&m[392])|(~m[355]&m[356]&~m[357]&~m[358]&m[392])|(~m[355]&~m[356]&m[357]&~m[358]&m[392])|(m[355]&m[356]&~m[357]&m[358]&m[392])|(m[355]&~m[356]&m[357]&m[358]&m[392])|(~m[355]&m[356]&m[357]&m[358]&m[392]))&~BiasedRNG[246])|((m[355]&m[356]&~m[357]&~m[358]&~m[392])|(m[355]&~m[356]&m[357]&~m[358]&~m[392])|(~m[355]&m[356]&m[357]&~m[358]&~m[392])|(m[355]&m[356]&m[357]&~m[358]&~m[392])|(m[355]&m[356]&m[357]&m[358]&~m[392])|(m[355]&m[356]&~m[357]&~m[358]&m[392])|(m[355]&~m[356]&m[357]&~m[358]&m[392])|(~m[355]&m[356]&m[357]&~m[358]&m[392])|(m[355]&m[356]&m[357]&~m[358]&m[392])|(m[355]&m[356]&m[357]&m[358]&m[392]));
    m[364] = (((m[360]&~m[361]&~m[362]&~m[363]&~m[397])|(~m[360]&m[361]&~m[362]&~m[363]&~m[397])|(~m[360]&~m[361]&m[362]&~m[363]&~m[397])|(m[360]&m[361]&~m[362]&m[363]&~m[397])|(m[360]&~m[361]&m[362]&m[363]&~m[397])|(~m[360]&m[361]&m[362]&m[363]&~m[397]))&BiasedRNG[247])|(((m[360]&~m[361]&~m[362]&~m[363]&m[397])|(~m[360]&m[361]&~m[362]&~m[363]&m[397])|(~m[360]&~m[361]&m[362]&~m[363]&m[397])|(m[360]&m[361]&~m[362]&m[363]&m[397])|(m[360]&~m[361]&m[362]&m[363]&m[397])|(~m[360]&m[361]&m[362]&m[363]&m[397]))&~BiasedRNG[247])|((m[360]&m[361]&~m[362]&~m[363]&~m[397])|(m[360]&~m[361]&m[362]&~m[363]&~m[397])|(~m[360]&m[361]&m[362]&~m[363]&~m[397])|(m[360]&m[361]&m[362]&~m[363]&~m[397])|(m[360]&m[361]&m[362]&m[363]&~m[397])|(m[360]&m[361]&~m[362]&~m[363]&m[397])|(m[360]&~m[361]&m[362]&~m[363]&m[397])|(~m[360]&m[361]&m[362]&~m[363]&m[397])|(m[360]&m[361]&m[362]&~m[363]&m[397])|(m[360]&m[361]&m[362]&m[363]&m[397]));
    m[369] = (((m[365]&~m[366]&~m[367]&~m[368]&~m[402])|(~m[365]&m[366]&~m[367]&~m[368]&~m[402])|(~m[365]&~m[366]&m[367]&~m[368]&~m[402])|(m[365]&m[366]&~m[367]&m[368]&~m[402])|(m[365]&~m[366]&m[367]&m[368]&~m[402])|(~m[365]&m[366]&m[367]&m[368]&~m[402]))&BiasedRNG[248])|(((m[365]&~m[366]&~m[367]&~m[368]&m[402])|(~m[365]&m[366]&~m[367]&~m[368]&m[402])|(~m[365]&~m[366]&m[367]&~m[368]&m[402])|(m[365]&m[366]&~m[367]&m[368]&m[402])|(m[365]&~m[366]&m[367]&m[368]&m[402])|(~m[365]&m[366]&m[367]&m[368]&m[402]))&~BiasedRNG[248])|((m[365]&m[366]&~m[367]&~m[368]&~m[402])|(m[365]&~m[366]&m[367]&~m[368]&~m[402])|(~m[365]&m[366]&m[367]&~m[368]&~m[402])|(m[365]&m[366]&m[367]&~m[368]&~m[402])|(m[365]&m[366]&m[367]&m[368]&~m[402])|(m[365]&m[366]&~m[367]&~m[368]&m[402])|(m[365]&~m[366]&m[367]&~m[368]&m[402])|(~m[365]&m[366]&m[367]&~m[368]&m[402])|(m[365]&m[366]&m[367]&~m[368]&m[402])|(m[365]&m[366]&m[367]&m[368]&m[402]));
    m[374] = (((m[370]&~m[371]&~m[372]&~m[373]&~m[407])|(~m[370]&m[371]&~m[372]&~m[373]&~m[407])|(~m[370]&~m[371]&m[372]&~m[373]&~m[407])|(m[370]&m[371]&~m[372]&m[373]&~m[407])|(m[370]&~m[371]&m[372]&m[373]&~m[407])|(~m[370]&m[371]&m[372]&m[373]&~m[407]))&BiasedRNG[249])|(((m[370]&~m[371]&~m[372]&~m[373]&m[407])|(~m[370]&m[371]&~m[372]&~m[373]&m[407])|(~m[370]&~m[371]&m[372]&~m[373]&m[407])|(m[370]&m[371]&~m[372]&m[373]&m[407])|(m[370]&~m[371]&m[372]&m[373]&m[407])|(~m[370]&m[371]&m[372]&m[373]&m[407]))&~BiasedRNG[249])|((m[370]&m[371]&~m[372]&~m[373]&~m[407])|(m[370]&~m[371]&m[372]&~m[373]&~m[407])|(~m[370]&m[371]&m[372]&~m[373]&~m[407])|(m[370]&m[371]&m[372]&~m[373]&~m[407])|(m[370]&m[371]&m[372]&m[373]&~m[407])|(m[370]&m[371]&~m[372]&~m[373]&m[407])|(m[370]&~m[371]&m[372]&~m[373]&m[407])|(~m[370]&m[371]&m[372]&~m[373]&m[407])|(m[370]&m[371]&m[372]&~m[373]&m[407])|(m[370]&m[371]&m[372]&m[373]&m[407]));
    m[379] = (((m[375]&~m[376]&~m[377]&~m[378]&~m[412])|(~m[375]&m[376]&~m[377]&~m[378]&~m[412])|(~m[375]&~m[376]&m[377]&~m[378]&~m[412])|(m[375]&m[376]&~m[377]&m[378]&~m[412])|(m[375]&~m[376]&m[377]&m[378]&~m[412])|(~m[375]&m[376]&m[377]&m[378]&~m[412]))&BiasedRNG[250])|(((m[375]&~m[376]&~m[377]&~m[378]&m[412])|(~m[375]&m[376]&~m[377]&~m[378]&m[412])|(~m[375]&~m[376]&m[377]&~m[378]&m[412])|(m[375]&m[376]&~m[377]&m[378]&m[412])|(m[375]&~m[376]&m[377]&m[378]&m[412])|(~m[375]&m[376]&m[377]&m[378]&m[412]))&~BiasedRNG[250])|((m[375]&m[376]&~m[377]&~m[378]&~m[412])|(m[375]&~m[376]&m[377]&~m[378]&~m[412])|(~m[375]&m[376]&m[377]&~m[378]&~m[412])|(m[375]&m[376]&m[377]&~m[378]&~m[412])|(m[375]&m[376]&m[377]&m[378]&~m[412])|(m[375]&m[376]&~m[377]&~m[378]&m[412])|(m[375]&~m[376]&m[377]&~m[378]&m[412])|(~m[375]&m[376]&m[377]&~m[378]&m[412])|(m[375]&m[376]&m[377]&~m[378]&m[412])|(m[375]&m[376]&m[377]&m[378]&m[412]));
    m[384] = (((m[380]&~m[381]&~m[382]&~m[383]&~m[415])|(~m[380]&m[381]&~m[382]&~m[383]&~m[415])|(~m[380]&~m[381]&m[382]&~m[383]&~m[415])|(m[380]&m[381]&~m[382]&m[383]&~m[415])|(m[380]&~m[381]&m[382]&m[383]&~m[415])|(~m[380]&m[381]&m[382]&m[383]&~m[415]))&BiasedRNG[251])|(((m[380]&~m[381]&~m[382]&~m[383]&m[415])|(~m[380]&m[381]&~m[382]&~m[383]&m[415])|(~m[380]&~m[381]&m[382]&~m[383]&m[415])|(m[380]&m[381]&~m[382]&m[383]&m[415])|(m[380]&~m[381]&m[382]&m[383]&m[415])|(~m[380]&m[381]&m[382]&m[383]&m[415]))&~BiasedRNG[251])|((m[380]&m[381]&~m[382]&~m[383]&~m[415])|(m[380]&~m[381]&m[382]&~m[383]&~m[415])|(~m[380]&m[381]&m[382]&~m[383]&~m[415])|(m[380]&m[381]&m[382]&~m[383]&~m[415])|(m[380]&m[381]&m[382]&m[383]&~m[415])|(m[380]&m[381]&~m[382]&~m[383]&m[415])|(m[380]&~m[381]&m[382]&~m[383]&m[415])|(~m[380]&m[381]&m[382]&~m[383]&m[415])|(m[380]&m[381]&m[382]&~m[383]&m[415])|(m[380]&m[381]&m[382]&m[383]&m[415]));
    m[389] = (((m[385]&~m[386]&~m[387]&~m[388]&~m[417])|(~m[385]&m[386]&~m[387]&~m[388]&~m[417])|(~m[385]&~m[386]&m[387]&~m[388]&~m[417])|(m[385]&m[386]&~m[387]&m[388]&~m[417])|(m[385]&~m[386]&m[387]&m[388]&~m[417])|(~m[385]&m[386]&m[387]&m[388]&~m[417]))&BiasedRNG[252])|(((m[385]&~m[386]&~m[387]&~m[388]&m[417])|(~m[385]&m[386]&~m[387]&~m[388]&m[417])|(~m[385]&~m[386]&m[387]&~m[388]&m[417])|(m[385]&m[386]&~m[387]&m[388]&m[417])|(m[385]&~m[386]&m[387]&m[388]&m[417])|(~m[385]&m[386]&m[387]&m[388]&m[417]))&~BiasedRNG[252])|((m[385]&m[386]&~m[387]&~m[388]&~m[417])|(m[385]&~m[386]&m[387]&~m[388]&~m[417])|(~m[385]&m[386]&m[387]&~m[388]&~m[417])|(m[385]&m[386]&m[387]&~m[388]&~m[417])|(m[385]&m[386]&m[387]&m[388]&~m[417])|(m[385]&m[386]&~m[387]&~m[388]&m[417])|(m[385]&~m[386]&m[387]&~m[388]&m[417])|(~m[385]&m[386]&m[387]&~m[388]&m[417])|(m[385]&m[386]&m[387]&~m[388]&m[417])|(m[385]&m[386]&m[387]&m[388]&m[417]));
    m[394] = (((m[390]&~m[391]&~m[392]&~m[393]&~m[422])|(~m[390]&m[391]&~m[392]&~m[393]&~m[422])|(~m[390]&~m[391]&m[392]&~m[393]&~m[422])|(m[390]&m[391]&~m[392]&m[393]&~m[422])|(m[390]&~m[391]&m[392]&m[393]&~m[422])|(~m[390]&m[391]&m[392]&m[393]&~m[422]))&BiasedRNG[253])|(((m[390]&~m[391]&~m[392]&~m[393]&m[422])|(~m[390]&m[391]&~m[392]&~m[393]&m[422])|(~m[390]&~m[391]&m[392]&~m[393]&m[422])|(m[390]&m[391]&~m[392]&m[393]&m[422])|(m[390]&~m[391]&m[392]&m[393]&m[422])|(~m[390]&m[391]&m[392]&m[393]&m[422]))&~BiasedRNG[253])|((m[390]&m[391]&~m[392]&~m[393]&~m[422])|(m[390]&~m[391]&m[392]&~m[393]&~m[422])|(~m[390]&m[391]&m[392]&~m[393]&~m[422])|(m[390]&m[391]&m[392]&~m[393]&~m[422])|(m[390]&m[391]&m[392]&m[393]&~m[422])|(m[390]&m[391]&~m[392]&~m[393]&m[422])|(m[390]&~m[391]&m[392]&~m[393]&m[422])|(~m[390]&m[391]&m[392]&~m[393]&m[422])|(m[390]&m[391]&m[392]&~m[393]&m[422])|(m[390]&m[391]&m[392]&m[393]&m[422]));
    m[399] = (((m[395]&~m[396]&~m[397]&~m[398]&~m[427])|(~m[395]&m[396]&~m[397]&~m[398]&~m[427])|(~m[395]&~m[396]&m[397]&~m[398]&~m[427])|(m[395]&m[396]&~m[397]&m[398]&~m[427])|(m[395]&~m[396]&m[397]&m[398]&~m[427])|(~m[395]&m[396]&m[397]&m[398]&~m[427]))&BiasedRNG[254])|(((m[395]&~m[396]&~m[397]&~m[398]&m[427])|(~m[395]&m[396]&~m[397]&~m[398]&m[427])|(~m[395]&~m[396]&m[397]&~m[398]&m[427])|(m[395]&m[396]&~m[397]&m[398]&m[427])|(m[395]&~m[396]&m[397]&m[398]&m[427])|(~m[395]&m[396]&m[397]&m[398]&m[427]))&~BiasedRNG[254])|((m[395]&m[396]&~m[397]&~m[398]&~m[427])|(m[395]&~m[396]&m[397]&~m[398]&~m[427])|(~m[395]&m[396]&m[397]&~m[398]&~m[427])|(m[395]&m[396]&m[397]&~m[398]&~m[427])|(m[395]&m[396]&m[397]&m[398]&~m[427])|(m[395]&m[396]&~m[397]&~m[398]&m[427])|(m[395]&~m[396]&m[397]&~m[398]&m[427])|(~m[395]&m[396]&m[397]&~m[398]&m[427])|(m[395]&m[396]&m[397]&~m[398]&m[427])|(m[395]&m[396]&m[397]&m[398]&m[427]));
    m[404] = (((m[400]&~m[401]&~m[402]&~m[403]&~m[432])|(~m[400]&m[401]&~m[402]&~m[403]&~m[432])|(~m[400]&~m[401]&m[402]&~m[403]&~m[432])|(m[400]&m[401]&~m[402]&m[403]&~m[432])|(m[400]&~m[401]&m[402]&m[403]&~m[432])|(~m[400]&m[401]&m[402]&m[403]&~m[432]))&BiasedRNG[255])|(((m[400]&~m[401]&~m[402]&~m[403]&m[432])|(~m[400]&m[401]&~m[402]&~m[403]&m[432])|(~m[400]&~m[401]&m[402]&~m[403]&m[432])|(m[400]&m[401]&~m[402]&m[403]&m[432])|(m[400]&~m[401]&m[402]&m[403]&m[432])|(~m[400]&m[401]&m[402]&m[403]&m[432]))&~BiasedRNG[255])|((m[400]&m[401]&~m[402]&~m[403]&~m[432])|(m[400]&~m[401]&m[402]&~m[403]&~m[432])|(~m[400]&m[401]&m[402]&~m[403]&~m[432])|(m[400]&m[401]&m[402]&~m[403]&~m[432])|(m[400]&m[401]&m[402]&m[403]&~m[432])|(m[400]&m[401]&~m[402]&~m[403]&m[432])|(m[400]&~m[401]&m[402]&~m[403]&m[432])|(~m[400]&m[401]&m[402]&~m[403]&m[432])|(m[400]&m[401]&m[402]&~m[403]&m[432])|(m[400]&m[401]&m[402]&m[403]&m[432]));
    m[409] = (((m[405]&~m[406]&~m[407]&~m[408]&~m[437])|(~m[405]&m[406]&~m[407]&~m[408]&~m[437])|(~m[405]&~m[406]&m[407]&~m[408]&~m[437])|(m[405]&m[406]&~m[407]&m[408]&~m[437])|(m[405]&~m[406]&m[407]&m[408]&~m[437])|(~m[405]&m[406]&m[407]&m[408]&~m[437]))&BiasedRNG[256])|(((m[405]&~m[406]&~m[407]&~m[408]&m[437])|(~m[405]&m[406]&~m[407]&~m[408]&m[437])|(~m[405]&~m[406]&m[407]&~m[408]&m[437])|(m[405]&m[406]&~m[407]&m[408]&m[437])|(m[405]&~m[406]&m[407]&m[408]&m[437])|(~m[405]&m[406]&m[407]&m[408]&m[437]))&~BiasedRNG[256])|((m[405]&m[406]&~m[407]&~m[408]&~m[437])|(m[405]&~m[406]&m[407]&~m[408]&~m[437])|(~m[405]&m[406]&m[407]&~m[408]&~m[437])|(m[405]&m[406]&m[407]&~m[408]&~m[437])|(m[405]&m[406]&m[407]&m[408]&~m[437])|(m[405]&m[406]&~m[407]&~m[408]&m[437])|(m[405]&~m[406]&m[407]&~m[408]&m[437])|(~m[405]&m[406]&m[407]&~m[408]&m[437])|(m[405]&m[406]&m[407]&~m[408]&m[437])|(m[405]&m[406]&m[407]&m[408]&m[437]));
    m[414] = (((m[410]&~m[411]&~m[412]&~m[413]&~m[442])|(~m[410]&m[411]&~m[412]&~m[413]&~m[442])|(~m[410]&~m[411]&m[412]&~m[413]&~m[442])|(m[410]&m[411]&~m[412]&m[413]&~m[442])|(m[410]&~m[411]&m[412]&m[413]&~m[442])|(~m[410]&m[411]&m[412]&m[413]&~m[442]))&BiasedRNG[257])|(((m[410]&~m[411]&~m[412]&~m[413]&m[442])|(~m[410]&m[411]&~m[412]&~m[413]&m[442])|(~m[410]&~m[411]&m[412]&~m[413]&m[442])|(m[410]&m[411]&~m[412]&m[413]&m[442])|(m[410]&~m[411]&m[412]&m[413]&m[442])|(~m[410]&m[411]&m[412]&m[413]&m[442]))&~BiasedRNG[257])|((m[410]&m[411]&~m[412]&~m[413]&~m[442])|(m[410]&~m[411]&m[412]&~m[413]&~m[442])|(~m[410]&m[411]&m[412]&~m[413]&~m[442])|(m[410]&m[411]&m[412]&~m[413]&~m[442])|(m[410]&m[411]&m[412]&m[413]&~m[442])|(m[410]&m[411]&~m[412]&~m[413]&m[442])|(m[410]&~m[411]&m[412]&~m[413]&m[442])|(~m[410]&m[411]&m[412]&~m[413]&m[442])|(m[410]&m[411]&m[412]&~m[413]&m[442])|(m[410]&m[411]&m[412]&m[413]&m[442]));
    m[419] = (((m[415]&~m[416]&~m[417]&~m[418]&~m[445])|(~m[415]&m[416]&~m[417]&~m[418]&~m[445])|(~m[415]&~m[416]&m[417]&~m[418]&~m[445])|(m[415]&m[416]&~m[417]&m[418]&~m[445])|(m[415]&~m[416]&m[417]&m[418]&~m[445])|(~m[415]&m[416]&m[417]&m[418]&~m[445]))&BiasedRNG[258])|(((m[415]&~m[416]&~m[417]&~m[418]&m[445])|(~m[415]&m[416]&~m[417]&~m[418]&m[445])|(~m[415]&~m[416]&m[417]&~m[418]&m[445])|(m[415]&m[416]&~m[417]&m[418]&m[445])|(m[415]&~m[416]&m[417]&m[418]&m[445])|(~m[415]&m[416]&m[417]&m[418]&m[445]))&~BiasedRNG[258])|((m[415]&m[416]&~m[417]&~m[418]&~m[445])|(m[415]&~m[416]&m[417]&~m[418]&~m[445])|(~m[415]&m[416]&m[417]&~m[418]&~m[445])|(m[415]&m[416]&m[417]&~m[418]&~m[445])|(m[415]&m[416]&m[417]&m[418]&~m[445])|(m[415]&m[416]&~m[417]&~m[418]&m[445])|(m[415]&~m[416]&m[417]&~m[418]&m[445])|(~m[415]&m[416]&m[417]&~m[418]&m[445])|(m[415]&m[416]&m[417]&~m[418]&m[445])|(m[415]&m[416]&m[417]&m[418]&m[445]));
    m[424] = (((m[420]&~m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&m[421]&~m[422]&~m[423]&~m[447])|(~m[420]&~m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&~m[422]&m[423]&~m[447])|(m[420]&~m[421]&m[422]&m[423]&~m[447])|(~m[420]&m[421]&m[422]&m[423]&~m[447]))&BiasedRNG[259])|(((m[420]&~m[421]&~m[422]&~m[423]&m[447])|(~m[420]&m[421]&~m[422]&~m[423]&m[447])|(~m[420]&~m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&~m[422]&m[423]&m[447])|(m[420]&~m[421]&m[422]&m[423]&m[447])|(~m[420]&m[421]&m[422]&m[423]&m[447]))&~BiasedRNG[259])|((m[420]&m[421]&~m[422]&~m[423]&~m[447])|(m[420]&~m[421]&m[422]&~m[423]&~m[447])|(~m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&~m[423]&~m[447])|(m[420]&m[421]&m[422]&m[423]&~m[447])|(m[420]&m[421]&~m[422]&~m[423]&m[447])|(m[420]&~m[421]&m[422]&~m[423]&m[447])|(~m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&~m[423]&m[447])|(m[420]&m[421]&m[422]&m[423]&m[447]));
    m[429] = (((m[425]&~m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&m[426]&~m[427]&~m[428]&~m[452])|(~m[425]&~m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&~m[427]&m[428]&~m[452])|(m[425]&~m[426]&m[427]&m[428]&~m[452])|(~m[425]&m[426]&m[427]&m[428]&~m[452]))&BiasedRNG[260])|(((m[425]&~m[426]&~m[427]&~m[428]&m[452])|(~m[425]&m[426]&~m[427]&~m[428]&m[452])|(~m[425]&~m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&~m[427]&m[428]&m[452])|(m[425]&~m[426]&m[427]&m[428]&m[452])|(~m[425]&m[426]&m[427]&m[428]&m[452]))&~BiasedRNG[260])|((m[425]&m[426]&~m[427]&~m[428]&~m[452])|(m[425]&~m[426]&m[427]&~m[428]&~m[452])|(~m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&~m[428]&~m[452])|(m[425]&m[426]&m[427]&m[428]&~m[452])|(m[425]&m[426]&~m[427]&~m[428]&m[452])|(m[425]&~m[426]&m[427]&~m[428]&m[452])|(~m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&~m[428]&m[452])|(m[425]&m[426]&m[427]&m[428]&m[452]));
    m[434] = (((m[430]&~m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&m[431]&~m[432]&~m[433]&~m[457])|(~m[430]&~m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&~m[432]&m[433]&~m[457])|(m[430]&~m[431]&m[432]&m[433]&~m[457])|(~m[430]&m[431]&m[432]&m[433]&~m[457]))&BiasedRNG[261])|(((m[430]&~m[431]&~m[432]&~m[433]&m[457])|(~m[430]&m[431]&~m[432]&~m[433]&m[457])|(~m[430]&~m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&~m[432]&m[433]&m[457])|(m[430]&~m[431]&m[432]&m[433]&m[457])|(~m[430]&m[431]&m[432]&m[433]&m[457]))&~BiasedRNG[261])|((m[430]&m[431]&~m[432]&~m[433]&~m[457])|(m[430]&~m[431]&m[432]&~m[433]&~m[457])|(~m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&~m[433]&~m[457])|(m[430]&m[431]&m[432]&m[433]&~m[457])|(m[430]&m[431]&~m[432]&~m[433]&m[457])|(m[430]&~m[431]&m[432]&~m[433]&m[457])|(~m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&~m[433]&m[457])|(m[430]&m[431]&m[432]&m[433]&m[457]));
    m[439] = (((m[435]&~m[436]&~m[437]&~m[438]&~m[462])|(~m[435]&m[436]&~m[437]&~m[438]&~m[462])|(~m[435]&~m[436]&m[437]&~m[438]&~m[462])|(m[435]&m[436]&~m[437]&m[438]&~m[462])|(m[435]&~m[436]&m[437]&m[438]&~m[462])|(~m[435]&m[436]&m[437]&m[438]&~m[462]))&BiasedRNG[262])|(((m[435]&~m[436]&~m[437]&~m[438]&m[462])|(~m[435]&m[436]&~m[437]&~m[438]&m[462])|(~m[435]&~m[436]&m[437]&~m[438]&m[462])|(m[435]&m[436]&~m[437]&m[438]&m[462])|(m[435]&~m[436]&m[437]&m[438]&m[462])|(~m[435]&m[436]&m[437]&m[438]&m[462]))&~BiasedRNG[262])|((m[435]&m[436]&~m[437]&~m[438]&~m[462])|(m[435]&~m[436]&m[437]&~m[438]&~m[462])|(~m[435]&m[436]&m[437]&~m[438]&~m[462])|(m[435]&m[436]&m[437]&~m[438]&~m[462])|(m[435]&m[436]&m[437]&m[438]&~m[462])|(m[435]&m[436]&~m[437]&~m[438]&m[462])|(m[435]&~m[436]&m[437]&~m[438]&m[462])|(~m[435]&m[436]&m[437]&~m[438]&m[462])|(m[435]&m[436]&m[437]&~m[438]&m[462])|(m[435]&m[436]&m[437]&m[438]&m[462]));
    m[444] = (((m[440]&~m[441]&~m[442]&~m[443]&~m[467])|(~m[440]&m[441]&~m[442]&~m[443]&~m[467])|(~m[440]&~m[441]&m[442]&~m[443]&~m[467])|(m[440]&m[441]&~m[442]&m[443]&~m[467])|(m[440]&~m[441]&m[442]&m[443]&~m[467])|(~m[440]&m[441]&m[442]&m[443]&~m[467]))&BiasedRNG[263])|(((m[440]&~m[441]&~m[442]&~m[443]&m[467])|(~m[440]&m[441]&~m[442]&~m[443]&m[467])|(~m[440]&~m[441]&m[442]&~m[443]&m[467])|(m[440]&m[441]&~m[442]&m[443]&m[467])|(m[440]&~m[441]&m[442]&m[443]&m[467])|(~m[440]&m[441]&m[442]&m[443]&m[467]))&~BiasedRNG[263])|((m[440]&m[441]&~m[442]&~m[443]&~m[467])|(m[440]&~m[441]&m[442]&~m[443]&~m[467])|(~m[440]&m[441]&m[442]&~m[443]&~m[467])|(m[440]&m[441]&m[442]&~m[443]&~m[467])|(m[440]&m[441]&m[442]&m[443]&~m[467])|(m[440]&m[441]&~m[442]&~m[443]&m[467])|(m[440]&~m[441]&m[442]&~m[443]&m[467])|(~m[440]&m[441]&m[442]&~m[443]&m[467])|(m[440]&m[441]&m[442]&~m[443]&m[467])|(m[440]&m[441]&m[442]&m[443]&m[467]));
    m[449] = (((m[445]&~m[446]&~m[447]&~m[448]&~m[470])|(~m[445]&m[446]&~m[447]&~m[448]&~m[470])|(~m[445]&~m[446]&m[447]&~m[448]&~m[470])|(m[445]&m[446]&~m[447]&m[448]&~m[470])|(m[445]&~m[446]&m[447]&m[448]&~m[470])|(~m[445]&m[446]&m[447]&m[448]&~m[470]))&BiasedRNG[264])|(((m[445]&~m[446]&~m[447]&~m[448]&m[470])|(~m[445]&m[446]&~m[447]&~m[448]&m[470])|(~m[445]&~m[446]&m[447]&~m[448]&m[470])|(m[445]&m[446]&~m[447]&m[448]&m[470])|(m[445]&~m[446]&m[447]&m[448]&m[470])|(~m[445]&m[446]&m[447]&m[448]&m[470]))&~BiasedRNG[264])|((m[445]&m[446]&~m[447]&~m[448]&~m[470])|(m[445]&~m[446]&m[447]&~m[448]&~m[470])|(~m[445]&m[446]&m[447]&~m[448]&~m[470])|(m[445]&m[446]&m[447]&~m[448]&~m[470])|(m[445]&m[446]&m[447]&m[448]&~m[470])|(m[445]&m[446]&~m[447]&~m[448]&m[470])|(m[445]&~m[446]&m[447]&~m[448]&m[470])|(~m[445]&m[446]&m[447]&~m[448]&m[470])|(m[445]&m[446]&m[447]&~m[448]&m[470])|(m[445]&m[446]&m[447]&m[448]&m[470]));
    m[454] = (((m[450]&~m[451]&~m[452]&~m[453]&~m[472])|(~m[450]&m[451]&~m[452]&~m[453]&~m[472])|(~m[450]&~m[451]&m[452]&~m[453]&~m[472])|(m[450]&m[451]&~m[452]&m[453]&~m[472])|(m[450]&~m[451]&m[452]&m[453]&~m[472])|(~m[450]&m[451]&m[452]&m[453]&~m[472]))&BiasedRNG[265])|(((m[450]&~m[451]&~m[452]&~m[453]&m[472])|(~m[450]&m[451]&~m[452]&~m[453]&m[472])|(~m[450]&~m[451]&m[452]&~m[453]&m[472])|(m[450]&m[451]&~m[452]&m[453]&m[472])|(m[450]&~m[451]&m[452]&m[453]&m[472])|(~m[450]&m[451]&m[452]&m[453]&m[472]))&~BiasedRNG[265])|((m[450]&m[451]&~m[452]&~m[453]&~m[472])|(m[450]&~m[451]&m[452]&~m[453]&~m[472])|(~m[450]&m[451]&m[452]&~m[453]&~m[472])|(m[450]&m[451]&m[452]&~m[453]&~m[472])|(m[450]&m[451]&m[452]&m[453]&~m[472])|(m[450]&m[451]&~m[452]&~m[453]&m[472])|(m[450]&~m[451]&m[452]&~m[453]&m[472])|(~m[450]&m[451]&m[452]&~m[453]&m[472])|(m[450]&m[451]&m[452]&~m[453]&m[472])|(m[450]&m[451]&m[452]&m[453]&m[472]));
    m[459] = (((m[455]&~m[456]&~m[457]&~m[458]&~m[477])|(~m[455]&m[456]&~m[457]&~m[458]&~m[477])|(~m[455]&~m[456]&m[457]&~m[458]&~m[477])|(m[455]&m[456]&~m[457]&m[458]&~m[477])|(m[455]&~m[456]&m[457]&m[458]&~m[477])|(~m[455]&m[456]&m[457]&m[458]&~m[477]))&BiasedRNG[266])|(((m[455]&~m[456]&~m[457]&~m[458]&m[477])|(~m[455]&m[456]&~m[457]&~m[458]&m[477])|(~m[455]&~m[456]&m[457]&~m[458]&m[477])|(m[455]&m[456]&~m[457]&m[458]&m[477])|(m[455]&~m[456]&m[457]&m[458]&m[477])|(~m[455]&m[456]&m[457]&m[458]&m[477]))&~BiasedRNG[266])|((m[455]&m[456]&~m[457]&~m[458]&~m[477])|(m[455]&~m[456]&m[457]&~m[458]&~m[477])|(~m[455]&m[456]&m[457]&~m[458]&~m[477])|(m[455]&m[456]&m[457]&~m[458]&~m[477])|(m[455]&m[456]&m[457]&m[458]&~m[477])|(m[455]&m[456]&~m[457]&~m[458]&m[477])|(m[455]&~m[456]&m[457]&~m[458]&m[477])|(~m[455]&m[456]&m[457]&~m[458]&m[477])|(m[455]&m[456]&m[457]&~m[458]&m[477])|(m[455]&m[456]&m[457]&m[458]&m[477]));
    m[464] = (((m[460]&~m[461]&~m[462]&~m[463]&~m[482])|(~m[460]&m[461]&~m[462]&~m[463]&~m[482])|(~m[460]&~m[461]&m[462]&~m[463]&~m[482])|(m[460]&m[461]&~m[462]&m[463]&~m[482])|(m[460]&~m[461]&m[462]&m[463]&~m[482])|(~m[460]&m[461]&m[462]&m[463]&~m[482]))&BiasedRNG[267])|(((m[460]&~m[461]&~m[462]&~m[463]&m[482])|(~m[460]&m[461]&~m[462]&~m[463]&m[482])|(~m[460]&~m[461]&m[462]&~m[463]&m[482])|(m[460]&m[461]&~m[462]&m[463]&m[482])|(m[460]&~m[461]&m[462]&m[463]&m[482])|(~m[460]&m[461]&m[462]&m[463]&m[482]))&~BiasedRNG[267])|((m[460]&m[461]&~m[462]&~m[463]&~m[482])|(m[460]&~m[461]&m[462]&~m[463]&~m[482])|(~m[460]&m[461]&m[462]&~m[463]&~m[482])|(m[460]&m[461]&m[462]&~m[463]&~m[482])|(m[460]&m[461]&m[462]&m[463]&~m[482])|(m[460]&m[461]&~m[462]&~m[463]&m[482])|(m[460]&~m[461]&m[462]&~m[463]&m[482])|(~m[460]&m[461]&m[462]&~m[463]&m[482])|(m[460]&m[461]&m[462]&~m[463]&m[482])|(m[460]&m[461]&m[462]&m[463]&m[482]));
    m[469] = (((m[465]&~m[466]&~m[467]&~m[468]&~m[487])|(~m[465]&m[466]&~m[467]&~m[468]&~m[487])|(~m[465]&~m[466]&m[467]&~m[468]&~m[487])|(m[465]&m[466]&~m[467]&m[468]&~m[487])|(m[465]&~m[466]&m[467]&m[468]&~m[487])|(~m[465]&m[466]&m[467]&m[468]&~m[487]))&BiasedRNG[268])|(((m[465]&~m[466]&~m[467]&~m[468]&m[487])|(~m[465]&m[466]&~m[467]&~m[468]&m[487])|(~m[465]&~m[466]&m[467]&~m[468]&m[487])|(m[465]&m[466]&~m[467]&m[468]&m[487])|(m[465]&~m[466]&m[467]&m[468]&m[487])|(~m[465]&m[466]&m[467]&m[468]&m[487]))&~BiasedRNG[268])|((m[465]&m[466]&~m[467]&~m[468]&~m[487])|(m[465]&~m[466]&m[467]&~m[468]&~m[487])|(~m[465]&m[466]&m[467]&~m[468]&~m[487])|(m[465]&m[466]&m[467]&~m[468]&~m[487])|(m[465]&m[466]&m[467]&m[468]&~m[487])|(m[465]&m[466]&~m[467]&~m[468]&m[487])|(m[465]&~m[466]&m[467]&~m[468]&m[487])|(~m[465]&m[466]&m[467]&~m[468]&m[487])|(m[465]&m[466]&m[467]&~m[468]&m[487])|(m[465]&m[466]&m[467]&m[468]&m[487]));
    m[474] = (((m[470]&~m[471]&~m[472]&~m[473]&~m[490])|(~m[470]&m[471]&~m[472]&~m[473]&~m[490])|(~m[470]&~m[471]&m[472]&~m[473]&~m[490])|(m[470]&m[471]&~m[472]&m[473]&~m[490])|(m[470]&~m[471]&m[472]&m[473]&~m[490])|(~m[470]&m[471]&m[472]&m[473]&~m[490]))&BiasedRNG[269])|(((m[470]&~m[471]&~m[472]&~m[473]&m[490])|(~m[470]&m[471]&~m[472]&~m[473]&m[490])|(~m[470]&~m[471]&m[472]&~m[473]&m[490])|(m[470]&m[471]&~m[472]&m[473]&m[490])|(m[470]&~m[471]&m[472]&m[473]&m[490])|(~m[470]&m[471]&m[472]&m[473]&m[490]))&~BiasedRNG[269])|((m[470]&m[471]&~m[472]&~m[473]&~m[490])|(m[470]&~m[471]&m[472]&~m[473]&~m[490])|(~m[470]&m[471]&m[472]&~m[473]&~m[490])|(m[470]&m[471]&m[472]&~m[473]&~m[490])|(m[470]&m[471]&m[472]&m[473]&~m[490])|(m[470]&m[471]&~m[472]&~m[473]&m[490])|(m[470]&~m[471]&m[472]&~m[473]&m[490])|(~m[470]&m[471]&m[472]&~m[473]&m[490])|(m[470]&m[471]&m[472]&~m[473]&m[490])|(m[470]&m[471]&m[472]&m[473]&m[490]));
    m[479] = (((m[475]&~m[476]&~m[477]&~m[478]&~m[492])|(~m[475]&m[476]&~m[477]&~m[478]&~m[492])|(~m[475]&~m[476]&m[477]&~m[478]&~m[492])|(m[475]&m[476]&~m[477]&m[478]&~m[492])|(m[475]&~m[476]&m[477]&m[478]&~m[492])|(~m[475]&m[476]&m[477]&m[478]&~m[492]))&BiasedRNG[270])|(((m[475]&~m[476]&~m[477]&~m[478]&m[492])|(~m[475]&m[476]&~m[477]&~m[478]&m[492])|(~m[475]&~m[476]&m[477]&~m[478]&m[492])|(m[475]&m[476]&~m[477]&m[478]&m[492])|(m[475]&~m[476]&m[477]&m[478]&m[492])|(~m[475]&m[476]&m[477]&m[478]&m[492]))&~BiasedRNG[270])|((m[475]&m[476]&~m[477]&~m[478]&~m[492])|(m[475]&~m[476]&m[477]&~m[478]&~m[492])|(~m[475]&m[476]&m[477]&~m[478]&~m[492])|(m[475]&m[476]&m[477]&~m[478]&~m[492])|(m[475]&m[476]&m[477]&m[478]&~m[492])|(m[475]&m[476]&~m[477]&~m[478]&m[492])|(m[475]&~m[476]&m[477]&~m[478]&m[492])|(~m[475]&m[476]&m[477]&~m[478]&m[492])|(m[475]&m[476]&m[477]&~m[478]&m[492])|(m[475]&m[476]&m[477]&m[478]&m[492]));
    m[484] = (((m[480]&~m[481]&~m[482]&~m[483]&~m[497])|(~m[480]&m[481]&~m[482]&~m[483]&~m[497])|(~m[480]&~m[481]&m[482]&~m[483]&~m[497])|(m[480]&m[481]&~m[482]&m[483]&~m[497])|(m[480]&~m[481]&m[482]&m[483]&~m[497])|(~m[480]&m[481]&m[482]&m[483]&~m[497]))&BiasedRNG[271])|(((m[480]&~m[481]&~m[482]&~m[483]&m[497])|(~m[480]&m[481]&~m[482]&~m[483]&m[497])|(~m[480]&~m[481]&m[482]&~m[483]&m[497])|(m[480]&m[481]&~m[482]&m[483]&m[497])|(m[480]&~m[481]&m[482]&m[483]&m[497])|(~m[480]&m[481]&m[482]&m[483]&m[497]))&~BiasedRNG[271])|((m[480]&m[481]&~m[482]&~m[483]&~m[497])|(m[480]&~m[481]&m[482]&~m[483]&~m[497])|(~m[480]&m[481]&m[482]&~m[483]&~m[497])|(m[480]&m[481]&m[482]&~m[483]&~m[497])|(m[480]&m[481]&m[482]&m[483]&~m[497])|(m[480]&m[481]&~m[482]&~m[483]&m[497])|(m[480]&~m[481]&m[482]&~m[483]&m[497])|(~m[480]&m[481]&m[482]&~m[483]&m[497])|(m[480]&m[481]&m[482]&~m[483]&m[497])|(m[480]&m[481]&m[482]&m[483]&m[497]));
    m[489] = (((m[485]&~m[486]&~m[487]&~m[488]&~m[502])|(~m[485]&m[486]&~m[487]&~m[488]&~m[502])|(~m[485]&~m[486]&m[487]&~m[488]&~m[502])|(m[485]&m[486]&~m[487]&m[488]&~m[502])|(m[485]&~m[486]&m[487]&m[488]&~m[502])|(~m[485]&m[486]&m[487]&m[488]&~m[502]))&BiasedRNG[272])|(((m[485]&~m[486]&~m[487]&~m[488]&m[502])|(~m[485]&m[486]&~m[487]&~m[488]&m[502])|(~m[485]&~m[486]&m[487]&~m[488]&m[502])|(m[485]&m[486]&~m[487]&m[488]&m[502])|(m[485]&~m[486]&m[487]&m[488]&m[502])|(~m[485]&m[486]&m[487]&m[488]&m[502]))&~BiasedRNG[272])|((m[485]&m[486]&~m[487]&~m[488]&~m[502])|(m[485]&~m[486]&m[487]&~m[488]&~m[502])|(~m[485]&m[486]&m[487]&~m[488]&~m[502])|(m[485]&m[486]&m[487]&~m[488]&~m[502])|(m[485]&m[486]&m[487]&m[488]&~m[502])|(m[485]&m[486]&~m[487]&~m[488]&m[502])|(m[485]&~m[486]&m[487]&~m[488]&m[502])|(~m[485]&m[486]&m[487]&~m[488]&m[502])|(m[485]&m[486]&m[487]&~m[488]&m[502])|(m[485]&m[486]&m[487]&m[488]&m[502]));
    m[494] = (((m[490]&~m[491]&~m[492]&~m[493]&~m[505])|(~m[490]&m[491]&~m[492]&~m[493]&~m[505])|(~m[490]&~m[491]&m[492]&~m[493]&~m[505])|(m[490]&m[491]&~m[492]&m[493]&~m[505])|(m[490]&~m[491]&m[492]&m[493]&~m[505])|(~m[490]&m[491]&m[492]&m[493]&~m[505]))&BiasedRNG[273])|(((m[490]&~m[491]&~m[492]&~m[493]&m[505])|(~m[490]&m[491]&~m[492]&~m[493]&m[505])|(~m[490]&~m[491]&m[492]&~m[493]&m[505])|(m[490]&m[491]&~m[492]&m[493]&m[505])|(m[490]&~m[491]&m[492]&m[493]&m[505])|(~m[490]&m[491]&m[492]&m[493]&m[505]))&~BiasedRNG[273])|((m[490]&m[491]&~m[492]&~m[493]&~m[505])|(m[490]&~m[491]&m[492]&~m[493]&~m[505])|(~m[490]&m[491]&m[492]&~m[493]&~m[505])|(m[490]&m[491]&m[492]&~m[493]&~m[505])|(m[490]&m[491]&m[492]&m[493]&~m[505])|(m[490]&m[491]&~m[492]&~m[493]&m[505])|(m[490]&~m[491]&m[492]&~m[493]&m[505])|(~m[490]&m[491]&m[492]&~m[493]&m[505])|(m[490]&m[491]&m[492]&~m[493]&m[505])|(m[490]&m[491]&m[492]&m[493]&m[505]));
    m[499] = (((m[495]&~m[496]&~m[497]&~m[498]&~m[507])|(~m[495]&m[496]&~m[497]&~m[498]&~m[507])|(~m[495]&~m[496]&m[497]&~m[498]&~m[507])|(m[495]&m[496]&~m[497]&m[498]&~m[507])|(m[495]&~m[496]&m[497]&m[498]&~m[507])|(~m[495]&m[496]&m[497]&m[498]&~m[507]))&BiasedRNG[274])|(((m[495]&~m[496]&~m[497]&~m[498]&m[507])|(~m[495]&m[496]&~m[497]&~m[498]&m[507])|(~m[495]&~m[496]&m[497]&~m[498]&m[507])|(m[495]&m[496]&~m[497]&m[498]&m[507])|(m[495]&~m[496]&m[497]&m[498]&m[507])|(~m[495]&m[496]&m[497]&m[498]&m[507]))&~BiasedRNG[274])|((m[495]&m[496]&~m[497]&~m[498]&~m[507])|(m[495]&~m[496]&m[497]&~m[498]&~m[507])|(~m[495]&m[496]&m[497]&~m[498]&~m[507])|(m[495]&m[496]&m[497]&~m[498]&~m[507])|(m[495]&m[496]&m[497]&m[498]&~m[507])|(m[495]&m[496]&~m[497]&~m[498]&m[507])|(m[495]&~m[496]&m[497]&~m[498]&m[507])|(~m[495]&m[496]&m[497]&~m[498]&m[507])|(m[495]&m[496]&m[497]&~m[498]&m[507])|(m[495]&m[496]&m[497]&m[498]&m[507]));
    m[504] = (((m[500]&~m[501]&~m[502]&~m[503]&~m[512])|(~m[500]&m[501]&~m[502]&~m[503]&~m[512])|(~m[500]&~m[501]&m[502]&~m[503]&~m[512])|(m[500]&m[501]&~m[502]&m[503]&~m[512])|(m[500]&~m[501]&m[502]&m[503]&~m[512])|(~m[500]&m[501]&m[502]&m[503]&~m[512]))&BiasedRNG[275])|(((m[500]&~m[501]&~m[502]&~m[503]&m[512])|(~m[500]&m[501]&~m[502]&~m[503]&m[512])|(~m[500]&~m[501]&m[502]&~m[503]&m[512])|(m[500]&m[501]&~m[502]&m[503]&m[512])|(m[500]&~m[501]&m[502]&m[503]&m[512])|(~m[500]&m[501]&m[502]&m[503]&m[512]))&~BiasedRNG[275])|((m[500]&m[501]&~m[502]&~m[503]&~m[512])|(m[500]&~m[501]&m[502]&~m[503]&~m[512])|(~m[500]&m[501]&m[502]&~m[503]&~m[512])|(m[500]&m[501]&m[502]&~m[503]&~m[512])|(m[500]&m[501]&m[502]&m[503]&~m[512])|(m[500]&m[501]&~m[502]&~m[503]&m[512])|(m[500]&~m[501]&m[502]&~m[503]&m[512])|(~m[500]&m[501]&m[502]&~m[503]&m[512])|(m[500]&m[501]&m[502]&~m[503]&m[512])|(m[500]&m[501]&m[502]&m[503]&m[512]));
    m[509] = (((m[505]&~m[506]&~m[507]&~m[508]&~m[515])|(~m[505]&m[506]&~m[507]&~m[508]&~m[515])|(~m[505]&~m[506]&m[507]&~m[508]&~m[515])|(m[505]&m[506]&~m[507]&m[508]&~m[515])|(m[505]&~m[506]&m[507]&m[508]&~m[515])|(~m[505]&m[506]&m[507]&m[508]&~m[515]))&BiasedRNG[276])|(((m[505]&~m[506]&~m[507]&~m[508]&m[515])|(~m[505]&m[506]&~m[507]&~m[508]&m[515])|(~m[505]&~m[506]&m[507]&~m[508]&m[515])|(m[505]&m[506]&~m[507]&m[508]&m[515])|(m[505]&~m[506]&m[507]&m[508]&m[515])|(~m[505]&m[506]&m[507]&m[508]&m[515]))&~BiasedRNG[276])|((m[505]&m[506]&~m[507]&~m[508]&~m[515])|(m[505]&~m[506]&m[507]&~m[508]&~m[515])|(~m[505]&m[506]&m[507]&~m[508]&~m[515])|(m[505]&m[506]&m[507]&~m[508]&~m[515])|(m[505]&m[506]&m[507]&m[508]&~m[515])|(m[505]&m[506]&~m[507]&~m[508]&m[515])|(m[505]&~m[506]&m[507]&~m[508]&m[515])|(~m[505]&m[506]&m[507]&~m[508]&m[515])|(m[505]&m[506]&m[507]&~m[508]&m[515])|(m[505]&m[506]&m[507]&m[508]&m[515]));
    m[514] = (((m[510]&~m[511]&~m[512]&~m[513]&~m[517])|(~m[510]&m[511]&~m[512]&~m[513]&~m[517])|(~m[510]&~m[511]&m[512]&~m[513]&~m[517])|(m[510]&m[511]&~m[512]&m[513]&~m[517])|(m[510]&~m[511]&m[512]&m[513]&~m[517])|(~m[510]&m[511]&m[512]&m[513]&~m[517]))&BiasedRNG[277])|(((m[510]&~m[511]&~m[512]&~m[513]&m[517])|(~m[510]&m[511]&~m[512]&~m[513]&m[517])|(~m[510]&~m[511]&m[512]&~m[513]&m[517])|(m[510]&m[511]&~m[512]&m[513]&m[517])|(m[510]&~m[511]&m[512]&m[513]&m[517])|(~m[510]&m[511]&m[512]&m[513]&m[517]))&~BiasedRNG[277])|((m[510]&m[511]&~m[512]&~m[513]&~m[517])|(m[510]&~m[511]&m[512]&~m[513]&~m[517])|(~m[510]&m[511]&m[512]&~m[513]&~m[517])|(m[510]&m[511]&m[512]&~m[513]&~m[517])|(m[510]&m[511]&m[512]&m[513]&~m[517])|(m[510]&m[511]&~m[512]&~m[513]&m[517])|(m[510]&~m[511]&m[512]&~m[513]&m[517])|(~m[510]&m[511]&m[512]&~m[513]&m[517])|(m[510]&m[511]&m[512]&~m[513]&m[517])|(m[510]&m[511]&m[512]&m[513]&m[517]));
end

//Update the registered value of RNGs one shifted clock before its needed:
always @(posedge sample_clk) begin
    BiasedRNG[0] = (LFSRcolor0[148]&LFSRcolor0[157]&LFSRcolor0[210]&LFSRcolor0[66]);
    BiasedRNG[1] = (LFSRcolor0[137]&LFSRcolor0[7]&LFSRcolor0[57]&LFSRcolor0[176]);
    BiasedRNG[2] = (LFSRcolor0[152]&LFSRcolor0[135]&LFSRcolor0[88]&LFSRcolor0[299]);
    BiasedRNG[3] = (LFSRcolor0[268]&LFSRcolor0[76]&LFSRcolor0[171]&LFSRcolor0[6]);
    BiasedRNG[4] = (LFSRcolor0[308]&LFSRcolor0[125]&LFSRcolor0[357]&LFSRcolor0[240]);
    BiasedRNG[5] = (LFSRcolor0[146]&LFSRcolor0[204]&LFSRcolor0[134]&LFSRcolor0[366]);
    BiasedRNG[6] = (LFSRcolor0[64]&LFSRcolor0[321]&LFSRcolor0[212]&LFSRcolor0[127]);
    BiasedRNG[7] = (LFSRcolor0[332]&LFSRcolor0[346]&LFSRcolor0[260]&LFSRcolor0[233]);
    BiasedRNG[8] = (LFSRcolor0[274]&LFSRcolor0[87]&LFSRcolor0[360]&LFSRcolor0[323]);
    BiasedRNG[9] = (LFSRcolor0[337]&LFSRcolor0[291]&LFSRcolor0[23]&LFSRcolor0[255]);
    BiasedRNG[10] = (LFSRcolor0[231]&LFSRcolor0[170]&LFSRcolor0[33]&LFSRcolor0[328]);
    BiasedRNG[11] = (LFSRcolor0[197]&LFSRcolor0[201]&LFSRcolor0[191]&LFSRcolor0[249]);
    BiasedRNG[12] = (LFSRcolor0[211]&LFSRcolor0[116]&LFSRcolor0[71]&LFSRcolor0[257]);
    BiasedRNG[13] = (LFSRcolor0[39]&LFSRcolor0[19]&LFSRcolor0[215]&LFSRcolor0[330]);
    BiasedRNG[14] = (LFSRcolor0[235]&LFSRcolor0[98]&LFSRcolor0[142]&LFSRcolor0[27]);
    BiasedRNG[15] = (LFSRcolor0[149]&LFSRcolor0[45]&LFSRcolor0[304]&LFSRcolor0[158]);
    BiasedRNG[16] = (LFSRcolor0[258]&LFSRcolor0[62]&LFSRcolor0[342]&LFSRcolor0[243]);
    BiasedRNG[17] = (LFSRcolor0[77]&LFSRcolor0[95]&LFSRcolor0[109]&LFSRcolor0[266]);
    BiasedRNG[18] = (LFSRcolor0[165]&LFSRcolor0[322]&LFSRcolor0[248]&LFSRcolor0[261]);
    BiasedRNG[19] = (LFSRcolor0[47]&LFSRcolor0[340]&LFSRcolor0[349]&LFSRcolor0[105]);
    BiasedRNG[20] = (LFSRcolor0[297]&LFSRcolor0[24]&LFSRcolor0[208]&LFSRcolor0[173]);
    BiasedRNG[21] = (LFSRcolor0[315]&LFSRcolor0[75]&LFSRcolor0[59]&LFSRcolor0[344]);
    BiasedRNG[22] = (LFSRcolor0[138]&LFSRcolor0[287]&LFSRcolor0[97]&LFSRcolor0[194]);
    BiasedRNG[23] = (LFSRcolor0[167]&LFSRcolor0[151]&LFSRcolor0[254]&LFSRcolor0[162]);
    BiasedRNG[24] = (LFSRcolor0[296]&LFSRcolor0[16]&LFSRcolor0[273]&LFSRcolor0[301]);
    BiasedRNG[25] = (LFSRcolor0[169]&LFSRcolor0[123]&LFSRcolor0[65]&LFSRcolor0[22]);
    BiasedRNG[26] = (LFSRcolor0[367]&LFSRcolor0[292]&LFSRcolor0[300]&LFSRcolor0[5]);
    BiasedRNG[27] = (LFSRcolor0[164]&LFSRcolor0[61]&LFSRcolor0[269]&LFSRcolor0[128]);
    BiasedRNG[28] = (LFSRcolor0[354]&LFSRcolor0[32]&LFSRcolor0[102]&LFSRcolor0[43]);
    BiasedRNG[29] = (LFSRcolor0[285]&LFSRcolor0[316]&LFSRcolor0[154]&LFSRcolor0[0]);
    BiasedRNG[30] = (LFSRcolor0[70]&LFSRcolor0[136]&LFSRcolor0[347]&LFSRcolor0[253]);
    BiasedRNG[31] = (LFSRcolor0[34]&LFSRcolor0[68]&LFSRcolor0[195]&LFSRcolor0[50]);
    BiasedRNG[32] = (LFSRcolor0[294]&LFSRcolor0[153]&LFSRcolor0[60]&LFSRcolor0[21]);
    BiasedRNG[33] = (LFSRcolor0[84]&LFSRcolor0[187]&LFSRcolor0[29]&LFSRcolor0[317]);
    BiasedRNG[34] = (LFSRcolor0[214]&LFSRcolor0[168]&LFSRcolor0[166]&LFSRcolor0[90]);
    BiasedRNG[35] = (LFSRcolor0[227]&LFSRcolor0[126]&LFSRcolor0[241]&LFSRcolor0[236]);
    BiasedRNG[36] = (LFSRcolor0[250]&LFSRcolor0[103]&LFSRcolor0[172]&LFSRcolor0[271]);
    BiasedRNG[37] = (LFSRcolor0[184]&LFSRcolor0[229]&LFSRcolor0[363]&LFSRcolor0[188]);
    BiasedRNG[38] = (LFSRcolor0[139]&LFSRcolor0[55]&LFSRcolor0[264]&LFSRcolor0[107]);
    BiasedRNG[39] = (LFSRcolor0[272]&LFSRcolor0[53]&LFSRcolor0[113]&LFSRcolor0[237]);
    BiasedRNG[40] = (LFSRcolor0[18]&LFSRcolor0[267]&LFSRcolor0[179]&LFSRcolor0[339]);
    BiasedRNG[41] = (LFSRcolor0[155]&LFSRcolor0[49]&LFSRcolor0[336]&LFSRcolor0[12]);
    BiasedRNG[42] = (LFSRcolor0[234]&LFSRcolor0[92]&LFSRcolor0[85]&LFSRcolor0[331]);
    BiasedRNG[43] = (LFSRcolor0[358]&LFSRcolor0[230]&LFSRcolor0[140]&LFSRcolor0[48]);
    BiasedRNG[44] = (LFSRcolor0[40]&LFSRcolor0[15]&LFSRcolor0[198]&LFSRcolor0[101]);
    BiasedRNG[45] = (LFSRcolor0[289]&LFSRcolor0[190]&LFSRcolor0[312]&LFSRcolor0[112]);
    BiasedRNG[46] = (LFSRcolor0[96]&LFSRcolor0[180]&LFSRcolor0[110]&LFSRcolor0[192]);
    BiasedRNG[47] = (LFSRcolor0[20]&LFSRcolor0[334]&LFSRcolor0[51]&LFSRcolor0[44]);
    BiasedRNG[48] = (LFSRcolor0[247]&LFSRcolor0[83]&LFSRcolor0[238]&LFSRcolor0[183]);
    BiasedRNG[49] = (LFSRcolor0[259]&LFSRcolor0[338]&LFSRcolor0[293]&LFSRcolor0[246]);
    BiasedRNG[50] = (LFSRcolor0[262]&LFSRcolor0[228]&LFSRcolor0[277]&LFSRcolor0[120]);
    BiasedRNG[51] = (LFSRcolor0[104]&LFSRcolor0[320]&LFSRcolor0[163]&LFSRcolor0[144]);
    BiasedRNG[52] = (LFSRcolor0[333]&LFSRcolor0[80]&LFSRcolor0[226]&LFSRcolor0[3]);
    BiasedRNG[53] = (LFSRcolor0[161]&LFSRcolor0[220]&LFSRcolor0[41]&LFSRcolor0[122]);
    BiasedRNG[54] = (LFSRcolor0[82]&LFSRcolor0[270]&LFSRcolor0[223]&LFSRcolor0[206]);
    BiasedRNG[55] = (LFSRcolor0[79]&LFSRcolor0[245]&LFSRcolor0[200]&LFSRcolor0[359]);
    BiasedRNG[56] = (LFSRcolor0[58]&LFSRcolor0[251]&LFSRcolor0[324]&LFSRcolor0[78]);
    BiasedRNG[57] = (LFSRcolor0[263]&LFSRcolor0[199]&LFSRcolor0[94]&LFSRcolor0[17]);
    BiasedRNG[58] = (LFSRcolor0[106]&LFSRcolor0[37]&LFSRcolor0[46]&LFSRcolor0[31]);
    BiasedRNG[59] = (LFSRcolor0[91]&LFSRcolor0[302]&LFSRcolor0[219]&LFSRcolor0[265]);
    BiasedRNG[60] = (LFSRcolor0[26]&LFSRcolor0[283]&LFSRcolor0[362]&LFSRcolor0[352]);
    BiasedRNG[61] = (LFSRcolor0[295]&LFSRcolor0[307]&LFSRcolor0[356]&LFSRcolor0[327]);
    BiasedRNG[62] = (LFSRcolor0[117]&LFSRcolor0[203]&LFSRcolor0[114]&LFSRcolor0[326]);
    BiasedRNG[63] = (LFSRcolor0[305]&LFSRcolor0[9]&LFSRcolor0[56]&LFSRcolor0[256]);
    UnbiasedRNG[0] = LFSRcolor0[288];
    UnbiasedRNG[1] = LFSRcolor0[181];
    UnbiasedRNG[2] = LFSRcolor0[14];
    UnbiasedRNG[3] = LFSRcolor0[132];
    UnbiasedRNG[4] = LFSRcolor0[290];
    UnbiasedRNG[5] = LFSRcolor0[209];
    UnbiasedRNG[6] = LFSRcolor0[115];
    UnbiasedRNG[7] = LFSRcolor0[318];
    UnbiasedRNG[8] = LFSRcolor0[244];
    UnbiasedRNG[9] = LFSRcolor0[282];
    UnbiasedRNG[10] = LFSRcolor0[72];
    UnbiasedRNG[11] = LFSRcolor0[310];
    UnbiasedRNG[12] = LFSRcolor0[186];
    UnbiasedRNG[13] = LFSRcolor0[129];
    UnbiasedRNG[14] = LFSRcolor0[232];
    UnbiasedRNG[15] = LFSRcolor0[225];
    UnbiasedRNG[16] = LFSRcolor0[196];
    UnbiasedRNG[17] = LFSRcolor0[11];
    UnbiasedRNG[18] = LFSRcolor0[100];
    UnbiasedRNG[19] = LFSRcolor0[141];
    UnbiasedRNG[20] = LFSRcolor0[239];
    UnbiasedRNG[21] = LFSRcolor0[145];
    UnbiasedRNG[22] = LFSRcolor0[216];
    UnbiasedRNG[23] = LFSRcolor0[311];
    UnbiasedRNG[24] = LFSRcolor0[52];
    UnbiasedRNG[25] = LFSRcolor0[281];
    UnbiasedRNG[26] = LFSRcolor0[364];
    UnbiasedRNG[27] = LFSRcolor0[130];
    UnbiasedRNG[28] = LFSRcolor0[276];
    UnbiasedRNG[29] = LFSRcolor0[361];
    UnbiasedRNG[30] = LFSRcolor0[118];
    UnbiasedRNG[31] = LFSRcolor0[279];
    UnbiasedRNG[32] = LFSRcolor0[86];
    UnbiasedRNG[33] = LFSRcolor0[329];
    UnbiasedRNG[34] = LFSRcolor0[341];
    UnbiasedRNG[35] = LFSRcolor0[36];
    UnbiasedRNG[36] = LFSRcolor0[217];
    UnbiasedRNG[37] = LFSRcolor0[81];
    UnbiasedRNG[38] = LFSRcolor0[242];
    UnbiasedRNG[39] = LFSRcolor0[284];
    UnbiasedRNG[40] = LFSRcolor0[178];
    UnbiasedRNG[41] = LFSRcolor0[353];
    UnbiasedRNG[42] = LFSRcolor0[351];
    UnbiasedRNG[43] = LFSRcolor0[159];
    UnbiasedRNG[44] = LFSRcolor0[174];
    UnbiasedRNG[45] = LFSRcolor0[177];
    UnbiasedRNG[46] = LFSRcolor0[207];
    UnbiasedRNG[47] = LFSRcolor0[124];
    UnbiasedRNG[48] = LFSRcolor0[63];
    UnbiasedRNG[49] = LFSRcolor0[42];
    UnbiasedRNG[50] = LFSRcolor0[4];
    UnbiasedRNG[51] = LFSRcolor0[275];
    UnbiasedRNG[52] = LFSRcolor0[278];
    UnbiasedRNG[53] = LFSRcolor0[67];
    UnbiasedRNG[54] = LFSRcolor0[30];
    UnbiasedRNG[55] = LFSRcolor0[69];
    UnbiasedRNG[56] = LFSRcolor0[286];
    UnbiasedRNG[57] = LFSRcolor0[224];
    UnbiasedRNG[58] = LFSRcolor0[147];
    UnbiasedRNG[59] = LFSRcolor0[343];
    UnbiasedRNG[60] = LFSRcolor0[108];
    UnbiasedRNG[61] = LFSRcolor0[222];
    UnbiasedRNG[62] = LFSRcolor0[185];
    UnbiasedRNG[63] = LFSRcolor0[365];
    UnbiasedRNG[64] = LFSRcolor0[218];
    UnbiasedRNG[65] = LFSRcolor0[313];
    UnbiasedRNG[66] = LFSRcolor0[221];
    UnbiasedRNG[67] = LFSRcolor0[355];
    UnbiasedRNG[68] = LFSRcolor0[111];
    UnbiasedRNG[69] = LFSRcolor0[8];
    UnbiasedRNG[70] = LFSRcolor0[28];
end

always @(posedge color0_clk) begin
    BiasedRNG[64] = (LFSRcolor1[410]&LFSRcolor1[343]&LFSRcolor1[41]&LFSRcolor1[42]);
    BiasedRNG[65] = (LFSRcolor1[215]&LFSRcolor1[161]&LFSRcolor1[332]&LFSRcolor1[288]);
    BiasedRNG[66] = (LFSRcolor1[258]&LFSRcolor1[301]&LFSRcolor1[200]&LFSRcolor1[389]);
    BiasedRNG[67] = (LFSRcolor1[220]&LFSRcolor1[212]&LFSRcolor1[251]&LFSRcolor1[62]);
    BiasedRNG[68] = (LFSRcolor1[394]&LFSRcolor1[276]&LFSRcolor1[79]&LFSRcolor1[299]);
    BiasedRNG[69] = (LFSRcolor1[208]&LFSRcolor1[35]&LFSRcolor1[402]&LFSRcolor1[346]);
    BiasedRNG[70] = (LFSRcolor1[264]&LFSRcolor1[131]&LFSRcolor1[175]&LFSRcolor1[305]);
    BiasedRNG[71] = (LFSRcolor1[67]&LFSRcolor1[45]&LFSRcolor1[368]&LFSRcolor1[164]);
    BiasedRNG[72] = (LFSRcolor1[113]&LFSRcolor1[304]&LFSRcolor1[433]&LFSRcolor1[82]);
    BiasedRNG[73] = (LFSRcolor1[441]&LFSRcolor1[380]&LFSRcolor1[431]&LFSRcolor1[22]);
    BiasedRNG[74] = (LFSRcolor1[125]&LFSRcolor1[330]&LFSRcolor1[140]&LFSRcolor1[255]);
    BiasedRNG[75] = (LFSRcolor1[442]&LFSRcolor1[154]&LFSRcolor1[158]&LFSRcolor1[457]);
    BiasedRNG[76] = (LFSRcolor1[438]&LFSRcolor1[60]&LFSRcolor1[393]&LFSRcolor1[311]);
    BiasedRNG[77] = (LFSRcolor1[138]&LFSRcolor1[53]&LFSRcolor1[443]&LFSRcolor1[253]);
    BiasedRNG[78] = (LFSRcolor1[152]&LFSRcolor1[223]&LFSRcolor1[271]&LFSRcolor1[318]);
    BiasedRNG[79] = (LFSRcolor1[249]&LFSRcolor1[278]&LFSRcolor1[427]&LFSRcolor1[216]);
    BiasedRNG[80] = (LFSRcolor1[214]&LFSRcolor1[183]&LFSRcolor1[219]&LFSRcolor1[172]);
    BiasedRNG[81] = (LFSRcolor1[87]&LFSRcolor1[123]&LFSRcolor1[121]&LFSRcolor1[171]);
    BiasedRNG[82] = (LFSRcolor1[458]&LFSRcolor1[279]&LFSRcolor1[73]&LFSRcolor1[344]);
    BiasedRNG[83] = (LFSRcolor1[50]&LFSRcolor1[241]&LFSRcolor1[282]&LFSRcolor1[358]);
    BiasedRNG[84] = (LFSRcolor1[116]&LFSRcolor1[334]&LFSRcolor1[198]&LFSRcolor1[14]);
    BiasedRNG[85] = (LFSRcolor1[61]&LFSRcolor1[272]&LFSRcolor1[371]&LFSRcolor1[341]);
    BiasedRNG[86] = (LFSRcolor1[89]&LFSRcolor1[379]&LFSRcolor1[303]&LFSRcolor1[376]);
    BiasedRNG[87] = (LFSRcolor1[3]&LFSRcolor1[27]&LFSRcolor1[136]&LFSRcolor1[205]);
    BiasedRNG[88] = (LFSRcolor1[298]&LFSRcolor1[201]&LFSRcolor1[401]&LFSRcolor1[286]);
    BiasedRNG[89] = (LFSRcolor1[197]&LFSRcolor1[254]&LFSRcolor1[246]&LFSRcolor1[235]);
    BiasedRNG[90] = (LFSRcolor1[34]&LFSRcolor1[115]&LFSRcolor1[177]&LFSRcolor1[356]);
    BiasedRNG[91] = (LFSRcolor1[156]&LFSRcolor1[347]&LFSRcolor1[186]&LFSRcolor1[207]);
    BiasedRNG[92] = (LFSRcolor1[385]&LFSRcolor1[367]&LFSRcolor1[147]&LFSRcolor1[193]);
    BiasedRNG[93] = (LFSRcolor1[59]&LFSRcolor1[267]&LFSRcolor1[374]&LFSRcolor1[316]);
    BiasedRNG[94] = (LFSRcolor1[391]&LFSRcolor1[233]&LFSRcolor1[218]&LFSRcolor1[29]);
    BiasedRNG[95] = (LFSRcolor1[132]&LFSRcolor1[65]&LFSRcolor1[155]&LFSRcolor1[144]);
    BiasedRNG[96] = (LFSRcolor1[403]&LFSRcolor1[129]&LFSRcolor1[49]&LFSRcolor1[232]);
    BiasedRNG[97] = (LFSRcolor1[317]&LFSRcolor1[117]&LFSRcolor1[43]&LFSRcolor1[203]);
    BiasedRNG[98] = (LFSRcolor1[323]&LFSRcolor1[238]&LFSRcolor1[151]&LFSRcolor1[99]);
    BiasedRNG[99] = (LFSRcolor1[237]&LFSRcolor1[274]&LFSRcolor1[256]&LFSRcolor1[6]);
    BiasedRNG[100] = (LFSRcolor1[395]&LFSRcolor1[122]&LFSRcolor1[265]&LFSRcolor1[103]);
    BiasedRNG[101] = (LFSRcolor1[39]&LFSRcolor1[64]&LFSRcolor1[292]&LFSRcolor1[135]);
    BiasedRNG[102] = (LFSRcolor1[225]&LFSRcolor1[439]&LFSRcolor1[133]&LFSRcolor1[108]);
    BiasedRNG[103] = (LFSRcolor1[333]&LFSRcolor1[196]&LFSRcolor1[96]&LFSRcolor1[242]);
    BiasedRNG[104] = (LFSRcolor1[437]&LFSRcolor1[114]&LFSRcolor1[70]&LFSRcolor1[357]);
    BiasedRNG[105] = (LFSRcolor1[362]&LFSRcolor1[406]&LFSRcolor1[90]&LFSRcolor1[206]);
    BiasedRNG[106] = (LFSRcolor1[7]&LFSRcolor1[454]&LFSRcolor1[263]&LFSRcolor1[436]);
    BiasedRNG[107] = (LFSRcolor1[310]&LFSRcolor1[210]&LFSRcolor1[157]&LFSRcolor1[243]);
    BiasedRNG[108] = (LFSRcolor1[52]&LFSRcolor1[338]&LFSRcolor1[349]&LFSRcolor1[328]);
    BiasedRNG[109] = (LFSRcolor1[8]&LFSRcolor1[359]&LFSRcolor1[100]&LFSRcolor1[13]);
    BiasedRNG[110] = (LFSRcolor1[363]&LFSRcolor1[409]&LFSRcolor1[153]&LFSRcolor1[425]);
    BiasedRNG[111] = (LFSRcolor1[86]&LFSRcolor1[38]&LFSRcolor1[455]&LFSRcolor1[421]);
    BiasedRNG[112] = (LFSRcolor1[234]&LFSRcolor1[32]&LFSRcolor1[308]&LFSRcolor1[190]);
    BiasedRNG[113] = (LFSRcolor1[199]&LFSRcolor1[163]&LFSRcolor1[295]&LFSRcolor1[174]);
    BiasedRNG[114] = (LFSRcolor1[134]&LFSRcolor1[259]&LFSRcolor1[284]&LFSRcolor1[400]);
    BiasedRNG[115] = (LFSRcolor1[266]&LFSRcolor1[297]&LFSRcolor1[350]&LFSRcolor1[83]);
    BiasedRNG[116] = (LFSRcolor1[54]&LFSRcolor1[18]&LFSRcolor1[168]&LFSRcolor1[10]);
    BiasedRNG[117] = (LFSRcolor1[451]&LFSRcolor1[289]&LFSRcolor1[227]&LFSRcolor1[329]);
    BiasedRNG[118] = (LFSRcolor1[84]&LFSRcolor1[76]&LFSRcolor1[326]&LFSRcolor1[381]);
    BiasedRNG[119] = (LFSRcolor1[187]&LFSRcolor1[137]&LFSRcolor1[105]&LFSRcolor1[104]);
    BiasedRNG[120] = (LFSRcolor1[435]&LFSRcolor1[194]&LFSRcolor1[85]&LFSRcolor1[33]);
    BiasedRNG[121] = (LFSRcolor1[262]&LFSRcolor1[107]&LFSRcolor1[399]&LFSRcolor1[19]);
    BiasedRNG[122] = (LFSRcolor1[98]&LFSRcolor1[360]&LFSRcolor1[300]&LFSRcolor1[51]);
    BiasedRNG[123] = (LFSRcolor1[378]&LFSRcolor1[26]&LFSRcolor1[257]&LFSRcolor1[307]);
    BiasedRNG[124] = (LFSRcolor1[320]&LFSRcolor1[423]&LFSRcolor1[159]&LFSRcolor1[434]);
    BiasedRNG[125] = (LFSRcolor1[324]&LFSRcolor1[250]&LFSRcolor1[74]&LFSRcolor1[63]);
    BiasedRNG[126] = (LFSRcolor1[229]&LFSRcolor1[424]&LFSRcolor1[48]&LFSRcolor1[112]);
    BiasedRNG[127] = (LFSRcolor1[459]&LFSRcolor1[81]&LFSRcolor1[209]&LFSRcolor1[93]);
    BiasedRNG[128] = (LFSRcolor1[31]&LFSRcolor1[327]&LFSRcolor1[407]&LFSRcolor1[179]);
    BiasedRNG[129] = (LFSRcolor1[184]&LFSRcolor1[321]&LFSRcolor1[339]&LFSRcolor1[322]);
    BiasedRNG[130] = (LFSRcolor1[118]&LFSRcolor1[354]&LFSRcolor1[188]&LFSRcolor1[245]);
    BiasedRNG[131] = (LFSRcolor1[335]&LFSRcolor1[432]&LFSRcolor1[240]&LFSRcolor1[4]);
    BiasedRNG[132] = (LFSRcolor1[191]&LFSRcolor1[146]&LFSRcolor1[302]&LFSRcolor1[440]);
    BiasedRNG[133] = (LFSRcolor1[69]&LFSRcolor1[375]&LFSRcolor1[148]&LFSRcolor1[236]);
    BiasedRNG[134] = (LFSRcolor1[287]&LFSRcolor1[77]&LFSRcolor1[384]&LFSRcolor1[72]);
    BiasedRNG[135] = (LFSRcolor1[55]&LFSRcolor1[97]&LFSRcolor1[352]&LFSRcolor1[170]);
    BiasedRNG[136] = (LFSRcolor1[426]&LFSRcolor1[24]&LFSRcolor1[355]&LFSRcolor1[396]);
    BiasedRNG[137] = (LFSRcolor1[370]&LFSRcolor1[75]&LFSRcolor1[12]&LFSRcolor1[110]);
    BiasedRNG[138] = (LFSRcolor1[269]&LFSRcolor1[192]&LFSRcolor1[248]&LFSRcolor1[331]);
    BiasedRNG[139] = (LFSRcolor1[291]&LFSRcolor1[221]&LFSRcolor1[275]&LFSRcolor1[345]);
    BiasedRNG[140] = (LFSRcolor1[173]&LFSRcolor1[351]&LFSRcolor1[340]&LFSRcolor1[15]);
    BiasedRNG[141] = (LFSRcolor1[449]&LFSRcolor1[239]&LFSRcolor1[377]&LFSRcolor1[430]);
    BiasedRNG[142] = (LFSRcolor1[78]&LFSRcolor1[418]&LFSRcolor1[119]&LFSRcolor1[36]);
    BiasedRNG[143] = (LFSRcolor1[169]&LFSRcolor1[181]&LFSRcolor1[270]&LFSRcolor1[260]);
    BiasedRNG[144] = (LFSRcolor1[261]&LFSRcolor1[111]&LFSRcolor1[416]&LFSRcolor1[95]);
    BiasedRNG[145] = (LFSRcolor1[165]&LFSRcolor1[143]&LFSRcolor1[456]&LFSRcolor1[195]);
    BiasedRNG[146] = (LFSRcolor1[386]&LFSRcolor1[353]&LFSRcolor1[180]&LFSRcolor1[16]);
    BiasedRNG[147] = (LFSRcolor1[88]&LFSRcolor1[127]&LFSRcolor1[211]&LFSRcolor1[213]);
    BiasedRNG[148] = (LFSRcolor1[319]&LFSRcolor1[293]&LFSRcolor1[224]&LFSRcolor1[139]);
    BiasedRNG[149] = (LFSRcolor1[160]&LFSRcolor1[387]&LFSRcolor1[417]&LFSRcolor1[25]);
    BiasedRNG[150] = (LFSRcolor1[128]&LFSRcolor1[9]&LFSRcolor1[313]&LFSRcolor1[408]);
    BiasedRNG[151] = (LFSRcolor1[365]&LFSRcolor1[231]&LFSRcolor1[342]&LFSRcolor1[189]);
    BiasedRNG[152] = (LFSRcolor1[142]&LFSRcolor1[404]&LFSRcolor1[281]&LFSRcolor1[80]);
    BiasedRNG[153] = (LFSRcolor1[411]&LFSRcolor1[420]&LFSRcolor1[182]&LFSRcolor1[294]);
    BiasedRNG[154] = (LFSRcolor1[230]&LFSRcolor1[102]&LFSRcolor1[314]&LFSRcolor1[419]);
    BiasedRNG[155] = (LFSRcolor1[222]&LFSRcolor1[68]&LFSRcolor1[452]&LFSRcolor1[30]);
    BiasedRNG[156] = (LFSRcolor1[94]&LFSRcolor1[398]&LFSRcolor1[141]&LFSRcolor1[412]);
    BiasedRNG[157] = (LFSRcolor1[290]&LFSRcolor1[185]&LFSRcolor1[92]&LFSRcolor1[364]);
    BiasedRNG[158] = (LFSRcolor1[247]&LFSRcolor1[306]&LFSRcolor1[178]&LFSRcolor1[20]);
    UnbiasedRNG[71] = LFSRcolor1[149];
    UnbiasedRNG[72] = LFSRcolor1[315];
    UnbiasedRNG[73] = LFSRcolor1[414];
    UnbiasedRNG[74] = LFSRcolor1[283];
    UnbiasedRNG[75] = LFSRcolor1[309];
    UnbiasedRNG[76] = LFSRcolor1[167];
    UnbiasedRNG[77] = LFSRcolor1[21];
    UnbiasedRNG[78] = LFSRcolor1[337];
    UnbiasedRNG[79] = LFSRcolor1[348];
    UnbiasedRNG[80] = LFSRcolor1[273];
    UnbiasedRNG[81] = LFSRcolor1[106];
    UnbiasedRNG[82] = LFSRcolor1[390];
    UnbiasedRNG[83] = LFSRcolor1[268];
    UnbiasedRNG[84] = LFSRcolor1[145];
    UnbiasedRNG[85] = LFSRcolor1[228];
    UnbiasedRNG[86] = LFSRcolor1[150];
    UnbiasedRNG[87] = LFSRcolor1[5];
    UnbiasedRNG[88] = LFSRcolor1[336];
    UnbiasedRNG[89] = LFSRcolor1[382];
    UnbiasedRNG[90] = LFSRcolor1[296];
    UnbiasedRNG[91] = LFSRcolor1[413];
    UnbiasedRNG[92] = LFSRcolor1[450];
    UnbiasedRNG[93] = LFSRcolor1[130];
    UnbiasedRNG[94] = LFSRcolor1[57];
    UnbiasedRNG[95] = LFSRcolor1[166];
    UnbiasedRNG[96] = LFSRcolor1[2];
    UnbiasedRNG[97] = LFSRcolor1[226];
    UnbiasedRNG[98] = LFSRcolor1[217];
    UnbiasedRNG[99] = LFSRcolor1[47];
    UnbiasedRNG[100] = LFSRcolor1[120];
    UnbiasedRNG[101] = LFSRcolor1[17];
    UnbiasedRNG[102] = LFSRcolor1[285];
    UnbiasedRNG[103] = LFSRcolor1[176];
    UnbiasedRNG[104] = LFSRcolor1[397];
    UnbiasedRNG[105] = LFSRcolor1[280];
    UnbiasedRNG[106] = LFSRcolor1[58];
    UnbiasedRNG[107] = LFSRcolor1[448];
    UnbiasedRNG[108] = LFSRcolor1[444];
    UnbiasedRNG[109] = LFSRcolor1[46];
    UnbiasedRNG[110] = LFSRcolor1[388];
    UnbiasedRNG[111] = LFSRcolor1[428];
    UnbiasedRNG[112] = LFSRcolor1[361];
    UnbiasedRNG[113] = LFSRcolor1[202];
    UnbiasedRNG[114] = LFSRcolor1[372];
    UnbiasedRNG[115] = LFSRcolor1[366];
    UnbiasedRNG[116] = LFSRcolor1[28];
    UnbiasedRNG[117] = LFSRcolor1[124];
    UnbiasedRNG[118] = LFSRcolor1[56];
    UnbiasedRNG[119] = LFSRcolor1[405];
end

always @(posedge color1_clk) begin
    BiasedRNG[159] = (LFSRcolor2[161]&LFSRcolor2[94]&LFSRcolor2[26]&LFSRcolor2[236]);
    BiasedRNG[160] = (LFSRcolor2[155]&LFSRcolor2[256]&LFSRcolor2[60]&LFSRcolor2[95]);
    BiasedRNG[161] = (LFSRcolor2[159]&LFSRcolor2[131]&LFSRcolor2[261]&LFSRcolor2[109]);
    BiasedRNG[162] = (LFSRcolor2[183]&LFSRcolor2[137]&LFSRcolor2[118]&LFSRcolor2[186]);
    BiasedRNG[163] = (LFSRcolor2[280]&LFSRcolor2[304]&LFSRcolor2[82]&LFSRcolor2[4]);
    BiasedRNG[164] = (LFSRcolor2[37]&LFSRcolor2[58]&LFSRcolor2[185]&LFSRcolor2[107]);
    BiasedRNG[165] = (LFSRcolor2[285]&LFSRcolor2[264]&LFSRcolor2[105]&LFSRcolor2[213]);
    BiasedRNG[166] = (LFSRcolor2[210]&LFSRcolor2[63]&LFSRcolor2[312]&LFSRcolor2[194]);
    BiasedRNG[167] = (LFSRcolor2[75]&LFSRcolor2[52]&LFSRcolor2[262]&LFSRcolor2[190]);
    BiasedRNG[168] = (LFSRcolor2[1]&LFSRcolor2[54]&LFSRcolor2[86]&LFSRcolor2[253]);
    BiasedRNG[169] = (LFSRcolor2[8]&LFSRcolor2[101]&LFSRcolor2[315]&LFSRcolor2[189]);
    BiasedRNG[170] = (LFSRcolor2[196]&LFSRcolor2[222]&LFSRcolor2[13]&LFSRcolor2[44]);
    BiasedRNG[171] = (LFSRcolor2[188]&LFSRcolor2[65]&LFSRcolor2[59]&LFSRcolor2[15]);
    BiasedRNG[172] = (LFSRcolor2[226]&LFSRcolor2[90]&LFSRcolor2[132]&LFSRcolor2[124]);
    BiasedRNG[173] = (LFSRcolor2[181]&LFSRcolor2[284]&LFSRcolor2[76]&LFSRcolor2[271]);
    BiasedRNG[174] = (LFSRcolor2[249]&LFSRcolor2[127]&LFSRcolor2[64]&LFSRcolor2[53]);
    BiasedRNG[175] = (LFSRcolor2[140]&LFSRcolor2[164]&LFSRcolor2[307]&LFSRcolor2[129]);
    BiasedRNG[176] = (LFSRcolor2[88]&LFSRcolor2[252]&LFSRcolor2[278]&LFSRcolor2[80]);
    BiasedRNG[177] = (LFSRcolor2[51]&LFSRcolor2[250]&LFSRcolor2[247]&LFSRcolor2[23]);
    BiasedRNG[178] = (LFSRcolor2[138]&LFSRcolor2[299]&LFSRcolor2[153]&LFSRcolor2[254]);
    BiasedRNG[179] = (LFSRcolor2[235]&LFSRcolor2[33]&LFSRcolor2[231]&LFSRcolor2[43]);
    BiasedRNG[180] = (LFSRcolor2[106]&LFSRcolor2[176]&LFSRcolor2[120]&LFSRcolor2[108]);
    BiasedRNG[181] = (LFSRcolor2[30]&LFSRcolor2[220]&LFSRcolor2[147]&LFSRcolor2[19]);
    BiasedRNG[182] = (LFSRcolor2[232]&LFSRcolor2[163]&LFSRcolor2[204]&LFSRcolor2[300]);
    BiasedRNG[183] = (LFSRcolor2[289]&LFSRcolor2[263]&LFSRcolor2[303]&LFSRcolor2[22]);
    BiasedRNG[184] = (LFSRcolor2[265]&LFSRcolor2[158]&LFSRcolor2[230]&LFSRcolor2[21]);
    BiasedRNG[185] = (LFSRcolor2[55]&LFSRcolor2[260]&LFSRcolor2[218]&LFSRcolor2[211]);
    BiasedRNG[186] = (LFSRcolor2[184]&LFSRcolor2[170]&LFSRcolor2[84]&LFSRcolor2[255]);
    BiasedRNG[187] = (LFSRcolor2[234]&LFSRcolor2[114]&LFSRcolor2[97]&LFSRcolor2[244]);
    BiasedRNG[188] = (LFSRcolor2[67]&LFSRcolor2[141]&LFSRcolor2[296]&LFSRcolor2[133]);
    BiasedRNG[189] = (LFSRcolor2[116]&LFSRcolor2[45]&LFSRcolor2[245]&LFSRcolor2[273]);
    BiasedRNG[190] = (LFSRcolor2[100]&LFSRcolor2[178]&LFSRcolor2[294]&LFSRcolor2[119]);
    BiasedRNG[191] = (LFSRcolor2[0]&LFSRcolor2[20]&LFSRcolor2[34]&LFSRcolor2[301]);
    BiasedRNG[192] = (LFSRcolor2[279]&LFSRcolor2[206]&LFSRcolor2[156]&LFSRcolor2[12]);
    BiasedRNG[193] = (LFSRcolor2[113]&LFSRcolor2[168]&LFSRcolor2[25]&LFSRcolor2[275]);
    BiasedRNG[194] = (LFSRcolor2[175]&LFSRcolor2[111]&LFSRcolor2[180]&LFSRcolor2[302]);
    BiasedRNG[195] = (LFSRcolor2[251]&LFSRcolor2[126]&LFSRcolor2[229]&LFSRcolor2[172]);
    BiasedRNG[196] = (LFSRcolor2[208]&LFSRcolor2[74]&LFSRcolor2[306]&LFSRcolor2[233]);
    BiasedRNG[197] = (LFSRcolor2[56]&LFSRcolor2[215]&LFSRcolor2[195]&LFSRcolor2[297]);
    BiasedRNG[198] = (LFSRcolor2[154]&LFSRcolor2[121]&LFSRcolor2[32]&LFSRcolor2[203]);
    BiasedRNG[199] = (LFSRcolor2[320]&LFSRcolor2[242]&LFSRcolor2[267]&LFSRcolor2[243]);
    BiasedRNG[200] = (LFSRcolor2[3]&LFSRcolor2[157]&LFSRcolor2[14]&LFSRcolor2[200]);
    BiasedRNG[201] = (LFSRcolor2[290]&LFSRcolor2[179]&LFSRcolor2[202]&LFSRcolor2[217]);
    BiasedRNG[202] = (LFSRcolor2[192]&LFSRcolor2[98]&LFSRcolor2[177]&LFSRcolor2[146]);
    BiasedRNG[203] = (LFSRcolor2[187]&LFSRcolor2[17]&LFSRcolor2[295]&LFSRcolor2[16]);
    BiasedRNG[204] = (LFSRcolor2[221]&LFSRcolor2[216]&LFSRcolor2[123]&LFSRcolor2[42]);
    BiasedRNG[205] = (LFSRcolor2[36]&LFSRcolor2[5]&LFSRcolor2[115]&LFSRcolor2[35]);
    BiasedRNG[206] = (LFSRcolor2[281]&LFSRcolor2[151]&LFSRcolor2[197]&LFSRcolor2[148]);
    BiasedRNG[207] = (LFSRcolor2[7]&LFSRcolor2[167]&LFSRcolor2[292]&LFSRcolor2[135]);
    BiasedRNG[208] = (LFSRcolor2[87]&LFSRcolor2[104]&LFSRcolor2[237]&LFSRcolor2[169]);
    BiasedRNG[209] = (LFSRcolor2[39]&LFSRcolor2[50]&LFSRcolor2[40]&LFSRcolor2[162]);
    BiasedRNG[210] = (LFSRcolor2[57]&LFSRcolor2[11]&LFSRcolor2[191]&LFSRcolor2[166]);
    BiasedRNG[211] = (LFSRcolor2[228]&LFSRcolor2[112]&LFSRcolor2[72]&LFSRcolor2[246]);
    BiasedRNG[212] = (LFSRcolor2[287]&LFSRcolor2[6]&LFSRcolor2[81]&LFSRcolor2[199]);
    BiasedRNG[213] = (LFSRcolor2[139]&LFSRcolor2[9]&LFSRcolor2[38]&LFSRcolor2[298]);
    BiasedRNG[214] = (LFSRcolor2[93]&LFSRcolor2[136]&LFSRcolor2[313]&LFSRcolor2[102]);
    BiasedRNG[215] = (LFSRcolor2[149]&LFSRcolor2[78]&LFSRcolor2[61]&LFSRcolor2[259]);
    BiasedRNG[216] = (LFSRcolor2[83]&LFSRcolor2[18]&LFSRcolor2[68]&LFSRcolor2[282]);
    BiasedRNG[217] = (LFSRcolor2[142]&LFSRcolor2[91]&LFSRcolor2[239]&LFSRcolor2[171]);
    BiasedRNG[218] = (LFSRcolor2[117]&LFSRcolor2[205]&LFSRcolor2[103]&LFSRcolor2[225]);
    BiasedRNG[219] = (LFSRcolor2[160]&LFSRcolor2[209]&LFSRcolor2[122]&LFSRcolor2[277]);
    BiasedRNG[220] = (LFSRcolor2[310]&LFSRcolor2[2]&LFSRcolor2[311]&LFSRcolor2[48]);
    BiasedRNG[221] = (LFSRcolor2[268]&LFSRcolor2[71]&LFSRcolor2[27]&LFSRcolor2[316]);
    BiasedRNG[222] = (LFSRcolor2[305]&LFSRcolor2[165]&LFSRcolor2[309]&LFSRcolor2[291]);
    UnbiasedRNG[120] = LFSRcolor2[219];
    UnbiasedRNG[121] = LFSRcolor2[152];
    UnbiasedRNG[122] = LFSRcolor2[173];
    UnbiasedRNG[123] = LFSRcolor2[223];
    UnbiasedRNG[124] = LFSRcolor2[134];
    UnbiasedRNG[125] = LFSRcolor2[70];
    UnbiasedRNG[126] = LFSRcolor2[66];
    UnbiasedRNG[127] = LFSRcolor2[110];
    UnbiasedRNG[128] = LFSRcolor2[257];
    UnbiasedRNG[129] = LFSRcolor2[269];
    UnbiasedRNG[130] = LFSRcolor2[41];
    UnbiasedRNG[131] = LFSRcolor2[79];
    UnbiasedRNG[132] = LFSRcolor2[212];
    UnbiasedRNG[133] = LFSRcolor2[150];
    UnbiasedRNG[134] = LFSRcolor2[224];
    UnbiasedRNG[135] = LFSRcolor2[276];
    UnbiasedRNG[136] = LFSRcolor2[130];
    UnbiasedRNG[137] = LFSRcolor2[193];
    UnbiasedRNG[138] = LFSRcolor2[10];
    UnbiasedRNG[139] = LFSRcolor2[318];
    UnbiasedRNG[140] = LFSRcolor2[214];
    UnbiasedRNG[141] = LFSRcolor2[125];
    UnbiasedRNG[142] = LFSRcolor2[241];
    UnbiasedRNG[143] = LFSRcolor2[240];
    UnbiasedRNG[144] = LFSRcolor2[248];
    UnbiasedRNG[145] = LFSRcolor2[288];
    UnbiasedRNG[146] = LFSRcolor2[238];
    UnbiasedRNG[147] = LFSRcolor2[49];
    UnbiasedRNG[148] = LFSRcolor2[293];
    UnbiasedRNG[149] = LFSRcolor2[321];
    UnbiasedRNG[150] = LFSRcolor2[227];
    UnbiasedRNG[151] = LFSRcolor2[89];
    UnbiasedRNG[152] = LFSRcolor2[77];
    UnbiasedRNG[153] = LFSRcolor2[182];
    UnbiasedRNG[154] = LFSRcolor2[47];
    UnbiasedRNG[155] = LFSRcolor2[201];
    UnbiasedRNG[156] = LFSRcolor2[283];
    UnbiasedRNG[157] = LFSRcolor2[319];
    UnbiasedRNG[158] = LFSRcolor2[308];
    UnbiasedRNG[159] = LFSRcolor2[24];
    UnbiasedRNG[160] = LFSRcolor2[314];
    UnbiasedRNG[161] = LFSRcolor2[144];
    UnbiasedRNG[162] = LFSRcolor2[286];
    UnbiasedRNG[163] = LFSRcolor2[274];
    UnbiasedRNG[164] = LFSRcolor2[270];
    UnbiasedRNG[165] = LFSRcolor2[69];
    UnbiasedRNG[166] = LFSRcolor2[207];
    UnbiasedRNG[167] = LFSRcolor2[92];
    UnbiasedRNG[168] = LFSRcolor2[62];
    UnbiasedRNG[169] = LFSRcolor2[272];
    UnbiasedRNG[170] = LFSRcolor2[46];
    UnbiasedRNG[171] = LFSRcolor2[99];
    UnbiasedRNG[172] = LFSRcolor2[143];
    UnbiasedRNG[173] = LFSRcolor2[145];
    UnbiasedRNG[174] = LFSRcolor2[29];
    UnbiasedRNG[175] = LFSRcolor2[174];
end

always @(posedge color2_clk) begin
    UnbiasedRNG[176] = LFSRcolor3[30];
    UnbiasedRNG[177] = LFSRcolor3[20];
    UnbiasedRNG[178] = LFSRcolor3[4];
    UnbiasedRNG[179] = LFSRcolor3[34];
    UnbiasedRNG[180] = LFSRcolor3[40];
    UnbiasedRNG[181] = LFSRcolor3[17];
    UnbiasedRNG[182] = LFSRcolor3[12];
    UnbiasedRNG[183] = LFSRcolor3[23];
    UnbiasedRNG[184] = LFSRcolor3[26];
    UnbiasedRNG[185] = LFSRcolor3[29];
    UnbiasedRNG[186] = LFSRcolor3[25];
    UnbiasedRNG[187] = LFSRcolor3[1];
    UnbiasedRNG[188] = LFSRcolor3[5];
    UnbiasedRNG[189] = LFSRcolor3[14];
    UnbiasedRNG[190] = LFSRcolor3[24];
    UnbiasedRNG[191] = LFSRcolor3[0];
    UnbiasedRNG[192] = LFSRcolor3[15];
    UnbiasedRNG[193] = LFSRcolor3[28];
    UnbiasedRNG[194] = LFSRcolor3[22];
    UnbiasedRNG[195] = LFSRcolor3[43];
    UnbiasedRNG[196] = LFSRcolor3[3];
    UnbiasedRNG[197] = LFSRcolor3[32];
    UnbiasedRNG[198] = LFSRcolor3[45];
    UnbiasedRNG[199] = LFSRcolor3[44];
    UnbiasedRNG[200] = LFSRcolor3[33];
    UnbiasedRNG[201] = LFSRcolor3[19];
    UnbiasedRNG[202] = LFSRcolor3[10];
    UnbiasedRNG[203] = LFSRcolor3[38];
    UnbiasedRNG[204] = LFSRcolor3[6];
    UnbiasedRNG[205] = LFSRcolor3[16];
    UnbiasedRNG[206] = LFSRcolor3[21];
    UnbiasedRNG[207] = LFSRcolor3[27];
    UnbiasedRNG[208] = LFSRcolor3[7];
    UnbiasedRNG[209] = LFSRcolor3[11];
    UnbiasedRNG[210] = LFSRcolor3[9];
    UnbiasedRNG[211] = LFSRcolor3[35];
    UnbiasedRNG[212] = LFSRcolor3[41];
    UnbiasedRNG[213] = LFSRcolor3[36];
    UnbiasedRNG[214] = LFSRcolor3[42];
    UnbiasedRNG[215] = LFSRcolor3[13];
    UnbiasedRNG[216] = LFSRcolor3[39];
    UnbiasedRNG[217] = LFSRcolor3[8];
end

always @(posedge color3_clk) begin
    BiasedRNG[223] = (LFSRcolor4[28]&LFSRcolor4[198]&LFSRcolor4[221]&LFSRcolor4[115]);
    BiasedRNG[224] = (LFSRcolor4[175]&LFSRcolor4[188]&LFSRcolor4[13]&LFSRcolor4[124]);
    BiasedRNG[225] = (LFSRcolor4[213]&LFSRcolor4[136]&LFSRcolor4[155]&LFSRcolor4[19]);
    BiasedRNG[226] = (LFSRcolor4[129]&LFSRcolor4[167]&LFSRcolor4[184]&LFSRcolor4[45]);
    BiasedRNG[227] = (LFSRcolor4[39]&LFSRcolor4[171]&LFSRcolor4[50]&LFSRcolor4[154]);
    BiasedRNG[228] = (LFSRcolor4[201]&LFSRcolor4[212]&LFSRcolor4[25]&LFSRcolor4[86]);
    BiasedRNG[229] = (LFSRcolor4[111]&LFSRcolor4[177]&LFSRcolor4[31]&LFSRcolor4[169]);
    BiasedRNG[230] = (LFSRcolor4[40]&LFSRcolor4[87]&LFSRcolor4[137]&LFSRcolor4[220]);
    BiasedRNG[231] = (LFSRcolor4[69]&LFSRcolor4[22]&LFSRcolor4[227]&LFSRcolor4[71]);
    BiasedRNG[232] = (LFSRcolor4[8]&LFSRcolor4[36]&LFSRcolor4[110]&LFSRcolor4[17]);
    BiasedRNG[233] = (LFSRcolor4[214]&LFSRcolor4[24]&LFSRcolor4[53]&LFSRcolor4[215]);
    BiasedRNG[234] = (LFSRcolor4[104]&LFSRcolor4[95]&LFSRcolor4[209]&LFSRcolor4[162]);
    BiasedRNG[235] = (LFSRcolor4[186]&LFSRcolor4[52]&LFSRcolor4[49]&LFSRcolor4[11]);
    BiasedRNG[236] = (LFSRcolor4[119]&LFSRcolor4[163]&LFSRcolor4[191]&LFSRcolor4[2]);
    BiasedRNG[237] = (LFSRcolor4[108]&LFSRcolor4[127]&LFSRcolor4[208]&LFSRcolor4[189]);
    BiasedRNG[238] = (LFSRcolor4[168]&LFSRcolor4[66]&LFSRcolor4[126]&LFSRcolor4[12]);
    BiasedRNG[239] = (LFSRcolor4[6]&LFSRcolor4[105]&LFSRcolor4[123]&LFSRcolor4[113]);
    BiasedRNG[240] = (LFSRcolor4[112]&LFSRcolor4[157]&LFSRcolor4[100]&LFSRcolor4[196]);
    BiasedRNG[241] = (LFSRcolor4[204]&LFSRcolor4[161]&LFSRcolor4[197]&LFSRcolor4[121]);
    BiasedRNG[242] = (LFSRcolor4[183]&LFSRcolor4[203]&LFSRcolor4[29]&LFSRcolor4[134]);
    BiasedRNG[243] = (LFSRcolor4[77]&LFSRcolor4[97]&LFSRcolor4[120]&LFSRcolor4[225]);
    BiasedRNG[244] = (LFSRcolor4[10]&LFSRcolor4[192]&LFSRcolor4[141]&LFSRcolor4[190]);
    BiasedRNG[245] = (LFSRcolor4[159]&LFSRcolor4[68]&LFSRcolor4[145]&LFSRcolor4[47]);
    BiasedRNG[246] = (LFSRcolor4[199]&LFSRcolor4[207]&LFSRcolor4[74]&LFSRcolor4[33]);
    BiasedRNG[247] = (LFSRcolor4[179]&LFSRcolor4[57]&LFSRcolor4[224]&LFSRcolor4[229]);
    BiasedRNG[248] = (LFSRcolor4[23]&LFSRcolor4[20]&LFSRcolor4[65]&LFSRcolor4[181]);
    BiasedRNG[249] = (LFSRcolor4[58]&LFSRcolor4[0]&LFSRcolor4[210]&LFSRcolor4[165]);
    BiasedRNG[250] = (LFSRcolor4[34]&LFSRcolor4[139]&LFSRcolor4[200]&LFSRcolor4[143]);
    BiasedRNG[251] = (LFSRcolor4[89]&LFSRcolor4[195]&LFSRcolor4[35]&LFSRcolor4[4]);
    BiasedRNG[252] = (LFSRcolor4[106]&LFSRcolor4[14]&LFSRcolor4[142]&LFSRcolor4[44]);
    BiasedRNG[253] = (LFSRcolor4[5]&LFSRcolor4[122]&LFSRcolor4[90]&LFSRcolor4[101]);
    BiasedRNG[254] = (LFSRcolor4[178]&LFSRcolor4[144]&LFSRcolor4[135]&LFSRcolor4[222]);
    BiasedRNG[255] = (LFSRcolor4[153]&LFSRcolor4[173]&LFSRcolor4[116]&LFSRcolor4[67]);
    BiasedRNG[256] = (LFSRcolor4[117]&LFSRcolor4[60]&LFSRcolor4[48]&LFSRcolor4[193]);
    BiasedRNG[257] = (LFSRcolor4[194]&LFSRcolor4[41]&LFSRcolor4[55]&LFSRcolor4[73]);
    BiasedRNG[258] = (LFSRcolor4[64]&LFSRcolor4[103]&LFSRcolor4[150]&LFSRcolor4[174]);
    BiasedRNG[259] = (LFSRcolor4[131]&LFSRcolor4[76]&LFSRcolor4[170]&LFSRcolor4[205]);
    BiasedRNG[260] = (LFSRcolor4[78]&LFSRcolor4[125]&LFSRcolor4[216]&LFSRcolor4[43]);
    BiasedRNG[261] = (LFSRcolor4[38]&LFSRcolor4[80]&LFSRcolor4[109]&LFSRcolor4[27]);
    BiasedRNG[262] = (LFSRcolor4[217]&LFSRcolor4[30]&LFSRcolor4[211]&LFSRcolor4[54]);
    BiasedRNG[263] = (LFSRcolor4[62]&LFSRcolor4[7]&LFSRcolor4[46]&LFSRcolor4[83]);
    BiasedRNG[264] = (LFSRcolor4[93]&LFSRcolor4[96]&LFSRcolor4[61]&LFSRcolor4[51]);
    BiasedRNG[265] = (LFSRcolor4[42]&LFSRcolor4[21]&LFSRcolor4[59]&LFSRcolor4[152]);
    BiasedRNG[266] = (LFSRcolor4[56]&LFSRcolor4[148]&LFSRcolor4[16]&LFSRcolor4[146]);
    BiasedRNG[267] = (LFSRcolor4[156]&LFSRcolor4[223]&LFSRcolor4[133]&LFSRcolor4[187]);
    BiasedRNG[268] = (LFSRcolor4[202]&LFSRcolor4[226]&LFSRcolor4[15]&LFSRcolor4[138]);
    BiasedRNG[269] = (LFSRcolor4[1]&LFSRcolor4[160]&LFSRcolor4[164]&LFSRcolor4[102]);
    BiasedRNG[270] = (LFSRcolor4[63]&LFSRcolor4[147]&LFSRcolor4[72]&LFSRcolor4[79]);
    BiasedRNG[271] = (LFSRcolor4[82]&LFSRcolor4[151]&LFSRcolor4[99]&LFSRcolor4[9]);
    BiasedRNG[272] = (LFSRcolor4[182]&LFSRcolor4[218]&LFSRcolor4[88]&LFSRcolor4[75]);
    BiasedRNG[273] = (LFSRcolor4[128]&LFSRcolor4[172]&LFSRcolor4[180]&LFSRcolor4[140]);
    BiasedRNG[274] = (LFSRcolor4[37]&LFSRcolor4[98]&LFSRcolor4[149]&LFSRcolor4[228]);
    BiasedRNG[275] = (LFSRcolor4[166]&LFSRcolor4[92]&LFSRcolor4[206]&LFSRcolor4[118]);
    BiasedRNG[276] = (LFSRcolor4[26]&LFSRcolor4[18]&LFSRcolor4[91]&LFSRcolor4[185]);
    BiasedRNG[277] = (LFSRcolor4[84]&LFSRcolor4[81]&LFSRcolor4[94]&LFSRcolor4[219]);
end

//Generate the 40MHz shifted clocks:
clk_wiz_0 myPLL(.clk_out1(sample_clk),.clk_out2(color0_clk),.clk_out3(color1_clk),.clk_out4(color2_clk),.clk_out5(color3_clk),.clk_out6(color4_clk),.clk_in1_p(SYS_CLK_100M_P),.clk_in1_n(SYS_CLK_100M_N));

endmodule

//Module for generating LFSR:
module lfsr #(parameter seed = 46'b1) (output reg[45:0] LFSRregister, input clk);

//Set it to the seed to begin:
initial begin
    LFSRregister = seed;
end

//Shift and replace zeroth bit:
always @(negedge clk) begin
    LFSRregister[45:0] = {LFSRregister[44:0],(LFSRregister[45] ^ LFSRregister[39] ^ LFSRregister[38] ^ LFSRregister[37])};
end
endmodule